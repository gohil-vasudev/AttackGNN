module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n106_, keyIn_0_26 );
not g001 ( new_n107_, N1 );
not g002 ( new_n108_, keyIn_0_18 );
not g003 ( new_n109_, keyIn_0_13 );
not g004 ( new_n110_, keyIn_0_11 );
not g005 ( new_n111_, keyIn_0_7 );
or g006 ( new_n112_, N33, N37 );
and g007 ( new_n113_, N33, N37 );
not g008 ( new_n114_, new_n113_ );
and g009 ( new_n115_, new_n114_, new_n112_ );
or g010 ( new_n116_, new_n115_, keyIn_0_2 );
and g011 ( new_n117_, new_n114_, keyIn_0_2, new_n112_ );
not g012 ( new_n118_, new_n117_ );
and g013 ( new_n119_, new_n116_, new_n118_ );
not g014 ( new_n120_, keyIn_0_3 );
or g015 ( new_n121_, N41, N45 );
and g016 ( new_n122_, N41, N45 );
not g017 ( new_n123_, new_n122_ );
and g018 ( new_n124_, new_n123_, new_n121_ );
or g019 ( new_n125_, new_n124_, new_n120_ );
and g020 ( new_n126_, new_n123_, new_n120_, new_n121_ );
not g021 ( new_n127_, new_n126_ );
and g022 ( new_n128_, new_n125_, new_n127_ );
or g023 ( new_n129_, new_n119_, new_n128_ );
and g024 ( new_n130_, new_n116_, new_n125_, new_n118_, new_n127_ );
not g025 ( new_n131_, new_n130_ );
and g026 ( new_n132_, new_n129_, new_n131_ );
or g027 ( new_n133_, new_n132_, new_n111_ );
and g028 ( new_n134_, new_n129_, new_n111_, new_n131_ );
not g029 ( new_n135_, new_n134_ );
and g030 ( new_n136_, new_n133_, new_n135_ );
not g031 ( new_n137_, keyIn_0_8 );
or g032 ( new_n138_, N49, N53 );
and g033 ( new_n139_, N49, N53 );
not g034 ( new_n140_, new_n139_ );
and g035 ( new_n141_, new_n140_, new_n138_ );
or g036 ( new_n142_, new_n141_, keyIn_0_4 );
and g037 ( new_n143_, new_n140_, keyIn_0_4, new_n138_ );
not g038 ( new_n144_, new_n143_ );
and g039 ( new_n145_, new_n142_, new_n144_ );
not g040 ( new_n146_, keyIn_0_5 );
or g041 ( new_n147_, N57, N61 );
and g042 ( new_n148_, N57, N61 );
not g043 ( new_n149_, new_n148_ );
and g044 ( new_n150_, new_n149_, new_n147_ );
or g045 ( new_n151_, new_n150_, new_n146_ );
and g046 ( new_n152_, new_n149_, new_n146_, new_n147_ );
not g047 ( new_n153_, new_n152_ );
and g048 ( new_n154_, new_n151_, new_n153_ );
or g049 ( new_n155_, new_n145_, new_n154_ );
and g050 ( new_n156_, new_n142_, new_n151_, new_n144_, new_n153_ );
not g051 ( new_n157_, new_n156_ );
and g052 ( new_n158_, new_n155_, new_n157_ );
or g053 ( new_n159_, new_n158_, new_n137_ );
and g054 ( new_n160_, new_n155_, new_n137_, new_n157_ );
not g055 ( new_n161_, new_n160_ );
and g056 ( new_n162_, new_n159_, new_n161_ );
or g057 ( new_n163_, new_n136_, new_n162_ );
and g058 ( new_n164_, new_n133_, new_n159_, new_n135_, new_n161_ );
not g059 ( new_n165_, new_n164_ );
and g060 ( new_n166_, new_n163_, new_n165_ );
or g061 ( new_n167_, new_n166_, keyIn_0_9 );
and g062 ( new_n168_, new_n163_, keyIn_0_9, new_n165_ );
not g063 ( new_n169_, new_n168_ );
and g064 ( new_n170_, new_n167_, new_n169_ );
and g065 ( new_n171_, N134, N137 );
not g066 ( new_n172_, new_n171_ );
or g067 ( new_n173_, new_n170_, new_n172_ );
and g068 ( new_n174_, new_n167_, new_n169_, new_n172_ );
not g069 ( new_n175_, new_n174_ );
and g070 ( new_n176_, new_n173_, new_n175_ );
or g071 ( new_n177_, new_n176_, new_n110_ );
and g072 ( new_n178_, new_n173_, new_n110_, new_n175_ );
not g073 ( new_n179_, new_n178_ );
and g074 ( new_n180_, new_n177_, new_n179_ );
not g075 ( new_n181_, N69 );
not g076 ( new_n182_, N85 );
and g077 ( new_n183_, new_n181_, new_n182_ );
and g078 ( new_n184_, N69, N85 );
or g079 ( new_n185_, new_n183_, new_n184_ );
not g080 ( new_n186_, N101 );
not g081 ( new_n187_, N117 );
and g082 ( new_n188_, new_n186_, new_n187_ );
and g083 ( new_n189_, N101, N117 );
or g084 ( new_n190_, new_n188_, new_n189_ );
and g085 ( new_n191_, new_n185_, new_n190_ );
not g086 ( new_n192_, new_n185_ );
not g087 ( new_n193_, new_n190_ );
and g088 ( new_n194_, new_n192_, new_n193_ );
or g089 ( new_n195_, new_n194_, new_n191_ );
or g090 ( new_n196_, new_n180_, new_n195_ );
and g091 ( new_n197_, new_n177_, new_n179_, new_n195_ );
not g092 ( new_n198_, new_n197_ );
and g093 ( new_n199_, new_n196_, new_n198_ );
or g094 ( new_n200_, new_n199_, new_n109_ );
and g095 ( new_n201_, new_n196_, new_n109_, new_n198_ );
not g096 ( new_n202_, new_n201_ );
and g097 ( new_n203_, new_n200_, new_n202_ );
or g098 ( new_n204_, new_n203_, keyIn_0_15 );
and g099 ( new_n205_, new_n200_, keyIn_0_15, new_n202_ );
not g100 ( new_n206_, new_n205_ );
and g101 ( new_n207_, new_n204_, new_n206_ );
not g102 ( new_n208_, keyIn_0_6 );
or g103 ( new_n209_, N1, N5 );
not g104 ( new_n210_, new_n209_ );
and g105 ( new_n211_, N1, N5 );
or g106 ( new_n212_, new_n210_, new_n211_ );
and g107 ( new_n213_, new_n212_, keyIn_0_0 );
not g108 ( new_n214_, keyIn_0_0 );
not g109 ( new_n215_, new_n211_ );
and g110 ( new_n216_, new_n215_, new_n214_, new_n209_ );
or g111 ( new_n217_, new_n213_, new_n216_ );
not g112 ( new_n218_, keyIn_0_1 );
or g113 ( new_n219_, N9, N13 );
not g114 ( new_n220_, new_n219_ );
and g115 ( new_n221_, N9, N13 );
or g116 ( new_n222_, new_n220_, new_n221_ );
and g117 ( new_n223_, new_n222_, new_n218_ );
not g118 ( new_n224_, new_n221_ );
and g119 ( new_n225_, new_n224_, keyIn_0_1, new_n219_ );
or g120 ( new_n226_, new_n223_, new_n225_ );
and g121 ( new_n227_, new_n217_, new_n226_ );
and g122 ( new_n228_, new_n215_, new_n209_ );
or g123 ( new_n229_, new_n228_, new_n214_ );
not g124 ( new_n230_, new_n216_ );
and g125 ( new_n231_, new_n229_, new_n230_ );
and g126 ( new_n232_, new_n224_, new_n219_ );
or g127 ( new_n233_, new_n232_, keyIn_0_1 );
not g128 ( new_n234_, new_n225_ );
and g129 ( new_n235_, new_n233_, new_n234_ );
and g130 ( new_n236_, new_n231_, new_n235_ );
or g131 ( new_n237_, new_n227_, new_n236_ );
and g132 ( new_n238_, new_n237_, new_n208_ );
or g133 ( new_n239_, new_n231_, new_n235_ );
not g134 ( new_n240_, new_n236_ );
and g135 ( new_n241_, new_n240_, new_n239_ );
and g136 ( new_n242_, new_n241_, keyIn_0_6 );
or g137 ( new_n243_, new_n242_, new_n238_ );
not g138 ( new_n244_, N17 );
not g139 ( new_n245_, N21 );
and g140 ( new_n246_, new_n244_, new_n245_ );
and g141 ( new_n247_, N17, N21 );
or g142 ( new_n248_, new_n246_, new_n247_ );
not g143 ( new_n249_, N25 );
not g144 ( new_n250_, N29 );
and g145 ( new_n251_, new_n249_, new_n250_ );
and g146 ( new_n252_, N25, N29 );
or g147 ( new_n253_, new_n251_, new_n252_ );
and g148 ( new_n254_, new_n248_, new_n253_ );
not g149 ( new_n255_, new_n248_ );
not g150 ( new_n256_, new_n253_ );
and g151 ( new_n257_, new_n255_, new_n256_ );
or g152 ( new_n258_, new_n257_, new_n254_ );
and g153 ( new_n259_, new_n243_, new_n258_ );
or g154 ( new_n260_, new_n241_, keyIn_0_6 );
or g155 ( new_n261_, new_n237_, new_n208_ );
and g156 ( new_n262_, new_n260_, new_n261_ );
not g157 ( new_n263_, new_n258_ );
and g158 ( new_n264_, new_n262_, new_n263_ );
or g159 ( new_n265_, new_n259_, new_n264_ );
and g160 ( new_n266_, N133, N137 );
or g161 ( new_n267_, new_n265_, new_n266_ );
and g162 ( new_n268_, new_n265_, new_n266_ );
not g163 ( new_n269_, new_n268_ );
and g164 ( new_n270_, new_n269_, new_n267_ );
not g165 ( new_n271_, new_n270_ );
not g166 ( new_n272_, N81 );
and g167 ( new_n273_, new_n272_, N65 );
not g168 ( new_n274_, N65 );
and g169 ( new_n275_, new_n274_, N81 );
or g170 ( new_n276_, new_n273_, new_n275_ );
not g171 ( new_n277_, N97 );
not g172 ( new_n278_, N113 );
and g173 ( new_n279_, new_n277_, new_n278_ );
and g174 ( new_n280_, N97, N113 );
or g175 ( new_n281_, new_n279_, new_n280_ );
and g176 ( new_n282_, new_n276_, new_n281_ );
not g177 ( new_n283_, new_n276_ );
not g178 ( new_n284_, new_n281_ );
and g179 ( new_n285_, new_n283_, new_n284_ );
or g180 ( new_n286_, new_n285_, new_n282_ );
and g181 ( new_n287_, new_n271_, new_n286_ );
not g182 ( new_n288_, new_n287_ );
or g183 ( new_n289_, new_n271_, new_n286_ );
and g184 ( new_n290_, new_n288_, new_n289_ );
not g185 ( new_n291_, new_n290_ );
not g186 ( new_n292_, keyIn_0_14 );
not g187 ( new_n293_, keyIn_0_12 );
or g188 ( new_n294_, new_n262_, new_n136_ );
and g189 ( new_n295_, new_n262_, new_n136_ );
not g190 ( new_n296_, new_n295_ );
and g191 ( new_n297_, new_n296_, new_n294_ );
or g192 ( new_n298_, new_n297_, keyIn_0_10 );
not g193 ( new_n299_, keyIn_0_10 );
not g194 ( new_n300_, keyIn_0_2 );
not g195 ( new_n301_, N33 );
not g196 ( new_n302_, N37 );
and g197 ( new_n303_, new_n301_, new_n302_ );
or g198 ( new_n304_, new_n303_, new_n113_ );
and g199 ( new_n305_, new_n304_, new_n300_ );
or g200 ( new_n306_, new_n305_, new_n117_ );
not g201 ( new_n307_, N41 );
not g202 ( new_n308_, N45 );
and g203 ( new_n309_, new_n307_, new_n308_ );
or g204 ( new_n310_, new_n309_, new_n122_ );
and g205 ( new_n311_, new_n310_, keyIn_0_3 );
or g206 ( new_n312_, new_n311_, new_n126_ );
and g207 ( new_n313_, new_n306_, new_n312_ );
or g208 ( new_n314_, new_n313_, new_n130_ );
and g209 ( new_n315_, new_n314_, keyIn_0_7 );
or g210 ( new_n316_, new_n315_, new_n134_ );
and g211 ( new_n317_, new_n243_, new_n316_ );
or g212 ( new_n318_, new_n317_, new_n295_ );
or g213 ( new_n319_, new_n318_, new_n299_ );
and g214 ( new_n320_, new_n298_, new_n319_ );
and g215 ( new_n321_, N135, N137 );
or g216 ( new_n322_, new_n320_, new_n321_ );
and g217 ( new_n323_, new_n318_, new_n299_ );
and g218 ( new_n324_, new_n297_, keyIn_0_10 );
or g219 ( new_n325_, new_n324_, new_n323_ );
not g220 ( new_n326_, new_n321_ );
or g221 ( new_n327_, new_n325_, new_n326_ );
and g222 ( new_n328_, new_n322_, new_n327_ );
or g223 ( new_n329_, new_n328_, new_n293_ );
and g224 ( new_n330_, new_n325_, new_n326_ );
and g225 ( new_n331_, new_n320_, new_n321_ );
or g226 ( new_n332_, new_n330_, new_n331_, keyIn_0_12 );
and g227 ( new_n333_, new_n329_, new_n332_ );
not g228 ( new_n334_, N73 );
not g229 ( new_n335_, N89 );
and g230 ( new_n336_, new_n334_, new_n335_ );
and g231 ( new_n337_, N73, N89 );
or g232 ( new_n338_, new_n336_, new_n337_ );
not g233 ( new_n339_, N105 );
not g234 ( new_n340_, N121 );
and g235 ( new_n341_, new_n339_, new_n340_ );
and g236 ( new_n342_, N105, N121 );
or g237 ( new_n343_, new_n341_, new_n342_ );
and g238 ( new_n344_, new_n338_, new_n343_ );
not g239 ( new_n345_, new_n338_ );
not g240 ( new_n346_, new_n343_ );
and g241 ( new_n347_, new_n345_, new_n346_ );
or g242 ( new_n348_, new_n347_, new_n344_ );
not g243 ( new_n349_, new_n348_ );
or g244 ( new_n350_, new_n333_, new_n349_ );
or g245 ( new_n351_, new_n330_, new_n331_ );
and g246 ( new_n352_, new_n351_, keyIn_0_12 );
not g247 ( new_n353_, new_n332_ );
or g248 ( new_n354_, new_n352_, new_n353_, new_n348_ );
and g249 ( new_n355_, new_n350_, new_n354_ );
or g250 ( new_n356_, new_n355_, new_n292_ );
or g251 ( new_n357_, new_n352_, new_n353_ );
and g252 ( new_n358_, new_n357_, new_n348_ );
not g253 ( new_n359_, new_n354_ );
or g254 ( new_n360_, new_n358_, new_n359_, keyIn_0_14 );
and g255 ( new_n361_, new_n356_, new_n360_ );
not g256 ( new_n362_, keyIn_0_17 );
or g257 ( new_n363_, new_n274_, N69 );
or g258 ( new_n364_, new_n181_, N65 );
and g259 ( new_n365_, new_n363_, new_n364_ );
or g260 ( new_n366_, N73, N77 );
and g261 ( new_n367_, N73, N77 );
not g262 ( new_n368_, new_n367_ );
and g263 ( new_n369_, new_n368_, new_n366_ );
or g264 ( new_n370_, new_n365_, new_n369_ );
and g265 ( new_n371_, new_n365_, new_n369_ );
not g266 ( new_n372_, new_n371_ );
and g267 ( new_n373_, new_n372_, new_n370_ );
not g268 ( new_n374_, new_n373_ );
and g269 ( new_n375_, new_n186_, N97 );
and g270 ( new_n376_, new_n277_, N101 );
or g271 ( new_n377_, new_n375_, new_n376_ );
not g272 ( new_n378_, new_n377_ );
or g273 ( new_n379_, N105, N109 );
and g274 ( new_n380_, N105, N109 );
not g275 ( new_n381_, new_n380_ );
and g276 ( new_n382_, new_n381_, new_n379_ );
or g277 ( new_n383_, new_n378_, new_n382_ );
and g278 ( new_n384_, new_n378_, new_n382_ );
not g279 ( new_n385_, new_n384_ );
and g280 ( new_n386_, new_n385_, new_n383_ );
and g281 ( new_n387_, new_n386_, new_n374_ );
not g282 ( new_n388_, new_n386_ );
and g283 ( new_n389_, new_n388_, new_n373_ );
or g284 ( new_n390_, new_n389_, new_n387_ );
not g285 ( new_n391_, new_n390_ );
and g286 ( new_n392_, N131, N137 );
or g287 ( new_n393_, new_n391_, new_n392_ );
not g288 ( new_n394_, new_n393_ );
and g289 ( new_n395_, new_n391_, new_n392_ );
or g290 ( new_n396_, new_n394_, new_n395_ );
and g291 ( new_n397_, new_n249_, N9 );
not g292 ( new_n398_, N9 );
and g293 ( new_n399_, new_n398_, N25 );
or g294 ( new_n400_, new_n397_, new_n399_ );
not g295 ( new_n401_, N57 );
and g296 ( new_n402_, new_n307_, new_n401_ );
and g297 ( new_n403_, N41, N57 );
or g298 ( new_n404_, new_n402_, new_n403_ );
and g299 ( new_n405_, new_n400_, new_n404_ );
not g300 ( new_n406_, new_n400_ );
not g301 ( new_n407_, new_n404_ );
and g302 ( new_n408_, new_n406_, new_n407_ );
or g303 ( new_n409_, new_n408_, new_n405_ );
and g304 ( new_n410_, new_n396_, new_n409_ );
not g305 ( new_n411_, new_n395_ );
not g306 ( new_n412_, new_n409_ );
and g307 ( new_n413_, new_n411_, new_n393_, new_n412_ );
or g308 ( new_n414_, new_n410_, new_n413_ );
not g309 ( new_n415_, new_n414_ );
or g310 ( new_n416_, new_n272_, N85 );
or g311 ( new_n417_, new_n182_, N81 );
and g312 ( new_n418_, new_n416_, new_n417_ );
or g313 ( new_n419_, N89, N93 );
and g314 ( new_n420_, N89, N93 );
not g315 ( new_n421_, new_n420_ );
and g316 ( new_n422_, new_n421_, new_n419_ );
or g317 ( new_n423_, new_n418_, new_n422_ );
and g318 ( new_n424_, new_n418_, new_n422_ );
not g319 ( new_n425_, new_n424_ );
and g320 ( new_n426_, new_n425_, new_n423_ );
and g321 ( new_n427_, new_n374_, new_n426_ );
not g322 ( new_n428_, new_n426_ );
and g323 ( new_n429_, new_n428_, new_n373_ );
or g324 ( new_n430_, new_n427_, new_n429_ );
not g325 ( new_n431_, new_n430_ );
and g326 ( new_n432_, N129, N137 );
or g327 ( new_n433_, new_n431_, new_n432_ );
not g328 ( new_n434_, new_n433_ );
and g329 ( new_n435_, new_n431_, new_n432_ );
or g330 ( new_n436_, new_n434_, new_n435_ );
and g331 ( new_n437_, new_n107_, new_n244_ );
and g332 ( new_n438_, N1, N17 );
or g333 ( new_n439_, new_n437_, new_n438_ );
not g334 ( new_n440_, N49 );
and g335 ( new_n441_, new_n301_, new_n440_ );
and g336 ( new_n442_, N33, N49 );
or g337 ( new_n443_, new_n441_, new_n442_ );
and g338 ( new_n444_, new_n439_, new_n443_ );
not g339 ( new_n445_, new_n439_ );
not g340 ( new_n446_, new_n443_ );
and g341 ( new_n447_, new_n445_, new_n446_ );
or g342 ( new_n448_, new_n447_, new_n444_ );
and g343 ( new_n449_, new_n436_, new_n448_ );
not g344 ( new_n450_, new_n435_ );
and g345 ( new_n451_, new_n450_, new_n433_ );
not g346 ( new_n452_, new_n448_ );
and g347 ( new_n453_, new_n451_, new_n452_ );
or g348 ( new_n454_, new_n449_, new_n453_ );
and g349 ( new_n455_, new_n187_, N113 );
and g350 ( new_n456_, new_n278_, N117 );
or g351 ( new_n457_, new_n455_, new_n456_ );
not g352 ( new_n458_, new_n457_ );
or g353 ( new_n459_, N121, N125 );
and g354 ( new_n460_, N121, N125 );
not g355 ( new_n461_, new_n460_ );
and g356 ( new_n462_, new_n461_, new_n459_ );
or g357 ( new_n463_, new_n458_, new_n462_ );
and g358 ( new_n464_, new_n458_, new_n462_ );
not g359 ( new_n465_, new_n464_ );
and g360 ( new_n466_, new_n465_, new_n463_ );
and g361 ( new_n467_, new_n388_, new_n466_ );
not g362 ( new_n468_, new_n466_ );
and g363 ( new_n469_, new_n468_, new_n386_ );
or g364 ( new_n470_, new_n467_, new_n469_ );
and g365 ( new_n471_, N130, N137 );
not g366 ( new_n472_, new_n471_ );
and g367 ( new_n473_, new_n470_, new_n472_ );
not g368 ( new_n474_, new_n467_ );
not g369 ( new_n475_, new_n469_ );
and g370 ( new_n476_, new_n474_, new_n475_ );
and g371 ( new_n477_, new_n476_, new_n471_ );
or g372 ( new_n478_, new_n477_, new_n473_ );
not g373 ( new_n479_, N5 );
and g374 ( new_n480_, new_n479_, new_n245_ );
and g375 ( new_n481_, N5, N21 );
or g376 ( new_n482_, new_n480_, new_n481_ );
not g377 ( new_n483_, N53 );
and g378 ( new_n484_, new_n302_, new_n483_ );
and g379 ( new_n485_, N37, N53 );
or g380 ( new_n486_, new_n484_, new_n485_ );
and g381 ( new_n487_, new_n482_, new_n486_ );
not g382 ( new_n488_, new_n482_ );
not g383 ( new_n489_, new_n486_ );
and g384 ( new_n490_, new_n488_, new_n489_ );
or g385 ( new_n491_, new_n490_, new_n487_ );
and g386 ( new_n492_, new_n478_, new_n491_ );
not g387 ( new_n493_, new_n492_ );
not g388 ( new_n494_, new_n473_ );
not g389 ( new_n495_, new_n477_ );
not g390 ( new_n496_, new_n491_ );
and g391 ( new_n497_, new_n495_, new_n494_, new_n496_ );
not g392 ( new_n498_, new_n497_ );
and g393 ( new_n499_, new_n493_, new_n498_ );
or g394 ( new_n500_, new_n415_, new_n454_, new_n499_ );
or g395 ( new_n501_, new_n451_, new_n452_ );
not g396 ( new_n502_, new_n453_ );
and g397 ( new_n503_, new_n502_, new_n501_ );
or g398 ( new_n504_, new_n492_, new_n497_ );
or g399 ( new_n505_, new_n415_, new_n503_, new_n504_ );
and g400 ( new_n506_, new_n500_, new_n505_ );
and g401 ( new_n507_, new_n466_, new_n428_ );
and g402 ( new_n508_, new_n468_, new_n426_ );
or g403 ( new_n509_, new_n508_, new_n507_ );
not g404 ( new_n510_, new_n509_ );
and g405 ( new_n511_, N132, N137 );
or g406 ( new_n512_, new_n510_, new_n511_ );
and g407 ( new_n513_, new_n510_, new_n511_ );
not g408 ( new_n514_, new_n513_ );
and g409 ( new_n515_, new_n514_, new_n512_ );
and g410 ( new_n516_, new_n250_, N13 );
not g411 ( new_n517_, N13 );
and g412 ( new_n518_, new_n517_, N29 );
or g413 ( new_n519_, new_n516_, new_n518_ );
not g414 ( new_n520_, N61 );
and g415 ( new_n521_, new_n308_, new_n520_ );
and g416 ( new_n522_, N45, N61 );
or g417 ( new_n523_, new_n521_, new_n522_ );
and g418 ( new_n524_, new_n519_, new_n523_ );
not g419 ( new_n525_, new_n519_ );
not g420 ( new_n526_, new_n523_ );
and g421 ( new_n527_, new_n525_, new_n526_ );
or g422 ( new_n528_, new_n527_, new_n524_ );
not g423 ( new_n529_, new_n528_ );
or g424 ( new_n530_, new_n515_, new_n529_ );
and g425 ( new_n531_, new_n515_, new_n529_ );
not g426 ( new_n532_, new_n531_ );
and g427 ( new_n533_, new_n532_, new_n530_ );
or g428 ( new_n534_, new_n506_, new_n533_ );
or g429 ( new_n535_, new_n533_, new_n414_ );
and g430 ( new_n536_, new_n533_, new_n414_ );
not g431 ( new_n537_, new_n536_ );
and g432 ( new_n538_, new_n537_, new_n535_ );
or g433 ( new_n539_, new_n538_, new_n454_, new_n504_ );
and g434 ( new_n540_, new_n534_, new_n539_ );
or g435 ( new_n541_, new_n540_, new_n362_ );
and g436 ( new_n542_, new_n503_, new_n504_ );
and g437 ( new_n543_, new_n542_, new_n414_ );
and g438 ( new_n544_, new_n499_, new_n454_ );
and g439 ( new_n545_, new_n544_, new_n414_ );
or g440 ( new_n546_, new_n543_, new_n545_ );
not g441 ( new_n547_, new_n530_ );
or g442 ( new_n548_, new_n547_, new_n531_ );
and g443 ( new_n549_, new_n546_, new_n548_ );
not g444 ( new_n550_, new_n535_ );
or g445 ( new_n551_, new_n550_, new_n536_ );
and g446 ( new_n552_, new_n551_, new_n503_, new_n499_ );
or g447 ( new_n553_, new_n552_, new_n549_, keyIn_0_17 );
and g448 ( new_n554_, new_n541_, new_n553_ );
not g449 ( new_n555_, keyIn_0_4 );
and g450 ( new_n556_, new_n440_, new_n483_ );
or g451 ( new_n557_, new_n556_, new_n139_ );
and g452 ( new_n558_, new_n557_, new_n555_ );
or g453 ( new_n559_, new_n558_, new_n143_ );
and g454 ( new_n560_, new_n401_, new_n520_ );
or g455 ( new_n561_, new_n560_, new_n148_ );
and g456 ( new_n562_, new_n561_, keyIn_0_5 );
or g457 ( new_n563_, new_n562_, new_n152_ );
and g458 ( new_n564_, new_n559_, new_n563_ );
or g459 ( new_n565_, new_n564_, new_n156_ );
and g460 ( new_n566_, new_n565_, keyIn_0_8 );
or g461 ( new_n567_, new_n566_, new_n160_ );
and g462 ( new_n568_, new_n567_, new_n263_ );
and g463 ( new_n569_, new_n162_, new_n258_ );
or g464 ( new_n570_, new_n568_, new_n569_ );
not g465 ( new_n571_, new_n570_ );
and g466 ( new_n572_, N136, N137 );
or g467 ( new_n573_, new_n571_, new_n572_ );
and g468 ( new_n574_, new_n571_, new_n572_ );
not g469 ( new_n575_, new_n574_ );
and g470 ( new_n576_, new_n575_, new_n573_ );
not g471 ( new_n577_, new_n576_ );
not g472 ( new_n578_, N93 );
and g473 ( new_n579_, new_n578_, N77 );
not g474 ( new_n580_, N77 );
and g475 ( new_n581_, new_n580_, N93 );
or g476 ( new_n582_, new_n579_, new_n581_ );
not g477 ( new_n583_, N109 );
not g478 ( new_n584_, N125 );
and g479 ( new_n585_, new_n583_, new_n584_ );
and g480 ( new_n586_, N109, N125 );
or g481 ( new_n587_, new_n585_, new_n586_ );
and g482 ( new_n588_, new_n582_, new_n587_ );
not g483 ( new_n589_, new_n582_ );
not g484 ( new_n590_, new_n587_ );
and g485 ( new_n591_, new_n589_, new_n590_ );
or g486 ( new_n592_, new_n591_, new_n588_ );
and g487 ( new_n593_, new_n577_, new_n592_ );
not g488 ( new_n594_, new_n593_ );
or g489 ( new_n595_, new_n577_, new_n592_ );
and g490 ( new_n596_, new_n594_, new_n595_ );
or g491 ( new_n597_, new_n554_, new_n596_ );
or g492 ( new_n598_, new_n361_, new_n291_, new_n597_ );
or g493 ( new_n599_, new_n207_, new_n598_ );
and g494 ( new_n600_, new_n599_, new_n108_ );
not g495 ( new_n601_, keyIn_0_15 );
not g496 ( new_n602_, keyIn_0_9 );
and g497 ( new_n603_, new_n316_, new_n567_ );
or g498 ( new_n604_, new_n603_, new_n164_ );
and g499 ( new_n605_, new_n604_, new_n602_ );
or g500 ( new_n606_, new_n605_, new_n168_ );
and g501 ( new_n607_, new_n606_, new_n171_ );
or g502 ( new_n608_, new_n607_, new_n174_ );
and g503 ( new_n609_, new_n608_, keyIn_0_11 );
or g504 ( new_n610_, new_n609_, new_n178_ );
not g505 ( new_n611_, new_n195_ );
and g506 ( new_n612_, new_n610_, new_n611_ );
or g507 ( new_n613_, new_n612_, new_n197_ );
and g508 ( new_n614_, new_n613_, keyIn_0_13 );
or g509 ( new_n615_, new_n614_, new_n201_ );
and g510 ( new_n616_, new_n615_, new_n601_ );
or g511 ( new_n617_, new_n616_, new_n205_ );
or g512 ( new_n618_, new_n358_, new_n359_ );
and g513 ( new_n619_, new_n618_, keyIn_0_14 );
not g514 ( new_n620_, new_n360_ );
or g515 ( new_n621_, new_n619_, new_n620_ );
not g516 ( new_n622_, new_n597_ );
and g517 ( new_n623_, new_n621_, new_n622_, new_n290_ );
and g518 ( new_n624_, new_n617_, keyIn_0_18, new_n623_ );
or g519 ( new_n625_, new_n624_, new_n503_ );
or g520 ( new_n626_, new_n625_, new_n600_ );
and g521 ( new_n627_, new_n626_, keyIn_0_20 );
not g522 ( new_n628_, keyIn_0_20 );
not g523 ( new_n629_, new_n600_ );
not g524 ( new_n630_, new_n624_ );
and g525 ( new_n631_, new_n629_, new_n628_, new_n454_, new_n630_ );
or g526 ( new_n632_, new_n627_, new_n631_ );
and g527 ( new_n633_, new_n632_, new_n107_ );
not g528 ( new_n634_, new_n627_ );
not g529 ( new_n635_, new_n631_ );
and g530 ( new_n636_, new_n634_, new_n635_, N1 );
or g531 ( new_n637_, new_n633_, new_n636_ );
and g532 ( new_n638_, new_n637_, new_n106_ );
not g533 ( new_n639_, new_n633_ );
not g534 ( new_n640_, new_n636_ );
and g535 ( new_n641_, new_n639_, new_n640_, keyIn_0_26 );
or g536 ( N724, new_n638_, new_n641_ );
not g537 ( new_n643_, keyIn_0_27 );
or g538 ( new_n644_, new_n624_, new_n499_ );
or g539 ( new_n645_, new_n644_, new_n600_ );
and g540 ( new_n646_, new_n645_, keyIn_0_21 );
not g541 ( new_n647_, keyIn_0_21 );
and g542 ( new_n648_, new_n629_, new_n647_, new_n504_, new_n630_ );
or g543 ( new_n649_, new_n646_, new_n648_ );
and g544 ( new_n650_, new_n649_, N5 );
not g545 ( new_n651_, new_n646_ );
not g546 ( new_n652_, new_n648_ );
and g547 ( new_n653_, new_n651_, new_n652_, new_n479_ );
or g548 ( new_n654_, new_n650_, new_n653_ );
and g549 ( new_n655_, new_n654_, new_n643_ );
not g550 ( new_n656_, new_n650_ );
not g551 ( new_n657_, new_n653_ );
and g552 ( new_n658_, new_n656_, new_n657_, keyIn_0_27 );
or g553 ( N725, new_n655_, new_n658_ );
or g554 ( new_n660_, new_n624_, new_n414_ );
or g555 ( new_n661_, new_n660_, new_n600_ );
and g556 ( new_n662_, new_n661_, keyIn_0_22 );
not g557 ( new_n663_, keyIn_0_22 );
and g558 ( new_n664_, new_n629_, new_n663_, new_n415_, new_n630_ );
or g559 ( new_n665_, new_n662_, new_n664_ );
and g560 ( new_n666_, new_n665_, new_n398_ );
not g561 ( new_n667_, new_n662_ );
not g562 ( new_n668_, new_n664_ );
and g563 ( new_n669_, new_n667_, new_n668_, N9 );
or g564 ( new_n670_, new_n666_, new_n669_ );
and g565 ( new_n671_, new_n670_, keyIn_0_28 );
not g566 ( new_n672_, keyIn_0_28 );
not g567 ( new_n673_, new_n666_ );
not g568 ( new_n674_, new_n669_ );
and g569 ( new_n675_, new_n673_, new_n674_, new_n672_ );
or g570 ( N726, new_n671_, new_n675_ );
not g571 ( new_n677_, keyIn_0_29 );
or g572 ( new_n678_, new_n624_, new_n548_ );
or g573 ( new_n679_, new_n678_, new_n600_ );
and g574 ( new_n680_, new_n679_, keyIn_0_23 );
not g575 ( new_n681_, keyIn_0_23 );
and g576 ( new_n682_, new_n629_, new_n681_, new_n533_, new_n630_ );
or g577 ( new_n683_, new_n680_, new_n682_ );
and g578 ( new_n684_, new_n683_, new_n517_ );
not g579 ( new_n685_, new_n680_ );
not g580 ( new_n686_, new_n682_ );
and g581 ( new_n687_, new_n685_, new_n686_, N13 );
or g582 ( new_n688_, new_n684_, new_n687_ );
and g583 ( new_n689_, new_n688_, new_n677_ );
not g584 ( new_n690_, new_n684_ );
not g585 ( new_n691_, new_n687_ );
and g586 ( new_n692_, new_n690_, new_n691_, keyIn_0_29 );
or g587 ( N727, new_n689_, new_n692_ );
not g588 ( new_n694_, keyIn_0_19 );
and g589 ( new_n695_, new_n615_, new_n290_ );
not g590 ( new_n696_, new_n554_ );
and g591 ( new_n697_, new_n696_, new_n596_ );
and g592 ( new_n698_, new_n695_, new_n361_, new_n697_ );
and g593 ( new_n699_, new_n698_, new_n694_ );
not g594 ( new_n700_, new_n699_ );
or g595 ( new_n701_, new_n698_, new_n694_ );
and g596 ( new_n702_, new_n700_, new_n454_, new_n701_ );
not g597 ( new_n703_, new_n702_ );
and g598 ( new_n704_, new_n703_, N17 );
and g599 ( new_n705_, new_n702_, new_n244_ );
or g600 ( N728, new_n704_, new_n705_ );
not g601 ( new_n707_, keyIn_0_30 );
and g602 ( new_n708_, new_n700_, new_n504_, new_n701_ );
or g603 ( new_n709_, new_n708_, keyIn_0_24 );
not g604 ( new_n710_, new_n709_ );
and g605 ( new_n711_, new_n708_, keyIn_0_24 );
or g606 ( new_n712_, new_n710_, new_n711_ );
and g607 ( new_n713_, new_n712_, new_n245_ );
not g608 ( new_n714_, new_n711_ );
and g609 ( new_n715_, new_n714_, new_n709_ );
and g610 ( new_n716_, new_n715_, N21 );
or g611 ( new_n717_, new_n713_, new_n716_ );
and g612 ( new_n718_, new_n717_, new_n707_ );
not g613 ( new_n719_, new_n713_ );
not g614 ( new_n720_, new_n716_ );
and g615 ( new_n721_, new_n719_, keyIn_0_30, new_n720_ );
or g616 ( N729, new_n718_, new_n721_ );
and g617 ( new_n723_, new_n700_, new_n415_, new_n701_ );
not g618 ( new_n724_, new_n723_ );
and g619 ( new_n725_, new_n724_, N25 );
and g620 ( new_n726_, new_n723_, new_n249_ );
or g621 ( N730, new_n725_, new_n726_ );
not g622 ( new_n728_, keyIn_0_31 );
and g623 ( new_n729_, new_n700_, new_n533_, new_n701_ );
or g624 ( new_n730_, new_n729_, keyIn_0_25 );
not g625 ( new_n731_, new_n730_ );
and g626 ( new_n732_, new_n729_, keyIn_0_25 );
or g627 ( new_n733_, new_n731_, new_n732_ );
and g628 ( new_n734_, new_n733_, new_n250_ );
not g629 ( new_n735_, new_n732_ );
and g630 ( new_n736_, new_n735_, new_n730_ );
and g631 ( new_n737_, new_n736_, N29 );
or g632 ( new_n738_, new_n734_, new_n737_ );
and g633 ( new_n739_, new_n738_, new_n728_ );
not g634 ( new_n740_, new_n734_ );
not g635 ( new_n741_, new_n737_ );
and g636 ( new_n742_, new_n740_, keyIn_0_31, new_n741_ );
or g637 ( N731, new_n739_, new_n742_ );
and g638 ( new_n744_, new_n203_, new_n291_ );
and g639 ( new_n745_, new_n744_, new_n621_, new_n622_ );
and g640 ( new_n746_, new_n745_, new_n454_ );
not g641 ( new_n747_, new_n746_ );
and g642 ( new_n748_, new_n747_, N33 );
and g643 ( new_n749_, new_n746_, new_n301_ );
or g644 ( N732, new_n748_, new_n749_ );
and g645 ( new_n751_, new_n745_, new_n504_ );
not g646 ( new_n752_, new_n751_ );
and g647 ( new_n753_, new_n752_, N37 );
and g648 ( new_n754_, new_n751_, new_n302_ );
or g649 ( N733, new_n753_, new_n754_ );
and g650 ( new_n756_, new_n745_, new_n415_ );
not g651 ( new_n757_, new_n756_ );
and g652 ( new_n758_, new_n757_, N41 );
and g653 ( new_n759_, new_n756_, new_n307_ );
or g654 ( N734, new_n758_, new_n759_ );
and g655 ( new_n761_, new_n745_, new_n533_ );
not g656 ( new_n762_, new_n761_ );
and g657 ( new_n763_, new_n762_, N45 );
and g658 ( new_n764_, new_n761_, new_n308_ );
or g659 ( N735, new_n763_, new_n764_ );
and g660 ( new_n766_, new_n744_, new_n361_ );
and g661 ( new_n767_, new_n766_, new_n697_ );
and g662 ( new_n768_, new_n767_, new_n454_ );
not g663 ( new_n769_, new_n768_ );
and g664 ( new_n770_, new_n769_, N49 );
and g665 ( new_n771_, new_n768_, new_n440_ );
or g666 ( N736, new_n770_, new_n771_ );
and g667 ( new_n773_, new_n767_, new_n504_ );
not g668 ( new_n774_, new_n773_ );
and g669 ( new_n775_, new_n774_, N53 );
and g670 ( new_n776_, new_n773_, new_n483_ );
or g671 ( N737, new_n775_, new_n776_ );
and g672 ( new_n778_, new_n767_, new_n415_ );
not g673 ( new_n779_, new_n778_ );
and g674 ( new_n780_, new_n779_, N57 );
and g675 ( new_n781_, new_n778_, new_n401_ );
or g676 ( N738, new_n780_, new_n781_ );
and g677 ( new_n783_, new_n767_, new_n533_ );
not g678 ( new_n784_, new_n783_ );
and g679 ( new_n785_, new_n784_, N61 );
and g680 ( new_n786_, new_n783_, new_n520_ );
or g681 ( N739, new_n785_, new_n786_ );
not g682 ( new_n788_, new_n766_ );
not g683 ( new_n789_, keyIn_0_16 );
and g684 ( new_n790_, new_n361_, new_n789_ );
and g685 ( new_n791_, new_n621_, keyIn_0_16 );
or g686 ( new_n792_, new_n791_, new_n790_, new_n203_, new_n291_ );
and g687 ( new_n793_, new_n792_, new_n788_ );
or g688 ( new_n794_, new_n793_, new_n596_ );
and g689 ( new_n795_, new_n361_, new_n596_ );
not g690 ( new_n796_, new_n596_ );
and g691 ( new_n797_, new_n621_, new_n796_ );
or g692 ( new_n798_, new_n797_, new_n795_ );
and g693 ( new_n799_, new_n798_, new_n615_, new_n291_ );
not g694 ( new_n800_, new_n799_ );
and g695 ( new_n801_, new_n794_, new_n800_ );
and g696 ( new_n802_, new_n550_, new_n544_ );
not g697 ( new_n803_, new_n802_ );
or g698 ( new_n804_, new_n801_, new_n803_ );
or g699 ( new_n805_, new_n804_, new_n291_ );
and g700 ( new_n806_, new_n805_, N65 );
not g701 ( new_n807_, new_n804_ );
and g702 ( new_n808_, new_n807_, new_n274_, new_n290_ );
or g703 ( N740, new_n806_, new_n808_ );
or g704 ( new_n810_, new_n804_, new_n615_ );
and g705 ( new_n811_, new_n810_, N69 );
and g706 ( new_n812_, new_n807_, new_n181_, new_n203_ );
or g707 ( N741, new_n811_, new_n812_ );
or g708 ( new_n814_, new_n804_, new_n361_ );
and g709 ( new_n815_, new_n814_, N73 );
and g710 ( new_n816_, new_n807_, new_n334_, new_n621_ );
or g711 ( N742, new_n815_, new_n816_ );
or g712 ( new_n818_, new_n804_, new_n796_ );
and g713 ( new_n819_, new_n818_, N77 );
and g714 ( new_n820_, new_n807_, new_n580_, new_n596_ );
or g715 ( N743, new_n819_, new_n820_ );
or g716 ( new_n822_, new_n801_, new_n505_, new_n548_ );
or g717 ( new_n823_, new_n822_, new_n291_ );
and g718 ( new_n824_, new_n823_, N81 );
not g719 ( new_n825_, new_n822_ );
and g720 ( new_n826_, new_n825_, new_n272_, new_n290_ );
or g721 ( N744, new_n824_, new_n826_ );
or g722 ( new_n828_, new_n822_, new_n615_ );
and g723 ( new_n829_, new_n828_, N85 );
and g724 ( new_n830_, new_n825_, new_n182_, new_n203_ );
or g725 ( N745, new_n829_, new_n830_ );
or g726 ( new_n832_, new_n822_, new_n361_ );
and g727 ( new_n833_, new_n832_, N89 );
and g728 ( new_n834_, new_n825_, new_n335_, new_n621_ );
or g729 ( N746, new_n833_, new_n834_ );
or g730 ( new_n836_, new_n822_, new_n796_ );
and g731 ( new_n837_, new_n836_, N93 );
and g732 ( new_n838_, new_n825_, new_n578_, new_n596_ );
or g733 ( N747, new_n837_, new_n838_ );
and g734 ( new_n840_, new_n550_, new_n542_ );
not g735 ( new_n841_, new_n840_ );
or g736 ( new_n842_, new_n801_, new_n841_ );
or g737 ( new_n843_, new_n842_, new_n291_ );
and g738 ( new_n844_, new_n843_, N97 );
not g739 ( new_n845_, new_n842_ );
and g740 ( new_n846_, new_n845_, new_n277_, new_n290_ );
or g741 ( N748, new_n844_, new_n846_ );
or g742 ( new_n848_, new_n842_, new_n615_ );
and g743 ( new_n849_, new_n848_, N101 );
and g744 ( new_n850_, new_n845_, new_n186_, new_n203_ );
or g745 ( N749, new_n849_, new_n850_ );
or g746 ( new_n852_, new_n842_, new_n361_ );
and g747 ( new_n853_, new_n852_, N105 );
and g748 ( new_n854_, new_n845_, new_n339_, new_n621_ );
or g749 ( N750, new_n853_, new_n854_ );
or g750 ( new_n856_, new_n842_, new_n796_ );
and g751 ( new_n857_, new_n856_, N109 );
and g752 ( new_n858_, new_n845_, new_n583_, new_n596_ );
or g753 ( N751, new_n857_, new_n858_ );
or g754 ( new_n860_, new_n801_, new_n500_, new_n548_ );
or g755 ( new_n861_, new_n860_, new_n291_ );
and g756 ( new_n862_, new_n861_, N113 );
not g757 ( new_n863_, new_n860_ );
and g758 ( new_n864_, new_n863_, new_n278_, new_n290_ );
or g759 ( N752, new_n862_, new_n864_ );
or g760 ( new_n866_, new_n860_, new_n615_ );
and g761 ( new_n867_, new_n866_, N117 );
and g762 ( new_n868_, new_n863_, new_n187_, new_n203_ );
or g763 ( N753, new_n867_, new_n868_ );
or g764 ( new_n870_, new_n860_, new_n361_ );
and g765 ( new_n871_, new_n870_, N121 );
and g766 ( new_n872_, new_n863_, new_n340_, new_n621_ );
or g767 ( N754, new_n871_, new_n872_ );
or g768 ( new_n874_, new_n860_, new_n796_ );
and g769 ( new_n875_, new_n874_, N125 );
and g770 ( new_n876_, new_n863_, new_n584_, new_n596_ );
or g771 ( N755, new_n875_, new_n876_ );
endmodule