module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n155_, new_n384_, new_n595_, new_n410_, new_n445_, new_n236_, new_n238_, new_n479_, new_n543_, new_n250_, new_n113_, new_n501_, new_n288_, new_n371_, new_n509_, new_n454_, new_n421_, new_n202_, new_n296_, new_n308_, new_n368_, new_n232_, new_n258_, new_n439_, new_n176_, new_n283_, new_n223_, new_n390_, new_n156_, new_n306_, new_n366_, new_n494_, new_n291_, new_n241_, new_n261_, new_n309_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n323_, new_n401_, new_n389_, new_n259_, new_n362_, new_n514_, new_n556_, new_n227_, new_n416_, new_n222_, new_n456_, new_n170_, new_n246_, new_n571_, new_n400_, new_n328_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n130_, new_n505_, new_n419_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n214_, new_n451_, new_n424_, new_n138_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n240_, new_n413_, new_n526_, new_n352_, new_n442_, new_n575_, new_n485_, new_n525_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n578_, new_n126_, new_n462_, new_n564_, new_n177_, new_n547_, new_n264_, new_n379_, new_n500_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n317_, new_n344_, new_n143_, new_n520_, new_n287_, new_n125_, new_n145_, new_n253_, new_n504_, new_n403_, new_n475_, new_n237_, new_n427_, new_n234_, new_n532_, new_n149_, new_n472_, new_n557_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n106_, new_n411_, new_n215_, new_n152_, new_n157_, new_n107_, new_n182_, new_n407_, new_n153_, new_n480_, new_n133_, new_n257_, new_n481_, new_n212_, new_n151_, new_n513_, new_n592_, new_n364_, new_n449_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n272_, new_n282_, new_n522_, new_n588_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n110_, new_n315_, new_n302_, new_n191_, new_n124_, new_n326_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n387_, new_n544_, new_n476_, new_n112_, new_n248_, new_n350_, new_n117_, new_n121_, new_n415_, new_n167_, new_n537_, new_n221_, new_n385_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n461_, new_n459_, new_n569_, new_n555_, new_n174_, new_n297_, new_n361_, new_n565_, new_n468_, new_n150_, new_n354_, new_n392_, new_n444_, new_n518_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n340_, new_n147_, new_n510_, new_n285_, new_n502_, new_n351_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n590_, new_n517_, new_n325_, new_n417_, new_n591_, new_n180_, new_n530_, new_n332_, new_n318_, new_n453_, new_n516_, new_n163_, new_n563_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n531_, new_n111_, new_n158_, new_n252_, new_n486_, new_n491_, new_n549_, new_n262_, new_n160_, new_n312_, new_n271_, new_n535_, new_n274_, new_n372_, new_n242_, new_n503_, new_n527_, new_n218_, new_n115_, new_n307_, new_n190_, new_n305_, new_n420_, new_n408_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n213_, new_n134_, new_n433_, new_n435_, new_n206_, new_n109_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n265_, new_n506_, new_n370_, new_n256_, new_n584_, new_n452_, new_n278_, new_n304_, new_n381_, new_n523_, new_n388_, new_n217_, new_n269_, new_n508_, new_n512_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n129_, new_n142_, new_n139_, new_n314_, new_n582_, new_n118_, new_n363_, new_n412_, new_n165_, new_n477_, new_n327_, new_n216_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n280_, new_n574_, new_n426_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n338_, new_n207_, new_n267_, new_n473_, new_n140_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n587_, new_n465_, new_n195_, new_n567_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n245_, new_n402_, new_n579_, new_n467_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n490_, new_n560_, new_n346_, new_n396_, new_n198_, new_n438_, new_n128_, new_n358_, new_n208_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n528_, new_n179_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n185_, new_n399_, new_n596_, new_n373_, new_n171_, new_n559_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n233_, new_n136_, new_n469_, new_n284_, new_n119_, new_n391_, new_n293_, new_n178_, new_n437_, new_n551_, new_n168_, new_n279_, new_n295_, new_n359_, new_n132_, new_n120_, new_n521_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n406_, new_n356_, new_n333_, new_n229_, new_n536_, new_n290_, new_n464_, new_n204_, new_n369_, new_n181_, new_n135_, new_n573_, new_n276_, new_n405_;

not g000 ( new_n106_, N81 );
not g001 ( new_n107_, N85 );
nand g002 ( new_n108_, new_n106_, new_n107_ );
nand g003 ( new_n109_, N81, N85 );
nand g004 ( new_n110_, new_n108_, new_n109_ );
not g005 ( new_n111_, N89 );
not g006 ( new_n112_, N93 );
nand g007 ( new_n113_, new_n111_, new_n112_ );
nand g008 ( new_n114_, N89, N93 );
nand g009 ( new_n115_, new_n113_, new_n114_ );
nand g010 ( new_n116_, new_n110_, new_n115_ );
nand g011 ( new_n117_, new_n108_, new_n113_, new_n109_, new_n114_ );
nand g012 ( new_n118_, new_n116_, new_n117_ );
nand g013 ( new_n119_, new_n118_, keyIn_0_5 );
not g014 ( new_n120_, keyIn_0_5 );
nand g015 ( new_n121_, new_n116_, new_n120_, new_n117_ );
nand g016 ( new_n122_, new_n119_, new_n121_ );
not g017 ( new_n123_, keyIn_0_7 );
not g018 ( new_n124_, N113 );
not g019 ( new_n125_, N117 );
nand g020 ( new_n126_, new_n124_, new_n125_ );
nand g021 ( new_n127_, N113, N117 );
nand g022 ( new_n128_, new_n126_, new_n127_ );
not g023 ( new_n129_, N121 );
not g024 ( new_n130_, N125 );
nand g025 ( new_n131_, new_n129_, new_n130_ );
nand g026 ( new_n132_, N121, N125 );
nand g027 ( new_n133_, new_n131_, new_n132_ );
nand g028 ( new_n134_, new_n128_, new_n133_ );
nand g029 ( new_n135_, new_n126_, new_n131_, new_n127_, new_n132_ );
nand g030 ( new_n136_, new_n134_, new_n135_ );
nand g031 ( new_n137_, new_n136_, new_n123_ );
nand g032 ( new_n138_, new_n134_, keyIn_0_7, new_n135_ );
nand g033 ( new_n139_, new_n137_, new_n138_ );
nand g034 ( new_n140_, new_n122_, new_n139_ );
nand g035 ( new_n141_, new_n119_, new_n137_, new_n121_, new_n138_ );
nand g036 ( new_n142_, new_n140_, new_n141_ );
nand g037 ( new_n143_, new_n142_, keyIn_0_23 );
not g038 ( new_n144_, keyIn_0_23 );
nand g039 ( new_n145_, new_n140_, new_n144_, new_n141_ );
nand g040 ( new_n146_, new_n143_, new_n145_ );
nand g041 ( new_n147_, N132, N137 );
not g042 ( new_n148_, new_n147_ );
nand g043 ( new_n149_, new_n146_, new_n148_ );
nand g044 ( new_n150_, new_n143_, new_n145_, new_n147_ );
nand g045 ( new_n151_, new_n149_, new_n150_ );
nand g046 ( new_n152_, new_n151_, keyIn_0_27 );
not g047 ( new_n153_, keyIn_0_27 );
nand g048 ( new_n154_, new_n149_, new_n153_, new_n150_ );
nand g049 ( new_n155_, new_n152_, new_n154_ );
xnor g050 ( new_n156_, N13, N29 );
xnor g051 ( new_n157_, N45, N61 );
xnor g052 ( new_n158_, new_n156_, new_n157_ );
xor g053 ( new_n159_, new_n158_, keyIn_0_11 );
not g054 ( new_n160_, new_n159_ );
nand g055 ( new_n161_, new_n155_, new_n160_ );
nand g056 ( new_n162_, new_n152_, new_n154_, new_n159_ );
nand g057 ( new_n163_, new_n161_, new_n162_ );
not g058 ( new_n164_, N65 );
not g059 ( new_n165_, N69 );
nand g060 ( new_n166_, new_n164_, new_n165_ );
nand g061 ( new_n167_, N65, N69 );
nand g062 ( new_n168_, new_n166_, new_n167_ );
xnor g063 ( new_n169_, N73, N77 );
nand g064 ( new_n170_, new_n168_, new_n169_ );
not g065 ( new_n171_, N73 );
not g066 ( new_n172_, N77 );
nand g067 ( new_n173_, new_n171_, new_n172_ );
nand g068 ( new_n174_, N73, N77 );
nand g069 ( new_n175_, new_n166_, new_n173_, new_n167_, new_n174_ );
nand g070 ( new_n176_, new_n170_, new_n175_ );
nand g071 ( new_n177_, new_n176_, keyIn_0_4 );
not g072 ( new_n178_, keyIn_0_4 );
nand g073 ( new_n179_, new_n170_, new_n178_, new_n175_ );
nand g074 ( new_n180_, new_n177_, new_n179_ );
not g075 ( new_n181_, keyIn_0_6 );
not g076 ( new_n182_, N97 );
not g077 ( new_n183_, N101 );
nand g078 ( new_n184_, new_n182_, new_n183_ );
nand g079 ( new_n185_, N97, N101 );
nand g080 ( new_n186_, new_n184_, new_n185_ );
xnor g081 ( new_n187_, N105, N109 );
nand g082 ( new_n188_, new_n186_, new_n187_ );
not g083 ( new_n189_, N105 );
not g084 ( new_n190_, N109 );
nand g085 ( new_n191_, new_n189_, new_n190_ );
nand g086 ( new_n192_, N105, N109 );
nand g087 ( new_n193_, new_n184_, new_n191_, new_n185_, new_n192_ );
nand g088 ( new_n194_, new_n188_, new_n193_ );
nand g089 ( new_n195_, new_n194_, new_n181_ );
nand g090 ( new_n196_, new_n188_, keyIn_0_6, new_n193_ );
nand g091 ( new_n197_, new_n195_, new_n196_ );
nand g092 ( new_n198_, new_n180_, new_n197_ );
nand g093 ( new_n199_, new_n177_, new_n195_, new_n179_, new_n196_ );
nand g094 ( new_n200_, new_n198_, new_n199_ );
nand g095 ( new_n201_, new_n200_, keyIn_0_22 );
not g096 ( new_n202_, keyIn_0_22 );
nand g097 ( new_n203_, new_n198_, new_n202_, new_n199_ );
nand g098 ( new_n204_, new_n201_, new_n203_ );
nand g099 ( new_n205_, N131, N137 );
not g100 ( new_n206_, new_n205_ );
nand g101 ( new_n207_, new_n204_, new_n206_ );
nand g102 ( new_n208_, new_n201_, new_n203_, new_n205_ );
nand g103 ( new_n209_, new_n207_, new_n208_ );
nand g104 ( new_n210_, new_n209_, keyIn_0_26 );
not g105 ( new_n211_, keyIn_0_26 );
nand g106 ( new_n212_, new_n207_, new_n211_, new_n208_ );
nand g107 ( new_n213_, new_n210_, new_n212_ );
xor g108 ( new_n214_, N9, N25 );
xnor g109 ( new_n215_, N41, N57 );
xnor g110 ( new_n216_, new_n214_, new_n215_ );
xor g111 ( new_n217_, new_n216_, keyIn_0_10 );
not g112 ( new_n218_, new_n217_ );
nand g113 ( new_n219_, new_n213_, new_n218_ );
nand g114 ( new_n220_, new_n210_, new_n212_, new_n217_ );
nand g115 ( new_n221_, new_n219_, new_n220_ );
nand g116 ( new_n222_, new_n122_, new_n180_ );
nand g117 ( new_n223_, new_n119_, new_n177_, new_n121_, new_n179_ );
nand g118 ( new_n224_, new_n222_, new_n223_ );
nand g119 ( new_n225_, new_n224_, keyIn_0_20 );
not g120 ( new_n226_, keyIn_0_20 );
nand g121 ( new_n227_, new_n222_, new_n226_, new_n223_ );
nand g122 ( new_n228_, new_n225_, new_n227_ );
nand g123 ( new_n229_, N129, N137 );
not g124 ( new_n230_, new_n229_ );
nand g125 ( new_n231_, new_n228_, new_n230_ );
nand g126 ( new_n232_, new_n225_, new_n227_, new_n229_ );
nand g127 ( new_n233_, new_n231_, new_n232_ );
nand g128 ( new_n234_, new_n233_, keyIn_0_24 );
not g129 ( new_n235_, keyIn_0_24 );
nand g130 ( new_n236_, new_n231_, new_n235_, new_n232_ );
nand g131 ( new_n237_, new_n234_, new_n236_ );
xnor g132 ( new_n238_, N1, N17 );
xnor g133 ( new_n239_, N33, N49 );
xnor g134 ( new_n240_, new_n238_, new_n239_ );
xnor g135 ( new_n241_, new_n240_, keyIn_0_8 );
not g136 ( new_n242_, new_n241_ );
nand g137 ( new_n243_, new_n237_, new_n242_ );
nand g138 ( new_n244_, new_n234_, new_n236_, new_n241_ );
nand g139 ( new_n245_, new_n243_, new_n244_ );
nand g140 ( new_n246_, new_n139_, new_n197_ );
nand g141 ( new_n247_, new_n137_, new_n195_, new_n138_, new_n196_ );
nand g142 ( new_n248_, new_n246_, new_n247_ );
nand g143 ( new_n249_, new_n248_, keyIn_0_21 );
not g144 ( new_n250_, keyIn_0_21 );
nand g145 ( new_n251_, new_n246_, new_n250_, new_n247_ );
nand g146 ( new_n252_, new_n249_, new_n251_ );
nand g147 ( new_n253_, N130, N137 );
not g148 ( new_n254_, new_n253_ );
nand g149 ( new_n255_, new_n252_, new_n254_ );
nand g150 ( new_n256_, new_n249_, new_n251_, new_n253_ );
nand g151 ( new_n257_, new_n255_, new_n256_ );
nand g152 ( new_n258_, new_n257_, keyIn_0_25 );
not g153 ( new_n259_, keyIn_0_25 );
nand g154 ( new_n260_, new_n255_, new_n259_, new_n256_ );
nand g155 ( new_n261_, new_n258_, new_n260_ );
xnor g156 ( new_n262_, N5, N21 );
xnor g157 ( new_n263_, N37, N53 );
xnor g158 ( new_n264_, new_n262_, new_n263_ );
xor g159 ( new_n265_, new_n264_, keyIn_0_9 );
nand g160 ( new_n266_, new_n261_, new_n265_ );
not g161 ( new_n267_, new_n265_ );
nand g162 ( new_n268_, new_n258_, new_n260_, new_n267_ );
nand g163 ( new_n269_, new_n266_, new_n268_ );
and g164 ( new_n270_, new_n163_, new_n221_, new_n245_, new_n269_ );
not g165 ( new_n271_, keyIn_0_1 );
not g166 ( new_n272_, N17 );
not g167 ( new_n273_, N21 );
nand g168 ( new_n274_, new_n272_, new_n273_ );
nand g169 ( new_n275_, N17, N21 );
nand g170 ( new_n276_, new_n274_, new_n275_ );
not g171 ( new_n277_, N25 );
not g172 ( new_n278_, N29 );
nand g173 ( new_n279_, new_n277_, new_n278_ );
nand g174 ( new_n280_, N25, N29 );
nand g175 ( new_n281_, new_n279_, new_n280_ );
nand g176 ( new_n282_, new_n276_, new_n281_ );
nand g177 ( new_n283_, new_n274_, new_n279_, new_n275_, new_n280_ );
nand g178 ( new_n284_, new_n282_, new_n283_ );
nand g179 ( new_n285_, new_n284_, new_n271_ );
nand g180 ( new_n286_, new_n282_, keyIn_0_1, new_n283_ );
nand g181 ( new_n287_, new_n285_, new_n286_ );
not g182 ( new_n288_, N49 );
not g183 ( new_n289_, N53 );
nand g184 ( new_n290_, new_n288_, new_n289_ );
nand g185 ( new_n291_, N49, N53 );
nand g186 ( new_n292_, new_n290_, new_n291_ );
not g187 ( new_n293_, N57 );
not g188 ( new_n294_, N61 );
nand g189 ( new_n295_, new_n293_, new_n294_ );
nand g190 ( new_n296_, N57, N61 );
nand g191 ( new_n297_, new_n295_, new_n296_ );
nand g192 ( new_n298_, new_n292_, new_n297_ );
nand g193 ( new_n299_, new_n290_, new_n295_, new_n291_, new_n296_ );
nand g194 ( new_n300_, new_n298_, new_n299_ );
nand g195 ( new_n301_, new_n300_, keyIn_0_3 );
not g196 ( new_n302_, keyIn_0_3 );
nand g197 ( new_n303_, new_n298_, new_n302_, new_n299_ );
nand g198 ( new_n304_, new_n301_, new_n303_ );
nand g199 ( new_n305_, new_n287_, new_n304_ );
nand g200 ( new_n306_, new_n285_, new_n301_, new_n286_, new_n303_ );
nand g201 ( new_n307_, new_n305_, new_n306_ );
nand g202 ( new_n308_, new_n307_, keyIn_0_19 );
not g203 ( new_n309_, keyIn_0_19 );
nand g204 ( new_n310_, new_n305_, new_n309_, new_n306_ );
nand g205 ( new_n311_, new_n308_, new_n310_ );
nand g206 ( new_n312_, N136, N137 );
nand g207 ( new_n313_, new_n311_, new_n312_ );
nand g208 ( new_n314_, new_n308_, N136, N137, new_n310_ );
nand g209 ( new_n315_, new_n313_, new_n314_ );
nand g210 ( new_n316_, new_n315_, keyIn_0_31 );
not g211 ( new_n317_, keyIn_0_31 );
nand g212 ( new_n318_, new_n313_, new_n317_, new_n314_ );
nand g213 ( new_n319_, new_n316_, new_n318_ );
xor g214 ( new_n320_, N77, N93 );
xnor g215 ( new_n321_, N109, N125 );
xnor g216 ( new_n322_, new_n320_, new_n321_ );
xor g217 ( new_n323_, new_n322_, keyIn_0_15 );
not g218 ( new_n324_, new_n323_ );
nand g219 ( new_n325_, new_n319_, new_n324_ );
nand g220 ( new_n326_, new_n316_, new_n318_, new_n323_ );
nand g221 ( new_n327_, new_n325_, new_n326_ );
not g222 ( new_n328_, keyIn_0_0 );
not g223 ( new_n329_, N1 );
not g224 ( new_n330_, N5 );
nand g225 ( new_n331_, new_n329_, new_n330_ );
nand g226 ( new_n332_, N1, N5 );
nand g227 ( new_n333_, new_n331_, new_n332_ );
xnor g228 ( new_n334_, N9, N13 );
nand g229 ( new_n335_, new_n333_, new_n334_ );
not g230 ( new_n336_, N9 );
not g231 ( new_n337_, N13 );
nand g232 ( new_n338_, new_n336_, new_n337_ );
nand g233 ( new_n339_, N9, N13 );
nand g234 ( new_n340_, new_n331_, new_n338_, new_n332_, new_n339_ );
nand g235 ( new_n341_, new_n335_, new_n340_ );
nand g236 ( new_n342_, new_n341_, new_n328_ );
nand g237 ( new_n343_, new_n335_, keyIn_0_0, new_n340_ );
nand g238 ( new_n344_, new_n342_, new_n343_ );
not g239 ( new_n345_, keyIn_0_2 );
not g240 ( new_n346_, N33 );
not g241 ( new_n347_, N37 );
nand g242 ( new_n348_, new_n346_, new_n347_ );
nand g243 ( new_n349_, N33, N37 );
nand g244 ( new_n350_, new_n348_, new_n349_ );
xnor g245 ( new_n351_, N41, N45 );
nand g246 ( new_n352_, new_n350_, new_n351_ );
not g247 ( new_n353_, N41 );
not g248 ( new_n354_, N45 );
nand g249 ( new_n355_, new_n353_, new_n354_ );
nand g250 ( new_n356_, N41, N45 );
nand g251 ( new_n357_, new_n348_, new_n355_, new_n349_, new_n356_ );
nand g252 ( new_n358_, new_n352_, new_n357_ );
nand g253 ( new_n359_, new_n358_, new_n345_ );
nand g254 ( new_n360_, new_n352_, keyIn_0_2, new_n357_ );
nand g255 ( new_n361_, new_n359_, new_n360_ );
nand g256 ( new_n362_, new_n344_, new_n361_ );
nand g257 ( new_n363_, new_n342_, new_n359_, new_n343_, new_n360_ );
nand g258 ( new_n364_, new_n362_, new_n363_ );
nand g259 ( new_n365_, new_n364_, keyIn_0_18 );
not g260 ( new_n366_, keyIn_0_18 );
nand g261 ( new_n367_, new_n362_, new_n366_, new_n363_ );
nand g262 ( new_n368_, new_n365_, new_n367_ );
nand g263 ( new_n369_, N135, N137 );
not g264 ( new_n370_, new_n369_ );
nand g265 ( new_n371_, new_n368_, new_n370_ );
nand g266 ( new_n372_, new_n365_, new_n367_, new_n369_ );
nand g267 ( new_n373_, new_n371_, new_n372_ );
nand g268 ( new_n374_, new_n373_, keyIn_0_30 );
not g269 ( new_n375_, keyIn_0_30 );
nand g270 ( new_n376_, new_n371_, new_n375_, new_n372_ );
nand g271 ( new_n377_, new_n374_, new_n376_ );
xnor g272 ( new_n378_, N73, N89 );
xnor g273 ( new_n379_, N105, N121 );
xnor g274 ( new_n380_, new_n378_, new_n379_ );
xnor g275 ( new_n381_, new_n380_, keyIn_0_14 );
not g276 ( new_n382_, new_n381_ );
nand g277 ( new_n383_, new_n377_, new_n382_ );
nand g278 ( new_n384_, new_n374_, new_n376_, new_n381_ );
nand g279 ( new_n385_, new_n383_, new_n384_ );
and g280 ( new_n386_, new_n327_, new_n385_ );
nand g281 ( new_n387_, new_n287_, new_n344_ );
nand g282 ( new_n388_, new_n285_, new_n342_, new_n286_, new_n343_ );
nand g283 ( new_n389_, new_n387_, new_n388_ );
nand g284 ( new_n390_, new_n389_, keyIn_0_16 );
not g285 ( new_n391_, keyIn_0_16 );
nand g286 ( new_n392_, new_n387_, new_n391_, new_n388_ );
nand g287 ( new_n393_, new_n390_, new_n392_ );
nand g288 ( new_n394_, N133, N137 );
not g289 ( new_n395_, new_n394_ );
nand g290 ( new_n396_, new_n393_, new_n395_ );
nand g291 ( new_n397_, new_n390_, new_n392_, new_n394_ );
nand g292 ( new_n398_, new_n396_, new_n397_ );
nand g293 ( new_n399_, new_n398_, keyIn_0_28 );
not g294 ( new_n400_, keyIn_0_28 );
nand g295 ( new_n401_, new_n396_, new_n400_, new_n397_ );
nand g296 ( new_n402_, new_n399_, new_n401_ );
xnor g297 ( new_n403_, N65, N81 );
xnor g298 ( new_n404_, N97, N113 );
xnor g299 ( new_n405_, new_n403_, new_n404_ );
xor g300 ( new_n406_, new_n405_, keyIn_0_12 );
not g301 ( new_n407_, new_n406_ );
nand g302 ( new_n408_, new_n402_, new_n407_ );
nand g303 ( new_n409_, new_n399_, new_n401_, new_n406_ );
nand g304 ( new_n410_, new_n408_, new_n409_ );
nand g305 ( new_n411_, new_n304_, new_n361_ );
nand g306 ( new_n412_, new_n301_, new_n359_, new_n303_, new_n360_ );
nand g307 ( new_n413_, new_n411_, new_n412_ );
nand g308 ( new_n414_, new_n413_, keyIn_0_17 );
not g309 ( new_n415_, keyIn_0_17 );
nand g310 ( new_n416_, new_n411_, new_n415_, new_n412_ );
nand g311 ( new_n417_, new_n414_, new_n416_ );
nand g312 ( new_n418_, N134, N137 );
not g313 ( new_n419_, new_n418_ );
nand g314 ( new_n420_, new_n417_, new_n419_ );
nand g315 ( new_n421_, new_n414_, new_n416_, new_n418_ );
nand g316 ( new_n422_, new_n420_, new_n421_ );
nand g317 ( new_n423_, new_n422_, keyIn_0_29 );
not g318 ( new_n424_, keyIn_0_29 );
nand g319 ( new_n425_, new_n420_, new_n424_, new_n421_ );
nand g320 ( new_n426_, new_n423_, new_n425_ );
xnor g321 ( new_n427_, N69, N85 );
xnor g322 ( new_n428_, N101, N117 );
xnor g323 ( new_n429_, new_n427_, new_n428_ );
xor g324 ( new_n430_, new_n429_, keyIn_0_13 );
not g325 ( new_n431_, new_n430_ );
nand g326 ( new_n432_, new_n426_, new_n431_ );
nand g327 ( new_n433_, new_n423_, new_n425_, new_n430_ );
nand g328 ( new_n434_, new_n432_, new_n433_ );
nor g329 ( new_n435_, new_n410_, new_n434_ );
nand g330 ( new_n436_, new_n270_, new_n386_, new_n435_ );
nand g331 ( new_n437_, new_n436_, N1 );
nand g332 ( new_n438_, new_n327_, new_n385_ );
nor g333 ( new_n439_, new_n438_, new_n410_, new_n434_ );
nand g334 ( new_n440_, new_n439_, new_n329_, new_n270_ );
nand g335 ( N724, new_n437_, new_n440_ );
and g336 ( new_n442_, new_n219_, new_n220_ );
nand g337 ( new_n443_, new_n243_, new_n266_, new_n244_, new_n268_ );
nor g338 ( new_n444_, new_n443_, new_n442_ );
nand g339 ( new_n445_, new_n444_, new_n163_, new_n386_, new_n435_ );
nand g340 ( new_n446_, new_n445_, N5 );
nand g341 ( new_n447_, new_n439_, new_n330_, new_n163_, new_n444_ );
nand g342 ( N725, new_n446_, new_n447_ );
and g343 ( new_n449_, new_n269_, new_n243_, new_n244_ );
and g344 ( new_n450_, new_n161_, new_n162_ );
nor g345 ( new_n451_, new_n450_, new_n221_ );
nand g346 ( new_n452_, new_n451_, new_n449_, new_n386_, new_n435_ );
nand g347 ( new_n453_, new_n452_, N9 );
nand g348 ( new_n454_, new_n439_, new_n336_, new_n449_, new_n451_ );
nand g349 ( N726, new_n453_, new_n454_ );
nor g350 ( new_n456_, new_n442_, new_n163_ );
nand g351 ( new_n457_, new_n449_, new_n456_, new_n386_, new_n435_ );
nand g352 ( new_n458_, new_n457_, N13 );
nand g353 ( new_n459_, new_n439_, new_n337_, new_n449_, new_n456_ );
nand g354 ( N727, new_n458_, new_n459_ );
nand g355 ( new_n461_, new_n325_, new_n383_, new_n326_, new_n384_ );
nor g356 ( new_n462_, new_n461_, new_n410_, new_n434_ );
nand g357 ( new_n463_, new_n270_, new_n462_ );
nand g358 ( new_n464_, new_n463_, N17 );
nand g359 ( new_n465_, new_n270_, new_n462_, new_n272_ );
nand g360 ( N728, new_n464_, new_n465_ );
nand g361 ( new_n467_, new_n462_, new_n163_, new_n444_ );
nand g362 ( new_n468_, new_n467_, N21 );
nand g363 ( new_n469_, new_n462_, new_n273_, new_n444_, new_n163_ );
nand g364 ( N729, new_n468_, new_n469_ );
nand g365 ( new_n471_, new_n462_, new_n449_, new_n451_ );
nand g366 ( new_n472_, new_n471_, N25 );
nand g367 ( new_n473_, new_n462_, new_n277_, new_n449_, new_n451_ );
nand g368 ( N730, new_n472_, new_n473_ );
nand g369 ( new_n475_, new_n462_, new_n449_, new_n456_ );
nand g370 ( new_n476_, new_n475_, N29 );
nand g371 ( new_n477_, new_n462_, new_n278_, new_n449_, new_n456_ );
nand g372 ( N731, new_n476_, new_n477_ );
nand g373 ( new_n479_, new_n410_, new_n434_ );
nor g374 ( new_n480_, new_n438_, new_n479_ );
nand g375 ( new_n481_, new_n480_, new_n270_ );
nand g376 ( new_n482_, new_n481_, N33 );
nand g377 ( new_n483_, new_n480_, new_n270_, new_n346_ );
nand g378 ( N732, new_n482_, new_n483_ );
and g379 ( new_n485_, new_n410_, new_n434_ );
nand g380 ( new_n486_, new_n444_, new_n163_, new_n386_, new_n485_ );
nand g381 ( new_n487_, new_n486_, N37 );
nand g382 ( new_n488_, new_n480_, new_n347_, new_n163_, new_n444_ );
nand g383 ( N733, new_n487_, new_n488_ );
nand g384 ( new_n490_, new_n451_, new_n449_, new_n386_, new_n485_ );
nand g385 ( new_n491_, new_n490_, N41 );
nand g386 ( new_n492_, new_n480_, new_n353_, new_n449_, new_n451_ );
nand g387 ( N734, new_n491_, new_n492_ );
nand g388 ( new_n494_, new_n449_, new_n456_, new_n386_, new_n485_ );
nand g389 ( new_n495_, new_n494_, N45 );
nand g390 ( new_n496_, new_n480_, new_n354_, new_n449_, new_n456_ );
nand g391 ( N735, new_n495_, new_n496_ );
and g392 ( new_n498_, new_n221_, new_n245_, new_n269_ );
and g393 ( new_n499_, new_n408_, new_n409_ );
nor g394 ( new_n500_, new_n461_, new_n499_ );
not g395 ( new_n501_, new_n434_ );
nor g396 ( new_n502_, new_n501_, new_n450_ );
nand g397 ( new_n503_, new_n502_, new_n500_, new_n498_ );
nand g398 ( new_n504_, new_n503_, N49 );
nor g399 ( new_n505_, new_n479_, new_n461_ );
nand g400 ( new_n506_, new_n270_, new_n505_, new_n288_ );
nand g401 ( N736, new_n504_, new_n506_ );
nand g402 ( new_n508_, new_n502_, new_n444_, new_n500_ );
nand g403 ( new_n509_, new_n508_, N53 );
nand g404 ( new_n510_, new_n505_, new_n289_, new_n444_, new_n163_ );
nand g405 ( N737, new_n509_, new_n510_ );
nand g406 ( new_n512_, new_n500_, new_n451_, new_n449_, new_n434_ );
nand g407 ( new_n513_, new_n512_, N57 );
nand g408 ( new_n514_, new_n505_, new_n293_, new_n449_, new_n451_ );
nand g409 ( N738, new_n513_, new_n514_ );
nand g410 ( new_n516_, new_n500_, new_n449_, new_n456_, new_n434_ );
nand g411 ( new_n517_, new_n516_, N61 );
nand g412 ( new_n518_, new_n505_, new_n294_, new_n449_, new_n456_ );
nand g413 ( N739, new_n517_, new_n518_ );
nand g414 ( new_n520_, new_n245_, new_n269_ );
not g415 ( new_n521_, new_n520_ );
and g416 ( new_n522_, new_n325_, new_n326_ );
nor g417 ( new_n523_, new_n522_, new_n385_ );
nand g418 ( new_n524_, new_n451_, new_n523_, new_n521_, new_n435_ );
nand g419 ( new_n525_, new_n524_, N65 );
nor g420 ( new_n526_, new_n520_, new_n450_, new_n221_ );
nor g421 ( new_n527_, new_n522_, new_n385_, new_n410_, new_n434_ );
nand g422 ( new_n528_, new_n527_, new_n164_, new_n526_ );
nand g423 ( N740, new_n525_, new_n528_ );
nand g424 ( new_n530_, new_n451_, new_n523_, new_n521_, new_n485_ );
nand g425 ( new_n531_, new_n530_, N69 );
nor g426 ( new_n532_, new_n479_, new_n522_, new_n385_ );
nand g427 ( new_n533_, new_n526_, new_n532_, new_n165_ );
nand g428 ( N741, new_n531_, new_n533_ );
nor g429 ( new_n535_, new_n499_, new_n434_ );
nand g430 ( new_n536_, new_n521_, new_n451_, new_n535_, new_n386_ );
nand g431 ( new_n537_, new_n536_, N73 );
nor g432 ( new_n538_, new_n438_, new_n499_, new_n434_ );
nand g433 ( new_n539_, new_n526_, new_n538_, new_n171_ );
nand g434 ( N742, new_n537_, new_n539_ );
nand g435 ( new_n541_, new_n500_, new_n451_, new_n521_, new_n501_ );
nand g436 ( new_n542_, new_n541_, N77 );
nor g437 ( new_n543_, new_n461_, new_n499_, new_n434_ );
nand g438 ( new_n544_, new_n526_, new_n543_, new_n172_ );
nand g439 ( N743, new_n542_, new_n544_ );
nand g440 ( new_n546_, new_n498_, new_n523_, new_n450_, new_n435_ );
nand g441 ( new_n547_, new_n546_, N81 );
nor g442 ( new_n548_, new_n520_, new_n163_, new_n442_ );
nand g443 ( new_n549_, new_n527_, new_n106_, new_n548_ );
nand g444 ( N744, new_n547_, new_n549_ );
nand g445 ( new_n551_, new_n498_, new_n523_, new_n485_, new_n450_ );
nand g446 ( new_n552_, new_n551_, N85 );
nand g447 ( new_n553_, new_n532_, new_n548_, new_n107_ );
nand g448 ( N745, new_n552_, new_n553_ );
nand g449 ( new_n555_, new_n498_, new_n535_, new_n386_, new_n450_ );
nand g450 ( new_n556_, new_n555_, N89 );
nand g451 ( new_n557_, new_n538_, new_n548_, new_n111_ );
nand g452 ( N746, new_n556_, new_n557_ );
nand g453 ( new_n559_, new_n500_, new_n498_, new_n450_, new_n501_ );
nand g454 ( new_n560_, new_n559_, N93 );
nand g455 ( new_n561_, new_n548_, new_n543_, new_n112_ );
nand g456 ( N747, new_n560_, new_n561_ );
not g457 ( new_n563_, new_n443_ );
nand g458 ( new_n564_, new_n451_, new_n523_, new_n435_, new_n563_ );
nand g459 ( new_n565_, new_n564_, N97 );
nor g460 ( new_n566_, new_n443_, new_n450_, new_n221_ );
nand g461 ( new_n567_, new_n527_, new_n566_, new_n182_ );
nand g462 ( N748, new_n565_, new_n567_ );
nand g463 ( new_n569_, new_n451_, new_n523_, new_n485_, new_n563_ );
nand g464 ( new_n570_, new_n569_, N101 );
nand g465 ( new_n571_, new_n532_, new_n566_, new_n183_ );
nand g466 ( N749, new_n570_, new_n571_ );
nand g467 ( new_n573_, new_n451_, new_n535_, new_n386_, new_n563_ );
nand g468 ( new_n574_, new_n573_, N105 );
nand g469 ( new_n575_, new_n538_, new_n566_, new_n189_ );
nand g470 ( N750, new_n574_, new_n575_ );
nand g471 ( new_n577_, new_n500_, new_n451_, new_n501_, new_n563_ );
nand g472 ( new_n578_, new_n577_, N109 );
nand g473 ( new_n579_, new_n566_, new_n543_, new_n190_ );
nand g474 ( N751, new_n578_, new_n579_ );
nand g475 ( new_n581_, new_n444_, new_n523_, new_n450_, new_n435_ );
nand g476 ( new_n582_, new_n581_, N113 );
nor g477 ( new_n583_, new_n443_, new_n442_, new_n163_ );
nand g478 ( new_n584_, new_n527_, new_n583_, new_n124_ );
nand g479 ( N752, new_n582_, new_n584_ );
nand g480 ( new_n586_, new_n444_, new_n523_, new_n450_, new_n485_ );
nand g481 ( new_n587_, new_n586_, N117 );
nand g482 ( new_n588_, new_n532_, new_n583_, new_n125_ );
nand g483 ( N753, new_n587_, new_n588_ );
nand g484 ( new_n590_, new_n444_, new_n535_, new_n386_, new_n450_ );
nand g485 ( new_n591_, new_n590_, N121 );
nand g486 ( new_n592_, new_n538_, new_n583_, new_n129_ );
nand g487 ( N754, new_n591_, new_n592_ );
nand g488 ( new_n594_, new_n444_, new_n500_, new_n450_, new_n501_ );
nand g489 ( new_n595_, new_n594_, N125 );
nand g490 ( new_n596_, new_n543_, new_n583_, new_n130_ );
nand g491 ( N755, new_n595_, new_n596_ );
endmodule