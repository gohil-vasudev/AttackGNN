module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n368_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n844_, new_n482_, new_n849_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n851_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n825_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n480_, new_n625_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n148_, new_n662_, new_n440_, new_n733_, new_n531_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n435_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n138_, N1 );
not g001 ( new_n139_, keyIn_0_41 );
not g002 ( new_n140_, N81 );
not g003 ( new_n141_, N85 );
nand g004 ( new_n142_, new_n140_, new_n141_ );
nand g005 ( new_n143_, N81, N85 );
nand g006 ( new_n144_, new_n142_, new_n143_ );
not g007 ( new_n145_, N89 );
not g008 ( new_n146_, N93 );
nand g009 ( new_n147_, new_n145_, new_n146_ );
nand g010 ( new_n148_, N89, N93 );
nand g011 ( new_n149_, new_n147_, new_n148_ );
nand g012 ( new_n150_, new_n144_, new_n149_ );
nand g013 ( new_n151_, new_n142_, new_n147_, new_n143_, new_n148_ );
nand g014 ( new_n152_, new_n150_, new_n151_ );
not g015 ( new_n153_, new_n152_ );
nor g016 ( new_n154_, N73, N77 );
not g017 ( new_n155_, new_n154_ );
nand g018 ( new_n156_, N73, N77 );
nand g019 ( new_n157_, new_n155_, new_n156_ );
not g020 ( new_n158_, N65 );
not g021 ( new_n159_, N69 );
nand g022 ( new_n160_, new_n158_, new_n159_ );
nand g023 ( new_n161_, N65, N69 );
not g024 ( new_n162_, keyIn_0_6 );
nand g025 ( new_n163_, new_n162_, keyIn_0_5 );
not g026 ( new_n164_, keyIn_0_5 );
nand g027 ( new_n165_, new_n164_, keyIn_0_6 );
nand g028 ( new_n166_, new_n160_, new_n163_, new_n165_, new_n161_ );
nand g029 ( new_n167_, new_n160_, new_n161_ );
nand g030 ( new_n168_, new_n163_, new_n165_ );
nand g031 ( new_n169_, new_n167_, new_n168_ );
nand g032 ( new_n170_, new_n169_, new_n157_, new_n166_ );
nand g033 ( new_n171_, new_n169_, new_n166_ );
nand g034 ( new_n172_, new_n171_, new_n155_, new_n156_ );
nand g035 ( new_n173_, new_n172_, new_n170_ );
nand g036 ( new_n174_, new_n173_, new_n153_ );
not g037 ( new_n175_, new_n173_ );
nand g038 ( new_n176_, new_n175_, new_n152_ );
nand g039 ( new_n177_, new_n176_, new_n174_ );
nand g040 ( new_n178_, N129, N137 );
nand g041 ( new_n179_, new_n177_, new_n178_ );
nand g042 ( new_n180_, new_n176_, N129, N137, new_n174_ );
not g043 ( new_n181_, N17 );
nand g044 ( new_n182_, new_n181_, N1 );
nand g045 ( new_n183_, new_n138_, N17 );
nand g046 ( new_n184_, new_n182_, new_n183_ );
not g047 ( new_n185_, N33 );
not g048 ( new_n186_, N49 );
nand g049 ( new_n187_, new_n185_, new_n186_ );
nand g050 ( new_n188_, N33, N49 );
nand g051 ( new_n189_, new_n187_, new_n188_ );
nand g052 ( new_n190_, new_n184_, new_n189_ );
nand g053 ( new_n191_, new_n187_, new_n182_, new_n183_, new_n188_ );
nand g054 ( new_n192_, new_n190_, new_n191_ );
nand g055 ( new_n193_, new_n179_, new_n180_, new_n192_ );
nand g056 ( new_n194_, new_n179_, new_n180_ );
nand g057 ( new_n195_, new_n194_, new_n190_, new_n191_ );
nand g058 ( new_n196_, new_n195_, new_n193_ );
not g059 ( new_n197_, N117 );
nand g060 ( new_n198_, new_n197_, N113 );
not g061 ( new_n199_, N113 );
nand g062 ( new_n200_, new_n199_, N117 );
nand g063 ( new_n201_, new_n198_, new_n200_ );
nand g064 ( new_n202_, new_n201_, keyIn_0_7 );
not g065 ( new_n203_, keyIn_0_7 );
nand g066 ( new_n204_, new_n198_, new_n200_, new_n203_ );
nand g067 ( new_n205_, new_n202_, new_n204_ );
not g068 ( new_n206_, N121 );
not g069 ( new_n207_, N125 );
nand g070 ( new_n208_, new_n206_, new_n207_ );
nand g071 ( new_n209_, N121, N125 );
nand g072 ( new_n210_, new_n208_, new_n209_ );
nand g073 ( new_n211_, new_n205_, new_n210_ );
nand g074 ( new_n212_, new_n202_, new_n204_, new_n208_, new_n209_ );
nand g075 ( new_n213_, new_n211_, new_n212_ );
nand g076 ( new_n214_, new_n213_, keyIn_0_19 );
not g077 ( new_n215_, keyIn_0_19 );
nand g078 ( new_n216_, new_n211_, new_n215_, new_n212_ );
not g079 ( new_n217_, N101 );
nand g080 ( new_n218_, new_n217_, N97 );
not g081 ( new_n219_, N97 );
nand g082 ( new_n220_, new_n219_, N101 );
nand g083 ( new_n221_, new_n218_, new_n220_ );
not g084 ( new_n222_, N105 );
not g085 ( new_n223_, N109 );
nand g086 ( new_n224_, new_n222_, new_n223_ );
nand g087 ( new_n225_, N105, N109 );
nand g088 ( new_n226_, new_n224_, new_n225_ );
nand g089 ( new_n227_, new_n221_, new_n226_ );
nand g090 ( new_n228_, new_n224_, new_n218_, new_n220_, new_n225_ );
nand g091 ( new_n229_, new_n227_, new_n228_ );
nand g092 ( new_n230_, new_n229_, keyIn_0_18 );
not g093 ( new_n231_, keyIn_0_18 );
nand g094 ( new_n232_, new_n227_, new_n231_, new_n228_ );
nand g095 ( new_n233_, new_n230_, new_n232_ );
not g096 ( new_n234_, new_n233_ );
nand g097 ( new_n235_, new_n214_, new_n234_, new_n216_ );
nand g098 ( new_n236_, new_n214_, new_n216_ );
nand g099 ( new_n237_, new_n236_, new_n233_ );
nand g100 ( new_n238_, new_n237_, new_n235_ );
nand g101 ( new_n239_, new_n238_, keyIn_0_22 );
not g102 ( new_n240_, keyIn_0_22 );
nand g103 ( new_n241_, new_n237_, new_n240_, new_n235_ );
nand g104 ( new_n242_, new_n239_, new_n241_ );
nand g105 ( new_n243_, new_n242_, keyIn_0_8 );
not g106 ( new_n244_, keyIn_0_8 );
nand g107 ( new_n245_, new_n239_, new_n244_, new_n241_ );
nand g108 ( new_n246_, new_n243_, new_n245_ );
nand g109 ( new_n247_, N130, N137 );
nand g110 ( new_n248_, new_n246_, new_n247_ );
nand g111 ( new_n249_, new_n243_, N130, N137, new_n245_ );
not g112 ( new_n250_, N21 );
nand g113 ( new_n251_, new_n250_, N5 );
not g114 ( new_n252_, N5 );
nand g115 ( new_n253_, new_n252_, N21 );
nand g116 ( new_n254_, new_n251_, new_n253_ );
nand g117 ( new_n255_, new_n254_, keyIn_0_12 );
not g118 ( new_n256_, keyIn_0_12 );
nand g119 ( new_n257_, new_n251_, new_n253_, new_n256_ );
nand g120 ( new_n258_, new_n255_, new_n257_ );
not g121 ( new_n259_, N53 );
nand g122 ( new_n260_, new_n259_, N37 );
not g123 ( new_n261_, N37 );
nand g124 ( new_n262_, new_n261_, N53 );
nand g125 ( new_n263_, new_n260_, new_n262_ );
nand g126 ( new_n264_, new_n263_, keyIn_0_13 );
not g127 ( new_n265_, keyIn_0_13 );
nand g128 ( new_n266_, new_n260_, new_n262_, new_n265_ );
nand g129 ( new_n267_, new_n264_, new_n266_ );
nand g130 ( new_n268_, new_n258_, new_n267_ );
nand g131 ( new_n269_, new_n255_, new_n264_, new_n257_, new_n266_ );
nand g132 ( new_n270_, new_n248_, new_n249_, new_n268_, new_n269_ );
nand g133 ( new_n271_, new_n248_, new_n249_ );
nand g134 ( new_n272_, new_n268_, new_n269_ );
nand g135 ( new_n273_, new_n271_, new_n272_ );
nand g136 ( new_n274_, new_n273_, new_n196_, new_n270_ );
not g137 ( new_n275_, new_n274_ );
not g138 ( new_n276_, keyIn_0_9 );
nand g139 ( new_n277_, new_n236_, new_n152_ );
nand g140 ( new_n278_, new_n214_, new_n153_, new_n216_ );
nand g141 ( new_n279_, new_n277_, new_n276_, new_n278_ );
nand g142 ( new_n280_, new_n277_, new_n278_ );
nand g143 ( new_n281_, new_n280_, keyIn_0_9 );
nand g144 ( new_n282_, new_n281_, new_n279_ );
nand g145 ( new_n283_, N132, N137 );
nand g146 ( new_n284_, new_n282_, new_n283_ );
nand g147 ( new_n285_, new_n281_, N132, N137, new_n279_ );
nand g148 ( new_n286_, new_n284_, new_n285_ );
nand g149 ( new_n287_, new_n286_, keyIn_0_23 );
not g150 ( new_n288_, keyIn_0_23 );
nand g151 ( new_n289_, new_n284_, new_n288_, new_n285_ );
not g152 ( new_n290_, N29 );
nand g153 ( new_n291_, new_n290_, N13 );
not g154 ( new_n292_, N13 );
nand g155 ( new_n293_, new_n292_, N29 );
nand g156 ( new_n294_, new_n291_, new_n293_ );
nand g157 ( new_n295_, new_n294_, keyIn_0_14 );
not g158 ( new_n296_, keyIn_0_14 );
nand g159 ( new_n297_, new_n291_, new_n293_, new_n296_ );
nand g160 ( new_n298_, new_n295_, new_n297_ );
not g161 ( new_n299_, N45 );
nor g162 ( new_n300_, new_n299_, N61 );
not g163 ( new_n301_, N61 );
nor g164 ( new_n302_, new_n301_, N45 );
nor g165 ( new_n303_, new_n300_, new_n302_ );
not g166 ( new_n304_, new_n303_ );
nand g167 ( new_n305_, new_n298_, new_n304_ );
nand g168 ( new_n306_, new_n295_, new_n297_, new_n303_ );
nand g169 ( new_n307_, new_n287_, new_n289_, new_n305_, new_n306_ );
nand g170 ( new_n308_, new_n287_, new_n289_ );
nand g171 ( new_n309_, new_n305_, new_n306_ );
nand g172 ( new_n310_, new_n308_, new_n309_ );
nand g173 ( new_n311_, new_n310_, new_n307_ );
not g174 ( new_n312_, keyIn_0_26 );
nand g175 ( new_n313_, new_n234_, new_n173_ );
nand g176 ( new_n314_, new_n175_, new_n233_ );
nand g177 ( new_n315_, new_n314_, new_n313_ );
nand g178 ( new_n316_, N131, N137 );
nand g179 ( new_n317_, new_n315_, new_n316_ );
nand g180 ( new_n318_, new_n314_, new_n313_, N131, N137 );
nand g181 ( new_n319_, new_n317_, new_n318_ );
not g182 ( new_n320_, N9 );
not g183 ( new_n321_, N25 );
nand g184 ( new_n322_, new_n320_, new_n321_ );
nand g185 ( new_n323_, N9, N25 );
nand g186 ( new_n324_, new_n322_, new_n323_ );
not g187 ( new_n325_, N41 );
not g188 ( new_n326_, N57 );
nand g189 ( new_n327_, new_n325_, new_n326_ );
nand g190 ( new_n328_, N41, N57 );
nand g191 ( new_n329_, new_n327_, new_n328_ );
nand g192 ( new_n330_, new_n324_, new_n329_ );
nand g193 ( new_n331_, new_n322_, new_n327_, new_n323_, new_n328_ );
nand g194 ( new_n332_, new_n330_, new_n331_ );
nand g195 ( new_n333_, new_n319_, new_n332_ );
nand g196 ( new_n334_, new_n317_, new_n318_, new_n330_, new_n331_ );
nand g197 ( new_n335_, new_n333_, new_n334_ );
nand g198 ( new_n336_, new_n335_, keyIn_0_24 );
not g199 ( new_n337_, keyIn_0_24 );
nand g200 ( new_n338_, new_n333_, new_n337_, new_n334_ );
nand g201 ( new_n339_, new_n336_, new_n312_, new_n338_ );
nand g202 ( new_n340_, new_n336_, new_n338_ );
nand g203 ( new_n341_, new_n340_, keyIn_0_26 );
nand g204 ( new_n342_, new_n341_, new_n339_ );
nor g205 ( new_n343_, new_n311_, new_n342_ );
nand g206 ( new_n344_, new_n343_, new_n275_, keyIn_0_36 );
not g207 ( new_n345_, keyIn_0_36 );
nand g208 ( new_n346_, new_n343_, new_n275_ );
nand g209 ( new_n347_, new_n346_, new_n345_ );
nand g210 ( new_n348_, new_n347_, new_n344_ );
not g211 ( new_n349_, new_n311_ );
nand g212 ( new_n350_, new_n273_, new_n270_ );
not g213 ( new_n351_, new_n196_ );
nand g214 ( new_n352_, new_n340_, new_n351_ );
not g215 ( new_n353_, new_n352_ );
nand g216 ( new_n354_, new_n350_, new_n353_ );
not g217 ( new_n355_, new_n350_ );
not g218 ( new_n356_, new_n340_ );
nand g219 ( new_n357_, new_n351_, keyIn_0_25 );
not g220 ( new_n358_, keyIn_0_25 );
nand g221 ( new_n359_, new_n196_, new_n358_ );
nand g222 ( new_n360_, new_n357_, new_n359_ );
not g223 ( new_n361_, new_n360_ );
nand g224 ( new_n362_, new_n355_, new_n356_, new_n361_ );
nand g225 ( new_n363_, new_n362_, new_n354_ );
nand g226 ( new_n364_, new_n363_, new_n349_ );
nand g227 ( new_n365_, new_n355_, new_n311_, new_n353_ );
nand g228 ( new_n366_, new_n348_, new_n364_, new_n365_ );
not g229 ( new_n367_, keyIn_0_21 );
not g230 ( new_n368_, keyIn_0_17 );
nand g231 ( new_n369_, new_n185_, keyIn_0_2 );
not g232 ( new_n370_, keyIn_0_2 );
nand g233 ( new_n371_, new_n370_, N33 );
nand g234 ( new_n372_, new_n369_, new_n371_ );
nand g235 ( new_n373_, new_n372_, new_n261_ );
nand g236 ( new_n374_, new_n369_, new_n371_, N37 );
nand g237 ( new_n375_, new_n373_, new_n374_ );
nor g238 ( new_n376_, N41, N45 );
not g239 ( new_n377_, new_n376_ );
nand g240 ( new_n378_, N41, N45 );
nand g241 ( new_n379_, new_n377_, new_n378_ );
nand g242 ( new_n380_, new_n379_, keyIn_0_3 );
not g243 ( new_n381_, keyIn_0_3 );
nand g244 ( new_n382_, new_n377_, new_n381_, new_n378_ );
nand g245 ( new_n383_, new_n380_, new_n382_ );
nand g246 ( new_n384_, new_n383_, new_n375_ );
nand g247 ( new_n385_, new_n380_, new_n373_, new_n374_, new_n382_ );
nand g248 ( new_n386_, new_n384_, new_n385_ );
nand g249 ( new_n387_, new_n386_, new_n368_ );
nand g250 ( new_n388_, new_n384_, keyIn_0_17, new_n385_ );
nand g251 ( new_n389_, new_n387_, new_n388_ );
not g252 ( new_n390_, keyIn_0_16 );
nand g253 ( new_n391_, new_n252_, N1 );
nand g254 ( new_n392_, new_n138_, N5 );
nand g255 ( new_n393_, new_n391_, new_n392_ );
nand g256 ( new_n394_, new_n320_, new_n292_ );
nand g257 ( new_n395_, N9, N13 );
nand g258 ( new_n396_, new_n394_, new_n395_ );
nand g259 ( new_n397_, new_n393_, new_n396_ );
nand g260 ( new_n398_, new_n394_, new_n391_, new_n392_, new_n395_ );
nand g261 ( new_n399_, new_n397_, new_n390_, new_n398_ );
nand g262 ( new_n400_, new_n397_, new_n398_ );
nand g263 ( new_n401_, new_n400_, keyIn_0_16 );
nand g264 ( new_n402_, new_n401_, new_n399_ );
not g265 ( new_n403_, new_n402_ );
nand g266 ( new_n404_, new_n389_, new_n403_ );
nand g267 ( new_n405_, new_n387_, new_n388_, new_n402_ );
nand g268 ( new_n406_, new_n404_, new_n405_ );
nand g269 ( new_n407_, new_n406_, new_n367_ );
nand g270 ( new_n408_, new_n404_, keyIn_0_21, new_n405_ );
nand g271 ( new_n409_, new_n407_, new_n408_ );
not g272 ( new_n410_, keyIn_0_10 );
nand g273 ( new_n411_, new_n410_, N135, N137 );
nand g274 ( new_n412_, N135, N137 );
nand g275 ( new_n413_, new_n412_, keyIn_0_10 );
nand g276 ( new_n414_, new_n413_, new_n411_ );
nand g277 ( new_n415_, new_n409_, new_n414_ );
nand g278 ( new_n416_, new_n407_, new_n408_, new_n411_, new_n413_ );
nand g279 ( new_n417_, new_n415_, new_n416_ );
not g280 ( new_n418_, keyIn_0_20 );
nand g281 ( new_n419_, new_n145_, N73 );
not g282 ( new_n420_, N73 );
nand g283 ( new_n421_, new_n420_, N89 );
nand g284 ( new_n422_, new_n419_, new_n421_ );
nand g285 ( new_n423_, new_n222_, new_n206_ );
nand g286 ( new_n424_, N105, N121 );
nand g287 ( new_n425_, new_n423_, new_n424_ );
nand g288 ( new_n426_, new_n422_, new_n425_ );
nand g289 ( new_n427_, new_n423_, new_n419_, new_n421_, new_n424_ );
nand g290 ( new_n428_, new_n426_, new_n427_ );
nand g291 ( new_n429_, new_n428_, new_n418_ );
nand g292 ( new_n430_, new_n426_, keyIn_0_20, new_n427_ );
nand g293 ( new_n431_, new_n429_, new_n430_ );
nand g294 ( new_n432_, new_n417_, new_n431_ );
nand g295 ( new_n433_, new_n415_, new_n416_, new_n429_, new_n430_ );
nand g296 ( new_n434_, new_n432_, new_n433_ );
nor g297 ( new_n435_, N49, N53 );
not g298 ( new_n436_, new_n435_ );
nand g299 ( new_n437_, N49, N53 );
nand g300 ( new_n438_, new_n436_, new_n437_ );
nand g301 ( new_n439_, new_n438_, keyIn_0_4 );
not g302 ( new_n440_, keyIn_0_4 );
nand g303 ( new_n441_, new_n436_, new_n440_, new_n437_ );
nand g304 ( new_n442_, new_n439_, new_n441_ );
nor g305 ( new_n443_, N57, N61 );
not g306 ( new_n444_, new_n443_ );
nand g307 ( new_n445_, N57, N61 );
nand g308 ( new_n446_, new_n444_, new_n445_ );
nand g309 ( new_n447_, new_n442_, new_n446_ );
nand g310 ( new_n448_, new_n439_, new_n441_, new_n444_, new_n445_ );
nand g311 ( new_n449_, new_n447_, new_n448_ );
nand g312 ( new_n450_, new_n389_, new_n449_ );
nand g313 ( new_n451_, new_n387_, new_n388_, new_n447_, new_n448_ );
nand g314 ( new_n452_, new_n450_, new_n451_ );
nand g315 ( new_n453_, N134, N137 );
nand g316 ( new_n454_, new_n452_, new_n453_ );
nand g317 ( new_n455_, new_n450_, N134, N137, new_n451_ );
nand g318 ( new_n456_, new_n159_, new_n141_ );
nand g319 ( new_n457_, N69, N85 );
nand g320 ( new_n458_, new_n456_, new_n457_ );
nand g321 ( new_n459_, new_n217_, new_n197_ );
nand g322 ( new_n460_, N101, N117 );
nand g323 ( new_n461_, new_n459_, new_n460_ );
nand g324 ( new_n462_, new_n458_, new_n461_ );
nand g325 ( new_n463_, new_n456_, new_n459_, new_n457_, new_n460_ );
nand g326 ( new_n464_, new_n454_, new_n455_, new_n462_, new_n463_ );
nand g327 ( new_n465_, new_n454_, new_n455_ );
nand g328 ( new_n466_, new_n462_, new_n463_ );
nand g329 ( new_n467_, new_n465_, new_n466_ );
nand g330 ( new_n468_, new_n467_, new_n464_ );
not g331 ( new_n469_, new_n468_ );
nor g332 ( new_n470_, N25, N29 );
not g333 ( new_n471_, new_n470_ );
nand g334 ( new_n472_, N25, N29 );
nand g335 ( new_n473_, new_n471_, new_n472_ );
nand g336 ( new_n474_, new_n473_, keyIn_0_1 );
not g337 ( new_n475_, keyIn_0_1 );
nand g338 ( new_n476_, new_n471_, new_n475_, new_n472_ );
nor g339 ( new_n477_, N17, N21 );
not g340 ( new_n478_, new_n477_ );
nand g341 ( new_n479_, N17, N21 );
nand g342 ( new_n480_, new_n478_, new_n479_ );
nand g343 ( new_n481_, new_n480_, keyIn_0_0 );
not g344 ( new_n482_, keyIn_0_0 );
nand g345 ( new_n483_, new_n478_, new_n482_, new_n479_ );
nand g346 ( new_n484_, new_n474_, new_n481_, new_n476_, new_n483_ );
nand g347 ( new_n485_, new_n474_, new_n476_ );
nand g348 ( new_n486_, new_n481_, new_n483_ );
nand g349 ( new_n487_, new_n485_, new_n486_ );
nand g350 ( new_n488_, new_n402_, new_n484_, new_n487_ );
nand g351 ( new_n489_, new_n487_, new_n484_ );
nand g352 ( new_n490_, new_n403_, new_n489_ );
nand g353 ( new_n491_, new_n490_, new_n488_ );
nand g354 ( new_n492_, N133, N137 );
nand g355 ( new_n493_, new_n491_, new_n492_ );
nand g356 ( new_n494_, new_n490_, new_n488_, N133, N137 );
nand g357 ( new_n495_, new_n493_, new_n494_ );
nor g358 ( new_n496_, N97, N113 );
not g359 ( new_n497_, new_n496_ );
nand g360 ( new_n498_, N97, N113 );
nand g361 ( new_n499_, new_n497_, new_n498_ );
nand g362 ( new_n500_, new_n499_, keyIn_0_15 );
not g363 ( new_n501_, new_n500_ );
nor g364 ( new_n502_, new_n499_, keyIn_0_15 );
nor g365 ( new_n503_, new_n501_, new_n502_ );
not g366 ( new_n504_, new_n503_ );
nor g367 ( new_n505_, N65, N81 );
nand g368 ( new_n506_, N65, N81 );
not g369 ( new_n507_, new_n506_ );
nor g370 ( new_n508_, new_n507_, new_n505_ );
not g371 ( new_n509_, new_n508_ );
nand g372 ( new_n510_, new_n504_, new_n509_ );
nand g373 ( new_n511_, new_n503_, new_n508_ );
nand g374 ( new_n512_, new_n510_, new_n511_ );
nand g375 ( new_n513_, new_n495_, new_n512_ );
nand g376 ( new_n514_, new_n493_, new_n494_, new_n510_, new_n511_ );
nand g377 ( new_n515_, new_n513_, new_n514_ );
nand g378 ( new_n516_, new_n489_, new_n449_ );
nand g379 ( new_n517_, new_n487_, new_n447_, new_n448_, new_n484_ );
nand g380 ( new_n518_, new_n516_, new_n517_ );
nand g381 ( new_n519_, new_n518_, keyIn_0_11 );
not g382 ( new_n520_, keyIn_0_11 );
nand g383 ( new_n521_, new_n516_, new_n520_, new_n517_ );
nand g384 ( new_n522_, new_n519_, new_n521_ );
nand g385 ( new_n523_, N136, N137 );
nand g386 ( new_n524_, new_n522_, new_n523_ );
nand g387 ( new_n525_, new_n519_, N136, N137, new_n521_ );
not g388 ( new_n526_, N77 );
nand g389 ( new_n527_, new_n526_, new_n146_ );
nand g390 ( new_n528_, N77, N93 );
nand g391 ( new_n529_, new_n527_, new_n528_ );
nand g392 ( new_n530_, new_n223_, new_n207_ );
nand g393 ( new_n531_, N109, N125 );
nand g394 ( new_n532_, new_n530_, new_n531_ );
nand g395 ( new_n533_, new_n529_, new_n532_ );
nand g396 ( new_n534_, new_n527_, new_n530_, new_n528_, new_n531_ );
nand g397 ( new_n535_, new_n533_, new_n534_ );
nand g398 ( new_n536_, new_n524_, new_n525_, new_n535_ );
nand g399 ( new_n537_, new_n524_, new_n525_ );
nand g400 ( new_n538_, new_n537_, new_n533_, new_n534_ );
nand g401 ( new_n539_, new_n538_, new_n536_ );
not g402 ( new_n540_, new_n539_ );
nand g403 ( new_n541_, new_n434_, new_n469_, new_n515_, new_n540_ );
not g404 ( new_n542_, new_n541_ );
nand g405 ( new_n543_, new_n366_, new_n196_, new_n542_ );
nand g406 ( new_n544_, new_n543_, new_n139_ );
nand g407 ( new_n545_, new_n366_, keyIn_0_41, new_n196_, new_n542_ );
nand g408 ( new_n546_, new_n544_, new_n138_, new_n545_ );
nand g409 ( new_n547_, new_n544_, new_n545_ );
nand g410 ( new_n548_, new_n547_, N1 );
nand g411 ( N724, new_n548_, new_n546_ );
not g412 ( new_n550_, keyIn_0_42 );
nand g413 ( new_n551_, new_n366_, new_n350_, new_n542_ );
nand g414 ( new_n552_, new_n551_, new_n550_ );
nand g415 ( new_n553_, new_n366_, keyIn_0_42, new_n350_, new_n542_ );
nand g416 ( new_n554_, new_n552_, N5, new_n553_ );
nand g417 ( new_n555_, new_n552_, new_n553_ );
nand g418 ( new_n556_, new_n555_, new_n252_ );
nand g419 ( N725, new_n556_, new_n554_ );
nand g420 ( new_n558_, new_n366_, new_n542_ );
nor g421 ( new_n559_, new_n558_, new_n340_ );
not g422 ( new_n560_, new_n559_ );
nand g423 ( new_n561_, new_n560_, N9 );
nand g424 ( new_n562_, new_n559_, new_n320_ );
nand g425 ( N726, new_n561_, new_n562_ );
nor g426 ( new_n564_, new_n558_, new_n349_ );
not g427 ( new_n565_, new_n564_ );
nand g428 ( new_n566_, new_n565_, N13 );
nand g429 ( new_n567_, new_n564_, new_n292_ );
nand g430 ( N727, new_n566_, new_n567_ );
not g431 ( new_n569_, keyIn_0_54 );
not g432 ( new_n570_, new_n515_ );
nor g433 ( new_n571_, new_n434_, new_n468_, new_n540_, new_n570_ );
nand g434 ( new_n572_, new_n366_, new_n196_, new_n571_ );
nand g435 ( new_n573_, new_n572_, N17 );
nand g436 ( new_n574_, new_n366_, new_n181_, new_n196_, new_n571_ );
nand g437 ( new_n575_, new_n573_, new_n569_, new_n574_ );
nand g438 ( new_n576_, new_n573_, new_n574_ );
nand g439 ( new_n577_, new_n576_, keyIn_0_54 );
nand g440 ( N728, new_n577_, new_n575_ );
not g441 ( new_n579_, keyIn_0_55 );
nand g442 ( new_n580_, new_n366_, new_n350_, new_n571_ );
nand g443 ( new_n581_, new_n580_, N21 );
nand g444 ( new_n582_, new_n366_, new_n250_, new_n350_, new_n571_ );
nand g445 ( new_n583_, new_n581_, new_n579_, new_n582_ );
nand g446 ( new_n584_, new_n581_, new_n582_ );
nand g447 ( new_n585_, new_n584_, keyIn_0_55 );
nand g448 ( N729, new_n585_, new_n583_ );
not g449 ( new_n587_, new_n571_ );
nand g450 ( new_n588_, new_n366_, new_n356_ );
nor g451 ( new_n589_, new_n588_, new_n587_ );
not g452 ( new_n590_, new_n589_ );
nand g453 ( new_n591_, new_n590_, N25 );
nand g454 ( new_n592_, new_n589_, new_n321_ );
nand g455 ( N730, new_n591_, new_n592_ );
not g456 ( new_n594_, keyIn_0_43 );
nand g457 ( new_n595_, new_n366_, new_n311_, new_n571_ );
nand g458 ( new_n596_, new_n595_, new_n594_ );
nand g459 ( new_n597_, new_n366_, keyIn_0_43, new_n311_, new_n571_ );
nand g460 ( new_n598_, new_n596_, new_n290_, new_n597_ );
nand g461 ( new_n599_, new_n596_, new_n597_ );
nand g462 ( new_n600_, new_n599_, N29 );
nand g463 ( N731, new_n600_, new_n598_ );
not g464 ( new_n602_, keyIn_0_56 );
nor g465 ( new_n603_, new_n469_, new_n539_, new_n515_ );
nand g466 ( new_n604_, new_n603_, new_n434_ );
not g467 ( new_n605_, new_n604_ );
nand g468 ( new_n606_, new_n366_, new_n196_, new_n605_ );
nand g469 ( new_n607_, new_n606_, N33 );
nand g470 ( new_n608_, new_n366_, new_n185_, new_n196_, new_n605_ );
nand g471 ( new_n609_, new_n607_, new_n602_, new_n608_ );
nand g472 ( new_n610_, new_n607_, new_n608_ );
nand g473 ( new_n611_, new_n610_, keyIn_0_56 );
nand g474 ( N732, new_n611_, new_n609_ );
not g475 ( new_n613_, keyIn_0_57 );
nand g476 ( new_n614_, new_n366_, new_n350_, new_n605_ );
nand g477 ( new_n615_, new_n614_, new_n261_ );
nand g478 ( new_n616_, new_n366_, N37, new_n350_, new_n605_ );
nand g479 ( new_n617_, new_n615_, new_n613_, new_n616_ );
nand g480 ( new_n618_, new_n615_, new_n616_ );
nand g481 ( new_n619_, new_n618_, keyIn_0_57 );
nand g482 ( N733, new_n619_, new_n617_ );
not g483 ( new_n621_, keyIn_0_44 );
nand g484 ( new_n622_, new_n366_, new_n356_, new_n605_ );
nand g485 ( new_n623_, new_n622_, new_n621_ );
nand g486 ( new_n624_, new_n366_, keyIn_0_44, new_n356_, new_n605_ );
nand g487 ( new_n625_, new_n623_, new_n325_, new_n624_ );
nand g488 ( new_n626_, new_n623_, new_n624_ );
nand g489 ( new_n627_, new_n626_, N41 );
nand g490 ( N734, new_n627_, new_n625_ );
not g491 ( new_n629_, keyIn_0_45 );
nand g492 ( new_n630_, new_n366_, new_n311_, new_n605_ );
nand g493 ( new_n631_, new_n630_, new_n629_ );
nand g494 ( new_n632_, new_n366_, keyIn_0_45, new_n311_, new_n605_ );
nand g495 ( new_n633_, new_n631_, new_n632_ );
nand g496 ( new_n634_, new_n633_, N45 );
nand g497 ( new_n635_, new_n631_, new_n299_, new_n632_ );
nand g498 ( new_n636_, new_n634_, new_n635_ );
nand g499 ( new_n637_, new_n636_, keyIn_0_58 );
not g500 ( new_n638_, keyIn_0_58 );
nand g501 ( new_n639_, new_n634_, new_n638_, new_n635_ );
nand g502 ( N735, new_n637_, new_n639_ );
nand g503 ( new_n641_, new_n434_, keyIn_0_27 );
not g504 ( new_n642_, keyIn_0_27 );
not g505 ( new_n643_, new_n434_ );
nand g506 ( new_n644_, new_n643_, new_n642_ );
nand g507 ( new_n645_, new_n644_, new_n641_ );
nand g508 ( new_n646_, new_n645_, new_n468_, new_n570_, new_n539_ );
not g509 ( new_n647_, new_n646_ );
nand g510 ( new_n648_, new_n366_, keyIn_0_39, new_n647_ );
not g511 ( new_n649_, keyIn_0_39 );
nand g512 ( new_n650_, new_n366_, new_n647_ );
nand g513 ( new_n651_, new_n650_, new_n649_ );
nand g514 ( new_n652_, new_n651_, new_n648_ );
nand g515 ( new_n653_, new_n652_, new_n196_ );
nand g516 ( new_n654_, new_n653_, N49 );
nand g517 ( new_n655_, new_n652_, new_n186_, new_n196_ );
nand g518 ( new_n656_, new_n654_, new_n655_ );
nand g519 ( new_n657_, new_n656_, keyIn_0_59 );
not g520 ( new_n658_, keyIn_0_59 );
nand g521 ( new_n659_, new_n654_, new_n658_, new_n655_ );
nand g522 ( N736, new_n657_, new_n659_ );
nand g523 ( new_n661_, new_n652_, new_n350_ );
nand g524 ( new_n662_, new_n661_, keyIn_0_46 );
not g525 ( new_n663_, keyIn_0_46 );
nand g526 ( new_n664_, new_n652_, new_n663_, new_n350_ );
nand g527 ( new_n665_, new_n662_, new_n664_ );
nand g528 ( new_n666_, new_n665_, N53 );
nand g529 ( new_n667_, new_n662_, new_n259_, new_n664_ );
nand g530 ( N737, new_n666_, new_n667_ );
nand g531 ( new_n669_, new_n652_, new_n356_ );
nand g532 ( new_n670_, new_n669_, N57 );
nand g533 ( new_n671_, new_n652_, new_n326_, new_n356_ );
nand g534 ( N738, new_n670_, new_n671_ );
nand g535 ( new_n673_, new_n652_, new_n311_ );
nand g536 ( new_n674_, new_n673_, N61 );
nand g537 ( new_n675_, new_n652_, new_n301_, new_n311_ );
nand g538 ( N739, new_n674_, new_n675_ );
not g539 ( new_n677_, keyIn_0_40 );
not g540 ( new_n678_, keyIn_0_37 );
not g541 ( new_n679_, keyIn_0_31 );
nand g542 ( new_n680_, new_n432_, new_n679_, new_n433_ );
nand g543 ( new_n681_, new_n434_, keyIn_0_31 );
nand g544 ( new_n682_, new_n681_, new_n678_, new_n603_, new_n680_ );
nand g545 ( new_n683_, new_n681_, new_n603_, new_n680_ );
nand g546 ( new_n684_, new_n683_, keyIn_0_37 );
not g547 ( new_n685_, keyIn_0_32 );
nand g548 ( new_n686_, new_n643_, new_n685_ );
nand g549 ( new_n687_, new_n434_, keyIn_0_32 );
nand g550 ( new_n688_, new_n538_, keyIn_0_33, new_n536_ );
not g551 ( new_n689_, keyIn_0_33 );
nand g552 ( new_n690_, new_n539_, new_n689_ );
nand g553 ( new_n691_, new_n690_, new_n469_, new_n515_, new_n688_ );
not g554 ( new_n692_, new_n691_ );
nand g555 ( new_n693_, new_n686_, new_n692_, new_n687_ );
not g556 ( new_n694_, keyIn_0_30 );
nand g557 ( new_n695_, new_n539_, new_n694_ );
nand g558 ( new_n696_, new_n538_, keyIn_0_30, new_n536_ );
nand g559 ( new_n697_, new_n695_, new_n696_ );
not g560 ( new_n698_, keyIn_0_29 );
nand g561 ( new_n699_, new_n570_, new_n698_ );
nand g562 ( new_n700_, new_n515_, keyIn_0_29 );
nand g563 ( new_n701_, new_n699_, new_n700_ );
nor g564 ( new_n702_, new_n701_, new_n468_ );
nand g565 ( new_n703_, new_n702_, new_n434_, new_n697_ );
nand g566 ( new_n704_, new_n468_, keyIn_0_28 );
not g567 ( new_n705_, keyIn_0_28 );
nand g568 ( new_n706_, new_n469_, new_n705_ );
nand g569 ( new_n707_, new_n706_, new_n704_ );
nand g570 ( new_n708_, new_n643_, new_n707_, new_n570_, new_n539_ );
nand g571 ( new_n709_, new_n708_, new_n703_ );
not g572 ( new_n710_, new_n709_ );
nand g573 ( new_n711_, new_n710_, new_n682_, new_n684_, new_n693_ );
nand g574 ( new_n712_, new_n711_, keyIn_0_38 );
not g575 ( new_n713_, keyIn_0_38 );
not g576 ( new_n714_, new_n693_ );
nor g577 ( new_n715_, new_n714_, new_n709_ );
nand g578 ( new_n716_, new_n715_, new_n713_, new_n682_, new_n684_ );
nand g579 ( new_n717_, new_n349_, new_n356_ );
nor g580 ( new_n718_, new_n717_, new_n274_ );
nand g581 ( new_n719_, new_n712_, new_n716_, new_n677_, new_n718_ );
nand g582 ( new_n720_, new_n712_, new_n716_, new_n718_ );
nand g583 ( new_n721_, new_n720_, keyIn_0_40 );
nand g584 ( new_n722_, new_n721_, new_n719_ );
nand g585 ( new_n723_, new_n722_, new_n515_ );
nand g586 ( new_n724_, new_n723_, keyIn_0_47 );
not g587 ( new_n725_, keyIn_0_47 );
nand g588 ( new_n726_, new_n722_, new_n725_, new_n515_ );
nand g589 ( new_n727_, new_n724_, new_n726_ );
nand g590 ( new_n728_, new_n727_, new_n158_ );
nand g591 ( new_n729_, new_n724_, N65, new_n726_ );
nand g592 ( N740, new_n728_, new_n729_ );
nand g593 ( new_n731_, new_n722_, new_n468_ );
nand g594 ( new_n732_, new_n731_, keyIn_0_48 );
not g595 ( new_n733_, keyIn_0_48 );
nand g596 ( new_n734_, new_n722_, new_n733_, new_n468_ );
nand g597 ( new_n735_, new_n732_, new_n734_ );
nand g598 ( new_n736_, new_n735_, new_n159_ );
nand g599 ( new_n737_, new_n732_, N69, new_n734_ );
nand g600 ( N741, new_n736_, new_n737_ );
nand g601 ( new_n739_, new_n722_, new_n434_ );
nand g602 ( new_n740_, new_n739_, N73 );
nand g603 ( new_n741_, new_n722_, new_n420_, new_n434_ );
nand g604 ( N742, new_n740_, new_n741_ );
nand g605 ( new_n743_, new_n722_, new_n539_ );
nand g606 ( new_n744_, new_n743_, N77 );
nand g607 ( new_n745_, new_n722_, new_n526_, new_n539_ );
nand g608 ( new_n746_, new_n744_, new_n745_ );
nand g609 ( new_n747_, new_n746_, keyIn_0_60 );
not g610 ( new_n748_, keyIn_0_60 );
nand g611 ( new_n749_, new_n744_, new_n748_, new_n745_ );
nand g612 ( N743, new_n747_, new_n749_ );
nand g613 ( new_n751_, new_n712_, new_n716_ );
not g614 ( new_n752_, new_n751_ );
not g615 ( new_n753_, keyIn_0_34 );
nand g616 ( new_n754_, new_n355_, new_n753_ );
nand g617 ( new_n755_, new_n350_, keyIn_0_34 );
nand g618 ( new_n756_, new_n340_, new_n196_ );
not g619 ( new_n757_, new_n756_ );
nand g620 ( new_n758_, new_n754_, new_n311_, new_n755_, new_n757_ );
not g621 ( new_n759_, new_n758_ );
nand g622 ( new_n760_, new_n752_, new_n759_ );
not g623 ( new_n761_, new_n760_ );
nand g624 ( new_n762_, new_n761_, new_n515_ );
nand g625 ( new_n763_, new_n762_, N81 );
nand g626 ( new_n764_, new_n761_, new_n140_, new_n515_ );
nand g627 ( N744, new_n763_, new_n764_ );
nand g628 ( new_n766_, new_n752_, new_n468_, new_n759_ );
nand g629 ( new_n767_, new_n766_, keyIn_0_49 );
not g630 ( new_n768_, keyIn_0_49 );
nand g631 ( new_n769_, new_n752_, new_n468_ );
not g632 ( new_n770_, new_n769_ );
nand g633 ( new_n771_, new_n770_, new_n768_, new_n759_ );
nand g634 ( new_n772_, new_n771_, new_n141_, new_n767_ );
nand g635 ( new_n773_, new_n771_, new_n767_ );
nand g636 ( new_n774_, new_n773_, N85 );
nand g637 ( N745, new_n774_, new_n772_ );
not g638 ( new_n776_, keyIn_0_61 );
nand g639 ( new_n777_, new_n752_, new_n434_, new_n759_ );
nand g640 ( new_n778_, new_n777_, N89 );
nand g641 ( new_n779_, new_n752_, new_n145_, new_n434_, new_n759_ );
nand g642 ( new_n780_, new_n778_, new_n776_, new_n779_ );
nand g643 ( new_n781_, new_n778_, new_n779_ );
nand g644 ( new_n782_, new_n781_, keyIn_0_61 );
nand g645 ( N746, new_n782_, new_n780_ );
nand g646 ( new_n784_, new_n761_, new_n539_ );
nand g647 ( new_n785_, new_n784_, N93 );
nand g648 ( new_n786_, new_n761_, new_n146_, new_n539_ );
nand g649 ( N747, new_n785_, new_n786_ );
nand g650 ( new_n788_, new_n351_, keyIn_0_35 );
not g651 ( new_n789_, keyIn_0_35 );
nand g652 ( new_n790_, new_n196_, new_n789_ );
nand g653 ( new_n791_, new_n350_, new_n788_, new_n790_ );
nor g654 ( new_n792_, new_n717_, new_n791_ );
nand g655 ( new_n793_, new_n752_, new_n792_ );
not g656 ( new_n794_, new_n793_ );
nand g657 ( new_n795_, new_n794_, new_n515_ );
nand g658 ( new_n796_, new_n795_, N97 );
nand g659 ( new_n797_, new_n794_, new_n219_, new_n515_ );
nand g660 ( N748, new_n796_, new_n797_ );
nand g661 ( new_n799_, new_n752_, new_n468_, new_n792_ );
nand g662 ( new_n800_, new_n799_, keyIn_0_50 );
not g663 ( new_n801_, keyIn_0_50 );
nand g664 ( new_n802_, new_n770_, new_n801_, new_n792_ );
nand g665 ( new_n803_, new_n802_, new_n217_, new_n800_ );
nand g666 ( new_n804_, new_n802_, new_n800_ );
nand g667 ( new_n805_, new_n804_, N101 );
nand g668 ( N749, new_n805_, new_n803_ );
nand g669 ( new_n807_, new_n794_, new_n434_ );
nand g670 ( new_n808_, new_n807_, N105 );
nand g671 ( new_n809_, new_n794_, new_n222_, new_n434_ );
nand g672 ( N750, new_n808_, new_n809_ );
nand g673 ( new_n811_, new_n794_, new_n539_ );
nand g674 ( new_n812_, new_n811_, N109 );
nand g675 ( new_n813_, new_n794_, new_n223_, new_n539_ );
nand g676 ( N751, new_n812_, new_n813_ );
nand g677 ( new_n815_, new_n350_, new_n311_, new_n353_ );
not g678 ( new_n816_, new_n815_ );
nand g679 ( new_n817_, new_n752_, new_n816_ );
not g680 ( new_n818_, new_n817_ );
nand g681 ( new_n819_, new_n818_, new_n515_ );
nand g682 ( new_n820_, new_n819_, N113 );
nand g683 ( new_n821_, new_n818_, new_n199_, new_n515_ );
nand g684 ( N752, new_n820_, new_n821_ );
nand g685 ( new_n823_, new_n752_, new_n468_, new_n816_ );
nand g686 ( new_n824_, new_n823_, keyIn_0_51 );
not g687 ( new_n825_, keyIn_0_51 );
nand g688 ( new_n826_, new_n770_, new_n825_, new_n816_ );
nand g689 ( new_n827_, new_n826_, N117, new_n824_ );
nand g690 ( new_n828_, new_n826_, new_n824_ );
nand g691 ( new_n829_, new_n828_, new_n197_ );
nand g692 ( N753, new_n829_, new_n827_ );
not g693 ( new_n831_, keyIn_0_62 );
nand g694 ( new_n832_, new_n712_, new_n716_, new_n434_, new_n816_ );
nand g695 ( new_n833_, new_n832_, keyIn_0_52 );
not g696 ( new_n834_, keyIn_0_52 );
nand g697 ( new_n835_, new_n752_, new_n834_, new_n434_, new_n816_ );
nand g698 ( new_n836_, new_n835_, new_n833_ );
nand g699 ( new_n837_, new_n836_, new_n206_ );
nand g700 ( new_n838_, new_n835_, N121, new_n833_ );
nand g701 ( new_n839_, new_n837_, new_n838_ );
nand g702 ( new_n840_, new_n839_, new_n831_ );
nand g703 ( new_n841_, new_n837_, keyIn_0_62, new_n838_ );
nand g704 ( N754, new_n840_, new_n841_ );
not g705 ( new_n843_, keyIn_0_63 );
nand g706 ( new_n844_, new_n712_, new_n716_, new_n539_, new_n816_ );
nand g707 ( new_n845_, new_n844_, keyIn_0_53 );
not g708 ( new_n846_, keyIn_0_53 );
nand g709 ( new_n847_, new_n752_, new_n846_, new_n539_, new_n816_ );
nand g710 ( new_n848_, new_n847_, new_n845_ );
nand g711 ( new_n849_, new_n848_, N125 );
nand g712 ( new_n850_, new_n847_, new_n207_, new_n845_ );
nand g713 ( new_n851_, new_n849_, new_n850_ );
nand g714 ( new_n852_, new_n851_, new_n843_ );
nand g715 ( new_n853_, new_n849_, keyIn_0_63, new_n850_ );
nand g716 ( N755, new_n852_, new_n853_ );
endmodule