module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n155_, new_n384_, new_n410_, new_n445_, new_n236_, new_n238_, new_n479_, new_n92_, new_n79_, new_n543_, new_n250_, new_n113_, new_n501_, new_n288_, new_n371_, new_n509_, new_n97_, new_n454_, new_n421_, new_n202_, new_n296_, new_n308_, new_n368_, new_n232_, new_n258_, new_n76_, new_n439_, new_n176_, new_n283_, new_n223_, new_n390_, new_n156_, new_n306_, new_n366_, new_n494_, new_n291_, new_n241_, new_n261_, new_n309_, new_n186_, new_n365_, new_n339_, new_n197_, new_n529_, new_n386_, new_n82_, new_n401_, new_n323_, new_n259_, new_n362_, new_n514_, new_n227_, new_n416_, new_n222_, new_n456_, new_n170_, new_n400_, new_n328_, new_n460_, new_n266_, new_n367_, new_n542_, new_n173_, new_n220_, new_n130_, new_n505_, new_n419_, new_n471_, new_n268_, new_n374_, new_n534_, new_n376_, new_n380_, new_n214_, new_n451_, new_n489_, new_n424_, new_n138_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n240_, new_n413_, new_n526_, new_n352_, new_n442_, new_n485_, new_n525_, new_n211_, new_n123_, new_n127_, new_n342_, new_n126_, new_n462_, new_n177_, new_n493_, new_n264_, new_n379_, new_n500_, new_n273_, new_n224_, new_n270_, new_n317_, new_n102_, new_n344_, new_n143_, new_n287_, new_n125_, new_n145_, new_n253_, new_n504_, new_n403_, new_n475_, new_n90_, new_n237_, new_n427_, new_n234_, new_n532_, new_n149_, new_n472_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n106_, new_n411_, new_n215_, new_n507_, new_n152_, new_n157_, new_n182_, new_n93_, new_n407_, new_n153_, new_n81_, new_n480_, new_n133_, new_n257_, new_n481_, new_n212_, new_n151_, new_n513_, new_n364_, new_n449_, new_n484_, new_n219_, new_n231_, new_n313_, new_n78_, new_n239_, new_n272_, new_n282_, new_n382_, new_n522_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n146_, new_n88_, new_n487_, new_n360_, new_n98_, new_n110_, new_n315_, new_n302_, new_n191_, new_n124_, new_n326_, new_n95_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n87_, new_n387_, new_n103_, new_n476_, new_n112_, new_n248_, new_n350_, new_n117_, new_n121_, new_n415_, new_n167_, new_n537_, new_n221_, new_n385_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n478_, new_n461_, new_n459_, new_n174_, new_n297_, new_n361_, new_n468_, new_n150_, new_n354_, new_n392_, new_n444_, new_n518_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n105_, new_n340_, new_n147_, new_n510_, new_n285_, new_n502_, new_n80_, new_n351_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n517_, new_n325_, new_n417_, new_n180_, new_n515_, new_n530_, new_n332_, new_n318_, new_n453_, new_n163_, new_n519_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n531_, new_n111_, new_n158_, new_n252_, new_n486_, new_n491_, new_n466_, new_n262_, new_n160_, new_n312_, new_n271_, new_n535_, new_n274_, new_n372_, new_n100_, new_n242_, new_n503_, new_n218_, new_n497_, new_n115_, new_n307_, new_n190_, new_n305_, new_n420_, new_n408_, new_n470_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n213_, new_n134_, new_n433_, new_n435_, new_n206_, new_n109_, new_n254_, new_n429_, new_n355_, new_n353_, new_n85_, new_n432_, new_n265_, new_n506_, new_n370_, new_n256_, new_n452_, new_n278_, new_n304_, new_n381_, new_n523_, new_n388_, new_n217_, new_n101_, new_n269_, new_n508_, new_n512_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n129_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n412_, new_n165_, new_n441_, new_n477_, new_n327_, new_n216_, new_n495_, new_n431_, new_n77_, new_n196_, new_n280_, new_n426_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n338_, new_n207_, new_n267_, new_n473_, new_n140_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n86_, new_n465_, new_n84_, new_n195_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n245_, new_n402_, new_n474_, new_n89_, new_n467_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n490_, new_n91_, new_n346_, new_n396_, new_n198_, new_n438_, new_n128_, new_n358_, new_n208_, new_n348_, new_n159_, new_n83_, new_n322_, new_n228_, new_n289_, new_n528_, new_n179_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n104_, new_n185_, new_n399_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n99_, new_n329_, new_n249_, new_n233_, new_n136_, new_n469_, new_n284_, new_n119_, new_n391_, new_n293_, new_n96_, new_n178_, new_n437_, new_n168_, new_n279_, new_n455_, new_n295_, new_n359_, new_n132_, new_n120_, new_n521_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n406_, new_n356_, new_n333_, new_n229_, new_n536_, new_n290_, new_n464_, new_n94_, new_n204_, new_n369_, new_n181_, new_n135_, new_n448_, new_n276_, new_n405_;

not g000 ( new_n76_, N102 );
and g001 ( new_n77_, new_n76_, N108 );
or g002 ( new_n78_, new_n77_, keyIn_0_4 );
and g003 ( new_n79_, new_n76_, keyIn_0_4 );
and g004 ( new_n80_, new_n79_, N108 );
not g005 ( new_n81_, new_n80_ );
and g006 ( new_n82_, new_n81_, new_n78_ );
not g007 ( new_n83_, N56 );
or g008 ( new_n84_, new_n83_, N50 );
not g009 ( new_n85_, N69 );
or g010 ( new_n86_, new_n85_, N63 );
and g011 ( new_n87_, new_n84_, new_n86_ );
not g012 ( new_n88_, N82 );
or g013 ( new_n89_, new_n88_, N76 );
not g014 ( new_n90_, N95 );
or g015 ( new_n91_, new_n90_, N89 );
and g016 ( new_n92_, new_n89_, new_n91_ );
and g017 ( new_n93_, new_n87_, new_n92_ );
not g018 ( new_n94_, N4 );
or g019 ( new_n95_, new_n94_, N1 );
not g020 ( new_n96_, N17 );
or g021 ( new_n97_, new_n96_, N11 );
and g022 ( new_n98_, new_n95_, new_n97_ );
not g023 ( new_n99_, N30 );
or g024 ( new_n100_, new_n99_, N24 );
not g025 ( new_n101_, N43 );
or g026 ( new_n102_, new_n101_, N37 );
and g027 ( new_n103_, new_n100_, new_n102_ );
and g028 ( new_n104_, new_n98_, new_n103_ );
and g029 ( new_n105_, new_n93_, new_n104_ );
and g030 ( new_n106_, new_n105_, new_n82_ );
not g031 ( N223, new_n106_ );
not g032 ( new_n108_, keyIn_0_18 );
not g033 ( new_n109_, new_n82_ );
or g034 ( new_n110_, new_n105_, new_n109_ );
and g035 ( new_n111_, new_n110_, keyIn_0_14 );
not g036 ( new_n112_, new_n111_ );
or g037 ( new_n113_, new_n110_, keyIn_0_14 );
and g038 ( new_n114_, new_n112_, new_n113_ );
not g039 ( new_n115_, N112 );
not g040 ( new_n116_, N108 );
and g041 ( new_n117_, new_n116_, keyIn_0_3 );
not g042 ( new_n118_, new_n117_ );
or g043 ( new_n119_, new_n116_, keyIn_0_3 );
and g044 ( new_n120_, new_n118_, new_n119_ );
and g045 ( new_n121_, new_n120_, new_n115_ );
and g046 ( new_n122_, new_n114_, new_n121_ );
and g047 ( new_n123_, new_n122_, new_n108_ );
not g048 ( new_n124_, new_n123_ );
and g049 ( new_n125_, new_n106_, new_n84_ );
not g050 ( new_n126_, new_n125_ );
or g051 ( new_n127_, new_n106_, new_n84_ );
and g052 ( new_n128_, new_n126_, new_n127_ );
or g053 ( new_n129_, new_n128_, new_n83_ );
or g054 ( new_n130_, new_n129_, N60 );
not g055 ( new_n131_, keyIn_0_17 );
and g056 ( new_n132_, N223, new_n91_ );
not g057 ( new_n133_, new_n132_ );
not g058 ( new_n134_, N99 );
and g059 ( new_n135_, keyIn_0_2, N95 );
not g060 ( new_n136_, new_n135_ );
or g061 ( new_n137_, keyIn_0_2, N95 );
and g062 ( new_n138_, new_n136_, new_n137_ );
and g063 ( new_n139_, new_n138_, new_n134_ );
and g064 ( new_n140_, new_n133_, new_n139_ );
or g065 ( new_n141_, new_n140_, new_n131_ );
and g066 ( new_n142_, new_n140_, new_n131_ );
not g067 ( new_n143_, new_n142_ );
and g068 ( new_n144_, new_n143_, new_n141_ );
and g069 ( new_n145_, new_n144_, new_n130_ );
and g070 ( new_n146_, new_n145_, new_n124_ );
not g071 ( new_n147_, keyIn_0_10 );
or g072 ( new_n148_, new_n106_, new_n97_ );
and g073 ( new_n149_, new_n106_, new_n97_ );
not g074 ( new_n150_, new_n149_ );
and g075 ( new_n151_, new_n150_, new_n148_ );
or g076 ( new_n152_, new_n151_, new_n147_ );
not g077 ( new_n153_, N11 );
and g078 ( new_n154_, new_n153_, N17 );
and g079 ( new_n155_, N223, new_n154_ );
or g080 ( new_n156_, new_n155_, new_n149_ );
or g081 ( new_n157_, new_n156_, keyIn_0_10 );
and g082 ( new_n158_, new_n157_, new_n152_ );
not g083 ( new_n159_, N21 );
and g084 ( new_n160_, keyIn_0_1, N17 );
not g085 ( new_n161_, new_n160_ );
or g086 ( new_n162_, keyIn_0_1, N17 );
and g087 ( new_n163_, new_n161_, new_n162_ );
not g088 ( new_n164_, new_n163_ );
and g089 ( new_n165_, new_n164_, new_n159_ );
not g090 ( new_n166_, new_n165_ );
or g091 ( new_n167_, new_n158_, new_n166_ );
or g092 ( new_n168_, new_n122_, new_n108_ );
not g093 ( new_n169_, N86 );
not g094 ( new_n170_, N76 );
and g095 ( new_n171_, new_n170_, N82 );
or g096 ( new_n172_, new_n106_, new_n171_ );
and g097 ( new_n173_, new_n172_, N82 );
and g098 ( new_n174_, new_n173_, new_n169_ );
not g099 ( new_n175_, new_n174_ );
and g100 ( new_n176_, new_n106_, new_n95_ );
not g101 ( new_n177_, new_n176_ );
or g102 ( new_n178_, new_n106_, new_n95_ );
and g103 ( new_n179_, new_n177_, new_n178_ );
and g104 ( new_n180_, keyIn_0_0, N4 );
not g105 ( new_n181_, new_n180_ );
or g106 ( new_n182_, keyIn_0_0, N4 );
and g107 ( new_n183_, new_n181_, new_n182_ );
not g108 ( new_n184_, new_n183_ );
or g109 ( new_n185_, new_n184_, N8 );
or g110 ( new_n186_, new_n179_, new_n185_ );
and g111 ( new_n187_, new_n175_, new_n186_ );
and g112 ( new_n188_, new_n168_, new_n187_ );
and g113 ( new_n189_, new_n167_, new_n188_ );
not g114 ( new_n190_, keyIn_0_12 );
and g115 ( new_n191_, new_n106_, new_n102_ );
not g116 ( new_n192_, N37 );
and g117 ( new_n193_, new_n192_, N43 );
and g118 ( new_n194_, N223, new_n193_ );
or g119 ( new_n195_, new_n194_, new_n191_ );
and g120 ( new_n196_, new_n195_, new_n190_ );
not g121 ( new_n197_, new_n191_ );
or g122 ( new_n198_, new_n106_, new_n102_ );
and g123 ( new_n199_, new_n197_, new_n198_ );
and g124 ( new_n200_, new_n199_, keyIn_0_12 );
or g125 ( new_n201_, new_n196_, new_n200_ );
not g126 ( new_n202_, N47 );
and g127 ( new_n203_, new_n202_, N43 );
not g128 ( new_n204_, new_n203_ );
and g129 ( new_n205_, new_n204_, keyIn_0_6 );
not g130 ( new_n206_, new_n205_ );
or g131 ( new_n207_, new_n204_, keyIn_0_6 );
and g132 ( new_n208_, new_n206_, new_n207_ );
not g133 ( new_n209_, new_n208_ );
or g134 ( new_n210_, new_n201_, new_n209_ );
not g135 ( new_n211_, N63 );
and g136 ( new_n212_, new_n211_, N69 );
and g137 ( new_n213_, N223, new_n212_ );
and g138 ( new_n214_, new_n106_, new_n86_ );
or g139 ( new_n215_, new_n213_, new_n214_ );
and g140 ( new_n216_, new_n215_, keyIn_0_13 );
or g141 ( new_n217_, new_n216_, new_n85_ );
not g142 ( new_n218_, keyIn_0_13 );
or g143 ( new_n219_, new_n106_, new_n86_ );
not g144 ( new_n220_, new_n214_ );
and g145 ( new_n221_, new_n220_, new_n219_ );
and g146 ( new_n222_, new_n221_, new_n218_ );
or g147 ( new_n223_, new_n222_, N73 );
or g148 ( new_n224_, new_n217_, new_n223_ );
and g149 ( new_n225_, new_n210_, new_n224_ );
and g150 ( new_n226_, new_n225_, new_n189_ );
and g151 ( new_n227_, new_n226_, new_n146_ );
not g152 ( new_n228_, keyIn_0_16 );
not g153 ( new_n229_, keyIn_0_11 );
and g154 ( new_n230_, new_n106_, new_n100_ );
not g155 ( new_n231_, new_n230_ );
or g156 ( new_n232_, new_n106_, new_n100_ );
and g157 ( new_n233_, new_n231_, new_n232_ );
not g158 ( new_n234_, new_n233_ );
and g159 ( new_n235_, new_n234_, new_n229_ );
and g160 ( new_n236_, new_n233_, keyIn_0_11 );
or g161 ( new_n237_, new_n235_, new_n236_ );
not g162 ( new_n238_, N34 );
and g163 ( new_n239_, new_n238_, N30 );
and g164 ( new_n240_, new_n237_, new_n239_ );
or g165 ( new_n241_, new_n240_, new_n228_ );
and g166 ( new_n242_, new_n240_, new_n228_ );
not g167 ( new_n243_, new_n242_ );
and g168 ( new_n244_, new_n243_, new_n241_ );
and g169 ( new_n245_, new_n227_, new_n244_ );
not g170 ( N329, new_n245_ );
not g171 ( new_n247_, new_n178_ );
or g172 ( new_n248_, new_n247_, new_n176_ );
not g173 ( new_n249_, new_n185_ );
and g174 ( new_n250_, new_n248_, new_n249_ );
and g175 ( new_n251_, N329, new_n250_ );
and g176 ( new_n252_, new_n245_, new_n186_ );
or g177 ( new_n253_, new_n251_, new_n252_ );
not g178 ( new_n254_, new_n253_ );
and g179 ( new_n255_, new_n254_, keyIn_0_22 );
not g180 ( new_n256_, keyIn_0_22 );
and g181 ( new_n257_, new_n253_, new_n256_ );
or g182 ( new_n258_, new_n184_, N14 );
or g183 ( new_n259_, new_n179_, new_n258_ );
or g184 ( new_n260_, new_n257_, new_n259_ );
or g185 ( new_n261_, new_n260_, new_n255_ );
not g186 ( new_n262_, new_n261_ );
or g187 ( new_n263_, new_n199_, keyIn_0_12 );
or g188 ( new_n264_, new_n195_, new_n190_ );
and g189 ( new_n265_, new_n264_, new_n263_ );
and g190 ( new_n266_, new_n265_, new_n208_ );
or g191 ( new_n267_, new_n245_, new_n266_ );
not g192 ( new_n268_, N53 );
and g193 ( new_n269_, new_n268_, N43 );
not g194 ( new_n270_, new_n269_ );
and g195 ( new_n271_, new_n270_, keyIn_0_7 );
not g196 ( new_n272_, new_n271_ );
or g197 ( new_n273_, new_n270_, keyIn_0_7 );
and g198 ( new_n274_, new_n272_, new_n273_ );
and g199 ( new_n275_, new_n265_, new_n274_ );
and g200 ( new_n276_, new_n267_, new_n275_ );
not g201 ( new_n277_, new_n130_ );
or g202 ( new_n278_, new_n245_, new_n277_ );
not g203 ( new_n279_, N66 );
not g204 ( new_n280_, new_n129_ );
and g205 ( new_n281_, new_n280_, new_n279_ );
not g206 ( new_n282_, new_n281_ );
and g207 ( new_n283_, new_n282_, keyIn_0_21 );
not g208 ( new_n284_, new_n283_ );
or g209 ( new_n285_, new_n282_, keyIn_0_21 );
and g210 ( new_n286_, new_n284_, new_n285_ );
and g211 ( new_n287_, new_n278_, new_n286_ );
or g212 ( new_n288_, new_n276_, new_n287_ );
and g213 ( new_n289_, new_n124_, new_n168_ );
not g214 ( new_n290_, new_n289_ );
or g215 ( new_n291_, new_n245_, new_n290_ );
not g216 ( new_n292_, N115 );
and g217 ( new_n293_, new_n120_, new_n292_ );
and g218 ( new_n294_, new_n114_, new_n293_ );
and g219 ( new_n295_, new_n294_, keyIn_0_19 );
not g220 ( new_n296_, new_n295_ );
or g221 ( new_n297_, new_n294_, keyIn_0_19 );
and g222 ( new_n298_, new_n296_, new_n297_ );
not g223 ( new_n299_, new_n298_ );
and g224 ( new_n300_, new_n291_, new_n299_ );
or g225 ( new_n301_, new_n245_, new_n169_ );
not g226 ( new_n302_, N92 );
and g227 ( new_n303_, new_n173_, new_n302_ );
and g228 ( new_n304_, new_n301_, new_n303_ );
or g229 ( new_n305_, new_n300_, new_n304_ );
or g230 ( new_n306_, new_n288_, new_n305_ );
not g231 ( new_n307_, keyIn_0_23 );
not g232 ( new_n308_, new_n146_ );
and g233 ( new_n309_, new_n156_, keyIn_0_10 );
and g234 ( new_n310_, new_n151_, new_n147_ );
or g235 ( new_n311_, new_n309_, new_n310_ );
and g236 ( new_n312_, new_n311_, new_n165_ );
not g237 ( new_n313_, keyIn_0_14 );
not g238 ( new_n314_, new_n105_ );
and g239 ( new_n315_, new_n314_, new_n82_ );
and g240 ( new_n316_, new_n315_, new_n313_ );
or g241 ( new_n317_, new_n316_, new_n111_ );
not g242 ( new_n318_, new_n121_ );
or g243 ( new_n319_, new_n317_, new_n318_ );
and g244 ( new_n320_, new_n319_, keyIn_0_18 );
or g245 ( new_n321_, new_n250_, new_n174_ );
or g246 ( new_n322_, new_n321_, new_n320_ );
or g247 ( new_n323_, new_n322_, new_n312_ );
or g248 ( new_n324_, new_n221_, new_n218_ );
and g249 ( new_n325_, new_n324_, N69 );
not g250 ( new_n326_, N73 );
or g251 ( new_n327_, new_n215_, keyIn_0_13 );
and g252 ( new_n328_, new_n327_, new_n326_ );
and g253 ( new_n329_, new_n328_, new_n325_ );
or g254 ( new_n330_, new_n266_, new_n329_ );
or g255 ( new_n331_, new_n323_, new_n330_ );
or g256 ( new_n332_, new_n331_, new_n308_ );
and g257 ( new_n333_, new_n332_, new_n244_ );
and g258 ( new_n334_, new_n333_, new_n307_ );
not g259 ( new_n335_, new_n334_ );
not g260 ( new_n336_, N40 );
and g261 ( new_n337_, new_n336_, N30 );
and g262 ( new_n338_, new_n337_, keyIn_0_5 );
not g263 ( new_n339_, new_n338_ );
or g264 ( new_n340_, new_n337_, keyIn_0_5 );
and g265 ( new_n341_, new_n339_, new_n340_ );
and g266 ( new_n342_, new_n237_, new_n341_ );
not g267 ( new_n343_, new_n342_ );
and g268 ( new_n344_, new_n343_, keyIn_0_20 );
not g269 ( new_n345_, new_n344_ );
or g270 ( new_n346_, new_n343_, keyIn_0_20 );
and g271 ( new_n347_, new_n345_, new_n346_ );
not g272 ( new_n348_, new_n347_ );
or g273 ( new_n349_, new_n333_, new_n307_ );
and g274 ( new_n350_, new_n349_, new_n348_ );
and g275 ( new_n351_, new_n350_, new_n335_ );
not g276 ( new_n352_, new_n141_ );
or g277 ( new_n353_, new_n352_, new_n142_ );
or g278 ( new_n354_, new_n245_, new_n353_ );
not g279 ( new_n355_, keyIn_0_8 );
not g280 ( new_n356_, N105 );
and g281 ( new_n357_, new_n138_, new_n356_ );
not g282 ( new_n358_, new_n357_ );
and g283 ( new_n359_, new_n358_, new_n355_ );
and g284 ( new_n360_, new_n357_, keyIn_0_8 );
or g285 ( new_n361_, new_n359_, new_n360_ );
and g286 ( new_n362_, new_n133_, new_n361_ );
and g287 ( new_n363_, new_n354_, new_n362_ );
or g288 ( new_n364_, new_n245_, new_n329_ );
not g289 ( new_n365_, N79 );
and g290 ( new_n366_, new_n327_, new_n365_ );
and g291 ( new_n367_, new_n366_, new_n325_ );
and g292 ( new_n368_, new_n364_, new_n367_ );
or g293 ( new_n369_, new_n363_, new_n368_ );
or g294 ( new_n370_, new_n351_, new_n369_ );
or g295 ( new_n371_, new_n370_, new_n306_ );
not g296 ( new_n372_, keyIn_0_26 );
or g297 ( new_n373_, new_n245_, new_n167_ );
and g298 ( new_n374_, new_n245_, new_n167_ );
not g299 ( new_n375_, new_n374_ );
and g300 ( new_n376_, new_n375_, new_n373_ );
not g301 ( new_n377_, N27 );
and g302 ( new_n378_, new_n164_, new_n377_ );
and g303 ( new_n379_, new_n311_, new_n378_ );
not g304 ( new_n380_, new_n379_ );
or g305 ( new_n381_, new_n376_, new_n380_ );
and g306 ( new_n382_, new_n381_, new_n372_ );
and g307 ( new_n383_, N329, new_n312_ );
or g308 ( new_n384_, new_n383_, new_n374_ );
and g309 ( new_n385_, new_n384_, new_n379_ );
and g310 ( new_n386_, new_n385_, keyIn_0_26 );
or g311 ( new_n387_, new_n382_, new_n386_ );
or g312 ( new_n388_, new_n387_, new_n371_ );
or g313 ( N370, new_n388_, new_n262_ );
and g314 ( new_n390_, N370, N27 );
and g315 ( new_n391_, N329, N21 );
and g316 ( new_n392_, N223, keyIn_0_9 );
not g317 ( new_n393_, keyIn_0_9 );
and g318 ( new_n394_, new_n106_, new_n393_ );
or g319 ( new_n395_, new_n392_, new_n394_ );
not g320 ( new_n396_, new_n395_ );
and g321 ( new_n397_, new_n396_, N11 );
or g322 ( new_n398_, new_n397_, new_n96_ );
or g323 ( new_n399_, new_n391_, new_n398_ );
or g324 ( new_n400_, new_n390_, new_n399_ );
and g325 ( new_n401_, N370, N40 );
and g326 ( new_n402_, N329, N34 );
and g327 ( new_n403_, new_n396_, N24 );
or g328 ( new_n404_, new_n403_, new_n99_ );
or g329 ( new_n405_, new_n402_, new_n404_ );
or g330 ( new_n406_, new_n401_, new_n405_ );
and g331 ( new_n407_, new_n406_, keyIn_0_28 );
not g332 ( new_n408_, new_n407_ );
or g333 ( new_n409_, new_n406_, keyIn_0_28 );
and g334 ( new_n410_, new_n408_, new_n409_ );
not g335 ( new_n411_, new_n288_ );
not g336 ( new_n412_, new_n300_ );
not g337 ( new_n413_, new_n304_ );
and g338 ( new_n414_, new_n412_, new_n413_ );
and g339 ( new_n415_, new_n411_, new_n414_ );
not g340 ( new_n416_, new_n244_ );
or g341 ( new_n417_, new_n416_, new_n227_ );
and g342 ( new_n418_, new_n417_, keyIn_0_23 );
or g343 ( new_n419_, new_n418_, new_n347_ );
or g344 ( new_n420_, new_n419_, new_n334_ );
not g345 ( new_n421_, new_n363_ );
not g346 ( new_n422_, new_n368_ );
and g347 ( new_n423_, new_n421_, new_n422_ );
and g348 ( new_n424_, new_n423_, new_n420_ );
and g349 ( new_n425_, new_n415_, new_n424_ );
or g350 ( new_n426_, new_n385_, keyIn_0_26 );
or g351 ( new_n427_, new_n381_, new_n372_ );
and g352 ( new_n428_, new_n426_, new_n427_ );
and g353 ( new_n429_, new_n425_, new_n428_ );
and g354 ( new_n430_, new_n429_, new_n261_ );
or g355 ( new_n431_, new_n430_, new_n279_ );
and g356 ( new_n432_, N329, N60 );
and g357 ( new_n433_, new_n396_, N50 );
or g358 ( new_n434_, new_n433_, new_n83_ );
or g359 ( new_n435_, new_n432_, new_n434_ );
not g360 ( new_n436_, new_n435_ );
and g361 ( new_n437_, new_n431_, new_n436_ );
or g362 ( new_n438_, new_n430_, new_n268_ );
and g363 ( new_n439_, N329, N47 );
and g364 ( new_n440_, new_n396_, N37 );
or g365 ( new_n441_, new_n440_, new_n101_ );
or g366 ( new_n442_, new_n439_, new_n441_ );
not g367 ( new_n443_, new_n442_ );
and g368 ( new_n444_, new_n438_, new_n443_ );
or g369 ( new_n445_, new_n437_, new_n444_ );
not g370 ( new_n446_, new_n445_ );
and g371 ( new_n447_, new_n410_, new_n446_ );
and g372 ( new_n448_, new_n447_, new_n400_ );
not g373 ( new_n449_, new_n448_ );
not g374 ( new_n450_, keyIn_0_27 );
or g375 ( new_n451_, new_n430_, new_n365_ );
and g376 ( new_n452_, new_n451_, new_n450_ );
and g377 ( new_n453_, N370, N79 );
and g378 ( new_n454_, new_n453_, keyIn_0_27 );
or g379 ( new_n455_, new_n454_, new_n452_ );
and g380 ( new_n456_, N329, N73 );
not g381 ( new_n457_, new_n456_ );
and g382 ( new_n458_, new_n457_, keyIn_0_24 );
not g383 ( new_n459_, new_n458_ );
or g384 ( new_n460_, new_n457_, keyIn_0_24 );
and g385 ( new_n461_, new_n396_, N63 );
or g386 ( new_n462_, new_n461_, new_n85_ );
not g387 ( new_n463_, new_n462_ );
and g388 ( new_n464_, new_n460_, new_n463_ );
and g389 ( new_n465_, new_n464_, new_n459_ );
and g390 ( new_n466_, new_n455_, new_n465_ );
or g391 ( new_n467_, new_n466_, keyIn_0_29 );
not g392 ( new_n468_, keyIn_0_29 );
or g393 ( new_n469_, new_n453_, keyIn_0_27 );
or g394 ( new_n470_, new_n451_, new_n450_ );
and g395 ( new_n471_, new_n469_, new_n470_ );
not g396 ( new_n472_, new_n465_ );
or g397 ( new_n473_, new_n471_, new_n472_ );
or g398 ( new_n474_, new_n473_, new_n468_ );
and g399 ( new_n475_, new_n474_, new_n467_ );
and g400 ( new_n476_, N370, N92 );
not g401 ( new_n477_, new_n476_ );
and g402 ( new_n478_, new_n396_, N76 );
not g403 ( new_n479_, new_n478_ );
and g404 ( new_n480_, new_n479_, keyIn_0_15 );
not g405 ( new_n481_, new_n480_ );
or g406 ( new_n482_, new_n479_, keyIn_0_15 );
and g407 ( new_n483_, new_n482_, N82 );
and g408 ( new_n484_, new_n483_, new_n481_ );
and g409 ( new_n485_, new_n301_, new_n484_ );
and g410 ( new_n486_, new_n477_, new_n485_ );
or g411 ( new_n487_, new_n430_, new_n292_ );
or g412 ( new_n488_, new_n245_, new_n115_ );
or g413 ( new_n489_, new_n395_, new_n76_ );
and g414 ( new_n490_, new_n489_, N108 );
and g415 ( new_n491_, new_n488_, new_n490_ );
and g416 ( new_n492_, new_n487_, new_n491_ );
and g417 ( new_n493_, N370, N105 );
not g418 ( new_n494_, new_n493_ );
not g419 ( new_n495_, keyIn_0_25 );
and g420 ( new_n496_, N329, N99 );
not g421 ( new_n497_, new_n496_ );
and g422 ( new_n498_, new_n497_, new_n495_ );
and g423 ( new_n499_, new_n496_, keyIn_0_25 );
or g424 ( new_n500_, new_n498_, new_n499_ );
and g425 ( new_n501_, new_n396_, N89 );
or g426 ( new_n502_, new_n501_, new_n90_ );
not g427 ( new_n503_, new_n502_ );
and g428 ( new_n504_, new_n500_, new_n503_ );
and g429 ( new_n505_, new_n494_, new_n504_ );
or g430 ( new_n506_, new_n505_, new_n492_ );
or g431 ( new_n507_, new_n506_, new_n486_ );
or g432 ( new_n508_, new_n475_, new_n507_ );
or g433 ( new_n509_, new_n508_, new_n449_ );
and g434 ( new_n510_, N370, N14 );
and g435 ( new_n511_, N329, N8 );
and g436 ( new_n512_, new_n396_, N1 );
or g437 ( new_n513_, new_n512_, new_n94_ );
or g438 ( new_n514_, new_n511_, new_n513_ );
or g439 ( new_n515_, new_n510_, new_n514_ );
and g440 ( N421, new_n509_, new_n515_ );
and g441 ( new_n517_, new_n449_, keyIn_0_30 );
not g442 ( new_n518_, keyIn_0_30 );
and g443 ( new_n519_, new_n448_, new_n518_ );
or g444 ( N430, new_n517_, new_n519_ );
not g445 ( new_n521_, new_n400_ );
and g446 ( new_n522_, new_n475_, new_n447_ );
or g447 ( new_n523_, new_n522_, new_n521_ );
not g448 ( new_n524_, new_n410_ );
and g449 ( new_n525_, new_n446_, new_n486_ );
or g450 ( new_n526_, new_n524_, new_n525_ );
or g451 ( N431, new_n523_, new_n526_ );
not g452 ( new_n528_, keyIn_0_31 );
not g453 ( new_n529_, new_n486_ );
and g454 ( new_n530_, new_n529_, new_n505_ );
or g455 ( new_n531_, new_n530_, new_n444_ );
and g456 ( new_n532_, new_n531_, new_n410_ );
or g457 ( new_n533_, new_n523_, new_n532_ );
and g458 ( new_n534_, new_n533_, new_n528_ );
not g459 ( new_n535_, new_n447_ );
and g460 ( new_n536_, new_n473_, new_n468_ );
and g461 ( new_n537_, new_n466_, keyIn_0_29 );
or g462 ( new_n538_, new_n536_, new_n537_ );
or g463 ( new_n539_, new_n538_, new_n535_ );
and g464 ( new_n540_, new_n539_, new_n400_ );
not g465 ( new_n541_, new_n532_ );
and g466 ( new_n542_, new_n540_, new_n541_ );
and g467 ( new_n543_, new_n542_, keyIn_0_31 );
or g468 ( N432, new_n534_, new_n543_ );
endmodule