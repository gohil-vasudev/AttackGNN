module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n368_, new_n369_, new_n371_, new_n372_, new_n374_, new_n375_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n396_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n407_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n418_, new_n419_, new_n421_, new_n423_, new_n424_, new_n426_, new_n427_, new_n429_, new_n431_, new_n433_, new_n434_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n462_, new_n463_, new_n465_, new_n466_, new_n468_, new_n469_, new_n471_, new_n472_, new_n473_, new_n475_, new_n476_, new_n477_, new_n479_, new_n481_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n507_, new_n509_, new_n510_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n523_, new_n524_, new_n525_, new_n527_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_;
  INV_X1 g000 ( .A(G1GAT), .ZN(new_n138_) );
  XNOR2_X1 g001 ( .A(G155GAT), .B(KEYINPUT3), .ZN(new_n139_) );
  XNOR2_X1 g002 ( .A(G141GAT), .B(KEYINPUT2), .ZN(new_n140_) );
  XNOR2_X1 g003 ( .A(new_n139_), .B(new_n140_), .ZN(new_n141_) );
  XOR2_X1 g004 ( .A(G57GAT), .B(KEYINPUT1), .Z(new_n142_) );
  NAND2_X1 g005 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n143_) );
  XNOR2_X1 g006 ( .A(new_n142_), .B(new_n143_), .ZN(new_n144_) );
  XNOR2_X1 g007 ( .A(new_n144_), .B(new_n141_), .ZN(new_n145_) );
  XNOR2_X1 g008 ( .A(G120GAT), .B(G127GAT), .ZN(new_n146_) );
  XNOR2_X1 g009 ( .A(G113GAT), .B(KEYINPUT0), .ZN(new_n147_) );
  XNOR2_X1 g010 ( .A(new_n146_), .B(new_n147_), .ZN(new_n148_) );
  XNOR2_X1 g011 ( .A(new_n148_), .B(G1GAT), .ZN(new_n149_) );
  XNOR2_X1 g012 ( .A(new_n145_), .B(new_n149_), .ZN(new_n150_) );
  XNOR2_X1 g013 ( .A(G29GAT), .B(G134GAT), .ZN(new_n151_) );
  XNOR2_X1 g014 ( .A(new_n150_), .B(new_n151_), .ZN(new_n152_) );
  XNOR2_X1 g015 ( .A(G85GAT), .B(G162GAT), .ZN(new_n153_) );
  XOR2_X1 g016 ( .A(new_n152_), .B(new_n153_), .Z(new_n154_) );
  XNOR2_X1 g017 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(new_n155_) );
  XNOR2_X1 g018 ( .A(G148GAT), .B(KEYINPUT6), .ZN(new_n156_) );
  XNOR2_X1 g019 ( .A(new_n155_), .B(new_n156_), .ZN(new_n157_) );
  XNOR2_X1 g020 ( .A(new_n154_), .B(new_n157_), .ZN(new_n158_) );
  INV_X1 g021 ( .A(new_n158_), .ZN(new_n159_) );
  INV_X1 g022 ( .A(G15GAT), .ZN(new_n160_) );
  XNOR2_X1 g023 ( .A(new_n148_), .B(new_n160_), .ZN(new_n161_) );
  NAND2_X1 g024 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n162_) );
  NAND2_X1 g025 ( .A1(new_n161_), .A2(new_n162_), .ZN(new_n163_) );
  OR2_X1 g026 ( .A1(new_n161_), .A2(new_n162_), .ZN(new_n164_) );
  NAND2_X1 g027 ( .A1(new_n164_), .A2(new_n163_), .ZN(new_n165_) );
  XNOR2_X1 g028 ( .A(G176GAT), .B(G183GAT), .ZN(new_n166_) );
  XNOR2_X1 g029 ( .A(G71GAT), .B(KEYINPUT20), .ZN(new_n167_) );
  XOR2_X1 g030 ( .A(new_n166_), .B(new_n167_), .Z(new_n168_) );
  INV_X1 g031 ( .A(new_n168_), .ZN(new_n169_) );
  NAND2_X1 g032 ( .A1(new_n165_), .A2(new_n169_), .ZN(new_n170_) );
  NAND3_X1 g033 ( .A1(new_n164_), .A2(new_n163_), .A3(new_n168_), .ZN(new_n171_) );
  NAND2_X1 g034 ( .A1(new_n170_), .A2(new_n171_), .ZN(new_n172_) );
  XOR2_X1 g035 ( .A(G134GAT), .B(G190GAT), .Z(new_n173_) );
  XNOR2_X1 g036 ( .A(G43GAT), .B(G99GAT), .ZN(new_n174_) );
  XNOR2_X1 g037 ( .A(new_n173_), .B(new_n174_), .ZN(new_n175_) );
  XNOR2_X1 g038 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(new_n176_) );
  XNOR2_X1 g039 ( .A(G169GAT), .B(KEYINPUT19), .ZN(new_n177_) );
  XNOR2_X1 g040 ( .A(new_n176_), .B(new_n177_), .ZN(new_n178_) );
  INV_X1 g041 ( .A(new_n178_), .ZN(new_n179_) );
  XNOR2_X1 g042 ( .A(new_n179_), .B(new_n175_), .ZN(new_n180_) );
  INV_X1 g043 ( .A(new_n180_), .ZN(new_n181_) );
  NAND2_X1 g044 ( .A1(new_n172_), .A2(new_n181_), .ZN(new_n182_) );
  NAND3_X1 g045 ( .A1(new_n170_), .A2(new_n171_), .A3(new_n180_), .ZN(new_n183_) );
  NAND2_X1 g046 ( .A1(new_n182_), .A2(new_n183_), .ZN(new_n184_) );
  INV_X1 g047 ( .A(G197GAT), .ZN(new_n185_) );
  XNOR2_X1 g048 ( .A(G211GAT), .B(G218GAT), .ZN(new_n186_) );
  XNOR2_X1 g049 ( .A(G204GAT), .B(KEYINPUT21), .ZN(new_n187_) );
  XNOR2_X1 g050 ( .A(new_n186_), .B(new_n187_), .ZN(new_n188_) );
  XNOR2_X1 g051 ( .A(new_n188_), .B(new_n185_), .ZN(new_n189_) );
  NAND2_X1 g052 ( .A1(new_n189_), .A2(new_n141_), .ZN(new_n190_) );
  INV_X1 g053 ( .A(new_n141_), .ZN(new_n191_) );
  NAND2_X1 g054 ( .A1(new_n188_), .A2(new_n185_), .ZN(new_n192_) );
  OR2_X1 g055 ( .A1(new_n188_), .A2(new_n185_), .ZN(new_n193_) );
  NAND3_X1 g056 ( .A1(new_n193_), .A2(new_n191_), .A3(new_n192_), .ZN(new_n194_) );
  NAND2_X1 g057 ( .A1(new_n190_), .A2(new_n194_), .ZN(new_n195_) );
  NAND2_X1 g058 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n196_) );
  OR2_X1 g059 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n197_) );
  NAND2_X1 g060 ( .A1(new_n197_), .A2(new_n196_), .ZN(new_n198_) );
  NAND2_X1 g061 ( .A1(new_n198_), .A2(G148GAT), .ZN(new_n199_) );
  INV_X1 g062 ( .A(G148GAT), .ZN(new_n200_) );
  NAND3_X1 g063 ( .A1(new_n197_), .A2(new_n200_), .A3(new_n196_), .ZN(new_n201_) );
  NAND2_X1 g064 ( .A1(new_n199_), .A2(new_n201_), .ZN(new_n202_) );
  XNOR2_X1 g065 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(new_n203_) );
  XNOR2_X1 g066 ( .A(G22GAT), .B(KEYINPUT22), .ZN(new_n204_) );
  XNOR2_X1 g067 ( .A(new_n203_), .B(new_n204_), .ZN(new_n205_) );
  XOR2_X1 g068 ( .A(new_n205_), .B(new_n202_), .Z(new_n206_) );
  INV_X1 g069 ( .A(new_n206_), .ZN(new_n207_) );
  NAND2_X1 g070 ( .A1(new_n195_), .A2(new_n207_), .ZN(new_n208_) );
  NAND3_X1 g071 ( .A1(new_n190_), .A2(new_n194_), .A3(new_n206_), .ZN(new_n209_) );
  NAND2_X1 g072 ( .A1(new_n208_), .A2(new_n209_), .ZN(new_n210_) );
  XNOR2_X1 g073 ( .A(G50GAT), .B(G162GAT), .ZN(new_n211_) );
  INV_X1 g074 ( .A(new_n211_), .ZN(new_n212_) );
  NAND2_X1 g075 ( .A1(new_n210_), .A2(new_n212_), .ZN(new_n213_) );
  NAND3_X1 g076 ( .A1(new_n208_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n214_) );
  NAND2_X1 g077 ( .A1(new_n213_), .A2(new_n214_), .ZN(new_n215_) );
  NAND2_X1 g078 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n216_) );
  INV_X1 g079 ( .A(new_n216_), .ZN(new_n217_) );
  NAND2_X1 g080 ( .A1(new_n215_), .A2(new_n217_), .ZN(new_n218_) );
  NAND3_X1 g081 ( .A1(new_n213_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n219_) );
  NAND4_X1 g082 ( .A1(new_n218_), .A2(new_n184_), .A3(KEYINPUT26), .A4(new_n219_), .ZN(new_n220_) );
  INV_X1 g083 ( .A(KEYINPUT26), .ZN(new_n221_) );
  NAND3_X1 g084 ( .A1(new_n218_), .A2(new_n184_), .A3(new_n219_), .ZN(new_n222_) );
  NAND2_X1 g085 ( .A1(new_n222_), .A2(new_n221_), .ZN(new_n223_) );
  NAND2_X1 g086 ( .A1(new_n223_), .A2(new_n220_), .ZN(new_n224_) );
  INV_X1 g087 ( .A(KEYINPUT27), .ZN(new_n225_) );
  XNOR2_X1 g088 ( .A(G64GAT), .B(G176GAT), .ZN(new_n226_) );
  XNOR2_X1 g089 ( .A(new_n226_), .B(G92GAT), .ZN(new_n227_) );
  NAND2_X1 g090 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n228_) );
  XNOR2_X1 g091 ( .A(new_n227_), .B(new_n228_), .ZN(new_n229_) );
  XNOR2_X1 g092 ( .A(G8GAT), .B(G183GAT), .ZN(new_n230_) );
  XNOR2_X1 g093 ( .A(new_n229_), .B(new_n230_), .ZN(new_n231_) );
  XOR2_X1 g094 ( .A(G36GAT), .B(G190GAT), .Z(new_n232_) );
  XNOR2_X1 g095 ( .A(new_n189_), .B(new_n232_), .ZN(new_n233_) );
  XNOR2_X1 g096 ( .A(new_n233_), .B(new_n231_), .ZN(new_n234_) );
  XNOR2_X1 g097 ( .A(new_n234_), .B(new_n179_), .ZN(new_n235_) );
  NAND2_X1 g098 ( .A1(new_n235_), .A2(new_n225_), .ZN(new_n236_) );
  XNOR2_X1 g099 ( .A(new_n234_), .B(new_n178_), .ZN(new_n237_) );
  NAND2_X1 g100 ( .A1(new_n237_), .A2(KEYINPUT27), .ZN(new_n238_) );
  NAND2_X1 g101 ( .A1(new_n236_), .A2(new_n238_), .ZN(new_n239_) );
  NAND2_X1 g102 ( .A1(new_n224_), .A2(new_n239_), .ZN(new_n240_) );
  INV_X1 g103 ( .A(KEYINPUT25), .ZN(new_n241_) );
  NAND2_X1 g104 ( .A1(new_n218_), .A2(new_n219_), .ZN(new_n242_) );
  INV_X1 g105 ( .A(new_n184_), .ZN(new_n243_) );
  NAND2_X1 g106 ( .A1(new_n237_), .A2(new_n243_), .ZN(new_n244_) );
  NAND3_X1 g107 ( .A1(new_n244_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n245_) );
  NAND2_X1 g108 ( .A1(new_n244_), .A2(new_n242_), .ZN(new_n246_) );
  NAND2_X1 g109 ( .A1(new_n246_), .A2(KEYINPUT25), .ZN(new_n247_) );
  NAND3_X1 g110 ( .A1(new_n240_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_) );
  NAND2_X1 g111 ( .A1(new_n248_), .A2(new_n159_), .ZN(new_n249_) );
  XNOR2_X1 g112 ( .A(new_n242_), .B(KEYINPUT28), .ZN(new_n250_) );
  NAND4_X1 g113 ( .A1(new_n158_), .A2(new_n184_), .A3(new_n239_), .A4(new_n250_), .ZN(new_n251_) );
  NAND2_X1 g114 ( .A1(new_n249_), .A2(new_n251_), .ZN(new_n252_) );
  INV_X1 g115 ( .A(new_n232_), .ZN(new_n253_) );
  NAND2_X1 g116 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n254_) );
  OR2_X1 g117 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n255_) );
  NAND2_X1 g118 ( .A1(new_n255_), .A2(new_n254_), .ZN(new_n256_) );
  NAND2_X1 g119 ( .A1(new_n256_), .A2(KEYINPUT7), .ZN(new_n257_) );
  INV_X1 g120 ( .A(KEYINPUT7), .ZN(new_n258_) );
  NAND3_X1 g121 ( .A1(new_n255_), .A2(new_n258_), .A3(new_n254_), .ZN(new_n259_) );
  NAND2_X1 g122 ( .A1(new_n257_), .A2(new_n259_), .ZN(new_n260_) );
  XNOR2_X1 g123 ( .A(G85GAT), .B(G99GAT), .ZN(new_n261_) );
  NAND2_X1 g124 ( .A1(new_n261_), .A2(G92GAT), .ZN(new_n262_) );
  INV_X1 g125 ( .A(G92GAT), .ZN(new_n263_) );
  NAND2_X1 g126 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n264_) );
  OR2_X1 g127 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n265_) );
  NAND3_X1 g128 ( .A1(new_n265_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n266_) );
  NAND2_X1 g129 ( .A1(new_n262_), .A2(new_n266_), .ZN(new_n267_) );
  NAND2_X1 g130 ( .A1(new_n260_), .A2(new_n267_), .ZN(new_n268_) );
  NAND4_X1 g131 ( .A1(new_n257_), .A2(new_n262_), .A3(new_n259_), .A4(new_n266_), .ZN(new_n269_) );
  NAND2_X1 g132 ( .A1(new_n268_), .A2(new_n269_), .ZN(new_n270_) );
  XNOR2_X1 g133 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(new_n271_) );
  NAND2_X1 g134 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n272_) );
  INV_X1 g135 ( .A(new_n272_), .ZN(new_n273_) );
  NAND2_X1 g136 ( .A1(new_n271_), .A2(new_n273_), .ZN(new_n274_) );
  NAND2_X1 g137 ( .A1(KEYINPUT11), .A2(KEYINPUT10), .ZN(new_n275_) );
  OR2_X1 g138 ( .A1(KEYINPUT11), .A2(KEYINPUT10), .ZN(new_n276_) );
  NAND3_X1 g139 ( .A1(new_n276_), .A2(new_n275_), .A3(new_n272_), .ZN(new_n277_) );
  NAND2_X1 g140 ( .A1(new_n274_), .A2(new_n277_), .ZN(new_n278_) );
  NAND2_X1 g141 ( .A1(new_n278_), .A2(KEYINPUT9), .ZN(new_n279_) );
  INV_X1 g142 ( .A(KEYINPUT9), .ZN(new_n280_) );
  NAND3_X1 g143 ( .A1(new_n274_), .A2(new_n280_), .A3(new_n277_), .ZN(new_n281_) );
  NAND2_X1 g144 ( .A1(new_n279_), .A2(new_n281_), .ZN(new_n282_) );
  NAND2_X1 g145 ( .A1(new_n270_), .A2(new_n282_), .ZN(new_n283_) );
  NAND4_X1 g146 ( .A1(new_n268_), .A2(new_n279_), .A3(new_n269_), .A4(new_n281_), .ZN(new_n284_) );
  NAND2_X1 g147 ( .A1(new_n283_), .A2(new_n284_), .ZN(new_n285_) );
  XNOR2_X1 g148 ( .A(G106GAT), .B(G218GAT), .ZN(new_n286_) );
  XOR2_X1 g149 ( .A(new_n151_), .B(new_n286_), .Z(new_n287_) );
  INV_X1 g150 ( .A(new_n287_), .ZN(new_n288_) );
  NAND2_X1 g151 ( .A1(new_n285_), .A2(new_n288_), .ZN(new_n289_) );
  NAND3_X1 g152 ( .A1(new_n283_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n290_) );
  NAND2_X1 g153 ( .A1(new_n289_), .A2(new_n290_), .ZN(new_n291_) );
  NAND2_X1 g154 ( .A1(new_n291_), .A2(new_n212_), .ZN(new_n292_) );
  NAND3_X1 g155 ( .A1(new_n289_), .A2(new_n211_), .A3(new_n290_), .ZN(new_n293_) );
  NAND2_X1 g156 ( .A1(new_n292_), .A2(new_n293_), .ZN(new_n294_) );
  NAND2_X1 g157 ( .A1(new_n294_), .A2(new_n253_), .ZN(new_n295_) );
  NAND3_X1 g158 ( .A1(new_n292_), .A2(new_n232_), .A3(new_n293_), .ZN(new_n296_) );
  NAND2_X1 g159 ( .A1(new_n295_), .A2(new_n296_), .ZN(new_n297_) );
  INV_X1 g160 ( .A(new_n297_), .ZN(new_n298_) );
  XNOR2_X1 g161 ( .A(G57GAT), .B(G71GAT), .ZN(new_n299_) );
  XOR2_X1 g162 ( .A(new_n299_), .B(KEYINPUT13), .Z(new_n300_) );
  XNOR2_X1 g163 ( .A(G15GAT), .B(G22GAT), .ZN(new_n301_) );
  XNOR2_X1 g164 ( .A(new_n301_), .B(new_n138_), .ZN(new_n302_) );
  XNOR2_X1 g165 ( .A(new_n300_), .B(new_n302_), .ZN(new_n303_) );
  XNOR2_X1 g166 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(new_n304_) );
  XNOR2_X1 g167 ( .A(G64GAT), .B(KEYINPUT15), .ZN(new_n305_) );
  XNOR2_X1 g168 ( .A(new_n304_), .B(new_n305_), .ZN(new_n306_) );
  XNOR2_X1 g169 ( .A(G78GAT), .B(G155GAT), .ZN(new_n307_) );
  XNOR2_X1 g170 ( .A(G127GAT), .B(G211GAT), .ZN(new_n308_) );
  XNOR2_X1 g171 ( .A(new_n307_), .B(new_n308_), .ZN(new_n309_) );
  XNOR2_X1 g172 ( .A(new_n306_), .B(new_n309_), .ZN(new_n310_) );
  XNOR2_X1 g173 ( .A(new_n303_), .B(new_n310_), .ZN(new_n311_) );
  XNOR2_X1 g174 ( .A(new_n311_), .B(new_n230_), .ZN(new_n312_) );
  NAND2_X1 g175 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n313_) );
  INV_X1 g176 ( .A(new_n313_), .ZN(new_n314_) );
  XNOR2_X1 g177 ( .A(new_n312_), .B(new_n314_), .ZN(new_n315_) );
  NAND2_X1 g178 ( .A1(new_n315_), .A2(new_n298_), .ZN(new_n316_) );
  XOR2_X1 g179 ( .A(new_n316_), .B(KEYINPUT16), .Z(new_n317_) );
  AND2_X1 g180 ( .A1(new_n252_), .A2(new_n317_), .ZN(new_n318_) );
  XOR2_X1 g181 ( .A(new_n302_), .B(new_n260_), .Z(new_n319_) );
  XNOR2_X1 g182 ( .A(G113GAT), .B(G197GAT), .ZN(new_n320_) );
  XNOR2_X1 g183 ( .A(G29GAT), .B(G141GAT), .ZN(new_n321_) );
  XNOR2_X1 g184 ( .A(new_n320_), .B(new_n321_), .ZN(new_n322_) );
  XNOR2_X1 g185 ( .A(G8GAT), .B(G169GAT), .ZN(new_n323_) );
  XNOR2_X1 g186 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(new_n324_) );
  XNOR2_X1 g187 ( .A(new_n323_), .B(new_n324_), .ZN(new_n325_) );
  XNOR2_X1 g188 ( .A(new_n322_), .B(new_n325_), .ZN(new_n326_) );
  XNOR2_X1 g189 ( .A(new_n319_), .B(new_n326_), .ZN(new_n327_) );
  XNOR2_X1 g190 ( .A(G36GAT), .B(G50GAT), .ZN(new_n328_) );
  NAND2_X1 g191 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n329_) );
  XNOR2_X1 g192 ( .A(new_n328_), .B(new_n329_), .ZN(new_n330_) );
  XOR2_X1 g193 ( .A(new_n327_), .B(new_n330_), .Z(new_n331_) );
  XOR2_X1 g194 ( .A(G120GAT), .B(G204GAT), .Z(new_n332_) );
  INV_X1 g195 ( .A(new_n332_), .ZN(new_n333_) );
  NAND2_X1 g196 ( .A1(new_n202_), .A2(new_n267_), .ZN(new_n334_) );
  NAND4_X1 g197 ( .A1(new_n199_), .A2(new_n262_), .A3(new_n201_), .A4(new_n266_), .ZN(new_n335_) );
  NAND2_X1 g198 ( .A1(new_n334_), .A2(new_n335_), .ZN(new_n336_) );
  XNOR2_X1 g199 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(new_n337_) );
  NAND2_X1 g200 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n338_) );
  INV_X1 g201 ( .A(new_n338_), .ZN(new_n339_) );
  NAND2_X1 g202 ( .A1(new_n337_), .A2(new_n339_), .ZN(new_n340_) );
  NAND2_X1 g203 ( .A1(KEYINPUT33), .A2(KEYINPUT31), .ZN(new_n341_) );
  OR2_X1 g204 ( .A1(KEYINPUT33), .A2(KEYINPUT31), .ZN(new_n342_) );
  NAND3_X1 g205 ( .A1(new_n342_), .A2(new_n341_), .A3(new_n338_), .ZN(new_n343_) );
  NAND2_X1 g206 ( .A1(new_n340_), .A2(new_n343_), .ZN(new_n344_) );
  NAND2_X1 g207 ( .A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n345_) );
  INV_X1 g208 ( .A(KEYINPUT32), .ZN(new_n346_) );
  NAND3_X1 g209 ( .A1(new_n340_), .A2(new_n346_), .A3(new_n343_), .ZN(new_n347_) );
  NAND2_X1 g210 ( .A1(new_n345_), .A2(new_n347_), .ZN(new_n348_) );
  NAND2_X1 g211 ( .A1(new_n336_), .A2(new_n348_), .ZN(new_n349_) );
  NAND4_X1 g212 ( .A1(new_n334_), .A2(new_n345_), .A3(new_n335_), .A4(new_n347_), .ZN(new_n350_) );
  NAND2_X1 g213 ( .A1(new_n349_), .A2(new_n350_), .ZN(new_n351_) );
  NAND2_X1 g214 ( .A1(new_n351_), .A2(new_n226_), .ZN(new_n352_) );
  INV_X1 g215 ( .A(new_n226_), .ZN(new_n353_) );
  NAND3_X1 g216 ( .A1(new_n349_), .A2(new_n353_), .A3(new_n350_), .ZN(new_n354_) );
  NAND3_X1 g217 ( .A1(new_n352_), .A2(new_n333_), .A3(new_n354_), .ZN(new_n355_) );
  NAND2_X1 g218 ( .A1(new_n352_), .A2(new_n354_), .ZN(new_n356_) );
  NAND2_X1 g219 ( .A1(new_n356_), .A2(new_n332_), .ZN(new_n357_) );
  NAND2_X1 g220 ( .A1(new_n357_), .A2(new_n355_), .ZN(new_n358_) );
  NAND2_X1 g221 ( .A1(new_n358_), .A2(new_n300_), .ZN(new_n359_) );
  INV_X1 g222 ( .A(new_n300_), .ZN(new_n360_) );
  NAND3_X1 g223 ( .A1(new_n357_), .A2(new_n360_), .A3(new_n355_), .ZN(new_n361_) );
  NAND2_X1 g224 ( .A1(new_n359_), .A2(new_n361_), .ZN(new_n362_) );
  AND2_X1 g225 ( .A1(new_n362_), .A2(new_n331_), .ZN(new_n363_) );
  NAND2_X1 g226 ( .A1(new_n318_), .A2(new_n363_), .ZN(new_n364_) );
  NOR2_X1 g227 ( .A1(new_n364_), .A2(new_n159_), .ZN(new_n365_) );
  XNOR2_X1 g228 ( .A(new_n365_), .B(KEYINPUT34), .ZN(new_n366_) );
  XNOR2_X1 g229 ( .A(new_n366_), .B(new_n138_), .ZN(G1324GAT) );
  INV_X1 g230 ( .A(new_n364_), .ZN(new_n368_) );
  NAND2_X1 g231 ( .A1(new_n368_), .A2(new_n237_), .ZN(new_n369_) );
  XNOR2_X1 g232 ( .A(new_n369_), .B(G8GAT), .ZN(G1325GAT) );
  NOR2_X1 g233 ( .A1(new_n364_), .A2(new_n184_), .ZN(new_n371_) );
  XNOR2_X1 g234 ( .A(G15GAT), .B(KEYINPUT35), .ZN(new_n372_) );
  XNOR2_X1 g235 ( .A(new_n371_), .B(new_n372_), .ZN(G1326GAT) );
  INV_X1 g236 ( .A(new_n250_), .ZN(new_n374_) );
  NAND2_X1 g237 ( .A1(new_n368_), .A2(new_n374_), .ZN(new_n375_) );
  XNOR2_X1 g238 ( .A(new_n375_), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 g239 ( .A(KEYINPUT37), .ZN(new_n377_) );
  NAND2_X1 g240 ( .A1(new_n297_), .A2(KEYINPUT36), .ZN(new_n378_) );
  INV_X1 g241 ( .A(KEYINPUT36), .ZN(new_n379_) );
  NAND3_X1 g242 ( .A1(new_n295_), .A2(new_n379_), .A3(new_n296_), .ZN(new_n380_) );
  NAND2_X1 g243 ( .A1(new_n378_), .A2(new_n380_), .ZN(new_n381_) );
  INV_X1 g244 ( .A(new_n381_), .ZN(new_n382_) );
  NOR2_X1 g245 ( .A1(new_n382_), .A2(new_n315_), .ZN(new_n383_) );
  NAND3_X1 g246 ( .A1(new_n252_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n384_) );
  NAND2_X1 g247 ( .A1(new_n252_), .A2(new_n383_), .ZN(new_n385_) );
  NAND2_X1 g248 ( .A1(new_n385_), .A2(KEYINPUT37), .ZN(new_n386_) );
  NAND2_X1 g249 ( .A1(new_n386_), .A2(new_n384_), .ZN(new_n387_) );
  NAND3_X1 g250 ( .A1(new_n387_), .A2(KEYINPUT38), .A3(new_n363_), .ZN(new_n388_) );
  INV_X1 g251 ( .A(KEYINPUT38), .ZN(new_n389_) );
  NAND2_X1 g252 ( .A1(new_n387_), .A2(new_n363_), .ZN(new_n390_) );
  NAND2_X1 g253 ( .A1(new_n390_), .A2(new_n389_), .ZN(new_n391_) );
  NAND2_X1 g254 ( .A1(new_n391_), .A2(new_n388_), .ZN(new_n392_) );
  NAND2_X1 g255 ( .A1(new_n392_), .A2(new_n158_), .ZN(new_n393_) );
  XOR2_X1 g256 ( .A(G29GAT), .B(KEYINPUT39), .Z(new_n394_) );
  XNOR2_X1 g257 ( .A(new_n393_), .B(new_n394_), .ZN(G1328GAT) );
  NAND2_X1 g258 ( .A1(new_n392_), .A2(new_n237_), .ZN(new_n396_) );
  XNOR2_X1 g259 ( .A(new_n396_), .B(G36GAT), .ZN(G1329GAT) );
  INV_X1 g260 ( .A(G43GAT), .ZN(new_n398_) );
  NAND3_X1 g261 ( .A1(new_n392_), .A2(KEYINPUT40), .A3(new_n243_), .ZN(new_n399_) );
  INV_X1 g262 ( .A(KEYINPUT40), .ZN(new_n400_) );
  NAND2_X1 g263 ( .A1(new_n392_), .A2(new_n243_), .ZN(new_n401_) );
  NAND2_X1 g264 ( .A1(new_n401_), .A2(new_n400_), .ZN(new_n402_) );
  NAND2_X1 g265 ( .A1(new_n402_), .A2(new_n399_), .ZN(new_n403_) );
  NAND2_X1 g266 ( .A1(new_n403_), .A2(new_n398_), .ZN(new_n404_) );
  NAND3_X1 g267 ( .A1(new_n402_), .A2(G43GAT), .A3(new_n399_), .ZN(new_n405_) );
  NAND2_X1 g268 ( .A1(new_n404_), .A2(new_n405_), .ZN(G1330GAT) );
  NAND2_X1 g269 ( .A1(new_n392_), .A2(new_n374_), .ZN(new_n407_) );
  XNOR2_X1 g270 ( .A(new_n407_), .B(G50GAT), .ZN(G1331GAT) );
  NAND3_X1 g271 ( .A1(new_n359_), .A2(KEYINPUT41), .A3(new_n361_), .ZN(new_n409_) );
  INV_X1 g272 ( .A(KEYINPUT41), .ZN(new_n410_) );
  NAND2_X1 g273 ( .A1(new_n362_), .A2(new_n410_), .ZN(new_n411_) );
  NAND2_X1 g274 ( .A1(new_n411_), .A2(new_n409_), .ZN(new_n412_) );
  NOR2_X1 g275 ( .A1(new_n412_), .A2(new_n331_), .ZN(new_n413_) );
  NAND2_X1 g276 ( .A1(new_n318_), .A2(new_n413_), .ZN(new_n414_) );
  NOR2_X1 g277 ( .A1(new_n414_), .A2(new_n159_), .ZN(new_n415_) );
  XOR2_X1 g278 ( .A(G57GAT), .B(KEYINPUT42), .Z(new_n416_) );
  XNOR2_X1 g279 ( .A(new_n415_), .B(new_n416_), .ZN(G1332GAT) );
  INV_X1 g280 ( .A(new_n414_), .ZN(new_n418_) );
  NAND2_X1 g281 ( .A1(new_n418_), .A2(new_n237_), .ZN(new_n419_) );
  XNOR2_X1 g282 ( .A(new_n419_), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 g283 ( .A1(new_n418_), .A2(new_n243_), .ZN(new_n421_) );
  XNOR2_X1 g284 ( .A(new_n421_), .B(G71GAT), .ZN(G1334GAT) );
  NOR2_X1 g285 ( .A1(new_n414_), .A2(new_n250_), .ZN(new_n423_) );
  XNOR2_X1 g286 ( .A(G78GAT), .B(KEYINPUT43), .ZN(new_n424_) );
  XNOR2_X1 g287 ( .A(new_n423_), .B(new_n424_), .ZN(G1335GAT) );
  AND2_X1 g288 ( .A1(new_n387_), .A2(new_n413_), .ZN(new_n426_) );
  NAND2_X1 g289 ( .A1(new_n426_), .A2(new_n158_), .ZN(new_n427_) );
  XNOR2_X1 g290 ( .A(new_n427_), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 g291 ( .A1(new_n426_), .A2(new_n237_), .ZN(new_n429_) );
  XNOR2_X1 g292 ( .A(new_n429_), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 g293 ( .A1(new_n426_), .A2(new_n243_), .ZN(new_n431_) );
  XNOR2_X1 g294 ( .A(new_n431_), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 g295 ( .A1(new_n426_), .A2(new_n374_), .ZN(new_n433_) );
  XNOR2_X1 g296 ( .A(new_n433_), .B(KEYINPUT44), .ZN(new_n434_) );
  XNOR2_X1 g297 ( .A(new_n434_), .B(G106GAT), .ZN(G1339GAT) );
  INV_X1 g298 ( .A(KEYINPUT47), .ZN(new_n436_) );
  NAND4_X1 g299 ( .A1(new_n411_), .A2(KEYINPUT46), .A3(new_n331_), .A4(new_n409_), .ZN(new_n437_) );
  INV_X1 g300 ( .A(KEYINPUT46), .ZN(new_n438_) );
  NAND3_X1 g301 ( .A1(new_n411_), .A2(new_n331_), .A3(new_n409_), .ZN(new_n439_) );
  NAND2_X1 g302 ( .A1(new_n439_), .A2(new_n438_), .ZN(new_n440_) );
  NOR2_X1 g303 ( .A1(new_n315_), .A2(new_n297_), .ZN(new_n441_) );
  NAND4_X1 g304 ( .A1(new_n440_), .A2(new_n436_), .A3(new_n437_), .A4(new_n441_), .ZN(new_n442_) );
  NAND2_X1 g305 ( .A1(new_n381_), .A2(new_n315_), .ZN(new_n443_) );
  NAND2_X1 g306 ( .A1(new_n443_), .A2(KEYINPUT45), .ZN(new_n444_) );
  INV_X1 g307 ( .A(KEYINPUT45), .ZN(new_n445_) );
  NAND3_X1 g308 ( .A1(new_n381_), .A2(new_n445_), .A3(new_n315_), .ZN(new_n446_) );
  INV_X1 g309 ( .A(new_n362_), .ZN(new_n447_) );
  NOR2_X1 g310 ( .A1(new_n447_), .A2(new_n331_), .ZN(new_n448_) );
  NAND3_X1 g311 ( .A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_) );
  NAND3_X1 g312 ( .A1(new_n440_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n450_) );
  NAND2_X1 g313 ( .A1(new_n450_), .A2(KEYINPUT47), .ZN(new_n451_) );
  NAND4_X1 g314 ( .A1(new_n451_), .A2(new_n449_), .A3(KEYINPUT48), .A4(new_n442_), .ZN(new_n452_) );
  INV_X1 g315 ( .A(KEYINPUT48), .ZN(new_n453_) );
  NAND3_X1 g316 ( .A1(new_n451_), .A2(new_n442_), .A3(new_n449_), .ZN(new_n454_) );
  NAND2_X1 g317 ( .A1(new_n454_), .A2(new_n453_), .ZN(new_n455_) );
  AND4_X1 g318 ( .A1(new_n158_), .A2(new_n455_), .A3(new_n239_), .A4(new_n452_), .ZN(new_n456_) );
  NOR2_X1 g319 ( .A1(new_n374_), .A2(new_n184_), .ZN(new_n457_) );
  NAND2_X1 g320 ( .A1(new_n456_), .A2(new_n457_), .ZN(new_n458_) );
  INV_X1 g321 ( .A(new_n458_), .ZN(new_n459_) );
  NAND2_X1 g322 ( .A1(new_n459_), .A2(new_n331_), .ZN(new_n460_) );
  XNOR2_X1 g323 ( .A(new_n460_), .B(G113GAT), .ZN(G1340GAT) );
  NOR2_X1 g324 ( .A1(new_n458_), .A2(new_n412_), .ZN(new_n462_) );
  XNOR2_X1 g325 ( .A(G120GAT), .B(KEYINPUT49), .ZN(new_n463_) );
  XNOR2_X1 g326 ( .A(new_n462_), .B(new_n463_), .ZN(G1341GAT) );
  NAND2_X1 g327 ( .A1(new_n459_), .A2(new_n315_), .ZN(new_n465_) );
  XNOR2_X1 g328 ( .A(new_n465_), .B(KEYINPUT50), .ZN(new_n466_) );
  XNOR2_X1 g329 ( .A(new_n466_), .B(G127GAT), .ZN(G1342GAT) );
  NOR2_X1 g330 ( .A1(new_n458_), .A2(new_n298_), .ZN(new_n468_) );
  XNOR2_X1 g331 ( .A(G134GAT), .B(KEYINPUT51), .ZN(new_n469_) );
  XNOR2_X1 g332 ( .A(new_n468_), .B(new_n469_), .ZN(G1343GAT) );
  NAND2_X1 g333 ( .A1(new_n456_), .A2(new_n224_), .ZN(new_n471_) );
  INV_X1 g334 ( .A(new_n471_), .ZN(new_n472_) );
  NAND2_X1 g335 ( .A1(new_n472_), .A2(new_n331_), .ZN(new_n473_) );
  XNOR2_X1 g336 ( .A(new_n473_), .B(G141GAT), .ZN(G1344GAT) );
  NOR2_X1 g337 ( .A1(new_n471_), .A2(new_n412_), .ZN(new_n475_) );
  XOR2_X1 g338 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(new_n476_) );
  XNOR2_X1 g339 ( .A(new_n475_), .B(new_n476_), .ZN(new_n477_) );
  XNOR2_X1 g340 ( .A(new_n477_), .B(new_n200_), .ZN(G1345GAT) );
  NAND2_X1 g341 ( .A1(new_n472_), .A2(new_n315_), .ZN(new_n479_) );
  XNOR2_X1 g342 ( .A(new_n479_), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 g343 ( .A1(new_n472_), .A2(new_n297_), .ZN(new_n481_) );
  XNOR2_X1 g344 ( .A(new_n481_), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 g345 ( .A(KEYINPUT55), .ZN(new_n483_) );
  NAND3_X1 g346 ( .A1(new_n455_), .A2(new_n237_), .A3(new_n452_), .ZN(new_n484_) );
  NAND2_X1 g347 ( .A1(new_n484_), .A2(KEYINPUT54), .ZN(new_n485_) );
  INV_X1 g348 ( .A(KEYINPUT54), .ZN(new_n486_) );
  NAND4_X1 g349 ( .A1(new_n455_), .A2(new_n486_), .A3(new_n237_), .A4(new_n452_), .ZN(new_n487_) );
  AND2_X1 g350 ( .A1(new_n487_), .A2(new_n242_), .ZN(new_n488_) );
  NAND4_X1 g351 ( .A1(new_n488_), .A2(new_n483_), .A3(new_n159_), .A4(new_n485_), .ZN(new_n489_) );
  NAND4_X1 g352 ( .A1(new_n485_), .A2(new_n159_), .A3(new_n242_), .A4(new_n487_), .ZN(new_n490_) );
  NAND2_X1 g353 ( .A1(new_n490_), .A2(KEYINPUT55), .ZN(new_n491_) );
  NAND2_X1 g354 ( .A1(new_n491_), .A2(new_n489_), .ZN(new_n492_) );
  AND2_X1 g355 ( .A1(new_n492_), .A2(new_n243_), .ZN(new_n493_) );
  NAND2_X1 g356 ( .A1(new_n493_), .A2(new_n331_), .ZN(new_n494_) );
  XNOR2_X1 g357 ( .A(new_n494_), .B(G169GAT), .ZN(G1348GAT) );
  INV_X1 g358 ( .A(G176GAT), .ZN(new_n496_) );
  INV_X1 g359 ( .A(new_n412_), .ZN(new_n497_) );
  XNOR2_X1 g360 ( .A(KEYINPUT57), .B(KEYINPUT56), .ZN(new_n498_) );
  INV_X1 g361 ( .A(new_n498_), .ZN(new_n499_) );
  NAND4_X1 g362 ( .A1(new_n492_), .A2(new_n243_), .A3(new_n497_), .A4(new_n499_), .ZN(new_n500_) );
  NAND3_X1 g363 ( .A1(new_n492_), .A2(new_n243_), .A3(new_n497_), .ZN(new_n501_) );
  NAND2_X1 g364 ( .A1(new_n501_), .A2(new_n498_), .ZN(new_n502_) );
  NAND2_X1 g365 ( .A1(new_n502_), .A2(new_n500_), .ZN(new_n503_) );
  NAND2_X1 g366 ( .A1(new_n503_), .A2(new_n496_), .ZN(new_n504_) );
  NAND3_X1 g367 ( .A1(new_n502_), .A2(G176GAT), .A3(new_n500_), .ZN(new_n505_) );
  NAND2_X1 g368 ( .A1(new_n504_), .A2(new_n505_), .ZN(G1349GAT) );
  NAND2_X1 g369 ( .A1(new_n493_), .A2(new_n315_), .ZN(new_n507_) );
  XNOR2_X1 g370 ( .A(new_n507_), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 g371 ( .A1(new_n493_), .A2(new_n297_), .ZN(new_n509_) );
  XNOR2_X1 g372 ( .A(G190GAT), .B(KEYINPUT58), .ZN(new_n510_) );
  XNOR2_X1 g373 ( .A(new_n509_), .B(new_n510_), .ZN(G1351GAT) );
  AND2_X1 g374 ( .A1(new_n485_), .A2(new_n159_), .ZN(new_n512_) );
  AND2_X1 g375 ( .A1(new_n487_), .A2(new_n224_), .ZN(new_n513_) );
  AND2_X1 g376 ( .A1(new_n512_), .A2(new_n513_), .ZN(new_n514_) );
  NAND2_X1 g377 ( .A1(new_n514_), .A2(new_n331_), .ZN(new_n515_) );
  XNOR2_X1 g378 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(new_n516_) );
  XNOR2_X1 g379 ( .A(new_n515_), .B(new_n516_), .ZN(new_n517_) );
  NAND2_X1 g380 ( .A1(new_n517_), .A2(new_n185_), .ZN(new_n518_) );
  OR2_X1 g381 ( .A1(new_n515_), .A2(new_n516_), .ZN(new_n519_) );
  NAND2_X1 g382 ( .A1(new_n515_), .A2(new_n516_), .ZN(new_n520_) );
  NAND3_X1 g383 ( .A1(new_n519_), .A2(G197GAT), .A3(new_n520_), .ZN(new_n521_) );
  NAND2_X1 g384 ( .A1(new_n518_), .A2(new_n521_), .ZN(G1352GAT) );
  NAND2_X1 g385 ( .A1(new_n512_), .A2(new_n513_), .ZN(new_n523_) );
  NOR2_X1 g386 ( .A1(new_n523_), .A2(new_n362_), .ZN(new_n524_) );
  XNOR2_X1 g387 ( .A(G204GAT), .B(KEYINPUT61), .ZN(new_n525_) );
  XNOR2_X1 g388 ( .A(new_n524_), .B(new_n525_), .ZN(G1353GAT) );
  NAND2_X1 g389 ( .A1(new_n514_), .A2(new_n315_), .ZN(new_n527_) );
  XNOR2_X1 g390 ( .A(new_n527_), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 g391 ( .A(G218GAT), .ZN(new_n529_) );
  NOR2_X1 g392 ( .A1(new_n523_), .A2(new_n382_), .ZN(new_n530_) );
  NAND2_X1 g393 ( .A1(new_n530_), .A2(KEYINPUT62), .ZN(new_n531_) );
  OR2_X1 g394 ( .A1(new_n530_), .A2(KEYINPUT62), .ZN(new_n532_) );
  NAND2_X1 g395 ( .A1(new_n532_), .A2(new_n531_), .ZN(new_n533_) );
  NAND2_X1 g396 ( .A1(new_n533_), .A2(new_n529_), .ZN(new_n534_) );
  NAND3_X1 g397 ( .A1(new_n532_), .A2(G218GAT), .A3(new_n531_), .ZN(new_n535_) );
  NAND2_X1 g398 ( .A1(new_n534_), .A2(new_n535_), .ZN(G1355GAT) );
endmodule


