module s38417 ( CK, g1249, g16297, g16355, g16399, g16437, g16496, g1943, 
        g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g2637, 
        g27380, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, 
        g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, 
        g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, 
        g4450, g4590, g51, g5388, g5437, g5472, g5511, g5549, g5555, g5595, 
        g5612, g5629, g563, g5637, g5648, g5657, g5686, g5695, g5738, g5747, 
        g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, 
        g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, 
        g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, 
        g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, 
        g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, 
        g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, 
        g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, test_se, 
        test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, 
        test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, 
        test_si8, test_so8, test_si9, test_so9, test_si10, test_so10, 
        test_si11, test_so11, test_si12, test_so12, test_si13, test_so13, 
        test_si14, test_so14, test_si15, test_so15, test_si16, test_so16, 
        test_si17, test_so17, test_si18, test_so18, test_si19, test_so19, 
        test_si20, test_so20, test_si21, test_so21, test_si22, test_so22, 
        test_si23, test_so23, test_si24, test_so24, test_si25, test_so25, 
        test_si26, test_so26, test_si27, test_so27, test_si28, test_so28, 
        test_si29, test_so29, test_si30, test_so30, test_si31, test_so31, 
        test_si32, test_so32, test_si33, test_so33, test_si34, test_so34, 
        test_si35, test_so35, test_si36, test_so36, test_si37, test_so37, 
        test_si38, test_so38, test_si39, test_so39, test_si40, test_so40, 
        test_si41, test_so41, test_si42, test_so42, test_si43, test_so43, 
        test_si44, test_so44, test_si45, test_so45, test_si46, test_so46, 
        test_si47, test_so47, test_si48, test_so48, test_si49, test_so49, 
        test_si50, test_so50, test_si51, test_so51, test_si52, test_so52, 
        test_si53, test_so53, test_si54, test_so54, test_si55, test_so55, 
        test_si56, test_so56, test_si57, test_so57, test_si58, test_so58, 
        test_si59, test_so59, test_si60, test_so60, test_si61, test_so61, 
        test_si62, test_so62, test_si63, test_so63, test_si64, test_so64, 
        test_si65, test_so65, test_si66, test_so66, test_si67, test_so67, 
        test_si68, test_so68, test_si69, test_so69, test_si70, test_so70, 
        test_si71, test_so71, test_si72, test_so72, test_si73, test_so73, 
        test_si74, test_so74, test_si75, test_so75, test_si76, test_so76, 
        test_si77, test_so77, test_si78, test_so78, test_si79, test_so79, 
        test_si80, test_so80, test_si81, test_so81, test_si82, test_so82, 
        test_si83, test_so83, test_si84, test_so84, test_si85, test_so85, 
        test_si86, test_so86, test_si87, test_so87, test_si88, test_so88, 
        test_si89, test_so89, test_si90, test_so90, test_si91, test_so91, 
        test_si92, test_so92, test_si93, test_so93, test_si94, test_so94, 
        test_si95, test_so95, test_si96, test_so96, test_si97, test_so97, 
        test_si98, test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217,
         g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227,
         g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;
  output g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275,
         test_so1, test_so2, test_so3, test_so4, test_so5, test_so6, test_so7,
         test_so8, test_so9, test_so10, test_so11, test_so12, test_so13,
         test_so14, test_so15, test_so16, test_so17, test_so18, test_so19,
         test_so20, test_so21, test_so22, test_so23, test_so24, test_so25,
         test_so26, test_so27, test_so28, test_so29, test_so30, test_so31,
         test_so32, test_so33, test_so34, test_so35, test_so36, test_so37,
         test_so38, test_so39, test_so40, test_so41, test_so42, test_so43,
         test_so44, test_so45, test_so46, test_so47, test_so48, test_so49,
         test_so50, test_so51, test_so52, test_so53, test_so54, test_so55,
         test_so56, test_so57, test_so58, test_so59, test_so60, test_so61,
         test_so62, test_so63, test_so64, test_so65, test_so66, test_so67,
         test_so68, test_so69, test_so70, test_so71, test_so72, test_so73,
         test_so74, test_so75, test_so76, test_so77, test_so78, test_so79,
         test_so80, test_so81, test_so82, test_so83, test_so84, test_so85,
         test_so86, test_so87, test_so88, test_so89, test_so90, test_so91,
         test_so92, test_so93, test_so94, test_so95, test_so96, test_so97,
         test_so98, test_so99, test_so100;
  wire   test_so3, test_so4, test_so5, test_so23, test_so57, test_so63,
         test_so73, test_so99, test_so100, n2230, n2217, n2231, n2374, n2361,
         n2375, DFF_2_n1, n4264, n2445, n2446, n2440, n2426, n2670, n2671,
         n2669, n2685, n2686, n2684, n2718, n2719, n2717, n2982, g2124, n2981,
         n2985, g1430, n2984, n2988, g744, n2987, n2991, g56, n2990, n3742,
         n3741, n8104, g16802, n8103, DFF_1_n1, g16823, n8102, g2950, n4423,
         n4274, g2883, n4330, g22026, g2888, g23358, g2896, n4431, g24473,
         g2892, g25201, g2903, n4305, g26037, g2900, n4291, g26798, g2908,
         n4355, n4273, g2912, n4482, g23357, g2917, n4479, g24476, g2924,
         n4349, g25199, g2920, n4280, DFF_15_n1, n4281, n8099, DFF_16_n1,
         n8098, DFF_18_n1, n4279, g2879, n4351, g2934, g2935, g2938, g2941,
         g2944, g2947, g2953, g2956, g2959, g2962, g2963, g2969, g2972, g2975,
         g2978, g2981, g2874, g18754, g1506, n4288, g18781, g1501, n4565,
         g18803, g1496, n4557, g18821, g1491, n4326, g18835, g1486, n4390,
         g18852, g1481, n4320, g18866, g1476, n4374, g18883, g1471, n4378,
         g21880, g2877, g19154, g813, n4289, g19163, g809, n4567, g19173, g805,
         n4559, g19184, g801, n4327, g20310, g797, n4391, g20343, g793, n4321,
         g20376, g789, n4375, g20417, g785, n4379, g21878, g2873, g19153, g125,
         n4290, g19162, g121, n4569, g19172, g117, n4561, g19144, g113, n4328,
         g19149, g109, n4392, g19157, g105, n4322, g19167, g101, n4376, g19178,
         g97, n4380, g20874, g2857, g18885, g2200, n4287, g18975, g2195, n4563,
         g18968, g2190, n4555, g18942, g2185, n4325, g18906, g2180, n4389,
         g18867, g2175, n4319, g18836, g2170, n4373, g18957, g2165, n4377,
         g21882, g2878, n4598, n4382, n4383, g3109, n4494, g18669, g18719,
         g3211, g18782, g3084, n4445, g17222, g3085, g17225, g3086, g17234,
         g3087, n4344, g17224, g3091, n4448, g17228, g3092, n4451, g17246,
         g3093, g17226, g3094, g17235, g3095, g17269, g3096, g25450, g3097,
         g25451, g3098, g25452, g3099, n4443, g28420, g3100, n4342, g28421,
         g28425, g3102, n4343, g29936, g3103, n4447, g29939, g3104, n4452,
         g29941, g3105, g30796, g3106, n4438, g30798, g3107, g30801, g3108,
         n4334, g17229, g3155, g17247, g3158, g17302, g3161, n4444, g17236,
         g3164, g17270, g3167, g17340, g3170, n4441, g17248, g3173, n4338,
         g17303, g3176, n4450, g17383, g17271, g3182, g17341, g3185, g17429,
         g3088, n8090, DFF_131_n1, n8089, DFF_132_n1, g3197, n8088, DFF_134_n1,
         g3201, n4406, g3204, g3207, n4329, g3188, n4405, g3133, n8087,
         DFF_140_n1, g3128, n8086, n8084, DFF_144_n1, g3124, n8083, DFF_146_n1,
         n8082, n8081, n8080, DFF_149_n1, g3112, g3110, g3111, n8079, n8078,
         n8077, DFF_155_n1, n8076, DFF_156_n1, g3151, n4424, g3142, n4301,
         g185, n4318, n4512, g165, n4369, g22100, g130, g22122, g131, g22141,
         g129, g22123, g133, g22142, g134, g22161, g132, g22025, g142, g22027,
         g143, g22030, g141, g22028, g145, g22031, g146, g22037, g22032, g148,
         g22038, g149, g22047, g147, g22039, g151, g22048, g152, g22063, g150,
         g22049, g154, g22064, g155, g22079, g153, g22065, g157, g22080, g158,
         g22101, g156, g22081, g160, g22102, g161, g22124, g159, g22103,
         g22125, g164, g22143, g162, g25204, g169, g25206, g170, g25211, g168,
         g25207, g172, g25212, g173, g25218, g171, g25213, g175, g25219, g176,
         g25228, g174, g25220, g178, g25229, g179, g25239, g177, g30261, g186,
         g30267, g30275, g192, g30637, g231, g30640, g234, g30645, g237,
         g30668, g195, g30674, g198, g30680, g201, g30641, g240, g30646, g243,
         g30653, g246, g30276, g204, g30284, g207, g30292, g210, g30254, g249,
         g30257, g252, g30262, g30245, g213, g30246, g216, g30248, g219,
         g30258, g258, g30263, g261, g30268, g264, g30635, g222, g30636, g225,
         g30639, g228, g30661, g267, g30669, g270, g30675, g273, g25027, g92,
         g25932, g88, g26529, g83, g27120, g27594, g74, g28145, g70, g28634,
         g65, g29109, g61, g29353, g29579, g52, g180, g181, n4506, g309, n4388,
         g27253, g354, g27255, g343, g27258, g27256, g369, g27259, g358,
         g27265, g361, g27260, g384, g27266, g373, g27277, g376, g27267, g398,
         g27278, g388, g27293, g391, g28732, g408, g28735, g411, g28744, g414,
         g29194, g417, g29197, g420, g29201, g423, g28736, g28745, g428,
         g28754, g426, g26803, g429, g26804, g432, g26807, g435, g26805, g438,
         g26808, g441, g26812, g444, g27759, g448, g27760, g449, g27762, g447,
         g29606, g312, g29608, g313, g29611, g314, g30699, g315, g30700,
         g30702, g317, g30455, g318, g30468, g319, g30482, g320, g29167, g322,
         g29169, g323, g29172, g321, g26655, g403, g26659, g404, g26664, g402,
         g450, n8066, DFF_299_n1, g452, n8065, DFF_301_n1, g454, DFF_303_n1,
         g280, n8062, DFF_305_n1, g282, n8061, DFF_307_n1, g284, n8060,
         DFF_309_n1, g286, n8059, DFF_311_n1, g288, n8058, DFF_313_n1, g290,
         n8057, n4485, n4282, n8056, g21346, g305, n4278, n8055, DFF_328_n1,
         g349, g350, g351, g352, g353, g357, g364, g365, g366, g367, g368,
         g372, g379, g380, g381, g383, g387, g394, g395, g396, g397, g324,
         g337, n4298, n4372, g550, n4313, g554, g18678, g557, n4360, g18726,
         g513, g523, g524, g455, g564, g569, g458, g570, g571, g461, g572,
         g573, g465, g574, g565, g566, g567, g471, g568, g489, n4461, g485,
         n4466, g23067, g486, g23093, g487, g23117, g488, g23385, g23399,
         g24174, g24178, g477, g24207, g478, g24216, g479, g23092, g480,
         g23000, g484, g23022, g464, g24206, g24215, g24228, g528, g535, g542,
         g13149, g543, g544, g21851, g548, g13111, g549, g499, n4541, g13160,
         g558, g559, g27261, g576, g27268, g577, g27279, g575, g27269, g579,
         g27280, g27294, g578, g27281, g582, g27295, g583, g27311, g581,
         g27296, g585, g27312, g586, g27327, g584, g24491, g587, g24498, g590,
         g24507, g593, g24499, g596, g24508, g599, g24519, g602, g28345, g614,
         g28349, g617, g28353, g28342, g605, g28344, g608, g28348, g611,
         g26541, g490, g26545, g493, g26553, g496, g506, n4570, g22578, n4571,
         g525, n8047, DFF_444_n1, n8046, DFF_445_n1, n8045, DFF_446_n1, n8044,
         DFF_447_n1, n8043, DFF_448_n1, DFF_449_n1, g536, g537, g24059, g538,
         n4492, n8040, n4359, g629, n4295, g16654, g630, g20314, g659, n4429,
         g20682, g640, n4404, g633, n4478, g23324, g653, n4422, g24426, g646,
         n4414, g25185, g660, n4403, g672, n4413, g26776, g27672, g679, n4477,
         g28199, g686, n4396, g28668, g692, n4418, g20875, g699, g20879, g700,
         g20891, g698, g20880, g702, g20892, g703, g20901, g701, g20893, g705,
         g20902, g706, g20921, g704, g20903, g708, g20922, g709, g20944, g707,
         g20923, g20945, g712, g20966, g710, g20946, g714, g20967, g715,
         g20989, g713, g20968, g717, g20990, g718, g21009, g716, g20991, g720,
         g21010, g721, g21031, g719, g21011, g723, g21032, g724, g21051, g722,
         g20876, g726, g20881, g20894, g725, g20924, g729, g20947, g730,
         g20969, g728, g20948, g732, g20970, g733, g20992, g731, g25260, g735,
         g25262, g736, g25266, g734, g22218, g738, g739, g22242, g737, n4323,
         n4312, g22126, g818, g22145, g819, g22162, g817, g22146, g821, g22163,
         g822, g22177, g820, g22029, g830, g22033, g831, g22040, g829, g22034,
         g833, g22041, g834, g22054, g832, g22042, g836, g22055, g837, g22066,
         g835, g22056, g22067, g840, g22087, g838, g22068, g842, g22088, g843,
         g22104, g841, g22089, g845, g22105, g846, g22127, g844, g22106, g848,
         g22128, g849, g22147, g847, g22129, g851, g22148, g852, g22164, g850,
         g25209, g857, g25214, g25221, g856, g25215, g860, g25222, g861,
         g25230, g859, g25223, g863, g25231, g864, g25240, g862, g25232, g866,
         g25241, g867, g25248, g865, g30269, g873, g30277, g876, g30285, g879,
         g30643, g918, g30648, g921, g30654, g30676, g882, g30681, g885,
         g30687, g888, g30649, g927, g30655, g930, g30662, g933, g30286, g891,
         g30293, g894, g30298, g897, g30259, g936, g30264, g939, g30270, g942,
         g30247, g900, g30249, g903, g30251, g906, g30265, g30271, g948,
         g30278, g951, g30638, g909, g30642, g912, g30647, g915, g30670, g954,
         g30677, g957, g30682, g960, g25042, g780, g25935, g776, g26530, g771,
         g27123, g767, g27603, g762, g28146, g758, g28635, g753, g29110,
         g29354, g29580, g740, g868, g869, n4363, n4364, g1088, n4381, g996,
         n4387, g27257, g1041, g27262, g1030, g27270, g1033, g27263, g1056,
         g27271, g1045, g27282, g1048, g27272, g27283, g1060, g27297, g1063,
         g27284, g1085, g27298, g1075, g27313, g1078, g28738, g1095, g28746,
         g1098, g28758, g1101, g29198, g1104, g29204, g1107, g29209, g1110,
         g28747, g1114, g28759, g1115, g28767, g1113, g26806, g1116, g26809,
         g26813, g1122, g26810, g1125, g26814, g1128, g26818, g1131, g27761,
         g1135, g27763, g1136, g27765, g1134, g29609, g999, g29612, g1000,
         g29616, g1001, g30701, g1002, g30703, g1003, g30705, g1004, g30470,
         g1005, g30485, g1006, g30500, g29170, g1009, g29173, g1010, g29179,
         g1008, g26661, g1090, g26665, g1091, g26669, g1089, g1137, n8027,
         DFF_649_n1, g1139, n8026, DFF_651_n1, g1141, n8025, DFF_653_n1, g967,
         n8024, DFF_655_n1, g969, DFF_657_n1, g971, n8021, DFF_659_n1, g973,
         n8020, DFF_661_n1, g975, n8019, DFF_663_n1, g977, n8018, n4486, n4283,
         g986, n4432, g992, n4277, n8017, g1029, g1036, g1037, g1038, g1040,
         g1044, g1051, g1052, g1053, g1054, g1055, g1059, g1066, g1067, g1068,
         g1069, g1070, g1074, g1081, g1083, g1084, g1011, g1024, n4371, n4316,
         g1236, n4300, g1240, g18707, g1243, n4353, g18763, g1196, n4304,
         g1199, g1209, g1210, g1142, g1255, g1145, g1256, g1257, g1148, g1258,
         g1259, g1152, g1260, g1251, g1155, g1252, g1253, g1158, g1254, g1176,
         n4460, n4459, g1172, n4465, g23081, g1173, g23111, g23126, g1175,
         g23392, g23406, g24179, g24181, g1164, g24213, g1165, g24223, g1166,
         g23110, g1167, g23014, g1171, g23039, g1151, g24212, g24222, g24235,
         g1214, g1221, g13155, g1229, n4549, n4361, g13124, g1235, g1186,
         n4548, g13171, g1244, g1245, g27273, g1262, g27285, g1263, g27299,
         g1261, g27286, g1265, g27300, g1266, g27314, g1264, g27301, g1268,
         g27315, g1269, g27328, g27316, g1271, g27329, g1272, g27339, g1270,
         g24501, g1273, g24510, g1276, g24521, g1279, g24511, g1282, g24522,
         g1285, g24532, g1288, g28351, g1300, g28355, g1303, g28360, g1306,
         g28346, g1291, g28350, g1294, g28354, g1297, g26547, g26557, g1180,
         g26569, g1183, g1192, n4454, g22615, n8009, DFF_783_n1, DFF_792_n1,
         g1211, n8008, DFF_794_n1, n8007, DFF_795_n1, n8006, DFF_796_n1, n8005,
         DFF_797_n1, n8004, DFF_798_n1, n8003, DFF_799_n1, g1222, g1223,
         g24072, g1224, n4489, n4358, g1315, n4294, g16671, g1316, g20333,
         g1345, n4428, g20717, g1326, n4402, g1319, n4476, g23329, g1339,
         n4421, g24430, g1332, n4412, g25189, g1346, n4401, g1358, n4411,
         g26781, g1352, n4469, g27678, g1365, n4475, g27718, g1372, n4395,
         g28321, g1378, n4417, g20882, g20896, g1386, g20910, g1384, g20897,
         g1388, g20911, g1389, g20925, g1387, g20912, g1391, g20926, g1392,
         g20949, g1390, g20927, g1394, g20950, g1395, g20972, g1393, g20951,
         g1397, g20973, g1398, g20993, g1396, g20974, g1400, g20994, g21015,
         g1399, g20995, g1403, g21016, g1404, g21033, g1402, g21017, g1406,
         g21034, g1407, g21052, g1405, g21035, g1409, g21053, g1410, g21070,
         g1408, g20883, g1412, g20898, g1413, g20913, g1411, g20952, g1415,
         g20975, g1416, g20996, g20976, g1418, g20997, g1419, g21018, g1417,
         g25263, g1421, g25267, g1422, g25270, g1420, g22234, g1424, g1425,
         g22263, g1423, n4317, n4515, g1547, n4368, g22149, g1512, g22166,
         g1513, g22178, g1511, g22167, g22179, g1516, g22191, g1514, g22035,
         g1524, g22043, g1525, g22057, g1523, g22044, g1527, g22058, g1528,
         g22073, g1526, g22059, g1530, g22074, g1531, g22090, g1529, g22075,
         g1533, g22091, g1534, g22112, g1532, g22092, g1536, g22113, g22130,
         g1535, g22114, g1539, g22131, g1540, g22150, g1538, g22132, g1542,
         g22151, g1543, g22168, g1541, g22152, g1545, g22169, g1546, g22180,
         g1544, g25217, g1551, g25224, g1552, g25233, g1550, g25225, g1554,
         g25234, g1555, g25242, g25235, g1557, g25243, g1558, g25249, g1556,
         g25244, g1560, g25250, g1561, g25255, g1559, g30279, g1567, g30287,
         g1570, g30294, g1573, g30651, g1612, g30657, g1615, g30663, g1618,
         g30683, g1576, g30688, g1579, g30692, g1582, g30658, g30664, g1624,
         g30671, g1627, g30295, g1585, g30299, g1588, g30302, g1591, g30266,
         g1630, g30272, g1633, g30280, g1636, g30250, g1594, g30252, g1597,
         g30255, g1600, g30273, g1639, g30281, g1642, g30288, g1645, g30644,
         g1603, g30650, g30656, g1609, g30678, g1648, g30684, g1651, g30689,
         g1654, g25056, g1466, g25938, g1462, g26531, g1457, g27129, g1453,
         g27612, g1448, g28147, g1444, g28636, g1439, g29111, g1435, g29355,
         g29581, g1426, g1562, g1563, n4518, g1690, n4386, g27264, g1735,
         g27274, g1724, g27287, g1727, g27275, g1750, g27288, g1739, g27302,
         g1742, g27289, g1765, g27303, g1754, g27317, g1757, g27304, g1779,
         g27318, g27330, g1772, g28749, g1789, g28760, g1792, g28771, g1795,
         g29205, g1798, g29212, g1801, g29218, g1804, g28761, g1808, g28772,
         g1809, g28778, g1807, g26811, g1810, g26815, g1813, g26820, g1816,
         g26816, g1819, g26821, g1822, g26824, g27764, g1829, g27766, g1830,
         g27768, g1828, g29613, g1693, g29617, g1694, g29620, g1695, g30704,
         g1696, g30706, g1697, g30708, g1698, g30487, g1699, g30503, g1700,
         g30338, g1701, g29178, g1703, g29181, g1704, g29184, g1702, g26667,
         g26670, g1785, g26675, g1783, g1831, n7988, DFF_999_n1, g1833, n7987,
         DFF_1001_n1, g1835, n7986, DFF_1003_n1, g1661, n7985, DFF_1005_n1,
         g1663, n7984, DFF_1007_n1, g1665, n7983, DFF_1009_n1, g1667,
         DFF_1011_n1, g1669, n7980, DFF_1013_n1, g1671, n7979, n4484, n4284,
         g1680, n4488, g1686, n4276, n7978, g1723, g1730, g1731, g1732, g1733,
         g1734, g1738, g1745, g1747, g1748, g1749, g1753, g1760, g1761, g1762,
         g1763, g1764, g1768, g1775, g1776, g1777, g1778, g1705, g1718, n4296,
         n4315, g1930, n4366, g1934, g18743, g1937, n4311, g18794, g1890,
         n4297, g1893, g1903, g1904, g1836, g1944, g1949, g1950, g1951, g1842,
         g1953, g1846, g1954, g1945, g1849, g1946, g1947, g1852, g1948, g1870,
         n4458, n4457, g1866, n4464, g23097, g1867, g23124, g1868, g23137,
         g1869, g23400, g23413, g24182, g24208, g1858, g24219, g1859, g24231,
         g1860, g23123, g1861, g23030, g1865, g23058, g1845, g24218, g24230,
         g24243, g1908, g1915, g1922, g13164, g1923, DFF_1099_n1, n7971,
         g13135, g1929, g1880, n4545, g13182, g1938, g1939, g27290, g1956,
         g27305, g1957, g27319, g1955, g27306, g1959, g27320, g1960, g27331,
         g1958, g27321, g1962, g27332, g1963, g27340, g1961, g27333, g27341,
         g1966, g27346, g1964, g24513, g1967, g24524, g1970, g24534, g1973,
         g24525, g1976, g24535, g1979, g24545, g1982, g28357, g1994, g28362,
         g1997, g28366, g2000, g28352, g1985, g28356, g1988, g28361, g1991,
         g26559, g26573, g1874, g26592, g1877, g1886, n4493, g22651, n7968,
         DFF_1133_n1, DFF_1142_n1, g1905, n7967, DFF_1144_n1, n7966,
         DFF_1145_n1, n7965, DFF_1146_n1, n7964, DFF_1147_n1, n7963,
         DFF_1148_n1, n7962, DFF_1149_n1, g1916, g1917, g24083, n7960, n4357,
         g2009, n4293, g16692, g2010, g20353, g2039, n4427, g20752, g2020,
         n4400, g2013, n4474, g23339, g2033, n4420, g24434, g2026, n4410,
         g25194, g2040, n4399, g2052, n4409, g26789, g2046, n4468, g27682,
         g2059, n4473, g27722, g28325, g2072, n4416, g20899, g2079, g20915,
         g2080, g20934, g2078, g20916, g2082, g20935, g2083, g20953, g2081,
         g20936, g2085, g20954, g2086, g20977, g2084, g20955, g2088, g20978,
         g2089, g20999, g2087, g20979, g2091, g21000, g21019, g2090, g21001,
         g2094, g21020, g2095, g21039, g2093, g21021, g2097, g21040, g2098,
         g21054, g2096, g21041, g2100, g21055, g2101, g21071, g2099, g21056,
         g2103, g21072, g2104, g21080, g2102, g20900, g2106, g20917, g20937,
         g2105, g20980, g2109, g21002, g2110, g21022, g2108, g21003, g2112,
         g21023, g2113, g21042, g2111, g25268, g2115, g25271, g2116, g25279,
         g2114, g22249, g2118, g2119, g22280, g2117, n4324, g2241, n4367,
         g22170, g2206, g22182, g2207, g22192, g2205, g22183, g2209, g22193,
         g2210, g22200, g2208, g22045, g2218, g22060, g2219, g22076, g2217,
         g22061, g2221, g22077, g2222, g22097, g2220, g22078, g2224, g22098,
         g22115, g2223, g22099, g2227, g22116, g2228, g22138, g2226, g22117,
         g2230, g22139, g2231, g22153, g2229, g22140, g2233, g22154, g2234,
         g22171, g2232, g22155, g2236, g22172, g2237, g22184, g2235, g22173,
         g2239, g22185, g22194, g2238, g25227, g2245, g25236, g2246, g25245,
         g2244, g25237, g2248, g25246, g2249, g25251, g2247, g25247, g2251,
         g25252, g2252, g25256, g2250, g25253, g2254, g25257, g2255, g25259,
         g2253, g30289, g2261, g30296, g30300, g2267, g30660, g2306, g30666,
         g2309, g30672, g2312, g30690, g2270, g30693, g2273, g30695, g2276,
         g30667, g2315, g30673, g2318, g30679, g2321, g30301, g2279, g30303,
         g2282, g30304, g2285, g30274, g2324, g30282, g30290, g2330, g30253,
         g2288, g30256, g2291, g30260, g2294, g30283, g2333, g30291, g2336,
         g30297, g2339, g30652, g2297, g30659, g2300, g30665, g2303, g30686,
         g2342, g30691, g2345, g30694, g2348, g25067, g2160, g25940, g26532,
         g2151, g27131, g2147, g27621, g2142, g28148, g2138, g28637, g2133,
         g29112, g2129, g29357, g29582, g2120, g2256, g2257, n4516, g27276,
         g2429, g27291, g2418, g27307, g2421, g27292, g2444, g27308, g2433,
         g27322, g2436, g27309, g2459, g27323, g2448, g27334, g2451, g27324,
         g2473, g27335, g2463, g27342, g2466, g28763, g2483, g28773, g2486,
         g28782, g29213, g2492, g29221, g2495, g29226, g2498, g28774, g2502,
         g28783, g2503, g28788, g2501, g26817, g2504, g26822, g2507, g26825,
         g2510, g26823, g2513, g26826, g2516, g26827, g2519, g27767, g2523,
         g27769, g2524, g27771, g29618, g2387, g29621, g2388, g29623, g2389,
         g30707, g2390, g30709, g2391, g30566, g2392, g30505, g2393, g30341,
         g2394, g30356, g2395, g29182, g2397, g29185, g2398, g29187, g2396,
         g26672, g2478, g26676, g2479, g26025, g2525, n7946, DFF_1349_n1,
         g2527, n7945, DFF_1351_n1, g2529, n7944, DFF_1353_n1, g2355, n7943,
         DFF_1355_n1, g2357, n7942, DFF_1357_n1, g2359, n7941, DFF_1359_n1,
         g2361, n7940, DFF_1361_n1, n7938, DFF_1363_n1, g2365, n7937, n4483,
         n4285, g2374, n4487, g30055, g2380, n4275, n7936, DFF_1378_n1, g2417,
         g2424, g2425, g2426, g2427, g2428, g2432, g2439, g2441, g2442, g2443,
         g2447, g2454, g2455, g2456, g2457, g2458, g2462, g2469, g2470, g2471,
         g2472, g2412, n4314, n4370, g2624, n4299, g2628, g18780, g2631, n4352,
         g18820, g2584, n4303, g2587, g2597, g2598, g2530, g2638, g2643, g2533,
         g2645, g2536, g2646, g2647, g2540, g2648, g2639, g2543, g2640, g2641,
         g2546, g2642, g2564, n4456, n4455, g2560, n4463, g23114, g2561,
         g23133, g2562, g21970, g23407, g23418, g24209, g24214, g2552, g24226,
         g2553, g24238, g2554, g23132, g2555, g23047, g2559, g23076, g2539,
         g24225, g24237, g24250, g2602, g2609, g13175, g2617, n7930, g30072,
         n7929, g13143, g2623, g2574, n4543, g13194, g2632, g2633, g27310,
         g2650, g27325, g2651, g27336, g2649, g27326, g2653, g27337, g2654,
         g27343, g2652, g27338, g2656, g27344, g27347, g2655, g27345, g2659,
         g27348, g2660, g27354, g2658, g24527, g2661, g24537, g2664, g24547,
         g2667, g24538, g2670, g24548, g2673, g24557, g2676, g28364, g2688,
         g28368, g2691, g28371, g2694, g28358, g2679, g28363, g28367, g2685,
         g26575, g2565, g26596, g2568, g26616, g2571, g2580, g22687, n7926,
         g30061, g2599, n7925, DFF_1494_n1, n7924, DFF_1495_n1, n7923,
         DFF_1496_n1, n7922, DFF_1497_n1, n7921, DFF_1498_n1, n7920,
         DFF_1499_n1, g2611, g24092, g2612, n4490, n7918, g2703, n4292, g16718,
         g2704, g20375, g2733, n4426, g20789, g2714, n4398, g2707, n4472,
         g23348, g2727, n4419, g24438, g2720, n4408, g25197, g2734, n4397,
         g2746, n4407, g26795, g27243, g2753, n4471, g27724, g2760, n4393,
         g28328, g2766, n4415, g20918, g2773, g20939, g2774, g20962, g2772,
         g20940, g2776, g20963, g2777, g20981, g2775, g20964, g2779, g20982,
         g2780, g21004, g2778, g20983, g2782, g21005, g2783, g21025, g21006,
         g2785, g21026, g2786, g21043, g2784, g21027, g2788, g21044, g2789,
         g21060, g2787, g21045, g2791, g21061, g2792, g21073, g2790, g21062,
         g2794, g21074, g2795, g21081, g2793, g21075, g2797, g21082, g2798,
         g21094, g20919, g2800, g20941, g2801, g20965, g2799, g21007, g2803,
         g21028, g2804, g21046, g2802, g21029, g2806, g21047, g2807, g21063,
         g2805, g25272, g2809, g25280, g2810, g25288, g2808, g22269, g2812,
         g22284, g2813, g22299, g20877, n7913, DFF_1561_n1, g20884, n7912,
         DFF_1562_n1, n4263, n4269, g3043, n4268, g3044, n4267, g3045, n4266,
         g3046, n4265, g3047, n4272, g3048, n4271, g3049, n4270, g3050, n4259,
         g3051, n4236, g3052, n4239, g3053, n4237, n4234, g3056, n4233, g3057,
         n4238, g3058, n4235, g3059, n4240, g3060, n4232, g3061, n4245, g3062,
         n4248, g3063, n4246, g3064, n4243, g3065, n4242, g3066, n4247, g3067,
         n4244, g3068, n4249, g3069, n4241, n4254, g3071, n4257, g3072, n4255,
         g3073, n4252, g3074, n4251, g3075, n4256, g3076, n4253, g3077, n4258,
         g3078, n4250, g2997, g25265, g2993, g26048, n7909, g3006, g24445,
         g3002, g25191, g3013, g26031, g26786, g3024, n4262, g3018, n4481,
         g3028, n4350, g24446, g3036, n4480, g25202, g3032, n7907, DFF_1612_n1,
         g2987, n4365, g16824, g16844, g16853, g16860, g16803, g16835, g16851,
         g16857, g16866, g3083, n4261, N995, n4577, g16845, g16854, g16861,
         g16880, g18755, g18804, g18837, g18868, g18907, g2990, N690, n4578,
         n4260, n4309, n4308, n4307, n4306, n4524, n4525, n4511, n4509, n4499,
         n4520, n3683, n3887, n3686, n3890, n3692, n3896, n4513, n3897, n3424,
         n3427, n3433, n4529, n4530, n4522, n4523, n4521, n3171, n3159, n3163,
         n3893, n3690, n3689, n3431, n3430, n3168, n3160, n3164, n3172, n4527,
         n4528, n4526, n3167, n3894, n3888, n3891, n2302, n2289, n2303, n2275,
         n4066, n4065, n4606, n4618, n4640, n2568, n3196, n3212, n3225, n3237,
         n3936, n4034, n4033, n4037, n4038, n4043, n4046, n3252, n3254, n3038,
         n3070, n3102, n3130, n2800, n2798, n2616, n2594, n3940, n3705, n3933,
         n3939, n3445, n3457, n3469, n3478, n3700, n4058, n4101, n3938, n4182,
         n4073, n3417, n4057, n4122, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4,
         Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         Tj_Trigger, RingOscENable1, RingOscENable2, RingOscENable3,
         RingOscENable, Out29, Out1, Out2, Out3, Out4, Out5, Out6, Out7, Out8,
         Out9, Out10, Out11, Out12, Out13, Out14, Out15, Out16, Out17, Out18,
         Out19, Out20, Out21, Out22, Out23, Out24, Out25, Out26, Out27, Out28,
         n10, n19, n91, n148, n244, n266, n270, n279, n309, n437, n438, n453,
         n475, n497, n498, n499, n512, n513, n514, n515, n520, n567, n596,
         n597, n653, n808, n822, n826, n872, n901, n902, n959, n1114, n1137,
         n1141, n1186, n1214, n1215, n1261, n1392, n1402, n1423, n1427, n1502,
         n1503, n1538, n1540, n1543, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7406, n7429, n7430, n7431, n7432, n7433, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7615, n7617, n7618, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7705,
         n7706, n7707, n7708, n7709, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7908, n7910, n7911,
         n7914, n7915, n7916, n7917, n7919, n7927, n7928, n7931, n7932, n7933,
         n7934, n7935, n7939, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7961, n7969, n7970, n7972,
         n7973, n7974, n7975, n7976, n7977, n7981, n7982, n7989, n7990, n7991,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8001, n8002, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8022, n8023, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8042, n8048, n8049, n8050, n8051, n8053, n8054, n8063, n8064, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8085, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8100, n8101, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, U3772_n1, U3776_n1, U3777_n1,
         U3778_n1, U3779_n1, U3780_n1, U3781_n1, U3782_n1, U3783_n1, U3784_n1,
         U3785_n1, U3786_n1, U3787_n1, U3901_n1, U3902_n1, U4467_n1, U4904_n1,
         U4930_n1, U5128_n1, U5141_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1,
         U5753_n1, U5754_n1, U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1,
         U5760_n1, U5761_n1, U5762_n1, U5763_n1, U5764_n1, U5882_n1, U5939_n1,
         U5940_n1, U5941_n1, U5942_n1, U6140_n1, U6460_n1, U6470_n1, U6562_n1,
         U6563_n1, U6718_n1, U7116_n1, U7118_n1, U7293_n1;
  assign g8251 = test_so3;
  assign g7519 = test_so4;
  assign g4450 = test_so5;
  assign g7909 = test_so23;
  assign g5612 = test_so57;
  assign g5695 = test_so63;
  assign g7084 = test_so73;
  assign g8270 = test_so99;
  assign g8258 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(g51), .SI(test_si1), .SE(n8133), .CLK(n8320), .Q(
        n8104), .QN(n14350) );
  SDFFX1 DFF_1_Q_reg ( .D(g16802), .SI(n8104), .SE(n8133), .CLK(n8320), .Q(
        n8103), .QN(DFF_1_n1) );
  SDFFX1 DFF_2_Q_reg ( .D(g16823), .SI(n8103), .SE(n8133), .CLK(n8320), .Q(
        n8102), .QN(DFF_2_n1) );
  SDFFX1 DFF_3_Q_reg ( .D(n4264), .SI(n8102), .SE(n8133), .CLK(n8320), .Q(
        g2950), .QN(n4423) );
  SDFFX1 DFF_4_Q_reg ( .D(n4274), .SI(g2950), .SE(n8134), .CLK(n8321), .Q(
        g2883), .QN(n4330) );
  SDFFX1 DFF_5_Q_reg ( .D(g22026), .SI(g2883), .SE(n8134), .CLK(n8321), .Q(
        g2888), .QN(n8016) );
  SDFFX1 DFF_6_Q_reg ( .D(g23358), .SI(g2888), .SE(n8134), .CLK(n8321), .Q(
        g2896), .QN(n4431) );
  SDFFX1 DFF_7_Q_reg ( .D(g24473), .SI(g2896), .SE(n8134), .CLK(n8321), .Q(
        g2892), .QN(n7752) );
  SDFFX1 DFF_8_Q_reg ( .D(g25201), .SI(g2892), .SE(n8134), .CLK(n8321), .Q(
        g2903), .QN(n4305) );
  SDFFX1 DFF_9_Q_reg ( .D(g26037), .SI(g2903), .SE(n8134), .CLK(n8321), .Q(
        g2900), .QN(n4291) );
  SDFFX1 DFF_10_Q_reg ( .D(g26798), .SI(g2900), .SE(n8134), .CLK(n8321), .Q(
        g2908), .QN(n4355) );
  SDFFX1 DFF_11_Q_reg ( .D(n4273), .SI(g2908), .SE(n8134), .CLK(n8321), .Q(
        g2912), .QN(n4482) );
  SDFFX1 DFF_12_Q_reg ( .D(g23357), .SI(g2912), .SE(n8134), .CLK(n8321), .Q(
        g2917), .QN(n4479) );
  SDFFX1 DFF_13_Q_reg ( .D(g24476), .SI(g2917), .SE(n8134), .CLK(n8321), .Q(
        g2924), .QN(n4349) );
  SDFFX1 DFF_14_Q_reg ( .D(g25199), .SI(g2924), .SE(n8134), .CLK(n8321), .Q(
        g2920), .QN(n7703) );
  SDFFX1 DFF_15_Q_reg ( .D(n4280), .SI(g2920), .SE(n8134), .CLK(n8321), .Q(
        test_so1), .QN(DFF_15_n1) );
  SDFFX1 DFF_16_Q_reg ( .D(n4281), .SI(test_si2), .SE(n8131), .CLK(n8318), .Q(
        n8099), .QN(DFF_16_n1) );
  SDFFX1 DFF_17_Q_reg ( .D(g51), .SI(n8099), .SE(n8131), .CLK(n8318), .Q(g8021) );
  SDFFX1 DFF_18_Q_reg ( .D(g8021), .SI(g8021), .SE(n8131), .CLK(n8318), .Q(
        n8098), .QN(DFF_18_n1) );
  SDFFX1 DFF_19_Q_reg ( .D(n4279), .SI(n8098), .SE(n8131), .CLK(n8318), .Q(
        g2879), .QN(n4351) );
  SDFFX1 DFF_20_Q_reg ( .D(g3212), .SI(g2879), .SE(n8131), .CLK(n8318), .Q(
        g2934), .QN(n8014) );
  SDFFX1 DFF_21_Q_reg ( .D(g3228), .SI(g2934), .SE(n8131), .CLK(n8318), .Q(
        g2935), .QN(n7982) );
  SDFFX1 DFF_22_Q_reg ( .D(g3227), .SI(g2935), .SE(n8132), .CLK(n8319), .Q(
        g2938), .QN(n7989) );
  SDFFX1 DFF_23_Q_reg ( .D(g3226), .SI(g2938), .SE(n8132), .CLK(n8319), .Q(
        g2941), .QN(n7977) );
  SDFFX1 DFF_24_Q_reg ( .D(g3225), .SI(g2941), .SE(n8132), .CLK(n8319), .Q(
        g2944) );
  SDFFX1 DFF_25_Q_reg ( .D(g3224), .SI(g2944), .SE(n8132), .CLK(n8319), .Q(
        g2947), .QN(n7990) );
  SDFFX1 DFF_26_Q_reg ( .D(g3223), .SI(g2947), .SE(n8132), .CLK(n8319), .Q(
        g2953), .QN(n7991) );
  SDFFX1 DFF_27_Q_reg ( .D(g3222), .SI(g2953), .SE(n8132), .CLK(n8319), .Q(
        g2956), .QN(n7993) );
  SDFFX1 DFF_28_Q_reg ( .D(g3221), .SI(g2956), .SE(n8132), .CLK(n8319), .Q(
        g2959), .QN(n7981) );
  SDFFX1 DFF_29_Q_reg ( .D(g3232), .SI(g2959), .SE(n8132), .CLK(n8319), .Q(
        g2962), .QN(n8012) );
  SDFFX1 DFF_30_Q_reg ( .D(g3220), .SI(g2962), .SE(n8132), .CLK(n8319), .Q(
        g2963), .QN(n7996) );
  SDFFX1 DFF_31_Q_reg ( .D(g3219), .SI(g2963), .SE(n8132), .CLK(n8319), .Q(
        test_so2) );
  SDFFX1 DFF_32_Q_reg ( .D(g3218), .SI(test_si3), .SE(n8131), .CLK(n8318), .Q(
        g2969), .QN(n7999) );
  SDFFX1 DFF_33_Q_reg ( .D(g3217), .SI(g2969), .SE(n8131), .CLK(n8318), .Q(
        g2972), .QN(n7997) );
  SDFFX1 DFF_34_Q_reg ( .D(g3216), .SI(g2972), .SE(n8131), .CLK(n8318), .Q(
        g2975), .QN(n7998) );
  SDFFX1 DFF_35_Q_reg ( .D(g3215), .SI(g2975), .SE(n8131), .CLK(n8318), .Q(
        g2978), .QN(n7994) );
  SDFFX1 DFF_36_Q_reg ( .D(g3214), .SI(g2978), .SE(n8131), .CLK(n8318), .Q(
        g2981) );
  SDFFX1 DFF_37_Q_reg ( .D(g3213), .SI(g2981), .SE(n8131), .CLK(n8318), .Q(
        g2874), .QN(n7995) );
  SDFFX1 DFF_38_Q_reg ( .D(g18754), .SI(g2874), .SE(n8132), .CLK(n8319), .Q(
        g1506), .QN(n4288) );
  SDFFX1 DFF_39_Q_reg ( .D(g18781), .SI(g1506), .SE(n8132), .CLK(n8319), .Q(
        g1501), .QN(n4565) );
  SDFFX1 DFF_40_Q_reg ( .D(g18803), .SI(g1501), .SE(n8133), .CLK(n8320), .Q(
        g1496), .QN(n4557) );
  SDFFX1 DFF_41_Q_reg ( .D(g18821), .SI(g1496), .SE(n8133), .CLK(n8320), .Q(
        g1491), .QN(n4326) );
  SDFFX1 DFF_42_Q_reg ( .D(g18835), .SI(g1491), .SE(n8133), .CLK(n8320), .Q(
        g1486), .QN(n4390) );
  SDFFX1 DFF_43_Q_reg ( .D(g18852), .SI(g1486), .SE(n8133), .CLK(n8320), .Q(
        g1481), .QN(n4320) );
  SDFFX1 DFF_44_Q_reg ( .D(g18866), .SI(g1481), .SE(n8133), .CLK(n8320), .Q(
        g1476), .QN(n4374) );
  SDFFX1 DFF_45_Q_reg ( .D(g18883), .SI(g1476), .SE(n8133), .CLK(n8320), .Q(
        g1471), .QN(n4378) );
  SDFFX1 DFF_46_Q_reg ( .D(g21880), .SI(g1471), .SE(n8138), .CLK(n8325), .Q(
        g2877) );
  SDFFX1 DFF_47_Q_reg ( .D(g19154), .SI(g2877), .SE(n8138), .CLK(n8325), .Q(
        test_so3) );
  SDFFX1 DFF_48_Q_reg ( .D(test_so3), .SI(test_si4), .SE(n8138), .CLK(n8325), 
        .Q(g813), .QN(n4289) );
  SDFFX1 DFF_49_Q_reg ( .D(g19163), .SI(g813), .SE(n8138), .CLK(n8325), .Q(
        g4090) );
  SDFFX1 DFF_50_Q_reg ( .D(g4090), .SI(g4090), .SE(n8138), .CLK(n8325), .Q(
        g809), .QN(n4567) );
  SDFFX1 DFF_51_Q_reg ( .D(g19173), .SI(g809), .SE(n8139), .CLK(n8326), .Q(
        g4323) );
  SDFFX1 DFF_52_Q_reg ( .D(g4323), .SI(g4323), .SE(n8139), .CLK(n8326), .Q(
        g805), .QN(n4559) );
  SDFFX1 DFF_53_Q_reg ( .D(g19184), .SI(g805), .SE(n8139), .CLK(n8326), .Q(
        g4590) );
  SDFFX1 DFF_54_Q_reg ( .D(g4590), .SI(g4590), .SE(n8139), .CLK(n8326), .Q(
        g801), .QN(n4327) );
  SDFFX1 DFF_55_Q_reg ( .D(g20310), .SI(g801), .SE(n8139), .CLK(n8326), .Q(
        g6225) );
  SDFFX1 DFF_56_Q_reg ( .D(g6225), .SI(g6225), .SE(n8139), .CLK(n8326), .Q(
        g797), .QN(n4391) );
  SDFFX1 DFF_57_Q_reg ( .D(g20343), .SI(g797), .SE(n8139), .CLK(n8326), .Q(
        g6442) );
  SDFFX1 DFF_58_Q_reg ( .D(g6442), .SI(g6442), .SE(n8139), .CLK(n8326), .Q(
        g793), .QN(n4321) );
  SDFFX1 DFF_59_Q_reg ( .D(g20376), .SI(g793), .SE(n8139), .CLK(n8326), .Q(
        g6895) );
  SDFFX1 DFF_60_Q_reg ( .D(g6895), .SI(g6895), .SE(n8139), .CLK(n8326), .Q(
        g789), .QN(n4375) );
  SDFFX1 DFF_61_Q_reg ( .D(g20417), .SI(g789), .SE(n8139), .CLK(n8326), .Q(
        g7334) );
  SDFFX1 DFF_62_Q_reg ( .D(g7334), .SI(g7334), .SE(n8139), .CLK(n8326), .Q(
        g785), .QN(n4379) );
  SDFFX1 DFF_63_Q_reg ( .D(g21878), .SI(g785), .SE(n8140), .CLK(n8327), .Q(
        test_so4) );
  SDFFX1 DFF_64_Q_reg ( .D(test_so4), .SI(test_si5), .SE(n8140), .CLK(n8327), 
        .Q(g2873) );
  SDFFX1 DFF_65_Q_reg ( .D(g19153), .SI(g2873), .SE(n8140), .CLK(n8327), .Q(
        g8249) );
  SDFFX1 DFF_66_Q_reg ( .D(g8249), .SI(g8249), .SE(n8140), .CLK(n8327), .Q(
        g125), .QN(n4290) );
  SDFFX1 DFF_67_Q_reg ( .D(g19162), .SI(g125), .SE(n8141), .CLK(n8328), .Q(
        g4088) );
  SDFFX1 DFF_68_Q_reg ( .D(g4088), .SI(g4088), .SE(n8141), .CLK(n8328), .Q(
        g121), .QN(n4569) );
  SDFFX1 DFF_69_Q_reg ( .D(g19172), .SI(g121), .SE(n8141), .CLK(n8328), .Q(
        g4321) );
  SDFFX1 DFF_70_Q_reg ( .D(g4321), .SI(g4321), .SE(n8141), .CLK(n8328), .Q(
        g117), .QN(n4561) );
  SDFFX1 DFF_71_Q_reg ( .D(g19144), .SI(g117), .SE(n8141), .CLK(n8328), .Q(
        g8023) );
  SDFFX1 DFF_72_Q_reg ( .D(g8023), .SI(g8023), .SE(n8141), .CLK(n8328), .Q(
        g113), .QN(n4328) );
  SDFFX1 DFF_73_Q_reg ( .D(g19149), .SI(g113), .SE(n8141), .CLK(n8328), .Q(
        g8175) );
  SDFFX1 DFF_74_Q_reg ( .D(g8175), .SI(g8175), .SE(n8141), .CLK(n8328), .Q(
        g109), .QN(n4392) );
  SDFFX1 DFF_75_Q_reg ( .D(g19157), .SI(g109), .SE(n8141), .CLK(n8328), .Q(
        g3993) );
  SDFFX1 DFF_76_Q_reg ( .D(g3993), .SI(g3993), .SE(n8141), .CLK(n8328), .Q(
        g105), .QN(n4322) );
  SDFFX1 DFF_77_Q_reg ( .D(g19167), .SI(g105), .SE(n8141), .CLK(n8328), .Q(
        g4200) );
  SDFFX1 DFF_78_Q_reg ( .D(g4200), .SI(g4200), .SE(n8141), .CLK(n8328), .Q(
        g101), .QN(n4376) );
  SDFFX1 DFF_79_Q_reg ( .D(g19178), .SI(g101), .SE(n8142), .CLK(n8329), .Q(
        test_so5) );
  SDFFX1 DFF_80_Q_reg ( .D(test_so5), .SI(test_si6), .SE(n8142), .CLK(n8329), 
        .Q(g97), .QN(n4380) );
  SDFFX1 DFF_81_Q_reg ( .D(g20874), .SI(g97), .SE(n8142), .CLK(n8329), .Q(
        g8096) );
  SDFFX1 DFF_82_Q_reg ( .D(g8096), .SI(g8096), .SE(n8142), .CLK(n8329), .Q(
        g2857) );
  SDFFX1 DFF_83_Q_reg ( .D(g18885), .SI(g2857), .SE(n8142), .CLK(n8329), .Q(
        g2200), .QN(n4287) );
  SDFFX1 DFF_84_Q_reg ( .D(g18975), .SI(g2200), .SE(n8142), .CLK(n8329), .Q(
        g2195), .QN(n4563) );
  SDFFX1 DFF_85_Q_reg ( .D(g18968), .SI(g2195), .SE(n8142), .CLK(n8329), .Q(
        g2190), .QN(n4555) );
  SDFFX1 DFF_86_Q_reg ( .D(g18942), .SI(g2190), .SE(n8142), .CLK(n8329), .Q(
        g2185), .QN(n4325) );
  SDFFX1 DFF_87_Q_reg ( .D(g18906), .SI(g2185), .SE(n8142), .CLK(n8329), .Q(
        g2180), .QN(n4389) );
  SDFFX1 DFF_88_Q_reg ( .D(g18867), .SI(g2180), .SE(n8142), .CLK(n8329), .Q(
        g2175), .QN(n4319) );
  SDFFX1 DFF_89_Q_reg ( .D(g18836), .SI(g2175), .SE(n8142), .CLK(n8329), .Q(
        g2170), .QN(n4373) );
  SDFFX1 DFF_90_Q_reg ( .D(g18957), .SI(g2170), .SE(n8142), .CLK(n8329), .Q(
        g2165), .QN(n4377) );
  SDFFX1 DFF_91_Q_reg ( .D(g21882), .SI(g2165), .SE(n8164), .CLK(n8351), .Q(
        g2878) );
  SDFFX1 DFF_92_Q_reg ( .D(n4598), .SI(g2878), .SE(n8256), .CLK(n8443), .Q(
        g8106), .QN(n4382) );
  SDFFX1 DFF_93_Q_reg ( .D(g8106), .SI(g8106), .SE(n8256), .CLK(n8443), .Q(
        g8030), .QN(n4383) );
  SDFFX1 DFF_94_Q_reg ( .D(g8030), .SI(g8030), .SE(n8256), .CLK(n8443), .Q(
        g3109), .QN(n4494) );
  SDFFX1 DFF_95_Q_reg ( .D(g18669), .SI(g3109), .SE(n8257), .CLK(n8444), .Q(
        test_so6) );
  SDFFX1 DFF_96_Q_reg ( .D(g18719), .SI(test_si7), .SE(n8257), .CLK(n8444), 
        .Q(g3211) );
  SDFFX1 DFF_97_Q_reg ( .D(g18782), .SI(g3211), .SE(n8257), .CLK(n8444), .Q(
        g3084), .QN(n4445) );
  SDFFX1 DFF_98_Q_reg ( .D(g17222), .SI(g3084), .SE(n8259), .CLK(n8446), .Q(
        g3085) );
  SDFFX1 DFF_99_Q_reg ( .D(g17225), .SI(g3085), .SE(n8259), .CLK(n8446), .Q(
        g3086) );
  SDFFX1 DFF_100_Q_reg ( .D(g17234), .SI(g3086), .SE(n8259), .CLK(n8446), .Q(
        g3087), .QN(n4344) );
  SDFFX1 DFF_101_Q_reg ( .D(g17224), .SI(g3087), .SE(n8259), .CLK(n8446), .Q(
        g3091), .QN(n4448) );
  SDFFX1 DFF_102_Q_reg ( .D(g17228), .SI(g3091), .SE(n8259), .CLK(n8446), .Q(
        g3092), .QN(n4451) );
  SDFFX1 DFF_103_Q_reg ( .D(g17246), .SI(g3092), .SE(n8259), .CLK(n8446), .Q(
        g3093) );
  SDFFX1 DFF_104_Q_reg ( .D(g17226), .SI(g3093), .SE(n8259), .CLK(n8446), .Q(
        g3094) );
  SDFFX1 DFF_105_Q_reg ( .D(g17235), .SI(g3094), .SE(n8259), .CLK(n8446), .Q(
        g3095) );
  SDFFX1 DFF_106_Q_reg ( .D(g17269), .SI(g3095), .SE(n8135), .CLK(n8322), .Q(
        g3096) );
  SDFFX1 DFF_107_Q_reg ( .D(g25450), .SI(g3096), .SE(n8257), .CLK(n8444), .Q(
        g3097) );
  SDFFX1 DFF_108_Q_reg ( .D(g25451), .SI(g3097), .SE(n8257), .CLK(n8444), .Q(
        g3098) );
  SDFFX1 DFF_109_Q_reg ( .D(g25452), .SI(g3098), .SE(n8257), .CLK(n8444), .Q(
        g3099), .QN(n4443) );
  SDFFX1 DFF_110_Q_reg ( .D(g28420), .SI(g3099), .SE(n8257), .CLK(n8444), .Q(
        g3100), .QN(n4342) );
  SDFFX1 DFF_111_Q_reg ( .D(g28421), .SI(g3100), .SE(n8258), .CLK(n8445), .Q(
        test_so7) );
  SDFFX1 DFF_112_Q_reg ( .D(g28425), .SI(test_si8), .SE(n8257), .CLK(n8444), 
        .Q(g3102), .QN(n4343) );
  SDFFX1 DFF_113_Q_reg ( .D(g29936), .SI(g3102), .SE(n8258), .CLK(n8445), .Q(
        g3103), .QN(n4447) );
  SDFFX1 DFF_114_Q_reg ( .D(g29939), .SI(g3103), .SE(n8258), .CLK(n8445), .Q(
        g3104), .QN(n4452) );
  SDFFX1 DFF_115_Q_reg ( .D(g29941), .SI(g3104), .SE(n8258), .CLK(n8445), .Q(
        g3105) );
  SDFFX1 DFF_116_Q_reg ( .D(g30796), .SI(g3105), .SE(n8258), .CLK(n8445), .Q(
        g3106), .QN(n4438) );
  SDFFX1 DFF_117_Q_reg ( .D(g30798), .SI(g3106), .SE(n8258), .CLK(n8445), .Q(
        g3107) );
  SDFFX1 DFF_118_Q_reg ( .D(g30801), .SI(g3107), .SE(n8258), .CLK(n8445), .Q(
        g3108), .QN(n4334) );
  SDFFX1 DFF_119_Q_reg ( .D(g17229), .SI(g3108), .SE(n8258), .CLK(n8445), .Q(
        g3155) );
  SDFFX1 DFF_120_Q_reg ( .D(g17247), .SI(g3155), .SE(n8258), .CLK(n8445), .Q(
        g3158) );
  SDFFX1 DFF_121_Q_reg ( .D(g17302), .SI(g3158), .SE(n8258), .CLK(n8445), .Q(
        g3161), .QN(n4444) );
  SDFFX1 DFF_122_Q_reg ( .D(g17236), .SI(g3161), .SE(n8258), .CLK(n8445), .Q(
        g3164) );
  SDFFX1 DFF_123_Q_reg ( .D(g17270), .SI(g3164), .SE(n8258), .CLK(n8445), .Q(
        g3167) );
  SDFFX1 DFF_124_Q_reg ( .D(g17340), .SI(g3167), .SE(n8259), .CLK(n8446), .Q(
        g3170), .QN(n4441) );
  SDFFX1 DFF_125_Q_reg ( .D(g17248), .SI(g3170), .SE(n8259), .CLK(n8446), .Q(
        g3173), .QN(n4338) );
  SDFFX1 DFF_126_Q_reg ( .D(g17303), .SI(g3173), .SE(n8259), .CLK(n8446), .Q(
        g3176), .QN(n4450) );
  SDFFX1 DFF_127_Q_reg ( .D(g17383), .SI(g3176), .SE(n8259), .CLK(n8446), .Q(
        test_so8) );
  SDFFX1 DFF_128_Q_reg ( .D(g17271), .SI(test_si9), .SE(n8257), .CLK(n8444), 
        .Q(g3182) );
  SDFFX1 DFF_129_Q_reg ( .D(g17341), .SI(g3182), .SE(n8257), .CLK(n8444), .Q(
        g3185) );
  SDFFX1 DFF_130_Q_reg ( .D(g17429), .SI(g3185), .SE(n8257), .CLK(n8444), .Q(
        g3088) );
  SDFFX1 DFF_131_Q_reg ( .D(g24734), .SI(g3088), .SE(n8257), .CLK(n8444), .Q(
        n8090), .QN(DFF_131_n1) );
  SDFFX1 DFF_132_Q_reg ( .D(g25442), .SI(n8090), .SE(n8136), .CLK(n8323), .Q(
        n8089), .QN(DFF_132_n1) );
  SDFFX1 DFF_133_Q_reg ( .D(g25435), .SI(n8089), .SE(n8260), .CLK(n8447), .Q(
        g3197) );
  SDFFX1 DFF_134_Q_reg ( .D(g25420), .SI(g3197), .SE(n8260), .CLK(n8447), .Q(
        n8088), .QN(DFF_134_n1) );
  SDFFX1 DFF_135_Q_reg ( .D(g26149), .SI(n8088), .SE(n8135), .CLK(n8322), .Q(
        g3201), .QN(n4406) );
  SDFFX1 DFF_136_Q_reg ( .D(g26135), .SI(g3201), .SE(n8135), .CLK(n8322), .Q(
        g3204), .QN(n8015) );
  SDFFX1 DFF_137_Q_reg ( .D(g26104), .SI(g3204), .SE(n8135), .CLK(n8322), .Q(
        g3207), .QN(n4329) );
  SDFFX1 DFF_138_Q_reg ( .D(g27380), .SI(g3207), .SE(n8136), .CLK(n8323), .Q(
        g3188), .QN(n4405) );
  SDFFX1 DFF_139_Q_reg ( .D(n91), .SI(g3188), .SE(n8136), .CLK(n8323), .Q(
        g3133), .QN(n7430) );
  SDFFX1 DFF_140_Q_reg ( .D(g26104), .SI(g3133), .SE(n8136), .CLK(n8323), .Q(
        n8087), .QN(DFF_140_n1) );
  SDFFX1 DFF_141_Q_reg ( .D(n244), .SI(n8087), .SE(n8136), .CLK(n8323), .Q(
        g3128) );
  SDFFX1 DFF_142_Q_reg ( .D(g26149), .SI(g3128), .SE(n8136), .CLK(n8323), .Q(
        n8086) );
  SDFFX1 DFF_143_Q_reg ( .D(g25420), .SI(n8086), .SE(n8137), .CLK(n8324), .Q(
        test_so9) );
  SDFFX1 DFF_144_Q_reg ( .D(n270), .SI(test_si10), .SE(n8136), .CLK(n8323), 
        .Q(n8084), .QN(DFF_144_n1) );
  SDFFX1 DFF_145_Q_reg ( .D(g25442), .SI(n8084), .SE(n8136), .CLK(n8323), .Q(
        g3124) );
  SDFFX1 DFF_146_Q_reg ( .D(n279), .SI(g3124), .SE(n8136), .CLK(n8323), .Q(
        n8083), .QN(DFF_146_n1) );
  SDFFX1 DFF_147_Q_reg ( .D(g26104), .SI(n8083), .SE(n8136), .CLK(n8323), .Q(
        n8082), .QN(n14349) );
  SDFFX1 DFF_148_Q_reg ( .D(g26135), .SI(n8082), .SE(n8137), .CLK(n8324), .Q(
        n8081), .QN(n14351) );
  SDFFX1 DFF_149_Q_reg ( .D(g26149), .SI(n8081), .SE(n8137), .CLK(n8324), .Q(
        n8080), .QN(DFF_149_n1) );
  SDFFX1 DFF_150_Q_reg ( .D(g25420), .SI(n8080), .SE(n8137), .CLK(n8324), .Q(
        g3112) );
  SDFFX1 DFF_151_Q_reg ( .D(g25435), .SI(g3112), .SE(n8137), .CLK(n8324), .Q(
        g3110) );
  SDFFX1 DFF_152_Q_reg ( .D(g25442), .SI(g3110), .SE(n8137), .CLK(n8324), .Q(
        g3111) );
  SDFFX1 DFF_153_Q_reg ( .D(g27380), .SI(g3111), .SE(n8137), .CLK(n8324), .Q(
        n8079), .QN(n14352) );
  SDFFX1 DFF_154_Q_reg ( .D(g26104), .SI(n8079), .SE(n8137), .CLK(n8324), .Q(
        n8078), .QN(n14353) );
  SDFFX1 DFF_155_Q_reg ( .D(g26135), .SI(n8078), .SE(n8137), .CLK(n8324), .Q(
        n8077), .QN(DFF_155_n1) );
  SDFFX1 DFF_156_Q_reg ( .D(g26149), .SI(n8077), .SE(n8137), .CLK(n8324), .Q(
        n8076), .QN(DFF_156_n1) );
  SDFFX1 DFF_157_Q_reg ( .D(g27380), .SI(n8076), .SE(n8137), .CLK(n8324), .Q(
        g3151), .QN(n4424) );
  SDFFX1 DFF_158_Q_reg ( .D(g26104), .SI(g3151), .SE(n8137), .CLK(n8324), .Q(
        g3142), .QN(n4301) );
  SDFFX1 DFF_159_Q_reg ( .D(g26135), .SI(g3142), .SE(n8138), .CLK(n8325), .Q(
        test_so10), .QN(n8095) );
  SDFFX1 DFF_160_Q_reg ( .D(n91), .SI(test_si11), .SE(n8135), .CLK(n8322), .Q(
        g185) );
  SDFFX1 DFF_161_Q_reg ( .D(g2950), .SI(g185), .SE(n8135), .CLK(n8322), .Q(
        g6231), .QN(n4318) );
  SDFFX1 DFF_162_Q_reg ( .D(g6231), .SI(g6231), .SE(n8136), .CLK(n8323), .Q(
        g6313), .QN(n4512) );
  SDFFX1 DFF_163_Q_reg ( .D(g6313), .SI(g6313), .SE(n8136), .CLK(n8323), .Q(
        g165), .QN(n4369) );
  SDFFX1 DFF_164_Q_reg ( .D(g22100), .SI(g165), .SE(n8149), .CLK(n8336), .Q(
        g130), .QN(n7952) );
  SDFFX1 DFF_165_Q_reg ( .D(g22122), .SI(g130), .SE(n8149), .CLK(n8336), .Q(
        g131), .QN(n7951) );
  SDFFX1 DFF_166_Q_reg ( .D(g22141), .SI(g131), .SE(n8150), .CLK(n8337), .Q(
        g129), .QN(n7554) );
  SDFFX1 DFF_167_Q_reg ( .D(g22123), .SI(g129), .SE(n8150), .CLK(n8337), .Q(
        g133), .QN(n7950) );
  SDFFX1 DFF_168_Q_reg ( .D(g22142), .SI(g133), .SE(n8150), .CLK(n8337), .Q(
        g134), .QN(n7949) );
  SDFFX1 DFF_169_Q_reg ( .D(g22161), .SI(g134), .SE(n8150), .CLK(n8337), .Q(
        g132), .QN(n7553) );
  SDFFX1 DFF_170_Q_reg ( .D(g22025), .SI(g132), .SE(n8150), .CLK(n8337), .Q(
        g142), .QN(n7948) );
  SDFFX1 DFF_171_Q_reg ( .D(g22027), .SI(g142), .SE(n8150), .CLK(n8337), .Q(
        g143), .QN(n7947) );
  SDFFX1 DFF_172_Q_reg ( .D(g22030), .SI(g143), .SE(n8150), .CLK(n8337), .Q(
        g141), .QN(n7552) );
  SDFFX1 DFF_173_Q_reg ( .D(g22028), .SI(g141), .SE(n8150), .CLK(n8337), .Q(
        g145), .QN(n7939) );
  SDFFX1 DFF_174_Q_reg ( .D(g22031), .SI(g145), .SE(n8150), .CLK(n8337), .Q(
        g146), .QN(n7935) );
  SDFFX1 DFF_175_Q_reg ( .D(g22037), .SI(g146), .SE(n8150), .CLK(n8337), .Q(
        test_so11), .QN(n8115) );
  SDFFX1 DFF_176_Q_reg ( .D(g22032), .SI(test_si12), .SE(n8148), .CLK(n8335), 
        .Q(g148), .QN(n7934) );
  SDFFX1 DFF_177_Q_reg ( .D(g22038), .SI(g148), .SE(n8148), .CLK(n8335), .Q(
        g149), .QN(n7933) );
  SDFFX1 DFF_178_Q_reg ( .D(g22047), .SI(g149), .SE(n8149), .CLK(n8336), .Q(
        g147), .QN(n7551) );
  SDFFX1 DFF_179_Q_reg ( .D(g22039), .SI(g147), .SE(n8149), .CLK(n8336), .Q(
        g151), .QN(n7932) );
  SDFFX1 DFF_180_Q_reg ( .D(g22048), .SI(g151), .SE(n8149), .CLK(n8336), .Q(
        g152), .QN(n7931) );
  SDFFX1 DFF_181_Q_reg ( .D(g22063), .SI(g152), .SE(n8149), .CLK(n8336), .Q(
        g150), .QN(n7550) );
  SDFFX1 DFF_182_Q_reg ( .D(g22049), .SI(g150), .SE(n8149), .CLK(n8336), .Q(
        g154), .QN(n7928) );
  SDFFX1 DFF_183_Q_reg ( .D(g22064), .SI(g154), .SE(n8149), .CLK(n8336), .Q(
        g155), .QN(n7927) );
  SDFFX1 DFF_184_Q_reg ( .D(g22079), .SI(g155), .SE(n8149), .CLK(n8336), .Q(
        g153), .QN(n7549) );
  SDFFX1 DFF_185_Q_reg ( .D(g22065), .SI(g153), .SE(n8145), .CLK(n8332), .Q(
        g157), .QN(n7919) );
  SDFFX1 DFF_186_Q_reg ( .D(g22080), .SI(g157), .SE(n8147), .CLK(n8334), .Q(
        g158), .QN(n7917) );
  SDFFX1 DFF_187_Q_reg ( .D(g22101), .SI(g158), .SE(n8147), .CLK(n8334), .Q(
        g156), .QN(n7548) );
  SDFFX1 DFF_188_Q_reg ( .D(g22081), .SI(g156), .SE(n8149), .CLK(n8336), .Q(
        g160), .QN(n7510) );
  SDFFX1 DFF_189_Q_reg ( .D(g22102), .SI(g160), .SE(n8149), .CLK(n8336), .Q(
        g161), .QN(n7509) );
  SDFFX1 DFF_190_Q_reg ( .D(g22124), .SI(g161), .SE(n8149), .CLK(n8336), .Q(
        g159), .QN(n7508) );
  SDFFX1 DFF_191_Q_reg ( .D(g22103), .SI(g159), .SE(n8150), .CLK(n8337), .Q(
        test_so12), .QN(n8114) );
  SDFFX1 DFF_192_Q_reg ( .D(g22125), .SI(test_si13), .SE(n8147), .CLK(n8334), 
        .Q(g164), .QN(n7547) );
  SDFFX1 DFF_193_Q_reg ( .D(g22143), .SI(g164), .SE(n8147), .CLK(n8334), .Q(
        g162), .QN(n7546) );
  SDFFX1 DFF_194_Q_reg ( .D(g25204), .SI(g162), .SE(n8147), .CLK(n8334), .Q(
        g169), .QN(n7612) );
  SDFFX1 DFF_195_Q_reg ( .D(g25206), .SI(g169), .SE(n8147), .CLK(n8334), .Q(
        g170), .QN(n7611) );
  SDFFX1 DFF_196_Q_reg ( .D(g25211), .SI(g170), .SE(n8148), .CLK(n8335), .Q(
        g168), .QN(n7610) );
  SDFFX1 DFF_197_Q_reg ( .D(g25207), .SI(g168), .SE(n8148), .CLK(n8335), .Q(
        g172), .QN(n7609) );
  SDFFX1 DFF_198_Q_reg ( .D(g25212), .SI(g172), .SE(n8148), .CLK(n8335), .Q(
        g173), .QN(n7608) );
  SDFFX1 DFF_199_Q_reg ( .D(g25218), .SI(g173), .SE(n8148), .CLK(n8335), .Q(
        g171), .QN(n7607) );
  SDFFX1 DFF_200_Q_reg ( .D(g25213), .SI(g171), .SE(n8148), .CLK(n8335), .Q(
        g175), .QN(n7606) );
  SDFFX1 DFF_201_Q_reg ( .D(g25219), .SI(g175), .SE(n8148), .CLK(n8335), .Q(
        g176), .QN(n7605) );
  SDFFX1 DFF_202_Q_reg ( .D(g25228), .SI(g176), .SE(n8148), .CLK(n8335), .Q(
        g174), .QN(n7604) );
  SDFFX1 DFF_203_Q_reg ( .D(g25220), .SI(g174), .SE(n8148), .CLK(n8335), .Q(
        g178), .QN(n7603) );
  SDFFX1 DFF_204_Q_reg ( .D(g25229), .SI(g178), .SE(n8148), .CLK(n8335), .Q(
        g179), .QN(n7602) );
  SDFFX1 DFF_205_Q_reg ( .D(g25239), .SI(g179), .SE(n8148), .CLK(n8335), .Q(
        g177), .QN(n7601) );
  SDFFX1 DFF_206_Q_reg ( .D(g30261), .SI(g177), .SE(n8155), .CLK(n8342), .Q(
        g186) );
  SDFFX1 DFF_207_Q_reg ( .D(g30267), .SI(g186), .SE(n8155), .CLK(n8342), .Q(
        test_so13) );
  SDFFX1 DFF_208_Q_reg ( .D(g30275), .SI(test_si14), .SE(n8155), .CLK(n8342), 
        .Q(g192) );
  SDFFX1 DFF_209_Q_reg ( .D(g30637), .SI(g192), .SE(n8155), .CLK(n8342), .Q(
        g231) );
  SDFFX1 DFF_210_Q_reg ( .D(g30640), .SI(g231), .SE(n8156), .CLK(n8343), .Q(
        g234) );
  SDFFX1 DFF_211_Q_reg ( .D(g30645), .SI(g234), .SE(n8156), .CLK(n8343), .Q(
        g237) );
  SDFFX1 DFF_212_Q_reg ( .D(g30668), .SI(g237), .SE(n8156), .CLK(n8343), .Q(
        g195) );
  SDFFX1 DFF_213_Q_reg ( .D(g30674), .SI(g195), .SE(n8156), .CLK(n8343), .Q(
        g198) );
  SDFFX1 DFF_214_Q_reg ( .D(g30680), .SI(g198), .SE(n8151), .CLK(n8338), .Q(
        g201) );
  SDFFX1 DFF_215_Q_reg ( .D(g30641), .SI(g201), .SE(n8151), .CLK(n8338), .Q(
        g240) );
  SDFFX1 DFF_216_Q_reg ( .D(g30646), .SI(g240), .SE(n8151), .CLK(n8338), .Q(
        g243) );
  SDFFX1 DFF_217_Q_reg ( .D(g30653), .SI(g243), .SE(n8150), .CLK(n8337), .Q(
        g246) );
  SDFFX1 DFF_218_Q_reg ( .D(g30276), .SI(g246), .SE(n8151), .CLK(n8338), .Q(
        g204) );
  SDFFX1 DFF_219_Q_reg ( .D(g30284), .SI(g204), .SE(n8151), .CLK(n8338), .Q(
        g207) );
  SDFFX1 DFF_220_Q_reg ( .D(g30292), .SI(g207), .SE(n8151), .CLK(n8338), .Q(
        g210) );
  SDFFX1 DFF_221_Q_reg ( .D(g30254), .SI(g210), .SE(n8154), .CLK(n8341), .Q(
        g249) );
  SDFFX1 DFF_222_Q_reg ( .D(g30257), .SI(g249), .SE(n8154), .CLK(n8341), .Q(
        g252) );
  SDFFX1 DFF_223_Q_reg ( .D(g30262), .SI(g252), .SE(n8154), .CLK(n8341), .Q(
        test_so14) );
  SDFFX1 DFF_224_Q_reg ( .D(g30245), .SI(test_si15), .SE(n8154), .CLK(n8341), 
        .Q(g213) );
  SDFFX1 DFF_225_Q_reg ( .D(g30246), .SI(g213), .SE(n8154), .CLK(n8341), .Q(
        g216) );
  SDFFX1 DFF_226_Q_reg ( .D(g30248), .SI(g216), .SE(n8154), .CLK(n8341), .Q(
        g219) );
  SDFFX1 DFF_227_Q_reg ( .D(g30258), .SI(g219), .SE(n8155), .CLK(n8342), .Q(
        g258) );
  SDFFX1 DFF_228_Q_reg ( .D(g30263), .SI(g258), .SE(n8155), .CLK(n8342), .Q(
        g261) );
  SDFFX1 DFF_229_Q_reg ( .D(g30268), .SI(g261), .SE(n8155), .CLK(n8342), .Q(
        g264) );
  SDFFX1 DFF_230_Q_reg ( .D(g30635), .SI(g264), .SE(n8155), .CLK(n8342), .Q(
        g222) );
  SDFFX1 DFF_231_Q_reg ( .D(g30636), .SI(g222), .SE(n8155), .CLK(n8342), .Q(
        g225) );
  SDFFX1 DFF_232_Q_reg ( .D(g30639), .SI(g225), .SE(n8155), .CLK(n8342), .Q(
        g228) );
  SDFFX1 DFF_233_Q_reg ( .D(g30661), .SI(g228), .SE(n8155), .CLK(n8342), .Q(
        g267) );
  SDFFX1 DFF_234_Q_reg ( .D(g30669), .SI(g267), .SE(n8155), .CLK(n8342), .Q(
        g270) );
  SDFFX1 DFF_235_Q_reg ( .D(g30675), .SI(g270), .SE(n8145), .CLK(n8332), .Q(
        g273) );
  SDFFX1 DFF_236_Q_reg ( .D(g25027), .SI(g273), .SE(n8145), .CLK(n8332), .Q(
        g92), .QN(n7702) );
  SDFFX1 DFF_237_Q_reg ( .D(g25932), .SI(g92), .SE(n8146), .CLK(n8333), .Q(g88) );
  SDFFX1 DFF_238_Q_reg ( .D(g26529), .SI(g88), .SE(n8146), .CLK(n8333), .Q(g83), .QN(n7701) );
  SDFFX1 DFF_239_Q_reg ( .D(g27120), .SI(g83), .SE(n8146), .CLK(n8333), .Q(
        test_so15) );
  SDFFX1 DFF_240_Q_reg ( .D(g27594), .SI(test_si16), .SE(n8146), .CLK(n8333), 
        .Q(g74), .QN(n7700) );
  SDFFX1 DFF_241_Q_reg ( .D(g28145), .SI(g74), .SE(n8146), .CLK(n8333), .Q(g70), .QN(n8067) );
  SDFFX1 DFF_242_Q_reg ( .D(g28634), .SI(g70), .SE(n8146), .CLK(n8333), .Q(g65), .QN(n7699) );
  SDFFX1 DFF_243_Q_reg ( .D(g29109), .SI(g65), .SE(n8146), .CLK(n8333), .Q(g61), .QN(n8048) );
  SDFFX1 DFF_244_Q_reg ( .D(g29353), .SI(g61), .SE(n8146), .CLK(n8333), .Q(g56), .QN(n7325) );
  SDFFX1 DFF_245_Q_reg ( .D(g29579), .SI(g56), .SE(n8146), .CLK(n8333), .Q(g52), .QN(n7164) );
  SDFFX1 DFF_246_Q_reg ( .D(n19), .SI(g52), .SE(n8146), .CLK(n8333), .Q(g180)
         );
  SDFFX1 DFF_247_Q_reg ( .D(g180), .SI(g180), .SE(n8146), .CLK(n8333), .Q(
        g5549) );
  SDFFX1 DFF_248_Q_reg ( .D(g5549), .SI(g5549), .SE(n8146), .CLK(n8333), .Q(
        g181), .QN(n7709) );
  SDFFX1 DFF_251_Q_reg ( .D(g6447), .SI(g6447), .SE(n8147), .CLK(n8334), .Q(
        n4640), .QN(n4506) );
  SDFFX1 DFF_252_Q_reg ( .D(g5549), .SI(n4640), .SE(n8147), .CLK(n8334), .Q(
        g309), .QN(n4388) );
  SDFFX1 DFF_253_Q_reg ( .D(g27253), .SI(g309), .SE(n8153), .CLK(n8340), .Q(
        g354), .QN(n7653) );
  SDFFX1 DFF_254_Q_reg ( .D(g27255), .SI(g354), .SE(n8153), .CLK(n8340), .Q(
        g343), .QN(n7652) );
  SDFFX1 DFF_255_Q_reg ( .D(g27258), .SI(g343), .SE(n8153), .CLK(n8340), .Q(
        test_so16), .QN(n8100) );
  SDFFX1 DFF_256_Q_reg ( .D(g27256), .SI(test_si17), .SE(n8153), .CLK(n8340), 
        .Q(g369), .QN(n7631) );
  SDFFX1 DFF_257_Q_reg ( .D(g27259), .SI(g369), .SE(n8154), .CLK(n8341), .Q(
        g358), .QN(n7630) );
  SDFFX1 DFF_258_Q_reg ( .D(g27265), .SI(g358), .SE(n8154), .CLK(n8341), .Q(
        g361), .QN(n7629) );
  SDFFX1 DFF_259_Q_reg ( .D(g27260), .SI(g361), .SE(n8154), .CLK(n8341), .Q(
        g384), .QN(n7379) );
  SDFFX1 DFF_260_Q_reg ( .D(g27266), .SI(g384), .SE(n8154), .CLK(n8341), .Q(
        g373), .QN(n7381) );
  SDFFX1 DFF_261_Q_reg ( .D(g27277), .SI(g373), .SE(n8153), .CLK(n8340), .Q(
        g376), .QN(n7380) );
  SDFFX1 DFF_262_Q_reg ( .D(g27267), .SI(g376), .SE(n8154), .CLK(n8341), .Q(
        g398), .QN(n7642) );
  SDFFX1 DFF_263_Q_reg ( .D(g27278), .SI(g398), .SE(n8154), .CLK(n8341), .Q(
        g388), .QN(n7641) );
  SDFFX1 DFF_264_Q_reg ( .D(g27293), .SI(g388), .SE(n8151), .CLK(n8338), .Q(
        g391), .QN(n7640) );
  SDFFX1 DFF_265_Q_reg ( .D(g28732), .SI(g391), .SE(n8151), .CLK(n8338), .Q(
        g408) );
  SDFFX1 DFF_266_Q_reg ( .D(g28735), .SI(g408), .SE(n8153), .CLK(n8340), .Q(
        g411) );
  SDFFX1 DFF_267_Q_reg ( .D(g28744), .SI(g411), .SE(n8153), .CLK(n8340), .Q(
        g414) );
  SDFFX1 DFF_268_Q_reg ( .D(g29194), .SI(g414), .SE(n8153), .CLK(n8340), .Q(
        g417) );
  SDFFX1 DFF_269_Q_reg ( .D(g29197), .SI(g417), .SE(n8153), .CLK(n8340), .Q(
        g420) );
  SDFFX1 DFF_270_Q_reg ( .D(g29201), .SI(g420), .SE(n8151), .CLK(n8338), .Q(
        g423) );
  SDFFX1 DFF_271_Q_reg ( .D(g28736), .SI(g423), .SE(n8152), .CLK(n8339), .Q(
        test_so17), .QN(n8106) );
  SDFFX1 DFF_272_Q_reg ( .D(g28745), .SI(test_si18), .SE(n8152), .CLK(n8339), 
        .Q(g428), .QN(n7685) );
  SDFFX1 DFF_273_Q_reg ( .D(g28754), .SI(g428), .SE(n8152), .CLK(n8339), .Q(
        g426), .QN(n7684) );
  SDFFX1 DFF_274_Q_reg ( .D(g26803), .SI(g426), .SE(n8152), .CLK(n8339), .Q(
        g429) );
  SDFFX1 DFF_275_Q_reg ( .D(g26804), .SI(g429), .SE(n8152), .CLK(n8339), .Q(
        g432) );
  SDFFX1 DFF_276_Q_reg ( .D(g26807), .SI(g432), .SE(n8152), .CLK(n8339), .Q(
        g435) );
  SDFFX1 DFF_277_Q_reg ( .D(g26805), .SI(g435), .SE(n8152), .CLK(n8339), .Q(
        g438) );
  SDFFX1 DFF_278_Q_reg ( .D(g26808), .SI(g438), .SE(n8152), .CLK(n8339), .Q(
        g441) );
  SDFFX1 DFF_279_Q_reg ( .D(g26812), .SI(g441), .SE(n8152), .CLK(n8339), .Q(
        g444) );
  SDFFX1 DFF_280_Q_reg ( .D(g27759), .SI(g444), .SE(n8153), .CLK(n8340), .Q(
        g448), .QN(n7683) );
  SDFFX1 DFF_281_Q_reg ( .D(g27760), .SI(g448), .SE(n8153), .CLK(n8340), .Q(
        g449), .QN(n7682) );
  SDFFX1 DFF_282_Q_reg ( .D(g27762), .SI(g449), .SE(n8152), .CLK(n8339), .Q(
        g447), .QN(n7681) );
  SDFFX1 DFF_283_Q_reg ( .D(g29606), .SI(g447), .SE(n8152), .CLK(n8339), .Q(
        g312), .QN(n7289) );
  SDFFX1 DFF_284_Q_reg ( .D(g29608), .SI(g312), .SE(n8152), .CLK(n8339), .Q(
        g313), .QN(n7288) );
  SDFFX1 DFF_285_Q_reg ( .D(g29611), .SI(g313), .SE(n8151), .CLK(n8338), .Q(
        g314), .QN(n7287) );
  SDFFX1 DFF_286_Q_reg ( .D(g30699), .SI(g314), .SE(n8151), .CLK(n8338), .Q(
        g315), .QN(n7286) );
  SDFFX1 DFF_287_Q_reg ( .D(g30700), .SI(g315), .SE(n8151), .CLK(n8338), .Q(
        test_so18), .QN(n8128) );
  SDFFX1 DFF_288_Q_reg ( .D(g30702), .SI(test_si19), .SE(n8145), .CLK(n8332), 
        .Q(g317), .QN(n7285) );
  SDFFX1 DFF_289_Q_reg ( .D(g30455), .SI(g317), .SE(n8147), .CLK(n8334), .Q(
        g318), .QN(n7284) );
  SDFFX1 DFF_290_Q_reg ( .D(g30468), .SI(g318), .SE(n8147), .CLK(n8334), .Q(
        g319), .QN(n7283) );
  SDFFX1 DFF_291_Q_reg ( .D(g30482), .SI(g319), .SE(n8145), .CLK(n8332), .Q(
        g320), .QN(n7282) );
  SDFFX1 DFF_292_Q_reg ( .D(g29167), .SI(g320), .SE(n8156), .CLK(n8343), .Q(
        g322), .QN(n7321) );
  SDFFX1 DFF_293_Q_reg ( .D(g29169), .SI(g322), .SE(n8156), .CLK(n8343), .Q(
        g323), .QN(n7320) );
  SDFFX1 DFF_294_Q_reg ( .D(g29172), .SI(g323), .SE(n8156), .CLK(n8343), .Q(
        g321), .QN(n7319) );
  SDFFX1 DFF_295_Q_reg ( .D(g26655), .SI(g321), .SE(n8156), .CLK(n8343), .Q(
        g403), .QN(n7680) );
  SDFFX1 DFF_296_Q_reg ( .D(g26659), .SI(g403), .SE(n8156), .CLK(n8343), .Q(
        g404), .QN(n7679) );
  SDFFX1 DFF_297_Q_reg ( .D(g26664), .SI(g404), .SE(n8156), .CLK(n8343), .Q(
        g402), .QN(n7678) );
  SDFFX1 DFF_298_Q_reg ( .D(n4290), .SI(g402), .SE(n8163), .CLK(n8350), .Q(
        g450) );
  SDFFX1 DFF_299_Q_reg ( .D(g450), .SI(g450), .SE(n8163), .CLK(n8350), .Q(
        n8066), .QN(DFF_299_n1) );
  SDFFX1 DFF_300_Q_reg ( .D(n4569), .SI(n8066), .SE(n8163), .CLK(n8350), .Q(
        g452) );
  SDFFX1 DFF_301_Q_reg ( .D(g452), .SI(g452), .SE(n8163), .CLK(n8350), .Q(
        n8065), .QN(DFF_301_n1) );
  SDFFX1 DFF_302_Q_reg ( .D(n4561), .SI(n8065), .SE(n8163), .CLK(n8350), .Q(
        g454) );
  SDFFX1 DFF_303_Q_reg ( .D(g454), .SI(g454), .SE(n8163), .CLK(n8350), .Q(
        test_so19), .QN(DFF_303_n1) );
  SDFFX1 DFF_304_Q_reg ( .D(n4328), .SI(test_si20), .SE(n8144), .CLK(n8331), 
        .Q(g280) );
  SDFFX1 DFF_305_Q_reg ( .D(g280), .SI(g280), .SE(n8144), .CLK(n8331), .Q(
        n8062), .QN(DFF_305_n1) );
  SDFFX1 DFF_306_Q_reg ( .D(n4392), .SI(n8062), .SE(n8144), .CLK(n8331), .Q(
        g282) );
  SDFFX1 DFF_307_Q_reg ( .D(g282), .SI(g282), .SE(n8144), .CLK(n8331), .Q(
        n8061), .QN(DFF_307_n1) );
  SDFFX1 DFF_308_Q_reg ( .D(n4322), .SI(n8061), .SE(n8144), .CLK(n8331), .Q(
        g284) );
  SDFFX1 DFF_309_Q_reg ( .D(g284), .SI(g284), .SE(n8144), .CLK(n8331), .Q(
        n8060), .QN(DFF_309_n1) );
  SDFFX1 DFF_310_Q_reg ( .D(n4376), .SI(n8060), .SE(n8144), .CLK(n8331), .Q(
        g286) );
  SDFFX1 DFF_311_Q_reg ( .D(g286), .SI(g286), .SE(n8145), .CLK(n8332), .Q(
        n8059), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(n4380), .SI(n8059), .SE(n8145), .CLK(n8332), .Q(
        g288) );
  SDFFX1 DFF_313_Q_reg ( .D(g288), .SI(g288), .SE(n8145), .CLK(n8332), .Q(
        n8058), .QN(DFF_313_n1) );
  SDFFX1 DFF_314_Q_reg ( .D(g2857), .SI(n8058), .SE(n8145), .CLK(n8332), .Q(
        g290) );
  SDFFX1 DFF_315_Q_reg ( .D(g290), .SI(g290), .SE(n8145), .CLK(n8332), .Q(
        n8057), .QN(n4485) );
  SDFFX1 DFF_316_Q_reg ( .D(n4282), .SI(n8057), .SE(n8153), .CLK(n8340), .Q(
        n8056), .QN(n14355) );
  SDFFX1 DFF_317_Q_reg ( .D(g21346), .SI(n8056), .SE(n8163), .CLK(n8350), .Q(
        g305), .QN(n7433) );
  SDFFX1 DFF_328_Q_reg ( .D(n4278), .SI(g305), .SE(n8156), .CLK(n8343), .Q(
        n8055), .QN(DFF_328_n1) );
  SDFFX1 DFF_329_Q_reg ( .D(g354), .SI(n8055), .SE(n8156), .CLK(n8343), .Q(
        test_so20) );
  SDFFX1 DFF_330_Q_reg ( .D(test_so20), .SI(test_si21), .SE(n8157), .CLK(n8344), .Q(g349) );
  SDFFX1 DFF_331_Q_reg ( .D(g343), .SI(g349), .SE(n8157), .CLK(n8344), .Q(g350) );
  SDFFX1 DFF_332_Q_reg ( .D(g350), .SI(g350), .SE(n8157), .CLK(n8344), .Q(g351) );
  SDFFX1 DFF_333_Q_reg ( .D(test_so16), .SI(g351), .SE(n8157), .CLK(n8344), 
        .Q(g352) );
  SDFFX1 DFF_334_Q_reg ( .D(g352), .SI(g352), .SE(n8157), .CLK(n8344), .Q(g353) );
  SDFFX1 DFF_335_Q_reg ( .D(g369), .SI(g353), .SE(n8157), .CLK(n8344), .Q(g357) );
  SDFFX1 DFF_336_Q_reg ( .D(g357), .SI(g357), .SE(n8157), .CLK(n8344), .Q(g364) );
  SDFFX1 DFF_337_Q_reg ( .D(g358), .SI(g364), .SE(n8157), .CLK(n8344), .Q(g365) );
  SDFFX1 DFF_338_Q_reg ( .D(g365), .SI(g365), .SE(n8157), .CLK(n8344), .Q(g366) );
  SDFFX1 DFF_339_Q_reg ( .D(g361), .SI(g366), .SE(n8157), .CLK(n8344), .Q(g367) );
  SDFFX1 DFF_340_Q_reg ( .D(g367), .SI(g367), .SE(n8157), .CLK(n8344), .Q(g368) );
  SDFFX1 DFF_341_Q_reg ( .D(g384), .SI(g368), .SE(n8157), .CLK(n8344), .Q(g372) );
  SDFFX1 DFF_342_Q_reg ( .D(g372), .SI(g372), .SE(n8158), .CLK(n8345), .Q(g379) );
  SDFFX1 DFF_343_Q_reg ( .D(g373), .SI(g379), .SE(n8158), .CLK(n8345), .Q(g380) );
  SDFFX1 DFF_344_Q_reg ( .D(g380), .SI(g380), .SE(n8158), .CLK(n8345), .Q(g381) );
  SDFFX1 DFF_345_Q_reg ( .D(g376), .SI(g381), .SE(n8158), .CLK(n8345), .Q(
        test_so21) );
  SDFFX1 DFF_346_Q_reg ( .D(test_so21), .SI(test_si22), .SE(n8158), .CLK(n8345), .Q(g383) );
  SDFFX1 DFF_347_Q_reg ( .D(g398), .SI(g383), .SE(n8158), .CLK(n8345), .Q(g387) );
  SDFFX1 DFF_348_Q_reg ( .D(g387), .SI(g387), .SE(n8158), .CLK(n8345), .Q(g394) );
  SDFFX1 DFF_349_Q_reg ( .D(g388), .SI(g394), .SE(n8158), .CLK(n8345), .Q(g395) );
  SDFFX1 DFF_350_Q_reg ( .D(g395), .SI(g395), .SE(n8158), .CLK(n8345), .Q(g396) );
  SDFFX1 DFF_351_Q_reg ( .D(g391), .SI(g396), .SE(n8158), .CLK(n8345), .Q(g397) );
  SDFFX1 DFF_352_Q_reg ( .D(g397), .SI(g397), .SE(n8158), .CLK(n8345), .Q(g324) );
  SDFFX1 DFF_353_Q_reg ( .D(n4598), .SI(g324), .SE(n8158), .CLK(n8345), .Q(
        g5629) );
  SDFFX1 DFF_354_Q_reg ( .D(g5629), .SI(g5629), .SE(n8159), .CLK(n8346), .Q(
        g5648) );
  SDFFX1 DFF_355_Q_reg ( .D(g5648), .SI(g5648), .SE(n8159), .CLK(n8346), .Q(
        g337) );
  SDFFX1 DFF_356_Q_reg ( .D(n4598), .SI(g337), .SE(n8159), .CLK(n8346), .Q(
        g6485), .QN(n4298) );
  SDFFX1 DFF_357_Q_reg ( .D(g6485), .SI(g6485), .SE(n8159), .CLK(n8346), .Q(
        g6642), .QN(n4372) );
  SDFFX1 DFF_358_Q_reg ( .D(g6642), .SI(g6642), .SE(n8159), .CLK(n8346), .Q(
        g550), .QN(n4313) );
  SDFFX1 DFF_359_Q_reg ( .D(n520), .SI(g550), .SE(n8165), .CLK(n8352), .Q(g554), .QN(n7972) );
  SDFFX1 DFF_360_Q_reg ( .D(g18678), .SI(g554), .SE(n8165), .CLK(n8352), .Q(
        g557), .QN(n4360) );
  SDFFX1 DFF_361_Q_reg ( .D(g18726), .SI(g557), .SE(n8166), .CLK(n8353), .Q(
        test_so22), .QN(n8091) );
  SDFFX1 DFF_362_Q_reg ( .D(n515), .SI(test_si23), .SE(n8159), .CLK(n8346), 
        .Q(g513) );
  SDFFX1 DFF_363_Q_reg ( .D(g513), .SI(g513), .SE(n8159), .CLK(n8346), .Q(g523) );
  SDFFX1 DFF_364_Q_reg ( .D(g523), .SI(g523), .SE(n8159), .CLK(n8346), .Q(g524) );
  SDFFX1 DFF_365_Q_reg ( .D(g455), .SI(g524), .SE(n8159), .CLK(n8346), .Q(g564) );
  SDFFX1 DFF_366_Q_reg ( .D(g564), .SI(g564), .SE(n8159), .CLK(n8346), .Q(g569) );
  SDFFX1 DFF_367_Q_reg ( .D(g458), .SI(g569), .SE(n8159), .CLK(n8346), .Q(g570) );
  SDFFX1 DFF_368_Q_reg ( .D(g570), .SI(g570), .SE(n8159), .CLK(n8346), .Q(g571) );
  SDFFX1 DFF_369_Q_reg ( .D(g461), .SI(g571), .SE(n8160), .CLK(n8347), .Q(g572) );
  SDFFX1 DFF_370_Q_reg ( .D(g572), .SI(g572), .SE(n8160), .CLK(n8347), .Q(g573) );
  SDFFX1 DFF_371_Q_reg ( .D(g465), .SI(g573), .SE(n8160), .CLK(n8347), .Q(g574) );
  SDFFX1 DFF_372_Q_reg ( .D(g574), .SI(g574), .SE(n8160), .CLK(n8347), .Q(g565) );
  SDFFX1 DFF_373_Q_reg ( .D(test_so24), .SI(g565), .SE(n8160), .CLK(n8347), 
        .Q(g566) );
  SDFFX1 DFF_374_Q_reg ( .D(g566), .SI(g566), .SE(n8160), .CLK(n8347), .Q(g567) );
  SDFFX1 DFF_375_Q_reg ( .D(g471), .SI(g567), .SE(n8160), .CLK(n8347), .Q(g568) );
  SDFFX1 DFF_376_Q_reg ( .D(g568), .SI(g568), .SE(n8160), .CLK(n8347), .Q(g489) );
  SDFFX1 DFF_377_Q_reg ( .D(g2950), .SI(g489), .SE(n8160), .CLK(n8347), .Q(
        test_so23), .QN(n8072) );
  SDFFX1 DFF_378_Q_reg ( .D(test_so23), .SI(test_si24), .SE(n8160), .CLK(n8347), .Q(g7956), .QN(n4461) );
  SDFFX1 DFF_379_Q_reg ( .D(g7956), .SI(g7956), .SE(n8160), .CLK(n8347), .Q(
        g485), .QN(n4466) );
  SDFFX1 DFF_380_Q_reg ( .D(g23067), .SI(g485), .SE(n8160), .CLK(n8347), .Q(
        g486) );
  SDFFX1 DFF_381_Q_reg ( .D(g23093), .SI(g486), .SE(n8161), .CLK(n8348), .Q(
        g487) );
  SDFFX1 DFF_382_Q_reg ( .D(g23117), .SI(g487), .SE(n8161), .CLK(n8348), .Q(
        g488) );
  SDFFX1 DFF_383_Q_reg ( .D(g23385), .SI(g488), .SE(n8161), .CLK(n8348), .Q(
        g455) );
  SDFFX1 DFF_384_Q_reg ( .D(g23399), .SI(g455), .SE(n8161), .CLK(n8348), .Q(
        g458) );
  SDFFX1 DFF_385_Q_reg ( .D(g24174), .SI(g458), .SE(n8161), .CLK(n8348), .Q(
        g461) );
  SDFFX1 DFF_386_Q_reg ( .D(g24178), .SI(g461), .SE(n8161), .CLK(n8348), .Q(
        g477) );
  SDFFX1 DFF_387_Q_reg ( .D(g24207), .SI(g477), .SE(n8161), .CLK(n8348), .Q(
        g478) );
  SDFFX1 DFF_388_Q_reg ( .D(g24216), .SI(g478), .SE(n8161), .CLK(n8348), .Q(
        g479) );
  SDFFX1 DFF_389_Q_reg ( .D(g23092), .SI(g479), .SE(n8161), .CLK(n8348), .Q(
        g480) );
  SDFFX1 DFF_390_Q_reg ( .D(g23000), .SI(g480), .SE(n8161), .CLK(n8348), .Q(
        g484) );
  SDFFX1 DFF_391_Q_reg ( .D(g23022), .SI(g484), .SE(n8161), .CLK(n8348), .Q(
        g464) );
  SDFFX1 DFF_392_Q_reg ( .D(g24206), .SI(g464), .SE(n8162), .CLK(n8349), .Q(
        g465) );
  SDFFX1 DFF_393_Q_reg ( .D(g24215), .SI(g465), .SE(n8162), .CLK(n8349), .Q(
        test_so24) );
  SDFFX1 DFF_394_Q_reg ( .D(g24228), .SI(test_si25), .SE(n8161), .CLK(n8348), 
        .Q(g471) );
  SDFFX1 DFF_395_Q_reg ( .D(n499), .SI(g471), .SE(n8162), .CLK(n8349), .Q(g528) );
  SDFFX1 DFF_396_Q_reg ( .D(g528), .SI(g528), .SE(n8162), .CLK(n8349), .Q(g535) );
  SDFFX1 DFF_397_Q_reg ( .D(g535), .SI(g535), .SE(n8162), .CLK(n8349), .Q(g542) );
  SDFFX1 DFF_398_Q_reg ( .D(g13149), .SI(g542), .SE(n8162), .CLK(n8349), .Q(
        g543) );
  SDFFX1 DFF_399_Q_reg ( .D(g543), .SI(g543), .SE(n8162), .CLK(n8349), .Q(g544) );
  SDFFX1 DFF_400_Q_reg ( .D(g21851), .SI(g544), .SE(n8162), .CLK(n8349), .Q(
        g548) );
  SDFFX1 DFF_401_Q_reg ( .D(g13111), .SI(g548), .SE(n8162), .CLK(n8349), .Q(
        g549) );
  SDFFX1 DFF_402_Q_reg ( .D(g549), .SI(g549), .SE(n8162), .CLK(n8349), .Q(g499), .QN(n4541) );
  SDFFX1 DFF_403_Q_reg ( .D(g13160), .SI(g499), .SE(n8162), .CLK(n8349), .Q(
        g558) );
  SDFFX1 DFF_404_Q_reg ( .D(g558), .SI(g558), .SE(n8162), .CLK(n8349), .Q(g559), .QN(n7744) );
  SDFFX1 DFF_405_Q_reg ( .D(g27261), .SI(g559), .SE(n8168), .CLK(n8355), .Q(
        g576), .QN(n7335) );
  SDFFX1 DFF_406_Q_reg ( .D(g27268), .SI(g576), .SE(n8168), .CLK(n8355), .Q(
        g577), .QN(n7337) );
  SDFFX1 DFF_407_Q_reg ( .D(g27279), .SI(g577), .SE(n8168), .CLK(n8355), .Q(
        g575), .QN(n7336) );
  SDFFX1 DFF_408_Q_reg ( .D(g27269), .SI(g575), .SE(n8169), .CLK(n8356), .Q(
        g579), .QN(n7347) );
  SDFFX1 DFF_409_Q_reg ( .D(g27280), .SI(g579), .SE(n8169), .CLK(n8356), .Q(
        test_so25), .QN(n8109) );
  SDFFX1 DFF_410_Q_reg ( .D(g27294), .SI(test_si26), .SE(n8169), .CLK(n8356), 
        .Q(g578), .QN(n7348) );
  SDFFX1 DFF_411_Q_reg ( .D(g27281), .SI(g578), .SE(n8169), .CLK(n8356), .Q(
        g582), .QN(n7172) );
  SDFFX1 DFF_412_Q_reg ( .D(g27295), .SI(g582), .SE(n8169), .CLK(n8356), .Q(
        g583), .QN(n7174) );
  SDFFX1 DFF_413_Q_reg ( .D(g27311), .SI(g583), .SE(n8168), .CLK(n8355), .Q(
        g581), .QN(n7173) );
  SDFFX1 DFF_414_Q_reg ( .D(g27296), .SI(g581), .SE(n8168), .CLK(n8355), .Q(
        g585), .QN(n7357) );
  SDFFX1 DFF_415_Q_reg ( .D(g27312), .SI(g585), .SE(n8169), .CLK(n8356), .Q(
        g586), .QN(n7359) );
  SDFFX1 DFF_416_Q_reg ( .D(g27327), .SI(g586), .SE(n8169), .CLK(n8356), .Q(
        g584), .QN(n7358) );
  SDFFX1 DFF_417_Q_reg ( .D(g24491), .SI(g584), .SE(n8169), .CLK(n8356), .Q(
        g587) );
  SDFFX1 DFF_418_Q_reg ( .D(g24498), .SI(g587), .SE(n8169), .CLK(n8356), .Q(
        g590) );
  SDFFX1 DFF_419_Q_reg ( .D(g24507), .SI(g590), .SE(n8169), .CLK(n8356), .Q(
        g593) );
  SDFFX1 DFF_420_Q_reg ( .D(g24499), .SI(g593), .SE(n8169), .CLK(n8356), .Q(
        g596) );
  SDFFX1 DFF_421_Q_reg ( .D(g24508), .SI(g596), .SE(n8169), .CLK(n8356), .Q(
        g599) );
  SDFFX1 DFF_422_Q_reg ( .D(g24519), .SI(g599), .SE(n8170), .CLK(n8357), .Q(
        g602) );
  SDFFX1 DFF_423_Q_reg ( .D(g28345), .SI(g602), .SE(n8170), .CLK(n8357), .Q(
        g614) );
  SDFFX1 DFF_424_Q_reg ( .D(g28349), .SI(g614), .SE(n8170), .CLK(n8357), .Q(
        g617) );
  SDFFX1 DFF_425_Q_reg ( .D(g28353), .SI(g617), .SE(n8168), .CLK(n8355), .Q(
        test_so26) );
  SDFFX1 DFF_426_Q_reg ( .D(g28342), .SI(test_si27), .SE(n8170), .CLK(n8357), 
        .Q(g605) );
  SDFFX1 DFF_427_Q_reg ( .D(g28344), .SI(g605), .SE(n8170), .CLK(n8357), .Q(
        g608) );
  SDFFX1 DFF_428_Q_reg ( .D(g28348), .SI(g608), .SE(n8170), .CLK(n8357), .Q(
        g611) );
  SDFFX1 DFF_429_Q_reg ( .D(g26541), .SI(g611), .SE(n8170), .CLK(n8357), .Q(
        g490) );
  SDFFX1 DFF_430_Q_reg ( .D(g26545), .SI(g490), .SE(n8170), .CLK(n8357), .Q(
        g493) );
  SDFFX1 DFF_431_Q_reg ( .D(g26553), .SI(g493), .SE(n8168), .CLK(n8355), .Q(
        g496) );
  SDFFX1 DFF_432_Q_reg ( .D(g499), .SI(g496), .SE(n8168), .CLK(n8355), .Q(g506), .QN(n4570) );
  SDFFX1 DFF_433_Q_reg ( .D(g22578), .SI(g506), .SE(n8170), .CLK(n8357), .Q(
        n4571), .QN(n7406) );
  SDFFX1 DFF_442_Q_reg ( .D(n514), .SI(n4571), .SE(n8170), .CLK(n8357), .Q(
        g16297), .QN(n8030) );
  SDFFX1 DFF_443_Q_reg ( .D(g16297), .SI(g16297), .SE(n8170), .CLK(n8357), .Q(
        g525), .QN(n8036) );
  SDFFX1 DFF_444_Q_reg ( .D(DFF_299_n1), .SI(g525), .SE(n8170), .CLK(n8357), 
        .Q(n8047), .QN(DFF_444_n1) );
  SDFFX1 DFF_445_Q_reg ( .D(DFF_301_n1), .SI(n8047), .SE(n8171), .CLK(n8358), 
        .Q(n8046), .QN(DFF_445_n1) );
  SDFFX1 DFF_446_Q_reg ( .D(DFF_303_n1), .SI(n8046), .SE(n8171), .CLK(n8358), 
        .Q(n8045), .QN(DFF_446_n1) );
  SDFFX1 DFF_447_Q_reg ( .D(DFF_305_n1), .SI(n8045), .SE(n8171), .CLK(n8358), 
        .Q(n8044), .QN(DFF_447_n1) );
  SDFFX1 DFF_448_Q_reg ( .D(DFF_307_n1), .SI(n8044), .SE(n8171), .CLK(n8358), 
        .Q(n8043), .QN(DFF_448_n1) );
  SDFFX1 DFF_449_Q_reg ( .D(DFF_309_n1), .SI(n8043), .SE(n8171), .CLK(n8358), 
        .Q(test_so27), .QN(DFF_449_n1) );
  SDFFX1 DFF_450_Q_reg ( .D(DFF_311_n1), .SI(test_si28), .SE(n8145), .CLK(
        n8332), .Q(g536), .QN(n7143) );
  SDFFX1 DFF_451_Q_reg ( .D(DFF_313_n1), .SI(g536), .SE(n8145), .CLK(n8332), 
        .Q(g537), .QN(n7142) );
  SDFFX1 DFF_452_Q_reg ( .D(g24059), .SI(g537), .SE(n8163), .CLK(n8350), .Q(
        g538), .QN(n4492) );
  SDFFX1 DFF_453_Q_reg ( .D(n4485), .SI(g538), .SE(n8163), .CLK(n8350), .Q(
        n8040), .QN(n14345) );
  SDFFX1 DFF_455_Q_reg ( .D(g6677), .SI(g6677), .SE(n8163), .CLK(n8350), .Q(
        g6911), .QN(n4359) );
  SDFFX1 DFF_456_Q_reg ( .D(g6911), .SI(g6911), .SE(n8163), .CLK(n8350), .Q(
        g629), .QN(n4295) );
  SDFFX1 DFF_457_Q_reg ( .D(g16654), .SI(g629), .SE(n8166), .CLK(n8353), .Q(
        g630), .QN(n7748) );
  SDFFX1 DFF_458_Q_reg ( .D(g20314), .SI(g630), .SE(n8166), .CLK(n8353), .Q(
        g659), .QN(n4429) );
  SDFFX1 DFF_459_Q_reg ( .D(g20682), .SI(g659), .SE(n8166), .CLK(n8353), .Q(
        g640), .QN(n4404) );
  SDFFX1 DFF_460_Q_reg ( .D(n596), .SI(g640), .SE(n8166), .CLK(n8353), .Q(g633), .QN(n4478) );
  SDFFX1 DFF_461_Q_reg ( .D(g23324), .SI(g633), .SE(n8166), .CLK(n8353), .Q(
        g653), .QN(n4422) );
  SDFFX1 DFF_462_Q_reg ( .D(g24426), .SI(g653), .SE(n8166), .CLK(n8353), .Q(
        g646), .QN(n4414) );
  SDFFX1 DFF_463_Q_reg ( .D(g25185), .SI(g646), .SE(n8166), .CLK(n8353), .Q(
        g660), .QN(n4403) );
  SDFFX1 DFF_464_Q_reg ( .D(n597), .SI(g660), .SE(n8166), .CLK(n8353), .Q(g672), .QN(n4413) );
  SDFFX1 DFF_465_Q_reg ( .D(g26776), .SI(g672), .SE(n8166), .CLK(n8353), .Q(
        test_so28), .QN(n8074) );
  SDFFX1 DFF_466_Q_reg ( .D(g27672), .SI(test_si29), .SE(n8166), .CLK(n8353), 
        .Q(g679), .QN(n4477) );
  SDFFX1 DFF_467_Q_reg ( .D(g28199), .SI(g679), .SE(n8166), .CLK(n8353), .Q(
        g686), .QN(n4396) );
  SDFFX1 DFF_468_Q_reg ( .D(g28668), .SI(g686), .SE(n8167), .CLK(n8354), .Q(
        g692), .QN(n4418) );
  SDFFX1 DFF_469_Q_reg ( .D(g20875), .SI(g692), .SE(n8171), .CLK(n8358), .Q(
        g699), .QN(n7826) );
  SDFFX1 DFF_470_Q_reg ( .D(g20879), .SI(g699), .SE(n8171), .CLK(n8358), .Q(
        g700), .QN(n7825) );
  SDFFX1 DFF_471_Q_reg ( .D(g20891), .SI(g700), .SE(n8171), .CLK(n8358), .Q(
        g698), .QN(n7864) );
  SDFFX1 DFF_472_Q_reg ( .D(g20880), .SI(g698), .SE(n8171), .CLK(n8358), .Q(
        g702), .QN(n7824) );
  SDFFX1 DFF_473_Q_reg ( .D(g20892), .SI(g702), .SE(n8171), .CLK(n8358), .Q(
        g703), .QN(n7823) );
  SDFFX1 DFF_474_Q_reg ( .D(g20901), .SI(g703), .SE(n8172), .CLK(n8359), .Q(
        g701), .QN(n7863) );
  SDFFX1 DFF_475_Q_reg ( .D(g20893), .SI(g701), .SE(n8172), .CLK(n8359), .Q(
        g705), .QN(n7822) );
  SDFFX1 DFF_476_Q_reg ( .D(g20902), .SI(g705), .SE(n8172), .CLK(n8359), .Q(
        g706), .QN(n7821) );
  SDFFX1 DFF_477_Q_reg ( .D(g20921), .SI(g706), .SE(n8172), .CLK(n8359), .Q(
        g704), .QN(n7862) );
  SDFFX1 DFF_478_Q_reg ( .D(g20903), .SI(g704), .SE(n8172), .CLK(n8359), .Q(
        g708), .QN(n7820) );
  SDFFX1 DFF_479_Q_reg ( .D(g20922), .SI(g708), .SE(n8172), .CLK(n8359), .Q(
        g709), .QN(n7819) );
  SDFFX1 DFF_480_Q_reg ( .D(g20944), .SI(g709), .SE(n8173), .CLK(n8360), .Q(
        g707), .QN(n7861) );
  SDFFX1 DFF_481_Q_reg ( .D(g20923), .SI(g707), .SE(n8173), .CLK(n8360), .Q(
        test_so29), .QN(n8125) );
  SDFFX1 DFF_482_Q_reg ( .D(g20945), .SI(test_si30), .SE(n8171), .CLK(n8358), 
        .Q(g712), .QN(n7818) );
  SDFFX1 DFF_483_Q_reg ( .D(g20966), .SI(g712), .SE(n8173), .CLK(n8360), .Q(
        g710), .QN(n7860) );
  SDFFX1 DFF_484_Q_reg ( .D(g20946), .SI(g710), .SE(n8173), .CLK(n8360), .Q(
        g714), .QN(n7817) );
  SDFFX1 DFF_485_Q_reg ( .D(g20967), .SI(g714), .SE(n8173), .CLK(n8360), .Q(
        g715), .QN(n7816) );
  SDFFX1 DFF_486_Q_reg ( .D(g20989), .SI(g715), .SE(n8173), .CLK(n8360), .Q(
        g713), .QN(n7859) );
  SDFFX1 DFF_487_Q_reg ( .D(g20968), .SI(g713), .SE(n8173), .CLK(n8360), .Q(
        g717), .QN(n7815) );
  SDFFX1 DFF_488_Q_reg ( .D(g20990), .SI(g717), .SE(n8173), .CLK(n8360), .Q(
        g718), .QN(n7814) );
  SDFFX1 DFF_489_Q_reg ( .D(g21009), .SI(g718), .SE(n8173), .CLK(n8360), .Q(
        g716), .QN(n7858) );
  SDFFX1 DFF_490_Q_reg ( .D(g20991), .SI(g716), .SE(n8173), .CLK(n8360), .Q(
        g720), .QN(n7813) );
  SDFFX1 DFF_491_Q_reg ( .D(g21010), .SI(g720), .SE(n8173), .CLK(n8360), .Q(
        g721), .QN(n7812) );
  SDFFX1 DFF_492_Q_reg ( .D(g21031), .SI(g721), .SE(n8173), .CLK(n8360), .Q(
        g719), .QN(n7857) );
  SDFFX1 DFF_493_Q_reg ( .D(g21011), .SI(g719), .SE(n8174), .CLK(n8361), .Q(
        g723), .QN(n7811) );
  SDFFX1 DFF_494_Q_reg ( .D(g21032), .SI(g723), .SE(n8174), .CLK(n8361), .Q(
        g724), .QN(n7810) );
  SDFFX1 DFF_495_Q_reg ( .D(g21051), .SI(g724), .SE(n8174), .CLK(n8361), .Q(
        g722), .QN(n7856) );
  SDFFX1 DFF_496_Q_reg ( .D(g20876), .SI(g722), .SE(n8174), .CLK(n8361), .Q(
        g726), .QN(n7809) );
  SDFFX1 DFF_497_Q_reg ( .D(g20881), .SI(g726), .SE(n8174), .CLK(n8361), .Q(
        test_so30), .QN(n8126) );
  SDFFX1 DFF_498_Q_reg ( .D(g20894), .SI(test_si31), .SE(n8171), .CLK(n8358), 
        .Q(g725), .QN(n7855) );
  SDFFX1 DFF_499_Q_reg ( .D(g20924), .SI(g725), .SE(n8172), .CLK(n8359), .Q(
        g729), .QN(n8022) );
  SDFFX1 DFF_500_Q_reg ( .D(g20947), .SI(g729), .SE(n8172), .CLK(n8359), .Q(
        g730), .QN(n7562) );
  SDFFX1 DFF_501_Q_reg ( .D(g20969), .SI(g730), .SE(n8172), .CLK(n8359), .Q(
        g728) );
  SDFFX1 DFF_502_Q_reg ( .D(g20948), .SI(g728), .SE(n8172), .CLK(n8359), .Q(
        g732), .QN(n7566) );
  SDFFX1 DFF_503_Q_reg ( .D(g20970), .SI(g732), .SE(n8172), .CLK(n8359), .Q(
        g733), .QN(n7561) );
  SDFFX1 DFF_504_Q_reg ( .D(g20992), .SI(g733), .SE(n8172), .CLK(n8359), .Q(
        g731), .QN(n7618) );
  SDFFX1 DFF_505_Q_reg ( .D(g25260), .SI(g731), .SE(n8174), .CLK(n8361), .Q(
        g735), .QN(n7497) );
  SDFFX1 DFF_506_Q_reg ( .D(g25262), .SI(g735), .SE(n8174), .CLK(n8361), .Q(
        g736), .QN(n7496) );
  SDFFX1 DFF_507_Q_reg ( .D(g25266), .SI(g736), .SE(n8174), .CLK(n8361), .Q(
        g734), .QN(n7501) );
  SDFFX1 DFF_508_Q_reg ( .D(g22218), .SI(g734), .SE(n8174), .CLK(n8361), .Q(
        g738), .QN(n7868) );
  SDFFX1 DFF_509_Q_reg ( .D(n567), .SI(g738), .SE(n8174), .CLK(n8361), .Q(g739), .QN(n7956) );
  SDFFX1 DFF_510_Q_reg ( .D(g22242), .SI(g739), .SE(n8174), .CLK(n8361), .Q(
        g737), .QN(n7959) );
  SDFFX1 DFF_511_Q_reg ( .D(g2950), .SI(g737), .SE(n8174), .CLK(n8361), .Q(
        g6368), .QN(n4323) );
  SDFFX1 DFF_512_Q_reg ( .D(g6368), .SI(g6368), .SE(n8175), .CLK(n8362), .Q(
        g6518), .QN(n4312) );
  SDFFX1 DFF_513_Q_reg ( .D(g6518), .SI(g6518), .SE(n8175), .CLK(n8362), .Q(
        test_so31), .QN(n8071) );
  SDFFX1 DFF_514_Q_reg ( .D(g22126), .SI(test_si32), .SE(n8176), .CLK(n8363), 
        .Q(g818), .QN(n7916) );
  SDFFX1 DFF_515_Q_reg ( .D(g22145), .SI(g818), .SE(n8179), .CLK(n8366), .Q(
        g819), .QN(n7915) );
  SDFFX1 DFF_516_Q_reg ( .D(g22162), .SI(g819), .SE(n8179), .CLK(n8366), .Q(
        g817), .QN(n7545) );
  SDFFX1 DFF_517_Q_reg ( .D(g22146), .SI(g817), .SE(n8176), .CLK(n8363), .Q(
        g821), .QN(n7914) );
  SDFFX1 DFF_518_Q_reg ( .D(g22163), .SI(g821), .SE(n8179), .CLK(n8366), .Q(
        g822), .QN(n7911) );
  SDFFX1 DFF_519_Q_reg ( .D(g22177), .SI(g822), .SE(n8180), .CLK(n8367), .Q(
        g820), .QN(n7544) );
  SDFFX1 DFF_520_Q_reg ( .D(g22029), .SI(g820), .SE(n8180), .CLK(n8367), .Q(
        g830), .QN(n7910) );
  SDFFX1 DFF_521_Q_reg ( .D(g22033), .SI(g830), .SE(n8180), .CLK(n8367), .Q(
        g831), .QN(n7908) );
  SDFFX1 DFF_522_Q_reg ( .D(g22040), .SI(g831), .SE(n8180), .CLK(n8367), .Q(
        g829), .QN(n7543) );
  SDFFX1 DFF_523_Q_reg ( .D(g22034), .SI(g829), .SE(n8180), .CLK(n8367), .Q(
        g833), .QN(n7906) );
  SDFFX1 DFF_524_Q_reg ( .D(g22041), .SI(g833), .SE(n8180), .CLK(n8367), .Q(
        g834), .QN(n7905) );
  SDFFX1 DFF_525_Q_reg ( .D(g22054), .SI(g834), .SE(n8180), .CLK(n8367), .Q(
        g832), .QN(n7542) );
  SDFFX1 DFF_526_Q_reg ( .D(g22042), .SI(g832), .SE(n8180), .CLK(n8367), .Q(
        g836), .QN(n7904) );
  SDFFX1 DFF_527_Q_reg ( .D(g22055), .SI(g836), .SE(n8180), .CLK(n8367), .Q(
        g837), .QN(n7903) );
  SDFFX1 DFF_528_Q_reg ( .D(g22066), .SI(g837), .SE(n8180), .CLK(n8367), .Q(
        g835), .QN(n7541) );
  SDFFX1 DFF_529_Q_reg ( .D(g22056), .SI(g835), .SE(n8180), .CLK(n8367), .Q(
        test_so32), .QN(n8113) );
  SDFFX1 DFF_530_Q_reg ( .D(g22067), .SI(test_si33), .SE(n8178), .CLK(n8365), 
        .Q(g840), .QN(n7902) );
  SDFFX1 DFF_531_Q_reg ( .D(g22087), .SI(g840), .SE(n8178), .CLK(n8365), .Q(
        g838), .QN(n7540) );
  SDFFX1 DFF_532_Q_reg ( .D(g22068), .SI(g838), .SE(n8178), .CLK(n8365), .Q(
        g842), .QN(n7901) );
  SDFFX1 DFF_533_Q_reg ( .D(g22088), .SI(g842), .SE(n8178), .CLK(n8365), .Q(
        g843), .QN(n7900) );
  SDFFX1 DFF_534_Q_reg ( .D(g22104), .SI(g843), .SE(n8178), .CLK(n8365), .Q(
        g841), .QN(n7539) );
  SDFFX1 DFF_535_Q_reg ( .D(g22089), .SI(g841), .SE(n8178), .CLK(n8365), .Q(
        g845), .QN(n7899) );
  SDFFX1 DFF_536_Q_reg ( .D(g22105), .SI(g845), .SE(n8178), .CLK(n8365), .Q(
        g846), .QN(n7898) );
  SDFFX1 DFF_537_Q_reg ( .D(g22127), .SI(g846), .SE(n8179), .CLK(n8366), .Q(
        g844), .QN(n7538) );
  SDFFX1 DFF_538_Q_reg ( .D(g22106), .SI(g844), .SE(n8179), .CLK(n8366), .Q(
        g848), .QN(n7537) );
  SDFFX1 DFF_539_Q_reg ( .D(g22128), .SI(g848), .SE(n8179), .CLK(n8366), .Q(
        g849), .QN(n7536) );
  SDFFX1 DFF_540_Q_reg ( .D(g22147), .SI(g849), .SE(n8179), .CLK(n8366), .Q(
        g847), .QN(n7535) );
  SDFFX1 DFF_541_Q_reg ( .D(g22129), .SI(g847), .SE(n8179), .CLK(n8366), .Q(
        g851), .QN(n7534) );
  SDFFX1 DFF_542_Q_reg ( .D(g22148), .SI(g851), .SE(n8179), .CLK(n8366), .Q(
        g852), .QN(n7533) );
  SDFFX1 DFF_543_Q_reg ( .D(g22164), .SI(g852), .SE(n8179), .CLK(n8366), .Q(
        g850), .QN(n7532) );
  SDFFX1 DFF_544_Q_reg ( .D(g25209), .SI(g850), .SE(n8179), .CLK(n8366), .Q(
        g857), .QN(n7600) );
  SDFFX1 DFF_545_Q_reg ( .D(g25214), .SI(g857), .SE(n8179), .CLK(n8366), .Q(
        test_so33), .QN(n8105) );
  SDFFX1 DFF_546_Q_reg ( .D(g25221), .SI(test_si34), .SE(n8175), .CLK(n8362), 
        .Q(g856), .QN(n7599) );
  SDFFX1 DFF_547_Q_reg ( .D(g25215), .SI(g856), .SE(n8175), .CLK(n8362), .Q(
        g860), .QN(n7598) );
  SDFFX1 DFF_548_Q_reg ( .D(g25222), .SI(g860), .SE(n8175), .CLK(n8362), .Q(
        g861), .QN(n7597) );
  SDFFX1 DFF_549_Q_reg ( .D(g25230), .SI(g861), .SE(n8175), .CLK(n8362), .Q(
        g859), .QN(n7596) );
  SDFFX1 DFF_550_Q_reg ( .D(g25223), .SI(g859), .SE(n8175), .CLK(n8362), .Q(
        g863), .QN(n7595) );
  SDFFX1 DFF_551_Q_reg ( .D(g25231), .SI(g863), .SE(n8175), .CLK(n8362), .Q(
        g864), .QN(n7594) );
  SDFFX1 DFF_552_Q_reg ( .D(g25240), .SI(g864), .SE(n8175), .CLK(n8362), .Q(
        g862), .QN(n7593) );
  SDFFX1 DFF_553_Q_reg ( .D(g25232), .SI(g862), .SE(n8175), .CLK(n8362), .Q(
        g866), .QN(n7592) );
  SDFFX1 DFF_554_Q_reg ( .D(g25241), .SI(g866), .SE(n8175), .CLK(n8362), .Q(
        g867), .QN(n7591) );
  SDFFX1 DFF_555_Q_reg ( .D(g25248), .SI(g867), .SE(n8175), .CLK(n8362), .Q(
        g865), .QN(n7590) );
  SDFFX1 DFF_556_Q_reg ( .D(g30269), .SI(g865), .SE(n8186), .CLK(n8373), .Q(
        g873) );
  SDFFX1 DFF_557_Q_reg ( .D(g30277), .SI(g873), .SE(n8186), .CLK(n8373), .Q(
        g876) );
  SDFFX1 DFF_558_Q_reg ( .D(g30285), .SI(g876), .SE(n8186), .CLK(n8373), .Q(
        g879) );
  SDFFX1 DFF_559_Q_reg ( .D(g30643), .SI(g879), .SE(n8186), .CLK(n8373), .Q(
        g918) );
  SDFFX1 DFF_560_Q_reg ( .D(g30648), .SI(g918), .SE(n8187), .CLK(n8374), .Q(
        g921) );
  SDFFX1 DFF_561_Q_reg ( .D(g30654), .SI(g921), .SE(n8182), .CLK(n8369), .Q(
        test_so34) );
  SDFFX1 DFF_562_Q_reg ( .D(g30676), .SI(test_si35), .SE(n8176), .CLK(n8363), 
        .Q(g882) );
  SDFFX1 DFF_563_Q_reg ( .D(g30681), .SI(g882), .SE(n8176), .CLK(n8363), .Q(
        g885) );
  SDFFX1 DFF_564_Q_reg ( .D(g30687), .SI(g885), .SE(n8176), .CLK(n8363), .Q(
        g888) );
  SDFFX1 DFF_565_Q_reg ( .D(g30649), .SI(g888), .SE(n8180), .CLK(n8367), .Q(
        g927) );
  SDFFX1 DFF_566_Q_reg ( .D(g30655), .SI(g927), .SE(n8181), .CLK(n8368), .Q(
        g930) );
  SDFFX1 DFF_567_Q_reg ( .D(g30662), .SI(g930), .SE(n8181), .CLK(n8368), .Q(
        g933) );
  SDFFX1 DFF_568_Q_reg ( .D(g30286), .SI(g933), .SE(n8181), .CLK(n8368), .Q(
        g891) );
  SDFFX1 DFF_569_Q_reg ( .D(g30293), .SI(g891), .SE(n8181), .CLK(n8368), .Q(
        g894) );
  SDFFX1 DFF_570_Q_reg ( .D(g30298), .SI(g894), .SE(n8181), .CLK(n8368), .Q(
        g897) );
  SDFFX1 DFF_571_Q_reg ( .D(g30259), .SI(g897), .SE(n8181), .CLK(n8368), .Q(
        g936) );
  SDFFX1 DFF_572_Q_reg ( .D(g30264), .SI(g936), .SE(n8181), .CLK(n8368), .Q(
        g939) );
  SDFFX1 DFF_573_Q_reg ( .D(g30270), .SI(g939), .SE(n8181), .CLK(n8368), .Q(
        g942) );
  SDFFX1 DFF_574_Q_reg ( .D(g30247), .SI(g942), .SE(n8181), .CLK(n8368), .Q(
        g900) );
  SDFFX1 DFF_575_Q_reg ( .D(g30249), .SI(g900), .SE(n8182), .CLK(n8369), .Q(
        g903) );
  SDFFX1 DFF_576_Q_reg ( .D(g30251), .SI(g903), .SE(n8182), .CLK(n8369), .Q(
        g906) );
  SDFFX1 DFF_577_Q_reg ( .D(g30265), .SI(g906), .SE(n8182), .CLK(n8369), .Q(
        test_so35) );
  SDFFX1 DFF_578_Q_reg ( .D(g30271), .SI(test_si36), .SE(n8182), .CLK(n8369), 
        .Q(g948) );
  SDFFX1 DFF_579_Q_reg ( .D(g30278), .SI(g948), .SE(n8182), .CLK(n8369), .Q(
        g951) );
  SDFFX1 DFF_580_Q_reg ( .D(g30638), .SI(g951), .SE(n8182), .CLK(n8369), .Q(
        g909) );
  SDFFX1 DFF_581_Q_reg ( .D(g30642), .SI(g909), .SE(n8182), .CLK(n8369), .Q(
        g912) );
  SDFFX1 DFF_582_Q_reg ( .D(g30647), .SI(g912), .SE(n8181), .CLK(n8368), .Q(
        g915) );
  SDFFX1 DFF_583_Q_reg ( .D(g30670), .SI(g915), .SE(n8181), .CLK(n8368), .Q(
        g954) );
  SDFFX1 DFF_584_Q_reg ( .D(g30677), .SI(g954), .SE(n8181), .CLK(n8368), .Q(
        g957) );
  SDFFX1 DFF_585_Q_reg ( .D(g30682), .SI(g957), .SE(n8176), .CLK(n8363), .Q(
        g960) );
  SDFFX1 DFF_586_Q_reg ( .D(g25042), .SI(g960), .SE(n8176), .CLK(n8363), .Q(
        g780), .QN(n7698) );
  SDFFX1 DFF_587_Q_reg ( .D(g25935), .SI(g780), .SE(n8176), .CLK(n8363), .Q(
        g776), .QN(n8054) );
  SDFFX1 DFF_588_Q_reg ( .D(g26530), .SI(g776), .SE(n8176), .CLK(n8363), .Q(
        g771), .QN(n7697) );
  SDFFX1 DFF_589_Q_reg ( .D(g27123), .SI(g771), .SE(n8176), .CLK(n8363), .Q(
        g767), .QN(n8063) );
  SDFFX1 DFF_590_Q_reg ( .D(g27603), .SI(g767), .SE(n8177), .CLK(n8364), .Q(
        g762), .QN(n7696) );
  SDFFX1 DFF_591_Q_reg ( .D(g28146), .SI(g762), .SE(n8177), .CLK(n8364), .Q(
        g758), .QN(n8064) );
  SDFFX1 DFF_592_Q_reg ( .D(g28635), .SI(g758), .SE(n8177), .CLK(n8364), .Q(
        g753), .QN(n7695) );
  SDFFX1 DFF_593_Q_reg ( .D(g29110), .SI(g753), .SE(n8177), .CLK(n8364), .Q(
        test_so36) );
  SDFFX1 DFF_594_Q_reg ( .D(g29354), .SI(test_si37), .SE(n8177), .CLK(n8364), 
        .Q(g744), .QN(n7324) );
  SDFFX1 DFF_595_Q_reg ( .D(g29580), .SI(g744), .SE(n8177), .CLK(n8364), .Q(
        g740), .QN(n7163) );
  SDFFX1 DFF_596_Q_reg ( .D(n19), .SI(g740), .SE(n8177), .CLK(n8364), .Q(g868)
         );
  SDFFX1 DFF_597_Q_reg ( .D(g868), .SI(g868), .SE(n8177), .CLK(n8364), .Q(
        g5595) );
  SDFFX1 DFF_598_Q_reg ( .D(g5595), .SI(g5595), .SE(n8177), .CLK(n8364), .Q(
        g869), .QN(n7708) );
  SDFFX1 DFF_599_Q_reg ( .D(g2950), .SI(g869), .SE(n8177), .CLK(n8364), .Q(
        g5472), .QN(n4363) );
  SDFFX1 DFF_600_Q_reg ( .D(g5472), .SI(g5472), .SE(n8177), .CLK(n8364), .Q(
        g6712), .QN(n4364) );
  SDFFX1 DFF_601_Q_reg ( .D(g6712), .SI(g6712), .SE(n8177), .CLK(n8364), .Q(
        g1088), .QN(n4381) );
  SDFFX1 DFF_602_Q_reg ( .D(g5595), .SI(g1088), .SE(n8178), .CLK(n8365), .Q(
        g996), .QN(n4387) );
  SDFFX1 DFF_603_Q_reg ( .D(g27257), .SI(g996), .SE(n8185), .CLK(n8372), .Q(
        g1041), .QN(n7651) );
  SDFFX1 DFF_604_Q_reg ( .D(g27262), .SI(g1041), .SE(n8185), .CLK(n8372), .Q(
        g1030), .QN(n7650) );
  SDFFX1 DFF_605_Q_reg ( .D(g27270), .SI(g1030), .SE(n8185), .CLK(n8372), .Q(
        g1033), .QN(n7649) );
  SDFFX1 DFF_606_Q_reg ( .D(g27263), .SI(g1033), .SE(n8186), .CLK(n8373), .Q(
        g1056), .QN(n7628) );
  SDFFX1 DFF_607_Q_reg ( .D(g27271), .SI(g1056), .SE(n8186), .CLK(n8373), .Q(
        g1045), .QN(n7627) );
  SDFFX1 DFF_608_Q_reg ( .D(g27282), .SI(g1045), .SE(n8186), .CLK(n8373), .Q(
        g1048), .QN(n7626) );
  SDFFX1 DFF_609_Q_reg ( .D(g27272), .SI(g1048), .SE(n8186), .CLK(n8373), .Q(
        test_so37), .QN(n8097) );
  SDFFX1 DFF_610_Q_reg ( .D(g27283), .SI(test_si38), .SE(n8186), .CLK(n8373), 
        .Q(g1060), .QN(n7377) );
  SDFFX1 DFF_611_Q_reg ( .D(g27297), .SI(g1060), .SE(n8186), .CLK(n8373), .Q(
        g1063), .QN(n7378) );
  SDFFX1 DFF_612_Q_reg ( .D(g27284), .SI(g1063), .SE(n8186), .CLK(n8373), .Q(
        g1085), .QN(n7639) );
  SDFFX1 DFF_613_Q_reg ( .D(g27298), .SI(g1085), .SE(n8186), .CLK(n8373), .Q(
        g1075), .QN(n7638) );
  SDFFX1 DFF_614_Q_reg ( .D(g27313), .SI(g1075), .SE(n8183), .CLK(n8370), .Q(
        g1078), .QN(n7637) );
  SDFFX1 DFF_615_Q_reg ( .D(g28738), .SI(g1078), .SE(n8184), .CLK(n8371), .Q(
        g1095) );
  SDFFX1 DFF_616_Q_reg ( .D(g28746), .SI(g1095), .SE(n8185), .CLK(n8372), .Q(
        g1098) );
  SDFFX1 DFF_617_Q_reg ( .D(g28758), .SI(g1098), .SE(n8185), .CLK(n8372), .Q(
        g1101) );
  SDFFX1 DFF_618_Q_reg ( .D(g29198), .SI(g1101), .SE(n8185), .CLK(n8372), .Q(
        g1104) );
  SDFFX1 DFF_619_Q_reg ( .D(g29204), .SI(g1104), .SE(n8185), .CLK(n8372), .Q(
        g1107) );
  SDFFX1 DFF_620_Q_reg ( .D(g29209), .SI(g1107), .SE(n8184), .CLK(n8371), .Q(
        g1110) );
  SDFFX1 DFF_621_Q_reg ( .D(g28747), .SI(g1110), .SE(n8184), .CLK(n8371), .Q(
        g1114), .QN(n7677) );
  SDFFX1 DFF_622_Q_reg ( .D(g28759), .SI(g1114), .SE(n8184), .CLK(n8371), .Q(
        g1115), .QN(n7662) );
  SDFFX1 DFF_623_Q_reg ( .D(g28767), .SI(g1115), .SE(n8184), .CLK(n8371), .Q(
        g1113), .QN(n7676) );
  SDFFX1 DFF_624_Q_reg ( .D(g26806), .SI(g1113), .SE(n8184), .CLK(n8371), .Q(
        g1116) );
  SDFFX1 DFF_625_Q_reg ( .D(g26809), .SI(g1116), .SE(n8184), .CLK(n8371), .Q(
        test_so38) );
  SDFFX1 DFF_626_Q_reg ( .D(g26813), .SI(test_si39), .SE(n8184), .CLK(n8371), 
        .Q(g1122) );
  SDFFX1 DFF_627_Q_reg ( .D(g26810), .SI(g1122), .SE(n8184), .CLK(n8371), .Q(
        g1125) );
  SDFFX1 DFF_628_Q_reg ( .D(g26814), .SI(g1125), .SE(n8185), .CLK(n8372), .Q(
        g1128) );
  SDFFX1 DFF_629_Q_reg ( .D(g26818), .SI(g1128), .SE(n8185), .CLK(n8372), .Q(
        g1131) );
  SDFFX1 DFF_630_Q_reg ( .D(g27761), .SI(g1131), .SE(n8185), .CLK(n8372), .Q(
        g1135), .QN(n7675) );
  SDFFX1 DFF_631_Q_reg ( .D(g27763), .SI(g1135), .SE(n8185), .CLK(n8372), .Q(
        g1136), .QN(n7661) );
  SDFFX1 DFF_632_Q_reg ( .D(g27765), .SI(g1136), .SE(n8184), .CLK(n8371), .Q(
        g1134), .QN(n7674) );
  SDFFX1 DFF_633_Q_reg ( .D(g29609), .SI(g1134), .SE(n8184), .CLK(n8371), .Q(
        g999), .QN(n7281) );
  SDFFX1 DFF_634_Q_reg ( .D(g29612), .SI(g999), .SE(n8184), .CLK(n8371), .Q(
        g1000), .QN(n7264) );
  SDFFX1 DFF_635_Q_reg ( .D(g29616), .SI(g1000), .SE(n8183), .CLK(n8370), .Q(
        g1001), .QN(n7280) );
  SDFFX1 DFF_636_Q_reg ( .D(g30701), .SI(g1001), .SE(n8176), .CLK(n8363), .Q(
        g1002), .QN(n7279) );
  SDFFX1 DFF_637_Q_reg ( .D(g30703), .SI(g1002), .SE(n8178), .CLK(n8365), .Q(
        g1003), .QN(n7263) );
  SDFFX1 DFF_638_Q_reg ( .D(g30705), .SI(g1003), .SE(n8178), .CLK(n8365), .Q(
        g1004), .QN(n7278) );
  SDFFX1 DFF_639_Q_reg ( .D(g30470), .SI(g1004), .SE(n8176), .CLK(n8363), .Q(
        g1005), .QN(n7277) );
  SDFFX1 DFF_640_Q_reg ( .D(g30485), .SI(g1005), .SE(n8178), .CLK(n8365), .Q(
        g1006), .QN(n7262) );
  SDFFX1 DFF_641_Q_reg ( .D(g30500), .SI(g1006), .SE(n8178), .CLK(n8365), .Q(
        test_so39), .QN(n8127) );
  SDFFX1 DFF_642_Q_reg ( .D(g29170), .SI(test_si40), .SE(n8187), .CLK(n8374), 
        .Q(g1009), .QN(n7318) );
  SDFFX1 DFF_643_Q_reg ( .D(g29173), .SI(g1009), .SE(n8187), .CLK(n8374), .Q(
        g1010), .QN(n7312) );
  SDFFX1 DFF_644_Q_reg ( .D(g29179), .SI(g1010), .SE(n8182), .CLK(n8369), .Q(
        g1008), .QN(n7317) );
  SDFFX1 DFF_645_Q_reg ( .D(g26661), .SI(g1008), .SE(n8182), .CLK(n8369), .Q(
        g1090), .QN(n7673) );
  SDFFX1 DFF_646_Q_reg ( .D(g26665), .SI(g1090), .SE(n8182), .CLK(n8369), .Q(
        g1091), .QN(n7660) );
  SDFFX1 DFF_647_Q_reg ( .D(g26669), .SI(g1091), .SE(n8182), .CLK(n8369), .Q(
        g1089), .QN(n7672) );
  SDFFX1 DFF_648_Q_reg ( .D(n4289), .SI(g1089), .SE(n8183), .CLK(n8370), .Q(
        g1137) );
  SDFFX1 DFF_649_Q_reg ( .D(g1137), .SI(g1137), .SE(n8183), .CLK(n8370), .Q(
        n8027), .QN(DFF_649_n1) );
  SDFFX1 DFF_650_Q_reg ( .D(n4567), .SI(n8027), .SE(n8183), .CLK(n8370), .Q(
        g1139) );
  SDFFX1 DFF_651_Q_reg ( .D(g1139), .SI(g1139), .SE(n8183), .CLK(n8370), .Q(
        n8026), .QN(DFF_651_n1) );
  SDFFX1 DFF_652_Q_reg ( .D(n4559), .SI(n8026), .SE(n8183), .CLK(n8370), .Q(
        g1141) );
  SDFFX1 DFF_653_Q_reg ( .D(g1141), .SI(g1141), .SE(n8183), .CLK(n8370), .Q(
        n8025), .QN(DFF_653_n1) );
  SDFFX1 DFF_654_Q_reg ( .D(n4327), .SI(n8025), .SE(n8183), .CLK(n8370), .Q(
        g967) );
  SDFFX1 DFF_655_Q_reg ( .D(g967), .SI(g967), .SE(n8183), .CLK(n8370), .Q(
        n8024), .QN(DFF_655_n1) );
  SDFFX1 DFF_656_Q_reg ( .D(n4391), .SI(n8024), .SE(n8183), .CLK(n8370), .Q(
        g969) );
  SDFFX1 DFF_657_Q_reg ( .D(g969), .SI(g969), .SE(n8183), .CLK(n8370), .Q(
        test_so40), .QN(DFF_657_n1) );
  SDFFX1 DFF_658_Q_reg ( .D(n4321), .SI(test_si41), .SE(n8140), .CLK(n8327), 
        .Q(g971) );
  SDFFX1 DFF_659_Q_reg ( .D(g971), .SI(g971), .SE(n8140), .CLK(n8327), .Q(
        n8021), .QN(DFF_659_n1) );
  SDFFX1 DFF_660_Q_reg ( .D(n4375), .SI(n8021), .SE(n8140), .CLK(n8327), .Q(
        g973) );
  SDFFX1 DFF_661_Q_reg ( .D(g973), .SI(g973), .SE(n8140), .CLK(n8327), .Q(
        n8020), .QN(DFF_661_n1) );
  SDFFX1 DFF_662_Q_reg ( .D(n4379), .SI(n8020), .SE(n8140), .CLK(n8327), .Q(
        g975) );
  SDFFX1 DFF_663_Q_reg ( .D(g975), .SI(g975), .SE(n8140), .CLK(n8327), .Q(
        n8019), .QN(DFF_663_n1) );
  SDFFX1 DFF_664_Q_reg ( .D(g2873), .SI(n8019), .SE(n8140), .CLK(n8327), .Q(
        g977) );
  SDFFX1 DFF_665_Q_reg ( .D(g977), .SI(g977), .SE(n8140), .CLK(n8327), .Q(
        n8018), .QN(n4486) );
  SDFFX1 DFF_666_Q_reg ( .D(n4283), .SI(n8018), .SE(n8185), .CLK(n8372), .Q(
        g986), .QN(n4432) );
  SDFFX1 DFF_667_Q_reg ( .D(n438), .SI(g986), .SE(n8187), .CLK(n8374), .Q(g992), .QN(n7705) );
  SDFFX1 DFF_678_Q_reg ( .D(n4277), .SI(g992), .SE(n8187), .CLK(n8374), .Q(
        n8017) );
  SDFFX1 DFF_679_Q_reg ( .D(g1041), .SI(n8017), .SE(n8187), .CLK(n8374), .Q(
        g1029) );
  SDFFX1 DFF_680_Q_reg ( .D(g1029), .SI(g1029), .SE(n8187), .CLK(n8374), .Q(
        g1036) );
  SDFFX1 DFF_681_Q_reg ( .D(g1030), .SI(g1036), .SE(n8187), .CLK(n8374), .Q(
        g1037) );
  SDFFX1 DFF_682_Q_reg ( .D(g1037), .SI(g1037), .SE(n8187), .CLK(n8374), .Q(
        g1038) );
  SDFFX1 DFF_683_Q_reg ( .D(g1033), .SI(g1038), .SE(n8187), .CLK(n8374), .Q(
        test_so41) );
  SDFFX1 DFF_684_Q_reg ( .D(test_so41), .SI(test_si42), .SE(n8187), .CLK(n8374), .Q(g1040) );
  SDFFX1 DFF_685_Q_reg ( .D(g1056), .SI(g1040), .SE(n8187), .CLK(n8374), .Q(
        g1044) );
  SDFFX1 DFF_686_Q_reg ( .D(g1044), .SI(g1044), .SE(n8188), .CLK(n8375), .Q(
        g1051) );
  SDFFX1 DFF_687_Q_reg ( .D(g1045), .SI(g1051), .SE(n8188), .CLK(n8375), .Q(
        g1052) );
  SDFFX1 DFF_688_Q_reg ( .D(g1052), .SI(g1052), .SE(n8188), .CLK(n8375), .Q(
        g1053) );
  SDFFX1 DFF_689_Q_reg ( .D(g1048), .SI(g1053), .SE(n8188), .CLK(n8375), .Q(
        g1054) );
  SDFFX1 DFF_690_Q_reg ( .D(g1054), .SI(g1054), .SE(n8188), .CLK(n8375), .Q(
        g1055) );
  SDFFX1 DFF_691_Q_reg ( .D(test_so37), .SI(g1055), .SE(n8188), .CLK(n8375), 
        .Q(g1059) );
  SDFFX1 DFF_692_Q_reg ( .D(g1059), .SI(g1059), .SE(n8188), .CLK(n8375), .Q(
        g1066) );
  SDFFX1 DFF_693_Q_reg ( .D(g1060), .SI(g1066), .SE(n8188), .CLK(n8375), .Q(
        g1067) );
  SDFFX1 DFF_694_Q_reg ( .D(g1067), .SI(g1067), .SE(n8188), .CLK(n8375), .Q(
        g1068) );
  SDFFX1 DFF_695_Q_reg ( .D(g1063), .SI(g1068), .SE(n8188), .CLK(n8375), .Q(
        g1069) );
  SDFFX1 DFF_696_Q_reg ( .D(g1069), .SI(g1069), .SE(n8188), .CLK(n8375), .Q(
        g1070) );
  SDFFX1 DFF_697_Q_reg ( .D(g1085), .SI(g1070), .SE(n8188), .CLK(n8375), .Q(
        g1074) );
  SDFFX1 DFF_698_Q_reg ( .D(g1074), .SI(g1074), .SE(n8189), .CLK(n8376), .Q(
        g1081) );
  SDFFX1 DFF_699_Q_reg ( .D(g1075), .SI(g1081), .SE(n8189), .CLK(n8376), .Q(
        test_so42) );
  SDFFX1 DFF_700_Q_reg ( .D(test_so42), .SI(test_si43), .SE(n8189), .CLK(n8376), .Q(g1083) );
  SDFFX1 DFF_701_Q_reg ( .D(g1078), .SI(g1083), .SE(n8189), .CLK(n8376), .Q(
        g1084) );
  SDFFX1 DFF_702_Q_reg ( .D(g1084), .SI(g1084), .SE(n8189), .CLK(n8376), .Q(
        g1011) );
  SDFFX1 DFF_703_Q_reg ( .D(n4598), .SI(g1011), .SE(n8189), .CLK(n8376), .Q(
        g5657) );
  SDFFX1 DFF_704_Q_reg ( .D(g5657), .SI(g5657), .SE(n8189), .CLK(n8376), .Q(
        g5686) );
  SDFFX1 DFF_705_Q_reg ( .D(g5686), .SI(g5686), .SE(n8189), .CLK(n8376), .Q(
        g1024) );
  SDFFX1 DFF_706_Q_reg ( .D(n4598), .SI(g1024), .SE(n8189), .CLK(n8376), .Q(
        g6750), .QN(n4371) );
  SDFFX1 DFF_707_Q_reg ( .D(g6750), .SI(g6750), .SE(n8189), .CLK(n8376), .Q(
        g6944), .QN(n4316) );
  SDFFX1 DFF_708_Q_reg ( .D(g6944), .SI(g6944), .SE(n8189), .CLK(n8376), .Q(
        g1236), .QN(n4300) );
  SDFFX1 DFF_709_Q_reg ( .D(n826), .SI(g1236), .SE(n8189), .CLK(n8376), .Q(
        g1240), .QN(n7970) );
  SDFFX1 DFF_710_Q_reg ( .D(g18707), .SI(g1240), .SE(n8190), .CLK(n8377), .Q(
        g1243), .QN(n4353) );
  SDFFX1 DFF_711_Q_reg ( .D(g18763), .SI(g1243), .SE(n8190), .CLK(n8377), .Q(
        g1196), .QN(n4304) );
  SDFFX1 DFF_712_Q_reg ( .D(n808), .SI(g1196), .SE(n8191), .CLK(n8378), .Q(
        g1199) );
  SDFFX1 DFF_713_Q_reg ( .D(g1199), .SI(g1199), .SE(n8191), .CLK(n8378), .Q(
        g1209) );
  SDFFX1 DFF_714_Q_reg ( .D(g1209), .SI(g1209), .SE(n8191), .CLK(n8378), .Q(
        g1210) );
  SDFFX1 DFF_715_Q_reg ( .D(g1142), .SI(g1210), .SE(n8191), .CLK(n8378), .Q(
        test_so43) );
  SDFFX1 DFF_716_Q_reg ( .D(test_so43), .SI(test_si44), .SE(n8191), .CLK(n8378), .Q(g1255) );
  SDFFX1 DFF_717_Q_reg ( .D(g1145), .SI(g1255), .SE(n8191), .CLK(n8378), .Q(
        g1256) );
  SDFFX1 DFF_718_Q_reg ( .D(g1256), .SI(g1256), .SE(n8191), .CLK(n8378), .Q(
        g1257) );
  SDFFX1 DFF_719_Q_reg ( .D(g1148), .SI(g1257), .SE(n8191), .CLK(n8378), .Q(
        g1258) );
  SDFFX1 DFF_720_Q_reg ( .D(g1258), .SI(g1258), .SE(n8191), .CLK(n8378), .Q(
        g1259) );
  SDFFX1 DFF_721_Q_reg ( .D(g1152), .SI(g1259), .SE(n8191), .CLK(n8378), .Q(
        g1260) );
  SDFFX1 DFF_722_Q_reg ( .D(g1260), .SI(g1260), .SE(n8192), .CLK(n8379), .Q(
        g1251) );
  SDFFX1 DFF_723_Q_reg ( .D(g1155), .SI(g1251), .SE(n8192), .CLK(n8379), .Q(
        g1252) );
  SDFFX1 DFF_724_Q_reg ( .D(g1252), .SI(g1252), .SE(n8192), .CLK(n8379), .Q(
        g1253) );
  SDFFX1 DFF_725_Q_reg ( .D(g1158), .SI(g1253), .SE(n8192), .CLK(n8379), .Q(
        g1254) );
  SDFFX1 DFF_726_Q_reg ( .D(g1254), .SI(g1254), .SE(n8192), .CLK(n8379), .Q(
        g1176) );
  SDFFX1 DFF_727_Q_reg ( .D(g2950), .SI(g1176), .SE(n8192), .CLK(n8379), .Q(
        g7961), .QN(n4460) );
  SDFFX1 DFF_728_Q_reg ( .D(g7961), .SI(g7961), .SE(n8192), .CLK(n8379), .Q(
        g8007), .QN(n4459) );
  SDFFX1 DFF_729_Q_reg ( .D(g8007), .SI(g8007), .SE(n8192), .CLK(n8379), .Q(
        g1172), .QN(n4465) );
  SDFFX1 DFF_730_Q_reg ( .D(g23081), .SI(g1172), .SE(n8192), .CLK(n8379), .Q(
        g1173) );
  SDFFX1 DFF_731_Q_reg ( .D(g23111), .SI(g1173), .SE(n8192), .CLK(n8379), .Q(
        test_so44) );
  SDFFX1 DFF_732_Q_reg ( .D(g23126), .SI(test_si45), .SE(n8192), .CLK(n8379), 
        .Q(g1175) );
  SDFFX1 DFF_733_Q_reg ( .D(g23392), .SI(g1175), .SE(n8192), .CLK(n8379), .Q(
        g1142) );
  SDFFX1 DFF_734_Q_reg ( .D(g23406), .SI(g1142), .SE(n8193), .CLK(n8380), .Q(
        g1145) );
  SDFFX1 DFF_735_Q_reg ( .D(g24179), .SI(g1145), .SE(n8193), .CLK(n8380), .Q(
        g1148) );
  SDFFX1 DFF_736_Q_reg ( .D(g24181), .SI(g1148), .SE(n8193), .CLK(n8380), .Q(
        g1164) );
  SDFFX1 DFF_737_Q_reg ( .D(g24213), .SI(g1164), .SE(n8193), .CLK(n8380), .Q(
        g1165) );
  SDFFX1 DFF_738_Q_reg ( .D(g24223), .SI(g1165), .SE(n8193), .CLK(n8380), .Q(
        g1166) );
  SDFFX1 DFF_739_Q_reg ( .D(g23110), .SI(g1166), .SE(n8193), .CLK(n8380), .Q(
        g1167) );
  SDFFX1 DFF_740_Q_reg ( .D(g23014), .SI(g1167), .SE(n8193), .CLK(n8380), .Q(
        g1171) );
  SDFFX1 DFF_741_Q_reg ( .D(g23039), .SI(g1171), .SE(n8193), .CLK(n8380), .Q(
        g1151) );
  SDFFX1 DFF_742_Q_reg ( .D(g24212), .SI(g1151), .SE(n8193), .CLK(n8380), .Q(
        g1152) );
  SDFFX1 DFF_743_Q_reg ( .D(g24222), .SI(g1152), .SE(n8193), .CLK(n8380), .Q(
        g1155) );
  SDFFX1 DFF_744_Q_reg ( .D(g24235), .SI(g1155), .SE(n8193), .CLK(n8380), .Q(
        g1158) );
  SDFFX1 DFF_745_Q_reg ( .D(n822), .SI(g1158), .SE(n8193), .CLK(n8380), .Q(
        g1214) );
  SDFFX1 DFF_746_Q_reg ( .D(g1214), .SI(g1214), .SE(n8194), .CLK(n8381), .Q(
        g1221) );
  SDFFX1 DFF_747_Q_reg ( .D(g1221), .SI(g1221), .SE(n8194), .CLK(n8381), .Q(
        test_so45) );
  SDFFX1 DFF_748_Q_reg ( .D(g13155), .SI(test_si46), .SE(n8194), .CLK(n8381), 
        .Q(g1229) );
  SDFFX1 DFF_749_Q_reg ( .D(g1229), .SI(g1229), .SE(n8194), .CLK(n8381), .Q(
        n4549), .QN(n7141) );
  SDFFX1 DFF_750_Q_reg ( .D(n498), .SI(n4549), .SE(n8194), .CLK(n8381), .Q(
        n4361) );
  SDFFX1 DFF_751_Q_reg ( .D(g13124), .SI(n4361), .SE(n8194), .CLK(n8381), .Q(
        g1235) );
  SDFFX1 DFF_752_Q_reg ( .D(g1235), .SI(g1235), .SE(n8194), .CLK(n8381), .Q(
        g1186), .QN(n4548) );
  SDFFX1 DFF_753_Q_reg ( .D(g13171), .SI(g1186), .SE(n8194), .CLK(n8381), .Q(
        g1244) );
  SDFFX1 DFF_754_Q_reg ( .D(g1244), .SI(g1244), .SE(n8194), .CLK(n8381), .Q(
        g1245), .QN(n7751) );
  SDFFX1 DFF_755_Q_reg ( .D(g27273), .SI(g1245), .SE(n8195), .CLK(n8382), .Q(
        g1262), .QN(n7332) );
  SDFFX1 DFF_756_Q_reg ( .D(g27285), .SI(g1262), .SE(n8196), .CLK(n8383), .Q(
        g1263), .QN(n7334) );
  SDFFX1 DFF_757_Q_reg ( .D(g27299), .SI(g1263), .SE(n8196), .CLK(n8383), .Q(
        g1261), .QN(n7333) );
  SDFFX1 DFF_758_Q_reg ( .D(g27286), .SI(g1261), .SE(n8196), .CLK(n8383), .Q(
        g1265), .QN(n7344) );
  SDFFX1 DFF_759_Q_reg ( .D(g27300), .SI(g1265), .SE(n8196), .CLK(n8383), .Q(
        g1266), .QN(n7346) );
  SDFFX1 DFF_760_Q_reg ( .D(g27314), .SI(g1266), .SE(n8196), .CLK(n8383), .Q(
        g1264), .QN(n7345) );
  SDFFX1 DFF_761_Q_reg ( .D(g27301), .SI(g1264), .SE(n8196), .CLK(n8383), .Q(
        g1268), .QN(n7170) );
  SDFFX1 DFF_762_Q_reg ( .D(g27315), .SI(g1268), .SE(n8196), .CLK(n8383), .Q(
        g1269), .QN(n7171) );
  SDFFX1 DFF_763_Q_reg ( .D(g27328), .SI(g1269), .SE(n8196), .CLK(n8383), .Q(
        test_so46), .QN(n8108) );
  SDFFX1 DFF_764_Q_reg ( .D(g27316), .SI(test_si47), .SE(n8195), .CLK(n8382), 
        .Q(g1271), .QN(n7354) );
  SDFFX1 DFF_765_Q_reg ( .D(g27329), .SI(g1271), .SE(n8196), .CLK(n8383), .Q(
        g1272), .QN(n7356) );
  SDFFX1 DFF_766_Q_reg ( .D(g27339), .SI(g1272), .SE(n8196), .CLK(n8383), .Q(
        g1270), .QN(n7355) );
  SDFFX1 DFF_767_Q_reg ( .D(g24501), .SI(g1270), .SE(n8196), .CLK(n8383), .Q(
        g1273) );
  SDFFX1 DFF_768_Q_reg ( .D(g24510), .SI(g1273), .SE(n8196), .CLK(n8383), .Q(
        g1276) );
  SDFFX1 DFF_769_Q_reg ( .D(g24521), .SI(g1276), .SE(n8197), .CLK(n8384), .Q(
        g1279) );
  SDFFX1 DFF_770_Q_reg ( .D(g24511), .SI(g1279), .SE(n8197), .CLK(n8384), .Q(
        g1282) );
  SDFFX1 DFF_771_Q_reg ( .D(g24522), .SI(g1282), .SE(n8197), .CLK(n8384), .Q(
        g1285) );
  SDFFX1 DFF_772_Q_reg ( .D(g24532), .SI(g1285), .SE(n8197), .CLK(n8384), .Q(
        g1288) );
  SDFFX1 DFF_773_Q_reg ( .D(g28351), .SI(g1288), .SE(n8197), .CLK(n8384), .Q(
        g1300) );
  SDFFX1 DFF_774_Q_reg ( .D(g28355), .SI(g1300), .SE(n8197), .CLK(n8384), .Q(
        g1303) );
  SDFFX1 DFF_775_Q_reg ( .D(g28360), .SI(g1303), .SE(n8195), .CLK(n8382), .Q(
        g1306) );
  SDFFX1 DFF_776_Q_reg ( .D(g28346), .SI(g1306), .SE(n8197), .CLK(n8384), .Q(
        g1291) );
  SDFFX1 DFF_777_Q_reg ( .D(g28350), .SI(g1291), .SE(n8197), .CLK(n8384), .Q(
        g1294) );
  SDFFX1 DFF_778_Q_reg ( .D(g28354), .SI(g1294), .SE(n8197), .CLK(n8384), .Q(
        g1297) );
  SDFFX1 DFF_779_Q_reg ( .D(g26547), .SI(g1297), .SE(n8197), .CLK(n8384), .Q(
        test_so47) );
  SDFFX1 DFF_780_Q_reg ( .D(g26557), .SI(test_si48), .SE(n8195), .CLK(n8382), 
        .Q(g1180) );
  SDFFX1 DFF_781_Q_reg ( .D(g26569), .SI(g1180), .SE(n8195), .CLK(n8382), .Q(
        g1183) );
  SDFFX1 DFF_782_Q_reg ( .D(g1186), .SI(g1183), .SE(n8195), .CLK(n8382), .Q(
        g1192), .QN(n4454) );
  SDFFX1 DFF_783_Q_reg ( .D(g22615), .SI(g1192), .SE(n8198), .CLK(n8385), .Q(
        n8009), .QN(DFF_783_n1) );
  SDFFX1 DFF_792_Q_reg ( .D(n513), .SI(n8009), .SE(n8198), .CLK(n8385), .Q(
        g16355), .QN(DFF_792_n1) );
  SDFFX1 DFF_793_Q_reg ( .D(g16355), .SI(g16355), .SE(n8198), .CLK(n8385), .Q(
        g1211), .QN(n8037) );
  SDFFX1 DFF_794_Q_reg ( .D(DFF_649_n1), .SI(g1211), .SE(n8198), .CLK(n8385), 
        .Q(n8008), .QN(DFF_794_n1) );
  SDFFX1 DFF_795_Q_reg ( .D(DFF_651_n1), .SI(n8008), .SE(n8198), .CLK(n8385), 
        .Q(n8007), .QN(DFF_795_n1) );
  SDFFX1 DFF_796_Q_reg ( .D(DFF_653_n1), .SI(n8007), .SE(n8198), .CLK(n8385), 
        .Q(n8006), .QN(DFF_796_n1) );
  SDFFX1 DFF_797_Q_reg ( .D(DFF_655_n1), .SI(n8006), .SE(n8198), .CLK(n8385), 
        .Q(n8005), .QN(DFF_797_n1) );
  SDFFX1 DFF_798_Q_reg ( .D(DFF_657_n1), .SI(n8005), .SE(n8198), .CLK(n8385), 
        .Q(n8004), .QN(DFF_798_n1) );
  SDFFX1 DFF_799_Q_reg ( .D(DFF_659_n1), .SI(n8004), .SE(n8198), .CLK(n8385), 
        .Q(n8003), .QN(DFF_799_n1) );
  SDFFX1 DFF_800_Q_reg ( .D(DFF_661_n1), .SI(n8003), .SE(n8198), .CLK(n8385), 
        .Q(g1222), .QN(n7149) );
  SDFFX1 DFF_801_Q_reg ( .D(DFF_663_n1), .SI(g1222), .SE(n8198), .CLK(n8385), 
        .Q(g1223), .QN(n7148) );
  SDFFX1 DFF_802_Q_reg ( .D(g24072), .SI(g1223), .SE(n8199), .CLK(n8386), .Q(
        g1224), .QN(n4489) );
  SDFFX1 DFF_803_Q_reg ( .D(n4486), .SI(g1224), .SE(n8199), .CLK(n8386), .Q(
        test_so48), .QN(n14348) );
  SDFFX1 DFF_805_Q_reg ( .D(g6979), .SI(g6979), .SE(n8130), .CLK(n8317), .Q(
        g7161), .QN(n4358) );
  SDFFX1 DFF_806_Q_reg ( .D(g7161), .SI(g7161), .SE(n8130), .CLK(n8317), .Q(
        g1315), .QN(n4294) );
  SDFFX1 DFF_807_Q_reg ( .D(g16671), .SI(g1315), .SE(n8190), .CLK(n8377), .Q(
        g1316), .QN(n7747) );
  SDFFX1 DFF_808_Q_reg ( .D(g20333), .SI(g1316), .SE(n8190), .CLK(n8377), .Q(
        g1345), .QN(n4428) );
  SDFFX1 DFF_809_Q_reg ( .D(g20717), .SI(g1345), .SE(n8190), .CLK(n8377), .Q(
        g1326), .QN(n4402) );
  SDFFX1 DFF_810_Q_reg ( .D(n901), .SI(g1326), .SE(n8190), .CLK(n8377), .Q(
        g1319), .QN(n4476) );
  SDFFX1 DFF_811_Q_reg ( .D(g23329), .SI(g1319), .SE(n8190), .CLK(n8377), .Q(
        g1339), .QN(n4421) );
  SDFFX1 DFF_812_Q_reg ( .D(g24430), .SI(g1339), .SE(n8190), .CLK(n8377), .Q(
        g1332), .QN(n4412) );
  SDFFX1 DFF_813_Q_reg ( .D(g25189), .SI(g1332), .SE(n8190), .CLK(n8377), .Q(
        g1346), .QN(n4401) );
  SDFFX1 DFF_814_Q_reg ( .D(n902), .SI(g1346), .SE(n8190), .CLK(n8377), .Q(
        g1358), .QN(n4411) );
  SDFFX1 DFF_815_Q_reg ( .D(g26781), .SI(g1358), .SE(n8190), .CLK(n8377), .Q(
        g1352), .QN(n4469) );
  SDFFX1 DFF_816_Q_reg ( .D(g27678), .SI(g1352), .SE(n8190), .CLK(n8377), .Q(
        g1365), .QN(n4475) );
  SDFFX1 DFF_817_Q_reg ( .D(g27718), .SI(g1365), .SE(n8191), .CLK(n8378), .Q(
        g1372), .QN(n4395) );
  SDFFX1 DFF_818_Q_reg ( .D(g28321), .SI(g1372), .SE(n8191), .CLK(n8378), .Q(
        g1378), .QN(n4417) );
  SDFFX1 DFF_819_Q_reg ( .D(g20882), .SI(g1378), .SE(n8199), .CLK(n8386), .Q(
        test_so49), .QN(n8124) );
  SDFFX1 DFF_820_Q_reg ( .D(g20896), .SI(test_si50), .SE(n8199), .CLK(n8386), 
        .Q(g1386), .QN(n7808) );
  SDFFX1 DFF_821_Q_reg ( .D(g20910), .SI(g1386), .SE(n8199), .CLK(n8386), .Q(
        g1384), .QN(n7854) );
  SDFFX1 DFF_822_Q_reg ( .D(g20897), .SI(g1384), .SE(n8199), .CLK(n8386), .Q(
        g1388), .QN(n7807) );
  SDFFX1 DFF_823_Q_reg ( .D(g20911), .SI(g1388), .SE(n8199), .CLK(n8386), .Q(
        g1389), .QN(n7806) );
  SDFFX1 DFF_824_Q_reg ( .D(g20925), .SI(g1389), .SE(n8199), .CLK(n8386), .Q(
        g1387), .QN(n7853) );
  SDFFX1 DFF_825_Q_reg ( .D(g20912), .SI(g1387), .SE(n8199), .CLK(n8386), .Q(
        g1391), .QN(n7805) );
  SDFFX1 DFF_826_Q_reg ( .D(g20926), .SI(g1391), .SE(n8199), .CLK(n8386), .Q(
        g1392), .QN(n7804) );
  SDFFX1 DFF_827_Q_reg ( .D(g20949), .SI(g1392), .SE(n8199), .CLK(n8386), .Q(
        g1390), .QN(n7852) );
  SDFFX1 DFF_828_Q_reg ( .D(g20927), .SI(g1390), .SE(n8199), .CLK(n8386), .Q(
        g1394), .QN(n7803) );
  SDFFX1 DFF_829_Q_reg ( .D(g20950), .SI(g1394), .SE(n8200), .CLK(n8387), .Q(
        g1395), .QN(n7802) );
  SDFFX1 DFF_830_Q_reg ( .D(g20972), .SI(g1395), .SE(n8200), .CLK(n8387), .Q(
        g1393), .QN(n7851) );
  SDFFX1 DFF_831_Q_reg ( .D(g20951), .SI(g1393), .SE(n8200), .CLK(n8387), .Q(
        g1397), .QN(n7801) );
  SDFFX1 DFF_832_Q_reg ( .D(g20973), .SI(g1397), .SE(n8200), .CLK(n8387), .Q(
        g1398), .QN(n7800) );
  SDFFX1 DFF_833_Q_reg ( .D(g20993), .SI(g1398), .SE(n8200), .CLK(n8387), .Q(
        g1396), .QN(n7850) );
  SDFFX1 DFF_834_Q_reg ( .D(g20974), .SI(g1396), .SE(n8200), .CLK(n8387), .Q(
        g1400), .QN(n7799) );
  SDFFX1 DFF_835_Q_reg ( .D(g20994), .SI(g1400), .SE(n8200), .CLK(n8387), .Q(
        test_so50), .QN(n8123) );
  SDFFX1 DFF_836_Q_reg ( .D(g21015), .SI(test_si51), .SE(n8200), .CLK(n8387), 
        .Q(g1399), .QN(n7849) );
  SDFFX1 DFF_837_Q_reg ( .D(g20995), .SI(g1399), .SE(n8200), .CLK(n8387), .Q(
        g1403), .QN(n7798) );
  SDFFX1 DFF_838_Q_reg ( .D(g21016), .SI(g1403), .SE(n8200), .CLK(n8387), .Q(
        g1404), .QN(n7797) );
  SDFFX1 DFF_839_Q_reg ( .D(g21033), .SI(g1404), .SE(n8200), .CLK(n8387), .Q(
        g1402), .QN(n7848) );
  SDFFX1 DFF_840_Q_reg ( .D(g21017), .SI(g1402), .SE(n8200), .CLK(n8387), .Q(
        g1406), .QN(n7796) );
  SDFFX1 DFF_841_Q_reg ( .D(g21034), .SI(g1406), .SE(n8201), .CLK(n8388), .Q(
        g1407), .QN(n7795) );
  SDFFX1 DFF_842_Q_reg ( .D(g21052), .SI(g1407), .SE(n8201), .CLK(n8388), .Q(
        g1405), .QN(n7847) );
  SDFFX1 DFF_843_Q_reg ( .D(g21035), .SI(g1405), .SE(n8201), .CLK(n8388), .Q(
        g1409), .QN(n7794) );
  SDFFX1 DFF_844_Q_reg ( .D(g21053), .SI(g1409), .SE(n8201), .CLK(n8388), .Q(
        g1410), .QN(n7793) );
  SDFFX1 DFF_845_Q_reg ( .D(g21070), .SI(g1410), .SE(n8201), .CLK(n8388), .Q(
        g1408), .QN(n7846) );
  SDFFX1 DFF_846_Q_reg ( .D(g20883), .SI(g1408), .SE(n8201), .CLK(n8388), .Q(
        g1412), .QN(n7792) );
  SDFFX1 DFF_847_Q_reg ( .D(g20898), .SI(g1412), .SE(n8201), .CLK(n8388), .Q(
        g1413), .QN(n7791) );
  SDFFX1 DFF_848_Q_reg ( .D(g20913), .SI(g1413), .SE(n8201), .CLK(n8388), .Q(
        g1411), .QN(n7845) );
  SDFFX1 DFF_849_Q_reg ( .D(g20952), .SI(g1411), .SE(n8201), .CLK(n8388), .Q(
        g1415), .QN(n8023) );
  SDFFX1 DFF_850_Q_reg ( .D(g20975), .SI(g1415), .SE(n8201), .CLK(n8388), .Q(
        g1416), .QN(n7560) );
  SDFFX1 DFF_851_Q_reg ( .D(g20996), .SI(g1416), .SE(n8201), .CLK(n8388), .Q(
        test_so51) );
  SDFFX1 DFF_852_Q_reg ( .D(g20976), .SI(test_si52), .SE(n8197), .CLK(n8384), 
        .Q(g1418), .QN(n7565) );
  SDFFX1 DFF_853_Q_reg ( .D(g20997), .SI(g1418), .SE(n8197), .CLK(n8384), .Q(
        g1419), .QN(n7559) );
  SDFFX1 DFF_854_Q_reg ( .D(g21018), .SI(g1419), .SE(n8198), .CLK(n8385), .Q(
        g1417), .QN(n7617) );
  SDFFX1 DFF_855_Q_reg ( .D(g25263), .SI(g1417), .SE(n8201), .CLK(n8388), .Q(
        g1421), .QN(n7495) );
  SDFFX1 DFF_856_Q_reg ( .D(g25267), .SI(g1421), .SE(n8202), .CLK(n8389), .Q(
        g1422), .QN(n7494) );
  SDFFX1 DFF_857_Q_reg ( .D(g25270), .SI(g1422), .SE(n8202), .CLK(n8389), .Q(
        g1420), .QN(n7500) );
  SDFFX1 DFF_858_Q_reg ( .D(g22234), .SI(g1420), .SE(n8202), .CLK(n8389), .Q(
        g1424), .QN(n7867) );
  SDFFX1 DFF_859_Q_reg ( .D(n872), .SI(g1424), .SE(n8202), .CLK(n8389), .Q(
        g1425), .QN(n7955) );
  SDFFX1 DFF_860_Q_reg ( .D(g22263), .SI(g1425), .SE(n8202), .CLK(n8389), .Q(
        g1423), .QN(n7958) );
  SDFFX1 DFF_861_Q_reg ( .D(g2950), .SI(g1423), .SE(n8202), .CLK(n8389), .Q(
        g6573), .QN(n4317) );
  SDFFX1 DFF_862_Q_reg ( .D(g6573), .SI(g6573), .SE(n8202), .CLK(n8389), .Q(
        g6782), .QN(n4515) );
  SDFFX1 DFF_863_Q_reg ( .D(g6782), .SI(g6782), .SE(n8202), .CLK(n8389), .Q(
        g1547), .QN(n4368) );
  SDFFX1 DFF_864_Q_reg ( .D(g22149), .SI(g1547), .SE(n8203), .CLK(n8390), .Q(
        g1512), .QN(n7897) );
  SDFFX1 DFF_865_Q_reg ( .D(g22166), .SI(g1512), .SE(n8205), .CLK(n8392), .Q(
        g1513), .QN(n7896) );
  SDFFX1 DFF_866_Q_reg ( .D(g22178), .SI(g1513), .SE(n8205), .CLK(n8392), .Q(
        g1511), .QN(n7531) );
  SDFFX1 DFF_867_Q_reg ( .D(g22167), .SI(g1511), .SE(n8203), .CLK(n8390), .Q(
        test_so52), .QN(n8093) );
  SDFFX1 DFF_868_Q_reg ( .D(g22179), .SI(test_si53), .SE(n8206), .CLK(n8393), 
        .Q(g1516), .QN(n7895) );
  SDFFX1 DFF_869_Q_reg ( .D(g22191), .SI(g1516), .SE(n8206), .CLK(n8393), .Q(
        g1514), .QN(n7530) );
  SDFFX1 DFF_870_Q_reg ( .D(g22035), .SI(g1514), .SE(n8206), .CLK(n8393), .Q(
        g1524), .QN(n7894) );
  SDFFX1 DFF_871_Q_reg ( .D(g22043), .SI(g1524), .SE(n8206), .CLK(n8393), .Q(
        g1525), .QN(n7893) );
  SDFFX1 DFF_872_Q_reg ( .D(g22057), .SI(g1525), .SE(n8207), .CLK(n8394), .Q(
        g1523), .QN(n7529) );
  SDFFX1 DFF_873_Q_reg ( .D(g22044), .SI(g1523), .SE(n8207), .CLK(n8394), .Q(
        g1527), .QN(n7892) );
  SDFFX1 DFF_874_Q_reg ( .D(g22058), .SI(g1527), .SE(n8207), .CLK(n8394), .Q(
        g1528), .QN(n7891) );
  SDFFX1 DFF_875_Q_reg ( .D(g22073), .SI(g1528), .SE(n8207), .CLK(n8394), .Q(
        g1526), .QN(n7528) );
  SDFFX1 DFF_876_Q_reg ( .D(g22059), .SI(g1526), .SE(n8207), .CLK(n8394), .Q(
        g1530), .QN(n7890) );
  SDFFX1 DFF_877_Q_reg ( .D(g22074), .SI(g1530), .SE(n8207), .CLK(n8394), .Q(
        g1531), .QN(n7889) );
  SDFFX1 DFF_878_Q_reg ( .D(g22090), .SI(g1531), .SE(n8207), .CLK(n8394), .Q(
        g1529), .QN(n7527) );
  SDFFX1 DFF_879_Q_reg ( .D(g22075), .SI(g1529), .SE(n8207), .CLK(n8394), .Q(
        g1533), .QN(n7888) );
  SDFFX1 DFF_880_Q_reg ( .D(g22091), .SI(g1533), .SE(n8207), .CLK(n8394), .Q(
        g1534), .QN(n7887) );
  SDFFX1 DFF_881_Q_reg ( .D(g22112), .SI(g1534), .SE(n8207), .CLK(n8394), .Q(
        g1532), .QN(n7526) );
  SDFFX1 DFF_882_Q_reg ( .D(g22092), .SI(g1532), .SE(n8207), .CLK(n8394), .Q(
        g1536), .QN(n7886) );
  SDFFX1 DFF_883_Q_reg ( .D(g22113), .SI(g1536), .SE(n8207), .CLK(n8394), .Q(
        test_so53), .QN(n8112) );
  SDFFX1 DFF_884_Q_reg ( .D(g22130), .SI(test_si54), .SE(n8205), .CLK(n8392), 
        .Q(g1535), .QN(n7525) );
  SDFFX1 DFF_885_Q_reg ( .D(g22114), .SI(g1535), .SE(n8205), .CLK(n8392), .Q(
        g1539), .QN(n7885) );
  SDFFX1 DFF_886_Q_reg ( .D(g22131), .SI(g1539), .SE(n8205), .CLK(n8392), .Q(
        g1540), .QN(n7884) );
  SDFFX1 DFF_887_Q_reg ( .D(g22150), .SI(g1540), .SE(n8205), .CLK(n8392), .Q(
        g1538), .QN(n7524) );
  SDFFX1 DFF_888_Q_reg ( .D(g22132), .SI(g1538), .SE(n8205), .CLK(n8392), .Q(
        g1542), .QN(n7507) );
  SDFFX1 DFF_889_Q_reg ( .D(g22151), .SI(g1542), .SE(n8205), .CLK(n8392), .Q(
        g1543), .QN(n7506) );
  SDFFX1 DFF_890_Q_reg ( .D(g22168), .SI(g1543), .SE(n8205), .CLK(n8392), .Q(
        g1541), .QN(n7505) );
  SDFFX1 DFF_891_Q_reg ( .D(g22152), .SI(g1541), .SE(n8206), .CLK(n8393), .Q(
        g1545), .QN(n7523) );
  SDFFX1 DFF_892_Q_reg ( .D(g22169), .SI(g1545), .SE(n8205), .CLK(n8392), .Q(
        g1546), .QN(n7522) );
  SDFFX1 DFF_893_Q_reg ( .D(g22180), .SI(g1546), .SE(n8206), .CLK(n8393), .Q(
        g1544), .QN(n7521) );
  SDFFX1 DFF_894_Q_reg ( .D(g25217), .SI(g1544), .SE(n8206), .CLK(n8393), .Q(
        g1551), .QN(n7589) );
  SDFFX1 DFF_895_Q_reg ( .D(g25224), .SI(g1551), .SE(n8206), .CLK(n8393), .Q(
        g1552), .QN(n7588) );
  SDFFX1 DFF_896_Q_reg ( .D(g25233), .SI(g1552), .SE(n8206), .CLK(n8393), .Q(
        g1550), .QN(n7587) );
  SDFFX1 DFF_897_Q_reg ( .D(g25225), .SI(g1550), .SE(n8206), .CLK(n8393), .Q(
        g1554), .QN(n7586) );
  SDFFX1 DFF_898_Q_reg ( .D(g25234), .SI(g1554), .SE(n8206), .CLK(n8393), .Q(
        g1555), .QN(n7585) );
  SDFFX1 DFF_899_Q_reg ( .D(g25242), .SI(g1555), .SE(n8206), .CLK(n8393), .Q(
        test_so54), .QN(n8129) );
  SDFFX1 DFF_900_Q_reg ( .D(g25235), .SI(test_si55), .SE(n8202), .CLK(n8389), 
        .Q(g1557), .QN(n7584) );
  SDFFX1 DFF_901_Q_reg ( .D(g25243), .SI(g1557), .SE(n8202), .CLK(n8389), .Q(
        g1558), .QN(n7583) );
  SDFFX1 DFF_902_Q_reg ( .D(g25249), .SI(g1558), .SE(n8202), .CLK(n8389), .Q(
        g1556), .QN(n7582) );
  SDFFX1 DFF_903_Q_reg ( .D(g25244), .SI(g1556), .SE(n8202), .CLK(n8389), .Q(
        g1560), .QN(n7581) );
  SDFFX1 DFF_904_Q_reg ( .D(g25250), .SI(g1560), .SE(n8203), .CLK(n8390), .Q(
        g1561), .QN(n7580) );
  SDFFX1 DFF_905_Q_reg ( .D(g25255), .SI(g1561), .SE(n8203), .CLK(n8390), .Q(
        g1559), .QN(n7579) );
  SDFFX1 DFF_906_Q_reg ( .D(g30279), .SI(g1559), .SE(n8212), .CLK(n8399), .Q(
        g1567) );
  SDFFX1 DFF_907_Q_reg ( .D(g30287), .SI(g1567), .SE(n8212), .CLK(n8399), .Q(
        g1570) );
  SDFFX1 DFF_908_Q_reg ( .D(g30294), .SI(g1570), .SE(n8212), .CLK(n8399), .Q(
        g1573) );
  SDFFX1 DFF_909_Q_reg ( .D(g30651), .SI(g1573), .SE(n8213), .CLK(n8400), .Q(
        g1612) );
  SDFFX1 DFF_910_Q_reg ( .D(g30657), .SI(g1612), .SE(n8213), .CLK(n8400), .Q(
        g1615) );
  SDFFX1 DFF_911_Q_reg ( .D(g30663), .SI(g1615), .SE(n8213), .CLK(n8400), .Q(
        g1618) );
  SDFFX1 DFF_912_Q_reg ( .D(g30683), .SI(g1618), .SE(n8213), .CLK(n8400), .Q(
        g1576) );
  SDFFX1 DFF_913_Q_reg ( .D(g30688), .SI(g1576), .SE(n8213), .CLK(n8400), .Q(
        g1579) );
  SDFFX1 DFF_914_Q_reg ( .D(g30692), .SI(g1579), .SE(n8208), .CLK(n8395), .Q(
        g1582) );
  SDFFX1 DFF_915_Q_reg ( .D(g30658), .SI(g1582), .SE(n8208), .CLK(n8395), .Q(
        test_so55) );
  SDFFX1 DFF_916_Q_reg ( .D(g30664), .SI(test_si56), .SE(n8208), .CLK(n8395), 
        .Q(g1624) );
  SDFFX1 DFF_917_Q_reg ( .D(g30671), .SI(g1624), .SE(n8208), .CLK(n8395), .Q(
        g1627) );
  SDFFX1 DFF_918_Q_reg ( .D(g30295), .SI(g1627), .SE(n8208), .CLK(n8395), .Q(
        g1585) );
  SDFFX1 DFF_919_Q_reg ( .D(g30299), .SI(g1585), .SE(n8208), .CLK(n8395), .Q(
        g1588) );
  SDFFX1 DFF_920_Q_reg ( .D(g30302), .SI(g1588), .SE(n8208), .CLK(n8395), .Q(
        g1591) );
  SDFFX1 DFF_921_Q_reg ( .D(g30266), .SI(g1591), .SE(n8208), .CLK(n8395), .Q(
        g1630) );
  SDFFX1 DFF_922_Q_reg ( .D(g30272), .SI(g1630), .SE(n8208), .CLK(n8395), .Q(
        g1633) );
  SDFFX1 DFF_923_Q_reg ( .D(g30280), .SI(g1633), .SE(n8208), .CLK(n8395), .Q(
        g1636) );
  SDFFX1 DFF_924_Q_reg ( .D(g30250), .SI(g1636), .SE(n8212), .CLK(n8399), .Q(
        g1594) );
  SDFFX1 DFF_925_Q_reg ( .D(g30252), .SI(g1594), .SE(n8212), .CLK(n8399), .Q(
        g1597) );
  SDFFX1 DFF_926_Q_reg ( .D(g30255), .SI(g1597), .SE(n8212), .CLK(n8399), .Q(
        g1600) );
  SDFFX1 DFF_927_Q_reg ( .D(g30273), .SI(g1600), .SE(n8212), .CLK(n8399), .Q(
        g1639) );
  SDFFX1 DFF_928_Q_reg ( .D(g30281), .SI(g1639), .SE(n8212), .CLK(n8399), .Q(
        g1642) );
  SDFFX1 DFF_929_Q_reg ( .D(g30288), .SI(g1642), .SE(n8212), .CLK(n8399), .Q(
        g1645) );
  SDFFX1 DFF_930_Q_reg ( .D(g30644), .SI(g1645), .SE(n8212), .CLK(n8399), .Q(
        g1603) );
  SDFFX1 DFF_931_Q_reg ( .D(g30650), .SI(g1603), .SE(n8212), .CLK(n8399), .Q(
        test_so56) );
  SDFFX1 DFF_932_Q_reg ( .D(g30656), .SI(test_si57), .SE(n8208), .CLK(n8395), 
        .Q(g1609) );
  SDFFX1 DFF_933_Q_reg ( .D(g30678), .SI(g1609), .SE(n8208), .CLK(n8395), .Q(
        g1648) );
  SDFFX1 DFF_934_Q_reg ( .D(g30684), .SI(g1648), .SE(n8209), .CLK(n8396), .Q(
        g1651) );
  SDFFX1 DFF_935_Q_reg ( .D(g30689), .SI(g1651), .SE(n8203), .CLK(n8390), .Q(
        g1654) );
  SDFFX1 DFF_936_Q_reg ( .D(g25056), .SI(g1654), .SE(n8203), .CLK(n8390), .Q(
        g1466), .QN(n7694) );
  SDFFX1 DFF_937_Q_reg ( .D(g25938), .SI(g1466), .SE(n8203), .CLK(n8390), .Q(
        g1462), .QN(n8042) );
  SDFFX1 DFF_938_Q_reg ( .D(g26531), .SI(g1462), .SE(n8203), .CLK(n8390), .Q(
        g1457), .QN(n7693) );
  SDFFX1 DFF_939_Q_reg ( .D(g27129), .SI(g1457), .SE(n8203), .CLK(n8390), .Q(
        g1453) );
  SDFFX1 DFF_940_Q_reg ( .D(g27612), .SI(g1453), .SE(n8203), .CLK(n8390), .Q(
        g1448), .QN(n7692) );
  SDFFX1 DFF_941_Q_reg ( .D(g28147), .SI(g1448), .SE(n8204), .CLK(n8391), .Q(
        g1444), .QN(n8068) );
  SDFFX1 DFF_942_Q_reg ( .D(g28636), .SI(g1444), .SE(n8204), .CLK(n8391), .Q(
        g1439), .QN(n7691) );
  SDFFX1 DFF_943_Q_reg ( .D(g29111), .SI(g1439), .SE(n8204), .CLK(n8391), .Q(
        g1435), .QN(n8049) );
  SDFFX1 DFF_944_Q_reg ( .D(g29355), .SI(g1435), .SE(n8204), .CLK(n8391), .Q(
        g1430), .QN(n7323) );
  SDFFX1 DFF_945_Q_reg ( .D(g29581), .SI(g1430), .SE(n8204), .CLK(n8391), .Q(
        g1426), .QN(n7162) );
  SDFFX1 DFF_946_Q_reg ( .D(n19), .SI(g1426), .SE(n8204), .CLK(n8391), .Q(
        g1562) );
  SDFFX1 DFF_947_Q_reg ( .D(g1562), .SI(g1562), .SE(n8204), .CLK(n8391), .Q(
        test_so57) );
  SDFFX1 DFF_948_Q_reg ( .D(test_so57), .SI(test_si58), .SE(n8204), .CLK(n8391), .Q(g1563), .QN(n7707) );
  SDFFX1 DFF_949_Q_reg ( .D(g2950), .SI(g1563), .SE(n8204), .CLK(n8391), .Q(
        g5511), .QN(n4518) );
  SDFFX1 DFF_952_Q_reg ( .D(test_so57), .SI(n4618), .SE(n8204), .CLK(n8391), 
        .Q(g1690), .QN(n4386) );
  SDFFX1 DFF_953_Q_reg ( .D(g27264), .SI(g1690), .SE(n8211), .CLK(n8398), .Q(
        g1735), .QN(n7648) );
  SDFFX1 DFF_954_Q_reg ( .D(g27274), .SI(g1735), .SE(n8211), .CLK(n8398), .Q(
        g1724), .QN(n7647) );
  SDFFX1 DFF_955_Q_reg ( .D(g27287), .SI(g1724), .SE(n8211), .CLK(n8398), .Q(
        g1727), .QN(n7646) );
  SDFFX1 DFF_956_Q_reg ( .D(g27275), .SI(g1727), .SE(n8211), .CLK(n8398), .Q(
        g1750), .QN(n7625) );
  SDFFX1 DFF_957_Q_reg ( .D(g27288), .SI(g1750), .SE(n8211), .CLK(n8398), .Q(
        g1739), .QN(n7624) );
  SDFFX1 DFF_958_Q_reg ( .D(g27302), .SI(g1739), .SE(n8211), .CLK(n8398), .Q(
        g1742), .QN(n7623) );
  SDFFX1 DFF_959_Q_reg ( .D(g27289), .SI(g1742), .SE(n8211), .CLK(n8398), .Q(
        g1765), .QN(n7374) );
  SDFFX1 DFF_960_Q_reg ( .D(g27303), .SI(g1765), .SE(n8211), .CLK(n8398), .Q(
        g1754), .QN(n7376) );
  SDFFX1 DFF_961_Q_reg ( .D(g27317), .SI(g1754), .SE(n8211), .CLK(n8398), .Q(
        g1757), .QN(n7375) );
  SDFFX1 DFF_962_Q_reg ( .D(g27304), .SI(g1757), .SE(n8211), .CLK(n8398), .Q(
        g1779), .QN(n7636) );
  SDFFX1 DFF_963_Q_reg ( .D(g27318), .SI(g1779), .SE(n8212), .CLK(n8399), .Q(
        test_so58), .QN(n8096) );
  SDFFX1 DFF_964_Q_reg ( .D(g27330), .SI(test_si59), .SE(n8209), .CLK(n8396), 
        .Q(g1772), .QN(n7635) );
  SDFFX1 DFF_965_Q_reg ( .D(g28749), .SI(g1772), .SE(n8209), .CLK(n8396), .Q(
        g1789) );
  SDFFX1 DFF_966_Q_reg ( .D(g28760), .SI(g1789), .SE(n8210), .CLK(n8397), .Q(
        g1792) );
  SDFFX1 DFF_967_Q_reg ( .D(g28771), .SI(g1792), .SE(n8210), .CLK(n8397), .Q(
        g1795) );
  SDFFX1 DFF_968_Q_reg ( .D(g29205), .SI(g1795), .SE(n8210), .CLK(n8397), .Q(
        g1798) );
  SDFFX1 DFF_969_Q_reg ( .D(g29212), .SI(g1798), .SE(n8211), .CLK(n8398), .Q(
        g1801) );
  SDFFX1 DFF_970_Q_reg ( .D(g29218), .SI(g1801), .SE(n8209), .CLK(n8396), .Q(
        g1804) );
  SDFFX1 DFF_971_Q_reg ( .D(g28761), .SI(g1804), .SE(n8209), .CLK(n8396), .Q(
        g1808), .QN(n7671) );
  SDFFX1 DFF_972_Q_reg ( .D(g28772), .SI(g1808), .SE(n8209), .CLK(n8396), .Q(
        g1809), .QN(n7659) );
  SDFFX1 DFF_973_Q_reg ( .D(g28778), .SI(g1809), .SE(n8209), .CLK(n8396), .Q(
        g1807), .QN(n7670) );
  SDFFX1 DFF_974_Q_reg ( .D(g26811), .SI(g1807), .SE(n8209), .CLK(n8396), .Q(
        g1810) );
  SDFFX1 DFF_975_Q_reg ( .D(g26815), .SI(g1810), .SE(n8209), .CLK(n8396), .Q(
        g1813) );
  SDFFX1 DFF_976_Q_reg ( .D(g26820), .SI(g1813), .SE(n8210), .CLK(n8397), .Q(
        g1816) );
  SDFFX1 DFF_977_Q_reg ( .D(g26816), .SI(g1816), .SE(n8210), .CLK(n8397), .Q(
        g1819) );
  SDFFX1 DFF_978_Q_reg ( .D(g26821), .SI(g1819), .SE(n8210), .CLK(n8397), .Q(
        g1822) );
  SDFFX1 DFF_979_Q_reg ( .D(g26824), .SI(g1822), .SE(n8210), .CLK(n8397), .Q(
        test_so59) );
  SDFFX1 DFF_980_Q_reg ( .D(g27764), .SI(test_si60), .SE(n8210), .CLK(n8397), 
        .Q(g1829), .QN(n7669) );
  SDFFX1 DFF_981_Q_reg ( .D(g27766), .SI(g1829), .SE(n8210), .CLK(n8397), .Q(
        g1830), .QN(n7658) );
  SDFFX1 DFF_982_Q_reg ( .D(g27768), .SI(g1830), .SE(n8210), .CLK(n8397), .Q(
        g1828), .QN(n7668) );
  SDFFX1 DFF_983_Q_reg ( .D(g29613), .SI(g1828), .SE(n8210), .CLK(n8397), .Q(
        g1693), .QN(n7276) );
  SDFFX1 DFF_984_Q_reg ( .D(g29617), .SI(g1693), .SE(n8210), .CLK(n8397), .Q(
        g1694), .QN(n7261) );
  SDFFX1 DFF_985_Q_reg ( .D(g29620), .SI(g1694), .SE(n8209), .CLK(n8396), .Q(
        g1695), .QN(n7275) );
  SDFFX1 DFF_986_Q_reg ( .D(g30704), .SI(g1695), .SE(n8209), .CLK(n8396), .Q(
        g1696), .QN(n7274) );
  SDFFX1 DFF_987_Q_reg ( .D(g30706), .SI(g1696), .SE(n8209), .CLK(n8396), .Q(
        g1697), .QN(n7260) );
  SDFFX1 DFF_988_Q_reg ( .D(g30708), .SI(g1697), .SE(n8203), .CLK(n8390), .Q(
        g1698), .QN(n7273) );
  SDFFX1 DFF_989_Q_reg ( .D(g30487), .SI(g1698), .SE(n8205), .CLK(n8392), .Q(
        g1699), .QN(n7272) );
  SDFFX1 DFF_990_Q_reg ( .D(g30503), .SI(g1699), .SE(n8203), .CLK(n8390), .Q(
        g1700), .QN(n7259) );
  SDFFX1 DFF_991_Q_reg ( .D(g30338), .SI(g1700), .SE(n8205), .CLK(n8392), .Q(
        g1701), .QN(n7271) );
  SDFFX1 DFF_992_Q_reg ( .D(g29178), .SI(g1701), .SE(n8213), .CLK(n8400), .Q(
        g1703), .QN(n7316) );
  SDFFX1 DFF_993_Q_reg ( .D(g29181), .SI(g1703), .SE(n8213), .CLK(n8400), .Q(
        g1704), .QN(n7311) );
  SDFFX1 DFF_994_Q_reg ( .D(g29184), .SI(g1704), .SE(n8213), .CLK(n8400), .Q(
        g1702), .QN(n7315) );
  SDFFX1 DFF_995_Q_reg ( .D(g26667), .SI(g1702), .SE(n8213), .CLK(n8400), .Q(
        test_so60), .QN(n8111) );
  SDFFX1 DFF_996_Q_reg ( .D(g26670), .SI(test_si61), .SE(n8213), .CLK(n8400), 
        .Q(g1785), .QN(n7657) );
  SDFFX1 DFF_997_Q_reg ( .D(g26675), .SI(g1785), .SE(n8213), .CLK(n8400), .Q(
        g1783), .QN(n7667) );
  SDFFX1 DFF_998_Q_reg ( .D(n4288), .SI(g1783), .SE(n8213), .CLK(n8400), .Q(
        g1831) );
  SDFFX1 DFF_999_Q_reg ( .D(g1831), .SI(g1831), .SE(n8214), .CLK(n8401), .Q(
        n7988), .QN(DFF_999_n1) );
  SDFFX1 DFF_1000_Q_reg ( .D(n4565), .SI(n7988), .SE(n8214), .CLK(n8401), .Q(
        g1833) );
  SDFFX1 DFF_1001_Q_reg ( .D(g1833), .SI(g1833), .SE(n8214), .CLK(n8401), .Q(
        n7987), .QN(DFF_1001_n1) );
  SDFFX1 DFF_1002_Q_reg ( .D(n4557), .SI(n7987), .SE(n8214), .CLK(n8401), .Q(
        g1835) );
  SDFFX1 DFF_1003_Q_reg ( .D(g1835), .SI(g1835), .SE(n8214), .CLK(n8401), .Q(
        n7986), .QN(DFF_1003_n1) );
  SDFFX1 DFF_1004_Q_reg ( .D(n4326), .SI(n7986), .SE(n8214), .CLK(n8401), .Q(
        g1661) );
  SDFFX1 DFF_1005_Q_reg ( .D(g1661), .SI(g1661), .SE(n8214), .CLK(n8401), .Q(
        n7985), .QN(DFF_1005_n1) );
  SDFFX1 DFF_1006_Q_reg ( .D(n4390), .SI(n7985), .SE(n8214), .CLK(n8401), .Q(
        g1663) );
  SDFFX1 DFF_1007_Q_reg ( .D(g1663), .SI(g1663), .SE(n8214), .CLK(n8401), .Q(
        n7984), .QN(DFF_1007_n1) );
  SDFFX1 DFF_1008_Q_reg ( .D(n4320), .SI(n7984), .SE(n8214), .CLK(n8401), .Q(
        g1665) );
  SDFFX1 DFF_1009_Q_reg ( .D(g1665), .SI(g1665), .SE(n8214), .CLK(n8401), .Q(
        n7983), .QN(DFF_1009_n1) );
  SDFFX1 DFF_1010_Q_reg ( .D(n4374), .SI(n7983), .SE(n8214), .CLK(n8401), .Q(
        g1667) );
  SDFFX1 DFF_1011_Q_reg ( .D(g1667), .SI(g1667), .SE(n8215), .CLK(n8402), .Q(
        test_so61), .QN(DFF_1011_n1) );
  SDFFX1 DFF_1012_Q_reg ( .D(n4378), .SI(test_si62), .SE(n8133), .CLK(n8320), 
        .Q(g1669) );
  SDFFX1 DFF_1013_Q_reg ( .D(g1669), .SI(g1669), .SE(n8133), .CLK(n8320), .Q(
        n7980), .QN(DFF_1013_n1) );
  SDFFX1 DFF_1014_Q_reg ( .D(g2877), .SI(n7980), .SE(n8138), .CLK(n8325), .Q(
        g1671) );
  SDFFX1 DFF_1015_Q_reg ( .D(g1671), .SI(g1671), .SE(n8138), .CLK(n8325), .Q(
        n7979), .QN(n4484) );
  SDFFX1 DFF_1016_Q_reg ( .D(n4284), .SI(n7979), .SE(n8211), .CLK(n8398), .Q(
        g1680), .QN(n4488) );
  SDFFX1 DFF_1017_Q_reg ( .D(n437), .SI(g1680), .SE(n8215), .CLK(n8402), .Q(
        g1686) );
  SDFFX1 DFF_1028_Q_reg ( .D(n4276), .SI(g1686), .SE(n8215), .CLK(n8402), .Q(
        n7978) );
  SDFFX1 DFF_1029_Q_reg ( .D(g1735), .SI(n7978), .SE(n8215), .CLK(n8402), .Q(
        g1723) );
  SDFFX1 DFF_1030_Q_reg ( .D(g1723), .SI(g1723), .SE(n8215), .CLK(n8402), .Q(
        g1730) );
  SDFFX1 DFF_1031_Q_reg ( .D(g1724), .SI(g1730), .SE(n8215), .CLK(n8402), .Q(
        g1731) );
  SDFFX1 DFF_1032_Q_reg ( .D(g1731), .SI(g1731), .SE(n8215), .CLK(n8402), .Q(
        g1732) );
  SDFFX1 DFF_1033_Q_reg ( .D(g1727), .SI(g1732), .SE(n8215), .CLK(n8402), .Q(
        g1733) );
  SDFFX1 DFF_1034_Q_reg ( .D(g1733), .SI(g1733), .SE(n8215), .CLK(n8402), .Q(
        g1734) );
  SDFFX1 DFF_1035_Q_reg ( .D(g1750), .SI(g1734), .SE(n8215), .CLK(n8402), .Q(
        g1738) );
  SDFFX1 DFF_1036_Q_reg ( .D(g1738), .SI(g1738), .SE(n8215), .CLK(n8402), .Q(
        g1745) );
  SDFFX1 DFF_1037_Q_reg ( .D(g1739), .SI(g1745), .SE(n8215), .CLK(n8402), .Q(
        test_so62) );
  SDFFX1 DFF_1038_Q_reg ( .D(test_so62), .SI(test_si63), .SE(n8216), .CLK(
        n8403), .Q(g1747) );
  SDFFX1 DFF_1039_Q_reg ( .D(g1742), .SI(g1747), .SE(n8216), .CLK(n8403), .Q(
        g1748) );
  SDFFX1 DFF_1040_Q_reg ( .D(g1748), .SI(g1748), .SE(n8216), .CLK(n8403), .Q(
        g1749) );
  SDFFX1 DFF_1041_Q_reg ( .D(g1765), .SI(g1749), .SE(n8216), .CLK(n8403), .Q(
        g1753) );
  SDFFX1 DFF_1042_Q_reg ( .D(g1753), .SI(g1753), .SE(n8216), .CLK(n8403), .Q(
        g1760) );
  SDFFX1 DFF_1043_Q_reg ( .D(g1754), .SI(g1760), .SE(n8216), .CLK(n8403), .Q(
        g1761) );
  SDFFX1 DFF_1044_Q_reg ( .D(g1761), .SI(g1761), .SE(n8216), .CLK(n8403), .Q(
        g1762) );
  SDFFX1 DFF_1045_Q_reg ( .D(g1757), .SI(g1762), .SE(n8216), .CLK(n8403), .Q(
        g1763) );
  SDFFX1 DFF_1046_Q_reg ( .D(g1763), .SI(g1763), .SE(n8216), .CLK(n8403), .Q(
        g1764) );
  SDFFX1 DFF_1047_Q_reg ( .D(g1779), .SI(g1764), .SE(n8216), .CLK(n8403), .Q(
        g1768) );
  SDFFX1 DFF_1048_Q_reg ( .D(g1768), .SI(g1768), .SE(n8216), .CLK(n8403), .Q(
        g1775) );
  SDFFX1 DFF_1049_Q_reg ( .D(test_so58), .SI(g1775), .SE(n8216), .CLK(n8403), 
        .Q(g1776) );
  SDFFX1 DFF_1050_Q_reg ( .D(g1776), .SI(g1776), .SE(n8217), .CLK(n8404), .Q(
        g1777) );
  SDFFX1 DFF_1051_Q_reg ( .D(g1772), .SI(g1777), .SE(n8217), .CLK(n8404), .Q(
        g1778) );
  SDFFX1 DFF_1052_Q_reg ( .D(g1778), .SI(g1778), .SE(n8217), .CLK(n8404), .Q(
        g1705) );
  SDFFX1 DFF_1053_Q_reg ( .D(n4598), .SI(g1705), .SE(n8217), .CLK(n8404), .Q(
        test_so63) );
  SDFFX1 DFF_1054_Q_reg ( .D(test_so63), .SI(test_si64), .SE(n8217), .CLK(
        n8404), .Q(g5738) );
  SDFFX1 DFF_1055_Q_reg ( .D(g5738), .SI(g5738), .SE(n8217), .CLK(n8404), .Q(
        g1718) );
  SDFFX1 DFF_1056_Q_reg ( .D(n4598), .SI(g1718), .SE(n8217), .CLK(n8404), .Q(
        g7052), .QN(n4296) );
  SDFFX1 DFF_1057_Q_reg ( .D(g7052), .SI(g7052), .SE(n8217), .CLK(n8404), .Q(
        g7194), .QN(n4315) );
  SDFFX1 DFF_1058_Q_reg ( .D(g7194), .SI(g7194), .SE(n8217), .CLK(n8404), .Q(
        g1930), .QN(n4366) );
  SDFFX1 DFF_1059_Q_reg ( .D(n1141), .SI(g1930), .SE(n8217), .CLK(n8404), .Q(
        g1934), .QN(n7969) );
  SDFFX1 DFF_1060_Q_reg ( .D(g18743), .SI(g1934), .SE(n8217), .CLK(n8404), .Q(
        g1937), .QN(n4311) );
  SDFFX1 DFF_1061_Q_reg ( .D(g18794), .SI(g1937), .SE(n8217), .CLK(n8404), .Q(
        g1890), .QN(n4297) );
  SDFFX1 DFF_1062_Q_reg ( .D(n1137), .SI(g1890), .SE(n8219), .CLK(n8406), .Q(
        g1893) );
  SDFFX1 DFF_1063_Q_reg ( .D(g1893), .SI(g1893), .SE(n8219), .CLK(n8406), .Q(
        g1903) );
  SDFFX1 DFF_1064_Q_reg ( .D(g1903), .SI(g1903), .SE(n8219), .CLK(n8406), .Q(
        g1904) );
  SDFFX1 DFF_1065_Q_reg ( .D(g1836), .SI(g1904), .SE(n8219), .CLK(n8406), .Q(
        g1944) );
  SDFFX1 DFF_1066_Q_reg ( .D(g1944), .SI(g1944), .SE(n8219), .CLK(n8406), .Q(
        g1949) );
  SDFFX1 DFF_1067_Q_reg ( .D(test_so65), .SI(g1949), .SE(n8219), .CLK(n8406), 
        .Q(g1950) );
  SDFFX1 DFF_1068_Q_reg ( .D(g1950), .SI(g1950), .SE(n8219), .CLK(n8406), .Q(
        g1951) );
  SDFFX1 DFF_1069_Q_reg ( .D(g1842), .SI(g1951), .SE(n8219), .CLK(n8406), .Q(
        test_so64) );
  SDFFX1 DFF_1070_Q_reg ( .D(test_so64), .SI(test_si65), .SE(n8219), .CLK(
        n8406), .Q(g1953) );
  SDFFX1 DFF_1071_Q_reg ( .D(g1846), .SI(g1953), .SE(n8219), .CLK(n8406), .Q(
        g1954) );
  SDFFX1 DFF_1072_Q_reg ( .D(g1954), .SI(g1954), .SE(n8219), .CLK(n8406), .Q(
        g1945) );
  SDFFX1 DFF_1073_Q_reg ( .D(g1849), .SI(g1945), .SE(n8219), .CLK(n8406), .Q(
        g1946) );
  SDFFX1 DFF_1074_Q_reg ( .D(g1946), .SI(g1946), .SE(n8220), .CLK(n8407), .Q(
        g1947) );
  SDFFX1 DFF_1075_Q_reg ( .D(g1852), .SI(g1947), .SE(n8220), .CLK(n8407), .Q(
        g1948) );
  SDFFX1 DFF_1076_Q_reg ( .D(g1948), .SI(g1948), .SE(n8220), .CLK(n8407), .Q(
        g1870) );
  SDFFX1 DFF_1077_Q_reg ( .D(g2950), .SI(g1870), .SE(n8220), .CLK(n8407), .Q(
        g8012), .QN(n4458) );
  SDFFX1 DFF_1078_Q_reg ( .D(g8012), .SI(g8012), .SE(n8220), .CLK(n8407), .Q(
        g8082), .QN(n4457) );
  SDFFX1 DFF_1079_Q_reg ( .D(g8082), .SI(g8082), .SE(n8220), .CLK(n8407), .Q(
        g1866), .QN(n4464) );
  SDFFX1 DFF_1080_Q_reg ( .D(g23097), .SI(g1866), .SE(n8220), .CLK(n8407), .Q(
        g1867) );
  SDFFX1 DFF_1081_Q_reg ( .D(g23124), .SI(g1867), .SE(n8220), .CLK(n8407), .Q(
        g1868) );
  SDFFX1 DFF_1082_Q_reg ( .D(g23137), .SI(g1868), .SE(n8220), .CLK(n8407), .Q(
        g1869) );
  SDFFX1 DFF_1083_Q_reg ( .D(g23400), .SI(g1869), .SE(n8220), .CLK(n8407), .Q(
        g1836) );
  SDFFX1 DFF_1084_Q_reg ( .D(g23413), .SI(g1836), .SE(n8220), .CLK(n8407), .Q(
        test_so65) );
  SDFFX1 DFF_1085_Q_reg ( .D(g24182), .SI(test_si66), .SE(n8220), .CLK(n8407), 
        .Q(g1842) );
  SDFFX1 DFF_1086_Q_reg ( .D(g24208), .SI(g1842), .SE(n8221), .CLK(n8408), .Q(
        g1858) );
  SDFFX1 DFF_1087_Q_reg ( .D(g24219), .SI(g1858), .SE(n8221), .CLK(n8408), .Q(
        g1859) );
  SDFFX1 DFF_1088_Q_reg ( .D(g24231), .SI(g1859), .SE(n8221), .CLK(n8408), .Q(
        g1860) );
  SDFFX1 DFF_1089_Q_reg ( .D(g23123), .SI(g1860), .SE(n8221), .CLK(n8408), .Q(
        g1861) );
  SDFFX1 DFF_1090_Q_reg ( .D(g23030), .SI(g1861), .SE(n8221), .CLK(n8408), .Q(
        g1865) );
  SDFFX1 DFF_1091_Q_reg ( .D(g23058), .SI(g1865), .SE(n8221), .CLK(n8408), .Q(
        g1845) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24218), .SI(g1845), .SE(n8221), .CLK(n8408), .Q(
        g1846) );
  SDFFX1 DFF_1093_Q_reg ( .D(g24230), .SI(g1846), .SE(n8221), .CLK(n8408), .Q(
        g1849) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24243), .SI(g1849), .SE(n8221), .CLK(n8408), .Q(
        g1852) );
  SDFFX1 DFF_1095_Q_reg ( .D(n1114), .SI(g1852), .SE(n8221), .CLK(n8408), .Q(
        g1908) );
  SDFFX1 DFF_1096_Q_reg ( .D(g1908), .SI(g1908), .SE(n8221), .CLK(n8408), .Q(
        g1915) );
  SDFFX1 DFF_1097_Q_reg ( .D(g1915), .SI(g1915), .SE(n8221), .CLK(n8408), .Q(
        g1922) );
  SDFFX1 DFF_1098_Q_reg ( .D(g13164), .SI(g1922), .SE(n8222), .CLK(n8409), .Q(
        g1923) );
  SDFFX1 DFF_1099_Q_reg ( .D(g1923), .SI(g1923), .SE(n8222), .CLK(n8409), .Q(
        test_so66), .QN(DFF_1099_n1) );
  SDFFX1 DFF_1100_Q_reg ( .D(n497), .SI(test_si67), .SE(n8222), .CLK(n8409), 
        .Q(n7971) );
  SDFFX1 DFF_1101_Q_reg ( .D(g13135), .SI(n7971), .SE(n8222), .CLK(n8409), .Q(
        g1929) );
  SDFFX1 DFF_1102_Q_reg ( .D(g1929), .SI(g1929), .SE(n8222), .CLK(n8409), .Q(
        g1880), .QN(n4545) );
  SDFFX1 DFF_1103_Q_reg ( .D(g13182), .SI(g1880), .SE(n8222), .CLK(n8409), .Q(
        g1938) );
  SDFFX1 DFF_1104_Q_reg ( .D(g1938), .SI(g1938), .SE(n8222), .CLK(n8409), .Q(
        g1939), .QN(n7750) );
  SDFFX1 DFF_1105_Q_reg ( .D(g27290), .SI(g1939), .SE(n8224), .CLK(n8411), .Q(
        g1956), .QN(n7329) );
  SDFFX1 DFF_1106_Q_reg ( .D(g27305), .SI(g1956), .SE(n8224), .CLK(n8411), .Q(
        g1957), .QN(n7331) );
  SDFFX1 DFF_1107_Q_reg ( .D(g27319), .SI(g1957), .SE(n8224), .CLK(n8411), .Q(
        g1955), .QN(n7330) );
  SDFFX1 DFF_1108_Q_reg ( .D(g27306), .SI(g1955), .SE(n8224), .CLK(n8411), .Q(
        g1959), .QN(n7341) );
  SDFFX1 DFF_1109_Q_reg ( .D(g27320), .SI(g1959), .SE(n8224), .CLK(n8411), .Q(
        g1960), .QN(n7343) );
  SDFFX1 DFF_1110_Q_reg ( .D(g27331), .SI(g1960), .SE(n8224), .CLK(n8411), .Q(
        g1958), .QN(n7342) );
  SDFFX1 DFF_1111_Q_reg ( .D(g27321), .SI(g1958), .SE(n8225), .CLK(n8412), .Q(
        g1962), .QN(n7167) );
  SDFFX1 DFF_1112_Q_reg ( .D(g27332), .SI(g1962), .SE(n8225), .CLK(n8412), .Q(
        g1963), .QN(n7169) );
  SDFFX1 DFF_1113_Q_reg ( .D(g27340), .SI(g1963), .SE(n8224), .CLK(n8411), .Q(
        g1961), .QN(n7168) );
  SDFFX1 DFF_1114_Q_reg ( .D(g27333), .SI(g1961), .SE(n8225), .CLK(n8412), .Q(
        test_so67), .QN(n8092) );
  SDFFX1 DFF_1115_Q_reg ( .D(g27341), .SI(test_si68), .SE(n8225), .CLK(n8412), 
        .Q(g1966), .QN(n7353) );
  SDFFX1 DFF_1116_Q_reg ( .D(g27346), .SI(g1966), .SE(n8223), .CLK(n8410), .Q(
        g1964), .QN(n7352) );
  SDFFX1 DFF_1117_Q_reg ( .D(g24513), .SI(g1964), .SE(n8223), .CLK(n8410), .Q(
        g1967) );
  SDFFX1 DFF_1118_Q_reg ( .D(g24524), .SI(g1967), .SE(n8223), .CLK(n8410), .Q(
        g1970) );
  SDFFX1 DFF_1119_Q_reg ( .D(g24534), .SI(g1970), .SE(n8223), .CLK(n8410), .Q(
        g1973) );
  SDFFX1 DFF_1120_Q_reg ( .D(g24525), .SI(g1973), .SE(n8224), .CLK(n8411), .Q(
        g1976) );
  SDFFX1 DFF_1121_Q_reg ( .D(g24535), .SI(g1976), .SE(n8224), .CLK(n8411), .Q(
        g1979) );
  SDFFX1 DFF_1122_Q_reg ( .D(g24545), .SI(g1979), .SE(n8224), .CLK(n8411), .Q(
        g1982) );
  SDFFX1 DFF_1123_Q_reg ( .D(g28357), .SI(g1982), .SE(n8224), .CLK(n8411), .Q(
        g1994) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28362), .SI(g1994), .SE(n8224), .CLK(n8411), .Q(
        g1997) );
  SDFFX1 DFF_1125_Q_reg ( .D(g28366), .SI(g1997), .SE(n8223), .CLK(n8410), .Q(
        g2000) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28352), .SI(g2000), .SE(n8225), .CLK(n8412), .Q(
        g1985) );
  SDFFX1 DFF_1127_Q_reg ( .D(g28356), .SI(g1985), .SE(n8225), .CLK(n8412), .Q(
        g1988) );
  SDFFX1 DFF_1128_Q_reg ( .D(g28361), .SI(g1988), .SE(n8225), .CLK(n8412), .Q(
        g1991) );
  SDFFX1 DFF_1129_Q_reg ( .D(g26559), .SI(g1991), .SE(n8225), .CLK(n8412), .Q(
        test_so68) );
  SDFFX1 DFF_1130_Q_reg ( .D(g26573), .SI(test_si69), .SE(n8223), .CLK(n8410), 
        .Q(g1874) );
  SDFFX1 DFF_1131_Q_reg ( .D(g26592), .SI(g1874), .SE(n8223), .CLK(n8410), .Q(
        g1877) );
  SDFFX1 DFF_1132_Q_reg ( .D(g1880), .SI(g1877), .SE(n8223), .CLK(n8410), .Q(
        g1886), .QN(n4493) );
  SDFFX1 DFF_1133_Q_reg ( .D(g22651), .SI(g1886), .SE(n8225), .CLK(n8412), .Q(
        n7968), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(n512), .SI(n7968), .SE(n8225), .CLK(n8412), .Q(
        g16399), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(g16399), .SI(g16399), .SE(n8225), .CLK(n8412), 
        .Q(g1905), .QN(n8038) );
  SDFFX1 DFF_1144_Q_reg ( .D(DFF_999_n1), .SI(g1905), .SE(n8225), .CLK(n8412), 
        .Q(n7967), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(DFF_1001_n1), .SI(n7967), .SE(n8226), .CLK(n8413), 
        .Q(n7966), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(DFF_1003_n1), .SI(n7966), .SE(n8226), .CLK(n8413), 
        .Q(n7965), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(DFF_1005_n1), .SI(n7965), .SE(n8226), .CLK(n8413), 
        .Q(n7964), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(DFF_1007_n1), .SI(n7964), .SE(n8226), .CLK(n8413), 
        .Q(n7963), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(DFF_1009_n1), .SI(n7963), .SE(n8226), .CLK(n8413), 
        .Q(n7962), .QN(DFF_1149_n1) );
  SDFFX1 DFF_1150_Q_reg ( .D(DFF_1011_n1), .SI(n7962), .SE(n8226), .CLK(n8413), 
        .Q(g1916), .QN(n7147) );
  SDFFX1 DFF_1151_Q_reg ( .D(DFF_1013_n1), .SI(g1916), .SE(n8226), .CLK(n8413), 
        .Q(g1917), .QN(n7146) );
  SDFFX1 DFF_1152_Q_reg ( .D(g24083), .SI(g1917), .SE(n8226), .CLK(n8413), .Q(
        test_so69), .QN(n8094) );
  SDFFX1 DFF_1153_Q_reg ( .D(n4484), .SI(test_si70), .SE(n8138), .CLK(n8325), 
        .Q(n7960), .QN(n14347) );
  SDFFX1 DFF_1155_Q_reg ( .D(g7229), .SI(g7229), .SE(n8138), .CLK(n8325), .Q(
        g7357), .QN(n4357) );
  SDFFX1 DFF_1156_Q_reg ( .D(g7357), .SI(g7357), .SE(n8138), .CLK(n8325), .Q(
        g2009), .QN(n4293) );
  SDFFX1 DFF_1157_Q_reg ( .D(g16692), .SI(g2009), .SE(n8218), .CLK(n8405), .Q(
        g2010), .QN(n7746) );
  SDFFX1 DFF_1158_Q_reg ( .D(g20353), .SI(g2010), .SE(n8218), .CLK(n8405), .Q(
        g2039), .QN(n4427) );
  SDFFX1 DFF_1159_Q_reg ( .D(g20752), .SI(g2039), .SE(n8218), .CLK(n8405), .Q(
        g2020), .QN(n4400) );
  SDFFX1 DFF_1160_Q_reg ( .D(n1214), .SI(g2020), .SE(n8218), .CLK(n8405), .Q(
        g2013), .QN(n4474) );
  SDFFX1 DFF_1161_Q_reg ( .D(g23339), .SI(g2013), .SE(n8218), .CLK(n8405), .Q(
        g2033), .QN(n4420) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24434), .SI(g2033), .SE(n8218), .CLK(n8405), .Q(
        g2026), .QN(n4410) );
  SDFFX1 DFF_1163_Q_reg ( .D(g25194), .SI(g2026), .SE(n8218), .CLK(n8405), .Q(
        g2040), .QN(n4399) );
  SDFFX1 DFF_1164_Q_reg ( .D(n1215), .SI(g2040), .SE(n8218), .CLK(n8405), .Q(
        g2052), .QN(n4409) );
  SDFFX1 DFF_1165_Q_reg ( .D(g26789), .SI(g2052), .SE(n8218), .CLK(n8405), .Q(
        g2046), .QN(n4468) );
  SDFFX1 DFF_1166_Q_reg ( .D(g27682), .SI(g2046), .SE(n8218), .CLK(n8405), .Q(
        g2059), .QN(n4473) );
  SDFFX1 DFF_1167_Q_reg ( .D(g27722), .SI(g2059), .SE(n8218), .CLK(n8405), .Q(
        test_so70), .QN(n8085) );
  SDFFX1 DFF_1168_Q_reg ( .D(g28325), .SI(test_si71), .SE(n8218), .CLK(n8405), 
        .Q(g2072), .QN(n4416) );
  SDFFX1 DFF_1169_Q_reg ( .D(g20899), .SI(g2072), .SE(n8226), .CLK(n8413), .Q(
        g2079), .QN(n7790) );
  SDFFX1 DFF_1170_Q_reg ( .D(g20915), .SI(g2079), .SE(n8226), .CLK(n8413), .Q(
        g2080), .QN(n7789) );
  SDFFX1 DFF_1171_Q_reg ( .D(g20934), .SI(g2080), .SE(n8226), .CLK(n8413), .Q(
        g2078), .QN(n7844) );
  SDFFX1 DFF_1172_Q_reg ( .D(g20916), .SI(g2078), .SE(n8226), .CLK(n8413), .Q(
        g2082), .QN(n7788) );
  SDFFX1 DFF_1173_Q_reg ( .D(g20935), .SI(g2082), .SE(n8227), .CLK(n8414), .Q(
        g2083), .QN(n7787) );
  SDFFX1 DFF_1174_Q_reg ( .D(g20953), .SI(g2083), .SE(n8227), .CLK(n8414), .Q(
        g2081), .QN(n7843) );
  SDFFX1 DFF_1175_Q_reg ( .D(g20936), .SI(g2081), .SE(n8227), .CLK(n8414), .Q(
        g2085), .QN(n7786) );
  SDFFX1 DFF_1176_Q_reg ( .D(g20954), .SI(g2085), .SE(n8227), .CLK(n8414), .Q(
        g2086), .QN(n7785) );
  SDFFX1 DFF_1177_Q_reg ( .D(g20977), .SI(g2086), .SE(n8227), .CLK(n8414), .Q(
        g2084), .QN(n7842) );
  SDFFX1 DFF_1178_Q_reg ( .D(g20955), .SI(g2084), .SE(n8228), .CLK(n8415), .Q(
        g2088), .QN(n7784) );
  SDFFX1 DFF_1179_Q_reg ( .D(g20978), .SI(g2088), .SE(n8228), .CLK(n8415), .Q(
        g2089), .QN(n7783) );
  SDFFX1 DFF_1180_Q_reg ( .D(g20999), .SI(g2089), .SE(n8228), .CLK(n8415), .Q(
        g2087), .QN(n7841) );
  SDFFX1 DFF_1181_Q_reg ( .D(g20979), .SI(g2087), .SE(n8228), .CLK(n8415), .Q(
        g2091), .QN(n7782) );
  SDFFX1 DFF_1182_Q_reg ( .D(g21000), .SI(g2091), .SE(n8228), .CLK(n8415), .Q(
        test_so71), .QN(n8121) );
  SDFFX1 DFF_1183_Q_reg ( .D(g21019), .SI(test_si72), .SE(n8228), .CLK(n8415), 
        .Q(g2090), .QN(n7840) );
  SDFFX1 DFF_1184_Q_reg ( .D(g21001), .SI(g2090), .SE(n8228), .CLK(n8415), .Q(
        g2094), .QN(n7781) );
  SDFFX1 DFF_1185_Q_reg ( .D(g21020), .SI(g2094), .SE(n8228), .CLK(n8415), .Q(
        g2095), .QN(n7780) );
  SDFFX1 DFF_1186_Q_reg ( .D(g21039), .SI(g2095), .SE(n8228), .CLK(n8415), .Q(
        g2093), .QN(n7839) );
  SDFFX1 DFF_1187_Q_reg ( .D(g21021), .SI(g2093), .SE(n8228), .CLK(n8415), .Q(
        g2097), .QN(n7779) );
  SDFFX1 DFF_1188_Q_reg ( .D(g21040), .SI(g2097), .SE(n8228), .CLK(n8415), .Q(
        g2098), .QN(n7778) );
  SDFFX1 DFF_1189_Q_reg ( .D(g21054), .SI(g2098), .SE(n8228), .CLK(n8415), .Q(
        g2096), .QN(n7838) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21041), .SI(g2096), .SE(n8229), .CLK(n8416), .Q(
        g2100), .QN(n7777) );
  SDFFX1 DFF_1191_Q_reg ( .D(g21055), .SI(g2100), .SE(n8229), .CLK(n8416), .Q(
        g2101), .QN(n7776) );
  SDFFX1 DFF_1192_Q_reg ( .D(g21071), .SI(g2101), .SE(n8229), .CLK(n8416), .Q(
        g2099), .QN(n7837) );
  SDFFX1 DFF_1193_Q_reg ( .D(g21056), .SI(g2099), .SE(n8229), .CLK(n8416), .Q(
        g2103), .QN(n7775) );
  SDFFX1 DFF_1194_Q_reg ( .D(g21072), .SI(g2103), .SE(n8229), .CLK(n8416), .Q(
        g2104), .QN(n7774) );
  SDFFX1 DFF_1195_Q_reg ( .D(g21080), .SI(g2104), .SE(n8229), .CLK(n8416), .Q(
        g2102), .QN(n7836) );
  SDFFX1 DFF_1196_Q_reg ( .D(g20900), .SI(g2102), .SE(n8229), .CLK(n8416), .Q(
        g2106), .QN(n7773) );
  SDFFX1 DFF_1197_Q_reg ( .D(g20917), .SI(g2106), .SE(n8229), .CLK(n8416), .Q(
        test_so72), .QN(n8122) );
  SDFFX1 DFF_1198_Q_reg ( .D(g20937), .SI(test_si73), .SE(n8227), .CLK(n8414), 
        .Q(g2105), .QN(n7835) );
  SDFFX1 DFF_1199_Q_reg ( .D(g20980), .SI(g2105), .SE(n8227), .CLK(n8414), .Q(
        g2109), .QN(n8028) );
  SDFFX1 DFF_1200_Q_reg ( .D(g21002), .SI(g2109), .SE(n8227), .CLK(n8414), .Q(
        g2110), .QN(n7558) );
  SDFFX1 DFF_1201_Q_reg ( .D(g21022), .SI(g2110), .SE(n8227), .CLK(n8414), .Q(
        g2108) );
  SDFFX1 DFF_1202_Q_reg ( .D(g21003), .SI(g2108), .SE(n8227), .CLK(n8414), .Q(
        g2112), .QN(n7564) );
  SDFFX1 DFF_1203_Q_reg ( .D(g21023), .SI(g2112), .SE(n8227), .CLK(n8414), .Q(
        g2113), .QN(n7557) );
  SDFFX1 DFF_1204_Q_reg ( .D(g21042), .SI(g2113), .SE(n8227), .CLK(n8414), .Q(
        g2111), .QN(n7615) );
  SDFFX1 DFF_1205_Q_reg ( .D(g25268), .SI(g2111), .SE(n8229), .CLK(n8416), .Q(
        g2115), .QN(n7493) );
  SDFFX1 DFF_1206_Q_reg ( .D(g25271), .SI(g2115), .SE(n8229), .CLK(n8416), .Q(
        g2116), .QN(n7492) );
  SDFFX1 DFF_1207_Q_reg ( .D(g25279), .SI(g2116), .SE(n8229), .CLK(n8416), .Q(
        g2114), .QN(n7499) );
  SDFFX1 DFF_1208_Q_reg ( .D(g22249), .SI(g2114), .SE(n8229), .CLK(n8416), .Q(
        g2118), .QN(n7866) );
  SDFFX1 DFF_1209_Q_reg ( .D(n1186), .SI(g2118), .SE(n8230), .CLK(n8417), .Q(
        g2119), .QN(n7954) );
  SDFFX1 DFF_1210_Q_reg ( .D(g22280), .SI(g2119), .SE(n8230), .CLK(n8417), .Q(
        g2117), .QN(n7957) );
  SDFFX1 DFF_1211_Q_reg ( .D(g2950), .SI(g2117), .SE(n8230), .CLK(n8417), .Q(
        g6837), .QN(n4324) );
  SDFFX1 DFF_1212_Q_reg ( .D(g6837), .SI(g6837), .SE(n8230), .CLK(n8417), .Q(
        test_so73), .QN(n8070) );
  SDFFX1 DFF_1213_Q_reg ( .D(test_so73), .SI(test_si74), .SE(n8230), .CLK(
        n8417), .Q(g2241), .QN(n4367) );
  SDFFX1 DFF_1214_Q_reg ( .D(g22170), .SI(g2241), .SE(n8230), .CLK(n8417), .Q(
        g2206), .QN(n7883) );
  SDFFX1 DFF_1215_Q_reg ( .D(g22182), .SI(g2206), .SE(n8234), .CLK(n8421), .Q(
        g2207), .QN(n7882) );
  SDFFX1 DFF_1216_Q_reg ( .D(g22192), .SI(g2207), .SE(n8234), .CLK(n8421), .Q(
        g2205), .QN(n7520) );
  SDFFX1 DFF_1217_Q_reg ( .D(g22183), .SI(g2205), .SE(n8230), .CLK(n8417), .Q(
        g2209), .QN(n7881) );
  SDFFX1 DFF_1218_Q_reg ( .D(g22193), .SI(g2209), .SE(n8234), .CLK(n8421), .Q(
        g2210), .QN(n7880) );
  SDFFX1 DFF_1219_Q_reg ( .D(g22200), .SI(g2210), .SE(n8235), .CLK(n8422), .Q(
        g2208), .QN(n7519) );
  SDFFX1 DFF_1220_Q_reg ( .D(g22045), .SI(g2208), .SE(n8235), .CLK(n8422), .Q(
        g2218), .QN(n7879) );
  SDFFX1 DFF_1221_Q_reg ( .D(g22060), .SI(g2218), .SE(n8235), .CLK(n8422), .Q(
        g2219), .QN(n7878) );
  SDFFX1 DFF_1222_Q_reg ( .D(g22076), .SI(g2219), .SE(n8235), .CLK(n8422), .Q(
        g2217), .QN(n7518) );
  SDFFX1 DFF_1223_Q_reg ( .D(g22061), .SI(g2217), .SE(n8235), .CLK(n8422), .Q(
        g2221), .QN(n7877) );
  SDFFX1 DFF_1224_Q_reg ( .D(g22077), .SI(g2221), .SE(n8235), .CLK(n8422), .Q(
        g2222), .QN(n7876) );
  SDFFX1 DFF_1225_Q_reg ( .D(g22097), .SI(g2222), .SE(n8235), .CLK(n8422), .Q(
        g2220), .QN(n7517) );
  SDFFX1 DFF_1226_Q_reg ( .D(g22078), .SI(g2220), .SE(n8235), .CLK(n8422), .Q(
        g2224), .QN(n7875) );
  SDFFX1 DFF_1227_Q_reg ( .D(g22098), .SI(g2224), .SE(n8235), .CLK(n8422), .Q(
        test_so74), .QN(n8118) );
  SDFFX1 DFF_1228_Q_reg ( .D(g22115), .SI(test_si75), .SE(n8232), .CLK(n8419), 
        .Q(g2223), .QN(n7516) );
  SDFFX1 DFF_1229_Q_reg ( .D(g22099), .SI(g2223), .SE(n8232), .CLK(n8419), .Q(
        g2227), .QN(n7874) );
  SDFFX1 DFF_1230_Q_reg ( .D(g22116), .SI(g2227), .SE(n8233), .CLK(n8420), .Q(
        g2228), .QN(n7873) );
  SDFFX1 DFF_1231_Q_reg ( .D(g22138), .SI(g2228), .SE(n8233), .CLK(n8420), .Q(
        g2226), .QN(n7515) );
  SDFFX1 DFF_1232_Q_reg ( .D(g22117), .SI(g2226), .SE(n8233), .CLK(n8420), .Q(
        g2230), .QN(n7872) );
  SDFFX1 DFF_1233_Q_reg ( .D(g22139), .SI(g2230), .SE(n8233), .CLK(n8420), .Q(
        g2231), .QN(n7871) );
  SDFFX1 DFF_1234_Q_reg ( .D(g22153), .SI(g2231), .SE(n8234), .CLK(n8421), .Q(
        g2229), .QN(n7514) );
  SDFFX1 DFF_1235_Q_reg ( .D(g22140), .SI(g2229), .SE(n8234), .CLK(n8421), .Q(
        g2233), .QN(n7870) );
  SDFFX1 DFF_1236_Q_reg ( .D(g22154), .SI(g2233), .SE(n8234), .CLK(n8421), .Q(
        g2234), .QN(n7869) );
  SDFFX1 DFF_1237_Q_reg ( .D(g22171), .SI(g2234), .SE(n8234), .CLK(n8421), .Q(
        g2232), .QN(n7513) );
  SDFFX1 DFF_1238_Q_reg ( .D(g22155), .SI(g2232), .SE(n8234), .CLK(n8421), .Q(
        g2236), .QN(n7504) );
  SDFFX1 DFF_1239_Q_reg ( .D(g22172), .SI(g2236), .SE(n8234), .CLK(n8421), .Q(
        g2237), .QN(n7503) );
  SDFFX1 DFF_1240_Q_reg ( .D(g22184), .SI(g2237), .SE(n8234), .CLK(n8421), .Q(
        g2235), .QN(n7502) );
  SDFFX1 DFF_1241_Q_reg ( .D(g22173), .SI(g2235), .SE(n8234), .CLK(n8421), .Q(
        g2239), .QN(n7512) );
  SDFFX1 DFF_1242_Q_reg ( .D(g22185), .SI(g2239), .SE(n8234), .CLK(n8421), .Q(
        test_so75), .QN(n8117) );
  SDFFX1 DFF_1243_Q_reg ( .D(g22194), .SI(test_si76), .SE(n8232), .CLK(n8419), 
        .Q(g2238), .QN(n7511) );
  SDFFX1 DFF_1244_Q_reg ( .D(g25227), .SI(g2238), .SE(n8232), .CLK(n8419), .Q(
        g2245), .QN(n7578) );
  SDFFX1 DFF_1245_Q_reg ( .D(g25236), .SI(g2245), .SE(n8232), .CLK(n8419), .Q(
        g2246), .QN(n7577) );
  SDFFX1 DFF_1246_Q_reg ( .D(g25245), .SI(g2246), .SE(n8232), .CLK(n8419), .Q(
        g2244), .QN(n7576) );
  SDFFX1 DFF_1247_Q_reg ( .D(g25237), .SI(g2244), .SE(n8233), .CLK(n8420), .Q(
        g2248), .QN(n7575) );
  SDFFX1 DFF_1248_Q_reg ( .D(g25246), .SI(g2248), .SE(n8233), .CLK(n8420), .Q(
        g2249), .QN(n7574) );
  SDFFX1 DFF_1249_Q_reg ( .D(g25251), .SI(g2249), .SE(n8233), .CLK(n8420), .Q(
        g2247), .QN(n7573) );
  SDFFX1 DFF_1250_Q_reg ( .D(g25247), .SI(g2247), .SE(n8233), .CLK(n8420), .Q(
        g2251), .QN(n7572) );
  SDFFX1 DFF_1251_Q_reg ( .D(g25252), .SI(g2251), .SE(n8233), .CLK(n8420), .Q(
        g2252), .QN(n7571) );
  SDFFX1 DFF_1252_Q_reg ( .D(g25256), .SI(g2252), .SE(n8233), .CLK(n8420), .Q(
        g2250), .QN(n7570) );
  SDFFX1 DFF_1253_Q_reg ( .D(g25253), .SI(g2250), .SE(n8233), .CLK(n8420), .Q(
        g2254), .QN(n7569) );
  SDFFX1 DFF_1254_Q_reg ( .D(g25257), .SI(g2254), .SE(n8233), .CLK(n8420), .Q(
        g2255), .QN(n7568) );
  SDFFX1 DFF_1255_Q_reg ( .D(g25259), .SI(g2255), .SE(n8135), .CLK(n8322), .Q(
        g2253), .QN(n7567) );
  SDFFX1 DFF_1256_Q_reg ( .D(g30289), .SI(g2253), .SE(n8243), .CLK(n8430), .Q(
        g2261) );
  SDFFX1 DFF_1257_Q_reg ( .D(g30296), .SI(g2261), .SE(n8243), .CLK(n8430), .Q(
        test_so76) );
  SDFFX1 DFF_1258_Q_reg ( .D(g30300), .SI(test_si77), .SE(n8243), .CLK(n8430), 
        .Q(g2267) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30660), .SI(g2267), .SE(n8243), .CLK(n8430), .Q(
        g2306) );
  SDFFX1 DFF_1260_Q_reg ( .D(g30666), .SI(g2306), .SE(n8243), .CLK(n8430), .Q(
        g2309) );
  SDFFX1 DFF_1261_Q_reg ( .D(g30672), .SI(g2309), .SE(n8243), .CLK(n8430), .Q(
        g2312) );
  SDFFX1 DFF_1262_Q_reg ( .D(g30690), .SI(g2312), .SE(n8243), .CLK(n8430), .Q(
        g2270) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30693), .SI(g2270), .SE(n8244), .CLK(n8431), .Q(
        g2273) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30695), .SI(g2273), .SE(n8235), .CLK(n8422), .Q(
        g2276) );
  SDFFX1 DFF_1265_Q_reg ( .D(g30667), .SI(g2276), .SE(n8235), .CLK(n8422), .Q(
        g2315) );
  SDFFX1 DFF_1266_Q_reg ( .D(g30673), .SI(g2315), .SE(n8235), .CLK(n8422), .Q(
        g2318) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30679), .SI(g2318), .SE(n8236), .CLK(n8423), .Q(
        g2321) );
  SDFFX1 DFF_1268_Q_reg ( .D(g30301), .SI(g2321), .SE(n8236), .CLK(n8423), .Q(
        g2279) );
  SDFFX1 DFF_1269_Q_reg ( .D(g30303), .SI(g2279), .SE(n8236), .CLK(n8423), .Q(
        g2282) );
  SDFFX1 DFF_1270_Q_reg ( .D(g30304), .SI(g2282), .SE(n8236), .CLK(n8423), .Q(
        g2285) );
  SDFFX1 DFF_1271_Q_reg ( .D(g30274), .SI(g2285), .SE(n8236), .CLK(n8423), .Q(
        g2324) );
  SDFFX1 DFF_1272_Q_reg ( .D(g30282), .SI(g2324), .SE(n8236), .CLK(n8423), .Q(
        test_so77) );
  SDFFX1 DFF_1273_Q_reg ( .D(g30290), .SI(test_si78), .SE(n8236), .CLK(n8423), 
        .Q(g2330) );
  SDFFX1 DFF_1274_Q_reg ( .D(g30253), .SI(g2330), .SE(n8242), .CLK(n8429), .Q(
        g2288) );
  SDFFX1 DFF_1275_Q_reg ( .D(g30256), .SI(g2288), .SE(n8242), .CLK(n8429), .Q(
        g2291) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30260), .SI(g2291), .SE(n8242), .CLK(n8429), .Q(
        g2294) );
  SDFFX1 DFF_1277_Q_reg ( .D(g30283), .SI(g2294), .SE(n8243), .CLK(n8430), .Q(
        g2333) );
  SDFFX1 DFF_1278_Q_reg ( .D(g30291), .SI(g2333), .SE(n8243), .CLK(n8430), .Q(
        g2336) );
  SDFFX1 DFF_1279_Q_reg ( .D(g30297), .SI(g2336), .SE(n8243), .CLK(n8430), .Q(
        g2339) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30652), .SI(g2339), .SE(n8243), .CLK(n8430), .Q(
        g2297) );
  SDFFX1 DFF_1281_Q_reg ( .D(g30659), .SI(g2297), .SE(n8243), .CLK(n8430), .Q(
        g2300) );
  SDFFX1 DFF_1282_Q_reg ( .D(g30665), .SI(g2300), .SE(n8236), .CLK(n8423), .Q(
        g2303) );
  SDFFX1 DFF_1283_Q_reg ( .D(g30686), .SI(g2303), .SE(n8236), .CLK(n8423), .Q(
        g2342) );
  SDFFX1 DFF_1284_Q_reg ( .D(g30691), .SI(g2342), .SE(n8236), .CLK(n8423), .Q(
        g2345) );
  SDFFX1 DFF_1285_Q_reg ( .D(g30694), .SI(g2345), .SE(n8230), .CLK(n8417), .Q(
        g2348) );
  SDFFX1 DFF_1286_Q_reg ( .D(g25067), .SI(g2348), .SE(n8230), .CLK(n8417), .Q(
        g2160), .QN(n7690) );
  SDFFX1 DFF_1287_Q_reg ( .D(g25940), .SI(g2160), .SE(n8230), .CLK(n8417), .Q(
        test_so78) );
  SDFFX1 DFF_1288_Q_reg ( .D(g26532), .SI(test_si79), .SE(n8231), .CLK(n8418), 
        .Q(g2151), .QN(n7689) );
  SDFFX1 DFF_1289_Q_reg ( .D(g27131), .SI(g2151), .SE(n8231), .CLK(n8418), .Q(
        g2147), .QN(n8053) );
  SDFFX1 DFF_1290_Q_reg ( .D(g27621), .SI(g2147), .SE(n8231), .CLK(n8418), .Q(
        g2142), .QN(n7688) );
  SDFFX1 DFF_1291_Q_reg ( .D(g28148), .SI(g2142), .SE(n8231), .CLK(n8418), .Q(
        g2138), .QN(n8069) );
  SDFFX1 DFF_1292_Q_reg ( .D(g28637), .SI(g2138), .SE(n8231), .CLK(n8418), .Q(
        g2133), .QN(n7687) );
  SDFFX1 DFF_1293_Q_reg ( .D(g29112), .SI(g2133), .SE(n8231), .CLK(n8418), .Q(
        g2129), .QN(n8050) );
  SDFFX1 DFF_1294_Q_reg ( .D(g29357), .SI(g2129), .SE(n8231), .CLK(n8418), .Q(
        g2124), .QN(n7322) );
  SDFFX1 DFF_1295_Q_reg ( .D(g29582), .SI(g2124), .SE(n8231), .CLK(n8418), .Q(
        g2120), .QN(n7161) );
  SDFFX1 DFF_1296_Q_reg ( .D(n19), .SI(g2120), .SE(n8231), .CLK(n8418), .Q(
        g2256) );
  SDFFX1 DFF_1297_Q_reg ( .D(g2256), .SI(g2256), .SE(n8231), .CLK(n8418), .Q(
        g5637) );
  SDFFX1 DFF_1298_Q_reg ( .D(g5637), .SI(g5637), .SE(n8231), .CLK(n8418), .Q(
        g2257), .QN(n7706) );
  SDFFX1 DFF_1299_Q_reg ( .D(g2950), .SI(g2257), .SE(n8231), .CLK(n8418), .Q(
        g5555), .QN(n4516) );
  SDFFX1 DFF_1302_Q_reg ( .D(g5637), .SI(n4606), .SE(n8232), .CLK(n8419), .Q(
        test_so79), .QN(n8075) );
  SDFFX1 DFF_1303_Q_reg ( .D(g27276), .SI(test_si80), .SE(n8241), .CLK(n8428), 
        .Q(g2429), .QN(n7645) );
  SDFFX1 DFF_1304_Q_reg ( .D(g27291), .SI(g2429), .SE(n8241), .CLK(n8428), .Q(
        g2418), .QN(n7644) );
  SDFFX1 DFF_1305_Q_reg ( .D(g27307), .SI(g2418), .SE(n8242), .CLK(n8429), .Q(
        g2421), .QN(n7643) );
  SDFFX1 DFF_1306_Q_reg ( .D(g27292), .SI(g2421), .SE(n8242), .CLK(n8429), .Q(
        g2444), .QN(n7622) );
  SDFFX1 DFF_1307_Q_reg ( .D(g27308), .SI(g2444), .SE(n8242), .CLK(n8429), .Q(
        g2433), .QN(n7621) );
  SDFFX1 DFF_1308_Q_reg ( .D(g27322), .SI(g2433), .SE(n8242), .CLK(n8429), .Q(
        g2436), .QN(n7620) );
  SDFFX1 DFF_1309_Q_reg ( .D(g27309), .SI(g2436), .SE(n8242), .CLK(n8429), .Q(
        g2459), .QN(n7371) );
  SDFFX1 DFF_1310_Q_reg ( .D(g27323), .SI(g2459), .SE(n8242), .CLK(n8429), .Q(
        g2448), .QN(n7373) );
  SDFFX1 DFF_1311_Q_reg ( .D(g27334), .SI(g2448), .SE(n8242), .CLK(n8429), .Q(
        g2451), .QN(n7372) );
  SDFFX1 DFF_1312_Q_reg ( .D(g27324), .SI(g2451), .SE(n8242), .CLK(n8429), .Q(
        g2473), .QN(n7634) );
  SDFFX1 DFF_1313_Q_reg ( .D(g27335), .SI(g2473), .SE(n8242), .CLK(n8429), .Q(
        g2463), .QN(n7633) );
  SDFFX1 DFF_1314_Q_reg ( .D(g27342), .SI(g2463), .SE(n8237), .CLK(n8424), .Q(
        g2466), .QN(n7632) );
  SDFFX1 DFF_1315_Q_reg ( .D(g28763), .SI(g2466), .SE(n8237), .CLK(n8424), .Q(
        g2483) );
  SDFFX1 DFF_1316_Q_reg ( .D(g28773), .SI(g2483), .SE(n8241), .CLK(n8428), .Q(
        g2486) );
  SDFFX1 DFF_1317_Q_reg ( .D(g28782), .SI(g2486), .SE(n8241), .CLK(n8428), .Q(
        test_so80) );
  SDFFX1 DFF_1318_Q_reg ( .D(g29213), .SI(test_si81), .SE(n8237), .CLK(n8424), 
        .Q(g2492) );
  SDFFX1 DFF_1319_Q_reg ( .D(g29221), .SI(g2492), .SE(n8237), .CLK(n8424), .Q(
        g2495) );
  SDFFX1 DFF_1320_Q_reg ( .D(g29226), .SI(g2495), .SE(n8237), .CLK(n8424), .Q(
        g2498) );
  SDFFX1 DFF_1321_Q_reg ( .D(g28774), .SI(g2498), .SE(n8240), .CLK(n8427), .Q(
        g2502), .QN(n7666) );
  SDFFX1 DFF_1322_Q_reg ( .D(g28783), .SI(g2502), .SE(n8241), .CLK(n8428), .Q(
        g2503), .QN(n7656) );
  SDFFX1 DFF_1323_Q_reg ( .D(g28788), .SI(g2503), .SE(n8241), .CLK(n8428), .Q(
        g2501), .QN(n7665) );
  SDFFX1 DFF_1324_Q_reg ( .D(g26817), .SI(g2501), .SE(n8241), .CLK(n8428), .Q(
        g2504) );
  SDFFX1 DFF_1325_Q_reg ( .D(g26822), .SI(g2504), .SE(n8241), .CLK(n8428), .Q(
        g2507) );
  SDFFX1 DFF_1326_Q_reg ( .D(g26825), .SI(g2507), .SE(n8241), .CLK(n8428), .Q(
        g2510) );
  SDFFX1 DFF_1327_Q_reg ( .D(g26823), .SI(g2510), .SE(n8241), .CLK(n8428), .Q(
        g2513) );
  SDFFX1 DFF_1328_Q_reg ( .D(g26826), .SI(g2513), .SE(n8241), .CLK(n8428), .Q(
        g2516) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26827), .SI(g2516), .SE(n8135), .CLK(n8322), .Q(
        g2519) );
  SDFFX1 DFF_1330_Q_reg ( .D(g27767), .SI(g2519), .SE(n8260), .CLK(n8447), .Q(
        g2523), .QN(n7664) );
  SDFFX1 DFF_1331_Q_reg ( .D(g27769), .SI(g2523), .SE(n8260), .CLK(n8447), .Q(
        g2524), .QN(n7655) );
  SDFFX1 DFF_1332_Q_reg ( .D(g27771), .SI(g2524), .SE(n8135), .CLK(n8322), .Q(
        test_so81), .QN(n8110) );
  SDFFX1 DFF_1333_Q_reg ( .D(g29618), .SI(test_si82), .SE(n8236), .CLK(n8423), 
        .Q(g2387), .QN(n7270) );
  SDFFX1 DFF_1334_Q_reg ( .D(g29621), .SI(g2387), .SE(n8236), .CLK(n8423), .Q(
        g2388), .QN(n7258) );
  SDFFX1 DFF_1335_Q_reg ( .D(g29623), .SI(g2388), .SE(n8237), .CLK(n8424), .Q(
        g2389), .QN(n7269) );
  SDFFX1 DFF_1336_Q_reg ( .D(g30707), .SI(g2389), .SE(n8237), .CLK(n8424), .Q(
        g2390), .QN(n7268) );
  SDFFX1 DFF_1337_Q_reg ( .D(g30709), .SI(g2390), .SE(n8230), .CLK(n8417), .Q(
        g2391), .QN(n7257) );
  SDFFX1 DFF_1338_Q_reg ( .D(g30566), .SI(g2391), .SE(n8232), .CLK(n8419), .Q(
        g2392), .QN(n7267) );
  SDFFX1 DFF_1339_Q_reg ( .D(g30505), .SI(g2392), .SE(n8230), .CLK(n8417), .Q(
        g2393), .QN(n7266) );
  SDFFX1 DFF_1340_Q_reg ( .D(g30341), .SI(g2393), .SE(n8232), .CLK(n8419), .Q(
        g2394), .QN(n7256) );
  SDFFX1 DFF_1341_Q_reg ( .D(g30356), .SI(g2394), .SE(n8232), .CLK(n8419), .Q(
        g2395), .QN(n7265) );
  SDFFX1 DFF_1342_Q_reg ( .D(g29182), .SI(g2395), .SE(n8244), .CLK(n8431), .Q(
        g2397), .QN(n7314) );
  SDFFX1 DFF_1343_Q_reg ( .D(g29185), .SI(g2397), .SE(n8244), .CLK(n8431), .Q(
        g2398), .QN(n7310) );
  SDFFX1 DFF_1344_Q_reg ( .D(g29187), .SI(g2398), .SE(n8244), .CLK(n8431), .Q(
        g2396), .QN(n7313) );
  SDFFX1 DFF_1345_Q_reg ( .D(g26672), .SI(g2396), .SE(n8244), .CLK(n8431), .Q(
        g2478), .QN(n7663) );
  SDFFX1 DFF_1346_Q_reg ( .D(g26676), .SI(g2478), .SE(n8244), .CLK(n8431), .Q(
        g2479), .QN(n7654) );
  SDFFX1 DFF_1347_Q_reg ( .D(g26025), .SI(g2479), .SE(n8244), .CLK(n8431), .Q(
        test_so82), .QN(n8116) );
  SDFFX1 DFF_1348_Q_reg ( .D(n4287), .SI(test_si83), .SE(n8143), .CLK(n8330), 
        .Q(g2525) );
  SDFFX1 DFF_1349_Q_reg ( .D(g2525), .SI(g2525), .SE(n8143), .CLK(n8330), .Q(
        n7946), .QN(DFF_1349_n1) );
  SDFFX1 DFF_1350_Q_reg ( .D(n4563), .SI(n7946), .SE(n8143), .CLK(n8330), .Q(
        g2527) );
  SDFFX1 DFF_1351_Q_reg ( .D(g2527), .SI(g2527), .SE(n8143), .CLK(n8330), .Q(
        n7945), .QN(DFF_1351_n1) );
  SDFFX1 DFF_1352_Q_reg ( .D(n4555), .SI(n7945), .SE(n8143), .CLK(n8330), .Q(
        g2529) );
  SDFFX1 DFF_1353_Q_reg ( .D(g2529), .SI(g2529), .SE(n8143), .CLK(n8330), .Q(
        n7944), .QN(DFF_1353_n1) );
  SDFFX1 DFF_1354_Q_reg ( .D(n4325), .SI(n7944), .SE(n8143), .CLK(n8330), .Q(
        g2355) );
  SDFFX1 DFF_1355_Q_reg ( .D(g2355), .SI(g2355), .SE(n8143), .CLK(n8330), .Q(
        n7943), .QN(DFF_1355_n1) );
  SDFFX1 DFF_1356_Q_reg ( .D(n4389), .SI(n7943), .SE(n8143), .CLK(n8330), .Q(
        g2357) );
  SDFFX1 DFF_1357_Q_reg ( .D(g2357), .SI(g2357), .SE(n8143), .CLK(n8330), .Q(
        n7942), .QN(DFF_1357_n1) );
  SDFFX1 DFF_1358_Q_reg ( .D(n4319), .SI(n7942), .SE(n8143), .CLK(n8330), .Q(
        g2359) );
  SDFFX1 DFF_1359_Q_reg ( .D(g2359), .SI(g2359), .SE(n8143), .CLK(n8330), .Q(
        n7941), .QN(DFF_1359_n1) );
  SDFFX1 DFF_1360_Q_reg ( .D(n4373), .SI(n7941), .SE(n8144), .CLK(n8331), .Q(
        g2361) );
  SDFFX1 DFF_1361_Q_reg ( .D(g2361), .SI(g2361), .SE(n8144), .CLK(n8331), .Q(
        n7940), .QN(DFF_1361_n1) );
  SDFFX1 DFF_1362_Q_reg ( .D(n4377), .SI(n7940), .SE(n8144), .CLK(n8331), .Q(
        test_so83) );
  SDFFX1 DFF_1363_Q_reg ( .D(test_so83), .SI(test_si84), .SE(n8144), .CLK(
        n8331), .Q(n7938), .QN(DFF_1363_n1) );
  SDFFX1 DFF_1364_Q_reg ( .D(g2878), .SI(n7938), .SE(n8164), .CLK(n8351), .Q(
        g2365) );
  SDFFX1 DFF_1365_Q_reg ( .D(g2365), .SI(g2365), .SE(n8164), .CLK(n8351), .Q(
        n7937), .QN(n4483) );
  SDFFX1 DFF_1366_Q_reg ( .D(n4285), .SI(n7937), .SE(n8241), .CLK(n8428), .Q(
        g2374), .QN(n4487) );
  SDFFX1 DFF_1367_Q_reg ( .D(g30055), .SI(g2374), .SE(n8246), .CLK(n8433), .Q(
        g2380) );
  SDFFX1 DFF_1378_Q_reg ( .D(n4275), .SI(g2380), .SE(n8244), .CLK(n8431), .Q(
        n7936), .QN(DFF_1378_n1) );
  SDFFX1 DFF_1379_Q_reg ( .D(g2429), .SI(n7936), .SE(n8244), .CLK(n8431), .Q(
        g2417) );
  SDFFX1 DFF_1380_Q_reg ( .D(g2417), .SI(g2417), .SE(n8244), .CLK(n8431), .Q(
        g2424) );
  SDFFX1 DFF_1381_Q_reg ( .D(g2418), .SI(g2424), .SE(n8244), .CLK(n8431), .Q(
        g2425) );
  SDFFX1 DFF_1382_Q_reg ( .D(g2425), .SI(g2425), .SE(n8244), .CLK(n8431), .Q(
        g2426) );
  SDFFX1 DFF_1383_Q_reg ( .D(g2421), .SI(g2426), .SE(n8245), .CLK(n8432), .Q(
        g2427) );
  SDFFX1 DFF_1384_Q_reg ( .D(g2427), .SI(g2427), .SE(n8245), .CLK(n8432), .Q(
        g2428) );
  SDFFX1 DFF_1385_Q_reg ( .D(g2444), .SI(g2428), .SE(n8245), .CLK(n8432), .Q(
        g2432) );
  SDFFX1 DFF_1386_Q_reg ( .D(g2432), .SI(g2432), .SE(n8245), .CLK(n8432), .Q(
        g2439) );
  SDFFX1 DFF_1387_Q_reg ( .D(g2433), .SI(g2439), .SE(n8245), .CLK(n8432), .Q(
        test_so84) );
  SDFFX1 DFF_1388_Q_reg ( .D(test_so84), .SI(test_si85), .SE(n8245), .CLK(
        n8432), .Q(g2441) );
  SDFFX1 DFF_1389_Q_reg ( .D(g2436), .SI(g2441), .SE(n8245), .CLK(n8432), .Q(
        g2442) );
  SDFFX1 DFF_1390_Q_reg ( .D(g2442), .SI(g2442), .SE(n8245), .CLK(n8432), .Q(
        g2443) );
  SDFFX1 DFF_1391_Q_reg ( .D(g2459), .SI(g2443), .SE(n8245), .CLK(n8432), .Q(
        g2447) );
  SDFFX1 DFF_1392_Q_reg ( .D(g2447), .SI(g2447), .SE(n8245), .CLK(n8432), .Q(
        g2454) );
  SDFFX1 DFF_1393_Q_reg ( .D(g2448), .SI(g2454), .SE(n8245), .CLK(n8432), .Q(
        g2455) );
  SDFFX1 DFF_1394_Q_reg ( .D(g2455), .SI(g2455), .SE(n8245), .CLK(n8432), .Q(
        g2456) );
  SDFFX1 DFF_1395_Q_reg ( .D(g2451), .SI(g2456), .SE(n8246), .CLK(n8433), .Q(
        g2457) );
  SDFFX1 DFF_1396_Q_reg ( .D(g2457), .SI(g2457), .SE(n8246), .CLK(n8433), .Q(
        g2458) );
  SDFFX1 DFF_1397_Q_reg ( .D(g2473), .SI(g2458), .SE(n8246), .CLK(n8433), .Q(
        g2462) );
  SDFFX1 DFF_1398_Q_reg ( .D(g2462), .SI(g2462), .SE(n8246), .CLK(n8433), .Q(
        g2469) );
  SDFFX1 DFF_1399_Q_reg ( .D(g2463), .SI(g2469), .SE(n8246), .CLK(n8433), .Q(
        g2470) );
  SDFFX1 DFF_1400_Q_reg ( .D(g2470), .SI(g2470), .SE(n8246), .CLK(n8433), .Q(
        g2471) );
  SDFFX1 DFF_1401_Q_reg ( .D(g2466), .SI(g2471), .SE(n8246), .CLK(n8433), .Q(
        g2472) );
  SDFFX1 DFF_1402_Q_reg ( .D(g2472), .SI(g2472), .SE(n8246), .CLK(n8433), .Q(
        test_so85) );
  SDFFX1 DFF_1403_Q_reg ( .D(n4598), .SI(test_si86), .SE(n8130), .CLK(n8317), 
        .Q(g5747) );
  SDFFX1 DFF_1404_Q_reg ( .D(g5747), .SI(g5747), .SE(n8130), .CLK(n8317), .Q(
        g5796) );
  SDFFX1 DFF_1405_Q_reg ( .D(g5796), .SI(g5796), .SE(n8130), .CLK(n8317), .Q(
        g2412) );
  SDFFX1 DFF_1406_Q_reg ( .D(n4598), .SI(g2412), .SE(n8130), .CLK(n8317), .Q(
        g7302), .QN(n4314) );
  SDFFX1 DFF_1407_Q_reg ( .D(g7302), .SI(g7302), .SE(n8130), .CLK(n8317), .Q(
        g7390), .QN(n4370) );
  SDFFX1 DFF_1408_Q_reg ( .D(g7390), .SI(g7390), .SE(n8130), .CLK(n8317), .Q(
        g2624), .QN(n4299) );
  SDFFX1 DFF_1409_Q_reg ( .D(n1427), .SI(g2624), .SE(n8167), .CLK(n8354), .Q(
        g2628), .QN(n7961) );
  SDFFX1 DFF_1410_Q_reg ( .D(g18780), .SI(g2628), .SE(n8167), .CLK(n8354), .Q(
        g2631), .QN(n4352) );
  SDFFX1 DFF_1411_Q_reg ( .D(g18820), .SI(g2631), .SE(n8167), .CLK(n8354), .Q(
        g2584), .QN(n4303) );
  SDFFX1 DFF_1412_Q_reg ( .D(n1423), .SI(g2584), .SE(n8240), .CLK(n8427), .Q(
        g2587) );
  SDFFX1 DFF_1413_Q_reg ( .D(g2587), .SI(g2587), .SE(n8240), .CLK(n8427), .Q(
        g2597) );
  SDFFX1 DFF_1414_Q_reg ( .D(g2597), .SI(g2597), .SE(n8240), .CLK(n8427), .Q(
        g2598) );
  SDFFX1 DFF_1415_Q_reg ( .D(g2530), .SI(g2598), .SE(n8239), .CLK(n8426), .Q(
        g2638) );
  SDFFX1 DFF_1416_Q_reg ( .D(g2638), .SI(g2638), .SE(n8239), .CLK(n8426), .Q(
        g2643) );
  SDFFX1 DFF_1417_Q_reg ( .D(g2533), .SI(g2643), .SE(n8239), .CLK(n8426), .Q(
        test_so86) );
  SDFFX1 DFF_1418_Q_reg ( .D(test_so86), .SI(test_si87), .SE(n8239), .CLK(
        n8426), .Q(g2645) );
  SDFFX1 DFF_1419_Q_reg ( .D(g2536), .SI(g2645), .SE(n8239), .CLK(n8426), .Q(
        g2646) );
  SDFFX1 DFF_1420_Q_reg ( .D(g2646), .SI(g2646), .SE(n8239), .CLK(n8426), .Q(
        g2647) );
  SDFFX1 DFF_1421_Q_reg ( .D(g2540), .SI(g2647), .SE(n8237), .CLK(n8424), .Q(
        g2648) );
  SDFFX1 DFF_1422_Q_reg ( .D(g2648), .SI(g2648), .SE(n8238), .CLK(n8425), .Q(
        g2639) );
  SDFFX1 DFF_1423_Q_reg ( .D(g2543), .SI(g2639), .SE(n8238), .CLK(n8425), .Q(
        g2640) );
  SDFFX1 DFF_1424_Q_reg ( .D(g2640), .SI(g2640), .SE(n8238), .CLK(n8425), .Q(
        g2641) );
  SDFFX1 DFF_1425_Q_reg ( .D(g2546), .SI(g2641), .SE(n8238), .CLK(n8425), .Q(
        g2642) );
  SDFFX1 DFF_1426_Q_reg ( .D(g2642), .SI(g2642), .SE(n8238), .CLK(n8425), .Q(
        g2564) );
  SDFFX1 DFF_1427_Q_reg ( .D(g2950), .SI(g2564), .SE(n8238), .CLK(n8425), .Q(
        g8087), .QN(n4456) );
  SDFFX1 DFF_1428_Q_reg ( .D(g8087), .SI(g8087), .SE(n8238), .CLK(n8425), .Q(
        g8167), .QN(n4455) );
  SDFFX1 DFF_1429_Q_reg ( .D(g8167), .SI(g8167), .SE(n8238), .CLK(n8425), .Q(
        g2560), .QN(n4463) );
  SDFFX1 DFF_1430_Q_reg ( .D(g23114), .SI(g2560), .SE(n8239), .CLK(n8426), .Q(
        g2561) );
  SDFFX1 DFF_1431_Q_reg ( .D(g23133), .SI(g2561), .SE(n8135), .CLK(n8322), .Q(
        g2562) );
  SDFFX1 DFF_1432_Q_reg ( .D(g21970), .SI(g2562), .SE(n8238), .CLK(n8425), .Q(
        test_so87) );
  SDFFX1 DFF_1433_Q_reg ( .D(g23407), .SI(test_si88), .SE(n8239), .CLK(n8426), 
        .Q(g2530) );
  SDFFX1 DFF_1434_Q_reg ( .D(g23418), .SI(g2530), .SE(n8239), .CLK(n8426), .Q(
        g2533) );
  SDFFX1 DFF_1435_Q_reg ( .D(g24209), .SI(g2533), .SE(n8239), .CLK(n8426), .Q(
        g2536) );
  SDFFX1 DFF_1436_Q_reg ( .D(g24214), .SI(g2536), .SE(n8240), .CLK(n8427), .Q(
        g2552) );
  SDFFX1 DFF_1437_Q_reg ( .D(g24226), .SI(g2552), .SE(n8240), .CLK(n8427), .Q(
        g2553) );
  SDFFX1 DFF_1438_Q_reg ( .D(g24238), .SI(g2553), .SE(n8240), .CLK(n8427), .Q(
        g2554) );
  SDFFX1 DFF_1439_Q_reg ( .D(g23132), .SI(g2554), .SE(n8237), .CLK(n8424), .Q(
        g2555) );
  SDFFX1 DFF_1440_Q_reg ( .D(g23047), .SI(g2555), .SE(n8237), .CLK(n8424), .Q(
        g2559) );
  SDFFX1 DFF_1441_Q_reg ( .D(g23076), .SI(g2559), .SE(n8237), .CLK(n8424), .Q(
        g2539) );
  SDFFX1 DFF_1442_Q_reg ( .D(g24225), .SI(g2539), .SE(n8237), .CLK(n8424), .Q(
        g2540) );
  SDFFX1 DFF_1443_Q_reg ( .D(g24237), .SI(g2540), .SE(n8238), .CLK(n8425), .Q(
        g2543) );
  SDFFX1 DFF_1444_Q_reg ( .D(g24250), .SI(g2543), .SE(n8238), .CLK(n8425), .Q(
        g2546) );
  SDFFX1 DFF_1445_Q_reg ( .D(n1402), .SI(g2546), .SE(n8238), .CLK(n8425), .Q(
        g2602) );
  SDFFX1 DFF_1446_Q_reg ( .D(g2602), .SI(g2602), .SE(n8239), .CLK(n8426), .Q(
        g2609) );
  SDFFX1 DFF_1447_Q_reg ( .D(g2609), .SI(g2609), .SE(n8239), .CLK(n8426), .Q(
        test_so88) );
  SDFFX1 DFF_1448_Q_reg ( .D(g13175), .SI(test_si89), .SE(n8240), .CLK(n8427), 
        .Q(g2617) );
  SDFFX1 DFF_1449_Q_reg ( .D(g2617), .SI(g2617), .SE(n8240), .CLK(n8427), .Q(
        n7930) );
  SDFFX1 DFF_1450_Q_reg ( .D(g30072), .SI(n7930), .SE(n8240), .CLK(n8427), .Q(
        n7929) );
  SDFFX1 DFF_1451_Q_reg ( .D(g13143), .SI(n7929), .SE(n8240), .CLK(n8427), .Q(
        g2623) );
  SDFFX1 DFF_1452_Q_reg ( .D(g2623), .SI(g2623), .SE(n8240), .CLK(n8427), .Q(
        g2574), .QN(n4543) );
  SDFFX1 DFF_1453_Q_reg ( .D(g13194), .SI(g2574), .SE(n8135), .CLK(n8322), .Q(
        g2632) );
  SDFFX1 DFF_1454_Q_reg ( .D(g2632), .SI(g2632), .SE(n8135), .CLK(n8322), .Q(
        g2633), .QN(n7749) );
  SDFFX1 DFF_1455_Q_reg ( .D(g27310), .SI(g2633), .SE(n8249), .CLK(n8436), .Q(
        g2650), .QN(n7326) );
  SDFFX1 DFF_1456_Q_reg ( .D(g27325), .SI(g2650), .SE(n8249), .CLK(n8436), .Q(
        g2651), .QN(n7328) );
  SDFFX1 DFF_1457_Q_reg ( .D(g27336), .SI(g2651), .SE(n8249), .CLK(n8436), .Q(
        g2649), .QN(n7327) );
  SDFFX1 DFF_1458_Q_reg ( .D(g27326), .SI(g2649), .SE(n8249), .CLK(n8436), .Q(
        g2653), .QN(n7338) );
  SDFFX1 DFF_1459_Q_reg ( .D(g27337), .SI(g2653), .SE(n8249), .CLK(n8436), .Q(
        g2654), .QN(n7340) );
  SDFFX1 DFF_1460_Q_reg ( .D(g27343), .SI(g2654), .SE(n8250), .CLK(n8437), .Q(
        g2652), .QN(n7339) );
  SDFFX1 DFF_1461_Q_reg ( .D(g27338), .SI(g2652), .SE(n8250), .CLK(n8437), .Q(
        g2656), .QN(n7165) );
  SDFFX1 DFF_1462_Q_reg ( .D(g27344), .SI(g2656), .SE(n8250), .CLK(n8437), .Q(
        test_so89), .QN(n8107) );
  SDFFX1 DFF_1463_Q_reg ( .D(g27347), .SI(test_si90), .SE(n8249), .CLK(n8436), 
        .Q(g2655), .QN(n7166) );
  SDFFX1 DFF_1464_Q_reg ( .D(g27345), .SI(g2655), .SE(n8250), .CLK(n8437), .Q(
        g2659), .QN(n7349) );
  SDFFX1 DFF_1465_Q_reg ( .D(g27348), .SI(g2659), .SE(n8250), .CLK(n8437), .Q(
        g2660), .QN(n7351) );
  SDFFX1 DFF_1466_Q_reg ( .D(g27354), .SI(g2660), .SE(n8248), .CLK(n8435), .Q(
        g2658), .QN(n7350) );
  SDFFX1 DFF_1467_Q_reg ( .D(g24527), .SI(g2658), .SE(n8248), .CLK(n8435), .Q(
        g2661) );
  SDFFX1 DFF_1468_Q_reg ( .D(g24537), .SI(g2661), .SE(n8248), .CLK(n8435), .Q(
        g2664) );
  SDFFX1 DFF_1469_Q_reg ( .D(g24547), .SI(g2664), .SE(n8249), .CLK(n8436), .Q(
        g2667) );
  SDFFX1 DFF_1470_Q_reg ( .D(g24538), .SI(g2667), .SE(n8249), .CLK(n8436), .Q(
        g2670) );
  SDFFX1 DFF_1471_Q_reg ( .D(g24548), .SI(g2670), .SE(n8249), .CLK(n8436), .Q(
        g2673) );
  SDFFX1 DFF_1472_Q_reg ( .D(g24557), .SI(g2673), .SE(n8249), .CLK(n8436), .Q(
        g2676) );
  SDFFX1 DFF_1473_Q_reg ( .D(g28364), .SI(g2676), .SE(n8249), .CLK(n8436), .Q(
        g2688) );
  SDFFX1 DFF_1474_Q_reg ( .D(g28368), .SI(g2688), .SE(n8249), .CLK(n8436), .Q(
        g2691) );
  SDFFX1 DFF_1475_Q_reg ( .D(g28371), .SI(g2691), .SE(n8248), .CLK(n8435), .Q(
        g2694) );
  SDFFX1 DFF_1476_Q_reg ( .D(g28358), .SI(g2694), .SE(n8250), .CLK(n8437), .Q(
        g2679) );
  SDFFX1 DFF_1477_Q_reg ( .D(g28363), .SI(g2679), .SE(n8250), .CLK(n8437), .Q(
        test_so90) );
  SDFFX1 DFF_1478_Q_reg ( .D(g28367), .SI(test_si91), .SE(n8250), .CLK(n8437), 
        .Q(g2685) );
  SDFFX1 DFF_1479_Q_reg ( .D(g26575), .SI(g2685), .SE(n8250), .CLK(n8437), .Q(
        g2565) );
  SDFFX1 DFF_1480_Q_reg ( .D(g26596), .SI(g2565), .SE(n8250), .CLK(n8437), .Q(
        g2568) );
  SDFFX1 DFF_1481_Q_reg ( .D(g26616), .SI(g2568), .SE(n8248), .CLK(n8435), .Q(
        g2571) );
  SDFFX1 DFF_1482_Q_reg ( .D(g2574), .SI(g2571), .SE(n8248), .CLK(n8435), .Q(
        g2580), .QN(n7489) );
  SDFFX1 DFF_1483_Q_reg ( .D(g22687), .SI(g2580), .SE(n8250), .CLK(n8437), .Q(
        n7926) );
  SDFFX1 DFF_1492_Q_reg ( .D(g30061), .SI(n7926), .SE(n8250), .CLK(n8437), .Q(
        g16437) );
  SDFFX1 DFF_1493_Q_reg ( .D(g16437), .SI(g16437), .SE(n8251), .CLK(n8438), 
        .Q(g2599), .QN(n8039) );
  SDFFX1 DFF_1494_Q_reg ( .D(DFF_1349_n1), .SI(g2599), .SE(n8251), .CLK(n8438), 
        .Q(n7925), .QN(DFF_1494_n1) );
  SDFFX1 DFF_1495_Q_reg ( .D(DFF_1351_n1), .SI(n7925), .SE(n8251), .CLK(n8438), 
        .Q(n7924), .QN(DFF_1495_n1) );
  SDFFX1 DFF_1496_Q_reg ( .D(DFF_1353_n1), .SI(n7924), .SE(n8251), .CLK(n8438), 
        .Q(n7923), .QN(DFF_1496_n1) );
  SDFFX1 DFF_1497_Q_reg ( .D(DFF_1355_n1), .SI(n7923), .SE(n8251), .CLK(n8438), 
        .Q(n7922), .QN(DFF_1497_n1) );
  SDFFX1 DFF_1498_Q_reg ( .D(DFF_1357_n1), .SI(n7922), .SE(n8251), .CLK(n8438), 
        .Q(n7921), .QN(DFF_1498_n1) );
  SDFFX1 DFF_1499_Q_reg ( .D(DFF_1359_n1), .SI(n7921), .SE(n8251), .CLK(n8438), 
        .Q(n7920), .QN(DFF_1499_n1) );
  SDFFX1 DFF_1500_Q_reg ( .D(DFF_1361_n1), .SI(n7920), .SE(n8251), .CLK(n8438), 
        .Q(test_so91), .QN(n7145) );
  SDFFX1 DFF_1501_Q_reg ( .D(DFF_1363_n1), .SI(test_si92), .SE(n8144), .CLK(
        n8331), .Q(g2611), .QN(n7144) );
  SDFFX1 DFF_1502_Q_reg ( .D(g24092), .SI(g2611), .SE(n8246), .CLK(n8433), .Q(
        g2612), .QN(n4490) );
  SDFFX1 DFF_1503_Q_reg ( .D(n4483), .SI(g2612), .SE(n8164), .CLK(n8351), .Q(
        n7918), .QN(n14346) );
  SDFFX1 DFF_1505_Q_reg ( .D(g7425), .SI(g7425), .SE(n8164), .CLK(n8351), .Q(
        g7487) );
  SDFFX1 DFF_1506_Q_reg ( .D(g7487), .SI(g7487), .SE(n8164), .CLK(n8351), .Q(
        g2703), .QN(n4292) );
  SDFFX1 DFF_1507_Q_reg ( .D(g16718), .SI(g2703), .SE(n8167), .CLK(n8354), .Q(
        g2704), .QN(n7745) );
  SDFFX1 DFF_1508_Q_reg ( .D(g20375), .SI(g2704), .SE(n8167), .CLK(n8354), .Q(
        g2733), .QN(n4426) );
  SDFFX1 DFF_1509_Q_reg ( .D(g20789), .SI(g2733), .SE(n8167), .CLK(n8354), .Q(
        g2714), .QN(n4398) );
  SDFFX1 DFF_1510_Q_reg ( .D(n1502), .SI(g2714), .SE(n8167), .CLK(n8354), .Q(
        g2707), .QN(n4472) );
  SDFFX1 DFF_1511_Q_reg ( .D(g23348), .SI(g2707), .SE(n8167), .CLK(n8354), .Q(
        g2727), .QN(n4419) );
  SDFFX1 DFF_1512_Q_reg ( .D(g24438), .SI(g2727), .SE(n8167), .CLK(n8354), .Q(
        g2720), .QN(n4408) );
  SDFFX1 DFF_1513_Q_reg ( .D(g25197), .SI(g2720), .SE(n8167), .CLK(n8354), .Q(
        g2734), .QN(n4397) );
  SDFFX1 DFF_1514_Q_reg ( .D(n1503), .SI(g2734), .SE(n8167), .CLK(n8354), .Q(
        g2746), .QN(n4407) );
  SDFFX1 DFF_1515_Q_reg ( .D(g26795), .SI(g2746), .SE(n8168), .CLK(n8355), .Q(
        test_so92), .QN(n8073) );
  SDFFX1 DFF_1516_Q_reg ( .D(g27243), .SI(test_si93), .SE(n8168), .CLK(n8355), 
        .Q(g2753), .QN(n4471) );
  SDFFX1 DFF_1517_Q_reg ( .D(g27724), .SI(g2753), .SE(n8168), .CLK(n8355), .Q(
        g2760), .QN(n4393) );
  SDFFX1 DFF_1518_Q_reg ( .D(g28328), .SI(g2760), .SE(n8168), .CLK(n8355), .Q(
        g2766), .QN(n4415) );
  SDFFX1 DFF_1519_Q_reg ( .D(g20918), .SI(g2766), .SE(n8251), .CLK(n8438), .Q(
        g2773), .QN(n7772) );
  SDFFX1 DFF_1520_Q_reg ( .D(g20939), .SI(g2773), .SE(n8251), .CLK(n8438), .Q(
        g2774), .QN(n7771) );
  SDFFX1 DFF_1521_Q_reg ( .D(g20962), .SI(g2774), .SE(n8252), .CLK(n8439), .Q(
        g2772), .QN(n7834) );
  SDFFX1 DFF_1522_Q_reg ( .D(g20940), .SI(g2772), .SE(n8252), .CLK(n8439), .Q(
        g2776), .QN(n7770) );
  SDFFX1 DFF_1523_Q_reg ( .D(g20963), .SI(g2776), .SE(n8252), .CLK(n8439), .Q(
        g2777), .QN(n7769) );
  SDFFX1 DFF_1524_Q_reg ( .D(g20981), .SI(g2777), .SE(n8253), .CLK(n8440), .Q(
        g2775), .QN(n7833) );
  SDFFX1 DFF_1525_Q_reg ( .D(g20964), .SI(g2775), .SE(n8253), .CLK(n8440), .Q(
        g2779), .QN(n7768) );
  SDFFX1 DFF_1526_Q_reg ( .D(g20982), .SI(g2779), .SE(n8253), .CLK(n8440), .Q(
        g2780), .QN(n7767) );
  SDFFX1 DFF_1527_Q_reg ( .D(g21004), .SI(g2780), .SE(n8253), .CLK(n8440), .Q(
        g2778), .QN(n7832) );
  SDFFX1 DFF_1528_Q_reg ( .D(g20983), .SI(g2778), .SE(n8253), .CLK(n8440), .Q(
        g2782), .QN(n7766) );
  SDFFX1 DFF_1529_Q_reg ( .D(g21005), .SI(g2782), .SE(n8253), .CLK(n8440), .Q(
        g2783), .QN(n7765) );
  SDFFX1 DFF_1530_Q_reg ( .D(g21025), .SI(g2783), .SE(n8253), .CLK(n8440), .Q(
        test_so93), .QN(n8119) );
  SDFFX1 DFF_1531_Q_reg ( .D(g21006), .SI(test_si94), .SE(n8251), .CLK(n8438), 
        .Q(g2785), .QN(n7764) );
  SDFFX1 DFF_1532_Q_reg ( .D(g21026), .SI(g2785), .SE(n8252), .CLK(n8439), .Q(
        g2786), .QN(n7763) );
  SDFFX1 DFF_1533_Q_reg ( .D(g21043), .SI(g2786), .SE(n8253), .CLK(n8440), .Q(
        g2784), .QN(n7831) );
  SDFFX1 DFF_1534_Q_reg ( .D(g21027), .SI(g2784), .SE(n8253), .CLK(n8440), .Q(
        g2788), .QN(n7762) );
  SDFFX1 DFF_1535_Q_reg ( .D(g21044), .SI(g2788), .SE(n8253), .CLK(n8440), .Q(
        g2789), .QN(n7761) );
  SDFFX1 DFF_1536_Q_reg ( .D(g21060), .SI(g2789), .SE(n8253), .CLK(n8440), .Q(
        g2787), .QN(n7830) );
  SDFFX1 DFF_1537_Q_reg ( .D(g21045), .SI(g2787), .SE(n8253), .CLK(n8440), .Q(
        g2791), .QN(n7760) );
  SDFFX1 DFF_1538_Q_reg ( .D(g21061), .SI(g2791), .SE(n8254), .CLK(n8441), .Q(
        g2792), .QN(n7759) );
  SDFFX1 DFF_1539_Q_reg ( .D(g21073), .SI(g2792), .SE(n8254), .CLK(n8441), .Q(
        g2790), .QN(n7829) );
  SDFFX1 DFF_1540_Q_reg ( .D(g21062), .SI(g2790), .SE(n8254), .CLK(n8441), .Q(
        g2794), .QN(n7758) );
  SDFFX1 DFF_1541_Q_reg ( .D(g21074), .SI(g2794), .SE(n8254), .CLK(n8441), .Q(
        g2795), .QN(n7757) );
  SDFFX1 DFF_1542_Q_reg ( .D(g21081), .SI(g2795), .SE(n8254), .CLK(n8441), .Q(
        g2793), .QN(n7828) );
  SDFFX1 DFF_1543_Q_reg ( .D(g21075), .SI(g2793), .SE(n8254), .CLK(n8441), .Q(
        g2797), .QN(n7756) );
  SDFFX1 DFF_1544_Q_reg ( .D(g21082), .SI(g2797), .SE(n8254), .CLK(n8441), .Q(
        g2798), .QN(n7755) );
  SDFFX1 DFF_1545_Q_reg ( .D(g21094), .SI(g2798), .SE(n8254), .CLK(n8441), .Q(
        test_so94), .QN(n8120) );
  SDFFX1 DFF_1546_Q_reg ( .D(g20919), .SI(test_si95), .SE(n8251), .CLK(n8438), 
        .Q(g2800), .QN(n7754) );
  SDFFX1 DFF_1547_Q_reg ( .D(g20941), .SI(g2800), .SE(n8252), .CLK(n8439), .Q(
        g2801), .QN(n7753) );
  SDFFX1 DFF_1548_Q_reg ( .D(g20965), .SI(g2801), .SE(n8252), .CLK(n8439), .Q(
        g2799), .QN(n7827) );
  SDFFX1 DFF_1549_Q_reg ( .D(g21007), .SI(g2799), .SE(n8252), .CLK(n8439), .Q(
        g2803), .QN(n8029) );
  SDFFX1 DFF_1550_Q_reg ( .D(g21028), .SI(g2803), .SE(n8252), .CLK(n8439), .Q(
        g2804), .QN(n7556) );
  SDFFX1 DFF_1551_Q_reg ( .D(g21046), .SI(g2804), .SE(n8252), .CLK(n8439), .Q(
        g2802) );
  SDFFX1 DFF_1552_Q_reg ( .D(g21029), .SI(g2802), .SE(n8252), .CLK(n8439), .Q(
        g2806), .QN(n7563) );
  SDFFX1 DFF_1553_Q_reg ( .D(g21047), .SI(g2806), .SE(n8252), .CLK(n8439), .Q(
        g2807), .QN(n7555) );
  SDFFX1 DFF_1554_Q_reg ( .D(g21063), .SI(g2807), .SE(n8252), .CLK(n8439), .Q(
        g2805), .QN(n7613) );
  SDFFX1 DFF_1555_Q_reg ( .D(g25272), .SI(g2805), .SE(n8254), .CLK(n8441), .Q(
        g2809), .QN(n7491) );
  SDFFX1 DFF_1556_Q_reg ( .D(g25280), .SI(g2809), .SE(n8254), .CLK(n8441), .Q(
        g2810), .QN(n7490) );
  SDFFX1 DFF_1557_Q_reg ( .D(g25288), .SI(g2810), .SE(n8254), .CLK(n8441), .Q(
        g2808), .QN(n7498) );
  SDFFX1 DFF_1558_Q_reg ( .D(g22269), .SI(g2808), .SE(n8254), .CLK(n8441), .Q(
        g2812), .QN(n7865) );
  SDFFX1 DFF_1559_Q_reg ( .D(g22284), .SI(g2812), .SE(n8255), .CLK(n8442), .Q(
        g2813), .QN(n7953) );
  SDFFX1 DFF_1560_Q_reg ( .D(g22299), .SI(g2813), .SE(n8255), .CLK(n8442), .Q(
        test_so95), .QN(n8101) );
  SDFFX1 DFF_1561_Q_reg ( .D(g20877), .SI(test_si96), .SE(n8130), .CLK(n8317), 
        .Q(n7913), .QN(DFF_1561_n1) );
  SDFFX1 DFF_1562_Q_reg ( .D(g20884), .SI(n7913), .SE(n8130), .CLK(n8317), .Q(
        n7912), .QN(DFF_1562_n1) );
  SDFFX1 DFF_1563_Q_reg ( .D(n4263), .SI(n7912), .SE(n8130), .CLK(n8317), .Q(
        n4598), .QN(n8031) );
  SDFFX1 DFF_1564_Q_reg ( .D(n4269), .SI(n4598), .SE(n8194), .CLK(n8381), .Q(
        g3043) );
  SDFFX1 DFF_1565_Q_reg ( .D(n4268), .SI(g3043), .SE(n8194), .CLK(n8381), .Q(
        g3044) );
  SDFFX1 DFF_1566_Q_reg ( .D(n4267), .SI(g3044), .SE(n8194), .CLK(n8381), .Q(
        g3045) );
  SDFFX1 DFF_1567_Q_reg ( .D(n4266), .SI(g3045), .SE(n8195), .CLK(n8382), .Q(
        g3046) );
  SDFFX1 DFF_1568_Q_reg ( .D(n4265), .SI(g3046), .SE(n8195), .CLK(n8382), .Q(
        g3047) );
  SDFFX1 DFF_1569_Q_reg ( .D(n4272), .SI(g3047), .SE(n8195), .CLK(n8382), .Q(
        g3048) );
  SDFFX1 DFF_1570_Q_reg ( .D(n4271), .SI(g3048), .SE(n8195), .CLK(n8382), .Q(
        g3049) );
  SDFFX1 DFF_1571_Q_reg ( .D(n4270), .SI(g3049), .SE(n8195), .CLK(n8382), .Q(
        g3050) );
  SDFFX1 DFF_1572_Q_reg ( .D(n4259), .SI(g3050), .SE(n8195), .CLK(n8382), .Q(
        g3051) );
  SDFFX1 DFF_1573_Q_reg ( .D(n4236), .SI(g3051), .SE(n8222), .CLK(n8409), .Q(
        g3052) );
  SDFFX1 DFF_1574_Q_reg ( .D(n4239), .SI(g3052), .SE(n8222), .CLK(n8409), .Q(
        g3053) );
  SDFFX1 DFF_1575_Q_reg ( .D(n4237), .SI(g3053), .SE(n8222), .CLK(n8409), .Q(
        test_so96) );
  SDFFX1 DFF_1576_Q_reg ( .D(n4234), .SI(test_si97), .SE(n8222), .CLK(n8409), 
        .Q(g3056) );
  SDFFX1 DFF_1577_Q_reg ( .D(n4233), .SI(g3056), .SE(n8222), .CLK(n8409), .Q(
        g3057) );
  SDFFX1 DFF_1578_Q_reg ( .D(n4238), .SI(g3057), .SE(n8223), .CLK(n8410), .Q(
        g3058) );
  SDFFX1 DFF_1579_Q_reg ( .D(n4235), .SI(g3058), .SE(n8223), .CLK(n8410), .Q(
        g3059) );
  SDFFX1 DFF_1580_Q_reg ( .D(n4240), .SI(g3059), .SE(n8223), .CLK(n8410), .Q(
        g3060) );
  SDFFX1 DFF_1581_Q_reg ( .D(n4232), .SI(g3060), .SE(n8223), .CLK(n8410), .Q(
        g3061) );
  SDFFX1 DFF_1582_Q_reg ( .D(n4245), .SI(g3061), .SE(n8246), .CLK(n8433), .Q(
        g3062) );
  SDFFX1 DFF_1583_Q_reg ( .D(n4248), .SI(g3062), .SE(n8247), .CLK(n8434), .Q(
        g3063) );
  SDFFX1 DFF_1584_Q_reg ( .D(n4246), .SI(g3063), .SE(n8247), .CLK(n8434), .Q(
        g3064) );
  SDFFX1 DFF_1585_Q_reg ( .D(n4243), .SI(g3064), .SE(n8247), .CLK(n8434), .Q(
        g3065) );
  SDFFX1 DFF_1586_Q_reg ( .D(n4242), .SI(g3065), .SE(n8247), .CLK(n8434), .Q(
        g3066) );
  SDFFX1 DFF_1587_Q_reg ( .D(n4247), .SI(g3066), .SE(n8247), .CLK(n8434), .Q(
        g3067) );
  SDFFX1 DFF_1588_Q_reg ( .D(n4244), .SI(g3067), .SE(n8247), .CLK(n8434), .Q(
        g3068) );
  SDFFX1 DFF_1589_Q_reg ( .D(n4249), .SI(g3068), .SE(n8248), .CLK(n8435), .Q(
        g3069) );
  SDFFX1 DFF_1590_Q_reg ( .D(n4241), .SI(g3069), .SE(n8248), .CLK(n8435), .Q(
        test_so97) );
  SDFFX1 DFF_1591_Q_reg ( .D(n4254), .SI(test_si98), .SE(n8255), .CLK(n8442), 
        .Q(g3071) );
  SDFFX1 DFF_1592_Q_reg ( .D(n4257), .SI(g3071), .SE(n8255), .CLK(n8442), .Q(
        g3072) );
  SDFFX1 DFF_1593_Q_reg ( .D(n4255), .SI(g3072), .SE(n8255), .CLK(n8442), .Q(
        g3073) );
  SDFFX1 DFF_1594_Q_reg ( .D(n4252), .SI(g3073), .SE(n8255), .CLK(n8442), .Q(
        g3074) );
  SDFFX1 DFF_1595_Q_reg ( .D(n4251), .SI(g3074), .SE(n8255), .CLK(n8442), .Q(
        g3075) );
  SDFFX1 DFF_1596_Q_reg ( .D(n4256), .SI(g3075), .SE(n8256), .CLK(n8443), .Q(
        g3076) );
  SDFFX1 DFF_1597_Q_reg ( .D(n4253), .SI(g3076), .SE(n8256), .CLK(n8443), .Q(
        g3077) );
  SDFFX1 DFF_1598_Q_reg ( .D(n4258), .SI(g3077), .SE(n8256), .CLK(n8443), .Q(
        g3078) );
  SDFFX1 DFF_1599_Q_reg ( .D(n4250), .SI(g3078), .SE(n8164), .CLK(n8351), .Q(
        g2997) );
  SDFFX1 DFF_1600_Q_reg ( .D(g25265), .SI(g2997), .SE(n8164), .CLK(n8351), .Q(
        g2993), .QN(n8032) );
  SDFFX1 DFF_1601_Q_reg ( .D(g26048), .SI(g2993), .SE(n8164), .CLK(n8351), .Q(
        n7909), .QN(n14354) );
  SDFFX1 DFF_1602_Q_reg ( .D(n1538), .SI(n7909), .SE(n8164), .CLK(n8351), .Q(
        g3006), .QN(n8035) );
  SDFFX1 DFF_1603_Q_reg ( .D(g24445), .SI(g3006), .SE(n8164), .CLK(n8351), .Q(
        g3002), .QN(n8034) );
  SDFFX1 DFF_1604_Q_reg ( .D(g25191), .SI(g3002), .SE(n8165), .CLK(n8352), .Q(
        g3013), .QN(n8051) );
  SDFFX1 DFF_1605_Q_reg ( .D(g26031), .SI(g3013), .SE(n8165), .CLK(n8352), .Q(
        test_so98) );
  SDFFX1 DFF_1606_Q_reg ( .D(g26786), .SI(test_si99), .SE(n8165), .CLK(n8352), 
        .Q(g3024), .QN(n8033) );
  SDFFX1 DFF_1607_Q_reg ( .D(n4262), .SI(g3024), .SE(n8165), .CLK(n8352), .Q(
        g3018), .QN(n4481) );
  SDFFX1 DFF_1608_Q_reg ( .D(n1540), .SI(g3018), .SE(n8165), .CLK(n8352), .Q(
        g3028), .QN(n4350) );
  SDFFX1 DFF_1609_Q_reg ( .D(g24446), .SI(g3028), .SE(n8165), .CLK(n8352), .Q(
        g3036), .QN(n4480) );
  SDFFX1 DFF_1610_Q_reg ( .D(g25202), .SI(g3036), .SE(n8165), .CLK(n8352), .Q(
        g3032), .QN(n7429) );
  SDFFX1 DFF_1611_Q_reg ( .D(g3234), .SI(g3032), .SE(n8165), .CLK(n8352), .Q(
        g5388) );
  SDFFX1 DFF_1612_Q_reg ( .D(g5388), .SI(g5388), .SE(n8165), .CLK(n8352), .Q(
        n7907), .QN(DFF_1612_n1) );
  SDFFX1 DFF_1613_Q_reg ( .D(g16496), .SI(n7907), .SE(n8165), .CLK(n8352), .Q(
        g2987), .QN(n4365) );
  SDFFX1 DFF_1614_Q_reg ( .D(g16824), .SI(g2987), .SE(n8246), .CLK(n8433), .Q(
        g8275) );
  SDFFX1 DFF_1615_Q_reg ( .D(g16844), .SI(g8275), .SE(n8247), .CLK(n8434), .Q(
        g8274), .QN(n8002) );
  SDFFX1 DFF_1616_Q_reg ( .D(g16853), .SI(g8274), .SE(n8247), .CLK(n8434), .Q(
        g8273), .QN(n14358) );
  SDFFX1 DFF_1617_Q_reg ( .D(g16860), .SI(g8273), .SE(n8247), .CLK(n8434), .Q(
        g8272), .QN(n14357) );
  SDFFX1 DFF_1618_Q_reg ( .D(g16803), .SI(g8272), .SE(n8247), .CLK(n8434), .Q(
        g8268), .QN(n14356) );
  SDFFX1 DFF_1619_Q_reg ( .D(g16835), .SI(g8268), .SE(n8247), .CLK(n8434), .Q(
        g8269), .QN(n8010) );
  SDFFX1 DFF_1620_Q_reg ( .D(g16851), .SI(g8269), .SE(n8247), .CLK(n8434), .Q(
        test_so99) );
  SDFFX1 DFF_1621_Q_reg ( .D(g16857), .SI(test_si100), .SE(n8248), .CLK(n8435), 
        .Q(g8271), .QN(n8001) );
  SDFFX1 DFF_1622_Q_reg ( .D(g16866), .SI(g8271), .SE(n8248), .CLK(n8435), .Q(
        g3083), .QN(n8013) );
  SDFFX1 DFF_1623_Q_reg ( .D(n4261), .SI(g3083), .SE(n8248), .CLK(n8435), .Q(
        g8267) );
  SDFFX1 DFF_1624_Q_reg ( .D(N995), .SI(g8267), .SE(n8248), .CLK(n8435), .Q(
        n4577), .QN(n7432) );
  SDFFX1 DFF_1625_Q_reg ( .D(g16845), .SI(n4577), .SE(n8255), .CLK(n8442), .Q(
        g8266), .QN(n14361) );
  SDFFX1 DFF_1626_Q_reg ( .D(g16854), .SI(g8266), .SE(n8255), .CLK(n8442), .Q(
        g8265), .QN(n14360) );
  SDFFX1 DFF_1627_Q_reg ( .D(g16861), .SI(g8265), .SE(n8255), .CLK(n8442), .Q(
        g8264), .QN(n7975) );
  SDFFX1 DFF_1628_Q_reg ( .D(g16880), .SI(g8264), .SE(n8255), .CLK(n8442), .Q(
        g8262) );
  SDFFX1 DFF_1629_Q_reg ( .D(g18755), .SI(g8262), .SE(n8255), .CLK(n8442), .Q(
        g8263), .QN(n7976) );
  SDFFX1 DFF_1630_Q_reg ( .D(g18804), .SI(g8263), .SE(n8256), .CLK(n8443), .Q(
        g8260), .QN(n7973) );
  SDFFX1 DFF_1631_Q_reg ( .D(g18837), .SI(g8260), .SE(n8256), .CLK(n8443), .Q(
        g8261), .QN(n14359) );
  SDFFX1 DFF_1632_Q_reg ( .D(g18868), .SI(g8261), .SE(n8256), .CLK(n8443), .Q(
        g8259), .QN(n7974) );
  SDFFX1 DFF_1633_Q_reg ( .D(g18907), .SI(g8259), .SE(n8256), .CLK(n8443), .Q(
        g2990), .QN(n8011) );
  SDFFX1 DFF_1634_Q_reg ( .D(N690), .SI(g2990), .SE(n8256), .CLK(n8443), .Q(
        n4578), .QN(n7431) );
  SDFFX1 DFF_1635_Q_reg ( .D(n4260), .SI(n4578), .SE(n8256), .CLK(n8443), .Q(
        test_so100) );
  SDFFX1 DFF_454_Q_reg ( .D(n4598), .SI(n8040), .SE(n8163), .CLK(n8350), .Q(
        g6677), .QN(n4309) );
  SDFFX1 DFF_804_Q_reg ( .D(n4598), .SI(test_si49), .SE(n8130), .CLK(n8317), 
        .Q(g6979), .QN(n4308) );
  SDFFX1 DFF_1154_Q_reg ( .D(n4598), .SI(n7960), .SE(n8138), .CLK(n8325), .Q(
        g7229), .QN(n4307) );
  SDFFX1 DFF_1504_Q_reg ( .D(n4598), .SI(n7918), .SE(n8164), .CLK(n8351), .Q(
        g7425), .QN(n4306) );
  SDFFX1 DFF_1300_Q_reg ( .D(g5555), .SI(g5555), .SE(n8232), .CLK(n8419), .Q(
        g7264), .QN(n4524) );
  SDFFX1 DFF_950_Q_reg ( .D(g5511), .SI(g5511), .SE(n8204), .CLK(n8391), .Q(
        g7014), .QN(n4525) );
  SDFFX1 DFF_951_Q_reg ( .D(g7014), .SI(g7014), .SE(n8204), .CLK(n8391), .Q(
        n4618), .QN(n4511) );
  SDFFX1 DFF_1301_Q_reg ( .D(g7264), .SI(g7264), .SE(n8232), .CLK(n8419), .Q(
        n4606), .QN(n4509) );
  SDFFX1 DFF_250_Q_reg ( .D(g5437), .SI(g5437), .SE(n8147), .CLK(n8334), .Q(
        g6447), .QN(n4499) );
  SDFFX1 DFF_249_Q_reg ( .D(g2950), .SI(g181), .SE(n8147), .CLK(n8334), .Q(
        g5437), .QN(n4520) );
  NOR2X0 Trojan1 ( .IN1(n4037), .IN2(n4043), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(n4034), .IN2(n4033), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(n4046), .IN2(n4038), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(n2568), .IN2(n3457), .QN(Tj_OUT4) );
  NOR4X0 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .QN(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(n3478), .IN2(n3469), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n3445), .IN2(n3212), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(n3237), .IN2(n3225), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(n3196), .IN2(n3417), .QN(Tj_OUT8) );
  NOR4X0 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .QN(Tj_OUT5678) );
  AND2X1 Trojan_CLK_NOT ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .Q(Tj_Trigger)
         );
  DFFX2 Trojan_Payload1 ( .D(1'b1), .CLK(Tj_Trigger), .Q(RingOscENable1) );
  DFFX2 Trojan_Payload2 ( .D(1'b0), .CLK(Tj_Trigger), .QN(RingOscENable2) );
  DFFX2 Trojan_Payload3 ( .D(1'b1), .CLK(Tj_Trigger), .Q(RingOscENable3) );
  AND3X4 Trojan_Payload ( .IN1(RingOscENable1), .IN2(RingOscENable2), .IN3(
        RingOscENable3), .Q(RingOscENable) );
  NAND3X1 TrojanEnableGATE ( .IN1(Out29), .IN2(RingOscENable), .IN3(g16692), 
        .QN(Out1) );
  INVX8 Trojan_Inv1 ( .INP(Out1), .ZN(Out2) );
  INVX8 Trojan_Inv2 ( .INP(Out2), .ZN(Out3) );
  INVX8 Trojan_Inv3 ( .INP(Out3), .ZN(Out4) );
  INVX8 Trojan_Inv4 ( .INP(Out4), .ZN(Out5) );
  INVX8 Trojan_Inv5 ( .INP(Out5), .ZN(Out6) );
  INVX8 Trojan_Inv6 ( .INP(Out6), .ZN(Out7) );
  INVX8 Trojan_Inv7 ( .INP(Out7), .ZN(Out8) );
  INVX8 Trojan_Inv8 ( .INP(Out8), .ZN(Out9) );
  INVX8 Trojan_Inv9 ( .INP(Out9), .ZN(Out10) );
  INVX8 Trojan_Inv10 ( .INP(Out10), .ZN(Out11) );
  INVX8 Trojan_Inv11 ( .INP(Out11), .ZN(Out12) );
  INVX8 Trojan_Inv12 ( .INP(Out12), .ZN(Out13) );
  INVX8 Trojan_Inv13 ( .INP(Out13), .ZN(Out14) );
  INVX8 Trojan_Inv14 ( .INP(Out14), .ZN(Out15) );
  INVX8 Trojan_Inv15 ( .INP(Out15), .ZN(Out16) );
  INVX8 Trojan_Inv16 ( .INP(Out16), .ZN(Out17) );
  INVX8 Trojan_Inv17 ( .INP(Out17), .ZN(Out18) );
  INVX8 Trojan_Inv18 ( .INP(Out18), .ZN(Out19) );
  INVX8 Trojan_Inv19 ( .INP(Out19), .ZN(Out20) );
  INVX8 Trojan_Inv20 ( .INP(Out20), .ZN(Out21) );
  INVX8 Trojan_Inv21 ( .INP(Out21), .ZN(Out22) );
  INVX8 Trojan_Inv22 ( .INP(Out22), .ZN(Out23) );
  INVX8 Trojan_Inv23 ( .INP(Out23), .ZN(Out24) );
  INVX8 Trojan_Inv24 ( .INP(Out24), .ZN(Out25) );
  INVX8 Trojan_Inv25 ( .INP(Out25), .ZN(Out26) );
  INVX8 Trojan_Inv26 ( .INP(Out26), .ZN(Out27) );
  INVX8 Trojan_Inv27 ( .INP(Out27), .ZN(Out28) );
  INVX8 Trojan_Inv28 ( .INP(Out28), .ZN(Out29) );
  NBUFFX2 U7966 ( .INP(n8304), .Z(n8130) );
  NBUFFX2 U7967 ( .INP(n8304), .Z(n8131) );
  NBUFFX2 U7968 ( .INP(n8265), .Z(n8247) );
  NBUFFX2 U7969 ( .INP(n8262), .Z(n8255) );
  NBUFFX2 U7970 ( .INP(n8263), .Z(n8254) );
  NBUFFX2 U7971 ( .INP(n8263), .Z(n8253) );
  NBUFFX2 U7972 ( .INP(n8263), .Z(n8252) );
  NBUFFX2 U7973 ( .INP(n8264), .Z(n8251) );
  NBUFFX2 U7974 ( .INP(n8265), .Z(n8248) );
  NBUFFX2 U7975 ( .INP(n8264), .Z(n8250) );
  NBUFFX2 U7976 ( .INP(n8264), .Z(n8249) );
  NBUFFX2 U7977 ( .INP(n8268), .Z(n8238) );
  NBUFFX2 U7978 ( .INP(n8268), .Z(n8239) );
  NBUFFX2 U7979 ( .INP(n8266), .Z(n8245) );
  NBUFFX2 U7980 ( .INP(n8265), .Z(n8246) );
  NBUFFX2 U7981 ( .INP(n8300), .Z(n8143) );
  NBUFFX2 U7982 ( .INP(n8267), .Z(n8240) );
  NBUFFX2 U7983 ( .INP(n8268), .Z(n8237) );
  NBUFFX2 U7984 ( .INP(n8267), .Z(n8241) );
  NBUFFX2 U7985 ( .INP(n8270), .Z(n8231) );
  NBUFFX2 U7986 ( .INP(n8267), .Z(n8242) );
  NBUFFX2 U7987 ( .INP(n8269), .Z(n8236) );
  NBUFFX2 U7988 ( .INP(n8266), .Z(n8244) );
  NBUFFX2 U7989 ( .INP(n8266), .Z(n8243) );
  NBUFFX2 U7990 ( .INP(n8270), .Z(n8233) );
  NBUFFX2 U7991 ( .INP(n8270), .Z(n8232) );
  NBUFFX2 U7992 ( .INP(n8269), .Z(n8235) );
  NBUFFX2 U7993 ( .INP(n8269), .Z(n8234) );
  NBUFFX2 U7994 ( .INP(n8271), .Z(n8230) );
  NBUFFX2 U7995 ( .INP(n8271), .Z(n8229) );
  NBUFFX2 U7996 ( .INP(n8271), .Z(n8228) );
  NBUFFX2 U7997 ( .INP(n8272), .Z(n8227) );
  NBUFFX2 U7998 ( .INP(n8275), .Z(n8218) );
  NBUFFX2 U7999 ( .INP(n8272), .Z(n8226) );
  NBUFFX2 U8000 ( .INP(n8273), .Z(n8223) );
  NBUFFX2 U8001 ( .INP(n8272), .Z(n8225) );
  NBUFFX2 U8002 ( .INP(n8273), .Z(n8224) );
  NBUFFX2 U8003 ( .INP(n8273), .Z(n8222) );
  NBUFFX2 U8004 ( .INP(n8274), .Z(n8221) );
  NBUFFX2 U8005 ( .INP(n8274), .Z(n8220) );
  NBUFFX2 U8006 ( .INP(n8274), .Z(n8219) );
  NBUFFX2 U8007 ( .INP(n8275), .Z(n8217) );
  NBUFFX2 U8008 ( .INP(n8275), .Z(n8216) );
  NBUFFX2 U8009 ( .INP(n8276), .Z(n8215) );
  NBUFFX2 U8010 ( .INP(n8276), .Z(n8214) );
  NBUFFX2 U8011 ( .INP(n8277), .Z(n8210) );
  NBUFFX2 U8012 ( .INP(n8277), .Z(n8211) );
  NBUFFX2 U8013 ( .INP(n8279), .Z(n8204) );
  NBUFFX2 U8014 ( .INP(n8278), .Z(n8209) );
  NBUFFX2 U8015 ( .INP(n8278), .Z(n8208) );
  NBUFFX2 U8016 ( .INP(n8276), .Z(n8213) );
  NBUFFX2 U8017 ( .INP(n8277), .Z(n8212) );
  NBUFFX2 U8018 ( .INP(n8278), .Z(n8207) );
  NBUFFX2 U8019 ( .INP(n8279), .Z(n8206) );
  NBUFFX2 U8020 ( .INP(n8279), .Z(n8205) );
  NBUFFX2 U8021 ( .INP(n8280), .Z(n8203) );
  NBUFFX2 U8022 ( .INP(n8280), .Z(n8202) );
  NBUFFX2 U8023 ( .INP(n8280), .Z(n8201) );
  NBUFFX2 U8024 ( .INP(n8281), .Z(n8200) );
  NBUFFX2 U8025 ( .INP(n8281), .Z(n8199) );
  NBUFFX2 U8026 ( .INP(n8281), .Z(n8198) );
  NBUFFX2 U8027 ( .INP(n8282), .Z(n8197) );
  NBUFFX2 U8028 ( .INP(n8282), .Z(n8196) );
  NBUFFX2 U8029 ( .INP(n8282), .Z(n8195) );
  NBUFFX2 U8030 ( .INP(n8283), .Z(n8194) );
  NBUFFX2 U8031 ( .INP(n8283), .Z(n8193) );
  NBUFFX2 U8032 ( .INP(n8283), .Z(n8192) );
  NBUFFX2 U8033 ( .INP(n8284), .Z(n8191) );
  NBUFFX2 U8034 ( .INP(n8284), .Z(n8190) );
  NBUFFX2 U8035 ( .INP(n8284), .Z(n8189) );
  NBUFFX2 U8036 ( .INP(n8285), .Z(n8188) );
  NBUFFX2 U8037 ( .INP(n8286), .Z(n8184) );
  NBUFFX2 U8038 ( .INP(n8286), .Z(n8183) );
  NBUFFX2 U8039 ( .INP(n8286), .Z(n8185) );
  NBUFFX2 U8040 ( .INP(n8288), .Z(n8177) );
  NBUFFX2 U8041 ( .INP(n8287), .Z(n8181) );
  NBUFFX2 U8042 ( .INP(n8287), .Z(n8182) );
  NBUFFX2 U8043 ( .INP(n8285), .Z(n8187) );
  NBUFFX2 U8044 ( .INP(n8285), .Z(n8186) );
  NBUFFX2 U8045 ( .INP(n8288), .Z(n8178) );
  NBUFFX2 U8046 ( .INP(n8287), .Z(n8180) );
  NBUFFX2 U8047 ( .INP(n8288), .Z(n8179) );
  NBUFFX2 U8048 ( .INP(n8289), .Z(n8176) );
  NBUFFX2 U8049 ( .INP(n8289), .Z(n8175) );
  NBUFFX2 U8050 ( .INP(n8289), .Z(n8174) );
  NBUFFX2 U8051 ( .INP(n8290), .Z(n8173) );
  NBUFFX2 U8052 ( .INP(n8290), .Z(n8172) );
  NBUFFX2 U8053 ( .INP(n8292), .Z(n8167) );
  NBUFFX2 U8054 ( .INP(n8290), .Z(n8171) );
  NBUFFX2 U8055 ( .INP(n8291), .Z(n8170) );
  NBUFFX2 U8056 ( .INP(n8291), .Z(n8169) );
  NBUFFX2 U8057 ( .INP(n8291), .Z(n8168) );
  NBUFFX2 U8058 ( .INP(n8293), .Z(n8162) );
  NBUFFX2 U8059 ( .INP(n8294), .Z(n8161) );
  NBUFFX2 U8060 ( .INP(n8294), .Z(n8160) );
  NBUFFX2 U8061 ( .INP(n8292), .Z(n8166) );
  NBUFFX2 U8062 ( .INP(n8292), .Z(n8165) );
  NBUFFX2 U8063 ( .INP(n8294), .Z(n8159) );
  NBUFFX2 U8064 ( .INP(n8295), .Z(n8158) );
  NBUFFX2 U8065 ( .INP(n8295), .Z(n8157) );
  NBUFFX2 U8066 ( .INP(n8299), .Z(n8144) );
  NBUFFX2 U8067 ( .INP(n8293), .Z(n8163) );
  NBUFFX2 U8068 ( .INP(n8297), .Z(n8152) );
  NBUFFX2 U8069 ( .INP(n8296), .Z(n8153) );
  NBUFFX2 U8070 ( .INP(n8299), .Z(n8146) );
  NBUFFX2 U8071 ( .INP(n8296), .Z(n8154) );
  NBUFFX2 U8072 ( .INP(n8297), .Z(n8151) );
  NBUFFX2 U8073 ( .INP(n8295), .Z(n8156) );
  NBUFFX2 U8074 ( .INP(n8296), .Z(n8155) );
  NBUFFX2 U8075 ( .INP(n8298), .Z(n8147) );
  NBUFFX2 U8076 ( .INP(n8299), .Z(n8145) );
  NBUFFX2 U8077 ( .INP(n8298), .Z(n8148) );
  NBUFFX2 U8078 ( .INP(n8297), .Z(n8150) );
  NBUFFX2 U8079 ( .INP(n8298), .Z(n8149) );
  NBUFFX2 U8080 ( .INP(n8302), .Z(n8137) );
  NBUFFX2 U8081 ( .INP(n8302), .Z(n8136) );
  NBUFFX2 U8082 ( .INP(n8261), .Z(n8258) );
  NBUFFX2 U8083 ( .INP(n8302), .Z(n8135) );
  NBUFFX2 U8084 ( .INP(n8261), .Z(n8259) );
  NBUFFX2 U8085 ( .INP(n8262), .Z(n8257) );
  NBUFFX2 U8086 ( .INP(n8262), .Z(n8256) );
  NBUFFX2 U8087 ( .INP(n8293), .Z(n8164) );
  NBUFFX2 U8088 ( .INP(n8300), .Z(n8142) );
  NBUFFX2 U8089 ( .INP(n8300), .Z(n8141) );
  NBUFFX2 U8090 ( .INP(n8301), .Z(n8140) );
  NBUFFX2 U8091 ( .INP(n8301), .Z(n8139) );
  NBUFFX2 U8092 ( .INP(n8301), .Z(n8138) );
  NBUFFX2 U8093 ( .INP(n8303), .Z(n8132) );
  NBUFFX2 U8094 ( .INP(n8303), .Z(n8134) );
  NBUFFX2 U8095 ( .INP(n8303), .Z(n8133) );
  NBUFFX2 U8096 ( .INP(n8491), .Z(n8317) );
  NBUFFX2 U8097 ( .INP(n8491), .Z(n8318) );
  NBUFFX2 U8098 ( .INP(n8452), .Z(n8434) );
  NBUFFX2 U8099 ( .INP(n8449), .Z(n8442) );
  NBUFFX2 U8100 ( .INP(n8450), .Z(n8441) );
  NBUFFX2 U8101 ( .INP(n8450), .Z(n8440) );
  NBUFFX2 U8102 ( .INP(n8450), .Z(n8439) );
  NBUFFX2 U8103 ( .INP(n8451), .Z(n8438) );
  NBUFFX2 U8104 ( .INP(n8452), .Z(n8435) );
  NBUFFX2 U8105 ( .INP(n8451), .Z(n8437) );
  NBUFFX2 U8106 ( .INP(n8451), .Z(n8436) );
  NBUFFX2 U8107 ( .INP(n8455), .Z(n8425) );
  NBUFFX2 U8108 ( .INP(n8455), .Z(n8426) );
  NBUFFX2 U8109 ( .INP(n8453), .Z(n8432) );
  NBUFFX2 U8110 ( .INP(n8452), .Z(n8433) );
  NBUFFX2 U8111 ( .INP(n8487), .Z(n8330) );
  NBUFFX2 U8112 ( .INP(n8454), .Z(n8427) );
  NBUFFX2 U8113 ( .INP(n8455), .Z(n8424) );
  NBUFFX2 U8114 ( .INP(n8454), .Z(n8428) );
  NBUFFX2 U8115 ( .INP(n8457), .Z(n8418) );
  NBUFFX2 U8116 ( .INP(n8454), .Z(n8429) );
  NBUFFX2 U8117 ( .INP(n8456), .Z(n8423) );
  NBUFFX2 U8118 ( .INP(n8453), .Z(n8431) );
  NBUFFX2 U8119 ( .INP(n8453), .Z(n8430) );
  NBUFFX2 U8120 ( .INP(n8457), .Z(n8420) );
  NBUFFX2 U8121 ( .INP(n8457), .Z(n8419) );
  NBUFFX2 U8122 ( .INP(n8456), .Z(n8422) );
  NBUFFX2 U8123 ( .INP(n8456), .Z(n8421) );
  NBUFFX2 U8124 ( .INP(n8458), .Z(n8417) );
  NBUFFX2 U8125 ( .INP(n8458), .Z(n8416) );
  NBUFFX2 U8126 ( .INP(n8458), .Z(n8415) );
  NBUFFX2 U8127 ( .INP(n8459), .Z(n8414) );
  NBUFFX2 U8128 ( .INP(n8462), .Z(n8405) );
  NBUFFX2 U8129 ( .INP(n8459), .Z(n8413) );
  NBUFFX2 U8130 ( .INP(n8460), .Z(n8410) );
  NBUFFX2 U8131 ( .INP(n8459), .Z(n8412) );
  NBUFFX2 U8132 ( .INP(n8460), .Z(n8411) );
  NBUFFX2 U8133 ( .INP(n8460), .Z(n8409) );
  NBUFFX2 U8134 ( .INP(n8461), .Z(n8408) );
  NBUFFX2 U8135 ( .INP(n8461), .Z(n8407) );
  NBUFFX2 U8136 ( .INP(n8461), .Z(n8406) );
  NBUFFX2 U8137 ( .INP(n8462), .Z(n8404) );
  NBUFFX2 U8138 ( .INP(n8462), .Z(n8403) );
  NBUFFX2 U8139 ( .INP(n8463), .Z(n8402) );
  NBUFFX2 U8140 ( .INP(n8463), .Z(n8401) );
  NBUFFX2 U8141 ( .INP(n8464), .Z(n8397) );
  NBUFFX2 U8142 ( .INP(n8464), .Z(n8398) );
  NBUFFX2 U8143 ( .INP(n8466), .Z(n8391) );
  NBUFFX2 U8144 ( .INP(n8465), .Z(n8396) );
  NBUFFX2 U8145 ( .INP(n8465), .Z(n8395) );
  NBUFFX2 U8146 ( .INP(n8463), .Z(n8400) );
  NBUFFX2 U8147 ( .INP(n8464), .Z(n8399) );
  NBUFFX2 U8148 ( .INP(n8465), .Z(n8394) );
  NBUFFX2 U8149 ( .INP(n8466), .Z(n8393) );
  NBUFFX2 U8150 ( .INP(n8466), .Z(n8392) );
  NBUFFX2 U8151 ( .INP(n8467), .Z(n8390) );
  NBUFFX2 U8152 ( .INP(n8467), .Z(n8389) );
  NBUFFX2 U8153 ( .INP(n8467), .Z(n8388) );
  NBUFFX2 U8154 ( .INP(n8468), .Z(n8387) );
  NBUFFX2 U8155 ( .INP(n8468), .Z(n8386) );
  NBUFFX2 U8156 ( .INP(n8468), .Z(n8385) );
  NBUFFX2 U8157 ( .INP(n8469), .Z(n8384) );
  NBUFFX2 U8158 ( .INP(n8469), .Z(n8383) );
  NBUFFX2 U8159 ( .INP(n8469), .Z(n8382) );
  NBUFFX2 U8160 ( .INP(n8470), .Z(n8381) );
  NBUFFX2 U8161 ( .INP(n8470), .Z(n8380) );
  NBUFFX2 U8162 ( .INP(n8470), .Z(n8379) );
  NBUFFX2 U8163 ( .INP(n8471), .Z(n8378) );
  NBUFFX2 U8164 ( .INP(n8471), .Z(n8377) );
  NBUFFX2 U8165 ( .INP(n8471), .Z(n8376) );
  NBUFFX2 U8166 ( .INP(n8472), .Z(n8375) );
  NBUFFX2 U8167 ( .INP(n8473), .Z(n8371) );
  NBUFFX2 U8168 ( .INP(n8473), .Z(n8370) );
  NBUFFX2 U8169 ( .INP(n8473), .Z(n8372) );
  NBUFFX2 U8170 ( .INP(n8475), .Z(n8364) );
  NBUFFX2 U8171 ( .INP(n8474), .Z(n8368) );
  NBUFFX2 U8172 ( .INP(n8474), .Z(n8369) );
  NBUFFX2 U8173 ( .INP(n8472), .Z(n8374) );
  NBUFFX2 U8174 ( .INP(n8472), .Z(n8373) );
  NBUFFX2 U8175 ( .INP(n8475), .Z(n8365) );
  NBUFFX2 U8176 ( .INP(n8474), .Z(n8367) );
  NBUFFX2 U8177 ( .INP(n8475), .Z(n8366) );
  NBUFFX2 U8178 ( .INP(n8476), .Z(n8363) );
  NBUFFX2 U8179 ( .INP(n8476), .Z(n8362) );
  NBUFFX2 U8180 ( .INP(n8476), .Z(n8361) );
  NBUFFX2 U8181 ( .INP(n8477), .Z(n8360) );
  NBUFFX2 U8182 ( .INP(n8477), .Z(n8359) );
  NBUFFX2 U8183 ( .INP(n8479), .Z(n8354) );
  NBUFFX2 U8184 ( .INP(n8477), .Z(n8358) );
  NBUFFX2 U8185 ( .INP(n8478), .Z(n8357) );
  NBUFFX2 U8186 ( .INP(n8478), .Z(n8356) );
  NBUFFX2 U8187 ( .INP(n8478), .Z(n8355) );
  NBUFFX2 U8188 ( .INP(n8480), .Z(n8349) );
  NBUFFX2 U8189 ( .INP(n8481), .Z(n8348) );
  NBUFFX2 U8190 ( .INP(n8481), .Z(n8347) );
  NBUFFX2 U8191 ( .INP(n8479), .Z(n8353) );
  NBUFFX2 U8192 ( .INP(n8479), .Z(n8352) );
  NBUFFX2 U8193 ( .INP(n8481), .Z(n8346) );
  NBUFFX2 U8194 ( .INP(n8482), .Z(n8345) );
  NBUFFX2 U8195 ( .INP(n8482), .Z(n8344) );
  NBUFFX2 U8196 ( .INP(n8486), .Z(n8331) );
  NBUFFX2 U8197 ( .INP(n8480), .Z(n8350) );
  NBUFFX2 U8198 ( .INP(n8484), .Z(n8339) );
  NBUFFX2 U8199 ( .INP(n8483), .Z(n8340) );
  NBUFFX2 U8200 ( .INP(n8486), .Z(n8333) );
  NBUFFX2 U8201 ( .INP(n8483), .Z(n8341) );
  NBUFFX2 U8202 ( .INP(n8484), .Z(n8338) );
  NBUFFX2 U8203 ( .INP(n8482), .Z(n8343) );
  NBUFFX2 U8204 ( .INP(n8483), .Z(n8342) );
  NBUFFX2 U8205 ( .INP(n8485), .Z(n8334) );
  NBUFFX2 U8206 ( .INP(n8486), .Z(n8332) );
  NBUFFX2 U8207 ( .INP(n8485), .Z(n8335) );
  NBUFFX2 U8208 ( .INP(n8484), .Z(n8337) );
  NBUFFX2 U8209 ( .INP(n8485), .Z(n8336) );
  NBUFFX2 U8210 ( .INP(n8489), .Z(n8324) );
  NBUFFX2 U8211 ( .INP(n8489), .Z(n8323) );
  NBUFFX2 U8212 ( .INP(n8448), .Z(n8445) );
  NBUFFX2 U8213 ( .INP(n8489), .Z(n8322) );
  NBUFFX2 U8214 ( .INP(n8448), .Z(n8446) );
  NBUFFX2 U8215 ( .INP(n8449), .Z(n8444) );
  NBUFFX2 U8216 ( .INP(n8449), .Z(n8443) );
  NBUFFX2 U8217 ( .INP(n8480), .Z(n8351) );
  NBUFFX2 U8218 ( .INP(n8487), .Z(n8329) );
  NBUFFX2 U8219 ( .INP(n8487), .Z(n8328) );
  NBUFFX2 U8220 ( .INP(n8488), .Z(n8327) );
  NBUFFX2 U8221 ( .INP(n8488), .Z(n8326) );
  NBUFFX2 U8222 ( .INP(n8488), .Z(n8325) );
  NBUFFX2 U8223 ( .INP(n8490), .Z(n8319) );
  NBUFFX2 U8224 ( .INP(n8490), .Z(n8321) );
  NBUFFX2 U8225 ( .INP(n8490), .Z(n8320) );
  NBUFFX2 U8226 ( .INP(n8261), .Z(n8260) );
  NBUFFX2 U8227 ( .INP(n8448), .Z(n8447) );
  NBUFFX2 U8228 ( .INP(n8500), .Z(n8450) );
  NBUFFX2 U8229 ( .INP(n8313), .Z(n8263) );
  NBUFFX2 U8230 ( .INP(n8500), .Z(n8451) );
  NBUFFX2 U8231 ( .INP(n8313), .Z(n8264) );
  NBUFFX2 U8232 ( .INP(n8500), .Z(n8448) );
  NBUFFX2 U8233 ( .INP(n8313), .Z(n8261) );
  NBUFFX2 U8234 ( .INP(n8500), .Z(n8449) );
  NBUFFX2 U8235 ( .INP(n8313), .Z(n8262) );
  NBUFFX2 U8236 ( .INP(n8499), .Z(n8452) );
  NBUFFX2 U8237 ( .INP(n8312), .Z(n8265) );
  NBUFFX2 U8238 ( .INP(n8499), .Z(n8455) );
  NBUFFX2 U8239 ( .INP(n8312), .Z(n8268) );
  NBUFFX2 U8240 ( .INP(n8499), .Z(n8454) );
  NBUFFX2 U8241 ( .INP(n8312), .Z(n8267) );
  NBUFFX2 U8242 ( .INP(n8499), .Z(n8453) );
  NBUFFX2 U8243 ( .INP(n8312), .Z(n8266) );
  NBUFFX2 U8244 ( .INP(n8498), .Z(n8457) );
  NBUFFX2 U8245 ( .INP(n8311), .Z(n8270) );
  NBUFFX2 U8246 ( .INP(n8499), .Z(n8456) );
  NBUFFX2 U8247 ( .INP(n8312), .Z(n8269) );
  NBUFFX2 U8248 ( .INP(n8498), .Z(n8458) );
  NBUFFX2 U8249 ( .INP(n8311), .Z(n8271) );
  NBUFFX2 U8250 ( .INP(n8498), .Z(n8459) );
  NBUFFX2 U8251 ( .INP(n8311), .Z(n8272) );
  NBUFFX2 U8252 ( .INP(n8498), .Z(n8460) );
  NBUFFX2 U8253 ( .INP(n8311), .Z(n8273) );
  NBUFFX2 U8254 ( .INP(n8498), .Z(n8461) );
  NBUFFX2 U8255 ( .INP(n8311), .Z(n8274) );
  NBUFFX2 U8256 ( .INP(n8497), .Z(n8462) );
  NBUFFX2 U8257 ( .INP(n8310), .Z(n8275) );
  NBUFFX2 U8258 ( .INP(n8497), .Z(n8463) );
  NBUFFX2 U8259 ( .INP(n8310), .Z(n8276) );
  NBUFFX2 U8260 ( .INP(n8497), .Z(n8464) );
  NBUFFX2 U8261 ( .INP(n8310), .Z(n8277) );
  NBUFFX2 U8262 ( .INP(n8497), .Z(n8465) );
  NBUFFX2 U8263 ( .INP(n8310), .Z(n8278) );
  NBUFFX2 U8264 ( .INP(n8497), .Z(n8466) );
  NBUFFX2 U8265 ( .INP(n8310), .Z(n8279) );
  NBUFFX2 U8266 ( .INP(n8496), .Z(n8467) );
  NBUFFX2 U8267 ( .INP(n8309), .Z(n8280) );
  NBUFFX2 U8268 ( .INP(n8496), .Z(n8468) );
  NBUFFX2 U8269 ( .INP(n8309), .Z(n8281) );
  NBUFFX2 U8270 ( .INP(n8496), .Z(n8469) );
  NBUFFX2 U8271 ( .INP(n8309), .Z(n8282) );
  NBUFFX2 U8272 ( .INP(n8496), .Z(n8470) );
  NBUFFX2 U8273 ( .INP(n8309), .Z(n8283) );
  NBUFFX2 U8274 ( .INP(n8496), .Z(n8471) );
  NBUFFX2 U8275 ( .INP(n8309), .Z(n8284) );
  NBUFFX2 U8276 ( .INP(n8495), .Z(n8473) );
  NBUFFX2 U8277 ( .INP(n8308), .Z(n8286) );
  NBUFFX2 U8278 ( .INP(n8495), .Z(n8472) );
  NBUFFX2 U8279 ( .INP(n8308), .Z(n8285) );
  NBUFFX2 U8280 ( .INP(n8495), .Z(n8474) );
  NBUFFX2 U8281 ( .INP(n8308), .Z(n8287) );
  NBUFFX2 U8282 ( .INP(n8495), .Z(n8475) );
  NBUFFX2 U8283 ( .INP(n8308), .Z(n8288) );
  NBUFFX2 U8284 ( .INP(n8495), .Z(n8476) );
  NBUFFX2 U8285 ( .INP(n8308), .Z(n8289) );
  NBUFFX2 U8286 ( .INP(n8494), .Z(n8477) );
  NBUFFX2 U8287 ( .INP(n8307), .Z(n8290) );
  NBUFFX2 U8288 ( .INP(n8494), .Z(n8478) );
  NBUFFX2 U8289 ( .INP(n8307), .Z(n8291) );
  NBUFFX2 U8290 ( .INP(n8494), .Z(n8479) );
  NBUFFX2 U8291 ( .INP(n8307), .Z(n8292) );
  NBUFFX2 U8292 ( .INP(n8494), .Z(n8481) );
  NBUFFX2 U8293 ( .INP(n8307), .Z(n8294) );
  NBUFFX2 U8294 ( .INP(n8493), .Z(n8482) );
  NBUFFX2 U8295 ( .INP(n8306), .Z(n8295) );
  NBUFFX2 U8296 ( .INP(n8493), .Z(n8483) );
  NBUFFX2 U8297 ( .INP(n8306), .Z(n8296) );
  NBUFFX2 U8298 ( .INP(n8493), .Z(n8486) );
  NBUFFX2 U8299 ( .INP(n8306), .Z(n8299) );
  NBUFFX2 U8300 ( .INP(n8493), .Z(n8484) );
  NBUFFX2 U8301 ( .INP(n8306), .Z(n8297) );
  NBUFFX2 U8302 ( .INP(n8493), .Z(n8485) );
  NBUFFX2 U8303 ( .INP(n8306), .Z(n8298) );
  NBUFFX2 U8304 ( .INP(n8492), .Z(n8489) );
  NBUFFX2 U8305 ( .INP(n8305), .Z(n8302) );
  NBUFFX2 U8306 ( .INP(n8494), .Z(n8480) );
  NBUFFX2 U8307 ( .INP(n8307), .Z(n8293) );
  NBUFFX2 U8308 ( .INP(n8492), .Z(n8487) );
  NBUFFX2 U8309 ( .INP(n8305), .Z(n8300) );
  NBUFFX2 U8310 ( .INP(n8492), .Z(n8488) );
  NBUFFX2 U8311 ( .INP(n8305), .Z(n8301) );
  NBUFFX2 U8312 ( .INP(n8492), .Z(n8490) );
  NBUFFX2 U8313 ( .INP(n8305), .Z(n8303) );
  NBUFFX2 U8314 ( .INP(n8492), .Z(n8491) );
  NBUFFX2 U8315 ( .INP(n8305), .Z(n8304) );
  NBUFFX2 U8316 ( .INP(n8316), .Z(n8305) );
  NBUFFX2 U8317 ( .INP(n8316), .Z(n8306) );
  NBUFFX2 U8318 ( .INP(n8316), .Z(n8307) );
  NBUFFX2 U8319 ( .INP(n8315), .Z(n8308) );
  NBUFFX2 U8320 ( .INP(n8315), .Z(n8309) );
  NBUFFX2 U8321 ( .INP(n8315), .Z(n8310) );
  NBUFFX2 U8322 ( .INP(n8314), .Z(n8311) );
  NBUFFX2 U8323 ( .INP(n8314), .Z(n8312) );
  NBUFFX2 U8324 ( .INP(n8314), .Z(n8313) );
  NBUFFX2 U8325 ( .INP(test_se), .Z(n8314) );
  NBUFFX2 U8326 ( .INP(test_se), .Z(n8315) );
  NBUFFX2 U8327 ( .INP(test_se), .Z(n8316) );
  NBUFFX2 U8328 ( .INP(n8503), .Z(n8492) );
  NBUFFX2 U8329 ( .INP(n8503), .Z(n8493) );
  NBUFFX2 U8330 ( .INP(n8503), .Z(n8494) );
  NBUFFX2 U8331 ( .INP(n8502), .Z(n8495) );
  NBUFFX2 U8332 ( .INP(n8502), .Z(n8496) );
  NBUFFX2 U8333 ( .INP(n8502), .Z(n8497) );
  NBUFFX2 U8334 ( .INP(n8501), .Z(n8498) );
  NBUFFX2 U8335 ( .INP(n8501), .Z(n8499) );
  NBUFFX2 U8336 ( .INP(n8501), .Z(n8500) );
  NBUFFX2 U8337 ( .INP(CK), .Z(n8501) );
  NBUFFX2 U8338 ( .INP(CK), .Z(n8502) );
  NBUFFX2 U8339 ( .INP(CK), .Z(n8503) );
  INVX0 U8340 ( .INP(n8504), .ZN(n959) );
  INVX0 U8341 ( .INP(g27380), .ZN(n91) );
  INVX0 U8342 ( .INP(n8505), .ZN(n902) );
  NAND3X0 U8343 ( .IN1(n8506), .IN2(n8507), .IN3(n8508), .QN(n8505) );
  NAND2X0 U8344 ( .IN1(n8509), .IN2(n4411), .QN(n8506) );
  NAND2X0 U8345 ( .IN1(g1346), .IN2(n8510), .QN(n8509) );
  NOR3X0 U8346 ( .IN1(n8511), .IN2(n8512), .IN3(n8513), .QN(n901) );
  NOR2X0 U8347 ( .IN1(n8514), .IN2(g1319), .QN(n8511) );
  NOR2X0 U8348 ( .IN1(n4402), .IN2(n8515), .QN(n8514) );
  NOR2X0 U8349 ( .IN1(n8512), .IN2(n8516), .QN(n872) );
  INVX0 U8350 ( .INP(n8517), .ZN(n8516) );
  NAND2X0 U8351 ( .IN1(n8518), .IN2(n7955), .QN(n8517) );
  INVX0 U8352 ( .INP(n8519), .ZN(n826) );
  NOR2X0 U8353 ( .IN1(n8520), .IN2(n8521), .QN(n8519) );
  NOR2X0 U8354 ( .IN1(g1236), .IN2(n7970), .QN(n8521) );
  INVX0 U8355 ( .INP(n8522), .ZN(n822) );
  INVX0 U8356 ( .INP(n8523), .ZN(n808) );
  INVX0 U8357 ( .INP(n8524), .ZN(n653) );
  INVX0 U8358 ( .INP(n8525), .ZN(n597) );
  NAND3X0 U8359 ( .IN1(n8526), .IN2(n8527), .IN3(n8528), .QN(n8525) );
  NAND2X0 U8360 ( .IN1(n8529), .IN2(n4413), .QN(n8526) );
  NAND2X0 U8361 ( .IN1(g660), .IN2(n8530), .QN(n8529) );
  INVX0 U8362 ( .INP(n8531), .ZN(n596) );
  NAND3X0 U8363 ( .IN1(n8532), .IN2(n8527), .IN3(n8533), .QN(n8531) );
  NAND2X0 U8364 ( .IN1(n8534), .IN2(n4478), .QN(n8532) );
  NAND2X0 U8365 ( .IN1(g640), .IN2(n8535), .QN(n8534) );
  NOR2X0 U8366 ( .IN1(n8536), .IN2(n8537), .QN(n567) );
  INVX0 U8367 ( .INP(n8538), .ZN(n8537) );
  NAND2X0 U8368 ( .IN1(n8539), .IN2(n7956), .QN(n8538) );
  INVX0 U8369 ( .INP(n8540), .ZN(n520) );
  NOR2X0 U8370 ( .IN1(n8541), .IN2(n8542), .QN(n8540) );
  NOR2X0 U8371 ( .IN1(g550), .IN2(n7972), .QN(n8542) );
  INVX0 U8372 ( .INP(n8543), .ZN(n515) );
  INVX0 U8373 ( .INP(n8544), .ZN(n514) );
  INVX0 U8374 ( .INP(n8545), .ZN(n513) );
  INVX0 U8375 ( .INP(n8546), .ZN(n499) );
  INVX0 U8376 ( .INP(n8547), .ZN(n475) );
  INVX0 U8377 ( .INP(n8548), .ZN(n453) );
  XNOR2X1 U8378 ( .IN1(n8012), .IN2(n8549), .Q(n4281) );
  XOR2X1 U8379 ( .IN1(n8550), .IN2(n8014), .Q(n4280) );
  NAND2X0 U8380 ( .IN1(g2879), .IN2(n8551), .QN(n4279) );
  NAND2X0 U8381 ( .IN1(DFF_18_n1), .IN2(g8021), .QN(n8551) );
  NOR2X0 U8382 ( .IN1(n8552), .IN2(n8553), .QN(n4278) );
  NOR2X0 U8383 ( .IN1(n2568), .IN2(n8554), .QN(n8553) );
  INVX0 U8384 ( .INP(n8555), .ZN(n8554) );
  NOR4X0 U8385 ( .IN1(n8556), .IN2(n8557), .IN3(n8558), .IN4(n8559), .QN(n8552) );
  NAND3X0 U8386 ( .IN1(n8560), .IN2(n8561), .IN3(n8562), .QN(n8559) );
  XOR2X1 U8387 ( .IN1(n7164), .IN2(n8563), .Q(n8562) );
  XOR2X1 U8388 ( .IN1(n8067), .IN2(n8564), .Q(n8561) );
  XOR2X1 U8389 ( .IN1(n8048), .IN2(n8565), .Q(n8560) );
  NAND3X0 U8390 ( .IN1(n8566), .IN2(n8567), .IN3(n8568), .QN(n8558) );
  XOR2X1 U8391 ( .IN1(n7699), .IN2(n8569), .Q(n8568) );
  XOR2X1 U8392 ( .IN1(g88), .IN2(n8570), .Q(n8567) );
  XOR2X1 U8393 ( .IN1(n7325), .IN2(n8571), .Q(n8566) );
  NAND3X0 U8394 ( .IN1(n8572), .IN2(n8573), .IN3(n8574), .QN(n8557) );
  XOR2X1 U8395 ( .IN1(n7700), .IN2(n8575), .Q(n8574) );
  XOR2X1 U8396 ( .IN1(n7701), .IN2(n8576), .Q(n8573) );
  XOR2X1 U8397 ( .IN1(n7702), .IN2(n8577), .Q(n8572) );
  NAND3X0 U8398 ( .IN1(n8578), .IN2(n8579), .IN3(n8580), .QN(n8556) );
  XOR2X1 U8399 ( .IN1(test_so15), .IN2(n8581), .Q(n8580) );
  NOR2X0 U8400 ( .IN1(n8582), .IN2(n8583), .QN(n4277) );
  NOR2X0 U8401 ( .IN1(n8584), .IN2(n8585), .QN(n8583) );
  NOR4X0 U8402 ( .IN1(n8586), .IN2(n8587), .IN3(n8588), .IN4(n8589), .QN(n8582) );
  NAND3X0 U8403 ( .IN1(n8590), .IN2(n8591), .IN3(n8592), .QN(n8589) );
  XOR2X1 U8404 ( .IN1(n8593), .IN2(n8054), .Q(n8592) );
  XOR2X1 U8405 ( .IN1(n8594), .IN2(n7695), .Q(n8591) );
  XOR2X1 U8406 ( .IN1(n8595), .IN2(n8063), .Q(n8590) );
  NAND3X0 U8407 ( .IN1(n8596), .IN2(n8597), .IN3(n8598), .QN(n8588) );
  XOR2X1 U8408 ( .IN1(n8599), .IN2(n7697), .Q(n8598) );
  XOR2X1 U8409 ( .IN1(n8600), .IN2(n7698), .Q(n8597) );
  XOR2X1 U8410 ( .IN1(n8601), .IN2(n8064), .Q(n8596) );
  NAND3X0 U8411 ( .IN1(n8602), .IN2(n8603), .IN3(n8604), .QN(n8587) );
  XOR2X1 U8412 ( .IN1(n8605), .IN2(n7163), .Q(n8604) );
  XOR2X1 U8413 ( .IN1(n8606), .IN2(n7696), .Q(n8603) );
  XOR2X1 U8414 ( .IN1(n8607), .IN2(n7324), .Q(n8602) );
  NAND3X0 U8415 ( .IN1(n8608), .IN2(n8578), .IN3(n8609), .QN(n8586) );
  XNOR2X1 U8416 ( .IN1(test_so36), .IN2(n8610), .Q(n8609) );
  NOR2X0 U8417 ( .IN1(n8611), .IN2(n8612), .QN(n4276) );
  NOR2X0 U8418 ( .IN1(n8613), .IN2(n8614), .QN(n8612) );
  INVX0 U8419 ( .INP(n8615), .ZN(n8614) );
  NOR2X0 U8420 ( .IN1(n8616), .IN2(n8617), .QN(n8611) );
  NAND4X0 U8421 ( .IN1(n8618), .IN2(n8619), .IN3(n8620), .IN4(n8621), .QN(
        n8617) );
  NOR3X0 U8422 ( .IN1(n8622), .IN2(n8623), .IN3(n8624), .QN(n8621) );
  XOR2X1 U8423 ( .IN1(n7691), .IN2(n8625), .Q(n8624) );
  XOR2X1 U8424 ( .IN1(n8049), .IN2(n8626), .Q(n8623) );
  XOR2X1 U8425 ( .IN1(n8042), .IN2(n8627), .Q(n8622) );
  XOR2X1 U8426 ( .IN1(g1453), .IN2(n8628), .Q(n8620) );
  XOR2X1 U8427 ( .IN1(n8068), .IN2(n8629), .Q(n8619) );
  XOR2X1 U8428 ( .IN1(n7162), .IN2(n8630), .Q(n8618) );
  NAND4X0 U8429 ( .IN1(n8631), .IN2(n8578), .IN3(n8632), .IN4(n8633), .QN(
        n8616) );
  NOR3X0 U8430 ( .IN1(n8634), .IN2(n8635), .IN3(n8636), .QN(n8633) );
  XNOR2X1 U8431 ( .IN1(n7693), .IN2(n8637), .Q(n8636) );
  XNOR2X1 U8432 ( .IN1(n7694), .IN2(n8638), .Q(n8635) );
  XOR2X1 U8433 ( .IN1(n7323), .IN2(n8639), .Q(n8634) );
  XOR2X1 U8434 ( .IN1(n7692), .IN2(n8640), .Q(n8632) );
  NOR2X0 U8435 ( .IN1(n8641), .IN2(n8642), .QN(n4275) );
  NOR2X0 U8436 ( .IN1(n8643), .IN2(n8644), .QN(n8642) );
  NOR4X0 U8437 ( .IN1(n8645), .IN2(n8646), .IN3(n8647), .IN4(n8648), .QN(n8641) );
  NAND3X0 U8438 ( .IN1(n8649), .IN2(n8650), .IN3(n8651), .QN(n8648) );
  XOR2X1 U8439 ( .IN1(n8652), .IN2(n8053), .Q(n8651) );
  XOR2X1 U8440 ( .IN1(n8653), .IN2(n8069), .Q(n8650) );
  XOR2X1 U8441 ( .IN1(n8654), .IN2(n7161), .Q(n8649) );
  NAND3X0 U8442 ( .IN1(n8655), .IN2(n8656), .IN3(n8657), .QN(n8647) );
  XOR2X1 U8443 ( .IN1(n8658), .IN2(n7687), .Q(n8657) );
  XOR2X1 U8444 ( .IN1(n8659), .IN2(n8050), .Q(n8656) );
  XOR2X1 U8445 ( .IN1(n8660), .IN2(n7690), .Q(n8655) );
  NAND3X0 U8446 ( .IN1(n8661), .IN2(n8662), .IN3(n8663), .QN(n8646) );
  XOR2X1 U8447 ( .IN1(n8664), .IN2(n7689), .Q(n8663) );
  XOR2X1 U8448 ( .IN1(n8665), .IN2(n7322), .Q(n8662) );
  XOR2X1 U8449 ( .IN1(n8666), .IN2(n7688), .Q(n8661) );
  NAND3X0 U8450 ( .IN1(n8667), .IN2(n8578), .IN3(n8668), .QN(n8645) );
  XOR2X1 U8451 ( .IN1(test_so78), .IN2(n8669), .Q(n8668) );
  NAND2X0 U8452 ( .IN1(n8670), .IN2(n8671), .QN(n4274) );
  INVX0 U8453 ( .INP(n8672), .ZN(n8671) );
  XNOR2X1 U8454 ( .IN1(n4330), .IN2(n4423), .Q(n8670) );
  NAND2X0 U8455 ( .IN1(n8673), .IN2(n8674), .QN(n4273) );
  NAND2X0 U8456 ( .IN1(n8675), .IN2(n8676), .QN(n8674) );
  NAND2X0 U8457 ( .IN1(n4482), .IN2(n8677), .QN(n8675) );
  NAND2X0 U8458 ( .IN1(n2426), .IN2(n8678), .QN(n4272) );
  NAND3X0 U8459 ( .IN1(n8679), .IN2(n8680), .IN3(n8681), .QN(n8678) );
  NAND2X0 U8460 ( .IN1(n8682), .IN2(n8683), .QN(n8680) );
  INVX0 U8461 ( .INP(n8684), .ZN(n8682) );
  NAND2X0 U8462 ( .IN1(n8685), .IN2(DFF_449_n1), .QN(n8679) );
  NAND2X0 U8463 ( .IN1(n8686), .IN2(n8687), .QN(n4271) );
  NAND2X0 U8464 ( .IN1(n2446), .IN2(n8688), .QN(n8687) );
  NAND3X0 U8465 ( .IN1(n8689), .IN2(n8690), .IN3(n8681), .QN(n8686) );
  NAND2X0 U8466 ( .IN1(n8691), .IN2(n8683), .QN(n8690) );
  INVX0 U8467 ( .INP(n8692), .ZN(n8691) );
  NAND2X0 U8468 ( .IN1(n7143), .IN2(n8685), .QN(n8689) );
  NAND2X0 U8469 ( .IN1(n8693), .IN2(n8694), .QN(n4270) );
  NAND2X0 U8470 ( .IN1(n2446), .IN2(n8695), .QN(n8694) );
  NAND3X0 U8471 ( .IN1(n8696), .IN2(n8697), .IN3(n8681), .QN(n8693) );
  NAND2X0 U8472 ( .IN1(n8698), .IN2(n8683), .QN(n8697) );
  NAND2X0 U8473 ( .IN1(n7142), .IN2(n8685), .QN(n8696) );
  NAND2X0 U8474 ( .IN1(n8699), .IN2(n8700), .QN(n4269) );
  NAND3X0 U8475 ( .IN1(n8701), .IN2(n8702), .IN3(n8681), .QN(n8700) );
  NAND2X0 U8476 ( .IN1(n8703), .IN2(n8683), .QN(n8702) );
  INVX0 U8477 ( .INP(n8704), .ZN(n8703) );
  NAND2X0 U8478 ( .IN1(n8685), .IN2(DFF_444_n1), .QN(n8701) );
  NAND3X0 U8479 ( .IN1(n2426), .IN2(n8705), .IN3(n2440), .QN(n4268) );
  NAND3X0 U8480 ( .IN1(n8706), .IN2(n8707), .IN3(n8681), .QN(n8705) );
  NAND2X0 U8481 ( .IN1(n8708), .IN2(n8683), .QN(n8707) );
  INVX0 U8482 ( .INP(n8709), .ZN(n8708) );
  NAND2X0 U8483 ( .IN1(n8685), .IN2(DFF_445_n1), .QN(n8706) );
  NAND3X0 U8484 ( .IN1(n2426), .IN2(n8710), .IN3(n2440), .QN(n4267) );
  NAND3X0 U8485 ( .IN1(n8711), .IN2(n8712), .IN3(n8681), .QN(n8710) );
  NAND2X0 U8486 ( .IN1(n8713), .IN2(n8683), .QN(n8712) );
  INVX0 U8487 ( .INP(n8714), .ZN(n8713) );
  NAND2X0 U8488 ( .IN1(n8685), .IN2(DFF_446_n1), .QN(n8711) );
  NAND2X0 U8489 ( .IN1(n8699), .IN2(n8715), .QN(n4266) );
  NAND3X0 U8490 ( .IN1(n8716), .IN2(n8717), .IN3(n8681), .QN(n8715) );
  NAND2X0 U8491 ( .IN1(n8718), .IN2(n8683), .QN(n8717) );
  NAND2X0 U8492 ( .IN1(n8685), .IN2(DFF_447_n1), .QN(n8716) );
  INVX0 U8493 ( .INP(n8719), .ZN(n8699) );
  NAND2X0 U8494 ( .IN1(n2426), .IN2(n8720), .QN(n8719) );
  NAND2X0 U8495 ( .IN1(n2446), .IN2(n2445), .QN(n8720) );
  NAND2X0 U8496 ( .IN1(n2426), .IN2(n8721), .QN(n4265) );
  NAND3X0 U8497 ( .IN1(n8722), .IN2(n8723), .IN3(n8681), .QN(n8721) );
  NAND2X0 U8498 ( .IN1(n8724), .IN2(n8683), .QN(n8723) );
  INVX0 U8499 ( .INP(n8725), .ZN(n8724) );
  NAND2X0 U8500 ( .IN1(n8685), .IN2(DFF_448_n1), .QN(n8722) );
  NAND2X0 U8501 ( .IN1(DFF_1562_n1), .IN2(n8726), .QN(n4263) );
  NAND2X0 U8502 ( .IN1(n8727), .IN2(n8728), .QN(n4262) );
  XOR2X1 U8503 ( .IN1(n4481), .IN2(n8729), .Q(n8727) );
  XNOR2X1 U8504 ( .IN1(n8730), .IN2(n8731), .Q(n4261) );
  XOR2X1 U8505 ( .IN1(n8731), .IN2(n8732), .Q(n4260) );
  INVX0 U8506 ( .INP(n8733), .ZN(n8732) );
  NOR2X0 U8507 ( .IN1(g3231), .IN2(n14353), .QN(n8731) );
  NAND3X0 U8508 ( .IN1(n8734), .IN2(n8735), .IN3(n8736), .QN(n4259) );
  NAND2X0 U8509 ( .IN1(test_so22), .IN2(n8737), .QN(n8736) );
  XOR2X1 U8510 ( .IN1(n8738), .IN2(n8739), .Q(n8737) );
  XNOR3X1 U8511 ( .IN1(n8725), .IN2(n8718), .IN3(n8740), .Q(n8739) );
  XNOR2X1 U8512 ( .IN1(n8709), .IN2(n8714), .Q(n8740) );
  NAND3X0 U8513 ( .IN1(n8741), .IN2(n8742), .IN3(n8743), .QN(n8714) );
  NAND2X0 U8514 ( .IN1(n8744), .IN2(n8745), .QN(n8742) );
  NAND2X0 U8515 ( .IN1(n8746), .IN2(n8747), .QN(n8741) );
  NAND3X0 U8516 ( .IN1(n8748), .IN2(n8749), .IN3(n8743), .QN(n8709) );
  NAND2X0 U8517 ( .IN1(n8750), .IN2(n8751), .QN(n8749) );
  NAND2X0 U8518 ( .IN1(n8752), .IN2(n8753), .QN(n8748) );
  INVX0 U8519 ( .INP(n8754), .ZN(n8718) );
  NAND3X0 U8520 ( .IN1(n8755), .IN2(n8756), .IN3(n8743), .QN(n8754) );
  NAND2X0 U8521 ( .IN1(n8757), .IN2(n8751), .QN(n8756) );
  NAND2X0 U8522 ( .IN1(n8752), .IN2(n8758), .QN(n8755) );
  NAND3X0 U8523 ( .IN1(n8759), .IN2(n8760), .IN3(n8761), .QN(n8725) );
  NAND2X0 U8524 ( .IN1(n8762), .IN2(n8745), .QN(n8760) );
  NAND2X0 U8525 ( .IN1(n8746), .IN2(n8763), .QN(n8759) );
  XNOR3X1 U8526 ( .IN1(n8704), .IN2(n8698), .IN3(n8764), .Q(n8738) );
  XNOR2X1 U8527 ( .IN1(n8684), .IN2(n8692), .Q(n8764) );
  NAND3X0 U8528 ( .IN1(n8765), .IN2(n8766), .IN3(n8761), .QN(n8692) );
  NAND2X0 U8529 ( .IN1(n8767), .IN2(n8745), .QN(n8766) );
  NAND2X0 U8530 ( .IN1(n8746), .IN2(n8768), .QN(n8765) );
  NAND3X0 U8531 ( .IN1(n8769), .IN2(n8770), .IN3(n8771), .QN(n8684) );
  NAND2X0 U8532 ( .IN1(n8772), .IN2(n8751), .QN(n8770) );
  NAND2X0 U8533 ( .IN1(n8752), .IN2(n8773), .QN(n8769) );
  INVX0 U8534 ( .INP(n8774), .ZN(n8698) );
  NAND3X0 U8535 ( .IN1(n8775), .IN2(n8776), .IN3(n8743), .QN(n8774) );
  NAND2X0 U8536 ( .IN1(n8777), .IN2(n8751), .QN(n8776) );
  NAND2X0 U8537 ( .IN1(n8752), .IN2(n8778), .QN(n8775) );
  NAND3X0 U8538 ( .IN1(n8779), .IN2(n8780), .IN3(n8743), .QN(n8704) );
  NAND2X0 U8539 ( .IN1(n8781), .IN2(n8745), .QN(n8780) );
  NAND2X0 U8540 ( .IN1(n8746), .IN2(n8782), .QN(n8779) );
  NAND4X0 U8541 ( .IN1(n8681), .IN2(n8685), .IN3(n8783), .IN4(n8784), .QN(
        n8735) );
  NAND2X0 U8542 ( .IN1(n14345), .IN2(n8785), .QN(n8784) );
  NAND2X0 U8543 ( .IN1(n4492), .IN2(g3229), .QN(n8783) );
  NOR2X0 U8544 ( .IN1(n8683), .IN2(n8548), .QN(n8685) );
  NAND2X0 U8545 ( .IN1(n8786), .IN2(g557), .QN(n8734) );
  XOR2X1 U8546 ( .IN1(n8688), .IN2(n8695), .Q(n8786) );
  NAND3X0 U8547 ( .IN1(n8787), .IN2(n8788), .IN3(n8771), .QN(n8695) );
  INVX0 U8548 ( .INP(n8789), .ZN(n8771) );
  NAND2X0 U8549 ( .IN1(n8743), .IN2(n8790), .QN(n8789) );
  NAND2X0 U8550 ( .IN1(n8791), .IN2(n8751), .QN(n8790) );
  NAND2X0 U8551 ( .IN1(n8792), .IN2(n8751), .QN(n8788) );
  NAND2X0 U8552 ( .IN1(n8752), .IN2(n8793), .QN(n8787) );
  NOR2X0 U8553 ( .IN1(n8751), .IN2(n8791), .QN(n8752) );
  NAND3X0 U8554 ( .IN1(n8794), .IN2(n8795), .IN3(n8761), .QN(n8688) );
  INVX0 U8555 ( .INP(n8796), .ZN(n8761) );
  NAND2X0 U8556 ( .IN1(n8743), .IN2(n8797), .QN(n8796) );
  NAND2X0 U8557 ( .IN1(n8791), .IN2(n8745), .QN(n8797) );
  NOR2X0 U8558 ( .IN1(n8548), .IN2(n4541), .QN(n8743) );
  NAND3X0 U8559 ( .IN1(n8798), .IN2(n7744), .IN3(n8799), .QN(n8548) );
  NOR2X0 U8560 ( .IN1(g563), .IN2(n8800), .QN(n8799) );
  NOR2X0 U8561 ( .IN1(n4298), .IN2(g499), .QN(n8800) );
  INVX0 U8562 ( .INP(g21851), .ZN(n8798) );
  NAND2X0 U8563 ( .IN1(n8801), .IN2(n8745), .QN(n8795) );
  NAND2X0 U8564 ( .IN1(n8746), .IN2(n8802), .QN(n8794) );
  NOR2X0 U8565 ( .IN1(n8745), .IN2(n8791), .QN(n8746) );
  INVX0 U8566 ( .INP(n8803), .ZN(n8791) );
  NAND2X0 U8567 ( .IN1(n8804), .IN2(n8805), .QN(n4258) );
  NAND2X0 U8568 ( .IN1(n2361), .IN2(n8806), .QN(n8805) );
  NAND3X0 U8569 ( .IN1(n8807), .IN2(n8808), .IN3(n8809), .QN(n8804) );
  NAND2X0 U8570 ( .IN1(n8810), .IN2(n8811), .QN(n8808) );
  NAND2X0 U8571 ( .IN1(n7144), .IN2(n8812), .QN(n8807) );
  NAND3X0 U8572 ( .IN1(n8813), .IN2(n8814), .IN3(n2375), .QN(n4257) );
  NAND3X0 U8573 ( .IN1(n8815), .IN2(n8816), .IN3(n8809), .QN(n8813) );
  NAND2X0 U8574 ( .IN1(n8817), .IN2(n8811), .QN(n8816) );
  INVX0 U8575 ( .INP(n8818), .ZN(n8817) );
  NAND2X0 U8576 ( .IN1(n8812), .IN2(DFF_1495_n1), .QN(n8815) );
  NAND2X0 U8577 ( .IN1(n8814), .IN2(n8819), .QN(n4256) );
  NAND3X0 U8578 ( .IN1(n8820), .IN2(n8821), .IN3(n8809), .QN(n8819) );
  NAND2X0 U8579 ( .IN1(n8822), .IN2(n8811), .QN(n8821) );
  NAND2X0 U8580 ( .IN1(n8812), .IN2(DFF_1499_n1), .QN(n8820) );
  NAND3X0 U8581 ( .IN1(n8823), .IN2(n8814), .IN3(n2375), .QN(n4255) );
  NAND3X0 U8582 ( .IN1(n8824), .IN2(n8825), .IN3(n8809), .QN(n8823) );
  NAND2X0 U8583 ( .IN1(n8826), .IN2(n8811), .QN(n8825) );
  NAND2X0 U8584 ( .IN1(n8812), .IN2(DFF_1496_n1), .QN(n8824) );
  NAND2X0 U8585 ( .IN1(n8827), .IN2(n8828), .QN(n4254) );
  NAND3X0 U8586 ( .IN1(n8829), .IN2(n8830), .IN3(n8809), .QN(n8828) );
  NAND2X0 U8587 ( .IN1(n8831), .IN2(n8811), .QN(n8830) );
  NAND2X0 U8588 ( .IN1(n8812), .IN2(DFF_1494_n1), .QN(n8829) );
  NAND2X0 U8589 ( .IN1(n8832), .IN2(n8833), .QN(n4253) );
  NAND2X0 U8590 ( .IN1(n2361), .IN2(n8834), .QN(n8833) );
  NAND3X0 U8591 ( .IN1(n8835), .IN2(n8836), .IN3(n8809), .QN(n8832) );
  NAND2X0 U8592 ( .IN1(n8837), .IN2(n8811), .QN(n8836) );
  INVX0 U8593 ( .INP(n8838), .ZN(n8837) );
  NAND2X0 U8594 ( .IN1(n8812), .IN2(n7145), .QN(n8835) );
  NAND2X0 U8595 ( .IN1(n8827), .IN2(n8839), .QN(n4252) );
  NAND3X0 U8596 ( .IN1(n8840), .IN2(n8841), .IN3(n8809), .QN(n8839) );
  NAND2X0 U8597 ( .IN1(n8842), .IN2(n8811), .QN(n8841) );
  INVX0 U8598 ( .INP(n8843), .ZN(n8842) );
  NAND2X0 U8599 ( .IN1(n8812), .IN2(DFF_1497_n1), .QN(n8840) );
  INVX0 U8600 ( .INP(n8844), .ZN(n8827) );
  NAND2X0 U8601 ( .IN1(n8814), .IN2(n8845), .QN(n8844) );
  NAND2X0 U8602 ( .IN1(n2361), .IN2(n2374), .QN(n8845) );
  NAND2X0 U8603 ( .IN1(n8814), .IN2(n8846), .QN(n4251) );
  NAND3X0 U8604 ( .IN1(n8847), .IN2(n8848), .IN3(n8809), .QN(n8846) );
  NAND2X0 U8605 ( .IN1(n8849), .IN2(n8811), .QN(n8848) );
  INVX0 U8606 ( .INP(n8850), .ZN(n8849) );
  NAND2X0 U8607 ( .IN1(n8812), .IN2(DFF_1498_n1), .QN(n8847) );
  NAND2X0 U8608 ( .IN1(n2361), .IN2(n8851), .QN(n8814) );
  NAND3X0 U8609 ( .IN1(n8852), .IN2(n8853), .IN3(n8854), .QN(n4250) );
  NAND2X0 U8610 ( .IN1(n8855), .IN2(g2584), .QN(n8854) );
  XOR3X1 U8611 ( .IN1(n8856), .IN2(n8857), .IN3(n8858), .Q(n8855) );
  XOR3X1 U8612 ( .IN1(n8850), .IN2(n8843), .IN3(n8859), .Q(n8858) );
  XOR2X1 U8613 ( .IN1(n8838), .IN2(n8831), .Q(n8859) );
  INVX0 U8614 ( .INP(n8860), .ZN(n8831) );
  NAND3X0 U8615 ( .IN1(n8861), .IN2(n8862), .IN3(n8863), .QN(n8860) );
  NAND2X0 U8616 ( .IN1(n8864), .IN2(n8865), .QN(n8862) );
  NAND2X0 U8617 ( .IN1(n8866), .IN2(n8867), .QN(n8861) );
  NAND3X0 U8618 ( .IN1(n8868), .IN2(n8869), .IN3(n8870), .QN(n8838) );
  NAND2X0 U8619 ( .IN1(n8871), .IN2(n8865), .QN(n8869) );
  NAND2X0 U8620 ( .IN1(n8866), .IN2(n8872), .QN(n8868) );
  NAND3X0 U8621 ( .IN1(n8873), .IN2(n8874), .IN3(n8863), .QN(n8843) );
  NAND2X0 U8622 ( .IN1(n8875), .IN2(n8876), .QN(n8874) );
  NAND2X0 U8623 ( .IN1(n8877), .IN2(n8878), .QN(n8873) );
  NAND3X0 U8624 ( .IN1(n8879), .IN2(n8880), .IN3(n8870), .QN(n8850) );
  NAND2X0 U8625 ( .IN1(n8881), .IN2(n8865), .QN(n8880) );
  NAND2X0 U8626 ( .IN1(n8866), .IN2(n8882), .QN(n8879) );
  XOR2X1 U8627 ( .IN1(n8818), .IN2(n8810), .Q(n8857) );
  INVX0 U8628 ( .INP(n8883), .ZN(n8810) );
  NAND3X0 U8629 ( .IN1(n8884), .IN2(n8885), .IN3(n8863), .QN(n8883) );
  NAND2X0 U8630 ( .IN1(n8886), .IN2(n8876), .QN(n8885) );
  NAND2X0 U8631 ( .IN1(n8877), .IN2(n8887), .QN(n8884) );
  NAND3X0 U8632 ( .IN1(n8888), .IN2(n8889), .IN3(n8863), .QN(n8818) );
  NAND2X0 U8633 ( .IN1(n8890), .IN2(n8876), .QN(n8889) );
  NAND2X0 U8634 ( .IN1(n8877), .IN2(n8891), .QN(n8888) );
  XOR2X1 U8635 ( .IN1(n8822), .IN2(n8826), .Q(n8856) );
  INVX0 U8636 ( .INP(n8892), .ZN(n8826) );
  NAND3X0 U8637 ( .IN1(n8893), .IN2(n8894), .IN3(n8863), .QN(n8892) );
  NAND2X0 U8638 ( .IN1(n8895), .IN2(n8865), .QN(n8894) );
  NAND2X0 U8639 ( .IN1(n8866), .IN2(n8896), .QN(n8893) );
  NOR3X0 U8640 ( .IN1(n8897), .IN2(n8898), .IN3(n8899), .QN(n8822) );
  NOR2X0 U8641 ( .IN1(n8900), .IN2(n8901), .QN(n8898) );
  INVX0 U8642 ( .INP(n8902), .ZN(n8897) );
  NAND2X0 U8643 ( .IN1(n8877), .IN2(n8900), .QN(n8902) );
  NAND4X0 U8644 ( .IN1(n8809), .IN2(n8812), .IN3(n8903), .IN4(n8904), .QN(
        n8853) );
  NAND2X0 U8645 ( .IN1(n14346), .IN2(n8785), .QN(n8904) );
  NAND2X0 U8646 ( .IN1(n4490), .IN2(g3229), .QN(n8903) );
  NOR2X0 U8647 ( .IN1(n8851), .IN2(n8811), .QN(n8812) );
  NAND2X0 U8648 ( .IN1(n8905), .IN2(g2631), .QN(n8852) );
  XOR2X1 U8649 ( .IN1(n8806), .IN2(n8834), .Q(n8905) );
  NAND3X0 U8650 ( .IN1(n8906), .IN2(n8907), .IN3(n8870), .QN(n8834) );
  INVX0 U8651 ( .INP(n8908), .ZN(n8870) );
  NAND2X0 U8652 ( .IN1(n8863), .IN2(n8909), .QN(n8908) );
  NAND2X0 U8653 ( .IN1(n8910), .IN2(n8865), .QN(n8909) );
  NAND2X0 U8654 ( .IN1(n8911), .IN2(n8865), .QN(n8907) );
  NAND2X0 U8655 ( .IN1(n8866), .IN2(n8912), .QN(n8906) );
  NOR2X0 U8656 ( .IN1(n8865), .IN2(n8910), .QN(n8866) );
  NAND3X0 U8657 ( .IN1(n8913), .IN2(n8914), .IN3(n8915), .QN(n8806) );
  INVX0 U8658 ( .INP(n8899), .ZN(n8915) );
  NAND2X0 U8659 ( .IN1(n8863), .IN2(n8916), .QN(n8899) );
  NAND2X0 U8660 ( .IN1(n8910), .IN2(n8876), .QN(n8916) );
  NOR2X0 U8661 ( .IN1(n8851), .IN2(n4543), .QN(n8863) );
  NAND2X0 U8662 ( .IN1(n8917), .IN2(n7749), .QN(n8851) );
  NOR2X0 U8663 ( .IN1(g2637), .IN2(g30072), .QN(n8917) );
  NAND2X0 U8664 ( .IN1(n8918), .IN2(n8876), .QN(n8914) );
  NAND2X0 U8665 ( .IN1(n8877), .IN2(n8919), .QN(n8913) );
  NOR2X0 U8666 ( .IN1(n8876), .IN2(n8910), .QN(n8877) );
  INVX0 U8667 ( .INP(n8920), .ZN(n8910) );
  NAND2X0 U8668 ( .IN1(n8921), .IN2(n8922), .QN(n4249) );
  NAND2X0 U8669 ( .IN1(n2289), .IN2(n8923), .QN(n8922) );
  NAND3X0 U8670 ( .IN1(n8924), .IN2(n8925), .IN3(n8926), .QN(n8921) );
  NAND2X0 U8671 ( .IN1(n8927), .IN2(n8928), .QN(n8925) );
  NAND2X0 U8672 ( .IN1(n7146), .IN2(n8929), .QN(n8924) );
  NAND3X0 U8673 ( .IN1(n2275), .IN2(n8930), .IN3(n2303), .QN(n4248) );
  NAND3X0 U8674 ( .IN1(n8931), .IN2(n8932), .IN3(n8926), .QN(n8930) );
  NAND2X0 U8675 ( .IN1(n8933), .IN2(n8928), .QN(n8932) );
  INVX0 U8676 ( .INP(n8934), .ZN(n8933) );
  NAND2X0 U8677 ( .IN1(n8929), .IN2(DFF_1145_n1), .QN(n8931) );
  NAND2X0 U8678 ( .IN1(n2275), .IN2(n8935), .QN(n4247) );
  NAND3X0 U8679 ( .IN1(n8936), .IN2(n8937), .IN3(n8926), .QN(n8935) );
  NAND2X0 U8680 ( .IN1(n8938), .IN2(n8928), .QN(n8937) );
  NAND2X0 U8681 ( .IN1(n8929), .IN2(DFF_1149_n1), .QN(n8936) );
  NAND3X0 U8682 ( .IN1(n2275), .IN2(n8939), .IN3(n2303), .QN(n4246) );
  NAND3X0 U8683 ( .IN1(n8940), .IN2(n8941), .IN3(n8926), .QN(n8939) );
  NAND2X0 U8684 ( .IN1(n8942), .IN2(n8928), .QN(n8941) );
  NAND2X0 U8685 ( .IN1(n8929), .IN2(DFF_1146_n1), .QN(n8940) );
  NAND2X0 U8686 ( .IN1(n8943), .IN2(n8944), .QN(n4245) );
  NAND3X0 U8687 ( .IN1(n8945), .IN2(n8946), .IN3(n8926), .QN(n8944) );
  NAND2X0 U8688 ( .IN1(n8947), .IN2(n8928), .QN(n8946) );
  NAND2X0 U8689 ( .IN1(n8929), .IN2(DFF_1144_n1), .QN(n8945) );
  NAND2X0 U8690 ( .IN1(n8948), .IN2(n8949), .QN(n4244) );
  NAND2X0 U8691 ( .IN1(n2289), .IN2(n8950), .QN(n8949) );
  NAND3X0 U8692 ( .IN1(n8951), .IN2(n8952), .IN3(n8926), .QN(n8948) );
  NAND2X0 U8693 ( .IN1(n8953), .IN2(n8928), .QN(n8952) );
  INVX0 U8694 ( .INP(n8954), .ZN(n8953) );
  NAND2X0 U8695 ( .IN1(n7147), .IN2(n8929), .QN(n8951) );
  NAND2X0 U8696 ( .IN1(n8943), .IN2(n8955), .QN(n4243) );
  NAND3X0 U8697 ( .IN1(n8956), .IN2(n8957), .IN3(n8926), .QN(n8955) );
  NAND2X0 U8698 ( .IN1(n8958), .IN2(n8928), .QN(n8957) );
  INVX0 U8699 ( .INP(n8959), .ZN(n8958) );
  NAND2X0 U8700 ( .IN1(n8929), .IN2(DFF_1147_n1), .QN(n8956) );
  INVX0 U8701 ( .INP(n8960), .ZN(n8943) );
  NAND2X0 U8702 ( .IN1(n2275), .IN2(n8961), .QN(n8960) );
  NAND2X0 U8703 ( .IN1(n2289), .IN2(n2302), .QN(n8961) );
  NAND2X0 U8704 ( .IN1(n2275), .IN2(n8962), .QN(n4242) );
  NAND3X0 U8705 ( .IN1(n8963), .IN2(n8964), .IN3(n8926), .QN(n8962) );
  NAND2X0 U8706 ( .IN1(n8965), .IN2(n8928), .QN(n8964) );
  INVX0 U8707 ( .INP(n8966), .ZN(n8965) );
  NAND2X0 U8708 ( .IN1(n8929), .IN2(DFF_1148_n1), .QN(n8963) );
  NAND3X0 U8709 ( .IN1(n8967), .IN2(n8968), .IN3(n8969), .QN(n4241) );
  NAND2X0 U8710 ( .IN1(n8970), .IN2(g1890), .QN(n8969) );
  XOR3X1 U8711 ( .IN1(n8971), .IN2(n8972), .IN3(n8973), .Q(n8970) );
  XOR3X1 U8712 ( .IN1(n8966), .IN2(n8959), .IN3(n8974), .Q(n8973) );
  XOR2X1 U8713 ( .IN1(n8954), .IN2(n8947), .Q(n8974) );
  INVX0 U8714 ( .INP(n8975), .ZN(n8947) );
  NAND3X0 U8715 ( .IN1(n8976), .IN2(n8977), .IN3(n8978), .QN(n8975) );
  NAND2X0 U8716 ( .IN1(n8979), .IN2(n8980), .QN(n8977) );
  NAND2X0 U8717 ( .IN1(n8981), .IN2(n8982), .QN(n8976) );
  NAND3X0 U8718 ( .IN1(n8983), .IN2(n8984), .IN3(n8985), .QN(n8954) );
  NAND2X0 U8719 ( .IN1(n8986), .IN2(n8980), .QN(n8984) );
  NAND2X0 U8720 ( .IN1(n8981), .IN2(n8987), .QN(n8983) );
  NAND3X0 U8721 ( .IN1(n8988), .IN2(n8989), .IN3(n8978), .QN(n8959) );
  INVX0 U8722 ( .INP(n8990), .ZN(n8989) );
  NOR2X0 U8723 ( .IN1(n8991), .IN2(n8992), .QN(n8990) );
  NAND2X0 U8724 ( .IN1(n8993), .IN2(n8991), .QN(n8988) );
  NAND3X0 U8725 ( .IN1(n8994), .IN2(n8995), .IN3(n8985), .QN(n8966) );
  NAND2X0 U8726 ( .IN1(n8996), .IN2(n8980), .QN(n8995) );
  NAND2X0 U8727 ( .IN1(n8981), .IN2(n8997), .QN(n8994) );
  XOR2X1 U8728 ( .IN1(n8934), .IN2(n8927), .Q(n8972) );
  INVX0 U8729 ( .INP(n8998), .ZN(n8927) );
  NAND3X0 U8730 ( .IN1(n8999), .IN2(n9000), .IN3(n8978), .QN(n8998) );
  NAND2X0 U8731 ( .IN1(n9001), .IN2(n9002), .QN(n9000) );
  NAND2X0 U8732 ( .IN1(n8993), .IN2(n9003), .QN(n8999) );
  NAND3X0 U8733 ( .IN1(n9004), .IN2(n9005), .IN3(n8978), .QN(n8934) );
  NAND2X0 U8734 ( .IN1(n9006), .IN2(n9002), .QN(n9005) );
  NAND2X0 U8735 ( .IN1(n8993), .IN2(n9007), .QN(n9004) );
  XOR2X1 U8736 ( .IN1(n8938), .IN2(n8942), .Q(n8971) );
  INVX0 U8737 ( .INP(n9008), .ZN(n8942) );
  NAND3X0 U8738 ( .IN1(n9009), .IN2(n9010), .IN3(n8978), .QN(n9008) );
  NAND2X0 U8739 ( .IN1(n9011), .IN2(n8980), .QN(n9010) );
  NAND2X0 U8740 ( .IN1(n8981), .IN2(n9012), .QN(n9009) );
  NOR3X0 U8741 ( .IN1(n9013), .IN2(n9014), .IN3(n9015), .QN(n8938) );
  NOR2X0 U8742 ( .IN1(n9016), .IN2(n8992), .QN(n9014) );
  INVX0 U8743 ( .INP(n9017), .ZN(n9013) );
  NAND2X0 U8744 ( .IN1(n8993), .IN2(n9016), .QN(n9017) );
  NAND4X0 U8745 ( .IN1(n8926), .IN2(n8929), .IN3(n9018), .IN4(n9019), .QN(
        n8968) );
  NAND2X0 U8746 ( .IN1(g3229), .IN2(n8094), .QN(n9019) );
  NAND2X0 U8747 ( .IN1(n14347), .IN2(n8785), .QN(n9018) );
  NOR2X0 U8748 ( .IN1(n8547), .IN2(n8928), .QN(n8929) );
  NAND2X0 U8749 ( .IN1(n9020), .IN2(g1937), .QN(n8967) );
  XOR2X1 U8750 ( .IN1(n8923), .IN2(n8950), .Q(n9020) );
  NAND3X0 U8751 ( .IN1(n9021), .IN2(n9022), .IN3(n8985), .QN(n8950) );
  INVX0 U8752 ( .INP(n9023), .ZN(n8985) );
  NAND2X0 U8753 ( .IN1(n8978), .IN2(n9024), .QN(n9023) );
  NAND2X0 U8754 ( .IN1(n9025), .IN2(n8980), .QN(n9024) );
  NAND2X0 U8755 ( .IN1(n9026), .IN2(n8980), .QN(n9022) );
  NAND2X0 U8756 ( .IN1(n8981), .IN2(n9027), .QN(n9021) );
  NOR2X0 U8757 ( .IN1(n8980), .IN2(n9025), .QN(n8981) );
  NAND3X0 U8758 ( .IN1(n9028), .IN2(n9029), .IN3(n9030), .QN(n8923) );
  INVX0 U8759 ( .INP(n9015), .ZN(n9030) );
  NAND2X0 U8760 ( .IN1(n8978), .IN2(n9031), .QN(n9015) );
  NAND2X0 U8761 ( .IN1(n9025), .IN2(n9002), .QN(n9031) );
  NOR2X0 U8762 ( .IN1(n8547), .IN2(n4545), .QN(n8978) );
  NAND2X0 U8763 ( .IN1(n9032), .IN2(n7750), .QN(n8547) );
  NOR2X0 U8764 ( .IN1(g1943), .IN2(n497), .QN(n9032) );
  NAND2X0 U8765 ( .IN1(n9033), .IN2(n9002), .QN(n9029) );
  NAND2X0 U8766 ( .IN1(n8993), .IN2(n9034), .QN(n9028) );
  NOR2X0 U8767 ( .IN1(n9002), .IN2(n9025), .QN(n8993) );
  INVX0 U8768 ( .INP(n9035), .ZN(n9025) );
  NAND2X0 U8769 ( .IN1(n9036), .IN2(n9037), .QN(n4240) );
  NAND2X0 U8770 ( .IN1(n2217), .IN2(n9038), .QN(n9037) );
  NAND3X0 U8771 ( .IN1(n9039), .IN2(n9040), .IN3(n9041), .QN(n9036) );
  NAND2X0 U8772 ( .IN1(n9042), .IN2(n9043), .QN(n9040) );
  NAND2X0 U8773 ( .IN1(n7148), .IN2(n9044), .QN(n9039) );
  NAND3X0 U8774 ( .IN1(n9045), .IN2(n9046), .IN3(n2231), .QN(n4239) );
  NAND3X0 U8775 ( .IN1(n9047), .IN2(n9048), .IN3(n9041), .QN(n9045) );
  NAND2X0 U8776 ( .IN1(n9049), .IN2(n9043), .QN(n9048) );
  INVX0 U8777 ( .INP(n9050), .ZN(n9049) );
  NAND2X0 U8778 ( .IN1(n9044), .IN2(DFF_795_n1), .QN(n9047) );
  NAND2X0 U8779 ( .IN1(n9046), .IN2(n9051), .QN(n4238) );
  NAND3X0 U8780 ( .IN1(n9052), .IN2(n9053), .IN3(n9041), .QN(n9051) );
  NAND2X0 U8781 ( .IN1(n9054), .IN2(n9043), .QN(n9053) );
  NAND2X0 U8782 ( .IN1(n9044), .IN2(DFF_799_n1), .QN(n9052) );
  NAND3X0 U8783 ( .IN1(n9055), .IN2(n9046), .IN3(n2231), .QN(n4237) );
  NAND3X0 U8784 ( .IN1(n9056), .IN2(n9057), .IN3(n9041), .QN(n9055) );
  NAND2X0 U8785 ( .IN1(n9058), .IN2(n9043), .QN(n9057) );
  NAND2X0 U8786 ( .IN1(n9044), .IN2(DFF_796_n1), .QN(n9056) );
  NAND2X0 U8787 ( .IN1(n9059), .IN2(n9060), .QN(n4236) );
  NAND3X0 U8788 ( .IN1(n9061), .IN2(n9062), .IN3(n9041), .QN(n9060) );
  NAND2X0 U8789 ( .IN1(n9063), .IN2(n9043), .QN(n9062) );
  NAND2X0 U8790 ( .IN1(n9044), .IN2(DFF_794_n1), .QN(n9061) );
  NAND2X0 U8791 ( .IN1(n9064), .IN2(n9065), .QN(n4235) );
  NAND2X0 U8792 ( .IN1(n2217), .IN2(n9066), .QN(n9065) );
  NAND3X0 U8793 ( .IN1(n9067), .IN2(n9068), .IN3(n9041), .QN(n9064) );
  NAND2X0 U8794 ( .IN1(n9069), .IN2(n9043), .QN(n9068) );
  INVX0 U8795 ( .INP(n9070), .ZN(n9069) );
  NAND2X0 U8796 ( .IN1(n7149), .IN2(n9044), .QN(n9067) );
  NAND2X0 U8797 ( .IN1(n9059), .IN2(n9071), .QN(n4234) );
  NAND3X0 U8798 ( .IN1(n9072), .IN2(n9073), .IN3(n9041), .QN(n9071) );
  NAND2X0 U8799 ( .IN1(n9074), .IN2(n9043), .QN(n9073) );
  INVX0 U8800 ( .INP(n9075), .ZN(n9074) );
  NAND2X0 U8801 ( .IN1(n9044), .IN2(DFF_797_n1), .QN(n9072) );
  INVX0 U8802 ( .INP(n9076), .ZN(n9059) );
  NAND2X0 U8803 ( .IN1(n9046), .IN2(n9077), .QN(n9076) );
  NAND2X0 U8804 ( .IN1(n2217), .IN2(n2230), .QN(n9077) );
  NAND2X0 U8805 ( .IN1(n9046), .IN2(n9078), .QN(n4233) );
  NAND3X0 U8806 ( .IN1(n9079), .IN2(n9080), .IN3(n9041), .QN(n9078) );
  NAND2X0 U8807 ( .IN1(n9081), .IN2(n9043), .QN(n9080) );
  INVX0 U8808 ( .INP(n9082), .ZN(n9081) );
  NAND2X0 U8809 ( .IN1(n9044), .IN2(DFF_798_n1), .QN(n9079) );
  NAND2X0 U8810 ( .IN1(n2217), .IN2(n9083), .QN(n9046) );
  NAND3X0 U8811 ( .IN1(n9084), .IN2(n9085), .IN3(n9086), .QN(n4232) );
  NAND2X0 U8812 ( .IN1(n9087), .IN2(g1196), .QN(n9086) );
  XOR3X1 U8813 ( .IN1(n9088), .IN2(n9089), .IN3(n9090), .Q(n9087) );
  XOR3X1 U8814 ( .IN1(n9082), .IN2(n9075), .IN3(n9091), .Q(n9090) );
  XOR2X1 U8815 ( .IN1(n9070), .IN2(n9063), .Q(n9091) );
  INVX0 U8816 ( .INP(n9092), .ZN(n9063) );
  NAND3X0 U8817 ( .IN1(n9093), .IN2(n9094), .IN3(n9095), .QN(n9092) );
  NAND2X0 U8818 ( .IN1(n9096), .IN2(n9097), .QN(n9094) );
  NAND2X0 U8819 ( .IN1(n9098), .IN2(n9099), .QN(n9093) );
  NAND3X0 U8820 ( .IN1(n9100), .IN2(n9101), .IN3(n9102), .QN(n9070) );
  NAND2X0 U8821 ( .IN1(n9103), .IN2(n9097), .QN(n9101) );
  NAND2X0 U8822 ( .IN1(n9098), .IN2(n9104), .QN(n9100) );
  NAND3X0 U8823 ( .IN1(n9105), .IN2(n9106), .IN3(n9095), .QN(n9075) );
  NAND2X0 U8824 ( .IN1(n9107), .IN2(n9108), .QN(n9106) );
  NAND2X0 U8825 ( .IN1(n9109), .IN2(n9110), .QN(n9105) );
  NAND3X0 U8826 ( .IN1(n9111), .IN2(n9112), .IN3(n9102), .QN(n9082) );
  NAND2X0 U8827 ( .IN1(n9113), .IN2(n9097), .QN(n9112) );
  NAND2X0 U8828 ( .IN1(n9098), .IN2(n9114), .QN(n9111) );
  XOR2X1 U8829 ( .IN1(n9050), .IN2(n9042), .Q(n9089) );
  INVX0 U8830 ( .INP(n9115), .ZN(n9042) );
  NAND3X0 U8831 ( .IN1(n9116), .IN2(n9117), .IN3(n9095), .QN(n9115) );
  INVX0 U8832 ( .INP(n9118), .ZN(n9117) );
  NOR2X0 U8833 ( .IN1(n9119), .IN2(n9120), .QN(n9118) );
  NAND2X0 U8834 ( .IN1(n9109), .IN2(n9119), .QN(n9116) );
  NAND3X0 U8835 ( .IN1(n9121), .IN2(n9122), .IN3(n9095), .QN(n9050) );
  NAND2X0 U8836 ( .IN1(n9123), .IN2(n9108), .QN(n9122) );
  NAND2X0 U8837 ( .IN1(n9109), .IN2(n9124), .QN(n9121) );
  XOR2X1 U8838 ( .IN1(n9054), .IN2(n9058), .Q(n9088) );
  INVX0 U8839 ( .INP(n9125), .ZN(n9058) );
  NAND3X0 U8840 ( .IN1(n9126), .IN2(n9127), .IN3(n9095), .QN(n9125) );
  NAND2X0 U8841 ( .IN1(n9128), .IN2(n9097), .QN(n9127) );
  NAND2X0 U8842 ( .IN1(n9098), .IN2(n9129), .QN(n9126) );
  NOR3X0 U8843 ( .IN1(n9130), .IN2(n9131), .IN3(n9132), .QN(n9054) );
  NOR2X0 U8844 ( .IN1(n9133), .IN2(n9120), .QN(n9131) );
  INVX0 U8845 ( .INP(n9134), .ZN(n9130) );
  NAND2X0 U8846 ( .IN1(n9109), .IN2(n9133), .QN(n9134) );
  NAND4X0 U8847 ( .IN1(n9041), .IN2(n9044), .IN3(n9135), .IN4(n9136), .QN(
        n9085) );
  NAND2X0 U8848 ( .IN1(n4489), .IN2(g3229), .QN(n9136) );
  NAND2X0 U8849 ( .IN1(n8785), .IN2(n14348), .QN(n9135) );
  NOR2X0 U8850 ( .IN1(n9083), .IN2(n9043), .QN(n9044) );
  NAND2X0 U8851 ( .IN1(n9137), .IN2(g1243), .QN(n9084) );
  XOR2X1 U8852 ( .IN1(n9038), .IN2(n9066), .Q(n9137) );
  NAND3X0 U8853 ( .IN1(n9138), .IN2(n9139), .IN3(n9102), .QN(n9066) );
  INVX0 U8854 ( .INP(n9140), .ZN(n9102) );
  NAND2X0 U8855 ( .IN1(n9095), .IN2(n9141), .QN(n9140) );
  NAND2X0 U8856 ( .IN1(n9142), .IN2(n9097), .QN(n9141) );
  NAND2X0 U8857 ( .IN1(n9143), .IN2(n9097), .QN(n9139) );
  NAND2X0 U8858 ( .IN1(n9098), .IN2(n9144), .QN(n9138) );
  NOR2X0 U8859 ( .IN1(n9097), .IN2(n9142), .QN(n9098) );
  NAND3X0 U8860 ( .IN1(n9145), .IN2(n9146), .IN3(n9147), .QN(n9038) );
  INVX0 U8861 ( .INP(n9132), .ZN(n9147) );
  NAND2X0 U8862 ( .IN1(n9095), .IN2(n9148), .QN(n9132) );
  NAND2X0 U8863 ( .IN1(n9142), .IN2(n9108), .QN(n9148) );
  NOR2X0 U8864 ( .IN1(n9083), .IN2(n4548), .QN(n9095) );
  NAND2X0 U8865 ( .IN1(n9149), .IN2(n7751), .QN(n9083) );
  NOR2X0 U8866 ( .IN1(g1249), .IN2(n498), .QN(n9149) );
  NAND2X0 U8867 ( .IN1(n9150), .IN2(n9108), .QN(n9146) );
  NAND2X0 U8868 ( .IN1(n9109), .IN2(n9151), .QN(n9145) );
  NOR2X0 U8869 ( .IN1(n9108), .IN2(n9142), .QN(n9109) );
  INVX0 U8870 ( .INP(n9152), .ZN(n9142) );
  INVX0 U8871 ( .INP(n9153), .ZN(n3938) );
  NAND2X0 U8872 ( .IN1(n3896), .IN2(g88), .QN(n4528) );
  NAND2X0 U8873 ( .IN1(n3890), .IN2(g1462), .QN(n4527) );
  NAND2X0 U8874 ( .IN1(n3887), .IN2(test_so78), .QN(n4526) );
  NAND3X0 U8875 ( .IN1(n9154), .IN2(n9155), .IN3(n9156), .QN(n3478) );
  NAND3X0 U8876 ( .IN1(n9157), .IN2(n9158), .IN3(n9159), .QN(n3469) );
  NAND3X0 U8877 ( .IN1(n9160), .IN2(n9161), .IN3(n9162), .QN(n3457) );
  NAND3X0 U8878 ( .IN1(n9163), .IN2(n9164), .IN3(n9165), .QN(n3445) );
  NAND2X0 U8879 ( .IN1(n3692), .IN2(test_so15), .QN(n4521) );
  NAND2X0 U8880 ( .IN1(n3686), .IN2(g1453), .QN(n4523) );
  NAND2X0 U8881 ( .IN1(n3683), .IN2(g2147), .QN(n4522) );
  NAND2X0 U8882 ( .IN1(n9166), .IN2(n9167), .QN(n3254) );
  NAND2X0 U8883 ( .IN1(n9168), .IN2(n9169), .QN(n9166) );
  INVX0 U8884 ( .INP(n9170), .ZN(n9168) );
  INVX0 U8885 ( .INP(n9171), .ZN(n309) );
  XOR2X1 U8886 ( .IN1(n9172), .IN2(n9173), .Q(n2800) );
  NAND2X0 U8887 ( .IN1(n9174), .IN2(n9175), .QN(n9172) );
  NAND2X0 U8888 ( .IN1(n9173), .IN2(n9176), .QN(n9175) );
  NAND3X0 U8889 ( .IN1(n9177), .IN2(n9178), .IN3(n9179), .QN(n9176) );
  NAND2X0 U8890 ( .IN1(n9180), .IN2(n9181), .QN(n9178) );
  NAND3X0 U8891 ( .IN1(n9182), .IN2(g996), .IN3(n9183), .QN(n9177) );
  NAND3X0 U8892 ( .IN1(n9184), .IN2(n9179), .IN3(n9185), .QN(n9174) );
  INVX0 U8893 ( .INP(g24734), .ZN(n279) );
  XOR2X1 U8894 ( .IN1(n8571), .IN2(n9186), .Q(n2719) );
  INVX0 U8895 ( .INP(g25435), .ZN(n270) );
  XOR2X1 U8896 ( .IN1(n9187), .IN2(n9188), .Q(n2686) );
  XOR2X1 U8897 ( .IN1(n8665), .IN2(n9189), .Q(n2671) );
  XOR2X1 U8898 ( .IN1(n9181), .IN2(n9190), .Q(n2616) );
  NAND2X0 U8899 ( .IN1(n9191), .IN2(n9192), .QN(n9190) );
  NAND2X0 U8900 ( .IN1(n9193), .IN2(n9194), .QN(n9192) );
  NAND4X0 U8901 ( .IN1(n9195), .IN2(n9196), .IN3(n9197), .IN4(n9179), .QN(
        n9191) );
  NAND3X0 U8902 ( .IN1(n9173), .IN2(n9198), .IN3(n9184), .QN(n9197) );
  NOR3X0 U8903 ( .IN1(n9199), .IN2(n9183), .IN3(n9200), .QN(n9184) );
  NAND2X0 U8904 ( .IN1(n9201), .IN2(n9181), .QN(n9196) );
  NAND2X0 U8905 ( .IN1(n9202), .IN2(n9183), .QN(n9195) );
  NAND2X0 U8906 ( .IN1(n9203), .IN2(n9204), .QN(n9202) );
  NAND2X0 U8907 ( .IN1(n9173), .IN2(n9205), .QN(n9204) );
  NAND3X0 U8908 ( .IN1(n9206), .IN2(n9198), .IN3(n9207), .QN(n9205) );
  INVX0 U8909 ( .INP(n9180), .ZN(n9207) );
  NAND2X0 U8910 ( .IN1(n9208), .IN2(n9209), .QN(n9180) );
  NAND2X0 U8911 ( .IN1(n9199), .IN2(n3102), .QN(n9209) );
  INVX0 U8912 ( .INP(n9210), .ZN(n9199) );
  NAND2X0 U8913 ( .IN1(n9211), .IN2(n9212), .QN(n9206) );
  NAND2X0 U8914 ( .IN1(n9213), .IN2(n9185), .QN(n9203) );
  NAND2X0 U8915 ( .IN1(n9214), .IN2(n9208), .QN(n9213) );
  NOR2X0 U8916 ( .IN1(n8683), .IN2(n8681), .QN(n2446) );
  NOR2X0 U8917 ( .IN1(g557), .IN2(n9215), .QN(n8681) );
  INVX0 U8918 ( .INP(n9216), .ZN(n9215) );
  NAND2X0 U8919 ( .IN1(n8036), .IN2(n8091), .QN(n9216) );
  NAND2X0 U8920 ( .IN1(n8091), .IN2(n9217), .QN(n8683) );
  NAND2X0 U8921 ( .IN1(n4360), .IN2(n8036), .QN(n9217) );
  NAND2X0 U8922 ( .IN1(g499), .IN2(n9218), .QN(n2445) );
  NAND4X0 U8923 ( .IN1(n9219), .IN2(n9220), .IN3(n9221), .IN4(n8803), .QN(
        n9218) );
  NAND4X0 U8924 ( .IN1(n9222), .IN2(n8768), .IN3(n9223), .IN4(n9224), .QN(
        n8803) );
  NOR4X0 U8925 ( .IN1(n9225), .IN2(n8747), .IN3(n8782), .IN4(n8753), .QN(n9224) );
  NAND3X0 U8926 ( .IN1(n8757), .IN2(n9226), .IN3(n8777), .QN(n9225) );
  NAND3X0 U8927 ( .IN1(n9227), .IN2(n9228), .IN3(n9229), .QN(n9226) );
  NAND2X0 U8928 ( .IN1(n7956), .IN2(g6911), .QN(n9229) );
  NAND2X0 U8929 ( .IN1(n7959), .IN2(g629), .QN(n9228) );
  NAND2X0 U8930 ( .IN1(n7868), .IN2(g6677), .QN(n9227) );
  NOR3X0 U8931 ( .IN1(n8762), .IN2(n8772), .IN3(n9230), .QN(n9223) );
  NOR2X0 U8932 ( .IN1(n8801), .IN2(n8792), .QN(n9222) );
  INVX0 U8933 ( .INP(n8802), .ZN(n8801) );
  NAND2X0 U8934 ( .IN1(n7501), .IN2(g629), .QN(n9221) );
  NAND2X0 U8935 ( .IN1(n7497), .IN2(g6677), .QN(n9220) );
  NAND2X0 U8936 ( .IN1(n7496), .IN2(g6911), .QN(n9219) );
  INVX0 U8937 ( .INP(g26135), .ZN(n244) );
  NAND2X0 U8938 ( .IN1(g2574), .IN2(n9231), .QN(n2374) );
  NAND4X0 U8939 ( .IN1(n9232), .IN2(n9233), .IN3(n9234), .IN4(n8920), .QN(
        n9231) );
  NAND4X0 U8940 ( .IN1(n9235), .IN2(n8900), .IN3(n9236), .IN4(n9237), .QN(
        n8920) );
  NOR4X0 U8941 ( .IN1(n9238), .IN2(n8896), .IN3(n8867), .IN4(n8891), .QN(n9237) );
  NAND3X0 U8942 ( .IN1(n8875), .IN2(n9239), .IN3(n8886), .QN(n9238) );
  NAND3X0 U8943 ( .IN1(n9240), .IN2(n9241), .IN3(n9242), .QN(n9239) );
  NAND2X0 U8944 ( .IN1(n7953), .IN2(g7487), .QN(n9242) );
  NAND2X0 U8945 ( .IN1(g2703), .IN2(n8101), .QN(n9241) );
  NAND2X0 U8946 ( .IN1(n7865), .IN2(g7425), .QN(n9240) );
  NOR3X0 U8947 ( .IN1(n8881), .IN2(n8918), .IN3(n9243), .QN(n9236) );
  NOR2X0 U8948 ( .IN1(n8911), .IN2(n8871), .QN(n9235) );
  INVX0 U8949 ( .INP(n8912), .ZN(n8911) );
  NAND2X0 U8950 ( .IN1(n7498), .IN2(g2703), .QN(n9234) );
  NAND2X0 U8951 ( .IN1(n7491), .IN2(g7425), .QN(n9233) );
  NAND2X0 U8952 ( .IN1(n7490), .IN2(g7487), .QN(n9232) );
  NOR2X0 U8953 ( .IN1(n8811), .IN2(n8809), .QN(n2361) );
  NOR2X0 U8954 ( .IN1(g2631), .IN2(n9244), .QN(n8809) );
  INVX0 U8955 ( .INP(n9245), .ZN(n9244) );
  NAND2X0 U8956 ( .IN1(n8039), .IN2(n4303), .QN(n9245) );
  NAND2X0 U8957 ( .IN1(n4303), .IN2(n9246), .QN(n8811) );
  NAND2X0 U8958 ( .IN1(n4352), .IN2(n8039), .QN(n9246) );
  NAND2X0 U8959 ( .IN1(g1880), .IN2(n9247), .QN(n2302) );
  NAND4X0 U8960 ( .IN1(n9248), .IN2(n9249), .IN3(n9250), .IN4(n9035), .QN(
        n9247) );
  NAND4X0 U8961 ( .IN1(n9251), .IN2(n9016), .IN3(n9252), .IN4(n9253), .QN(
        n9035) );
  NOR4X0 U8962 ( .IN1(n9254), .IN2(n9003), .IN3(n8991), .IN4(n9012), .QN(n9253) );
  NAND3X0 U8963 ( .IN1(n9006), .IN2(n9255), .IN3(n8979), .QN(n9254) );
  NAND3X0 U8964 ( .IN1(n9256), .IN2(n9257), .IN3(n9258), .QN(n9255) );
  NAND2X0 U8965 ( .IN1(n7954), .IN2(g7357), .QN(n9258) );
  NAND2X0 U8966 ( .IN1(n7957), .IN2(g2009), .QN(n9257) );
  NAND2X0 U8967 ( .IN1(n7866), .IN2(g7229), .QN(n9256) );
  INVX0 U8968 ( .INP(n9007), .ZN(n9006) );
  NOR3X0 U8969 ( .IN1(n8996), .IN2(n9033), .IN3(n9259), .QN(n9252) );
  NOR2X0 U8970 ( .IN1(n9026), .IN2(n8986), .QN(n9251) );
  INVX0 U8971 ( .INP(n9027), .ZN(n9026) );
  NAND2X0 U8972 ( .IN1(n7499), .IN2(g2009), .QN(n9250) );
  NAND2X0 U8973 ( .IN1(n7493), .IN2(g7229), .QN(n9249) );
  NAND2X0 U8974 ( .IN1(n7492), .IN2(g7357), .QN(n9248) );
  NOR2X0 U8975 ( .IN1(n8928), .IN2(n8926), .QN(n2289) );
  NOR2X0 U8976 ( .IN1(g1937), .IN2(n9260), .QN(n8926) );
  INVX0 U8977 ( .INP(n9261), .ZN(n9260) );
  NAND2X0 U8978 ( .IN1(n8038), .IN2(n4297), .QN(n9261) );
  NAND2X0 U8979 ( .IN1(n4297), .IN2(n9262), .QN(n8928) );
  NAND2X0 U8980 ( .IN1(n4311), .IN2(n8038), .QN(n9262) );
  NAND2X0 U8981 ( .IN1(g1186), .IN2(n9263), .QN(n2230) );
  NAND4X0 U8982 ( .IN1(n9264), .IN2(n9265), .IN3(n9266), .IN4(n9152), .QN(
        n9263) );
  NAND4X0 U8983 ( .IN1(n9267), .IN2(n9133), .IN3(n9268), .IN4(n9269), .QN(
        n9152) );
  NOR4X0 U8984 ( .IN1(n9270), .IN2(n9119), .IN3(n9110), .IN4(n9129), .QN(n9269) );
  NAND3X0 U8985 ( .IN1(n9123), .IN2(n9271), .IN3(n9096), .QN(n9270) );
  NAND3X0 U8986 ( .IN1(n9272), .IN2(n9273), .IN3(n9274), .QN(n9271) );
  NAND2X0 U8987 ( .IN1(n7955), .IN2(g7161), .QN(n9274) );
  NAND2X0 U8988 ( .IN1(n7958), .IN2(g1315), .QN(n9273) );
  NAND2X0 U8989 ( .IN1(n7867), .IN2(g6979), .QN(n9272) );
  INVX0 U8990 ( .INP(n9124), .ZN(n9123) );
  NOR3X0 U8991 ( .IN1(n9113), .IN2(n9150), .IN3(n9275), .QN(n9268) );
  NOR2X0 U8992 ( .IN1(n9143), .IN2(n9103), .QN(n9267) );
  NAND2X0 U8993 ( .IN1(n7500), .IN2(g1315), .QN(n9266) );
  NAND2X0 U8994 ( .IN1(n7495), .IN2(g6979), .QN(n9265) );
  NAND2X0 U8995 ( .IN1(n7494), .IN2(g7161), .QN(n9264) );
  NOR2X0 U8996 ( .IN1(n9043), .IN2(n9041), .QN(n2217) );
  NOR2X0 U8997 ( .IN1(g1243), .IN2(n9276), .QN(n9041) );
  INVX0 U8998 ( .INP(n9277), .ZN(n9276) );
  NAND2X0 U8999 ( .IN1(n8037), .IN2(n4304), .QN(n9277) );
  NAND2X0 U9000 ( .IN1(n4304), .IN2(n9278), .QN(n9043) );
  NAND2X0 U9001 ( .IN1(n4353), .IN2(n8037), .QN(n9278) );
  INVX0 U9002 ( .INP(n9279), .ZN(n1540) );
  NAND3X0 U9003 ( .IN1(n9280), .IN2(n1543), .IN3(n8728), .QN(n9279) );
  NAND2X0 U9004 ( .IN1(n9281), .IN2(n4350), .QN(n9280) );
  NAND2X0 U9005 ( .IN1(g3018), .IN2(n8729), .QN(n9281) );
  INVX0 U9006 ( .INP(n9282), .ZN(n1538) );
  NAND3X0 U9007 ( .IN1(n9283), .IN2(n4066), .IN3(n9284), .QN(n9282) );
  NAND2X0 U9008 ( .IN1(n9285), .IN2(n8035), .QN(n9284) );
  NAND2X0 U9009 ( .IN1(n7909), .IN2(n9286), .QN(n9285) );
  INVX0 U9010 ( .INP(n9287), .ZN(n1503) );
  NAND3X0 U9011 ( .IN1(n9288), .IN2(n9289), .IN3(n9290), .QN(n9287) );
  NAND2X0 U9012 ( .IN1(n9291), .IN2(n4407), .QN(n9288) );
  NAND2X0 U9013 ( .IN1(g2734), .IN2(n9292), .QN(n9291) );
  INVX0 U9014 ( .INP(n9293), .ZN(n1502) );
  NAND3X0 U9015 ( .IN1(n9294), .IN2(n9289), .IN3(n9295), .QN(n9293) );
  NAND2X0 U9016 ( .IN1(n9296), .IN2(n4472), .QN(n9294) );
  NAND2X0 U9017 ( .IN1(g2714), .IN2(n9297), .QN(n9296) );
  INVX0 U9018 ( .INP(n9298), .ZN(n1427) );
  NOR2X0 U9019 ( .IN1(n9299), .IN2(n9300), .QN(n9298) );
  NOR2X0 U9020 ( .IN1(g2624), .IN2(n7961), .QN(n9300) );
  INVX0 U9021 ( .INP(n9301), .ZN(n1423) );
  INVX0 U9022 ( .INP(n9302), .ZN(n1402) );
  INVX0 U9023 ( .INP(n9303), .ZN(n1261) );
  NOR3X0 U9024 ( .IN1(n9304), .IN2(n9305), .IN3(n9306), .QN(n1215) );
  NOR2X0 U9025 ( .IN1(n9307), .IN2(g2052), .QN(n9304) );
  NOR2X0 U9026 ( .IN1(n4399), .IN2(n9308), .QN(n9307) );
  INVX0 U9027 ( .INP(n9309), .ZN(n1214) );
  NAND3X0 U9028 ( .IN1(n9310), .IN2(n9311), .IN3(n9312), .QN(n9309) );
  NAND2X0 U9029 ( .IN1(n9313), .IN2(n4474), .QN(n9310) );
  NAND2X0 U9030 ( .IN1(g2020), .IN2(n9314), .QN(n9313) );
  NOR2X0 U9031 ( .IN1(n9305), .IN2(n9315), .QN(n1186) );
  INVX0 U9032 ( .INP(n9316), .ZN(n9315) );
  NAND2X0 U9033 ( .IN1(n9317), .IN2(n7954), .QN(n9316) );
  INVX0 U9034 ( .INP(n9318), .ZN(n1141) );
  NOR2X0 U9035 ( .IN1(n9319), .IN2(n9320), .QN(n9318) );
  NOR2X0 U9036 ( .IN1(g1930), .IN2(n7969), .QN(n9320) );
  INVX0 U9037 ( .INP(n9321), .ZN(n1137) );
  INVX0 U9038 ( .INP(n9322), .ZN(n1114) );
  NAND2X0 U9039 ( .IN1(n9323), .IN2(n9324), .QN(g30801) );
  INVX0 U9040 ( .INP(n9325), .ZN(n9324) );
  NOR2X0 U9041 ( .IN1(g3109), .IN2(n4334), .QN(n9325) );
  NAND2X0 U9042 ( .IN1(g30072), .IN2(g3109), .QN(n9323) );
  NAND2X0 U9043 ( .IN1(n9326), .IN2(n9327), .QN(g30798) );
  NAND2X0 U9044 ( .IN1(n4383), .IN2(g3107), .QN(n9327) );
  NAND2X0 U9045 ( .IN1(g30072), .IN2(g8030), .QN(n9326) );
  NAND2X0 U9046 ( .IN1(n9328), .IN2(n9329), .QN(g30796) );
  NAND2X0 U9047 ( .IN1(n4382), .IN2(g3106), .QN(n9329) );
  NAND2X0 U9048 ( .IN1(g30072), .IN2(g8106), .QN(n9328) );
  NAND2X0 U9049 ( .IN1(n9330), .IN2(n9331), .QN(g30709) );
  NAND2X0 U9050 ( .IN1(n9332), .IN2(g7264), .QN(n9331) );
  NAND2X0 U9051 ( .IN1(n4524), .IN2(g2391), .QN(n9330) );
  NAND2X0 U9052 ( .IN1(n9333), .IN2(n9334), .QN(g30708) );
  NAND2X0 U9053 ( .IN1(n9335), .IN2(n4618), .QN(n9334) );
  NAND2X0 U9054 ( .IN1(n4511), .IN2(g1698), .QN(n9333) );
  NAND2X0 U9055 ( .IN1(n9336), .IN2(n9337), .QN(g30707) );
  NAND2X0 U9056 ( .IN1(n9332), .IN2(g5555), .QN(n9337) );
  NAND2X0 U9057 ( .IN1(n4516), .IN2(g2390), .QN(n9336) );
  NAND2X0 U9058 ( .IN1(n9338), .IN2(n9339), .QN(g30706) );
  NAND2X0 U9059 ( .IN1(n9335), .IN2(g7014), .QN(n9339) );
  NAND2X0 U9060 ( .IN1(n4525), .IN2(g1697), .QN(n9338) );
  NAND2X0 U9061 ( .IN1(n9340), .IN2(n9341), .QN(g30705) );
  NAND2X0 U9062 ( .IN1(n4381), .IN2(g1004), .QN(n9341) );
  NAND2X0 U9063 ( .IN1(n2594), .IN2(g1088), .QN(n9340) );
  NAND2X0 U9064 ( .IN1(n9342), .IN2(n9343), .QN(g30704) );
  NAND2X0 U9065 ( .IN1(n9335), .IN2(g5511), .QN(n9343) );
  INVX0 U9066 ( .INP(n9344), .ZN(n9335) );
  NAND2X0 U9067 ( .IN1(n9345), .IN2(n9346), .QN(n9344) );
  XOR2X1 U9068 ( .IN1(n9347), .IN2(n9348), .Q(n9345) );
  NAND2X0 U9069 ( .IN1(n9349), .IN2(n9350), .QN(n9348) );
  NAND2X0 U9070 ( .IN1(n9351), .IN2(n9352), .QN(n9350) );
  NAND4X0 U9071 ( .IN1(n9353), .IN2(n9354), .IN3(n9355), .IN4(n9356), .QN(
        n9349) );
  NAND3X0 U9072 ( .IN1(n9357), .IN2(n9358), .IN3(n9359), .QN(n9355) );
  NAND2X0 U9073 ( .IN1(n9360), .IN2(n9347), .QN(n9354) );
  INVX0 U9074 ( .INP(n9361), .ZN(n9360) );
  NAND2X0 U9075 ( .IN1(n9362), .IN2(n9363), .QN(n9353) );
  NAND2X0 U9076 ( .IN1(n9364), .IN2(n9365), .QN(n9362) );
  NAND2X0 U9077 ( .IN1(n9357), .IN2(n9366), .QN(n9365) );
  NAND3X0 U9078 ( .IN1(n9367), .IN2(n9358), .IN3(n9368), .QN(n9366) );
  INVX0 U9079 ( .INP(n9369), .ZN(n9368) );
  NAND2X0 U9080 ( .IN1(n9370), .IN2(n9361), .QN(n9367) );
  NAND2X0 U9081 ( .IN1(n9371), .IN2(n9372), .QN(n9364) );
  NAND2X0 U9082 ( .IN1(n9373), .IN2(n9374), .QN(n9371) );
  NAND2X0 U9083 ( .IN1(n4518), .IN2(g1696), .QN(n9342) );
  NAND2X0 U9084 ( .IN1(n9375), .IN2(n9376), .QN(g30703) );
  NAND2X0 U9085 ( .IN1(n4364), .IN2(g1003), .QN(n9376) );
  NAND2X0 U9086 ( .IN1(n2594), .IN2(g6712), .QN(n9375) );
  NAND2X0 U9087 ( .IN1(n9377), .IN2(n9378), .QN(g30702) );
  NAND2X0 U9088 ( .IN1(n9379), .IN2(n4640), .QN(n9378) );
  NAND2X0 U9089 ( .IN1(n4506), .IN2(g317), .QN(n9377) );
  NAND2X0 U9090 ( .IN1(n9380), .IN2(n9381), .QN(g30701) );
  NAND2X0 U9091 ( .IN1(n4363), .IN2(g1002), .QN(n9381) );
  NAND2X0 U9092 ( .IN1(n2594), .IN2(g5472), .QN(n9380) );
  NAND2X0 U9093 ( .IN1(n9382), .IN2(n9383), .QN(g30700) );
  NAND2X0 U9094 ( .IN1(n9379), .IN2(g6447), .QN(n9383) );
  NAND2X0 U9095 ( .IN1(test_so18), .IN2(n4499), .QN(n9382) );
  NAND2X0 U9096 ( .IN1(n9384), .IN2(n9385), .QN(g30699) );
  NAND2X0 U9097 ( .IN1(n9379), .IN2(g5437), .QN(n9385) );
  INVX0 U9098 ( .INP(n9386), .ZN(n9379) );
  NAND2X0 U9099 ( .IN1(n9387), .IN2(n9388), .QN(n9386) );
  XOR2X1 U9100 ( .IN1(n9389), .IN2(n9390), .Q(n9387) );
  NAND2X0 U9101 ( .IN1(n9391), .IN2(n9392), .QN(n9390) );
  NAND2X0 U9102 ( .IN1(n9393), .IN2(n9394), .QN(n9392) );
  NAND4X0 U9103 ( .IN1(n9395), .IN2(n9396), .IN3(n9397), .IN4(n9398), .QN(
        n9391) );
  NAND3X0 U9104 ( .IN1(n9399), .IN2(n9400), .IN3(n9401), .QN(n9397) );
  NAND2X0 U9105 ( .IN1(n9402), .IN2(n9389), .QN(n9396) );
  INVX0 U9106 ( .INP(n9403), .ZN(n9402) );
  NAND2X0 U9107 ( .IN1(n9404), .IN2(n9405), .QN(n9395) );
  NAND2X0 U9108 ( .IN1(n9406), .IN2(n9407), .QN(n9404) );
  NAND2X0 U9109 ( .IN1(n9399), .IN2(n9408), .QN(n9407) );
  NAND3X0 U9110 ( .IN1(n9409), .IN2(n9400), .IN3(n9410), .QN(n9408) );
  INVX0 U9111 ( .INP(n9411), .ZN(n9410) );
  NAND2X0 U9112 ( .IN1(n9412), .IN2(n9403), .QN(n9409) );
  NAND2X0 U9113 ( .IN1(n9413), .IN2(n9414), .QN(n9406) );
  NAND2X0 U9114 ( .IN1(n9415), .IN2(n9416), .QN(n9413) );
  NAND2X0 U9115 ( .IN1(n4520), .IN2(g315), .QN(n9384) );
  NAND2X0 U9116 ( .IN1(n9417), .IN2(n9418), .QN(g30695) );
  NAND2X0 U9117 ( .IN1(n4367), .IN2(g2276), .QN(n9418) );
  NAND2X0 U9118 ( .IN1(n9419), .IN2(g2241), .QN(n9417) );
  NAND2X0 U9119 ( .IN1(n9420), .IN2(n9421), .QN(g30694) );
  NAND2X0 U9120 ( .IN1(n4367), .IN2(g2348), .QN(n9421) );
  NAND2X0 U9121 ( .IN1(n9422), .IN2(g2241), .QN(n9420) );
  NAND2X0 U9122 ( .IN1(n9423), .IN2(n9424), .QN(g30693) );
  NAND2X0 U9123 ( .IN1(g2273), .IN2(n8070), .QN(n9424) );
  NAND2X0 U9124 ( .IN1(test_so73), .IN2(n9419), .QN(n9423) );
  NAND2X0 U9125 ( .IN1(n9425), .IN2(n9426), .QN(g30692) );
  NAND2X0 U9126 ( .IN1(n4368), .IN2(g1582), .QN(n9426) );
  NAND2X0 U9127 ( .IN1(n9427), .IN2(g1547), .QN(n9425) );
  NAND2X0 U9128 ( .IN1(n9428), .IN2(n9429), .QN(g30691) );
  NAND2X0 U9129 ( .IN1(g2345), .IN2(n8070), .QN(n9429) );
  NAND2X0 U9130 ( .IN1(n9422), .IN2(test_so73), .QN(n9428) );
  NAND2X0 U9131 ( .IN1(n9430), .IN2(n9431), .QN(g30690) );
  NAND2X0 U9132 ( .IN1(n4324), .IN2(g2270), .QN(n9431) );
  NAND2X0 U9133 ( .IN1(n9419), .IN2(g6837), .QN(n9430) );
  NAND3X0 U9134 ( .IN1(n9432), .IN2(n9433), .IN3(n9434), .QN(n9419) );
  NAND2X0 U9135 ( .IN1(n9435), .IN2(n9436), .QN(n9433) );
  XOR2X1 U9136 ( .IN1(n9437), .IN2(n9438), .Q(n9435) );
  NAND2X0 U9137 ( .IN1(n9439), .IN2(g2175), .QN(n9432) );
  NAND2X0 U9138 ( .IN1(n9440), .IN2(n9441), .QN(g30689) );
  NAND2X0 U9139 ( .IN1(n4368), .IN2(g1654), .QN(n9441) );
  NAND2X0 U9140 ( .IN1(n9442), .IN2(g1547), .QN(n9440) );
  NAND2X0 U9141 ( .IN1(n9443), .IN2(n9444), .QN(g30688) );
  NAND2X0 U9142 ( .IN1(n4515), .IN2(g1579), .QN(n9444) );
  NAND2X0 U9143 ( .IN1(n9427), .IN2(g6782), .QN(n9443) );
  NAND2X0 U9144 ( .IN1(n9445), .IN2(n9446), .QN(g30687) );
  NAND2X0 U9145 ( .IN1(g888), .IN2(n8071), .QN(n9446) );
  NAND2X0 U9146 ( .IN1(test_so31), .IN2(n9447), .QN(n9445) );
  NAND2X0 U9147 ( .IN1(n9448), .IN2(n9449), .QN(g30686) );
  NAND2X0 U9148 ( .IN1(n4324), .IN2(g2342), .QN(n9449) );
  NAND2X0 U9149 ( .IN1(n9422), .IN2(g6837), .QN(n9448) );
  INVX0 U9150 ( .INP(n9450), .ZN(n9422) );
  NAND3X0 U9151 ( .IN1(n9451), .IN2(n9452), .IN3(n9453), .QN(n9450) );
  NAND2X0 U9152 ( .IN1(n9439), .IN2(n9454), .QN(n9453) );
  NAND2X0 U9153 ( .IN1(n9455), .IN2(n9436), .QN(n9451) );
  XOR2X1 U9154 ( .IN1(n8654), .IN2(n2669), .Q(n9455) );
  NAND2X0 U9155 ( .IN1(n9456), .IN2(n9457), .QN(g30684) );
  NAND2X0 U9156 ( .IN1(n4515), .IN2(g1651), .QN(n9457) );
  NAND2X0 U9157 ( .IN1(n9442), .IN2(g6782), .QN(n9456) );
  NAND2X0 U9158 ( .IN1(n9458), .IN2(n9459), .QN(g30683) );
  NAND2X0 U9159 ( .IN1(n4317), .IN2(g1576), .QN(n9459) );
  NAND2X0 U9160 ( .IN1(n9427), .IN2(g6573), .QN(n9458) );
  NAND3X0 U9161 ( .IN1(n9460), .IN2(n9461), .IN3(n9462), .QN(n9427) );
  NAND2X0 U9162 ( .IN1(n9463), .IN2(n9464), .QN(n9461) );
  XNOR2X1 U9163 ( .IN1(n9465), .IN2(n8637), .Q(n9463) );
  NAND2X0 U9164 ( .IN1(n9466), .IN2(g1481), .QN(n9460) );
  NAND2X0 U9165 ( .IN1(n9467), .IN2(n9468), .QN(g30682) );
  NAND2X0 U9166 ( .IN1(g960), .IN2(n8071), .QN(n9468) );
  NAND2X0 U9167 ( .IN1(n9469), .IN2(test_so31), .QN(n9467) );
  NAND2X0 U9168 ( .IN1(n9470), .IN2(n9471), .QN(g30681) );
  NAND2X0 U9169 ( .IN1(n4312), .IN2(g885), .QN(n9471) );
  NAND2X0 U9170 ( .IN1(n9447), .IN2(g6518), .QN(n9470) );
  NAND2X0 U9171 ( .IN1(n9472), .IN2(n9473), .QN(g30680) );
  NAND2X0 U9172 ( .IN1(n4369), .IN2(g201), .QN(n9473) );
  NAND2X0 U9173 ( .IN1(n9474), .IN2(g165), .QN(n9472) );
  NAND2X0 U9174 ( .IN1(n9475), .IN2(n9476), .QN(g30679) );
  NAND2X0 U9175 ( .IN1(n4367), .IN2(g2321), .QN(n9476) );
  NAND2X0 U9176 ( .IN1(n9477), .IN2(g2241), .QN(n9475) );
  NAND2X0 U9177 ( .IN1(n9478), .IN2(n9479), .QN(g30678) );
  NAND2X0 U9178 ( .IN1(n4317), .IN2(g1648), .QN(n9479) );
  NAND2X0 U9179 ( .IN1(n9442), .IN2(g6573), .QN(n9478) );
  INVX0 U9180 ( .INP(n9480), .ZN(n9442) );
  NAND3X0 U9181 ( .IN1(n9481), .IN2(n9482), .IN3(n9483), .QN(n9480) );
  NAND2X0 U9182 ( .IN1(n9466), .IN2(n9484), .QN(n9483) );
  NAND2X0 U9183 ( .IN1(n9485), .IN2(n9464), .QN(n9481) );
  XOR2X1 U9184 ( .IN1(n8630), .IN2(n2684), .Q(n9485) );
  NAND2X0 U9185 ( .IN1(n9486), .IN2(n9487), .QN(g30677) );
  NAND2X0 U9186 ( .IN1(n4312), .IN2(g957), .QN(n9487) );
  NAND2X0 U9187 ( .IN1(n9469), .IN2(g6518), .QN(n9486) );
  NAND2X0 U9188 ( .IN1(n9488), .IN2(n9489), .QN(g30676) );
  NAND2X0 U9189 ( .IN1(n4323), .IN2(g882), .QN(n9489) );
  NAND2X0 U9190 ( .IN1(n9447), .IN2(g6368), .QN(n9488) );
  NAND3X0 U9191 ( .IN1(n9490), .IN2(n9491), .IN3(n9492), .QN(n9447) );
  NAND2X0 U9192 ( .IN1(n9493), .IN2(g793), .QN(n9492) );
  NAND2X0 U9193 ( .IN1(n9494), .IN2(n9495), .QN(n9490) );
  XNOR2X1 U9194 ( .IN1(n9496), .IN2(n8599), .Q(n9494) );
  NAND2X0 U9195 ( .IN1(n9497), .IN2(n9498), .QN(g30675) );
  NAND2X0 U9196 ( .IN1(n4369), .IN2(g273), .QN(n9498) );
  NAND2X0 U9197 ( .IN1(n9499), .IN2(g165), .QN(n9497) );
  NAND2X0 U9198 ( .IN1(n9500), .IN2(n9501), .QN(g30674) );
  NAND2X0 U9199 ( .IN1(n4512), .IN2(g198), .QN(n9501) );
  NAND2X0 U9200 ( .IN1(n9474), .IN2(g6313), .QN(n9500) );
  NAND2X0 U9201 ( .IN1(n9502), .IN2(n9503), .QN(g30673) );
  NAND2X0 U9202 ( .IN1(g2318), .IN2(n8070), .QN(n9503) );
  NAND2X0 U9203 ( .IN1(n9477), .IN2(test_so73), .QN(n9502) );
  NAND2X0 U9204 ( .IN1(n9504), .IN2(n9505), .QN(g30672) );
  NAND2X0 U9205 ( .IN1(n4367), .IN2(g2312), .QN(n9505) );
  NAND2X0 U9206 ( .IN1(n9506), .IN2(g2241), .QN(n9504) );
  NAND2X0 U9207 ( .IN1(n9507), .IN2(n9508), .QN(g30671) );
  NAND2X0 U9208 ( .IN1(n4368), .IN2(g1627), .QN(n9508) );
  NAND2X0 U9209 ( .IN1(n9509), .IN2(g1547), .QN(n9507) );
  NAND2X0 U9210 ( .IN1(n9510), .IN2(n9511), .QN(g30670) );
  NAND2X0 U9211 ( .IN1(n4323), .IN2(g954), .QN(n9511) );
  NAND2X0 U9212 ( .IN1(n9469), .IN2(g6368), .QN(n9510) );
  INVX0 U9213 ( .INP(n9512), .ZN(n9469) );
  NAND3X0 U9214 ( .IN1(n9513), .IN2(n9514), .IN3(n9515), .QN(n9512) );
  NAND2X0 U9215 ( .IN1(n9516), .IN2(n9493), .QN(n9515) );
  NAND2X0 U9216 ( .IN1(n9495), .IN2(n9517), .QN(n9513) );
  XNOR2X1 U9217 ( .IN1(n8605), .IN2(n9518), .Q(n9517) );
  NOR2X0 U9218 ( .IN1(n9519), .IN2(n9520), .QN(n9518) );
  XOR2X1 U9219 ( .IN1(n9521), .IN2(n8607), .Q(n9519) );
  NAND2X0 U9220 ( .IN1(n9522), .IN2(n9523), .QN(g30669) );
  NAND2X0 U9221 ( .IN1(n4512), .IN2(g270), .QN(n9523) );
  NAND2X0 U9222 ( .IN1(n9499), .IN2(g6313), .QN(n9522) );
  NAND2X0 U9223 ( .IN1(n9524), .IN2(n9525), .QN(g30668) );
  NAND2X0 U9224 ( .IN1(n4318), .IN2(g195), .QN(n9525) );
  NAND2X0 U9225 ( .IN1(n9474), .IN2(g6231), .QN(n9524) );
  NAND3X0 U9226 ( .IN1(n9526), .IN2(n9527), .IN3(n9528), .QN(n9474) );
  NAND2X0 U9227 ( .IN1(n9529), .IN2(g105), .QN(n9528) );
  NAND2X0 U9228 ( .IN1(n9530), .IN2(n9531), .QN(n9526) );
  XNOR2X1 U9229 ( .IN1(n9532), .IN2(n8576), .Q(n9530) );
  NAND2X0 U9230 ( .IN1(n9533), .IN2(n9534), .QN(g30667) );
  NAND2X0 U9231 ( .IN1(n4324), .IN2(g2315), .QN(n9534) );
  NAND2X0 U9232 ( .IN1(n9477), .IN2(g6837), .QN(n9533) );
  INVX0 U9233 ( .INP(n9535), .ZN(n9477) );
  NAND3X0 U9234 ( .IN1(n9536), .IN2(n9452), .IN3(n9537), .QN(n9535) );
  NAND2X0 U9235 ( .IN1(n9439), .IN2(n4389), .QN(n9537) );
  NAND2X0 U9236 ( .IN1(n9436), .IN2(n9538), .QN(n9536) );
  XOR2X1 U9237 ( .IN1(n9539), .IN2(n9540), .Q(n9538) );
  NAND2X0 U9238 ( .IN1(n9541), .IN2(n9542), .QN(g30666) );
  NAND2X0 U9239 ( .IN1(g2309), .IN2(n8070), .QN(n9542) );
  NAND2X0 U9240 ( .IN1(n9506), .IN2(test_so73), .QN(n9541) );
  NAND2X0 U9241 ( .IN1(n9543), .IN2(n9544), .QN(g30665) );
  NAND2X0 U9242 ( .IN1(n4367), .IN2(g2303), .QN(n9544) );
  NAND2X0 U9243 ( .IN1(n9545), .IN2(g2241), .QN(n9543) );
  NAND2X0 U9244 ( .IN1(n9546), .IN2(n9547), .QN(g30664) );
  NAND2X0 U9245 ( .IN1(n4515), .IN2(g1624), .QN(n9547) );
  NAND2X0 U9246 ( .IN1(n9509), .IN2(g6782), .QN(n9546) );
  NAND2X0 U9247 ( .IN1(n9548), .IN2(n9549), .QN(g30663) );
  NAND2X0 U9248 ( .IN1(n4368), .IN2(g1618), .QN(n9549) );
  NAND2X0 U9249 ( .IN1(n9550), .IN2(g1547), .QN(n9548) );
  NAND2X0 U9250 ( .IN1(n9551), .IN2(n9552), .QN(g30662) );
  NAND2X0 U9251 ( .IN1(g933), .IN2(n8071), .QN(n9552) );
  NAND2X0 U9252 ( .IN1(n9553), .IN2(test_so31), .QN(n9551) );
  NAND2X0 U9253 ( .IN1(n9554), .IN2(n9555), .QN(g30661) );
  NAND2X0 U9254 ( .IN1(n4318), .IN2(g267), .QN(n9555) );
  NAND2X0 U9255 ( .IN1(n9499), .IN2(g6231), .QN(n9554) );
  INVX0 U9256 ( .INP(n9556), .ZN(n9499) );
  NAND3X0 U9257 ( .IN1(n9557), .IN2(n9558), .IN3(n9559), .QN(n9556) );
  NAND2X0 U9258 ( .IN1(n9560), .IN2(n9529), .QN(n9559) );
  NAND2X0 U9259 ( .IN1(n9561), .IN2(n9531), .QN(n9557) );
  XOR2X1 U9260 ( .IN1(n8563), .IN2(n2717), .Q(n9561) );
  NAND2X0 U9261 ( .IN1(n9562), .IN2(n9563), .QN(g30660) );
  NAND2X0 U9262 ( .IN1(n4324), .IN2(g2306), .QN(n9563) );
  NAND2X0 U9263 ( .IN1(n9506), .IN2(g6837), .QN(n9562) );
  INVX0 U9264 ( .INP(n9564), .ZN(n9506) );
  NAND3X0 U9265 ( .IN1(n9565), .IN2(n9452), .IN3(n9566), .QN(n9564) );
  NAND2X0 U9266 ( .IN1(n9439), .IN2(n4373), .QN(n9566) );
  NAND2X0 U9267 ( .IN1(n9567), .IN2(n4529), .QN(n9452) );
  NAND2X0 U9268 ( .IN1(n9436), .IN2(n9568), .QN(n9565) );
  XOR2X1 U9269 ( .IN1(n8669), .IN2(n9569), .Q(n9568) );
  INVX0 U9270 ( .INP(n9570), .ZN(n8669) );
  NAND2X0 U9271 ( .IN1(n9571), .IN2(n9572), .QN(g30659) );
  NAND2X0 U9272 ( .IN1(g2300), .IN2(n8070), .QN(n9572) );
  NAND2X0 U9273 ( .IN1(test_so73), .IN2(n9545), .QN(n9571) );
  NAND2X0 U9274 ( .IN1(n9573), .IN2(n9574), .QN(g30658) );
  NAND2X0 U9275 ( .IN1(n9509), .IN2(g6573), .QN(n9574) );
  INVX0 U9276 ( .INP(n9575), .ZN(n9509) );
  NAND3X0 U9277 ( .IN1(n9576), .IN2(n9482), .IN3(n9577), .QN(n9575) );
  NAND2X0 U9278 ( .IN1(n9466), .IN2(n4390), .QN(n9577) );
  NAND2X0 U9279 ( .IN1(n9464), .IN2(n9578), .QN(n9576) );
  XOR2X1 U9280 ( .IN1(n9579), .IN2(n8628), .Q(n9578) );
  NAND2X0 U9281 ( .IN1(test_so55), .IN2(n4317), .QN(n9573) );
  NAND2X0 U9282 ( .IN1(n9580), .IN2(n9581), .QN(g30657) );
  NAND2X0 U9283 ( .IN1(n4515), .IN2(g1615), .QN(n9581) );
  NAND2X0 U9284 ( .IN1(n9550), .IN2(g6782), .QN(n9580) );
  NAND2X0 U9285 ( .IN1(n9582), .IN2(n9583), .QN(g30656) );
  NAND2X0 U9286 ( .IN1(n4368), .IN2(g1609), .QN(n9583) );
  NAND2X0 U9287 ( .IN1(n9584), .IN2(g1547), .QN(n9582) );
  NAND2X0 U9288 ( .IN1(n9585), .IN2(n9586), .QN(g30655) );
  NAND2X0 U9289 ( .IN1(n4312), .IN2(g930), .QN(n9586) );
  NAND2X0 U9290 ( .IN1(n9553), .IN2(g6518), .QN(n9585) );
  NAND2X0 U9291 ( .IN1(n9587), .IN2(n9588), .QN(g30654) );
  NAND2X0 U9292 ( .IN1(test_so34), .IN2(n8071), .QN(n9588) );
  NAND2X0 U9293 ( .IN1(n9589), .IN2(test_so31), .QN(n9587) );
  NAND2X0 U9294 ( .IN1(n9590), .IN2(n9591), .QN(g30653) );
  NAND2X0 U9295 ( .IN1(n4369), .IN2(g246), .QN(n9591) );
  NAND2X0 U9296 ( .IN1(n9592), .IN2(g165), .QN(n9590) );
  NAND2X0 U9297 ( .IN1(n9593), .IN2(n9594), .QN(g30652) );
  NAND2X0 U9298 ( .IN1(n4324), .IN2(g2297), .QN(n9594) );
  NAND2X0 U9299 ( .IN1(n9545), .IN2(g6837), .QN(n9593) );
  NAND3X0 U9300 ( .IN1(n9595), .IN2(n9596), .IN3(n9434), .QN(n9545) );
  NAND2X0 U9301 ( .IN1(n9567), .IN2(n9597), .QN(n9434) );
  NAND2X0 U9302 ( .IN1(n9598), .IN2(n9436), .QN(n9596) );
  XNOR2X1 U9303 ( .IN1(n2670), .IN2(n8665), .Q(n9598) );
  NAND2X0 U9304 ( .IN1(n9599), .IN2(n9600), .QN(n2670) );
  XOR2X1 U9305 ( .IN1(n8659), .IN2(n9189), .Q(n9600) );
  NAND2X0 U9306 ( .IN1(n9439), .IN2(n9601), .QN(n9595) );
  NAND2X0 U9307 ( .IN1(n9602), .IN2(n9603), .QN(g30651) );
  NAND2X0 U9308 ( .IN1(n4317), .IN2(g1612), .QN(n9603) );
  NAND2X0 U9309 ( .IN1(n9550), .IN2(g6573), .QN(n9602) );
  INVX0 U9310 ( .INP(n9604), .ZN(n9550) );
  NAND3X0 U9311 ( .IN1(n9605), .IN2(n9482), .IN3(n9606), .QN(n9604) );
  NAND2X0 U9312 ( .IN1(n9466), .IN2(n4374), .QN(n9606) );
  NAND2X0 U9313 ( .IN1(n9607), .IN2(n4530), .QN(n9482) );
  NAND2X0 U9314 ( .IN1(n9464), .IN2(n9608), .QN(n9605) );
  XOR2X1 U9315 ( .IN1(n8627), .IN2(n9609), .Q(n9608) );
  NAND2X0 U9316 ( .IN1(n9610), .IN2(n9611), .QN(g30650) );
  NAND2X0 U9317 ( .IN1(test_so56), .IN2(n4515), .QN(n9611) );
  NAND2X0 U9318 ( .IN1(n9584), .IN2(g6782), .QN(n9610) );
  NAND2X0 U9319 ( .IN1(n9612), .IN2(n9613), .QN(g30649) );
  NAND2X0 U9320 ( .IN1(n4323), .IN2(g927), .QN(n9613) );
  NAND2X0 U9321 ( .IN1(n9553), .IN2(g6368), .QN(n9612) );
  INVX0 U9322 ( .INP(n9614), .ZN(n9553) );
  NAND3X0 U9323 ( .IN1(n9615), .IN2(n9514), .IN3(n9616), .QN(n9614) );
  NAND2X0 U9324 ( .IN1(n4391), .IN2(n9493), .QN(n9616) );
  NAND2X0 U9325 ( .IN1(n9495), .IN2(n9617), .QN(n9615) );
  XOR2X1 U9326 ( .IN1(n9618), .IN2(n9619), .Q(n9617) );
  NAND2X0 U9327 ( .IN1(n9620), .IN2(n9621), .QN(g30648) );
  NAND2X0 U9328 ( .IN1(n4312), .IN2(g921), .QN(n9621) );
  NAND2X0 U9329 ( .IN1(n9589), .IN2(g6518), .QN(n9620) );
  NAND2X0 U9330 ( .IN1(n9622), .IN2(n9623), .QN(g30647) );
  NAND2X0 U9331 ( .IN1(g915), .IN2(n8071), .QN(n9623) );
  NAND2X0 U9332 ( .IN1(test_so31), .IN2(n9624), .QN(n9622) );
  NAND2X0 U9333 ( .IN1(n9625), .IN2(n9626), .QN(g30646) );
  NAND2X0 U9334 ( .IN1(n4512), .IN2(g243), .QN(n9626) );
  NAND2X0 U9335 ( .IN1(n9592), .IN2(g6313), .QN(n9625) );
  NAND2X0 U9336 ( .IN1(n9627), .IN2(n9628), .QN(g30645) );
  NAND2X0 U9337 ( .IN1(n4369), .IN2(g237), .QN(n9628) );
  NAND2X0 U9338 ( .IN1(n9629), .IN2(g165), .QN(n9627) );
  NAND2X0 U9339 ( .IN1(n9630), .IN2(n9631), .QN(g30644) );
  NAND2X0 U9340 ( .IN1(n4317), .IN2(g1603), .QN(n9631) );
  NAND2X0 U9341 ( .IN1(n9584), .IN2(g6573), .QN(n9630) );
  NAND3X0 U9342 ( .IN1(n9632), .IN2(n9633), .IN3(n9462), .QN(n9584) );
  NAND2X0 U9343 ( .IN1(n9607), .IN2(n9634), .QN(n9462) );
  NAND2X0 U9344 ( .IN1(n9635), .IN2(n9464), .QN(n9633) );
  XOR2X1 U9345 ( .IN1(n2685), .IN2(n8639), .Q(n9635) );
  NAND2X0 U9346 ( .IN1(n9636), .IN2(n9637), .QN(n2685) );
  XOR2X1 U9347 ( .IN1(n9638), .IN2(n9188), .Q(n9637) );
  NAND2X0 U9348 ( .IN1(n9466), .IN2(n9639), .QN(n9632) );
  NAND2X0 U9349 ( .IN1(n9640), .IN2(n9641), .QN(g30643) );
  NAND2X0 U9350 ( .IN1(n4323), .IN2(g918), .QN(n9641) );
  NAND2X0 U9351 ( .IN1(n9589), .IN2(g6368), .QN(n9640) );
  INVX0 U9352 ( .INP(n9642), .ZN(n9589) );
  NAND3X0 U9353 ( .IN1(n9643), .IN2(n9514), .IN3(n9644), .QN(n9642) );
  NAND2X0 U9354 ( .IN1(n4375), .IN2(n9493), .QN(n9644) );
  NAND3X0 U9355 ( .IN1(n9645), .IN2(n9521), .IN3(n9646), .QN(n9514) );
  NAND2X0 U9356 ( .IN1(n9495), .IN2(n9647), .QN(n9643) );
  XOR2X1 U9357 ( .IN1(n9648), .IN2(n9649), .Q(n9647) );
  NAND2X0 U9358 ( .IN1(n9650), .IN2(n9651), .QN(g30642) );
  NAND2X0 U9359 ( .IN1(n4312), .IN2(g912), .QN(n9651) );
  NAND2X0 U9360 ( .IN1(n9624), .IN2(g6518), .QN(n9650) );
  NAND2X0 U9361 ( .IN1(n9652), .IN2(n9653), .QN(g30641) );
  NAND2X0 U9362 ( .IN1(n4318), .IN2(g240), .QN(n9653) );
  NAND2X0 U9363 ( .IN1(n9592), .IN2(g6231), .QN(n9652) );
  INVX0 U9364 ( .INP(n9654), .ZN(n9592) );
  NAND3X0 U9365 ( .IN1(n9655), .IN2(n9558), .IN3(n9656), .QN(n9654) );
  NAND2X0 U9366 ( .IN1(n4392), .IN2(n9529), .QN(n9656) );
  NAND2X0 U9367 ( .IN1(n9531), .IN2(n9657), .QN(n9655) );
  XOR2X1 U9368 ( .IN1(n8581), .IN2(n9658), .Q(n9657) );
  NAND2X0 U9369 ( .IN1(n9659), .IN2(n9660), .QN(g30640) );
  NAND2X0 U9370 ( .IN1(n4512), .IN2(g234), .QN(n9660) );
  NAND2X0 U9371 ( .IN1(n9629), .IN2(g6313), .QN(n9659) );
  NAND2X0 U9372 ( .IN1(n9661), .IN2(n9662), .QN(g30639) );
  NAND2X0 U9373 ( .IN1(n4369), .IN2(g228), .QN(n9662) );
  NAND2X0 U9374 ( .IN1(n9663), .IN2(g165), .QN(n9661) );
  NAND2X0 U9375 ( .IN1(n9664), .IN2(n9665), .QN(g30638) );
  NAND2X0 U9376 ( .IN1(n4323), .IN2(g909), .QN(n9665) );
  NAND2X0 U9377 ( .IN1(n9624), .IN2(g6368), .QN(n9664) );
  NAND3X0 U9378 ( .IN1(n9666), .IN2(n9491), .IN3(n9667), .QN(n9624) );
  NAND2X0 U9379 ( .IN1(n9493), .IN2(n9668), .QN(n9667) );
  NAND3X0 U9380 ( .IN1(n9645), .IN2(n9669), .IN3(n9646), .QN(n9491) );
  NAND2X0 U9381 ( .IN1(n9670), .IN2(n9495), .QN(n9666) );
  XNOR2X1 U9382 ( .IN1(n9520), .IN2(n8607), .Q(n9670) );
  NAND2X0 U9383 ( .IN1(n9671), .IN2(n9672), .QN(n9520) );
  XOR2X1 U9384 ( .IN1(n8610), .IN2(n9669), .Q(n9672) );
  NAND2X0 U9385 ( .IN1(n9673), .IN2(n9674), .QN(g30637) );
  NAND2X0 U9386 ( .IN1(n4318), .IN2(g231), .QN(n9674) );
  NAND2X0 U9387 ( .IN1(n9629), .IN2(g6231), .QN(n9673) );
  INVX0 U9388 ( .INP(n9675), .ZN(n9629) );
  NAND3X0 U9389 ( .IN1(n9676), .IN2(n9558), .IN3(n9677), .QN(n9675) );
  NAND2X0 U9390 ( .IN1(n4376), .IN2(n9529), .QN(n9677) );
  NAND3X0 U9391 ( .IN1(n9678), .IN2(n9679), .IN3(n9680), .QN(n9558) );
  NAND2X0 U9392 ( .IN1(n9531), .IN2(n9681), .QN(n9676) );
  XOR2X1 U9393 ( .IN1(n8570), .IN2(n9682), .Q(n9681) );
  NAND2X0 U9394 ( .IN1(n9683), .IN2(n9684), .QN(g30636) );
  NAND2X0 U9395 ( .IN1(n4512), .IN2(g225), .QN(n9684) );
  NAND2X0 U9396 ( .IN1(n9663), .IN2(g6313), .QN(n9683) );
  NAND2X0 U9397 ( .IN1(n9685), .IN2(n9686), .QN(g30635) );
  NAND2X0 U9398 ( .IN1(n4318), .IN2(g222), .QN(n9686) );
  NAND2X0 U9399 ( .IN1(n9663), .IN2(g6231), .QN(n9685) );
  NAND3X0 U9400 ( .IN1(n9687), .IN2(n9527), .IN3(n9688), .QN(n9663) );
  NAND2X0 U9401 ( .IN1(n9529), .IN2(n9689), .QN(n9688) );
  NAND3X0 U9402 ( .IN1(n9678), .IN2(n9186), .IN3(n9680), .QN(n9527) );
  NAND2X0 U9403 ( .IN1(n9690), .IN2(n9531), .QN(n9687) );
  XOR2X1 U9404 ( .IN1(n2718), .IN2(n9691), .Q(n9690) );
  NAND2X0 U9405 ( .IN1(n9692), .IN2(n9693), .QN(n2718) );
  XOR2X1 U9406 ( .IN1(n8565), .IN2(n9186), .Q(n9693) );
  NAND2X0 U9407 ( .IN1(n9694), .IN2(n9695), .QN(g30566) );
  NAND2X0 U9408 ( .IN1(n9332), .IN2(n4606), .QN(n9695) );
  INVX0 U9409 ( .INP(n9696), .ZN(n9332) );
  NAND2X0 U9410 ( .IN1(n9697), .IN2(n9698), .QN(n9696) );
  XOR2X1 U9411 ( .IN1(n9699), .IN2(n9700), .Q(n9697) );
  NAND2X0 U9412 ( .IN1(n9701), .IN2(n9702), .QN(n9700) );
  NAND2X0 U9413 ( .IN1(n9703), .IN2(n9704), .QN(n9702) );
  NAND4X0 U9414 ( .IN1(n9705), .IN2(n9706), .IN3(n9707), .IN4(n9708), .QN(
        n9701) );
  NAND3X0 U9415 ( .IN1(n9709), .IN2(n9710), .IN3(n9711), .QN(n9707) );
  NAND2X0 U9416 ( .IN1(n9712), .IN2(n9699), .QN(n9706) );
  INVX0 U9417 ( .INP(n9713), .ZN(n9712) );
  NAND2X0 U9418 ( .IN1(n9714), .IN2(n9715), .QN(n9705) );
  NAND2X0 U9419 ( .IN1(n9716), .IN2(n9717), .QN(n9714) );
  NAND2X0 U9420 ( .IN1(n9709), .IN2(n9718), .QN(n9717) );
  NAND3X0 U9421 ( .IN1(n9719), .IN2(n9710), .IN3(n9720), .QN(n9718) );
  INVX0 U9422 ( .INP(n9721), .ZN(n9720) );
  NAND2X0 U9423 ( .IN1(n9722), .IN2(n9713), .QN(n9719) );
  NAND2X0 U9424 ( .IN1(n9723), .IN2(n9724), .QN(n9716) );
  NAND2X0 U9425 ( .IN1(n9725), .IN2(n9726), .QN(n9723) );
  NAND2X0 U9426 ( .IN1(n4509), .IN2(g2392), .QN(n9694) );
  NAND2X0 U9427 ( .IN1(n9727), .IN2(n9728), .QN(g30505) );
  NAND2X0 U9428 ( .IN1(n9729), .IN2(g5555), .QN(n9728) );
  NAND2X0 U9429 ( .IN1(n4516), .IN2(g2393), .QN(n9727) );
  NAND2X0 U9430 ( .IN1(n9730), .IN2(n9731), .QN(g30503) );
  NAND2X0 U9431 ( .IN1(n9732), .IN2(g7014), .QN(n9731) );
  NAND2X0 U9432 ( .IN1(n4525), .IN2(g1700), .QN(n9730) );
  NAND2X0 U9433 ( .IN1(n9733), .IN2(n9734), .QN(g30500) );
  NAND2X0 U9434 ( .IN1(n2798), .IN2(g1088), .QN(n9734) );
  NAND2X0 U9435 ( .IN1(test_so39), .IN2(n4381), .QN(n9733) );
  NAND2X0 U9436 ( .IN1(n9735), .IN2(n9736), .QN(g30487) );
  NAND2X0 U9437 ( .IN1(n9732), .IN2(g5511), .QN(n9736) );
  NAND2X0 U9438 ( .IN1(n4518), .IN2(g1699), .QN(n9735) );
  NAND2X0 U9439 ( .IN1(n9737), .IN2(n9738), .QN(g30485) );
  NAND2X0 U9440 ( .IN1(n4364), .IN2(g1006), .QN(n9738) );
  NAND2X0 U9441 ( .IN1(n2798), .IN2(g6712), .QN(n9737) );
  NAND2X0 U9442 ( .IN1(n9739), .IN2(n9740), .QN(g30482) );
  NAND2X0 U9443 ( .IN1(n9741), .IN2(n4640), .QN(n9740) );
  NAND2X0 U9444 ( .IN1(n4506), .IN2(g320), .QN(n9739) );
  NAND2X0 U9445 ( .IN1(n9742), .IN2(n9743), .QN(g30470) );
  NAND2X0 U9446 ( .IN1(n4363), .IN2(g1005), .QN(n9743) );
  NAND2X0 U9447 ( .IN1(n2798), .IN2(g5472), .QN(n9742) );
  NAND2X0 U9448 ( .IN1(n9744), .IN2(n9745), .QN(g30468) );
  NAND2X0 U9449 ( .IN1(n9741), .IN2(g6447), .QN(n9745) );
  NAND2X0 U9450 ( .IN1(n4499), .IN2(g319), .QN(n9744) );
  NAND2X0 U9451 ( .IN1(n9746), .IN2(n9747), .QN(g30455) );
  NAND2X0 U9452 ( .IN1(n9741), .IN2(g5437), .QN(n9747) );
  INVX0 U9453 ( .INP(n9748), .ZN(n9741) );
  NAND2X0 U9454 ( .IN1(n9749), .IN2(n9388), .QN(n9748) );
  XOR2X1 U9455 ( .IN1(n9750), .IN2(n9399), .Q(n9749) );
  NAND2X0 U9456 ( .IN1(n9751), .IN2(n9752), .QN(n9750) );
  NAND2X0 U9457 ( .IN1(n9399), .IN2(n9753), .QN(n9752) );
  NAND3X0 U9458 ( .IN1(n9754), .IN2(n9755), .IN3(n9398), .QN(n9753) );
  NAND2X0 U9459 ( .IN1(n9411), .IN2(n9389), .QN(n9755) );
  NAND2X0 U9460 ( .IN1(n9416), .IN2(n9756), .QN(n9411) );
  NAND2X0 U9461 ( .IN1(n9757), .IN2(n3130), .QN(n9756) );
  INVX0 U9462 ( .INP(n9758), .ZN(n9757) );
  NAND3X0 U9463 ( .IN1(n9759), .IN2(g309), .IN3(n9405), .QN(n9754) );
  NAND3X0 U9464 ( .IN1(n9401), .IN2(n9398), .IN3(n9414), .QN(n9751) );
  INVX0 U9465 ( .INP(n9760), .ZN(n9401) );
  NAND3X0 U9466 ( .IN1(n9758), .IN2(n9389), .IN3(n3130), .QN(n9760) );
  NAND2X0 U9467 ( .IN1(n4520), .IN2(g318), .QN(n9746) );
  NAND2X0 U9468 ( .IN1(n9761), .IN2(n9762), .QN(g30356) );
  NAND2X0 U9469 ( .IN1(n9729), .IN2(n4606), .QN(n9762) );
  NAND2X0 U9470 ( .IN1(n4509), .IN2(g2395), .QN(n9761) );
  NAND2X0 U9471 ( .IN1(n9763), .IN2(n9764), .QN(g30341) );
  NAND2X0 U9472 ( .IN1(n9729), .IN2(g7264), .QN(n9764) );
  INVX0 U9473 ( .INP(n9765), .ZN(n9729) );
  NAND2X0 U9474 ( .IN1(n9766), .IN2(n9698), .QN(n9765) );
  XOR2X1 U9475 ( .IN1(n9767), .IN2(n9709), .Q(n9766) );
  NAND2X0 U9476 ( .IN1(n9768), .IN2(n9769), .QN(n9767) );
  NAND2X0 U9477 ( .IN1(n9709), .IN2(n9770), .QN(n9769) );
  NAND3X0 U9478 ( .IN1(n9771), .IN2(n9772), .IN3(n9708), .QN(n9770) );
  NAND2X0 U9479 ( .IN1(n9721), .IN2(n9699), .QN(n9772) );
  NAND2X0 U9480 ( .IN1(n9726), .IN2(n9773), .QN(n9721) );
  NAND2X0 U9481 ( .IN1(n9774), .IN2(n3038), .QN(n9773) );
  INVX0 U9482 ( .INP(n9775), .ZN(n9774) );
  NAND3X0 U9483 ( .IN1(test_so79), .IN2(n9776), .IN3(n9715), .QN(n9771) );
  NAND3X0 U9484 ( .IN1(n9711), .IN2(n9708), .IN3(n9724), .QN(n9768) );
  INVX0 U9485 ( .INP(n9777), .ZN(n9711) );
  NAND3X0 U9486 ( .IN1(n9775), .IN2(n9699), .IN3(n3038), .QN(n9777) );
  NAND2X0 U9487 ( .IN1(n4524), .IN2(g2394), .QN(n9763) );
  NAND2X0 U9488 ( .IN1(n9778), .IN2(n9779), .QN(g30338) );
  NAND2X0 U9489 ( .IN1(n9732), .IN2(n4618), .QN(n9779) );
  INVX0 U9490 ( .INP(n9780), .ZN(n9732) );
  NAND2X0 U9491 ( .IN1(n9781), .IN2(n9346), .QN(n9780) );
  XOR2X1 U9492 ( .IN1(n9782), .IN2(n9357), .Q(n9781) );
  NAND2X0 U9493 ( .IN1(n9783), .IN2(n9784), .QN(n9782) );
  NAND2X0 U9494 ( .IN1(n9357), .IN2(n9785), .QN(n9784) );
  NAND3X0 U9495 ( .IN1(n9786), .IN2(n9787), .IN3(n9356), .QN(n9785) );
  NAND2X0 U9496 ( .IN1(n9369), .IN2(n9347), .QN(n9787) );
  NAND2X0 U9497 ( .IN1(n9374), .IN2(n9788), .QN(n9369) );
  NAND2X0 U9498 ( .IN1(n9789), .IN2(n3070), .QN(n9788) );
  INVX0 U9499 ( .INP(n9790), .ZN(n9789) );
  NAND3X0 U9500 ( .IN1(n9791), .IN2(g1690), .IN3(n9363), .QN(n9786) );
  NAND3X0 U9501 ( .IN1(n9359), .IN2(n9356), .IN3(n9372), .QN(n9783) );
  INVX0 U9502 ( .INP(n9792), .ZN(n9359) );
  NAND3X0 U9503 ( .IN1(n9790), .IN2(n9347), .IN3(n3070), .QN(n9792) );
  NAND2X0 U9504 ( .IN1(n4511), .IN2(g1701), .QN(n9778) );
  NAND2X0 U9505 ( .IN1(n9793), .IN2(n9794), .QN(g30304) );
  NAND2X0 U9506 ( .IN1(n4367), .IN2(g2285), .QN(n9794) );
  NAND2X0 U9507 ( .IN1(n9795), .IN2(g2241), .QN(n9793) );
  NAND2X0 U9508 ( .IN1(n9796), .IN2(n9797), .QN(g30303) );
  NAND2X0 U9509 ( .IN1(g2282), .IN2(n8070), .QN(n9797) );
  NAND2X0 U9510 ( .IN1(test_so73), .IN2(n9795), .QN(n9796) );
  NAND2X0 U9511 ( .IN1(n9798), .IN2(n9799), .QN(g30302) );
  NAND2X0 U9512 ( .IN1(n4368), .IN2(g1591), .QN(n9799) );
  NAND2X0 U9513 ( .IN1(n9800), .IN2(g1547), .QN(n9798) );
  NAND2X0 U9514 ( .IN1(n9801), .IN2(n9802), .QN(g30301) );
  NAND2X0 U9515 ( .IN1(n4324), .IN2(g2279), .QN(n9802) );
  NAND2X0 U9516 ( .IN1(n9795), .IN2(g6837), .QN(n9801) );
  NAND2X0 U9517 ( .IN1(n9803), .IN2(n9804), .QN(n9795) );
  NAND2X0 U9518 ( .IN1(n9805), .IN2(n9436), .QN(n9804) );
  XOR2X1 U9519 ( .IN1(n9806), .IN2(n9807), .Q(n9805) );
  NAND2X0 U9520 ( .IN1(n9439), .IN2(g2185), .QN(n9803) );
  NAND2X0 U9521 ( .IN1(n9808), .IN2(n9809), .QN(g30300) );
  NAND2X0 U9522 ( .IN1(n4367), .IN2(g2267), .QN(n9809) );
  NAND2X0 U9523 ( .IN1(n9810), .IN2(g2241), .QN(n9808) );
  NAND2X0 U9524 ( .IN1(n9811), .IN2(n9812), .QN(g30299) );
  NAND2X0 U9525 ( .IN1(n4515), .IN2(g1588), .QN(n9812) );
  NAND2X0 U9526 ( .IN1(n9800), .IN2(g6782), .QN(n9811) );
  NAND2X0 U9527 ( .IN1(n9813), .IN2(n9814), .QN(g30298) );
  NAND2X0 U9528 ( .IN1(g897), .IN2(n8071), .QN(n9814) );
  NAND2X0 U9529 ( .IN1(test_so31), .IN2(n9815), .QN(n9813) );
  NAND2X0 U9530 ( .IN1(n9816), .IN2(n9817), .QN(g30297) );
  NAND2X0 U9531 ( .IN1(n4367), .IN2(g2339), .QN(n9817) );
  NAND2X0 U9532 ( .IN1(n9818), .IN2(g2241), .QN(n9816) );
  NAND2X0 U9533 ( .IN1(n9819), .IN2(n9820), .QN(g30296) );
  NAND2X0 U9534 ( .IN1(test_so76), .IN2(n8070), .QN(n9820) );
  NAND2X0 U9535 ( .IN1(test_so73), .IN2(n9810), .QN(n9819) );
  NAND2X0 U9536 ( .IN1(n9821), .IN2(n9822), .QN(g30295) );
  NAND2X0 U9537 ( .IN1(n4317), .IN2(g1585), .QN(n9822) );
  NAND2X0 U9538 ( .IN1(n9800), .IN2(g6573), .QN(n9821) );
  NAND2X0 U9539 ( .IN1(n9823), .IN2(n9824), .QN(n9800) );
  NAND2X0 U9540 ( .IN1(n9825), .IN2(n9464), .QN(n9824) );
  XNOR2X1 U9541 ( .IN1(n9826), .IN2(n8640), .Q(n9825) );
  NAND2X0 U9542 ( .IN1(n9466), .IN2(g1491), .QN(n9823) );
  NAND2X0 U9543 ( .IN1(n9827), .IN2(n9828), .QN(g30294) );
  NAND2X0 U9544 ( .IN1(n4368), .IN2(g1573), .QN(n9828) );
  NAND2X0 U9545 ( .IN1(n9829), .IN2(g1547), .QN(n9827) );
  NAND2X0 U9546 ( .IN1(n9830), .IN2(n9831), .QN(g30293) );
  NAND2X0 U9547 ( .IN1(n4312), .IN2(g894), .QN(n9831) );
  NAND2X0 U9548 ( .IN1(n9815), .IN2(g6518), .QN(n9830) );
  NAND2X0 U9549 ( .IN1(n9832), .IN2(n9833), .QN(g30292) );
  NAND2X0 U9550 ( .IN1(n4369), .IN2(g210), .QN(n9833) );
  NAND2X0 U9551 ( .IN1(n9834), .IN2(g165), .QN(n9832) );
  NAND2X0 U9552 ( .IN1(n9835), .IN2(n9836), .QN(g30291) );
  NAND2X0 U9553 ( .IN1(g2336), .IN2(n8070), .QN(n9836) );
  NAND2X0 U9554 ( .IN1(test_so73), .IN2(n9818), .QN(n9835) );
  NAND2X0 U9555 ( .IN1(n9837), .IN2(n9838), .QN(g30290) );
  NAND2X0 U9556 ( .IN1(n4367), .IN2(g2330), .QN(n9838) );
  NAND2X0 U9557 ( .IN1(n9839), .IN2(g2241), .QN(n9837) );
  NAND2X0 U9558 ( .IN1(n9840), .IN2(n9841), .QN(g30289) );
  NAND2X0 U9559 ( .IN1(n4324), .IN2(g2261), .QN(n9841) );
  NAND2X0 U9560 ( .IN1(n9810), .IN2(g6837), .QN(n9840) );
  NAND2X0 U9561 ( .IN1(n9842), .IN2(n9843), .QN(n9810) );
  NAND2X0 U9562 ( .IN1(n9436), .IN2(n9844), .QN(n9843) );
  XOR2X1 U9563 ( .IN1(n9845), .IN2(n9846), .Q(n9844) );
  NAND2X0 U9564 ( .IN1(n9439), .IN2(g2165), .QN(n9842) );
  NAND2X0 U9565 ( .IN1(n9847), .IN2(n9848), .QN(g30288) );
  NAND2X0 U9566 ( .IN1(n4368), .IN2(g1645), .QN(n9848) );
  NAND2X0 U9567 ( .IN1(n9849), .IN2(g1547), .QN(n9847) );
  NAND2X0 U9568 ( .IN1(n9850), .IN2(n9851), .QN(g30287) );
  NAND2X0 U9569 ( .IN1(n4515), .IN2(g1570), .QN(n9851) );
  NAND2X0 U9570 ( .IN1(n9829), .IN2(g6782), .QN(n9850) );
  NAND2X0 U9571 ( .IN1(n9852), .IN2(n9853), .QN(g30286) );
  NAND2X0 U9572 ( .IN1(n4323), .IN2(g891), .QN(n9853) );
  NAND2X0 U9573 ( .IN1(n9815), .IN2(g6368), .QN(n9852) );
  NAND2X0 U9574 ( .IN1(n9854), .IN2(n9855), .QN(n9815) );
  NAND2X0 U9575 ( .IN1(n9856), .IN2(n9495), .QN(n9855) );
  XNOR2X1 U9576 ( .IN1(n9857), .IN2(n8606), .Q(n9856) );
  INVX0 U9577 ( .INP(n9858), .ZN(n9854) );
  NOR2X0 U9578 ( .IN1(n9646), .IN2(n4327), .QN(n9858) );
  NAND2X0 U9579 ( .IN1(n9859), .IN2(n9860), .QN(g30285) );
  NAND2X0 U9580 ( .IN1(g879), .IN2(n8071), .QN(n9860) );
  NAND2X0 U9581 ( .IN1(test_so31), .IN2(n9861), .QN(n9859) );
  NAND2X0 U9582 ( .IN1(n9862), .IN2(n9863), .QN(g30284) );
  NAND2X0 U9583 ( .IN1(n4512), .IN2(g207), .QN(n9863) );
  NAND2X0 U9584 ( .IN1(n9834), .IN2(g6313), .QN(n9862) );
  NAND2X0 U9585 ( .IN1(n9864), .IN2(n9865), .QN(g30283) );
  NAND2X0 U9586 ( .IN1(n4324), .IN2(g2333), .QN(n9865) );
  NAND2X0 U9587 ( .IN1(n9818), .IN2(g6837), .QN(n9864) );
  NAND2X0 U9588 ( .IN1(n9866), .IN2(n9867), .QN(n9818) );
  NAND3X0 U9589 ( .IN1(n9436), .IN2(n9868), .IN3(n9869), .QN(n9867) );
  XOR2X1 U9590 ( .IN1(n8659), .IN2(n9599), .Q(n9869) );
  NOR2X0 U9591 ( .IN1(n9870), .IN2(n9871), .QN(n9599) );
  XOR2X1 U9592 ( .IN1(n9872), .IN2(n9189), .Q(n9871) );
  NAND2X0 U9593 ( .IN1(n9439), .IN2(g2200), .QN(n9866) );
  NAND2X0 U9594 ( .IN1(n9873), .IN2(n9874), .QN(g30282) );
  NAND2X0 U9595 ( .IN1(test_so77), .IN2(n8070), .QN(n9874) );
  NAND2X0 U9596 ( .IN1(test_so73), .IN2(n9839), .QN(n9873) );
  NAND2X0 U9597 ( .IN1(n9875), .IN2(n9876), .QN(g30281) );
  NAND2X0 U9598 ( .IN1(n4515), .IN2(g1642), .QN(n9876) );
  NAND2X0 U9599 ( .IN1(n9849), .IN2(g6782), .QN(n9875) );
  NAND2X0 U9600 ( .IN1(n9877), .IN2(n9878), .QN(g30280) );
  NAND2X0 U9601 ( .IN1(n4368), .IN2(g1636), .QN(n9878) );
  NAND2X0 U9602 ( .IN1(n9879), .IN2(g1547), .QN(n9877) );
  NAND2X0 U9603 ( .IN1(n9880), .IN2(n9881), .QN(g30279) );
  NAND2X0 U9604 ( .IN1(n4317), .IN2(g1567), .QN(n9881) );
  NAND2X0 U9605 ( .IN1(n9829), .IN2(g6573), .QN(n9880) );
  NAND2X0 U9606 ( .IN1(n9882), .IN2(n9883), .QN(n9829) );
  NAND2X0 U9607 ( .IN1(n9464), .IN2(n9884), .QN(n9883) );
  XOR2X1 U9608 ( .IN1(n8638), .IN2(n9885), .Q(n9884) );
  NAND2X0 U9609 ( .IN1(n9466), .IN2(g1471), .QN(n9882) );
  NAND2X0 U9610 ( .IN1(n9886), .IN2(n9887), .QN(g30278) );
  NAND2X0 U9611 ( .IN1(g951), .IN2(n8071), .QN(n9887) );
  NAND2X0 U9612 ( .IN1(test_so31), .IN2(n9888), .QN(n9886) );
  NAND2X0 U9613 ( .IN1(n9889), .IN2(n9890), .QN(g30277) );
  NAND2X0 U9614 ( .IN1(n4312), .IN2(g876), .QN(n9890) );
  NAND2X0 U9615 ( .IN1(n9861), .IN2(g6518), .QN(n9889) );
  NAND2X0 U9616 ( .IN1(n9891), .IN2(n9892), .QN(g30276) );
  NAND2X0 U9617 ( .IN1(n4318), .IN2(g204), .QN(n9892) );
  NAND2X0 U9618 ( .IN1(n9834), .IN2(g6231), .QN(n9891) );
  NAND2X0 U9619 ( .IN1(n9893), .IN2(n9894), .QN(n9834) );
  NAND2X0 U9620 ( .IN1(n9895), .IN2(n9531), .QN(n9894) );
  XNOR2X1 U9621 ( .IN1(n9896), .IN2(n8575), .Q(n9895) );
  NAND2X0 U9622 ( .IN1(n9529), .IN2(g113), .QN(n9893) );
  NAND2X0 U9623 ( .IN1(n9897), .IN2(n9898), .QN(g30275) );
  NAND2X0 U9624 ( .IN1(n4369), .IN2(g192), .QN(n9898) );
  NAND2X0 U9625 ( .IN1(n9899), .IN2(g165), .QN(n9897) );
  NAND2X0 U9626 ( .IN1(n9900), .IN2(n9901), .QN(g30274) );
  NAND2X0 U9627 ( .IN1(n4324), .IN2(g2324), .QN(n9901) );
  NAND2X0 U9628 ( .IN1(n9839), .IN2(g6837), .QN(n9900) );
  NAND2X0 U9629 ( .IN1(n9902), .IN2(n9903), .QN(n9839) );
  NAND3X0 U9630 ( .IN1(n9436), .IN2(n9868), .IN3(n9904), .QN(n9903) );
  XOR2X1 U9631 ( .IN1(n8653), .IN2(n9905), .Q(n9904) );
  INVX0 U9632 ( .INP(n9567), .ZN(n9868) );
  NAND2X0 U9633 ( .IN1(n9439), .IN2(g2190), .QN(n9902) );
  NAND2X0 U9634 ( .IN1(n9906), .IN2(n9907), .QN(g30273) );
  NAND2X0 U9635 ( .IN1(n4317), .IN2(g1639), .QN(n9907) );
  NAND2X0 U9636 ( .IN1(n9849), .IN2(g6573), .QN(n9906) );
  NAND2X0 U9637 ( .IN1(n9908), .IN2(n9909), .QN(n9849) );
  NAND3X0 U9638 ( .IN1(n9464), .IN2(n9910), .IN3(n9911), .QN(n9909) );
  XOR2X1 U9639 ( .IN1(n9638), .IN2(n9636), .Q(n9911) );
  NOR2X0 U9640 ( .IN1(n9912), .IN2(n9913), .QN(n9636) );
  XOR2X1 U9641 ( .IN1(n8625), .IN2(n9188), .Q(n9913) );
  NAND2X0 U9642 ( .IN1(n9466), .IN2(g1506), .QN(n9908) );
  NAND2X0 U9643 ( .IN1(n9914), .IN2(n9915), .QN(g30272) );
  NAND2X0 U9644 ( .IN1(n4515), .IN2(g1633), .QN(n9915) );
  NAND2X0 U9645 ( .IN1(n9879), .IN2(g6782), .QN(n9914) );
  NAND2X0 U9646 ( .IN1(n9916), .IN2(n9917), .QN(g30271) );
  NAND2X0 U9647 ( .IN1(n4312), .IN2(g948), .QN(n9917) );
  NAND2X0 U9648 ( .IN1(n9888), .IN2(g6518), .QN(n9916) );
  NAND2X0 U9649 ( .IN1(n9918), .IN2(n9919), .QN(g30270) );
  NAND2X0 U9650 ( .IN1(g942), .IN2(n8071), .QN(n9919) );
  NAND2X0 U9651 ( .IN1(test_so31), .IN2(n9920), .QN(n9918) );
  NAND2X0 U9652 ( .IN1(n9921), .IN2(n9922), .QN(g30269) );
  NAND2X0 U9653 ( .IN1(n4323), .IN2(g873), .QN(n9922) );
  NAND2X0 U9654 ( .IN1(n9861), .IN2(g6368), .QN(n9921) );
  NAND2X0 U9655 ( .IN1(n9923), .IN2(n9924), .QN(n9861) );
  NAND2X0 U9656 ( .IN1(n9495), .IN2(n9925), .QN(n9924) );
  XOR2X1 U9657 ( .IN1(n9926), .IN2(n9927), .Q(n9925) );
  INVX0 U9658 ( .INP(n9928), .ZN(n9923) );
  NOR2X0 U9659 ( .IN1(n9646), .IN2(n4379), .QN(n9928) );
  NAND2X0 U9660 ( .IN1(n9929), .IN2(n9930), .QN(g30268) );
  NAND2X0 U9661 ( .IN1(n4369), .IN2(g264), .QN(n9930) );
  NAND2X0 U9662 ( .IN1(n9931), .IN2(g165), .QN(n9929) );
  NAND2X0 U9663 ( .IN1(n9932), .IN2(n9933), .QN(g30267) );
  NAND2X0 U9664 ( .IN1(test_so13), .IN2(n4512), .QN(n9933) );
  NAND2X0 U9665 ( .IN1(n9899), .IN2(g6313), .QN(n9932) );
  NAND2X0 U9666 ( .IN1(n9934), .IN2(n9935), .QN(g30266) );
  NAND2X0 U9667 ( .IN1(n4317), .IN2(g1630), .QN(n9935) );
  NAND2X0 U9668 ( .IN1(n9879), .IN2(g6573), .QN(n9934) );
  NAND2X0 U9669 ( .IN1(n9936), .IN2(n9937), .QN(n9879) );
  NAND3X0 U9670 ( .IN1(n9464), .IN2(n9910), .IN3(n9938), .QN(n9937) );
  XOR2X1 U9671 ( .IN1(n8629), .IN2(n9939), .Q(n9938) );
  INVX0 U9672 ( .INP(n9607), .ZN(n9910) );
  NAND2X0 U9673 ( .IN1(n9466), .IN2(g1496), .QN(n9936) );
  NAND2X0 U9674 ( .IN1(n9940), .IN2(n9941), .QN(g30265) );
  NAND2X0 U9675 ( .IN1(test_so35), .IN2(n4323), .QN(n9941) );
  NAND2X0 U9676 ( .IN1(n9888), .IN2(g6368), .QN(n9940) );
  NAND2X0 U9677 ( .IN1(n9942), .IN2(n9943), .QN(n9888) );
  NAND2X0 U9678 ( .IN1(n9944), .IN2(n9495), .QN(n9943) );
  XOR2X1 U9679 ( .IN1(n8610), .IN2(n9671), .Q(n9944) );
  NOR2X0 U9680 ( .IN1(n9945), .IN2(n9946), .QN(n9671) );
  XOR2X1 U9681 ( .IN1(n9947), .IN2(n9669), .Q(n9946) );
  NAND2X0 U9682 ( .IN1(n9493), .IN2(g813), .QN(n9942) );
  NAND2X0 U9683 ( .IN1(n9948), .IN2(n9949), .QN(g30264) );
  NAND2X0 U9684 ( .IN1(n4312), .IN2(g939), .QN(n9949) );
  NAND2X0 U9685 ( .IN1(n9920), .IN2(g6518), .QN(n9948) );
  NAND2X0 U9686 ( .IN1(n9950), .IN2(n9951), .QN(g30263) );
  NAND2X0 U9687 ( .IN1(n4512), .IN2(g261), .QN(n9951) );
  NAND2X0 U9688 ( .IN1(n9931), .IN2(g6313), .QN(n9950) );
  NAND2X0 U9689 ( .IN1(n9952), .IN2(n9953), .QN(g30262) );
  NAND2X0 U9690 ( .IN1(n4369), .IN2(test_so14), .QN(n9953) );
  NAND2X0 U9691 ( .IN1(n9954), .IN2(g165), .QN(n9952) );
  NAND2X0 U9692 ( .IN1(n9955), .IN2(n9956), .QN(g30261) );
  NAND2X0 U9693 ( .IN1(n4318), .IN2(g186), .QN(n9956) );
  NAND2X0 U9694 ( .IN1(n9899), .IN2(g6231), .QN(n9955) );
  NAND2X0 U9695 ( .IN1(n9957), .IN2(n9958), .QN(n9899) );
  NAND2X0 U9696 ( .IN1(n9531), .IN2(n9959), .QN(n9958) );
  XOR2X1 U9697 ( .IN1(n4513), .IN2(n9960), .Q(n9959) );
  NAND2X0 U9698 ( .IN1(n9529), .IN2(g97), .QN(n9957) );
  NAND2X0 U9699 ( .IN1(n9961), .IN2(n9962), .QN(g30260) );
  NAND2X0 U9700 ( .IN1(n4367), .IN2(g2294), .QN(n9962) );
  NAND2X0 U9701 ( .IN1(n9963), .IN2(g2241), .QN(n9961) );
  NAND2X0 U9702 ( .IN1(n9964), .IN2(n9965), .QN(g30259) );
  NAND2X0 U9703 ( .IN1(n4323), .IN2(g936), .QN(n9965) );
  NAND2X0 U9704 ( .IN1(n9920), .IN2(g6368), .QN(n9964) );
  NAND2X0 U9705 ( .IN1(n9966), .IN2(n9967), .QN(n9920) );
  NAND2X0 U9706 ( .IN1(n9968), .IN2(n9495), .QN(n9967) );
  XOR2X1 U9707 ( .IN1(n8601), .IN2(n9969), .Q(n9968) );
  NAND2X0 U9708 ( .IN1(n9493), .IN2(g805), .QN(n9966) );
  NAND2X0 U9709 ( .IN1(n9970), .IN2(n9971), .QN(g30258) );
  NAND2X0 U9710 ( .IN1(n4318), .IN2(g258), .QN(n9971) );
  NAND2X0 U9711 ( .IN1(n9931), .IN2(g6231), .QN(n9970) );
  NAND2X0 U9712 ( .IN1(n9972), .IN2(n9973), .QN(n9931) );
  NAND2X0 U9713 ( .IN1(n9974), .IN2(n9531), .QN(n9973) );
  XOR2X1 U9714 ( .IN1(n8565), .IN2(n9692), .Q(n9974) );
  NOR2X0 U9715 ( .IN1(n9975), .IN2(n9976), .QN(n9692) );
  XOR2X1 U9716 ( .IN1(n8569), .IN2(n9679), .Q(n9976) );
  NAND2X0 U9717 ( .IN1(n9529), .IN2(g125), .QN(n9972) );
  NAND2X0 U9718 ( .IN1(n9977), .IN2(n9978), .QN(g30257) );
  NAND2X0 U9719 ( .IN1(n4512), .IN2(g252), .QN(n9978) );
  NAND2X0 U9720 ( .IN1(n9954), .IN2(g6313), .QN(n9977) );
  NAND2X0 U9721 ( .IN1(n9979), .IN2(n9980), .QN(g30256) );
  NAND2X0 U9722 ( .IN1(g2291), .IN2(n8070), .QN(n9980) );
  NAND2X0 U9723 ( .IN1(test_so73), .IN2(n9963), .QN(n9979) );
  NAND2X0 U9724 ( .IN1(n9981), .IN2(n9982), .QN(g30255) );
  NAND2X0 U9725 ( .IN1(n4368), .IN2(g1600), .QN(n9982) );
  NAND2X0 U9726 ( .IN1(n9983), .IN2(g1547), .QN(n9981) );
  NAND2X0 U9727 ( .IN1(n9984), .IN2(n9985), .QN(g30254) );
  NAND2X0 U9728 ( .IN1(n4318), .IN2(g249), .QN(n9985) );
  NAND2X0 U9729 ( .IN1(n9954), .IN2(g6231), .QN(n9984) );
  NAND2X0 U9730 ( .IN1(n9986), .IN2(n9987), .QN(n9954) );
  NAND2X0 U9731 ( .IN1(n9988), .IN2(n9531), .QN(n9987) );
  XOR2X1 U9732 ( .IN1(n8564), .IN2(n9989), .Q(n9988) );
  NAND2X0 U9733 ( .IN1(n9529), .IN2(g117), .QN(n9986) );
  NAND2X0 U9734 ( .IN1(n9990), .IN2(n9991), .QN(g30253) );
  NAND2X0 U9735 ( .IN1(n4324), .IN2(g2288), .QN(n9991) );
  NAND2X0 U9736 ( .IN1(n9963), .IN2(g6837), .QN(n9990) );
  NAND2X0 U9737 ( .IN1(n9992), .IN2(n9993), .QN(n9963) );
  NAND2X0 U9738 ( .IN1(n9994), .IN2(n9436), .QN(n9993) );
  XOR2X1 U9739 ( .IN1(n9870), .IN2(n9872), .Q(n9994) );
  NAND2X0 U9740 ( .IN1(n9905), .IN2(n9995), .QN(n9870) );
  XOR2X1 U9741 ( .IN1(n8653), .IN2(n9189), .Q(n9995) );
  NOR2X0 U9742 ( .IN1(n9806), .IN2(n9996), .QN(n9905) );
  XOR2X1 U9743 ( .IN1(n9807), .IN2(n9189), .Q(n9996) );
  INVX0 U9744 ( .INP(n8666), .ZN(n9807) );
  NAND2X0 U9745 ( .IN1(n9539), .IN2(n9997), .QN(n9806) );
  XOR2X1 U9746 ( .IN1(n8652), .IN2(n9189), .Q(n9997) );
  NOR2X0 U9747 ( .IN1(n9437), .IN2(n9998), .QN(n9539) );
  XOR2X1 U9748 ( .IN1(n9438), .IN2(n9189), .Q(n9998) );
  NAND2X0 U9749 ( .IN1(n9569), .IN2(n9999), .QN(n9437) );
  XOR2X1 U9750 ( .IN1(n9570), .IN2(n9189), .Q(n9999) );
  NOR2X0 U9751 ( .IN1(n10000), .IN2(n9846), .QN(n9569) );
  XOR2X1 U9752 ( .IN1(n9845), .IN2(n9189), .Q(n10000) );
  NAND2X0 U9753 ( .IN1(n9439), .IN2(g2195), .QN(n9992) );
  NOR2X0 U9754 ( .IN1(n9567), .IN2(n9436), .QN(n9439) );
  NOR2X0 U9755 ( .IN1(n10001), .IN2(n10002), .QN(n9436) );
  NOR2X0 U9756 ( .IN1(n10003), .IN2(n10004), .QN(n10002) );
  NOR2X0 U9757 ( .IN1(n9597), .IN2(n10005), .QN(n10004) );
  NOR2X0 U9758 ( .IN1(n10001), .IN2(n10003), .QN(n9567) );
  NAND2X0 U9759 ( .IN1(n10006), .IN2(n10007), .QN(n10003) );
  NAND2X0 U9760 ( .IN1(n10008), .IN2(n8643), .QN(n10007) );
  NAND4X0 U9761 ( .IN1(n9540), .IN2(n10009), .IN3(n10010), .IN4(n10011), .QN(
        n8643) );
  NOR3X0 U9762 ( .IN1(n8664), .IN2(n9570), .IN3(n8665), .QN(n10011) );
  INVX0 U9763 ( .INP(n10012), .ZN(n10010) );
  INVX0 U9764 ( .INP(n8654), .ZN(n10009) );
  INVX0 U9765 ( .INP(n8652), .ZN(n9540) );
  INVX0 U9766 ( .INP(n10005), .ZN(n10008) );
  NOR4X0 U9767 ( .IN1(n10012), .IN2(n9438), .IN3(n9597), .IN4(n10013), .QN(
        n10005) );
  NAND4X0 U9768 ( .IN1(n8652), .IN2(n8654), .IN3(n9570), .IN4(n8665), .QN(
        n10013) );
  INVX0 U9769 ( .INP(n4529), .ZN(n9597) );
  INVX0 U9770 ( .INP(n8664), .ZN(n9438) );
  NAND4X0 U9771 ( .IN1(n10014), .IN2(n9872), .IN3(n10015), .IN4(n9845), .QN(
        n10012) );
  INVX0 U9772 ( .INP(n8660), .ZN(n9845) );
  NOR2X0 U9773 ( .IN1(n8666), .IN2(n8659), .QN(n10015) );
  INVX0 U9774 ( .INP(n8658), .ZN(n9872) );
  INVX0 U9775 ( .INP(n8653), .ZN(n10014) );
  INVX0 U9776 ( .INP(n9846), .ZN(n10006) );
  NOR2X0 U9777 ( .IN1(n10016), .IN2(n4529), .QN(n9846) );
  INVX0 U9778 ( .INP(n9189), .ZN(n4529) );
  NAND3X0 U9779 ( .IN1(n10017), .IN2(n9698), .IN3(n10018), .QN(n10001) );
  NAND2X0 U9780 ( .IN1(n10019), .IN2(n9722), .QN(n10018) );
  NAND2X0 U9781 ( .IN1(n10020), .IN2(n9708), .QN(n10017) );
  NAND2X0 U9782 ( .IN1(n9726), .IN2(n10021), .QN(n10020) );
  NAND3X0 U9783 ( .IN1(n9722), .IN2(n9715), .IN3(n9776), .QN(n10021) );
  INVX0 U9784 ( .INP(n9725), .ZN(n9722) );
  NAND2X0 U9785 ( .IN1(n10022), .IN2(n10023), .QN(n9725) );
  NAND3X0 U9786 ( .IN1(n10024), .IN2(n10025), .IN3(n10026), .QN(n10023) );
  NAND2X0 U9787 ( .IN1(n7310), .IN2(n10027), .QN(n10026) );
  NAND2X0 U9788 ( .IN1(n7313), .IN2(n10028), .QN(n10025) );
  NAND2X0 U9789 ( .IN1(n7314), .IN2(n10029), .QN(n10024) );
  NAND2X0 U9790 ( .IN1(n10030), .IN2(n10031), .QN(g30252) );
  NAND2X0 U9791 ( .IN1(n4515), .IN2(g1597), .QN(n10031) );
  NAND2X0 U9792 ( .IN1(n9983), .IN2(g6782), .QN(n10030) );
  NAND2X0 U9793 ( .IN1(n10032), .IN2(n10033), .QN(g30251) );
  NAND2X0 U9794 ( .IN1(g906), .IN2(n8071), .QN(n10033) );
  NAND2X0 U9795 ( .IN1(test_so31), .IN2(n10034), .QN(n10032) );
  NAND2X0 U9796 ( .IN1(n10035), .IN2(n10036), .QN(g30250) );
  NAND2X0 U9797 ( .IN1(n4317), .IN2(g1594), .QN(n10036) );
  NAND2X0 U9798 ( .IN1(n9983), .IN2(g6573), .QN(n10035) );
  NAND2X0 U9799 ( .IN1(n10037), .IN2(n10038), .QN(n9983) );
  NAND2X0 U9800 ( .IN1(n10039), .IN2(n9464), .QN(n10038) );
  XOR2X1 U9801 ( .IN1(n9912), .IN2(n8625), .Q(n10039) );
  NAND2X0 U9802 ( .IN1(n9939), .IN2(n10040), .QN(n9912) );
  XOR2X1 U9803 ( .IN1(n8629), .IN2(n9188), .Q(n10040) );
  NOR2X0 U9804 ( .IN1(n9826), .IN2(n10041), .QN(n9939) );
  XNOR2X1 U9805 ( .IN1(n8640), .IN2(n9188), .Q(n10041) );
  NAND2X0 U9806 ( .IN1(n9579), .IN2(n10042), .QN(n9826) );
  XOR2X1 U9807 ( .IN1(n10043), .IN2(n9188), .Q(n10042) );
  NOR2X0 U9808 ( .IN1(n9465), .IN2(n10044), .QN(n9579) );
  XOR2X1 U9809 ( .IN1(n8637), .IN2(n4530), .Q(n10044) );
  NAND2X0 U9810 ( .IN1(n9609), .IN2(n10045), .QN(n9465) );
  XOR2X1 U9811 ( .IN1(n10046), .IN2(n9188), .Q(n10045) );
  NOR2X0 U9812 ( .IN1(n10047), .IN2(n10048), .QN(n9609) );
  XOR2X1 U9813 ( .IN1(n8638), .IN2(n4530), .Q(n10047) );
  NAND2X0 U9814 ( .IN1(n9466), .IN2(g1501), .QN(n10037) );
  NOR2X0 U9815 ( .IN1(n9607), .IN2(n9464), .QN(n9466) );
  NOR2X0 U9816 ( .IN1(n10049), .IN2(n10050), .QN(n9464) );
  NOR2X0 U9817 ( .IN1(n10051), .IN2(n10052), .QN(n10050) );
  NOR2X0 U9818 ( .IN1(n9634), .IN2(n10053), .QN(n10052) );
  INVX0 U9819 ( .INP(n10054), .ZN(n10053) );
  INVX0 U9820 ( .INP(n4530), .ZN(n9634) );
  NOR2X0 U9821 ( .IN1(n10049), .IN2(n10051), .QN(n9607) );
  NAND2X0 U9822 ( .IN1(n9885), .IN2(n10055), .QN(n10051) );
  NAND2X0 U9823 ( .IN1(n10054), .IN2(n8613), .QN(n10055) );
  NAND4X0 U9824 ( .IN1(n8628), .IN2(n10056), .IN3(n10057), .IN4(n10058), .QN(
        n8613) );
  NOR3X0 U9825 ( .IN1(n10046), .IN2(n8637), .IN3(n9187), .QN(n10058) );
  NAND4X0 U9826 ( .IN1(n10057), .IN2(n8637), .IN3(n4530), .IN4(n10059), .QN(
        n10054) );
  NOR4X0 U9827 ( .IN1(n8628), .IN2(n10056), .IN3(n8627), .IN4(n8639), .QN(
        n10059) );
  INVX0 U9828 ( .INP(n10043), .ZN(n8628) );
  INVX0 U9829 ( .INP(n10060), .ZN(n10057) );
  NAND4X0 U9830 ( .IN1(n10061), .IN2(n8625), .IN3(n10062), .IN4(n8626), .QN(
        n10060) );
  NOR2X0 U9831 ( .IN1(n8640), .IN2(n8638), .QN(n10062) );
  INVX0 U9832 ( .INP(n10063), .ZN(n8625) );
  INVX0 U9833 ( .INP(n10048), .ZN(n9885) );
  NOR2X0 U9834 ( .IN1(n8615), .IN2(n4530), .QN(n10048) );
  INVX0 U9835 ( .INP(n9188), .ZN(n4530) );
  NAND3X0 U9836 ( .IN1(n10064), .IN2(n9346), .IN3(n10065), .QN(n10049) );
  NAND2X0 U9837 ( .IN1(n10066), .IN2(n9370), .QN(n10065) );
  NAND2X0 U9838 ( .IN1(n10067), .IN2(n9356), .QN(n10064) );
  NAND2X0 U9839 ( .IN1(n9374), .IN2(n10068), .QN(n10067) );
  NAND3X0 U9840 ( .IN1(n9370), .IN2(n9363), .IN3(n9791), .QN(n10068) );
  INVX0 U9841 ( .INP(n9373), .ZN(n9370) );
  NAND2X0 U9842 ( .IN1(n10069), .IN2(n10070), .QN(n9373) );
  NAND3X0 U9843 ( .IN1(n10071), .IN2(n10072), .IN3(n10073), .QN(n10070) );
  NAND2X0 U9844 ( .IN1(n7311), .IN2(n10074), .QN(n10073) );
  NAND2X0 U9845 ( .IN1(n7315), .IN2(n10075), .QN(n10072) );
  NAND2X0 U9846 ( .IN1(n7316), .IN2(n10076), .QN(n10071) );
  NAND2X0 U9847 ( .IN1(n10077), .IN2(n10078), .QN(g30249) );
  NAND2X0 U9848 ( .IN1(n4312), .IN2(g903), .QN(n10078) );
  NAND2X0 U9849 ( .IN1(n10034), .IN2(g6518), .QN(n10077) );
  NAND2X0 U9850 ( .IN1(n10079), .IN2(n10080), .QN(g30248) );
  NAND2X0 U9851 ( .IN1(n4369), .IN2(g219), .QN(n10080) );
  NAND2X0 U9852 ( .IN1(n10081), .IN2(g165), .QN(n10079) );
  NAND2X0 U9853 ( .IN1(n10082), .IN2(n10083), .QN(g30247) );
  NAND2X0 U9854 ( .IN1(n4323), .IN2(g900), .QN(n10083) );
  NAND2X0 U9855 ( .IN1(n10034), .IN2(g6368), .QN(n10082) );
  NAND2X0 U9856 ( .IN1(n10084), .IN2(n10085), .QN(n10034) );
  NAND2X0 U9857 ( .IN1(n10086), .IN2(n9495), .QN(n10085) );
  INVX0 U9858 ( .INP(n10087), .ZN(n9495) );
  NAND2X0 U9859 ( .IN1(n9646), .IN2(n10088), .QN(n10087) );
  NAND2X0 U9860 ( .IN1(n9645), .IN2(n10089), .QN(n10088) );
  NAND2X0 U9861 ( .IN1(n9521), .IN2(n10090), .QN(n10089) );
  NOR2X0 U9862 ( .IN1(n9927), .IN2(n10091), .QN(n9645) );
  INVX0 U9863 ( .INP(n10092), .ZN(n10091) );
  NAND2X0 U9864 ( .IN1(n10090), .IN2(n8584), .QN(n10092) );
  NAND4X0 U9865 ( .IN1(n9648), .IN2(n9618), .IN3(n10093), .IN4(n10094), .QN(
        n8584) );
  NOR3X0 U9866 ( .IN1(n8599), .IN2(n8607), .IN3(n8605), .QN(n10094) );
  INVX0 U9867 ( .INP(n8595), .ZN(n9618) );
  INVX0 U9868 ( .INP(n8593), .ZN(n9648) );
  NAND4X0 U9869 ( .IN1(n10093), .IN2(n8607), .IN3(n9521), .IN4(n10095), .QN(
        n10090) );
  INVX0 U9870 ( .INP(n10096), .ZN(n10095) );
  NAND4X0 U9871 ( .IN1(n8593), .IN2(n8595), .IN3(n8599), .IN4(n8605), .QN(
        n10096) );
  INVX0 U9872 ( .INP(n10097), .ZN(n10093) );
  NAND4X0 U9873 ( .IN1(n9947), .IN2(n10098), .IN3(n10099), .IN4(n9926), .QN(
        n10097) );
  NOR2X0 U9874 ( .IN1(n8610), .IN2(n8606), .QN(n10099) );
  INVX0 U9875 ( .INP(n8601), .ZN(n10098) );
  INVX0 U9876 ( .INP(n9493), .ZN(n9646) );
  XOR2X1 U9877 ( .IN1(n9945), .IN2(n9947), .Q(n10086) );
  INVX0 U9878 ( .INP(n8594), .ZN(n9947) );
  NAND2X0 U9879 ( .IN1(n9969), .IN2(n10100), .QN(n9945) );
  XOR2X1 U9880 ( .IN1(n8601), .IN2(n9669), .Q(n10100) );
  NOR2X0 U9881 ( .IN1(n9857), .IN2(n10101), .QN(n9969) );
  XNOR2X1 U9882 ( .IN1(n8606), .IN2(n9669), .Q(n10101) );
  NAND2X0 U9883 ( .IN1(n9619), .IN2(n10102), .QN(n9857) );
  XOR2X1 U9884 ( .IN1(n8595), .IN2(n9669), .Q(n10102) );
  NOR2X0 U9885 ( .IN1(n9496), .IN2(n10103), .QN(n9619) );
  XOR2X1 U9886 ( .IN1(n8599), .IN2(n9521), .Q(n10103) );
  NAND2X0 U9887 ( .IN1(n9649), .IN2(n10104), .QN(n9496) );
  XOR2X1 U9888 ( .IN1(n8593), .IN2(n9669), .Q(n10104) );
  NOR2X0 U9889 ( .IN1(n10105), .IN2(n9927), .QN(n9649) );
  NOR2X0 U9890 ( .IN1(n10106), .IN2(n9521), .QN(n9927) );
  XOR2X1 U9891 ( .IN1(n9926), .IN2(n9669), .Q(n10105) );
  INVX0 U9892 ( .INP(n8600), .ZN(n9926) );
  NAND2X0 U9893 ( .IN1(n9493), .IN2(g809), .QN(n10084) );
  NAND3X0 U9894 ( .IN1(n10107), .IN2(n10108), .IN3(n10109), .QN(n9493) );
  NAND2X0 U9895 ( .IN1(n10110), .IN2(n9211), .QN(n10109) );
  NAND2X0 U9896 ( .IN1(n10111), .IN2(n9179), .QN(n10107) );
  NAND2X0 U9897 ( .IN1(n9208), .IN2(n10112), .QN(n10111) );
  NAND3X0 U9898 ( .IN1(n9182), .IN2(n9183), .IN3(n9211), .QN(n10112) );
  INVX0 U9899 ( .INP(n9214), .ZN(n9211) );
  NAND2X0 U9900 ( .IN1(n10113), .IN2(n10114), .QN(n9214) );
  NAND3X0 U9901 ( .IN1(n10115), .IN2(n10116), .IN3(n10117), .QN(n10114) );
  NAND2X0 U9902 ( .IN1(n7317), .IN2(g1088), .QN(n10117) );
  NAND2X0 U9903 ( .IN1(n7318), .IN2(g5472), .QN(n10116) );
  NAND2X0 U9904 ( .IN1(n7312), .IN2(g6712), .QN(n10115) );
  NAND2X0 U9905 ( .IN1(n10118), .IN2(n10119), .QN(g30246) );
  NAND2X0 U9906 ( .IN1(n4512), .IN2(g216), .QN(n10119) );
  NAND2X0 U9907 ( .IN1(n10081), .IN2(g6313), .QN(n10118) );
  NAND2X0 U9908 ( .IN1(n10120), .IN2(n10121), .QN(g30245) );
  NAND2X0 U9909 ( .IN1(n4318), .IN2(g213), .QN(n10121) );
  NAND2X0 U9910 ( .IN1(n10081), .IN2(g6231), .QN(n10120) );
  NAND2X0 U9911 ( .IN1(n10122), .IN2(n10123), .QN(n10081) );
  NAND2X0 U9912 ( .IN1(n10124), .IN2(n9531), .QN(n10123) );
  INVX0 U9913 ( .INP(n10125), .ZN(n9531) );
  NAND2X0 U9914 ( .IN1(n9680), .IN2(n10126), .QN(n10125) );
  NAND2X0 U9915 ( .IN1(n9678), .IN2(n10127), .QN(n10126) );
  NAND2X0 U9916 ( .IN1(n9679), .IN2(n10128), .QN(n10127) );
  NOR2X0 U9917 ( .IN1(n9960), .IN2(n10129), .QN(n9678) );
  INVX0 U9918 ( .INP(n10130), .ZN(n10129) );
  NAND2X0 U9919 ( .IN1(n10128), .IN2(n2568), .QN(n10130) );
  NAND4X0 U9920 ( .IN1(n10131), .IN2(n9691), .IN3(n10132), .IN4(n10133), .QN(
        n2568) );
  NOR3X0 U9921 ( .IN1(n10134), .IN2(n10135), .IN3(n8576), .QN(n10133) );
  NAND4X0 U9922 ( .IN1(n10132), .IN2(n8576), .IN3(n9679), .IN4(n10136), .QN(
        n10128) );
  NOR4X0 U9923 ( .IN1(n8581), .IN2(n10131), .IN3(n8570), .IN4(n9691), .QN(
        n10136) );
  NOR4X0 U9924 ( .IN1(n8569), .IN2(n8575), .IN3(n8564), .IN4(n10137), .QN(
        n10132) );
  NAND2X0 U9925 ( .IN1(n10138), .IN2(n4513), .QN(n10137) );
  INVX0 U9926 ( .INP(n9529), .ZN(n9680) );
  XNOR2X1 U9927 ( .IN1(n9975), .IN2(n8569), .Q(n10124) );
  NAND2X0 U9928 ( .IN1(n9989), .IN2(n10139), .QN(n9975) );
  XOR2X1 U9929 ( .IN1(n8564), .IN2(n9186), .Q(n10139) );
  NOR2X0 U9930 ( .IN1(n9896), .IN2(n10140), .QN(n9989) );
  XNOR2X1 U9931 ( .IN1(n8575), .IN2(n9186), .Q(n10140) );
  NAND2X0 U9932 ( .IN1(n9658), .IN2(n10141), .QN(n9896) );
  XOR2X1 U9933 ( .IN1(n10135), .IN2(n9186), .Q(n10141) );
  NOR2X0 U9934 ( .IN1(n9532), .IN2(n10142), .QN(n9658) );
  XNOR2X1 U9935 ( .IN1(n8576), .IN2(n9186), .Q(n10142) );
  NAND2X0 U9936 ( .IN1(n9682), .IN2(n10143), .QN(n9532) );
  XOR2X1 U9937 ( .IN1(n10134), .IN2(n9186), .Q(n10143) );
  NOR2X0 U9938 ( .IN1(n10144), .IN2(n9960), .QN(n9682) );
  NOR2X0 U9939 ( .IN1(n8555), .IN2(n9679), .QN(n9960) );
  INVX0 U9940 ( .INP(n9186), .ZN(n9679) );
  XOR2X1 U9941 ( .IN1(n4513), .IN2(n9186), .Q(n10144) );
  INVX0 U9942 ( .INP(n8577), .ZN(n4513) );
  NAND3X0 U9943 ( .IN1(n10145), .IN2(n10146), .IN3(n10147), .QN(n8577) );
  NAND2X0 U9944 ( .IN1(test_so13), .IN2(g6313), .QN(n10147) );
  NAND2X0 U9945 ( .IN1(g6231), .IN2(g186), .QN(n10146) );
  NAND2X0 U9946 ( .IN1(g165), .IN2(g192), .QN(n10145) );
  NAND2X0 U9947 ( .IN1(n9529), .IN2(g121), .QN(n10122) );
  NAND3X0 U9948 ( .IN1(n10148), .IN2(n9388), .IN3(n10149), .QN(n9529) );
  NAND2X0 U9949 ( .IN1(n10150), .IN2(n9412), .QN(n10149) );
  NAND2X0 U9950 ( .IN1(n10151), .IN2(n9398), .QN(n10148) );
  NAND2X0 U9951 ( .IN1(n9416), .IN2(n10152), .QN(n10151) );
  NAND3X0 U9952 ( .IN1(n9412), .IN2(n9405), .IN3(n9759), .QN(n10152) );
  INVX0 U9953 ( .INP(n9415), .ZN(n9412) );
  NAND2X0 U9954 ( .IN1(n10153), .IN2(n10154), .QN(n9415) );
  NAND3X0 U9955 ( .IN1(n10155), .IN2(n10156), .IN3(n10157), .QN(n10154) );
  NAND2X0 U9956 ( .IN1(n7321), .IN2(n10158), .QN(n10157) );
  NAND2X0 U9957 ( .IN1(n7320), .IN2(n10159), .QN(n10156) );
  NAND2X0 U9958 ( .IN1(n7319), .IN2(n10160), .QN(n10155) );
  NAND2X0 U9959 ( .IN1(n10161), .IN2(n10162), .QN(g30072) );
  NAND2X0 U9960 ( .IN1(g2574), .IN2(n7930), .QN(n10162) );
  NAND2X0 U9961 ( .IN1(n4543), .IN2(n10163), .QN(n10161) );
  NAND2X0 U9962 ( .IN1(n10164), .IN2(n10165), .QN(n10163) );
  NAND2X0 U9963 ( .IN1(n497), .IN2(n10166), .QN(n10165) );
  NAND2X0 U9964 ( .IN1(n10167), .IN2(n7929), .QN(n10164) );
  NAND2X0 U9965 ( .IN1(n10168), .IN2(n10169), .QN(g30061) );
  NAND2X0 U9966 ( .IN1(g2580), .IN2(n7926), .QN(n10169) );
  NAND2X0 U9967 ( .IN1(n7489), .IN2(n10170), .QN(n10168) );
  NAND2X0 U9968 ( .IN1(n10171), .IN2(n10172), .QN(n10170) );
  NAND2X0 U9969 ( .IN1(n4370), .IN2(g16437), .QN(n10172) );
  NAND2X0 U9970 ( .IN1(n512), .IN2(g7390), .QN(n10171) );
  INVX0 U9971 ( .INP(n10173), .ZN(n512) );
  NAND2X0 U9972 ( .IN1(n10174), .IN2(n10175), .QN(n10173) );
  NAND2X0 U9973 ( .IN1(g1886), .IN2(DFF_1133_n1), .QN(n10175) );
  NAND2X0 U9974 ( .IN1(n4493), .IN2(n10176), .QN(n10174) );
  NAND2X0 U9975 ( .IN1(n10177), .IN2(n10178), .QN(n10176) );
  NAND2X0 U9976 ( .IN1(n4315), .IN2(DFF_1142_n1), .QN(n10178) );
  NAND2X0 U9977 ( .IN1(n8545), .IN2(g7194), .QN(n10177) );
  NAND2X0 U9978 ( .IN1(n10179), .IN2(n10180), .QN(n8545) );
  NAND2X0 U9979 ( .IN1(g1192), .IN2(DFF_783_n1), .QN(n10180) );
  NAND2X0 U9980 ( .IN1(n4454), .IN2(n10181), .QN(n10179) );
  NAND2X0 U9981 ( .IN1(n10182), .IN2(n10183), .QN(n10181) );
  NAND2X0 U9982 ( .IN1(n4316), .IN2(DFF_792_n1), .QN(n10183) );
  NAND2X0 U9983 ( .IN1(n8544), .IN2(g6944), .QN(n10182) );
  NAND2X0 U9984 ( .IN1(n10184), .IN2(n10185), .QN(n8544) );
  NAND2X0 U9985 ( .IN1(n7406), .IN2(g506), .QN(n10185) );
  NAND3X0 U9986 ( .IN1(n8030), .IN2(n4372), .IN3(n4570), .QN(n10184) );
  NAND2X0 U9987 ( .IN1(n10186), .IN2(n10187), .QN(g30055) );
  NAND2X0 U9988 ( .IN1(n4487), .IN2(DFF_1378_n1), .QN(n10187) );
  NAND2X0 U9989 ( .IN1(n10188), .IN2(g2374), .QN(n10186) );
  NAND2X0 U9990 ( .IN1(n10189), .IN2(n10190), .QN(n10188) );
  NAND2X0 U9991 ( .IN1(n437), .IN2(g7264), .QN(n10190) );
  INVX0 U9992 ( .INP(n10191), .ZN(n437) );
  NAND2X0 U9993 ( .IN1(n10192), .IN2(n10193), .QN(n10191) );
  NAND2X0 U9994 ( .IN1(n4488), .IN2(n7978), .QN(n10193) );
  NAND3X0 U9995 ( .IN1(n10194), .IN2(n10195), .IN3(g1680), .QN(n10192) );
  NAND2X0 U9996 ( .IN1(g7014), .IN2(n438), .QN(n10195) );
  INVX0 U9997 ( .INP(n10196), .ZN(n438) );
  NAND2X0 U9998 ( .IN1(n10197), .IN2(n10198), .QN(n10196) );
  NAND2X0 U9999 ( .IN1(n4432), .IN2(n8017), .QN(n10198) );
  NAND2X0 U10000 ( .IN1(n10199), .IN2(g986), .QN(n10197) );
  NAND2X0 U10001 ( .IN1(n10200), .IN2(n10201), .QN(n10199) );
  NAND2X0 U10002 ( .IN1(n4364), .IN2(n7705), .QN(n10201) );
  INVX0 U10003 ( .INP(n10202), .ZN(n10200) );
  NOR2X0 U10004 ( .IN1(g21346), .IN2(n4364), .QN(n10202) );
  NAND2X0 U10005 ( .IN1(n4525), .IN2(g1686), .QN(n10194) );
  NAND2X0 U10006 ( .IN1(n4524), .IN2(g2380), .QN(n10189) );
  NAND2X0 U10007 ( .IN1(n10203), .IN2(n10204), .QN(g29941) );
  NAND2X0 U10008 ( .IN1(n4494), .IN2(g3105), .QN(n10204) );
  NAND2X0 U10009 ( .IN1(n497), .IN2(g3109), .QN(n10203) );
  NAND2X0 U10010 ( .IN1(n10205), .IN2(n10206), .QN(g29939) );
  NAND2X0 U10011 ( .IN1(n4383), .IN2(g3104), .QN(n10206) );
  NAND2X0 U10012 ( .IN1(n497), .IN2(g8030), .QN(n10205) );
  NAND2X0 U10013 ( .IN1(n10207), .IN2(n10208), .QN(g29936) );
  NAND2X0 U10014 ( .IN1(n4382), .IN2(g3103), .QN(n10208) );
  NAND2X0 U10015 ( .IN1(n497), .IN2(g8106), .QN(n10207) );
  INVX0 U10016 ( .INP(n10209), .ZN(n497) );
  NAND2X0 U10017 ( .IN1(n10210), .IN2(n10211), .QN(n10209) );
  NAND2X0 U10018 ( .IN1(g1880), .IN2(DFF_1099_n1), .QN(n10211) );
  NAND3X0 U10019 ( .IN1(n10212), .IN2(n10213), .IN3(n4545), .QN(n10210) );
  NAND2X0 U10020 ( .IN1(n498), .IN2(n10214), .QN(n10213) );
  NAND2X0 U10021 ( .IN1(n10215), .IN2(n7971), .QN(n10212) );
  NAND2X0 U10022 ( .IN1(n10216), .IN2(n10217), .QN(g29623) );
  NAND2X0 U10023 ( .IN1(n10218), .IN2(n4606), .QN(n10217) );
  NAND2X0 U10024 ( .IN1(n4509), .IN2(g2389), .QN(n10216) );
  NAND2X0 U10025 ( .IN1(n10219), .IN2(n10220), .QN(g29621) );
  NAND2X0 U10026 ( .IN1(n10218), .IN2(g7264), .QN(n10220) );
  NAND2X0 U10027 ( .IN1(n4524), .IN2(g2388), .QN(n10219) );
  NAND2X0 U10028 ( .IN1(n10221), .IN2(n10222), .QN(g29620) );
  NAND2X0 U10029 ( .IN1(n10223), .IN2(n4618), .QN(n10222) );
  NAND2X0 U10030 ( .IN1(n4511), .IN2(g1695), .QN(n10221) );
  NAND2X0 U10031 ( .IN1(n10224), .IN2(n10225), .QN(g29618) );
  NAND2X0 U10032 ( .IN1(n10218), .IN2(g5555), .QN(n10225) );
  INVX0 U10033 ( .INP(n10226), .ZN(n10218) );
  NAND2X0 U10034 ( .IN1(n9698), .IN2(n10227), .QN(n10226) );
  NAND2X0 U10035 ( .IN1(n10228), .IN2(n9189), .QN(n10227) );
  NAND3X0 U10036 ( .IN1(n9703), .IN2(n9699), .IN3(n9709), .QN(n9189) );
  NAND3X0 U10037 ( .IN1(n9708), .IN2(n10229), .IN3(n10230), .QN(n10228) );
  NAND2X0 U10038 ( .IN1(n10022), .IN2(n10231), .QN(n9698) );
  NAND2X0 U10039 ( .IN1(n4516), .IN2(g2387), .QN(n10224) );
  NAND2X0 U10040 ( .IN1(n10232), .IN2(n10233), .QN(g29617) );
  NAND2X0 U10041 ( .IN1(n10223), .IN2(g7014), .QN(n10233) );
  NAND2X0 U10042 ( .IN1(n4525), .IN2(g1694), .QN(n10232) );
  NAND2X0 U10043 ( .IN1(n10234), .IN2(n10235), .QN(g29616) );
  NAND2X0 U10044 ( .IN1(n4381), .IN2(g1001), .QN(n10235) );
  NAND2X0 U10045 ( .IN1(n10236), .IN2(g1088), .QN(n10234) );
  NAND2X0 U10046 ( .IN1(n10237), .IN2(n10238), .QN(g29613) );
  NAND2X0 U10047 ( .IN1(n10223), .IN2(g5511), .QN(n10238) );
  INVX0 U10048 ( .INP(n10239), .ZN(n10223) );
  NAND2X0 U10049 ( .IN1(n9346), .IN2(n10240), .QN(n10239) );
  NAND2X0 U10050 ( .IN1(n10241), .IN2(n9188), .QN(n10240) );
  NAND3X0 U10051 ( .IN1(n9351), .IN2(n9347), .IN3(n9357), .QN(n9188) );
  NAND3X0 U10052 ( .IN1(n9356), .IN2(n10242), .IN3(n10243), .QN(n10241) );
  NAND2X0 U10053 ( .IN1(n10069), .IN2(n10244), .QN(n9346) );
  NAND2X0 U10054 ( .IN1(n4518), .IN2(g1693), .QN(n10237) );
  NAND2X0 U10055 ( .IN1(n10245), .IN2(n10246), .QN(g29612) );
  NAND2X0 U10056 ( .IN1(n4364), .IN2(g1000), .QN(n10246) );
  NAND2X0 U10057 ( .IN1(n10236), .IN2(g6712), .QN(n10245) );
  NAND2X0 U10058 ( .IN1(n10247), .IN2(n10248), .QN(g29611) );
  NAND2X0 U10059 ( .IN1(n10249), .IN2(n4640), .QN(n10248) );
  NAND2X0 U10060 ( .IN1(n4506), .IN2(g314), .QN(n10247) );
  NAND2X0 U10061 ( .IN1(n10250), .IN2(n10251), .QN(g29609) );
  NAND2X0 U10062 ( .IN1(n4363), .IN2(g999), .QN(n10251) );
  NAND2X0 U10063 ( .IN1(n10236), .IN2(g5472), .QN(n10250) );
  NOR2X0 U10064 ( .IN1(n10252), .IN2(n148), .QN(n10236) );
  INVX0 U10065 ( .INP(n10108), .ZN(n148) );
  NAND2X0 U10066 ( .IN1(n10113), .IN2(n10253), .QN(n10108) );
  NOR2X0 U10067 ( .IN1(n9521), .IN2(n10254), .QN(n10252) );
  NOR3X0 U10068 ( .IN1(n9182), .IN2(n9193), .IN3(n10110), .QN(n10254) );
  INVX0 U10069 ( .INP(n9669), .ZN(n9521) );
  NAND3X0 U10070 ( .IN1(n9193), .IN2(n9181), .IN3(n9173), .QN(n9669) );
  NAND2X0 U10071 ( .IN1(n10255), .IN2(n10256), .QN(g29608) );
  NAND2X0 U10072 ( .IN1(n10249), .IN2(g6447), .QN(n10256) );
  NAND2X0 U10073 ( .IN1(n4499), .IN2(g313), .QN(n10255) );
  NAND2X0 U10074 ( .IN1(n10257), .IN2(n10258), .QN(g29606) );
  NAND2X0 U10075 ( .IN1(n10249), .IN2(g5437), .QN(n10258) );
  INVX0 U10076 ( .INP(n10259), .ZN(n10249) );
  NAND2X0 U10077 ( .IN1(n9388), .IN2(n10260), .QN(n10259) );
  NAND2X0 U10078 ( .IN1(n10261), .IN2(n9186), .QN(n10260) );
  NAND3X0 U10079 ( .IN1(n9393), .IN2(n9389), .IN3(n9399), .QN(n9186) );
  NAND3X0 U10080 ( .IN1(n9398), .IN2(n10262), .IN3(n10263), .QN(n10261) );
  NAND2X0 U10081 ( .IN1(n10153), .IN2(n10264), .QN(n9388) );
  NAND2X0 U10082 ( .IN1(n4520), .IN2(g312), .QN(n10257) );
  NOR2X0 U10083 ( .IN1(n10265), .IN2(n10266), .QN(g29582) );
  XNOR2X1 U10084 ( .IN1(n7161), .IN2(n2981), .Q(n10266) );
  NOR2X0 U10085 ( .IN1(n10267), .IN2(n10268), .QN(g29581) );
  XNOR2X1 U10086 ( .IN1(n7162), .IN2(n2984), .Q(n10268) );
  NOR2X0 U10087 ( .IN1(n10269), .IN2(n10270), .QN(g29580) );
  XNOR2X1 U10088 ( .IN1(n7163), .IN2(n2987), .Q(n10270) );
  NOR2X0 U10089 ( .IN1(n10271), .IN2(n10272), .QN(g29579) );
  XNOR2X1 U10090 ( .IN1(n7164), .IN2(n2990), .Q(n10272) );
  NOR2X0 U10091 ( .IN1(n10265), .IN2(n10273), .QN(g29357) );
  XNOR2X1 U10092 ( .IN1(n7322), .IN2(n2982), .Q(n10273) );
  NAND2X0 U10093 ( .IN1(n3159), .IN2(g2129), .QN(n2982) );
  NOR2X0 U10094 ( .IN1(n10267), .IN2(n10274), .QN(g29355) );
  XNOR2X1 U10095 ( .IN1(n7323), .IN2(n2985), .Q(n10274) );
  NAND2X0 U10096 ( .IN1(n3163), .IN2(g1435), .QN(n2985) );
  NOR2X0 U10097 ( .IN1(n10269), .IN2(n10275), .QN(g29354) );
  XNOR2X1 U10098 ( .IN1(n7324), .IN2(n2988), .Q(n10275) );
  NAND2X0 U10099 ( .IN1(n3167), .IN2(test_so36), .QN(n2988) );
  NOR2X0 U10100 ( .IN1(n10271), .IN2(n10276), .QN(g29353) );
  XNOR2X1 U10101 ( .IN1(n7325), .IN2(n2991), .Q(n10276) );
  NAND2X0 U10102 ( .IN1(n3171), .IN2(g61), .QN(n2991) );
  NAND2X0 U10103 ( .IN1(n10277), .IN2(n10278), .QN(g29226) );
  NAND2X0 U10104 ( .IN1(n10279), .IN2(n4606), .QN(n10278) );
  NAND2X0 U10105 ( .IN1(n4509), .IN2(g2498), .QN(n10277) );
  NAND2X0 U10106 ( .IN1(n10280), .IN2(n10281), .QN(g29221) );
  NAND2X0 U10107 ( .IN1(n10279), .IN2(g7264), .QN(n10281) );
  NAND2X0 U10108 ( .IN1(n4524), .IN2(g2495), .QN(n10280) );
  NAND2X0 U10109 ( .IN1(n10282), .IN2(n10283), .QN(g29218) );
  NAND2X0 U10110 ( .IN1(n10284), .IN2(n4618), .QN(n10283) );
  NAND2X0 U10111 ( .IN1(n4511), .IN2(g1804), .QN(n10282) );
  NAND2X0 U10112 ( .IN1(n10285), .IN2(n10286), .QN(g29213) );
  NAND2X0 U10113 ( .IN1(n10279), .IN2(g5555), .QN(n10286) );
  XOR2X1 U10114 ( .IN1(n10287), .IN2(n10288), .Q(n10279) );
  NAND3X0 U10115 ( .IN1(test_so79), .IN2(n10289), .IN3(n10290), .QN(n10287) );
  XOR2X1 U10116 ( .IN1(n10291), .IN2(n10288), .Q(n10290) );
  NAND2X0 U10117 ( .IN1(n10292), .IN2(n10293), .QN(n10289) );
  NAND2X0 U10118 ( .IN1(n10294), .IN2(n10288), .QN(n10293) );
  NAND2X0 U10119 ( .IN1(n10295), .IN2(n10296), .QN(n10292) );
  NAND2X0 U10120 ( .IN1(n4516), .IN2(g2492), .QN(n10285) );
  NAND2X0 U10121 ( .IN1(n10297), .IN2(n10298), .QN(g29212) );
  NAND2X0 U10122 ( .IN1(n10284), .IN2(g7014), .QN(n10298) );
  NAND2X0 U10123 ( .IN1(n4525), .IN2(g1801), .QN(n10297) );
  NAND2X0 U10124 ( .IN1(n10299), .IN2(n10300), .QN(g29209) );
  NAND2X0 U10125 ( .IN1(n4381), .IN2(g1110), .QN(n10300) );
  NAND2X0 U10126 ( .IN1(n10301), .IN2(g1088), .QN(n10299) );
  NAND2X0 U10127 ( .IN1(n10302), .IN2(n10303), .QN(g29205) );
  NAND2X0 U10128 ( .IN1(n10284), .IN2(g5511), .QN(n10303) );
  XOR2X1 U10129 ( .IN1(n10304), .IN2(n10305), .Q(n10284) );
  NAND3X0 U10130 ( .IN1(n10306), .IN2(g1690), .IN3(n10307), .QN(n10304) );
  XOR2X1 U10131 ( .IN1(n4284), .IN2(n10308), .Q(n10307) );
  NAND2X0 U10132 ( .IN1(n10309), .IN2(n10310), .QN(n10306) );
  NAND2X0 U10133 ( .IN1(n10311), .IN2(n10305), .QN(n10310) );
  NAND2X0 U10134 ( .IN1(n10312), .IN2(n10313), .QN(n10309) );
  NAND2X0 U10135 ( .IN1(n4518), .IN2(g1798), .QN(n10302) );
  NAND2X0 U10136 ( .IN1(n10314), .IN2(n10315), .QN(g29204) );
  NAND2X0 U10137 ( .IN1(n4364), .IN2(g1107), .QN(n10315) );
  NAND2X0 U10138 ( .IN1(n10301), .IN2(g6712), .QN(n10314) );
  NAND2X0 U10139 ( .IN1(n10316), .IN2(n10317), .QN(g29201) );
  NAND2X0 U10140 ( .IN1(n10318), .IN2(n4640), .QN(n10317) );
  NAND2X0 U10141 ( .IN1(n4506), .IN2(g423), .QN(n10316) );
  NAND2X0 U10142 ( .IN1(n10319), .IN2(n10320), .QN(g29198) );
  NAND2X0 U10143 ( .IN1(n4363), .IN2(g1104), .QN(n10320) );
  NAND2X0 U10144 ( .IN1(n10301), .IN2(g5472), .QN(n10319) );
  XOR2X1 U10145 ( .IN1(n10321), .IN2(n10322), .Q(n10301) );
  NAND3X0 U10146 ( .IN1(n10323), .IN2(g996), .IN3(n10324), .QN(n10321) );
  XOR2X1 U10147 ( .IN1(n10325), .IN2(n10322), .Q(n10324) );
  NAND2X0 U10148 ( .IN1(n10326), .IN2(n10327), .QN(n10323) );
  NAND2X0 U10149 ( .IN1(n10328), .IN2(n10322), .QN(n10327) );
  NAND2X0 U10150 ( .IN1(n10329), .IN2(n10330), .QN(n10326) );
  NAND2X0 U10151 ( .IN1(n10331), .IN2(n10332), .QN(g29197) );
  NAND2X0 U10152 ( .IN1(n10318), .IN2(g6447), .QN(n10332) );
  NAND2X0 U10153 ( .IN1(n4499), .IN2(g420), .QN(n10331) );
  NAND2X0 U10154 ( .IN1(n10333), .IN2(n10334), .QN(g29194) );
  NAND2X0 U10155 ( .IN1(n10318), .IN2(g5437), .QN(n10334) );
  XOR2X1 U10156 ( .IN1(n10335), .IN2(n10336), .Q(n10318) );
  NAND3X0 U10157 ( .IN1(n10337), .IN2(g309), .IN3(n10338), .QN(n10335) );
  XOR2X1 U10158 ( .IN1(n4282), .IN2(n10339), .Q(n10338) );
  NAND2X0 U10159 ( .IN1(n10340), .IN2(n10341), .QN(n10337) );
  NAND2X0 U10160 ( .IN1(n10342), .IN2(n10336), .QN(n10341) );
  NAND2X0 U10161 ( .IN1(n10343), .IN2(n10344), .QN(n10340) );
  NAND2X0 U10162 ( .IN1(n4520), .IN2(g417), .QN(n10333) );
  NAND2X0 U10163 ( .IN1(n10345), .IN2(n10346), .QN(g29187) );
  NAND2X0 U10164 ( .IN1(n10347), .IN2(g2396), .QN(n10346) );
  NAND2X0 U10165 ( .IN1(n10348), .IN2(n10028), .QN(n10347) );
  NAND2X0 U10166 ( .IN1(n10349), .IN2(n10028), .QN(n10345) );
  NAND2X0 U10167 ( .IN1(n10350), .IN2(n10351), .QN(g29185) );
  NAND2X0 U10168 ( .IN1(n10352), .IN2(g2398), .QN(n10351) );
  NAND2X0 U10169 ( .IN1(n10348), .IN2(n10027), .QN(n10352) );
  NAND2X0 U10170 ( .IN1(n10349), .IN2(n10027), .QN(n10350) );
  NAND2X0 U10171 ( .IN1(n10353), .IN2(n10354), .QN(g29184) );
  NAND2X0 U10172 ( .IN1(n10355), .IN2(g1702), .QN(n10354) );
  NAND2X0 U10173 ( .IN1(n10356), .IN2(n10075), .QN(n10355) );
  NAND2X0 U10174 ( .IN1(n10357), .IN2(n10075), .QN(n10353) );
  NAND2X0 U10175 ( .IN1(n10358), .IN2(n10359), .QN(g29182) );
  NAND2X0 U10176 ( .IN1(n10360), .IN2(g2397), .QN(n10359) );
  NAND2X0 U10177 ( .IN1(n10348), .IN2(n10029), .QN(n10360) );
  INVX0 U10178 ( .INP(n10361), .ZN(n10348) );
  NAND2X0 U10179 ( .IN1(n10349), .IN2(n10029), .QN(n10358) );
  INVX0 U10180 ( .INP(n10362), .ZN(n10349) );
  NAND2X0 U10181 ( .IN1(n10363), .IN2(n10361), .QN(n10362) );
  NAND3X0 U10182 ( .IN1(n10363), .IN2(n10364), .IN3(n10022), .QN(n10361) );
  INVX0 U10183 ( .INP(n10365), .ZN(n10022) );
  NAND2X0 U10184 ( .IN1(n10230), .IN2(n10366), .QN(n10364) );
  NAND3X0 U10185 ( .IN1(n9709), .IN2(n9708), .IN3(n9776), .QN(n10366) );
  INVX0 U10186 ( .INP(n10229), .ZN(n9776) );
  NAND2X0 U10187 ( .IN1(n9713), .IN2(n9710), .QN(n10229) );
  NAND2X0 U10188 ( .IN1(n3038), .IN2(n10367), .QN(n9710) );
  NAND3X0 U10189 ( .IN1(n10368), .IN2(n10369), .IN3(n10370), .QN(n10367) );
  NAND3X0 U10190 ( .IN1(n10371), .IN2(n10372), .IN3(n10373), .QN(n10370) );
  NAND2X0 U10191 ( .IN1(n10374), .IN2(n10375), .QN(n10371) );
  NAND3X0 U10192 ( .IN1(n10376), .IN2(n10377), .IN3(n10378), .QN(n10369) );
  NAND2X0 U10193 ( .IN1(n10379), .IN2(n10380), .QN(n10377) );
  NAND2X0 U10194 ( .IN1(n10381), .IN2(n10374), .QN(n10376) );
  NAND3X0 U10195 ( .IN1(n10382), .IN2(n10383), .IN3(n10384), .QN(n10368) );
  NAND2X0 U10196 ( .IN1(n10380), .IN2(n10374), .QN(n10383) );
  INVX0 U10197 ( .INP(n10385), .ZN(n10374) );
  INVX0 U10198 ( .INP(n10373), .ZN(n10380) );
  NAND2X0 U10199 ( .IN1(n10379), .IN2(n10375), .QN(n10382) );
  INVX0 U10200 ( .INP(n10378), .ZN(n10375) );
  NAND2X0 U10201 ( .IN1(n3038), .IN2(n10386), .QN(n9713) );
  NAND3X0 U10202 ( .IN1(n10387), .IN2(n10388), .IN3(n10389), .QN(n10386) );
  NAND3X0 U10203 ( .IN1(n10390), .IN2(n10391), .IN3(n10392), .QN(n10389) );
  NAND2X0 U10204 ( .IN1(n10393), .IN2(n10394), .QN(n10391) );
  NAND2X0 U10205 ( .IN1(n10395), .IN2(n10396), .QN(n10390) );
  NAND3X0 U10206 ( .IN1(n10397), .IN2(n10398), .IN3(n10399), .QN(n10388) );
  NAND2X0 U10207 ( .IN1(n10395), .IN2(n10394), .QN(n10398) );
  NAND2X0 U10208 ( .IN1(n10400), .IN2(n10396), .QN(n10397) );
  NAND3X0 U10209 ( .IN1(n10401), .IN2(n10402), .IN3(n10403), .QN(n10387) );
  INVX0 U10210 ( .INP(n10395), .ZN(n10403) );
  NAND2X0 U10211 ( .IN1(n10393), .IN2(n10396), .QN(n10402) );
  INVX0 U10212 ( .INP(n10404), .ZN(n10396) );
  NAND2X0 U10213 ( .IN1(n10394), .IN2(n10400), .QN(n10401) );
  INVX0 U10214 ( .INP(n10392), .ZN(n10400) );
  INVX0 U10215 ( .INP(n10405), .ZN(n10394) );
  NAND2X0 U10216 ( .IN1(n10406), .IN2(n10407), .QN(n10363) );
  NAND3X0 U10217 ( .IN1(n3038), .IN2(n9775), .IN3(n10230), .QN(n10407) );
  NAND4X0 U10218 ( .IN1(n10395), .IN2(n10393), .IN3(n10408), .IN4(n10409), 
        .QN(n9775) );
  NOR4X0 U10219 ( .IN1(n10372), .IN2(n10373), .IN3(n10385), .IN4(n10378), .QN(
        n10409) );
  XNOR2X1 U10220 ( .IN1(n8653), .IN2(n4555), .Q(n10378) );
  NAND3X0 U10221 ( .IN1(n10410), .IN2(n10411), .IN3(n10412), .QN(n8653) );
  NAND2X0 U10222 ( .IN1(test_so77), .IN2(test_so73), .QN(n10412) );
  NAND2X0 U10223 ( .IN1(g6837), .IN2(g2324), .QN(n10411) );
  NAND2X0 U10224 ( .IN1(g2241), .IN2(g2330), .QN(n10410) );
  XNOR2X1 U10225 ( .IN1(n8652), .IN2(n4389), .Q(n10385) );
  NAND3X0 U10226 ( .IN1(n10413), .IN2(n10414), .IN3(n10415), .QN(n8652) );
  NAND2X0 U10227 ( .IN1(test_so73), .IN2(g2318), .QN(n10415) );
  NAND2X0 U10228 ( .IN1(g6837), .IN2(g2315), .QN(n10414) );
  NAND2X0 U10229 ( .IN1(g2241), .IN2(g2321), .QN(n10413) );
  XNOR2X1 U10230 ( .IN1(n9570), .IN2(n4373), .Q(n10373) );
  NAND3X0 U10231 ( .IN1(n10416), .IN2(n10417), .IN3(n10418), .QN(n9570) );
  NAND2X0 U10232 ( .IN1(test_so73), .IN2(g2309), .QN(n10418) );
  NAND2X0 U10233 ( .IN1(g6837), .IN2(g2306), .QN(n10417) );
  NAND2X0 U10234 ( .IN1(g2241), .IN2(g2312), .QN(n10416) );
  NAND2X0 U10235 ( .IN1(n10381), .IN2(n10379), .QN(n10372) );
  XOR2X1 U10236 ( .IN1(n8659), .IN2(n4287), .Q(n10379) );
  NAND3X0 U10237 ( .IN1(n10419), .IN2(n10420), .IN3(n10421), .QN(n8659) );
  NAND2X0 U10238 ( .IN1(test_so73), .IN2(g2336), .QN(n10421) );
  NAND2X0 U10239 ( .IN1(g6837), .IN2(g2333), .QN(n10420) );
  NAND2X0 U10240 ( .IN1(g2241), .IN2(g2339), .QN(n10419) );
  INVX0 U10241 ( .INP(n10384), .ZN(n10381) );
  XNOR2X1 U10242 ( .IN1(n8654), .IN2(n9454), .Q(n10384) );
  NAND3X0 U10243 ( .IN1(n10422), .IN2(n10423), .IN3(n10424), .QN(n8654) );
  NAND2X0 U10244 ( .IN1(test_so73), .IN2(g2345), .QN(n10424) );
  NAND2X0 U10245 ( .IN1(g6837), .IN2(g2342), .QN(n10423) );
  NAND2X0 U10246 ( .IN1(g2241), .IN2(g2348), .QN(n10422) );
  NOR3X0 U10247 ( .IN1(n10405), .IN2(n10404), .IN3(n10392), .QN(n10408) );
  XNOR2X1 U10248 ( .IN1(n8660), .IN2(n4377), .Q(n10392) );
  NAND3X0 U10249 ( .IN1(n10425), .IN2(n10426), .IN3(n10427), .QN(n8660) );
  NAND2X0 U10250 ( .IN1(test_so76), .IN2(test_so73), .QN(n10427) );
  NAND2X0 U10251 ( .IN1(g6837), .IN2(g2261), .QN(n10426) );
  NAND2X0 U10252 ( .IN1(g2241), .IN2(g2267), .QN(n10425) );
  XNOR2X1 U10253 ( .IN1(n8658), .IN2(n4563), .Q(n10404) );
  NAND3X0 U10254 ( .IN1(n10428), .IN2(n10429), .IN3(n10430), .QN(n8658) );
  NAND2X0 U10255 ( .IN1(test_so73), .IN2(g2291), .QN(n10430) );
  NAND2X0 U10256 ( .IN1(g6837), .IN2(g2288), .QN(n10429) );
  NAND2X0 U10257 ( .IN1(g2241), .IN2(g2294), .QN(n10428) );
  XNOR2X1 U10258 ( .IN1(n8664), .IN2(n4319), .Q(n10405) );
  NAND3X0 U10259 ( .IN1(n10431), .IN2(n10432), .IN3(n10433), .QN(n8664) );
  NAND2X0 U10260 ( .IN1(test_so73), .IN2(g2273), .QN(n10433) );
  NAND2X0 U10261 ( .IN1(g6837), .IN2(g2270), .QN(n10432) );
  NAND2X0 U10262 ( .IN1(g2241), .IN2(g2276), .QN(n10431) );
  INVX0 U10263 ( .INP(n10399), .ZN(n10393) );
  XNOR2X1 U10264 ( .IN1(n8666), .IN2(n4325), .Q(n10399) );
  NAND3X0 U10265 ( .IN1(n10434), .IN2(n10435), .IN3(n10436), .QN(n8666) );
  NAND2X0 U10266 ( .IN1(test_so73), .IN2(g2282), .QN(n10436) );
  NAND2X0 U10267 ( .IN1(g6837), .IN2(g2279), .QN(n10435) );
  NAND2X0 U10268 ( .IN1(g2241), .IN2(g2285), .QN(n10434) );
  XOR2X1 U10269 ( .IN1(n8665), .IN2(n10437), .Q(n10395) );
  NAND3X0 U10270 ( .IN1(n10438), .IN2(n10439), .IN3(n10440), .QN(n8665) );
  NAND2X0 U10271 ( .IN1(test_so73), .IN2(g2300), .QN(n10440) );
  NAND2X0 U10272 ( .IN1(g6837), .IN2(g2297), .QN(n10439) );
  NAND2X0 U10273 ( .IN1(g2241), .IN2(g2303), .QN(n10438) );
  NAND2X0 U10274 ( .IN1(test_so79), .IN2(n10019), .QN(n10406) );
  NAND2X0 U10275 ( .IN1(n10441), .IN2(n10442), .QN(g29181) );
  NAND2X0 U10276 ( .IN1(n10443), .IN2(g1704), .QN(n10442) );
  NAND2X0 U10277 ( .IN1(n10356), .IN2(n10074), .QN(n10443) );
  NAND2X0 U10278 ( .IN1(n10357), .IN2(n10074), .QN(n10441) );
  NAND2X0 U10279 ( .IN1(n10444), .IN2(n10445), .QN(g29179) );
  NAND2X0 U10280 ( .IN1(n10446), .IN2(g1008), .QN(n10445) );
  NAND2X0 U10281 ( .IN1(n10447), .IN2(g1088), .QN(n10446) );
  NAND2X0 U10282 ( .IN1(n10448), .IN2(g1088), .QN(n10444) );
  NAND2X0 U10283 ( .IN1(n10449), .IN2(n10450), .QN(g29178) );
  NAND2X0 U10284 ( .IN1(n10451), .IN2(g1703), .QN(n10450) );
  NAND2X0 U10285 ( .IN1(n10356), .IN2(n10076), .QN(n10451) );
  INVX0 U10286 ( .INP(n10452), .ZN(n10356) );
  NAND2X0 U10287 ( .IN1(n10357), .IN2(n10076), .QN(n10449) );
  INVX0 U10288 ( .INP(n10453), .ZN(n10357) );
  NAND2X0 U10289 ( .IN1(n10454), .IN2(n10452), .QN(n10453) );
  NAND3X0 U10290 ( .IN1(n10454), .IN2(n10455), .IN3(n10069), .QN(n10452) );
  INVX0 U10291 ( .INP(n10456), .ZN(n10069) );
  NAND2X0 U10292 ( .IN1(n10243), .IN2(n10457), .QN(n10455) );
  NAND3X0 U10293 ( .IN1(n9357), .IN2(n9356), .IN3(n9791), .QN(n10457) );
  INVX0 U10294 ( .INP(n10242), .ZN(n9791) );
  NAND2X0 U10295 ( .IN1(n9361), .IN2(n9358), .QN(n10242) );
  NAND2X0 U10296 ( .IN1(n3070), .IN2(n10458), .QN(n9358) );
  NAND3X0 U10297 ( .IN1(n10459), .IN2(n10460), .IN3(n10461), .QN(n10458) );
  NAND3X0 U10298 ( .IN1(n10462), .IN2(n10463), .IN3(n10464), .QN(n10461) );
  NAND2X0 U10299 ( .IN1(n10465), .IN2(n10466), .QN(n10463) );
  NAND3X0 U10300 ( .IN1(n10467), .IN2(n10468), .IN3(n10469), .QN(n10460) );
  NAND2X0 U10301 ( .IN1(n10466), .IN2(n10470), .QN(n10468) );
  NAND2X0 U10302 ( .IN1(n10465), .IN2(n10471), .QN(n10467) );
  INVX0 U10303 ( .INP(n10472), .ZN(n10465) );
  NAND3X0 U10304 ( .IN1(n10473), .IN2(n10474), .IN3(n10472), .QN(n10459) );
  NAND2X0 U10305 ( .IN1(n10470), .IN2(n10471), .QN(n10474) );
  INVX0 U10306 ( .INP(n10464), .ZN(n10470) );
  NAND2X0 U10307 ( .IN1(n10466), .IN2(n10475), .QN(n10473) );
  INVX0 U10308 ( .INP(n10476), .ZN(n10466) );
  NAND2X0 U10309 ( .IN1(n3070), .IN2(n10477), .QN(n9361) );
  NAND3X0 U10310 ( .IN1(n10478), .IN2(n10479), .IN3(n10480), .QN(n10477) );
  NAND3X0 U10311 ( .IN1(n10481), .IN2(n10482), .IN3(n10483), .QN(n10480) );
  NAND2X0 U10312 ( .IN1(n10484), .IN2(n10485), .QN(n10482) );
  NAND2X0 U10313 ( .IN1(n10486), .IN2(n10487), .QN(n10481) );
  NAND3X0 U10314 ( .IN1(n10488), .IN2(n10489), .IN3(n10490), .QN(n10479) );
  NAND2X0 U10315 ( .IN1(n10486), .IN2(n10485), .QN(n10489) );
  NAND2X0 U10316 ( .IN1(n10491), .IN2(n10487), .QN(n10488) );
  NAND3X0 U10317 ( .IN1(n10492), .IN2(n10493), .IN3(n10494), .QN(n10478) );
  NAND2X0 U10318 ( .IN1(n10484), .IN2(n10487), .QN(n10493) );
  NAND2X0 U10319 ( .IN1(n10485), .IN2(n10491), .QN(n10492) );
  NAND2X0 U10320 ( .IN1(n10495), .IN2(n10496), .QN(n10454) );
  NAND2X0 U10321 ( .IN1(n10066), .IN2(g1690), .QN(n10496) );
  NAND3X0 U10322 ( .IN1(n3070), .IN2(n9790), .IN3(n10243), .QN(n10495) );
  NAND4X0 U10323 ( .IN1(n10486), .IN2(n10484), .IN3(n10497), .IN4(n10498), 
        .QN(n9790) );
  NOR4X0 U10324 ( .IN1(n10464), .IN2(n10462), .IN3(n10476), .IN4(n10472), .QN(
        n10498) );
  XNOR2X1 U10325 ( .IN1(n10499), .IN2(n10056), .Q(n10472) );
  INVX0 U10326 ( .INP(n8630), .ZN(n10056) );
  NAND3X0 U10327 ( .IN1(n10500), .IN2(n10501), .IN3(n10502), .QN(n8630) );
  NAND2X0 U10328 ( .IN1(g6782), .IN2(g1651), .QN(n10502) );
  NAND2X0 U10329 ( .IN1(g6573), .IN2(g1648), .QN(n10501) );
  NAND2X0 U10330 ( .IN1(g1547), .IN2(g1654), .QN(n10500) );
  XNOR2X1 U10331 ( .IN1(g1506), .IN2(n8626), .Q(n10476) );
  INVX0 U10332 ( .INP(n9638), .ZN(n8626) );
  NAND3X0 U10333 ( .IN1(n10503), .IN2(n10504), .IN3(n10505), .QN(n9638) );
  NAND2X0 U10334 ( .IN1(g6782), .IN2(g1642), .QN(n10505) );
  NAND2X0 U10335 ( .IN1(g6573), .IN2(g1639), .QN(n10504) );
  NAND2X0 U10336 ( .IN1(g1547), .IN2(g1645), .QN(n10503) );
  NAND2X0 U10337 ( .IN1(n10475), .IN2(n10471), .QN(n10462) );
  XOR2X1 U10338 ( .IN1(n4390), .IN2(n10043), .Q(n10471) );
  NAND3X0 U10339 ( .IN1(n10506), .IN2(n10507), .IN3(n10508), .QN(n10043) );
  NAND2X0 U10340 ( .IN1(g6782), .IN2(g1624), .QN(n10508) );
  NAND2X0 U10341 ( .IN1(test_so55), .IN2(g6573), .QN(n10507) );
  NAND2X0 U10342 ( .IN1(g1547), .IN2(g1627), .QN(n10506) );
  INVX0 U10343 ( .INP(n10469), .ZN(n10475) );
  XNOR2X1 U10344 ( .IN1(g1496), .IN2(n10061), .Q(n10469) );
  INVX0 U10345 ( .INP(n8629), .ZN(n10061) );
  NAND3X0 U10346 ( .IN1(n10509), .IN2(n10510), .IN3(n10511), .QN(n8629) );
  NAND2X0 U10347 ( .IN1(g6782), .IN2(g1633), .QN(n10511) );
  NAND2X0 U10348 ( .IN1(g6573), .IN2(g1630), .QN(n10510) );
  NAND2X0 U10349 ( .IN1(g1547), .IN2(g1636), .QN(n10509) );
  XOR2X1 U10350 ( .IN1(n4374), .IN2(n8627), .Q(n10464) );
  INVX0 U10351 ( .INP(n10046), .ZN(n8627) );
  NAND3X0 U10352 ( .IN1(n10512), .IN2(n10513), .IN3(n10514), .QN(n10046) );
  NAND2X0 U10353 ( .IN1(g6782), .IN2(g1615), .QN(n10514) );
  NAND2X0 U10354 ( .IN1(g6573), .IN2(g1612), .QN(n10513) );
  NAND2X0 U10355 ( .IN1(g1547), .IN2(g1618), .QN(n10512) );
  INVX0 U10356 ( .INP(n10515), .ZN(n10497) );
  NAND3X0 U10357 ( .IN1(n10485), .IN2(n10487), .IN3(n10491), .QN(n10515) );
  INVX0 U10358 ( .INP(n10483), .ZN(n10491) );
  XOR2X1 U10359 ( .IN1(g1471), .IN2(n8638), .Q(n10483) );
  NAND3X0 U10360 ( .IN1(n10516), .IN2(n10517), .IN3(n10518), .QN(n8638) );
  NAND2X0 U10361 ( .IN1(g6782), .IN2(g1570), .QN(n10518) );
  NAND2X0 U10362 ( .IN1(g6573), .IN2(g1567), .QN(n10517) );
  NAND2X0 U10363 ( .IN1(g1547), .IN2(g1573), .QN(n10516) );
  XOR2X1 U10364 ( .IN1(n4565), .IN2(n10063), .Q(n10487) );
  NAND3X0 U10365 ( .IN1(n10519), .IN2(n10520), .IN3(n10521), .QN(n10063) );
  NAND2X0 U10366 ( .IN1(g6782), .IN2(g1597), .QN(n10521) );
  NAND2X0 U10367 ( .IN1(g6573), .IN2(g1594), .QN(n10520) );
  NAND2X0 U10368 ( .IN1(g1547), .IN2(g1600), .QN(n10519) );
  XNOR2X1 U10369 ( .IN1(g1481), .IN2(n8637), .Q(n10485) );
  NAND3X0 U10370 ( .IN1(n10522), .IN2(n10523), .IN3(n10524), .QN(n8637) );
  NAND2X0 U10371 ( .IN1(g6782), .IN2(g1579), .QN(n10524) );
  NAND2X0 U10372 ( .IN1(g6573), .IN2(g1576), .QN(n10523) );
  NAND2X0 U10373 ( .IN1(g1547), .IN2(g1582), .QN(n10522) );
  INVX0 U10374 ( .INP(n10490), .ZN(n10484) );
  XOR2X1 U10375 ( .IN1(g1491), .IN2(n8640), .Q(n10490) );
  NAND3X0 U10376 ( .IN1(n10525), .IN2(n10526), .IN3(n10527), .QN(n8640) );
  NAND2X0 U10377 ( .IN1(g6782), .IN2(g1588), .QN(n10527) );
  NAND2X0 U10378 ( .IN1(g6573), .IN2(g1585), .QN(n10526) );
  NAND2X0 U10379 ( .IN1(g1547), .IN2(g1591), .QN(n10525) );
  INVX0 U10380 ( .INP(n10494), .ZN(n10486) );
  XNOR2X1 U10381 ( .IN1(n9639), .IN2(n8639), .Q(n10494) );
  INVX0 U10382 ( .INP(n9187), .ZN(n8639) );
  NAND3X0 U10383 ( .IN1(n10528), .IN2(n10529), .IN3(n10530), .QN(n9187) );
  NAND2X0 U10384 ( .IN1(test_so56), .IN2(g6782), .QN(n10530) );
  NAND2X0 U10385 ( .IN1(g6573), .IN2(g1603), .QN(n10529) );
  NAND2X0 U10386 ( .IN1(g1547), .IN2(g1609), .QN(n10528) );
  NAND2X0 U10387 ( .IN1(n10531), .IN2(n10532), .QN(g29173) );
  NAND2X0 U10388 ( .IN1(n10533), .IN2(g1010), .QN(n10532) );
  NAND2X0 U10389 ( .IN1(n10447), .IN2(g6712), .QN(n10533) );
  NAND2X0 U10390 ( .IN1(n10448), .IN2(g6712), .QN(n10531) );
  NAND2X0 U10391 ( .IN1(n10534), .IN2(n10535), .QN(g29172) );
  NAND2X0 U10392 ( .IN1(n10536), .IN2(g321), .QN(n10535) );
  NAND2X0 U10393 ( .IN1(n10537), .IN2(n10160), .QN(n10536) );
  NAND2X0 U10394 ( .IN1(n10538), .IN2(n10160), .QN(n10534) );
  NAND2X0 U10395 ( .IN1(n10539), .IN2(n10540), .QN(g29170) );
  NAND2X0 U10396 ( .IN1(n10541), .IN2(g1009), .QN(n10540) );
  NAND2X0 U10397 ( .IN1(n10447), .IN2(g5472), .QN(n10541) );
  INVX0 U10398 ( .INP(n10542), .ZN(n10447) );
  NAND2X0 U10399 ( .IN1(n10448), .IN2(g5472), .QN(n10539) );
  INVX0 U10400 ( .INP(n10543), .ZN(n10448) );
  NAND2X0 U10401 ( .IN1(n10544), .IN2(n10542), .QN(n10543) );
  NAND3X0 U10402 ( .IN1(n10544), .IN2(n10545), .IN3(n10113), .QN(n10542) );
  INVX0 U10403 ( .INP(n10546), .ZN(n10113) );
  NAND2X0 U10404 ( .IN1(n10547), .IN2(n10548), .QN(n10545) );
  NAND3X0 U10405 ( .IN1(n9173), .IN2(n9179), .IN3(n9182), .QN(n10548) );
  NOR2X0 U10406 ( .IN1(n10549), .IN2(n9201), .QN(n9182) );
  INVX0 U10407 ( .INP(n9212), .ZN(n9201) );
  NAND2X0 U10408 ( .IN1(n3102), .IN2(n10550), .QN(n9212) );
  NAND3X0 U10409 ( .IN1(n10551), .IN2(n10552), .IN3(n10553), .QN(n10550) );
  NAND3X0 U10410 ( .IN1(n10554), .IN2(n10555), .IN3(n10556), .QN(n10553) );
  NAND2X0 U10411 ( .IN1(n10557), .IN2(n10558), .QN(n10555) );
  NAND2X0 U10412 ( .IN1(n10559), .IN2(n10560), .QN(n10554) );
  NAND3X0 U10413 ( .IN1(n10561), .IN2(n10562), .IN3(n10563), .QN(n10552) );
  INVX0 U10414 ( .INP(n10559), .ZN(n10563) );
  NAND2X0 U10415 ( .IN1(n10557), .IN2(n10560), .QN(n10562) );
  NAND2X0 U10416 ( .IN1(n10564), .IN2(n10558), .QN(n10561) );
  NAND3X0 U10417 ( .IN1(n10565), .IN2(n10566), .IN3(n10567), .QN(n10551) );
  INVX0 U10418 ( .INP(n10557), .ZN(n10567) );
  NAND2X0 U10419 ( .IN1(n10559), .IN2(n10558), .QN(n10566) );
  INVX0 U10420 ( .INP(n10568), .ZN(n10558) );
  NAND2X0 U10421 ( .IN1(n10560), .IN2(n10564), .QN(n10565) );
  INVX0 U10422 ( .INP(n9198), .ZN(n10549) );
  NAND2X0 U10423 ( .IN1(n3102), .IN2(n10569), .QN(n9198) );
  NAND3X0 U10424 ( .IN1(n10570), .IN2(n10571), .IN3(n10572), .QN(n10569) );
  NAND3X0 U10425 ( .IN1(n10573), .IN2(n10574), .IN3(n10575), .QN(n10572) );
  NAND2X0 U10426 ( .IN1(n10576), .IN2(n10577), .QN(n10574) );
  NAND2X0 U10427 ( .IN1(n10578), .IN2(n10579), .QN(n10573) );
  NAND3X0 U10428 ( .IN1(n10580), .IN2(n10581), .IN3(n10582), .QN(n10571) );
  NAND2X0 U10429 ( .IN1(n10576), .IN2(n10579), .QN(n10581) );
  NAND2X0 U10430 ( .IN1(n10577), .IN2(n10583), .QN(n10580) );
  NAND3X0 U10431 ( .IN1(n10584), .IN2(n10585), .IN3(n10586), .QN(n10570) );
  INVX0 U10432 ( .INP(n10576), .ZN(n10586) );
  NAND2X0 U10433 ( .IN1(n10578), .IN2(n10577), .QN(n10585) );
  NAND2X0 U10434 ( .IN1(n10579), .IN2(n10583), .QN(n10584) );
  NAND2X0 U10435 ( .IN1(n10587), .IN2(n10588), .QN(n10544) );
  NAND2X0 U10436 ( .IN1(n10110), .IN2(g996), .QN(n10588) );
  NAND3X0 U10437 ( .IN1(n3102), .IN2(n9210), .IN3(n10547), .QN(n10587) );
  NAND4X0 U10438 ( .IN1(n10559), .IN2(n10557), .IN3(n10589), .IN4(n10590), 
        .QN(n9210) );
  NOR4X0 U10439 ( .IN1(n10591), .IN2(n10592), .IN3(n10568), .IN4(n10575), .QN(
        n10590) );
  INVX0 U10440 ( .INP(n10583), .ZN(n10575) );
  XOR2X1 U10441 ( .IN1(n8593), .IN2(n4375), .Q(n10583) );
  NAND3X0 U10442 ( .IN1(n10593), .IN2(n10594), .IN3(n10595), .QN(n8593) );
  NAND2X0 U10443 ( .IN1(test_so34), .IN2(test_so31), .QN(n10595) );
  NAND2X0 U10444 ( .IN1(g6518), .IN2(g921), .QN(n10594) );
  NAND2X0 U10445 ( .IN1(g6368), .IN2(g918), .QN(n10593) );
  XNOR2X1 U10446 ( .IN1(n8594), .IN2(n4567), .Q(n10568) );
  NAND3X0 U10447 ( .IN1(n10596), .IN2(n10597), .IN3(n10598), .QN(n8594) );
  NAND2X0 U10448 ( .IN1(test_so31), .IN2(g906), .QN(n10598) );
  NAND2X0 U10449 ( .IN1(g6518), .IN2(g903), .QN(n10597) );
  NAND2X0 U10450 ( .IN1(g6368), .IN2(g900), .QN(n10596) );
  INVX0 U10451 ( .INP(n10579), .ZN(n10592) );
  XOR2X1 U10452 ( .IN1(n8595), .IN2(n4391), .Q(n10579) );
  NAND3X0 U10453 ( .IN1(n10599), .IN2(n10600), .IN3(n10601), .QN(n8595) );
  NAND2X0 U10454 ( .IN1(test_so31), .IN2(g933), .QN(n10601) );
  NAND2X0 U10455 ( .IN1(g6518), .IN2(g930), .QN(n10600) );
  NAND2X0 U10456 ( .IN1(g6368), .IN2(g927), .QN(n10599) );
  NAND2X0 U10457 ( .IN1(n10577), .IN2(n10564), .QN(n10591) );
  INVX0 U10458 ( .INP(n10556), .ZN(n10564) );
  XNOR2X1 U10459 ( .IN1(n8600), .IN2(n4379), .Q(n10556) );
  NAND3X0 U10460 ( .IN1(n10602), .IN2(n10603), .IN3(n10604), .QN(n8600) );
  NAND2X0 U10461 ( .IN1(test_so31), .IN2(g879), .QN(n10604) );
  NAND2X0 U10462 ( .IN1(g6518), .IN2(g876), .QN(n10603) );
  NAND2X0 U10463 ( .IN1(g6368), .IN2(g873), .QN(n10602) );
  XOR2X1 U10464 ( .IN1(n8610), .IN2(n4289), .Q(n10577) );
  NAND3X0 U10465 ( .IN1(n10605), .IN2(n10606), .IN3(n10607), .QN(n8610) );
  NAND2X0 U10466 ( .IN1(test_so31), .IN2(g951), .QN(n10607) );
  NAND2X0 U10467 ( .IN1(g6518), .IN2(g948), .QN(n10606) );
  NAND2X0 U10468 ( .IN1(test_so35), .IN2(g6368), .QN(n10605) );
  INVX0 U10469 ( .INP(n10608), .ZN(n10589) );
  NAND3X0 U10470 ( .IN1(n10576), .IN2(n10560), .IN3(n10578), .QN(n10608) );
  INVX0 U10471 ( .INP(n10582), .ZN(n10578) );
  XNOR2X1 U10472 ( .IN1(n8601), .IN2(n4559), .Q(n10582) );
  NAND3X0 U10473 ( .IN1(n10609), .IN2(n10610), .IN3(n10611), .QN(n8601) );
  NAND2X0 U10474 ( .IN1(test_so31), .IN2(g942), .QN(n10611) );
  NAND2X0 U10475 ( .IN1(g6518), .IN2(g939), .QN(n10610) );
  NAND2X0 U10476 ( .IN1(g6368), .IN2(g936), .QN(n10609) );
  XOR2X1 U10477 ( .IN1(n8599), .IN2(n4321), .Q(n10560) );
  NAND3X0 U10478 ( .IN1(n10612), .IN2(n10613), .IN3(n10614), .QN(n8599) );
  NAND2X0 U10479 ( .IN1(test_so31), .IN2(g888), .QN(n10614) );
  NAND2X0 U10480 ( .IN1(g6518), .IN2(g885), .QN(n10613) );
  NAND2X0 U10481 ( .IN1(g6368), .IN2(g882), .QN(n10612) );
  XOR2X1 U10482 ( .IN1(n8605), .IN2(n9516), .Q(n10576) );
  NAND3X0 U10483 ( .IN1(n10615), .IN2(n10616), .IN3(n10617), .QN(n8605) );
  NAND2X0 U10484 ( .IN1(test_so31), .IN2(g960), .QN(n10617) );
  NAND2X0 U10485 ( .IN1(g6518), .IN2(g957), .QN(n10616) );
  NAND2X0 U10486 ( .IN1(g6368), .IN2(g954), .QN(n10615) );
  XOR2X1 U10487 ( .IN1(n8607), .IN2(n10618), .Q(n10557) );
  NAND3X0 U10488 ( .IN1(n10619), .IN2(n10620), .IN3(n10621), .QN(n8607) );
  NAND2X0 U10489 ( .IN1(test_so31), .IN2(g915), .QN(n10621) );
  NAND2X0 U10490 ( .IN1(g6518), .IN2(g912), .QN(n10620) );
  NAND2X0 U10491 ( .IN1(g6368), .IN2(g909), .QN(n10619) );
  XOR2X1 U10492 ( .IN1(n8606), .IN2(n4327), .Q(n10559) );
  NAND3X0 U10493 ( .IN1(n10622), .IN2(n10623), .IN3(n10624), .QN(n8606) );
  NAND2X0 U10494 ( .IN1(test_so31), .IN2(g897), .QN(n10624) );
  NAND2X0 U10495 ( .IN1(g6518), .IN2(g894), .QN(n10623) );
  NAND2X0 U10496 ( .IN1(g6368), .IN2(g891), .QN(n10622) );
  NAND2X0 U10497 ( .IN1(n10625), .IN2(n10626), .QN(g29169) );
  NAND2X0 U10498 ( .IN1(n10627), .IN2(g323), .QN(n10626) );
  NAND2X0 U10499 ( .IN1(n10537), .IN2(n10159), .QN(n10627) );
  NAND2X0 U10500 ( .IN1(n10538), .IN2(n10159), .QN(n10625) );
  NAND2X0 U10501 ( .IN1(n10628), .IN2(n10629), .QN(g29167) );
  NAND2X0 U10502 ( .IN1(n10630), .IN2(g322), .QN(n10629) );
  NAND2X0 U10503 ( .IN1(n10537), .IN2(n10158), .QN(n10630) );
  INVX0 U10504 ( .INP(n10631), .ZN(n10537) );
  NAND2X0 U10505 ( .IN1(n10538), .IN2(n10158), .QN(n10628) );
  INVX0 U10506 ( .INP(n10632), .ZN(n10538) );
  NAND2X0 U10507 ( .IN1(n10633), .IN2(n10631), .QN(n10632) );
  NAND3X0 U10508 ( .IN1(n10633), .IN2(n10634), .IN3(n10153), .QN(n10631) );
  INVX0 U10509 ( .INP(n10635), .ZN(n10153) );
  NAND2X0 U10510 ( .IN1(n10263), .IN2(n10636), .QN(n10634) );
  NAND3X0 U10511 ( .IN1(n9399), .IN2(n9398), .IN3(n9759), .QN(n10636) );
  INVX0 U10512 ( .INP(n10262), .ZN(n9759) );
  NAND2X0 U10513 ( .IN1(n9403), .IN2(n9400), .QN(n10262) );
  NAND2X0 U10514 ( .IN1(n3130), .IN2(n10637), .QN(n9400) );
  NAND3X0 U10515 ( .IN1(n10638), .IN2(n10639), .IN3(n10640), .QN(n10637) );
  NAND3X0 U10516 ( .IN1(n10641), .IN2(n10642), .IN3(n10643), .QN(n10640) );
  NAND2X0 U10517 ( .IN1(n10644), .IN2(n10645), .QN(n10642) );
  NAND2X0 U10518 ( .IN1(n10646), .IN2(n10647), .QN(n10641) );
  NAND3X0 U10519 ( .IN1(n10648), .IN2(n10649), .IN3(n10650), .QN(n10639) );
  INVX0 U10520 ( .INP(n10647), .ZN(n10650) );
  NAND2X0 U10521 ( .IN1(n10645), .IN2(n10651), .QN(n10649) );
  NAND2X0 U10522 ( .IN1(n10644), .IN2(n10646), .QN(n10648) );
  NAND3X0 U10523 ( .IN1(n10652), .IN2(n10653), .IN3(n10654), .QN(n10638) );
  NAND2X0 U10524 ( .IN1(n10651), .IN2(n10646), .QN(n10653) );
  NAND2X0 U10525 ( .IN1(n10645), .IN2(n10647), .QN(n10652) );
  NAND2X0 U10526 ( .IN1(n3130), .IN2(n10655), .QN(n9403) );
  NAND3X0 U10527 ( .IN1(n10656), .IN2(n10657), .IN3(n10658), .QN(n10655) );
  NAND3X0 U10528 ( .IN1(n10659), .IN2(n10660), .IN3(n10661), .QN(n10658) );
  NAND2X0 U10529 ( .IN1(n10662), .IN2(n10663), .QN(n10660) );
  NAND2X0 U10530 ( .IN1(n10664), .IN2(n10665), .QN(n10659) );
  NAND3X0 U10531 ( .IN1(n10666), .IN2(n10667), .IN3(n10668), .QN(n10657) );
  NAND2X0 U10532 ( .IN1(n10664), .IN2(n10663), .QN(n10667) );
  INVX0 U10533 ( .INP(n10669), .ZN(n10664) );
  NAND3X0 U10534 ( .IN1(n10670), .IN2(n10671), .IN3(n10669), .QN(n10656) );
  NAND2X0 U10535 ( .IN1(n10662), .IN2(n10665), .QN(n10671) );
  INVX0 U10536 ( .INP(n10668), .ZN(n10662) );
  NAND2X0 U10537 ( .IN1(n10663), .IN2(n10672), .QN(n10670) );
  INVX0 U10538 ( .INP(n10673), .ZN(n10663) );
  NAND2X0 U10539 ( .IN1(n10674), .IN2(n10675), .QN(n10633) );
  NAND2X0 U10540 ( .IN1(n10150), .IN2(g309), .QN(n10675) );
  NAND3X0 U10541 ( .IN1(n3130), .IN2(n9758), .IN3(n10263), .QN(n10674) );
  NAND4X0 U10542 ( .IN1(n10644), .IN2(n10645), .IN3(n10676), .IN4(n10677), 
        .QN(n9758) );
  NOR4X0 U10543 ( .IN1(n10673), .IN2(n10666), .IN3(n10668), .IN4(n10669), .QN(
        n10677) );
  XNOR2X1 U10544 ( .IN1(n9689), .IN2(n9691), .Q(n10669) );
  INVX0 U10545 ( .INP(n8571), .ZN(n9691) );
  NAND3X0 U10546 ( .IN1(n10678), .IN2(n10679), .IN3(n10680), .QN(n8571) );
  NAND2X0 U10547 ( .IN1(g6313), .IN2(g225), .QN(n10680) );
  NAND2X0 U10548 ( .IN1(g6231), .IN2(g222), .QN(n10679) );
  NAND2X0 U10549 ( .IN1(g165), .IN2(g228), .QN(n10678) );
  XOR2X1 U10550 ( .IN1(g113), .IN2(n8575), .Q(n10668) );
  NAND3X0 U10551 ( .IN1(n10681), .IN2(n10682), .IN3(n10683), .QN(n8575) );
  NAND2X0 U10552 ( .IN1(g6313), .IN2(g207), .QN(n10683) );
  NAND2X0 U10553 ( .IN1(g6231), .IN2(g204), .QN(n10682) );
  NAND2X0 U10554 ( .IN1(g165), .IN2(g210), .QN(n10681) );
  NAND2X0 U10555 ( .IN1(n10672), .IN2(n10665), .QN(n10666) );
  XOR2X1 U10556 ( .IN1(n4569), .IN2(n8569), .Q(n10665) );
  NAND3X0 U10557 ( .IN1(n10684), .IN2(n10685), .IN3(n10686), .QN(n8569) );
  NAND2X0 U10558 ( .IN1(g6313), .IN2(g216), .QN(n10686) );
  NAND2X0 U10559 ( .IN1(g6231), .IN2(g213), .QN(n10685) );
  NAND2X0 U10560 ( .IN1(g165), .IN2(g219), .QN(n10684) );
  INVX0 U10561 ( .INP(n10661), .ZN(n10672) );
  XOR2X1 U10562 ( .IN1(n4513), .IN2(n4380), .Q(n10661) );
  XOR2X1 U10563 ( .IN1(g105), .IN2(n8576), .Q(n10673) );
  NAND3X0 U10564 ( .IN1(n10687), .IN2(n10688), .IN3(n10689), .QN(n8576) );
  NAND2X0 U10565 ( .IN1(g6313), .IN2(g198), .QN(n10689) );
  NAND2X0 U10566 ( .IN1(g6231), .IN2(g195), .QN(n10688) );
  NAND2X0 U10567 ( .IN1(g165), .IN2(g201), .QN(n10687) );
  INVX0 U10568 ( .INP(n10690), .ZN(n10676) );
  NAND3X0 U10569 ( .IN1(n10651), .IN2(n10646), .IN3(n10647), .QN(n10690) );
  XNOR2X1 U10570 ( .IN1(n4561), .IN2(n10691), .Q(n10647) );
  INVX0 U10571 ( .INP(n8564), .ZN(n10691) );
  NAND3X0 U10572 ( .IN1(n10692), .IN2(n10693), .IN3(n10694), .QN(n8564) );
  NAND2X0 U10573 ( .IN1(g6313), .IN2(g252), .QN(n10694) );
  NAND2X0 U10574 ( .IN1(g6231), .IN2(g249), .QN(n10693) );
  NAND2X0 U10575 ( .IN1(test_so14), .IN2(g165), .QN(n10692) );
  XNOR2X1 U10576 ( .IN1(n4392), .IN2(n8581), .Q(n10646) );
  INVX0 U10577 ( .INP(n10135), .ZN(n8581) );
  NAND3X0 U10578 ( .IN1(n10695), .IN2(n10696), .IN3(n10697), .QN(n10135) );
  NAND2X0 U10579 ( .IN1(g6313), .IN2(g243), .QN(n10697) );
  NAND2X0 U10580 ( .IN1(g6231), .IN2(g240), .QN(n10696) );
  NAND2X0 U10581 ( .IN1(g165), .IN2(g246), .QN(n10695) );
  INVX0 U10582 ( .INP(n10643), .ZN(n10651) );
  XOR2X1 U10583 ( .IN1(n4376), .IN2(n8570), .Q(n10643) );
  INVX0 U10584 ( .INP(n10134), .ZN(n8570) );
  NAND3X0 U10585 ( .IN1(n10698), .IN2(n10699), .IN3(n10700), .QN(n10134) );
  NAND2X0 U10586 ( .IN1(g6313), .IN2(g234), .QN(n10700) );
  NAND2X0 U10587 ( .IN1(g6231), .IN2(g231), .QN(n10699) );
  NAND2X0 U10588 ( .IN1(g165), .IN2(g237), .QN(n10698) );
  XOR2X1 U10589 ( .IN1(g125), .IN2(n10138), .Q(n10645) );
  INVX0 U10590 ( .INP(n8565), .ZN(n10138) );
  NAND3X0 U10591 ( .IN1(n10701), .IN2(n10702), .IN3(n10703), .QN(n8565) );
  NAND2X0 U10592 ( .IN1(g6313), .IN2(g261), .QN(n10703) );
  NAND2X0 U10593 ( .IN1(g6231), .IN2(g258), .QN(n10702) );
  NAND2X0 U10594 ( .IN1(g165), .IN2(g264), .QN(n10701) );
  INVX0 U10595 ( .INP(n10654), .ZN(n10644) );
  XNOR2X1 U10596 ( .IN1(n10704), .IN2(n10131), .Q(n10654) );
  INVX0 U10597 ( .INP(n8563), .ZN(n10131) );
  NAND3X0 U10598 ( .IN1(n10705), .IN2(n10706), .IN3(n10707), .QN(n8563) );
  NAND2X0 U10599 ( .IN1(g6313), .IN2(g270), .QN(n10707) );
  NAND2X0 U10600 ( .IN1(g6231), .IN2(g267), .QN(n10706) );
  NAND2X0 U10601 ( .IN1(g165), .IN2(g273), .QN(n10705) );
  NOR2X0 U10602 ( .IN1(n10265), .IN2(n10708), .QN(g29112) );
  XOR2X1 U10603 ( .IN1(n8050), .IN2(n3159), .Q(n10708) );
  NOR2X0 U10604 ( .IN1(n10267), .IN2(n10709), .QN(g29111) );
  XOR2X1 U10605 ( .IN1(n8049), .IN2(n3163), .Q(n10709) );
  NOR2X0 U10606 ( .IN1(n10269), .IN2(n10710), .QN(g29110) );
  XNOR2X1 U10607 ( .IN1(n3167), .IN2(test_so36), .Q(n10710) );
  NOR2X0 U10608 ( .IN1(n10271), .IN2(n10711), .QN(g29109) );
  XOR2X1 U10609 ( .IN1(n8048), .IN2(n3171), .Q(n10711) );
  NAND2X0 U10610 ( .IN1(n10712), .IN2(n10713), .QN(g28788) );
  NAND2X0 U10611 ( .IN1(n10714), .IN2(g2501), .QN(n10713) );
  NAND2X0 U10612 ( .IN1(n10715), .IN2(n10028), .QN(n10714) );
  NAND2X0 U10613 ( .IN1(n10716), .IN2(n10028), .QN(n10712) );
  NAND2X0 U10614 ( .IN1(n10717), .IN2(n10718), .QN(g28783) );
  NAND2X0 U10615 ( .IN1(n10719), .IN2(g2503), .QN(n10718) );
  NAND2X0 U10616 ( .IN1(n10715), .IN2(n10027), .QN(n10719) );
  NAND2X0 U10617 ( .IN1(n10716), .IN2(n10027), .QN(n10717) );
  NAND2X0 U10618 ( .IN1(n10720), .IN2(n10721), .QN(g28782) );
  NAND2X0 U10619 ( .IN1(n4606), .IN2(n10722), .QN(n10721) );
  NAND2X0 U10620 ( .IN1(test_so80), .IN2(n4509), .QN(n10720) );
  NAND2X0 U10621 ( .IN1(n10723), .IN2(n10724), .QN(g28778) );
  NAND2X0 U10622 ( .IN1(n10725), .IN2(g1807), .QN(n10724) );
  NAND2X0 U10623 ( .IN1(n10726), .IN2(n10075), .QN(n10725) );
  NAND2X0 U10624 ( .IN1(n10727), .IN2(n10075), .QN(n10723) );
  NAND2X0 U10625 ( .IN1(n10728), .IN2(n10729), .QN(g28774) );
  NAND2X0 U10626 ( .IN1(n10730), .IN2(g2502), .QN(n10729) );
  NAND2X0 U10627 ( .IN1(n10715), .IN2(n10029), .QN(n10730) );
  INVX0 U10628 ( .INP(n10731), .ZN(n10715) );
  NAND3X0 U10629 ( .IN1(test_so79), .IN2(n10732), .IN3(n10733), .QN(n10731) );
  NAND2X0 U10630 ( .IN1(n10716), .IN2(n10029), .QN(n10728) );
  INVX0 U10631 ( .INP(n10734), .ZN(n10716) );
  NAND2X0 U10632 ( .IN1(n10735), .IN2(n10736), .QN(g28773) );
  NAND2X0 U10633 ( .IN1(g7264), .IN2(n10722), .QN(n10736) );
  NAND2X0 U10634 ( .IN1(n4524), .IN2(g2486), .QN(n10735) );
  NAND2X0 U10635 ( .IN1(n10737), .IN2(n10738), .QN(g28772) );
  NAND2X0 U10636 ( .IN1(n10739), .IN2(g1809), .QN(n10738) );
  NAND2X0 U10637 ( .IN1(n10726), .IN2(n10074), .QN(n10739) );
  NAND2X0 U10638 ( .IN1(n10727), .IN2(n10074), .QN(n10737) );
  NAND2X0 U10639 ( .IN1(n10740), .IN2(n10741), .QN(g28771) );
  NAND2X0 U10640 ( .IN1(n4618), .IN2(n10742), .QN(n10741) );
  NAND2X0 U10641 ( .IN1(n4511), .IN2(g1795), .QN(n10740) );
  NAND2X0 U10642 ( .IN1(n10743), .IN2(n10744), .QN(g28767) );
  NAND2X0 U10643 ( .IN1(n10745), .IN2(g1113), .QN(n10744) );
  NAND2X0 U10644 ( .IN1(n10746), .IN2(g1088), .QN(n10745) );
  NAND2X0 U10645 ( .IN1(n10747), .IN2(g1088), .QN(n10743) );
  NAND2X0 U10646 ( .IN1(n10748), .IN2(n10749), .QN(g28763) );
  NAND2X0 U10647 ( .IN1(g5555), .IN2(n10722), .QN(n10749) );
  NAND2X0 U10648 ( .IN1(n10734), .IN2(n10750), .QN(n10722) );
  NAND2X0 U10649 ( .IN1(n10751), .IN2(n10296), .QN(n10750) );
  NAND2X0 U10650 ( .IN1(test_so79), .IN2(n10752), .QN(n10751) );
  NAND2X0 U10651 ( .IN1(n10733), .IN2(n10732), .QN(n10752) );
  INVX0 U10652 ( .INP(n10295), .ZN(n10733) );
  NAND3X0 U10653 ( .IN1(n10753), .IN2(n10754), .IN3(n10755), .QN(n10295) );
  NAND2X0 U10654 ( .IN1(n7656), .IN2(n10027), .QN(n10755) );
  NAND2X0 U10655 ( .IN1(n7665), .IN2(n10028), .QN(n10754) );
  NAND2X0 U10656 ( .IN1(n7666), .IN2(n10029), .QN(n10753) );
  NAND3X0 U10657 ( .IN1(test_so79), .IN2(n10732), .IN3(n10756), .QN(n10734) );
  INVX0 U10658 ( .INP(n10296), .ZN(n10756) );
  NAND3X0 U10659 ( .IN1(n10757), .IN2(n10758), .IN3(n10759), .QN(n10296) );
  NAND2X0 U10660 ( .IN1(g5555), .IN2(g2483), .QN(n10759) );
  NAND2X0 U10661 ( .IN1(test_so80), .IN2(n4606), .QN(n10758) );
  NAND2X0 U10662 ( .IN1(g7264), .IN2(g2486), .QN(n10757) );
  NAND2X0 U10663 ( .IN1(n3196), .IN2(n10760), .QN(n10732) );
  NAND2X0 U10664 ( .IN1(n10291), .IN2(n4285), .QN(n10760) );
  NAND3X0 U10665 ( .IN1(n9726), .IN2(n10288), .IN3(n10761), .QN(n3196) );
  INVX0 U10666 ( .INP(n10291), .ZN(n10761) );
  NAND3X0 U10667 ( .IN1(n10762), .IN2(n9601), .IN3(n10763), .QN(n10291) );
  INVX0 U10668 ( .INP(n10294), .ZN(n9726) );
  NOR2X0 U10669 ( .IN1(n9303), .IN2(n7706), .QN(n10294) );
  NAND3X0 U10670 ( .IN1(n10764), .IN2(n10765), .IN3(n10766), .QN(n9303) );
  NAND2X0 U10671 ( .IN1(n7577), .IN2(test_so73), .QN(n10766) );
  NAND2X0 U10672 ( .IN1(n7578), .IN2(g6837), .QN(n10765) );
  NAND2X0 U10673 ( .IN1(n7576), .IN2(g2241), .QN(n10764) );
  NAND2X0 U10674 ( .IN1(n4516), .IN2(g2483), .QN(n10748) );
  NAND2X0 U10675 ( .IN1(n10767), .IN2(n10768), .QN(g28761) );
  NAND2X0 U10676 ( .IN1(n10769), .IN2(g1808), .QN(n10768) );
  NAND2X0 U10677 ( .IN1(n10726), .IN2(n10076), .QN(n10769) );
  INVX0 U10678 ( .INP(n10770), .ZN(n10726) );
  NAND3X0 U10679 ( .IN1(n10771), .IN2(g1690), .IN3(n10772), .QN(n10770) );
  NAND2X0 U10680 ( .IN1(n10727), .IN2(n10076), .QN(n10767) );
  INVX0 U10681 ( .INP(n10773), .ZN(n10727) );
  NAND2X0 U10682 ( .IN1(n10774), .IN2(n10775), .QN(g28760) );
  NAND2X0 U10683 ( .IN1(g7014), .IN2(n10742), .QN(n10775) );
  NAND2X0 U10684 ( .IN1(n4525), .IN2(g1792), .QN(n10774) );
  NAND2X0 U10685 ( .IN1(n10776), .IN2(n10777), .QN(g28759) );
  NAND2X0 U10686 ( .IN1(n10778), .IN2(g1115), .QN(n10777) );
  NAND2X0 U10687 ( .IN1(n10746), .IN2(g6712), .QN(n10778) );
  NAND2X0 U10688 ( .IN1(n10747), .IN2(g6712), .QN(n10776) );
  NAND2X0 U10689 ( .IN1(n10779), .IN2(n10780), .QN(g28758) );
  NAND2X0 U10690 ( .IN1(n4381), .IN2(g1101), .QN(n10780) );
  NAND2X0 U10691 ( .IN1(n10781), .IN2(g1088), .QN(n10779) );
  NAND2X0 U10692 ( .IN1(n10782), .IN2(n10783), .QN(g28754) );
  NAND2X0 U10693 ( .IN1(n10784), .IN2(g426), .QN(n10783) );
  NAND2X0 U10694 ( .IN1(n10785), .IN2(n10160), .QN(n10784) );
  NAND2X0 U10695 ( .IN1(n10786), .IN2(n10160), .QN(n10782) );
  NAND2X0 U10696 ( .IN1(n10787), .IN2(n10788), .QN(g28749) );
  NAND2X0 U10697 ( .IN1(g5511), .IN2(n10742), .QN(n10788) );
  NAND2X0 U10698 ( .IN1(n10773), .IN2(n10789), .QN(n10742) );
  NAND2X0 U10699 ( .IN1(n10790), .IN2(n10313), .QN(n10789) );
  NAND2X0 U10700 ( .IN1(g1690), .IN2(n10791), .QN(n10790) );
  NAND2X0 U10701 ( .IN1(n10772), .IN2(n10771), .QN(n10791) );
  INVX0 U10702 ( .INP(n10312), .ZN(n10772) );
  NAND3X0 U10703 ( .IN1(n10792), .IN2(n10793), .IN3(n10794), .QN(n10312) );
  NAND2X0 U10704 ( .IN1(n7659), .IN2(n10074), .QN(n10794) );
  NAND2X0 U10705 ( .IN1(n7670), .IN2(n10075), .QN(n10793) );
  NAND2X0 U10706 ( .IN1(n7671), .IN2(n10076), .QN(n10792) );
  NAND3X0 U10707 ( .IN1(n10771), .IN2(g1690), .IN3(n10795), .QN(n10773) );
  INVX0 U10708 ( .INP(n10313), .ZN(n10795) );
  NAND3X0 U10709 ( .IN1(n10796), .IN2(n10797), .IN3(n10798), .QN(n10313) );
  NAND2X0 U10710 ( .IN1(g5511), .IN2(g1789), .QN(n10798) );
  NAND2X0 U10711 ( .IN1(n4618), .IN2(g1795), .QN(n10797) );
  NAND2X0 U10712 ( .IN1(g7014), .IN2(g1792), .QN(n10796) );
  NAND2X0 U10713 ( .IN1(n3212), .IN2(n10799), .QN(n10771) );
  NAND2X0 U10714 ( .IN1(n10800), .IN2(n4284), .QN(n10799) );
  NAND3X0 U10715 ( .IN1(n9374), .IN2(n10305), .IN3(n10308), .QN(n3212) );
  INVX0 U10716 ( .INP(n10800), .ZN(n10308) );
  NAND3X0 U10717 ( .IN1(n10499), .IN2(n9639), .IN3(n10801), .QN(n10800) );
  INVX0 U10718 ( .INP(n10311), .ZN(n9374) );
  NOR2X0 U10719 ( .IN1(n8504), .IN2(n7707), .QN(n10311) );
  NAND3X0 U10720 ( .IN1(n10802), .IN2(n10803), .IN3(n10804), .QN(n8504) );
  NAND2X0 U10721 ( .IN1(n7588), .IN2(g6782), .QN(n10804) );
  NAND2X0 U10722 ( .IN1(n7589), .IN2(g6573), .QN(n10803) );
  NAND2X0 U10723 ( .IN1(n7587), .IN2(g1547), .QN(n10802) );
  NAND2X0 U10724 ( .IN1(n4518), .IN2(g1789), .QN(n10787) );
  NAND2X0 U10725 ( .IN1(n10805), .IN2(n10806), .QN(g28747) );
  NAND2X0 U10726 ( .IN1(n10807), .IN2(g1114), .QN(n10806) );
  NAND2X0 U10727 ( .IN1(n10746), .IN2(g5472), .QN(n10807) );
  INVX0 U10728 ( .INP(n10808), .ZN(n10746) );
  NAND3X0 U10729 ( .IN1(n10809), .IN2(g996), .IN3(n10810), .QN(n10808) );
  NAND2X0 U10730 ( .IN1(n10747), .IN2(g5472), .QN(n10805) );
  INVX0 U10731 ( .INP(n10811), .ZN(n10747) );
  NAND2X0 U10732 ( .IN1(n10812), .IN2(n10813), .QN(g28746) );
  NAND2X0 U10733 ( .IN1(n4364), .IN2(g1098), .QN(n10813) );
  NAND2X0 U10734 ( .IN1(n10781), .IN2(g6712), .QN(n10812) );
  NAND2X0 U10735 ( .IN1(n10814), .IN2(n10815), .QN(g28745) );
  NAND2X0 U10736 ( .IN1(n10816), .IN2(g428), .QN(n10815) );
  NAND2X0 U10737 ( .IN1(n10785), .IN2(n10159), .QN(n10816) );
  NAND2X0 U10738 ( .IN1(n10786), .IN2(n10159), .QN(n10814) );
  NAND2X0 U10739 ( .IN1(n10817), .IN2(n10818), .QN(g28744) );
  NAND2X0 U10740 ( .IN1(n4640), .IN2(n10819), .QN(n10818) );
  NAND2X0 U10741 ( .IN1(n4506), .IN2(g414), .QN(n10817) );
  NAND2X0 U10742 ( .IN1(n10820), .IN2(n10821), .QN(g28738) );
  NAND2X0 U10743 ( .IN1(n4363), .IN2(g1095), .QN(n10821) );
  NAND2X0 U10744 ( .IN1(n10781), .IN2(g5472), .QN(n10820) );
  NAND2X0 U10745 ( .IN1(n10811), .IN2(n10822), .QN(n10781) );
  NAND2X0 U10746 ( .IN1(n10823), .IN2(n10330), .QN(n10822) );
  NAND2X0 U10747 ( .IN1(g996), .IN2(n10824), .QN(n10823) );
  NAND2X0 U10748 ( .IN1(n10810), .IN2(n10809), .QN(n10824) );
  INVX0 U10749 ( .INP(n10329), .ZN(n10810) );
  NAND3X0 U10750 ( .IN1(n10825), .IN2(n10826), .IN3(n10827), .QN(n10329) );
  NAND2X0 U10751 ( .IN1(n7676), .IN2(g1088), .QN(n10827) );
  NAND2X0 U10752 ( .IN1(n7677), .IN2(g5472), .QN(n10826) );
  NAND2X0 U10753 ( .IN1(n7662), .IN2(g6712), .QN(n10825) );
  NAND3X0 U10754 ( .IN1(n10809), .IN2(g996), .IN3(n10828), .QN(n10811) );
  INVX0 U10755 ( .INP(n10330), .ZN(n10828) );
  NAND3X0 U10756 ( .IN1(n10829), .IN2(n10830), .IN3(n10831), .QN(n10330) );
  NAND2X0 U10757 ( .IN1(g1088), .IN2(g1101), .QN(n10831) );
  NAND2X0 U10758 ( .IN1(g5472), .IN2(g1095), .QN(n10830) );
  NAND2X0 U10759 ( .IN1(g6712), .IN2(g1098), .QN(n10829) );
  NAND2X0 U10760 ( .IN1(n3225), .IN2(n10832), .QN(n10809) );
  NAND2X0 U10761 ( .IN1(n10325), .IN2(n4283), .QN(n10832) );
  NAND3X0 U10762 ( .IN1(n9208), .IN2(n10322), .IN3(n10833), .QN(n3225) );
  INVX0 U10763 ( .INP(n10325), .ZN(n10833) );
  NAND3X0 U10764 ( .IN1(n10834), .IN2(n9668), .IN3(n10835), .QN(n10325) );
  INVX0 U10765 ( .INP(n10328), .ZN(n9208) );
  NOR2X0 U10766 ( .IN1(n8524), .IN2(n7708), .QN(n10328) );
  NAND3X0 U10767 ( .IN1(n10836), .IN2(n10837), .IN3(n10838), .QN(n8524) );
  NAND2X0 U10768 ( .IN1(test_so31), .IN2(n7599), .QN(n10838) );
  NAND2X0 U10769 ( .IN1(g6518), .IN2(n8105), .QN(n10837) );
  NAND2X0 U10770 ( .IN1(n7600), .IN2(g6368), .QN(n10836) );
  NAND2X0 U10771 ( .IN1(n10839), .IN2(n10840), .QN(g28736) );
  NAND2X0 U10772 ( .IN1(test_so17), .IN2(n10841), .QN(n10840) );
  NAND2X0 U10773 ( .IN1(n10785), .IN2(n10158), .QN(n10841) );
  INVX0 U10774 ( .INP(n10842), .ZN(n10785) );
  NAND3X0 U10775 ( .IN1(n10843), .IN2(g309), .IN3(n10844), .QN(n10842) );
  NAND2X0 U10776 ( .IN1(n10786), .IN2(n10158), .QN(n10839) );
  INVX0 U10777 ( .INP(n10845), .ZN(n10786) );
  NAND2X0 U10778 ( .IN1(n10846), .IN2(n10847), .QN(g28735) );
  NAND2X0 U10779 ( .IN1(g6447), .IN2(n10819), .QN(n10847) );
  NAND2X0 U10780 ( .IN1(n4499), .IN2(g411), .QN(n10846) );
  NAND2X0 U10781 ( .IN1(n10848), .IN2(n10849), .QN(g28732) );
  NAND2X0 U10782 ( .IN1(g5437), .IN2(n10819), .QN(n10849) );
  NAND2X0 U10783 ( .IN1(n10845), .IN2(n10850), .QN(n10819) );
  NAND2X0 U10784 ( .IN1(n10851), .IN2(n10344), .QN(n10850) );
  NAND2X0 U10785 ( .IN1(g309), .IN2(n10852), .QN(n10851) );
  NAND2X0 U10786 ( .IN1(n10844), .IN2(n10843), .QN(n10852) );
  INVX0 U10787 ( .INP(n10343), .ZN(n10844) );
  NAND3X0 U10788 ( .IN1(n10853), .IN2(n10854), .IN3(n10855), .QN(n10343) );
  NAND2X0 U10789 ( .IN1(n10158), .IN2(n8106), .QN(n10855) );
  NAND2X0 U10790 ( .IN1(n7685), .IN2(n10159), .QN(n10854) );
  NAND2X0 U10791 ( .IN1(n7684), .IN2(n10160), .QN(n10853) );
  NAND3X0 U10792 ( .IN1(n10843), .IN2(g309), .IN3(n10856), .QN(n10845) );
  INVX0 U10793 ( .INP(n10344), .ZN(n10856) );
  NAND3X0 U10794 ( .IN1(n10857), .IN2(n10858), .IN3(n10859), .QN(n10344) );
  NAND2X0 U10795 ( .IN1(g5437), .IN2(g408), .QN(n10859) );
  NAND2X0 U10796 ( .IN1(n4640), .IN2(g414), .QN(n10858) );
  NAND2X0 U10797 ( .IN1(g6447), .IN2(g411), .QN(n10857) );
  NAND2X0 U10798 ( .IN1(n3237), .IN2(n10860), .QN(n10843) );
  NAND2X0 U10799 ( .IN1(n10861), .IN2(n4282), .QN(n10860) );
  NAND3X0 U10800 ( .IN1(n9416), .IN2(n10336), .IN3(n10339), .QN(n3237) );
  INVX0 U10801 ( .INP(n10861), .ZN(n10339) );
  NAND3X0 U10802 ( .IN1(n10704), .IN2(n9689), .IN3(n10862), .QN(n10861) );
  INVX0 U10803 ( .INP(n10342), .ZN(n9416) );
  NOR2X0 U10804 ( .IN1(n9171), .IN2(n7709), .QN(n10342) );
  NAND3X0 U10805 ( .IN1(n10863), .IN2(n10864), .IN3(n10865), .QN(n9171) );
  NAND2X0 U10806 ( .IN1(n7611), .IN2(g6313), .QN(n10865) );
  NAND2X0 U10807 ( .IN1(n7612), .IN2(g6231), .QN(n10864) );
  NAND2X0 U10808 ( .IN1(n7610), .IN2(g165), .QN(n10863) );
  NAND2X0 U10809 ( .IN1(n4520), .IN2(g408), .QN(n10848) );
  NOR2X0 U10810 ( .IN1(n8536), .IN2(n10866), .QN(g28668) );
  XNOR2X1 U10811 ( .IN1(n4418), .IN2(n10867), .Q(n10866) );
  NAND2X0 U10812 ( .IN1(n10868), .IN2(g686), .QN(n10867) );
  NOR2X0 U10813 ( .IN1(n10265), .IN2(n10869), .QN(g28637) );
  XNOR2X1 U10814 ( .IN1(n7687), .IN2(n3160), .Q(n10869) );
  NAND2X0 U10815 ( .IN1(n3424), .IN2(g2138), .QN(n3160) );
  NOR2X0 U10816 ( .IN1(n10267), .IN2(n10870), .QN(g28636) );
  XNOR2X1 U10817 ( .IN1(n7691), .IN2(n3164), .Q(n10870) );
  NAND2X0 U10818 ( .IN1(n3427), .IN2(g1444), .QN(n3164) );
  NOR2X0 U10819 ( .IN1(n10269), .IN2(n10871), .QN(g28635) );
  XNOR2X1 U10820 ( .IN1(n7695), .IN2(n3168), .Q(n10871) );
  NAND2X0 U10821 ( .IN1(n3430), .IN2(g758), .QN(n3168) );
  NOR2X0 U10822 ( .IN1(n10271), .IN2(n10872), .QN(g28634) );
  XNOR2X1 U10823 ( .IN1(n7699), .IN2(n3172), .Q(n10872) );
  NAND2X0 U10824 ( .IN1(n3433), .IN2(g70), .QN(n3172) );
  NAND2X0 U10825 ( .IN1(n10873), .IN2(n10874), .QN(g28425) );
  NAND2X0 U10826 ( .IN1(n4494), .IN2(g3102), .QN(n10874) );
  NAND2X0 U10827 ( .IN1(n498), .IN2(g3109), .QN(n10873) );
  NAND2X0 U10828 ( .IN1(n10875), .IN2(n10876), .QN(g28421) );
  NAND2X0 U10829 ( .IN1(n4383), .IN2(test_so7), .QN(n10876) );
  NAND2X0 U10830 ( .IN1(n498), .IN2(g8030), .QN(n10875) );
  NAND2X0 U10831 ( .IN1(n10877), .IN2(n10878), .QN(g28420) );
  INVX0 U10832 ( .INP(n10879), .ZN(n10878) );
  NOR2X0 U10833 ( .IN1(g8106), .IN2(n4342), .QN(n10879) );
  NAND2X0 U10834 ( .IN1(n498), .IN2(g8106), .QN(n10877) );
  INVX0 U10835 ( .INP(n10880), .ZN(n498) );
  NAND2X0 U10836 ( .IN1(n10881), .IN2(n10882), .QN(n10880) );
  NAND2X0 U10837 ( .IN1(n7141), .IN2(g1186), .QN(n10882) );
  NAND3X0 U10838 ( .IN1(n10883), .IN2(n10884), .IN3(n4548), .QN(n10881) );
  NAND2X0 U10839 ( .IN1(g6750), .IN2(g21851), .QN(n10884) );
  NAND2X0 U10840 ( .IN1(n4371), .IN2(n4361), .QN(n10883) );
  NAND2X0 U10841 ( .IN1(n10885), .IN2(n10886), .QN(g28371) );
  NAND2X0 U10842 ( .IN1(n4299), .IN2(g2694), .QN(n10886) );
  NAND2X0 U10843 ( .IN1(n10887), .IN2(g2624), .QN(n10885) );
  NAND2X0 U10844 ( .IN1(n10888), .IN2(n10889), .QN(g28368) );
  NAND2X0 U10845 ( .IN1(n4370), .IN2(g2691), .QN(n10889) );
  NAND2X0 U10846 ( .IN1(n10887), .IN2(g7390), .QN(n10888) );
  NAND2X0 U10847 ( .IN1(n10890), .IN2(n10891), .QN(g28367) );
  NAND2X0 U10848 ( .IN1(n4299), .IN2(g2685), .QN(n10891) );
  NAND2X0 U10849 ( .IN1(n10892), .IN2(g2624), .QN(n10890) );
  NAND2X0 U10850 ( .IN1(n10893), .IN2(n10894), .QN(g28366) );
  NAND2X0 U10851 ( .IN1(n4366), .IN2(g2000), .QN(n10894) );
  NAND2X0 U10852 ( .IN1(n10895), .IN2(g1930), .QN(n10893) );
  NAND2X0 U10853 ( .IN1(n10896), .IN2(n10897), .QN(g28364) );
  NAND2X0 U10854 ( .IN1(n4314), .IN2(g2688), .QN(n10897) );
  NAND2X0 U10855 ( .IN1(n10887), .IN2(n10166), .QN(n10896) );
  NAND2X0 U10856 ( .IN1(n10898), .IN2(n10899), .QN(n10887) );
  NAND2X0 U10857 ( .IN1(n3252), .IN2(n10900), .QN(n10899) );
  NAND2X0 U10858 ( .IN1(n8876), .IN2(n10901), .QN(n10898) );
  NAND2X0 U10859 ( .IN1(n10902), .IN2(n10903), .QN(g28363) );
  NAND2X0 U10860 ( .IN1(n10892), .IN2(g7390), .QN(n10903) );
  NAND2X0 U10861 ( .IN1(n4370), .IN2(test_so90), .QN(n10902) );
  NAND2X0 U10862 ( .IN1(n10904), .IN2(n10905), .QN(g28362) );
  NAND2X0 U10863 ( .IN1(n4315), .IN2(g1997), .QN(n10905) );
  NAND2X0 U10864 ( .IN1(n10895), .IN2(g7194), .QN(n10904) );
  NAND2X0 U10865 ( .IN1(n10906), .IN2(n10907), .QN(g28361) );
  NAND2X0 U10866 ( .IN1(n4366), .IN2(g1991), .QN(n10907) );
  NAND2X0 U10867 ( .IN1(n10908), .IN2(g1930), .QN(n10906) );
  NAND2X0 U10868 ( .IN1(n10909), .IN2(n10910), .QN(g28360) );
  NAND2X0 U10869 ( .IN1(n4300), .IN2(g1306), .QN(n10910) );
  NAND2X0 U10870 ( .IN1(n10911), .IN2(g1236), .QN(n10909) );
  NAND2X0 U10871 ( .IN1(n10912), .IN2(n10913), .QN(g28358) );
  NAND2X0 U10872 ( .IN1(g7302), .IN2(n10892), .QN(n10913) );
  NAND2X0 U10873 ( .IN1(n10914), .IN2(n10915), .QN(n10892) );
  NAND2X0 U10874 ( .IN1(n8865), .IN2(n10901), .QN(n10915) );
  NAND4X0 U10875 ( .IN1(n10916), .IN2(n9167), .IN3(n9169), .IN4(n10900), .QN(
        n10914) );
  INVX0 U10876 ( .INP(n10917), .ZN(n9169) );
  NAND3X0 U10877 ( .IN1(n10918), .IN2(n10919), .IN3(n10920), .QN(n10917) );
  NAND3X0 U10878 ( .IN1(n10921), .IN2(n10922), .IN3(n10923), .QN(n10920) );
  NAND2X0 U10879 ( .IN1(n10924), .IN2(n10925), .QN(n10923) );
  NAND2X0 U10880 ( .IN1(n10926), .IN2(n10927), .QN(n10925) );
  NAND2X0 U10881 ( .IN1(n10928), .IN2(n10929), .QN(n10922) );
  NAND2X0 U10882 ( .IN1(n10930), .IN2(n10931), .QN(n10921) );
  NAND2X0 U10883 ( .IN1(n10932), .IN2(n10933), .QN(n10930) );
  NAND2X0 U10884 ( .IN1(n10934), .IN2(n10927), .QN(n10919) );
  NAND2X0 U10885 ( .IN1(n10935), .IN2(n10936), .QN(n10934) );
  NAND2X0 U10886 ( .IN1(n10937), .IN2(n10938), .QN(n10936) );
  NAND2X0 U10887 ( .IN1(n10939), .IN2(n10940), .QN(n10937) );
  NAND2X0 U10888 ( .IN1(n10941), .IN2(n10942), .QN(n10940) );
  NAND2X0 U10889 ( .IN1(n10943), .IN2(n10944), .QN(n10935) );
  NAND2X0 U10890 ( .IN1(n10945), .IN2(n10946), .QN(n10918) );
  NAND2X0 U10891 ( .IN1(n10947), .IN2(n10948), .QN(n10946) );
  NAND2X0 U10892 ( .IN1(n10949), .IN2(n10950), .QN(n10948) );
  NAND2X0 U10893 ( .IN1(n10951), .IN2(n10952), .QN(n10950) );
  NAND3X0 U10894 ( .IN1(n10924), .IN2(n10953), .IN3(n10941), .QN(n10952) );
  INVX0 U10895 ( .INP(n10943), .ZN(n10951) );
  NAND2X0 U10896 ( .IN1(n10954), .IN2(n10955), .QN(n10943) );
  NAND2X0 U10897 ( .IN1(n10932), .IN2(n10931), .QN(n10955) );
  NAND2X0 U10898 ( .IN1(n10956), .IN2(n10928), .QN(n10954) );
  NAND2X0 U10899 ( .IN1(n10957), .IN2(n10958), .QN(n10947) );
  NAND2X0 U10900 ( .IN1(n10933), .IN2(n10959), .QN(n10957) );
  NAND2X0 U10901 ( .IN1(n10929), .IN2(n10931), .QN(n10959) );
  NAND2X0 U10902 ( .IN1(n9170), .IN2(n10960), .QN(n9167) );
  NAND2X0 U10903 ( .IN1(n1392), .IN2(n10961), .QN(n10916) );
  INVX0 U10904 ( .INP(n10960), .ZN(n10961) );
  INVX0 U10905 ( .INP(n10962), .ZN(n1392) );
  NAND3X0 U10906 ( .IN1(n10963), .IN2(n10964), .IN3(n10965), .QN(n10962) );
  NAND2X0 U10907 ( .IN1(n10966), .IN2(n10931), .QN(n10965) );
  NAND2X0 U10908 ( .IN1(n10967), .IN2(n10968), .QN(n10966) );
  NAND3X0 U10909 ( .IN1(n10949), .IN2(n10924), .IN3(n10969), .QN(n10968) );
  INVX0 U10910 ( .INP(n10929), .ZN(n10969) );
  NAND2X0 U10911 ( .IN1(n10945), .IN2(n10970), .QN(n10967) );
  NAND3X0 U10912 ( .IN1(n10971), .IN2(n10972), .IN3(n10973), .QN(n10970) );
  NAND2X0 U10913 ( .IN1(n10941), .IN2(n10938), .QN(n10973) );
  NAND3X0 U10914 ( .IN1(n10953), .IN2(n10944), .IN3(n10929), .QN(n10972) );
  NAND2X0 U10915 ( .IN1(n10974), .IN2(n10956), .QN(n10971) );
  NAND3X0 U10916 ( .IN1(n10975), .IN2(n10938), .IN3(n10932), .QN(n10964) );
  NAND2X0 U10917 ( .IN1(n10976), .IN2(n10977), .QN(n10975) );
  NAND2X0 U10918 ( .IN1(n10928), .IN2(n10933), .QN(n10977) );
  NAND2X0 U10919 ( .IN1(n10945), .IN2(n10924), .QN(n10976) );
  INVX0 U10920 ( .INP(n10927), .ZN(n10945) );
  NAND2X0 U10921 ( .IN1(n10978), .IN2(n10927), .QN(n10963) );
  NAND3X0 U10922 ( .IN1(n10979), .IN2(n10980), .IN3(n10981), .QN(n10927) );
  NAND2X0 U10923 ( .IN1(g5796), .IN2(g2426), .QN(n10981) );
  NAND2X0 U10924 ( .IN1(g5747), .IN2(g2424), .QN(n10980) );
  NAND2X0 U10925 ( .IN1(g2412), .IN2(g2428), .QN(n10979) );
  NAND2X0 U10926 ( .IN1(n10982), .IN2(n10983), .QN(n10978) );
  NAND2X0 U10927 ( .IN1(n10956), .IN2(n10958), .QN(n10983) );
  NOR2X0 U10928 ( .IN1(n10941), .IN2(n10932), .QN(n10956) );
  NAND2X0 U10929 ( .IN1(n10928), .IN2(n10984), .QN(n10982) );
  NAND3X0 U10930 ( .IN1(n10942), .IN2(n10985), .IN3(n10986), .QN(n10984) );
  NAND2X0 U10931 ( .IN1(n10974), .IN2(n10941), .QN(n10986) );
  INVX0 U10932 ( .INP(n10933), .ZN(n10941) );
  NAND3X0 U10933 ( .IN1(n10987), .IN2(n10988), .IN3(n10989), .QN(n10933) );
  NAND2X0 U10934 ( .IN1(g5796), .IN2(g2456), .QN(n10989) );
  NAND2X0 U10935 ( .IN1(g5747), .IN2(g2454), .QN(n10988) );
  NAND2X0 U10936 ( .IN1(g2412), .IN2(g2458), .QN(n10987) );
  NAND2X0 U10937 ( .IN1(n10990), .IN2(n10949), .QN(n10985) );
  INVX0 U10938 ( .INP(n10939), .ZN(n10990) );
  NAND3X0 U10939 ( .IN1(n10929), .IN2(n10953), .IN3(n10924), .QN(n10939) );
  NAND3X0 U10940 ( .IN1(n10991), .IN2(n10992), .IN3(n10993), .QN(n10929) );
  NAND2X0 U10941 ( .IN1(g5796), .IN2(g2471), .QN(n10993) );
  NAND2X0 U10942 ( .IN1(g5747), .IN2(g2469), .QN(n10992) );
  NAND2X0 U10943 ( .IN1(test_so85), .IN2(g2412), .QN(n10991) );
  NAND2X0 U10944 ( .IN1(n10932), .IN2(n10944), .QN(n10942) );
  INVX0 U10945 ( .INP(n10953), .ZN(n10932) );
  NAND3X0 U10946 ( .IN1(n10994), .IN2(n10995), .IN3(n10996), .QN(n10953) );
  NAND2X0 U10947 ( .IN1(g5796), .IN2(g2441), .QN(n10996) );
  NAND2X0 U10948 ( .IN1(g5747), .IN2(g2439), .QN(n10995) );
  NAND2X0 U10949 ( .IN1(g2412), .IN2(g2443), .QN(n10994) );
  NAND2X0 U10950 ( .IN1(n4314), .IN2(g2679), .QN(n10912) );
  NAND2X0 U10951 ( .IN1(n10997), .IN2(n10998), .QN(g28357) );
  NAND2X0 U10952 ( .IN1(n4296), .IN2(g1994), .QN(n10998) );
  NAND2X0 U10953 ( .IN1(n10895), .IN2(n10214), .QN(n10997) );
  NAND2X0 U10954 ( .IN1(n10999), .IN2(n11000), .QN(n10895) );
  NAND2X0 U10955 ( .IN1(n9002), .IN2(n10901), .QN(n11000) );
  NAND4X0 U10956 ( .IN1(n11001), .IN2(n11002), .IN3(n11003), .IN4(n10900), 
        .QN(n10999) );
  NAND2X0 U10957 ( .IN1(n11004), .IN2(n11005), .QN(n11001) );
  INVX0 U10958 ( .INP(n11006), .ZN(n11004) );
  NAND2X0 U10959 ( .IN1(n11007), .IN2(n11008), .QN(g28356) );
  NAND2X0 U10960 ( .IN1(n4315), .IN2(g1988), .QN(n11008) );
  NAND2X0 U10961 ( .IN1(n10908), .IN2(g7194), .QN(n11007) );
  NAND2X0 U10962 ( .IN1(n11009), .IN2(n11010), .QN(g28355) );
  NAND2X0 U10963 ( .IN1(n4316), .IN2(g1303), .QN(n11010) );
  NAND2X0 U10964 ( .IN1(n10911), .IN2(g6944), .QN(n11009) );
  NAND2X0 U10965 ( .IN1(n11011), .IN2(n11012), .QN(g28354) );
  NAND2X0 U10966 ( .IN1(n4300), .IN2(g1297), .QN(n11012) );
  NAND2X0 U10967 ( .IN1(n11013), .IN2(g1236), .QN(n11011) );
  NAND2X0 U10968 ( .IN1(n11014), .IN2(n11015), .QN(g28353) );
  NAND2X0 U10969 ( .IN1(n11016), .IN2(g550), .QN(n11015) );
  NAND2X0 U10970 ( .IN1(test_so26), .IN2(n4313), .QN(n11014) );
  NAND2X0 U10971 ( .IN1(n11017), .IN2(n11018), .QN(g28352) );
  NAND2X0 U10972 ( .IN1(g7052), .IN2(n10908), .QN(n11018) );
  NAND2X0 U10973 ( .IN1(n11019), .IN2(n11020), .QN(n10908) );
  NAND2X0 U10974 ( .IN1(n8980), .IN2(n10901), .QN(n11020) );
  NAND4X0 U10975 ( .IN1(n11002), .IN2(n11021), .IN3(n11005), .IN4(n10900), 
        .QN(n11019) );
  INVX0 U10976 ( .INP(n11022), .ZN(n11005) );
  NAND4X0 U10977 ( .IN1(n11023), .IN2(n11024), .IN3(n11025), .IN4(n11026), 
        .QN(n11022) );
  NAND2X0 U10978 ( .IN1(n11027), .IN2(n11028), .QN(n11026) );
  NAND2X0 U10979 ( .IN1(n11029), .IN2(n11030), .QN(n11028) );
  NAND2X0 U10980 ( .IN1(n11031), .IN2(n11032), .QN(n11030) );
  INVX0 U10981 ( .INP(n11033), .ZN(n11032) );
  NAND2X0 U10982 ( .IN1(n11034), .IN2(n11035), .QN(n11029) );
  NAND3X0 U10983 ( .IN1(n11036), .IN2(n11037), .IN3(n11038), .QN(n11025) );
  NAND2X0 U10984 ( .IN1(n11033), .IN2(n11039), .QN(n11037) );
  NAND2X0 U10985 ( .IN1(n11035), .IN2(n11040), .QN(n11039) );
  NAND2X0 U10986 ( .IN1(n11041), .IN2(n11042), .QN(n11035) );
  NAND2X0 U10987 ( .IN1(n11043), .IN2(n11044), .QN(n11042) );
  NOR2X0 U10988 ( .IN1(n11045), .IN2(n11046), .QN(n11033) );
  NOR2X0 U10989 ( .IN1(n11047), .IN2(n11044), .QN(n11046) );
  NOR2X0 U10990 ( .IN1(n11041), .IN2(n11048), .QN(n11045) );
  NAND2X0 U10991 ( .IN1(n11048), .IN2(n11049), .QN(n11024) );
  NAND2X0 U10992 ( .IN1(n11050), .IN2(n11051), .QN(n11049) );
  NAND3X0 U10993 ( .IN1(n11052), .IN2(n11053), .IN3(n11054), .QN(n11051) );
  NAND2X0 U10994 ( .IN1(n11055), .IN2(n11056), .QN(n11050) );
  NAND2X0 U10995 ( .IN1(n11040), .IN2(n11057), .QN(n11055) );
  NAND2X0 U10996 ( .IN1(n11058), .IN2(n11038), .QN(n11057) );
  NAND3X0 U10997 ( .IN1(n11059), .IN2(n11047), .IN3(n11044), .QN(n11023) );
  NAND2X0 U10998 ( .IN1(n11060), .IN2(n11061), .QN(n11059) );
  NAND2X0 U10999 ( .IN1(n11041), .IN2(n11062), .QN(n11061) );
  NAND2X0 U11000 ( .IN1(n11040), .IN2(n11063), .QN(n11062) );
  NAND2X0 U11001 ( .IN1(n11054), .IN2(n11053), .QN(n11060) );
  NAND2X0 U11002 ( .IN1(n11064), .IN2(n11003), .QN(n11021) );
  INVX0 U11003 ( .INP(n11065), .ZN(n11003) );
  NAND3X0 U11004 ( .IN1(n11066), .IN2(n11067), .IN3(n11068), .QN(n11065) );
  NAND2X0 U11005 ( .IN1(n11069), .IN2(n11038), .QN(n11068) );
  NAND2X0 U11006 ( .IN1(n11070), .IN2(n11071), .QN(n11069) );
  NAND2X0 U11007 ( .IN1(n11034), .IN2(n11052), .QN(n11071) );
  INVX0 U11008 ( .INP(n11058), .ZN(n11034) );
  NAND2X0 U11009 ( .IN1(n11048), .IN2(n11072), .QN(n11070) );
  NAND3X0 U11010 ( .IN1(n11073), .IN2(n11074), .IN3(n11075), .QN(n11072) );
  NAND2X0 U11011 ( .IN1(n11054), .IN2(n11047), .QN(n11075) );
  NAND2X0 U11012 ( .IN1(n11076), .IN2(n11077), .QN(n11074) );
  NAND2X0 U11013 ( .IN1(n11078), .IN2(n11031), .QN(n11073) );
  NAND3X0 U11014 ( .IN1(n11079), .IN2(n11047), .IN3(n11036), .QN(n11067) );
  NAND2X0 U11015 ( .IN1(n11080), .IN2(n11081), .QN(n11079) );
  NAND2X0 U11016 ( .IN1(n11027), .IN2(n11040), .QN(n11081) );
  NAND2X0 U11017 ( .IN1(n11048), .IN2(n11041), .QN(n11080) );
  INVX0 U11018 ( .INP(n11044), .ZN(n11048) );
  NAND2X0 U11019 ( .IN1(n11082), .IN2(n11044), .QN(n11066) );
  NAND3X0 U11020 ( .IN1(n11083), .IN2(n11084), .IN3(n11085), .QN(n11044) );
  NAND2X0 U11021 ( .IN1(test_so63), .IN2(g1730), .QN(n11085) );
  NAND2X0 U11022 ( .IN1(g1718), .IN2(g1734), .QN(n11084) );
  NAND2X0 U11023 ( .IN1(g5738), .IN2(g1732), .QN(n11083) );
  NAND2X0 U11024 ( .IN1(n11086), .IN2(n11087), .QN(n11082) );
  NAND2X0 U11025 ( .IN1(n11031), .IN2(n11056), .QN(n11087) );
  NOR2X0 U11026 ( .IN1(n11054), .IN2(n11036), .QN(n11031) );
  NAND2X0 U11027 ( .IN1(n11027), .IN2(n11088), .QN(n11086) );
  NAND3X0 U11028 ( .IN1(n11089), .IN2(n11090), .IN3(n11091), .QN(n11088) );
  NAND2X0 U11029 ( .IN1(n11078), .IN2(n11054), .QN(n11091) );
  INVX0 U11030 ( .INP(n11040), .ZN(n11054) );
  NAND3X0 U11031 ( .IN1(n11092), .IN2(n11093), .IN3(n11094), .QN(n11040) );
  NAND2X0 U11032 ( .IN1(test_so63), .IN2(g1760), .QN(n11094) );
  NAND2X0 U11033 ( .IN1(g1718), .IN2(g1764), .QN(n11093) );
  NAND2X0 U11034 ( .IN1(g5738), .IN2(g1762), .QN(n11092) );
  NAND2X0 U11035 ( .IN1(n11052), .IN2(n11076), .QN(n11090) );
  INVX0 U11036 ( .INP(n11063), .ZN(n11076) );
  NAND2X0 U11037 ( .IN1(n11058), .IN2(n11053), .QN(n11063) );
  NAND3X0 U11038 ( .IN1(n11095), .IN2(n11096), .IN3(n11097), .QN(n11058) );
  NAND2X0 U11039 ( .IN1(test_so63), .IN2(g1775), .QN(n11097) );
  NAND2X0 U11040 ( .IN1(g1718), .IN2(g1705), .QN(n11096) );
  NAND2X0 U11041 ( .IN1(g5738), .IN2(g1777), .QN(n11095) );
  NAND2X0 U11042 ( .IN1(n11036), .IN2(n11077), .QN(n11089) );
  INVX0 U11043 ( .INP(n11053), .ZN(n11036) );
  NAND3X0 U11044 ( .IN1(n11098), .IN2(n11099), .IN3(n11100), .QN(n11053) );
  NAND2X0 U11045 ( .IN1(test_so63), .IN2(g1745), .QN(n11100) );
  NAND2X0 U11046 ( .IN1(g1718), .IN2(g1749), .QN(n11099) );
  NAND2X0 U11047 ( .IN1(g5738), .IN2(g1747), .QN(n11098) );
  INVX0 U11048 ( .INP(n11101), .ZN(n11064) );
  NAND2X0 U11049 ( .IN1(n11006), .IN2(n11101), .QN(n11002) );
  NAND2X0 U11050 ( .IN1(n4296), .IN2(g1985), .QN(n11017) );
  NAND2X0 U11051 ( .IN1(n11102), .IN2(n11103), .QN(g28351) );
  NAND2X0 U11052 ( .IN1(n4371), .IN2(g1300), .QN(n11103) );
  NAND2X0 U11053 ( .IN1(n10911), .IN2(n11104), .QN(n11102) );
  NAND2X0 U11054 ( .IN1(n11105), .IN2(n11106), .QN(n10911) );
  NAND2X0 U11055 ( .IN1(n9108), .IN2(n10901), .QN(n11106) );
  NAND4X0 U11056 ( .IN1(n11107), .IN2(n11108), .IN3(n11109), .IN4(n10900), 
        .QN(n11105) );
  NAND2X0 U11057 ( .IN1(n11110), .IN2(n11111), .QN(n11107) );
  INVX0 U11058 ( .INP(n11112), .ZN(n11110) );
  NAND2X0 U11059 ( .IN1(n11113), .IN2(n11114), .QN(g28350) );
  NAND2X0 U11060 ( .IN1(n4316), .IN2(g1294), .QN(n11114) );
  NAND2X0 U11061 ( .IN1(n11013), .IN2(g6944), .QN(n11113) );
  NAND2X0 U11062 ( .IN1(n11115), .IN2(n11116), .QN(g28349) );
  NAND2X0 U11063 ( .IN1(n4372), .IN2(g617), .QN(n11116) );
  NAND2X0 U11064 ( .IN1(n11016), .IN2(g6642), .QN(n11115) );
  NAND2X0 U11065 ( .IN1(n11117), .IN2(n11118), .QN(g28348) );
  NAND2X0 U11066 ( .IN1(n4313), .IN2(g611), .QN(n11118) );
  NAND2X0 U11067 ( .IN1(n11119), .IN2(g550), .QN(n11117) );
  NAND2X0 U11068 ( .IN1(n11120), .IN2(n11121), .QN(g28346) );
  NAND2X0 U11069 ( .IN1(g6750), .IN2(n11013), .QN(n11121) );
  NAND2X0 U11070 ( .IN1(n11122), .IN2(n11123), .QN(n11013) );
  NAND2X0 U11071 ( .IN1(n9097), .IN2(n10901), .QN(n11123) );
  NAND4X0 U11072 ( .IN1(n11108), .IN2(n11124), .IN3(n11111), .IN4(n10900), 
        .QN(n11122) );
  INVX0 U11073 ( .INP(n11125), .ZN(n11111) );
  NAND4X0 U11074 ( .IN1(n11126), .IN2(n11127), .IN3(n11128), .IN4(n11129), 
        .QN(n11125) );
  NAND2X0 U11075 ( .IN1(n11130), .IN2(n11131), .QN(n11129) );
  NAND2X0 U11076 ( .IN1(n11132), .IN2(n11133), .QN(n11131) );
  NAND2X0 U11077 ( .IN1(n11134), .IN2(n11135), .QN(n11133) );
  INVX0 U11078 ( .INP(n11136), .ZN(n11135) );
  NAND2X0 U11079 ( .IN1(n11137), .IN2(n11138), .QN(n11132) );
  NAND3X0 U11080 ( .IN1(n11139), .IN2(n11140), .IN3(n11141), .QN(n11128) );
  NAND2X0 U11081 ( .IN1(n11136), .IN2(n11142), .QN(n11140) );
  NAND2X0 U11082 ( .IN1(n11138), .IN2(n11143), .QN(n11142) );
  NAND2X0 U11083 ( .IN1(n11144), .IN2(n11145), .QN(n11138) );
  NAND2X0 U11084 ( .IN1(n11146), .IN2(n11147), .QN(n11145) );
  NOR2X0 U11085 ( .IN1(n11148), .IN2(n11149), .QN(n11136) );
  NOR2X0 U11086 ( .IN1(n11150), .IN2(n11147), .QN(n11149) );
  NOR2X0 U11087 ( .IN1(n11144), .IN2(n11151), .QN(n11148) );
  NAND2X0 U11088 ( .IN1(n11151), .IN2(n11152), .QN(n11127) );
  NAND2X0 U11089 ( .IN1(n11153), .IN2(n11154), .QN(n11152) );
  NAND3X0 U11090 ( .IN1(n11155), .IN2(n11156), .IN3(n11157), .QN(n11154) );
  NAND2X0 U11091 ( .IN1(n11158), .IN2(n11159), .QN(n11153) );
  NAND2X0 U11092 ( .IN1(n11143), .IN2(n11160), .QN(n11158) );
  NAND2X0 U11093 ( .IN1(n11161), .IN2(n11141), .QN(n11160) );
  NAND3X0 U11094 ( .IN1(n11162), .IN2(n11150), .IN3(n11147), .QN(n11126) );
  NAND2X0 U11095 ( .IN1(n11163), .IN2(n11164), .QN(n11162) );
  NAND2X0 U11096 ( .IN1(n11144), .IN2(n11165), .QN(n11164) );
  NAND2X0 U11097 ( .IN1(n11143), .IN2(n11166), .QN(n11165) );
  NAND2X0 U11098 ( .IN1(n11157), .IN2(n11156), .QN(n11163) );
  NAND2X0 U11099 ( .IN1(n11167), .IN2(n11109), .QN(n11124) );
  INVX0 U11100 ( .INP(n11168), .ZN(n11109) );
  NAND3X0 U11101 ( .IN1(n11169), .IN2(n11170), .IN3(n11171), .QN(n11168) );
  NAND2X0 U11102 ( .IN1(n11172), .IN2(n11141), .QN(n11171) );
  NAND2X0 U11103 ( .IN1(n11173), .IN2(n11174), .QN(n11172) );
  NAND2X0 U11104 ( .IN1(n11137), .IN2(n11155), .QN(n11174) );
  INVX0 U11105 ( .INP(n11161), .ZN(n11137) );
  NAND2X0 U11106 ( .IN1(n11151), .IN2(n11175), .QN(n11173) );
  NAND3X0 U11107 ( .IN1(n11176), .IN2(n11177), .IN3(n11178), .QN(n11175) );
  NAND2X0 U11108 ( .IN1(n11157), .IN2(n11150), .QN(n11178) );
  NAND2X0 U11109 ( .IN1(n11179), .IN2(n11180), .QN(n11177) );
  NAND2X0 U11110 ( .IN1(n11181), .IN2(n11134), .QN(n11176) );
  NAND3X0 U11111 ( .IN1(n11182), .IN2(n11150), .IN3(n11139), .QN(n11170) );
  NAND2X0 U11112 ( .IN1(n11183), .IN2(n11184), .QN(n11182) );
  NAND2X0 U11113 ( .IN1(n11130), .IN2(n11143), .QN(n11184) );
  NAND2X0 U11114 ( .IN1(n11151), .IN2(n11144), .QN(n11183) );
  INVX0 U11115 ( .INP(n11147), .ZN(n11151) );
  NAND2X0 U11116 ( .IN1(n11185), .IN2(n11147), .QN(n11169) );
  NAND3X0 U11117 ( .IN1(n11186), .IN2(n11187), .IN3(n11188), .QN(n11147) );
  NAND2X0 U11118 ( .IN1(g5686), .IN2(g1038), .QN(n11188) );
  NAND2X0 U11119 ( .IN1(g5657), .IN2(g1036), .QN(n11187) );
  NAND2X0 U11120 ( .IN1(g1024), .IN2(g1040), .QN(n11186) );
  NAND2X0 U11121 ( .IN1(n11189), .IN2(n11190), .QN(n11185) );
  NAND2X0 U11122 ( .IN1(n11134), .IN2(n11159), .QN(n11190) );
  NOR2X0 U11123 ( .IN1(n11157), .IN2(n11139), .QN(n11134) );
  NAND2X0 U11124 ( .IN1(n11130), .IN2(n11191), .QN(n11189) );
  NAND3X0 U11125 ( .IN1(n11192), .IN2(n11193), .IN3(n11194), .QN(n11191) );
  NAND2X0 U11126 ( .IN1(n11181), .IN2(n11157), .QN(n11194) );
  INVX0 U11127 ( .INP(n11143), .ZN(n11157) );
  NAND3X0 U11128 ( .IN1(n11195), .IN2(n11196), .IN3(n11197), .QN(n11143) );
  NAND2X0 U11129 ( .IN1(g5686), .IN2(g1068), .QN(n11197) );
  NAND2X0 U11130 ( .IN1(g5657), .IN2(g1066), .QN(n11196) );
  NAND2X0 U11131 ( .IN1(g1024), .IN2(g1070), .QN(n11195) );
  NAND2X0 U11132 ( .IN1(n11155), .IN2(n11179), .QN(n11193) );
  INVX0 U11133 ( .INP(n11166), .ZN(n11179) );
  NAND2X0 U11134 ( .IN1(n11161), .IN2(n11156), .QN(n11166) );
  NAND3X0 U11135 ( .IN1(n11198), .IN2(n11199), .IN3(n11200), .QN(n11161) );
  NAND2X0 U11136 ( .IN1(g5686), .IN2(g1083), .QN(n11200) );
  NAND2X0 U11137 ( .IN1(g5657), .IN2(g1081), .QN(n11199) );
  NAND2X0 U11138 ( .IN1(g1024), .IN2(g1011), .QN(n11198) );
  NAND2X0 U11139 ( .IN1(n11139), .IN2(n11180), .QN(n11192) );
  INVX0 U11140 ( .INP(n11156), .ZN(n11139) );
  NAND3X0 U11141 ( .IN1(n11201), .IN2(n11202), .IN3(n11203), .QN(n11156) );
  NAND2X0 U11142 ( .IN1(g5686), .IN2(g1053), .QN(n11203) );
  NAND2X0 U11143 ( .IN1(g5657), .IN2(g1051), .QN(n11202) );
  NAND2X0 U11144 ( .IN1(g1024), .IN2(g1055), .QN(n11201) );
  INVX0 U11145 ( .INP(n11204), .ZN(n11167) );
  NAND2X0 U11146 ( .IN1(n11112), .IN2(n11204), .QN(n11108) );
  NAND2X0 U11147 ( .IN1(n4371), .IN2(g1291), .QN(n11120) );
  NAND2X0 U11148 ( .IN1(n11205), .IN2(n11206), .QN(g28345) );
  NAND2X0 U11149 ( .IN1(n4298), .IN2(g614), .QN(n11206) );
  NAND2X0 U11150 ( .IN1(n11016), .IN2(n11207), .QN(n11205) );
  NAND2X0 U11151 ( .IN1(n11208), .IN2(n11209), .QN(n11016) );
  NAND2X0 U11152 ( .IN1(n8751), .IN2(n10901), .QN(n11209) );
  NAND4X0 U11153 ( .IN1(n11210), .IN2(n11211), .IN3(n11212), .IN4(n10900), 
        .QN(n11208) );
  NAND2X0 U11154 ( .IN1(n11213), .IN2(n11214), .QN(n11210) );
  INVX0 U11155 ( .INP(n11215), .ZN(n11213) );
  NAND2X0 U11156 ( .IN1(n11216), .IN2(n11217), .QN(g28344) );
  NAND2X0 U11157 ( .IN1(n4372), .IN2(g608), .QN(n11217) );
  NAND2X0 U11158 ( .IN1(n11119), .IN2(g6642), .QN(n11216) );
  NAND2X0 U11159 ( .IN1(n11218), .IN2(n11219), .QN(g28342) );
  NAND2X0 U11160 ( .IN1(g6485), .IN2(n11119), .QN(n11219) );
  NAND2X0 U11161 ( .IN1(n11220), .IN2(n11221), .QN(n11119) );
  NAND2X0 U11162 ( .IN1(n8745), .IN2(n10901), .QN(n11221) );
  NAND4X0 U11163 ( .IN1(n11211), .IN2(n11222), .IN3(n11214), .IN4(n10900), 
        .QN(n11220) );
  INVX0 U11164 ( .INP(n11223), .ZN(n11214) );
  NAND4X0 U11165 ( .IN1(n11224), .IN2(n11225), .IN3(n11226), .IN4(n11227), 
        .QN(n11223) );
  NAND2X0 U11166 ( .IN1(n11228), .IN2(n11229), .QN(n11227) );
  NAND2X0 U11167 ( .IN1(n11230), .IN2(n11231), .QN(n11229) );
  NAND2X0 U11168 ( .IN1(n11232), .IN2(n11233), .QN(n11231) );
  INVX0 U11169 ( .INP(n11234), .ZN(n11233) );
  NAND2X0 U11170 ( .IN1(n11235), .IN2(n11236), .QN(n11230) );
  NAND3X0 U11171 ( .IN1(n11237), .IN2(n11238), .IN3(n11239), .QN(n11226) );
  NAND2X0 U11172 ( .IN1(n11234), .IN2(n11240), .QN(n11238) );
  NAND2X0 U11173 ( .IN1(n11236), .IN2(n11241), .QN(n11240) );
  NAND2X0 U11174 ( .IN1(n11242), .IN2(n11243), .QN(n11236) );
  NAND2X0 U11175 ( .IN1(n11244), .IN2(n11245), .QN(n11243) );
  NOR2X0 U11176 ( .IN1(n11246), .IN2(n11247), .QN(n11234) );
  NOR2X0 U11177 ( .IN1(n11248), .IN2(n11245), .QN(n11247) );
  NOR2X0 U11178 ( .IN1(n11242), .IN2(n11249), .QN(n11246) );
  NAND2X0 U11179 ( .IN1(n11249), .IN2(n11250), .QN(n11225) );
  NAND2X0 U11180 ( .IN1(n11251), .IN2(n11252), .QN(n11250) );
  NAND3X0 U11181 ( .IN1(n11253), .IN2(n11254), .IN3(n11255), .QN(n11252) );
  NAND2X0 U11182 ( .IN1(n11256), .IN2(n11257), .QN(n11251) );
  NAND2X0 U11183 ( .IN1(n11241), .IN2(n11258), .QN(n11256) );
  NAND2X0 U11184 ( .IN1(n11259), .IN2(n11239), .QN(n11258) );
  NAND3X0 U11185 ( .IN1(n11260), .IN2(n11248), .IN3(n11245), .QN(n11224) );
  NAND2X0 U11186 ( .IN1(n11261), .IN2(n11262), .QN(n11260) );
  NAND2X0 U11187 ( .IN1(n11242), .IN2(n11263), .QN(n11262) );
  NAND2X0 U11188 ( .IN1(n11241), .IN2(n11264), .QN(n11263) );
  NAND2X0 U11189 ( .IN1(n11255), .IN2(n11254), .QN(n11261) );
  NAND2X0 U11190 ( .IN1(n11265), .IN2(n11212), .QN(n11222) );
  INVX0 U11191 ( .INP(n11266), .ZN(n11212) );
  NAND3X0 U11192 ( .IN1(n11267), .IN2(n11268), .IN3(n11269), .QN(n11266) );
  NAND2X0 U11193 ( .IN1(n11270), .IN2(n11239), .QN(n11269) );
  NAND2X0 U11194 ( .IN1(n11271), .IN2(n11272), .QN(n11270) );
  NAND2X0 U11195 ( .IN1(n11235), .IN2(n11253), .QN(n11272) );
  INVX0 U11196 ( .INP(n11259), .ZN(n11235) );
  NAND2X0 U11197 ( .IN1(n11249), .IN2(n11273), .QN(n11271) );
  NAND3X0 U11198 ( .IN1(n11274), .IN2(n11275), .IN3(n11276), .QN(n11273) );
  NAND2X0 U11199 ( .IN1(n11255), .IN2(n11248), .QN(n11276) );
  NAND2X0 U11200 ( .IN1(n11277), .IN2(n11278), .QN(n11275) );
  NAND2X0 U11201 ( .IN1(n11279), .IN2(n11232), .QN(n11274) );
  NAND3X0 U11202 ( .IN1(n11280), .IN2(n11248), .IN3(n11237), .QN(n11268) );
  NAND2X0 U11203 ( .IN1(n11281), .IN2(n11282), .QN(n11280) );
  NAND2X0 U11204 ( .IN1(n11228), .IN2(n11241), .QN(n11282) );
  NAND2X0 U11205 ( .IN1(n11249), .IN2(n11242), .QN(n11281) );
  INVX0 U11206 ( .INP(n11245), .ZN(n11249) );
  NAND2X0 U11207 ( .IN1(n11283), .IN2(n11245), .QN(n11267) );
  NAND3X0 U11208 ( .IN1(n11284), .IN2(n11285), .IN3(n11286), .QN(n11245) );
  NAND2X0 U11209 ( .IN1(g5648), .IN2(g351), .QN(n11286) );
  NAND2X0 U11210 ( .IN1(g5629), .IN2(g349), .QN(n11285) );
  NAND2X0 U11211 ( .IN1(g337), .IN2(g353), .QN(n11284) );
  NAND2X0 U11212 ( .IN1(n11287), .IN2(n11288), .QN(n11283) );
  NAND2X0 U11213 ( .IN1(n11232), .IN2(n11257), .QN(n11288) );
  NOR2X0 U11214 ( .IN1(n11255), .IN2(n11237), .QN(n11232) );
  NAND2X0 U11215 ( .IN1(n11228), .IN2(n11289), .QN(n11287) );
  NAND3X0 U11216 ( .IN1(n11290), .IN2(n11291), .IN3(n11292), .QN(n11289) );
  NAND2X0 U11217 ( .IN1(n11279), .IN2(n11255), .QN(n11292) );
  INVX0 U11218 ( .INP(n11241), .ZN(n11255) );
  NAND3X0 U11219 ( .IN1(n11293), .IN2(n11294), .IN3(n11295), .QN(n11241) );
  NAND2X0 U11220 ( .IN1(g5648), .IN2(g381), .QN(n11295) );
  NAND2X0 U11221 ( .IN1(g5629), .IN2(g379), .QN(n11294) );
  NAND2X0 U11222 ( .IN1(g337), .IN2(g383), .QN(n11293) );
  NAND2X0 U11223 ( .IN1(n11253), .IN2(n11277), .QN(n11291) );
  INVX0 U11224 ( .INP(n11264), .ZN(n11277) );
  NAND2X0 U11225 ( .IN1(n11259), .IN2(n11254), .QN(n11264) );
  NAND3X0 U11226 ( .IN1(n11296), .IN2(n11297), .IN3(n11298), .QN(n11259) );
  NAND2X0 U11227 ( .IN1(g5648), .IN2(g396), .QN(n11298) );
  NAND2X0 U11228 ( .IN1(g5629), .IN2(g394), .QN(n11297) );
  NAND2X0 U11229 ( .IN1(g337), .IN2(g324), .QN(n11296) );
  NAND2X0 U11230 ( .IN1(n11237), .IN2(n11278), .QN(n11290) );
  INVX0 U11231 ( .INP(n11254), .ZN(n11237) );
  NAND3X0 U11232 ( .IN1(n11299), .IN2(n11300), .IN3(n11301), .QN(n11254) );
  NAND2X0 U11233 ( .IN1(g5648), .IN2(g366), .QN(n11301) );
  NAND2X0 U11234 ( .IN1(g5629), .IN2(g364), .QN(n11300) );
  NAND2X0 U11235 ( .IN1(g337), .IN2(g368), .QN(n11299) );
  INVX0 U11236 ( .INP(n11302), .ZN(n11265) );
  NAND2X0 U11237 ( .IN1(n11215), .IN2(n11302), .QN(n11211) );
  NAND2X0 U11238 ( .IN1(n4298), .IN2(g605), .QN(n11218) );
  NOR2X0 U11239 ( .IN1(n11303), .IN2(n11304), .QN(g28328) );
  XNOR2X1 U11240 ( .IN1(n4415), .IN2(n11305), .Q(n11304) );
  NAND2X0 U11241 ( .IN1(n11306), .IN2(g2760), .QN(n11305) );
  NOR2X0 U11242 ( .IN1(n9305), .IN2(n11307), .QN(g28325) );
  XOR2X1 U11243 ( .IN1(n4416), .IN2(n11308), .Q(n11307) );
  NOR2X0 U11244 ( .IN1(n8512), .IN2(n11309), .QN(g28321) );
  XNOR2X1 U11245 ( .IN1(n4417), .IN2(n11310), .Q(n11309) );
  NAND2X0 U11246 ( .IN1(n11311), .IN2(g1372), .QN(n11310) );
  NOR2X0 U11247 ( .IN1(n8536), .IN2(n11312), .QN(g28199) );
  XOR2X1 U11248 ( .IN1(n4396), .IN2(n10868), .Q(n11312) );
  NOR2X0 U11249 ( .IN1(n10265), .IN2(n11313), .QN(g28148) );
  XOR2X1 U11250 ( .IN1(n8069), .IN2(n3424), .Q(n11313) );
  NOR2X0 U11251 ( .IN1(n10267), .IN2(n11314), .QN(g28147) );
  XOR2X1 U11252 ( .IN1(n8068), .IN2(n3427), .Q(n11314) );
  NOR2X0 U11253 ( .IN1(n10269), .IN2(n11315), .QN(g28146) );
  XOR2X1 U11254 ( .IN1(n8064), .IN2(n3430), .Q(n11315) );
  NOR2X0 U11255 ( .IN1(n10271), .IN2(n11316), .QN(g28145) );
  XOR2X1 U11256 ( .IN1(n8067), .IN2(n3433), .Q(n11316) );
  NAND2X0 U11257 ( .IN1(n11317), .IN2(n11318), .QN(g27771) );
  NAND2X0 U11258 ( .IN1(test_so81), .IN2(n11319), .QN(n11318) );
  NAND2X0 U11259 ( .IN1(n11320), .IN2(n10028), .QN(n11319) );
  NAND2X0 U11260 ( .IN1(n11321), .IN2(n10028), .QN(n11317) );
  NAND2X0 U11261 ( .IN1(n11322), .IN2(n11323), .QN(g27769) );
  NAND2X0 U11262 ( .IN1(n11324), .IN2(g2524), .QN(n11323) );
  NAND2X0 U11263 ( .IN1(n11320), .IN2(n10027), .QN(n11324) );
  NAND2X0 U11264 ( .IN1(n11321), .IN2(n10027), .QN(n11322) );
  NAND2X0 U11265 ( .IN1(n11325), .IN2(n11326), .QN(g27768) );
  NAND2X0 U11266 ( .IN1(n11327), .IN2(g1828), .QN(n11326) );
  NAND2X0 U11267 ( .IN1(n11328), .IN2(n10075), .QN(n11327) );
  NAND2X0 U11268 ( .IN1(n11329), .IN2(n10075), .QN(n11325) );
  NAND2X0 U11269 ( .IN1(n11330), .IN2(n11331), .QN(g27767) );
  NAND2X0 U11270 ( .IN1(n11332), .IN2(g2523), .QN(n11331) );
  NAND2X0 U11271 ( .IN1(n11320), .IN2(n10029), .QN(n11332) );
  NOR2X0 U11272 ( .IN1(n11333), .IN2(n11334), .QN(n11320) );
  NAND2X0 U11273 ( .IN1(n11321), .IN2(n10029), .QN(n11330) );
  INVX0 U11274 ( .INP(n11335), .ZN(n11321) );
  NAND4X0 U11275 ( .IN1(test_so79), .IN2(n11336), .IN3(n11337), .IN4(n11338), 
        .QN(n11335) );
  NAND2X0 U11276 ( .IN1(n9164), .IN2(n11339), .QN(n11338) );
  NAND2X0 U11277 ( .IN1(n9163), .IN2(n11340), .QN(n11337) );
  NAND2X0 U11278 ( .IN1(n9165), .IN2(n11341), .QN(n11336) );
  NAND2X0 U11279 ( .IN1(n11342), .IN2(n11343), .QN(g27766) );
  NAND2X0 U11280 ( .IN1(n11344), .IN2(g1830), .QN(n11343) );
  NAND2X0 U11281 ( .IN1(n11328), .IN2(n10074), .QN(n11344) );
  NAND2X0 U11282 ( .IN1(n11329), .IN2(n10074), .QN(n11342) );
  NAND2X0 U11283 ( .IN1(n11345), .IN2(n11346), .QN(g27765) );
  NAND2X0 U11284 ( .IN1(n11347), .IN2(g1134), .QN(n11346) );
  NAND2X0 U11285 ( .IN1(n11348), .IN2(g1088), .QN(n11347) );
  NAND2X0 U11286 ( .IN1(n11349), .IN2(g1088), .QN(n11345) );
  NAND2X0 U11287 ( .IN1(n11350), .IN2(n11351), .QN(g27764) );
  NAND2X0 U11288 ( .IN1(n11352), .IN2(g1829), .QN(n11351) );
  NAND2X0 U11289 ( .IN1(n11328), .IN2(n10076), .QN(n11352) );
  NOR2X0 U11290 ( .IN1(n11353), .IN2(n11354), .QN(n11328) );
  NAND2X0 U11291 ( .IN1(n11329), .IN2(n10076), .QN(n11350) );
  INVX0 U11292 ( .INP(n11355), .ZN(n11329) );
  NAND4X0 U11293 ( .IN1(n11356), .IN2(g1690), .IN3(n11357), .IN4(n11358), .QN(
        n11355) );
  NAND2X0 U11294 ( .IN1(n9161), .IN2(n11359), .QN(n11358) );
  NAND2X0 U11295 ( .IN1(n9160), .IN2(n11360), .QN(n11357) );
  NAND2X0 U11296 ( .IN1(n9162), .IN2(n11361), .QN(n11356) );
  NAND2X0 U11297 ( .IN1(n11362), .IN2(n11363), .QN(g27763) );
  NAND2X0 U11298 ( .IN1(n11364), .IN2(g1136), .QN(n11363) );
  NAND2X0 U11299 ( .IN1(n11348), .IN2(g6712), .QN(n11364) );
  NAND2X0 U11300 ( .IN1(n11349), .IN2(g6712), .QN(n11362) );
  NAND2X0 U11301 ( .IN1(n11365), .IN2(n11366), .QN(g27762) );
  NAND2X0 U11302 ( .IN1(n11367), .IN2(g447), .QN(n11366) );
  NAND2X0 U11303 ( .IN1(n11368), .IN2(n10160), .QN(n11367) );
  NAND2X0 U11304 ( .IN1(n11369), .IN2(n10160), .QN(n11365) );
  NAND2X0 U11305 ( .IN1(n11370), .IN2(n11371), .QN(g27761) );
  NAND2X0 U11306 ( .IN1(n11372), .IN2(g1135), .QN(n11371) );
  NAND2X0 U11307 ( .IN1(n11348), .IN2(g5472), .QN(n11372) );
  NOR2X0 U11308 ( .IN1(n11373), .IN2(n11374), .QN(n11348) );
  NAND2X0 U11309 ( .IN1(n11349), .IN2(g5472), .QN(n11370) );
  INVX0 U11310 ( .INP(n11375), .ZN(n11349) );
  NAND4X0 U11311 ( .IN1(n11376), .IN2(g996), .IN3(n11377), .IN4(n11378), .QN(
        n11375) );
  NAND2X0 U11312 ( .IN1(n9158), .IN2(n11379), .QN(n11378) );
  NAND2X0 U11313 ( .IN1(n9157), .IN2(n11380), .QN(n11377) );
  NAND2X0 U11314 ( .IN1(n9159), .IN2(n11381), .QN(n11376) );
  NAND2X0 U11315 ( .IN1(n11382), .IN2(n11383), .QN(g27760) );
  NAND2X0 U11316 ( .IN1(n11384), .IN2(g449), .QN(n11383) );
  NAND2X0 U11317 ( .IN1(n11368), .IN2(n10159), .QN(n11384) );
  NAND2X0 U11318 ( .IN1(n11369), .IN2(n10159), .QN(n11382) );
  NAND2X0 U11319 ( .IN1(n11385), .IN2(n11386), .QN(g27759) );
  NAND2X0 U11320 ( .IN1(n11387), .IN2(g448), .QN(n11386) );
  NAND2X0 U11321 ( .IN1(n11368), .IN2(n10158), .QN(n11387) );
  NOR2X0 U11322 ( .IN1(n11388), .IN2(n11389), .QN(n11368) );
  NAND2X0 U11323 ( .IN1(n11369), .IN2(n10158), .QN(n11385) );
  INVX0 U11324 ( .INP(n11390), .ZN(n11369) );
  NAND4X0 U11325 ( .IN1(n11391), .IN2(g309), .IN3(n11392), .IN4(n11393), .QN(
        n11390) );
  NAND2X0 U11326 ( .IN1(n9155), .IN2(n11394), .QN(n11393) );
  NAND2X0 U11327 ( .IN1(n9154), .IN2(n11395), .QN(n11392) );
  NAND2X0 U11328 ( .IN1(n9156), .IN2(n11396), .QN(n11391) );
  NOR2X0 U11329 ( .IN1(n11303), .IN2(n11397), .QN(g27724) );
  XOR2X1 U11330 ( .IN1(n4393), .IN2(n11306), .Q(n11397) );
  NOR3X0 U11331 ( .IN1(n11398), .IN2(n9305), .IN3(n11308), .QN(g27722) );
  INVX0 U11332 ( .INP(n3417), .ZN(n11308) );
  NAND2X0 U11333 ( .IN1(test_so70), .IN2(n11399), .QN(n3417) );
  NOR2X0 U11334 ( .IN1(n11399), .IN2(test_so70), .QN(n11398) );
  NOR2X0 U11335 ( .IN1(n8512), .IN2(n11400), .QN(g27718) );
  XOR2X1 U11336 ( .IN1(n4395), .IN2(n11311), .Q(n11400) );
  NOR3X0 U11337 ( .IN1(n11401), .IN2(n9305), .IN3(n11399), .QN(g27682) );
  NOR3X0 U11338 ( .IN1(n4468), .IN2(n4473), .IN3(n11402), .QN(n11399) );
  NOR2X0 U11339 ( .IN1(n11403), .IN2(g2059), .QN(n11401) );
  NOR2X0 U11340 ( .IN1(n4468), .IN2(n11402), .QN(n11403) );
  INVX0 U11341 ( .INP(n9306), .ZN(n11402) );
  NOR3X0 U11342 ( .IN1(n11404), .IN2(n8512), .IN3(n11311), .QN(g27678) );
  NOR3X0 U11343 ( .IN1(n4469), .IN2(n4475), .IN3(n8508), .QN(n11311) );
  NOR2X0 U11344 ( .IN1(n11405), .IN2(g1365), .QN(n11404) );
  NOR2X0 U11345 ( .IN1(n4469), .IN2(n8508), .QN(n11405) );
  NOR3X0 U11346 ( .IN1(n11406), .IN2(n8536), .IN3(n10868), .QN(g27672) );
  NOR3X0 U11347 ( .IN1(n8528), .IN2(n4477), .IN3(n8074), .QN(n10868) );
  NOR2X0 U11348 ( .IN1(n11407), .IN2(g679), .QN(n11406) );
  NOR2X0 U11349 ( .IN1(n8528), .IN2(n8074), .QN(n11407) );
  NOR2X0 U11350 ( .IN1(n10265), .IN2(n11408), .QN(g27621) );
  XOR2X1 U11351 ( .IN1(n11409), .IN2(n7688), .Q(n11408) );
  NOR2X0 U11352 ( .IN1(n10267), .IN2(n11410), .QN(g27612) );
  XOR2X1 U11353 ( .IN1(n11411), .IN2(n7692), .Q(n11410) );
  NOR2X0 U11354 ( .IN1(n10269), .IN2(n11412), .QN(g27603) );
  XNOR2X1 U11355 ( .IN1(n7696), .IN2(n3431), .Q(n11412) );
  NAND2X0 U11356 ( .IN1(n3689), .IN2(g767), .QN(n3431) );
  NOR2X0 U11357 ( .IN1(n10271), .IN2(n11413), .QN(g27594) );
  XOR2X1 U11358 ( .IN1(n11414), .IN2(n7700), .Q(n11413) );
  NAND4X0 U11359 ( .IN1(n11415), .IN2(n11416), .IN3(n3700), .IN4(n11417), .QN(
        g27380) );
  NOR4X0 U11360 ( .IN1(n11418), .IN2(n11419), .IN3(n11420), .IN4(n11421), .QN(
        n11417) );
  NOR2X0 U11361 ( .IN1(n4424), .IN2(n11422), .QN(n11421) );
  NOR2X0 U11362 ( .IN1(n11423), .IN2(n11424), .QN(n11420) );
  NOR2X0 U11363 ( .IN1(n11425), .IN2(n3705), .QN(n11423) );
  NOR3X0 U11364 ( .IN1(g185), .IN2(n4405), .IN3(n11426), .QN(n11425) );
  NOR4X0 U11365 ( .IN1(n11427), .IN2(n11428), .IN3(n11426), .IN4(n11429), .QN(
        n11419) );
  NOR2X0 U11366 ( .IN1(n14351), .IN2(n11430), .QN(n11428) );
  NOR2X0 U11367 ( .IN1(n14349), .IN2(n11431), .QN(n11427) );
  INVX0 U11368 ( .INP(n11432), .ZN(n11416) );
  NOR2X0 U11369 ( .IN1(n11433), .IN2(n14352), .QN(n11432) );
  NAND2X0 U11370 ( .IN1(n7430), .IN2(n11434), .QN(n11415) );
  NAND2X0 U11371 ( .IN1(n11435), .IN2(n11436), .QN(g27354) );
  INVX0 U11372 ( .INP(n11437), .ZN(n11436) );
  NOR2X0 U11373 ( .IN1(n11438), .IN2(n7350), .QN(n11437) );
  NAND2X0 U11374 ( .IN1(n11438), .IN2(n11439), .QN(n11435) );
  NAND2X0 U11375 ( .IN1(n11440), .IN2(n11441), .QN(g27348) );
  NAND2X0 U11376 ( .IN1(n11442), .IN2(g2660), .QN(n11441) );
  NAND2X0 U11377 ( .IN1(n11443), .IN2(n11439), .QN(n11440) );
  NAND2X0 U11378 ( .IN1(n11444), .IN2(n11445), .QN(g27347) );
  INVX0 U11379 ( .INP(n11446), .ZN(n11445) );
  NOR2X0 U11380 ( .IN1(n11438), .IN2(n7166), .QN(n11446) );
  NAND2X0 U11381 ( .IN1(n11438), .IN2(n11447), .QN(n11444) );
  NAND2X0 U11382 ( .IN1(n11448), .IN2(n11449), .QN(g27346) );
  INVX0 U11383 ( .INP(n11450), .ZN(n11449) );
  NOR2X0 U11384 ( .IN1(n11451), .IN2(n7352), .QN(n11450) );
  NAND2X0 U11385 ( .IN1(n11451), .IN2(n11452), .QN(n11448) );
  NAND2X0 U11386 ( .IN1(n11453), .IN2(n11454), .QN(g27345) );
  INVX0 U11387 ( .INP(n11455), .ZN(n11454) );
  NOR2X0 U11388 ( .IN1(n11456), .IN2(n7349), .QN(n11455) );
  NAND2X0 U11389 ( .IN1(n11456), .IN2(n11439), .QN(n11453) );
  NAND3X0 U11390 ( .IN1(n10949), .IN2(n10924), .IN3(n11457), .QN(n11439) );
  INVX0 U11391 ( .INP(n10938), .ZN(n10949) );
  NAND2X0 U11392 ( .IN1(n11458), .IN2(n11459), .QN(g27344) );
  NAND2X0 U11393 ( .IN1(test_so89), .IN2(n11442), .QN(n11459) );
  NAND2X0 U11394 ( .IN1(n11443), .IN2(n11447), .QN(n11458) );
  NAND2X0 U11395 ( .IN1(n11460), .IN2(n11461), .QN(g27343) );
  INVX0 U11396 ( .INP(n11462), .ZN(n11461) );
  NOR2X0 U11397 ( .IN1(n11438), .IN2(n7339), .QN(n11462) );
  NAND2X0 U11398 ( .IN1(n11438), .IN2(n11463), .QN(n11460) );
  NAND2X0 U11399 ( .IN1(n11464), .IN2(n11465), .QN(g27342) );
  INVX0 U11400 ( .INP(n11466), .ZN(n11465) );
  NOR2X0 U11401 ( .IN1(n11467), .IN2(n7632), .QN(n11466) );
  NAND2X0 U11402 ( .IN1(n11467), .IN2(n11468), .QN(n11464) );
  NAND2X0 U11403 ( .IN1(n11469), .IN2(n11470), .QN(g27341) );
  INVX0 U11404 ( .INP(n11471), .ZN(n11470) );
  NOR2X0 U11405 ( .IN1(n11472), .IN2(n7353), .QN(n11471) );
  NAND2X0 U11406 ( .IN1(n11472), .IN2(n11452), .QN(n11469) );
  NAND2X0 U11407 ( .IN1(n11473), .IN2(n11474), .QN(g27340) );
  INVX0 U11408 ( .INP(n11475), .ZN(n11474) );
  NOR2X0 U11409 ( .IN1(n11451), .IN2(n7168), .QN(n11475) );
  NAND2X0 U11410 ( .IN1(n11451), .IN2(n11476), .QN(n11473) );
  NAND2X0 U11411 ( .IN1(n11477), .IN2(n11478), .QN(g27339) );
  NAND2X0 U11412 ( .IN1(n11479), .IN2(g1270), .QN(n11478) );
  NAND2X0 U11413 ( .IN1(n11480), .IN2(n11481), .QN(n11477) );
  NAND2X0 U11414 ( .IN1(n11482), .IN2(n11483), .QN(g27338) );
  INVX0 U11415 ( .INP(n11484), .ZN(n11483) );
  NOR2X0 U11416 ( .IN1(n11456), .IN2(n7165), .QN(n11484) );
  NAND2X0 U11417 ( .IN1(n11456), .IN2(n11447), .QN(n11482) );
  INVX0 U11418 ( .INP(n11485), .ZN(n11447) );
  NAND2X0 U11419 ( .IN1(n11486), .IN2(n11487), .QN(n11485) );
  NAND2X0 U11420 ( .IN1(n11488), .IN2(n10974), .QN(n11487) );
  NAND2X0 U11421 ( .IN1(n11457), .IN2(n10938), .QN(n11486) );
  INVX0 U11422 ( .INP(n11488), .ZN(n11457) );
  NAND2X0 U11423 ( .IN1(n11489), .IN2(n11490), .QN(g27337) );
  NAND2X0 U11424 ( .IN1(n11442), .IN2(g2654), .QN(n11490) );
  NAND2X0 U11425 ( .IN1(n11443), .IN2(n11463), .QN(n11489) );
  NAND2X0 U11426 ( .IN1(n11491), .IN2(n11492), .QN(g27336) );
  INVX0 U11427 ( .INP(n11493), .ZN(n11492) );
  NOR2X0 U11428 ( .IN1(n11438), .IN2(n7327), .QN(n11493) );
  NAND2X0 U11429 ( .IN1(n11438), .IN2(n11494), .QN(n11491) );
  NOR2X0 U11430 ( .IN1(n11495), .IN2(n4299), .QN(n11438) );
  NAND2X0 U11431 ( .IN1(n11496), .IN2(n11497), .QN(g27335) );
  INVX0 U11432 ( .INP(n11498), .ZN(n11497) );
  NOR2X0 U11433 ( .IN1(n11499), .IN2(n7633), .QN(n11498) );
  NAND2X0 U11434 ( .IN1(n11499), .IN2(n11468), .QN(n11496) );
  NAND2X0 U11435 ( .IN1(n11500), .IN2(n11501), .QN(g27334) );
  INVX0 U11436 ( .INP(n11502), .ZN(n11501) );
  NOR2X0 U11437 ( .IN1(n11467), .IN2(n7372), .QN(n11502) );
  NAND2X0 U11438 ( .IN1(n11467), .IN2(n11503), .QN(n11500) );
  NAND2X0 U11439 ( .IN1(n11504), .IN2(n11505), .QN(g27333) );
  NAND2X0 U11440 ( .IN1(n11506), .IN2(n11452), .QN(n11505) );
  NAND2X0 U11441 ( .IN1(n11507), .IN2(n11052), .QN(n11452) );
  NOR2X0 U11442 ( .IN1(n11047), .IN2(n11077), .QN(n11052) );
  INVX0 U11443 ( .INP(n11508), .ZN(n11504) );
  NOR2X0 U11444 ( .IN1(n8092), .IN2(n11506), .QN(n11508) );
  NAND2X0 U11445 ( .IN1(n11509), .IN2(n11510), .QN(g27332) );
  INVX0 U11446 ( .INP(n11511), .ZN(n11510) );
  NOR2X0 U11447 ( .IN1(n11472), .IN2(n7169), .QN(n11511) );
  NAND2X0 U11448 ( .IN1(n11472), .IN2(n11476), .QN(n11509) );
  NAND2X0 U11449 ( .IN1(n11512), .IN2(n11513), .QN(g27331) );
  INVX0 U11450 ( .INP(n11514), .ZN(n11513) );
  NOR2X0 U11451 ( .IN1(n11451), .IN2(n7342), .QN(n11514) );
  NAND2X0 U11452 ( .IN1(n11451), .IN2(n11515), .QN(n11512) );
  NAND2X0 U11453 ( .IN1(n11516), .IN2(n11517), .QN(g27330) );
  INVX0 U11454 ( .INP(n11518), .ZN(n11517) );
  NOR2X0 U11455 ( .IN1(n11519), .IN2(n7635), .QN(n11518) );
  NAND2X0 U11456 ( .IN1(n11519), .IN2(n11520), .QN(n11516) );
  NAND2X0 U11457 ( .IN1(n11521), .IN2(n11522), .QN(g27329) );
  NAND2X0 U11458 ( .IN1(n11523), .IN2(n11481), .QN(n11522) );
  INVX0 U11459 ( .INP(n11524), .ZN(n11521) );
  NOR2X0 U11460 ( .IN1(n11523), .IN2(n7356), .QN(n11524) );
  NAND2X0 U11461 ( .IN1(n11525), .IN2(n11526), .QN(g27328) );
  NAND2X0 U11462 ( .IN1(test_so46), .IN2(n11479), .QN(n11526) );
  NAND2X0 U11463 ( .IN1(n11480), .IN2(n11527), .QN(n11525) );
  NAND2X0 U11464 ( .IN1(n11528), .IN2(n11529), .QN(g27327) );
  INVX0 U11465 ( .INP(n11530), .ZN(n11529) );
  NOR2X0 U11466 ( .IN1(n11531), .IN2(n7358), .QN(n11530) );
  NAND2X0 U11467 ( .IN1(n11531), .IN2(n11532), .QN(n11528) );
  NAND2X0 U11468 ( .IN1(n11533), .IN2(n11534), .QN(g27326) );
  INVX0 U11469 ( .INP(n11535), .ZN(n11534) );
  NOR2X0 U11470 ( .IN1(n11456), .IN2(n7338), .QN(n11535) );
  NAND2X0 U11471 ( .IN1(n11456), .IN2(n11463), .QN(n11533) );
  INVX0 U11472 ( .INP(n11536), .ZN(n11463) );
  NAND2X0 U11473 ( .IN1(n11537), .IN2(n11538), .QN(n11536) );
  NAND2X0 U11474 ( .IN1(n11488), .IN2(n10944), .QN(n11537) );
  XNOR2X1 U11475 ( .IN1(n8785), .IN2(n10928), .Q(n11488) );
  NAND2X0 U11476 ( .IN1(n11539), .IN2(n11540), .QN(g27325) );
  NAND2X0 U11477 ( .IN1(n11442), .IN2(g2651), .QN(n11540) );
  INVX0 U11478 ( .INP(n11443), .ZN(n11442) );
  NAND2X0 U11479 ( .IN1(n11443), .IN2(n11494), .QN(n11539) );
  NOR2X0 U11480 ( .IN1(n11495), .IN2(n4370), .QN(n11443) );
  NAND2X0 U11481 ( .IN1(n11541), .IN2(n11542), .QN(g27324) );
  INVX0 U11482 ( .INP(n11543), .ZN(n11542) );
  NOR2X0 U11483 ( .IN1(n11544), .IN2(n7634), .QN(n11543) );
  NAND2X0 U11484 ( .IN1(n11544), .IN2(n11468), .QN(n11541) );
  NAND3X0 U11485 ( .IN1(n11545), .IN2(n11546), .IN3(n11547), .QN(n11468) );
  NAND2X0 U11486 ( .IN1(n11548), .IN2(n11549), .QN(g27323) );
  INVX0 U11487 ( .INP(n11550), .ZN(n11549) );
  NOR2X0 U11488 ( .IN1(n11499), .IN2(n7373), .QN(n11550) );
  NAND2X0 U11489 ( .IN1(n11499), .IN2(n11503), .QN(n11548) );
  NAND2X0 U11490 ( .IN1(n11551), .IN2(n11552), .QN(g27322) );
  INVX0 U11491 ( .INP(n11553), .ZN(n11552) );
  NOR2X0 U11492 ( .IN1(n11467), .IN2(n7620), .QN(n11553) );
  NAND2X0 U11493 ( .IN1(n11554), .IN2(n11467), .QN(n11551) );
  NAND2X0 U11494 ( .IN1(n11555), .IN2(n11556), .QN(g27321) );
  INVX0 U11495 ( .INP(n11557), .ZN(n11556) );
  NOR2X0 U11496 ( .IN1(n11506), .IN2(n7167), .QN(n11557) );
  NAND2X0 U11497 ( .IN1(n11506), .IN2(n11476), .QN(n11555) );
  INVX0 U11498 ( .INP(n11558), .ZN(n11476) );
  NAND2X0 U11499 ( .IN1(n11559), .IN2(n11560), .QN(n11558) );
  NAND2X0 U11500 ( .IN1(n11561), .IN2(n11078), .QN(n11560) );
  NAND2X0 U11501 ( .IN1(n11507), .IN2(n11047), .QN(n11559) );
  INVX0 U11502 ( .INP(n11561), .ZN(n11507) );
  NAND2X0 U11503 ( .IN1(n11562), .IN2(n11563), .QN(g27320) );
  INVX0 U11504 ( .INP(n11564), .ZN(n11563) );
  NOR2X0 U11505 ( .IN1(n11472), .IN2(n7343), .QN(n11564) );
  NAND2X0 U11506 ( .IN1(n11472), .IN2(n11515), .QN(n11562) );
  NAND2X0 U11507 ( .IN1(n11565), .IN2(n11566), .QN(g27319) );
  INVX0 U11508 ( .INP(n11567), .ZN(n11566) );
  NOR2X0 U11509 ( .IN1(n11451), .IN2(n7330), .QN(n11567) );
  NAND2X0 U11510 ( .IN1(n11451), .IN2(n11568), .QN(n11565) );
  NOR2X0 U11511 ( .IN1(n11569), .IN2(n4366), .QN(n11451) );
  NAND2X0 U11512 ( .IN1(n11570), .IN2(n11571), .QN(g27318) );
  NAND2X0 U11513 ( .IN1(n11572), .IN2(n11520), .QN(n11571) );
  NAND2X0 U11514 ( .IN1(test_so58), .IN2(n11573), .QN(n11570) );
  NAND2X0 U11515 ( .IN1(n11574), .IN2(n11575), .QN(g27317) );
  INVX0 U11516 ( .INP(n11576), .ZN(n11575) );
  NOR2X0 U11517 ( .IN1(n11519), .IN2(n7375), .QN(n11576) );
  NAND2X0 U11518 ( .IN1(n11519), .IN2(n11577), .QN(n11574) );
  NAND2X0 U11519 ( .IN1(n11578), .IN2(n11579), .QN(g27316) );
  NAND2X0 U11520 ( .IN1(n11580), .IN2(n11481), .QN(n11579) );
  NAND2X0 U11521 ( .IN1(n11581), .IN2(n11155), .QN(n11481) );
  NOR2X0 U11522 ( .IN1(n11150), .IN2(n11180), .QN(n11155) );
  NAND2X0 U11523 ( .IN1(n11582), .IN2(g1271), .QN(n11578) );
  NAND2X0 U11524 ( .IN1(n11583), .IN2(n11584), .QN(g27315) );
  INVX0 U11525 ( .INP(n11585), .ZN(n11584) );
  NOR2X0 U11526 ( .IN1(n11523), .IN2(n7171), .QN(n11585) );
  NAND2X0 U11527 ( .IN1(n11523), .IN2(n11527), .QN(n11583) );
  NAND2X0 U11528 ( .IN1(n11586), .IN2(n11587), .QN(g27314) );
  NAND2X0 U11529 ( .IN1(n11479), .IN2(g1264), .QN(n11587) );
  NAND2X0 U11530 ( .IN1(n11480), .IN2(n11588), .QN(n11586) );
  NAND2X0 U11531 ( .IN1(n11589), .IN2(n11590), .QN(g27313) );
  INVX0 U11532 ( .INP(n11591), .ZN(n11590) );
  NOR2X0 U11533 ( .IN1(n11592), .IN2(n7637), .QN(n11591) );
  NAND2X0 U11534 ( .IN1(n11592), .IN2(n11593), .QN(n11589) );
  NAND2X0 U11535 ( .IN1(n11594), .IN2(n11595), .QN(g27312) );
  NAND2X0 U11536 ( .IN1(n11596), .IN2(n11532), .QN(n11595) );
  NAND2X0 U11537 ( .IN1(n11597), .IN2(g586), .QN(n11594) );
  NAND2X0 U11538 ( .IN1(n11598), .IN2(n11599), .QN(g27311) );
  INVX0 U11539 ( .INP(n11600), .ZN(n11599) );
  NOR2X0 U11540 ( .IN1(n11531), .IN2(n7173), .QN(n11600) );
  NAND2X0 U11541 ( .IN1(n11531), .IN2(n11601), .QN(n11598) );
  NAND2X0 U11542 ( .IN1(n11602), .IN2(n11603), .QN(g27310) );
  INVX0 U11543 ( .INP(n11604), .ZN(n11603) );
  NOR2X0 U11544 ( .IN1(n11456), .IN2(n7326), .QN(n11604) );
  NAND2X0 U11545 ( .IN1(n11456), .IN2(n11494), .QN(n11602) );
  NOR2X0 U11546 ( .IN1(n11605), .IN2(n11606), .QN(n11494) );
  NOR2X0 U11547 ( .IN1(n11607), .IN2(g3229), .QN(n11606) );
  INVX0 U11548 ( .INP(n11608), .ZN(n11607) );
  NAND2X0 U11549 ( .IN1(n11538), .IN2(n11609), .QN(n11608) );
  NAND2X0 U11550 ( .IN1(n10926), .IN2(n10931), .QN(n11609) );
  INVX0 U11551 ( .INP(n10958), .ZN(n10926) );
  NAND2X0 U11552 ( .IN1(n10924), .IN2(n10938), .QN(n11538) );
  INVX0 U11553 ( .INP(n10944), .ZN(n10924) );
  NOR2X0 U11554 ( .IN1(n8785), .IN2(n11610), .QN(n11605) );
  NOR2X0 U11555 ( .IN1(n10958), .IN2(n11611), .QN(n11610) );
  NOR2X0 U11556 ( .IN1(n10928), .IN2(n11612), .QN(n11611) );
  NOR2X0 U11557 ( .IN1(n10944), .IN2(n10974), .QN(n11612) );
  NOR2X0 U11558 ( .IN1(n10938), .IN2(n10958), .QN(n10974) );
  NAND3X0 U11559 ( .IN1(n11613), .IN2(n11614), .IN3(n11615), .QN(n10938) );
  NAND2X0 U11560 ( .IN1(n7340), .IN2(g7390), .QN(n11615) );
  NAND2X0 U11561 ( .IN1(n7339), .IN2(g2624), .QN(n11614) );
  NAND2X0 U11562 ( .IN1(n7338), .IN2(n10166), .QN(n11613) );
  NAND3X0 U11563 ( .IN1(n11616), .IN2(n11617), .IN3(n11618), .QN(n10944) );
  NAND2X0 U11564 ( .IN1(g7390), .IN2(n8107), .QN(n11618) );
  NAND2X0 U11565 ( .IN1(n7166), .IN2(g2624), .QN(n11617) );
  NAND2X0 U11566 ( .IN1(n7165), .IN2(n10166), .QN(n11616) );
  INVX0 U11567 ( .INP(n10931), .ZN(n10928) );
  NAND3X0 U11568 ( .IN1(n11619), .IN2(n11620), .IN3(n11621), .QN(n10931) );
  NAND2X0 U11569 ( .IN1(n7328), .IN2(g7390), .QN(n11621) );
  NAND2X0 U11570 ( .IN1(n7327), .IN2(g2624), .QN(n11620) );
  NAND2X0 U11571 ( .IN1(n7326), .IN2(n10166), .QN(n11619) );
  NAND3X0 U11572 ( .IN1(n11622), .IN2(n11623), .IN3(n11624), .QN(n10958) );
  NAND2X0 U11573 ( .IN1(n7351), .IN2(g7390), .QN(n11624) );
  NAND2X0 U11574 ( .IN1(n7350), .IN2(g2624), .QN(n11623) );
  NAND2X0 U11575 ( .IN1(n7349), .IN2(n10166), .QN(n11622) );
  NOR2X0 U11576 ( .IN1(n10167), .IN2(n11495), .QN(n11456) );
  INVX0 U11577 ( .INP(g22687), .ZN(n11495) );
  INVX0 U11578 ( .INP(g7302), .ZN(n10167) );
  NAND2X0 U11579 ( .IN1(n11625), .IN2(n11626), .QN(g27309) );
  INVX0 U11580 ( .INP(n11627), .ZN(n11626) );
  NOR2X0 U11581 ( .IN1(n11544), .IN2(n7371), .QN(n11627) );
  NAND2X0 U11582 ( .IN1(n11544), .IN2(n11503), .QN(n11625) );
  INVX0 U11583 ( .INP(n11628), .ZN(n11503) );
  NAND2X0 U11584 ( .IN1(n11629), .IN2(n11630), .QN(n11628) );
  NAND2X0 U11585 ( .IN1(n11545), .IN2(n11631), .QN(n11630) );
  NAND3X0 U11586 ( .IN1(n11632), .IN2(n11633), .IN3(n11546), .QN(n11629) );
  NAND2X0 U11587 ( .IN1(n11634), .IN2(n11635), .QN(g27308) );
  INVX0 U11588 ( .INP(n11636), .ZN(n11635) );
  NOR2X0 U11589 ( .IN1(n11499), .IN2(n7621), .QN(n11636) );
  NAND2X0 U11590 ( .IN1(n11554), .IN2(n11499), .QN(n11634) );
  NAND2X0 U11591 ( .IN1(n11637), .IN2(n11638), .QN(g27307) );
  INVX0 U11592 ( .INP(n11639), .ZN(n11638) );
  NOR2X0 U11593 ( .IN1(n11467), .IN2(n7643), .QN(n11639) );
  NAND2X0 U11594 ( .IN1(n11640), .IN2(n11467), .QN(n11637) );
  NOR2X0 U11595 ( .IN1(n11641), .IN2(n4509), .QN(n11467) );
  NAND2X0 U11596 ( .IN1(n11642), .IN2(n11643), .QN(g27306) );
  INVX0 U11597 ( .INP(n11644), .ZN(n11643) );
  NOR2X0 U11598 ( .IN1(n11506), .IN2(n7341), .QN(n11644) );
  NAND2X0 U11599 ( .IN1(n11506), .IN2(n11515), .QN(n11642) );
  INVX0 U11600 ( .INP(n11645), .ZN(n11515) );
  NAND2X0 U11601 ( .IN1(n11646), .IN2(n11647), .QN(n11645) );
  NAND2X0 U11602 ( .IN1(n11561), .IN2(n11077), .QN(n11646) );
  XNOR2X1 U11603 ( .IN1(n8785), .IN2(n11027), .Q(n11561) );
  NAND2X0 U11604 ( .IN1(n11648), .IN2(n11649), .QN(g27305) );
  INVX0 U11605 ( .INP(n11650), .ZN(n11649) );
  NOR2X0 U11606 ( .IN1(n11472), .IN2(n7331), .QN(n11650) );
  NAND2X0 U11607 ( .IN1(n11472), .IN2(n11568), .QN(n11648) );
  NOR2X0 U11608 ( .IN1(n11569), .IN2(n4315), .QN(n11472) );
  NAND2X0 U11609 ( .IN1(n11651), .IN2(n11652), .QN(g27304) );
  NAND2X0 U11610 ( .IN1(n11653), .IN2(n11520), .QN(n11652) );
  NAND3X0 U11611 ( .IN1(n11654), .IN2(n11655), .IN3(n11656), .QN(n11520) );
  INVX0 U11612 ( .INP(n11657), .ZN(n11651) );
  NOR2X0 U11613 ( .IN1(n11653), .IN2(n7636), .QN(n11657) );
  NAND2X0 U11614 ( .IN1(n11658), .IN2(n11659), .QN(g27303) );
  NAND2X0 U11615 ( .IN1(n11573), .IN2(g1754), .QN(n11659) );
  NAND2X0 U11616 ( .IN1(n11572), .IN2(n11577), .QN(n11658) );
  NAND2X0 U11617 ( .IN1(n11660), .IN2(n11661), .QN(g27302) );
  INVX0 U11618 ( .INP(n11662), .ZN(n11661) );
  NOR2X0 U11619 ( .IN1(n11519), .IN2(n7623), .QN(n11662) );
  NAND2X0 U11620 ( .IN1(n11663), .IN2(n11519), .QN(n11660) );
  NAND2X0 U11621 ( .IN1(n11664), .IN2(n11665), .QN(g27301) );
  NAND2X0 U11622 ( .IN1(n11582), .IN2(g1268), .QN(n11665) );
  NAND2X0 U11623 ( .IN1(n11580), .IN2(n11527), .QN(n11664) );
  INVX0 U11624 ( .INP(n11666), .ZN(n11527) );
  NAND2X0 U11625 ( .IN1(n11667), .IN2(n11668), .QN(n11666) );
  NAND2X0 U11626 ( .IN1(n11669), .IN2(n11181), .QN(n11668) );
  NAND2X0 U11627 ( .IN1(n11581), .IN2(n11150), .QN(n11667) );
  INVX0 U11628 ( .INP(n11669), .ZN(n11581) );
  NAND2X0 U11629 ( .IN1(n11670), .IN2(n11671), .QN(g27300) );
  INVX0 U11630 ( .INP(n11672), .ZN(n11671) );
  NOR2X0 U11631 ( .IN1(n11523), .IN2(n7346), .QN(n11672) );
  NAND2X0 U11632 ( .IN1(n11523), .IN2(n11588), .QN(n11670) );
  NAND2X0 U11633 ( .IN1(n11673), .IN2(n11674), .QN(g27299) );
  NAND2X0 U11634 ( .IN1(n11479), .IN2(g1261), .QN(n11674) );
  NAND2X0 U11635 ( .IN1(n11480), .IN2(n11675), .QN(n11673) );
  INVX0 U11636 ( .INP(n11479), .ZN(n11480) );
  NAND2X0 U11637 ( .IN1(g1236), .IN2(g22615), .QN(n11479) );
  NAND2X0 U11638 ( .IN1(n11676), .IN2(n11677), .QN(g27298) );
  INVX0 U11639 ( .INP(n11678), .ZN(n11677) );
  NOR2X0 U11640 ( .IN1(n11679), .IN2(n7638), .QN(n11678) );
  NAND2X0 U11641 ( .IN1(n11679), .IN2(n11593), .QN(n11676) );
  NAND2X0 U11642 ( .IN1(n11680), .IN2(n11681), .QN(g27297) );
  INVX0 U11643 ( .INP(n11682), .ZN(n11681) );
  NOR2X0 U11644 ( .IN1(n11592), .IN2(n7378), .QN(n11682) );
  NAND2X0 U11645 ( .IN1(n11592), .IN2(n11683), .QN(n11680) );
  NAND2X0 U11646 ( .IN1(n11684), .IN2(n11685), .QN(g27296) );
  NAND2X0 U11647 ( .IN1(n11686), .IN2(n11532), .QN(n11685) );
  NAND2X0 U11648 ( .IN1(n11687), .IN2(n11253), .QN(n11532) );
  NOR2X0 U11649 ( .IN1(n11248), .IN2(n11278), .QN(n11253) );
  NAND2X0 U11650 ( .IN1(n11688), .IN2(g585), .QN(n11684) );
  NAND2X0 U11651 ( .IN1(n11689), .IN2(n11690), .QN(g27295) );
  NAND2X0 U11652 ( .IN1(n11597), .IN2(g583), .QN(n11690) );
  NAND2X0 U11653 ( .IN1(n11596), .IN2(n11601), .QN(n11689) );
  NAND2X0 U11654 ( .IN1(n11691), .IN2(n11692), .QN(g27294) );
  INVX0 U11655 ( .INP(n11693), .ZN(n11692) );
  NOR2X0 U11656 ( .IN1(n11531), .IN2(n7348), .QN(n11693) );
  NAND2X0 U11657 ( .IN1(n11531), .IN2(n11694), .QN(n11691) );
  NAND2X0 U11658 ( .IN1(n11695), .IN2(n11696), .QN(g27293) );
  NAND2X0 U11659 ( .IN1(n11697), .IN2(g391), .QN(n11696) );
  NAND2X0 U11660 ( .IN1(n11698), .IN2(n11699), .QN(n11695) );
  NAND2X0 U11661 ( .IN1(n11700), .IN2(n11701), .QN(g27292) );
  INVX0 U11662 ( .INP(n11702), .ZN(n11701) );
  NOR2X0 U11663 ( .IN1(n11544), .IN2(n7622), .QN(n11702) );
  NAND2X0 U11664 ( .IN1(n11554), .IN2(n11544), .QN(n11700) );
  NAND2X0 U11665 ( .IN1(n11703), .IN2(n11704), .QN(n11554) );
  NAND2X0 U11666 ( .IN1(n11547), .IN2(n11546), .QN(n11704) );
  INVX0 U11667 ( .INP(n11631), .ZN(n11546) );
  NAND2X0 U11668 ( .IN1(n11545), .IN2(n11705), .QN(n11703) );
  INVX0 U11669 ( .INP(n11633), .ZN(n11545) );
  XOR2X1 U11670 ( .IN1(n8785), .IN2(n11706), .Q(n11633) );
  NAND2X0 U11671 ( .IN1(n11707), .IN2(n11708), .QN(g27291) );
  INVX0 U11672 ( .INP(n11709), .ZN(n11708) );
  NOR2X0 U11673 ( .IN1(n11499), .IN2(n7644), .QN(n11709) );
  NAND2X0 U11674 ( .IN1(n11640), .IN2(n11499), .QN(n11707) );
  NOR2X0 U11675 ( .IN1(n11641), .IN2(n11710), .QN(n11499) );
  INVX0 U11676 ( .INP(g7264), .ZN(n11710) );
  NAND2X0 U11677 ( .IN1(n11711), .IN2(n11712), .QN(g27290) );
  INVX0 U11678 ( .INP(n11713), .ZN(n11712) );
  NOR2X0 U11679 ( .IN1(n11506), .IN2(n7329), .QN(n11713) );
  NAND2X0 U11680 ( .IN1(n11506), .IN2(n11568), .QN(n11711) );
  NOR2X0 U11681 ( .IN1(n11714), .IN2(n11715), .QN(n11568) );
  NOR2X0 U11682 ( .IN1(n11716), .IN2(g3229), .QN(n11715) );
  INVX0 U11683 ( .INP(n11717), .ZN(n11716) );
  NAND2X0 U11684 ( .IN1(n11647), .IN2(n11718), .QN(n11717) );
  NAND2X0 U11685 ( .IN1(n11043), .IN2(n11038), .QN(n11718) );
  INVX0 U11686 ( .INP(n11056), .ZN(n11043) );
  NAND2X0 U11687 ( .IN1(n11041), .IN2(n11047), .QN(n11647) );
  INVX0 U11688 ( .INP(n11077), .ZN(n11041) );
  NOR2X0 U11689 ( .IN1(n8785), .IN2(n11719), .QN(n11714) );
  NOR2X0 U11690 ( .IN1(n11056), .IN2(n11720), .QN(n11719) );
  NOR2X0 U11691 ( .IN1(n11027), .IN2(n11721), .QN(n11720) );
  NOR2X0 U11692 ( .IN1(n11077), .IN2(n11078), .QN(n11721) );
  NOR2X0 U11693 ( .IN1(n11056), .IN2(n11047), .QN(n11078) );
  NAND3X0 U11694 ( .IN1(n11722), .IN2(n11723), .IN3(n11724), .QN(n11047) );
  NAND2X0 U11695 ( .IN1(n7342), .IN2(g1930), .QN(n11724) );
  NAND2X0 U11696 ( .IN1(n7341), .IN2(n10214), .QN(n11723) );
  NAND2X0 U11697 ( .IN1(n7343), .IN2(g7194), .QN(n11722) );
  NAND3X0 U11698 ( .IN1(n11725), .IN2(n11726), .IN3(n11727), .QN(n11077) );
  NAND2X0 U11699 ( .IN1(n7168), .IN2(g1930), .QN(n11727) );
  NAND2X0 U11700 ( .IN1(n7167), .IN2(n10214), .QN(n11726) );
  NAND2X0 U11701 ( .IN1(n7169), .IN2(g7194), .QN(n11725) );
  INVX0 U11702 ( .INP(n11038), .ZN(n11027) );
  NAND3X0 U11703 ( .IN1(n11728), .IN2(n11729), .IN3(n11730), .QN(n11038) );
  NAND2X0 U11704 ( .IN1(n7330), .IN2(g1930), .QN(n11730) );
  NAND2X0 U11705 ( .IN1(n7329), .IN2(n10214), .QN(n11729) );
  NAND2X0 U11706 ( .IN1(n7331), .IN2(g7194), .QN(n11728) );
  NAND3X0 U11707 ( .IN1(n11731), .IN2(n11732), .IN3(n11733), .QN(n11056) );
  NAND2X0 U11708 ( .IN1(n7352), .IN2(g1930), .QN(n11733) );
  NAND2X0 U11709 ( .IN1(n10214), .IN2(n8092), .QN(n11732) );
  NAND2X0 U11710 ( .IN1(n7353), .IN2(g7194), .QN(n11731) );
  NOR2X0 U11711 ( .IN1(n10215), .IN2(n11569), .QN(n11506) );
  INVX0 U11712 ( .INP(g22651), .ZN(n11569) );
  INVX0 U11713 ( .INP(g7052), .ZN(n10215) );
  NAND2X0 U11714 ( .IN1(n11734), .IN2(n11735), .QN(g27289) );
  INVX0 U11715 ( .INP(n11736), .ZN(n11735) );
  NOR2X0 U11716 ( .IN1(n11653), .IN2(n7374), .QN(n11736) );
  NAND2X0 U11717 ( .IN1(n11653), .IN2(n11577), .QN(n11734) );
  INVX0 U11718 ( .INP(n11737), .ZN(n11577) );
  NAND2X0 U11719 ( .IN1(n11738), .IN2(n11739), .QN(n11737) );
  NAND2X0 U11720 ( .IN1(n11654), .IN2(n11740), .QN(n11739) );
  NAND3X0 U11721 ( .IN1(n11741), .IN2(n11742), .IN3(n11655), .QN(n11738) );
  NAND2X0 U11722 ( .IN1(n11743), .IN2(n11744), .QN(g27288) );
  NAND2X0 U11723 ( .IN1(n11573), .IN2(g1739), .QN(n11744) );
  NAND2X0 U11724 ( .IN1(n11663), .IN2(n11572), .QN(n11743) );
  NAND2X0 U11725 ( .IN1(n11745), .IN2(n11746), .QN(g27287) );
  INVX0 U11726 ( .INP(n11747), .ZN(n11746) );
  NOR2X0 U11727 ( .IN1(n11519), .IN2(n7646), .QN(n11747) );
  NAND2X0 U11728 ( .IN1(n11748), .IN2(n11519), .QN(n11745) );
  INVX0 U11729 ( .INP(n11749), .ZN(n11519) );
  NAND2X0 U11730 ( .IN1(n11750), .IN2(n10075), .QN(n11749) );
  NAND2X0 U11731 ( .IN1(n11751), .IN2(n11752), .QN(g27286) );
  NAND2X0 U11732 ( .IN1(n11582), .IN2(g1265), .QN(n11752) );
  NAND2X0 U11733 ( .IN1(n11580), .IN2(n11588), .QN(n11751) );
  INVX0 U11734 ( .INP(n11753), .ZN(n11588) );
  NAND2X0 U11735 ( .IN1(n11754), .IN2(n11755), .QN(n11753) );
  NAND2X0 U11736 ( .IN1(n11669), .IN2(n11180), .QN(n11754) );
  XNOR2X1 U11737 ( .IN1(n8785), .IN2(n11130), .Q(n11669) );
  NAND2X0 U11738 ( .IN1(n11756), .IN2(n11757), .QN(g27285) );
  INVX0 U11739 ( .INP(n11758), .ZN(n11757) );
  NOR2X0 U11740 ( .IN1(n11523), .IN2(n7334), .QN(n11758) );
  NAND2X0 U11741 ( .IN1(n11523), .IN2(n11675), .QN(n11756) );
  NOR2X0 U11742 ( .IN1(n4316), .IN2(n11759), .QN(n11523) );
  INVX0 U11743 ( .INP(g22615), .ZN(n11759) );
  NAND2X0 U11744 ( .IN1(n11760), .IN2(n11761), .QN(g27284) );
  NAND2X0 U11745 ( .IN1(n11762), .IN2(g1085), .QN(n11761) );
  NAND2X0 U11746 ( .IN1(n11763), .IN2(n11593), .QN(n11760) );
  NAND3X0 U11747 ( .IN1(n11764), .IN2(n11765), .IN3(n11766), .QN(n11593) );
  NAND2X0 U11748 ( .IN1(n11767), .IN2(n11768), .QN(g27283) );
  INVX0 U11749 ( .INP(n11769), .ZN(n11768) );
  NOR2X0 U11750 ( .IN1(n11679), .IN2(n7377), .QN(n11769) );
  NAND2X0 U11751 ( .IN1(n11679), .IN2(n11683), .QN(n11767) );
  NAND2X0 U11752 ( .IN1(n11770), .IN2(n11771), .QN(g27282) );
  INVX0 U11753 ( .INP(n11772), .ZN(n11771) );
  NOR2X0 U11754 ( .IN1(n11592), .IN2(n7626), .QN(n11772) );
  NAND2X0 U11755 ( .IN1(n11773), .IN2(n11592), .QN(n11770) );
  NAND2X0 U11756 ( .IN1(n11774), .IN2(n11775), .QN(g27281) );
  NAND2X0 U11757 ( .IN1(n11688), .IN2(g582), .QN(n11775) );
  NAND2X0 U11758 ( .IN1(n11686), .IN2(n11601), .QN(n11774) );
  INVX0 U11759 ( .INP(n11776), .ZN(n11601) );
  NAND2X0 U11760 ( .IN1(n11777), .IN2(n11778), .QN(n11776) );
  NAND2X0 U11761 ( .IN1(n11779), .IN2(n11279), .QN(n11778) );
  NAND2X0 U11762 ( .IN1(n11687), .IN2(n11248), .QN(n11777) );
  INVX0 U11763 ( .INP(n11779), .ZN(n11687) );
  NAND2X0 U11764 ( .IN1(n11780), .IN2(n11781), .QN(g27280) );
  NAND2X0 U11765 ( .IN1(test_so25), .IN2(n11597), .QN(n11781) );
  NAND2X0 U11766 ( .IN1(n11596), .IN2(n11694), .QN(n11780) );
  NAND2X0 U11767 ( .IN1(n11782), .IN2(n11783), .QN(g27279) );
  INVX0 U11768 ( .INP(n11784), .ZN(n11783) );
  NOR2X0 U11769 ( .IN1(n11531), .IN2(n7336), .QN(n11784) );
  NAND2X0 U11770 ( .IN1(n11531), .IN2(n11785), .QN(n11782) );
  NOR2X0 U11771 ( .IN1(n4313), .IN2(n11786), .QN(n11531) );
  NAND2X0 U11772 ( .IN1(n11787), .IN2(n11788), .QN(g27278) );
  NAND2X0 U11773 ( .IN1(n11789), .IN2(g388), .QN(n11788) );
  NAND2X0 U11774 ( .IN1(n11790), .IN2(n11699), .QN(n11787) );
  NAND2X0 U11775 ( .IN1(n11791), .IN2(n11792), .QN(g27277) );
  NAND2X0 U11776 ( .IN1(n11697), .IN2(g376), .QN(n11792) );
  NAND2X0 U11777 ( .IN1(n11698), .IN2(n11793), .QN(n11791) );
  NAND2X0 U11778 ( .IN1(n11794), .IN2(n11795), .QN(g27276) );
  INVX0 U11779 ( .INP(n11796), .ZN(n11795) );
  NOR2X0 U11780 ( .IN1(n11544), .IN2(n7645), .QN(n11796) );
  NAND2X0 U11781 ( .IN1(n11640), .IN2(n11544), .QN(n11794) );
  NOR2X0 U11782 ( .IN1(n11641), .IN2(n11797), .QN(n11544) );
  INVX0 U11783 ( .INP(g5555), .ZN(n11797) );
  NAND2X0 U11784 ( .IN1(n8667), .IN2(n11798), .QN(n11641) );
  NAND2X0 U11785 ( .IN1(n11799), .IN2(n8644), .QN(n11798) );
  INVX0 U11786 ( .INP(n10016), .ZN(n8644) );
  INVX0 U11787 ( .INP(n11800), .ZN(n11640) );
  NAND3X0 U11788 ( .IN1(n11801), .IN2(n11802), .IN3(n11803), .QN(n11800) );
  NAND2X0 U11789 ( .IN1(g3229), .IN2(n11804), .QN(n11803) );
  INVX0 U11790 ( .INP(n11805), .ZN(n11802) );
  NOR2X0 U11791 ( .IN1(n11806), .IN2(g3229), .QN(n11805) );
  NAND3X0 U11792 ( .IN1(n11632), .IN2(n11706), .IN3(n11806), .QN(n11801) );
  NAND2X0 U11793 ( .IN1(n11547), .IN2(n11631), .QN(n11806) );
  NAND3X0 U11794 ( .IN1(n11807), .IN2(n11808), .IN3(n11809), .QN(n11631) );
  NAND2X0 U11795 ( .IN1(n7621), .IN2(n10027), .QN(n11809) );
  NAND2X0 U11796 ( .IN1(n7620), .IN2(n10028), .QN(n11808) );
  NAND2X0 U11797 ( .IN1(n7622), .IN2(n10029), .QN(n11807) );
  INVX0 U11798 ( .INP(n11705), .ZN(n11547) );
  NAND3X0 U11799 ( .IN1(n11810), .IN2(n11811), .IN3(n11812), .QN(n11705) );
  NAND2X0 U11800 ( .IN1(n7373), .IN2(n10027), .QN(n11812) );
  NAND2X0 U11801 ( .IN1(n7372), .IN2(n10028), .QN(n11811) );
  NAND2X0 U11802 ( .IN1(n7371), .IN2(n10029), .QN(n11810) );
  NAND3X0 U11803 ( .IN1(n11813), .IN2(n11814), .IN3(n11815), .QN(n11706) );
  NAND2X0 U11804 ( .IN1(n7644), .IN2(n10027), .QN(n11815) );
  NAND2X0 U11805 ( .IN1(n7643), .IN2(n10028), .QN(n11814) );
  NAND2X0 U11806 ( .IN1(n7645), .IN2(n10029), .QN(n11813) );
  INVX0 U11807 ( .INP(n11804), .ZN(n11632) );
  NAND3X0 U11808 ( .IN1(n11816), .IN2(n11817), .IN3(n11818), .QN(n11804) );
  NAND2X0 U11809 ( .IN1(n7633), .IN2(n10027), .QN(n11818) );
  NAND2X0 U11810 ( .IN1(n7632), .IN2(n10028), .QN(n11817) );
  NAND2X0 U11811 ( .IN1(n7634), .IN2(n10029), .QN(n11816) );
  NAND2X0 U11812 ( .IN1(n11819), .IN2(n11820), .QN(g27275) );
  INVX0 U11813 ( .INP(n11821), .ZN(n11820) );
  NOR2X0 U11814 ( .IN1(n11653), .IN2(n7625), .QN(n11821) );
  NAND2X0 U11815 ( .IN1(n11663), .IN2(n11653), .QN(n11819) );
  NAND2X0 U11816 ( .IN1(n11822), .IN2(n11823), .QN(n11663) );
  NAND2X0 U11817 ( .IN1(n11656), .IN2(n11655), .QN(n11823) );
  INVX0 U11818 ( .INP(n11740), .ZN(n11655) );
  NAND2X0 U11819 ( .IN1(n11654), .IN2(n11824), .QN(n11822) );
  INVX0 U11820 ( .INP(n11742), .ZN(n11654) );
  XOR2X1 U11821 ( .IN1(n8785), .IN2(n11825), .Q(n11742) );
  NAND2X0 U11822 ( .IN1(n11826), .IN2(n11827), .QN(g27274) );
  NAND2X0 U11823 ( .IN1(n11573), .IN2(g1724), .QN(n11827) );
  NAND2X0 U11824 ( .IN1(n11748), .IN2(n11572), .QN(n11826) );
  INVX0 U11825 ( .INP(n11573), .ZN(n11572) );
  NAND2X0 U11826 ( .IN1(n11750), .IN2(g7014), .QN(n11573) );
  NAND2X0 U11827 ( .IN1(n11828), .IN2(n11829), .QN(g27273) );
  NAND2X0 U11828 ( .IN1(n11582), .IN2(g1262), .QN(n11829) );
  NAND2X0 U11829 ( .IN1(n11580), .IN2(n11675), .QN(n11828) );
  NOR2X0 U11830 ( .IN1(n11830), .IN2(n11831), .QN(n11675) );
  NOR2X0 U11831 ( .IN1(n11832), .IN2(g3229), .QN(n11831) );
  INVX0 U11832 ( .INP(n11833), .ZN(n11832) );
  NAND2X0 U11833 ( .IN1(n11755), .IN2(n11834), .QN(n11833) );
  NAND2X0 U11834 ( .IN1(n11146), .IN2(n11141), .QN(n11834) );
  INVX0 U11835 ( .INP(n11159), .ZN(n11146) );
  NAND2X0 U11836 ( .IN1(n11144), .IN2(n11150), .QN(n11755) );
  INVX0 U11837 ( .INP(n11180), .ZN(n11144) );
  NOR2X0 U11838 ( .IN1(n8785), .IN2(n11835), .QN(n11830) );
  NOR2X0 U11839 ( .IN1(n11159), .IN2(n11836), .QN(n11835) );
  NOR2X0 U11840 ( .IN1(n11130), .IN2(n11837), .QN(n11836) );
  NOR2X0 U11841 ( .IN1(n11180), .IN2(n11181), .QN(n11837) );
  NOR2X0 U11842 ( .IN1(n11159), .IN2(n11150), .QN(n11181) );
  NAND3X0 U11843 ( .IN1(n11838), .IN2(n11839), .IN3(n11840), .QN(n11150) );
  NAND2X0 U11844 ( .IN1(n7344), .IN2(n11104), .QN(n11840) );
  NAND2X0 U11845 ( .IN1(n7345), .IN2(g1236), .QN(n11839) );
  NAND2X0 U11846 ( .IN1(n7346), .IN2(g6944), .QN(n11838) );
  NAND3X0 U11847 ( .IN1(n11841), .IN2(n11842), .IN3(n11843), .QN(n11180) );
  NAND2X0 U11848 ( .IN1(n7170), .IN2(n11104), .QN(n11843) );
  NAND2X0 U11849 ( .IN1(g1236), .IN2(n8108), .QN(n11842) );
  NAND2X0 U11850 ( .IN1(n7171), .IN2(g6944), .QN(n11841) );
  INVX0 U11851 ( .INP(n11141), .ZN(n11130) );
  NAND3X0 U11852 ( .IN1(n11844), .IN2(n11845), .IN3(n11846), .QN(n11141) );
  NAND2X0 U11853 ( .IN1(n7332), .IN2(n11104), .QN(n11846) );
  NAND2X0 U11854 ( .IN1(n7333), .IN2(g1236), .QN(n11845) );
  NAND2X0 U11855 ( .IN1(n7334), .IN2(g6944), .QN(n11844) );
  NAND3X0 U11856 ( .IN1(n11847), .IN2(n11848), .IN3(n11849), .QN(n11159) );
  NAND2X0 U11857 ( .IN1(n7354), .IN2(n11104), .QN(n11849) );
  NAND2X0 U11858 ( .IN1(n7355), .IN2(g1236), .QN(n11848) );
  NAND2X0 U11859 ( .IN1(n7356), .IN2(g6944), .QN(n11847) );
  INVX0 U11860 ( .INP(n11582), .ZN(n11580) );
  NAND2X0 U11861 ( .IN1(g6750), .IN2(g22615), .QN(n11582) );
  NAND2X0 U11862 ( .IN1(n11850), .IN2(n11851), .QN(g27272) );
  NAND2X0 U11863 ( .IN1(test_so37), .IN2(n11762), .QN(n11851) );
  NAND2X0 U11864 ( .IN1(n11763), .IN2(n11683), .QN(n11850) );
  INVX0 U11865 ( .INP(n11852), .ZN(n11683) );
  NAND2X0 U11866 ( .IN1(n11853), .IN2(n11854), .QN(n11852) );
  NAND2X0 U11867 ( .IN1(n11764), .IN2(n11855), .QN(n11854) );
  NAND3X0 U11868 ( .IN1(n11856), .IN2(n11857), .IN3(n11765), .QN(n11853) );
  NAND2X0 U11869 ( .IN1(n11858), .IN2(n11859), .QN(g27271) );
  INVX0 U11870 ( .INP(n11860), .ZN(n11859) );
  NOR2X0 U11871 ( .IN1(n11679), .IN2(n7627), .QN(n11860) );
  NAND2X0 U11872 ( .IN1(n11773), .IN2(n11679), .QN(n11858) );
  NAND2X0 U11873 ( .IN1(n11861), .IN2(n11862), .QN(g27270) );
  INVX0 U11874 ( .INP(n11863), .ZN(n11862) );
  NOR2X0 U11875 ( .IN1(n11592), .IN2(n7649), .QN(n11863) );
  NAND2X0 U11876 ( .IN1(n11864), .IN2(n11592), .QN(n11861) );
  NOR2X0 U11877 ( .IN1(n11865), .IN2(n4381), .QN(n11592) );
  NAND2X0 U11878 ( .IN1(n11866), .IN2(n11867), .QN(g27269) );
  NAND2X0 U11879 ( .IN1(n11688), .IN2(g579), .QN(n11867) );
  NAND2X0 U11880 ( .IN1(n11686), .IN2(n11694), .QN(n11866) );
  INVX0 U11881 ( .INP(n11868), .ZN(n11694) );
  NAND2X0 U11882 ( .IN1(n11869), .IN2(n11870), .QN(n11868) );
  NAND2X0 U11883 ( .IN1(n11779), .IN2(n11278), .QN(n11869) );
  XNOR2X1 U11884 ( .IN1(n8785), .IN2(n11228), .Q(n11779) );
  NAND2X0 U11885 ( .IN1(n11871), .IN2(n11872), .QN(g27268) );
  NAND2X0 U11886 ( .IN1(n11597), .IN2(g577), .QN(n11872) );
  INVX0 U11887 ( .INP(n11596), .ZN(n11597) );
  NAND2X0 U11888 ( .IN1(n11596), .IN2(n11785), .QN(n11871) );
  NOR2X0 U11889 ( .IN1(n4372), .IN2(n11786), .QN(n11596) );
  INVX0 U11890 ( .INP(g22578), .ZN(n11786) );
  NAND2X0 U11891 ( .IN1(n11873), .IN2(n11874), .QN(g27267) );
  NAND2X0 U11892 ( .IN1(n11875), .IN2(g398), .QN(n11874) );
  NAND2X0 U11893 ( .IN1(n11876), .IN2(n11699), .QN(n11873) );
  NAND3X0 U11894 ( .IN1(n11877), .IN2(n11878), .IN3(n11879), .QN(n11699) );
  NAND2X0 U11895 ( .IN1(n11880), .IN2(n11881), .QN(g27266) );
  NAND2X0 U11896 ( .IN1(n11789), .IN2(g373), .QN(n11881) );
  NAND2X0 U11897 ( .IN1(n11790), .IN2(n11793), .QN(n11880) );
  NAND2X0 U11898 ( .IN1(n11882), .IN2(n11883), .QN(g27265) );
  NAND2X0 U11899 ( .IN1(n11697), .IN2(g361), .QN(n11883) );
  NAND2X0 U11900 ( .IN1(n11884), .IN2(n11698), .QN(n11882) );
  NAND2X0 U11901 ( .IN1(n11885), .IN2(n11886), .QN(g27264) );
  INVX0 U11902 ( .INP(n11887), .ZN(n11886) );
  NOR2X0 U11903 ( .IN1(n11653), .IN2(n7648), .QN(n11887) );
  NAND2X0 U11904 ( .IN1(n11748), .IN2(n11653), .QN(n11885) );
  INVX0 U11905 ( .INP(n11888), .ZN(n11653) );
  NAND2X0 U11906 ( .IN1(n11750), .IN2(g5511), .QN(n11888) );
  NOR2X0 U11907 ( .IN1(n11889), .IN2(n11890), .QN(n11750) );
  NOR2X0 U11908 ( .IN1(n8578), .IN2(n8615), .QN(n11890) );
  INVX0 U11909 ( .INP(n11891), .ZN(n11748) );
  NAND3X0 U11910 ( .IN1(n11892), .IN2(n11893), .IN3(n11894), .QN(n11891) );
  NAND2X0 U11911 ( .IN1(g3229), .IN2(n11895), .QN(n11894) );
  INVX0 U11912 ( .INP(n11896), .ZN(n11893) );
  NOR2X0 U11913 ( .IN1(n11897), .IN2(g3229), .QN(n11896) );
  NAND3X0 U11914 ( .IN1(n11741), .IN2(n11825), .IN3(n11897), .QN(n11892) );
  NAND2X0 U11915 ( .IN1(n11656), .IN2(n11740), .QN(n11897) );
  NAND3X0 U11916 ( .IN1(n11898), .IN2(n11899), .IN3(n11900), .QN(n11740) );
  NAND2X0 U11917 ( .IN1(n7624), .IN2(n10074), .QN(n11900) );
  NAND2X0 U11918 ( .IN1(n7623), .IN2(n10075), .QN(n11899) );
  NAND2X0 U11919 ( .IN1(n7625), .IN2(n10076), .QN(n11898) );
  INVX0 U11920 ( .INP(n11824), .ZN(n11656) );
  NAND3X0 U11921 ( .IN1(n11901), .IN2(n11902), .IN3(n11903), .QN(n11824) );
  NAND2X0 U11922 ( .IN1(n7376), .IN2(n10074), .QN(n11903) );
  NAND2X0 U11923 ( .IN1(n7375), .IN2(n10075), .QN(n11902) );
  NAND2X0 U11924 ( .IN1(n7374), .IN2(n10076), .QN(n11901) );
  NAND3X0 U11925 ( .IN1(n11904), .IN2(n11905), .IN3(n11906), .QN(n11825) );
  NAND2X0 U11926 ( .IN1(n7647), .IN2(n10074), .QN(n11906) );
  NAND2X0 U11927 ( .IN1(n7646), .IN2(n10075), .QN(n11905) );
  NAND2X0 U11928 ( .IN1(n7648), .IN2(n10076), .QN(n11904) );
  INVX0 U11929 ( .INP(n11895), .ZN(n11741) );
  NAND3X0 U11930 ( .IN1(n11907), .IN2(n11908), .IN3(n11909), .QN(n11895) );
  NAND2X0 U11931 ( .IN1(n10074), .IN2(n8096), .QN(n11909) );
  NAND2X0 U11932 ( .IN1(n7635), .IN2(n10075), .QN(n11908) );
  NAND2X0 U11933 ( .IN1(n7636), .IN2(n10076), .QN(n11907) );
  NAND2X0 U11934 ( .IN1(n11910), .IN2(n11911), .QN(g27263) );
  NAND2X0 U11935 ( .IN1(n11762), .IN2(g1056), .QN(n11911) );
  NAND2X0 U11936 ( .IN1(n11773), .IN2(n11763), .QN(n11910) );
  NAND2X0 U11937 ( .IN1(n11912), .IN2(n11913), .QN(n11773) );
  NAND2X0 U11938 ( .IN1(n11766), .IN2(n11765), .QN(n11913) );
  INVX0 U11939 ( .INP(n11855), .ZN(n11765) );
  NAND2X0 U11940 ( .IN1(n11764), .IN2(n11914), .QN(n11912) );
  INVX0 U11941 ( .INP(n11857), .ZN(n11764) );
  XOR2X1 U11942 ( .IN1(n8785), .IN2(n11915), .Q(n11857) );
  NAND2X0 U11943 ( .IN1(n11916), .IN2(n11917), .QN(g27262) );
  INVX0 U11944 ( .INP(n11918), .ZN(n11917) );
  NOR2X0 U11945 ( .IN1(n11679), .IN2(n7650), .QN(n11918) );
  NAND2X0 U11946 ( .IN1(n11864), .IN2(n11679), .QN(n11916) );
  NOR2X0 U11947 ( .IN1(n11865), .IN2(n4364), .QN(n11679) );
  NAND2X0 U11948 ( .IN1(n11919), .IN2(n11920), .QN(g27261) );
  NAND2X0 U11949 ( .IN1(n11688), .IN2(g576), .QN(n11920) );
  NAND2X0 U11950 ( .IN1(n11686), .IN2(n11785), .QN(n11919) );
  NOR2X0 U11951 ( .IN1(n11921), .IN2(n11922), .QN(n11785) );
  NOR2X0 U11952 ( .IN1(n11923), .IN2(g3229), .QN(n11922) );
  INVX0 U11953 ( .INP(n11924), .ZN(n11923) );
  NAND2X0 U11954 ( .IN1(n11870), .IN2(n11925), .QN(n11924) );
  NAND2X0 U11955 ( .IN1(n11244), .IN2(n11239), .QN(n11925) );
  INVX0 U11956 ( .INP(n11257), .ZN(n11244) );
  NAND2X0 U11957 ( .IN1(n11242), .IN2(n11248), .QN(n11870) );
  INVX0 U11958 ( .INP(n11278), .ZN(n11242) );
  NOR2X0 U11959 ( .IN1(n8785), .IN2(n11926), .QN(n11921) );
  NOR2X0 U11960 ( .IN1(n11257), .IN2(n11927), .QN(n11926) );
  NOR2X0 U11961 ( .IN1(n11228), .IN2(n11928), .QN(n11927) );
  NOR2X0 U11962 ( .IN1(n11278), .IN2(n11279), .QN(n11928) );
  NOR2X0 U11963 ( .IN1(n11257), .IN2(n11248), .QN(n11279) );
  NAND3X0 U11964 ( .IN1(n11929), .IN2(n11930), .IN3(n11931), .QN(n11248) );
  NAND2X0 U11965 ( .IN1(g6642), .IN2(n8109), .QN(n11931) );
  NAND2X0 U11966 ( .IN1(n7347), .IN2(n11207), .QN(n11930) );
  NAND2X0 U11967 ( .IN1(n7348), .IN2(g550), .QN(n11929) );
  NAND3X0 U11968 ( .IN1(n11932), .IN2(n11933), .IN3(n11934), .QN(n11278) );
  NAND2X0 U11969 ( .IN1(n7174), .IN2(g6642), .QN(n11934) );
  NAND2X0 U11970 ( .IN1(n7172), .IN2(n11207), .QN(n11933) );
  NAND2X0 U11971 ( .IN1(n7173), .IN2(g550), .QN(n11932) );
  INVX0 U11972 ( .INP(n11239), .ZN(n11228) );
  NAND3X0 U11973 ( .IN1(n11935), .IN2(n11936), .IN3(n11937), .QN(n11239) );
  NAND2X0 U11974 ( .IN1(n7337), .IN2(g6642), .QN(n11937) );
  NAND2X0 U11975 ( .IN1(n7335), .IN2(n11207), .QN(n11936) );
  NAND2X0 U11976 ( .IN1(n7336), .IN2(g550), .QN(n11935) );
  NAND3X0 U11977 ( .IN1(n11938), .IN2(n11939), .IN3(n11940), .QN(n11257) );
  NAND2X0 U11978 ( .IN1(n7359), .IN2(g6642), .QN(n11940) );
  NAND2X0 U11979 ( .IN1(n7357), .IN2(n11207), .QN(n11939) );
  NAND2X0 U11980 ( .IN1(n7358), .IN2(g550), .QN(n11938) );
  INVX0 U11981 ( .INP(n11688), .ZN(n11686) );
  NAND2X0 U11982 ( .IN1(g6485), .IN2(g22578), .QN(n11688) );
  NAND2X0 U11983 ( .IN1(n11941), .IN2(n11942), .QN(g27260) );
  NAND2X0 U11984 ( .IN1(n11875), .IN2(g384), .QN(n11942) );
  NAND2X0 U11985 ( .IN1(n11876), .IN2(n11793), .QN(n11941) );
  INVX0 U11986 ( .INP(n11943), .ZN(n11793) );
  NAND2X0 U11987 ( .IN1(n11944), .IN2(n11945), .QN(n11943) );
  NAND2X0 U11988 ( .IN1(n11877), .IN2(n11946), .QN(n11945) );
  NAND3X0 U11989 ( .IN1(n11947), .IN2(n11948), .IN3(n11878), .QN(n11944) );
  NAND2X0 U11990 ( .IN1(n11949), .IN2(n11950), .QN(g27259) );
  NAND2X0 U11991 ( .IN1(n11789), .IN2(g358), .QN(n11950) );
  NAND2X0 U11992 ( .IN1(n11884), .IN2(n11790), .QN(n11949) );
  NAND2X0 U11993 ( .IN1(n11951), .IN2(n11952), .QN(g27258) );
  NAND2X0 U11994 ( .IN1(test_so16), .IN2(n11697), .QN(n11952) );
  NAND2X0 U11995 ( .IN1(n11953), .IN2(n11698), .QN(n11951) );
  INVX0 U11996 ( .INP(n11697), .ZN(n11698) );
  NAND2X0 U11997 ( .IN1(n11954), .IN2(n10160), .QN(n11697) );
  NAND2X0 U11998 ( .IN1(n11955), .IN2(n11956), .QN(g27257) );
  NAND2X0 U11999 ( .IN1(n11762), .IN2(g1041), .QN(n11956) );
  INVX0 U12000 ( .INP(n11763), .ZN(n11762) );
  NAND2X0 U12001 ( .IN1(n11864), .IN2(n11763), .QN(n11955) );
  NOR2X0 U12002 ( .IN1(n11865), .IN2(n4363), .QN(n11763) );
  NAND2X0 U12003 ( .IN1(n8608), .IN2(n11957), .QN(n11865) );
  NAND2X0 U12004 ( .IN1(n11799), .IN2(n8585), .QN(n11957) );
  INVX0 U12005 ( .INP(n10106), .ZN(n8585) );
  INVX0 U12006 ( .INP(n11958), .ZN(n11864) );
  NAND3X0 U12007 ( .IN1(n11959), .IN2(n11960), .IN3(n11961), .QN(n11958) );
  NAND2X0 U12008 ( .IN1(g3229), .IN2(n11962), .QN(n11961) );
  INVX0 U12009 ( .INP(n11963), .ZN(n11960) );
  NOR2X0 U12010 ( .IN1(n11964), .IN2(g3229), .QN(n11963) );
  NAND3X0 U12011 ( .IN1(n11856), .IN2(n11915), .IN3(n11964), .QN(n11959) );
  NAND2X0 U12012 ( .IN1(n11766), .IN2(n11855), .QN(n11964) );
  NAND3X0 U12013 ( .IN1(n11965), .IN2(n11966), .IN3(n11967), .QN(n11855) );
  NAND2X0 U12014 ( .IN1(n7626), .IN2(g1088), .QN(n11967) );
  NAND2X0 U12015 ( .IN1(n7628), .IN2(g5472), .QN(n11966) );
  NAND2X0 U12016 ( .IN1(n7627), .IN2(g6712), .QN(n11965) );
  INVX0 U12017 ( .INP(n11914), .ZN(n11766) );
  NAND3X0 U12018 ( .IN1(n11968), .IN2(n11969), .IN3(n11970), .QN(n11914) );
  NAND2X0 U12019 ( .IN1(n7378), .IN2(g1088), .QN(n11970) );
  NAND2X0 U12020 ( .IN1(g5472), .IN2(n8097), .QN(n11969) );
  NAND2X0 U12021 ( .IN1(n7377), .IN2(g6712), .QN(n11968) );
  NAND3X0 U12022 ( .IN1(n11971), .IN2(n11972), .IN3(n11973), .QN(n11915) );
  NAND2X0 U12023 ( .IN1(n7649), .IN2(g1088), .QN(n11973) );
  NAND2X0 U12024 ( .IN1(n7651), .IN2(g5472), .QN(n11972) );
  NAND2X0 U12025 ( .IN1(n7650), .IN2(g6712), .QN(n11971) );
  INVX0 U12026 ( .INP(n11962), .ZN(n11856) );
  NAND3X0 U12027 ( .IN1(n11974), .IN2(n11975), .IN3(n11976), .QN(n11962) );
  NAND2X0 U12028 ( .IN1(n7637), .IN2(g1088), .QN(n11976) );
  NAND2X0 U12029 ( .IN1(n7639), .IN2(g5472), .QN(n11975) );
  NAND2X0 U12030 ( .IN1(n7638), .IN2(g6712), .QN(n11974) );
  NAND2X0 U12031 ( .IN1(n11977), .IN2(n11978), .QN(g27256) );
  NAND2X0 U12032 ( .IN1(n11875), .IN2(g369), .QN(n11978) );
  NAND2X0 U12033 ( .IN1(n11884), .IN2(n11876), .QN(n11977) );
  NAND2X0 U12034 ( .IN1(n11979), .IN2(n11980), .QN(n11884) );
  NAND2X0 U12035 ( .IN1(n11879), .IN2(n11878), .QN(n11980) );
  INVX0 U12036 ( .INP(n11946), .ZN(n11878) );
  NAND2X0 U12037 ( .IN1(n11877), .IN2(n11981), .QN(n11979) );
  INVX0 U12038 ( .INP(n11948), .ZN(n11877) );
  XOR2X1 U12039 ( .IN1(n8785), .IN2(n11982), .Q(n11948) );
  NAND2X0 U12040 ( .IN1(n11983), .IN2(n11984), .QN(g27255) );
  NAND2X0 U12041 ( .IN1(n11789), .IN2(g343), .QN(n11984) );
  NAND2X0 U12042 ( .IN1(n11953), .IN2(n11790), .QN(n11983) );
  INVX0 U12043 ( .INP(n11789), .ZN(n11790) );
  NAND2X0 U12044 ( .IN1(n11954), .IN2(g6447), .QN(n11789) );
  NAND2X0 U12045 ( .IN1(n11985), .IN2(n11986), .QN(g27253) );
  NAND2X0 U12046 ( .IN1(n11875), .IN2(g354), .QN(n11986) );
  NAND2X0 U12047 ( .IN1(n11953), .IN2(n11876), .QN(n11985) );
  INVX0 U12048 ( .INP(n11875), .ZN(n11876) );
  NAND2X0 U12049 ( .IN1(n11954), .IN2(g5437), .QN(n11875) );
  NOR2X0 U12050 ( .IN1(n11987), .IN2(n11988), .QN(n11954) );
  NOR2X0 U12051 ( .IN1(n8578), .IN2(n8555), .QN(n11988) );
  INVX0 U12052 ( .INP(n11989), .ZN(n11953) );
  NAND3X0 U12053 ( .IN1(n11990), .IN2(n11991), .IN3(n11992), .QN(n11989) );
  NAND2X0 U12054 ( .IN1(g3229), .IN2(n11993), .QN(n11992) );
  INVX0 U12055 ( .INP(n11994), .ZN(n11991) );
  NOR2X0 U12056 ( .IN1(n11995), .IN2(g3229), .QN(n11994) );
  NAND3X0 U12057 ( .IN1(n11947), .IN2(n11982), .IN3(n11995), .QN(n11990) );
  NAND2X0 U12058 ( .IN1(n11879), .IN2(n11946), .QN(n11995) );
  NAND3X0 U12059 ( .IN1(n11996), .IN2(n11997), .IN3(n11998), .QN(n11946) );
  NAND2X0 U12060 ( .IN1(n7631), .IN2(n10158), .QN(n11998) );
  NAND2X0 U12061 ( .IN1(n7630), .IN2(n10159), .QN(n11997) );
  NAND2X0 U12062 ( .IN1(n7629), .IN2(n10160), .QN(n11996) );
  INVX0 U12063 ( .INP(n11981), .ZN(n11879) );
  NAND3X0 U12064 ( .IN1(n11999), .IN2(n12000), .IN3(n12001), .QN(n11981) );
  NAND2X0 U12065 ( .IN1(n7379), .IN2(n10158), .QN(n12001) );
  NAND2X0 U12066 ( .IN1(n7381), .IN2(n10159), .QN(n12000) );
  NAND2X0 U12067 ( .IN1(n7380), .IN2(n10160), .QN(n11999) );
  NAND3X0 U12068 ( .IN1(n12002), .IN2(n12003), .IN3(n12004), .QN(n11982) );
  NAND2X0 U12069 ( .IN1(n7653), .IN2(n10158), .QN(n12004) );
  NAND2X0 U12070 ( .IN1(n7652), .IN2(n10159), .QN(n12003) );
  NAND2X0 U12071 ( .IN1(n10160), .IN2(n8100), .QN(n12002) );
  INVX0 U12072 ( .INP(n11993), .ZN(n11947) );
  NAND3X0 U12073 ( .IN1(n12005), .IN2(n12006), .IN3(n12007), .QN(n11993) );
  NAND2X0 U12074 ( .IN1(n7642), .IN2(n10158), .QN(n12007) );
  NAND2X0 U12075 ( .IN1(n7641), .IN2(n10159), .QN(n12006) );
  NAND2X0 U12076 ( .IN1(n7640), .IN2(n10160), .QN(n12005) );
  NOR3X0 U12077 ( .IN1(n12008), .IN2(n11303), .IN3(n11306), .QN(g27243) );
  NOR3X0 U12078 ( .IN1(n9290), .IN2(n4471), .IN3(n8073), .QN(n11306) );
  NOR2X0 U12079 ( .IN1(n12009), .IN2(g2753), .QN(n12008) );
  NOR2X0 U12080 ( .IN1(n9290), .IN2(n8073), .QN(n12009) );
  NOR3X0 U12081 ( .IN1(n11409), .IN2(n10265), .IN3(n12010), .QN(g27131) );
  NOR2X0 U12082 ( .IN1(n3683), .IN2(g2147), .QN(n12010) );
  INVX0 U12083 ( .INP(n4522), .ZN(n11409) );
  NOR3X0 U12084 ( .IN1(n11411), .IN2(n10267), .IN3(n12011), .QN(g27129) );
  NOR2X0 U12085 ( .IN1(n3686), .IN2(g1453), .QN(n12011) );
  INVX0 U12086 ( .INP(n4523), .ZN(n11411) );
  NOR2X0 U12087 ( .IN1(n10269), .IN2(n12012), .QN(g27123) );
  XOR2X1 U12088 ( .IN1(n8063), .IN2(n3689), .Q(n12012) );
  NOR3X0 U12089 ( .IN1(n11414), .IN2(n10271), .IN3(n12013), .QN(g27120) );
  NOR2X0 U12090 ( .IN1(n3692), .IN2(test_so15), .QN(n12013) );
  INVX0 U12091 ( .INP(n4521), .ZN(n11414) );
  NAND2X0 U12092 ( .IN1(n12014), .IN2(n12015), .QN(g26827) );
  NAND2X0 U12093 ( .IN1(n12016), .IN2(n4606), .QN(n12015) );
  NAND2X0 U12094 ( .IN1(n4509), .IN2(g2519), .QN(n12014) );
  NAND2X0 U12095 ( .IN1(n12017), .IN2(n12018), .QN(g26826) );
  NAND2X0 U12096 ( .IN1(n12016), .IN2(g7264), .QN(n12018) );
  NAND2X0 U12097 ( .IN1(n4524), .IN2(g2516), .QN(n12017) );
  NAND2X0 U12098 ( .IN1(n12019), .IN2(n12020), .QN(g26825) );
  NAND2X0 U12099 ( .IN1(n4606), .IN2(n12021), .QN(n12020) );
  NAND2X0 U12100 ( .IN1(n4509), .IN2(g2510), .QN(n12019) );
  NAND2X0 U12101 ( .IN1(n12022), .IN2(n12023), .QN(g26824) );
  NAND2X0 U12102 ( .IN1(n12024), .IN2(n4618), .QN(n12023) );
  NAND2X0 U12103 ( .IN1(n4511), .IN2(test_so59), .QN(n12022) );
  NAND2X0 U12104 ( .IN1(n12025), .IN2(n12026), .QN(g26823) );
  NAND2X0 U12105 ( .IN1(n12016), .IN2(g5555), .QN(n12026) );
  XOR2X1 U12106 ( .IN1(n11339), .IN2(n12027), .Q(n12016) );
  NOR2X0 U12107 ( .IN1(n12028), .IN2(n11334), .QN(n12027) );
  NAND3X0 U12108 ( .IN1(n12029), .IN2(n12030), .IN3(test_so79), .QN(n11334) );
  NAND2X0 U12109 ( .IN1(n12031), .IN2(n11341), .QN(n12030) );
  NAND2X0 U12110 ( .IN1(n9165), .IN2(n9164), .QN(n12031) );
  INVX0 U12111 ( .INP(n11339), .ZN(n9165) );
  NAND2X0 U12112 ( .IN1(n9163), .IN2(n12032), .QN(n12029) );
  NAND2X0 U12113 ( .IN1(n11340), .IN2(n11339), .QN(n12032) );
  INVX0 U12114 ( .INP(n11341), .ZN(n9163) );
  INVX0 U12115 ( .INP(n11333), .ZN(n12028) );
  NAND3X0 U12116 ( .IN1(n12033), .IN2(n12034), .IN3(n12035), .QN(n11333) );
  NAND2X0 U12117 ( .IN1(n7655), .IN2(n10027), .QN(n12035) );
  NAND2X0 U12118 ( .IN1(n10028), .IN2(n8110), .QN(n12034) );
  NAND2X0 U12119 ( .IN1(n7664), .IN2(n10029), .QN(n12033) );
  NAND2X0 U12120 ( .IN1(n4516), .IN2(g2513), .QN(n12025) );
  NAND2X0 U12121 ( .IN1(n12036), .IN2(n12037), .QN(g26822) );
  NAND2X0 U12122 ( .IN1(g7264), .IN2(n12021), .QN(n12037) );
  NAND2X0 U12123 ( .IN1(n4524), .IN2(g2507), .QN(n12036) );
  NAND2X0 U12124 ( .IN1(n12038), .IN2(n12039), .QN(g26821) );
  NAND2X0 U12125 ( .IN1(n12024), .IN2(g7014), .QN(n12039) );
  NAND2X0 U12126 ( .IN1(n4525), .IN2(g1822), .QN(n12038) );
  NAND2X0 U12127 ( .IN1(n12040), .IN2(n12041), .QN(g26820) );
  NAND2X0 U12128 ( .IN1(n4618), .IN2(n12042), .QN(n12041) );
  NAND2X0 U12129 ( .IN1(n4511), .IN2(g1816), .QN(n12040) );
  NAND2X0 U12130 ( .IN1(n12043), .IN2(n12044), .QN(g26818) );
  NAND2X0 U12131 ( .IN1(n4381), .IN2(g1131), .QN(n12044) );
  NAND2X0 U12132 ( .IN1(n12045), .IN2(g1088), .QN(n12043) );
  NAND2X0 U12133 ( .IN1(n12046), .IN2(n12047), .QN(g26817) );
  NAND2X0 U12134 ( .IN1(g5555), .IN2(n12021), .QN(n12047) );
  NAND2X0 U12135 ( .IN1(n12048), .IN2(n12049), .QN(n12021) );
  NAND2X0 U12136 ( .IN1(n11341), .IN2(n8075), .QN(n12049) );
  NAND3X0 U12137 ( .IN1(n12050), .IN2(n12051), .IN3(n12052), .QN(n11341) );
  NAND2X0 U12138 ( .IN1(g5555), .IN2(g2504), .QN(n12052) );
  NAND2X0 U12139 ( .IN1(n4606), .IN2(g2510), .QN(n12051) );
  NAND2X0 U12140 ( .IN1(g7264), .IN2(g2507), .QN(n12050) );
  NAND2X0 U12141 ( .IN1(test_so79), .IN2(n9164), .QN(n12048) );
  INVX0 U12142 ( .INP(n11340), .ZN(n9164) );
  NAND2X0 U12143 ( .IN1(n10763), .IN2(n12053), .QN(n11340) );
  NAND3X0 U12144 ( .IN1(n12054), .IN2(n12055), .IN3(n12056), .QN(n12053) );
  NAND2X0 U12145 ( .IN1(n7568), .IN2(test_so73), .QN(n12056) );
  NAND2X0 U12146 ( .IN1(n7569), .IN2(g6837), .QN(n12055) );
  NAND2X0 U12147 ( .IN1(n7567), .IN2(g2241), .QN(n12054) );
  INVX0 U12148 ( .INP(n12057), .ZN(n10763) );
  NAND2X0 U12149 ( .IN1(n4516), .IN2(g2504), .QN(n12046) );
  NAND2X0 U12150 ( .IN1(n12058), .IN2(n12059), .QN(g26816) );
  NAND2X0 U12151 ( .IN1(n12024), .IN2(g5511), .QN(n12059) );
  XOR2X1 U12152 ( .IN1(n11359), .IN2(n12060), .Q(n12024) );
  NOR2X0 U12153 ( .IN1(n12061), .IN2(n11354), .QN(n12060) );
  NAND3X0 U12154 ( .IN1(n12062), .IN2(n12063), .IN3(g1690), .QN(n11354) );
  NAND2X0 U12155 ( .IN1(n12064), .IN2(n11361), .QN(n12063) );
  NAND2X0 U12156 ( .IN1(n9162), .IN2(n9161), .QN(n12064) );
  INVX0 U12157 ( .INP(n11359), .ZN(n9162) );
  NAND2X0 U12158 ( .IN1(n9160), .IN2(n12065), .QN(n12062) );
  NAND2X0 U12159 ( .IN1(n11360), .IN2(n11359), .QN(n12065) );
  INVX0 U12160 ( .INP(n11361), .ZN(n9160) );
  INVX0 U12161 ( .INP(n11353), .ZN(n12061) );
  NAND3X0 U12162 ( .IN1(n12066), .IN2(n12067), .IN3(n12068), .QN(n11353) );
  NAND2X0 U12163 ( .IN1(n7658), .IN2(n10074), .QN(n12068) );
  NAND2X0 U12164 ( .IN1(n7668), .IN2(n10075), .QN(n12067) );
  NAND2X0 U12165 ( .IN1(n7669), .IN2(n10076), .QN(n12066) );
  NAND2X0 U12166 ( .IN1(n4518), .IN2(g1819), .QN(n12058) );
  NAND2X0 U12167 ( .IN1(n12069), .IN2(n12070), .QN(g26815) );
  NAND2X0 U12168 ( .IN1(g7014), .IN2(n12042), .QN(n12070) );
  NAND2X0 U12169 ( .IN1(n4525), .IN2(g1813), .QN(n12069) );
  NAND2X0 U12170 ( .IN1(n12071), .IN2(n12072), .QN(g26814) );
  NAND2X0 U12171 ( .IN1(n4364), .IN2(g1128), .QN(n12072) );
  NAND2X0 U12172 ( .IN1(n12045), .IN2(g6712), .QN(n12071) );
  NAND2X0 U12173 ( .IN1(n12073), .IN2(n12074), .QN(g26813) );
  NAND2X0 U12174 ( .IN1(n4381), .IN2(g1122), .QN(n12074) );
  NAND2X0 U12175 ( .IN1(n12075), .IN2(g1088), .QN(n12073) );
  NAND2X0 U12176 ( .IN1(n12076), .IN2(n12077), .QN(g26812) );
  NAND2X0 U12177 ( .IN1(n12078), .IN2(n4640), .QN(n12077) );
  NAND2X0 U12178 ( .IN1(n4506), .IN2(g444), .QN(n12076) );
  NAND2X0 U12179 ( .IN1(n12079), .IN2(n12080), .QN(g26811) );
  NAND2X0 U12180 ( .IN1(g5511), .IN2(n12042), .QN(n12080) );
  NAND2X0 U12181 ( .IN1(n12081), .IN2(n12082), .QN(n12042) );
  NAND2X0 U12182 ( .IN1(n4386), .IN2(n11361), .QN(n12082) );
  NAND3X0 U12183 ( .IN1(n12083), .IN2(n12084), .IN3(n12085), .QN(n11361) );
  NAND2X0 U12184 ( .IN1(g5511), .IN2(g1810), .QN(n12085) );
  NAND2X0 U12185 ( .IN1(n4618), .IN2(g1816), .QN(n12084) );
  NAND2X0 U12186 ( .IN1(g7014), .IN2(g1813), .QN(n12083) );
  NAND2X0 U12187 ( .IN1(n9161), .IN2(g1690), .QN(n12081) );
  INVX0 U12188 ( .INP(n11360), .ZN(n9161) );
  NAND2X0 U12189 ( .IN1(n10801), .IN2(n12086), .QN(n11360) );
  NAND3X0 U12190 ( .IN1(n12087), .IN2(n12088), .IN3(n12089), .QN(n12086) );
  NAND2X0 U12191 ( .IN1(n7580), .IN2(g6782), .QN(n12089) );
  NAND2X0 U12192 ( .IN1(n7581), .IN2(g6573), .QN(n12088) );
  NAND2X0 U12193 ( .IN1(n7579), .IN2(g1547), .QN(n12087) );
  INVX0 U12194 ( .INP(n12090), .ZN(n10801) );
  NAND2X0 U12195 ( .IN1(n4518), .IN2(g1810), .QN(n12079) );
  NAND2X0 U12196 ( .IN1(n12091), .IN2(n12092), .QN(g26810) );
  NAND2X0 U12197 ( .IN1(n4363), .IN2(g1125), .QN(n12092) );
  NAND2X0 U12198 ( .IN1(n12045), .IN2(g5472), .QN(n12091) );
  XOR2X1 U12199 ( .IN1(n11379), .IN2(n12093), .Q(n12045) );
  NOR2X0 U12200 ( .IN1(n12094), .IN2(n11374), .QN(n12093) );
  NAND3X0 U12201 ( .IN1(n12095), .IN2(n12096), .IN3(g996), .QN(n11374) );
  NAND2X0 U12202 ( .IN1(n12097), .IN2(n11381), .QN(n12096) );
  NAND2X0 U12203 ( .IN1(n9159), .IN2(n9158), .QN(n12097) );
  INVX0 U12204 ( .INP(n11379), .ZN(n9159) );
  NAND2X0 U12205 ( .IN1(n9157), .IN2(n12098), .QN(n12095) );
  NAND2X0 U12206 ( .IN1(n11380), .IN2(n11379), .QN(n12098) );
  INVX0 U12207 ( .INP(n11381), .ZN(n9157) );
  INVX0 U12208 ( .INP(n11373), .ZN(n12094) );
  NAND3X0 U12209 ( .IN1(n12099), .IN2(n12100), .IN3(n12101), .QN(n11373) );
  NAND2X0 U12210 ( .IN1(n7674), .IN2(g1088), .QN(n12101) );
  NAND2X0 U12211 ( .IN1(n7675), .IN2(g5472), .QN(n12100) );
  NAND2X0 U12212 ( .IN1(n7661), .IN2(g6712), .QN(n12099) );
  NAND2X0 U12213 ( .IN1(n12102), .IN2(n12103), .QN(g26809) );
  NAND2X0 U12214 ( .IN1(n12075), .IN2(g6712), .QN(n12103) );
  NAND2X0 U12215 ( .IN1(n4364), .IN2(test_so38), .QN(n12102) );
  NAND2X0 U12216 ( .IN1(n12104), .IN2(n12105), .QN(g26808) );
  NAND2X0 U12217 ( .IN1(n12078), .IN2(g6447), .QN(n12105) );
  NAND2X0 U12218 ( .IN1(n4499), .IN2(g441), .QN(n12104) );
  NAND2X0 U12219 ( .IN1(n12106), .IN2(n12107), .QN(g26807) );
  NAND2X0 U12220 ( .IN1(n4640), .IN2(n12108), .QN(n12107) );
  NAND2X0 U12221 ( .IN1(n4506), .IN2(g435), .QN(n12106) );
  NAND2X0 U12222 ( .IN1(n12109), .IN2(n12110), .QN(g26806) );
  NAND2X0 U12223 ( .IN1(n4363), .IN2(g1116), .QN(n12110) );
  NAND2X0 U12224 ( .IN1(n12075), .IN2(g5472), .QN(n12109) );
  NAND2X0 U12225 ( .IN1(n12111), .IN2(n12112), .QN(n12075) );
  NAND2X0 U12226 ( .IN1(n4387), .IN2(n11381), .QN(n12112) );
  NAND3X0 U12227 ( .IN1(n12113), .IN2(n12114), .IN3(n12115), .QN(n11381) );
  NAND2X0 U12228 ( .IN1(g1088), .IN2(g1122), .QN(n12115) );
  NAND2X0 U12229 ( .IN1(g5472), .IN2(g1116), .QN(n12114) );
  NAND2X0 U12230 ( .IN1(test_so38), .IN2(g6712), .QN(n12113) );
  NAND2X0 U12231 ( .IN1(n9158), .IN2(g996), .QN(n12111) );
  INVX0 U12232 ( .INP(n11380), .ZN(n9158) );
  NAND2X0 U12233 ( .IN1(n10835), .IN2(n12116), .QN(n11380) );
  NAND3X0 U12234 ( .IN1(n12117), .IN2(n12118), .IN3(n12119), .QN(n12116) );
  NAND2X0 U12235 ( .IN1(n7590), .IN2(test_so31), .QN(n12119) );
  NAND2X0 U12236 ( .IN1(n7591), .IN2(g6518), .QN(n12118) );
  NAND2X0 U12237 ( .IN1(n7592), .IN2(g6368), .QN(n12117) );
  INVX0 U12238 ( .INP(n12120), .ZN(n10835) );
  NAND2X0 U12239 ( .IN1(n12121), .IN2(n12122), .QN(g26805) );
  NAND2X0 U12240 ( .IN1(n12078), .IN2(g5437), .QN(n12122) );
  XOR2X1 U12241 ( .IN1(n11394), .IN2(n12123), .Q(n12078) );
  NOR2X0 U12242 ( .IN1(n12124), .IN2(n11389), .QN(n12123) );
  NAND3X0 U12243 ( .IN1(n12125), .IN2(n12126), .IN3(g309), .QN(n11389) );
  NAND2X0 U12244 ( .IN1(n12127), .IN2(n11396), .QN(n12126) );
  NAND2X0 U12245 ( .IN1(n9156), .IN2(n9155), .QN(n12127) );
  INVX0 U12246 ( .INP(n11394), .ZN(n9156) );
  NAND2X0 U12247 ( .IN1(n9154), .IN2(n12128), .QN(n12125) );
  NAND2X0 U12248 ( .IN1(n11395), .IN2(n11394), .QN(n12128) );
  INVX0 U12249 ( .INP(n11396), .ZN(n9154) );
  INVX0 U12250 ( .INP(n11388), .ZN(n12124) );
  NAND3X0 U12251 ( .IN1(n12129), .IN2(n12130), .IN3(n12131), .QN(n11388) );
  NAND2X0 U12252 ( .IN1(n7683), .IN2(n10158), .QN(n12131) );
  NAND2X0 U12253 ( .IN1(n7682), .IN2(n10159), .QN(n12130) );
  NAND2X0 U12254 ( .IN1(n7681), .IN2(n10160), .QN(n12129) );
  NAND2X0 U12255 ( .IN1(n4520), .IN2(g438), .QN(n12121) );
  NAND2X0 U12256 ( .IN1(n12132), .IN2(n12133), .QN(g26804) );
  NAND2X0 U12257 ( .IN1(g6447), .IN2(n12108), .QN(n12133) );
  NAND2X0 U12258 ( .IN1(n4499), .IN2(g432), .QN(n12132) );
  NAND2X0 U12259 ( .IN1(n12134), .IN2(n12135), .QN(g26803) );
  NAND2X0 U12260 ( .IN1(g5437), .IN2(n12108), .QN(n12135) );
  NAND2X0 U12261 ( .IN1(n12136), .IN2(n12137), .QN(n12108) );
  NAND2X0 U12262 ( .IN1(n4388), .IN2(n11396), .QN(n12137) );
  NAND3X0 U12263 ( .IN1(n12138), .IN2(n12139), .IN3(n12140), .QN(n11396) );
  NAND2X0 U12264 ( .IN1(g5437), .IN2(g429), .QN(n12140) );
  NAND2X0 U12265 ( .IN1(n4640), .IN2(g435), .QN(n12139) );
  NAND2X0 U12266 ( .IN1(g6447), .IN2(g432), .QN(n12138) );
  NAND2X0 U12267 ( .IN1(n9155), .IN2(g309), .QN(n12136) );
  INVX0 U12268 ( .INP(n11395), .ZN(n9155) );
  NAND2X0 U12269 ( .IN1(n10862), .IN2(n12141), .QN(n11395) );
  NAND3X0 U12270 ( .IN1(n12142), .IN2(n12143), .IN3(n12144), .QN(n12141) );
  NAND2X0 U12271 ( .IN1(n7602), .IN2(g6313), .QN(n12144) );
  NAND2X0 U12272 ( .IN1(n7603), .IN2(g6231), .QN(n12143) );
  NAND2X0 U12273 ( .IN1(n7601), .IN2(g165), .QN(n12142) );
  INVX0 U12274 ( .INP(n12145), .ZN(n10862) );
  NAND2X0 U12275 ( .IN1(n4520), .IN2(g429), .QN(n12134) );
  NOR2X0 U12276 ( .IN1(n8672), .IN2(n12146), .QN(g26798) );
  XNOR2X1 U12277 ( .IN1(n4355), .IN2(n12147), .Q(n12146) );
  NAND2X0 U12278 ( .IN1(n12148), .IN2(g2900), .QN(n12147) );
  NOR2X0 U12279 ( .IN1(n11303), .IN2(n12149), .QN(g26795) );
  XOR2X1 U12280 ( .IN1(n9290), .IN2(test_so92), .Q(n12149) );
  NAND3X0 U12281 ( .IN1(g2734), .IN2(g2746), .IN3(n9292), .QN(n9290) );
  NOR2X0 U12282 ( .IN1(n9305), .IN2(n12150), .QN(g26789) );
  XOR2X1 U12283 ( .IN1(n4468), .IN2(n9306), .Q(n12150) );
  NOR3X0 U12284 ( .IN1(n4399), .IN2(n4409), .IN3(n9308), .QN(n9306) );
  INVX0 U12285 ( .INP(n12151), .ZN(n9308) );
  NOR2X0 U12286 ( .IN1(n12152), .IN2(n12153), .QN(g26786) );
  XOR2X1 U12287 ( .IN1(g3024), .IN2(n3741), .Q(n12152) );
  NOR2X0 U12288 ( .IN1(n8512), .IN2(n12154), .QN(g26781) );
  XNOR2X1 U12289 ( .IN1(n4469), .IN2(n8508), .Q(n12154) );
  NAND3X0 U12290 ( .IN1(g1346), .IN2(g1358), .IN3(n8510), .QN(n8508) );
  NOR2X0 U12291 ( .IN1(n8536), .IN2(n12155), .QN(g26776) );
  XOR2X1 U12292 ( .IN1(n8528), .IN2(test_so28), .Q(n12155) );
  NAND3X0 U12293 ( .IN1(g660), .IN2(g672), .IN3(n8530), .QN(n8528) );
  NAND2X0 U12294 ( .IN1(n12156), .IN2(n12157), .QN(g26676) );
  NAND2X0 U12295 ( .IN1(n12158), .IN2(g2479), .QN(n12157) );
  NAND2X0 U12296 ( .IN1(n12159), .IN2(n10027), .QN(n12158) );
  NAND2X0 U12297 ( .IN1(n12160), .IN2(n10027), .QN(n12156) );
  NAND2X0 U12298 ( .IN1(n12161), .IN2(n12162), .QN(g26675) );
  NAND2X0 U12299 ( .IN1(n12163), .IN2(g1783), .QN(n12162) );
  NAND2X0 U12300 ( .IN1(n12164), .IN2(n10075), .QN(n12163) );
  NAND2X0 U12301 ( .IN1(n12165), .IN2(n10075), .QN(n12161) );
  NAND2X0 U12302 ( .IN1(n12166), .IN2(n12167), .QN(g26672) );
  NAND2X0 U12303 ( .IN1(n12168), .IN2(g2478), .QN(n12167) );
  NAND2X0 U12304 ( .IN1(n12159), .IN2(n10029), .QN(n12168) );
  NAND2X0 U12305 ( .IN1(n12160), .IN2(n10029), .QN(n12166) );
  NAND2X0 U12306 ( .IN1(n12169), .IN2(n12170), .QN(g26670) );
  NAND2X0 U12307 ( .IN1(n12171), .IN2(g1785), .QN(n12170) );
  NAND2X0 U12308 ( .IN1(n12164), .IN2(n10074), .QN(n12171) );
  NAND2X0 U12309 ( .IN1(n12165), .IN2(n10074), .QN(n12169) );
  NAND2X0 U12310 ( .IN1(n12172), .IN2(n12173), .QN(g26669) );
  NAND2X0 U12311 ( .IN1(n12174), .IN2(g1089), .QN(n12173) );
  NAND2X0 U12312 ( .IN1(n12175), .IN2(g1088), .QN(n12174) );
  NAND2X0 U12313 ( .IN1(n12176), .IN2(g1088), .QN(n12172) );
  NAND2X0 U12314 ( .IN1(n12177), .IN2(n12178), .QN(g26667) );
  NAND2X0 U12315 ( .IN1(test_so60), .IN2(n12179), .QN(n12178) );
  NAND2X0 U12316 ( .IN1(n12164), .IN2(n10076), .QN(n12179) );
  NAND2X0 U12317 ( .IN1(n12165), .IN2(n10076), .QN(n12177) );
  NOR2X0 U12318 ( .IN1(n12164), .IN2(n4386), .QN(n12165) );
  NOR3X0 U12319 ( .IN1(n10456), .IN2(n4386), .IN3(n10244), .QN(n12164) );
  NAND3X0 U12320 ( .IN1(n12180), .IN2(n12181), .IN3(n12182), .QN(n10244) );
  NAND2X0 U12321 ( .IN1(n7657), .IN2(n10074), .QN(n12182) );
  NAND2X0 U12322 ( .IN1(n7667), .IN2(n10075), .QN(n12181) );
  NAND2X0 U12323 ( .IN1(n10076), .IN2(n8111), .QN(n12180) );
  NAND4X0 U12324 ( .IN1(n12183), .IN2(n12184), .IN3(n12185), .IN4(n12186), 
        .QN(n10456) );
  NOR4X0 U12325 ( .IN1(n12187), .IN2(n12188), .IN3(n12189), .IN4(n12190), .QN(
        n12186) );
  XNOR2X1 U12326 ( .IN1(n4374), .IN2(n12191), .Q(n12190) );
  NAND3X0 U12327 ( .IN1(n12192), .IN2(n12193), .IN3(n12194), .QN(n12191) );
  NAND2X0 U12328 ( .IN1(n7895), .IN2(g6782), .QN(n12194) );
  NAND2X0 U12329 ( .IN1(g6573), .IN2(n8093), .QN(n12193) );
  NAND2X0 U12330 ( .IN1(n7530), .IN2(g1547), .QN(n12192) );
  XOR2X1 U12331 ( .IN1(g1481), .IN2(n12195), .Q(n12189) );
  NAND3X0 U12332 ( .IN1(n12196), .IN2(n12197), .IN3(n12198), .QN(n12195) );
  NAND2X0 U12333 ( .IN1(n7893), .IN2(g6782), .QN(n12198) );
  NAND2X0 U12334 ( .IN1(n7894), .IN2(g6573), .QN(n12197) );
  NAND2X0 U12335 ( .IN1(n7529), .IN2(g1547), .QN(n12196) );
  XOR2X1 U12336 ( .IN1(n9639), .IN2(n12199), .Q(n12188) );
  NAND3X0 U12337 ( .IN1(n12200), .IN2(n12201), .IN3(n12202), .QN(n12199) );
  NAND2X0 U12338 ( .IN1(n7506), .IN2(g6782), .QN(n12202) );
  NAND2X0 U12339 ( .IN1(n7507), .IN2(g6573), .QN(n12201) );
  NAND2X0 U12340 ( .IN1(n7505), .IN2(g1547), .QN(n12200) );
  NAND3X0 U12341 ( .IN1(n12203), .IN2(n3070), .IN3(n12204), .QN(n12187) );
  XOR2X1 U12342 ( .IN1(n12205), .IN2(n4378), .Q(n12204) );
  NAND3X0 U12343 ( .IN1(n12206), .IN2(n12207), .IN3(n12208), .QN(n12205) );
  NAND2X0 U12344 ( .IN1(n7896), .IN2(g6782), .QN(n12208) );
  NAND2X0 U12345 ( .IN1(n7897), .IN2(g6573), .QN(n12207) );
  NAND2X0 U12346 ( .IN1(n7531), .IN2(g1547), .QN(n12206) );
  XOR2X1 U12347 ( .IN1(n12209), .IN2(n9484), .Q(n12203) );
  NAND3X0 U12348 ( .IN1(n12210), .IN2(n12211), .IN3(n12212), .QN(n12209) );
  NAND2X0 U12349 ( .IN1(n7522), .IN2(g6782), .QN(n12212) );
  NAND2X0 U12350 ( .IN1(n7523), .IN2(g6573), .QN(n12211) );
  NAND2X0 U12351 ( .IN1(n7521), .IN2(g1547), .QN(n12210) );
  NOR3X0 U12352 ( .IN1(n12213), .IN2(n12214), .IN3(n12215), .QN(n12185) );
  XOR2X1 U12353 ( .IN1(g1501), .IN2(n12216), .Q(n12215) );
  NAND3X0 U12354 ( .IN1(n12217), .IN2(n12218), .IN3(n12219), .QN(n12216) );
  NAND2X0 U12355 ( .IN1(g6782), .IN2(n8112), .QN(n12219) );
  NAND2X0 U12356 ( .IN1(n7886), .IN2(g6573), .QN(n12218) );
  NAND2X0 U12357 ( .IN1(n7525), .IN2(g1547), .QN(n12217) );
  XOR2X1 U12358 ( .IN1(g1496), .IN2(n12220), .Q(n12214) );
  NAND3X0 U12359 ( .IN1(n12221), .IN2(n12222), .IN3(n12223), .QN(n12220) );
  NAND2X0 U12360 ( .IN1(n7887), .IN2(g6782), .QN(n12223) );
  NAND2X0 U12361 ( .IN1(n7888), .IN2(g6573), .QN(n12222) );
  NAND2X0 U12362 ( .IN1(n7526), .IN2(g1547), .QN(n12221) );
  XNOR2X1 U12363 ( .IN1(n4390), .IN2(n12224), .Q(n12213) );
  NAND3X0 U12364 ( .IN1(n12225), .IN2(n12226), .IN3(n12227), .QN(n12224) );
  NAND2X0 U12365 ( .IN1(n7891), .IN2(g6782), .QN(n12227) );
  NAND2X0 U12366 ( .IN1(n7892), .IN2(g6573), .QN(n12226) );
  NAND2X0 U12367 ( .IN1(n7528), .IN2(g1547), .QN(n12225) );
  XOR2X1 U12368 ( .IN1(n12228), .IN2(n4288), .Q(n12184) );
  NAND3X0 U12369 ( .IN1(n12229), .IN2(n12230), .IN3(n12231), .QN(n12228) );
  NAND2X0 U12370 ( .IN1(n7884), .IN2(g6782), .QN(n12231) );
  NAND2X0 U12371 ( .IN1(n7885), .IN2(g6573), .QN(n12230) );
  NAND2X0 U12372 ( .IN1(n7524), .IN2(g1547), .QN(n12229) );
  XOR2X1 U12373 ( .IN1(n12232), .IN2(n4326), .Q(n12183) );
  NAND3X0 U12374 ( .IN1(n12233), .IN2(n12234), .IN3(n12235), .QN(n12232) );
  NAND2X0 U12375 ( .IN1(n7889), .IN2(g6782), .QN(n12235) );
  NAND2X0 U12376 ( .IN1(n7890), .IN2(g6573), .QN(n12234) );
  NAND2X0 U12377 ( .IN1(n7527), .IN2(g1547), .QN(n12233) );
  NAND2X0 U12378 ( .IN1(n12236), .IN2(n12237), .QN(g26665) );
  NAND2X0 U12379 ( .IN1(n12238), .IN2(g1091), .QN(n12237) );
  NAND2X0 U12380 ( .IN1(n12175), .IN2(g6712), .QN(n12238) );
  NAND2X0 U12381 ( .IN1(n12176), .IN2(g6712), .QN(n12236) );
  NAND2X0 U12382 ( .IN1(n12239), .IN2(n12240), .QN(g26664) );
  NAND2X0 U12383 ( .IN1(n12241), .IN2(g402), .QN(n12240) );
  NAND2X0 U12384 ( .IN1(n12242), .IN2(n10160), .QN(n12241) );
  NAND2X0 U12385 ( .IN1(n12243), .IN2(n10160), .QN(n12239) );
  NAND2X0 U12386 ( .IN1(n12244), .IN2(n12245), .QN(g26661) );
  NAND2X0 U12387 ( .IN1(n12246), .IN2(g1090), .QN(n12245) );
  NAND2X0 U12388 ( .IN1(n12175), .IN2(g5472), .QN(n12246) );
  NAND2X0 U12389 ( .IN1(n12176), .IN2(g5472), .QN(n12244) );
  NOR2X0 U12390 ( .IN1(n12175), .IN2(n4387), .QN(n12176) );
  NOR3X0 U12391 ( .IN1(n10546), .IN2(n4387), .IN3(n10253), .QN(n12175) );
  NAND3X0 U12392 ( .IN1(n12247), .IN2(n12248), .IN3(n12249), .QN(n10253) );
  NAND2X0 U12393 ( .IN1(n7672), .IN2(g1088), .QN(n12249) );
  NAND2X0 U12394 ( .IN1(n7673), .IN2(g5472), .QN(n12248) );
  NAND2X0 U12395 ( .IN1(n7660), .IN2(g6712), .QN(n12247) );
  NAND4X0 U12396 ( .IN1(n12250), .IN2(n12251), .IN3(n12252), .IN4(n12253), 
        .QN(n10546) );
  NOR4X0 U12397 ( .IN1(n12254), .IN2(n12255), .IN3(n9200), .IN4(n12256), .QN(
        n12253) );
  XOR2X1 U12398 ( .IN1(n9668), .IN2(n12257), .Q(n12256) );
  NAND3X0 U12399 ( .IN1(n12258), .IN2(n12259), .IN3(n12260), .QN(n12257) );
  NAND2X0 U12400 ( .IN1(n7535), .IN2(test_so31), .QN(n12260) );
  NAND2X0 U12401 ( .IN1(n7536), .IN2(g6518), .QN(n12259) );
  NAND2X0 U12402 ( .IN1(n7537), .IN2(g6368), .QN(n12258) );
  INVX0 U12403 ( .INP(n3102), .ZN(n9200) );
  XOR2X1 U12404 ( .IN1(n10834), .IN2(n12261), .Q(n12255) );
  NAND3X0 U12405 ( .IN1(n12262), .IN2(n12263), .IN3(n12264), .QN(n12261) );
  NAND2X0 U12406 ( .IN1(n7532), .IN2(test_so31), .QN(n12264) );
  NAND2X0 U12407 ( .IN1(n7533), .IN2(g6518), .QN(n12263) );
  NAND2X0 U12408 ( .IN1(n7534), .IN2(g6368), .QN(n12262) );
  NAND3X0 U12409 ( .IN1(n12265), .IN2(n12266), .IN3(n12267), .QN(n12254) );
  XOR2X1 U12410 ( .IN1(n12268), .IN2(n4375), .Q(n12267) );
  NAND3X0 U12411 ( .IN1(n12269), .IN2(n12270), .IN3(n12271), .QN(n12268) );
  NAND2X0 U12412 ( .IN1(n7544), .IN2(test_so31), .QN(n12271) );
  NAND2X0 U12413 ( .IN1(n7911), .IN2(g6518), .QN(n12270) );
  NAND2X0 U12414 ( .IN1(n7914), .IN2(g6368), .QN(n12269) );
  XOR2X1 U12415 ( .IN1(n12272), .IN2(n4321), .Q(n12266) );
  NAND3X0 U12416 ( .IN1(n12273), .IN2(n12274), .IN3(n12275), .QN(n12272) );
  NAND2X0 U12417 ( .IN1(n7543), .IN2(test_so31), .QN(n12275) );
  NAND2X0 U12418 ( .IN1(n7908), .IN2(g6518), .QN(n12274) );
  NAND2X0 U12419 ( .IN1(n7910), .IN2(g6368), .QN(n12273) );
  XOR2X1 U12420 ( .IN1(n12276), .IN2(n4379), .Q(n12265) );
  NAND3X0 U12421 ( .IN1(n12277), .IN2(n12278), .IN3(n12279), .QN(n12276) );
  NAND2X0 U12422 ( .IN1(n7545), .IN2(test_so31), .QN(n12279) );
  NAND2X0 U12423 ( .IN1(n7915), .IN2(g6518), .QN(n12278) );
  NAND2X0 U12424 ( .IN1(n7916), .IN2(g6368), .QN(n12277) );
  NOR3X0 U12425 ( .IN1(n12280), .IN2(n12281), .IN3(n12282), .QN(n12252) );
  XOR2X1 U12426 ( .IN1(g809), .IN2(n12283), .Q(n12282) );
  NAND3X0 U12427 ( .IN1(n12284), .IN2(n12285), .IN3(n12286), .QN(n12283) );
  NAND2X0 U12428 ( .IN1(n7539), .IN2(test_so31), .QN(n12286) );
  NAND2X0 U12429 ( .IN1(n7900), .IN2(g6518), .QN(n12285) );
  NAND2X0 U12430 ( .IN1(n7901), .IN2(g6368), .QN(n12284) );
  XOR2X1 U12431 ( .IN1(g805), .IN2(n12287), .Q(n12281) );
  NAND3X0 U12432 ( .IN1(n12288), .IN2(n12289), .IN3(n12290), .QN(n12287) );
  NAND2X0 U12433 ( .IN1(n7540), .IN2(test_so31), .QN(n12290) );
  NAND2X0 U12434 ( .IN1(n7902), .IN2(g6518), .QN(n12289) );
  NAND2X0 U12435 ( .IN1(g6368), .IN2(n8113), .QN(n12288) );
  XNOR2X1 U12436 ( .IN1(n4391), .IN2(n12291), .Q(n12280) );
  NAND3X0 U12437 ( .IN1(n12292), .IN2(n12293), .IN3(n12294), .QN(n12291) );
  NAND2X0 U12438 ( .IN1(n7542), .IN2(test_so31), .QN(n12294) );
  NAND2X0 U12439 ( .IN1(n7905), .IN2(g6518), .QN(n12293) );
  NAND2X0 U12440 ( .IN1(n7906), .IN2(g6368), .QN(n12292) );
  XOR2X1 U12441 ( .IN1(n12295), .IN2(n4289), .Q(n12251) );
  NAND3X0 U12442 ( .IN1(n12296), .IN2(n12297), .IN3(n12298), .QN(n12295) );
  NAND2X0 U12443 ( .IN1(n7538), .IN2(test_so31), .QN(n12298) );
  NAND2X0 U12444 ( .IN1(n7898), .IN2(g6518), .QN(n12297) );
  NAND2X0 U12445 ( .IN1(n7899), .IN2(g6368), .QN(n12296) );
  XOR2X1 U12446 ( .IN1(n12299), .IN2(n4327), .Q(n12250) );
  NAND3X0 U12447 ( .IN1(n12300), .IN2(n12301), .IN3(n12302), .QN(n12299) );
  NAND2X0 U12448 ( .IN1(n7541), .IN2(test_so31), .QN(n12302) );
  NAND2X0 U12449 ( .IN1(n7903), .IN2(g6518), .QN(n12301) );
  NAND2X0 U12450 ( .IN1(n7904), .IN2(g6368), .QN(n12300) );
  NAND2X0 U12451 ( .IN1(n12303), .IN2(n12304), .QN(g26659) );
  NAND2X0 U12452 ( .IN1(n12305), .IN2(g404), .QN(n12304) );
  NAND2X0 U12453 ( .IN1(n12242), .IN2(n10159), .QN(n12305) );
  NAND2X0 U12454 ( .IN1(n12243), .IN2(n10159), .QN(n12303) );
  NAND2X0 U12455 ( .IN1(n12306), .IN2(n12307), .QN(g26655) );
  NAND2X0 U12456 ( .IN1(n12308), .IN2(g403), .QN(n12307) );
  NAND2X0 U12457 ( .IN1(n12242), .IN2(n10158), .QN(n12308) );
  NAND2X0 U12458 ( .IN1(n12243), .IN2(n10158), .QN(n12306) );
  NOR2X0 U12459 ( .IN1(n12242), .IN2(n4388), .QN(n12243) );
  NOR3X0 U12460 ( .IN1(n10635), .IN2(n4388), .IN3(n10264), .QN(n12242) );
  NAND3X0 U12461 ( .IN1(n12309), .IN2(n12310), .IN3(n12311), .QN(n10264) );
  NAND2X0 U12462 ( .IN1(n7680), .IN2(n10158), .QN(n12311) );
  NAND2X0 U12463 ( .IN1(n7679), .IN2(n10159), .QN(n12310) );
  NAND2X0 U12464 ( .IN1(n7678), .IN2(n10160), .QN(n12309) );
  NAND4X0 U12465 ( .IN1(n12312), .IN2(n12313), .IN3(n12314), .IN4(n12315), 
        .QN(n10635) );
  NOR4X0 U12466 ( .IN1(n12316), .IN2(n12317), .IN3(n12318), .IN4(n12319), .QN(
        n12315) );
  XNOR2X1 U12467 ( .IN1(n4376), .IN2(n12320), .Q(n12319) );
  NAND3X0 U12468 ( .IN1(n12321), .IN2(n12322), .IN3(n12323), .QN(n12320) );
  NAND2X0 U12469 ( .IN1(n7949), .IN2(g6313), .QN(n12323) );
  NAND2X0 U12470 ( .IN1(n7950), .IN2(g6231), .QN(n12322) );
  NAND2X0 U12471 ( .IN1(n7553), .IN2(g165), .QN(n12321) );
  XOR2X1 U12472 ( .IN1(g97), .IN2(n12324), .Q(n12318) );
  NAND3X0 U12473 ( .IN1(n12325), .IN2(n12326), .IN3(n12327), .QN(n12324) );
  NAND2X0 U12474 ( .IN1(n7951), .IN2(g6313), .QN(n12327) );
  NAND2X0 U12475 ( .IN1(n7952), .IN2(g6231), .QN(n12326) );
  NAND2X0 U12476 ( .IN1(n7554), .IN2(g165), .QN(n12325) );
  XOR2X1 U12477 ( .IN1(n10704), .IN2(n12328), .Q(n12317) );
  NAND3X0 U12478 ( .IN1(n12329), .IN2(n12330), .IN3(n12331), .QN(n12328) );
  NAND2X0 U12479 ( .IN1(n7547), .IN2(g6313), .QN(n12331) );
  NAND2X0 U12480 ( .IN1(g6231), .IN2(n8114), .QN(n12330) );
  NAND2X0 U12481 ( .IN1(n7546), .IN2(g165), .QN(n12329) );
  NAND3X0 U12482 ( .IN1(n12332), .IN2(n3130), .IN3(n12333), .QN(n12316) );
  XOR2X1 U12483 ( .IN1(n12334), .IN2(n4322), .Q(n12333) );
  NAND3X0 U12484 ( .IN1(n12335), .IN2(n12336), .IN3(n12337), .QN(n12334) );
  NAND2X0 U12485 ( .IN1(n7947), .IN2(g6313), .QN(n12337) );
  NAND2X0 U12486 ( .IN1(n7948), .IN2(g6231), .QN(n12336) );
  NAND2X0 U12487 ( .IN1(n7552), .IN2(g165), .QN(n12335) );
  XOR2X1 U12488 ( .IN1(n12338), .IN2(n12339), .Q(n12332) );
  NAND3X0 U12489 ( .IN1(n12340), .IN2(n12341), .IN3(n12342), .QN(n12338) );
  NAND2X0 U12490 ( .IN1(n7509), .IN2(g6313), .QN(n12342) );
  NAND2X0 U12491 ( .IN1(n7510), .IN2(g6231), .QN(n12341) );
  NAND2X0 U12492 ( .IN1(n7508), .IN2(g165), .QN(n12340) );
  NOR3X0 U12493 ( .IN1(n12343), .IN2(n12344), .IN3(n12345), .QN(n12314) );
  XNOR2X1 U12494 ( .IN1(n4569), .IN2(n12346), .Q(n12345) );
  NAND3X0 U12495 ( .IN1(n12347), .IN2(n12348), .IN3(n12349), .QN(n12346) );
  NAND2X0 U12496 ( .IN1(n7927), .IN2(g6313), .QN(n12349) );
  NAND2X0 U12497 ( .IN1(n7928), .IN2(g6231), .QN(n12348) );
  NAND2X0 U12498 ( .IN1(n7549), .IN2(g165), .QN(n12347) );
  XNOR2X1 U12499 ( .IN1(n4561), .IN2(n12350), .Q(n12344) );
  NAND3X0 U12500 ( .IN1(n12351), .IN2(n12352), .IN3(n12353), .QN(n12350) );
  NAND2X0 U12501 ( .IN1(n7931), .IN2(g6313), .QN(n12353) );
  NAND2X0 U12502 ( .IN1(n7932), .IN2(g6231), .QN(n12352) );
  NAND2X0 U12503 ( .IN1(n7550), .IN2(g165), .QN(n12351) );
  XNOR2X1 U12504 ( .IN1(n4392), .IN2(n12354), .Q(n12343) );
  NAND3X0 U12505 ( .IN1(n12355), .IN2(n12356), .IN3(n12357), .QN(n12354) );
  NAND2X0 U12506 ( .IN1(n7935), .IN2(g6313), .QN(n12357) );
  NAND2X0 U12507 ( .IN1(n7939), .IN2(g6231), .QN(n12356) );
  NAND2X0 U12508 ( .IN1(g165), .IN2(n8115), .QN(n12355) );
  XOR2X1 U12509 ( .IN1(n12358), .IN2(n4290), .Q(n12313) );
  NAND3X0 U12510 ( .IN1(n12359), .IN2(n12360), .IN3(n12361), .QN(n12358) );
  NAND2X0 U12511 ( .IN1(n7917), .IN2(g6313), .QN(n12361) );
  NAND2X0 U12512 ( .IN1(n7919), .IN2(g6231), .QN(n12360) );
  NAND2X0 U12513 ( .IN1(n7548), .IN2(g165), .QN(n12359) );
  XOR2X1 U12514 ( .IN1(n12362), .IN2(n4328), .Q(n12312) );
  NAND3X0 U12515 ( .IN1(n12363), .IN2(n12364), .IN3(n12365), .QN(n12362) );
  NAND2X0 U12516 ( .IN1(n7933), .IN2(g6313), .QN(n12365) );
  NAND2X0 U12517 ( .IN1(n7934), .IN2(g6231), .QN(n12364) );
  NAND2X0 U12518 ( .IN1(n7551), .IN2(g165), .QN(n12363) );
  NAND2X0 U12519 ( .IN1(n12366), .IN2(n12367), .QN(g26616) );
  NAND2X0 U12520 ( .IN1(n4299), .IN2(g2571), .QN(n12367) );
  NAND2X0 U12521 ( .IN1(n12368), .IN2(g2624), .QN(n12366) );
  NAND2X0 U12522 ( .IN1(n12369), .IN2(n12370), .QN(g26596) );
  NAND2X0 U12523 ( .IN1(n4370), .IN2(g2568), .QN(n12370) );
  NAND2X0 U12524 ( .IN1(n12368), .IN2(g7390), .QN(n12369) );
  NAND2X0 U12525 ( .IN1(n12371), .IN2(n12372), .QN(g26592) );
  NAND2X0 U12526 ( .IN1(n4366), .IN2(g1877), .QN(n12372) );
  NAND2X0 U12527 ( .IN1(n12373), .IN2(g1930), .QN(n12371) );
  NAND2X0 U12528 ( .IN1(n12374), .IN2(n12375), .QN(g26575) );
  NAND2X0 U12529 ( .IN1(n4314), .IN2(g2565), .QN(n12375) );
  NAND2X0 U12530 ( .IN1(n12368), .IN2(n10166), .QN(n12374) );
  NOR3X0 U12531 ( .IN1(n8876), .IN2(n4303), .IN3(n12376), .QN(n12368) );
  NAND2X0 U12532 ( .IN1(n12377), .IN2(n12378), .QN(g26573) );
  NAND2X0 U12533 ( .IN1(n4315), .IN2(g1874), .QN(n12378) );
  NAND2X0 U12534 ( .IN1(n12373), .IN2(g7194), .QN(n12377) );
  NAND2X0 U12535 ( .IN1(n12379), .IN2(n12380), .QN(g26569) );
  NAND2X0 U12536 ( .IN1(n4300), .IN2(g1183), .QN(n12380) );
  NAND2X0 U12537 ( .IN1(n12381), .IN2(g1236), .QN(n12379) );
  NAND2X0 U12538 ( .IN1(n12382), .IN2(n12383), .QN(g26559) );
  NAND2X0 U12539 ( .IN1(n12373), .IN2(n10214), .QN(n12383) );
  NOR3X0 U12540 ( .IN1(n9002), .IN2(n4297), .IN3(n12384), .QN(n12373) );
  NAND2X0 U12541 ( .IN1(test_so68), .IN2(n4296), .QN(n12382) );
  NAND2X0 U12542 ( .IN1(n12385), .IN2(n12386), .QN(g26557) );
  NAND2X0 U12543 ( .IN1(n4316), .IN2(g1180), .QN(n12386) );
  NAND2X0 U12544 ( .IN1(n12381), .IN2(g6944), .QN(n12385) );
  NAND2X0 U12545 ( .IN1(n12387), .IN2(n12388), .QN(g26553) );
  NAND2X0 U12546 ( .IN1(n4313), .IN2(g496), .QN(n12388) );
  NAND2X0 U12547 ( .IN1(n12389), .IN2(g550), .QN(n12387) );
  NAND2X0 U12548 ( .IN1(n12390), .IN2(n12391), .QN(g26547) );
  NAND2X0 U12549 ( .IN1(n12381), .IN2(n11104), .QN(n12391) );
  NOR3X0 U12550 ( .IN1(n9108), .IN2(n4304), .IN3(n12392), .QN(n12381) );
  NAND2X0 U12551 ( .IN1(test_so47), .IN2(n4371), .QN(n12390) );
  NAND2X0 U12552 ( .IN1(n12393), .IN2(n12394), .QN(g26545) );
  NAND2X0 U12553 ( .IN1(n4372), .IN2(g493), .QN(n12394) );
  NAND2X0 U12554 ( .IN1(n12389), .IN2(g6642), .QN(n12393) );
  NAND2X0 U12555 ( .IN1(n12395), .IN2(n12396), .QN(g26541) );
  NAND2X0 U12556 ( .IN1(n4298), .IN2(g490), .QN(n12396) );
  NAND2X0 U12557 ( .IN1(n12389), .IN2(n11207), .QN(n12395) );
  NOR3X0 U12558 ( .IN1(n8091), .IN2(n8751), .IN3(n12397), .QN(n12389) );
  NOR2X0 U12559 ( .IN1(n10265), .IN2(n12398), .QN(g26532) );
  XOR2X1 U12560 ( .IN1(n12399), .IN2(n7689), .Q(n12398) );
  NOR2X0 U12561 ( .IN1(n10267), .IN2(n12400), .QN(g26531) );
  XOR2X1 U12562 ( .IN1(n12401), .IN2(n7693), .Q(n12400) );
  NOR2X0 U12563 ( .IN1(n10269), .IN2(n12402), .QN(g26530) );
  XNOR2X1 U12564 ( .IN1(n7697), .IN2(n3690), .Q(n12402) );
  NAND2X0 U12565 ( .IN1(n3893), .IN2(g776), .QN(n3690) );
  NOR2X0 U12566 ( .IN1(n10271), .IN2(n12403), .QN(g26529) );
  XOR2X1 U12567 ( .IN1(n12404), .IN2(n7701), .Q(n12403) );
  NAND4X0 U12568 ( .IN1(n3700), .IN2(n12405), .IN3(n12406), .IN4(n12407), .QN(
        g26149) );
  NOR4X0 U12569 ( .IN1(n12408), .IN2(n12409), .IN3(n12410), .IN4(n12411), .QN(
        n12407) );
  NOR2X0 U12570 ( .IN1(n4441), .IN2(n12412), .QN(n12411) );
  NOR2X0 U12571 ( .IN1(n4338), .IN2(n12413), .QN(n12410) );
  NOR2X0 U12572 ( .IN1(n11433), .IN2(DFF_156_n1), .QN(n12409) );
  NAND3X0 U12573 ( .IN1(n12414), .IN2(n12415), .IN3(n12416), .QN(n12408) );
  NAND2X0 U12574 ( .IN1(n3936), .IN2(n12417), .QN(n12416) );
  NAND4X0 U12575 ( .IN1(n12418), .IN2(n12419), .IN3(n12420), .IN4(n12421), 
        .QN(n12417) );
  NAND2X0 U12576 ( .IN1(n12422), .IN2(g3088), .QN(n12421) );
  NAND2X0 U12577 ( .IN1(n12423), .IN2(g3164), .QN(n12420) );
  NAND2X0 U12578 ( .IN1(n12424), .IN2(g3158), .QN(n12419) );
  NAND2X0 U12579 ( .IN1(n12425), .IN2(g3182), .QN(n12418) );
  NAND2X0 U12580 ( .IN1(n12426), .IN2(g3167), .QN(n12415) );
  NAND2X0 U12581 ( .IN1(n3939), .IN2(n12427), .QN(n12414) );
  NAND3X0 U12582 ( .IN1(n12428), .IN2(n12429), .IN3(n12430), .QN(n12427) );
  NAND2X0 U12583 ( .IN1(n3940), .IN2(g3185), .QN(n12430) );
  NAND2X0 U12584 ( .IN1(test_so8), .IN2(n12431), .QN(n12429) );
  NAND2X0 U12585 ( .IN1(n12432), .IN2(g3155), .QN(n12428) );
  NOR3X0 U12586 ( .IN1(n12433), .IN2(n12434), .IN3(n12435), .QN(n12406) );
  NOR2X0 U12587 ( .IN1(n4444), .IN2(n12436), .QN(n12435) );
  NOR2X0 U12588 ( .IN1(n4450), .IN2(n12437), .QN(n12434) );
  NOR2X0 U12589 ( .IN1(n12438), .IN2(DFF_149_n1), .QN(n12433) );
  NAND2X0 U12590 ( .IN1(n11434), .IN2(n8086), .QN(n12405) );
  NAND4X0 U12591 ( .IN1(n12439), .IN2(n3700), .IN3(n12440), .IN4(n12441), .QN(
        g26135) );
  NOR4X0 U12592 ( .IN1(n12442), .IN2(n12443), .IN3(n12444), .IN4(n12445), .QN(
        n12441) );
  NOR2X0 U12593 ( .IN1(n4447), .IN2(n12413), .QN(n12445) );
  NOR2X0 U12594 ( .IN1(n12446), .IN2(n12447), .QN(n12444) );
  INVX0 U12595 ( .INP(n3936), .ZN(n12447) );
  NOR4X0 U12596 ( .IN1(n12448), .IN2(n12449), .IN3(n12450), .IN4(n12451), .QN(
        n12446) );
  NOR2X0 U12597 ( .IN1(n4438), .IN2(n11424), .QN(n12451) );
  INVX0 U12598 ( .INP(n12452), .ZN(n12450) );
  NAND2X0 U12599 ( .IN1(g3098), .IN2(n12424), .QN(n12452) );
  NOR2X0 U12600 ( .IN1(n4342), .IN2(n12453), .QN(n12449) );
  INVX0 U12601 ( .INP(n12423), .ZN(n12453) );
  NOR2X0 U12602 ( .IN1(n4334), .IN2(n12454), .QN(n12448) );
  INVX0 U12603 ( .INP(n12422), .ZN(n12454) );
  NOR2X0 U12604 ( .IN1(n4343), .IN2(n12412), .QN(n12443) );
  NAND4X0 U12605 ( .IN1(n12455), .IN2(n12456), .IN3(n12457), .IN4(n12458), 
        .QN(n12442) );
  NAND2X0 U12606 ( .IN1(test_so10), .IN2(n12459), .QN(n12458) );
  NAND2X0 U12607 ( .IN1(test_so7), .IN2(n12426), .QN(n12457) );
  NAND2X0 U12608 ( .IN1(n11418), .IN2(n12460), .QN(n12456) );
  INVX0 U12609 ( .INP(n12461), .ZN(n11418) );
  NAND2X0 U12610 ( .IN1(n3939), .IN2(n12462), .QN(n12455) );
  NAND3X0 U12611 ( .IN1(n12463), .IN2(n12464), .IN3(n12465), .QN(n12462) );
  NAND2X0 U12612 ( .IN1(n3940), .IN2(g3107), .QN(n12465) );
  NAND2X0 U12613 ( .IN1(n12431), .IN2(g3105), .QN(n12464) );
  NAND2X0 U12614 ( .IN1(n12432), .IN2(g3097), .QN(n12463) );
  NOR3X0 U12615 ( .IN1(n12466), .IN2(n12467), .IN3(n12468), .QN(n12440) );
  NOR2X0 U12616 ( .IN1(n4452), .IN2(n12437), .QN(n12468) );
  NOR2X0 U12617 ( .IN1(n11433), .IN2(DFF_155_n1), .QN(n12467) );
  NOR2X0 U12618 ( .IN1(n4443), .IN2(n12436), .QN(n12466) );
  NOR2X0 U12619 ( .IN1(n12469), .IN2(n12470), .QN(n12439) );
  NOR2X0 U12620 ( .IN1(n12471), .IN2(g3128), .QN(n12470) );
  NOR2X0 U12621 ( .IN1(n14351), .IN2(n12438), .QN(n12469) );
  NAND4X0 U12622 ( .IN1(n12472), .IN2(n3700), .IN3(n12473), .IN4(n12474), .QN(
        g26104) );
  NOR4X0 U12623 ( .IN1(n12475), .IN2(n12476), .IN3(n12477), .IN4(n12478), .QN(
        n12474) );
  NOR2X0 U12624 ( .IN1(n4448), .IN2(n12413), .QN(n12478) );
  NAND3X0 U12625 ( .IN1(n12479), .IN2(n4406), .IN3(n3933), .QN(n12413) );
  NOR2X0 U12626 ( .IN1(n11431), .IN2(n12461), .QN(n12477) );
  NAND2X0 U12627 ( .IN1(n3705), .IN2(n12432), .QN(n12461) );
  INVX0 U12628 ( .INP(n12480), .ZN(n11431) );
  NOR2X0 U12629 ( .IN1(n4344), .IN2(n12412), .QN(n12476) );
  NAND2X0 U12630 ( .IN1(n12481), .IN2(n4329), .QN(n12412) );
  NAND4X0 U12631 ( .IN1(n12482), .IN2(n12483), .IN3(n12484), .IN4(n12485), 
        .QN(n12475) );
  NAND2X0 U12632 ( .IN1(n12459), .IN2(g3142), .QN(n12485) );
  INVX0 U12633 ( .INP(n11422), .ZN(n12459) );
  NAND3X0 U12634 ( .IN1(n3940), .IN2(g3204), .IN3(n4073), .QN(n11422) );
  NAND2X0 U12635 ( .IN1(n12426), .IN2(g3086), .QN(n12484) );
  NOR2X0 U12636 ( .IN1(n11426), .IN2(n12486), .QN(n12426) );
  NAND2X0 U12637 ( .IN1(n3939), .IN2(n12487), .QN(n12483) );
  NAND3X0 U12638 ( .IN1(n12488), .IN2(n12489), .IN3(n12490), .QN(n12487) );
  NAND2X0 U12639 ( .IN1(n3940), .IN2(g3095), .QN(n12490) );
  NAND2X0 U12640 ( .IN1(n12431), .IN2(g3093), .QN(n12489) );
  NAND2X0 U12641 ( .IN1(test_so6), .IN2(n12432), .QN(n12488) );
  NAND2X0 U12642 ( .IN1(n3936), .IN2(n12491), .QN(n12482) );
  NAND4X0 U12643 ( .IN1(n12492), .IN2(n12493), .IN3(n12494), .IN4(n12495), 
        .QN(n12491) );
  NAND2X0 U12644 ( .IN1(n12422), .IN2(g3096), .QN(n12495) );
  NOR2X0 U12645 ( .IN1(n4329), .IN2(n4406), .QN(n12422) );
  NAND2X0 U12646 ( .IN1(n12423), .IN2(g3085), .QN(n12494) );
  NOR2X0 U12647 ( .IN1(g3201), .IN2(n4329), .QN(n12423) );
  NAND2X0 U12648 ( .IN1(n12424), .IN2(g3211), .QN(n12493) );
  NAND2X0 U12649 ( .IN1(n12425), .IN2(g3094), .QN(n12492) );
  NOR3X0 U12650 ( .IN1(n12496), .IN2(n12497), .IN3(n12498), .QN(n12473) );
  NOR2X0 U12651 ( .IN1(n4451), .IN2(n12437), .QN(n12498) );
  NAND2X0 U12652 ( .IN1(n12481), .IN2(g3207), .QN(n12437) );
  NOR3X0 U12653 ( .IN1(g3201), .IN2(n4405), .IN3(n11426), .QN(n12481) );
  INVX0 U12654 ( .INP(n12479), .ZN(n11426) );
  NOR2X0 U12655 ( .IN1(n9153), .IN2(n8015), .QN(n12479) );
  NAND2X0 U12656 ( .IN1(n266), .IN2(g3197), .QN(n9153) );
  INVX0 U12657 ( .INP(n12499), .ZN(n266) );
  NAND3X0 U12658 ( .IN1(DFF_132_n1), .IN2(DFF_131_n1), .IN3(DFF_134_n1), .QN(
        n12499) );
  NOR2X0 U12659 ( .IN1(n14353), .IN2(n11433), .QN(n12497) );
  NAND3X0 U12660 ( .IN1(n12431), .IN2(g3204), .IN3(n4073), .QN(n11433) );
  INVX0 U12661 ( .INP(n11429), .ZN(n12431) );
  NAND2X0 U12662 ( .IN1(n12425), .IN2(n4405), .QN(n11429) );
  INVX0 U12663 ( .INP(n11424), .ZN(n12425) );
  NAND2X0 U12664 ( .IN1(n4329), .IN2(g3201), .QN(n11424) );
  NOR2X0 U12665 ( .IN1(n4445), .IN2(n12436), .QN(n12496) );
  NAND3X0 U12666 ( .IN1(n3939), .IN2(n4406), .IN3(n3933), .QN(n12436) );
  NOR2X0 U12667 ( .IN1(g3188), .IN2(n4329), .QN(n3933) );
  NOR2X0 U12668 ( .IN1(n12500), .IN2(n12501), .QN(n12472) );
  NOR2X0 U12669 ( .IN1(n12471), .IN2(DFF_140_n1), .QN(n12501) );
  NOR2X0 U12670 ( .IN1(n14349), .IN2(n12438), .QN(n12500) );
  NAND2X0 U12671 ( .IN1(n8726), .IN2(n12502), .QN(g26048) );
  NAND2X0 U12672 ( .IN1(n12503), .IN2(n9283), .QN(n12502) );
  XOR2X1 U12673 ( .IN1(n7909), .IN2(n9286), .Q(n12503) );
  NOR2X0 U12674 ( .IN1(n8672), .IN2(n12504), .QN(g26037) );
  XOR2X1 U12675 ( .IN1(n4291), .IN2(n12148), .Q(n12504) );
  NOR2X0 U12676 ( .IN1(n12505), .IN2(n12153), .QN(g26031) );
  XOR2X1 U12677 ( .IN1(test_so98), .IN2(n3742), .Q(n12505) );
  NAND2X0 U12678 ( .IN1(n4065), .IN2(g3013), .QN(n3742) );
  NAND2X0 U12679 ( .IN1(n12506), .IN2(n12507), .QN(g26025) );
  NAND2X0 U12680 ( .IN1(test_so82), .IN2(n12508), .QN(n12507) );
  NAND2X0 U12681 ( .IN1(n12159), .IN2(n10028), .QN(n12508) );
  NAND2X0 U12682 ( .IN1(n12160), .IN2(n10028), .QN(n12506) );
  NOR2X0 U12683 ( .IN1(n8075), .IN2(n12159), .QN(n12160) );
  NOR3X0 U12684 ( .IN1(n8075), .IN2(n10365), .IN3(n10231), .QN(n12159) );
  NAND3X0 U12685 ( .IN1(n12509), .IN2(n12510), .IN3(n12511), .QN(n10231) );
  NAND2X0 U12686 ( .IN1(n7654), .IN2(n10027), .QN(n12511) );
  NAND2X0 U12687 ( .IN1(n10028), .IN2(n8116), .QN(n12510) );
  NAND2X0 U12688 ( .IN1(n7663), .IN2(n10029), .QN(n12509) );
  NAND4X0 U12689 ( .IN1(n12512), .IN2(n12513), .IN3(n12514), .IN4(n12515), 
        .QN(n10365) );
  NOR4X0 U12690 ( .IN1(n12516), .IN2(n12517), .IN3(n12518), .IN4(n12519), .QN(
        n12515) );
  XOR2X1 U12691 ( .IN1(g2170), .IN2(n12520), .Q(n12519) );
  NAND3X0 U12692 ( .IN1(n12521), .IN2(n12522), .IN3(n12523), .QN(n12520) );
  NAND2X0 U12693 ( .IN1(n7880), .IN2(test_so73), .QN(n12523) );
  NAND2X0 U12694 ( .IN1(n7881), .IN2(g6837), .QN(n12522) );
  NAND2X0 U12695 ( .IN1(n7519), .IN2(g2241), .QN(n12521) );
  XOR2X1 U12696 ( .IN1(g2165), .IN2(n12524), .Q(n12518) );
  NAND3X0 U12697 ( .IN1(n12525), .IN2(n12526), .IN3(n12527), .QN(n12524) );
  NAND2X0 U12698 ( .IN1(n7882), .IN2(test_so73), .QN(n12527) );
  NAND2X0 U12699 ( .IN1(n7883), .IN2(g6837), .QN(n12526) );
  NAND2X0 U12700 ( .IN1(n7520), .IN2(g2241), .QN(n12525) );
  XOR2X1 U12701 ( .IN1(n10762), .IN2(n12528), .Q(n12517) );
  NAND3X0 U12702 ( .IN1(n12529), .IN2(n12530), .IN3(n12531), .QN(n12528) );
  NAND2X0 U12703 ( .IN1(test_so73), .IN2(n8117), .QN(n12531) );
  NAND2X0 U12704 ( .IN1(n7512), .IN2(g6837), .QN(n12530) );
  NAND2X0 U12705 ( .IN1(n7511), .IN2(g2241), .QN(n12529) );
  NAND3X0 U12706 ( .IN1(n12532), .IN2(n3038), .IN3(n12533), .QN(n12516) );
  XOR2X1 U12707 ( .IN1(n12534), .IN2(n4319), .Q(n12533) );
  NAND3X0 U12708 ( .IN1(n12535), .IN2(n12536), .IN3(n12537), .QN(n12534) );
  NAND2X0 U12709 ( .IN1(n7878), .IN2(test_so73), .QN(n12537) );
  NAND2X0 U12710 ( .IN1(n7879), .IN2(g6837), .QN(n12536) );
  NAND2X0 U12711 ( .IN1(n7518), .IN2(g2241), .QN(n12535) );
  XOR2X1 U12712 ( .IN1(n12538), .IN2(n10437), .Q(n12532) );
  NAND3X0 U12713 ( .IN1(n12539), .IN2(n12540), .IN3(n12541), .QN(n12538) );
  NAND2X0 U12714 ( .IN1(n7503), .IN2(test_so73), .QN(n12541) );
  NAND2X0 U12715 ( .IN1(n7504), .IN2(g6837), .QN(n12540) );
  NAND2X0 U12716 ( .IN1(n7502), .IN2(g2241), .QN(n12539) );
  NOR3X0 U12717 ( .IN1(n12542), .IN2(n12543), .IN3(n12544), .QN(n12514) );
  XOR2X1 U12718 ( .IN1(g2195), .IN2(n12545), .Q(n12544) );
  NAND3X0 U12719 ( .IN1(n12546), .IN2(n12547), .IN3(n12548), .QN(n12545) );
  NAND2X0 U12720 ( .IN1(n7871), .IN2(test_so73), .QN(n12548) );
  NAND2X0 U12721 ( .IN1(n7872), .IN2(g6837), .QN(n12547) );
  NAND2X0 U12722 ( .IN1(n7514), .IN2(g2241), .QN(n12546) );
  XOR2X1 U12723 ( .IN1(g2190), .IN2(n12549), .Q(n12543) );
  NAND3X0 U12724 ( .IN1(n12550), .IN2(n12551), .IN3(n12552), .QN(n12549) );
  NAND2X0 U12725 ( .IN1(n7873), .IN2(test_so73), .QN(n12552) );
  NAND2X0 U12726 ( .IN1(n7874), .IN2(g6837), .QN(n12551) );
  NAND2X0 U12727 ( .IN1(n7515), .IN2(g2241), .QN(n12550) );
  XOR2X1 U12728 ( .IN1(g2180), .IN2(n12553), .Q(n12542) );
  NAND3X0 U12729 ( .IN1(n12554), .IN2(n12555), .IN3(n12556), .QN(n12553) );
  NAND2X0 U12730 ( .IN1(n7876), .IN2(test_so73), .QN(n12556) );
  NAND2X0 U12731 ( .IN1(n7877), .IN2(g6837), .QN(n12555) );
  NAND2X0 U12732 ( .IN1(n7517), .IN2(g2241), .QN(n12554) );
  XOR2X1 U12733 ( .IN1(n12557), .IN2(n4287), .Q(n12513) );
  NAND3X0 U12734 ( .IN1(n12558), .IN2(n12559), .IN3(n12560), .QN(n12557) );
  NAND2X0 U12735 ( .IN1(n7869), .IN2(test_so73), .QN(n12560) );
  NAND2X0 U12736 ( .IN1(n7870), .IN2(g6837), .QN(n12559) );
  NAND2X0 U12737 ( .IN1(n7513), .IN2(g2241), .QN(n12558) );
  XOR2X1 U12738 ( .IN1(n12561), .IN2(n4325), .Q(n12512) );
  NAND3X0 U12739 ( .IN1(n12562), .IN2(n12563), .IN3(n12564), .QN(n12561) );
  NAND2X0 U12740 ( .IN1(test_so73), .IN2(n8118), .QN(n12564) );
  NAND2X0 U12741 ( .IN1(n7875), .IN2(g6837), .QN(n12563) );
  NAND2X0 U12742 ( .IN1(n7516), .IN2(g2241), .QN(n12562) );
  NOR3X0 U12743 ( .IN1(n12399), .IN2(n10265), .IN3(n12565), .QN(g25940) );
  NOR2X0 U12744 ( .IN1(n3887), .IN2(test_so78), .QN(n12565) );
  INVX0 U12745 ( .INP(n4526), .ZN(n12399) );
  NOR3X0 U12746 ( .IN1(n12401), .IN2(n10267), .IN3(n12566), .QN(g25938) );
  NOR2X0 U12747 ( .IN1(n3890), .IN2(g1462), .QN(n12566) );
  INVX0 U12748 ( .INP(n4527), .ZN(n12401) );
  NOR2X0 U12749 ( .IN1(n10269), .IN2(n12567), .QN(g25935) );
  XOR2X1 U12750 ( .IN1(n8054), .IN2(n3893), .Q(n12567) );
  NOR3X0 U12751 ( .IN1(n12404), .IN2(n10271), .IN3(n12568), .QN(g25932) );
  NOR2X0 U12752 ( .IN1(n3896), .IN2(g88), .QN(n12568) );
  INVX0 U12753 ( .INP(n4528), .ZN(n12404) );
  NAND2X0 U12754 ( .IN1(n12569), .IN2(n12570), .QN(g25489) );
  NAND2X0 U12755 ( .IN1(n12571), .IN2(n8095), .QN(n12570) );
  NAND2X0 U12756 ( .IN1(n12572), .IN2(n12573), .QN(n12571) );
  NAND2X0 U12757 ( .IN1(n4424), .IN2(n12574), .QN(n12573) );
  NAND2X0 U12758 ( .IN1(n11430), .IN2(g3142), .QN(n12574) );
  INVX0 U12759 ( .INP(n12460), .ZN(n11430) );
  NAND2X0 U12760 ( .IN1(n7432), .IN2(n7431), .QN(n12460) );
  NAND2X0 U12761 ( .IN1(n4301), .IN2(n12480), .QN(n12572) );
  NAND2X0 U12762 ( .IN1(DFF_15_n1), .IN2(DFF_16_n1), .QN(n12480) );
  NAND4X0 U12763 ( .IN1(g3151), .IN2(g3097), .IN3(g3142), .IN4(test_so10), 
        .QN(n12569) );
  NAND2X0 U12764 ( .IN1(n12575), .IN2(n12576), .QN(g25452) );
  NAND2X0 U12765 ( .IN1(n4494), .IN2(g3099), .QN(n12576) );
  NAND2X0 U12766 ( .IN1(g21851), .IN2(g3109), .QN(n12575) );
  NAND2X0 U12767 ( .IN1(n12577), .IN2(n12578), .QN(g25451) );
  NAND2X0 U12768 ( .IN1(n4383), .IN2(g3098), .QN(n12578) );
  NAND2X0 U12769 ( .IN1(g21851), .IN2(g8030), .QN(n12577) );
  NAND2X0 U12770 ( .IN1(n12579), .IN2(n12580), .QN(g25450) );
  NAND2X0 U12771 ( .IN1(n4382), .IN2(g3097), .QN(n12580) );
  NAND2X0 U12772 ( .IN1(g21851), .IN2(g8106), .QN(n12579) );
  NAND3X0 U12773 ( .IN1(n12581), .IN2(n12582), .IN3(n3700), .QN(g25442) );
  NAND2X0 U12774 ( .IN1(n12583), .IN2(g3111), .QN(n12582) );
  NAND2X0 U12775 ( .IN1(n11434), .IN2(g3124), .QN(n12581) );
  NAND3X0 U12776 ( .IN1(n12584), .IN2(n12585), .IN3(n3700), .QN(g25435) );
  NAND2X0 U12777 ( .IN1(n12583), .IN2(g3110), .QN(n12585) );
  NAND2X0 U12778 ( .IN1(n11434), .IN2(DFF_144_n1), .QN(n12584) );
  NAND3X0 U12779 ( .IN1(n12586), .IN2(n12587), .IN3(n3700), .QN(g25420) );
  NAND2X0 U12780 ( .IN1(n12583), .IN2(g3112), .QN(n12587) );
  INVX0 U12781 ( .INP(n12438), .ZN(n12583) );
  NAND3X0 U12782 ( .IN1(n12432), .IN2(g3204), .IN3(n4073), .QN(n12438) );
  INVX0 U12783 ( .INP(n12486), .ZN(n12432) );
  NAND2X0 U12784 ( .IN1(n4405), .IN2(n12424), .QN(n12486) );
  NOR2X0 U12785 ( .IN1(g3201), .IN2(g3207), .QN(n12424) );
  NAND2X0 U12786 ( .IN1(test_so9), .IN2(n11434), .QN(n12586) );
  NAND2X0 U12787 ( .IN1(n12588), .IN2(n12589), .QN(g25288) );
  NAND2X0 U12788 ( .IN1(n12590), .IN2(g2808), .QN(n12589) );
  NAND2X0 U12789 ( .IN1(n12591), .IN2(n12592), .QN(n12588) );
  NAND2X0 U12790 ( .IN1(n12593), .IN2(n12594), .QN(g25280) );
  NAND2X0 U12791 ( .IN1(n12595), .IN2(g2810), .QN(n12594) );
  NAND2X0 U12792 ( .IN1(n12596), .IN2(n12591), .QN(n12593) );
  NAND2X0 U12793 ( .IN1(n12597), .IN2(n12598), .QN(g25279) );
  NAND2X0 U12794 ( .IN1(n12599), .IN2(g2114), .QN(n12598) );
  NAND2X0 U12795 ( .IN1(n12600), .IN2(n12601), .QN(n12597) );
  NAND2X0 U12796 ( .IN1(n12602), .IN2(n12603), .QN(g25272) );
  NAND2X0 U12797 ( .IN1(n12604), .IN2(g2809), .QN(n12603) );
  NAND2X0 U12798 ( .IN1(n12605), .IN2(n12591), .QN(n12602) );
  INVX0 U12799 ( .INP(n12606), .ZN(n12591) );
  NAND4X0 U12800 ( .IN1(n9243), .IN2(n12607), .IN3(n12608), .IN4(n12609), .QN(
        n12606) );
  NAND2X0 U12801 ( .IN1(n8029), .IN2(g7425), .QN(n12609) );
  NOR2X0 U12802 ( .IN1(n12610), .IN2(n12611), .QN(n12608) );
  NOR2X0 U12803 ( .IN1(n4292), .IN2(g2802), .QN(n12611) );
  NOR4X0 U12804 ( .IN1(n12612), .IN2(n12613), .IN3(n12614), .IN4(n12615), .QN(
        n12610) );
  XNOR2X1 U12805 ( .IN1(n4419), .IN2(n8900), .Q(n12615) );
  NAND3X0 U12806 ( .IN1(n12616), .IN2(n12617), .IN3(n12618), .QN(n8900) );
  NAND2X0 U12807 ( .IN1(n7767), .IN2(g7487), .QN(n12618) );
  NAND2X0 U12808 ( .IN1(n7832), .IN2(g2703), .QN(n12617) );
  NAND2X0 U12809 ( .IN1(n7768), .IN2(g7425), .QN(n12616) );
  XOR2X1 U12810 ( .IN1(n4471), .IN2(n8864), .Q(n12614) );
  INVX0 U12811 ( .INP(n8867), .ZN(n8864) );
  NAND3X0 U12812 ( .IN1(n12619), .IN2(n12620), .IN3(n12621), .QN(n8867) );
  NAND2X0 U12813 ( .IN1(n7757), .IN2(g7487), .QN(n12621) );
  NAND2X0 U12814 ( .IN1(n7828), .IN2(g2703), .QN(n12620) );
  NAND2X0 U12815 ( .IN1(n7758), .IN2(g7425), .QN(n12619) );
  NAND3X0 U12816 ( .IN1(n12622), .IN2(n12623), .IN3(n12624), .QN(n12613) );
  XOR2X1 U12817 ( .IN1(g2734), .IN2(n8875), .Q(n12624) );
  INVX0 U12818 ( .INP(n8878), .ZN(n8875) );
  NAND3X0 U12819 ( .IN1(n12625), .IN2(n12626), .IN3(n12627), .QN(n8878) );
  NAND2X0 U12820 ( .IN1(n7763), .IN2(g7487), .QN(n12627) );
  NAND2X0 U12821 ( .IN1(n7831), .IN2(g2703), .QN(n12626) );
  NAND2X0 U12822 ( .IN1(n7764), .IN2(g7425), .QN(n12625) );
  XOR2X1 U12823 ( .IN1(g2714), .IN2(n8886), .Q(n12623) );
  INVX0 U12824 ( .INP(n8887), .ZN(n8886) );
  NAND3X0 U12825 ( .IN1(n12628), .IN2(n12629), .IN3(n12630), .QN(n8887) );
  NAND2X0 U12826 ( .IN1(n7771), .IN2(g7487), .QN(n12630) );
  NAND2X0 U12827 ( .IN1(n7834), .IN2(g2703), .QN(n12629) );
  NAND2X0 U12828 ( .IN1(n7772), .IN2(g7425), .QN(n12628) );
  XOR2X1 U12829 ( .IN1(g2720), .IN2(n8881), .Q(n12622) );
  INVX0 U12830 ( .INP(n8882), .ZN(n8881) );
  NAND3X0 U12831 ( .IN1(n12631), .IN2(n12632), .IN3(n12633), .QN(n8882) );
  NAND2X0 U12832 ( .IN1(n7765), .IN2(g7487), .QN(n12633) );
  NAND2X0 U12833 ( .IN1(g2703), .IN2(n8119), .QN(n12632) );
  NAND2X0 U12834 ( .IN1(n7766), .IN2(g7425), .QN(n12631) );
  NAND4X0 U12835 ( .IN1(n12634), .IN2(n12635), .IN3(n12636), .IN4(n12637), 
        .QN(n12612) );
  XOR2X1 U12836 ( .IN1(g2707), .IN2(n8871), .Q(n12637) );
  INVX0 U12837 ( .INP(n8872), .ZN(n8871) );
  NAND3X0 U12838 ( .IN1(n12638), .IN2(n12639), .IN3(n12640), .QN(n8872) );
  NAND2X0 U12839 ( .IN1(n7769), .IN2(g7487), .QN(n12640) );
  NAND2X0 U12840 ( .IN1(n7833), .IN2(g2703), .QN(n12639) );
  NAND2X0 U12841 ( .IN1(n7770), .IN2(g7425), .QN(n12638) );
  NOR2X0 U12842 ( .IN1(n12641), .IN2(n12642), .QN(n12636) );
  XOR2X1 U12843 ( .IN1(n4393), .IN2(n8918), .Q(n12642) );
  INVX0 U12844 ( .INP(n8919), .ZN(n8918) );
  NAND3X0 U12845 ( .IN1(n12643), .IN2(n12644), .IN3(n12645), .QN(n8919) );
  NAND2X0 U12846 ( .IN1(n7755), .IN2(g7487), .QN(n12645) );
  NAND2X0 U12847 ( .IN1(g2703), .IN2(n8120), .QN(n12644) );
  NAND2X0 U12848 ( .IN1(n7756), .IN2(g7425), .QN(n12643) );
  XOR2X1 U12849 ( .IN1(n8073), .IN2(n8890), .Q(n12641) );
  INVX0 U12850 ( .INP(n8891), .ZN(n8890) );
  NAND3X0 U12851 ( .IN1(n12646), .IN2(n12647), .IN3(n12648), .QN(n8891) );
  NAND2X0 U12852 ( .IN1(n7759), .IN2(g7487), .QN(n12648) );
  NAND2X0 U12853 ( .IN1(n7829), .IN2(g2703), .QN(n12647) );
  NAND2X0 U12854 ( .IN1(n7760), .IN2(g7425), .QN(n12646) );
  XOR2X1 U12855 ( .IN1(n4415), .IN2(n8912), .Q(n12635) );
  NAND3X0 U12856 ( .IN1(n12649), .IN2(n12650), .IN3(n12651), .QN(n8912) );
  NAND2X0 U12857 ( .IN1(n7753), .IN2(g7487), .QN(n12651) );
  NAND2X0 U12858 ( .IN1(n7827), .IN2(g2703), .QN(n12650) );
  NAND2X0 U12859 ( .IN1(n7754), .IN2(g7425), .QN(n12649) );
  XOR2X1 U12860 ( .IN1(g2746), .IN2(n8895), .Q(n12634) );
  INVX0 U12861 ( .INP(n8896), .ZN(n8895) );
  NAND3X0 U12862 ( .IN1(n12652), .IN2(n12653), .IN3(n12654), .QN(n8896) );
  NAND2X0 U12863 ( .IN1(n7761), .IN2(g7487), .QN(n12654) );
  NAND2X0 U12864 ( .IN1(n7830), .IN2(g2703), .QN(n12653) );
  NAND2X0 U12865 ( .IN1(n7762), .IN2(g7425), .QN(n12652) );
  NAND2X0 U12866 ( .IN1(n7556), .IN2(g7487), .QN(n12607) );
  INVX0 U12867 ( .INP(n12655), .ZN(n9243) );
  NAND3X0 U12868 ( .IN1(n12656), .IN2(n12657), .IN3(n12658), .QN(n12655) );
  NAND2X0 U12869 ( .IN1(n7555), .IN2(g7487), .QN(n12658) );
  NAND2X0 U12870 ( .IN1(n7613), .IN2(g2703), .QN(n12657) );
  NAND2X0 U12871 ( .IN1(n7563), .IN2(g7425), .QN(n12656) );
  NAND2X0 U12872 ( .IN1(n12659), .IN2(n12660), .QN(g25271) );
  NAND2X0 U12873 ( .IN1(n9317), .IN2(g2116), .QN(n12660) );
  NAND2X0 U12874 ( .IN1(n12661), .IN2(n12600), .QN(n12659) );
  NAND2X0 U12875 ( .IN1(n12662), .IN2(n12663), .QN(g25270) );
  INVX0 U12876 ( .INP(n12664), .ZN(n12663) );
  NOR2X0 U12877 ( .IN1(n12665), .IN2(n7500), .QN(n12664) );
  NAND2X0 U12878 ( .IN1(n12666), .IN2(n12665), .QN(n12662) );
  NAND2X0 U12879 ( .IN1(n12667), .IN2(n12668), .QN(g25268) );
  NAND2X0 U12880 ( .IN1(n12669), .IN2(g2115), .QN(n12668) );
  NAND2X0 U12881 ( .IN1(n12670), .IN2(n12600), .QN(n12667) );
  INVX0 U12882 ( .INP(n12671), .ZN(n12600) );
  NAND4X0 U12883 ( .IN1(n9259), .IN2(n12672), .IN3(n12673), .IN4(n12674), .QN(
        n12671) );
  NAND2X0 U12884 ( .IN1(n8028), .IN2(g7229), .QN(n12674) );
  NOR2X0 U12885 ( .IN1(n12675), .IN2(n12676), .QN(n12673) );
  NOR2X0 U12886 ( .IN1(n4293), .IN2(g2108), .QN(n12676) );
  NOR4X0 U12887 ( .IN1(n12677), .IN2(n12678), .IN3(n12679), .IN4(n12680), .QN(
        n12675) );
  XNOR2X1 U12888 ( .IN1(n4420), .IN2(n9016), .Q(n12680) );
  NAND3X0 U12889 ( .IN1(n12681), .IN2(n12682), .IN3(n12683), .QN(n9016) );
  NAND2X0 U12890 ( .IN1(n7785), .IN2(g7357), .QN(n12683) );
  NAND2X0 U12891 ( .IN1(n7842), .IN2(g2009), .QN(n12682) );
  NAND2X0 U12892 ( .IN1(n7786), .IN2(g7229), .QN(n12681) );
  XNOR2X1 U12893 ( .IN1(n4399), .IN2(n8991), .Q(n12679) );
  NAND3X0 U12894 ( .IN1(n12684), .IN2(n12685), .IN3(n12686), .QN(n8991) );
  NAND2X0 U12895 ( .IN1(g7357), .IN2(n8121), .QN(n12686) );
  NAND2X0 U12896 ( .IN1(n7840), .IN2(g2009), .QN(n12685) );
  NAND2X0 U12897 ( .IN1(n7782), .IN2(g7229), .QN(n12684) );
  NAND3X0 U12898 ( .IN1(n12687), .IN2(n12688), .IN3(n12689), .QN(n12678) );
  XOR2X1 U12899 ( .IN1(n4468), .IN2(n9007), .Q(n12689) );
  NAND3X0 U12900 ( .IN1(n12690), .IN2(n12691), .IN3(n12692), .QN(n9007) );
  NAND2X0 U12901 ( .IN1(n7778), .IN2(g7357), .QN(n12692) );
  NAND2X0 U12902 ( .IN1(n7838), .IN2(g2009), .QN(n12691) );
  NAND2X0 U12903 ( .IN1(n7779), .IN2(g7229), .QN(n12690) );
  XOR2X1 U12904 ( .IN1(g2059), .IN2(n8979), .Q(n12688) );
  INVX0 U12905 ( .INP(n8982), .ZN(n8979) );
  NAND3X0 U12906 ( .IN1(n12693), .IN2(n12694), .IN3(n12695), .QN(n8982) );
  NAND2X0 U12907 ( .IN1(n7776), .IN2(g7357), .QN(n12695) );
  NAND2X0 U12908 ( .IN1(n7837), .IN2(g2009), .QN(n12694) );
  NAND2X0 U12909 ( .IN1(n7777), .IN2(g7229), .QN(n12693) );
  XOR2X1 U12910 ( .IN1(g2020), .IN2(n9001), .Q(n12687) );
  INVX0 U12911 ( .INP(n9003), .ZN(n9001) );
  NAND3X0 U12912 ( .IN1(n12696), .IN2(n12697), .IN3(n12698), .QN(n9003) );
  NAND2X0 U12913 ( .IN1(n7789), .IN2(g7357), .QN(n12698) );
  NAND2X0 U12914 ( .IN1(n7844), .IN2(g2009), .QN(n12697) );
  NAND2X0 U12915 ( .IN1(n7790), .IN2(g7229), .QN(n12696) );
  NAND4X0 U12916 ( .IN1(n12699), .IN2(n12700), .IN3(n12701), .IN4(n12702), 
        .QN(n12677) );
  XOR2X1 U12917 ( .IN1(g2013), .IN2(n8986), .Q(n12702) );
  INVX0 U12918 ( .INP(n8987), .ZN(n8986) );
  NAND3X0 U12919 ( .IN1(n12703), .IN2(n12704), .IN3(n12705), .QN(n8987) );
  NAND2X0 U12920 ( .IN1(n7787), .IN2(g7357), .QN(n12705) );
  NAND2X0 U12921 ( .IN1(n7843), .IN2(g2009), .QN(n12704) );
  NAND2X0 U12922 ( .IN1(n7788), .IN2(g7229), .QN(n12703) );
  NOR2X0 U12923 ( .IN1(n12706), .IN2(n12707), .QN(n12701) );
  XOR2X1 U12924 ( .IN1(n4409), .IN2(n9011), .Q(n12707) );
  INVX0 U12925 ( .INP(n9012), .ZN(n9011) );
  NAND3X0 U12926 ( .IN1(n12708), .IN2(n12709), .IN3(n12710), .QN(n9012) );
  NAND2X0 U12927 ( .IN1(n7780), .IN2(g7357), .QN(n12710) );
  NAND2X0 U12928 ( .IN1(n7839), .IN2(g2009), .QN(n12709) );
  NAND2X0 U12929 ( .IN1(n7781), .IN2(g7229), .QN(n12708) );
  XOR2X1 U12930 ( .IN1(n8085), .IN2(n9033), .Q(n12706) );
  INVX0 U12931 ( .INP(n9034), .ZN(n9033) );
  NAND3X0 U12932 ( .IN1(n12711), .IN2(n12712), .IN3(n12713), .QN(n9034) );
  NAND2X0 U12933 ( .IN1(n7774), .IN2(g7357), .QN(n12713) );
  NAND2X0 U12934 ( .IN1(n7836), .IN2(g2009), .QN(n12712) );
  NAND2X0 U12935 ( .IN1(n7775), .IN2(g7229), .QN(n12711) );
  XOR2X1 U12936 ( .IN1(n4416), .IN2(n9027), .Q(n12700) );
  NAND3X0 U12937 ( .IN1(n12714), .IN2(n12715), .IN3(n12716), .QN(n9027) );
  NAND2X0 U12938 ( .IN1(g7357), .IN2(n8122), .QN(n12716) );
  NAND2X0 U12939 ( .IN1(n7835), .IN2(g2009), .QN(n12715) );
  NAND2X0 U12940 ( .IN1(n7773), .IN2(g7229), .QN(n12714) );
  XOR2X1 U12941 ( .IN1(g2026), .IN2(n8996), .Q(n12699) );
  INVX0 U12942 ( .INP(n8997), .ZN(n8996) );
  NAND3X0 U12943 ( .IN1(n12717), .IN2(n12718), .IN3(n12719), .QN(n8997) );
  NAND2X0 U12944 ( .IN1(n7783), .IN2(g7357), .QN(n12719) );
  NAND2X0 U12945 ( .IN1(n7841), .IN2(g2009), .QN(n12718) );
  NAND2X0 U12946 ( .IN1(n7784), .IN2(g7229), .QN(n12717) );
  NAND2X0 U12947 ( .IN1(n7558), .IN2(g7357), .QN(n12672) );
  INVX0 U12948 ( .INP(n12720), .ZN(n9259) );
  NAND3X0 U12949 ( .IN1(n12721), .IN2(n12722), .IN3(n12723), .QN(n12720) );
  NAND2X0 U12950 ( .IN1(n7557), .IN2(g7357), .QN(n12723) );
  NAND2X0 U12951 ( .IN1(n7615), .IN2(g2009), .QN(n12722) );
  NAND2X0 U12952 ( .IN1(n7564), .IN2(g7229), .QN(n12721) );
  NAND2X0 U12953 ( .IN1(n12724), .IN2(n12725), .QN(g25267) );
  NAND2X0 U12954 ( .IN1(n8518), .IN2(g1422), .QN(n12725) );
  NAND2X0 U12955 ( .IN1(n12726), .IN2(n12666), .QN(n12724) );
  NAND2X0 U12956 ( .IN1(n12727), .IN2(n12728), .QN(g25266) );
  NAND2X0 U12957 ( .IN1(n12729), .IN2(g734), .QN(n12728) );
  NAND2X0 U12958 ( .IN1(n12730), .IN2(n12731), .QN(n12727) );
  NAND2X0 U12959 ( .IN1(n12732), .IN2(n12733), .QN(g25265) );
  NAND2X0 U12960 ( .IN1(n12153), .IN2(n8726), .QN(n12733) );
  NAND2X0 U12961 ( .IN1(n12734), .IN2(n9283), .QN(n12732) );
  XOR2X1 U12962 ( .IN1(n8032), .IN2(n8031), .Q(n12734) );
  NAND2X0 U12963 ( .IN1(n12735), .IN2(n12736), .QN(g25263) );
  NAND2X0 U12964 ( .IN1(n12737), .IN2(g1421), .QN(n12736) );
  NAND2X0 U12965 ( .IN1(n12738), .IN2(n12666), .QN(n12735) );
  INVX0 U12966 ( .INP(n12739), .ZN(n12666) );
  NAND4X0 U12967 ( .IN1(n9275), .IN2(n12740), .IN3(n12741), .IN4(n12742), .QN(
        n12739) );
  NAND2X0 U12968 ( .IN1(n8023), .IN2(g6979), .QN(n12742) );
  NOR2X0 U12969 ( .IN1(n12743), .IN2(n12744), .QN(n12741) );
  NOR2X0 U12970 ( .IN1(test_so51), .IN2(n4294), .QN(n12744) );
  NOR4X0 U12971 ( .IN1(n12745), .IN2(n12746), .IN3(n12747), .IN4(n12748), .QN(
        n12743) );
  XOR2X1 U12972 ( .IN1(n4412), .IN2(n9113), .Q(n12748) );
  INVX0 U12973 ( .INP(n9114), .ZN(n9113) );
  NAND3X0 U12974 ( .IN1(n12749), .IN2(n12750), .IN3(n12751), .QN(n9114) );
  NAND2X0 U12975 ( .IN1(n7802), .IN2(g7161), .QN(n12751) );
  NAND2X0 U12976 ( .IN1(n7851), .IN2(g1315), .QN(n12750) );
  NAND2X0 U12977 ( .IN1(n7803), .IN2(g6979), .QN(n12749) );
  XOR2X1 U12978 ( .IN1(n4417), .IN2(n9143), .Q(n12747) );
  INVX0 U12979 ( .INP(n9144), .ZN(n9143) );
  NAND3X0 U12980 ( .IN1(n12752), .IN2(n12753), .IN3(n12754), .QN(n9144) );
  NAND2X0 U12981 ( .IN1(n7791), .IN2(g7161), .QN(n12754) );
  NAND2X0 U12982 ( .IN1(n7845), .IN2(g1315), .QN(n12753) );
  NAND2X0 U12983 ( .IN1(n7792), .IN2(g6979), .QN(n12752) );
  NAND3X0 U12984 ( .IN1(n12755), .IN2(n12756), .IN3(n12757), .QN(n12746) );
  XOR2X1 U12985 ( .IN1(g1358), .IN2(n9128), .Q(n12757) );
  INVX0 U12986 ( .INP(n9129), .ZN(n9128) );
  NAND3X0 U12987 ( .IN1(n12758), .IN2(n12759), .IN3(n12760), .QN(n9129) );
  NAND2X0 U12988 ( .IN1(g7161), .IN2(n8123), .QN(n12760) );
  NAND2X0 U12989 ( .IN1(n7849), .IN2(g1315), .QN(n12759) );
  NAND2X0 U12990 ( .IN1(n7799), .IN2(g6979), .QN(n12758) );
  XOR2X1 U12991 ( .IN1(g1372), .IN2(n9150), .Q(n12756) );
  INVX0 U12992 ( .INP(n9151), .ZN(n9150) );
  NAND3X0 U12993 ( .IN1(n12761), .IN2(n12762), .IN3(n12763), .QN(n9151) );
  NAND2X0 U12994 ( .IN1(n7793), .IN2(g7161), .QN(n12763) );
  NAND2X0 U12995 ( .IN1(n7846), .IN2(g1315), .QN(n12762) );
  NAND2X0 U12996 ( .IN1(n7794), .IN2(g6979), .QN(n12761) );
  XOR2X1 U12997 ( .IN1(g1319), .IN2(n9103), .Q(n12755) );
  INVX0 U12998 ( .INP(n9104), .ZN(n9103) );
  NAND3X0 U12999 ( .IN1(n12764), .IN2(n12765), .IN3(n12766), .QN(n9104) );
  NAND2X0 U13000 ( .IN1(n7806), .IN2(g7161), .QN(n12766) );
  NAND2X0 U13001 ( .IN1(n7853), .IN2(g1315), .QN(n12765) );
  NAND2X0 U13002 ( .IN1(n7807), .IN2(g6979), .QN(n12764) );
  NAND4X0 U13003 ( .IN1(n12767), .IN2(n12768), .IN3(n12769), .IN4(n12770), 
        .QN(n12745) );
  XOR2X1 U13004 ( .IN1(n4469), .IN2(n9124), .Q(n12770) );
  NAND3X0 U13005 ( .IN1(n12771), .IN2(n12772), .IN3(n12773), .QN(n9124) );
  NAND2X0 U13006 ( .IN1(n7797), .IN2(g7161), .QN(n12773) );
  NAND2X0 U13007 ( .IN1(n7848), .IN2(g1315), .QN(n12772) );
  NAND2X0 U13008 ( .IN1(n7798), .IN2(g6979), .QN(n12771) );
  NOR2X0 U13009 ( .IN1(n12774), .IN2(n12775), .QN(n12769) );
  XNOR2X1 U13010 ( .IN1(n4402), .IN2(n9119), .Q(n12775) );
  NAND3X0 U13011 ( .IN1(n12776), .IN2(n12777), .IN3(n12778), .QN(n9119) );
  NAND2X0 U13012 ( .IN1(n7808), .IN2(g7161), .QN(n12778) );
  NAND2X0 U13013 ( .IN1(n7854), .IN2(g1315), .QN(n12777) );
  NAND2X0 U13014 ( .IN1(g6979), .IN2(n8124), .QN(n12776) );
  XOR2X1 U13015 ( .IN1(n4475), .IN2(n9096), .Q(n12774) );
  INVX0 U13016 ( .INP(n9099), .ZN(n9096) );
  NAND3X0 U13017 ( .IN1(n12779), .IN2(n12780), .IN3(n12781), .QN(n9099) );
  NAND2X0 U13018 ( .IN1(n7795), .IN2(g7161), .QN(n12781) );
  NAND2X0 U13019 ( .IN1(n7847), .IN2(g1315), .QN(n12780) );
  NAND2X0 U13020 ( .IN1(n7796), .IN2(g6979), .QN(n12779) );
  XOR2X1 U13021 ( .IN1(g1346), .IN2(n9107), .Q(n12768) );
  INVX0 U13022 ( .INP(n9110), .ZN(n9107) );
  NAND3X0 U13023 ( .IN1(n12782), .IN2(n12783), .IN3(n12784), .QN(n9110) );
  NAND2X0 U13024 ( .IN1(n7800), .IN2(g7161), .QN(n12784) );
  NAND2X0 U13025 ( .IN1(n7850), .IN2(g1315), .QN(n12783) );
  NAND2X0 U13026 ( .IN1(n7801), .IN2(g6979), .QN(n12782) );
  XOR2X1 U13027 ( .IN1(n4421), .IN2(n9133), .Q(n12767) );
  NAND3X0 U13028 ( .IN1(n12785), .IN2(n12786), .IN3(n12787), .QN(n9133) );
  NAND2X0 U13029 ( .IN1(n7804), .IN2(g7161), .QN(n12787) );
  NAND2X0 U13030 ( .IN1(n7852), .IN2(g1315), .QN(n12786) );
  NAND2X0 U13031 ( .IN1(n7805), .IN2(g6979), .QN(n12785) );
  NAND2X0 U13032 ( .IN1(n7560), .IN2(g7161), .QN(n12740) );
  INVX0 U13033 ( .INP(n12788), .ZN(n9275) );
  NAND3X0 U13034 ( .IN1(n12789), .IN2(n12790), .IN3(n12791), .QN(n12788) );
  NAND2X0 U13035 ( .IN1(n7559), .IN2(g7161), .QN(n12791) );
  NAND2X0 U13036 ( .IN1(n7617), .IN2(g1315), .QN(n12790) );
  NAND2X0 U13037 ( .IN1(n7565), .IN2(g6979), .QN(n12789) );
  NAND2X0 U13038 ( .IN1(n12792), .IN2(n12793), .QN(g25262) );
  NAND2X0 U13039 ( .IN1(n8539), .IN2(g736), .QN(n12793) );
  NAND2X0 U13040 ( .IN1(n12794), .IN2(n12730), .QN(n12792) );
  NAND2X0 U13041 ( .IN1(n12795), .IN2(n12796), .QN(g25260) );
  NAND2X0 U13042 ( .IN1(n12797), .IN2(g735), .QN(n12796) );
  NAND2X0 U13043 ( .IN1(n12798), .IN2(n12730), .QN(n12795) );
  INVX0 U13044 ( .INP(n12799), .ZN(n12730) );
  NAND4X0 U13045 ( .IN1(n9230), .IN2(n12800), .IN3(n12801), .IN4(n12802), .QN(
        n12799) );
  NAND2X0 U13046 ( .IN1(n8022), .IN2(g6677), .QN(n12802) );
  NOR2X0 U13047 ( .IN1(n12803), .IN2(n12804), .QN(n12801) );
  NOR2X0 U13048 ( .IN1(n4295), .IN2(g728), .QN(n12804) );
  NOR4X0 U13049 ( .IN1(n12805), .IN2(n12806), .IN3(n12807), .IN4(n12808), .QN(
        n12803) );
  XOR2X1 U13050 ( .IN1(n4422), .IN2(n8772), .Q(n12808) );
  INVX0 U13051 ( .INP(n8773), .ZN(n8772) );
  NAND3X0 U13052 ( .IN1(n12809), .IN2(n12810), .IN3(n12811), .QN(n8773) );
  NAND2X0 U13053 ( .IN1(n7821), .IN2(g6911), .QN(n12811) );
  NAND2X0 U13054 ( .IN1(n7862), .IN2(g629), .QN(n12810) );
  NAND2X0 U13055 ( .IN1(n7822), .IN2(g6677), .QN(n12809) );
  XOR2X1 U13056 ( .IN1(n4477), .IN2(n8781), .Q(n12807) );
  INVX0 U13057 ( .INP(n8782), .ZN(n8781) );
  NAND3X0 U13058 ( .IN1(n12812), .IN2(n12813), .IN3(n12814), .QN(n8782) );
  NAND2X0 U13059 ( .IN1(n7812), .IN2(g6911), .QN(n12814) );
  NAND2X0 U13060 ( .IN1(n7857), .IN2(g629), .QN(n12813) );
  NAND2X0 U13061 ( .IN1(n7813), .IN2(g6677), .QN(n12812) );
  NAND3X0 U13062 ( .IN1(n12815), .IN2(n12816), .IN3(n12817), .QN(n12806) );
  XOR2X1 U13063 ( .IN1(g660), .IN2(n8757), .Q(n12817) );
  INVX0 U13064 ( .INP(n8758), .ZN(n8757) );
  NAND3X0 U13065 ( .IN1(n12818), .IN2(n12819), .IN3(n12820), .QN(n8758) );
  NAND2X0 U13066 ( .IN1(n7818), .IN2(g6911), .QN(n12820) );
  NAND2X0 U13067 ( .IN1(n7860), .IN2(g629), .QN(n12819) );
  NAND2X0 U13068 ( .IN1(g6677), .IN2(n8125), .QN(n12818) );
  XOR2X1 U13069 ( .IN1(g640), .IN2(n8777), .Q(n12816) );
  INVX0 U13070 ( .INP(n8778), .ZN(n8777) );
  NAND3X0 U13071 ( .IN1(n12821), .IN2(n12822), .IN3(n12823), .QN(n8778) );
  NAND2X0 U13072 ( .IN1(n7825), .IN2(g6911), .QN(n12823) );
  NAND2X0 U13073 ( .IN1(n7864), .IN2(g629), .QN(n12822) );
  NAND2X0 U13074 ( .IN1(n7826), .IN2(g6677), .QN(n12821) );
  XOR2X1 U13075 ( .IN1(g646), .IN2(n8762), .Q(n12815) );
  INVX0 U13076 ( .INP(n8763), .ZN(n8762) );
  NAND3X0 U13077 ( .IN1(n12824), .IN2(n12825), .IN3(n12826), .QN(n8763) );
  NAND2X0 U13078 ( .IN1(n7819), .IN2(g6911), .QN(n12826) );
  NAND2X0 U13079 ( .IN1(n7861), .IN2(g629), .QN(n12825) );
  NAND2X0 U13080 ( .IN1(n7820), .IN2(g6677), .QN(n12824) );
  NAND4X0 U13081 ( .IN1(n12827), .IN2(n12828), .IN3(n12829), .IN4(n12830), 
        .QN(n12805) );
  XOR2X1 U13082 ( .IN1(g633), .IN2(n8767), .Q(n12830) );
  INVX0 U13083 ( .INP(n8768), .ZN(n8767) );
  NAND3X0 U13084 ( .IN1(n12831), .IN2(n12832), .IN3(n12833), .QN(n8768) );
  NAND2X0 U13085 ( .IN1(n7823), .IN2(g6911), .QN(n12833) );
  NAND2X0 U13086 ( .IN1(n7863), .IN2(g629), .QN(n12832) );
  NAND2X0 U13087 ( .IN1(n7824), .IN2(g6677), .QN(n12831) );
  NOR2X0 U13088 ( .IN1(n12834), .IN2(n12835), .QN(n12829) );
  XOR2X1 U13089 ( .IN1(n4396), .IN2(n8792), .Q(n12835) );
  INVX0 U13090 ( .INP(n8793), .ZN(n8792) );
  NAND3X0 U13091 ( .IN1(n12836), .IN2(n12837), .IN3(n12838), .QN(n8793) );
  NAND2X0 U13092 ( .IN1(n7810), .IN2(g6911), .QN(n12838) );
  NAND2X0 U13093 ( .IN1(n7856), .IN2(g629), .QN(n12837) );
  NAND2X0 U13094 ( .IN1(n7811), .IN2(g6677), .QN(n12836) );
  XOR2X1 U13095 ( .IN1(n8074), .IN2(n8750), .Q(n12834) );
  INVX0 U13096 ( .INP(n8753), .ZN(n8750) );
  NAND3X0 U13097 ( .IN1(n12839), .IN2(n12840), .IN3(n12841), .QN(n8753) );
  NAND2X0 U13098 ( .IN1(n7814), .IN2(g6911), .QN(n12841) );
  NAND2X0 U13099 ( .IN1(n7858), .IN2(g629), .QN(n12840) );
  NAND2X0 U13100 ( .IN1(n7815), .IN2(g6677), .QN(n12839) );
  XOR2X1 U13101 ( .IN1(n4418), .IN2(n8802), .Q(n12828) );
  NAND3X0 U13102 ( .IN1(n12842), .IN2(n12843), .IN3(n12844), .QN(n8802) );
  NAND2X0 U13103 ( .IN1(g6911), .IN2(n8126), .QN(n12844) );
  NAND2X0 U13104 ( .IN1(n7855), .IN2(g629), .QN(n12843) );
  NAND2X0 U13105 ( .IN1(n7809), .IN2(g6677), .QN(n12842) );
  XOR2X1 U13106 ( .IN1(g672), .IN2(n8744), .Q(n12827) );
  INVX0 U13107 ( .INP(n8747), .ZN(n8744) );
  NAND3X0 U13108 ( .IN1(n12845), .IN2(n12846), .IN3(n12847), .QN(n8747) );
  NAND2X0 U13109 ( .IN1(n7816), .IN2(g6911), .QN(n12847) );
  NAND2X0 U13110 ( .IN1(n7859), .IN2(g629), .QN(n12846) );
  NAND2X0 U13111 ( .IN1(n7817), .IN2(g6677), .QN(n12845) );
  NAND2X0 U13112 ( .IN1(n7562), .IN2(g6911), .QN(n12800) );
  INVX0 U13113 ( .INP(n12848), .ZN(n9230) );
  NAND3X0 U13114 ( .IN1(n12849), .IN2(n12850), .IN3(n12851), .QN(n12848) );
  NAND2X0 U13115 ( .IN1(n7561), .IN2(g6911), .QN(n12851) );
  NAND2X0 U13116 ( .IN1(n7618), .IN2(g629), .QN(n12850) );
  NAND2X0 U13117 ( .IN1(n7566), .IN2(g6677), .QN(n12849) );
  NAND2X0 U13118 ( .IN1(n12852), .IN2(n12853), .QN(g25259) );
  INVX0 U13119 ( .INP(n12854), .ZN(n12853) );
  NOR2X0 U13120 ( .IN1(n12855), .IN2(n7567), .QN(n12854) );
  NAND2X0 U13121 ( .IN1(n12855), .IN2(n12057), .QN(n12852) );
  NAND2X0 U13122 ( .IN1(n12856), .IN2(n12857), .QN(g25257) );
  INVX0 U13123 ( .INP(n12858), .ZN(n12857) );
  NOR2X0 U13124 ( .IN1(n12859), .IN2(n7568), .QN(n12858) );
  NAND2X0 U13125 ( .IN1(n12859), .IN2(n12057), .QN(n12856) );
  NAND2X0 U13126 ( .IN1(n12860), .IN2(n12861), .QN(g25256) );
  NAND2X0 U13127 ( .IN1(n12855), .IN2(n4377), .QN(n12861) );
  INVX0 U13128 ( .INP(n12862), .ZN(n12860) );
  NOR2X0 U13129 ( .IN1(n12855), .IN2(n7570), .QN(n12862) );
  NAND2X0 U13130 ( .IN1(n12863), .IN2(n12864), .QN(g25255) );
  NAND2X0 U13131 ( .IN1(n4033), .IN2(g1559), .QN(n12864) );
  NAND2X0 U13132 ( .IN1(n12090), .IN2(n12865), .QN(n12863) );
  NAND2X0 U13133 ( .IN1(n12866), .IN2(n12867), .QN(g25253) );
  NAND2X0 U13134 ( .IN1(n4034), .IN2(g2254), .QN(n12867) );
  NAND2X0 U13135 ( .IN1(n12057), .IN2(n12868), .QN(n12866) );
  NAND4X0 U13136 ( .IN1(g2200), .IN2(g2175), .IN3(n12869), .IN4(n12870), .QN(
        n12057) );
  NOR4X0 U13137 ( .IN1(n4563), .IN2(n4555), .IN3(n4389), .IN4(n4377), .QN(
        n12870) );
  NOR2X0 U13138 ( .IN1(n4373), .IN2(n4325), .QN(n12869) );
  NAND2X0 U13139 ( .IN1(n12871), .IN2(n12872), .QN(g25252) );
  NAND2X0 U13140 ( .IN1(n12859), .IN2(n4377), .QN(n12872) );
  INVX0 U13141 ( .INP(n12873), .ZN(n12871) );
  NOR2X0 U13142 ( .IN1(n12859), .IN2(n7571), .QN(n12873) );
  NAND2X0 U13143 ( .IN1(n12874), .IN2(n12875), .QN(g25251) );
  NAND2X0 U13144 ( .IN1(n12855), .IN2(n4373), .QN(n12875) );
  INVX0 U13145 ( .INP(n12876), .ZN(n12874) );
  NOR2X0 U13146 ( .IN1(n12855), .IN2(n7573), .QN(n12876) );
  NAND2X0 U13147 ( .IN1(n12877), .IN2(n12878), .QN(g25250) );
  NAND2X0 U13148 ( .IN1(n4037), .IN2(g1561), .QN(n12878) );
  NAND2X0 U13149 ( .IN1(n12090), .IN2(n12879), .QN(n12877) );
  NAND2X0 U13150 ( .IN1(n12880), .IN2(n12881), .QN(g25249) );
  NAND2X0 U13151 ( .IN1(n4378), .IN2(n12865), .QN(n12881) );
  NAND2X0 U13152 ( .IN1(n4033), .IN2(g1556), .QN(n12880) );
  NAND2X0 U13153 ( .IN1(n12882), .IN2(n12883), .QN(g25248) );
  NAND2X0 U13154 ( .IN1(n4038), .IN2(g865), .QN(n12883) );
  NAND2X0 U13155 ( .IN1(n12120), .IN2(n12884), .QN(n12882) );
  NAND2X0 U13156 ( .IN1(n12885), .IN2(n12886), .QN(g25247) );
  NAND2X0 U13157 ( .IN1(n4377), .IN2(n12868), .QN(n12886) );
  NAND2X0 U13158 ( .IN1(n4034), .IN2(g2251), .QN(n12885) );
  NAND2X0 U13159 ( .IN1(n12887), .IN2(n12888), .QN(g25246) );
  NAND2X0 U13160 ( .IN1(n12859), .IN2(n4373), .QN(n12888) );
  INVX0 U13161 ( .INP(n12889), .ZN(n12887) );
  NOR2X0 U13162 ( .IN1(n12859), .IN2(n7574), .QN(n12889) );
  NAND2X0 U13163 ( .IN1(n12890), .IN2(n12891), .QN(g25245) );
  NAND2X0 U13164 ( .IN1(n12892), .IN2(n12855), .QN(n12891) );
  INVX0 U13165 ( .INP(n12893), .ZN(n12890) );
  NOR2X0 U13166 ( .IN1(n12855), .IN2(n7576), .QN(n12893) );
  NOR2X0 U13167 ( .IN1(n12894), .IN2(n4367), .QN(n12855) );
  NAND2X0 U13168 ( .IN1(n12895), .IN2(n12896), .QN(g25244) );
  INVX0 U13169 ( .INP(n12897), .ZN(n12896) );
  NOR2X0 U13170 ( .IN1(n12898), .IN2(n7581), .QN(n12897) );
  NAND2X0 U13171 ( .IN1(n12898), .IN2(n12090), .QN(n12895) );
  NAND4X0 U13172 ( .IN1(g1506), .IN2(g1481), .IN3(n12899), .IN4(n12900), .QN(
        n12090) );
  NOR4X0 U13173 ( .IN1(n4565), .IN2(n4557), .IN3(n4390), .IN4(n4378), .QN(
        n12900) );
  NOR2X0 U13174 ( .IN1(n4374), .IN2(n4326), .QN(n12899) );
  NAND2X0 U13175 ( .IN1(n12901), .IN2(n12902), .QN(g25243) );
  NAND2X0 U13176 ( .IN1(n4378), .IN2(n12879), .QN(n12902) );
  NAND2X0 U13177 ( .IN1(n4037), .IN2(g1558), .QN(n12901) );
  NAND2X0 U13178 ( .IN1(n12903), .IN2(n12904), .QN(g25242) );
  NAND2X0 U13179 ( .IN1(test_so54), .IN2(n4033), .QN(n12904) );
  NAND2X0 U13180 ( .IN1(n4374), .IN2(n12865), .QN(n12903) );
  NAND2X0 U13181 ( .IN1(n12905), .IN2(n12906), .QN(g25241) );
  NAND2X0 U13182 ( .IN1(n4043), .IN2(g867), .QN(n12906) );
  NAND2X0 U13183 ( .IN1(n12120), .IN2(n12907), .QN(n12905) );
  NAND2X0 U13184 ( .IN1(n12908), .IN2(n12909), .QN(g25240) );
  NAND2X0 U13185 ( .IN1(n4379), .IN2(n12884), .QN(n12909) );
  NAND2X0 U13186 ( .IN1(n4038), .IN2(g862), .QN(n12908) );
  NAND2X0 U13187 ( .IN1(n12910), .IN2(n12911), .QN(g25239) );
  INVX0 U13188 ( .INP(n12912), .ZN(n12911) );
  NOR2X0 U13189 ( .IN1(n12913), .IN2(n7601), .QN(n12912) );
  NAND2X0 U13190 ( .IN1(n12913), .IN2(n12145), .QN(n12910) );
  NAND2X0 U13191 ( .IN1(n12914), .IN2(n12915), .QN(g25237) );
  NAND2X0 U13192 ( .IN1(n4373), .IN2(n12868), .QN(n12915) );
  NAND2X0 U13193 ( .IN1(n4034), .IN2(g2248), .QN(n12914) );
  NAND2X0 U13194 ( .IN1(n12916), .IN2(n12917), .QN(g25236) );
  NAND2X0 U13195 ( .IN1(n12892), .IN2(n12859), .QN(n12917) );
  INVX0 U13196 ( .INP(n12918), .ZN(n12916) );
  NOR2X0 U13197 ( .IN1(n12859), .IN2(n7577), .QN(n12918) );
  NOR2X0 U13198 ( .IN1(n12894), .IN2(n8070), .QN(n12859) );
  NAND2X0 U13199 ( .IN1(n12919), .IN2(n12920), .QN(g25235) );
  NAND2X0 U13200 ( .IN1(n12898), .IN2(n4378), .QN(n12920) );
  INVX0 U13201 ( .INP(n12921), .ZN(n12919) );
  NOR2X0 U13202 ( .IN1(n12898), .IN2(n7584), .QN(n12921) );
  NAND2X0 U13203 ( .IN1(n12922), .IN2(n12923), .QN(g25234) );
  NAND2X0 U13204 ( .IN1(n4374), .IN2(n12879), .QN(n12923) );
  NAND2X0 U13205 ( .IN1(n4037), .IN2(g1555), .QN(n12922) );
  NAND2X0 U13206 ( .IN1(n12924), .IN2(n12925), .QN(g25233) );
  NAND2X0 U13207 ( .IN1(n12926), .IN2(n12865), .QN(n12925) );
  INVX0 U13208 ( .INP(n4033), .ZN(n12865) );
  NAND2X0 U13209 ( .IN1(n4033), .IN2(g1550), .QN(n12924) );
  NAND2X0 U13210 ( .IN1(n19), .IN2(g1547), .QN(n4033) );
  NAND2X0 U13211 ( .IN1(n12927), .IN2(n12928), .QN(g25232) );
  NAND2X0 U13212 ( .IN1(n4046), .IN2(g866), .QN(n12928) );
  NAND2X0 U13213 ( .IN1(n12120), .IN2(n12929), .QN(n12927) );
  NAND4X0 U13214 ( .IN1(g813), .IN2(g793), .IN3(n12930), .IN4(n12931), .QN(
        n12120) );
  NOR4X0 U13215 ( .IN1(n4567), .IN2(n4559), .IN3(n4391), .IN4(n4379), .QN(
        n12931) );
  NOR2X0 U13216 ( .IN1(n4375), .IN2(n4327), .QN(n12930) );
  NAND2X0 U13217 ( .IN1(n12932), .IN2(n12933), .QN(g25231) );
  NAND2X0 U13218 ( .IN1(n4379), .IN2(n12907), .QN(n12933) );
  NAND2X0 U13219 ( .IN1(n4043), .IN2(g864), .QN(n12932) );
  NAND2X0 U13220 ( .IN1(n12934), .IN2(n12935), .QN(g25230) );
  NAND2X0 U13221 ( .IN1(n4375), .IN2(n12884), .QN(n12935) );
  NAND2X0 U13222 ( .IN1(n4038), .IN2(g859), .QN(n12934) );
  NAND2X0 U13223 ( .IN1(n12936), .IN2(n12937), .QN(g25229) );
  INVX0 U13224 ( .INP(n12938), .ZN(n12937) );
  NOR2X0 U13225 ( .IN1(n12939), .IN2(n7602), .QN(n12938) );
  NAND2X0 U13226 ( .IN1(n12939), .IN2(n12145), .QN(n12936) );
  NAND2X0 U13227 ( .IN1(n12940), .IN2(n12941), .QN(g25228) );
  NAND2X0 U13228 ( .IN1(n4380), .IN2(n12913), .QN(n12941) );
  INVX0 U13229 ( .INP(n12942), .ZN(n12940) );
  NOR2X0 U13230 ( .IN1(n12913), .IN2(n7604), .QN(n12942) );
  NAND2X0 U13231 ( .IN1(n12943), .IN2(n12944), .QN(g25227) );
  NAND2X0 U13232 ( .IN1(n12892), .IN2(n12868), .QN(n12944) );
  INVX0 U13233 ( .INP(n4034), .ZN(n12868) );
  NOR4X0 U13234 ( .IN1(g2195), .IN2(g2190), .IN3(n4287), .IN4(n4325), .QN(
        n12892) );
  NAND2X0 U13235 ( .IN1(n4034), .IN2(g2245), .QN(n12943) );
  NAND2X0 U13236 ( .IN1(n19), .IN2(g6837), .QN(n4034) );
  NAND2X0 U13237 ( .IN1(n12945), .IN2(n12946), .QN(g25225) );
  NAND2X0 U13238 ( .IN1(n12898), .IN2(n4374), .QN(n12946) );
  INVX0 U13239 ( .INP(n12947), .ZN(n12945) );
  NOR2X0 U13240 ( .IN1(n12898), .IN2(n7586), .QN(n12947) );
  NAND2X0 U13241 ( .IN1(n12948), .IN2(n12949), .QN(g25224) );
  NAND2X0 U13242 ( .IN1(n12926), .IN2(n12879), .QN(n12949) );
  INVX0 U13243 ( .INP(n4037), .ZN(n12879) );
  NAND2X0 U13244 ( .IN1(n4037), .IN2(g1552), .QN(n12948) );
  NAND2X0 U13245 ( .IN1(n19), .IN2(g6782), .QN(n4037) );
  NAND2X0 U13246 ( .IN1(n12950), .IN2(n12951), .QN(g25223) );
  NAND2X0 U13247 ( .IN1(n4379), .IN2(n12929), .QN(n12951) );
  NAND2X0 U13248 ( .IN1(n4046), .IN2(g863), .QN(n12950) );
  NAND2X0 U13249 ( .IN1(n12952), .IN2(n12953), .QN(g25222) );
  NAND2X0 U13250 ( .IN1(n4375), .IN2(n12907), .QN(n12953) );
  NAND2X0 U13251 ( .IN1(n4043), .IN2(g861), .QN(n12952) );
  NAND2X0 U13252 ( .IN1(n12954), .IN2(n12955), .QN(g25221) );
  NAND2X0 U13253 ( .IN1(n12956), .IN2(n12884), .QN(n12955) );
  INVX0 U13254 ( .INP(n4038), .ZN(n12884) );
  NAND2X0 U13255 ( .IN1(n4038), .IN2(g856), .QN(n12954) );
  NAND2X0 U13256 ( .IN1(n19), .IN2(test_so31), .QN(n4038) );
  NAND2X0 U13257 ( .IN1(n12957), .IN2(n12958), .QN(g25220) );
  INVX0 U13258 ( .INP(n12959), .ZN(n12958) );
  NOR2X0 U13259 ( .IN1(n12960), .IN2(n7603), .QN(n12959) );
  NAND2X0 U13260 ( .IN1(n12960), .IN2(n12145), .QN(n12957) );
  NAND4X0 U13261 ( .IN1(g125), .IN2(g105), .IN3(n12961), .IN4(n12962), .QN(
        n12145) );
  NOR4X0 U13262 ( .IN1(n4569), .IN2(n4561), .IN3(n4392), .IN4(n4380), .QN(
        n12962) );
  NOR2X0 U13263 ( .IN1(n4376), .IN2(n4328), .QN(n12961) );
  NAND2X0 U13264 ( .IN1(n12963), .IN2(n12964), .QN(g25219) );
  NAND2X0 U13265 ( .IN1(n4380), .IN2(n12939), .QN(n12964) );
  INVX0 U13266 ( .INP(n12965), .ZN(n12963) );
  NOR2X0 U13267 ( .IN1(n12939), .IN2(n7605), .QN(n12965) );
  NAND2X0 U13268 ( .IN1(n12966), .IN2(n12967), .QN(g25218) );
  NAND2X0 U13269 ( .IN1(n12913), .IN2(n4376), .QN(n12967) );
  INVX0 U13270 ( .INP(n12968), .ZN(n12966) );
  NOR2X0 U13271 ( .IN1(n12913), .IN2(n7607), .QN(n12968) );
  NAND2X0 U13272 ( .IN1(n12969), .IN2(n12970), .QN(g25217) );
  INVX0 U13273 ( .INP(n12971), .ZN(n12970) );
  NOR2X0 U13274 ( .IN1(n12898), .IN2(n7589), .QN(n12971) );
  NAND2X0 U13275 ( .IN1(n12926), .IN2(n12898), .QN(n12969) );
  NOR2X0 U13276 ( .IN1(n12894), .IN2(n4317), .QN(n12898) );
  NOR4X0 U13277 ( .IN1(g1501), .IN2(g1496), .IN3(n4288), .IN4(n4326), .QN(
        n12926) );
  NAND2X0 U13278 ( .IN1(n12972), .IN2(n12973), .QN(g25215) );
  NAND2X0 U13279 ( .IN1(n4375), .IN2(n12929), .QN(n12973) );
  NAND2X0 U13280 ( .IN1(n4046), .IN2(g860), .QN(n12972) );
  NAND2X0 U13281 ( .IN1(n12974), .IN2(n12975), .QN(g25214) );
  NAND2X0 U13282 ( .IN1(test_so33), .IN2(n4043), .QN(n12975) );
  NAND2X0 U13283 ( .IN1(n12956), .IN2(n12907), .QN(n12974) );
  INVX0 U13284 ( .INP(n4043), .ZN(n12907) );
  NAND2X0 U13285 ( .IN1(n19), .IN2(g6518), .QN(n4043) );
  NAND2X0 U13286 ( .IN1(n12976), .IN2(n12977), .QN(g25213) );
  NAND2X0 U13287 ( .IN1(n12960), .IN2(n4380), .QN(n12977) );
  INVX0 U13288 ( .INP(n12978), .ZN(n12976) );
  NOR2X0 U13289 ( .IN1(n12960), .IN2(n7606), .QN(n12978) );
  NAND2X0 U13290 ( .IN1(n12979), .IN2(n12980), .QN(g25212) );
  NAND2X0 U13291 ( .IN1(n12939), .IN2(n4376), .QN(n12980) );
  INVX0 U13292 ( .INP(n12981), .ZN(n12979) );
  NOR2X0 U13293 ( .IN1(n12939), .IN2(n7608), .QN(n12981) );
  NAND2X0 U13294 ( .IN1(n12982), .IN2(n12983), .QN(g25211) );
  NAND2X0 U13295 ( .IN1(n12984), .IN2(n12913), .QN(n12983) );
  INVX0 U13296 ( .INP(n12985), .ZN(n12982) );
  NOR2X0 U13297 ( .IN1(n12913), .IN2(n7610), .QN(n12985) );
  NOR2X0 U13298 ( .IN1(n12894), .IN2(n4369), .QN(n12913) );
  NAND2X0 U13299 ( .IN1(n12986), .IN2(n12987), .QN(g25209) );
  NAND2X0 U13300 ( .IN1(n12956), .IN2(n12929), .QN(n12987) );
  INVX0 U13301 ( .INP(n4046), .ZN(n12929) );
  NOR4X0 U13302 ( .IN1(g809), .IN2(g805), .IN3(n4289), .IN4(n4327), .QN(n12956) );
  NAND2X0 U13303 ( .IN1(n4046), .IN2(g857), .QN(n12986) );
  NAND2X0 U13304 ( .IN1(n19), .IN2(g6368), .QN(n4046) );
  INVX0 U13305 ( .INP(n12894), .ZN(n19) );
  NAND2X0 U13306 ( .IN1(n12988), .IN2(n12989), .QN(g25207) );
  NAND2X0 U13307 ( .IN1(n12960), .IN2(n4376), .QN(n12989) );
  INVX0 U13308 ( .INP(n12990), .ZN(n12988) );
  NOR2X0 U13309 ( .IN1(n12960), .IN2(n7609), .QN(n12990) );
  NAND2X0 U13310 ( .IN1(n12991), .IN2(n12992), .QN(g25206) );
  NAND2X0 U13311 ( .IN1(n12984), .IN2(n12939), .QN(n12992) );
  INVX0 U13312 ( .INP(n12993), .ZN(n12991) );
  NOR2X0 U13313 ( .IN1(n12939), .IN2(n7611), .QN(n12993) );
  NOR2X0 U13314 ( .IN1(n12894), .IN2(n4512), .QN(n12939) );
  NAND2X0 U13315 ( .IN1(n12994), .IN2(n12995), .QN(g25204) );
  INVX0 U13316 ( .INP(n12996), .ZN(n12995) );
  NOR2X0 U13317 ( .IN1(n12960), .IN2(n7612), .QN(n12996) );
  NAND2X0 U13318 ( .IN1(n12984), .IN2(n12960), .QN(n12994) );
  NOR2X0 U13319 ( .IN1(n12894), .IN2(n4318), .QN(n12960) );
  NAND4X0 U13320 ( .IN1(n7703), .IN2(n11799), .IN3(n8016), .IN4(n12997), .QN(
        n12894) );
  NOR4X0 U13321 ( .IN1(n4349), .IN2(n4330), .IN3(g2912), .IN4(g2917), .QN(
        n12997) );
  NOR4X0 U13322 ( .IN1(g121), .IN2(g117), .IN3(n4290), .IN4(n4328), .QN(n12984) );
  NOR2X0 U13323 ( .IN1(n12998), .IN2(n12999), .QN(g25202) );
  XOR2X1 U13324 ( .IN1(n7429), .IN2(n13000), .Q(n12999) );
  NOR3X0 U13325 ( .IN1(n8672), .IN2(n4057), .IN3(n12148), .QN(g25201) );
  NOR2X0 U13326 ( .IN1(n4058), .IN2(n4305), .QN(n12148) );
  NAND2X0 U13327 ( .IN1(n13001), .IN2(g2892), .QN(n4058) );
  NOR2X0 U13328 ( .IN1(n13002), .IN2(n13003), .QN(g25199) );
  XOR2X1 U13329 ( .IN1(n7703), .IN2(n13004), .Q(n13003) );
  NOR2X0 U13330 ( .IN1(n11303), .IN2(n13005), .QN(g25197) );
  XOR2X1 U13331 ( .IN1(n4397), .IN2(n9292), .Q(n13005) );
  NOR2X0 U13332 ( .IN1(n9305), .IN2(n13006), .QN(g25194) );
  XOR2X1 U13333 ( .IN1(n4399), .IN2(n12151), .Q(n13006) );
  NOR2X0 U13334 ( .IN1(n12153), .IN2(n13007), .QN(g25191) );
  XOR2X1 U13335 ( .IN1(n8051), .IN2(n4065), .Q(n13007) );
  NOR2X0 U13336 ( .IN1(n8512), .IN2(n13008), .QN(g25189) );
  XOR2X1 U13337 ( .IN1(n4401), .IN2(n8510), .Q(n13008) );
  NOR2X0 U13338 ( .IN1(n8536), .IN2(n13009), .QN(g25185) );
  XOR2X1 U13339 ( .IN1(n4403), .IN2(n8530), .Q(n13009) );
  NOR2X0 U13340 ( .IN1(n10265), .IN2(n13010), .QN(g25067) );
  XNOR2X1 U13341 ( .IN1(n7690), .IN2(n3888), .Q(n13010) );
  NAND2X0 U13342 ( .IN1(g2241), .IN2(n8578), .QN(n3888) );
  INVX0 U13343 ( .INP(n13011), .ZN(n10265) );
  NAND2X0 U13344 ( .IN1(n13012), .IN2(n11799), .QN(n13011) );
  NOR2X0 U13345 ( .IN1(n10267), .IN2(n13013), .QN(g25056) );
  XNOR2X1 U13346 ( .IN1(n7694), .IN2(n3891), .Q(n13013) );
  NAND2X0 U13347 ( .IN1(g1547), .IN2(n8578), .QN(n3891) );
  INVX0 U13348 ( .INP(n13014), .ZN(n10267) );
  NAND2X0 U13349 ( .IN1(n13015), .IN2(n11799), .QN(n13014) );
  NOR2X0 U13350 ( .IN1(n10269), .IN2(n13016), .QN(g25042) );
  XNOR2X1 U13351 ( .IN1(n7698), .IN2(n3894), .Q(n13016) );
  NAND2X0 U13352 ( .IN1(test_so31), .IN2(n8578), .QN(n3894) );
  INVX0 U13353 ( .INP(n13017), .ZN(n10269) );
  NAND2X0 U13354 ( .IN1(n13018), .IN2(n11799), .QN(n13017) );
  INVX0 U13355 ( .INP(n8578), .ZN(n11799) );
  NOR2X0 U13356 ( .IN1(n10271), .IN2(n13019), .QN(g25027) );
  XNOR2X1 U13357 ( .IN1(n7702), .IN2(n3897), .Q(n13019) );
  NAND2X0 U13358 ( .IN1(g165), .IN2(n8578), .QN(n3897) );
  NOR2X0 U13359 ( .IN1(n13020), .IN2(n8578), .QN(n10271) );
  NAND4X0 U13360 ( .IN1(n7752), .IN2(n4431), .IN3(n13021), .IN4(n4355), .QN(
        n8578) );
  INVX0 U13361 ( .INP(n13022), .ZN(n13021) );
  NAND2X0 U13362 ( .IN1(n4291), .IN2(n4305), .QN(n13022) );
  NAND2X0 U13363 ( .IN1(n3700), .IN2(n13023), .QN(g24734) );
  NAND2X0 U13364 ( .IN1(n11434), .IN2(DFF_146_n1), .QN(n13023) );
  INVX0 U13365 ( .INP(n12471), .ZN(n11434) );
  NAND2X0 U13366 ( .IN1(n3940), .IN2(n3705), .QN(n12471) );
  NAND2X0 U13367 ( .IN1(n13024), .IN2(n13025), .QN(g24557) );
  NAND2X0 U13368 ( .IN1(n9299), .IN2(n9170), .QN(n13025) );
  NAND2X0 U13369 ( .IN1(n4299), .IN2(g2676), .QN(n13024) );
  NAND2X0 U13370 ( .IN1(n13026), .IN2(n13027), .QN(g24548) );
  NAND2X0 U13371 ( .IN1(n4370), .IN2(g2673), .QN(n13027) );
  NAND3X0 U13372 ( .IN1(n9170), .IN2(n10901), .IN3(g7390), .QN(n13026) );
  NAND2X0 U13373 ( .IN1(n13028), .IN2(n13029), .QN(g24547) );
  NAND2X0 U13374 ( .IN1(n9299), .IN2(n10960), .QN(n13029) );
  NOR2X0 U13375 ( .IN1(n10900), .IN2(n4299), .QN(n9299) );
  NAND2X0 U13376 ( .IN1(n4299), .IN2(g2667), .QN(n13028) );
  NAND2X0 U13377 ( .IN1(n13030), .IN2(n13031), .QN(g24545) );
  NAND2X0 U13378 ( .IN1(n9319), .IN2(n11006), .QN(n13031) );
  NAND2X0 U13379 ( .IN1(n4366), .IN2(g1982), .QN(n13030) );
  NAND2X0 U13380 ( .IN1(n13032), .IN2(n13033), .QN(g24538) );
  NAND3X0 U13381 ( .IN1(n9170), .IN2(n10901), .IN3(g7302), .QN(n13033) );
  NAND4X0 U13382 ( .IN1(n13034), .IN2(n13035), .IN3(n13036), .IN4(n13037), 
        .QN(n9170) );
  NAND3X0 U13383 ( .IN1(n9302), .IN2(g185), .IN3(test_so88), .QN(n13037) );
  NAND3X0 U13384 ( .IN1(n13038), .IN2(n13039), .IN3(n13040), .QN(n9302) );
  NAND2X0 U13385 ( .IN1(g7390), .IN2(g2641), .QN(n13040) );
  NAND2X0 U13386 ( .IN1(g2624), .IN2(g2564), .QN(n13039) );
  NAND2X0 U13387 ( .IN1(n10166), .IN2(g2639), .QN(n13038) );
  NAND2X0 U13388 ( .IN1(g2624), .IN2(g2676), .QN(n13036) );
  NAND2X0 U13389 ( .IN1(n10166), .IN2(g2670), .QN(n13035) );
  NAND2X0 U13390 ( .IN1(g7390), .IN2(g2673), .QN(n13034) );
  NAND2X0 U13391 ( .IN1(n4314), .IN2(g2670), .QN(n13032) );
  NAND2X0 U13392 ( .IN1(n13041), .IN2(n13042), .QN(g24537) );
  NAND2X0 U13393 ( .IN1(n4370), .IN2(g2664), .QN(n13042) );
  NAND3X0 U13394 ( .IN1(n10960), .IN2(n10901), .IN3(g7390), .QN(n13041) );
  NAND2X0 U13395 ( .IN1(n13043), .IN2(n13044), .QN(g24535) );
  NAND2X0 U13396 ( .IN1(n4315), .IN2(g1979), .QN(n13044) );
  NAND3X0 U13397 ( .IN1(n11006), .IN2(n10901), .IN3(g7194), .QN(n13043) );
  NAND2X0 U13398 ( .IN1(n13045), .IN2(n13046), .QN(g24534) );
  NAND2X0 U13399 ( .IN1(n9319), .IN2(n11101), .QN(n13046) );
  NOR2X0 U13400 ( .IN1(n10900), .IN2(n4366), .QN(n9319) );
  NAND2X0 U13401 ( .IN1(n4366), .IN2(g1973), .QN(n13045) );
  NAND2X0 U13402 ( .IN1(n13047), .IN2(n13048), .QN(g24532) );
  NAND2X0 U13403 ( .IN1(n8520), .IN2(n11112), .QN(n13048) );
  NAND2X0 U13404 ( .IN1(n4300), .IN2(g1288), .QN(n13047) );
  NAND2X0 U13405 ( .IN1(n13049), .IN2(n13050), .QN(g24527) );
  NAND2X0 U13406 ( .IN1(n4314), .IN2(g2661), .QN(n13050) );
  NAND3X0 U13407 ( .IN1(n10960), .IN2(n10901), .IN3(n10166), .QN(n13049) );
  NAND4X0 U13408 ( .IN1(n13051), .IN2(n13052), .IN3(n13053), .IN4(n13054), 
        .QN(n10960) );
  NAND3X0 U13409 ( .IN1(g185), .IN2(g2598), .IN3(n9301), .QN(n13054) );
  NAND3X0 U13410 ( .IN1(n13055), .IN2(n13056), .IN3(n13057), .QN(n9301) );
  NAND2X0 U13411 ( .IN1(g7390), .IN2(g2645), .QN(n13057) );
  NAND2X0 U13412 ( .IN1(g7302), .IN2(g2643), .QN(n13056) );
  NAND2X0 U13413 ( .IN1(g2624), .IN2(g2647), .QN(n13055) );
  NAND2X0 U13414 ( .IN1(g7302), .IN2(g2661), .QN(n13053) );
  NAND2X0 U13415 ( .IN1(g2624), .IN2(g2667), .QN(n13052) );
  NAND2X0 U13416 ( .IN1(g7390), .IN2(g2664), .QN(n13051) );
  NAND2X0 U13417 ( .IN1(n13058), .IN2(n13059), .QN(g24525) );
  NAND3X0 U13418 ( .IN1(n11006), .IN2(n10901), .IN3(g7052), .QN(n13059) );
  NAND4X0 U13419 ( .IN1(n13060), .IN2(n13061), .IN3(n13062), .IN4(n13063), 
        .QN(n11006) );
  NAND3X0 U13420 ( .IN1(g185), .IN2(g1922), .IN3(n9322), .QN(n13063) );
  NAND3X0 U13421 ( .IN1(n13064), .IN2(n13065), .IN3(n13066), .QN(n9322) );
  NAND2X0 U13422 ( .IN1(g1930), .IN2(g1870), .QN(n13066) );
  NAND2X0 U13423 ( .IN1(n10214), .IN2(g1945), .QN(n13065) );
  NAND2X0 U13424 ( .IN1(g7194), .IN2(g1947), .QN(n13064) );
  NAND2X0 U13425 ( .IN1(n10214), .IN2(g1976), .QN(n13062) );
  NAND2X0 U13426 ( .IN1(g7194), .IN2(g1979), .QN(n13061) );
  NAND2X0 U13427 ( .IN1(g1930), .IN2(g1982), .QN(n13060) );
  NAND2X0 U13428 ( .IN1(n4296), .IN2(g1976), .QN(n13058) );
  NAND2X0 U13429 ( .IN1(n13067), .IN2(n13068), .QN(g24524) );
  NAND2X0 U13430 ( .IN1(n4315), .IN2(g1970), .QN(n13068) );
  NAND3X0 U13431 ( .IN1(n11101), .IN2(n10901), .IN3(g7194), .QN(n13067) );
  NAND2X0 U13432 ( .IN1(n13069), .IN2(n13070), .QN(g24522) );
  NAND2X0 U13433 ( .IN1(n4316), .IN2(g1285), .QN(n13070) );
  NAND3X0 U13434 ( .IN1(n11112), .IN2(n10901), .IN3(g6944), .QN(n13069) );
  NAND2X0 U13435 ( .IN1(n13071), .IN2(n13072), .QN(g24521) );
  NAND2X0 U13436 ( .IN1(n8520), .IN2(n11204), .QN(n13072) );
  NOR2X0 U13437 ( .IN1(n10900), .IN2(n4300), .QN(n8520) );
  NAND2X0 U13438 ( .IN1(n4300), .IN2(g1279), .QN(n13071) );
  NAND2X0 U13439 ( .IN1(n13073), .IN2(n13074), .QN(g24519) );
  NAND2X0 U13440 ( .IN1(n8541), .IN2(n11215), .QN(n13074) );
  NAND2X0 U13441 ( .IN1(n4313), .IN2(g602), .QN(n13073) );
  NAND2X0 U13442 ( .IN1(n13075), .IN2(n13076), .QN(g24513) );
  NAND2X0 U13443 ( .IN1(n4296), .IN2(g1967), .QN(n13076) );
  NAND3X0 U13444 ( .IN1(n11101), .IN2(n10901), .IN3(n10214), .QN(n13075) );
  NAND4X0 U13445 ( .IN1(n13077), .IN2(n13078), .IN3(n13079), .IN4(n13080), 
        .QN(n11101) );
  NAND3X0 U13446 ( .IN1(g185), .IN2(g1904), .IN3(n9321), .QN(n13080) );
  NAND3X0 U13447 ( .IN1(n13081), .IN2(n13082), .IN3(n13083), .QN(n9321) );
  NAND2X0 U13448 ( .IN1(g1930), .IN2(g1953), .QN(n13083) );
  NAND2X0 U13449 ( .IN1(g7052), .IN2(g1949), .QN(n13082) );
  NAND2X0 U13450 ( .IN1(g7194), .IN2(g1951), .QN(n13081) );
  NAND2X0 U13451 ( .IN1(g7052), .IN2(g1967), .QN(n13079) );
  NAND2X0 U13452 ( .IN1(g7194), .IN2(g1970), .QN(n13078) );
  NAND2X0 U13453 ( .IN1(g1930), .IN2(g1973), .QN(n13077) );
  NAND2X0 U13454 ( .IN1(n13084), .IN2(n13085), .QN(g24511) );
  NAND3X0 U13455 ( .IN1(n11112), .IN2(n10901), .IN3(g6750), .QN(n13085) );
  NAND4X0 U13456 ( .IN1(n13086), .IN2(n13087), .IN3(n13088), .IN4(n13089), 
        .QN(n11112) );
  NAND3X0 U13457 ( .IN1(n8522), .IN2(g185), .IN3(test_so45), .QN(n13089) );
  NAND3X0 U13458 ( .IN1(n13090), .IN2(n13091), .IN3(n13092), .QN(n8522) );
  NAND2X0 U13459 ( .IN1(g6944), .IN2(g1253), .QN(n13092) );
  NAND2X0 U13460 ( .IN1(g6750), .IN2(g1251), .QN(n13091) );
  NAND2X0 U13461 ( .IN1(g1236), .IN2(g1176), .QN(n13090) );
  NAND2X0 U13462 ( .IN1(g1236), .IN2(g1288), .QN(n13088) );
  NAND2X0 U13463 ( .IN1(g6944), .IN2(g1285), .QN(n13087) );
  NAND2X0 U13464 ( .IN1(n11104), .IN2(g1282), .QN(n13086) );
  NAND2X0 U13465 ( .IN1(n4371), .IN2(g1282), .QN(n13084) );
  NAND2X0 U13466 ( .IN1(n13093), .IN2(n13094), .QN(g24510) );
  NAND2X0 U13467 ( .IN1(n4316), .IN2(g1276), .QN(n13094) );
  NAND3X0 U13468 ( .IN1(n11204), .IN2(n10901), .IN3(g6944), .QN(n13093) );
  NAND2X0 U13469 ( .IN1(n13095), .IN2(n13096), .QN(g24508) );
  NAND2X0 U13470 ( .IN1(n4372), .IN2(g599), .QN(n13096) );
  NAND3X0 U13471 ( .IN1(n11215), .IN2(n10901), .IN3(g6642), .QN(n13095) );
  NAND2X0 U13472 ( .IN1(n13097), .IN2(n13098), .QN(g24507) );
  NAND2X0 U13473 ( .IN1(n8541), .IN2(n11302), .QN(n13098) );
  NOR2X0 U13474 ( .IN1(n10900), .IN2(n4313), .QN(n8541) );
  NAND2X0 U13475 ( .IN1(n4313), .IN2(g593), .QN(n13097) );
  NAND2X0 U13476 ( .IN1(n13099), .IN2(n13100), .QN(g24501) );
  NAND2X0 U13477 ( .IN1(n4371), .IN2(g1273), .QN(n13100) );
  NAND3X0 U13478 ( .IN1(n11204), .IN2(n10901), .IN3(n11104), .QN(n13099) );
  NAND4X0 U13479 ( .IN1(n13101), .IN2(n13102), .IN3(n13103), .IN4(n13104), 
        .QN(n11204) );
  NAND3X0 U13480 ( .IN1(g185), .IN2(g1210), .IN3(n8523), .QN(n13104) );
  NAND3X0 U13481 ( .IN1(n13105), .IN2(n13106), .IN3(n13107), .QN(n8523) );
  NAND2X0 U13482 ( .IN1(n11104), .IN2(g1255), .QN(n13107) );
  NAND2X0 U13483 ( .IN1(g1236), .IN2(g1259), .QN(n13106) );
  NAND2X0 U13484 ( .IN1(g6944), .IN2(g1257), .QN(n13105) );
  NAND2X0 U13485 ( .IN1(g6750), .IN2(g1273), .QN(n13103) );
  NAND2X0 U13486 ( .IN1(g1236), .IN2(g1279), .QN(n13102) );
  NAND2X0 U13487 ( .IN1(g6944), .IN2(g1276), .QN(n13101) );
  NAND2X0 U13488 ( .IN1(n13108), .IN2(n13109), .QN(g24499) );
  NAND3X0 U13489 ( .IN1(n11215), .IN2(n10901), .IN3(g6485), .QN(n13109) );
  NAND4X0 U13490 ( .IN1(n13110), .IN2(n13111), .IN3(n13112), .IN4(n13113), 
        .QN(n11215) );
  NAND3X0 U13491 ( .IN1(g185), .IN2(g542), .IN3(n8546), .QN(n13113) );
  NAND3X0 U13492 ( .IN1(n13114), .IN2(n13115), .IN3(n13116), .QN(n8546) );
  NAND2X0 U13493 ( .IN1(g6642), .IN2(g567), .QN(n13116) );
  NAND2X0 U13494 ( .IN1(n11207), .IN2(g565), .QN(n13115) );
  NAND2X0 U13495 ( .IN1(g550), .IN2(g489), .QN(n13114) );
  NAND2X0 U13496 ( .IN1(g6485), .IN2(g596), .QN(n13112) );
  NAND2X0 U13497 ( .IN1(g550), .IN2(g602), .QN(n13111) );
  NAND2X0 U13498 ( .IN1(g6642), .IN2(g599), .QN(n13110) );
  NAND2X0 U13499 ( .IN1(n4298), .IN2(g596), .QN(n13108) );
  NAND2X0 U13500 ( .IN1(n13117), .IN2(n13118), .QN(g24498) );
  NAND2X0 U13501 ( .IN1(n4372), .IN2(g590), .QN(n13118) );
  NAND3X0 U13502 ( .IN1(n11302), .IN2(n10901), .IN3(g6642), .QN(n13117) );
  NAND2X0 U13503 ( .IN1(n13119), .IN2(n13120), .QN(g24491) );
  NAND2X0 U13504 ( .IN1(n4298), .IN2(g587), .QN(n13120) );
  NAND3X0 U13505 ( .IN1(n11302), .IN2(n10901), .IN3(n11207), .QN(n13119) );
  INVX0 U13506 ( .INP(n10900), .ZN(n10901) );
  NOR4X0 U13507 ( .IN1(n4350), .IN2(n4481), .IN3(n13121), .IN4(n13122), .QN(
        n10900) );
  NAND2X0 U13508 ( .IN1(n4480), .IN2(n7429), .QN(n13122) );
  NAND4X0 U13509 ( .IN1(n13123), .IN2(n13124), .IN3(n13125), .IN4(n13126), 
        .QN(n11302) );
  NAND3X0 U13510 ( .IN1(g185), .IN2(g524), .IN3(n8543), .QN(n13126) );
  NAND3X0 U13511 ( .IN1(n13127), .IN2(n13128), .IN3(n13129), .QN(n8543) );
  NAND2X0 U13512 ( .IN1(g6642), .IN2(g571), .QN(n13129) );
  NAND2X0 U13513 ( .IN1(g6485), .IN2(g569), .QN(n13128) );
  NAND2X0 U13514 ( .IN1(g550), .IN2(g573), .QN(n13127) );
  NAND2X0 U13515 ( .IN1(n11207), .IN2(g587), .QN(n13125) );
  NAND2X0 U13516 ( .IN1(g550), .IN2(g593), .QN(n13124) );
  NAND2X0 U13517 ( .IN1(g6642), .IN2(g590), .QN(n13123) );
  NOR3X0 U13518 ( .IN1(n13130), .IN2(n13004), .IN3(n13002), .QN(g24476) );
  NOR3X0 U13519 ( .IN1(n4349), .IN2(n4479), .IN3(n8676), .QN(n13004) );
  NOR2X0 U13520 ( .IN1(n13131), .IN2(g2924), .QN(n13130) );
  NOR2X0 U13521 ( .IN1(n4479), .IN2(n8676), .QN(n13131) );
  NOR2X0 U13522 ( .IN1(n8672), .IN2(n13132), .QN(g24473) );
  XOR2X1 U13523 ( .IN1(n7752), .IN2(n13001), .Q(n13132) );
  NOR3X0 U13524 ( .IN1(n13000), .IN2(n4101), .IN3(n12998), .QN(g24446) );
  INVX0 U13525 ( .INP(n8728), .ZN(n12998) );
  NAND2X0 U13526 ( .IN1(n12153), .IN2(n13133), .QN(n8728) );
  NAND2X0 U13527 ( .IN1(n13134), .IN2(n8726), .QN(n13133) );
  INVX0 U13528 ( .INP(g3234), .ZN(n8726) );
  NAND4X0 U13529 ( .IN1(n4350), .IN2(n4480), .IN3(g3018), .IN4(g3032), .QN(
        n13134) );
  NOR2X0 U13530 ( .IN1(n1543), .IN2(n4480), .QN(n13000) );
  NAND3X0 U13531 ( .IN1(g3028), .IN2(g3018), .IN3(n8729), .QN(n1543) );
  NOR2X0 U13532 ( .IN1(n12153), .IN2(n13135), .QN(g24445) );
  XNOR2X1 U13533 ( .IN1(n8034), .IN2(n4066), .Q(n13135) );
  NAND3X0 U13534 ( .IN1(g3006), .IN2(n7909), .IN3(n9286), .QN(n4066) );
  NOR2X0 U13535 ( .IN1(n8032), .IN2(n8031), .QN(n9286) );
  INVX0 U13536 ( .INP(n9283), .ZN(n12153) );
  NOR2X0 U13537 ( .IN1(g3234), .IN2(n8729), .QN(n9283) );
  NOR2X0 U13538 ( .IN1(n13121), .IN2(n8031), .QN(n8729) );
  NAND4X0 U13539 ( .IN1(n8032), .IN2(g3024), .IN3(n8035), .IN4(n13136), .QN(
        n13121) );
  NOR4X0 U13540 ( .IN1(test_so98), .IN2(n14354), .IN3(n8051), .IN4(n8034), 
        .QN(n13136) );
  NOR3X0 U13541 ( .IN1(n13137), .IN2(n11303), .IN3(n9292), .QN(g24438) );
  NOR3X0 U13542 ( .IN1(n4408), .IN2(n4419), .IN3(n9295), .QN(n9292) );
  NOR2X0 U13543 ( .IN1(n13138), .IN2(g2720), .QN(n13137) );
  NOR2X0 U13544 ( .IN1(n4419), .IN2(n9295), .QN(n13138) );
  NOR3X0 U13545 ( .IN1(n13139), .IN2(n9305), .IN3(n12151), .QN(g24434) );
  NOR3X0 U13546 ( .IN1(n4410), .IN2(n4420), .IN3(n9312), .QN(n12151) );
  NOR2X0 U13547 ( .IN1(n13140), .IN2(g2026), .QN(n13139) );
  NOR2X0 U13548 ( .IN1(n4420), .IN2(n9312), .QN(n13140) );
  NOR3X0 U13549 ( .IN1(n13141), .IN2(n8512), .IN3(n8510), .QN(g24430) );
  NOR3X0 U13550 ( .IN1(n4412), .IN2(n4421), .IN3(n13142), .QN(n8510) );
  NOR2X0 U13551 ( .IN1(n13143), .IN2(g1332), .QN(n13141) );
  NOR2X0 U13552 ( .IN1(n4421), .IN2(n13142), .QN(n13143) );
  INVX0 U13553 ( .INP(n8513), .ZN(n13142) );
  NOR3X0 U13554 ( .IN1(n13144), .IN2(n8536), .IN3(n8530), .QN(g24426) );
  NOR3X0 U13555 ( .IN1(n4414), .IN2(n4422), .IN3(n8533), .QN(n8530) );
  NOR2X0 U13556 ( .IN1(n13145), .IN2(g646), .QN(n13144) );
  NOR2X0 U13557 ( .IN1(n4422), .IN2(n8533), .QN(n13145) );
  NAND2X0 U13558 ( .IN1(n13146), .IN2(n13147), .QN(g24250) );
  NAND2X0 U13559 ( .IN1(n4463), .IN2(g2546), .QN(n13147) );
  NAND2X0 U13560 ( .IN1(n10016), .IN2(g2560), .QN(n13146) );
  NAND2X0 U13561 ( .IN1(n13148), .IN2(n13149), .QN(g24243) );
  NAND2X0 U13562 ( .IN1(n4464), .IN2(g1852), .QN(n13149) );
  NAND2X0 U13563 ( .IN1(n8615), .IN2(g1866), .QN(n13148) );
  NAND2X0 U13564 ( .IN1(n13150), .IN2(n13151), .QN(g24238) );
  NAND2X0 U13565 ( .IN1(n4463), .IN2(g2554), .QN(n13151) );
  NAND2X0 U13566 ( .IN1(n10019), .IN2(g2560), .QN(n13150) );
  NAND2X0 U13567 ( .IN1(n13152), .IN2(n13153), .QN(g24237) );
  NAND2X0 U13568 ( .IN1(n4455), .IN2(g2543), .QN(n13153) );
  NAND2X0 U13569 ( .IN1(n10016), .IN2(g8167), .QN(n13152) );
  NAND2X0 U13570 ( .IN1(n13154), .IN2(n13155), .QN(g24235) );
  NAND2X0 U13571 ( .IN1(n4465), .IN2(g1158), .QN(n13155) );
  NAND2X0 U13572 ( .IN1(n10106), .IN2(g1172), .QN(n13154) );
  NAND2X0 U13573 ( .IN1(n13156), .IN2(n13157), .QN(g24231) );
  NAND2X0 U13574 ( .IN1(n4464), .IN2(g1860), .QN(n13157) );
  NAND2X0 U13575 ( .IN1(n10066), .IN2(g1866), .QN(n13156) );
  NAND2X0 U13576 ( .IN1(n13158), .IN2(n13159), .QN(g24230) );
  NAND2X0 U13577 ( .IN1(n4457), .IN2(g1849), .QN(n13159) );
  NAND2X0 U13578 ( .IN1(n8615), .IN2(g8082), .QN(n13158) );
  NAND2X0 U13579 ( .IN1(n13160), .IN2(n13161), .QN(g24228) );
  NAND2X0 U13580 ( .IN1(n4466), .IN2(g471), .QN(n13161) );
  NAND2X0 U13581 ( .IN1(n8555), .IN2(g485), .QN(n13160) );
  NAND2X0 U13582 ( .IN1(n13162), .IN2(n13163), .QN(g24226) );
  NAND2X0 U13583 ( .IN1(n4455), .IN2(g2553), .QN(n13163) );
  NAND2X0 U13584 ( .IN1(n10019), .IN2(g8167), .QN(n13162) );
  NAND2X0 U13585 ( .IN1(n13164), .IN2(n13165), .QN(g24225) );
  NAND2X0 U13586 ( .IN1(n4456), .IN2(g2540), .QN(n13165) );
  NAND2X0 U13587 ( .IN1(n10016), .IN2(g8087), .QN(n13164) );
  NOR2X0 U13588 ( .IN1(n9704), .IN2(n9708), .QN(n10016) );
  NAND2X0 U13589 ( .IN1(n9709), .IN2(n9715), .QN(n9704) );
  INVX0 U13590 ( .INP(n9724), .ZN(n9709) );
  NAND2X0 U13591 ( .IN1(n13166), .IN2(n13167), .QN(g24223) );
  NAND2X0 U13592 ( .IN1(n4465), .IN2(g1166), .QN(n13167) );
  NAND2X0 U13593 ( .IN1(n10110), .IN2(g1172), .QN(n13166) );
  NAND2X0 U13594 ( .IN1(n13168), .IN2(n13169), .QN(g24222) );
  NAND2X0 U13595 ( .IN1(n4459), .IN2(g1155), .QN(n13169) );
  NAND2X0 U13596 ( .IN1(n10106), .IN2(g8007), .QN(n13168) );
  NAND2X0 U13597 ( .IN1(n13170), .IN2(n13171), .QN(g24219) );
  NAND2X0 U13598 ( .IN1(n4457), .IN2(g1859), .QN(n13171) );
  NAND2X0 U13599 ( .IN1(n10066), .IN2(g8082), .QN(n13170) );
  NAND2X0 U13600 ( .IN1(n13172), .IN2(n13173), .QN(g24218) );
  NAND2X0 U13601 ( .IN1(n4458), .IN2(g1846), .QN(n13173) );
  NAND2X0 U13602 ( .IN1(n8615), .IN2(g8012), .QN(n13172) );
  NOR2X0 U13603 ( .IN1(n9352), .IN2(n9356), .QN(n8615) );
  NAND2X0 U13604 ( .IN1(n9357), .IN2(n9363), .QN(n9352) );
  INVX0 U13605 ( .INP(n9372), .ZN(n9357) );
  NAND2X0 U13606 ( .IN1(n13174), .IN2(n13175), .QN(g24216) );
  NAND2X0 U13607 ( .IN1(n4466), .IN2(g479), .QN(n13175) );
  NAND2X0 U13608 ( .IN1(n10150), .IN2(g485), .QN(n13174) );
  NAND2X0 U13609 ( .IN1(n13176), .IN2(n13177), .QN(g24215) );
  NAND2X0 U13610 ( .IN1(n8555), .IN2(g7956), .QN(n13177) );
  NAND2X0 U13611 ( .IN1(test_so24), .IN2(n4461), .QN(n13176) );
  NAND2X0 U13612 ( .IN1(n13178), .IN2(n13179), .QN(g24214) );
  NAND2X0 U13613 ( .IN1(n4456), .IN2(g2552), .QN(n13179) );
  NAND2X0 U13614 ( .IN1(n10019), .IN2(g8087), .QN(n13178) );
  INVX0 U13615 ( .INP(n10230), .ZN(n10019) );
  NAND3X0 U13616 ( .IN1(n9708), .IN2(n9724), .IN3(n9715), .QN(n10230) );
  INVX0 U13617 ( .INP(n9699), .ZN(n9715) );
  NAND2X0 U13618 ( .IN1(n13180), .IN2(n13181), .QN(g24213) );
  NAND2X0 U13619 ( .IN1(n4459), .IN2(g1165), .QN(n13181) );
  NAND2X0 U13620 ( .IN1(n10110), .IN2(g8007), .QN(n13180) );
  NAND2X0 U13621 ( .IN1(n13182), .IN2(n13183), .QN(g24212) );
  NAND2X0 U13622 ( .IN1(n4460), .IN2(g1152), .QN(n13183) );
  NAND2X0 U13623 ( .IN1(n10106), .IN2(g7961), .QN(n13182) );
  NOR2X0 U13624 ( .IN1(n9194), .IN2(n9179), .QN(n10106) );
  NAND2X0 U13625 ( .IN1(n9173), .IN2(n9183), .QN(n9194) );
  INVX0 U13626 ( .INP(n9185), .ZN(n9173) );
  NAND2X0 U13627 ( .IN1(n13184), .IN2(n13185), .QN(g24209) );
  NAND2X0 U13628 ( .IN1(n4463), .IN2(g2536), .QN(n13185) );
  NAND2X0 U13629 ( .IN1(n13186), .IN2(g2560), .QN(n13184) );
  NAND2X0 U13630 ( .IN1(n13187), .IN2(n13188), .QN(g24208) );
  NAND2X0 U13631 ( .IN1(n4458), .IN2(g1858), .QN(n13188) );
  NAND2X0 U13632 ( .IN1(n10066), .IN2(g8012), .QN(n13187) );
  INVX0 U13633 ( .INP(n10243), .ZN(n10066) );
  NAND3X0 U13634 ( .IN1(n9356), .IN2(n9372), .IN3(n9363), .QN(n10243) );
  INVX0 U13635 ( .INP(n9347), .ZN(n9363) );
  NAND2X0 U13636 ( .IN1(n13189), .IN2(n13190), .QN(g24207) );
  NAND2X0 U13637 ( .IN1(n4461), .IN2(g478), .QN(n13190) );
  NAND2X0 U13638 ( .IN1(n10150), .IN2(g7956), .QN(n13189) );
  NAND2X0 U13639 ( .IN1(n13191), .IN2(n13192), .QN(g24206) );
  NAND2X0 U13640 ( .IN1(g465), .IN2(n8072), .QN(n13192) );
  NAND2X0 U13641 ( .IN1(test_so23), .IN2(n8555), .QN(n13191) );
  NOR2X0 U13642 ( .IN1(n9394), .IN2(n9398), .QN(n8555) );
  NAND2X0 U13643 ( .IN1(n9399), .IN2(n9405), .QN(n9394) );
  INVX0 U13644 ( .INP(n9414), .ZN(n9399) );
  NAND2X0 U13645 ( .IN1(n13193), .IN2(n13194), .QN(g24182) );
  NAND2X0 U13646 ( .IN1(n4464), .IN2(g1842), .QN(n13194) );
  NAND2X0 U13647 ( .IN1(n11889), .IN2(g1866), .QN(n13193) );
  NAND2X0 U13648 ( .IN1(n13195), .IN2(n13196), .QN(g24181) );
  NAND2X0 U13649 ( .IN1(n4460), .IN2(g1164), .QN(n13196) );
  NAND2X0 U13650 ( .IN1(n10110), .IN2(g7961), .QN(n13195) );
  INVX0 U13651 ( .INP(n10547), .ZN(n10110) );
  NAND3X0 U13652 ( .IN1(n9179), .IN2(n9185), .IN3(n9183), .QN(n10547) );
  INVX0 U13653 ( .INP(n9181), .ZN(n9183) );
  NAND2X0 U13654 ( .IN1(n13197), .IN2(n13198), .QN(g24179) );
  NAND2X0 U13655 ( .IN1(n4465), .IN2(g1148), .QN(n13198) );
  NAND2X0 U13656 ( .IN1(n13199), .IN2(g1172), .QN(n13197) );
  NAND2X0 U13657 ( .IN1(n13200), .IN2(n13201), .QN(g24178) );
  NAND2X0 U13658 ( .IN1(g477), .IN2(n8072), .QN(n13201) );
  NAND2X0 U13659 ( .IN1(test_so23), .IN2(n10150), .QN(n13200) );
  INVX0 U13660 ( .INP(n10263), .ZN(n10150) );
  NAND3X0 U13661 ( .IN1(n9398), .IN2(n9414), .IN3(n9405), .QN(n10263) );
  INVX0 U13662 ( .INP(n9389), .ZN(n9405) );
  NAND2X0 U13663 ( .IN1(n13202), .IN2(n13203), .QN(g24174) );
  NAND2X0 U13664 ( .IN1(n4466), .IN2(g461), .QN(n13203) );
  NAND2X0 U13665 ( .IN1(n11987), .IN2(g485), .QN(n13202) );
  NAND2X0 U13666 ( .IN1(n13204), .IN2(n13205), .QN(g24092) );
  NAND2X0 U13667 ( .IN1(g3229), .IN2(n4483), .QN(n13205) );
  NAND2X0 U13668 ( .IN1(n8785), .IN2(g2380), .QN(n13204) );
  NAND2X0 U13669 ( .IN1(n13206), .IN2(n13207), .QN(g24083) );
  NAND2X0 U13670 ( .IN1(g3229), .IN2(n4484), .QN(n13207) );
  NAND2X0 U13671 ( .IN1(n8785), .IN2(g1686), .QN(n13206) );
  NAND2X0 U13672 ( .IN1(n13208), .IN2(n13209), .QN(g24072) );
  NAND2X0 U13673 ( .IN1(g3229), .IN2(n4486), .QN(n13209) );
  NAND2X0 U13674 ( .IN1(n8785), .IN2(g992), .QN(n13208) );
  NAND2X0 U13675 ( .IN1(n13210), .IN2(n13211), .QN(g24059) );
  NAND2X0 U13676 ( .IN1(g3229), .IN2(n4485), .QN(n13211) );
  NAND2X0 U13677 ( .IN1(n8785), .IN2(g305), .QN(n13210) );
  INVX0 U13678 ( .INP(g3229), .ZN(n8785) );
  NAND2X0 U13679 ( .IN1(n13212), .IN2(n13213), .QN(g23418) );
  NAND2X0 U13680 ( .IN1(n4455), .IN2(g2533), .QN(n13213) );
  NAND2X0 U13681 ( .IN1(n13186), .IN2(g8167), .QN(n13212) );
  NAND2X0 U13682 ( .IN1(n13214), .IN2(n13215), .QN(g23413) );
  NAND2X0 U13683 ( .IN1(n11889), .IN2(g8082), .QN(n13215) );
  NAND2X0 U13684 ( .IN1(test_so65), .IN2(n4457), .QN(n13214) );
  NAND2X0 U13685 ( .IN1(n13216), .IN2(n13217), .QN(g23407) );
  NAND2X0 U13686 ( .IN1(n4456), .IN2(g2530), .QN(n13217) );
  NAND2X0 U13687 ( .IN1(n13186), .IN2(g8087), .QN(n13216) );
  INVX0 U13688 ( .INP(n8667), .ZN(n13186) );
  NAND3X0 U13689 ( .IN1(n9699), .IN2(n9724), .IN3(n9703), .QN(n8667) );
  INVX0 U13690 ( .INP(n9708), .ZN(n9703) );
  NAND3X0 U13691 ( .IN1(n13218), .IN2(n13219), .IN3(n13220), .QN(n9708) );
  NAND2X0 U13692 ( .IN1(n7258), .IN2(n10027), .QN(n13220) );
  NAND2X0 U13693 ( .IN1(n7269), .IN2(n10028), .QN(n13219) );
  NAND2X0 U13694 ( .IN1(n7270), .IN2(n10029), .QN(n13218) );
  NAND3X0 U13695 ( .IN1(n13221), .IN2(n13222), .IN3(n13223), .QN(n9724) );
  NAND2X0 U13696 ( .IN1(n7256), .IN2(n10027), .QN(n13223) );
  NAND2X0 U13697 ( .IN1(n7265), .IN2(n10028), .QN(n13222) );
  NAND2X0 U13698 ( .IN1(n7266), .IN2(n10029), .QN(n13221) );
  NAND3X0 U13699 ( .IN1(n13224), .IN2(n13225), .IN3(n13226), .QN(n9699) );
  NAND2X0 U13700 ( .IN1(n7257), .IN2(n10027), .QN(n13226) );
  INVX0 U13701 ( .INP(n4524), .ZN(n10027) );
  NAND2X0 U13702 ( .IN1(n7267), .IN2(n10028), .QN(n13225) );
  INVX0 U13703 ( .INP(n4509), .ZN(n10028) );
  NAND2X0 U13704 ( .IN1(n7268), .IN2(n10029), .QN(n13224) );
  INVX0 U13705 ( .INP(n4516), .ZN(n10029) );
  NAND2X0 U13706 ( .IN1(n13227), .IN2(n13228), .QN(g23406) );
  NAND2X0 U13707 ( .IN1(n4459), .IN2(g1145), .QN(n13228) );
  NAND2X0 U13708 ( .IN1(n13199), .IN2(g8007), .QN(n13227) );
  NAND2X0 U13709 ( .IN1(n13229), .IN2(n13230), .QN(g23400) );
  NAND2X0 U13710 ( .IN1(n4458), .IN2(g1836), .QN(n13230) );
  NAND2X0 U13711 ( .IN1(n11889), .IN2(g8012), .QN(n13229) );
  INVX0 U13712 ( .INP(n8631), .ZN(n11889) );
  NAND3X0 U13713 ( .IN1(n9347), .IN2(n9372), .IN3(n9351), .QN(n8631) );
  INVX0 U13714 ( .INP(n9356), .ZN(n9351) );
  NAND3X0 U13715 ( .IN1(n13231), .IN2(n13232), .IN3(n13233), .QN(n9356) );
  NAND2X0 U13716 ( .IN1(n7261), .IN2(n10074), .QN(n13233) );
  NAND2X0 U13717 ( .IN1(n7275), .IN2(n10075), .QN(n13232) );
  NAND2X0 U13718 ( .IN1(n7276), .IN2(n10076), .QN(n13231) );
  NAND3X0 U13719 ( .IN1(n13234), .IN2(n13235), .IN3(n13236), .QN(n9372) );
  NAND2X0 U13720 ( .IN1(n7259), .IN2(n10074), .QN(n13236) );
  NAND2X0 U13721 ( .IN1(n7271), .IN2(n10075), .QN(n13235) );
  NAND2X0 U13722 ( .IN1(n7272), .IN2(n10076), .QN(n13234) );
  NAND3X0 U13723 ( .IN1(n13237), .IN2(n13238), .IN3(n13239), .QN(n9347) );
  NAND2X0 U13724 ( .IN1(n7260), .IN2(n10074), .QN(n13239) );
  INVX0 U13725 ( .INP(n4525), .ZN(n10074) );
  NAND2X0 U13726 ( .IN1(n7273), .IN2(n10075), .QN(n13238) );
  INVX0 U13727 ( .INP(n4511), .ZN(n10075) );
  NAND2X0 U13728 ( .IN1(n7274), .IN2(n10076), .QN(n13237) );
  INVX0 U13729 ( .INP(n4518), .ZN(n10076) );
  NAND2X0 U13730 ( .IN1(n13240), .IN2(n13241), .QN(g23399) );
  NAND2X0 U13731 ( .IN1(n4461), .IN2(g458), .QN(n13241) );
  NAND2X0 U13732 ( .IN1(n11987), .IN2(g7956), .QN(n13240) );
  NAND2X0 U13733 ( .IN1(n13242), .IN2(n13243), .QN(g23392) );
  NAND2X0 U13734 ( .IN1(n4460), .IN2(g1142), .QN(n13243) );
  NAND2X0 U13735 ( .IN1(n13199), .IN2(g7961), .QN(n13242) );
  INVX0 U13736 ( .INP(n8608), .ZN(n13199) );
  NAND3X0 U13737 ( .IN1(n9181), .IN2(n9185), .IN3(n9193), .QN(n8608) );
  INVX0 U13738 ( .INP(n9179), .ZN(n9193) );
  NAND3X0 U13739 ( .IN1(n13244), .IN2(n13245), .IN3(n13246), .QN(n9179) );
  NAND2X0 U13740 ( .IN1(n7280), .IN2(g1088), .QN(n13246) );
  NAND2X0 U13741 ( .IN1(n7281), .IN2(g5472), .QN(n13245) );
  NAND2X0 U13742 ( .IN1(n7264), .IN2(g6712), .QN(n13244) );
  NAND3X0 U13743 ( .IN1(n13247), .IN2(n13248), .IN3(n13249), .QN(n9185) );
  NAND2X0 U13744 ( .IN1(g1088), .IN2(n8127), .QN(n13249) );
  NAND2X0 U13745 ( .IN1(n7277), .IN2(g5472), .QN(n13248) );
  NAND2X0 U13746 ( .IN1(n7262), .IN2(g6712), .QN(n13247) );
  NAND3X0 U13747 ( .IN1(n13250), .IN2(n13251), .IN3(n13252), .QN(n9181) );
  NAND2X0 U13748 ( .IN1(n7278), .IN2(g1088), .QN(n13252) );
  NAND2X0 U13749 ( .IN1(n7279), .IN2(g5472), .QN(n13251) );
  NAND2X0 U13750 ( .IN1(n7263), .IN2(g6712), .QN(n13250) );
  NAND2X0 U13751 ( .IN1(n13253), .IN2(n13254), .QN(g23385) );
  NAND2X0 U13752 ( .IN1(g455), .IN2(n8072), .QN(n13254) );
  NAND2X0 U13753 ( .IN1(n11987), .IN2(test_so23), .QN(n13253) );
  INVX0 U13754 ( .INP(n8579), .ZN(n11987) );
  NAND3X0 U13755 ( .IN1(n9389), .IN2(n9414), .IN3(n9393), .QN(n8579) );
  INVX0 U13756 ( .INP(n9398), .ZN(n9393) );
  NAND3X0 U13757 ( .IN1(n13255), .IN2(n13256), .IN3(n13257), .QN(n9398) );
  NAND2X0 U13758 ( .IN1(n7289), .IN2(n10158), .QN(n13257) );
  NAND2X0 U13759 ( .IN1(n7288), .IN2(n10159), .QN(n13256) );
  NAND2X0 U13760 ( .IN1(n7287), .IN2(n10160), .QN(n13255) );
  NAND3X0 U13761 ( .IN1(n13258), .IN2(n13259), .IN3(n13260), .QN(n9414) );
  NAND2X0 U13762 ( .IN1(n7284), .IN2(n10158), .QN(n13260) );
  NAND2X0 U13763 ( .IN1(n7283), .IN2(n10159), .QN(n13259) );
  NAND2X0 U13764 ( .IN1(n7282), .IN2(n10160), .QN(n13258) );
  NAND3X0 U13765 ( .IN1(n13261), .IN2(n13262), .IN3(n13263), .QN(n9389) );
  NAND2X0 U13766 ( .IN1(n7286), .IN2(n10158), .QN(n13263) );
  INVX0 U13767 ( .INP(n4520), .ZN(n10158) );
  NAND2X0 U13768 ( .IN1(n10159), .IN2(n8128), .QN(n13262) );
  INVX0 U13769 ( .INP(n4499), .ZN(n10159) );
  NAND2X0 U13770 ( .IN1(n7285), .IN2(n10160), .QN(n13261) );
  INVX0 U13771 ( .INP(n4506), .ZN(n10160) );
  NOR3X0 U13772 ( .IN1(n8672), .IN2(n4122), .IN3(n13001), .QN(g23358) );
  NOR2X0 U13773 ( .IN1(n10), .IN2(n4431), .QN(n13001) );
  NAND2X0 U13774 ( .IN1(n13264), .IN2(g2888), .QN(n10) );
  NOR2X0 U13775 ( .IN1(n13002), .IN2(n13265), .QN(g23357) );
  XOR2X1 U13776 ( .IN1(g2917), .IN2(n8676), .Q(n13265) );
  NAND2X0 U13777 ( .IN1(n13266), .IN2(g2912), .QN(n8676) );
  INVX0 U13778 ( .INP(n8677), .ZN(n13266) );
  INVX0 U13779 ( .INP(n8673), .ZN(n13002) );
  NAND2X0 U13780 ( .IN1(n8672), .IN2(n13267), .QN(n8673) );
  NAND2X0 U13781 ( .IN1(n14350), .IN2(n13268), .QN(n13267) );
  NAND4X0 U13782 ( .IN1(n4479), .IN2(n4349), .IN3(g2912), .IN4(g2920), .QN(
        n13268) );
  NOR2X0 U13783 ( .IN1(n11303), .IN2(n13269), .QN(g23348) );
  XNOR2X1 U13784 ( .IN1(n4419), .IN2(n9295), .Q(n13269) );
  NAND3X0 U13785 ( .IN1(g2714), .IN2(g2707), .IN3(n9297), .QN(n9295) );
  NOR2X0 U13786 ( .IN1(n9305), .IN2(n13270), .QN(g23339) );
  XNOR2X1 U13787 ( .IN1(n4420), .IN2(n9312), .Q(n13270) );
  NAND3X0 U13788 ( .IN1(g2020), .IN2(g2013), .IN3(n9314), .QN(n9312) );
  NOR2X0 U13789 ( .IN1(n8512), .IN2(n13271), .QN(g23329) );
  XOR2X1 U13790 ( .IN1(n4421), .IN2(n8513), .Q(n13271) );
  NOR3X0 U13791 ( .IN1(n4402), .IN2(n4476), .IN3(n8515), .QN(n8513) );
  NOR2X0 U13792 ( .IN1(n8536), .IN2(n13272), .QN(g23324) );
  XNOR2X1 U13793 ( .IN1(n4422), .IN2(n8533), .Q(n13272) );
  NAND3X0 U13794 ( .IN1(g640), .IN2(g633), .IN3(n8535), .QN(n8533) );
  NAND2X0 U13795 ( .IN1(n13273), .IN2(n13274), .QN(g23137) );
  NAND2X0 U13796 ( .IN1(n4464), .IN2(g1869), .QN(n13274) );
  NAND2X0 U13797 ( .IN1(n11359), .IN2(g1866), .QN(n13273) );
  NAND2X0 U13798 ( .IN1(n13275), .IN2(n13276), .QN(g23133) );
  NAND2X0 U13799 ( .IN1(n4455), .IN2(g2562), .QN(n13276) );
  NAND2X0 U13800 ( .IN1(n11339), .IN2(g8167), .QN(n13275) );
  NAND2X0 U13801 ( .IN1(n13277), .IN2(n13278), .QN(g23132) );
  NAND2X0 U13802 ( .IN1(n4456), .IN2(g2555), .QN(n13278) );
  NAND2X0 U13803 ( .IN1(n10288), .IN2(g8087), .QN(n13277) );
  NAND2X0 U13804 ( .IN1(n13279), .IN2(n13280), .QN(g23126) );
  NAND2X0 U13805 ( .IN1(n4465), .IN2(g1175), .QN(n13280) );
  NAND2X0 U13806 ( .IN1(n11379), .IN2(g1172), .QN(n13279) );
  NAND2X0 U13807 ( .IN1(n13281), .IN2(n13282), .QN(g23124) );
  NAND2X0 U13808 ( .IN1(n4457), .IN2(g1868), .QN(n13282) );
  NAND2X0 U13809 ( .IN1(n11359), .IN2(g8082), .QN(n13281) );
  NAND2X0 U13810 ( .IN1(n13283), .IN2(n13284), .QN(g23123) );
  NAND2X0 U13811 ( .IN1(n4458), .IN2(g1861), .QN(n13284) );
  NAND2X0 U13812 ( .IN1(n10305), .IN2(g8012), .QN(n13283) );
  NAND2X0 U13813 ( .IN1(n13285), .IN2(n13286), .QN(g23117) );
  NAND2X0 U13814 ( .IN1(n4466), .IN2(g488), .QN(n13286) );
  NAND2X0 U13815 ( .IN1(n11394), .IN2(g485), .QN(n13285) );
  NAND2X0 U13816 ( .IN1(n13287), .IN2(n13288), .QN(g23114) );
  NAND2X0 U13817 ( .IN1(n4456), .IN2(g2561), .QN(n13288) );
  NAND2X0 U13818 ( .IN1(n11339), .IN2(g8087), .QN(n13287) );
  NAND2X0 U13819 ( .IN1(n13289), .IN2(n13290), .QN(g23111) );
  NAND2X0 U13820 ( .IN1(test_so44), .IN2(n4459), .QN(n13290) );
  NAND2X0 U13821 ( .IN1(n11379), .IN2(g8007), .QN(n13289) );
  NAND2X0 U13822 ( .IN1(n13291), .IN2(n13292), .QN(g23110) );
  NAND2X0 U13823 ( .IN1(n4460), .IN2(g1167), .QN(n13292) );
  NAND2X0 U13824 ( .IN1(n10322), .IN2(g7961), .QN(n13291) );
  NAND2X0 U13825 ( .IN1(n13293), .IN2(n13294), .QN(g23097) );
  NAND2X0 U13826 ( .IN1(n4458), .IN2(g1867), .QN(n13294) );
  NAND2X0 U13827 ( .IN1(n11359), .IN2(g8012), .QN(n13293) );
  NAND3X0 U13828 ( .IN1(n13295), .IN2(n13296), .IN3(n13297), .QN(n11359) );
  NAND2X0 U13829 ( .IN1(g5511), .IN2(g1819), .QN(n13297) );
  NAND2X0 U13830 ( .IN1(test_so59), .IN2(n4618), .QN(n13296) );
  NAND2X0 U13831 ( .IN1(g7014), .IN2(g1822), .QN(n13295) );
  NAND2X0 U13832 ( .IN1(n13298), .IN2(n13299), .QN(g23093) );
  NAND2X0 U13833 ( .IN1(n4461), .IN2(g487), .QN(n13299) );
  NAND2X0 U13834 ( .IN1(n11394), .IN2(g7956), .QN(n13298) );
  NAND2X0 U13835 ( .IN1(n13300), .IN2(n13301), .QN(g23092) );
  NAND2X0 U13836 ( .IN1(g480), .IN2(n8072), .QN(n13301) );
  NAND2X0 U13837 ( .IN1(test_so23), .IN2(n10336), .QN(n13300) );
  NAND2X0 U13838 ( .IN1(n13302), .IN2(n13303), .QN(g23081) );
  NAND2X0 U13839 ( .IN1(n4460), .IN2(g1173), .QN(n13303) );
  NAND2X0 U13840 ( .IN1(n11379), .IN2(g7961), .QN(n13302) );
  NAND3X0 U13841 ( .IN1(n13304), .IN2(n13305), .IN3(n13306), .QN(n11379) );
  NAND2X0 U13842 ( .IN1(g1088), .IN2(g1131), .QN(n13306) );
  NAND2X0 U13843 ( .IN1(g5472), .IN2(g1125), .QN(n13305) );
  NAND2X0 U13844 ( .IN1(g6712), .IN2(g1128), .QN(n13304) );
  NAND2X0 U13845 ( .IN1(n13307), .IN2(n13308), .QN(g23076) );
  NAND2X0 U13846 ( .IN1(n4463), .IN2(g2539), .QN(n13308) );
  NAND2X0 U13847 ( .IN1(n10288), .IN2(g2560), .QN(n13307) );
  NAND2X0 U13848 ( .IN1(n13309), .IN2(n13310), .QN(g23067) );
  NAND2X0 U13849 ( .IN1(g486), .IN2(n8072), .QN(n13310) );
  NAND2X0 U13850 ( .IN1(test_so23), .IN2(n11394), .QN(n13309) );
  NAND3X0 U13851 ( .IN1(n13311), .IN2(n13312), .IN3(n13313), .QN(n11394) );
  NAND2X0 U13852 ( .IN1(g5437), .IN2(g438), .QN(n13313) );
  NAND2X0 U13853 ( .IN1(n4640), .IN2(g444), .QN(n13312) );
  NAND2X0 U13854 ( .IN1(g6447), .IN2(g441), .QN(n13311) );
  NAND2X0 U13855 ( .IN1(n13314), .IN2(n13315), .QN(g23058) );
  NAND2X0 U13856 ( .IN1(n4464), .IN2(g1845), .QN(n13315) );
  NAND2X0 U13857 ( .IN1(n10305), .IN2(g1866), .QN(n13314) );
  NAND2X0 U13858 ( .IN1(n13316), .IN2(n13317), .QN(g23047) );
  NAND2X0 U13859 ( .IN1(n4455), .IN2(g2559), .QN(n13317) );
  NAND2X0 U13860 ( .IN1(n10288), .IN2(g8167), .QN(n13316) );
  INVX0 U13861 ( .INP(n4285), .ZN(n10288) );
  NAND3X0 U13862 ( .IN1(n13318), .IN2(n13319), .IN3(n13320), .QN(n4285) );
  NAND2X0 U13863 ( .IN1(g5555), .IN2(g2492), .QN(n13320) );
  NAND2X0 U13864 ( .IN1(n4606), .IN2(g2498), .QN(n13319) );
  NAND2X0 U13865 ( .IN1(g7264), .IN2(g2495), .QN(n13318) );
  NAND2X0 U13866 ( .IN1(n13321), .IN2(n13322), .QN(g23039) );
  NAND2X0 U13867 ( .IN1(n4465), .IN2(g1151), .QN(n13322) );
  NAND2X0 U13868 ( .IN1(n10322), .IN2(g1172), .QN(n13321) );
  NAND2X0 U13869 ( .IN1(n13323), .IN2(n13324), .QN(g23030) );
  NAND2X0 U13870 ( .IN1(n4457), .IN2(g1865), .QN(n13324) );
  NAND2X0 U13871 ( .IN1(n10305), .IN2(g8082), .QN(n13323) );
  INVX0 U13872 ( .INP(n4284), .ZN(n10305) );
  NAND3X0 U13873 ( .IN1(n13325), .IN2(n13326), .IN3(n13327), .QN(n4284) );
  NAND2X0 U13874 ( .IN1(g5511), .IN2(g1798), .QN(n13327) );
  NAND2X0 U13875 ( .IN1(n4618), .IN2(g1804), .QN(n13326) );
  NAND2X0 U13876 ( .IN1(g7014), .IN2(g1801), .QN(n13325) );
  NAND2X0 U13877 ( .IN1(n13328), .IN2(n13329), .QN(g23022) );
  NAND2X0 U13878 ( .IN1(n4466), .IN2(g464), .QN(n13329) );
  NAND2X0 U13879 ( .IN1(n10336), .IN2(g485), .QN(n13328) );
  NAND2X0 U13880 ( .IN1(n13330), .IN2(n13331), .QN(g23014) );
  NAND2X0 U13881 ( .IN1(n4459), .IN2(g1171), .QN(n13331) );
  NAND2X0 U13882 ( .IN1(n10322), .IN2(g8007), .QN(n13330) );
  INVX0 U13883 ( .INP(n4283), .ZN(n10322) );
  NAND3X0 U13884 ( .IN1(n13332), .IN2(n13333), .IN3(n13334), .QN(n4283) );
  NAND2X0 U13885 ( .IN1(g1088), .IN2(g1110), .QN(n13334) );
  NAND2X0 U13886 ( .IN1(g5472), .IN2(g1104), .QN(n13333) );
  NAND2X0 U13887 ( .IN1(g6712), .IN2(g1107), .QN(n13332) );
  NAND2X0 U13888 ( .IN1(n13335), .IN2(n13336), .QN(g23000) );
  NAND2X0 U13889 ( .IN1(n4461), .IN2(g484), .QN(n13336) );
  NAND2X0 U13890 ( .IN1(n10336), .IN2(g7956), .QN(n13335) );
  INVX0 U13891 ( .INP(n4282), .ZN(n10336) );
  NAND3X0 U13892 ( .IN1(n13337), .IN2(n13338), .IN3(n13339), .QN(n4282) );
  NAND2X0 U13893 ( .IN1(g5437), .IN2(g417), .QN(n13339) );
  NAND2X0 U13894 ( .IN1(n4640), .IN2(g423), .QN(n13338) );
  NAND2X0 U13895 ( .IN1(g6447), .IN2(g420), .QN(n13337) );
  NAND2X0 U13896 ( .IN1(n13340), .IN2(n13341), .QN(g22687) );
  NAND3X0 U13897 ( .IN1(n8876), .IN2(g2584), .IN3(n13342), .QN(n13341) );
  INVX0 U13898 ( .INP(n12376), .ZN(n13342) );
  NAND2X0 U13899 ( .IN1(n13343), .IN2(n13344), .QN(n13340) );
  NAND2X0 U13900 ( .IN1(n8865), .IN2(n12376), .QN(n13343) );
  NAND3X0 U13901 ( .IN1(n13345), .IN2(n13346), .IN3(n13347), .QN(n12376) );
  NAND2X0 U13902 ( .IN1(g7390), .IN2(g2568), .QN(n13347) );
  NAND2X0 U13903 ( .IN1(g2624), .IN2(g2571), .QN(n13346) );
  NAND2X0 U13904 ( .IN1(n10166), .IN2(g2565), .QN(n13345) );
  NAND2X0 U13905 ( .IN1(n13348), .IN2(n13349), .QN(g22651) );
  NAND3X0 U13906 ( .IN1(n9002), .IN2(g1890), .IN3(n13350), .QN(n13349) );
  INVX0 U13907 ( .INP(n12384), .ZN(n13350) );
  NAND2X0 U13908 ( .IN1(n13351), .IN2(n13344), .QN(n13348) );
  NAND2X0 U13909 ( .IN1(n8980), .IN2(n12384), .QN(n13351) );
  NAND3X0 U13910 ( .IN1(n13352), .IN2(n13353), .IN3(n13354), .QN(n12384) );
  NAND2X0 U13911 ( .IN1(g1930), .IN2(g1877), .QN(n13354) );
  NAND2X0 U13912 ( .IN1(test_so68), .IN2(n10214), .QN(n13353) );
  NAND2X0 U13913 ( .IN1(g7194), .IN2(g1874), .QN(n13352) );
  NAND2X0 U13914 ( .IN1(n13355), .IN2(n13356), .QN(g22615) );
  NAND3X0 U13915 ( .IN1(n9108), .IN2(g1196), .IN3(n13357), .QN(n13356) );
  INVX0 U13916 ( .INP(n12392), .ZN(n13357) );
  NAND2X0 U13917 ( .IN1(n13358), .IN2(n13344), .QN(n13355) );
  NAND2X0 U13918 ( .IN1(n9097), .IN2(n12392), .QN(n13358) );
  NAND3X0 U13919 ( .IN1(n13359), .IN2(n13360), .IN3(n13361), .QN(n12392) );
  NAND2X0 U13920 ( .IN1(test_so47), .IN2(n11104), .QN(n13361) );
  NAND2X0 U13921 ( .IN1(g1236), .IN2(g1183), .QN(n13360) );
  NAND2X0 U13922 ( .IN1(g6944), .IN2(g1180), .QN(n13359) );
  NAND2X0 U13923 ( .IN1(n13362), .IN2(n13363), .QN(g22578) );
  NAND3X0 U13924 ( .IN1(test_so22), .IN2(n8751), .IN3(n13364), .QN(n13363) );
  INVX0 U13925 ( .INP(n12397), .ZN(n13364) );
  NAND2X0 U13926 ( .IN1(n13365), .IN2(n13344), .QN(n13362) );
  NAND2X0 U13927 ( .IN1(n8745), .IN2(n12397), .QN(n13365) );
  NAND3X0 U13928 ( .IN1(n13366), .IN2(n13367), .IN3(n13368), .QN(n12397) );
  NAND2X0 U13929 ( .IN1(g6642), .IN2(g493), .QN(n13368) );
  NAND2X0 U13930 ( .IN1(g6485), .IN2(g490), .QN(n13367) );
  NAND2X0 U13931 ( .IN1(g550), .IN2(g496), .QN(n13366) );
  NOR2X0 U13932 ( .IN1(n13369), .IN2(n13370), .QN(g22299) );
  NOR2X0 U13933 ( .IN1(n12592), .IN2(test_so95), .QN(n13370) );
  NOR2X0 U13934 ( .IN1(n11303), .IN2(n13371), .QN(g22284) );
  INVX0 U13935 ( .INP(n13372), .ZN(n13371) );
  NAND2X0 U13936 ( .IN1(n12595), .IN2(n7953), .QN(n13372) );
  NOR2X0 U13937 ( .IN1(n13373), .IN2(n13374), .QN(g22280) );
  NOR2X0 U13938 ( .IN1(n12601), .IN2(g2117), .QN(n13374) );
  NOR2X0 U13939 ( .IN1(n13375), .IN2(n13376), .QN(g22269) );
  INVX0 U13940 ( .INP(n13377), .ZN(n13376) );
  NAND2X0 U13941 ( .IN1(n12604), .IN2(n7865), .QN(n13377) );
  NOR2X0 U13942 ( .IN1(n13378), .IN2(n13379), .QN(g22263) );
  NOR2X0 U13943 ( .IN1(n12665), .IN2(g1423), .QN(n13379) );
  NOR2X0 U13944 ( .IN1(n13380), .IN2(n13381), .QN(g22249) );
  INVX0 U13945 ( .INP(n13382), .ZN(n13381) );
  NAND2X0 U13946 ( .IN1(n12669), .IN2(n7866), .QN(n13382) );
  NOR2X0 U13947 ( .IN1(n13383), .IN2(n13384), .QN(g22242) );
  NOR2X0 U13948 ( .IN1(n12731), .IN2(g737), .QN(n13384) );
  NOR2X0 U13949 ( .IN1(n13385), .IN2(n13386), .QN(g22234) );
  INVX0 U13950 ( .INP(n13387), .ZN(n13386) );
  NAND2X0 U13951 ( .IN1(n12737), .IN2(n7867), .QN(n13387) );
  NOR2X0 U13952 ( .IN1(n13388), .IN2(n13389), .QN(g22218) );
  INVX0 U13953 ( .INP(n13390), .ZN(n13389) );
  NAND2X0 U13954 ( .IN1(n12797), .IN2(n7868), .QN(n13390) );
  NAND2X0 U13955 ( .IN1(n13391), .IN2(n13392), .QN(g22200) );
  NAND2X0 U13956 ( .IN1(n13012), .IN2(n4373), .QN(n13392) );
  INVX0 U13957 ( .INP(n13393), .ZN(n13391) );
  NOR2X0 U13958 ( .IN1(n13012), .IN2(n7519), .QN(n13393) );
  NAND2X0 U13959 ( .IN1(n13394), .IN2(n13395), .QN(g22194) );
  INVX0 U13960 ( .INP(n13396), .ZN(n13395) );
  NOR2X0 U13961 ( .IN1(n13012), .IN2(n7511), .QN(n13396) );
  NAND2X0 U13962 ( .IN1(n13012), .IN2(n9454), .QN(n13394) );
  NAND2X0 U13963 ( .IN1(n13397), .IN2(n13398), .QN(g22193) );
  NAND2X0 U13964 ( .IN1(n13399), .IN2(n4373), .QN(n13398) );
  NAND2X0 U13965 ( .IN1(n13400), .IN2(g2210), .QN(n13397) );
  NAND2X0 U13966 ( .IN1(n13401), .IN2(n13402), .QN(g22192) );
  NAND2X0 U13967 ( .IN1(n13012), .IN2(n4377), .QN(n13402) );
  INVX0 U13968 ( .INP(n13403), .ZN(n13401) );
  NOR2X0 U13969 ( .IN1(n13012), .IN2(n7520), .QN(n13403) );
  NAND2X0 U13970 ( .IN1(n13404), .IN2(n13405), .QN(g22191) );
  NAND2X0 U13971 ( .IN1(n13015), .IN2(n4374), .QN(n13405) );
  INVX0 U13972 ( .INP(n13406), .ZN(n13404) );
  NOR2X0 U13973 ( .IN1(n13015), .IN2(n7530), .QN(n13406) );
  NAND2X0 U13974 ( .IN1(n13407), .IN2(n13408), .QN(g22185) );
  NAND2X0 U13975 ( .IN1(test_so75), .IN2(n13400), .QN(n13408) );
  NAND2X0 U13976 ( .IN1(n13399), .IN2(n9454), .QN(n13407) );
  NAND2X0 U13977 ( .IN1(n13409), .IN2(n13410), .QN(g22184) );
  INVX0 U13978 ( .INP(n13411), .ZN(n13410) );
  NOR2X0 U13979 ( .IN1(n13012), .IN2(n7502), .QN(n13411) );
  NAND2X0 U13980 ( .IN1(n10437), .IN2(n13012), .QN(n13409) );
  NAND2X0 U13981 ( .IN1(n13412), .IN2(n13413), .QN(g22183) );
  NAND2X0 U13982 ( .IN1(n13414), .IN2(n4373), .QN(n13413) );
  INVX0 U13983 ( .INP(n13415), .ZN(n13412) );
  NOR2X0 U13984 ( .IN1(n13414), .IN2(n7881), .QN(n13415) );
  NAND2X0 U13985 ( .IN1(n13416), .IN2(n13417), .QN(g22182) );
  NAND2X0 U13986 ( .IN1(n13399), .IN2(n4377), .QN(n13417) );
  NAND2X0 U13987 ( .IN1(n13400), .IN2(g2207), .QN(n13416) );
  NAND2X0 U13988 ( .IN1(n13418), .IN2(n13419), .QN(g22180) );
  INVX0 U13989 ( .INP(n13420), .ZN(n13419) );
  NOR2X0 U13990 ( .IN1(n13015), .IN2(n7521), .QN(n13420) );
  NAND2X0 U13991 ( .IN1(n13015), .IN2(n9484), .QN(n13418) );
  NAND2X0 U13992 ( .IN1(n13421), .IN2(n13422), .QN(g22179) );
  NAND2X0 U13993 ( .IN1(n13423), .IN2(n4374), .QN(n13422) );
  NAND2X0 U13994 ( .IN1(n13424), .IN2(g1516), .QN(n13421) );
  NAND2X0 U13995 ( .IN1(n13425), .IN2(n13426), .QN(g22178) );
  NAND2X0 U13996 ( .IN1(n13015), .IN2(n4378), .QN(n13426) );
  INVX0 U13997 ( .INP(n13427), .ZN(n13425) );
  NOR2X0 U13998 ( .IN1(n13015), .IN2(n7531), .QN(n13427) );
  NAND2X0 U13999 ( .IN1(n13428), .IN2(n13429), .QN(g22177) );
  NAND2X0 U14000 ( .IN1(n13018), .IN2(n4375), .QN(n13429) );
  INVX0 U14001 ( .INP(n13430), .ZN(n13428) );
  NOR2X0 U14002 ( .IN1(n13018), .IN2(n7544), .QN(n13430) );
  NAND2X0 U14003 ( .IN1(n13431), .IN2(n13432), .QN(g22173) );
  INVX0 U14004 ( .INP(n13433), .ZN(n13432) );
  NOR2X0 U14005 ( .IN1(n13414), .IN2(n7512), .QN(n13433) );
  NAND2X0 U14006 ( .IN1(n13414), .IN2(n9454), .QN(n13431) );
  INVX0 U14007 ( .INP(n10762), .ZN(n9454) );
  NAND3X0 U14008 ( .IN1(n13434), .IN2(n13435), .IN3(n13436), .QN(n10762) );
  NAND2X0 U14009 ( .IN1(n7574), .IN2(test_so73), .QN(n13436) );
  NAND2X0 U14010 ( .IN1(n7575), .IN2(g6837), .QN(n13435) );
  NAND2X0 U14011 ( .IN1(n7573), .IN2(g2241), .QN(n13434) );
  NAND2X0 U14012 ( .IN1(n13437), .IN2(n13438), .QN(g22172) );
  NAND2X0 U14013 ( .IN1(n13400), .IN2(g2237), .QN(n13438) );
  NAND2X0 U14014 ( .IN1(n10437), .IN2(n13399), .QN(n13437) );
  NAND2X0 U14015 ( .IN1(n13439), .IN2(n13440), .QN(g22171) );
  NAND2X0 U14016 ( .IN1(n13012), .IN2(n4287), .QN(n13440) );
  INVX0 U14017 ( .INP(n13441), .ZN(n13439) );
  NOR2X0 U14018 ( .IN1(n13012), .IN2(n7513), .QN(n13441) );
  NAND2X0 U14019 ( .IN1(n13442), .IN2(n13443), .QN(g22170) );
  NAND2X0 U14020 ( .IN1(n13414), .IN2(n4377), .QN(n13443) );
  INVX0 U14021 ( .INP(n13444), .ZN(n13442) );
  NOR2X0 U14022 ( .IN1(n13414), .IN2(n7883), .QN(n13444) );
  NAND2X0 U14023 ( .IN1(n13445), .IN2(n13446), .QN(g22169) );
  NAND2X0 U14024 ( .IN1(n13424), .IN2(g1546), .QN(n13446) );
  NAND2X0 U14025 ( .IN1(n13423), .IN2(n9484), .QN(n13445) );
  NAND2X0 U14026 ( .IN1(n13447), .IN2(n13448), .QN(g22168) );
  INVX0 U14027 ( .INP(n13449), .ZN(n13448) );
  NOR2X0 U14028 ( .IN1(n13015), .IN2(n7505), .QN(n13449) );
  NAND2X0 U14029 ( .IN1(n13450), .IN2(n13015), .QN(n13447) );
  NAND2X0 U14030 ( .IN1(n13451), .IN2(n13452), .QN(g22167) );
  INVX0 U14031 ( .INP(n13453), .ZN(n13452) );
  NOR2X0 U14032 ( .IN1(n8093), .IN2(n13454), .QN(n13453) );
  NAND2X0 U14033 ( .IN1(n13454), .IN2(n4374), .QN(n13451) );
  NAND2X0 U14034 ( .IN1(n13455), .IN2(n13456), .QN(g22166) );
  NAND2X0 U14035 ( .IN1(n13423), .IN2(n4378), .QN(n13456) );
  NAND2X0 U14036 ( .IN1(n13424), .IN2(g1513), .QN(n13455) );
  NAND2X0 U14037 ( .IN1(n13457), .IN2(n13458), .QN(g22164) );
  INVX0 U14038 ( .INP(n13459), .ZN(n13458) );
  NOR2X0 U14039 ( .IN1(n13018), .IN2(n7532), .QN(n13459) );
  NAND2X0 U14040 ( .IN1(n13018), .IN2(n9516), .QN(n13457) );
  NAND2X0 U14041 ( .IN1(n13460), .IN2(n13461), .QN(g22163) );
  NAND2X0 U14042 ( .IN1(n13462), .IN2(n4375), .QN(n13461) );
  INVX0 U14043 ( .INP(n13463), .ZN(n13460) );
  NOR2X0 U14044 ( .IN1(n13462), .IN2(n7911), .QN(n13463) );
  NAND2X0 U14045 ( .IN1(n13464), .IN2(n13465), .QN(g22162) );
  NAND2X0 U14046 ( .IN1(n4379), .IN2(n13018), .QN(n13465) );
  INVX0 U14047 ( .INP(n13466), .ZN(n13464) );
  NOR2X0 U14048 ( .IN1(n13018), .IN2(n7545), .QN(n13466) );
  NAND2X0 U14049 ( .IN1(n13467), .IN2(n13468), .QN(g22161) );
  NAND2X0 U14050 ( .IN1(n13469), .IN2(n4376), .QN(n13468) );
  NAND2X0 U14051 ( .IN1(n13020), .IN2(g132), .QN(n13467) );
  NAND2X0 U14052 ( .IN1(n13470), .IN2(n13471), .QN(g22155) );
  INVX0 U14053 ( .INP(n13472), .ZN(n13471) );
  NOR2X0 U14054 ( .IN1(n13414), .IN2(n7504), .QN(n13472) );
  NAND2X0 U14055 ( .IN1(n13414), .IN2(n10437), .QN(n13470) );
  INVX0 U14056 ( .INP(n9601), .ZN(n10437) );
  NAND3X0 U14057 ( .IN1(n13473), .IN2(n13474), .IN3(n13475), .QN(n9601) );
  NAND2X0 U14058 ( .IN1(n7571), .IN2(test_so73), .QN(n13475) );
  NAND2X0 U14059 ( .IN1(n7572), .IN2(g6837), .QN(n13474) );
  NAND2X0 U14060 ( .IN1(n7570), .IN2(g2241), .QN(n13473) );
  NAND2X0 U14061 ( .IN1(n13476), .IN2(n13477), .QN(g22154) );
  NAND2X0 U14062 ( .IN1(n13399), .IN2(n4287), .QN(n13477) );
  NAND2X0 U14063 ( .IN1(n13400), .IN2(g2234), .QN(n13476) );
  NAND2X0 U14064 ( .IN1(n13478), .IN2(n13479), .QN(g22153) );
  NAND2X0 U14065 ( .IN1(n13012), .IN2(n4563), .QN(n13479) );
  INVX0 U14066 ( .INP(n13480), .ZN(n13478) );
  NOR2X0 U14067 ( .IN1(n13012), .IN2(n7514), .QN(n13480) );
  NAND2X0 U14068 ( .IN1(n13481), .IN2(n13482), .QN(g22152) );
  INVX0 U14069 ( .INP(n13483), .ZN(n13482) );
  NOR2X0 U14070 ( .IN1(n13454), .IN2(n7523), .QN(n13483) );
  NAND2X0 U14071 ( .IN1(n13454), .IN2(n9484), .QN(n13481) );
  INVX0 U14072 ( .INP(n10499), .ZN(n9484) );
  NAND3X0 U14073 ( .IN1(n13484), .IN2(n13485), .IN3(n13486), .QN(n10499) );
  NAND2X0 U14074 ( .IN1(n7585), .IN2(g6782), .QN(n13486) );
  NAND2X0 U14075 ( .IN1(n7586), .IN2(g6573), .QN(n13485) );
  NAND2X0 U14076 ( .IN1(g1547), .IN2(n8129), .QN(n13484) );
  NAND2X0 U14077 ( .IN1(n13487), .IN2(n13488), .QN(g22151) );
  NAND2X0 U14078 ( .IN1(n13424), .IN2(g1543), .QN(n13488) );
  NAND2X0 U14079 ( .IN1(n13450), .IN2(n13423), .QN(n13487) );
  NAND2X0 U14080 ( .IN1(n13489), .IN2(n13490), .QN(g22150) );
  NAND2X0 U14081 ( .IN1(n13015), .IN2(n4288), .QN(n13490) );
  INVX0 U14082 ( .INP(n13491), .ZN(n13489) );
  NOR2X0 U14083 ( .IN1(n13015), .IN2(n7524), .QN(n13491) );
  NAND2X0 U14084 ( .IN1(n13492), .IN2(n13493), .QN(g22149) );
  NAND2X0 U14085 ( .IN1(n13454), .IN2(n4378), .QN(n13493) );
  INVX0 U14086 ( .INP(n13494), .ZN(n13492) );
  NOR2X0 U14087 ( .IN1(n13454), .IN2(n7897), .QN(n13494) );
  NAND2X0 U14088 ( .IN1(n13495), .IN2(n13496), .QN(g22148) );
  INVX0 U14089 ( .INP(n13497), .ZN(n13496) );
  NOR2X0 U14090 ( .IN1(n13462), .IN2(n7533), .QN(n13497) );
  NAND2X0 U14091 ( .IN1(n13462), .IN2(n9516), .QN(n13495) );
  NAND2X0 U14092 ( .IN1(n13498), .IN2(n13499), .QN(g22147) );
  INVX0 U14093 ( .INP(n13500), .ZN(n13499) );
  NOR2X0 U14094 ( .IN1(n13018), .IN2(n7535), .QN(n13500) );
  NAND2X0 U14095 ( .IN1(n10618), .IN2(n13018), .QN(n13498) );
  NAND2X0 U14096 ( .IN1(n13501), .IN2(n13502), .QN(g22146) );
  NAND2X0 U14097 ( .IN1(n13503), .IN2(n4375), .QN(n13502) );
  NAND2X0 U14098 ( .IN1(n13504), .IN2(g821), .QN(n13501) );
  NAND2X0 U14099 ( .IN1(n13505), .IN2(n13506), .QN(g22145) );
  NAND2X0 U14100 ( .IN1(n13462), .IN2(n4379), .QN(n13506) );
  INVX0 U14101 ( .INP(n13507), .ZN(n13505) );
  NOR2X0 U14102 ( .IN1(n13462), .IN2(n7915), .QN(n13507) );
  NAND2X0 U14103 ( .IN1(n13508), .IN2(n13509), .QN(g22143) );
  NAND2X0 U14104 ( .IN1(n13020), .IN2(g162), .QN(n13509) );
  NAND2X0 U14105 ( .IN1(n13469), .IN2(n9560), .QN(n13508) );
  NAND2X0 U14106 ( .IN1(n13510), .IN2(n13511), .QN(g22142) );
  NAND2X0 U14107 ( .IN1(n13512), .IN2(n4376), .QN(n13511) );
  INVX0 U14108 ( .INP(n13513), .ZN(n13510) );
  NOR2X0 U14109 ( .IN1(n13512), .IN2(n7949), .QN(n13513) );
  NAND2X0 U14110 ( .IN1(n13514), .IN2(n13515), .QN(g22141) );
  NAND2X0 U14111 ( .IN1(n4380), .IN2(n13469), .QN(n13515) );
  NAND2X0 U14112 ( .IN1(n13020), .IN2(g129), .QN(n13514) );
  NAND2X0 U14113 ( .IN1(n13516), .IN2(n13517), .QN(g22140) );
  NAND2X0 U14114 ( .IN1(n13414), .IN2(n4287), .QN(n13517) );
  INVX0 U14115 ( .INP(n13518), .ZN(n13516) );
  NOR2X0 U14116 ( .IN1(n13414), .IN2(n7870), .QN(n13518) );
  NAND2X0 U14117 ( .IN1(n13519), .IN2(n13520), .QN(g22139) );
  NAND2X0 U14118 ( .IN1(n13399), .IN2(n4563), .QN(n13520) );
  NAND2X0 U14119 ( .IN1(n13400), .IN2(g2231), .QN(n13519) );
  NAND2X0 U14120 ( .IN1(n13521), .IN2(n13522), .QN(g22138) );
  NAND2X0 U14121 ( .IN1(n13012), .IN2(n4555), .QN(n13522) );
  INVX0 U14122 ( .INP(n13523), .ZN(n13521) );
  NOR2X0 U14123 ( .IN1(n13012), .IN2(n7515), .QN(n13523) );
  NAND2X0 U14124 ( .IN1(n13524), .IN2(n13525), .QN(g22132) );
  INVX0 U14125 ( .INP(n13526), .ZN(n13525) );
  NOR2X0 U14126 ( .IN1(n13454), .IN2(n7507), .QN(n13526) );
  NAND2X0 U14127 ( .IN1(n13454), .IN2(n13450), .QN(n13524) );
  INVX0 U14128 ( .INP(n9639), .ZN(n13450) );
  NAND3X0 U14129 ( .IN1(n13527), .IN2(n13528), .IN3(n13529), .QN(n9639) );
  NAND2X0 U14130 ( .IN1(n7583), .IN2(g6782), .QN(n13529) );
  NAND2X0 U14131 ( .IN1(n7584), .IN2(g6573), .QN(n13528) );
  NAND2X0 U14132 ( .IN1(n7582), .IN2(g1547), .QN(n13527) );
  NAND2X0 U14133 ( .IN1(n13530), .IN2(n13531), .QN(g22131) );
  NAND2X0 U14134 ( .IN1(n13423), .IN2(n4288), .QN(n13531) );
  NAND2X0 U14135 ( .IN1(n13424), .IN2(g1540), .QN(n13530) );
  NAND2X0 U14136 ( .IN1(n13532), .IN2(n13533), .QN(g22130) );
  NAND2X0 U14137 ( .IN1(n13015), .IN2(n4565), .QN(n13533) );
  INVX0 U14138 ( .INP(n13534), .ZN(n13532) );
  NOR2X0 U14139 ( .IN1(n13015), .IN2(n7525), .QN(n13534) );
  NAND2X0 U14140 ( .IN1(n13535), .IN2(n13536), .QN(g22129) );
  NAND2X0 U14141 ( .IN1(n13504), .IN2(g851), .QN(n13536) );
  NAND2X0 U14142 ( .IN1(n13503), .IN2(n9516), .QN(n13535) );
  INVX0 U14143 ( .INP(n10834), .ZN(n9516) );
  NAND3X0 U14144 ( .IN1(n13537), .IN2(n13538), .IN3(n13539), .QN(n10834) );
  NAND2X0 U14145 ( .IN1(n7596), .IN2(test_so31), .QN(n13539) );
  NAND2X0 U14146 ( .IN1(n7597), .IN2(g6518), .QN(n13538) );
  NAND2X0 U14147 ( .IN1(n7598), .IN2(g6368), .QN(n13537) );
  NAND2X0 U14148 ( .IN1(n13540), .IN2(n13541), .QN(g22128) );
  INVX0 U14149 ( .INP(n13542), .ZN(n13541) );
  NOR2X0 U14150 ( .IN1(n13462), .IN2(n7536), .QN(n13542) );
  NAND2X0 U14151 ( .IN1(n10618), .IN2(n13462), .QN(n13540) );
  NAND2X0 U14152 ( .IN1(n13543), .IN2(n13544), .QN(g22127) );
  NAND2X0 U14153 ( .IN1(n4289), .IN2(n13018), .QN(n13544) );
  INVX0 U14154 ( .INP(n13545), .ZN(n13543) );
  NOR2X0 U14155 ( .IN1(n13018), .IN2(n7538), .QN(n13545) );
  NAND2X0 U14156 ( .IN1(n13546), .IN2(n13547), .QN(g22126) );
  NAND2X0 U14157 ( .IN1(n13503), .IN2(n4379), .QN(n13547) );
  NAND2X0 U14158 ( .IN1(n13504), .IN2(g818), .QN(n13546) );
  NAND2X0 U14159 ( .IN1(n13548), .IN2(n13549), .QN(g22125) );
  INVX0 U14160 ( .INP(n13550), .ZN(n13549) );
  NOR2X0 U14161 ( .IN1(n13512), .IN2(n7547), .QN(n13550) );
  NAND2X0 U14162 ( .IN1(n13512), .IN2(n9560), .QN(n13548) );
  NAND2X0 U14163 ( .IN1(n13551), .IN2(n13552), .QN(g22124) );
  NAND2X0 U14164 ( .IN1(n13020), .IN2(g159), .QN(n13552) );
  NAND2X0 U14165 ( .IN1(n12339), .IN2(n13469), .QN(n13551) );
  NAND2X0 U14166 ( .IN1(n13553), .IN2(n13554), .QN(g22123) );
  NAND2X0 U14167 ( .IN1(n13555), .IN2(n4376), .QN(n13554) );
  NAND2X0 U14168 ( .IN1(n13556), .IN2(g133), .QN(n13553) );
  NAND2X0 U14169 ( .IN1(n13557), .IN2(n13558), .QN(g22122) );
  NAND2X0 U14170 ( .IN1(n13512), .IN2(n4380), .QN(n13558) );
  INVX0 U14171 ( .INP(n13559), .ZN(n13557) );
  NOR2X0 U14172 ( .IN1(n13512), .IN2(n7951), .QN(n13559) );
  NAND2X0 U14173 ( .IN1(n13560), .IN2(n13561), .QN(g22117) );
  NAND2X0 U14174 ( .IN1(n13414), .IN2(n4563), .QN(n13561) );
  INVX0 U14175 ( .INP(n13562), .ZN(n13560) );
  NOR2X0 U14176 ( .IN1(n13414), .IN2(n7872), .QN(n13562) );
  NAND2X0 U14177 ( .IN1(n13563), .IN2(n13564), .QN(g22116) );
  NAND2X0 U14178 ( .IN1(n13399), .IN2(n4555), .QN(n13564) );
  NAND2X0 U14179 ( .IN1(n13400), .IN2(g2228), .QN(n13563) );
  NAND2X0 U14180 ( .IN1(n13565), .IN2(n13566), .QN(g22115) );
  NAND2X0 U14181 ( .IN1(n13012), .IN2(n4325), .QN(n13566) );
  INVX0 U14182 ( .INP(n13567), .ZN(n13565) );
  NOR2X0 U14183 ( .IN1(n13012), .IN2(n7516), .QN(n13567) );
  NAND2X0 U14184 ( .IN1(n13568), .IN2(n13569), .QN(g22114) );
  NAND2X0 U14185 ( .IN1(n13454), .IN2(n4288), .QN(n13569) );
  INVX0 U14186 ( .INP(n13570), .ZN(n13568) );
  NOR2X0 U14187 ( .IN1(n13454), .IN2(n7885), .QN(n13570) );
  NAND2X0 U14188 ( .IN1(n13571), .IN2(n13572), .QN(g22113) );
  NAND2X0 U14189 ( .IN1(test_so53), .IN2(n13424), .QN(n13572) );
  NAND2X0 U14190 ( .IN1(n13423), .IN2(n4565), .QN(n13571) );
  NAND2X0 U14191 ( .IN1(n13573), .IN2(n13574), .QN(g22112) );
  NAND2X0 U14192 ( .IN1(n13015), .IN2(n4557), .QN(n13574) );
  INVX0 U14193 ( .INP(n13575), .ZN(n13573) );
  NOR2X0 U14194 ( .IN1(n13015), .IN2(n7526), .QN(n13575) );
  NAND2X0 U14195 ( .IN1(n13576), .IN2(n13577), .QN(g22106) );
  NAND2X0 U14196 ( .IN1(n13504), .IN2(g848), .QN(n13577) );
  NAND2X0 U14197 ( .IN1(n13503), .IN2(n10618), .QN(n13576) );
  INVX0 U14198 ( .INP(n9668), .ZN(n10618) );
  NAND3X0 U14199 ( .IN1(n13578), .IN2(n13579), .IN3(n13580), .QN(n9668) );
  NAND2X0 U14200 ( .IN1(n7593), .IN2(test_so31), .QN(n13580) );
  NAND2X0 U14201 ( .IN1(n7594), .IN2(g6518), .QN(n13579) );
  NAND2X0 U14202 ( .IN1(n7595), .IN2(g6368), .QN(n13578) );
  NAND2X0 U14203 ( .IN1(n13581), .IN2(n13582), .QN(g22105) );
  NAND2X0 U14204 ( .IN1(n4289), .IN2(n13462), .QN(n13582) );
  INVX0 U14205 ( .INP(n13583), .ZN(n13581) );
  NOR2X0 U14206 ( .IN1(n13462), .IN2(n7898), .QN(n13583) );
  NAND2X0 U14207 ( .IN1(n13584), .IN2(n13585), .QN(g22104) );
  NAND2X0 U14208 ( .IN1(n13018), .IN2(n4567), .QN(n13585) );
  INVX0 U14209 ( .INP(n13586), .ZN(n13584) );
  NOR2X0 U14210 ( .IN1(n13018), .IN2(n7539), .QN(n13586) );
  NAND2X0 U14211 ( .IN1(n13587), .IN2(n13588), .QN(g22103) );
  NAND2X0 U14212 ( .IN1(test_so12), .IN2(n13556), .QN(n13588) );
  NAND2X0 U14213 ( .IN1(n13555), .IN2(n9560), .QN(n13587) );
  INVX0 U14214 ( .INP(n10704), .ZN(n9560) );
  NAND3X0 U14215 ( .IN1(n13589), .IN2(n13590), .IN3(n13591), .QN(n10704) );
  NAND2X0 U14216 ( .IN1(n7608), .IN2(g6313), .QN(n13591) );
  NAND2X0 U14217 ( .IN1(n7609), .IN2(g6231), .QN(n13590) );
  NAND2X0 U14218 ( .IN1(n7607), .IN2(g165), .QN(n13589) );
  NAND2X0 U14219 ( .IN1(n13592), .IN2(n13593), .QN(g22102) );
  INVX0 U14220 ( .INP(n13594), .ZN(n13593) );
  NOR2X0 U14221 ( .IN1(n13512), .IN2(n7509), .QN(n13594) );
  NAND2X0 U14222 ( .IN1(n12339), .IN2(n13512), .QN(n13592) );
  NAND2X0 U14223 ( .IN1(n13595), .IN2(n13596), .QN(g22101) );
  NAND2X0 U14224 ( .IN1(n4290), .IN2(n13469), .QN(n13596) );
  NAND2X0 U14225 ( .IN1(n13020), .IN2(g156), .QN(n13595) );
  NAND2X0 U14226 ( .IN1(n13597), .IN2(n13598), .QN(g22100) );
  NAND2X0 U14227 ( .IN1(n13555), .IN2(n4380), .QN(n13598) );
  NAND2X0 U14228 ( .IN1(n13556), .IN2(g130), .QN(n13597) );
  NAND2X0 U14229 ( .IN1(n13599), .IN2(n13600), .QN(g22099) );
  NAND2X0 U14230 ( .IN1(n13414), .IN2(n4555), .QN(n13600) );
  INVX0 U14231 ( .INP(n13601), .ZN(n13599) );
  NOR2X0 U14232 ( .IN1(n13414), .IN2(n7874), .QN(n13601) );
  NAND2X0 U14233 ( .IN1(n13602), .IN2(n13603), .QN(g22098) );
  NAND2X0 U14234 ( .IN1(test_so74), .IN2(n13400), .QN(n13603) );
  NAND2X0 U14235 ( .IN1(n13399), .IN2(n4325), .QN(n13602) );
  NAND2X0 U14236 ( .IN1(n13604), .IN2(n13605), .QN(g22097) );
  NAND2X0 U14237 ( .IN1(n13012), .IN2(n4389), .QN(n13605) );
  INVX0 U14238 ( .INP(n13606), .ZN(n13604) );
  NOR2X0 U14239 ( .IN1(n13012), .IN2(n7517), .QN(n13606) );
  NAND2X0 U14240 ( .IN1(n13607), .IN2(n13608), .QN(g22092) );
  NAND2X0 U14241 ( .IN1(n13454), .IN2(n4565), .QN(n13608) );
  INVX0 U14242 ( .INP(n13609), .ZN(n13607) );
  NOR2X0 U14243 ( .IN1(n13454), .IN2(n7886), .QN(n13609) );
  NAND2X0 U14244 ( .IN1(n13610), .IN2(n13611), .QN(g22091) );
  NAND2X0 U14245 ( .IN1(n13423), .IN2(n4557), .QN(n13611) );
  NAND2X0 U14246 ( .IN1(n13424), .IN2(g1534), .QN(n13610) );
  NAND2X0 U14247 ( .IN1(n13612), .IN2(n13613), .QN(g22090) );
  NAND2X0 U14248 ( .IN1(n13015), .IN2(n4326), .QN(n13613) );
  INVX0 U14249 ( .INP(n13614), .ZN(n13612) );
  NOR2X0 U14250 ( .IN1(n13015), .IN2(n7527), .QN(n13614) );
  NAND2X0 U14251 ( .IN1(n13615), .IN2(n13616), .QN(g22089) );
  NAND2X0 U14252 ( .IN1(n4289), .IN2(n13503), .QN(n13616) );
  NAND2X0 U14253 ( .IN1(n13504), .IN2(g845), .QN(n13615) );
  NAND2X0 U14254 ( .IN1(n13617), .IN2(n13618), .QN(g22088) );
  NAND2X0 U14255 ( .IN1(n13462), .IN2(n4567), .QN(n13618) );
  INVX0 U14256 ( .INP(n13619), .ZN(n13617) );
  NOR2X0 U14257 ( .IN1(n13462), .IN2(n7900), .QN(n13619) );
  NAND2X0 U14258 ( .IN1(n13620), .IN2(n13621), .QN(g22087) );
  NAND2X0 U14259 ( .IN1(n13018), .IN2(n4559), .QN(n13621) );
  INVX0 U14260 ( .INP(n13622), .ZN(n13620) );
  NOR2X0 U14261 ( .IN1(n13018), .IN2(n7540), .QN(n13622) );
  NAND2X0 U14262 ( .IN1(n13623), .IN2(n13624), .QN(g22081) );
  NAND2X0 U14263 ( .IN1(n13556), .IN2(g160), .QN(n13624) );
  NAND2X0 U14264 ( .IN1(n13555), .IN2(n12339), .QN(n13623) );
  INVX0 U14265 ( .INP(n9689), .ZN(n12339) );
  NAND3X0 U14266 ( .IN1(n13625), .IN2(n13626), .IN3(n13627), .QN(n9689) );
  NAND2X0 U14267 ( .IN1(n7605), .IN2(g6313), .QN(n13627) );
  NAND2X0 U14268 ( .IN1(n7606), .IN2(g6231), .QN(n13626) );
  NAND2X0 U14269 ( .IN1(n7604), .IN2(g165), .QN(n13625) );
  NAND2X0 U14270 ( .IN1(n13628), .IN2(n13629), .QN(g22080) );
  NAND2X0 U14271 ( .IN1(n4290), .IN2(n13512), .QN(n13629) );
  INVX0 U14272 ( .INP(n13630), .ZN(n13628) );
  NOR2X0 U14273 ( .IN1(n13512), .IN2(n7917), .QN(n13630) );
  NAND2X0 U14274 ( .IN1(n13631), .IN2(n13632), .QN(g22079) );
  NAND2X0 U14275 ( .IN1(n13469), .IN2(n4569), .QN(n13632) );
  NAND2X0 U14276 ( .IN1(n13020), .IN2(g153), .QN(n13631) );
  NAND2X0 U14277 ( .IN1(n13633), .IN2(n13634), .QN(g22078) );
  NAND2X0 U14278 ( .IN1(n13414), .IN2(n4325), .QN(n13634) );
  INVX0 U14279 ( .INP(n13635), .ZN(n13633) );
  NOR2X0 U14280 ( .IN1(n13414), .IN2(n7875), .QN(n13635) );
  NAND2X0 U14281 ( .IN1(n13636), .IN2(n13637), .QN(g22077) );
  NAND2X0 U14282 ( .IN1(n13399), .IN2(n4389), .QN(n13637) );
  NAND2X0 U14283 ( .IN1(n13400), .IN2(g2222), .QN(n13636) );
  NAND2X0 U14284 ( .IN1(n13638), .IN2(n13639), .QN(g22076) );
  NAND2X0 U14285 ( .IN1(n13012), .IN2(n4319), .QN(n13639) );
  INVX0 U14286 ( .INP(n13640), .ZN(n13638) );
  NOR2X0 U14287 ( .IN1(n13012), .IN2(n7518), .QN(n13640) );
  NOR2X0 U14288 ( .IN1(n4367), .IN2(n7706), .QN(n13012) );
  NAND2X0 U14289 ( .IN1(n13641), .IN2(n13642), .QN(g22075) );
  NAND2X0 U14290 ( .IN1(n13454), .IN2(n4557), .QN(n13642) );
  INVX0 U14291 ( .INP(n13643), .ZN(n13641) );
  NOR2X0 U14292 ( .IN1(n13454), .IN2(n7888), .QN(n13643) );
  NAND2X0 U14293 ( .IN1(n13644), .IN2(n13645), .QN(g22074) );
  NAND2X0 U14294 ( .IN1(n13423), .IN2(n4326), .QN(n13645) );
  NAND2X0 U14295 ( .IN1(n13424), .IN2(g1531), .QN(n13644) );
  NAND2X0 U14296 ( .IN1(n13646), .IN2(n13647), .QN(g22073) );
  NAND2X0 U14297 ( .IN1(n13015), .IN2(n4390), .QN(n13647) );
  INVX0 U14298 ( .INP(n13648), .ZN(n13646) );
  NOR2X0 U14299 ( .IN1(n13015), .IN2(n7528), .QN(n13648) );
  NAND2X0 U14300 ( .IN1(n13649), .IN2(n13650), .QN(g22068) );
  NAND2X0 U14301 ( .IN1(n13503), .IN2(n4567), .QN(n13650) );
  NAND2X0 U14302 ( .IN1(n13504), .IN2(g842), .QN(n13649) );
  NAND2X0 U14303 ( .IN1(n13651), .IN2(n13652), .QN(g22067) );
  NAND2X0 U14304 ( .IN1(n13462), .IN2(n4559), .QN(n13652) );
  INVX0 U14305 ( .INP(n13653), .ZN(n13651) );
  NOR2X0 U14306 ( .IN1(n13462), .IN2(n7902), .QN(n13653) );
  NAND2X0 U14307 ( .IN1(n13654), .IN2(n13655), .QN(g22066) );
  NAND2X0 U14308 ( .IN1(n4327), .IN2(n13018), .QN(n13655) );
  INVX0 U14309 ( .INP(n13656), .ZN(n13654) );
  NOR2X0 U14310 ( .IN1(n13018), .IN2(n7541), .QN(n13656) );
  NAND2X0 U14311 ( .IN1(n13657), .IN2(n13658), .QN(g22065) );
  NAND2X0 U14312 ( .IN1(n4290), .IN2(n13555), .QN(n13658) );
  NAND2X0 U14313 ( .IN1(n13556), .IN2(g157), .QN(n13657) );
  NAND2X0 U14314 ( .IN1(n13659), .IN2(n13660), .QN(g22064) );
  NAND2X0 U14315 ( .IN1(n13512), .IN2(n4569), .QN(n13660) );
  INVX0 U14316 ( .INP(n13661), .ZN(n13659) );
  NOR2X0 U14317 ( .IN1(n13512), .IN2(n7927), .QN(n13661) );
  NAND2X0 U14318 ( .IN1(n13662), .IN2(n13663), .QN(g22063) );
  NAND2X0 U14319 ( .IN1(n13469), .IN2(n4561), .QN(n13663) );
  NAND2X0 U14320 ( .IN1(n13020), .IN2(g150), .QN(n13662) );
  NAND2X0 U14321 ( .IN1(n13664), .IN2(n13665), .QN(g22061) );
  NAND2X0 U14322 ( .IN1(n13414), .IN2(n4389), .QN(n13665) );
  INVX0 U14323 ( .INP(n13666), .ZN(n13664) );
  NOR2X0 U14324 ( .IN1(n13414), .IN2(n7877), .QN(n13666) );
  NAND2X0 U14325 ( .IN1(n13667), .IN2(n13668), .QN(g22060) );
  NAND2X0 U14326 ( .IN1(n13399), .IN2(n4319), .QN(n13668) );
  NAND2X0 U14327 ( .IN1(n13400), .IN2(g2219), .QN(n13667) );
  INVX0 U14328 ( .INP(n13399), .ZN(n13400) );
  NOR2X0 U14329 ( .IN1(n8070), .IN2(n7706), .QN(n13399) );
  NAND2X0 U14330 ( .IN1(n13669), .IN2(n13670), .QN(g22059) );
  NAND2X0 U14331 ( .IN1(n13454), .IN2(n4326), .QN(n13670) );
  INVX0 U14332 ( .INP(n13671), .ZN(n13669) );
  NOR2X0 U14333 ( .IN1(n13454), .IN2(n7890), .QN(n13671) );
  NAND2X0 U14334 ( .IN1(n13672), .IN2(n13673), .QN(g22058) );
  NAND2X0 U14335 ( .IN1(n13423), .IN2(n4390), .QN(n13673) );
  NAND2X0 U14336 ( .IN1(n13424), .IN2(g1528), .QN(n13672) );
  NAND2X0 U14337 ( .IN1(n13674), .IN2(n13675), .QN(g22057) );
  NAND2X0 U14338 ( .IN1(n13015), .IN2(n4320), .QN(n13675) );
  INVX0 U14339 ( .INP(n13676), .ZN(n13674) );
  NOR2X0 U14340 ( .IN1(n13015), .IN2(n7529), .QN(n13676) );
  NOR2X0 U14341 ( .IN1(n4368), .IN2(n7707), .QN(n13015) );
  NAND2X0 U14342 ( .IN1(n13677), .IN2(n13678), .QN(g22056) );
  NAND2X0 U14343 ( .IN1(test_so32), .IN2(n13504), .QN(n13678) );
  NAND2X0 U14344 ( .IN1(n13503), .IN2(n4559), .QN(n13677) );
  NAND2X0 U14345 ( .IN1(n13679), .IN2(n13680), .QN(g22055) );
  NAND2X0 U14346 ( .IN1(n4327), .IN2(n13462), .QN(n13680) );
  INVX0 U14347 ( .INP(n13681), .ZN(n13679) );
  NOR2X0 U14348 ( .IN1(n13462), .IN2(n7903), .QN(n13681) );
  NAND2X0 U14349 ( .IN1(n13682), .IN2(n13683), .QN(g22054) );
  NAND2X0 U14350 ( .IN1(n13018), .IN2(n4391), .QN(n13683) );
  INVX0 U14351 ( .INP(n13684), .ZN(n13682) );
  NOR2X0 U14352 ( .IN1(n13018), .IN2(n7542), .QN(n13684) );
  NAND2X0 U14353 ( .IN1(n13685), .IN2(n13686), .QN(g22049) );
  NAND2X0 U14354 ( .IN1(n13555), .IN2(n4569), .QN(n13686) );
  NAND2X0 U14355 ( .IN1(n13556), .IN2(g154), .QN(n13685) );
  NAND2X0 U14356 ( .IN1(n13687), .IN2(n13688), .QN(g22048) );
  NAND2X0 U14357 ( .IN1(n13512), .IN2(n4561), .QN(n13688) );
  INVX0 U14358 ( .INP(n13689), .ZN(n13687) );
  NOR2X0 U14359 ( .IN1(n13512), .IN2(n7931), .QN(n13689) );
  NAND2X0 U14360 ( .IN1(n13690), .IN2(n13691), .QN(g22047) );
  NAND2X0 U14361 ( .IN1(n4328), .IN2(n13469), .QN(n13691) );
  NAND2X0 U14362 ( .IN1(n13020), .IN2(g147), .QN(n13690) );
  NAND2X0 U14363 ( .IN1(n13692), .IN2(n13693), .QN(g22045) );
  NAND2X0 U14364 ( .IN1(n13414), .IN2(n4319), .QN(n13693) );
  INVX0 U14365 ( .INP(n13694), .ZN(n13692) );
  NOR2X0 U14366 ( .IN1(n13414), .IN2(n7879), .QN(n13694) );
  NOR2X0 U14367 ( .IN1(n4324), .IN2(n7706), .QN(n13414) );
  NAND2X0 U14368 ( .IN1(n13695), .IN2(n13696), .QN(g22044) );
  NAND2X0 U14369 ( .IN1(n13454), .IN2(n4390), .QN(n13696) );
  INVX0 U14370 ( .INP(n13697), .ZN(n13695) );
  NOR2X0 U14371 ( .IN1(n13454), .IN2(n7892), .QN(n13697) );
  NAND2X0 U14372 ( .IN1(n13698), .IN2(n13699), .QN(g22043) );
  NAND2X0 U14373 ( .IN1(n13423), .IN2(n4320), .QN(n13699) );
  NAND2X0 U14374 ( .IN1(n13424), .IN2(g1525), .QN(n13698) );
  INVX0 U14375 ( .INP(n13423), .ZN(n13424) );
  NOR2X0 U14376 ( .IN1(n4515), .IN2(n7707), .QN(n13423) );
  NAND2X0 U14377 ( .IN1(n13700), .IN2(n13701), .QN(g22042) );
  NAND2X0 U14378 ( .IN1(n4327), .IN2(n13503), .QN(n13701) );
  NAND2X0 U14379 ( .IN1(n13504), .IN2(g836), .QN(n13700) );
  NAND2X0 U14380 ( .IN1(n13702), .IN2(n13703), .QN(g22041) );
  NAND2X0 U14381 ( .IN1(n13462), .IN2(n4391), .QN(n13703) );
  INVX0 U14382 ( .INP(n13704), .ZN(n13702) );
  NOR2X0 U14383 ( .IN1(n13462), .IN2(n7905), .QN(n13704) );
  NAND2X0 U14384 ( .IN1(n13705), .IN2(n13706), .QN(g22040) );
  NAND2X0 U14385 ( .IN1(n4321), .IN2(n13018), .QN(n13706) );
  INVX0 U14386 ( .INP(n13707), .ZN(n13705) );
  NOR2X0 U14387 ( .IN1(n13018), .IN2(n7543), .QN(n13707) );
  NOR2X0 U14388 ( .IN1(n8071), .IN2(n7708), .QN(n13018) );
  NAND2X0 U14389 ( .IN1(n13708), .IN2(n13709), .QN(g22039) );
  NAND2X0 U14390 ( .IN1(n13555), .IN2(n4561), .QN(n13709) );
  NAND2X0 U14391 ( .IN1(n13556), .IN2(g151), .QN(n13708) );
  NAND2X0 U14392 ( .IN1(n13710), .IN2(n13711), .QN(g22038) );
  NAND2X0 U14393 ( .IN1(n4328), .IN2(n13512), .QN(n13711) );
  INVX0 U14394 ( .INP(n13712), .ZN(n13710) );
  NOR2X0 U14395 ( .IN1(n13512), .IN2(n7933), .QN(n13712) );
  NAND2X0 U14396 ( .IN1(n13713), .IN2(n13714), .QN(g22037) );
  NAND2X0 U14397 ( .IN1(test_so11), .IN2(n13020), .QN(n13714) );
  NAND2X0 U14398 ( .IN1(n13469), .IN2(n4392), .QN(n13713) );
  NAND2X0 U14399 ( .IN1(n13715), .IN2(n13716), .QN(g22035) );
  NAND2X0 U14400 ( .IN1(n13454), .IN2(n4320), .QN(n13716) );
  INVX0 U14401 ( .INP(n13717), .ZN(n13715) );
  NOR2X0 U14402 ( .IN1(n13454), .IN2(n7894), .QN(n13717) );
  NOR2X0 U14403 ( .IN1(n4317), .IN2(n7707), .QN(n13454) );
  NAND2X0 U14404 ( .IN1(n13718), .IN2(n13719), .QN(g22034) );
  NAND2X0 U14405 ( .IN1(n13503), .IN2(n4391), .QN(n13719) );
  NAND2X0 U14406 ( .IN1(n13504), .IN2(g833), .QN(n13718) );
  NAND2X0 U14407 ( .IN1(n13720), .IN2(n13721), .QN(g22033) );
  NAND2X0 U14408 ( .IN1(n4321), .IN2(n13462), .QN(n13721) );
  INVX0 U14409 ( .INP(n13722), .ZN(n13720) );
  NOR2X0 U14410 ( .IN1(n13462), .IN2(n7908), .QN(n13722) );
  NOR2X0 U14411 ( .IN1(n4312), .IN2(n7708), .QN(n13462) );
  NAND2X0 U14412 ( .IN1(n13723), .IN2(n13724), .QN(g22032) );
  NAND2X0 U14413 ( .IN1(n4328), .IN2(n13555), .QN(n13724) );
  NAND2X0 U14414 ( .IN1(n13556), .IN2(g148), .QN(n13723) );
  NAND2X0 U14415 ( .IN1(n13725), .IN2(n13726), .QN(g22031) );
  NAND2X0 U14416 ( .IN1(n13512), .IN2(n4392), .QN(n13726) );
  INVX0 U14417 ( .INP(n13727), .ZN(n13725) );
  NOR2X0 U14418 ( .IN1(n13512), .IN2(n7935), .QN(n13727) );
  NAND2X0 U14419 ( .IN1(n13728), .IN2(n13729), .QN(g22030) );
  NAND2X0 U14420 ( .IN1(n4322), .IN2(n13469), .QN(n13729) );
  NAND2X0 U14421 ( .IN1(n13020), .IN2(g141), .QN(n13728) );
  INVX0 U14422 ( .INP(n13469), .ZN(n13020) );
  NOR2X0 U14423 ( .IN1(n4369), .IN2(n7709), .QN(n13469) );
  NAND2X0 U14424 ( .IN1(n13730), .IN2(n13731), .QN(g22029) );
  NAND2X0 U14425 ( .IN1(n4321), .IN2(n13503), .QN(n13731) );
  NAND2X0 U14426 ( .IN1(n13504), .IN2(g830), .QN(n13730) );
  INVX0 U14427 ( .INP(n13503), .ZN(n13504) );
  NOR2X0 U14428 ( .IN1(n4323), .IN2(n7708), .QN(n13503) );
  NAND2X0 U14429 ( .IN1(n13732), .IN2(n13733), .QN(g22028) );
  NAND2X0 U14430 ( .IN1(n13555), .IN2(n4392), .QN(n13733) );
  NAND2X0 U14431 ( .IN1(n13556), .IN2(g145), .QN(n13732) );
  NAND2X0 U14432 ( .IN1(n13734), .IN2(n13735), .QN(g22027) );
  NAND2X0 U14433 ( .IN1(n4322), .IN2(n13512), .QN(n13735) );
  INVX0 U14434 ( .INP(n13736), .ZN(n13734) );
  NOR2X0 U14435 ( .IN1(n13512), .IN2(n7947), .QN(n13736) );
  NOR2X0 U14436 ( .IN1(n4512), .IN2(n7709), .QN(n13512) );
  NOR2X0 U14437 ( .IN1(n8672), .IN2(n13737), .QN(g22026) );
  XOR2X1 U14438 ( .IN1(n8016), .IN2(n13264), .Q(n13737) );
  NOR2X0 U14439 ( .IN1(n4423), .IN2(n4330), .QN(n13264) );
  NAND2X0 U14440 ( .IN1(n14350), .IN2(n8677), .QN(n8672) );
  NAND4X0 U14441 ( .IN1(n4182), .IN2(n4431), .IN3(n4330), .IN4(n13738), .QN(
        n8677) );
  NOR4X0 U14442 ( .IN1(n8016), .IN2(n4423), .IN3(n4355), .IN4(g2900), .QN(
        n13738) );
  NAND2X0 U14443 ( .IN1(n13739), .IN2(n13740), .QN(g22025) );
  NAND2X0 U14444 ( .IN1(n4322), .IN2(n13555), .QN(n13740) );
  NAND2X0 U14445 ( .IN1(n13556), .IN2(g142), .QN(n13739) );
  INVX0 U14446 ( .INP(n13555), .ZN(n13556) );
  NOR2X0 U14447 ( .IN1(n4318), .IN2(n7709), .QN(n13555) );
  NAND2X0 U14448 ( .IN1(n13741), .IN2(n13742), .QN(g21970) );
  NAND2X0 U14449 ( .IN1(test_so87), .IN2(n4463), .QN(n13742) );
  NAND2X0 U14450 ( .IN1(n11339), .IN2(g2560), .QN(n13741) );
  NAND3X0 U14451 ( .IN1(n13743), .IN2(n13744), .IN3(n13745), .QN(n11339) );
  NAND2X0 U14452 ( .IN1(g5555), .IN2(g2513), .QN(n13745) );
  NAND2X0 U14453 ( .IN1(n4606), .IN2(g2519), .QN(n13744) );
  NAND2X0 U14454 ( .IN1(g7264), .IN2(g2516), .QN(n13743) );
  NAND2X0 U14455 ( .IN1(n13746), .IN2(n13747), .QN(g21882) );
  NAND2X0 U14456 ( .IN1(n4351), .IN2(g2878), .QN(n13747) );
  NAND2X0 U14457 ( .IN1(n13748), .IN2(g2879), .QN(n13746) );
  NAND2X0 U14458 ( .IN1(n13749), .IN2(n13750), .QN(g21880) );
  NAND2X0 U14459 ( .IN1(n4351), .IN2(g2877), .QN(n13750) );
  NAND2X0 U14460 ( .IN1(n13751), .IN2(g2879), .QN(n13749) );
  NAND2X0 U14461 ( .IN1(n13752), .IN2(n13753), .QN(g21878) );
  NAND2X0 U14462 ( .IN1(test_so4), .IN2(g2879), .QN(n13753) );
  NAND2X0 U14463 ( .IN1(n13748), .IN2(n4351), .QN(n13752) );
  XNOR2X1 U14464 ( .IN1(n8549), .IN2(n13754), .Q(n13748) );
  XOR3X1 U14465 ( .IN1(n13755), .IN2(n13756), .IN3(n13757), .Q(n8549) );
  XOR3X1 U14466 ( .IN1(n7999), .IN2(n7998), .IN3(n13758), .Q(n13757) );
  XOR2X1 U14467 ( .IN1(g2981), .IN2(test_so2), .Q(n13758) );
  XOR2X1 U14468 ( .IN1(n7995), .IN2(n7994), .Q(n13756) );
  XOR2X1 U14469 ( .IN1(n7997), .IN2(n7996), .Q(n13755) );
  NAND2X0 U14470 ( .IN1(n13759), .IN2(n13760), .QN(g21851) );
  NAND2X0 U14471 ( .IN1(g499), .IN2(g544), .QN(n13760) );
  NAND3X0 U14472 ( .IN1(n4298), .IN2(g548), .IN3(n4541), .QN(n13759) );
  NAND2X0 U14473 ( .IN1(n13761), .IN2(n13762), .QN(g21346) );
  NAND2X0 U14474 ( .IN1(n14355), .IN2(DFF_328_n1), .QN(n13762) );
  INVX0 U14475 ( .INP(n13763), .ZN(n13761) );
  NOR3X0 U14476 ( .IN1(g6447), .IN2(n7433), .IN3(n14355), .QN(n13763) );
  NAND2X0 U14477 ( .IN1(n13764), .IN2(n13765), .QN(g21094) );
  NAND2X0 U14478 ( .IN1(test_so94), .IN2(n12590), .QN(n13765) );
  NAND2X0 U14479 ( .IN1(n4393), .IN2(n12592), .QN(n13764) );
  NAND2X0 U14480 ( .IN1(n13766), .IN2(n13767), .QN(g21082) );
  NAND2X0 U14481 ( .IN1(n4393), .IN2(n12596), .QN(n13767) );
  NAND2X0 U14482 ( .IN1(n12595), .IN2(g2798), .QN(n13766) );
  NAND2X0 U14483 ( .IN1(n13768), .IN2(n13769), .QN(g21081) );
  NAND2X0 U14484 ( .IN1(n12592), .IN2(n4471), .QN(n13769) );
  NAND2X0 U14485 ( .IN1(n12590), .IN2(g2793), .QN(n13768) );
  NAND2X0 U14486 ( .IN1(n13770), .IN2(n13771), .QN(g21080) );
  NAND2X0 U14487 ( .IN1(n12601), .IN2(n8085), .QN(n13771) );
  NAND2X0 U14488 ( .IN1(n12599), .IN2(g2102), .QN(n13770) );
  NAND2X0 U14489 ( .IN1(n13772), .IN2(n13773), .QN(g21075) );
  NAND2X0 U14490 ( .IN1(n4393), .IN2(n12605), .QN(n13773) );
  NAND2X0 U14491 ( .IN1(n12604), .IN2(g2797), .QN(n13772) );
  NAND2X0 U14492 ( .IN1(n13774), .IN2(n13775), .QN(g21074) );
  NAND2X0 U14493 ( .IN1(n12596), .IN2(n4471), .QN(n13775) );
  NAND2X0 U14494 ( .IN1(n12595), .IN2(g2795), .QN(n13774) );
  NAND2X0 U14495 ( .IN1(n13776), .IN2(n13777), .QN(g21073) );
  NAND2X0 U14496 ( .IN1(n12592), .IN2(n8073), .QN(n13777) );
  NAND2X0 U14497 ( .IN1(n12590), .IN2(g2790), .QN(n13776) );
  NAND2X0 U14498 ( .IN1(n13778), .IN2(n13779), .QN(g21072) );
  NAND2X0 U14499 ( .IN1(n12661), .IN2(n8085), .QN(n13779) );
  NAND2X0 U14500 ( .IN1(n9317), .IN2(g2104), .QN(n13778) );
  NAND2X0 U14501 ( .IN1(n13780), .IN2(n13781), .QN(g21071) );
  NAND2X0 U14502 ( .IN1(n12601), .IN2(n4473), .QN(n13781) );
  NAND2X0 U14503 ( .IN1(n12599), .IN2(g2099), .QN(n13780) );
  NAND2X0 U14504 ( .IN1(n13782), .IN2(n13783), .QN(g21070) );
  NAND2X0 U14505 ( .IN1(n4395), .IN2(n12665), .QN(n13783) );
  INVX0 U14506 ( .INP(n13784), .ZN(n13782) );
  NOR2X0 U14507 ( .IN1(n12665), .IN2(n7846), .QN(n13784) );
  NAND2X0 U14508 ( .IN1(n13785), .IN2(n13786), .QN(g21063) );
  NAND2X0 U14509 ( .IN1(n13787), .IN2(g2805), .QN(n13786) );
  NAND2X0 U14510 ( .IN1(n13369), .IN2(n13788), .QN(n13785) );
  NAND2X0 U14511 ( .IN1(n13789), .IN2(n13790), .QN(g21062) );
  NAND2X0 U14512 ( .IN1(n12605), .IN2(n4471), .QN(n13790) );
  NAND2X0 U14513 ( .IN1(n12604), .IN2(g2794), .QN(n13789) );
  NAND2X0 U14514 ( .IN1(n13791), .IN2(n13792), .QN(g21061) );
  NAND2X0 U14515 ( .IN1(n12596), .IN2(n8073), .QN(n13792) );
  NAND2X0 U14516 ( .IN1(n12595), .IN2(g2792), .QN(n13791) );
  NAND2X0 U14517 ( .IN1(n13793), .IN2(n13794), .QN(g21060) );
  NAND2X0 U14518 ( .IN1(n12592), .IN2(n4407), .QN(n13794) );
  NAND2X0 U14519 ( .IN1(n12590), .IN2(g2787), .QN(n13793) );
  NAND2X0 U14520 ( .IN1(n13795), .IN2(n13796), .QN(g21056) );
  NAND2X0 U14521 ( .IN1(n12670), .IN2(n8085), .QN(n13796) );
  NAND2X0 U14522 ( .IN1(n12669), .IN2(g2103), .QN(n13795) );
  NAND2X0 U14523 ( .IN1(n13797), .IN2(n13798), .QN(g21055) );
  NAND2X0 U14524 ( .IN1(n12661), .IN2(n4473), .QN(n13798) );
  NAND2X0 U14525 ( .IN1(n9317), .IN2(g2101), .QN(n13797) );
  NAND2X0 U14526 ( .IN1(n13799), .IN2(n13800), .QN(g21054) );
  NAND2X0 U14527 ( .IN1(n4468), .IN2(n12601), .QN(n13800) );
  NAND2X0 U14528 ( .IN1(n12599), .IN2(g2096), .QN(n13799) );
  NAND2X0 U14529 ( .IN1(n13801), .IN2(n13802), .QN(g21053) );
  NAND2X0 U14530 ( .IN1(n4395), .IN2(n12726), .QN(n13802) );
  NAND2X0 U14531 ( .IN1(n8518), .IN2(g1410), .QN(n13801) );
  NAND2X0 U14532 ( .IN1(n13803), .IN2(n13804), .QN(g21052) );
  NAND2X0 U14533 ( .IN1(n12665), .IN2(n4475), .QN(n13804) );
  INVX0 U14534 ( .INP(n13805), .ZN(n13803) );
  NOR2X0 U14535 ( .IN1(n12665), .IN2(n7847), .QN(n13805) );
  NAND2X0 U14536 ( .IN1(n13806), .IN2(n13807), .QN(g21051) );
  NAND2X0 U14537 ( .IN1(n4396), .IN2(n12731), .QN(n13807) );
  NAND2X0 U14538 ( .IN1(n12729), .IN2(g722), .QN(n13806) );
  NAND2X0 U14539 ( .IN1(n13808), .IN2(n13809), .QN(g21047) );
  NAND2X0 U14540 ( .IN1(n9289), .IN2(g2807), .QN(n13809) );
  NAND2X0 U14541 ( .IN1(n11303), .IN2(n13788), .QN(n13808) );
  NAND2X0 U14542 ( .IN1(n13810), .IN2(n13811), .QN(g21046) );
  NAND2X0 U14543 ( .IN1(n13787), .IN2(g2802), .QN(n13811) );
  NAND2X0 U14544 ( .IN1(n13369), .IN2(n8901), .QN(n13810) );
  INVX0 U14545 ( .INP(n13787), .ZN(n13369) );
  NAND2X0 U14546 ( .IN1(g2703), .IN2(g2704), .QN(n13787) );
  NAND2X0 U14547 ( .IN1(n13812), .IN2(n13813), .QN(g21045) );
  NAND2X0 U14548 ( .IN1(n12605), .IN2(n8073), .QN(n13813) );
  NAND2X0 U14549 ( .IN1(n12604), .IN2(g2791), .QN(n13812) );
  NAND2X0 U14550 ( .IN1(n13814), .IN2(n13815), .QN(g21044) );
  NAND2X0 U14551 ( .IN1(n12596), .IN2(n4407), .QN(n13815) );
  NAND2X0 U14552 ( .IN1(n12595), .IN2(g2789), .QN(n13814) );
  NAND2X0 U14553 ( .IN1(n13816), .IN2(n13817), .QN(g21043) );
  NAND2X0 U14554 ( .IN1(n4397), .IN2(n12592), .QN(n13817) );
  NAND2X0 U14555 ( .IN1(n12590), .IN2(g2784), .QN(n13816) );
  NAND2X0 U14556 ( .IN1(n13818), .IN2(n13819), .QN(g21042) );
  NAND2X0 U14557 ( .IN1(n13820), .IN2(g2111), .QN(n13819) );
  NAND2X0 U14558 ( .IN1(n13373), .IN2(n13821), .QN(n13818) );
  NAND2X0 U14559 ( .IN1(n13822), .IN2(n13823), .QN(g21041) );
  NAND2X0 U14560 ( .IN1(n12670), .IN2(n4473), .QN(n13823) );
  NAND2X0 U14561 ( .IN1(n12669), .IN2(g2100), .QN(n13822) );
  NAND2X0 U14562 ( .IN1(n13824), .IN2(n13825), .QN(g21040) );
  NAND2X0 U14563 ( .IN1(n4468), .IN2(n12661), .QN(n13825) );
  NAND2X0 U14564 ( .IN1(n9317), .IN2(g2098), .QN(n13824) );
  NAND2X0 U14565 ( .IN1(n13826), .IN2(n13827), .QN(g21039) );
  NAND2X0 U14566 ( .IN1(n12601), .IN2(n4409), .QN(n13827) );
  NAND2X0 U14567 ( .IN1(n12599), .IN2(g2093), .QN(n13826) );
  NAND2X0 U14568 ( .IN1(n13828), .IN2(n13829), .QN(g21035) );
  NAND2X0 U14569 ( .IN1(n4395), .IN2(n12738), .QN(n13829) );
  NAND2X0 U14570 ( .IN1(n12737), .IN2(g1409), .QN(n13828) );
  NAND2X0 U14571 ( .IN1(n13830), .IN2(n13831), .QN(g21034) );
  NAND2X0 U14572 ( .IN1(n12726), .IN2(n4475), .QN(n13831) );
  NAND2X0 U14573 ( .IN1(n8518), .IN2(g1407), .QN(n13830) );
  NAND2X0 U14574 ( .IN1(n13832), .IN2(n13833), .QN(g21033) );
  NAND2X0 U14575 ( .IN1(n4469), .IN2(n12665), .QN(n13833) );
  INVX0 U14576 ( .INP(n13834), .ZN(n13832) );
  NOR2X0 U14577 ( .IN1(n12665), .IN2(n7848), .QN(n13834) );
  NAND2X0 U14578 ( .IN1(n13835), .IN2(n13836), .QN(g21032) );
  NAND2X0 U14579 ( .IN1(n4396), .IN2(n12794), .QN(n13836) );
  NAND2X0 U14580 ( .IN1(n8539), .IN2(g724), .QN(n13835) );
  NAND2X0 U14581 ( .IN1(n13837), .IN2(n13838), .QN(g21031) );
  NAND2X0 U14582 ( .IN1(n12731), .IN2(n4477), .QN(n13838) );
  NAND2X0 U14583 ( .IN1(n12729), .IN2(g719), .QN(n13837) );
  NAND2X0 U14584 ( .IN1(n13839), .IN2(n13840), .QN(g21029) );
  INVX0 U14585 ( .INP(n13841), .ZN(n13840) );
  NOR2X0 U14586 ( .IN1(n13375), .IN2(n7563), .QN(n13841) );
  NAND2X0 U14587 ( .IN1(n13375), .IN2(n13788), .QN(n13839) );
  INVX0 U14588 ( .INP(n8865), .ZN(n13788) );
  NAND3X0 U14589 ( .IN1(n13842), .IN2(n13843), .IN3(n13844), .QN(n8865) );
  NAND2X0 U14590 ( .IN1(test_so90), .IN2(g7390), .QN(n13844) );
  NAND2X0 U14591 ( .IN1(g7302), .IN2(g2679), .QN(n13843) );
  NAND2X0 U14592 ( .IN1(g2624), .IN2(g2685), .QN(n13842) );
  NAND2X0 U14593 ( .IN1(n13845), .IN2(n13846), .QN(g21028) );
  NAND2X0 U14594 ( .IN1(n9289), .IN2(g2804), .QN(n13846) );
  NAND2X0 U14595 ( .IN1(n11303), .IN2(n8901), .QN(n13845) );
  NAND2X0 U14596 ( .IN1(n13847), .IN2(n13848), .QN(g21027) );
  NAND2X0 U14597 ( .IN1(n12605), .IN2(n4407), .QN(n13848) );
  NAND2X0 U14598 ( .IN1(n12604), .IN2(g2788), .QN(n13847) );
  NAND2X0 U14599 ( .IN1(n13849), .IN2(n13850), .QN(g21026) );
  NAND2X0 U14600 ( .IN1(n4397), .IN2(n12596), .QN(n13850) );
  NAND2X0 U14601 ( .IN1(n12595), .IN2(g2786), .QN(n13849) );
  NAND2X0 U14602 ( .IN1(n13851), .IN2(n13852), .QN(g21025) );
  NAND2X0 U14603 ( .IN1(test_so93), .IN2(n12590), .QN(n13852) );
  NAND2X0 U14604 ( .IN1(n12592), .IN2(n4408), .QN(n13851) );
  NAND2X0 U14605 ( .IN1(n13853), .IN2(n13854), .QN(g21023) );
  NAND2X0 U14606 ( .IN1(n9311), .IN2(g2113), .QN(n13854) );
  NAND2X0 U14607 ( .IN1(n9305), .IN2(n13821), .QN(n13853) );
  NAND2X0 U14608 ( .IN1(n13855), .IN2(n13856), .QN(g21022) );
  NAND2X0 U14609 ( .IN1(n13820), .IN2(g2108), .QN(n13856) );
  INVX0 U14610 ( .INP(n13373), .ZN(n13820) );
  NAND2X0 U14611 ( .IN1(n13373), .IN2(n8992), .QN(n13855) );
  NOR2X0 U14612 ( .IN1(n4293), .IN2(n7746), .QN(n13373) );
  NAND2X0 U14613 ( .IN1(n13857), .IN2(n13858), .QN(g21021) );
  NAND2X0 U14614 ( .IN1(n4468), .IN2(n12670), .QN(n13858) );
  NAND2X0 U14615 ( .IN1(n12669), .IN2(g2097), .QN(n13857) );
  NAND2X0 U14616 ( .IN1(n13859), .IN2(n13860), .QN(g21020) );
  NAND2X0 U14617 ( .IN1(n12661), .IN2(n4409), .QN(n13860) );
  NAND2X0 U14618 ( .IN1(n9317), .IN2(g2095), .QN(n13859) );
  NAND2X0 U14619 ( .IN1(n13861), .IN2(n13862), .QN(g21019) );
  NAND2X0 U14620 ( .IN1(n4399), .IN2(n12601), .QN(n13862) );
  NAND2X0 U14621 ( .IN1(n12599), .IN2(g2090), .QN(n13861) );
  NAND2X0 U14622 ( .IN1(n13863), .IN2(n13864), .QN(g21018) );
  NAND2X0 U14623 ( .IN1(n13865), .IN2(g1417), .QN(n13864) );
  NAND2X0 U14624 ( .IN1(n13378), .IN2(n13866), .QN(n13863) );
  NAND2X0 U14625 ( .IN1(n13867), .IN2(n13868), .QN(g21017) );
  NAND2X0 U14626 ( .IN1(n12738), .IN2(n4475), .QN(n13868) );
  NAND2X0 U14627 ( .IN1(n12737), .IN2(g1406), .QN(n13867) );
  NAND2X0 U14628 ( .IN1(n13869), .IN2(n13870), .QN(g21016) );
  NAND2X0 U14629 ( .IN1(n4469), .IN2(n12726), .QN(n13870) );
  NAND2X0 U14630 ( .IN1(n8518), .IN2(g1404), .QN(n13869) );
  NAND2X0 U14631 ( .IN1(n13871), .IN2(n13872), .QN(g21015) );
  NAND2X0 U14632 ( .IN1(n12665), .IN2(n4411), .QN(n13872) );
  INVX0 U14633 ( .INP(n13873), .ZN(n13871) );
  NOR2X0 U14634 ( .IN1(n12665), .IN2(n7849), .QN(n13873) );
  NAND2X0 U14635 ( .IN1(n13874), .IN2(n13875), .QN(g21011) );
  NAND2X0 U14636 ( .IN1(n4396), .IN2(n12798), .QN(n13875) );
  NAND2X0 U14637 ( .IN1(n12797), .IN2(g723), .QN(n13874) );
  NAND2X0 U14638 ( .IN1(n13876), .IN2(n13877), .QN(g21010) );
  NAND2X0 U14639 ( .IN1(n12794), .IN2(n4477), .QN(n13877) );
  NAND2X0 U14640 ( .IN1(n8539), .IN2(g721), .QN(n13876) );
  NAND2X0 U14641 ( .IN1(n13878), .IN2(n13879), .QN(g21009) );
  NAND2X0 U14642 ( .IN1(n12731), .IN2(n8074), .QN(n13879) );
  NAND2X0 U14643 ( .IN1(n12729), .IN2(g716), .QN(n13878) );
  NAND2X0 U14644 ( .IN1(n13880), .IN2(n13881), .QN(g21007) );
  INVX0 U14645 ( .INP(n13882), .ZN(n13881) );
  NOR2X0 U14646 ( .IN1(n13375), .IN2(n8029), .QN(n13882) );
  NAND2X0 U14647 ( .IN1(n13375), .IN2(n8901), .QN(n13880) );
  INVX0 U14648 ( .INP(n8876), .ZN(n8901) );
  NAND3X0 U14649 ( .IN1(n13883), .IN2(n13884), .IN3(n13885), .QN(n8876) );
  NAND2X0 U14650 ( .IN1(g7390), .IN2(g2691), .QN(n13885) );
  NAND2X0 U14651 ( .IN1(g2624), .IN2(g2694), .QN(n13884) );
  NAND2X0 U14652 ( .IN1(n10166), .IN2(g2688), .QN(n13883) );
  INVX0 U14653 ( .INP(n4314), .ZN(n10166) );
  NOR2X0 U14654 ( .IN1(n4306), .IN2(n7745), .QN(n13375) );
  NAND2X0 U14655 ( .IN1(n13886), .IN2(n13887), .QN(g21006) );
  NAND2X0 U14656 ( .IN1(n4397), .IN2(n12605), .QN(n13887) );
  NAND2X0 U14657 ( .IN1(n12604), .IN2(g2785), .QN(n13886) );
  NAND2X0 U14658 ( .IN1(n13888), .IN2(n13889), .QN(g21005) );
  NAND2X0 U14659 ( .IN1(n12596), .IN2(n4408), .QN(n13889) );
  NAND2X0 U14660 ( .IN1(n12595), .IN2(g2783), .QN(n13888) );
  NAND2X0 U14661 ( .IN1(n13890), .IN2(n13891), .QN(g21004) );
  NAND2X0 U14662 ( .IN1(n4419), .IN2(n12592), .QN(n13891) );
  NAND2X0 U14663 ( .IN1(n12590), .IN2(g2778), .QN(n13890) );
  NAND2X0 U14664 ( .IN1(n13892), .IN2(n13893), .QN(g21003) );
  INVX0 U14665 ( .INP(n13894), .ZN(n13893) );
  NOR2X0 U14666 ( .IN1(n13380), .IN2(n7564), .QN(n13894) );
  NAND2X0 U14667 ( .IN1(n13380), .IN2(n13821), .QN(n13892) );
  INVX0 U14668 ( .INP(n8980), .ZN(n13821) );
  NAND3X0 U14669 ( .IN1(n13895), .IN2(n13896), .IN3(n13897), .QN(n8980) );
  NAND2X0 U14670 ( .IN1(g1930), .IN2(g1991), .QN(n13897) );
  NAND2X0 U14671 ( .IN1(g7052), .IN2(g1985), .QN(n13896) );
  NAND2X0 U14672 ( .IN1(g7194), .IN2(g1988), .QN(n13895) );
  NAND2X0 U14673 ( .IN1(n13898), .IN2(n13899), .QN(g21002) );
  NAND2X0 U14674 ( .IN1(n9311), .IN2(g2110), .QN(n13899) );
  INVX0 U14675 ( .INP(n9305), .ZN(n9311) );
  NAND2X0 U14676 ( .IN1(n9305), .IN2(n8992), .QN(n13898) );
  NAND2X0 U14677 ( .IN1(n13900), .IN2(n13901), .QN(g21001) );
  NAND2X0 U14678 ( .IN1(n12670), .IN2(n4409), .QN(n13901) );
  NAND2X0 U14679 ( .IN1(n12669), .IN2(g2094), .QN(n13900) );
  NAND2X0 U14680 ( .IN1(n13902), .IN2(n13903), .QN(g21000) );
  NAND2X0 U14681 ( .IN1(test_so71), .IN2(n9317), .QN(n13903) );
  NAND2X0 U14682 ( .IN1(n4399), .IN2(n12661), .QN(n13902) );
  NAND2X0 U14683 ( .IN1(n13904), .IN2(n13905), .QN(g20999) );
  NAND2X0 U14684 ( .IN1(n12601), .IN2(n4410), .QN(n13905) );
  NAND2X0 U14685 ( .IN1(n12599), .IN2(g2087), .QN(n13904) );
  NAND2X0 U14686 ( .IN1(n13906), .IN2(n13907), .QN(g20997) );
  NAND2X0 U14687 ( .IN1(n8507), .IN2(g1419), .QN(n13907) );
  NAND2X0 U14688 ( .IN1(n8512), .IN2(n13866), .QN(n13906) );
  NAND2X0 U14689 ( .IN1(n13908), .IN2(n13909), .QN(g20996) );
  NAND2X0 U14690 ( .IN1(test_so51), .IN2(n13865), .QN(n13909) );
  INVX0 U14691 ( .INP(n13378), .ZN(n13865) );
  NAND2X0 U14692 ( .IN1(n13378), .IN2(n9120), .QN(n13908) );
  NOR2X0 U14693 ( .IN1(n4294), .IN2(n7747), .QN(n13378) );
  NAND2X0 U14694 ( .IN1(n13910), .IN2(n13911), .QN(g20995) );
  NAND2X0 U14695 ( .IN1(n4469), .IN2(n12738), .QN(n13911) );
  NAND2X0 U14696 ( .IN1(n12737), .IN2(g1403), .QN(n13910) );
  NAND2X0 U14697 ( .IN1(n13912), .IN2(n13913), .QN(g20994) );
  NAND2X0 U14698 ( .IN1(test_so50), .IN2(n8518), .QN(n13913) );
  NAND2X0 U14699 ( .IN1(n12726), .IN2(n4411), .QN(n13912) );
  NAND2X0 U14700 ( .IN1(n13914), .IN2(n13915), .QN(g20993) );
  NAND2X0 U14701 ( .IN1(n4401), .IN2(n12665), .QN(n13915) );
  INVX0 U14702 ( .INP(n13916), .ZN(n13914) );
  NOR2X0 U14703 ( .IN1(n12665), .IN2(n7850), .QN(n13916) );
  NAND2X0 U14704 ( .IN1(n13917), .IN2(n13918), .QN(g20992) );
  NAND2X0 U14705 ( .IN1(n13919), .IN2(g731), .QN(n13918) );
  NAND2X0 U14706 ( .IN1(n13383), .IN2(n13920), .QN(n13917) );
  NAND2X0 U14707 ( .IN1(n13921), .IN2(n13922), .QN(g20991) );
  NAND2X0 U14708 ( .IN1(n12798), .IN2(n4477), .QN(n13922) );
  NAND2X0 U14709 ( .IN1(n12797), .IN2(g720), .QN(n13921) );
  NAND2X0 U14710 ( .IN1(n13923), .IN2(n13924), .QN(g20990) );
  NAND2X0 U14711 ( .IN1(n12794), .IN2(n8074), .QN(n13924) );
  NAND2X0 U14712 ( .IN1(n8539), .IN2(g718), .QN(n13923) );
  NAND2X0 U14713 ( .IN1(n13925), .IN2(n13926), .QN(g20989) );
  NAND2X0 U14714 ( .IN1(n12731), .IN2(n4413), .QN(n13926) );
  NAND2X0 U14715 ( .IN1(n12729), .IN2(g713), .QN(n13925) );
  NAND2X0 U14716 ( .IN1(n13927), .IN2(n13928), .QN(g20983) );
  NAND2X0 U14717 ( .IN1(n12605), .IN2(n4408), .QN(n13928) );
  NAND2X0 U14718 ( .IN1(n12604), .IN2(g2782), .QN(n13927) );
  NAND2X0 U14719 ( .IN1(n13929), .IN2(n13930), .QN(g20982) );
  NAND2X0 U14720 ( .IN1(n4419), .IN2(n12596), .QN(n13930) );
  NAND2X0 U14721 ( .IN1(n12595), .IN2(g2780), .QN(n13929) );
  NAND2X0 U14722 ( .IN1(n13931), .IN2(n13932), .QN(g20981) );
  NAND2X0 U14723 ( .IN1(n12592), .IN2(n4472), .QN(n13932) );
  NAND2X0 U14724 ( .IN1(n12590), .IN2(g2775), .QN(n13931) );
  NAND2X0 U14725 ( .IN1(n13933), .IN2(n13934), .QN(g20980) );
  INVX0 U14726 ( .INP(n13935), .ZN(n13934) );
  NOR2X0 U14727 ( .IN1(n13380), .IN2(n8028), .QN(n13935) );
  NAND2X0 U14728 ( .IN1(n13380), .IN2(n8992), .QN(n13933) );
  INVX0 U14729 ( .INP(n9002), .ZN(n8992) );
  NAND3X0 U14730 ( .IN1(n13936), .IN2(n13937), .IN3(n13938), .QN(n9002) );
  NAND2X0 U14731 ( .IN1(g1930), .IN2(g2000), .QN(n13938) );
  NAND2X0 U14732 ( .IN1(n10214), .IN2(g1994), .QN(n13937) );
  INVX0 U14733 ( .INP(n4296), .ZN(n10214) );
  NAND2X0 U14734 ( .IN1(g7194), .IN2(g1997), .QN(n13936) );
  NOR2X0 U14735 ( .IN1(n4307), .IN2(n7746), .QN(n13380) );
  NAND2X0 U14736 ( .IN1(n13939), .IN2(n13940), .QN(g20979) );
  NAND2X0 U14737 ( .IN1(n4399), .IN2(n12670), .QN(n13940) );
  NAND2X0 U14738 ( .IN1(n12669), .IN2(g2091), .QN(n13939) );
  NAND2X0 U14739 ( .IN1(n13941), .IN2(n13942), .QN(g20978) );
  NAND2X0 U14740 ( .IN1(n12661), .IN2(n4410), .QN(n13942) );
  NAND2X0 U14741 ( .IN1(n9317), .IN2(g2089), .QN(n13941) );
  NAND2X0 U14742 ( .IN1(n13943), .IN2(n13944), .QN(g20977) );
  NAND2X0 U14743 ( .IN1(n4420), .IN2(n12601), .QN(n13944) );
  NAND2X0 U14744 ( .IN1(n12599), .IN2(g2084), .QN(n13943) );
  NAND2X0 U14745 ( .IN1(n13945), .IN2(n13946), .QN(g20976) );
  INVX0 U14746 ( .INP(n13947), .ZN(n13946) );
  NOR2X0 U14747 ( .IN1(n13385), .IN2(n7565), .QN(n13947) );
  NAND2X0 U14748 ( .IN1(n13385), .IN2(n13866), .QN(n13945) );
  INVX0 U14749 ( .INP(n9097), .ZN(n13866) );
  NAND3X0 U14750 ( .IN1(n13948), .IN2(n13949), .IN3(n13950), .QN(n9097) );
  NAND2X0 U14751 ( .IN1(g6944), .IN2(g1294), .QN(n13950) );
  NAND2X0 U14752 ( .IN1(g6750), .IN2(g1291), .QN(n13949) );
  NAND2X0 U14753 ( .IN1(g1236), .IN2(g1297), .QN(n13948) );
  NAND2X0 U14754 ( .IN1(n13951), .IN2(n13952), .QN(g20975) );
  NAND2X0 U14755 ( .IN1(n8507), .IN2(g1416), .QN(n13952) );
  INVX0 U14756 ( .INP(n8512), .ZN(n8507) );
  NAND2X0 U14757 ( .IN1(n8512), .IN2(n9120), .QN(n13951) );
  NAND2X0 U14758 ( .IN1(n13953), .IN2(n13954), .QN(g20974) );
  NAND2X0 U14759 ( .IN1(n12738), .IN2(n4411), .QN(n13954) );
  NAND2X0 U14760 ( .IN1(n12737), .IN2(g1400), .QN(n13953) );
  NAND2X0 U14761 ( .IN1(n13955), .IN2(n13956), .QN(g20973) );
  NAND2X0 U14762 ( .IN1(n4401), .IN2(n12726), .QN(n13956) );
  NAND2X0 U14763 ( .IN1(n8518), .IN2(g1398), .QN(n13955) );
  NAND2X0 U14764 ( .IN1(n13957), .IN2(n13958), .QN(g20972) );
  NAND2X0 U14765 ( .IN1(n12665), .IN2(n4412), .QN(n13958) );
  INVX0 U14766 ( .INP(n13959), .ZN(n13957) );
  NOR2X0 U14767 ( .IN1(n12665), .IN2(n7851), .QN(n13959) );
  NAND2X0 U14768 ( .IN1(n13960), .IN2(n13961), .QN(g20970) );
  NAND2X0 U14769 ( .IN1(n8527), .IN2(g733), .QN(n13961) );
  NAND2X0 U14770 ( .IN1(n8536), .IN2(n13920), .QN(n13960) );
  NAND2X0 U14771 ( .IN1(n13962), .IN2(n13963), .QN(g20969) );
  NAND2X0 U14772 ( .IN1(n13919), .IN2(g728), .QN(n13963) );
  INVX0 U14773 ( .INP(n13383), .ZN(n13919) );
  NAND2X0 U14774 ( .IN1(n13383), .IN2(n13964), .QN(n13962) );
  NOR2X0 U14775 ( .IN1(n4295), .IN2(n7748), .QN(n13383) );
  NAND2X0 U14776 ( .IN1(n13965), .IN2(n13966), .QN(g20968) );
  NAND2X0 U14777 ( .IN1(n12798), .IN2(n8074), .QN(n13966) );
  NAND2X0 U14778 ( .IN1(n12797), .IN2(g717), .QN(n13965) );
  NAND2X0 U14779 ( .IN1(n13967), .IN2(n13968), .QN(g20967) );
  NAND2X0 U14780 ( .IN1(n12794), .IN2(n4413), .QN(n13968) );
  NAND2X0 U14781 ( .IN1(n8539), .IN2(g715), .QN(n13967) );
  NAND2X0 U14782 ( .IN1(n13969), .IN2(n13970), .QN(g20966) );
  NAND2X0 U14783 ( .IN1(n4403), .IN2(n12731), .QN(n13970) );
  NAND2X0 U14784 ( .IN1(n12729), .IN2(g710), .QN(n13969) );
  NAND2X0 U14785 ( .IN1(n13971), .IN2(n13972), .QN(g20965) );
  NAND2X0 U14786 ( .IN1(n4415), .IN2(n12592), .QN(n13972) );
  NAND2X0 U14787 ( .IN1(n12590), .IN2(g2799), .QN(n13971) );
  NAND2X0 U14788 ( .IN1(n13973), .IN2(n13974), .QN(g20964) );
  NAND2X0 U14789 ( .IN1(n4419), .IN2(n12605), .QN(n13974) );
  NAND2X0 U14790 ( .IN1(n12604), .IN2(g2779), .QN(n13973) );
  NAND2X0 U14791 ( .IN1(n13975), .IN2(n13976), .QN(g20963) );
  NAND2X0 U14792 ( .IN1(n12596), .IN2(n4472), .QN(n13976) );
  NAND2X0 U14793 ( .IN1(n12595), .IN2(g2777), .QN(n13975) );
  NAND2X0 U14794 ( .IN1(n13977), .IN2(n13978), .QN(g20962) );
  NAND2X0 U14795 ( .IN1(n4398), .IN2(n12592), .QN(n13978) );
  INVX0 U14796 ( .INP(n12590), .ZN(n12592) );
  NAND2X0 U14797 ( .IN1(n12590), .IN2(g2772), .QN(n13977) );
  NAND2X0 U14798 ( .IN1(n13979), .IN2(n9297), .QN(n12590) );
  NAND2X0 U14799 ( .IN1(n13980), .IN2(n13981), .QN(g20955) );
  NAND2X0 U14800 ( .IN1(n12670), .IN2(n4410), .QN(n13981) );
  NAND2X0 U14801 ( .IN1(n12669), .IN2(g2088), .QN(n13980) );
  NAND2X0 U14802 ( .IN1(n13982), .IN2(n13983), .QN(g20954) );
  NAND2X0 U14803 ( .IN1(n4420), .IN2(n12661), .QN(n13983) );
  NAND2X0 U14804 ( .IN1(n9317), .IN2(g2086), .QN(n13982) );
  NAND2X0 U14805 ( .IN1(n13984), .IN2(n13985), .QN(g20953) );
  NAND2X0 U14806 ( .IN1(n12601), .IN2(n4474), .QN(n13985) );
  NAND2X0 U14807 ( .IN1(n12599), .IN2(g2081), .QN(n13984) );
  NAND2X0 U14808 ( .IN1(n13986), .IN2(n13987), .QN(g20952) );
  INVX0 U14809 ( .INP(n13988), .ZN(n13987) );
  NOR2X0 U14810 ( .IN1(n13385), .IN2(n8023), .QN(n13988) );
  NAND2X0 U14811 ( .IN1(n13385), .IN2(n9120), .QN(n13986) );
  INVX0 U14812 ( .INP(n9108), .ZN(n9120) );
  NAND3X0 U14813 ( .IN1(n13989), .IN2(n13990), .IN3(n13991), .QN(n9108) );
  NAND2X0 U14814 ( .IN1(n11104), .IN2(g1300), .QN(n13991) );
  INVX0 U14815 ( .INP(n4371), .ZN(n11104) );
  NAND2X0 U14816 ( .IN1(g1236), .IN2(g1306), .QN(n13990) );
  NAND2X0 U14817 ( .IN1(g6944), .IN2(g1303), .QN(n13989) );
  NOR2X0 U14818 ( .IN1(n4308), .IN2(n7747), .QN(n13385) );
  NAND2X0 U14819 ( .IN1(n13992), .IN2(n13993), .QN(g20951) );
  NAND2X0 U14820 ( .IN1(n4401), .IN2(n12738), .QN(n13993) );
  NAND2X0 U14821 ( .IN1(n12737), .IN2(g1397), .QN(n13992) );
  NAND2X0 U14822 ( .IN1(n13994), .IN2(n13995), .QN(g20950) );
  NAND2X0 U14823 ( .IN1(n12726), .IN2(n4412), .QN(n13995) );
  NAND2X0 U14824 ( .IN1(n8518), .IN2(g1395), .QN(n13994) );
  NAND2X0 U14825 ( .IN1(n13996), .IN2(n13997), .QN(g20949) );
  NAND2X0 U14826 ( .IN1(n4421), .IN2(n12665), .QN(n13997) );
  INVX0 U14827 ( .INP(n13998), .ZN(n13996) );
  NOR2X0 U14828 ( .IN1(n12665), .IN2(n7852), .QN(n13998) );
  NAND2X0 U14829 ( .IN1(n13999), .IN2(n14000), .QN(g20948) );
  INVX0 U14830 ( .INP(n14001), .ZN(n14000) );
  NOR2X0 U14831 ( .IN1(n13388), .IN2(n7566), .QN(n14001) );
  NAND2X0 U14832 ( .IN1(n13388), .IN2(n13920), .QN(n13999) );
  INVX0 U14833 ( .INP(n8745), .ZN(n13920) );
  NAND3X0 U14834 ( .IN1(n14002), .IN2(n14003), .IN3(n14004), .QN(n8745) );
  NAND2X0 U14835 ( .IN1(g6642), .IN2(g608), .QN(n14004) );
  NAND2X0 U14836 ( .IN1(n11207), .IN2(g605), .QN(n14003) );
  INVX0 U14837 ( .INP(n4298), .ZN(n11207) );
  NAND2X0 U14838 ( .IN1(g550), .IN2(g611), .QN(n14002) );
  NAND2X0 U14839 ( .IN1(n14005), .IN2(n14006), .QN(g20947) );
  NAND2X0 U14840 ( .IN1(n8527), .IN2(g730), .QN(n14006) );
  INVX0 U14841 ( .INP(n8536), .ZN(n8527) );
  NAND2X0 U14842 ( .IN1(n8536), .IN2(n13964), .QN(n14005) );
  NAND2X0 U14843 ( .IN1(n14007), .IN2(n14008), .QN(g20946) );
  NAND2X0 U14844 ( .IN1(n12798), .IN2(n4413), .QN(n14008) );
  NAND2X0 U14845 ( .IN1(n12797), .IN2(g714), .QN(n14007) );
  NAND2X0 U14846 ( .IN1(n14009), .IN2(n14010), .QN(g20945) );
  NAND2X0 U14847 ( .IN1(n4403), .IN2(n12794), .QN(n14010) );
  NAND2X0 U14848 ( .IN1(n8539), .IN2(g712), .QN(n14009) );
  NAND2X0 U14849 ( .IN1(n14011), .IN2(n14012), .QN(g20944) );
  NAND2X0 U14850 ( .IN1(n12731), .IN2(n4414), .QN(n14012) );
  NAND2X0 U14851 ( .IN1(n12729), .IN2(g707), .QN(n14011) );
  NAND2X0 U14852 ( .IN1(n14013), .IN2(n14014), .QN(g20941) );
  NAND2X0 U14853 ( .IN1(n4415), .IN2(n12596), .QN(n14014) );
  NAND2X0 U14854 ( .IN1(n12595), .IN2(g2801), .QN(n14013) );
  NAND2X0 U14855 ( .IN1(n14015), .IN2(n14016), .QN(g20940) );
  NAND2X0 U14856 ( .IN1(n12605), .IN2(n4472), .QN(n14016) );
  NAND2X0 U14857 ( .IN1(n12604), .IN2(g2776), .QN(n14015) );
  NAND2X0 U14858 ( .IN1(n14017), .IN2(n14018), .QN(g20939) );
  NAND2X0 U14859 ( .IN1(n4398), .IN2(n12596), .QN(n14018) );
  INVX0 U14860 ( .INP(n12595), .ZN(n12596) );
  NAND2X0 U14861 ( .IN1(n12595), .IN2(g2774), .QN(n14017) );
  NAND3X0 U14862 ( .IN1(n4426), .IN2(g7487), .IN3(n13979), .QN(n12595) );
  NAND2X0 U14863 ( .IN1(n14019), .IN2(n14020), .QN(g20937) );
  NAND2X0 U14864 ( .IN1(n4416), .IN2(n12601), .QN(n14020) );
  NAND2X0 U14865 ( .IN1(n12599), .IN2(g2105), .QN(n14019) );
  NAND2X0 U14866 ( .IN1(n14021), .IN2(n14022), .QN(g20936) );
  NAND2X0 U14867 ( .IN1(n4420), .IN2(n12670), .QN(n14022) );
  NAND2X0 U14868 ( .IN1(n12669), .IN2(g2085), .QN(n14021) );
  NAND2X0 U14869 ( .IN1(n14023), .IN2(n14024), .QN(g20935) );
  NAND2X0 U14870 ( .IN1(n12661), .IN2(n4474), .QN(n14024) );
  NAND2X0 U14871 ( .IN1(n9317), .IN2(g2083), .QN(n14023) );
  NAND2X0 U14872 ( .IN1(n14025), .IN2(n14026), .QN(g20934) );
  NAND2X0 U14873 ( .IN1(n4400), .IN2(n12601), .QN(n14026) );
  INVX0 U14874 ( .INP(n12599), .ZN(n12601) );
  NAND2X0 U14875 ( .IN1(n12599), .IN2(g2078), .QN(n14025) );
  NAND2X0 U14876 ( .IN1(n14027), .IN2(n9314), .QN(n12599) );
  NAND2X0 U14877 ( .IN1(n14028), .IN2(n14029), .QN(g20927) );
  NAND2X0 U14878 ( .IN1(n12738), .IN2(n4412), .QN(n14029) );
  NAND2X0 U14879 ( .IN1(n12737), .IN2(g1394), .QN(n14028) );
  NAND2X0 U14880 ( .IN1(n14030), .IN2(n14031), .QN(g20926) );
  NAND2X0 U14881 ( .IN1(n4421), .IN2(n12726), .QN(n14031) );
  NAND2X0 U14882 ( .IN1(n8518), .IN2(g1392), .QN(n14030) );
  NAND2X0 U14883 ( .IN1(n14032), .IN2(n14033), .QN(g20925) );
  NAND2X0 U14884 ( .IN1(n12665), .IN2(n4476), .QN(n14033) );
  INVX0 U14885 ( .INP(n14034), .ZN(n14032) );
  NOR2X0 U14886 ( .IN1(n12665), .IN2(n7853), .QN(n14034) );
  NAND2X0 U14887 ( .IN1(n14035), .IN2(n14036), .QN(g20924) );
  INVX0 U14888 ( .INP(n14037), .ZN(n14036) );
  NOR2X0 U14889 ( .IN1(n13388), .IN2(n8022), .QN(n14037) );
  NAND2X0 U14890 ( .IN1(n13388), .IN2(n13964), .QN(n14035) );
  INVX0 U14891 ( .INP(n8751), .ZN(n13964) );
  NAND3X0 U14892 ( .IN1(n14038), .IN2(n14039), .IN3(n14040), .QN(n8751) );
  NAND2X0 U14893 ( .IN1(g6642), .IN2(g617), .QN(n14040) );
  NAND2X0 U14894 ( .IN1(g6485), .IN2(g614), .QN(n14039) );
  NAND2X0 U14895 ( .IN1(test_so26), .IN2(g550), .QN(n14038) );
  NOR2X0 U14896 ( .IN1(n4309), .IN2(n7748), .QN(n13388) );
  NAND2X0 U14897 ( .IN1(n14041), .IN2(n14042), .QN(g20923) );
  NAND2X0 U14898 ( .IN1(test_so29), .IN2(n12797), .QN(n14042) );
  NAND2X0 U14899 ( .IN1(n4403), .IN2(n12798), .QN(n14041) );
  NAND2X0 U14900 ( .IN1(n14043), .IN2(n14044), .QN(g20922) );
  NAND2X0 U14901 ( .IN1(n12794), .IN2(n4414), .QN(n14044) );
  NAND2X0 U14902 ( .IN1(n8539), .IN2(g709), .QN(n14043) );
  NAND2X0 U14903 ( .IN1(n14045), .IN2(n14046), .QN(g20921) );
  NAND2X0 U14904 ( .IN1(n4422), .IN2(n12731), .QN(n14046) );
  NAND2X0 U14905 ( .IN1(n12729), .IN2(g704), .QN(n14045) );
  NAND2X0 U14906 ( .IN1(n14047), .IN2(n14048), .QN(g20919) );
  NAND2X0 U14907 ( .IN1(n4415), .IN2(n12605), .QN(n14048) );
  NAND2X0 U14908 ( .IN1(n12604), .IN2(g2800), .QN(n14047) );
  NAND2X0 U14909 ( .IN1(n14049), .IN2(n14050), .QN(g20918) );
  NAND2X0 U14910 ( .IN1(n4398), .IN2(n12605), .QN(n14050) );
  INVX0 U14911 ( .INP(n12604), .ZN(n12605) );
  NAND2X0 U14912 ( .IN1(n12604), .IN2(g2773), .QN(n14049) );
  NAND3X0 U14913 ( .IN1(n4426), .IN2(g7425), .IN3(n13979), .QN(n12604) );
  NOR2X0 U14914 ( .IN1(n4490), .IN2(n8039), .QN(n13979) );
  NAND2X0 U14915 ( .IN1(n14051), .IN2(n14052), .QN(g20917) );
  NAND2X0 U14916 ( .IN1(test_so72), .IN2(n9317), .QN(n14052) );
  NAND2X0 U14917 ( .IN1(n4416), .IN2(n12661), .QN(n14051) );
  NAND2X0 U14918 ( .IN1(n14053), .IN2(n14054), .QN(g20916) );
  NAND2X0 U14919 ( .IN1(n12670), .IN2(n4474), .QN(n14054) );
  NAND2X0 U14920 ( .IN1(n12669), .IN2(g2082), .QN(n14053) );
  NAND2X0 U14921 ( .IN1(n14055), .IN2(n14056), .QN(g20915) );
  NAND2X0 U14922 ( .IN1(n4400), .IN2(n12661), .QN(n14056) );
  INVX0 U14923 ( .INP(n9317), .ZN(n12661) );
  NAND2X0 U14924 ( .IN1(n9317), .IN2(g2080), .QN(n14055) );
  NAND3X0 U14925 ( .IN1(n4427), .IN2(g7357), .IN3(n14027), .QN(n9317) );
  NAND2X0 U14926 ( .IN1(n14057), .IN2(n14058), .QN(g20913) );
  NAND2X0 U14927 ( .IN1(n4417), .IN2(n12665), .QN(n14058) );
  INVX0 U14928 ( .INP(n14059), .ZN(n14057) );
  NOR2X0 U14929 ( .IN1(n12665), .IN2(n7845), .QN(n14059) );
  NAND2X0 U14930 ( .IN1(n14060), .IN2(n14061), .QN(g20912) );
  NAND2X0 U14931 ( .IN1(n4421), .IN2(n12738), .QN(n14061) );
  NAND2X0 U14932 ( .IN1(n12737), .IN2(g1391), .QN(n14060) );
  NAND2X0 U14933 ( .IN1(n14062), .IN2(n14063), .QN(g20911) );
  NAND2X0 U14934 ( .IN1(n12726), .IN2(n4476), .QN(n14063) );
  NAND2X0 U14935 ( .IN1(n8518), .IN2(g1389), .QN(n14062) );
  NAND2X0 U14936 ( .IN1(n14064), .IN2(n14065), .QN(g20910) );
  NAND2X0 U14937 ( .IN1(n4402), .IN2(n12665), .QN(n14065) );
  INVX0 U14938 ( .INP(n14066), .ZN(n14064) );
  NOR2X0 U14939 ( .IN1(n12665), .IN2(n7854), .QN(n14066) );
  NOR2X0 U14940 ( .IN1(n14067), .IN2(n8515), .QN(n12665) );
  INVX0 U14941 ( .INP(n14068), .ZN(n14067) );
  NAND2X0 U14942 ( .IN1(n14069), .IN2(n14070), .QN(g20903) );
  NAND2X0 U14943 ( .IN1(n12798), .IN2(n4414), .QN(n14070) );
  NAND2X0 U14944 ( .IN1(n12797), .IN2(g708), .QN(n14069) );
  NAND2X0 U14945 ( .IN1(n14071), .IN2(n14072), .QN(g20902) );
  NAND2X0 U14946 ( .IN1(n4422), .IN2(n12794), .QN(n14072) );
  NAND2X0 U14947 ( .IN1(n8539), .IN2(g706), .QN(n14071) );
  NAND2X0 U14948 ( .IN1(n14073), .IN2(n14074), .QN(g20901) );
  NAND2X0 U14949 ( .IN1(n12731), .IN2(n4478), .QN(n14074) );
  NAND2X0 U14950 ( .IN1(n12729), .IN2(g701), .QN(n14073) );
  NAND2X0 U14951 ( .IN1(n14075), .IN2(n14076), .QN(g20900) );
  NAND2X0 U14952 ( .IN1(n4416), .IN2(n12670), .QN(n14076) );
  NAND2X0 U14953 ( .IN1(n12669), .IN2(g2106), .QN(n14075) );
  NAND2X0 U14954 ( .IN1(n14077), .IN2(n14078), .QN(g20899) );
  NAND2X0 U14955 ( .IN1(n4400), .IN2(n12670), .QN(n14078) );
  INVX0 U14956 ( .INP(n12669), .ZN(n12670) );
  NAND2X0 U14957 ( .IN1(n12669), .IN2(g2079), .QN(n14077) );
  NAND3X0 U14958 ( .IN1(n4427), .IN2(g7229), .IN3(n14027), .QN(n12669) );
  NOR2X0 U14959 ( .IN1(n8094), .IN2(n8038), .QN(n14027) );
  NAND2X0 U14960 ( .IN1(n14079), .IN2(n14080), .QN(g20898) );
  NAND2X0 U14961 ( .IN1(n4417), .IN2(n12726), .QN(n14080) );
  NAND2X0 U14962 ( .IN1(n8518), .IN2(g1413), .QN(n14079) );
  NAND2X0 U14963 ( .IN1(n14081), .IN2(n14082), .QN(g20897) );
  NAND2X0 U14964 ( .IN1(n12738), .IN2(n4476), .QN(n14082) );
  NAND2X0 U14965 ( .IN1(n12737), .IN2(g1388), .QN(n14081) );
  NAND2X0 U14966 ( .IN1(n14083), .IN2(n14084), .QN(g20896) );
  NAND2X0 U14967 ( .IN1(n4402), .IN2(n12726), .QN(n14084) );
  INVX0 U14968 ( .INP(n8518), .ZN(n12726) );
  NAND2X0 U14969 ( .IN1(n8518), .IN2(g1386), .QN(n14083) );
  NAND3X0 U14970 ( .IN1(n4428), .IN2(g7161), .IN3(n14068), .QN(n8518) );
  NAND2X0 U14971 ( .IN1(n14085), .IN2(n14086), .QN(g20894) );
  NAND2X0 U14972 ( .IN1(n4418), .IN2(n12731), .QN(n14086) );
  NAND2X0 U14973 ( .IN1(n12729), .IN2(g725), .QN(n14085) );
  NAND2X0 U14974 ( .IN1(n14087), .IN2(n14088), .QN(g20893) );
  NAND2X0 U14975 ( .IN1(n4422), .IN2(n12798), .QN(n14088) );
  NAND2X0 U14976 ( .IN1(n12797), .IN2(g705), .QN(n14087) );
  NAND2X0 U14977 ( .IN1(n14089), .IN2(n14090), .QN(g20892) );
  NAND2X0 U14978 ( .IN1(n12794), .IN2(n4478), .QN(n14090) );
  NAND2X0 U14979 ( .IN1(n8539), .IN2(g703), .QN(n14089) );
  NAND2X0 U14980 ( .IN1(n14091), .IN2(n14092), .QN(g20891) );
  NAND2X0 U14981 ( .IN1(n4404), .IN2(n12731), .QN(n14092) );
  INVX0 U14982 ( .INP(n12729), .ZN(n12731) );
  NAND2X0 U14983 ( .IN1(n12729), .IN2(g698), .QN(n14091) );
  NAND2X0 U14984 ( .IN1(n14093), .IN2(n8535), .QN(n12729) );
  NOR2X0 U14985 ( .IN1(g3234), .IN2(DFF_1561_n1), .QN(g20884) );
  NAND2X0 U14986 ( .IN1(n14094), .IN2(n14095), .QN(g20883) );
  NAND2X0 U14987 ( .IN1(n4417), .IN2(n12738), .QN(n14095) );
  NAND2X0 U14988 ( .IN1(n12737), .IN2(g1412), .QN(n14094) );
  NAND2X0 U14989 ( .IN1(n14096), .IN2(n14097), .QN(g20882) );
  NAND2X0 U14990 ( .IN1(test_so49), .IN2(n12737), .QN(n14097) );
  NAND2X0 U14991 ( .IN1(n4402), .IN2(n12738), .QN(n14096) );
  INVX0 U14992 ( .INP(n12737), .ZN(n12738) );
  NAND3X0 U14993 ( .IN1(n4428), .IN2(g6979), .IN3(n14068), .QN(n12737) );
  NOR2X0 U14994 ( .IN1(n4489), .IN2(n8037), .QN(n14068) );
  NAND2X0 U14995 ( .IN1(n14098), .IN2(n14099), .QN(g20881) );
  NAND2X0 U14996 ( .IN1(test_so30), .IN2(n8539), .QN(n14099) );
  NAND2X0 U14997 ( .IN1(n4418), .IN2(n12794), .QN(n14098) );
  NAND2X0 U14998 ( .IN1(n14100), .IN2(n14101), .QN(g20880) );
  NAND2X0 U14999 ( .IN1(n12798), .IN2(n4478), .QN(n14101) );
  NAND2X0 U15000 ( .IN1(n12797), .IN2(g702), .QN(n14100) );
  NAND2X0 U15001 ( .IN1(n14102), .IN2(n14103), .QN(g20879) );
  NAND2X0 U15002 ( .IN1(n4404), .IN2(n12794), .QN(n14103) );
  INVX0 U15003 ( .INP(n8539), .ZN(n12794) );
  NAND2X0 U15004 ( .IN1(n8539), .IN2(g700), .QN(n14102) );
  NAND3X0 U15005 ( .IN1(n4429), .IN2(g6911), .IN3(n14093), .QN(n8539) );
  NAND2X0 U15006 ( .IN1(n14104), .IN2(n14105), .QN(g20876) );
  NAND2X0 U15007 ( .IN1(n4418), .IN2(n12798), .QN(n14105) );
  NAND2X0 U15008 ( .IN1(n12797), .IN2(g726), .QN(n14104) );
  NAND2X0 U15009 ( .IN1(n14106), .IN2(n14107), .QN(g20875) );
  NAND2X0 U15010 ( .IN1(n4404), .IN2(n12798), .QN(n14107) );
  INVX0 U15011 ( .INP(n12797), .ZN(n12798) );
  NAND2X0 U15012 ( .IN1(n12797), .IN2(g699), .QN(n14106) );
  NAND3X0 U15013 ( .IN1(n4429), .IN2(g6677), .IN3(n14093), .QN(n12797) );
  NOR2X0 U15014 ( .IN1(n4492), .IN2(n8036), .QN(n14093) );
  NAND2X0 U15015 ( .IN1(n14108), .IN2(n14109), .QN(g20874) );
  NAND2X0 U15016 ( .IN1(g2879), .IN2(g8096), .QN(n14109) );
  NAND2X0 U15017 ( .IN1(n4351), .IN2(n13751), .QN(n14108) );
  XOR2X1 U15018 ( .IN1(n8550), .IN2(n13754), .Q(n13751) );
  NOR2X0 U15019 ( .IN1(g3231), .IN2(n14352), .QN(n13754) );
  XOR3X1 U15020 ( .IN1(n14110), .IN2(n14111), .IN3(n14112), .Q(n8550) );
  XOR3X1 U15021 ( .IN1(n7991), .IN2(n7990), .IN3(n14113), .Q(n14112) );
  XOR2X1 U15022 ( .IN1(g2944), .IN2(n7993), .Q(n14113) );
  XOR2X1 U15023 ( .IN1(n7981), .IN2(n7977), .Q(n14111) );
  XOR2X1 U15024 ( .IN1(n7989), .IN2(n7982), .Q(n14110) );
  NOR2X0 U15025 ( .IN1(n11303), .IN2(n14114), .QN(g20789) );
  XOR2X1 U15026 ( .IN1(n4398), .IN2(n9297), .Q(n14114) );
  NOR2X0 U15027 ( .IN1(g2733), .IN2(n4292), .QN(n9297) );
  INVX0 U15028 ( .INP(n9289), .ZN(n11303) );
  NAND2X0 U15029 ( .IN1(g7487), .IN2(g2704), .QN(n9289) );
  NOR2X0 U15030 ( .IN1(n9305), .IN2(n14115), .QN(g20752) );
  XOR2X1 U15031 ( .IN1(n4400), .IN2(n9314), .Q(n14115) );
  NOR2X0 U15032 ( .IN1(g2039), .IN2(n4293), .QN(n9314) );
  NOR2X0 U15033 ( .IN1(n4357), .IN2(n7746), .QN(n9305) );
  NOR2X0 U15034 ( .IN1(n8512), .IN2(n14116), .QN(g20717) );
  XNOR2X1 U15035 ( .IN1(n4402), .IN2(n8515), .Q(n14116) );
  NAND2X0 U15036 ( .IN1(n4428), .IN2(g1315), .QN(n8515) );
  NOR2X0 U15037 ( .IN1(n4358), .IN2(n7747), .QN(n8512) );
  NOR2X0 U15038 ( .IN1(n8536), .IN2(n14117), .QN(g20682) );
  XOR2X1 U15039 ( .IN1(n4404), .IN2(n8535), .Q(n14117) );
  NOR2X0 U15040 ( .IN1(g659), .IN2(n4295), .QN(n8535) );
  NOR2X0 U15041 ( .IN1(n4359), .IN2(n7748), .QN(n8536) );
  NAND2X0 U15042 ( .IN1(n14118), .IN2(n14119), .QN(g20417) );
  NAND2X0 U15043 ( .IN1(n4351), .IN2(g2963), .QN(n14119) );
  NAND2X0 U15044 ( .IN1(g2879), .IN2(g7334), .QN(n14118) );
  NAND2X0 U15045 ( .IN1(n14120), .IN2(n14121), .QN(g20376) );
  NAND2X0 U15046 ( .IN1(test_so2), .IN2(n4351), .QN(n14121) );
  NAND2X0 U15047 ( .IN1(g2879), .IN2(g6895), .QN(n14120) );
  NAND2X0 U15048 ( .IN1(n14122), .IN2(n14123), .QN(g20375) );
  NAND2X0 U15049 ( .IN1(n4292), .IN2(g2733), .QN(n14123) );
  NAND2X0 U15050 ( .IN1(n14124), .IN2(g2703), .QN(n14122) );
  NAND2X0 U15051 ( .IN1(n14125), .IN2(n14126), .QN(g20353) );
  NAND2X0 U15052 ( .IN1(n4293), .IN2(g2039), .QN(n14126) );
  NAND2X0 U15053 ( .IN1(n14124), .IN2(g2009), .QN(n14125) );
  NAND2X0 U15054 ( .IN1(n14127), .IN2(n14128), .QN(g20343) );
  NAND2X0 U15055 ( .IN1(n4351), .IN2(g2969), .QN(n14128) );
  NAND2X0 U15056 ( .IN1(g2879), .IN2(g6442), .QN(n14127) );
  NAND2X0 U15057 ( .IN1(n14129), .IN2(n14130), .QN(g20333) );
  NAND2X0 U15058 ( .IN1(n4294), .IN2(g1345), .QN(n14130) );
  NAND2X0 U15059 ( .IN1(n14124), .IN2(g1315), .QN(n14129) );
  NAND2X0 U15060 ( .IN1(n14131), .IN2(n14132), .QN(g20314) );
  NAND2X0 U15061 ( .IN1(n4295), .IN2(g659), .QN(n14132) );
  NAND2X0 U15062 ( .IN1(n14124), .IN2(g629), .QN(n14131) );
  INVX0 U15063 ( .INP(n13344), .ZN(n14124) );
  NAND4X0 U15064 ( .IN1(n8051), .IN2(n8034), .IN3(n14133), .IN4(n8033), .QN(
        n13344) );
  NOR2X0 U15065 ( .IN1(test_so98), .IN2(g3006), .QN(n14133) );
  NAND2X0 U15066 ( .IN1(n14134), .IN2(n14135), .QN(g20310) );
  NAND2X0 U15067 ( .IN1(n4351), .IN2(g2972), .QN(n14135) );
  NAND2X0 U15068 ( .IN1(g2879), .IN2(g6225), .QN(n14134) );
  NAND2X0 U15069 ( .IN1(n14136), .IN2(n14137), .QN(g19184) );
  NAND2X0 U15070 ( .IN1(n4351), .IN2(g2975), .QN(n14137) );
  NAND2X0 U15071 ( .IN1(g2879), .IN2(g4590), .QN(n14136) );
  NAND2X0 U15072 ( .IN1(n14138), .IN2(n14139), .QN(g19178) );
  NAND2X0 U15073 ( .IN1(n4351), .IN2(g2935), .QN(n14139) );
  NAND2X0 U15074 ( .IN1(test_so5), .IN2(g2879), .QN(n14138) );
  NAND2X0 U15075 ( .IN1(n14140), .IN2(n14141), .QN(g19173) );
  NAND2X0 U15076 ( .IN1(n4351), .IN2(g2978), .QN(n14141) );
  NAND2X0 U15077 ( .IN1(g2879), .IN2(g4323), .QN(n14140) );
  NAND2X0 U15078 ( .IN1(n14142), .IN2(n14143), .QN(g19172) );
  NAND2X0 U15079 ( .IN1(n4351), .IN2(g2953), .QN(n14143) );
  NAND2X0 U15080 ( .IN1(g2879), .IN2(g4321), .QN(n14142) );
  NAND2X0 U15081 ( .IN1(n14144), .IN2(n14145), .QN(g19167) );
  NAND2X0 U15082 ( .IN1(n4351), .IN2(g2938), .QN(n14145) );
  NAND2X0 U15083 ( .IN1(g2879), .IN2(g4200), .QN(n14144) );
  NAND2X0 U15084 ( .IN1(n14146), .IN2(n14147), .QN(g19163) );
  NAND2X0 U15085 ( .IN1(n4351), .IN2(g2981), .QN(n14147) );
  NAND2X0 U15086 ( .IN1(g2879), .IN2(g4090), .QN(n14146) );
  NAND2X0 U15087 ( .IN1(n14148), .IN2(n14149), .QN(g19162) );
  NAND2X0 U15088 ( .IN1(n4351), .IN2(g2956), .QN(n14149) );
  NAND2X0 U15089 ( .IN1(g2879), .IN2(g4088), .QN(n14148) );
  NAND2X0 U15090 ( .IN1(n14150), .IN2(n14151), .QN(g19157) );
  NAND2X0 U15091 ( .IN1(n4351), .IN2(g2941), .QN(n14151) );
  NAND2X0 U15092 ( .IN1(g2879), .IN2(g3993), .QN(n14150) );
  NAND2X0 U15093 ( .IN1(n14152), .IN2(n14153), .QN(g19154) );
  NAND2X0 U15094 ( .IN1(n4351), .IN2(g2874), .QN(n14153) );
  NAND2X0 U15095 ( .IN1(test_so3), .IN2(g2879), .QN(n14152) );
  NAND2X0 U15096 ( .IN1(n14154), .IN2(n14155), .QN(g19153) );
  NAND2X0 U15097 ( .IN1(n4351), .IN2(g2959), .QN(n14155) );
  NAND2X0 U15098 ( .IN1(g2879), .IN2(g8249), .QN(n14154) );
  NAND2X0 U15099 ( .IN1(n14156), .IN2(n14157), .QN(g19149) );
  NAND2X0 U15100 ( .IN1(n4351), .IN2(g2944), .QN(n14157) );
  NAND2X0 U15101 ( .IN1(g2879), .IN2(g8175), .QN(n14156) );
  NAND2X0 U15102 ( .IN1(n14158), .IN2(n14159), .QN(g19144) );
  NAND2X0 U15103 ( .IN1(n4351), .IN2(g2947), .QN(n14159) );
  NAND2X0 U15104 ( .IN1(g2879), .IN2(g8023), .QN(n14158) );
  NAND2X0 U15105 ( .IN1(n14160), .IN2(n14161), .QN(g18975) );
  NAND2X0 U15106 ( .IN1(n4351), .IN2(g2195), .QN(n14161) );
  NAND2X0 U15107 ( .IN1(g2879), .IN2(g2981), .QN(n14160) );
  NAND2X0 U15108 ( .IN1(n14162), .IN2(n14163), .QN(g18968) );
  NAND2X0 U15109 ( .IN1(n4351), .IN2(g2190), .QN(n14163) );
  NAND2X0 U15110 ( .IN1(g2879), .IN2(g2978), .QN(n14162) );
  NAND2X0 U15111 ( .IN1(n14164), .IN2(n14165), .QN(g18957) );
  NAND2X0 U15112 ( .IN1(n4351), .IN2(g2165), .QN(n14165) );
  NAND2X0 U15113 ( .IN1(g2879), .IN2(g2963), .QN(n14164) );
  NAND2X0 U15114 ( .IN1(n14166), .IN2(n14167), .QN(g18942) );
  NAND2X0 U15115 ( .IN1(g2879), .IN2(g2975), .QN(n14167) );
  NAND2X0 U15116 ( .IN1(n4351), .IN2(g2185), .QN(n14166) );
  NAND2X0 U15117 ( .IN1(n14168), .IN2(n14169), .QN(g18907) );
  NAND2X0 U15118 ( .IN1(n4365), .IN2(g3061), .QN(n14169) );
  NAND2X0 U15119 ( .IN1(g2987), .IN2(g2997), .QN(n14168) );
  NAND2X0 U15120 ( .IN1(n14170), .IN2(n14171), .QN(g18906) );
  NAND2X0 U15121 ( .IN1(n4351), .IN2(g2180), .QN(n14171) );
  NAND2X0 U15122 ( .IN1(g2879), .IN2(g2972), .QN(n14170) );
  NAND2X0 U15123 ( .IN1(n14172), .IN2(n14173), .QN(g18885) );
  NAND2X0 U15124 ( .IN1(g2879), .IN2(g2874), .QN(n14173) );
  NAND2X0 U15125 ( .IN1(n4351), .IN2(g2200), .QN(n14172) );
  NAND2X0 U15126 ( .IN1(n14174), .IN2(n14175), .QN(g18883) );
  NAND2X0 U15127 ( .IN1(n4351), .IN2(g1471), .QN(n14175) );
  NAND2X0 U15128 ( .IN1(g2879), .IN2(g2935), .QN(n14174) );
  NAND2X0 U15129 ( .IN1(n14176), .IN2(n14177), .QN(g18868) );
  NAND2X0 U15130 ( .IN1(n4365), .IN2(g3060), .QN(n14177) );
  NAND2X0 U15131 ( .IN1(g2987), .IN2(g3078), .QN(n14176) );
  NAND2X0 U15132 ( .IN1(n14178), .IN2(n14179), .QN(g18867) );
  NAND2X0 U15133 ( .IN1(g2879), .IN2(g2969), .QN(n14179) );
  NAND2X0 U15134 ( .IN1(n4351), .IN2(g2175), .QN(n14178) );
  NAND2X0 U15135 ( .IN1(n14180), .IN2(n14181), .QN(g18866) );
  NAND2X0 U15136 ( .IN1(n4351), .IN2(g1476), .QN(n14181) );
  NAND2X0 U15137 ( .IN1(g2879), .IN2(g2938), .QN(n14180) );
  NAND2X0 U15138 ( .IN1(n14182), .IN2(n14183), .QN(g18852) );
  NAND2X0 U15139 ( .IN1(g2879), .IN2(g2941), .QN(n14183) );
  NAND2X0 U15140 ( .IN1(n4351), .IN2(g1481), .QN(n14182) );
  NAND2X0 U15141 ( .IN1(n14184), .IN2(n14185), .QN(g18837) );
  NAND2X0 U15142 ( .IN1(n4365), .IN2(g3059), .QN(n14185) );
  NAND2X0 U15143 ( .IN1(g2987), .IN2(g3077), .QN(n14184) );
  NAND2X0 U15144 ( .IN1(n14186), .IN2(n14187), .QN(g18836) );
  NAND2X0 U15145 ( .IN1(n4351), .IN2(g2170), .QN(n14187) );
  NAND2X0 U15146 ( .IN1(test_so2), .IN2(g2879), .QN(n14186) );
  NAND2X0 U15147 ( .IN1(n14188), .IN2(n14189), .QN(g18835) );
  NAND2X0 U15148 ( .IN1(n4351), .IN2(g1486), .QN(n14189) );
  NAND2X0 U15149 ( .IN1(g2879), .IN2(g2944), .QN(n14188) );
  NAND2X0 U15150 ( .IN1(n14190), .IN2(n14191), .QN(g18821) );
  NAND2X0 U15151 ( .IN1(g2879), .IN2(g2947), .QN(n14191) );
  NAND2X0 U15152 ( .IN1(n4351), .IN2(g1491), .QN(n14190) );
  NAND2X0 U15153 ( .IN1(n14192), .IN2(n14193), .QN(g18820) );
  NAND2X0 U15154 ( .IN1(n4299), .IN2(g2584), .QN(n14193) );
  NAND2X0 U15155 ( .IN1(g2624), .IN2(g2631), .QN(n14192) );
  NAND2X0 U15156 ( .IN1(n14194), .IN2(n14195), .QN(g18804) );
  NAND2X0 U15157 ( .IN1(n4365), .IN2(g3058), .QN(n14195) );
  NAND2X0 U15158 ( .IN1(g2987), .IN2(g3076), .QN(n14194) );
  NAND2X0 U15159 ( .IN1(n14196), .IN2(n14197), .QN(g18803) );
  NAND2X0 U15160 ( .IN1(n4351), .IN2(g1496), .QN(n14197) );
  NAND2X0 U15161 ( .IN1(g2879), .IN2(g2953), .QN(n14196) );
  NAND2X0 U15162 ( .IN1(n14198), .IN2(n14199), .QN(g18794) );
  NAND2X0 U15163 ( .IN1(g1937), .IN2(g1930), .QN(n14199) );
  NAND2X0 U15164 ( .IN1(n4366), .IN2(g1890), .QN(n14198) );
  NAND2X0 U15165 ( .IN1(n14200), .IN2(n14201), .QN(g18782) );
  NAND2X0 U15166 ( .IN1(g3109), .IN2(g559), .QN(n14201) );
  NAND2X0 U15167 ( .IN1(n4494), .IN2(g3084), .QN(n14200) );
  NAND2X0 U15168 ( .IN1(n14202), .IN2(n14203), .QN(g18781) );
  NAND2X0 U15169 ( .IN1(n4351), .IN2(g1501), .QN(n14203) );
  NAND2X0 U15170 ( .IN1(g2879), .IN2(g2956), .QN(n14202) );
  NAND2X0 U15171 ( .IN1(n14204), .IN2(n14205), .QN(g18780) );
  NAND2X0 U15172 ( .IN1(n4299), .IN2(g2631), .QN(n14205) );
  NAND2X0 U15173 ( .IN1(n7961), .IN2(g2624), .QN(n14204) );
  NAND2X0 U15174 ( .IN1(n14206), .IN2(n14207), .QN(g18763) );
  NAND2X0 U15175 ( .IN1(n4300), .IN2(g1196), .QN(n14207) );
  NAND2X0 U15176 ( .IN1(g1236), .IN2(g1243), .QN(n14206) );
  NAND2X0 U15177 ( .IN1(n14208), .IN2(n14209), .QN(g18755) );
  NAND2X0 U15178 ( .IN1(n4365), .IN2(g3057), .QN(n14209) );
  NAND2X0 U15179 ( .IN1(g2987), .IN2(g3075), .QN(n14208) );
  NAND2X0 U15180 ( .IN1(n14210), .IN2(n14211), .QN(g18754) );
  NAND2X0 U15181 ( .IN1(g2879), .IN2(g2959), .QN(n14211) );
  NAND2X0 U15182 ( .IN1(n4351), .IN2(g1506), .QN(n14210) );
  NAND2X0 U15183 ( .IN1(n14212), .IN2(n14213), .QN(g18743) );
  NAND2X0 U15184 ( .IN1(n7969), .IN2(g1930), .QN(n14213) );
  NAND2X0 U15185 ( .IN1(n4366), .IN2(g1937), .QN(n14212) );
  NAND2X0 U15186 ( .IN1(n14214), .IN2(n14215), .QN(g18726) );
  NAND2X0 U15187 ( .IN1(test_so22), .IN2(n4313), .QN(n14215) );
  NAND2X0 U15188 ( .IN1(g550), .IN2(g557), .QN(n14214) );
  NAND2X0 U15189 ( .IN1(n14216), .IN2(n14217), .QN(g18719) );
  NAND2X0 U15190 ( .IN1(n4383), .IN2(g3211), .QN(n14217) );
  NAND2X0 U15191 ( .IN1(g8030), .IN2(g559), .QN(n14216) );
  NAND2X0 U15192 ( .IN1(n14218), .IN2(n14219), .QN(g18707) );
  NAND2X0 U15193 ( .IN1(n4300), .IN2(g1243), .QN(n14219) );
  NAND2X0 U15194 ( .IN1(n7970), .IN2(g1236), .QN(n14218) );
  NAND2X0 U15195 ( .IN1(n14220), .IN2(n14221), .QN(g18678) );
  NAND2X0 U15196 ( .IN1(n4313), .IN2(g557), .QN(n14221) );
  NAND2X0 U15197 ( .IN1(n7972), .IN2(g550), .QN(n14220) );
  NAND2X0 U15198 ( .IN1(n14222), .IN2(n14223), .QN(g18669) );
  NAND2X0 U15199 ( .IN1(n4382), .IN2(test_so6), .QN(n14223) );
  NAND2X0 U15200 ( .IN1(g8106), .IN2(g559), .QN(n14222) );
  NAND2X0 U15201 ( .IN1(n14224), .IN2(n14225), .QN(g17429) );
  NAND2X0 U15202 ( .IN1(g3109), .IN2(g2574), .QN(n14225) );
  NAND2X0 U15203 ( .IN1(n4494), .IN2(g3088), .QN(n14224) );
  NAND2X0 U15204 ( .IN1(n14226), .IN2(n14227), .QN(g17383) );
  NAND2X0 U15205 ( .IN1(n4494), .IN2(test_so8), .QN(n14227) );
  NAND2X0 U15206 ( .IN1(g3109), .IN2(g1880), .QN(n14226) );
  NAND2X0 U15207 ( .IN1(n14228), .IN2(n14229), .QN(g17341) );
  NAND2X0 U15208 ( .IN1(n4383), .IN2(g3185), .QN(n14229) );
  NAND2X0 U15209 ( .IN1(g8030), .IN2(g2574), .QN(n14228) );
  NAND2X0 U15210 ( .IN1(n14230), .IN2(n14231), .QN(g17340) );
  NAND2X0 U15211 ( .IN1(g3109), .IN2(g1186), .QN(n14231) );
  NAND2X0 U15212 ( .IN1(n4494), .IN2(g3170), .QN(n14230) );
  NAND2X0 U15213 ( .IN1(n14232), .IN2(n14233), .QN(g17303) );
  NAND2X0 U15214 ( .IN1(n4383), .IN2(g3176), .QN(n14233) );
  NAND2X0 U15215 ( .IN1(g8030), .IN2(g1880), .QN(n14232) );
  NAND2X0 U15216 ( .IN1(n14234), .IN2(n14235), .QN(g17302) );
  NAND2X0 U15217 ( .IN1(g3109), .IN2(g499), .QN(n14235) );
  NAND2X0 U15218 ( .IN1(n4494), .IN2(g3161), .QN(n14234) );
  NAND2X0 U15219 ( .IN1(n14236), .IN2(n14237), .QN(g17271) );
  NAND2X0 U15220 ( .IN1(n4382), .IN2(g3182), .QN(n14237) );
  NAND2X0 U15221 ( .IN1(g8106), .IN2(g2574), .QN(n14236) );
  NAND2X0 U15222 ( .IN1(n14238), .IN2(n14239), .QN(g17270) );
  NAND2X0 U15223 ( .IN1(g8030), .IN2(g1186), .QN(n14239) );
  NAND2X0 U15224 ( .IN1(n4383), .IN2(g3167), .QN(n14238) );
  NAND2X0 U15225 ( .IN1(n14240), .IN2(n14241), .QN(g17269) );
  NAND2X0 U15226 ( .IN1(g3109), .IN2(g2633), .QN(n14241) );
  NAND2X0 U15227 ( .IN1(n4494), .IN2(g3096), .QN(n14240) );
  NAND2X0 U15228 ( .IN1(n14242), .IN2(n14243), .QN(g17248) );
  NAND2X0 U15229 ( .IN1(g8106), .IN2(g1880), .QN(n14243) );
  NAND2X0 U15230 ( .IN1(n4382), .IN2(g3173), .QN(n14242) );
  NAND2X0 U15231 ( .IN1(n14244), .IN2(n14245), .QN(g17247) );
  NAND2X0 U15232 ( .IN1(n4383), .IN2(g3158), .QN(n14245) );
  NAND2X0 U15233 ( .IN1(g8030), .IN2(g499), .QN(n14244) );
  NAND2X0 U15234 ( .IN1(n14246), .IN2(n14247), .QN(g17246) );
  NAND2X0 U15235 ( .IN1(g3109), .IN2(g1939), .QN(n14247) );
  NAND2X0 U15236 ( .IN1(n4494), .IN2(g3093), .QN(n14246) );
  NAND2X0 U15237 ( .IN1(n14248), .IN2(n14249), .QN(g17236) );
  NAND2X0 U15238 ( .IN1(g8106), .IN2(g1186), .QN(n14249) );
  NAND2X0 U15239 ( .IN1(n4382), .IN2(g3164), .QN(n14248) );
  NAND2X0 U15240 ( .IN1(n14250), .IN2(n14251), .QN(g17235) );
  NAND2X0 U15241 ( .IN1(n4383), .IN2(g3095), .QN(n14251) );
  NAND2X0 U15242 ( .IN1(g8030), .IN2(g2633), .QN(n14250) );
  NAND2X0 U15243 ( .IN1(n14252), .IN2(n14253), .QN(g17234) );
  NAND2X0 U15244 ( .IN1(g3109), .IN2(g1245), .QN(n14253) );
  NAND2X0 U15245 ( .IN1(n4494), .IN2(g3087), .QN(n14252) );
  NAND2X0 U15246 ( .IN1(n14254), .IN2(n14255), .QN(g17229) );
  NAND2X0 U15247 ( .IN1(n4382), .IN2(g3155), .QN(n14255) );
  NAND2X0 U15248 ( .IN1(g8106), .IN2(g499), .QN(n14254) );
  NAND2X0 U15249 ( .IN1(n14256), .IN2(n14257), .QN(g17228) );
  NAND2X0 U15250 ( .IN1(n4383), .IN2(g3092), .QN(n14257) );
  NAND2X0 U15251 ( .IN1(g8030), .IN2(g1939), .QN(n14256) );
  NAND2X0 U15252 ( .IN1(n14258), .IN2(n14259), .QN(g17226) );
  NAND2X0 U15253 ( .IN1(n4382), .IN2(g3094), .QN(n14259) );
  NAND2X0 U15254 ( .IN1(g8106), .IN2(g2633), .QN(n14258) );
  NAND2X0 U15255 ( .IN1(n14260), .IN2(n14261), .QN(g17225) );
  NAND2X0 U15256 ( .IN1(g8030), .IN2(g1245), .QN(n14261) );
  NAND2X0 U15257 ( .IN1(n4383), .IN2(g3086), .QN(n14260) );
  NAND2X0 U15258 ( .IN1(n14262), .IN2(n14263), .QN(g17224) );
  NAND2X0 U15259 ( .IN1(n4382), .IN2(g3091), .QN(n14263) );
  NAND2X0 U15260 ( .IN1(g8106), .IN2(g1939), .QN(n14262) );
  NAND2X0 U15261 ( .IN1(n14264), .IN2(n14265), .QN(g17222) );
  NAND2X0 U15262 ( .IN1(g8106), .IN2(g1245), .QN(n14265) );
  NAND2X0 U15263 ( .IN1(n4382), .IN2(g3085), .QN(n14264) );
  NAND2X0 U15264 ( .IN1(n14266), .IN2(n14267), .QN(g16880) );
  NAND2X0 U15265 ( .IN1(n4365), .IN2(g3056), .QN(n14267) );
  NAND2X0 U15266 ( .IN1(g2987), .IN2(g3074), .QN(n14266) );
  NAND2X0 U15267 ( .IN1(n14268), .IN2(n14269), .QN(g16866) );
  NAND2X0 U15268 ( .IN1(n4365), .IN2(g3051), .QN(n14269) );
  NAND2X0 U15269 ( .IN1(test_so97), .IN2(g2987), .QN(n14268) );
  NAND2X0 U15270 ( .IN1(n14270), .IN2(n14271), .QN(g16861) );
  NAND2X0 U15271 ( .IN1(test_so96), .IN2(n4365), .QN(n14271) );
  NAND2X0 U15272 ( .IN1(g2987), .IN2(g3073), .QN(n14270) );
  NAND2X0 U15273 ( .IN1(n14272), .IN2(n14273), .QN(g16860) );
  NAND2X0 U15274 ( .IN1(n4365), .IN2(g3046), .QN(n14273) );
  NAND2X0 U15275 ( .IN1(g2987), .IN2(g3065), .QN(n14272) );
  NAND2X0 U15276 ( .IN1(n14274), .IN2(n14275), .QN(g16857) );
  NAND2X0 U15277 ( .IN1(n4365), .IN2(g3050), .QN(n14275) );
  NAND2X0 U15278 ( .IN1(g2987), .IN2(g3069), .QN(n14274) );
  NAND2X0 U15279 ( .IN1(n14276), .IN2(n14277), .QN(g16854) );
  NAND2X0 U15280 ( .IN1(n4365), .IN2(g3053), .QN(n14277) );
  NAND2X0 U15281 ( .IN1(g2987), .IN2(g3072), .QN(n14276) );
  NAND2X0 U15282 ( .IN1(n14278), .IN2(n14279), .QN(g16853) );
  NAND2X0 U15283 ( .IN1(n4365), .IN2(g3045), .QN(n14279) );
  NAND2X0 U15284 ( .IN1(g2987), .IN2(g3064), .QN(n14278) );
  NAND2X0 U15285 ( .IN1(n14280), .IN2(n14281), .QN(g16851) );
  NAND2X0 U15286 ( .IN1(n4365), .IN2(g3049), .QN(n14281) );
  NAND2X0 U15287 ( .IN1(g2987), .IN2(g3068), .QN(n14280) );
  NAND2X0 U15288 ( .IN1(n14282), .IN2(n14283), .QN(g16845) );
  NAND2X0 U15289 ( .IN1(n4365), .IN2(g3052), .QN(n14283) );
  NAND2X0 U15290 ( .IN1(g2987), .IN2(g3071), .QN(n14282) );
  NAND2X0 U15291 ( .IN1(n14284), .IN2(n14285), .QN(g16844) );
  NAND2X0 U15292 ( .IN1(n4365), .IN2(g3044), .QN(n14285) );
  NAND2X0 U15293 ( .IN1(g2987), .IN2(g3063), .QN(n14284) );
  NAND2X0 U15294 ( .IN1(n14286), .IN2(n14287), .QN(g16835) );
  NAND2X0 U15295 ( .IN1(n4365), .IN2(g3048), .QN(n14287) );
  NAND2X0 U15296 ( .IN1(g2987), .IN2(g3067), .QN(n14286) );
  NAND2X0 U15297 ( .IN1(n14288), .IN2(n14289), .QN(g16824) );
  NAND2X0 U15298 ( .IN1(n4365), .IN2(g3043), .QN(n14289) );
  NAND2X0 U15299 ( .IN1(g2987), .IN2(g3062), .QN(n14288) );
  NOR2X0 U15300 ( .IN1(g51), .IN2(DFF_1_n1), .QN(g16823) );
  NAND2X0 U15301 ( .IN1(n14290), .IN2(n14291), .QN(g16803) );
  NAND2X0 U15302 ( .IN1(n4365), .IN2(g3047), .QN(n14291) );
  NAND2X0 U15303 ( .IN1(g2987), .IN2(g3066), .QN(n14290) );
  NOR2X0 U15304 ( .IN1(n4423), .IN2(g51), .QN(g16802) );
  NAND2X0 U15305 ( .IN1(n14292), .IN2(n14293), .QN(g16718) );
  NAND2X0 U15306 ( .IN1(n4292), .IN2(g2704), .QN(n14293) );
  NAND2X0 U15307 ( .IN1(g2703), .IN2(g2584), .QN(n14292) );
  NAND2X0 U15308 ( .IN1(n14294), .IN2(n14295), .QN(g16692) );
  NAND2X0 U15309 ( .IN1(n4293), .IN2(g2010), .QN(n14295) );
  NAND2X0 U15310 ( .IN1(g2009), .IN2(g1890), .QN(n14294) );
  NAND2X0 U15311 ( .IN1(n14296), .IN2(n14297), .QN(g16671) );
  NAND2X0 U15312 ( .IN1(n4294), .IN2(g1316), .QN(n14297) );
  NAND2X0 U15313 ( .IN1(g1315), .IN2(g1196), .QN(n14296) );
  NAND2X0 U15314 ( .IN1(n14298), .IN2(n14299), .QN(g16654) );
  NAND2X0 U15315 ( .IN1(n4295), .IN2(g630), .QN(n14299) );
  NAND2X0 U15316 ( .IN1(test_so22), .IN2(g629), .QN(n14298) );
  NAND2X0 U15317 ( .IN1(n14300), .IN2(g2987), .QN(g16496) );
  NAND2X0 U15318 ( .IN1(DFF_1612_n1), .IN2(g5388), .QN(n14300) );
  NOR3X0 U15319 ( .IN1(n14301), .IN2(n14302), .IN3(n14303), .QN(g13194) );
  NOR2X0 U15320 ( .IN1(n4314), .IN2(test_so87), .QN(n14303) );
  NOR2X0 U15321 ( .IN1(n4370), .IN2(g2561), .QN(n14302) );
  NOR2X0 U15322 ( .IN1(n4299), .IN2(g2562), .QN(n14301) );
  NOR3X0 U15323 ( .IN1(n14304), .IN2(n14305), .IN3(n14306), .QN(g13182) );
  NOR2X0 U15324 ( .IN1(n4366), .IN2(g1868), .QN(n14306) );
  NOR2X0 U15325 ( .IN1(n4296), .IN2(g1869), .QN(n14305) );
  NOR2X0 U15326 ( .IN1(n4315), .IN2(g1867), .QN(n14304) );
  NOR3X0 U15327 ( .IN1(n14307), .IN2(n14308), .IN3(n14309), .QN(g13175) );
  NOR2X0 U15328 ( .IN1(n4299), .IN2(g2553), .QN(n14309) );
  NOR2X0 U15329 ( .IN1(n4314), .IN2(g2554), .QN(n14308) );
  NOR2X0 U15330 ( .IN1(n4370), .IN2(g2552), .QN(n14307) );
  NOR3X0 U15331 ( .IN1(n14310), .IN2(n14311), .IN3(n14312), .QN(g13171) );
  NOR2X0 U15332 ( .IN1(n4300), .IN2(test_so44), .QN(n14312) );
  NOR2X0 U15333 ( .IN1(n4316), .IN2(g1173), .QN(n14311) );
  NOR2X0 U15334 ( .IN1(n4371), .IN2(g1175), .QN(n14310) );
  NOR3X0 U15335 ( .IN1(n14313), .IN2(n14314), .IN3(n14315), .QN(g13164) );
  NOR2X0 U15336 ( .IN1(n4366), .IN2(g1859), .QN(n14315) );
  NOR2X0 U15337 ( .IN1(n4296), .IN2(g1860), .QN(n14314) );
  NOR2X0 U15338 ( .IN1(n4315), .IN2(g1858), .QN(n14313) );
  NOR3X0 U15339 ( .IN1(n14316), .IN2(n14317), .IN3(n14318), .QN(g13160) );
  NOR2X0 U15340 ( .IN1(n4313), .IN2(g487), .QN(n14318) );
  NOR2X0 U15341 ( .IN1(n4298), .IN2(g488), .QN(n14317) );
  NOR2X0 U15342 ( .IN1(n4372), .IN2(g486), .QN(n14316) );
  NOR3X0 U15343 ( .IN1(n14319), .IN2(n14320), .IN3(n14321), .QN(g13155) );
  NOR2X0 U15344 ( .IN1(n4300), .IN2(g1165), .QN(n14321) );
  NOR2X0 U15345 ( .IN1(n4371), .IN2(g1166), .QN(n14320) );
  NOR2X0 U15346 ( .IN1(n4316), .IN2(g1164), .QN(n14319) );
  NOR3X0 U15347 ( .IN1(n14322), .IN2(n14323), .IN3(n14324), .QN(g13149) );
  NOR2X0 U15348 ( .IN1(n4313), .IN2(g478), .QN(n14324) );
  NOR2X0 U15349 ( .IN1(n4298), .IN2(g479), .QN(n14323) );
  NOR2X0 U15350 ( .IN1(n4372), .IN2(g477), .QN(n14322) );
  NOR3X0 U15351 ( .IN1(n14325), .IN2(n14326), .IN3(n14327), .QN(g13143) );
  NOR2X0 U15352 ( .IN1(n4299), .IN2(g2559), .QN(n14327) );
  NOR2X0 U15353 ( .IN1(n4314), .IN2(g2539), .QN(n14326) );
  NOR2X0 U15354 ( .IN1(n4370), .IN2(g2555), .QN(n14325) );
  NOR3X0 U15355 ( .IN1(n14328), .IN2(n14329), .IN3(n14330), .QN(g13135) );
  NOR2X0 U15356 ( .IN1(n4366), .IN2(g1865), .QN(n14330) );
  NOR2X0 U15357 ( .IN1(n4296), .IN2(g1845), .QN(n14329) );
  NOR2X0 U15358 ( .IN1(n4315), .IN2(g1861), .QN(n14328) );
  NOR3X0 U15359 ( .IN1(n14331), .IN2(n14332), .IN3(n14333), .QN(g13124) );
  NOR2X0 U15360 ( .IN1(n4300), .IN2(g1171), .QN(n14333) );
  NOR2X0 U15361 ( .IN1(n4371), .IN2(g1151), .QN(n14332) );
  NOR2X0 U15362 ( .IN1(n4316), .IN2(g1167), .QN(n14331) );
  NOR3X0 U15363 ( .IN1(n14334), .IN2(n14335), .IN3(n14336), .QN(g13111) );
  NOR2X0 U15364 ( .IN1(n4313), .IN2(g484), .QN(n14336) );
  NOR2X0 U15365 ( .IN1(n4298), .IN2(g464), .QN(n14335) );
  NOR2X0 U15366 ( .IN1(n4372), .IN2(g480), .QN(n14334) );
  XOR2X1 U15367 ( .IN1(n8013), .IN2(n8730), .Q(N995) );
  XNOR3X1 U15368 ( .IN1(n14337), .IN2(n14338), .IN3(n14339), .Q(n8730) );
  XOR3X1 U15369 ( .IN1(n14356), .IN2(n14357), .IN3(n14340), .Q(n14339) );
  XOR2X1 U15370 ( .IN1(g8275), .IN2(test_so99), .Q(n14340) );
  XOR2X1 U15371 ( .IN1(n8002), .IN2(n8001), .Q(n14338) );
  XOR2X1 U15372 ( .IN1(n14358), .IN2(n8010), .Q(n14337) );
  XOR2X1 U15373 ( .IN1(n8733), .IN2(n8011), .Q(N690) );
  XOR3X1 U15374 ( .IN1(n14341), .IN2(n14342), .IN3(n14343), .Q(n8733) );
  XOR3X1 U15375 ( .IN1(n14360), .IN2(n14361), .IN3(n14344), .Q(n14343) );
  XOR2X1 U15376 ( .IN1(g8262), .IN2(n14359), .Q(n14344) );
  XOR2X1 U15377 ( .IN1(n7974), .IN2(n7973), .Q(n14342) );
  XOR2X1 U15378 ( .IN1(n7976), .IN2(n7975), .Q(n14341) );
  NOR2X0 U3772_U2 ( .IN1(n2230), .IN2(n2217), .QN(U3772_n1) );
  INVX0 U3772_U1 ( .INP(U3772_n1), .ZN(n2231) );
  NOR2X0 U3776_U2 ( .IN1(n2374), .IN2(n2361), .QN(U3776_n1) );
  INVX0 U3776_U1 ( .INP(U3776_n1), .ZN(n2375) );
  NOR2X0 U3777_U2 ( .IN1(g51), .IN2(DFF_2_n1), .QN(U3777_n1) );
  INVX0 U3777_U1 ( .INP(U3777_n1), .ZN(n4264) );
  NOR2X0 U3778_U2 ( .IN1(n2445), .IN2(n2446), .QN(U3778_n1) );
  INVX0 U3778_U1 ( .INP(U3778_n1), .ZN(n2440) );
  NOR2X0 U3779_U2 ( .IN1(n453), .IN2(n2446), .QN(U3779_n1) );
  INVX0 U3779_U1 ( .INP(U3779_n1), .ZN(n2426) );
  NOR2X0 U3780_U2 ( .IN1(n2670), .IN2(n2671), .QN(U3780_n1) );
  INVX0 U3780_U1 ( .INP(U3780_n1), .ZN(n2669) );
  NOR2X0 U3781_U2 ( .IN1(n2685), .IN2(n2686), .QN(U3781_n1) );
  INVX0 U3781_U1 ( .INP(U3781_n1), .ZN(n2684) );
  NOR2X0 U3782_U2 ( .IN1(n2718), .IN2(n2719), .QN(U3782_n1) );
  INVX0 U3782_U1 ( .INP(U3782_n1), .ZN(n2717) );
  NOR2X0 U3783_U2 ( .IN1(n2982), .IN2(g2124), .QN(U3783_n1) );
  INVX0 U3783_U1 ( .INP(U3783_n1), .ZN(n2981) );
  NOR2X0 U3784_U2 ( .IN1(n2985), .IN2(g1430), .QN(U3784_n1) );
  INVX0 U3784_U1 ( .INP(U3784_n1), .ZN(n2984) );
  NOR2X0 U3785_U2 ( .IN1(n2988), .IN2(g744), .QN(U3785_n1) );
  INVX0 U3785_U1 ( .INP(U3785_n1), .ZN(n2987) );
  NOR2X0 U3786_U2 ( .IN1(n2991), .IN2(g56), .QN(U3786_n1) );
  INVX0 U3786_U1 ( .INP(U3786_n1), .ZN(n2990) );
  NOR2X0 U3787_U2 ( .IN1(n3742), .IN2(test_so98), .QN(U3787_n1) );
  INVX0 U3787_U1 ( .INP(U3787_n1), .ZN(n3741) );
  NOR2X0 U3901_U2 ( .IN1(n2302), .IN2(n2289), .QN(U3901_n1) );
  INVX0 U3901_U1 ( .INP(U3901_n1), .ZN(n2303) );
  NOR2X0 U3902_U2 ( .IN1(n475), .IN2(n2289), .QN(U3902_n1) );
  INVX0 U3902_U1 ( .INP(U3902_n1), .ZN(n2275) );
  INVX0 U4467_U2 ( .INP(n1392), .ZN(U4467_n1) );
  NOR2X0 U4467_U1 ( .IN1(n3254), .IN2(U4467_n1), .QN(n3252) );
  INVX0 U4904_U2 ( .INP(n2800), .ZN(U4904_n1) );
  NOR2X0 U4904_U1 ( .IN1(n148), .IN2(U4904_n1), .QN(n2798) );
  INVX0 U4930_U2 ( .INP(n2616), .ZN(U4930_n1) );
  NOR2X0 U4930_U1 ( .IN1(n148), .IN2(U4930_n1), .QN(n2594) );
  INVX0 U5128_U2 ( .INP(n3933), .ZN(U5128_n1) );
  NOR2X0 U5128_U1 ( .IN1(n4406), .IN2(U5128_n1), .QN(n3940) );
  INVX0 U5141_U2 ( .INP(n3939), .ZN(U5141_n1) );
  NOR2X0 U5141_U1 ( .IN1(n4405), .IN2(U5141_n1), .QN(n3936) );
  INVX0 U5749_U2 ( .INP(g2133), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n3160), .IN2(U5749_n1), .QN(n3159) );
  INVX0 U5750_U2 ( .INP(g1439), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n3164), .IN2(U5750_n1), .QN(n3163) );
  INVX0 U5751_U2 ( .INP(g753), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n3168), .IN2(U5751_n1), .QN(n3167) );
  INVX0 U5752_U2 ( .INP(g65), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n3172), .IN2(U5752_n1), .QN(n3171) );
  INVX0 U5753_U2 ( .INP(g2142), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n4522), .IN2(U5753_n1), .QN(n3424) );
  INVX0 U5754_U2 ( .INP(g2151), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n4526), .IN2(U5754_n1), .QN(n3683) );
  INVX0 U5755_U2 ( .INP(g2160), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n3888), .IN2(U5755_n1), .QN(n3887) );
  INVX0 U5756_U2 ( .INP(g1448), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n4523), .IN2(U5756_n1), .QN(n3427) );
  INVX0 U5757_U2 ( .INP(g1457), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n4527), .IN2(U5757_n1), .QN(n3686) );
  INVX0 U5758_U2 ( .INP(g1466), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n3891), .IN2(U5758_n1), .QN(n3890) );
  INVX0 U5759_U2 ( .INP(g762), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n3431), .IN2(U5759_n1), .QN(n3430) );
  INVX0 U5760_U2 ( .INP(g771), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n3690), .IN2(U5760_n1), .QN(n3689) );
  INVX0 U5761_U2 ( .INP(g780), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n3894), .IN2(U5761_n1), .QN(n3893) );
  INVX0 U5762_U2 ( .INP(g74), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n4521), .IN2(U5762_n1), .QN(n3433) );
  INVX0 U5763_U2 ( .INP(g83), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n4528), .IN2(U5763_n1), .QN(n3692) );
  INVX0 U5764_U2 ( .INP(g92), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n3897), .IN2(U5764_n1), .QN(n3896) );
  INVX0 U5882_U2 ( .INP(n1543), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(g3036), .IN2(U5882_n1), .QN(n4101) );
  INVX0 U5939_U2 ( .INP(g2257), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n1261), .IN2(U5939_n1), .QN(n3038) );
  INVX0 U5940_U2 ( .INP(g1563), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n959), .IN2(U5940_n1), .QN(n3070) );
  INVX0 U5941_U2 ( .INP(g869), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n653), .IN2(U5941_n1), .QN(n3102) );
  INVX0 U5942_U2 ( .INP(g181), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n309), .IN2(U5942_n1), .QN(n3130) );
  INVX0 U6140_U2 ( .INP(g3002), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n4066), .IN2(U6140_n1), .QN(n4065) );
  INVX0 U6460_U2 ( .INP(g3233), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(g3230), .IN2(U6460_n1), .QN(n3700) );
  INVX0 U6470_U2 ( .INP(g2892), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n4305), .IN2(U6470_n1), .QN(n4182) );
  INVX0 U6562_U2 ( .INP(n3938), .ZN(U6562_n1) );
  NOR2X0 U6562_U1 ( .IN1(g3204), .IN2(U6562_n1), .QN(n3939) );
  INVX0 U6563_U2 ( .INP(n4073), .ZN(U6563_n1) );
  NOR2X0 U6563_U1 ( .IN1(g3204), .IN2(U6563_n1), .QN(n3705) );
  INVX0 U6718_U2 ( .INP(n266), .ZN(U6718_n1) );
  NOR2X0 U6718_U1 ( .IN1(g3197), .IN2(U6718_n1), .QN(n4073) );
  INVX0 U7116_U2 ( .INP(n4058), .ZN(U7116_n1) );
  NOR2X0 U7116_U1 ( .IN1(g2903), .IN2(U7116_n1), .QN(n4057) );
  INVX0 U7118_U2 ( .INP(n10), .ZN(U7118_n1) );
  NOR2X0 U7118_U1 ( .IN1(g2896), .IN2(U7118_n1), .QN(n4122) );
  INVX0 U7293_U2 ( .INP(n4598), .ZN(U7293_n1) );
  NOR2X0 U7293_U1 ( .IN1(g3234), .IN2(U7293_n1), .QN(g20877) );
endmodule

