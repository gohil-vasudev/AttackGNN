module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n1359_, new_n595_, new_n1233_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n501_, new_n1157_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1433_, new_n1517_, new_n1575_, new_n1472_, new_n1048_, new_n885_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n1327_, new_n241_, new_n1535_, new_n566_, new_n641_, new_n339_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n1351_, new_n556_, new_n636_, new_n691_, new_n1024_, new_n670_, new_n456_, new_n1125_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n1568_, new_n728_, new_n1479_, new_n1071_, new_n1294_, new_n214_, new_n894_, new_n853_, new_n695_, new_n660_, new_n1311_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n706_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n1415_, new_n1390_, new_n721_, new_n504_, new_n1414_, new_n742_, new_n892_, new_n1368_, new_n234_, new_n472_, new_n873_, new_n1167_, new_n1530_, new_n1300_, new_n1490_, new_n774_, new_n792_, new_n953_, new_n257_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n1580_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n1447_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n983_, new_n822_, new_n1406_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n1054_, new_n655_, new_n1288_, new_n630_, new_n385_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n297_, new_n565_, new_n1196_, new_n1366_, new_n511_, new_n303_, new_n325_, new_n1285_, new_n1031_, new_n1216_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n324_, new_n960_, new_n1377_, new_n1522_, new_n549_, new_n491_, new_n676_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n1463_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1424_, new_n1062_, new_n680_, new_n981_, new_n506_, new_n872_, new_n1527_, new_n1275_, new_n1198_, new_n1428_, new_n1440_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n483_, new_n1004_, new_n1152_, new_n1558_, new_n299_, new_n394_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n363_, new_n1266_, new_n785_, new_n1501_, new_n441_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n1562_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n1576_, new_n301_, new_n1333_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n207_, new_n267_, new_n1395_, new_n473_, new_n1147_, new_n1373_, new_n1229_, new_n1422_, new_n1523_, new_n1468_, new_n969_, new_n334_, new_n331_, new_n1234_, new_n835_, new_n1360_, new_n378_, new_n1574_, new_n621_, new_n1423_, new_n244_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1321_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n1419_, new_n921_, new_n346_, new_n396_, new_n1003_, new_n696_, new_n208_, new_n1039_, new_n1507_, new_n1439_, new_n1365_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n729_, new_n1111_, new_n1413_, new_n1218_, new_n1385_, new_n1346_, new_n1201_, new_n559_, new_n1282_, new_n762_, new_n1349_, new_n1193_, new_n1547_, new_n1437_, new_n1187_, new_n1205_, new_n1154_, new_n1253_, new_n1546_, new_n295_, new_n1453_, new_n1256_, new_n628_, new_n1513_, new_n409_, new_n1090_, new_n745_, new_n1489_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n1573_, new_n369_, new_n1171_, new_n867_, new_n954_, new_n1032_, new_n1545_, new_n276_, new_n901_, new_n688_, new_n1255_, new_n410_, new_n985_, new_n851_, new_n1518_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n202_, new_n296_, new_n661_, new_n797_, new_n232_, new_n1358_, new_n724_, new_n1070_, new_n1416_, new_n1109_, new_n261_, new_n672_, new_n1496_, new_n1269_, new_n616_, new_n529_, new_n323_, new_n914_, new_n884_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n604_, new_n1461_, new_n1104_, new_n1511_, new_n571_, new_n1504_, new_n758_, new_n460_, new_n1267_, new_n328_, new_n268_, new_n1466_, new_n1516_, new_n1299_, new_n380_, new_n1477_, new_n1079_, new_n861_, new_n1564_, new_n1252_, new_n352_, new_n1553_, new_n931_, new_n575_, new_n1493_, new_n562_, new_n944_, new_n1542_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n1480_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n963_, new_n1481_, new_n1325_, new_n993_, new_n1191_, new_n1357_, new_n824_, new_n717_, new_n1455_, new_n403_, new_n868_, new_n1242_, new_n475_, new_n237_, new_n858_, new_n1384_, new_n1343_, new_n936_, new_n1459_, new_n1434_, new_n1438_, new_n1016_, new_n411_, new_n673_, new_n1144_, new_n1465_, new_n666_, new_n1290_, new_n407_, new_n1519_, new_n1407_, new_n879_, new_n1417_, new_n736_, new_n513_, new_n558_, new_n219_, new_n382_, new_n313_, new_n1370_, new_n239_, new_n718_, new_n1310_, new_n1398_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n302_, new_n755_, new_n1509_, new_n1559_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n345_, new_n499_, new_n533_, new_n255_, new_n1130_, new_n795_, new_n459_, new_n1441_, new_n1122_, new_n1185_, new_n1240_, new_n1510_, new_n354_, new_n1174_, new_n968_, new_n1464_, new_n613_, new_n1508_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n837_, new_n591_, new_n801_, new_n1458_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1521_, new_n1334_, new_n531_, new_n593_, new_n1543_, new_n974_, new_n1565_, new_n252_, new_n1248_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n1474_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n1430_, new_n470_, new_n213_, new_n769_, new_n433_, new_n871_, new_n1450_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n933_, new_n584_, new_n815_, new_n278_, new_n304_, new_n1052_, new_n1425_, new_n857_, new_n1379_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1471_, new_n1220_, new_n989_, new_n1117_, new_n1421_, new_n644_, new_n836_, new_n1116_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n1427_, new_n818_, new_n881_, new_n1268_, new_n1376_, new_n1381_, new_n1566_, new_n1534_, new_n684_, new_n640_, new_n1274_, new_n754_, new_n653_, new_n905_, new_n377_, new_n1539_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1391_, new_n1436_, new_n567_, new_n1353_, new_n1033_, new_n576_, new_n831_, new_n791_, new_n1153_, new_n357_, new_n1339_, new_n320_, new_n984_, new_n780_, new_n1183_, new_n245_, new_n643_, new_n1316_, new_n1194_, new_n1338_, new_n1460_, new_n1230_, new_n1027_, new_n348_, new_n610_, new_n1369_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1165_, new_n1401_, new_n1259_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n686_, new_n293_, new_n934_, new_n1567_, new_n770_, new_n1389_, new_n1400_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n1249_, new_n1354_, new_n955_, new_n847_, new_n250_, new_n888_, new_n1505_, new_n288_, new_n1340_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1361_, new_n941_, new_n1410_, new_n738_, new_n827_, new_n1356_, new_n1363_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n1211_, new_n1412_, new_n1207_, new_n1176_, new_n1374_, new_n601_, new_n842_, new_n1552_, new_n1057_, new_n682_, new_n812_, new_n1563_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1397_, new_n220_, new_n1402_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n804_, new_n1342_, new_n424_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n240_, new_n413_, new_n1544_, new_n1382_, new_n442_, new_n677_, new_n1487_, new_n642_, new_n211_, new_n1418_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n761_, new_n840_, new_n735_, new_n1283_, new_n898_, new_n799_, new_n1304_, new_n1537_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n1469_, new_n862_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n1585_, new_n1587_, new_n1264_, new_n215_, new_n1319_, new_n626_, new_n959_, new_n990_, new_n716_, new_n701_, new_n1238_, new_n1058_, new_n1162_, new_n212_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n414_, new_n1101_, new_n1250_, new_n315_, new_n1482_, new_n1050_, new_n554_, new_n230_, new_n844_, new_n1302_, new_n281_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n1297_, new_n829_, new_n1257_, new_n1306_, new_n988_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n1486_, new_n361_, new_n764_, new_n906_, new_n683_, new_n1409_, new_n1429_, new_n463_, new_n1372_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n1292_, new_n1426_, new_n517_, new_n609_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n1560_, new_n715_, new_n811_, new_n1445_, new_n1371_, new_n443_, new_n1086_, new_n763_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1452_, new_n1051_, new_n899_, new_n1053_, new_n1540_, new_n205_, new_n492_, new_n1200_, new_n1533_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1483_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n820_, new_n771_, new_n979_, new_n508_, new_n714_, new_n1280_, new_n1007_, new_n1241_, new_n882_, new_n1145_, new_n1557_, new_n929_, new_n986_, new_n1159_, new_n314_, new_n1584_, new_n1337_, new_n216_, new_n917_, new_n1555_, new_n1322_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n541_, new_n210_, new_n447_, new_n1388_, new_n1550_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n1247_, new_n1411_, new_n465_, new_n783_, new_n1380_, new_n739_, new_n263_, new_n341_, new_n996_, new_n1318_, new_n846_, new_n915_, new_n488_, new_n524_, new_n349_, new_n848_, new_n277_, new_n1245_, new_n663_, new_n1499_, new_n1497_, new_n579_, new_n286_, new_n1375_, new_n1254_, new_n438_, new_n1344_, new_n939_, new_n1393_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n1514_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n1526_, new_n397_, new_n1446_, new_n975_, new_n1199_, new_n399_, new_n1581_, new_n596_, new_n870_, new_n805_, new_n1420_, new_n1403_, new_n1115_, new_n1383_, new_n1231_, new_n948_, new_n1520_, new_n1055_, new_n1431_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n457_, new_n1301_, new_n1128_, new_n1582_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1329_, new_n1161_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n1000_, new_n308_, new_n633_, new_n784_, new_n1273_, new_n1396_, new_n1491_, new_n1554_, new_n258_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n1166_, new_n259_, new_n1536_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n1043_, new_n222_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n1272_, new_n693_, new_n1287_, new_n1485_, new_n505_, new_n1462_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1538_, new_n1579_, new_n1289_, new_n1561_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n1095_, new_n310_, new_n275_, new_n998_, new_n1056_, new_n1331_, new_n839_, new_n1030_, new_n485_, new_n578_, new_n525_, new_n918_, new_n1586_, new_n810_, new_n808_, new_n1284_, new_n1572_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n1387_, new_n719_, new_n869_, new_n1178_, new_n1525_, new_n270_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n520_, new_n1347_, new_n1001_, new_n253_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n1503_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n1286_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n1326_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n231_, new_n1080_, new_n583_, new_n617_, new_n1279_, new_n1467_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n916_, new_n428_, new_n487_, new_n675_, new_n1155_, new_n360_, new_n1186_, new_n1261_, new_n225_, new_n1246_, new_n1488_, new_n922_, new_n387_, new_n476_, new_n987_, new_n949_, new_n221_, new_n450_, new_n1394_, new_n243_, new_n1179_, new_n298_, new_n1088_, new_n1148_, new_n569_, new_n555_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n209_, new_n623_, new_n446_, new_n316_, new_n203_, new_n590_, new_n826_, new_n789_, new_n1476_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n1350_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n307_, new_n1378_, new_n1478_, new_n1181_, new_n1093_, new_n597_, new_n1451_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n435_, new_n1309_, new_n1010_, new_n776_, new_n687_, new_n1029_, new_n370_, new_n1515_, new_n638_, new_n523_, new_n909_, new_n1571_, new_n217_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1470_, new_n1112_, new_n711_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1475_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n1529_, new_n1541_, new_n645_, new_n1087_, new_n1096_, new_n723_, new_n756_, new_n823_, new_n1549_, new_n1577_, new_n574_, new_n1500_, new_n928_, new_n1548_, new_n1578_, new_n319_, new_n1008_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n1291_, new_n247_, new_n539_, new_n1399_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n1531_, new_n294_, new_n1295_, new_n1173_, new_n704_, new_n1432_, new_n1189_, new_n1197_, new_n1312_, new_n1502_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n467_, new_n404_, new_n1243_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n1506_, new_n1583_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n1556_, new_n947_, new_n994_, new_n982_, new_n1494_, new_n1449_, new_n964_, new_n1078_, new_n551_, new_n1408_, new_n279_, new_n455_, new_n1569_, new_n618_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n464_, new_n1498_, new_n204_, new_n1588_, new_n573_, new_n765_, new_n1314_, new_n1103_;

not g0000 ( new_n202_, keyIn_0_55 );
not g0001 ( new_n203_, keyIn_0_10 );
not g0002 ( new_n204_, N81 );
nor g0003 ( new_n205_, new_n204_, N85 );
not g0004 ( new_n206_, N85 );
nor g0005 ( new_n207_, new_n206_, N81 );
nor g0006 ( new_n208_, new_n205_, new_n207_ );
not g0007 ( new_n209_, new_n208_ );
nand g0008 ( new_n210_, new_n209_, new_n203_ );
not g0009 ( new_n211_, new_n210_ );
nor g0010 ( new_n212_, new_n209_, new_n203_ );
nor g0011 ( new_n213_, new_n211_, new_n212_ );
not g0012 ( new_n214_, new_n213_ );
not g0013 ( new_n215_, N89 );
nor g0014 ( new_n216_, new_n215_, N93 );
not g0015 ( new_n217_, N93 );
nor g0016 ( new_n218_, new_n217_, N89 );
nor g0017 ( new_n219_, new_n216_, new_n218_ );
not g0018 ( new_n220_, new_n219_ );
nand g0019 ( new_n221_, new_n220_, keyIn_0_11 );
not g0020 ( new_n222_, new_n221_ );
nor g0021 ( new_n223_, new_n220_, keyIn_0_11 );
nor g0022 ( new_n224_, new_n222_, new_n223_ );
not g0023 ( new_n225_, new_n224_ );
nand g0024 ( new_n226_, new_n214_, new_n225_ );
nand g0025 ( new_n227_, new_n213_, new_n224_ );
nand g0026 ( new_n228_, new_n226_, new_n227_ );
nand g0027 ( new_n229_, new_n228_, keyIn_0_33 );
not g0028 ( new_n230_, new_n229_ );
nor g0029 ( new_n231_, new_n228_, keyIn_0_33 );
nor g0030 ( new_n232_, new_n230_, new_n231_ );
not g0031 ( new_n233_, new_n232_ );
not g0032 ( new_n234_, keyIn_0_8 );
not g0033 ( new_n235_, N65 );
nor g0034 ( new_n236_, new_n235_, N69 );
not g0035 ( new_n237_, N69 );
nor g0036 ( new_n238_, new_n237_, N65 );
nor g0037 ( new_n239_, new_n236_, new_n238_ );
not g0038 ( new_n240_, new_n239_ );
nand g0039 ( new_n241_, new_n240_, new_n234_ );
not g0040 ( new_n242_, new_n241_ );
nor g0041 ( new_n243_, new_n240_, new_n234_ );
nor g0042 ( new_n244_, new_n242_, new_n243_ );
not g0043 ( new_n245_, new_n244_ );
not g0044 ( new_n246_, N73 );
nor g0045 ( new_n247_, new_n246_, N77 );
not g0046 ( new_n248_, N77 );
nor g0047 ( new_n249_, new_n248_, N73 );
nor g0048 ( new_n250_, new_n247_, new_n249_ );
not g0049 ( new_n251_, new_n250_ );
nand g0050 ( new_n252_, new_n251_, keyIn_0_9 );
not g0051 ( new_n253_, new_n252_ );
nor g0052 ( new_n254_, new_n251_, keyIn_0_9 );
nor g0053 ( new_n255_, new_n253_, new_n254_ );
not g0054 ( new_n256_, new_n255_ );
nand g0055 ( new_n257_, new_n245_, new_n256_ );
nand g0056 ( new_n258_, new_n244_, new_n255_ );
nand g0057 ( new_n259_, new_n257_, new_n258_ );
nand g0058 ( new_n260_, new_n259_, keyIn_0_32 );
not g0059 ( new_n261_, new_n260_ );
nor g0060 ( new_n262_, new_n259_, keyIn_0_32 );
nor g0061 ( new_n263_, new_n261_, new_n262_ );
nand g0062 ( new_n264_, new_n233_, new_n263_ );
not g0063 ( new_n265_, new_n263_ );
nand g0064 ( new_n266_, new_n265_, new_n232_ );
nand g0065 ( new_n267_, new_n264_, new_n266_ );
nand g0066 ( new_n268_, new_n267_, keyIn_0_43 );
not g0067 ( new_n269_, new_n268_ );
nor g0068 ( new_n270_, new_n267_, keyIn_0_43 );
nor g0069 ( new_n271_, new_n269_, new_n270_ );
not g0070 ( new_n272_, new_n271_ );
nand g0071 ( new_n273_, N129, N137 );
not g0072 ( new_n274_, new_n273_ );
nor g0073 ( new_n275_, new_n272_, new_n274_ );
not g0074 ( new_n276_, new_n275_ );
nor g0075 ( new_n277_, new_n271_, new_n273_ );
not g0076 ( new_n278_, new_n277_ );
nand g0077 ( new_n279_, new_n276_, new_n278_ );
nand g0078 ( new_n280_, new_n279_, keyIn_0_47 );
not g0079 ( new_n281_, new_n280_ );
nor g0080 ( new_n282_, new_n279_, keyIn_0_47 );
nor g0081 ( new_n283_, new_n281_, new_n282_ );
not g0082 ( new_n284_, N1 );
nor g0083 ( new_n285_, new_n284_, N17 );
not g0084 ( new_n286_, N17 );
nor g0085 ( new_n287_, new_n286_, N1 );
nor g0086 ( new_n288_, new_n285_, new_n287_ );
not g0087 ( new_n289_, new_n288_ );
nand g0088 ( new_n290_, N33, N49 );
not g0089 ( new_n291_, new_n290_ );
nor g0090 ( new_n292_, N33, N49 );
nor g0091 ( new_n293_, new_n291_, new_n292_ );
not g0092 ( new_n294_, new_n293_ );
nor g0093 ( new_n295_, new_n289_, new_n294_ );
nor g0094 ( new_n296_, new_n288_, new_n293_ );
nor g0095 ( new_n297_, new_n295_, new_n296_ );
nor g0096 ( new_n298_, new_n283_, new_n297_ );
not g0097 ( new_n299_, keyIn_0_47 );
not g0098 ( new_n300_, new_n279_ );
nand g0099 ( new_n301_, new_n300_, new_n299_ );
nand g0100 ( new_n302_, new_n301_, new_n280_ );
not g0101 ( new_n303_, new_n297_ );
nor g0102 ( new_n304_, new_n302_, new_n303_ );
nor g0103 ( new_n305_, new_n298_, new_n304_ );
nand g0104 ( new_n306_, new_n305_, new_n202_ );
nand g0105 ( new_n307_, new_n302_, new_n303_ );
nand g0106 ( new_n308_, new_n283_, new_n297_ );
nand g0107 ( new_n309_, new_n308_, new_n307_ );
nand g0108 ( new_n310_, new_n309_, keyIn_0_55 );
nand g0109 ( new_n311_, new_n306_, new_n310_ );
not g0110 ( new_n312_, new_n311_ );
not g0111 ( new_n313_, keyIn_0_58 );
not g0112 ( new_n314_, keyIn_0_46 );
not g0113 ( new_n315_, N113 );
nor g0114 ( new_n316_, new_n315_, N117 );
not g0115 ( new_n317_, N117 );
nor g0116 ( new_n318_, new_n317_, N113 );
nor g0117 ( new_n319_, new_n316_, new_n318_ );
not g0118 ( new_n320_, new_n319_ );
nand g0119 ( new_n321_, new_n320_, keyIn_0_14 );
not g0120 ( new_n322_, new_n321_ );
nor g0121 ( new_n323_, new_n320_, keyIn_0_14 );
nor g0122 ( new_n324_, new_n322_, new_n323_ );
not g0123 ( new_n325_, new_n324_ );
not g0124 ( new_n326_, N121 );
nor g0125 ( new_n327_, new_n326_, N125 );
not g0126 ( new_n328_, N125 );
nor g0127 ( new_n329_, new_n328_, N121 );
nor g0128 ( new_n330_, new_n327_, new_n329_ );
not g0129 ( new_n331_, new_n330_ );
nand g0130 ( new_n332_, new_n331_, keyIn_0_15 );
not g0131 ( new_n333_, new_n332_ );
nor g0132 ( new_n334_, new_n331_, keyIn_0_15 );
nor g0133 ( new_n335_, new_n333_, new_n334_ );
not g0134 ( new_n336_, new_n335_ );
nand g0135 ( new_n337_, new_n325_, new_n336_ );
nand g0136 ( new_n338_, new_n324_, new_n335_ );
nand g0137 ( new_n339_, new_n337_, new_n338_ );
nand g0138 ( new_n340_, new_n339_, keyIn_0_35 );
not g0139 ( new_n341_, new_n340_ );
nor g0140 ( new_n342_, new_n339_, keyIn_0_35 );
nor g0141 ( new_n343_, new_n341_, new_n342_ );
not g0142 ( new_n344_, new_n343_ );
nand g0143 ( new_n345_, new_n233_, new_n344_ );
nand g0144 ( new_n346_, new_n232_, new_n343_ );
nand g0145 ( new_n347_, new_n345_, new_n346_ );
nand g0146 ( new_n348_, new_n347_, new_n314_ );
not g0147 ( new_n349_, new_n348_ );
nor g0148 ( new_n350_, new_n347_, new_n314_ );
nor g0149 ( new_n351_, new_n349_, new_n350_ );
not g0150 ( new_n352_, new_n351_ );
nand g0151 ( new_n353_, N132, N137 );
not g0152 ( new_n354_, new_n353_ );
nand g0153 ( new_n355_, new_n352_, new_n354_ );
nand g0154 ( new_n356_, new_n351_, new_n353_ );
nand g0155 ( new_n357_, new_n355_, new_n356_ );
nand g0156 ( new_n358_, new_n357_, keyIn_0_50 );
not g0157 ( new_n359_, new_n358_ );
nor g0158 ( new_n360_, new_n357_, keyIn_0_50 );
nor g0159 ( new_n361_, new_n359_, new_n360_ );
nand g0160 ( new_n362_, N13, N29 );
not g0161 ( new_n363_, new_n362_ );
nor g0162 ( new_n364_, N13, N29 );
nor g0163 ( new_n365_, new_n363_, new_n364_ );
not g0164 ( new_n366_, new_n365_ );
nor g0165 ( new_n367_, new_n366_, keyIn_0_23 );
nand g0166 ( new_n368_, new_n366_, keyIn_0_23 );
not g0167 ( new_n369_, new_n368_ );
nor g0168 ( new_n370_, new_n369_, new_n367_ );
not g0169 ( new_n371_, new_n370_ );
not g0170 ( new_n372_, N45 );
nor g0171 ( new_n373_, new_n372_, N61 );
not g0172 ( new_n374_, N61 );
nor g0173 ( new_n375_, new_n374_, N45 );
nor g0174 ( new_n376_, new_n373_, new_n375_ );
not g0175 ( new_n377_, new_n376_ );
nor g0176 ( new_n378_, new_n371_, new_n377_ );
nor g0177 ( new_n379_, new_n370_, new_n376_ );
nor g0178 ( new_n380_, new_n378_, new_n379_ );
nor g0179 ( new_n381_, new_n361_, new_n380_ );
nand g0180 ( new_n382_, new_n361_, new_n380_ );
not g0181 ( new_n383_, new_n382_ );
nor g0182 ( new_n384_, new_n383_, new_n381_ );
nand g0183 ( new_n385_, new_n384_, new_n313_ );
not g0184 ( new_n386_, new_n381_ );
nand g0185 ( new_n387_, new_n386_, new_n382_ );
nand g0186 ( new_n388_, new_n387_, keyIn_0_58 );
nand g0187 ( new_n389_, new_n385_, new_n388_ );
not g0188 ( new_n390_, keyIn_0_57 );
not g0189 ( new_n391_, N97 );
nor g0190 ( new_n392_, new_n391_, N101 );
not g0191 ( new_n393_, N101 );
nor g0192 ( new_n394_, new_n393_, N97 );
nor g0193 ( new_n395_, new_n392_, new_n394_ );
not g0194 ( new_n396_, new_n395_ );
nand g0195 ( new_n397_, new_n396_, keyIn_0_12 );
not g0196 ( new_n398_, new_n397_ );
nor g0197 ( new_n399_, new_n396_, keyIn_0_12 );
nor g0198 ( new_n400_, new_n398_, new_n399_ );
not g0199 ( new_n401_, new_n400_ );
not g0200 ( new_n402_, N105 );
nor g0201 ( new_n403_, new_n402_, N109 );
not g0202 ( new_n404_, N109 );
nor g0203 ( new_n405_, new_n404_, N105 );
nor g0204 ( new_n406_, new_n403_, new_n405_ );
not g0205 ( new_n407_, new_n406_ );
nand g0206 ( new_n408_, new_n407_, keyIn_0_13 );
not g0207 ( new_n409_, new_n408_ );
nor g0208 ( new_n410_, new_n407_, keyIn_0_13 );
nor g0209 ( new_n411_, new_n409_, new_n410_ );
not g0210 ( new_n412_, new_n411_ );
nand g0211 ( new_n413_, new_n401_, new_n412_ );
nand g0212 ( new_n414_, new_n400_, new_n411_ );
nand g0213 ( new_n415_, new_n413_, new_n414_ );
nand g0214 ( new_n416_, new_n415_, keyIn_0_34 );
not g0215 ( new_n417_, new_n416_ );
nor g0216 ( new_n418_, new_n415_, keyIn_0_34 );
nor g0217 ( new_n419_, new_n417_, new_n418_ );
not g0218 ( new_n420_, new_n419_ );
nand g0219 ( new_n421_, new_n265_, new_n420_ );
nand g0220 ( new_n422_, new_n263_, new_n419_ );
nand g0221 ( new_n423_, new_n421_, new_n422_ );
nand g0222 ( new_n424_, new_n423_, keyIn_0_45 );
not g0223 ( new_n425_, new_n424_ );
nor g0224 ( new_n426_, new_n423_, keyIn_0_45 );
nor g0225 ( new_n427_, new_n425_, new_n426_ );
nand g0226 ( new_n428_, N131, N137 );
nand g0227 ( new_n429_, new_n428_, keyIn_0_16 );
not g0228 ( new_n430_, new_n429_ );
nor g0229 ( new_n431_, new_n428_, keyIn_0_16 );
nor g0230 ( new_n432_, new_n430_, new_n431_ );
nor g0231 ( new_n433_, new_n427_, new_n432_ );
not g0232 ( new_n434_, new_n433_ );
nand g0233 ( new_n435_, new_n427_, new_n432_ );
nand g0234 ( new_n436_, new_n434_, new_n435_ );
nand g0235 ( new_n437_, new_n436_, keyIn_0_49 );
not g0236 ( new_n438_, keyIn_0_49 );
not g0237 ( new_n439_, new_n435_ );
nor g0238 ( new_n440_, new_n439_, new_n433_ );
nand g0239 ( new_n441_, new_n440_, new_n438_ );
nand g0240 ( new_n442_, new_n441_, new_n437_ );
not g0241 ( new_n443_, N9 );
nor g0242 ( new_n444_, new_n443_, N25 );
not g0243 ( new_n445_, N25 );
nor g0244 ( new_n446_, new_n445_, N9 );
nor g0245 ( new_n447_, new_n444_, new_n446_ );
not g0246 ( new_n448_, new_n447_ );
nand g0247 ( new_n449_, new_n448_, keyIn_0_21 );
not g0248 ( new_n450_, new_n449_ );
nor g0249 ( new_n451_, new_n448_, keyIn_0_21 );
nor g0250 ( new_n452_, new_n450_, new_n451_ );
not g0251 ( new_n453_, N41 );
nor g0252 ( new_n454_, new_n453_, N57 );
not g0253 ( new_n455_, N57 );
nor g0254 ( new_n456_, new_n455_, N41 );
nor g0255 ( new_n457_, new_n454_, new_n456_ );
not g0256 ( new_n458_, new_n457_ );
nand g0257 ( new_n459_, new_n458_, keyIn_0_22 );
not g0258 ( new_n460_, new_n459_ );
nor g0259 ( new_n461_, new_n458_, keyIn_0_22 );
nor g0260 ( new_n462_, new_n460_, new_n461_ );
not g0261 ( new_n463_, new_n462_ );
nor g0262 ( new_n464_, new_n463_, new_n452_ );
nand g0263 ( new_n465_, new_n463_, new_n452_ );
not g0264 ( new_n466_, new_n465_ );
nor g0265 ( new_n467_, new_n466_, new_n464_ );
not g0266 ( new_n468_, new_n467_ );
nand g0267 ( new_n469_, new_n468_, keyIn_0_36 );
not g0268 ( new_n470_, new_n469_ );
nor g0269 ( new_n471_, new_n468_, keyIn_0_36 );
nor g0270 ( new_n472_, new_n470_, new_n471_ );
not g0271 ( new_n473_, new_n472_ );
nand g0272 ( new_n474_, new_n442_, new_n473_ );
not g0273 ( new_n475_, new_n474_ );
nor g0274 ( new_n476_, new_n442_, new_n473_ );
nor g0275 ( new_n477_, new_n475_, new_n476_ );
nand g0276 ( new_n478_, new_n477_, new_n390_ );
not g0277 ( new_n479_, new_n476_ );
nand g0278 ( new_n480_, new_n479_, new_n474_ );
nand g0279 ( new_n481_, new_n480_, keyIn_0_57 );
nand g0280 ( new_n482_, new_n478_, new_n481_ );
not g0281 ( new_n483_, keyIn_0_56 );
not g0282 ( new_n484_, keyIn_0_48 );
nand g0283 ( new_n485_, new_n344_, new_n420_ );
nand g0284 ( new_n486_, new_n343_, new_n419_ );
nand g0285 ( new_n487_, new_n485_, new_n486_ );
nand g0286 ( new_n488_, new_n487_, keyIn_0_44 );
not g0287 ( new_n489_, new_n488_ );
nor g0288 ( new_n490_, new_n487_, keyIn_0_44 );
nor g0289 ( new_n491_, new_n489_, new_n490_ );
nand g0290 ( new_n492_, N130, N137 );
nand g0291 ( new_n493_, new_n491_, new_n492_ );
not g0292 ( new_n494_, new_n493_ );
nor g0293 ( new_n495_, new_n491_, new_n492_ );
nor g0294 ( new_n496_, new_n494_, new_n495_ );
nand g0295 ( new_n497_, new_n496_, new_n484_ );
not g0296 ( new_n498_, new_n495_ );
nand g0297 ( new_n499_, new_n498_, new_n493_ );
nand g0298 ( new_n500_, new_n499_, keyIn_0_48 );
nand g0299 ( new_n501_, new_n497_, new_n500_ );
not g0300 ( new_n502_, N5 );
nor g0301 ( new_n503_, new_n502_, N21 );
not g0302 ( new_n504_, N21 );
nor g0303 ( new_n505_, new_n504_, N5 );
nor g0304 ( new_n506_, new_n503_, new_n505_ );
not g0305 ( new_n507_, new_n506_ );
nand g0306 ( new_n508_, N37, N53 );
not g0307 ( new_n509_, new_n508_ );
nor g0308 ( new_n510_, N37, N53 );
nor g0309 ( new_n511_, new_n509_, new_n510_ );
not g0310 ( new_n512_, new_n511_ );
nor g0311 ( new_n513_, new_n507_, new_n512_ );
nor g0312 ( new_n514_, new_n506_, new_n511_ );
nor g0313 ( new_n515_, new_n513_, new_n514_ );
not g0314 ( new_n516_, new_n515_ );
nand g0315 ( new_n517_, new_n501_, new_n516_ );
not g0316 ( new_n518_, new_n517_ );
nor g0317 ( new_n519_, new_n501_, new_n516_ );
nor g0318 ( new_n520_, new_n518_, new_n519_ );
nand g0319 ( new_n521_, new_n520_, new_n483_ );
not g0320 ( new_n522_, new_n501_ );
nand g0321 ( new_n523_, new_n522_, new_n515_ );
nand g0322 ( new_n524_, new_n523_, new_n517_ );
nand g0323 ( new_n525_, new_n524_, keyIn_0_56 );
nand g0324 ( new_n526_, new_n521_, new_n525_ );
nand g0325 ( new_n527_, new_n482_, new_n526_ );
nor g0326 ( new_n528_, new_n527_, new_n389_ );
not g0327 ( new_n529_, new_n528_ );
nand g0328 ( new_n530_, new_n527_, new_n389_ );
nor g0329 ( new_n531_, new_n482_, new_n526_ );
nor g0330 ( new_n532_, new_n531_, new_n311_ );
nand g0331 ( new_n533_, new_n532_, new_n530_ );
not g0332 ( new_n534_, new_n533_ );
nand g0333 ( new_n535_, new_n534_, new_n529_ );
not g0334 ( new_n536_, keyIn_0_63 );
not g0335 ( new_n537_, new_n482_ );
nand g0336 ( new_n538_, new_n537_, new_n536_ );
nand g0337 ( new_n539_, new_n482_, keyIn_0_63 );
nand g0338 ( new_n540_, new_n538_, new_n539_ );
nand g0339 ( new_n541_, new_n311_, new_n526_ );
nor g0340 ( new_n542_, new_n541_, new_n389_ );
nand g0341 ( new_n543_, new_n542_, new_n540_ );
nand g0342 ( new_n544_, new_n535_, new_n543_ );
not g0343 ( new_n545_, keyIn_0_42 );
nor g0344 ( new_n546_, N25, N29 );
not g0345 ( new_n547_, new_n546_ );
nand g0346 ( new_n548_, N25, N29 );
nand g0347 ( new_n549_, new_n547_, new_n548_ );
nand g0348 ( new_n550_, new_n549_, keyIn_0_3 );
not g0349 ( new_n551_, keyIn_0_3 );
not g0350 ( new_n552_, new_n548_ );
nor g0351 ( new_n553_, new_n552_, new_n546_ );
nand g0352 ( new_n554_, new_n553_, new_n551_ );
nand g0353 ( new_n555_, new_n550_, new_n554_ );
not g0354 ( new_n556_, keyIn_0_2 );
nand g0355 ( new_n557_, new_n286_, new_n504_ );
nand g0356 ( new_n558_, N17, N21 );
nand g0357 ( new_n559_, new_n557_, new_n558_ );
nand g0358 ( new_n560_, new_n559_, new_n556_ );
nor g0359 ( new_n561_, N17, N21 );
not g0360 ( new_n562_, new_n558_ );
nor g0361 ( new_n563_, new_n562_, new_n561_ );
nand g0362 ( new_n564_, new_n563_, keyIn_0_2 );
nand g0363 ( new_n565_, new_n564_, new_n560_ );
nand g0364 ( new_n566_, new_n555_, new_n565_ );
not g0365 ( new_n567_, new_n566_ );
nor g0366 ( new_n568_, new_n555_, new_n565_ );
nor g0367 ( new_n569_, new_n567_, new_n568_ );
nand g0368 ( new_n570_, new_n569_, keyIn_0_29 );
not g0369 ( new_n571_, keyIn_0_29 );
not g0370 ( new_n572_, new_n555_ );
not g0371 ( new_n573_, new_n565_ );
nand g0372 ( new_n574_, new_n572_, new_n573_ );
nand g0373 ( new_n575_, new_n574_, new_n566_ );
nand g0374 ( new_n576_, new_n575_, new_n571_ );
nand g0375 ( new_n577_, new_n570_, new_n576_ );
not g0376 ( new_n578_, keyIn_0_31 );
not g0377 ( new_n579_, keyIn_0_6 );
nand g0378 ( new_n580_, N49, N53 );
not g0379 ( new_n581_, new_n580_ );
nor g0380 ( new_n582_, N49, N53 );
nor g0381 ( new_n583_, new_n581_, new_n582_ );
nand g0382 ( new_n584_, new_n583_, new_n579_ );
not g0383 ( new_n585_, new_n582_ );
nand g0384 ( new_n586_, new_n585_, new_n580_ );
nand g0385 ( new_n587_, new_n586_, keyIn_0_6 );
nand g0386 ( new_n588_, new_n587_, new_n584_ );
not g0387 ( new_n589_, keyIn_0_7 );
nand g0388 ( new_n590_, N57, N61 );
not g0389 ( new_n591_, new_n590_ );
nor g0390 ( new_n592_, N57, N61 );
nor g0391 ( new_n593_, new_n591_, new_n592_ );
nand g0392 ( new_n594_, new_n593_, new_n589_ );
nand g0393 ( new_n595_, new_n455_, new_n374_ );
nand g0394 ( new_n596_, new_n595_, new_n590_ );
nand g0395 ( new_n597_, new_n596_, keyIn_0_7 );
nand g0396 ( new_n598_, new_n594_, new_n597_ );
nand g0397 ( new_n599_, new_n588_, new_n598_ );
not g0398 ( new_n600_, new_n599_ );
nor g0399 ( new_n601_, new_n588_, new_n598_ );
nor g0400 ( new_n602_, new_n600_, new_n601_ );
nand g0401 ( new_n603_, new_n602_, new_n578_ );
not g0402 ( new_n604_, new_n588_ );
not g0403 ( new_n605_, new_n598_ );
nand g0404 ( new_n606_, new_n604_, new_n605_ );
nand g0405 ( new_n607_, new_n606_, new_n599_ );
nand g0406 ( new_n608_, new_n607_, keyIn_0_31 );
nand g0407 ( new_n609_, new_n603_, new_n608_ );
nand g0408 ( new_n610_, new_n577_, new_n609_ );
not g0409 ( new_n611_, new_n610_ );
nor g0410 ( new_n612_, new_n577_, new_n609_ );
nor g0411 ( new_n613_, new_n611_, new_n612_ );
nand g0412 ( new_n614_, new_n613_, new_n545_ );
not g0413 ( new_n615_, new_n614_ );
nor g0414 ( new_n616_, new_n613_, new_n545_ );
nor g0415 ( new_n617_, new_n615_, new_n616_ );
not g0416 ( new_n618_, keyIn_0_20 );
nand g0417 ( new_n619_, N136, N137 );
nand g0418 ( new_n620_, new_n619_, new_n618_ );
not g0419 ( new_n621_, new_n620_ );
nor g0420 ( new_n622_, new_n619_, new_n618_ );
nor g0421 ( new_n623_, new_n621_, new_n622_ );
nand g0422 ( new_n624_, new_n617_, new_n623_ );
not g0423 ( new_n625_, new_n616_ );
nand g0424 ( new_n626_, new_n625_, new_n614_ );
not g0425 ( new_n627_, new_n623_ );
nand g0426 ( new_n628_, new_n626_, new_n627_ );
nand g0427 ( new_n629_, new_n624_, new_n628_ );
nand g0428 ( new_n630_, new_n629_, keyIn_0_54 );
nor g0429 ( new_n631_, new_n629_, keyIn_0_54 );
not g0430 ( new_n632_, new_n631_ );
nand g0431 ( new_n633_, new_n632_, new_n630_ );
nor g0432 ( new_n634_, new_n248_, N93 );
nor g0433 ( new_n635_, new_n217_, N77 );
nor g0434 ( new_n636_, new_n634_, new_n635_ );
not g0435 ( new_n637_, new_n636_ );
nand g0436 ( new_n638_, N109, N125 );
not g0437 ( new_n639_, new_n638_ );
nor g0438 ( new_n640_, N109, N125 );
nor g0439 ( new_n641_, new_n639_, new_n640_ );
not g0440 ( new_n642_, new_n641_ );
nor g0441 ( new_n643_, new_n637_, new_n642_ );
nor g0442 ( new_n644_, new_n636_, new_n641_ );
nor g0443 ( new_n645_, new_n643_, new_n644_ );
not g0444 ( new_n646_, new_n645_ );
nor g0445 ( new_n647_, new_n633_, new_n646_ );
not g0446 ( new_n648_, new_n630_ );
nor g0447 ( new_n649_, new_n648_, new_n631_ );
nor g0448 ( new_n650_, new_n649_, new_n645_ );
nor g0449 ( new_n651_, new_n650_, new_n647_ );
nand g0450 ( new_n652_, new_n651_, keyIn_0_62 );
not g0451 ( new_n653_, keyIn_0_62 );
nand g0452 ( new_n654_, new_n649_, new_n645_ );
nand g0453 ( new_n655_, new_n633_, new_n646_ );
nand g0454 ( new_n656_, new_n654_, new_n655_ );
nand g0455 ( new_n657_, new_n656_, new_n653_ );
nand g0456 ( new_n658_, new_n652_, new_n657_ );
not g0457 ( new_n659_, keyIn_0_30 );
not g0458 ( new_n660_, keyIn_0_5 );
nand g0459 ( new_n661_, new_n372_, N41 );
nand g0460 ( new_n662_, new_n453_, N45 );
nand g0461 ( new_n663_, new_n661_, new_n662_ );
nand g0462 ( new_n664_, new_n663_, new_n660_ );
not g0463 ( new_n665_, new_n664_ );
nor g0464 ( new_n666_, new_n663_, new_n660_ );
nor g0465 ( new_n667_, new_n665_, new_n666_ );
not g0466 ( new_n668_, keyIn_0_4 );
nand g0467 ( new_n669_, N33, N37 );
not g0468 ( new_n670_, new_n669_ );
nor g0469 ( new_n671_, N33, N37 );
nor g0470 ( new_n672_, new_n670_, new_n671_ );
nor g0471 ( new_n673_, new_n672_, new_n668_ );
not g0472 ( new_n674_, N33 );
not g0473 ( new_n675_, N37 );
nand g0474 ( new_n676_, new_n674_, new_n675_ );
nand g0475 ( new_n677_, new_n676_, new_n669_ );
nor g0476 ( new_n678_, new_n677_, keyIn_0_4 );
nor g0477 ( new_n679_, new_n673_, new_n678_ );
nor g0478 ( new_n680_, new_n667_, new_n679_ );
not g0479 ( new_n681_, new_n663_ );
nand g0480 ( new_n682_, new_n681_, keyIn_0_5 );
nand g0481 ( new_n683_, new_n682_, new_n664_ );
nand g0482 ( new_n684_, new_n677_, keyIn_0_4 );
nand g0483 ( new_n685_, new_n672_, new_n668_ );
nand g0484 ( new_n686_, new_n685_, new_n684_ );
nor g0485 ( new_n687_, new_n683_, new_n686_ );
nor g0486 ( new_n688_, new_n680_, new_n687_ );
nand g0487 ( new_n689_, new_n688_, new_n659_ );
nand g0488 ( new_n690_, new_n683_, new_n686_ );
nand g0489 ( new_n691_, new_n667_, new_n679_ );
nand g0490 ( new_n692_, new_n691_, new_n690_ );
nand g0491 ( new_n693_, new_n692_, keyIn_0_30 );
nand g0492 ( new_n694_, new_n689_, new_n693_ );
not g0493 ( new_n695_, keyIn_0_1 );
nand g0494 ( new_n696_, N9, N13 );
not g0495 ( new_n697_, new_n696_ );
nor g0496 ( new_n698_, N9, N13 );
nor g0497 ( new_n699_, new_n697_, new_n698_ );
nand g0498 ( new_n700_, new_n699_, new_n695_ );
not g0499 ( new_n701_, N13 );
nand g0500 ( new_n702_, new_n443_, new_n701_ );
nand g0501 ( new_n703_, new_n702_, new_n696_ );
nand g0502 ( new_n704_, new_n703_, keyIn_0_1 );
nand g0503 ( new_n705_, new_n700_, new_n704_ );
not g0504 ( new_n706_, keyIn_0_0 );
nand g0505 ( new_n707_, N1, N5 );
not g0506 ( new_n708_, new_n707_ );
nor g0507 ( new_n709_, N1, N5 );
nor g0508 ( new_n710_, new_n708_, new_n709_ );
nand g0509 ( new_n711_, new_n710_, new_n706_ );
nand g0510 ( new_n712_, new_n284_, new_n502_ );
nand g0511 ( new_n713_, new_n712_, new_n707_ );
nand g0512 ( new_n714_, new_n713_, keyIn_0_0 );
nand g0513 ( new_n715_, new_n711_, new_n714_ );
nand g0514 ( new_n716_, new_n705_, new_n715_ );
not g0515 ( new_n717_, new_n716_ );
nor g0516 ( new_n718_, new_n705_, new_n715_ );
nor g0517 ( new_n719_, new_n717_, new_n718_ );
nand g0518 ( new_n720_, new_n719_, keyIn_0_28 );
not g0519 ( new_n721_, keyIn_0_28 );
not g0520 ( new_n722_, new_n705_ );
not g0521 ( new_n723_, new_n715_ );
nand g0522 ( new_n724_, new_n722_, new_n723_ );
nand g0523 ( new_n725_, new_n724_, new_n716_ );
nand g0524 ( new_n726_, new_n725_, new_n721_ );
nand g0525 ( new_n727_, new_n720_, new_n726_ );
nand g0526 ( new_n728_, new_n694_, new_n727_ );
not g0527 ( new_n729_, new_n728_ );
nor g0528 ( new_n730_, new_n694_, new_n727_ );
nor g0529 ( new_n731_, new_n729_, new_n730_ );
nor g0530 ( new_n732_, new_n731_, keyIn_0_41 );
not g0531 ( new_n733_, keyIn_0_41 );
nor g0532 ( new_n734_, new_n692_, keyIn_0_30 );
not g0533 ( new_n735_, new_n693_ );
nor g0534 ( new_n736_, new_n735_, new_n734_ );
not g0535 ( new_n737_, new_n727_ );
nand g0536 ( new_n738_, new_n737_, new_n736_ );
nand g0537 ( new_n739_, new_n738_, new_n728_ );
nor g0538 ( new_n740_, new_n739_, new_n733_ );
nor g0539 ( new_n741_, new_n732_, new_n740_ );
nand g0540 ( new_n742_, N135, N137 );
nand g0541 ( new_n743_, new_n742_, keyIn_0_19 );
not g0542 ( new_n744_, new_n743_ );
nor g0543 ( new_n745_, new_n742_, keyIn_0_19 );
nor g0544 ( new_n746_, new_n744_, new_n745_ );
nor g0545 ( new_n747_, new_n741_, new_n746_ );
nand g0546 ( new_n748_, new_n739_, new_n733_ );
nand g0547 ( new_n749_, new_n731_, keyIn_0_41 );
nand g0548 ( new_n750_, new_n749_, new_n748_ );
not g0549 ( new_n751_, new_n746_ );
nor g0550 ( new_n752_, new_n750_, new_n751_ );
nor g0551 ( new_n753_, new_n747_, new_n752_ );
nor g0552 ( new_n754_, new_n753_, keyIn_0_53 );
not g0553 ( new_n755_, keyIn_0_53 );
nand g0554 ( new_n756_, new_n750_, new_n751_ );
nand g0555 ( new_n757_, new_n741_, new_n746_ );
nand g0556 ( new_n758_, new_n757_, new_n756_ );
nor g0557 ( new_n759_, new_n758_, new_n755_ );
nor g0558 ( new_n760_, new_n754_, new_n759_ );
not g0559 ( new_n761_, keyIn_0_38 );
nor g0560 ( new_n762_, new_n402_, N121 );
nor g0561 ( new_n763_, new_n326_, N105 );
nor g0562 ( new_n764_, new_n762_, new_n763_ );
not g0563 ( new_n765_, new_n764_ );
nand g0564 ( new_n766_, new_n765_, keyIn_0_27 );
not g0565 ( new_n767_, new_n766_ );
nor g0566 ( new_n768_, new_n765_, keyIn_0_27 );
nor g0567 ( new_n769_, new_n767_, new_n768_ );
not g0568 ( new_n770_, new_n769_ );
nand g0569 ( new_n771_, N73, N89 );
not g0570 ( new_n772_, new_n771_ );
nor g0571 ( new_n773_, N73, N89 );
nor g0572 ( new_n774_, new_n772_, new_n773_ );
not g0573 ( new_n775_, new_n774_ );
nor g0574 ( new_n776_, new_n775_, keyIn_0_26 );
nand g0575 ( new_n777_, new_n775_, keyIn_0_26 );
not g0576 ( new_n778_, new_n777_ );
nor g0577 ( new_n779_, new_n778_, new_n776_ );
not g0578 ( new_n780_, new_n779_ );
nor g0579 ( new_n781_, new_n770_, new_n780_ );
nor g0580 ( new_n782_, new_n769_, new_n779_ );
nor g0581 ( new_n783_, new_n781_, new_n782_ );
not g0582 ( new_n784_, new_n783_ );
nor g0583 ( new_n785_, new_n784_, new_n761_ );
nor g0584 ( new_n786_, new_n783_, keyIn_0_38 );
nor g0585 ( new_n787_, new_n785_, new_n786_ );
not g0586 ( new_n788_, new_n787_ );
nor g0587 ( new_n789_, new_n760_, new_n788_ );
nand g0588 ( new_n790_, new_n758_, new_n755_ );
nand g0589 ( new_n791_, new_n753_, keyIn_0_53 );
nand g0590 ( new_n792_, new_n791_, new_n790_ );
nor g0591 ( new_n793_, new_n792_, new_n787_ );
nor g0592 ( new_n794_, new_n789_, new_n793_ );
nand g0593 ( new_n795_, new_n794_, keyIn_0_61 );
not g0594 ( new_n796_, keyIn_0_61 );
nand g0595 ( new_n797_, new_n792_, new_n787_ );
nand g0596 ( new_n798_, new_n760_, new_n788_ );
nand g0597 ( new_n799_, new_n798_, new_n797_ );
nand g0598 ( new_n800_, new_n799_, new_n796_ );
nand g0599 ( new_n801_, new_n795_, new_n800_ );
nor g0600 ( new_n802_, new_n658_, new_n801_ );
nand g0601 ( new_n803_, new_n544_, new_n802_ );
not g0602 ( new_n804_, keyIn_0_40 );
nand g0603 ( new_n805_, new_n736_, new_n609_ );
nor g0604 ( new_n806_, new_n607_, keyIn_0_31 );
nor g0605 ( new_n807_, new_n602_, new_n578_ );
nor g0606 ( new_n808_, new_n807_, new_n806_ );
nand g0607 ( new_n809_, new_n808_, new_n694_ );
nand g0608 ( new_n810_, new_n805_, new_n809_ );
nand g0609 ( new_n811_, new_n810_, new_n804_ );
not g0610 ( new_n812_, new_n810_ );
nand g0611 ( new_n813_, new_n812_, keyIn_0_40 );
nand g0612 ( new_n814_, new_n813_, new_n811_ );
not g0613 ( new_n815_, keyIn_0_18 );
nand g0614 ( new_n816_, N134, N137 );
nand g0615 ( new_n817_, new_n816_, new_n815_ );
not g0616 ( new_n818_, new_n817_ );
nor g0617 ( new_n819_, new_n816_, new_n815_ );
nor g0618 ( new_n820_, new_n818_, new_n819_ );
nand g0619 ( new_n821_, new_n814_, new_n820_ );
not g0620 ( new_n822_, new_n811_ );
nor g0621 ( new_n823_, new_n810_, new_n804_ );
nor g0622 ( new_n824_, new_n822_, new_n823_ );
not g0623 ( new_n825_, new_n820_ );
nand g0624 ( new_n826_, new_n824_, new_n825_ );
nand g0625 ( new_n827_, new_n826_, new_n821_ );
nand g0626 ( new_n828_, new_n827_, keyIn_0_52 );
not g0627 ( new_n829_, keyIn_0_52 );
nor g0628 ( new_n830_, new_n824_, new_n825_ );
nor g0629 ( new_n831_, new_n814_, new_n820_ );
nor g0630 ( new_n832_, new_n830_, new_n831_ );
nand g0631 ( new_n833_, new_n832_, new_n829_ );
nand g0632 ( new_n834_, new_n833_, new_n828_ );
nor g0633 ( new_n835_, new_n237_, N85 );
nor g0634 ( new_n836_, new_n206_, N69 );
nor g0635 ( new_n837_, new_n835_, new_n836_ );
not g0636 ( new_n838_, new_n837_ );
nand g0637 ( new_n839_, new_n838_, keyIn_0_24 );
not g0638 ( new_n840_, new_n839_ );
nor g0639 ( new_n841_, new_n838_, keyIn_0_24 );
nor g0640 ( new_n842_, new_n840_, new_n841_ );
not g0641 ( new_n843_, new_n842_ );
nand g0642 ( new_n844_, N101, N117 );
not g0643 ( new_n845_, new_n844_ );
nor g0644 ( new_n846_, N101, N117 );
nor g0645 ( new_n847_, new_n845_, new_n846_ );
not g0646 ( new_n848_, new_n847_ );
nor g0647 ( new_n849_, new_n848_, keyIn_0_25 );
nand g0648 ( new_n850_, new_n848_, keyIn_0_25 );
not g0649 ( new_n851_, new_n850_ );
nor g0650 ( new_n852_, new_n851_, new_n849_ );
not g0651 ( new_n853_, new_n852_ );
nor g0652 ( new_n854_, new_n843_, new_n853_ );
nor g0653 ( new_n855_, new_n842_, new_n852_ );
nor g0654 ( new_n856_, new_n854_, new_n855_ );
not g0655 ( new_n857_, new_n856_ );
nor g0656 ( new_n858_, new_n857_, keyIn_0_37 );
nand g0657 ( new_n859_, new_n857_, keyIn_0_37 );
not g0658 ( new_n860_, new_n859_ );
nor g0659 ( new_n861_, new_n860_, new_n858_ );
not g0660 ( new_n862_, new_n861_ );
nand g0661 ( new_n863_, new_n834_, new_n862_ );
not g0662 ( new_n864_, new_n863_ );
nor g0663 ( new_n865_, new_n834_, new_n862_ );
nor g0664 ( new_n866_, new_n864_, new_n865_ );
nor g0665 ( new_n867_, new_n866_, keyIn_0_60 );
not g0666 ( new_n868_, keyIn_0_60 );
not g0667 ( new_n869_, new_n828_ );
nor g0668 ( new_n870_, new_n827_, keyIn_0_52 );
nor g0669 ( new_n871_, new_n869_, new_n870_ );
nand g0670 ( new_n872_, new_n871_, new_n861_ );
nand g0671 ( new_n873_, new_n872_, new_n863_ );
nor g0672 ( new_n874_, new_n873_, new_n868_ );
nor g0673 ( new_n875_, new_n867_, new_n874_ );
not g0674 ( new_n876_, keyIn_0_59 );
not g0675 ( new_n877_, keyIn_0_51 );
not g0676 ( new_n878_, keyIn_0_39 );
nand g0677 ( new_n879_, new_n577_, new_n727_ );
not g0678 ( new_n880_, new_n879_ );
nor g0679 ( new_n881_, new_n577_, new_n727_ );
nor g0680 ( new_n882_, new_n880_, new_n881_ );
nand g0681 ( new_n883_, new_n882_, new_n878_ );
not g0682 ( new_n884_, new_n577_ );
nand g0683 ( new_n885_, new_n884_, new_n737_ );
nand g0684 ( new_n886_, new_n885_, new_n879_ );
nand g0685 ( new_n887_, new_n886_, keyIn_0_39 );
nand g0686 ( new_n888_, new_n883_, new_n887_ );
not g0687 ( new_n889_, keyIn_0_17 );
nand g0688 ( new_n890_, N133, N137 );
nand g0689 ( new_n891_, new_n890_, new_n889_ );
not g0690 ( new_n892_, new_n891_ );
nor g0691 ( new_n893_, new_n890_, new_n889_ );
nor g0692 ( new_n894_, new_n892_, new_n893_ );
not g0693 ( new_n895_, new_n894_ );
nand g0694 ( new_n896_, new_n888_, new_n895_ );
nor g0695 ( new_n897_, new_n886_, keyIn_0_39 );
nor g0696 ( new_n898_, new_n882_, new_n878_ );
nor g0697 ( new_n899_, new_n898_, new_n897_ );
nand g0698 ( new_n900_, new_n899_, new_n894_ );
nand g0699 ( new_n901_, new_n900_, new_n896_ );
nor g0700 ( new_n902_, new_n901_, new_n877_ );
nor g0701 ( new_n903_, new_n899_, new_n894_ );
nor g0702 ( new_n904_, new_n888_, new_n895_ );
nor g0703 ( new_n905_, new_n903_, new_n904_ );
nor g0704 ( new_n906_, new_n905_, keyIn_0_51 );
nor g0705 ( new_n907_, new_n906_, new_n902_ );
nor g0706 ( new_n908_, new_n235_, N81 );
nor g0707 ( new_n909_, new_n204_, N65 );
nor g0708 ( new_n910_, new_n908_, new_n909_ );
not g0709 ( new_n911_, new_n910_ );
nand g0710 ( new_n912_, N97, N113 );
not g0711 ( new_n913_, new_n912_ );
nor g0712 ( new_n914_, N97, N113 );
nor g0713 ( new_n915_, new_n913_, new_n914_ );
not g0714 ( new_n916_, new_n915_ );
nor g0715 ( new_n917_, new_n911_, new_n916_ );
nor g0716 ( new_n918_, new_n910_, new_n915_ );
nor g0717 ( new_n919_, new_n917_, new_n918_ );
nor g0718 ( new_n920_, new_n907_, new_n919_ );
nand g0719 ( new_n921_, new_n905_, keyIn_0_51 );
nand g0720 ( new_n922_, new_n901_, new_n877_ );
nand g0721 ( new_n923_, new_n921_, new_n922_ );
not g0722 ( new_n924_, new_n919_ );
nor g0723 ( new_n925_, new_n923_, new_n924_ );
nor g0724 ( new_n926_, new_n920_, new_n925_ );
nand g0725 ( new_n927_, new_n926_, new_n876_ );
nand g0726 ( new_n928_, new_n923_, new_n924_ );
nand g0727 ( new_n929_, new_n907_, new_n919_ );
nand g0728 ( new_n930_, new_n929_, new_n928_ );
nand g0729 ( new_n931_, new_n930_, keyIn_0_59 );
nand g0730 ( new_n932_, new_n927_, new_n931_ );
nand g0731 ( new_n933_, new_n875_, new_n932_ );
nor g0732 ( new_n934_, new_n803_, new_n933_ );
not g0733 ( new_n935_, new_n934_ );
nor g0734 ( new_n936_, new_n935_, new_n312_ );
not g0735 ( new_n937_, new_n936_ );
nand g0736 ( new_n938_, new_n937_, N1 );
nand g0737 ( new_n939_, new_n936_, new_n284_ );
nand g0738 ( N724, new_n938_, new_n939_ );
nor g0739 ( new_n941_, new_n935_, new_n526_ );
not g0740 ( new_n942_, new_n941_ );
nand g0741 ( new_n943_, new_n942_, N5 );
nand g0742 ( new_n944_, new_n941_, new_n502_ );
nand g0743 ( N725, new_n943_, new_n944_ );
nor g0744 ( new_n946_, new_n935_, new_n482_ );
not g0745 ( new_n947_, new_n946_ );
nand g0746 ( new_n948_, new_n947_, N9 );
nand g0747 ( new_n949_, new_n946_, new_n443_ );
nand g0748 ( N726, new_n948_, new_n949_ );
not g0749 ( new_n951_, new_n389_ );
nor g0750 ( new_n952_, new_n935_, new_n951_ );
not g0751 ( new_n953_, new_n952_ );
nand g0752 ( new_n954_, new_n953_, N13 );
nand g0753 ( new_n955_, new_n952_, new_n701_ );
nand g0754 ( N727, new_n954_, new_n955_ );
not g0755 ( new_n957_, keyIn_0_105 );
not g0756 ( new_n958_, keyIn_0_82 );
nand g0757 ( new_n959_, new_n658_, new_n801_ );
not g0758 ( new_n960_, new_n959_ );
nand g0759 ( new_n961_, new_n544_, new_n960_ );
nor g0760 ( new_n962_, new_n961_, new_n933_ );
nand g0761 ( new_n963_, new_n962_, keyIn_0_76 );
not g0762 ( new_n964_, keyIn_0_76 );
nand g0763 ( new_n965_, new_n873_, new_n868_ );
nand g0764 ( new_n966_, new_n866_, keyIn_0_60 );
nand g0765 ( new_n967_, new_n966_, new_n965_ );
nor g0766 ( new_n968_, new_n930_, keyIn_0_59 );
nor g0767 ( new_n969_, new_n926_, new_n876_ );
nor g0768 ( new_n970_, new_n969_, new_n968_ );
nor g0769 ( new_n971_, new_n970_, new_n967_ );
nor g0770 ( new_n972_, new_n533_, new_n528_ );
not g0771 ( new_n973_, new_n543_ );
nor g0772 ( new_n974_, new_n973_, new_n972_ );
nor g0773 ( new_n975_, new_n974_, new_n959_ );
nand g0774 ( new_n976_, new_n975_, new_n971_ );
nand g0775 ( new_n977_, new_n976_, new_n964_ );
nand g0776 ( new_n978_, new_n963_, new_n977_ );
nand g0777 ( new_n979_, new_n978_, new_n311_ );
nand g0778 ( new_n980_, new_n979_, new_n958_ );
not g0779 ( new_n981_, new_n980_ );
nor g0780 ( new_n982_, new_n979_, new_n958_ );
nor g0781 ( new_n983_, new_n981_, new_n982_ );
nor g0782 ( new_n984_, new_n983_, N17 );
not g0783 ( new_n985_, new_n979_ );
nand g0784 ( new_n986_, new_n985_, keyIn_0_82 );
nand g0785 ( new_n987_, new_n986_, new_n980_ );
nor g0786 ( new_n988_, new_n987_, new_n286_ );
nor g0787 ( new_n989_, new_n984_, new_n988_ );
nand g0788 ( new_n990_, new_n989_, new_n957_ );
nand g0789 ( new_n991_, new_n987_, new_n286_ );
nand g0790 ( new_n992_, new_n983_, N17 );
nand g0791 ( new_n993_, new_n992_, new_n991_ );
nand g0792 ( new_n994_, new_n993_, keyIn_0_105 );
nand g0793 ( N728, new_n990_, new_n994_ );
not g0794 ( new_n996_, keyIn_0_106 );
not g0795 ( new_n997_, keyIn_0_83 );
not g0796 ( new_n998_, new_n526_ );
nand g0797 ( new_n999_, new_n978_, new_n998_ );
nand g0798 ( new_n1000_, new_n999_, new_n997_ );
not g0799 ( new_n1001_, new_n1000_ );
nor g0800 ( new_n1002_, new_n999_, new_n997_ );
nor g0801 ( new_n1003_, new_n1001_, new_n1002_ );
nor g0802 ( new_n1004_, new_n1003_, new_n504_ );
not g0803 ( new_n1005_, new_n999_ );
nand g0804 ( new_n1006_, new_n1005_, keyIn_0_83 );
nand g0805 ( new_n1007_, new_n1006_, new_n1000_ );
nor g0806 ( new_n1008_, new_n1007_, N21 );
nor g0807 ( new_n1009_, new_n1004_, new_n1008_ );
nand g0808 ( new_n1010_, new_n1009_, new_n996_ );
nand g0809 ( new_n1011_, new_n1007_, N21 );
nand g0810 ( new_n1012_, new_n1003_, new_n504_ );
nand g0811 ( new_n1013_, new_n1012_, new_n1011_ );
nand g0812 ( new_n1014_, new_n1013_, keyIn_0_106 );
nand g0813 ( N729, new_n1010_, new_n1014_ );
nand g0814 ( new_n1016_, new_n978_, new_n537_ );
not g0815 ( new_n1017_, new_n1016_ );
nand g0816 ( new_n1018_, new_n1017_, new_n445_ );
nand g0817 ( new_n1019_, new_n1016_, N25 );
nand g0818 ( N730, new_n1018_, new_n1019_ );
not g0819 ( new_n1021_, N29 );
not g0820 ( new_n1022_, keyIn_0_84 );
nand g0821 ( new_n1023_, new_n978_, new_n389_ );
nand g0822 ( new_n1024_, new_n1023_, new_n1022_ );
not g0823 ( new_n1025_, new_n1024_ );
nor g0824 ( new_n1026_, new_n1023_, new_n1022_ );
nor g0825 ( new_n1027_, new_n1025_, new_n1026_ );
nor g0826 ( new_n1028_, new_n1027_, new_n1021_ );
not g0827 ( new_n1029_, new_n1023_ );
nand g0828 ( new_n1030_, new_n1029_, keyIn_0_84 );
nand g0829 ( new_n1031_, new_n1030_, new_n1024_ );
nor g0830 ( new_n1032_, new_n1031_, N29 );
nor g0831 ( new_n1033_, new_n1028_, new_n1032_ );
nand g0832 ( new_n1034_, new_n1033_, keyIn_0_107 );
not g0833 ( new_n1035_, keyIn_0_107 );
nand g0834 ( new_n1036_, new_n1031_, N29 );
nand g0835 ( new_n1037_, new_n1027_, new_n1021_ );
nand g0836 ( new_n1038_, new_n1037_, new_n1036_ );
nand g0837 ( new_n1039_, new_n1038_, new_n1035_ );
nand g0838 ( N731, new_n1034_, new_n1039_ );
not g0839 ( new_n1041_, keyIn_0_108 );
not g0840 ( new_n1042_, keyIn_0_85 );
nand g0841 ( new_n1043_, new_n970_, new_n967_ );
nor g0842 ( new_n1044_, new_n803_, new_n1043_ );
nand g0843 ( new_n1045_, new_n1044_, keyIn_0_77 );
not g0844 ( new_n1046_, keyIn_0_77 );
nor g0845 ( new_n1047_, new_n656_, new_n653_ );
not g0846 ( new_n1048_, new_n657_ );
nor g0847 ( new_n1049_, new_n1048_, new_n1047_ );
nor g0848 ( new_n1050_, new_n799_, new_n796_ );
nor g0849 ( new_n1051_, new_n794_, keyIn_0_61 );
nor g0850 ( new_n1052_, new_n1051_, new_n1050_ );
nand g0851 ( new_n1053_, new_n1049_, new_n1052_ );
nor g0852 ( new_n1054_, new_n974_, new_n1053_ );
nor g0853 ( new_n1055_, new_n875_, new_n932_ );
nand g0854 ( new_n1056_, new_n1054_, new_n1055_ );
nand g0855 ( new_n1057_, new_n1056_, new_n1046_ );
nand g0856 ( new_n1058_, new_n1045_, new_n1057_ );
nand g0857 ( new_n1059_, new_n1058_, new_n311_ );
nand g0858 ( new_n1060_, new_n1059_, new_n1042_ );
not g0859 ( new_n1061_, new_n1060_ );
nor g0860 ( new_n1062_, new_n1059_, new_n1042_ );
nor g0861 ( new_n1063_, new_n1061_, new_n1062_ );
nor g0862 ( new_n1064_, new_n1063_, N33 );
not g0863 ( new_n1065_, new_n1059_ );
nand g0864 ( new_n1066_, new_n1065_, keyIn_0_85 );
nand g0865 ( new_n1067_, new_n1066_, new_n1060_ );
nor g0866 ( new_n1068_, new_n1067_, new_n674_ );
nor g0867 ( new_n1069_, new_n1064_, new_n1068_ );
nand g0868 ( new_n1070_, new_n1069_, new_n1041_ );
nand g0869 ( new_n1071_, new_n1067_, new_n674_ );
nand g0870 ( new_n1072_, new_n1063_, N33 );
nand g0871 ( new_n1073_, new_n1072_, new_n1071_ );
nand g0872 ( new_n1074_, new_n1073_, keyIn_0_108 );
nand g0873 ( N732, new_n1070_, new_n1074_ );
not g0874 ( new_n1076_, keyIn_0_86 );
nand g0875 ( new_n1077_, new_n1058_, new_n998_ );
nand g0876 ( new_n1078_, new_n1077_, new_n1076_ );
not g0877 ( new_n1079_, new_n1078_ );
nor g0878 ( new_n1080_, new_n1077_, new_n1076_ );
nor g0879 ( new_n1081_, new_n1079_, new_n1080_ );
nor g0880 ( new_n1082_, new_n1081_, new_n675_ );
not g0881 ( new_n1083_, new_n1077_ );
nand g0882 ( new_n1084_, new_n1083_, keyIn_0_86 );
nand g0883 ( new_n1085_, new_n1084_, new_n1078_ );
nor g0884 ( new_n1086_, new_n1085_, N37 );
nor g0885 ( new_n1087_, new_n1082_, new_n1086_ );
nand g0886 ( new_n1088_, new_n1087_, keyIn_0_109 );
not g0887 ( new_n1089_, keyIn_0_109 );
nand g0888 ( new_n1090_, new_n1085_, N37 );
nand g0889 ( new_n1091_, new_n1081_, new_n675_ );
nand g0890 ( new_n1092_, new_n1091_, new_n1090_ );
nand g0891 ( new_n1093_, new_n1092_, new_n1089_ );
nand g0892 ( N733, new_n1088_, new_n1093_ );
not g0893 ( new_n1095_, keyIn_0_110 );
not g0894 ( new_n1096_, keyIn_0_87 );
nand g0895 ( new_n1097_, new_n1058_, new_n537_ );
nand g0896 ( new_n1098_, new_n1097_, new_n1096_ );
not g0897 ( new_n1099_, new_n1098_ );
nor g0898 ( new_n1100_, new_n1097_, new_n1096_ );
nor g0899 ( new_n1101_, new_n1099_, new_n1100_ );
nor g0900 ( new_n1102_, new_n1101_, N41 );
not g0901 ( new_n1103_, new_n1097_ );
nand g0902 ( new_n1104_, new_n1103_, keyIn_0_87 );
nand g0903 ( new_n1105_, new_n1104_, new_n1098_ );
nor g0904 ( new_n1106_, new_n1105_, new_n453_ );
nor g0905 ( new_n1107_, new_n1102_, new_n1106_ );
nand g0906 ( new_n1108_, new_n1107_, new_n1095_ );
nand g0907 ( new_n1109_, new_n1105_, new_n453_ );
nand g0908 ( new_n1110_, new_n1101_, N41 );
nand g0909 ( new_n1111_, new_n1110_, new_n1109_ );
nand g0910 ( new_n1112_, new_n1111_, keyIn_0_110 );
nand g0911 ( N734, new_n1108_, new_n1112_ );
not g0912 ( new_n1114_, keyIn_0_111 );
not g0913 ( new_n1115_, keyIn_0_88 );
nand g0914 ( new_n1116_, new_n1058_, new_n389_ );
nand g0915 ( new_n1117_, new_n1116_, new_n1115_ );
not g0916 ( new_n1118_, new_n1117_ );
nor g0917 ( new_n1119_, new_n1116_, new_n1115_ );
nor g0918 ( new_n1120_, new_n1118_, new_n1119_ );
nor g0919 ( new_n1121_, new_n1120_, N45 );
not g0920 ( new_n1122_, new_n1116_ );
nand g0921 ( new_n1123_, new_n1122_, keyIn_0_88 );
nand g0922 ( new_n1124_, new_n1123_, new_n1117_ );
nor g0923 ( new_n1125_, new_n1124_, new_n372_ );
nor g0924 ( new_n1126_, new_n1121_, new_n1125_ );
nand g0925 ( new_n1127_, new_n1126_, new_n1114_ );
nand g0926 ( new_n1128_, new_n1124_, new_n372_ );
nand g0927 ( new_n1129_, new_n1120_, N45 );
nand g0928 ( new_n1130_, new_n1129_, new_n1128_ );
nand g0929 ( new_n1131_, new_n1130_, keyIn_0_111 );
nand g0930 ( N735, new_n1127_, new_n1131_ );
nor g0931 ( new_n1133_, new_n961_, new_n1043_ );
not g0932 ( new_n1134_, new_n1133_ );
nor g0933 ( new_n1135_, new_n1134_, new_n312_ );
not g0934 ( new_n1136_, new_n1135_ );
nand g0935 ( new_n1137_, new_n1136_, N49 );
not g0936 ( new_n1138_, N49 );
nand g0937 ( new_n1139_, new_n1135_, new_n1138_ );
nand g0938 ( N736, new_n1137_, new_n1139_ );
nor g0939 ( new_n1141_, new_n1134_, new_n526_ );
not g0940 ( new_n1142_, new_n1141_ );
nand g0941 ( new_n1143_, new_n1142_, N53 );
not g0942 ( new_n1144_, N53 );
nand g0943 ( new_n1145_, new_n1141_, new_n1144_ );
nand g0944 ( N737, new_n1143_, new_n1145_ );
nor g0945 ( new_n1147_, new_n1134_, new_n482_ );
not g0946 ( new_n1148_, new_n1147_ );
nand g0947 ( new_n1149_, new_n1148_, N57 );
nand g0948 ( new_n1150_, new_n1147_, new_n455_ );
nand g0949 ( N738, new_n1149_, new_n1150_ );
nor g0950 ( new_n1152_, new_n1134_, new_n951_ );
not g0951 ( new_n1153_, new_n1152_ );
nand g0952 ( new_n1154_, new_n1153_, N61 );
nand g0953 ( new_n1155_, new_n1152_, new_n374_ );
nand g0954 ( N739, new_n1154_, new_n1155_ );
not g0955 ( new_n1157_, keyIn_0_112 );
not g0956 ( new_n1158_, keyIn_0_78 );
not g0957 ( new_n1159_, keyIn_0_75 );
nor g0958 ( new_n1160_, new_n933_, new_n658_ );
not g0959 ( new_n1161_, keyIn_0_66 );
nor g0960 ( new_n1162_, new_n801_, new_n1161_ );
nand g0961 ( new_n1163_, new_n801_, new_n1161_ );
not g0962 ( new_n1164_, new_n1163_ );
nor g0963 ( new_n1165_, new_n1164_, new_n1162_ );
nand g0964 ( new_n1166_, new_n1165_, new_n1160_ );
nand g0965 ( new_n1167_, new_n1166_, keyIn_0_74 );
not g0966 ( new_n1168_, keyIn_0_74 );
nand g0967 ( new_n1169_, new_n971_, new_n1049_ );
nand g0968 ( new_n1170_, new_n1052_, keyIn_0_66 );
nand g0969 ( new_n1171_, new_n1170_, new_n1163_ );
nor g0970 ( new_n1172_, new_n1169_, new_n1171_ );
nand g0971 ( new_n1173_, new_n1172_, new_n1168_ );
nand g0972 ( new_n1174_, new_n1167_, new_n1173_ );
nor g0973 ( new_n1175_, new_n967_, new_n932_ );
nand g0974 ( new_n1176_, new_n802_, new_n1175_ );
nand g0975 ( new_n1177_, new_n1176_, keyIn_0_72 );
not g0976 ( new_n1178_, keyIn_0_72 );
not g0977 ( new_n1179_, new_n1176_ );
nand g0978 ( new_n1180_, new_n1179_, new_n1178_ );
nand g0979 ( new_n1181_, new_n1180_, new_n1177_ );
nand g0980 ( new_n1182_, new_n1174_, new_n1181_ );
not g0981 ( new_n1183_, new_n1182_ );
not g0982 ( new_n1184_, keyIn_0_71 );
not g0983 ( new_n1185_, keyIn_0_64 );
nand g0984 ( new_n1186_, new_n801_, new_n1185_ );
nand g0985 ( new_n1187_, new_n1186_, new_n658_ );
nand g0986 ( new_n1188_, new_n1052_, keyIn_0_64 );
nand g0987 ( new_n1189_, new_n1188_, new_n1175_ );
nor g0988 ( new_n1190_, new_n1189_, new_n1187_ );
nor g0989 ( new_n1191_, new_n1190_, new_n1184_ );
not g0990 ( new_n1192_, new_n1187_ );
nand g0991 ( new_n1193_, new_n875_, new_n970_ );
nor g0992 ( new_n1194_, new_n801_, new_n1185_ );
nor g0993 ( new_n1195_, new_n1193_, new_n1194_ );
nand g0994 ( new_n1196_, new_n1195_, new_n1192_ );
nor g0995 ( new_n1197_, new_n1196_, keyIn_0_71 );
nor g0996 ( new_n1198_, new_n1197_, new_n1191_ );
not g0997 ( new_n1199_, keyIn_0_73 );
nand g0998 ( new_n1200_, new_n801_, keyIn_0_65 );
not g0999 ( new_n1201_, keyIn_0_65 );
nand g1000 ( new_n1202_, new_n1052_, new_n1201_ );
nand g1001 ( new_n1203_, new_n1202_, new_n1200_ );
nor g1002 ( new_n1204_, new_n1043_, new_n658_ );
nand g1003 ( new_n1205_, new_n1204_, new_n1203_ );
nand g1004 ( new_n1206_, new_n1205_, new_n1199_ );
not g1005 ( new_n1207_, new_n1206_ );
nor g1006 ( new_n1208_, new_n1205_, new_n1199_ );
nor g1007 ( new_n1209_, new_n1207_, new_n1208_ );
nor g1008 ( new_n1210_, new_n1209_, new_n1198_ );
nand g1009 ( new_n1211_, new_n1210_, new_n1183_ );
nand g1010 ( new_n1212_, new_n1211_, new_n1159_ );
nand g1011 ( new_n1213_, new_n1196_, keyIn_0_71 );
nand g1012 ( new_n1214_, new_n1190_, new_n1184_ );
nand g1013 ( new_n1215_, new_n1213_, new_n1214_ );
not g1014 ( new_n1216_, new_n1200_ );
nor g1015 ( new_n1217_, new_n801_, keyIn_0_65 );
nor g1016 ( new_n1218_, new_n1216_, new_n1217_ );
nand g1017 ( new_n1219_, new_n1055_, new_n1049_ );
nor g1018 ( new_n1220_, new_n1218_, new_n1219_ );
nand g1019 ( new_n1221_, new_n1220_, keyIn_0_73 );
nand g1020 ( new_n1222_, new_n1221_, new_n1206_ );
nand g1021 ( new_n1223_, new_n1222_, new_n1215_ );
nor g1022 ( new_n1224_, new_n1223_, new_n1182_ );
nand g1023 ( new_n1225_, new_n1224_, keyIn_0_75 );
nand g1024 ( new_n1226_, new_n1212_, new_n1225_ );
not g1025 ( new_n1227_, keyIn_0_67 );
nor g1026 ( new_n1228_, new_n998_, new_n1227_ );
nor g1027 ( new_n1229_, new_n526_, keyIn_0_67 );
nor g1028 ( new_n1230_, new_n1228_, new_n1229_ );
nor g1029 ( new_n1231_, new_n312_, new_n389_ );
nand g1030 ( new_n1232_, new_n1231_, new_n537_ );
nor g1031 ( new_n1233_, new_n1232_, new_n1230_ );
nand g1032 ( new_n1234_, new_n1226_, new_n1233_ );
nand g1033 ( new_n1235_, new_n1234_, new_n1158_ );
not g1034 ( new_n1236_, new_n1235_ );
nor g1035 ( new_n1237_, new_n1234_, new_n1158_ );
nor g1036 ( new_n1238_, new_n1236_, new_n1237_ );
nor g1037 ( new_n1239_, new_n1238_, new_n970_ );
nor g1038 ( new_n1240_, new_n1239_, keyIn_0_89 );
not g1039 ( new_n1241_, keyIn_0_89 );
not g1040 ( new_n1242_, new_n1237_ );
nand g1041 ( new_n1243_, new_n1242_, new_n1235_ );
nand g1042 ( new_n1244_, new_n1243_, new_n932_ );
nor g1043 ( new_n1245_, new_n1244_, new_n1241_ );
nor g1044 ( new_n1246_, new_n1240_, new_n1245_ );
nor g1045 ( new_n1247_, new_n1246_, N65 );
nand g1046 ( new_n1248_, new_n1244_, new_n1241_ );
nand g1047 ( new_n1249_, new_n1239_, keyIn_0_89 );
nand g1048 ( new_n1250_, new_n1249_, new_n1248_ );
nor g1049 ( new_n1251_, new_n1250_, new_n235_ );
nor g1050 ( new_n1252_, new_n1247_, new_n1251_ );
nand g1051 ( new_n1253_, new_n1252_, new_n1157_ );
nand g1052 ( new_n1254_, new_n1250_, new_n235_ );
nand g1053 ( new_n1255_, new_n1246_, N65 );
nand g1054 ( new_n1256_, new_n1255_, new_n1254_ );
nand g1055 ( new_n1257_, new_n1256_, keyIn_0_112 );
nand g1056 ( N740, new_n1253_, new_n1257_ );
not g1057 ( new_n1259_, keyIn_0_113 );
nor g1058 ( new_n1260_, new_n1238_, new_n875_ );
nor g1059 ( new_n1261_, new_n1260_, keyIn_0_90 );
not g1060 ( new_n1262_, keyIn_0_90 );
nand g1061 ( new_n1263_, new_n1243_, new_n967_ );
nor g1062 ( new_n1264_, new_n1263_, new_n1262_ );
nor g1063 ( new_n1265_, new_n1261_, new_n1264_ );
nor g1064 ( new_n1266_, new_n1265_, N69 );
nand g1065 ( new_n1267_, new_n1263_, new_n1262_ );
nand g1066 ( new_n1268_, new_n1260_, keyIn_0_90 );
nand g1067 ( new_n1269_, new_n1268_, new_n1267_ );
nor g1068 ( new_n1270_, new_n1269_, new_n237_ );
nor g1069 ( new_n1271_, new_n1266_, new_n1270_ );
nand g1070 ( new_n1272_, new_n1271_, new_n1259_ );
nand g1071 ( new_n1273_, new_n1269_, new_n237_ );
nand g1072 ( new_n1274_, new_n1265_, N69 );
nand g1073 ( new_n1275_, new_n1274_, new_n1273_ );
nand g1074 ( new_n1276_, new_n1275_, keyIn_0_113 );
nand g1075 ( N741, new_n1272_, new_n1276_ );
nor g1076 ( new_n1278_, new_n1238_, new_n801_ );
nor g1077 ( new_n1279_, new_n1278_, keyIn_0_91 );
not g1078 ( new_n1280_, keyIn_0_91 );
nand g1079 ( new_n1281_, new_n1243_, new_n1052_ );
nor g1080 ( new_n1282_, new_n1281_, new_n1280_ );
nor g1081 ( new_n1283_, new_n1279_, new_n1282_ );
nor g1082 ( new_n1284_, new_n1283_, new_n246_ );
nand g1083 ( new_n1285_, new_n1281_, new_n1280_ );
nand g1084 ( new_n1286_, new_n1278_, keyIn_0_91 );
nand g1085 ( new_n1287_, new_n1286_, new_n1285_ );
nor g1086 ( new_n1288_, new_n1287_, N73 );
nor g1087 ( new_n1289_, new_n1284_, new_n1288_ );
nand g1088 ( new_n1290_, new_n1289_, keyIn_0_114 );
not g1089 ( new_n1291_, keyIn_0_114 );
nand g1090 ( new_n1292_, new_n1287_, N73 );
nand g1091 ( new_n1293_, new_n1283_, new_n246_ );
nand g1092 ( new_n1294_, new_n1293_, new_n1292_ );
nand g1093 ( new_n1295_, new_n1294_, new_n1291_ );
nand g1094 ( N742, new_n1290_, new_n1295_ );
not g1095 ( new_n1297_, keyIn_0_115 );
nor g1096 ( new_n1298_, new_n1238_, new_n1049_ );
nor g1097 ( new_n1299_, new_n1298_, keyIn_0_92 );
not g1098 ( new_n1300_, keyIn_0_92 );
nand g1099 ( new_n1301_, new_n1243_, new_n658_ );
nor g1100 ( new_n1302_, new_n1301_, new_n1300_ );
nor g1101 ( new_n1303_, new_n1299_, new_n1302_ );
nor g1102 ( new_n1304_, new_n1303_, new_n248_ );
nand g1103 ( new_n1305_, new_n1301_, new_n1300_ );
nand g1104 ( new_n1306_, new_n1298_, keyIn_0_92 );
nand g1105 ( new_n1307_, new_n1306_, new_n1305_ );
nor g1106 ( new_n1308_, new_n1307_, N77 );
nor g1107 ( new_n1309_, new_n1304_, new_n1308_ );
nand g1108 ( new_n1310_, new_n1309_, new_n1297_ );
nand g1109 ( new_n1311_, new_n1307_, N77 );
nand g1110 ( new_n1312_, new_n1303_, new_n248_ );
nand g1111 ( new_n1313_, new_n1312_, new_n1311_ );
nand g1112 ( new_n1314_, new_n1313_, keyIn_0_115 );
nand g1113 ( N743, new_n1310_, new_n1314_ );
not g1114 ( new_n1316_, keyIn_0_116 );
nand g1115 ( new_n1317_, new_n537_, keyIn_0_68 );
not g1116 ( new_n1318_, keyIn_0_68 );
nand g1117 ( new_n1319_, new_n482_, new_n1318_ );
nand g1118 ( new_n1320_, new_n1317_, new_n1319_ );
nor g1119 ( new_n1321_, new_n541_, new_n951_ );
nand g1120 ( new_n1322_, new_n1321_, new_n1320_ );
not g1121 ( new_n1323_, new_n1322_ );
nand g1122 ( new_n1324_, new_n1226_, new_n1323_ );
nand g1123 ( new_n1325_, new_n1324_, keyIn_0_79 );
not g1124 ( new_n1326_, new_n1325_ );
nor g1125 ( new_n1327_, new_n1324_, keyIn_0_79 );
nor g1126 ( new_n1328_, new_n1326_, new_n1327_ );
nor g1127 ( new_n1329_, new_n1328_, new_n970_ );
nor g1128 ( new_n1330_, new_n1329_, keyIn_0_93 );
not g1129 ( new_n1331_, keyIn_0_93 );
not g1130 ( new_n1332_, new_n1327_ );
nand g1131 ( new_n1333_, new_n1332_, new_n1325_ );
nand g1132 ( new_n1334_, new_n1333_, new_n932_ );
nor g1133 ( new_n1335_, new_n1334_, new_n1331_ );
nor g1134 ( new_n1336_, new_n1330_, new_n1335_ );
nor g1135 ( new_n1337_, new_n1336_, N81 );
nand g1136 ( new_n1338_, new_n1334_, new_n1331_ );
nand g1137 ( new_n1339_, new_n1329_, keyIn_0_93 );
nand g1138 ( new_n1340_, new_n1339_, new_n1338_ );
nor g1139 ( new_n1341_, new_n1340_, new_n204_ );
nor g1140 ( new_n1342_, new_n1337_, new_n1341_ );
nand g1141 ( new_n1343_, new_n1342_, new_n1316_ );
nand g1142 ( new_n1344_, new_n1340_, new_n204_ );
nand g1143 ( new_n1345_, new_n1336_, N81 );
nand g1144 ( new_n1346_, new_n1345_, new_n1344_ );
nand g1145 ( new_n1347_, new_n1346_, keyIn_0_116 );
nand g1146 ( N744, new_n1343_, new_n1347_ );
not g1147 ( new_n1349_, keyIn_0_117 );
not g1148 ( new_n1350_, keyIn_0_94 );
nor g1149 ( new_n1351_, new_n1328_, new_n875_ );
nor g1150 ( new_n1352_, new_n1351_, new_n1350_ );
nand g1151 ( new_n1353_, new_n1333_, new_n967_ );
nor g1152 ( new_n1354_, new_n1353_, keyIn_0_94 );
nor g1153 ( new_n1355_, new_n1352_, new_n1354_ );
nor g1154 ( new_n1356_, new_n1355_, N85 );
nand g1155 ( new_n1357_, new_n1353_, keyIn_0_94 );
nand g1156 ( new_n1358_, new_n1351_, new_n1350_ );
nand g1157 ( new_n1359_, new_n1358_, new_n1357_ );
nor g1158 ( new_n1360_, new_n1359_, new_n206_ );
nor g1159 ( new_n1361_, new_n1356_, new_n1360_ );
nand g1160 ( new_n1362_, new_n1361_, new_n1349_ );
nand g1161 ( new_n1363_, new_n1359_, new_n206_ );
nand g1162 ( new_n1364_, new_n1355_, N85 );
nand g1163 ( new_n1365_, new_n1364_, new_n1363_ );
nand g1164 ( new_n1366_, new_n1365_, keyIn_0_117 );
nand g1165 ( N745, new_n1362_, new_n1366_ );
nor g1166 ( new_n1368_, new_n1328_, new_n801_ );
nor g1167 ( new_n1369_, new_n1368_, keyIn_0_95 );
not g1168 ( new_n1370_, keyIn_0_95 );
nand g1169 ( new_n1371_, new_n1333_, new_n1052_ );
nor g1170 ( new_n1372_, new_n1371_, new_n1370_ );
nor g1171 ( new_n1373_, new_n1369_, new_n1372_ );
nor g1172 ( new_n1374_, new_n1373_, new_n215_ );
nand g1173 ( new_n1375_, new_n1371_, new_n1370_ );
nand g1174 ( new_n1376_, new_n1368_, keyIn_0_95 );
nand g1175 ( new_n1377_, new_n1376_, new_n1375_ );
nor g1176 ( new_n1378_, new_n1377_, N89 );
nor g1177 ( new_n1379_, new_n1374_, new_n1378_ );
nand g1178 ( new_n1380_, new_n1379_, keyIn_0_118 );
not g1179 ( new_n1381_, keyIn_0_118 );
nand g1180 ( new_n1382_, new_n1377_, N89 );
nand g1181 ( new_n1383_, new_n1373_, new_n215_ );
nand g1182 ( new_n1384_, new_n1383_, new_n1382_ );
nand g1183 ( new_n1385_, new_n1384_, new_n1381_ );
nand g1184 ( N746, new_n1380_, new_n1385_ );
nor g1185 ( new_n1387_, new_n1328_, new_n1049_ );
nor g1186 ( new_n1388_, new_n1387_, keyIn_0_96 );
not g1187 ( new_n1389_, keyIn_0_96 );
nand g1188 ( new_n1390_, new_n1333_, new_n658_ );
nor g1189 ( new_n1391_, new_n1390_, new_n1389_ );
nor g1190 ( new_n1392_, new_n1388_, new_n1391_ );
nor g1191 ( new_n1393_, new_n1392_, new_n217_ );
nand g1192 ( new_n1394_, new_n1390_, new_n1389_ );
nand g1193 ( new_n1395_, new_n1387_, keyIn_0_96 );
nand g1194 ( new_n1396_, new_n1395_, new_n1394_ );
nor g1195 ( new_n1397_, new_n1396_, N93 );
nor g1196 ( new_n1398_, new_n1393_, new_n1397_ );
nand g1197 ( new_n1399_, new_n1398_, keyIn_0_119 );
not g1198 ( new_n1400_, keyIn_0_119 );
nand g1199 ( new_n1401_, new_n1396_, N93 );
nand g1200 ( new_n1402_, new_n1392_, new_n217_ );
nand g1201 ( new_n1403_, new_n1402_, new_n1401_ );
nand g1202 ( new_n1404_, new_n1403_, new_n1400_ );
nand g1203 ( N747, new_n1399_, new_n1404_ );
not g1204 ( new_n1406_, keyIn_0_120 );
not g1205 ( new_n1407_, keyIn_0_80 );
nor g1206 ( new_n1408_, new_n311_, new_n389_ );
nand g1207 ( new_n1409_, new_n1408_, new_n531_ );
not g1208 ( new_n1410_, new_n1409_ );
nand g1209 ( new_n1411_, new_n1226_, new_n1410_ );
nand g1210 ( new_n1412_, new_n1411_, new_n1407_ );
not g1211 ( new_n1413_, new_n1412_ );
nor g1212 ( new_n1414_, new_n1411_, new_n1407_ );
nor g1213 ( new_n1415_, new_n1413_, new_n1414_ );
nor g1214 ( new_n1416_, new_n1415_, new_n970_ );
nor g1215 ( new_n1417_, new_n1416_, keyIn_0_97 );
not g1216 ( new_n1418_, keyIn_0_97 );
not g1217 ( new_n1419_, new_n1414_ );
nand g1218 ( new_n1420_, new_n1419_, new_n1412_ );
nand g1219 ( new_n1421_, new_n1420_, new_n932_ );
nor g1220 ( new_n1422_, new_n1421_, new_n1418_ );
nor g1221 ( new_n1423_, new_n1417_, new_n1422_ );
nor g1222 ( new_n1424_, new_n1423_, new_n391_ );
nand g1223 ( new_n1425_, new_n1421_, new_n1418_ );
nand g1224 ( new_n1426_, new_n1416_, keyIn_0_97 );
nand g1225 ( new_n1427_, new_n1426_, new_n1425_ );
nor g1226 ( new_n1428_, new_n1427_, N97 );
nor g1227 ( new_n1429_, new_n1424_, new_n1428_ );
nand g1228 ( new_n1430_, new_n1429_, new_n1406_ );
nand g1229 ( new_n1431_, new_n1427_, N97 );
nand g1230 ( new_n1432_, new_n1423_, new_n391_ );
nand g1231 ( new_n1433_, new_n1432_, new_n1431_ );
nand g1232 ( new_n1434_, new_n1433_, keyIn_0_120 );
nand g1233 ( N748, new_n1430_, new_n1434_ );
not g1234 ( new_n1436_, keyIn_0_121 );
not g1235 ( new_n1437_, keyIn_0_98 );
nor g1236 ( new_n1438_, new_n1415_, new_n875_ );
nor g1237 ( new_n1439_, new_n1438_, new_n1437_ );
nand g1238 ( new_n1440_, new_n1420_, new_n967_ );
nor g1239 ( new_n1441_, new_n1440_, keyIn_0_98 );
nor g1240 ( new_n1442_, new_n1439_, new_n1441_ );
nor g1241 ( new_n1443_, new_n1442_, N101 );
nand g1242 ( new_n1444_, new_n1440_, keyIn_0_98 );
nand g1243 ( new_n1445_, new_n1438_, new_n1437_ );
nand g1244 ( new_n1446_, new_n1445_, new_n1444_ );
nor g1245 ( new_n1447_, new_n1446_, new_n393_ );
nor g1246 ( new_n1448_, new_n1443_, new_n1447_ );
nand g1247 ( new_n1449_, new_n1448_, new_n1436_ );
nand g1248 ( new_n1450_, new_n1446_, new_n393_ );
nand g1249 ( new_n1451_, new_n1442_, N101 );
nand g1250 ( new_n1452_, new_n1451_, new_n1450_ );
nand g1251 ( new_n1453_, new_n1452_, keyIn_0_121 );
nand g1252 ( N749, new_n1449_, new_n1453_ );
not g1253 ( new_n1455_, keyIn_0_122 );
not g1254 ( new_n1456_, keyIn_0_99 );
nor g1255 ( new_n1457_, new_n1415_, new_n801_ );
nor g1256 ( new_n1458_, new_n1457_, new_n1456_ );
nand g1257 ( new_n1459_, new_n1420_, new_n1052_ );
nor g1258 ( new_n1460_, new_n1459_, keyIn_0_99 );
nor g1259 ( new_n1461_, new_n1458_, new_n1460_ );
nor g1260 ( new_n1462_, new_n1461_, new_n402_ );
nand g1261 ( new_n1463_, new_n1459_, keyIn_0_99 );
nand g1262 ( new_n1464_, new_n1457_, new_n1456_ );
nand g1263 ( new_n1465_, new_n1464_, new_n1463_ );
nor g1264 ( new_n1466_, new_n1465_, N105 );
nor g1265 ( new_n1467_, new_n1462_, new_n1466_ );
nand g1266 ( new_n1468_, new_n1467_, new_n1455_ );
nand g1267 ( new_n1469_, new_n1465_, N105 );
nand g1268 ( new_n1470_, new_n1461_, new_n402_ );
nand g1269 ( new_n1471_, new_n1470_, new_n1469_ );
nand g1270 ( new_n1472_, new_n1471_, keyIn_0_122 );
nand g1271 ( N750, new_n1468_, new_n1472_ );
not g1272 ( new_n1474_, keyIn_0_100 );
nor g1273 ( new_n1475_, new_n1415_, new_n1049_ );
nor g1274 ( new_n1476_, new_n1475_, new_n1474_ );
nand g1275 ( new_n1477_, new_n1420_, new_n658_ );
nor g1276 ( new_n1478_, new_n1477_, keyIn_0_100 );
nor g1277 ( new_n1479_, new_n1476_, new_n1478_ );
nor g1278 ( new_n1480_, new_n1479_, new_n404_ );
nand g1279 ( new_n1481_, new_n1477_, keyIn_0_100 );
nand g1280 ( new_n1482_, new_n1475_, new_n1474_ );
nand g1281 ( new_n1483_, new_n1482_, new_n1481_ );
nor g1282 ( new_n1484_, new_n1483_, N109 );
nor g1283 ( new_n1485_, new_n1480_, new_n1484_ );
nand g1284 ( new_n1486_, new_n1485_, keyIn_0_123 );
not g1285 ( new_n1487_, keyIn_0_123 );
nand g1286 ( new_n1488_, new_n1483_, N109 );
nand g1287 ( new_n1489_, new_n1479_, new_n404_ );
nand g1288 ( new_n1490_, new_n1489_, new_n1488_ );
nand g1289 ( new_n1491_, new_n1490_, new_n1487_ );
nand g1290 ( N751, new_n1486_, new_n1491_ );
not g1291 ( new_n1493_, keyIn_0_81 );
not g1292 ( new_n1494_, keyIn_0_69 );
nor g1293 ( new_n1495_, new_n312_, new_n1494_ );
not g1294 ( new_n1496_, new_n1495_ );
nor g1295 ( new_n1497_, new_n951_, new_n526_ );
nand g1296 ( new_n1498_, new_n1496_, new_n1497_ );
not g1297 ( new_n1499_, keyIn_0_70 );
nor g1298 ( new_n1500_, new_n537_, new_n1499_ );
not g1299 ( new_n1501_, new_n1500_ );
nor g1300 ( new_n1502_, new_n311_, keyIn_0_69 );
nor g1301 ( new_n1503_, new_n482_, keyIn_0_70 );
nor g1302 ( new_n1504_, new_n1502_, new_n1503_ );
nand g1303 ( new_n1505_, new_n1504_, new_n1501_ );
nor g1304 ( new_n1506_, new_n1498_, new_n1505_ );
nand g1305 ( new_n1507_, new_n1226_, new_n1506_ );
nand g1306 ( new_n1508_, new_n1507_, new_n1493_ );
not g1307 ( new_n1509_, new_n1508_ );
nor g1308 ( new_n1510_, new_n1507_, new_n1493_ );
nor g1309 ( new_n1511_, new_n1509_, new_n1510_ );
nor g1310 ( new_n1512_, new_n1511_, new_n970_ );
nor g1311 ( new_n1513_, new_n1512_, keyIn_0_101 );
not g1312 ( new_n1514_, keyIn_0_101 );
not g1313 ( new_n1515_, new_n1510_ );
nand g1314 ( new_n1516_, new_n1515_, new_n1508_ );
nand g1315 ( new_n1517_, new_n1516_, new_n932_ );
nor g1316 ( new_n1518_, new_n1517_, new_n1514_ );
nor g1317 ( new_n1519_, new_n1513_, new_n1518_ );
nor g1318 ( new_n1520_, new_n1519_, N113 );
nand g1319 ( new_n1521_, new_n1517_, new_n1514_ );
nand g1320 ( new_n1522_, new_n1512_, keyIn_0_101 );
nand g1321 ( new_n1523_, new_n1522_, new_n1521_ );
nor g1322 ( new_n1524_, new_n1523_, new_n315_ );
nor g1323 ( new_n1525_, new_n1520_, new_n1524_ );
nand g1324 ( new_n1526_, new_n1525_, keyIn_0_124 );
not g1325 ( new_n1527_, keyIn_0_124 );
nand g1326 ( new_n1528_, new_n1523_, new_n315_ );
nand g1327 ( new_n1529_, new_n1519_, N113 );
nand g1328 ( new_n1530_, new_n1529_, new_n1528_ );
nand g1329 ( new_n1531_, new_n1530_, new_n1527_ );
nand g1330 ( N752, new_n1526_, new_n1531_ );
nor g1331 ( new_n1533_, new_n1511_, new_n875_ );
nor g1332 ( new_n1534_, new_n1533_, keyIn_0_102 );
not g1333 ( new_n1535_, keyIn_0_102 );
nand g1334 ( new_n1536_, new_n1516_, new_n967_ );
nor g1335 ( new_n1537_, new_n1536_, new_n1535_ );
nor g1336 ( new_n1538_, new_n1534_, new_n1537_ );
nor g1337 ( new_n1539_, new_n1538_, new_n317_ );
nand g1338 ( new_n1540_, new_n1536_, new_n1535_ );
nand g1339 ( new_n1541_, new_n1533_, keyIn_0_102 );
nand g1340 ( new_n1542_, new_n1541_, new_n1540_ );
nor g1341 ( new_n1543_, new_n1542_, N117 );
nor g1342 ( new_n1544_, new_n1539_, new_n1543_ );
nand g1343 ( new_n1545_, new_n1544_, keyIn_0_125 );
not g1344 ( new_n1546_, keyIn_0_125 );
nand g1345 ( new_n1547_, new_n1542_, N117 );
nand g1346 ( new_n1548_, new_n1538_, new_n317_ );
nand g1347 ( new_n1549_, new_n1548_, new_n1547_ );
nand g1348 ( new_n1550_, new_n1549_, new_n1546_ );
nand g1349 ( N753, new_n1545_, new_n1550_ );
not g1350 ( new_n1552_, keyIn_0_126 );
nor g1351 ( new_n1553_, new_n1511_, new_n801_ );
nor g1352 ( new_n1554_, new_n1553_, keyIn_0_103 );
not g1353 ( new_n1555_, keyIn_0_103 );
nand g1354 ( new_n1556_, new_n1516_, new_n1052_ );
nor g1355 ( new_n1557_, new_n1556_, new_n1555_ );
nor g1356 ( new_n1558_, new_n1554_, new_n1557_ );
nor g1357 ( new_n1559_, new_n1558_, N121 );
nand g1358 ( new_n1560_, new_n1556_, new_n1555_ );
nand g1359 ( new_n1561_, new_n1553_, keyIn_0_103 );
nand g1360 ( new_n1562_, new_n1561_, new_n1560_ );
nor g1361 ( new_n1563_, new_n1562_, new_n326_ );
nor g1362 ( new_n1564_, new_n1559_, new_n1563_ );
nand g1363 ( new_n1565_, new_n1564_, new_n1552_ );
nand g1364 ( new_n1566_, new_n1562_, new_n326_ );
nand g1365 ( new_n1567_, new_n1558_, N121 );
nand g1366 ( new_n1568_, new_n1567_, new_n1566_ );
nand g1367 ( new_n1569_, new_n1568_, keyIn_0_126 );
nand g1368 ( N754, new_n1565_, new_n1569_ );
nor g1369 ( new_n1571_, new_n1511_, new_n1049_ );
nor g1370 ( new_n1572_, new_n1571_, keyIn_0_104 );
not g1371 ( new_n1573_, keyIn_0_104 );
nand g1372 ( new_n1574_, new_n1516_, new_n658_ );
nor g1373 ( new_n1575_, new_n1574_, new_n1573_ );
nor g1374 ( new_n1576_, new_n1572_, new_n1575_ );
nor g1375 ( new_n1577_, new_n1576_, new_n328_ );
nand g1376 ( new_n1578_, new_n1574_, new_n1573_ );
nand g1377 ( new_n1579_, new_n1571_, keyIn_0_104 );
nand g1378 ( new_n1580_, new_n1579_, new_n1578_ );
nor g1379 ( new_n1581_, new_n1580_, N125 );
nor g1380 ( new_n1582_, new_n1577_, new_n1581_ );
nand g1381 ( new_n1583_, new_n1582_, keyIn_0_127 );
not g1382 ( new_n1584_, keyIn_0_127 );
nand g1383 ( new_n1585_, new_n1580_, N125 );
nand g1384 ( new_n1586_, new_n1576_, new_n328_ );
nand g1385 ( new_n1587_, new_n1586_, new_n1585_ );
nand g1386 ( new_n1588_, new_n1587_, new_n1584_ );
nand g1387 ( N755, new_n1583_, new_n1588_ );
endmodule