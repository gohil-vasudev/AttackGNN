module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n976_, new_n1009_, new_n479_, new_n1105_, new_n955_, new_n608_, new_n888_, new_n847_, new_n501_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n390_, new_n743_, new_n779_, new_n1025_, new_n566_, new_n641_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n1125_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n660_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n481_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n635_, new_n685_, new_n1050_, new_n554_, new_n648_, new_n903_, new_n983_, new_n1151_, new_n844_, new_n430_, new_n822_, new_n482_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n1083_, new_n655_, new_n759_, new_n1054_, new_n630_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n565_, new_n361_, new_n764_, new_n906_, new_n683_, new_n511_, new_n510_, new_n966_, new_n351_, new_n517_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n883_, new_n1005_, new_n999_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n568_, new_n420_, new_n1051_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n429_, new_n355_, new_n926_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n1007_, new_n935_, new_n882_, new_n1145_, new_n657_, new_n1150_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1020_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n1041_, new_n917_, new_n426_, new_n1036_, new_n1133_, new_n398_, new_n646_, new_n1132_, new_n395_, new_n538_, new_n1026_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n1106_, new_n473_, new_n1147_, new_n790_, new_n1081_, new_n587_, new_n465_, new_n739_, new_n969_, new_n835_, new_n996_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n705_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n347_, new_n659_, new_n700_, new_n921_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n469_, new_n391_, new_n1154_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n1128_, new_n1002_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n661_, new_n1124_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n494_, new_n672_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n1104_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n460_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n1095_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n897_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n963_, new_n586_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n717_, new_n403_, new_n475_, new_n868_, new_n825_, new_n858_, new_n557_, new_n936_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n407_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n382_, new_n583_, new_n617_, new_n1080_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n755_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n450_, new_n345_, new_n499_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n692_, new_n502_, new_n613_, new_n623_, new_n446_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n585_, new_n751_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n503_, new_n772_, new_n852_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n732_, new_n687_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1052_, new_n638_, new_n523_, new_n909_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n1096_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n1008_, new_n640_, new_n684_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n377_, new_n539_, new_n905_, new_n803_, new_n727_, new_n375_, new_n962_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n780_, new_n984_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n610_, new_n843_, new_n545_, new_n611_, new_n703_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n866_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n686_, new_n934_, new_n551_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n889_, new_n536_, new_n464_, new_n1089_, new_n573_, new_n765_, new_n405_, new_n1103_;

nand g000 ( new_n343_, N29, N42, N75 );
xnor g001 ( N388, new_n343_, keyIn_0_5 );
nand g002 ( new_n345_, N29, N36, N80 );
xnor g003 ( N389, new_n345_, keyIn_0_6 );
nand g004 ( new_n347_, N29, N36, N42 );
not g005 ( N390, new_n347_ );
nand g006 ( new_n349_, N85, N86 );
xnor g007 ( N391, new_n349_, keyIn_0_11 );
nand g008 ( new_n351_, N1, N8, N13, N17 );
xor g009 ( new_n352_, new_n351_, keyIn_0_0 );
xnor g010 ( N418, new_n352_, keyIn_0_40 );
nand g011 ( new_n354_, N1, N13, N17, N26 );
xor g012 ( new_n355_, new_n354_, keyIn_0_1 );
xor g013 ( new_n356_, new_n347_, keyIn_0_2 );
nand g014 ( N419, new_n355_, new_n356_ );
nand g015 ( new_n358_, N59, N75, N80 );
xnor g016 ( new_n359_, new_n358_, keyIn_0_7 );
xnor g017 ( N420, new_n359_, keyIn_0_46 );
nand g018 ( new_n361_, N36, N59, N80 );
xor g019 ( new_n362_, new_n361_, keyIn_0_9 );
xnor g020 ( N421, new_n362_, keyIn_0_47 );
nand g021 ( new_n364_, N36, N42, N59 );
xor g022 ( new_n365_, new_n364_, keyIn_0_10 );
xnor g023 ( N422, new_n365_, keyIn_0_48 );
nor g024 ( new_n367_, N87, N88 );
xor g025 ( new_n368_, new_n367_, keyIn_0_12 );
nand g026 ( new_n369_, new_n368_, N90 );
xnor g027 ( N423, new_n369_, keyIn_0_50 );
xnor g028 ( new_n371_, new_n356_, keyIn_0_41 );
nand g029 ( new_n372_, new_n371_, new_n355_ );
xor g030 ( N446, new_n372_, keyIn_0_58 );
nand g031 ( new_n374_, N1, N26, N51 );
xnor g032 ( new_n375_, new_n374_, keyIn_0_43 );
xnor g033 ( N447, new_n375_, keyIn_0_60 );
nand g034 ( new_n377_, N1, N8, N13, N55 );
not g035 ( new_n378_, new_n377_ );
nand g036 ( new_n379_, new_n378_, N29, N68 );
xnor g037 ( N448, new_n379_, keyIn_0_62 );
nand g038 ( new_n381_, new_n378_, N59, N68, N74 );
xnor g039 ( new_n382_, new_n381_, keyIn_0_45 );
xnor g040 ( N449, new_n382_, keyIn_0_63 );
nand g041 ( new_n384_, new_n368_, N89 );
xor g042 ( N450, new_n384_, keyIn_0_49 );
not g043 ( new_n386_, N121 );
not g044 ( new_n387_, N126 );
nand g045 ( new_n388_, new_n386_, new_n387_ );
nand g046 ( new_n389_, new_n388_, keyIn_0_18 );
nand g047 ( new_n390_, N121, N126 );
not g048 ( new_n391_, keyIn_0_18 );
nand g049 ( new_n392_, new_n391_, new_n386_, new_n387_ );
nand g050 ( new_n393_, new_n389_, new_n390_, new_n392_ );
xnor g051 ( new_n394_, new_n393_, keyIn_0_53 );
xor g052 ( new_n395_, new_n394_, keyIn_0_68 );
nor g053 ( new_n396_, N111, N116 );
xor g054 ( new_n397_, new_n396_, keyIn_0_17 );
nand g055 ( new_n398_, N111, N116 );
xor g056 ( new_n399_, new_n398_, keyIn_0_16 );
nand g057 ( new_n400_, new_n397_, new_n399_ );
xnor g058 ( new_n401_, new_n400_, keyIn_0_52 );
xor g059 ( new_n402_, new_n401_, keyIn_0_67 );
nand g060 ( new_n403_, new_n402_, new_n395_ );
nand g061 ( new_n404_, new_n403_, keyIn_0_78 );
nand g062 ( new_n405_, new_n401_, new_n394_ );
xnor g063 ( new_n406_, new_n405_, keyIn_0_69 );
not g064 ( new_n407_, keyIn_0_78 );
nand g065 ( new_n408_, new_n402_, new_n407_, new_n395_ );
nand g066 ( new_n409_, new_n404_, new_n406_, new_n408_ );
xnor g067 ( new_n410_, new_n409_, keyIn_0_87 );
nand g068 ( new_n411_, new_n410_, N135 );
xor g069 ( new_n412_, new_n411_, keyIn_0_104 );
not g070 ( new_n413_, N135 );
not g071 ( new_n414_, new_n410_ );
nand g072 ( new_n415_, new_n414_, new_n413_ );
xnor g073 ( new_n416_, new_n415_, keyIn_0_105 );
nand g074 ( new_n417_, new_n416_, new_n412_ );
xnor g075 ( new_n418_, new_n417_, keyIn_0_123 );
xnor g076 ( new_n419_, new_n418_, keyIn_0_129 );
nor g077 ( new_n420_, N91, N96 );
xnor g078 ( new_n421_, new_n420_, keyIn_0_14 );
nand g079 ( new_n422_, N91, N96 );
xnor g080 ( new_n423_, new_n422_, keyIn_0_13 );
nand g081 ( new_n424_, new_n421_, new_n423_ );
xnor g082 ( new_n425_, new_n424_, keyIn_0_51 );
not g083 ( new_n426_, new_n425_ );
nand g084 ( new_n427_, new_n426_, keyIn_0_64 );
not g085 ( new_n428_, N101 );
not g086 ( new_n429_, N106 );
nand g087 ( new_n430_, new_n428_, new_n429_ );
nand g088 ( new_n431_, new_n430_, keyIn_0_15 );
nand g089 ( new_n432_, N101, N106 );
not g090 ( new_n433_, keyIn_0_15 );
nand g091 ( new_n434_, new_n433_, new_n428_, new_n429_ );
nand g092 ( new_n435_, new_n431_, new_n432_, new_n434_ );
xnor g093 ( new_n436_, new_n435_, keyIn_0_65 );
not g094 ( new_n437_, new_n436_ );
not g095 ( new_n438_, keyIn_0_64 );
nand g096 ( new_n439_, new_n425_, new_n438_ );
nand g097 ( new_n440_, new_n427_, new_n439_, new_n437_ );
nand g098 ( new_n441_, new_n440_, keyIn_0_77 );
nand g099 ( new_n442_, new_n426_, new_n435_ );
xor g100 ( new_n443_, new_n442_, keyIn_0_66 );
not g101 ( new_n444_, keyIn_0_77 );
nand g102 ( new_n445_, new_n427_, new_n444_, new_n437_, new_n439_ );
nand g103 ( new_n446_, new_n443_, new_n441_, new_n445_ );
xor g104 ( new_n447_, new_n446_, keyIn_0_86 );
nand g105 ( new_n448_, new_n447_, N130 );
xor g106 ( new_n449_, new_n448_, keyIn_0_102 );
not g107 ( new_n450_, N130 );
not g108 ( new_n451_, new_n447_ );
nand g109 ( new_n452_, new_n451_, new_n450_ );
xnor g110 ( new_n453_, new_n452_, keyIn_0_103 );
nand g111 ( new_n454_, new_n453_, new_n449_ );
xnor g112 ( new_n455_, new_n454_, keyIn_0_122 );
xnor g113 ( new_n456_, new_n455_, keyIn_0_128 );
nand g114 ( new_n457_, new_n419_, keyIn_0_138, new_n456_ );
nand g115 ( new_n458_, new_n418_, new_n455_ );
not g116 ( new_n459_, keyIn_0_138 );
nand g117 ( new_n460_, new_n419_, new_n456_ );
nand g118 ( new_n461_, new_n460_, new_n459_ );
nand g119 ( new_n462_, new_n461_, new_n457_, new_n458_ );
xor g120 ( N767, new_n462_, keyIn_0_156 );
not g121 ( new_n464_, keyIn_0_136 );
not g122 ( new_n465_, N171 );
not g123 ( new_n466_, N177 );
nand g124 ( new_n467_, new_n465_, new_n466_ );
xnor g125 ( new_n468_, new_n467_, keyIn_0_28 );
nand g126 ( new_n469_, N171, N177 );
xor g127 ( new_n470_, new_n469_, keyIn_0_27 );
nand g128 ( new_n471_, new_n468_, new_n470_ );
xor g129 ( new_n472_, new_n471_, keyIn_0_72 );
nor g130 ( new_n473_, N159, N165 );
xnor g131 ( new_n474_, new_n473_, keyIn_0_26 );
nand g132 ( new_n475_, N159, N165 );
xnor g133 ( new_n476_, new_n475_, keyIn_0_25 );
nand g134 ( new_n477_, new_n474_, new_n476_ );
xor g135 ( new_n478_, new_n477_, keyIn_0_71 );
nand g136 ( new_n479_, new_n472_, new_n478_ );
xor g137 ( new_n480_, new_n479_, keyIn_0_84 );
nand g138 ( new_n481_, new_n471_, new_n477_ );
nand g139 ( new_n482_, new_n480_, new_n481_ );
xor g140 ( new_n483_, new_n482_, keyIn_0_101 );
nand g141 ( new_n484_, new_n483_, new_n450_ );
xor g142 ( new_n485_, new_n484_, keyIn_0_115 );
not g143 ( new_n486_, new_n483_ );
nand g144 ( new_n487_, new_n486_, N130 );
xnor g145 ( new_n488_, new_n487_, keyIn_0_114 );
nand g146 ( new_n489_, new_n488_, new_n485_, new_n464_ );
nand g147 ( new_n490_, new_n488_, new_n485_ );
nand g148 ( new_n491_, new_n490_, keyIn_0_136 );
not g149 ( new_n492_, keyIn_0_73 );
nor g150 ( new_n493_, N195, N201 );
xnor g151 ( new_n494_, new_n493_, keyIn_0_31 );
nand g152 ( new_n495_, N195, N201 );
xnor g153 ( new_n496_, new_n495_, keyIn_0_30 );
nand g154 ( new_n497_, new_n494_, new_n496_ );
xor g155 ( new_n498_, new_n497_, keyIn_0_57 );
not g156 ( new_n499_, new_n498_ );
nand g157 ( new_n500_, new_n499_, new_n492_ );
not g158 ( new_n501_, N183 );
not g159 ( new_n502_, N189 );
nand g160 ( new_n503_, new_n501_, new_n502_ );
nand g161 ( new_n504_, new_n503_, keyIn_0_29 );
nand g162 ( new_n505_, N183, N189 );
not g163 ( new_n506_, keyIn_0_29 );
nand g164 ( new_n507_, new_n506_, new_n501_, new_n502_ );
nand g165 ( new_n508_, new_n504_, new_n505_, new_n507_ );
xor g166 ( new_n509_, new_n508_, keyIn_0_56 );
not g167 ( new_n510_, new_n509_ );
nand g168 ( new_n511_, new_n498_, keyIn_0_73 );
nand g169 ( new_n512_, new_n500_, new_n511_, new_n510_ );
xor g170 ( new_n513_, new_n512_, keyIn_0_85 );
nand g171 ( new_n514_, new_n499_, new_n509_ );
xnor g172 ( new_n515_, new_n514_, keyIn_0_74 );
nand g173 ( new_n516_, new_n513_, N207, new_n515_ );
xor g174 ( new_n517_, new_n516_, keyIn_0_116 );
not g175 ( new_n518_, N207 );
nand g176 ( new_n519_, new_n513_, new_n515_ );
nand g177 ( new_n520_, new_n519_, new_n518_ );
nand g178 ( new_n521_, new_n491_, new_n489_, new_n517_, new_n520_ );
xor g179 ( new_n522_, new_n521_, keyIn_0_139 );
nand g180 ( new_n523_, new_n517_, new_n520_ );
nand g181 ( new_n524_, new_n490_, new_n523_ );
xnor g182 ( new_n525_, new_n524_, keyIn_0_137 );
nand g183 ( new_n526_, new_n522_, new_n525_ );
xor g184 ( N768, new_n526_, keyIn_0_157 );
not g185 ( new_n528_, keyIn_0_209 );
not g186 ( new_n529_, keyIn_0_192 );
not g187 ( new_n530_, keyIn_0_82 );
not g188 ( new_n531_, keyIn_0_59 );
nand g189 ( new_n532_, keyIn_0_42, N1, N26, N51 );
not g190 ( new_n533_, keyIn_0_42 );
nand g191 ( new_n534_, new_n374_, new_n533_ );
nand g192 ( new_n535_, new_n534_, new_n532_ );
nand g193 ( new_n536_, new_n535_, new_n531_ );
nand g194 ( new_n537_, new_n534_, keyIn_0_59, new_n532_ );
nand g195 ( new_n538_, new_n536_, new_n537_ );
not g196 ( new_n539_, keyIn_0_24 );
nand g197 ( new_n540_, N17, N42 );
nand g198 ( new_n541_, new_n540_, new_n539_ );
nand g199 ( new_n542_, keyIn_0_24, N17, N42 );
nand g200 ( new_n543_, new_n541_, new_n542_ );
not g201 ( new_n544_, keyIn_0_23 );
not g202 ( new_n545_, N17 );
not g203 ( new_n546_, N42 );
nand g204 ( new_n547_, new_n545_, new_n546_ );
nand g205 ( new_n548_, new_n547_, new_n544_ );
nand g206 ( new_n549_, new_n545_, new_n546_, keyIn_0_23 );
nand g207 ( new_n550_, new_n543_, new_n548_, new_n549_ );
nand g208 ( new_n551_, new_n550_, keyIn_0_55 );
nand g209 ( new_n552_, N59, N156 );
not g210 ( new_n553_, new_n552_ );
not g211 ( new_n554_, keyIn_0_55 );
nand g212 ( new_n555_, new_n543_, new_n548_, new_n554_, new_n549_ );
nand g213 ( new_n556_, new_n538_, new_n551_, new_n553_, new_n555_ );
nand g214 ( new_n557_, new_n556_, new_n530_ );
nand g215 ( new_n558_, new_n555_, new_n553_ );
not g216 ( new_n559_, new_n558_ );
nand g217 ( new_n560_, new_n559_, keyIn_0_82, new_n538_, new_n551_ );
nand g218 ( new_n561_, new_n557_, new_n560_ );
nand g219 ( new_n562_, N1, N8, N17, N51 );
xnor g220 ( new_n563_, new_n562_, keyIn_0_3 );
nand g221 ( new_n564_, N42, N59, N75 );
xnor g222 ( new_n565_, new_n564_, keyIn_0_8 );
nand g223 ( new_n566_, new_n563_, new_n565_ );
xor g224 ( new_n567_, new_n566_, keyIn_0_70 );
nand g225 ( new_n568_, new_n561_, new_n567_ );
nand g226 ( new_n569_, new_n568_, keyIn_0_88 );
not g227 ( new_n570_, keyIn_0_88 );
nand g228 ( new_n571_, new_n561_, new_n570_, new_n567_ );
nand g229 ( new_n572_, new_n569_, new_n571_ );
nand g230 ( new_n573_, new_n572_, N126 );
not g231 ( new_n574_, keyIn_0_97 );
not g232 ( new_n575_, keyIn_0_22 );
nand g233 ( new_n576_, new_n552_, new_n575_ );
nand g234 ( new_n577_, keyIn_0_22, N59, N156 );
nand g235 ( new_n578_, new_n576_, new_n577_ );
nand g236 ( new_n579_, new_n578_, N17 );
not g237 ( new_n580_, new_n579_ );
nand g238 ( new_n581_, new_n538_, keyIn_0_83, new_n580_ );
not g239 ( new_n582_, keyIn_0_83 );
nand g240 ( new_n583_, new_n538_, new_n580_ );
nand g241 ( new_n584_, new_n583_, new_n582_ );
nand g242 ( new_n585_, new_n584_, N1, new_n581_ );
nand g243 ( new_n586_, new_n585_, new_n574_ );
nand g244 ( new_n587_, new_n584_, keyIn_0_97, N1, new_n581_ );
nand g245 ( new_n588_, new_n586_, new_n587_ );
nand g246 ( new_n589_, new_n588_, N153 );
nand g247 ( new_n590_, new_n573_, keyIn_0_127, new_n589_ );
nand g248 ( new_n591_, new_n538_, N29, N75, N80 );
not g249 ( new_n592_, new_n591_ );
nand g250 ( new_n593_, new_n592_, keyIn_0_81, N55 );
xnor g251 ( new_n594_, keyIn_0_19, N268 );
xor g252 ( new_n595_, new_n594_, keyIn_0_54 );
not g253 ( new_n596_, new_n595_ );
not g254 ( new_n597_, keyIn_0_81 );
nand g255 ( new_n598_, new_n592_, N55 );
nand g256 ( new_n599_, new_n598_, new_n597_ );
nand g257 ( new_n600_, new_n599_, new_n593_, new_n596_ );
not g258 ( new_n601_, keyIn_0_127 );
nand g259 ( new_n602_, new_n573_, new_n589_ );
nand g260 ( new_n603_, new_n602_, new_n601_ );
nand g261 ( new_n604_, new_n603_, new_n590_, new_n600_ );
nand g262 ( new_n605_, new_n604_, keyIn_0_135 );
not g263 ( new_n606_, keyIn_0_135 );
nand g264 ( new_n607_, new_n603_, new_n606_, new_n590_, new_n600_ );
nand g265 ( new_n608_, new_n605_, N201, new_n607_ );
not g266 ( new_n609_, keyIn_0_154 );
not g267 ( new_n610_, N201 );
nand g268 ( new_n611_, new_n605_, new_n607_ );
nand g269 ( new_n612_, new_n611_, new_n610_ );
nand g270 ( new_n613_, new_n612_, new_n609_ );
nand g271 ( new_n614_, new_n611_, keyIn_0_154, new_n610_ );
nand g272 ( new_n615_, new_n613_, new_n614_ );
nand g273 ( new_n616_, new_n615_, new_n608_ );
not g274 ( new_n617_, new_n616_ );
nand g275 ( new_n618_, new_n617_, new_n529_, N261 );
not g276 ( new_n619_, N261 );
nand g277 ( new_n620_, new_n616_, new_n619_ );
nand g278 ( new_n621_, new_n617_, N261 );
nand g279 ( new_n622_, new_n621_, keyIn_0_192 );
nand g280 ( new_n623_, new_n622_, new_n528_, new_n618_, new_n620_ );
nand g281 ( new_n624_, new_n622_, new_n618_, new_n620_ );
nand g282 ( new_n625_, new_n624_, keyIn_0_209 );
nand g283 ( new_n626_, new_n625_, N219, new_n623_ );
nand g284 ( new_n627_, new_n626_, keyIn_0_215 );
not g285 ( new_n628_, keyIn_0_215 );
nand g286 ( new_n629_, new_n625_, new_n628_, N219, new_n623_ );
not g287 ( new_n630_, keyIn_0_193 );
nand g288 ( new_n631_, new_n617_, new_n630_, N228 );
xnor g289 ( new_n632_, new_n608_, keyIn_0_172 );
nand g290 ( new_n633_, new_n632_, N237 );
xnor g291 ( new_n634_, new_n633_, keyIn_0_194 );
nand g292 ( new_n635_, new_n617_, N228 );
nand g293 ( new_n636_, new_n635_, keyIn_0_193 );
nand g294 ( new_n637_, new_n636_, new_n631_, new_n634_ );
xnor g295 ( new_n638_, new_n637_, keyIn_0_210 );
not g296 ( new_n639_, keyIn_0_173 );
not g297 ( new_n640_, keyIn_0_155 );
not g298 ( new_n641_, new_n611_ );
nand g299 ( new_n642_, new_n641_, N246 );
nand g300 ( new_n643_, new_n642_, new_n640_ );
nand g301 ( new_n644_, N255, N267 );
xnor g302 ( new_n645_, new_n644_, keyIn_0_39 );
not g303 ( new_n646_, new_n645_ );
nand g304 ( new_n647_, new_n641_, keyIn_0_155, N246 );
nand g305 ( new_n648_, new_n643_, new_n639_, new_n646_, new_n647_ );
nand g306 ( new_n649_, new_n643_, new_n646_, new_n647_ );
nand g307 ( new_n650_, new_n649_, keyIn_0_173 );
nand g308 ( new_n651_, N42, N59, N68, N72 );
xnor g309 ( new_n652_, new_n651_, keyIn_0_4 );
nand g310 ( new_n653_, new_n652_, new_n378_ );
xnor g311 ( new_n654_, new_n653_, keyIn_0_44 );
nand g312 ( new_n655_, new_n654_, N73 );
xnor g313 ( new_n656_, new_n655_, keyIn_0_61 );
xor g314 ( new_n657_, new_n656_, keyIn_0_76 );
nand g315 ( new_n658_, new_n657_, N201 );
nand g316 ( new_n659_, N121, N210 );
xor g317 ( new_n660_, new_n659_, keyIn_0_38 );
nand g318 ( new_n661_, new_n650_, new_n648_, new_n658_, new_n660_ );
not g319 ( new_n662_, new_n661_ );
nand g320 ( new_n663_, new_n627_, new_n629_, new_n638_, new_n662_ );
xnor g321 ( new_n664_, new_n663_, keyIn_0_223 );
xnor g322 ( new_n665_, new_n664_, keyIn_0_229 );
xnor g323 ( N850, new_n665_, keyIn_0_234 );
not g324 ( new_n667_, keyIn_0_238 );
not g325 ( new_n668_, keyIn_0_233 );
not g326 ( new_n669_, keyIn_0_226 );
not g327 ( new_n670_, keyIn_0_216 );
not g328 ( new_n671_, keyIn_0_211 );
not g329 ( new_n672_, keyIn_0_165 );
not g330 ( new_n673_, keyIn_0_149 );
nand g331 ( new_n674_, new_n572_, keyIn_0_111, N111 );
nand g332 ( new_n675_, new_n588_, N143 );
not g333 ( new_n676_, keyIn_0_111 );
nand g334 ( new_n677_, new_n572_, N111 );
nand g335 ( new_n678_, new_n677_, new_n676_ );
nand g336 ( new_n679_, new_n678_, new_n674_, new_n675_ );
xnor g337 ( new_n680_, new_n679_, keyIn_0_126 );
xor g338 ( new_n681_, new_n600_, keyIn_0_98 );
nand g339 ( new_n682_, new_n680_, new_n681_ );
xnor g340 ( new_n683_, new_n682_, keyIn_0_132 );
not g341 ( new_n684_, new_n683_ );
nand g342 ( new_n685_, new_n684_, N183 );
xnor g343 ( new_n686_, new_n685_, new_n673_ );
nand g344 ( new_n687_, new_n683_, new_n501_ );
xnor g345 ( new_n688_, new_n687_, keyIn_0_150 );
nand g346 ( new_n689_, new_n686_, new_n688_ );
xnor g347 ( new_n690_, new_n689_, new_n672_ );
not g348 ( new_n691_, keyIn_0_204 );
not g349 ( new_n692_, keyIn_0_176 );
nand g350 ( new_n693_, new_n572_, N116 );
nand g351 ( new_n694_, new_n588_, N146 );
xor g352 ( new_n695_, new_n600_, keyIn_0_99 );
nand g353 ( new_n696_, new_n695_, new_n693_, new_n694_ );
xnor g354 ( new_n697_, new_n696_, keyIn_0_133 );
nand g355 ( new_n698_, new_n697_, new_n502_ );
not g356 ( new_n699_, N195 );
not g357 ( new_n700_, keyIn_0_134 );
xnor g358 ( new_n701_, new_n600_, keyIn_0_100 );
nand g359 ( new_n702_, new_n572_, N121 );
nand g360 ( new_n703_, new_n702_, keyIn_0_113 );
nand g361 ( new_n704_, new_n588_, N149 );
nand g362 ( new_n705_, new_n704_, keyIn_0_112 );
not g363 ( new_n706_, keyIn_0_112 );
nand g364 ( new_n707_, new_n588_, new_n706_, N149 );
nand g365 ( new_n708_, new_n705_, new_n707_ );
not g366 ( new_n709_, keyIn_0_113 );
nand g367 ( new_n710_, new_n572_, new_n709_, N121 );
nand g368 ( new_n711_, new_n703_, new_n701_, new_n708_, new_n710_ );
nand g369 ( new_n712_, new_n711_, new_n700_ );
nand g370 ( new_n713_, new_n708_, new_n710_ );
not g371 ( new_n714_, new_n713_ );
nand g372 ( new_n715_, new_n714_, keyIn_0_134, new_n701_, new_n703_ );
nand g373 ( new_n716_, new_n715_, new_n712_ );
nand g374 ( new_n717_, new_n716_, new_n699_ );
nand g375 ( new_n718_, new_n717_, keyIn_0_152 );
not g376 ( new_n719_, keyIn_0_152 );
nand g377 ( new_n720_, new_n716_, new_n719_, new_n699_ );
nand g378 ( new_n721_, new_n718_, new_n720_ );
nand g379 ( new_n722_, new_n615_, N261, new_n721_, new_n698_ );
xnor g380 ( new_n723_, new_n722_, new_n692_ );
not g381 ( new_n724_, keyIn_0_197 );
nand g382 ( new_n725_, new_n632_, new_n721_, new_n698_ );
xnor g383 ( new_n726_, new_n725_, new_n724_ );
not g384 ( new_n727_, keyIn_0_169 );
nand g385 ( new_n728_, new_n715_, N195, new_n712_ );
nand g386 ( new_n729_, new_n728_, new_n727_ );
nand g387 ( new_n730_, new_n715_, keyIn_0_169, N195, new_n712_ );
nand g388 ( new_n731_, new_n729_, new_n730_ );
nand g389 ( new_n732_, new_n731_, new_n698_ );
nand g390 ( new_n733_, new_n732_, keyIn_0_196 );
not g391 ( new_n734_, keyIn_0_196 );
nand g392 ( new_n735_, new_n731_, new_n734_, new_n698_ );
nand g393 ( new_n736_, new_n733_, new_n735_ );
not g394 ( new_n737_, new_n697_ );
nand g395 ( new_n738_, new_n737_, N189 );
nand g396 ( new_n739_, new_n736_, new_n738_ );
not g397 ( new_n740_, new_n739_ );
nand g398 ( new_n741_, new_n723_, new_n726_, new_n740_ );
nand g399 ( new_n742_, new_n741_, new_n691_ );
nand g400 ( new_n743_, new_n723_, keyIn_0_204, new_n726_, new_n740_ );
nand g401 ( new_n744_, new_n742_, new_n743_ );
not g402 ( new_n745_, new_n744_ );
nand g403 ( new_n746_, new_n690_, new_n745_ );
nand g404 ( new_n747_, new_n746_, new_n671_ );
nand g405 ( new_n748_, new_n690_, new_n745_, keyIn_0_211 );
not g406 ( new_n749_, new_n690_ );
nand g407 ( new_n750_, new_n749_, new_n744_ );
nand g408 ( new_n751_, new_n747_, new_n670_, new_n748_, new_n750_ );
nand g409 ( new_n752_, new_n747_, new_n748_, new_n750_ );
nand g410 ( new_n753_, new_n752_, keyIn_0_216 );
nand g411 ( new_n754_, new_n753_, N219, new_n751_ );
xor g412 ( new_n755_, new_n754_, keyIn_0_220 );
nand g413 ( new_n756_, N106, N210 );
xor g414 ( new_n757_, new_n756_, keyIn_0_34 );
nand g415 ( new_n758_, new_n755_, new_n669_, new_n757_ );
nand g416 ( new_n759_, new_n755_, new_n757_ );
nand g417 ( new_n760_, new_n759_, keyIn_0_226 );
not g418 ( new_n761_, keyIn_0_205 );
nand g419 ( new_n762_, new_n749_, N228 );
not g420 ( new_n763_, new_n686_ );
nand g421 ( new_n764_, new_n763_, N237 );
xnor g422 ( new_n765_, new_n764_, keyIn_0_186 );
nand g423 ( new_n766_, new_n762_, new_n761_, new_n765_ );
nand g424 ( new_n767_, new_n762_, new_n765_ );
nand g425 ( new_n768_, new_n767_, keyIn_0_205 );
nand g426 ( new_n769_, new_n684_, N246 );
nand g427 ( new_n770_, new_n657_, N183 );
xnor g428 ( new_n771_, new_n770_, keyIn_0_121 );
nand g429 ( new_n772_, new_n769_, new_n771_ );
xnor g430 ( new_n773_, new_n772_, keyIn_0_166 );
nand g431 ( new_n774_, new_n768_, new_n766_, new_n773_ );
not g432 ( new_n775_, new_n774_ );
nand g433 ( new_n776_, new_n760_, new_n758_, new_n775_ );
nand g434 ( new_n777_, new_n776_, new_n668_ );
nand g435 ( new_n778_, new_n760_, keyIn_0_233, new_n758_, new_n775_ );
nand g436 ( new_n779_, new_n777_, new_n778_ );
nand g437 ( new_n780_, new_n779_, new_n667_ );
nand g438 ( new_n781_, new_n777_, keyIn_0_238, new_n778_ );
nand g439 ( new_n782_, new_n780_, new_n781_ );
xnor g440 ( N863, new_n782_, keyIn_0_245 );
not g441 ( new_n784_, keyIn_0_221 );
nand g442 ( new_n785_, new_n615_, N261, new_n721_ );
xnor g443 ( new_n786_, new_n785_, keyIn_0_175 );
not g444 ( new_n787_, keyIn_0_195 );
nand g445 ( new_n788_, new_n632_, new_n721_ );
nand g446 ( new_n789_, new_n788_, new_n787_ );
xor g447 ( new_n790_, new_n731_, keyIn_0_189 );
nand g448 ( new_n791_, new_n632_, new_n721_, keyIn_0_195 );
nand g449 ( new_n792_, new_n786_, new_n789_, new_n790_, new_n791_ );
xnor g450 ( new_n793_, new_n792_, keyIn_0_206 );
nand g451 ( new_n794_, new_n738_, new_n698_ );
xor g452 ( new_n795_, new_n794_, keyIn_0_167 );
not g453 ( new_n796_, new_n795_ );
nand g454 ( new_n797_, new_n793_, keyIn_0_212, new_n796_ );
not g455 ( new_n798_, keyIn_0_212 );
nand g456 ( new_n799_, new_n793_, new_n796_ );
nand g457 ( new_n800_, new_n799_, new_n798_ );
not g458 ( new_n801_, new_n793_ );
nand g459 ( new_n802_, new_n801_, new_n795_ );
nand g460 ( new_n803_, new_n802_, N219 );
not g461 ( new_n804_, new_n803_ );
nand g462 ( new_n805_, new_n804_, new_n797_, new_n800_ );
nand g463 ( new_n806_, new_n805_, new_n784_ );
nand g464 ( new_n807_, N111, N210 );
xor g465 ( new_n808_, new_n807_, keyIn_0_35 );
nand g466 ( new_n809_, new_n804_, keyIn_0_221, new_n797_, new_n800_ );
nand g467 ( new_n810_, new_n806_, new_n808_, new_n809_ );
xnor g468 ( new_n811_, new_n810_, keyIn_0_227 );
nand g469 ( new_n812_, new_n796_, N228 );
xnor g470 ( new_n813_, new_n812_, keyIn_0_187 );
nand g471 ( new_n814_, new_n737_, N246 );
xnor g472 ( new_n815_, new_n814_, keyIn_0_151 );
nand g473 ( new_n816_, N255, N259 );
xnor g474 ( new_n817_, new_n816_, keyIn_0_36 );
nand g475 ( new_n818_, new_n815_, keyIn_0_168, new_n817_ );
not g476 ( new_n819_, keyIn_0_168 );
nand g477 ( new_n820_, new_n815_, new_n817_ );
nand g478 ( new_n821_, new_n820_, new_n819_ );
not g479 ( new_n822_, keyIn_0_188 );
nand g480 ( new_n823_, new_n737_, N189, N237 );
nand g481 ( new_n824_, new_n823_, new_n822_ );
nand g482 ( new_n825_, new_n657_, N189 );
not g483 ( new_n826_, new_n825_ );
nor g484 ( new_n827_, new_n823_, new_n822_ );
nor g485 ( new_n828_, new_n827_, new_n826_ );
nand g486 ( new_n829_, new_n821_, new_n818_, new_n824_, new_n828_ );
not g487 ( new_n830_, new_n829_ );
nand g488 ( new_n831_, new_n811_, new_n813_, new_n830_ );
xor g489 ( new_n832_, new_n831_, keyIn_0_239 );
xnor g490 ( N864, new_n832_, keyIn_0_246 );
not g491 ( new_n834_, keyIn_0_228 );
not g492 ( new_n835_, keyIn_0_222 );
not g493 ( new_n836_, keyIn_0_213 );
nand g494 ( new_n837_, new_n721_, new_n728_ );
xor g495 ( new_n838_, new_n837_, keyIn_0_170 );
not g496 ( new_n839_, new_n632_ );
nand g497 ( new_n840_, new_n615_, N261 );
xor g498 ( new_n841_, new_n840_, keyIn_0_174 );
nand g499 ( new_n842_, new_n841_, new_n839_ );
xor g500 ( new_n843_, new_n842_, keyIn_0_207 );
not g501 ( new_n844_, new_n843_ );
nand g502 ( new_n845_, new_n844_, new_n838_ );
xnor g503 ( new_n846_, new_n845_, new_n836_ );
not g504 ( new_n847_, new_n838_ );
nand g505 ( new_n848_, new_n843_, new_n847_ );
xor g506 ( new_n849_, new_n848_, keyIn_0_214 );
nand g507 ( new_n850_, new_n846_, new_n849_, keyIn_0_217 );
not g508 ( new_n851_, keyIn_0_217 );
nand g509 ( new_n852_, new_n846_, new_n849_ );
nand g510 ( new_n853_, new_n852_, new_n851_ );
nand g511 ( new_n854_, new_n853_, N219, new_n850_ );
nand g512 ( new_n855_, new_n854_, new_n835_ );
nand g513 ( new_n856_, N116, N210 );
nand g514 ( new_n857_, new_n853_, keyIn_0_222, N219, new_n850_ );
nand g515 ( new_n858_, new_n855_, new_n856_, new_n857_ );
nand g516 ( new_n859_, new_n858_, new_n834_ );
nand g517 ( new_n860_, new_n855_, keyIn_0_228, new_n856_, new_n857_ );
nand g518 ( new_n861_, new_n847_, N228 );
nand g519 ( new_n862_, new_n861_, keyIn_0_190 );
nand g520 ( new_n863_, new_n731_, N237 );
xor g521 ( new_n864_, new_n863_, keyIn_0_191 );
not g522 ( new_n865_, new_n864_ );
not g523 ( new_n866_, keyIn_0_190 );
nand g524 ( new_n867_, new_n847_, new_n866_, N228 );
nand g525 ( new_n868_, new_n862_, keyIn_0_208, new_n865_, new_n867_ );
not g526 ( new_n869_, keyIn_0_208 );
nand g527 ( new_n870_, new_n862_, new_n865_, new_n867_ );
nand g528 ( new_n871_, new_n870_, new_n869_ );
not g529 ( new_n872_, keyIn_0_171 );
nand g530 ( new_n873_, new_n715_, N246, new_n712_ );
xnor g531 ( new_n874_, new_n873_, keyIn_0_153 );
nand g532 ( new_n875_, N255, N260 );
xor g533 ( new_n876_, new_n875_, keyIn_0_37 );
nand g534 ( new_n877_, new_n874_, new_n872_, new_n876_ );
nand g535 ( new_n878_, new_n657_, N195 );
nand g536 ( new_n879_, new_n874_, new_n876_ );
nand g537 ( new_n880_, new_n879_, keyIn_0_171 );
nand g538 ( new_n881_, new_n880_, new_n877_, new_n878_ );
not g539 ( new_n882_, new_n881_ );
nand g540 ( new_n883_, new_n871_, new_n868_, new_n882_ );
not g541 ( new_n884_, new_n883_ );
nand g542 ( new_n885_, new_n859_, new_n860_, new_n884_ );
xor g543 ( new_n886_, new_n885_, keyIn_0_240 );
xnor g544 ( N865, new_n886_, keyIn_0_247 );
not g545 ( new_n888_, keyIn_0_225 );
not g546 ( new_n889_, keyIn_0_80 );
nand g547 ( new_n890_, new_n592_, new_n889_, N17 );
nand g548 ( new_n891_, new_n592_, N17 );
nand g549 ( new_n892_, new_n891_, keyIn_0_80 );
nand g550 ( new_n893_, new_n892_, new_n594_, new_n890_ );
xor g551 ( new_n894_, new_n893_, keyIn_0_94 );
nand g552 ( new_n895_, new_n538_, N55, new_n578_ );
xor g553 ( new_n896_, new_n895_, keyIn_0_79 );
nand g554 ( new_n897_, new_n896_, N149 );
xnor g555 ( new_n898_, new_n897_, keyIn_0_93 );
nand g556 ( new_n899_, new_n894_, new_n898_ );
xor g557 ( new_n900_, new_n899_, keyIn_0_108 );
nand g558 ( new_n901_, new_n572_, N101 );
nand g559 ( new_n902_, N17, N138 );
xor g560 ( new_n903_, new_n902_, keyIn_0_21 );
nand g561 ( new_n904_, new_n901_, new_n903_ );
xnor g562 ( new_n905_, new_n904_, keyIn_0_124 );
nand g563 ( new_n906_, new_n900_, new_n905_ );
xnor g564 ( new_n907_, new_n906_, keyIn_0_131 );
nand g565 ( new_n908_, new_n907_, new_n465_ );
xnor g566 ( new_n909_, new_n908_, keyIn_0_145 );
not g567 ( new_n910_, N165 );
xor g568 ( new_n911_, new_n893_, keyIn_0_92 );
nand g569 ( new_n912_, new_n896_, N146 );
xnor g570 ( new_n913_, new_n912_, keyIn_0_91 );
nand g571 ( new_n914_, new_n911_, new_n913_ );
xnor g572 ( new_n915_, new_n914_, keyIn_0_107 );
not g573 ( new_n916_, keyIn_0_106 );
nand g574 ( new_n917_, new_n572_, new_n916_, N96 );
nand g575 ( new_n918_, N51, N138 );
xnor g576 ( new_n919_, new_n918_, keyIn_0_20 );
nand g577 ( new_n920_, new_n572_, N96 );
nand g578 ( new_n921_, new_n920_, keyIn_0_106 );
nand g579 ( new_n922_, new_n915_, new_n917_, new_n919_, new_n921_ );
xor g580 ( new_n923_, new_n922_, keyIn_0_130 );
nand g581 ( new_n924_, new_n923_, new_n910_ );
xor g582 ( new_n925_, new_n924_, keyIn_0_144 );
nand g583 ( new_n926_, new_n925_, new_n909_ );
not g584 ( new_n927_, new_n926_ );
nand g585 ( new_n928_, new_n744_, new_n688_ );
xor g586 ( new_n929_, new_n686_, keyIn_0_185 );
nand g587 ( new_n930_, new_n928_, new_n929_ );
nand g588 ( new_n931_, new_n572_, N106 );
nand g589 ( new_n932_, new_n931_, keyIn_0_109 );
nand g590 ( new_n933_, N138, N152 );
not g591 ( new_n934_, keyIn_0_109 );
nand g592 ( new_n935_, new_n572_, new_n934_, N106 );
nand g593 ( new_n936_, new_n932_, keyIn_0_125, new_n933_, new_n935_ );
not g594 ( new_n937_, keyIn_0_125 );
nand g595 ( new_n938_, new_n932_, new_n933_, new_n935_ );
nand g596 ( new_n939_, new_n938_, new_n937_ );
xnor g597 ( new_n940_, new_n893_, keyIn_0_96 );
nand g598 ( new_n941_, new_n896_, N153 );
xnor g599 ( new_n942_, new_n941_, keyIn_0_95 );
nand g600 ( new_n943_, new_n940_, new_n942_ );
xnor g601 ( new_n944_, new_n943_, keyIn_0_110 );
nand g602 ( new_n945_, new_n944_, new_n939_, new_n466_, new_n936_ );
xnor g603 ( new_n946_, new_n945_, keyIn_0_147 );
nand g604 ( new_n947_, new_n930_, new_n888_, new_n927_, new_n946_ );
nand g605 ( new_n948_, new_n930_, new_n927_, new_n946_ );
nand g606 ( new_n949_, new_n948_, keyIn_0_225 );
nand g607 ( new_n950_, new_n944_, new_n939_, new_n936_ );
nand g608 ( new_n951_, new_n950_, N177 );
xnor g609 ( new_n952_, new_n951_, keyIn_0_146 );
xor g610 ( new_n953_, new_n952_, keyIn_0_162 );
not g611 ( new_n954_, new_n953_ );
nand g612 ( new_n955_, new_n927_, new_n954_ );
nand g613 ( new_n956_, new_n955_, keyIn_0_200 );
not g614 ( new_n957_, new_n956_ );
not g615 ( new_n958_, keyIn_0_200 );
nand g616 ( new_n959_, new_n927_, new_n958_, new_n954_ );
not g617 ( new_n960_, new_n923_ );
nand g618 ( new_n961_, new_n960_, N165 );
xnor g619 ( new_n962_, new_n961_, keyIn_0_143 );
xnor g620 ( new_n963_, new_n962_, keyIn_0_179 );
not g621 ( new_n964_, keyIn_0_199 );
not g622 ( new_n965_, new_n907_ );
nand g623 ( new_n966_, new_n965_, N171 );
not g624 ( new_n967_, new_n966_ );
nand g625 ( new_n968_, new_n925_, new_n967_ );
xnor g626 ( new_n969_, new_n968_, new_n964_ );
nand g627 ( new_n970_, new_n969_, new_n959_, new_n963_ );
nor g628 ( new_n971_, new_n970_, new_n957_ );
nand g629 ( new_n972_, new_n949_, new_n947_, new_n971_ );
not g630 ( new_n973_, N159 );
nand g631 ( new_n974_, new_n572_, N91 );
xor g632 ( new_n975_, new_n893_, keyIn_0_90 );
not g633 ( new_n976_, keyIn_0_89 );
nand g634 ( new_n977_, new_n896_, new_n976_, N143 );
nand g635 ( new_n978_, N8, N138 );
nand g636 ( new_n979_, new_n896_, N143 );
nand g637 ( new_n980_, new_n979_, keyIn_0_89 );
nand g638 ( new_n981_, new_n980_, new_n977_, new_n978_ );
nor g639 ( new_n982_, new_n975_, new_n981_ );
nand g640 ( new_n983_, new_n982_, new_n973_, new_n974_ );
xor g641 ( new_n984_, new_n983_, keyIn_0_141 );
nand g642 ( new_n985_, new_n972_, keyIn_0_235, new_n984_ );
nand g643 ( new_n986_, new_n982_, new_n974_ );
nand g644 ( new_n987_, new_n986_, N159 );
xor g645 ( new_n988_, new_n987_, keyIn_0_140 );
xnor g646 ( new_n989_, new_n988_, keyIn_0_177 );
not g647 ( new_n990_, keyIn_0_235 );
nand g648 ( new_n991_, new_n972_, new_n984_ );
nand g649 ( new_n992_, new_n991_, new_n990_ );
nand g650 ( new_n993_, new_n992_, new_n985_, new_n989_ );
xor g651 ( new_n994_, new_n993_, keyIn_0_241 );
xnor g652 ( N866, new_n994_, keyIn_0_248 );
nand g653 ( new_n996_, new_n952_, new_n946_ );
xnor g654 ( new_n997_, new_n996_, keyIn_0_163 );
not g655 ( new_n998_, new_n997_ );
nand g656 ( new_n999_, new_n930_, new_n998_ );
xor g657 ( new_n1000_, new_n999_, keyIn_0_219 );
not g658 ( new_n1001_, new_n930_ );
nand g659 ( new_n1002_, new_n1001_, keyIn_0_218, new_n997_ );
not g660 ( new_n1003_, keyIn_0_218 );
nand g661 ( new_n1004_, new_n1001_, new_n997_ );
nand g662 ( new_n1005_, new_n1004_, new_n1003_ );
nand g663 ( new_n1006_, new_n1000_, new_n1002_, N219, new_n1005_ );
not g664 ( new_n1007_, keyIn_0_184 );
nand g665 ( new_n1008_, new_n998_, N228 );
nand g666 ( new_n1009_, new_n1008_, new_n1007_ );
nand g667 ( new_n1010_, new_n998_, keyIn_0_184, N228 );
nand g668 ( new_n1011_, new_n954_, N237 );
not g669 ( new_n1012_, new_n1011_ );
not g670 ( new_n1013_, keyIn_0_164 );
nand g671 ( new_n1014_, new_n950_, keyIn_0_148, N246 );
nand g672 ( new_n1015_, new_n657_, N177 );
xnor g673 ( new_n1016_, new_n1015_, keyIn_0_120 );
not g674 ( new_n1017_, keyIn_0_148 );
nand g675 ( new_n1018_, new_n950_, N246 );
nand g676 ( new_n1019_, new_n1018_, new_n1017_ );
nand g677 ( new_n1020_, new_n1019_, new_n1014_, new_n1016_ );
nand g678 ( new_n1021_, new_n1020_, new_n1013_ );
nand g679 ( new_n1022_, new_n1019_, keyIn_0_164, new_n1014_, new_n1016_ );
nand g680 ( new_n1023_, N101, N210 );
nand g681 ( new_n1024_, new_n1021_, new_n1022_, new_n1023_ );
nor g682 ( new_n1025_, new_n1012_, new_n1024_ );
nand g683 ( new_n1026_, new_n1006_, new_n1009_, new_n1010_, new_n1025_ );
xnor g684 ( new_n1027_, new_n1026_, keyIn_0_244 );
xnor g685 ( N874, new_n1027_, keyIn_0_253 );
not g686 ( new_n1029_, keyIn_0_251 );
not g687 ( new_n1030_, keyIn_0_249 );
not g688 ( new_n1031_, keyIn_0_236 );
nand g689 ( new_n1032_, new_n988_, new_n984_ );
xnor g690 ( new_n1033_, new_n1032_, keyIn_0_158 );
not g691 ( new_n1034_, new_n1033_ );
nand g692 ( new_n1035_, new_n972_, new_n1034_ );
nand g693 ( new_n1036_, new_n1035_, keyIn_0_230 );
not g694 ( new_n1037_, keyIn_0_230 );
nand g695 ( new_n1038_, new_n972_, new_n1037_, new_n1034_ );
nand g696 ( new_n1039_, new_n1036_, new_n1038_ );
nand g697 ( new_n1040_, new_n949_, new_n971_, new_n947_, new_n1033_ );
nand g698 ( new_n1041_, new_n1039_, new_n1031_, new_n1040_ );
nand g699 ( new_n1042_, new_n1039_, new_n1040_ );
nand g700 ( new_n1043_, new_n1042_, keyIn_0_236 );
nand g701 ( new_n1044_, new_n1043_, N219, new_n1041_ );
nand g702 ( new_n1045_, new_n595_, N210 );
xnor g703 ( new_n1046_, new_n1045_, keyIn_0_75 );
nand g704 ( new_n1047_, new_n1044_, new_n1046_ );
nand g705 ( new_n1048_, new_n1047_, new_n1030_ );
nand g706 ( new_n1049_, new_n1044_, keyIn_0_249, new_n1046_ );
nand g707 ( new_n1050_, new_n1048_, new_n1049_ );
nand g708 ( new_n1051_, new_n1034_, N228 );
xor g709 ( new_n1052_, new_n1051_, keyIn_0_178 );
not g710 ( new_n1053_, new_n988_ );
nand g711 ( new_n1054_, new_n1053_, N237 );
nand g712 ( new_n1055_, new_n1052_, keyIn_0_201, new_n1054_ );
not g713 ( new_n1056_, keyIn_0_201 );
nand g714 ( new_n1057_, new_n1052_, new_n1054_ );
nand g715 ( new_n1058_, new_n1057_, new_n1056_ );
nand g716 ( new_n1059_, new_n986_, keyIn_0_142, N246 );
not g717 ( new_n1060_, keyIn_0_142 );
nand g718 ( new_n1061_, new_n986_, N246 );
nand g719 ( new_n1062_, new_n1061_, new_n1060_ );
nand g720 ( new_n1063_, new_n657_, N159 );
xnor g721 ( new_n1064_, new_n1063_, keyIn_0_117 );
nand g722 ( new_n1065_, new_n1062_, new_n1064_, new_n1059_ );
not g723 ( new_n1066_, new_n1065_ );
nand g724 ( new_n1067_, new_n1058_, new_n1055_, new_n1066_ );
not g725 ( new_n1068_, new_n1067_ );
nand g726 ( new_n1069_, new_n1050_, new_n1068_ );
nand g727 ( new_n1070_, new_n1069_, new_n1029_ );
nand g728 ( new_n1071_, new_n1050_, keyIn_0_251, new_n1068_ );
nand g729 ( new_n1072_, new_n1070_, new_n1071_ );
nand g730 ( new_n1073_, new_n1072_, keyIn_0_254 );
not g731 ( new_n1074_, keyIn_0_254 );
nand g732 ( new_n1075_, new_n1070_, new_n1074_, new_n1071_ );
nand g733 ( N878, new_n1073_, new_n1075_ );
not g734 ( new_n1077_, keyIn_0_255 );
nand g735 ( new_n1078_, new_n930_, new_n946_ );
not g736 ( new_n1079_, new_n1078_ );
nand g737 ( new_n1080_, new_n1079_, keyIn_0_224, new_n909_ );
not g738 ( new_n1081_, keyIn_0_224 );
nand g739 ( new_n1082_, new_n1079_, new_n909_ );
nand g740 ( new_n1083_, new_n1082_, new_n1081_ );
not g741 ( new_n1084_, keyIn_0_198 );
nand g742 ( new_n1085_, new_n954_, new_n1084_, new_n909_ );
nand g743 ( new_n1086_, new_n954_, new_n909_ );
nand g744 ( new_n1087_, new_n1086_, keyIn_0_198 );
xnor g745 ( new_n1088_, new_n966_, keyIn_0_181 );
nand g746 ( new_n1089_, new_n1087_, new_n1085_, new_n1088_ );
not g747 ( new_n1090_, new_n1089_ );
not g748 ( new_n1091_, new_n962_ );
nand g749 ( new_n1092_, new_n1091_, new_n925_ );
xor g750 ( new_n1093_, new_n1092_, keyIn_0_159 );
nand g751 ( new_n1094_, new_n1083_, new_n1080_, new_n1090_, new_n1093_ );
nand g752 ( new_n1095_, new_n1083_, new_n1080_, new_n1090_ );
not g753 ( new_n1096_, new_n1093_ );
nand g754 ( new_n1097_, new_n1095_, new_n1096_ );
nand g755 ( new_n1098_, new_n1097_, N219, new_n1094_ );
xnor g756 ( new_n1099_, new_n1098_, keyIn_0_242 );
nand g757 ( new_n1100_, N91, N210 );
xor g758 ( new_n1101_, new_n1100_, keyIn_0_32 );
nand g759 ( new_n1102_, new_n1099_, new_n1101_ );
xor g760 ( new_n1103_, new_n1102_, keyIn_0_250 );
nand g761 ( new_n1104_, new_n1096_, keyIn_0_180, N228 );
nand g762 ( new_n1105_, new_n962_, N237 );
not g763 ( new_n1106_, keyIn_0_180 );
nand g764 ( new_n1107_, new_n1096_, N228 );
nand g765 ( new_n1108_, new_n1107_, new_n1106_ );
nand g766 ( new_n1109_, new_n1108_, keyIn_0_202, new_n1104_, new_n1105_ );
not g767 ( new_n1110_, keyIn_0_202 );
nand g768 ( new_n1111_, new_n1108_, new_n1104_, new_n1105_ );
nand g769 ( new_n1112_, new_n1111_, new_n1110_ );
nand g770 ( new_n1113_, new_n960_, N246 );
nand g771 ( new_n1114_, new_n657_, N165 );
xnor g772 ( new_n1115_, new_n1114_, keyIn_0_118 );
nand g773 ( new_n1116_, new_n1112_, new_n1109_, new_n1113_, new_n1115_ );
not g774 ( new_n1117_, new_n1116_ );
nand g775 ( new_n1118_, new_n1103_, new_n1117_ );
xnor g776 ( N879, new_n1118_, new_n1077_ );
not g777 ( new_n1120_, keyIn_0_237 );
nand g778 ( new_n1121_, new_n909_, new_n966_ );
xnor g779 ( new_n1122_, new_n1121_, keyIn_0_160 );
xor g780 ( new_n1123_, new_n953_, keyIn_0_183 );
nand g781 ( new_n1124_, new_n1078_, new_n1122_, new_n1123_ );
xnor g782 ( new_n1125_, new_n1124_, keyIn_0_231 );
not g783 ( new_n1126_, new_n1122_ );
nand g784 ( new_n1127_, new_n1078_, new_n1123_ );
nand g785 ( new_n1128_, new_n1127_, new_n1126_ );
xor g786 ( new_n1129_, new_n1128_, keyIn_0_232 );
nand g787 ( new_n1130_, new_n1129_, new_n1125_ );
nand g788 ( new_n1131_, new_n1130_, new_n1120_ );
nand g789 ( new_n1132_, new_n1129_, keyIn_0_237, new_n1125_ );
nand g790 ( new_n1133_, new_n1131_, N219, new_n1132_ );
nand g791 ( new_n1134_, new_n1133_, keyIn_0_243 );
not g792 ( new_n1135_, keyIn_0_243 );
nand g793 ( new_n1136_, new_n1131_, new_n1135_, N219, new_n1132_ );
not g794 ( new_n1137_, keyIn_0_203 );
nand g795 ( new_n1138_, new_n1126_, N228 );
nand g796 ( new_n1139_, new_n967_, N237 );
xnor g797 ( new_n1140_, new_n1139_, keyIn_0_182 );
nand g798 ( new_n1141_, new_n1138_, new_n1140_ );
nand g799 ( new_n1142_, new_n1141_, new_n1137_ );
nand g800 ( new_n1143_, new_n1138_, keyIn_0_203, new_n1140_ );
not g801 ( new_n1144_, keyIn_0_161 );
nand g802 ( new_n1145_, new_n965_, N246 );
nand g803 ( new_n1146_, new_n657_, N171 );
xnor g804 ( new_n1147_, new_n1146_, keyIn_0_119 );
nand g805 ( new_n1148_, new_n1145_, new_n1147_ );
nand g806 ( new_n1149_, new_n1148_, new_n1144_ );
nand g807 ( new_n1150_, new_n1145_, keyIn_0_161, new_n1147_ );
nand g808 ( new_n1151_, N96, N210 );
xor g809 ( new_n1152_, new_n1151_, keyIn_0_33 );
nand g810 ( new_n1153_, new_n1143_, new_n1149_, new_n1150_, new_n1152_ );
not g811 ( new_n1154_, new_n1153_ );
nand g812 ( new_n1155_, new_n1134_, new_n1136_, new_n1142_, new_n1154_ );
xnor g813 ( N880, new_n1155_, keyIn_0_252 );
endmodule