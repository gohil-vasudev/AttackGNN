module add_mul_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, 
        b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, 
        b_15_, operation, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077;

  AND2_X1 U3569 ( .A1(n3537), .A2(operation), .ZN(Result_9_) );
  AND2_X1 U3570 ( .A1(n3538), .A2(n3539), .ZN(n3537) );
  OR2_X1 U3571 ( .A1(n3540), .A2(n3541), .ZN(n3539) );
  INV_X1 U3572 ( .A(n3542), .ZN(n3538) );
  AND2_X1 U3573 ( .A1(n3541), .A2(n3540), .ZN(n3542) );
  OR2_X1 U3574 ( .A1(n3543), .A2(n3544), .ZN(n3540) );
  AND2_X1 U3575 ( .A1(n3545), .A2(n3546), .ZN(n3544) );
  AND2_X1 U3576 ( .A1(n3547), .A2(n3548), .ZN(n3543) );
  INV_X1 U3577 ( .A(n3546), .ZN(n3547) );
  AND2_X1 U3578 ( .A1(n3549), .A2(operation), .ZN(Result_8_) );
  AND2_X1 U3579 ( .A1(n3550), .A2(n3551), .ZN(n3549) );
  OR2_X1 U3580 ( .A1(n3552), .A2(n3553), .ZN(n3551) );
  OR2_X1 U3581 ( .A1(n3554), .A2(n3555), .ZN(n3553) );
  AND2_X1 U3582 ( .A1(n3556), .A2(n3557), .ZN(n3555) );
  AND2_X1 U3583 ( .A1(n3558), .A2(n3559), .ZN(n3554) );
  OR2_X1 U3584 ( .A1(n3559), .A2(n3560), .ZN(n3550) );
  AND2_X1 U3585 ( .A1(operation), .A2(n3561), .ZN(Result_7_) );
  OR2_X1 U3586 ( .A1(n3562), .A2(n3563), .ZN(n3561) );
  INV_X1 U3587 ( .A(n3564), .ZN(n3563) );
  OR2_X1 U3588 ( .A1(n3565), .A2(n3566), .ZN(n3564) );
  AND2_X1 U3589 ( .A1(n3566), .A2(n3565), .ZN(n3562) );
  OR2_X1 U3590 ( .A1(n3567), .A2(n3568), .ZN(n3565) );
  AND2_X1 U3591 ( .A1(n3569), .A2(n3570), .ZN(n3568) );
  OR2_X1 U3592 ( .A1(n3571), .A2(n3572), .ZN(n3570) );
  AND2_X1 U3593 ( .A1(n3573), .A2(operation), .ZN(Result_6_) );
  AND2_X1 U3594 ( .A1(n3574), .A2(n3575), .ZN(n3573) );
  INV_X1 U3595 ( .A(n3576), .ZN(n3575) );
  AND2_X1 U3596 ( .A1(n3577), .A2(n3578), .ZN(n3576) );
  OR2_X1 U3597 ( .A1(n3577), .A2(n3579), .ZN(n3574) );
  OR2_X1 U3598 ( .A1(n3580), .A2(n3581), .ZN(n3579) );
  AND2_X1 U3599 ( .A1(n3578), .A2(n3582), .ZN(n3581) );
  AND2_X1 U3600 ( .A1(n3583), .A2(n3584), .ZN(n3580) );
  AND2_X1 U3601 ( .A1(operation), .A2(n3585), .ZN(Result_5_) );
  OR2_X1 U3602 ( .A1(n3586), .A2(n3587), .ZN(n3585) );
  INV_X1 U3603 ( .A(n3588), .ZN(n3587) );
  OR2_X1 U3604 ( .A1(n3589), .A2(n3590), .ZN(n3588) );
  AND2_X1 U3605 ( .A1(n3590), .A2(n3589), .ZN(n3586) );
  OR2_X1 U3606 ( .A1(n3591), .A2(n3592), .ZN(n3589) );
  AND2_X1 U3607 ( .A1(n3593), .A2(n3594), .ZN(n3592) );
  OR2_X1 U3608 ( .A1(n3595), .A2(n3596), .ZN(n3594) );
  AND2_X1 U3609 ( .A1(n3597), .A2(operation), .ZN(Result_4_) );
  AND2_X1 U3610 ( .A1(n3598), .A2(n3599), .ZN(n3597) );
  INV_X1 U3611 ( .A(n3600), .ZN(n3599) );
  AND2_X1 U3612 ( .A1(n3601), .A2(n3602), .ZN(n3600) );
  OR2_X1 U3613 ( .A1(n3601), .A2(n3603), .ZN(n3598) );
  OR2_X1 U3614 ( .A1(n3604), .A2(n3605), .ZN(n3603) );
  AND2_X1 U3615 ( .A1(n3602), .A2(n3606), .ZN(n3605) );
  AND2_X1 U3616 ( .A1(n3607), .A2(n3608), .ZN(n3604) );
  AND2_X1 U3617 ( .A1(operation), .A2(n3609), .ZN(Result_3_) );
  OR2_X1 U3618 ( .A1(n3610), .A2(n3611), .ZN(n3609) );
  INV_X1 U3619 ( .A(n3612), .ZN(n3611) );
  OR2_X1 U3620 ( .A1(n3613), .A2(n3614), .ZN(n3612) );
  AND2_X1 U3621 ( .A1(n3614), .A2(n3613), .ZN(n3610) );
  OR2_X1 U3622 ( .A1(n3615), .A2(n3616), .ZN(n3613) );
  AND2_X1 U3623 ( .A1(n3617), .A2(n3618), .ZN(n3616) );
  OR2_X1 U3624 ( .A1(n3619), .A2(n3620), .ZN(n3618) );
  OR2_X1 U3625 ( .A1(n3621), .A2(n3622), .ZN(Result_31_) );
  AND2_X1 U3626 ( .A1(n3623), .A2(operation), .ZN(n3622) );
  AND2_X1 U3627 ( .A1(n3624), .A2(n3625), .ZN(n3621) );
  OR2_X1 U3628 ( .A1(n3626), .A2(n3627), .ZN(n3624) );
  AND2_X1 U3629 ( .A1(b_15_), .A2(n3628), .ZN(n3626) );
  OR2_X1 U3630 ( .A1(n3629), .A2(n3630), .ZN(Result_30_) );
  AND2_X1 U3631 ( .A1(n3631), .A2(n3625), .ZN(n3630) );
  OR2_X1 U3632 ( .A1(n3632), .A2(n3633), .ZN(n3631) );
  AND2_X1 U3633 ( .A1(n3634), .A2(n3635), .ZN(n3633) );
  INV_X1 U3634 ( .A(n3636), .ZN(n3632) );
  OR2_X1 U3635 ( .A1(n3635), .A2(n3634), .ZN(n3636) );
  OR2_X1 U3636 ( .A1(n3637), .A2(n3638), .ZN(n3634) );
  AND2_X1 U3637 ( .A1(b_14_), .A2(n3639), .ZN(n3637) );
  AND2_X1 U3638 ( .A1(operation), .A2(n3640), .ZN(n3629) );
  OR2_X1 U3639 ( .A1(n3641), .A2(n3642), .ZN(n3640) );
  AND2_X1 U3640 ( .A1(b_15_), .A2(n3643), .ZN(n3642) );
  OR2_X1 U3641 ( .A1(n3638), .A2(n3644), .ZN(n3643) );
  AND2_X1 U3642 ( .A1(a_14_), .A2(n3645), .ZN(n3638) );
  AND2_X1 U3643 ( .A1(b_14_), .A2(n3646), .ZN(n3641) );
  OR2_X1 U3644 ( .A1(n3627), .A2(n3647), .ZN(n3646) );
  AND2_X1 U3645 ( .A1(a_15_), .A2(n3648), .ZN(n3627) );
  AND2_X1 U3646 ( .A1(n3649), .A2(operation), .ZN(Result_2_) );
  AND2_X1 U3647 ( .A1(n3650), .A2(n3651), .ZN(n3649) );
  OR2_X1 U3648 ( .A1(n3652), .A2(n3653), .ZN(n3651) );
  OR2_X1 U3649 ( .A1(n3654), .A2(n3655), .ZN(n3650) );
  OR2_X1 U3650 ( .A1(n3656), .A2(n3657), .ZN(n3655) );
  INV_X1 U3651 ( .A(n3658), .ZN(n3657) );
  OR2_X1 U3652 ( .A1(n3653), .A2(n3659), .ZN(n3658) );
  AND2_X1 U3653 ( .A1(n3659), .A2(n3653), .ZN(n3656) );
  OR2_X1 U3654 ( .A1(n3660), .A2(n3661), .ZN(Result_29_) );
  AND2_X1 U3655 ( .A1(n3662), .A2(operation), .ZN(n3661) );
  OR2_X1 U3656 ( .A1(n3663), .A2(n3664), .ZN(n3662) );
  AND2_X1 U3657 ( .A1(n3665), .A2(n3666), .ZN(n3664) );
  INV_X1 U3658 ( .A(n3667), .ZN(n3663) );
  OR2_X1 U3659 ( .A1(n3666), .A2(n3665), .ZN(n3667) );
  AND2_X1 U3660 ( .A1(n3668), .A2(n3669), .ZN(n3665) );
  OR2_X1 U3661 ( .A1(n3670), .A2(n3671), .ZN(n3669) );
  OR2_X1 U3662 ( .A1(n3672), .A2(n3673), .ZN(n3668) );
  INV_X1 U3663 ( .A(n3671), .ZN(n3672) );
  AND2_X1 U3664 ( .A1(n3674), .A2(n3625), .ZN(n3660) );
  OR2_X1 U3665 ( .A1(n3675), .A2(n3676), .ZN(n3674) );
  AND2_X1 U3666 ( .A1(n3677), .A2(n3678), .ZN(n3676) );
  OR2_X1 U3667 ( .A1(n3679), .A2(n3680), .ZN(n3677) );
  AND2_X1 U3668 ( .A1(a_13_), .A2(n3681), .ZN(n3680) );
  AND2_X1 U3669 ( .A1(b_13_), .A2(n3682), .ZN(n3679) );
  AND2_X1 U3670 ( .A1(n3683), .A2(n3684), .ZN(n3675) );
  INV_X1 U3671 ( .A(n3678), .ZN(n3684) );
  OR2_X1 U3672 ( .A1(n3685), .A2(n3686), .ZN(n3683) );
  OR2_X1 U3673 ( .A1(n3687), .A2(n3688), .ZN(Result_28_) );
  AND2_X1 U3674 ( .A1(n3689), .A2(operation), .ZN(n3688) );
  AND2_X1 U3675 ( .A1(n3690), .A2(n3691), .ZN(n3689) );
  INV_X1 U3676 ( .A(n3692), .ZN(n3691) );
  AND2_X1 U3677 ( .A1(n3693), .A2(n3694), .ZN(n3692) );
  OR2_X1 U3678 ( .A1(n3694), .A2(n3693), .ZN(n3690) );
  AND2_X1 U3679 ( .A1(n3695), .A2(n3696), .ZN(n3693) );
  OR2_X1 U3680 ( .A1(n3697), .A2(n3698), .ZN(n3696) );
  INV_X1 U3681 ( .A(n3699), .ZN(n3698) );
  OR2_X1 U3682 ( .A1(n3699), .A2(n3700), .ZN(n3695) );
  INV_X1 U3683 ( .A(n3697), .ZN(n3700) );
  AND2_X1 U3684 ( .A1(n3701), .A2(n3625), .ZN(n3687) );
  OR2_X1 U3685 ( .A1(n3702), .A2(n3703), .ZN(n3701) );
  AND2_X1 U3686 ( .A1(n3704), .A2(n3705), .ZN(n3703) );
  INV_X1 U3687 ( .A(n3706), .ZN(n3705) );
  AND2_X1 U3688 ( .A1(n3707), .A2(n3708), .ZN(n3702) );
  OR2_X1 U3689 ( .A1(n3706), .A2(n3709), .ZN(n3708) );
  INV_X1 U3690 ( .A(n3710), .ZN(n3707) );
  OR2_X1 U3691 ( .A1(n3711), .A2(n3712), .ZN(Result_27_) );
  AND2_X1 U3692 ( .A1(n3713), .A2(operation), .ZN(n3712) );
  AND2_X1 U3693 ( .A1(n3714), .A2(n3715), .ZN(n3713) );
  INV_X1 U3694 ( .A(n3716), .ZN(n3715) );
  AND2_X1 U3695 ( .A1(n3717), .A2(n3718), .ZN(n3716) );
  OR2_X1 U3696 ( .A1(n3718), .A2(n3717), .ZN(n3714) );
  AND2_X1 U3697 ( .A1(n3719), .A2(n3720), .ZN(n3717) );
  INV_X1 U3698 ( .A(n3721), .ZN(n3720) );
  AND2_X1 U3699 ( .A1(n3722), .A2(n3723), .ZN(n3721) );
  OR2_X1 U3700 ( .A1(n3723), .A2(n3722), .ZN(n3719) );
  INV_X1 U3701 ( .A(n3724), .ZN(n3722) );
  AND2_X1 U3702 ( .A1(n3725), .A2(n3625), .ZN(n3711) );
  OR2_X1 U3703 ( .A1(n3726), .A2(n3727), .ZN(n3725) );
  OR2_X1 U3704 ( .A1(n3728), .A2(n3729), .ZN(n3727) );
  AND2_X1 U3705 ( .A1(n3730), .A2(n3731), .ZN(n3729) );
  OR2_X1 U3706 ( .A1(n3732), .A2(n3733), .ZN(n3730) );
  AND2_X1 U3707 ( .A1(n3734), .A2(n3735), .ZN(n3733) );
  AND2_X1 U3708 ( .A1(a_11_), .A2(n3736), .ZN(n3732) );
  AND2_X1 U3709 ( .A1(n3737), .A2(b_11_), .ZN(n3728) );
  AND2_X1 U3710 ( .A1(n3736), .A2(n3735), .ZN(n3737) );
  AND2_X1 U3711 ( .A1(n3734), .A2(n3738), .ZN(n3726) );
  INV_X1 U3712 ( .A(n3736), .ZN(n3734) );
  OR2_X1 U3713 ( .A1(n3739), .A2(n3740), .ZN(Result_26_) );
  AND2_X1 U3714 ( .A1(n3741), .A2(operation), .ZN(n3740) );
  AND2_X1 U3715 ( .A1(n3742), .A2(n3743), .ZN(n3741) );
  INV_X1 U3716 ( .A(n3744), .ZN(n3743) );
  AND2_X1 U3717 ( .A1(n3745), .A2(n3746), .ZN(n3744) );
  OR2_X1 U3718 ( .A1(n3746), .A2(n3745), .ZN(n3742) );
  AND2_X1 U3719 ( .A1(n3747), .A2(n3748), .ZN(n3745) );
  OR2_X1 U3720 ( .A1(n3749), .A2(n3750), .ZN(n3748) );
  INV_X1 U3721 ( .A(n3751), .ZN(n3747) );
  AND2_X1 U3722 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  INV_X1 U3723 ( .A(n3752), .ZN(n3750) );
  AND2_X1 U3724 ( .A1(n3753), .A2(n3625), .ZN(n3739) );
  OR2_X1 U3725 ( .A1(n3754), .A2(n3755), .ZN(n3753) );
  AND2_X1 U3726 ( .A1(n3756), .A2(n3757), .ZN(n3755) );
  INV_X1 U3727 ( .A(n3758), .ZN(n3756) );
  AND2_X1 U3728 ( .A1(n3759), .A2(n3758), .ZN(n3754) );
  OR2_X1 U3729 ( .A1(n3760), .A2(n3761), .ZN(n3758) );
  INV_X1 U3730 ( .A(n3757), .ZN(n3759) );
  OR2_X1 U3731 ( .A1(n3762), .A2(n3763), .ZN(Result_25_) );
  AND2_X1 U3732 ( .A1(n3764), .A2(operation), .ZN(n3763) );
  AND2_X1 U3733 ( .A1(n3765), .A2(n3766), .ZN(n3764) );
  INV_X1 U3734 ( .A(n3767), .ZN(n3766) );
  AND2_X1 U3735 ( .A1(n3768), .A2(n3769), .ZN(n3767) );
  OR2_X1 U3736 ( .A1(n3769), .A2(n3768), .ZN(n3765) );
  AND2_X1 U3737 ( .A1(n3770), .A2(n3771), .ZN(n3768) );
  OR2_X1 U3738 ( .A1(n3772), .A2(n3773), .ZN(n3771) );
  INV_X1 U3739 ( .A(n3774), .ZN(n3773) );
  OR2_X1 U3740 ( .A1(n3774), .A2(n3775), .ZN(n3770) );
  INV_X1 U3741 ( .A(n3772), .ZN(n3775) );
  AND2_X1 U3742 ( .A1(n3776), .A2(n3625), .ZN(n3762) );
  OR2_X1 U3743 ( .A1(n3777), .A2(n3778), .ZN(n3776) );
  OR2_X1 U3744 ( .A1(n3779), .A2(n3780), .ZN(n3778) );
  AND2_X1 U3745 ( .A1(n3781), .A2(n3782), .ZN(n3780) );
  OR2_X1 U3746 ( .A1(n3783), .A2(n3784), .ZN(n3781) );
  AND2_X1 U3747 ( .A1(n3785), .A2(n3786), .ZN(n3784) );
  AND2_X1 U3748 ( .A1(a_9_), .A2(n3787), .ZN(n3783) );
  AND2_X1 U3749 ( .A1(n3788), .A2(b_9_), .ZN(n3779) );
  AND2_X1 U3750 ( .A1(n3787), .A2(n3786), .ZN(n3788) );
  AND2_X1 U3751 ( .A1(n3785), .A2(n3789), .ZN(n3777) );
  INV_X1 U3752 ( .A(n3787), .ZN(n3785) );
  OR2_X1 U3753 ( .A1(n3790), .A2(n3791), .ZN(Result_24_) );
  AND2_X1 U3754 ( .A1(n3792), .A2(operation), .ZN(n3791) );
  AND2_X1 U3755 ( .A1(n3793), .A2(n3794), .ZN(n3792) );
  INV_X1 U3756 ( .A(n3795), .ZN(n3794) );
  AND2_X1 U3757 ( .A1(n3796), .A2(n3797), .ZN(n3795) );
  OR2_X1 U3758 ( .A1(n3797), .A2(n3796), .ZN(n3793) );
  AND2_X1 U3759 ( .A1(n3798), .A2(n3799), .ZN(n3796) );
  OR2_X1 U3760 ( .A1(n3800), .A2(n3801), .ZN(n3799) );
  INV_X1 U3761 ( .A(n3802), .ZN(n3801) );
  OR2_X1 U3762 ( .A1(n3802), .A2(n3803), .ZN(n3798) );
  INV_X1 U3763 ( .A(n3800), .ZN(n3803) );
  AND2_X1 U3764 ( .A1(n3804), .A2(n3625), .ZN(n3790) );
  OR2_X1 U3765 ( .A1(n3805), .A2(n3806), .ZN(n3804) );
  AND2_X1 U3766 ( .A1(n3807), .A2(n3808), .ZN(n3806) );
  INV_X1 U3767 ( .A(n3809), .ZN(n3805) );
  OR2_X1 U3768 ( .A1(n3808), .A2(n3807), .ZN(n3809) );
  AND2_X1 U3769 ( .A1(n3810), .A2(n3811), .ZN(n3807) );
  INV_X1 U3770 ( .A(n3812), .ZN(n3810) );
  OR2_X1 U3771 ( .A1(n3813), .A2(n3814), .ZN(Result_23_) );
  AND2_X1 U3772 ( .A1(n3815), .A2(operation), .ZN(n3814) );
  AND2_X1 U3773 ( .A1(n3816), .A2(n3817), .ZN(n3815) );
  INV_X1 U3774 ( .A(n3818), .ZN(n3817) );
  AND2_X1 U3775 ( .A1(n3819), .A2(n3820), .ZN(n3818) );
  OR2_X1 U3776 ( .A1(n3820), .A2(n3819), .ZN(n3816) );
  AND2_X1 U3777 ( .A1(n3821), .A2(n3822), .ZN(n3819) );
  OR2_X1 U3778 ( .A1(n3823), .A2(n3824), .ZN(n3822) );
  INV_X1 U3779 ( .A(n3825), .ZN(n3824) );
  OR2_X1 U3780 ( .A1(n3825), .A2(n3826), .ZN(n3821) );
  INV_X1 U3781 ( .A(n3823), .ZN(n3826) );
  AND2_X1 U3782 ( .A1(n3827), .A2(n3625), .ZN(n3813) );
  OR2_X1 U3783 ( .A1(n3828), .A2(n3829), .ZN(n3827) );
  OR2_X1 U3784 ( .A1(n3830), .A2(n3831), .ZN(n3829) );
  AND2_X1 U3785 ( .A1(n3832), .A2(n3833), .ZN(n3831) );
  OR2_X1 U3786 ( .A1(n3834), .A2(n3835), .ZN(n3832) );
  AND2_X1 U3787 ( .A1(n3836), .A2(n3837), .ZN(n3835) );
  AND2_X1 U3788 ( .A1(a_7_), .A2(n3838), .ZN(n3834) );
  AND2_X1 U3789 ( .A1(n3839), .A2(b_7_), .ZN(n3830) );
  AND2_X1 U3790 ( .A1(n3838), .A2(n3837), .ZN(n3839) );
  AND2_X1 U3791 ( .A1(n3836), .A2(n3840), .ZN(n3828) );
  INV_X1 U3792 ( .A(n3838), .ZN(n3836) );
  OR2_X1 U3793 ( .A1(n3841), .A2(n3842), .ZN(Result_22_) );
  AND2_X1 U3794 ( .A1(n3843), .A2(operation), .ZN(n3842) );
  AND2_X1 U3795 ( .A1(n3844), .A2(n3845), .ZN(n3843) );
  INV_X1 U3796 ( .A(n3846), .ZN(n3845) );
  AND2_X1 U3797 ( .A1(n3847), .A2(n3848), .ZN(n3846) );
  OR2_X1 U3798 ( .A1(n3848), .A2(n3847), .ZN(n3844) );
  AND2_X1 U3799 ( .A1(n3849), .A2(n3850), .ZN(n3847) );
  OR2_X1 U3800 ( .A1(n3851), .A2(n3852), .ZN(n3850) );
  INV_X1 U3801 ( .A(n3853), .ZN(n3852) );
  OR2_X1 U3802 ( .A1(n3853), .A2(n3854), .ZN(n3849) );
  INV_X1 U3803 ( .A(n3851), .ZN(n3854) );
  AND2_X1 U3804 ( .A1(n3855), .A2(n3625), .ZN(n3841) );
  OR2_X1 U3805 ( .A1(n3856), .A2(n3857), .ZN(n3855) );
  AND2_X1 U3806 ( .A1(n3858), .A2(n3859), .ZN(n3857) );
  INV_X1 U3807 ( .A(n3860), .ZN(n3856) );
  OR2_X1 U3808 ( .A1(n3859), .A2(n3858), .ZN(n3860) );
  AND2_X1 U3809 ( .A1(n3861), .A2(n3862), .ZN(n3858) );
  INV_X1 U3810 ( .A(n3863), .ZN(n3861) );
  OR2_X1 U3811 ( .A1(n3864), .A2(n3865), .ZN(Result_21_) );
  AND2_X1 U3812 ( .A1(n3866), .A2(operation), .ZN(n3865) );
  AND2_X1 U3813 ( .A1(n3867), .A2(n3868), .ZN(n3866) );
  INV_X1 U3814 ( .A(n3869), .ZN(n3868) );
  AND2_X1 U3815 ( .A1(n3870), .A2(n3871), .ZN(n3869) );
  OR2_X1 U3816 ( .A1(n3871), .A2(n3870), .ZN(n3867) );
  AND2_X1 U3817 ( .A1(n3872), .A2(n3873), .ZN(n3870) );
  OR2_X1 U3818 ( .A1(n3874), .A2(n3875), .ZN(n3873) );
  INV_X1 U3819 ( .A(n3876), .ZN(n3875) );
  OR2_X1 U3820 ( .A1(n3876), .A2(n3877), .ZN(n3872) );
  INV_X1 U3821 ( .A(n3874), .ZN(n3877) );
  AND2_X1 U3822 ( .A1(n3878), .A2(n3625), .ZN(n3864) );
  OR2_X1 U3823 ( .A1(n3879), .A2(n3880), .ZN(n3878) );
  OR2_X1 U3824 ( .A1(n3881), .A2(n3882), .ZN(n3880) );
  AND2_X1 U3825 ( .A1(n3883), .A2(n3884), .ZN(n3882) );
  OR2_X1 U3826 ( .A1(n3885), .A2(n3886), .ZN(n3883) );
  AND2_X1 U3827 ( .A1(n3887), .A2(n3888), .ZN(n3886) );
  AND2_X1 U3828 ( .A1(a_5_), .A2(n3889), .ZN(n3885) );
  AND2_X1 U3829 ( .A1(n3890), .A2(b_5_), .ZN(n3881) );
  AND2_X1 U3830 ( .A1(n3889), .A2(n3888), .ZN(n3890) );
  AND2_X1 U3831 ( .A1(n3887), .A2(n3891), .ZN(n3879) );
  INV_X1 U3832 ( .A(n3889), .ZN(n3887) );
  OR2_X1 U3833 ( .A1(n3892), .A2(n3893), .ZN(Result_20_) );
  AND2_X1 U3834 ( .A1(n3894), .A2(operation), .ZN(n3893) );
  AND2_X1 U3835 ( .A1(n3895), .A2(n3896), .ZN(n3894) );
  INV_X1 U3836 ( .A(n3897), .ZN(n3896) );
  AND2_X1 U3837 ( .A1(n3898), .A2(n3899), .ZN(n3897) );
  OR2_X1 U3838 ( .A1(n3899), .A2(n3898), .ZN(n3895) );
  AND2_X1 U3839 ( .A1(n3900), .A2(n3901), .ZN(n3898) );
  OR2_X1 U3840 ( .A1(n3902), .A2(n3903), .ZN(n3901) );
  INV_X1 U3841 ( .A(n3904), .ZN(n3903) );
  OR2_X1 U3842 ( .A1(n3904), .A2(n3905), .ZN(n3900) );
  INV_X1 U3843 ( .A(n3902), .ZN(n3905) );
  AND2_X1 U3844 ( .A1(n3906), .A2(n3625), .ZN(n3892) );
  OR2_X1 U3845 ( .A1(n3907), .A2(n3908), .ZN(n3906) );
  AND2_X1 U3846 ( .A1(n3909), .A2(n3910), .ZN(n3908) );
  INV_X1 U3847 ( .A(n3911), .ZN(n3907) );
  OR2_X1 U3848 ( .A1(n3910), .A2(n3909), .ZN(n3911) );
  AND2_X1 U3849 ( .A1(n3912), .A2(n3913), .ZN(n3909) );
  INV_X1 U3850 ( .A(n3914), .ZN(n3912) );
  AND2_X1 U3851 ( .A1(operation), .A2(n3915), .ZN(Result_1_) );
  OR2_X1 U3852 ( .A1(n3916), .A2(n3917), .ZN(n3915) );
  AND2_X1 U3853 ( .A1(n3918), .A2(n3919), .ZN(n3917) );
  AND2_X1 U3854 ( .A1(n3920), .A2(n3921), .ZN(n3916) );
  INV_X1 U3855 ( .A(n3918), .ZN(n3921) );
  AND2_X1 U3856 ( .A1(n3922), .A2(n3923), .ZN(n3918) );
  OR2_X1 U3857 ( .A1(n3924), .A2(n3925), .ZN(n3923) );
  INV_X1 U3858 ( .A(n3926), .ZN(n3922) );
  OR2_X1 U3859 ( .A1(n3927), .A2(n3928), .ZN(Result_19_) );
  AND2_X1 U3860 ( .A1(n3929), .A2(operation), .ZN(n3928) );
  AND2_X1 U3861 ( .A1(n3930), .A2(n3931), .ZN(n3929) );
  INV_X1 U3862 ( .A(n3932), .ZN(n3931) );
  AND2_X1 U3863 ( .A1(n3933), .A2(n3934), .ZN(n3932) );
  OR2_X1 U3864 ( .A1(n3934), .A2(n3933), .ZN(n3930) );
  AND2_X1 U3865 ( .A1(n3935), .A2(n3936), .ZN(n3933) );
  OR2_X1 U3866 ( .A1(n3937), .A2(n3938), .ZN(n3936) );
  INV_X1 U3867 ( .A(n3939), .ZN(n3938) );
  OR2_X1 U3868 ( .A1(n3939), .A2(n3940), .ZN(n3935) );
  INV_X1 U3869 ( .A(n3937), .ZN(n3940) );
  AND2_X1 U3870 ( .A1(n3941), .A2(n3625), .ZN(n3927) );
  OR2_X1 U3871 ( .A1(n3942), .A2(n3943), .ZN(n3941) );
  OR2_X1 U3872 ( .A1(n3944), .A2(n3945), .ZN(n3943) );
  AND2_X1 U3873 ( .A1(n3946), .A2(n3947), .ZN(n3945) );
  OR2_X1 U3874 ( .A1(n3948), .A2(n3949), .ZN(n3946) );
  AND2_X1 U3875 ( .A1(n3950), .A2(n3951), .ZN(n3949) );
  AND2_X1 U3876 ( .A1(a_3_), .A2(n3952), .ZN(n3948) );
  AND2_X1 U3877 ( .A1(n3953), .A2(b_3_), .ZN(n3944) );
  AND2_X1 U3878 ( .A1(n3952), .A2(n3951), .ZN(n3953) );
  AND2_X1 U3879 ( .A1(n3950), .A2(n3954), .ZN(n3942) );
  INV_X1 U3880 ( .A(n3952), .ZN(n3950) );
  OR2_X1 U3881 ( .A1(n3955), .A2(n3956), .ZN(Result_18_) );
  AND2_X1 U3882 ( .A1(n3957), .A2(operation), .ZN(n3956) );
  AND2_X1 U3883 ( .A1(n3958), .A2(n3959), .ZN(n3957) );
  INV_X1 U3884 ( .A(n3960), .ZN(n3959) );
  AND2_X1 U3885 ( .A1(n3961), .A2(n3962), .ZN(n3960) );
  OR2_X1 U3886 ( .A1(n3962), .A2(n3961), .ZN(n3958) );
  AND2_X1 U3887 ( .A1(n3963), .A2(n3964), .ZN(n3961) );
  OR2_X1 U3888 ( .A1(n3965), .A2(n3966), .ZN(n3964) );
  INV_X1 U3889 ( .A(n3967), .ZN(n3966) );
  OR2_X1 U3890 ( .A1(n3967), .A2(n3968), .ZN(n3963) );
  INV_X1 U3891 ( .A(n3965), .ZN(n3968) );
  AND2_X1 U3892 ( .A1(n3969), .A2(n3625), .ZN(n3955) );
  OR2_X1 U3893 ( .A1(n3970), .A2(n3971), .ZN(n3969) );
  AND2_X1 U3894 ( .A1(n3972), .A2(n3973), .ZN(n3971) );
  INV_X1 U3895 ( .A(n3974), .ZN(n3970) );
  OR2_X1 U3896 ( .A1(n3973), .A2(n3972), .ZN(n3974) );
  AND2_X1 U3897 ( .A1(n3975), .A2(n3976), .ZN(n3972) );
  INV_X1 U3898 ( .A(n3977), .ZN(n3975) );
  OR2_X1 U3899 ( .A1(n3978), .A2(n3979), .ZN(Result_17_) );
  AND2_X1 U3900 ( .A1(n3980), .A2(operation), .ZN(n3979) );
  AND2_X1 U3901 ( .A1(n3981), .A2(n3982), .ZN(n3980) );
  INV_X1 U3902 ( .A(n3983), .ZN(n3982) );
  AND2_X1 U3903 ( .A1(n3984), .A2(n3985), .ZN(n3983) );
  OR2_X1 U3904 ( .A1(n3985), .A2(n3984), .ZN(n3981) );
  AND2_X1 U3905 ( .A1(n3986), .A2(n3987), .ZN(n3984) );
  OR2_X1 U3906 ( .A1(n3988), .A2(n3989), .ZN(n3987) );
  INV_X1 U3907 ( .A(n3990), .ZN(n3989) );
  OR2_X1 U3908 ( .A1(n3990), .A2(n3991), .ZN(n3986) );
  INV_X1 U3909 ( .A(n3988), .ZN(n3991) );
  AND2_X1 U3910 ( .A1(n3992), .A2(n3625), .ZN(n3978) );
  OR2_X1 U3911 ( .A1(n3993), .A2(n3994), .ZN(n3992) );
  OR2_X1 U3912 ( .A1(n3995), .A2(n3996), .ZN(n3994) );
  AND2_X1 U3913 ( .A1(n3997), .A2(n3998), .ZN(n3996) );
  OR2_X1 U3914 ( .A1(n3999), .A2(n4000), .ZN(n3997) );
  AND2_X1 U3915 ( .A1(n4001), .A2(n4002), .ZN(n4000) );
  AND2_X1 U3916 ( .A1(a_1_), .A2(n4003), .ZN(n3999) );
  AND2_X1 U3917 ( .A1(n4004), .A2(b_1_), .ZN(n3995) );
  AND2_X1 U3918 ( .A1(n4003), .A2(n4002), .ZN(n4004) );
  AND2_X1 U3919 ( .A1(n4001), .A2(n4005), .ZN(n3993) );
  INV_X1 U3920 ( .A(n4003), .ZN(n4001) );
  OR2_X1 U3921 ( .A1(n4006), .A2(n4007), .ZN(Result_16_) );
  AND2_X1 U3922 ( .A1(n4008), .A2(operation), .ZN(n4007) );
  AND2_X1 U3923 ( .A1(n4009), .A2(n4010), .ZN(n4008) );
  INV_X1 U3924 ( .A(n4011), .ZN(n4010) );
  AND2_X1 U3925 ( .A1(n4012), .A2(n4013), .ZN(n4011) );
  OR2_X1 U3926 ( .A1(n4013), .A2(n4012), .ZN(n4009) );
  AND2_X1 U3927 ( .A1(n4014), .A2(n4015), .ZN(n4012) );
  OR2_X1 U3928 ( .A1(n4016), .A2(n4017), .ZN(n4015) );
  INV_X1 U3929 ( .A(n4018), .ZN(n4017) );
  OR2_X1 U3930 ( .A1(n4018), .A2(n4019), .ZN(n4014) );
  AND2_X1 U3931 ( .A1(n4020), .A2(n3625), .ZN(n4006) );
  INV_X1 U3932 ( .A(operation), .ZN(n3625) );
  OR2_X1 U3933 ( .A1(n4021), .A2(n4022), .ZN(n4020) );
  INV_X1 U3934 ( .A(n4023), .ZN(n4022) );
  OR2_X1 U3935 ( .A1(n4024), .A2(n4025), .ZN(n4023) );
  AND2_X1 U3936 ( .A1(n4025), .A2(n4024), .ZN(n4021) );
  AND2_X1 U3937 ( .A1(n4026), .A2(n4027), .ZN(n4024) );
  OR2_X1 U3938 ( .A1(n4028), .A2(b_0_), .ZN(n4027) );
  OR2_X1 U3939 ( .A1(n4029), .A2(a_0_), .ZN(n4026) );
  INV_X1 U3940 ( .A(n4030), .ZN(n4025) );
  OR2_X1 U3941 ( .A1(n4031), .A2(n4032), .ZN(n4030) );
  AND2_X1 U3942 ( .A1(n4002), .A2(n3998), .ZN(n4032) );
  AND2_X1 U3943 ( .A1(n4003), .A2(n4033), .ZN(n4031) );
  OR2_X1 U3944 ( .A1(n4034), .A2(n3977), .ZN(n4003) );
  AND2_X1 U3945 ( .A1(n4035), .A2(n4036), .ZN(n3977) );
  AND2_X1 U3946 ( .A1(n3973), .A2(n3976), .ZN(n4034) );
  OR2_X1 U3947 ( .A1(n4037), .A2(n4038), .ZN(n3973) );
  AND2_X1 U3948 ( .A1(n3951), .A2(n3947), .ZN(n4038) );
  AND2_X1 U3949 ( .A1(n3952), .A2(n4039), .ZN(n4037) );
  OR2_X1 U3950 ( .A1(n4040), .A2(n3914), .ZN(n3952) );
  AND2_X1 U3951 ( .A1(n4041), .A2(n4042), .ZN(n3914) );
  AND2_X1 U3952 ( .A1(n3910), .A2(n3913), .ZN(n4040) );
  OR2_X1 U3953 ( .A1(n4043), .A2(n4044), .ZN(n3910) );
  AND2_X1 U3954 ( .A1(n3888), .A2(n3884), .ZN(n4044) );
  AND2_X1 U3955 ( .A1(n3889), .A2(n4045), .ZN(n4043) );
  OR2_X1 U3956 ( .A1(n4046), .A2(n3863), .ZN(n3889) );
  AND2_X1 U3957 ( .A1(n4047), .A2(n4048), .ZN(n3863) );
  AND2_X1 U3958 ( .A1(n3859), .A2(n3862), .ZN(n4046) );
  OR2_X1 U3959 ( .A1(n4049), .A2(n4050), .ZN(n3859) );
  AND2_X1 U3960 ( .A1(n3837), .A2(n3833), .ZN(n4050) );
  AND2_X1 U3961 ( .A1(n3838), .A2(n4051), .ZN(n4049) );
  OR2_X1 U3962 ( .A1(n4052), .A2(n3812), .ZN(n3838) );
  AND2_X1 U3963 ( .A1(n4053), .A2(n4054), .ZN(n3812) );
  AND2_X1 U3964 ( .A1(n3808), .A2(n3811), .ZN(n4052) );
  OR2_X1 U3965 ( .A1(n4055), .A2(n4056), .ZN(n3808) );
  AND2_X1 U3966 ( .A1(n3786), .A2(n3782), .ZN(n4056) );
  AND2_X1 U3967 ( .A1(n3787), .A2(n4057), .ZN(n4055) );
  OR2_X1 U3968 ( .A1(n4058), .A2(n3760), .ZN(n3787) );
  AND2_X1 U3969 ( .A1(n4059), .A2(n4060), .ZN(n3760) );
  AND2_X1 U3970 ( .A1(n3757), .A2(n4061), .ZN(n4058) );
  OR2_X1 U3971 ( .A1(n4062), .A2(n4063), .ZN(n3757) );
  AND2_X1 U3972 ( .A1(n3735), .A2(n3731), .ZN(n4063) );
  AND2_X1 U3973 ( .A1(n4064), .A2(n3736), .ZN(n4062) );
  OR2_X1 U3974 ( .A1(n3706), .A2(n3704), .ZN(n3736) );
  AND2_X1 U3975 ( .A1(n3710), .A2(n4065), .ZN(n3704) );
  OR2_X1 U3976 ( .A1(n3686), .A2(n4066), .ZN(n3710) );
  AND2_X1 U3977 ( .A1(n3678), .A2(n4067), .ZN(n4066) );
  AND2_X1 U3978 ( .A1(n4068), .A2(n4069), .ZN(n3678) );
  OR2_X1 U3979 ( .A1(n3648), .A2(n4070), .ZN(n4069) );
  OR2_X1 U3980 ( .A1(n3645), .A2(n4071), .ZN(n4068) );
  AND2_X1 U3981 ( .A1(n3635), .A2(n3639), .ZN(n4071) );
  INV_X1 U3982 ( .A(n3623), .ZN(n3635) );
  AND2_X1 U3983 ( .A1(a_15_), .A2(b_15_), .ZN(n3623) );
  AND2_X1 U3984 ( .A1(n3682), .A2(n3681), .ZN(n3686) );
  AND2_X1 U3985 ( .A1(n4072), .A2(n4073), .ZN(n3706) );
  AND2_X1 U3986 ( .A1(operation), .A2(n4074), .ZN(Result_15_) );
  OR2_X1 U3987 ( .A1(n4075), .A2(n4076), .ZN(n4074) );
  AND2_X1 U3988 ( .A1(n4077), .A2(n4078), .ZN(n4076) );
  AND2_X1 U3989 ( .A1(n4079), .A2(n4080), .ZN(n4075) );
  AND2_X1 U3990 ( .A1(n4081), .A2(operation), .ZN(Result_14_) );
  AND2_X1 U3991 ( .A1(n4082), .A2(n4083), .ZN(n4081) );
  OR2_X1 U3992 ( .A1(n4084), .A2(n4085), .ZN(n4082) );
  AND2_X1 U3993 ( .A1(n4080), .A2(n4077), .ZN(n4084) );
  AND2_X1 U3994 ( .A1(operation), .A2(n4086), .ZN(Result_13_) );
  OR2_X1 U3995 ( .A1(n4087), .A2(n4088), .ZN(n4086) );
  AND2_X1 U3996 ( .A1(n4089), .A2(n4090), .ZN(n4088) );
  INV_X1 U3997 ( .A(n4091), .ZN(n4087) );
  OR2_X1 U3998 ( .A1(n4089), .A2(n4090), .ZN(n4091) );
  OR2_X1 U3999 ( .A1(n4092), .A2(n4093), .ZN(n4089) );
  AND2_X1 U4000 ( .A1(n4094), .A2(n4083), .ZN(n4093) );
  INV_X1 U4001 ( .A(n4095), .ZN(n4083) );
  AND2_X1 U4002 ( .A1(n4095), .A2(n4096), .ZN(n4092) );
  AND2_X1 U4003 ( .A1(n4097), .A2(operation), .ZN(Result_12_) );
  AND2_X1 U4004 ( .A1(n4098), .A2(n4099), .ZN(n4097) );
  OR2_X1 U4005 ( .A1(n4100), .A2(n4101), .ZN(n4099) );
  INV_X1 U4006 ( .A(n4102), .ZN(n4101) );
  OR2_X1 U4007 ( .A1(n4103), .A2(n4102), .ZN(n4098) );
  AND2_X1 U4008 ( .A1(n4104), .A2(n4105), .ZN(n4102) );
  INV_X1 U4009 ( .A(n4106), .ZN(n4105) );
  OR2_X1 U4010 ( .A1(n4107), .A2(n4108), .ZN(n4104) );
  AND2_X1 U4011 ( .A1(n4109), .A2(operation), .ZN(Result_11_) );
  AND2_X1 U4012 ( .A1(n4110), .A2(n4111), .ZN(n4109) );
  OR2_X1 U4013 ( .A1(n4112), .A2(n4113), .ZN(n4111) );
  INV_X1 U4014 ( .A(n4114), .ZN(n4113) );
  OR2_X1 U4015 ( .A1(n4115), .A2(n4114), .ZN(n4110) );
  AND2_X1 U4016 ( .A1(n4116), .A2(n4117), .ZN(n4114) );
  INV_X1 U4017 ( .A(n4118), .ZN(n4117) );
  OR2_X1 U4018 ( .A1(n4119), .A2(n4120), .ZN(n4116) );
  AND2_X1 U4019 ( .A1(n4121), .A2(operation), .ZN(Result_10_) );
  AND2_X1 U4020 ( .A1(n4122), .A2(n4123), .ZN(n4121) );
  OR2_X1 U4021 ( .A1(n4124), .A2(n4125), .ZN(n4123) );
  INV_X1 U4022 ( .A(n4126), .ZN(n4125) );
  OR2_X1 U4023 ( .A1(n4127), .A2(n4126), .ZN(n4122) );
  AND2_X1 U4024 ( .A1(n4128), .A2(n4129), .ZN(n4126) );
  INV_X1 U4025 ( .A(n4130), .ZN(n4129) );
  OR2_X1 U4026 ( .A1(n4131), .A2(n4132), .ZN(n4128) );
  AND2_X1 U4027 ( .A1(operation), .A2(n4133), .ZN(Result_0_) );
  OR2_X1 U4028 ( .A1(n4134), .A2(n4135), .ZN(n4133) );
  OR2_X1 U4029 ( .A1(n3926), .A2(n4136), .ZN(n4135) );
  AND2_X1 U4030 ( .A1(n3920), .A2(n3924), .ZN(n4136) );
  INV_X1 U4031 ( .A(n3919), .ZN(n3920) );
  OR2_X1 U4032 ( .A1(n4137), .A2(n3653), .ZN(n3919) );
  OR2_X1 U4033 ( .A1(n4138), .A2(n3925), .ZN(n3653) );
  AND2_X1 U4034 ( .A1(n4139), .A2(n4140), .ZN(n4138) );
  AND2_X1 U4035 ( .A1(n3652), .A2(n4141), .ZN(n4137) );
  INV_X1 U4036 ( .A(n3654), .ZN(n3652) );
  OR2_X1 U4037 ( .A1(n4142), .A2(n3615), .ZN(n3654) );
  AND2_X1 U4038 ( .A1(n4143), .A2(n4144), .ZN(n3615) );
  AND2_X1 U4039 ( .A1(n4145), .A2(n4146), .ZN(n4144) );
  AND2_X1 U4040 ( .A1(n3614), .A2(n4143), .ZN(n4142) );
  INV_X1 U4041 ( .A(n3617), .ZN(n4143) );
  OR2_X1 U4042 ( .A1(n3659), .A2(n4147), .ZN(n3617) );
  AND2_X1 U4043 ( .A1(n4148), .A2(n4149), .ZN(n4147) );
  INV_X1 U4044 ( .A(n4141), .ZN(n3659) );
  OR2_X1 U4045 ( .A1(n4148), .A2(n4149), .ZN(n4141) );
  OR2_X1 U4046 ( .A1(n4150), .A2(n4151), .ZN(n4149) );
  AND2_X1 U4047 ( .A1(n4152), .A2(n4153), .ZN(n4151) );
  AND2_X1 U4048 ( .A1(n4154), .A2(n4155), .ZN(n4150) );
  OR2_X1 U4049 ( .A1(n4153), .A2(n4152), .ZN(n4155) );
  INV_X1 U4050 ( .A(n4156), .ZN(n4152) );
  AND2_X1 U4051 ( .A1(n4157), .A2(n4158), .ZN(n4148) );
  OR2_X1 U4052 ( .A1(n4159), .A2(n4160), .ZN(n4158) );
  INV_X1 U4053 ( .A(n4161), .ZN(n4159) );
  OR2_X1 U4054 ( .A1(n4162), .A2(n4161), .ZN(n4157) );
  AND2_X1 U4055 ( .A1(n4163), .A2(n4164), .ZN(n4161) );
  OR2_X1 U4056 ( .A1(n4165), .A2(n4166), .ZN(n4164) );
  INV_X1 U4057 ( .A(n4167), .ZN(n4163) );
  AND2_X1 U4058 ( .A1(n4166), .A2(n4165), .ZN(n4167) );
  INV_X1 U4059 ( .A(n4168), .ZN(n4166) );
  AND2_X1 U4060 ( .A1(n4169), .A2(n3602), .ZN(n3614) );
  INV_X1 U4061 ( .A(n3608), .ZN(n3602) );
  AND2_X1 U4062 ( .A1(n4170), .A2(n4171), .ZN(n3608) );
  OR2_X1 U4063 ( .A1(n3619), .A2(n4146), .ZN(n4171) );
  INV_X1 U4064 ( .A(n3620), .ZN(n4146) );
  OR2_X1 U4065 ( .A1(n4145), .A2(n3620), .ZN(n4170) );
  OR2_X1 U4066 ( .A1(n4172), .A2(n4173), .ZN(n3620) );
  AND2_X1 U4067 ( .A1(n4174), .A2(n4175), .ZN(n4173) );
  AND2_X1 U4068 ( .A1(n4176), .A2(n4177), .ZN(n4172) );
  OR2_X1 U4069 ( .A1(n4175), .A2(n4174), .ZN(n4177) );
  INV_X1 U4070 ( .A(n3619), .ZN(n4145) );
  AND2_X1 U4071 ( .A1(n4178), .A2(n4179), .ZN(n3619) );
  INV_X1 U4072 ( .A(n4180), .ZN(n4179) );
  AND2_X1 U4073 ( .A1(n4181), .A2(n4154), .ZN(n4180) );
  OR2_X1 U4074 ( .A1(n4154), .A2(n4181), .ZN(n4178) );
  OR2_X1 U4075 ( .A1(n4182), .A2(n4183), .ZN(n4181) );
  AND2_X1 U4076 ( .A1(n4156), .A2(n4153), .ZN(n4183) );
  INV_X1 U4077 ( .A(n4184), .ZN(n4182) );
  OR2_X1 U4078 ( .A1(n4153), .A2(n4156), .ZN(n4184) );
  AND2_X1 U4079 ( .A1(b_3_), .A2(a_0_), .ZN(n4156) );
  OR2_X1 U4080 ( .A1(n4185), .A2(n4186), .ZN(n4153) );
  AND2_X1 U4081 ( .A1(n4187), .A2(n4188), .ZN(n4186) );
  AND2_X1 U4082 ( .A1(n4189), .A2(n4190), .ZN(n4185) );
  OR2_X1 U4083 ( .A1(n4188), .A2(n4187), .ZN(n4190) );
  AND2_X1 U4084 ( .A1(n4191), .A2(n4192), .ZN(n4154) );
  INV_X1 U4085 ( .A(n4193), .ZN(n4192) );
  AND2_X1 U4086 ( .A1(n4194), .A2(n4195), .ZN(n4193) );
  OR2_X1 U4087 ( .A1(n4195), .A2(n4194), .ZN(n4191) );
  OR2_X1 U4088 ( .A1(n4196), .A2(n4197), .ZN(n4194) );
  AND2_X1 U4089 ( .A1(n4198), .A2(n4199), .ZN(n4197) );
  INV_X1 U4090 ( .A(n4200), .ZN(n4198) );
  AND2_X1 U4091 ( .A1(n4201), .A2(n4200), .ZN(n4196) );
  INV_X1 U4092 ( .A(n4199), .ZN(n4201) );
  OR2_X1 U4093 ( .A1(n3601), .A2(n3607), .ZN(n4169) );
  OR2_X1 U4094 ( .A1(n4202), .A2(n3591), .ZN(n3601) );
  AND2_X1 U4095 ( .A1(n4203), .A2(n4204), .ZN(n3591) );
  AND2_X1 U4096 ( .A1(n4205), .A2(n4206), .ZN(n4204) );
  AND2_X1 U4097 ( .A1(n3590), .A2(n4203), .ZN(n4202) );
  INV_X1 U4098 ( .A(n3593), .ZN(n4203) );
  OR2_X1 U4099 ( .A1(n3607), .A2(n4207), .ZN(n3593) );
  AND2_X1 U4100 ( .A1(n4208), .A2(n4209), .ZN(n4207) );
  INV_X1 U4101 ( .A(n3606), .ZN(n3607) );
  OR2_X1 U4102 ( .A1(n4208), .A2(n4209), .ZN(n3606) );
  OR2_X1 U4103 ( .A1(n4210), .A2(n4211), .ZN(n4209) );
  AND2_X1 U4104 ( .A1(n4212), .A2(n4213), .ZN(n4211) );
  AND2_X1 U4105 ( .A1(n4214), .A2(n4215), .ZN(n4210) );
  OR2_X1 U4106 ( .A1(n4213), .A2(n4212), .ZN(n4215) );
  INV_X1 U4107 ( .A(n4216), .ZN(n4212) );
  AND2_X1 U4108 ( .A1(n4217), .A2(n4218), .ZN(n4208) );
  OR2_X1 U4109 ( .A1(n4219), .A2(n4176), .ZN(n4218) );
  INV_X1 U4110 ( .A(n4220), .ZN(n4219) );
  OR2_X1 U4111 ( .A1(n4221), .A2(n4220), .ZN(n4217) );
  AND2_X1 U4112 ( .A1(n4222), .A2(n4223), .ZN(n4220) );
  OR2_X1 U4113 ( .A1(n4174), .A2(n4224), .ZN(n4223) );
  INV_X1 U4114 ( .A(n4225), .ZN(n4222) );
  AND2_X1 U4115 ( .A1(n4224), .A2(n4174), .ZN(n4225) );
  OR2_X1 U4116 ( .A1(n4042), .A2(n4028), .ZN(n4174) );
  INV_X1 U4117 ( .A(n4175), .ZN(n4224) );
  OR2_X1 U4118 ( .A1(n4226), .A2(n4227), .ZN(n4175) );
  AND2_X1 U4119 ( .A1(n4228), .A2(n4229), .ZN(n4227) );
  AND2_X1 U4120 ( .A1(n4230), .A2(n4231), .ZN(n4226) );
  OR2_X1 U4121 ( .A1(n4229), .A2(n4228), .ZN(n4231) );
  INV_X1 U4122 ( .A(n4176), .ZN(n4221) );
  AND2_X1 U4123 ( .A1(n4232), .A2(n4233), .ZN(n4176) );
  INV_X1 U4124 ( .A(n4234), .ZN(n4233) );
  AND2_X1 U4125 ( .A1(n4235), .A2(n4189), .ZN(n4234) );
  OR2_X1 U4126 ( .A1(n4189), .A2(n4235), .ZN(n4232) );
  OR2_X1 U4127 ( .A1(n4236), .A2(n4237), .ZN(n4235) );
  AND2_X1 U4128 ( .A1(n4238), .A2(n4188), .ZN(n4237) );
  INV_X1 U4129 ( .A(n4187), .ZN(n4238) );
  AND2_X1 U4130 ( .A1(n4239), .A2(n4187), .ZN(n4236) );
  OR2_X1 U4131 ( .A1(n3947), .A2(n4002), .ZN(n4187) );
  INV_X1 U4132 ( .A(n4188), .ZN(n4239) );
  OR2_X1 U4133 ( .A1(n4240), .A2(n4241), .ZN(n4188) );
  AND2_X1 U4134 ( .A1(n4242), .A2(n4243), .ZN(n4241) );
  AND2_X1 U4135 ( .A1(n4244), .A2(n4245), .ZN(n4240) );
  OR2_X1 U4136 ( .A1(n4243), .A2(n4242), .ZN(n4245) );
  AND2_X1 U4137 ( .A1(n4246), .A2(n4247), .ZN(n4189) );
  INV_X1 U4138 ( .A(n4248), .ZN(n4247) );
  AND2_X1 U4139 ( .A1(n4249), .A2(n4250), .ZN(n4248) );
  OR2_X1 U4140 ( .A1(n4250), .A2(n4249), .ZN(n4246) );
  OR2_X1 U4141 ( .A1(n4251), .A2(n4252), .ZN(n4249) );
  AND2_X1 U4142 ( .A1(n4253), .A2(n4254), .ZN(n4252) );
  INV_X1 U4143 ( .A(n4255), .ZN(n4251) );
  OR2_X1 U4144 ( .A1(n4254), .A2(n4253), .ZN(n4255) );
  AND2_X1 U4145 ( .A1(n4256), .A2(n3578), .ZN(n3590) );
  INV_X1 U4146 ( .A(n3584), .ZN(n3578) );
  AND2_X1 U4147 ( .A1(n4257), .A2(n4258), .ZN(n3584) );
  OR2_X1 U4148 ( .A1(n3595), .A2(n4206), .ZN(n4258) );
  INV_X1 U4149 ( .A(n3596), .ZN(n4206) );
  OR2_X1 U4150 ( .A1(n4205), .A2(n3596), .ZN(n4257) );
  OR2_X1 U4151 ( .A1(n4259), .A2(n4260), .ZN(n3596) );
  AND2_X1 U4152 ( .A1(n4261), .A2(n4262), .ZN(n4260) );
  AND2_X1 U4153 ( .A1(n4263), .A2(n4264), .ZN(n4259) );
  OR2_X1 U4154 ( .A1(n4262), .A2(n4261), .ZN(n4264) );
  INV_X1 U4155 ( .A(n3595), .ZN(n4205) );
  AND2_X1 U4156 ( .A1(n4265), .A2(n4266), .ZN(n3595) );
  INV_X1 U4157 ( .A(n4267), .ZN(n4266) );
  AND2_X1 U4158 ( .A1(n4268), .A2(n4214), .ZN(n4267) );
  OR2_X1 U4159 ( .A1(n4214), .A2(n4268), .ZN(n4265) );
  OR2_X1 U4160 ( .A1(n4269), .A2(n4270), .ZN(n4268) );
  AND2_X1 U4161 ( .A1(n4216), .A2(n4213), .ZN(n4270) );
  INV_X1 U4162 ( .A(n4271), .ZN(n4269) );
  OR2_X1 U4163 ( .A1(n4213), .A2(n4216), .ZN(n4271) );
  AND2_X1 U4164 ( .A1(b_5_), .A2(a_0_), .ZN(n4216) );
  OR2_X1 U4165 ( .A1(n4272), .A2(n4273), .ZN(n4213) );
  AND2_X1 U4166 ( .A1(n4274), .A2(n4275), .ZN(n4273) );
  AND2_X1 U4167 ( .A1(n4276), .A2(n4277), .ZN(n4272) );
  OR2_X1 U4168 ( .A1(n4275), .A2(n4274), .ZN(n4277) );
  AND2_X1 U4169 ( .A1(n4278), .A2(n4279), .ZN(n4214) );
  INV_X1 U4170 ( .A(n4280), .ZN(n4279) );
  AND2_X1 U4171 ( .A1(n4281), .A2(n4230), .ZN(n4280) );
  OR2_X1 U4172 ( .A1(n4230), .A2(n4281), .ZN(n4278) );
  OR2_X1 U4173 ( .A1(n4282), .A2(n4283), .ZN(n4281) );
  AND2_X1 U4174 ( .A1(n4284), .A2(n4229), .ZN(n4283) );
  INV_X1 U4175 ( .A(n4228), .ZN(n4284) );
  AND2_X1 U4176 ( .A1(n4285), .A2(n4228), .ZN(n4282) );
  OR2_X1 U4177 ( .A1(n4042), .A2(n4002), .ZN(n4228) );
  INV_X1 U4178 ( .A(n4229), .ZN(n4285) );
  OR2_X1 U4179 ( .A1(n4286), .A2(n4287), .ZN(n4229) );
  AND2_X1 U4180 ( .A1(n4288), .A2(n4289), .ZN(n4287) );
  AND2_X1 U4181 ( .A1(n4290), .A2(n4291), .ZN(n4286) );
  OR2_X1 U4182 ( .A1(n4289), .A2(n4288), .ZN(n4291) );
  AND2_X1 U4183 ( .A1(n4292), .A2(n4293), .ZN(n4230) );
  INV_X1 U4184 ( .A(n4294), .ZN(n4293) );
  AND2_X1 U4185 ( .A1(n4295), .A2(n4244), .ZN(n4294) );
  OR2_X1 U4186 ( .A1(n4244), .A2(n4295), .ZN(n4292) );
  OR2_X1 U4187 ( .A1(n4296), .A2(n4297), .ZN(n4295) );
  AND2_X1 U4188 ( .A1(n4298), .A2(n4243), .ZN(n4297) );
  INV_X1 U4189 ( .A(n4242), .ZN(n4298) );
  AND2_X1 U4190 ( .A1(n4299), .A2(n4242), .ZN(n4296) );
  OR2_X1 U4191 ( .A1(n3947), .A2(n4035), .ZN(n4242) );
  INV_X1 U4192 ( .A(n4243), .ZN(n4299) );
  OR2_X1 U4193 ( .A1(n4300), .A2(n4301), .ZN(n4243) );
  AND2_X1 U4194 ( .A1(n4039), .A2(n4302), .ZN(n4301) );
  AND2_X1 U4195 ( .A1(n4303), .A2(n4304), .ZN(n4300) );
  OR2_X1 U4196 ( .A1(n4302), .A2(n4039), .ZN(n4304) );
  AND2_X1 U4197 ( .A1(n4305), .A2(n4306), .ZN(n4244) );
  INV_X1 U4198 ( .A(n4307), .ZN(n4306) );
  AND2_X1 U4199 ( .A1(n4308), .A2(n4309), .ZN(n4307) );
  OR2_X1 U4200 ( .A1(n4309), .A2(n4308), .ZN(n4305) );
  OR2_X1 U4201 ( .A1(n4310), .A2(n4311), .ZN(n4308) );
  AND2_X1 U4202 ( .A1(n4312), .A2(n4313), .ZN(n4311) );
  INV_X1 U4203 ( .A(n4314), .ZN(n4312) );
  AND2_X1 U4204 ( .A1(n4315), .A2(n4314), .ZN(n4310) );
  INV_X1 U4205 ( .A(n4313), .ZN(n4315) );
  OR2_X1 U4206 ( .A1(n3577), .A2(n3583), .ZN(n4256) );
  OR2_X1 U4207 ( .A1(n4316), .A2(n3567), .ZN(n3577) );
  AND2_X1 U4208 ( .A1(n4317), .A2(n4318), .ZN(n3567) );
  AND2_X1 U4209 ( .A1(n4319), .A2(n4320), .ZN(n4318) );
  AND2_X1 U4210 ( .A1(n3566), .A2(n4317), .ZN(n4316) );
  INV_X1 U4211 ( .A(n3569), .ZN(n4317) );
  OR2_X1 U4212 ( .A1(n3583), .A2(n4321), .ZN(n3569) );
  AND2_X1 U4213 ( .A1(n4322), .A2(n4323), .ZN(n4321) );
  INV_X1 U4214 ( .A(n3582), .ZN(n3583) );
  OR2_X1 U4215 ( .A1(n4322), .A2(n4323), .ZN(n3582) );
  OR2_X1 U4216 ( .A1(n4324), .A2(n4325), .ZN(n4323) );
  AND2_X1 U4217 ( .A1(n4326), .A2(n4327), .ZN(n4325) );
  AND2_X1 U4218 ( .A1(n4328), .A2(n4329), .ZN(n4324) );
  OR2_X1 U4219 ( .A1(n4327), .A2(n4326), .ZN(n4329) );
  INV_X1 U4220 ( .A(n4330), .ZN(n4326) );
  AND2_X1 U4221 ( .A1(n4331), .A2(n4332), .ZN(n4322) );
  OR2_X1 U4222 ( .A1(n4333), .A2(n4263), .ZN(n4332) );
  INV_X1 U4223 ( .A(n4334), .ZN(n4333) );
  OR2_X1 U4224 ( .A1(n4335), .A2(n4334), .ZN(n4331) );
  AND2_X1 U4225 ( .A1(n4336), .A2(n4337), .ZN(n4334) );
  OR2_X1 U4226 ( .A1(n4261), .A2(n4338), .ZN(n4337) );
  INV_X1 U4227 ( .A(n4339), .ZN(n4336) );
  AND2_X1 U4228 ( .A1(n4338), .A2(n4261), .ZN(n4339) );
  OR2_X1 U4229 ( .A1(n4048), .A2(n4028), .ZN(n4261) );
  INV_X1 U4230 ( .A(n4262), .ZN(n4338) );
  OR2_X1 U4231 ( .A1(n4340), .A2(n4341), .ZN(n4262) );
  AND2_X1 U4232 ( .A1(n4342), .A2(n4343), .ZN(n4341) );
  AND2_X1 U4233 ( .A1(n4344), .A2(n4345), .ZN(n4340) );
  OR2_X1 U4234 ( .A1(n4343), .A2(n4342), .ZN(n4345) );
  INV_X1 U4235 ( .A(n4263), .ZN(n4335) );
  AND2_X1 U4236 ( .A1(n4346), .A2(n4347), .ZN(n4263) );
  INV_X1 U4237 ( .A(n4348), .ZN(n4347) );
  AND2_X1 U4238 ( .A1(n4349), .A2(n4276), .ZN(n4348) );
  OR2_X1 U4239 ( .A1(n4276), .A2(n4349), .ZN(n4346) );
  OR2_X1 U4240 ( .A1(n4350), .A2(n4351), .ZN(n4349) );
  AND2_X1 U4241 ( .A1(n4352), .A2(n4275), .ZN(n4351) );
  INV_X1 U4242 ( .A(n4274), .ZN(n4352) );
  AND2_X1 U4243 ( .A1(n4353), .A2(n4274), .ZN(n4350) );
  OR2_X1 U4244 ( .A1(n3884), .A2(n4002), .ZN(n4274) );
  INV_X1 U4245 ( .A(n4275), .ZN(n4353) );
  OR2_X1 U4246 ( .A1(n4354), .A2(n4355), .ZN(n4275) );
  AND2_X1 U4247 ( .A1(n4356), .A2(n4357), .ZN(n4355) );
  AND2_X1 U4248 ( .A1(n4358), .A2(n4359), .ZN(n4354) );
  OR2_X1 U4249 ( .A1(n4357), .A2(n4356), .ZN(n4359) );
  AND2_X1 U4250 ( .A1(n4360), .A2(n4361), .ZN(n4276) );
  INV_X1 U4251 ( .A(n4362), .ZN(n4361) );
  AND2_X1 U4252 ( .A1(n4363), .A2(n4290), .ZN(n4362) );
  OR2_X1 U4253 ( .A1(n4290), .A2(n4363), .ZN(n4360) );
  OR2_X1 U4254 ( .A1(n4364), .A2(n4365), .ZN(n4363) );
  AND2_X1 U4255 ( .A1(n4366), .A2(n4289), .ZN(n4365) );
  INV_X1 U4256 ( .A(n4288), .ZN(n4366) );
  AND2_X1 U4257 ( .A1(n4367), .A2(n4288), .ZN(n4364) );
  OR2_X1 U4258 ( .A1(n4042), .A2(n4035), .ZN(n4288) );
  INV_X1 U4259 ( .A(n4289), .ZN(n4367) );
  OR2_X1 U4260 ( .A1(n4368), .A2(n4369), .ZN(n4289) );
  AND2_X1 U4261 ( .A1(n4370), .A2(n4371), .ZN(n4369) );
  AND2_X1 U4262 ( .A1(n4372), .A2(n4373), .ZN(n4368) );
  OR2_X1 U4263 ( .A1(n4371), .A2(n4370), .ZN(n4373) );
  AND2_X1 U4264 ( .A1(n4374), .A2(n4375), .ZN(n4290) );
  INV_X1 U4265 ( .A(n4376), .ZN(n4375) );
  AND2_X1 U4266 ( .A1(n4377), .A2(n4303), .ZN(n4376) );
  OR2_X1 U4267 ( .A1(n4303), .A2(n4377), .ZN(n4374) );
  OR2_X1 U4268 ( .A1(n4378), .A2(n4379), .ZN(n4377) );
  AND2_X1 U4269 ( .A1(n3954), .A2(n4302), .ZN(n4379) );
  INV_X1 U4270 ( .A(n4039), .ZN(n3954) );
  AND2_X1 U4271 ( .A1(n4380), .A2(n4039), .ZN(n4378) );
  OR2_X1 U4272 ( .A1(n3947), .A2(n3951), .ZN(n4039) );
  INV_X1 U4273 ( .A(n4302), .ZN(n4380) );
  OR2_X1 U4274 ( .A1(n4381), .A2(n4382), .ZN(n4302) );
  AND2_X1 U4275 ( .A1(n4383), .A2(n4384), .ZN(n4382) );
  AND2_X1 U4276 ( .A1(n4385), .A2(n4386), .ZN(n4381) );
  OR2_X1 U4277 ( .A1(n4384), .A2(n4383), .ZN(n4386) );
  AND2_X1 U4278 ( .A1(n4387), .A2(n4388), .ZN(n4303) );
  INV_X1 U4279 ( .A(n4389), .ZN(n4388) );
  AND2_X1 U4280 ( .A1(n4390), .A2(n4391), .ZN(n4389) );
  OR2_X1 U4281 ( .A1(n4391), .A2(n4390), .ZN(n4387) );
  OR2_X1 U4282 ( .A1(n4392), .A2(n4393), .ZN(n4390) );
  AND2_X1 U4283 ( .A1(n4394), .A2(n4395), .ZN(n4393) );
  INV_X1 U4284 ( .A(n4396), .ZN(n4394) );
  AND2_X1 U4285 ( .A1(n4397), .A2(n4396), .ZN(n4392) );
  INV_X1 U4286 ( .A(n4395), .ZN(n4397) );
  AND2_X1 U4287 ( .A1(n4398), .A2(n3556), .ZN(n3566) );
  INV_X1 U4288 ( .A(n3559), .ZN(n3556) );
  AND2_X1 U4289 ( .A1(n4399), .A2(n4400), .ZN(n3559) );
  OR2_X1 U4290 ( .A1(n3571), .A2(n4320), .ZN(n4400) );
  INV_X1 U4291 ( .A(n3572), .ZN(n4320) );
  OR2_X1 U4292 ( .A1(n4319), .A2(n3572), .ZN(n4399) );
  OR2_X1 U4293 ( .A1(n4401), .A2(n4402), .ZN(n3572) );
  AND2_X1 U4294 ( .A1(n4403), .A2(n4404), .ZN(n4402) );
  AND2_X1 U4295 ( .A1(n4405), .A2(n4406), .ZN(n4401) );
  OR2_X1 U4296 ( .A1(n4404), .A2(n4403), .ZN(n4406) );
  INV_X1 U4297 ( .A(n3571), .ZN(n4319) );
  AND2_X1 U4298 ( .A1(n4407), .A2(n4408), .ZN(n3571) );
  INV_X1 U4299 ( .A(n4409), .ZN(n4408) );
  AND2_X1 U4300 ( .A1(n4410), .A2(n4328), .ZN(n4409) );
  OR2_X1 U4301 ( .A1(n4328), .A2(n4410), .ZN(n4407) );
  OR2_X1 U4302 ( .A1(n4411), .A2(n4412), .ZN(n4410) );
  AND2_X1 U4303 ( .A1(n4330), .A2(n4327), .ZN(n4412) );
  INV_X1 U4304 ( .A(n4413), .ZN(n4411) );
  OR2_X1 U4305 ( .A1(n4327), .A2(n4330), .ZN(n4413) );
  AND2_X1 U4306 ( .A1(b_7_), .A2(a_0_), .ZN(n4330) );
  OR2_X1 U4307 ( .A1(n4414), .A2(n4415), .ZN(n4327) );
  AND2_X1 U4308 ( .A1(n4416), .A2(n4417), .ZN(n4415) );
  AND2_X1 U4309 ( .A1(n4418), .A2(n4419), .ZN(n4414) );
  OR2_X1 U4310 ( .A1(n4417), .A2(n4416), .ZN(n4419) );
  AND2_X1 U4311 ( .A1(n4420), .A2(n4421), .ZN(n4328) );
  INV_X1 U4312 ( .A(n4422), .ZN(n4421) );
  AND2_X1 U4313 ( .A1(n4423), .A2(n4344), .ZN(n4422) );
  OR2_X1 U4314 ( .A1(n4344), .A2(n4423), .ZN(n4420) );
  OR2_X1 U4315 ( .A1(n4424), .A2(n4425), .ZN(n4423) );
  AND2_X1 U4316 ( .A1(n4426), .A2(n4343), .ZN(n4425) );
  INV_X1 U4317 ( .A(n4342), .ZN(n4426) );
  AND2_X1 U4318 ( .A1(n4427), .A2(n4342), .ZN(n4424) );
  OR2_X1 U4319 ( .A1(n4048), .A2(n4002), .ZN(n4342) );
  INV_X1 U4320 ( .A(n4343), .ZN(n4427) );
  OR2_X1 U4321 ( .A1(n4428), .A2(n4429), .ZN(n4343) );
  AND2_X1 U4322 ( .A1(n4430), .A2(n4431), .ZN(n4429) );
  AND2_X1 U4323 ( .A1(n4432), .A2(n4433), .ZN(n4428) );
  OR2_X1 U4324 ( .A1(n4431), .A2(n4430), .ZN(n4433) );
  AND2_X1 U4325 ( .A1(n4434), .A2(n4435), .ZN(n4344) );
  INV_X1 U4326 ( .A(n4436), .ZN(n4435) );
  AND2_X1 U4327 ( .A1(n4437), .A2(n4358), .ZN(n4436) );
  OR2_X1 U4328 ( .A1(n4358), .A2(n4437), .ZN(n4434) );
  OR2_X1 U4329 ( .A1(n4438), .A2(n4439), .ZN(n4437) );
  AND2_X1 U4330 ( .A1(n4440), .A2(n4357), .ZN(n4439) );
  INV_X1 U4331 ( .A(n4356), .ZN(n4440) );
  AND2_X1 U4332 ( .A1(n4441), .A2(n4356), .ZN(n4438) );
  OR2_X1 U4333 ( .A1(n3884), .A2(n4035), .ZN(n4356) );
  INV_X1 U4334 ( .A(n4357), .ZN(n4441) );
  OR2_X1 U4335 ( .A1(n4442), .A2(n4443), .ZN(n4357) );
  AND2_X1 U4336 ( .A1(n4444), .A2(n4445), .ZN(n4443) );
  AND2_X1 U4337 ( .A1(n4446), .A2(n4447), .ZN(n4442) );
  OR2_X1 U4338 ( .A1(n4445), .A2(n4444), .ZN(n4447) );
  AND2_X1 U4339 ( .A1(n4448), .A2(n4449), .ZN(n4358) );
  INV_X1 U4340 ( .A(n4450), .ZN(n4449) );
  AND2_X1 U4341 ( .A1(n4451), .A2(n4372), .ZN(n4450) );
  OR2_X1 U4342 ( .A1(n4372), .A2(n4451), .ZN(n4448) );
  OR2_X1 U4343 ( .A1(n4452), .A2(n4453), .ZN(n4451) );
  AND2_X1 U4344 ( .A1(n4454), .A2(n4371), .ZN(n4453) );
  INV_X1 U4345 ( .A(n4370), .ZN(n4454) );
  AND2_X1 U4346 ( .A1(n4455), .A2(n4370), .ZN(n4452) );
  OR2_X1 U4347 ( .A1(n4042), .A2(n3951), .ZN(n4370) );
  INV_X1 U4348 ( .A(n4371), .ZN(n4455) );
  OR2_X1 U4349 ( .A1(n4456), .A2(n4457), .ZN(n4371) );
  AND2_X1 U4350 ( .A1(n3913), .A2(n4458), .ZN(n4457) );
  AND2_X1 U4351 ( .A1(n4459), .A2(n4460), .ZN(n4456) );
  OR2_X1 U4352 ( .A1(n4458), .A2(n3913), .ZN(n4460) );
  INV_X1 U4353 ( .A(n4461), .ZN(n3913) );
  AND2_X1 U4354 ( .A1(n4462), .A2(n4463), .ZN(n4372) );
  INV_X1 U4355 ( .A(n4464), .ZN(n4463) );
  AND2_X1 U4356 ( .A1(n4465), .A2(n4385), .ZN(n4464) );
  OR2_X1 U4357 ( .A1(n4385), .A2(n4465), .ZN(n4462) );
  OR2_X1 U4358 ( .A1(n4466), .A2(n4467), .ZN(n4465) );
  AND2_X1 U4359 ( .A1(n4468), .A2(n4384), .ZN(n4467) );
  INV_X1 U4360 ( .A(n4383), .ZN(n4468) );
  AND2_X1 U4361 ( .A1(n4469), .A2(n4383), .ZN(n4466) );
  OR2_X1 U4362 ( .A1(n3947), .A2(n4041), .ZN(n4383) );
  INV_X1 U4363 ( .A(n4384), .ZN(n4469) );
  OR2_X1 U4364 ( .A1(n4470), .A2(n4471), .ZN(n4384) );
  AND2_X1 U4365 ( .A1(n4472), .A2(n4473), .ZN(n4471) );
  AND2_X1 U4366 ( .A1(n4474), .A2(n4475), .ZN(n4470) );
  OR2_X1 U4367 ( .A1(n4473), .A2(n4472), .ZN(n4475) );
  AND2_X1 U4368 ( .A1(n4476), .A2(n4477), .ZN(n4385) );
  INV_X1 U4369 ( .A(n4478), .ZN(n4477) );
  AND2_X1 U4370 ( .A1(n4479), .A2(n4480), .ZN(n4478) );
  OR2_X1 U4371 ( .A1(n4480), .A2(n4479), .ZN(n4476) );
  OR2_X1 U4372 ( .A1(n4481), .A2(n4482), .ZN(n4479) );
  AND2_X1 U4373 ( .A1(n4483), .A2(n4484), .ZN(n4482) );
  INV_X1 U4374 ( .A(n4485), .ZN(n4483) );
  AND2_X1 U4375 ( .A1(n4486), .A2(n4485), .ZN(n4481) );
  INV_X1 U4376 ( .A(n4484), .ZN(n4486) );
  OR2_X1 U4377 ( .A1(n3558), .A2(n3552), .ZN(n4398) );
  INV_X1 U4378 ( .A(n3560), .ZN(n3552) );
  OR2_X1 U4379 ( .A1(n4487), .A2(n3546), .ZN(n3560) );
  OR2_X1 U4380 ( .A1(n3558), .A2(n4488), .ZN(n3546) );
  AND2_X1 U4381 ( .A1(n4489), .A2(n4490), .ZN(n4488) );
  AND2_X1 U4382 ( .A1(n3545), .A2(n3541), .ZN(n4487) );
  INV_X1 U4383 ( .A(n3548), .ZN(n3545) );
  OR2_X1 U4384 ( .A1(n4130), .A2(n4491), .ZN(n3548) );
  AND2_X1 U4385 ( .A1(n4127), .A2(n4132), .ZN(n4491) );
  INV_X1 U4386 ( .A(n4124), .ZN(n4127) );
  AND2_X1 U4387 ( .A1(n4132), .A2(n4131), .ZN(n4130) );
  OR2_X1 U4388 ( .A1(n4118), .A2(n4492), .ZN(n4131) );
  AND2_X1 U4389 ( .A1(n4115), .A2(n4120), .ZN(n4492) );
  INV_X1 U4390 ( .A(n4112), .ZN(n4115) );
  AND2_X1 U4391 ( .A1(n4120), .A2(n4119), .ZN(n4118) );
  OR2_X1 U4392 ( .A1(n4106), .A2(n4493), .ZN(n4119) );
  AND2_X1 U4393 ( .A1(n4103), .A2(n4108), .ZN(n4493) );
  AND2_X1 U4394 ( .A1(n4108), .A2(n4107), .ZN(n4106) );
  OR2_X1 U4395 ( .A1(n4494), .A2(n4495), .ZN(n4107) );
  INV_X1 U4396 ( .A(n4496), .ZN(n4495) );
  OR2_X1 U4397 ( .A1(n4090), .A2(n4096), .ZN(n4496) );
  AND2_X1 U4398 ( .A1(n4095), .A2(n4094), .ZN(n4494) );
  INV_X1 U4399 ( .A(n4096), .ZN(n4094) );
  OR2_X1 U4400 ( .A1(n4497), .A2(n4103), .ZN(n4096) );
  INV_X1 U4401 ( .A(n4100), .ZN(n4103) );
  OR2_X1 U4402 ( .A1(n4498), .A2(n4499), .ZN(n4100) );
  AND2_X1 U4403 ( .A1(n4498), .A2(n4499), .ZN(n4497) );
  OR2_X1 U4404 ( .A1(n4500), .A2(n4501), .ZN(n4499) );
  AND2_X1 U4405 ( .A1(n4502), .A2(n4503), .ZN(n4501) );
  AND2_X1 U4406 ( .A1(n4504), .A2(n4505), .ZN(n4500) );
  OR2_X1 U4407 ( .A1(n4503), .A2(n4502), .ZN(n4505) );
  AND2_X1 U4408 ( .A1(n4506), .A2(n4507), .ZN(n4498) );
  INV_X1 U4409 ( .A(n4508), .ZN(n4507) );
  AND2_X1 U4410 ( .A1(n4509), .A2(n4510), .ZN(n4508) );
  OR2_X1 U4411 ( .A1(n4510), .A2(n4509), .ZN(n4506) );
  OR2_X1 U4412 ( .A1(n4511), .A2(n4512), .ZN(n4509) );
  AND2_X1 U4413 ( .A1(n4513), .A2(n4514), .ZN(n4512) );
  INV_X1 U4414 ( .A(n4515), .ZN(n4511) );
  OR2_X1 U4415 ( .A1(n4514), .A2(n4513), .ZN(n4515) );
  AND2_X1 U4416 ( .A1(n4080), .A2(n4516), .ZN(n4095) );
  AND2_X1 U4417 ( .A1(n4085), .A2(n4077), .ZN(n4516) );
  INV_X1 U4418 ( .A(n4079), .ZN(n4077) );
  AND2_X1 U4419 ( .A1(n4517), .A2(n4518), .ZN(n4079) );
  INV_X1 U4420 ( .A(n4519), .ZN(n4518) );
  AND2_X1 U4421 ( .A1(n4520), .A2(n4521), .ZN(n4519) );
  OR2_X1 U4422 ( .A1(n4521), .A2(n4520), .ZN(n4517) );
  OR2_X1 U4423 ( .A1(n4522), .A2(n4523), .ZN(n4520) );
  AND2_X1 U4424 ( .A1(n4524), .A2(n4525), .ZN(n4523) );
  INV_X1 U4425 ( .A(n4526), .ZN(n4522) );
  OR2_X1 U4426 ( .A1(n4525), .A2(n4524), .ZN(n4526) );
  AND2_X1 U4427 ( .A1(n4090), .A2(n4527), .ZN(n4085) );
  INV_X1 U4428 ( .A(n4528), .ZN(n4527) );
  AND2_X1 U4429 ( .A1(n4529), .A2(n4530), .ZN(n4528) );
  OR2_X1 U4430 ( .A1(n4529), .A2(n4530), .ZN(n4090) );
  OR2_X1 U4431 ( .A1(n4531), .A2(n4532), .ZN(n4530) );
  AND2_X1 U4432 ( .A1(n4533), .A2(n4525), .ZN(n4532) );
  AND2_X1 U4433 ( .A1(n4521), .A2(n4534), .ZN(n4531) );
  OR2_X1 U4434 ( .A1(n4533), .A2(n4525), .ZN(n4534) );
  OR2_X1 U4435 ( .A1(n4535), .A2(n4536), .ZN(n4525) );
  AND2_X1 U4436 ( .A1(n4537), .A2(n4538), .ZN(n4536) );
  AND2_X1 U4437 ( .A1(n4539), .A2(n4540), .ZN(n4535) );
  OR2_X1 U4438 ( .A1(n4538), .A2(n4537), .ZN(n4540) );
  INV_X1 U4439 ( .A(n4524), .ZN(n4533) );
  AND2_X1 U4440 ( .A1(a_0_), .A2(b_14_), .ZN(n4524) );
  AND2_X1 U4441 ( .A1(n4541), .A2(n4542), .ZN(n4521) );
  INV_X1 U4442 ( .A(n4543), .ZN(n4542) );
  AND2_X1 U4443 ( .A1(n4544), .A2(n4545), .ZN(n4543) );
  OR2_X1 U4444 ( .A1(n4545), .A2(n4544), .ZN(n4541) );
  OR2_X1 U4445 ( .A1(n4546), .A2(n4547), .ZN(n4544) );
  AND2_X1 U4446 ( .A1(n4548), .A2(n4549), .ZN(n4547) );
  INV_X1 U4447 ( .A(n4550), .ZN(n4548) );
  AND2_X1 U4448 ( .A1(n4551), .A2(n4550), .ZN(n4546) );
  INV_X1 U4449 ( .A(n4549), .ZN(n4551) );
  OR2_X1 U4450 ( .A1(n4552), .A2(n4553), .ZN(n4529) );
  INV_X1 U4451 ( .A(n4554), .ZN(n4553) );
  OR2_X1 U4452 ( .A1(n4555), .A2(n4504), .ZN(n4554) );
  AND2_X1 U4453 ( .A1(n4504), .A2(n4555), .ZN(n4552) );
  AND2_X1 U4454 ( .A1(n4556), .A2(n4557), .ZN(n4555) );
  OR2_X1 U4455 ( .A1(n4502), .A2(n4558), .ZN(n4557) );
  INV_X1 U4456 ( .A(n4503), .ZN(n4558) );
  INV_X1 U4457 ( .A(n4559), .ZN(n4502) );
  OR2_X1 U4458 ( .A1(n4503), .A2(n4559), .ZN(n4556) );
  AND2_X1 U4459 ( .A1(a_0_), .A2(b_13_), .ZN(n4559) );
  OR2_X1 U4460 ( .A1(n4560), .A2(n4561), .ZN(n4503) );
  AND2_X1 U4461 ( .A1(n4550), .A2(n4549), .ZN(n4561) );
  AND2_X1 U4462 ( .A1(n4545), .A2(n4562), .ZN(n4560) );
  OR2_X1 U4463 ( .A1(n4549), .A2(n4550), .ZN(n4562) );
  OR2_X1 U4464 ( .A1(n4002), .A2(n3681), .ZN(n4550) );
  OR2_X1 U4465 ( .A1(n4563), .A2(n4564), .ZN(n4549) );
  AND2_X1 U4466 ( .A1(n4565), .A2(n4566), .ZN(n4564) );
  AND2_X1 U4467 ( .A1(n4567), .A2(n4568), .ZN(n4563) );
  OR2_X1 U4468 ( .A1(n4566), .A2(n4565), .ZN(n4568) );
  AND2_X1 U4469 ( .A1(n4569), .A2(n4570), .ZN(n4545) );
  INV_X1 U4470 ( .A(n4571), .ZN(n4570) );
  AND2_X1 U4471 ( .A1(n4572), .A2(n4573), .ZN(n4571) );
  OR2_X1 U4472 ( .A1(n4573), .A2(n4572), .ZN(n4569) );
  OR2_X1 U4473 ( .A1(n4574), .A2(n4575), .ZN(n4572) );
  AND2_X1 U4474 ( .A1(n4576), .A2(n4577), .ZN(n4575) );
  INV_X1 U4475 ( .A(n4578), .ZN(n4576) );
  AND2_X1 U4476 ( .A1(n4579), .A2(n4578), .ZN(n4574) );
  INV_X1 U4477 ( .A(n4577), .ZN(n4579) );
  OR2_X1 U4478 ( .A1(n4580), .A2(n4581), .ZN(n4504) );
  INV_X1 U4479 ( .A(n4582), .ZN(n4581) );
  OR2_X1 U4480 ( .A1(n4583), .A2(n4584), .ZN(n4582) );
  AND2_X1 U4481 ( .A1(n4584), .A2(n4583), .ZN(n4580) );
  AND2_X1 U4482 ( .A1(n4585), .A2(n4586), .ZN(n4583) );
  OR2_X1 U4483 ( .A1(n4587), .A2(n4588), .ZN(n4586) );
  INV_X1 U4484 ( .A(n4589), .ZN(n4588) );
  OR2_X1 U4485 ( .A1(n4589), .A2(n4590), .ZN(n4585) );
  INV_X1 U4486 ( .A(n4587), .ZN(n4590) );
  INV_X1 U4487 ( .A(n4078), .ZN(n4080) );
  OR2_X1 U4488 ( .A1(n4591), .A2(n4592), .ZN(n4078) );
  AND2_X1 U4489 ( .A1(n4016), .A2(n4018), .ZN(n4592) );
  AND2_X1 U4490 ( .A1(n4013), .A2(n4593), .ZN(n4591) );
  OR2_X1 U4491 ( .A1(n4016), .A2(n4018), .ZN(n4593) );
  OR2_X1 U4492 ( .A1(n4594), .A2(n4595), .ZN(n4018) );
  AND2_X1 U4493 ( .A1(n3988), .A2(n3990), .ZN(n4595) );
  AND2_X1 U4494 ( .A1(n3985), .A2(n4596), .ZN(n4594) );
  OR2_X1 U4495 ( .A1(n3988), .A2(n3990), .ZN(n4596) );
  OR2_X1 U4496 ( .A1(n4597), .A2(n4598), .ZN(n3990) );
  AND2_X1 U4497 ( .A1(n3965), .A2(n3967), .ZN(n4598) );
  AND2_X1 U4498 ( .A1(n3962), .A2(n4599), .ZN(n4597) );
  OR2_X1 U4499 ( .A1(n3965), .A2(n3967), .ZN(n4599) );
  OR2_X1 U4500 ( .A1(n4600), .A2(n4601), .ZN(n3967) );
  AND2_X1 U4501 ( .A1(n3937), .A2(n3939), .ZN(n4601) );
  AND2_X1 U4502 ( .A1(n3934), .A2(n4602), .ZN(n4600) );
  OR2_X1 U4503 ( .A1(n3937), .A2(n3939), .ZN(n4602) );
  OR2_X1 U4504 ( .A1(n4603), .A2(n4604), .ZN(n3939) );
  AND2_X1 U4505 ( .A1(n3902), .A2(n3904), .ZN(n4604) );
  AND2_X1 U4506 ( .A1(n3899), .A2(n4605), .ZN(n4603) );
  OR2_X1 U4507 ( .A1(n3902), .A2(n3904), .ZN(n4605) );
  OR2_X1 U4508 ( .A1(n4606), .A2(n4607), .ZN(n3904) );
  AND2_X1 U4509 ( .A1(n3874), .A2(n3876), .ZN(n4607) );
  AND2_X1 U4510 ( .A1(n3871), .A2(n4608), .ZN(n4606) );
  OR2_X1 U4511 ( .A1(n3874), .A2(n3876), .ZN(n4608) );
  OR2_X1 U4512 ( .A1(n4609), .A2(n4610), .ZN(n3876) );
  AND2_X1 U4513 ( .A1(n3851), .A2(n3853), .ZN(n4610) );
  AND2_X1 U4514 ( .A1(n3848), .A2(n4611), .ZN(n4609) );
  OR2_X1 U4515 ( .A1(n3851), .A2(n3853), .ZN(n4611) );
  OR2_X1 U4516 ( .A1(n4612), .A2(n4613), .ZN(n3853) );
  AND2_X1 U4517 ( .A1(n3823), .A2(n3825), .ZN(n4613) );
  AND2_X1 U4518 ( .A1(n3820), .A2(n4614), .ZN(n4612) );
  OR2_X1 U4519 ( .A1(n3823), .A2(n3825), .ZN(n4614) );
  OR2_X1 U4520 ( .A1(n4615), .A2(n4616), .ZN(n3825) );
  AND2_X1 U4521 ( .A1(n3800), .A2(n3802), .ZN(n4616) );
  AND2_X1 U4522 ( .A1(n3797), .A2(n4617), .ZN(n4615) );
  OR2_X1 U4523 ( .A1(n3800), .A2(n3802), .ZN(n4617) );
  OR2_X1 U4524 ( .A1(n4618), .A2(n4619), .ZN(n3802) );
  AND2_X1 U4525 ( .A1(n3772), .A2(n3774), .ZN(n4619) );
  AND2_X1 U4526 ( .A1(n3769), .A2(n4620), .ZN(n4618) );
  OR2_X1 U4527 ( .A1(n3772), .A2(n3774), .ZN(n4620) );
  OR2_X1 U4528 ( .A1(n4621), .A2(n4622), .ZN(n3774) );
  AND2_X1 U4529 ( .A1(n3749), .A2(n3752), .ZN(n4622) );
  AND2_X1 U4530 ( .A1(n3746), .A2(n4623), .ZN(n4621) );
  OR2_X1 U4531 ( .A1(n3749), .A2(n3752), .ZN(n4623) );
  OR2_X1 U4532 ( .A1(n4624), .A2(n4625), .ZN(n3752) );
  AND2_X1 U4533 ( .A1(n3724), .A2(n3723), .ZN(n4625) );
  AND2_X1 U4534 ( .A1(n3718), .A2(n4626), .ZN(n4624) );
  OR2_X1 U4535 ( .A1(n3724), .A2(n3723), .ZN(n4626) );
  OR2_X1 U4536 ( .A1(n4627), .A2(n4628), .ZN(n3723) );
  AND2_X1 U4537 ( .A1(n3697), .A2(n3699), .ZN(n4628) );
  AND2_X1 U4538 ( .A1(n3694), .A2(n4629), .ZN(n4627) );
  OR2_X1 U4539 ( .A1(n3697), .A2(n3699), .ZN(n4629) );
  OR2_X1 U4540 ( .A1(n4630), .A2(n4631), .ZN(n3699) );
  AND2_X1 U4541 ( .A1(n3673), .A2(n3671), .ZN(n4631) );
  AND2_X1 U4542 ( .A1(n4632), .A2(n4633), .ZN(n4630) );
  OR2_X1 U4543 ( .A1(n3673), .A2(n3671), .ZN(n4633) );
  OR2_X1 U4544 ( .A1(n3648), .A2(n4634), .ZN(n3671) );
  OR2_X1 U4545 ( .A1(n4070), .A2(n3645), .ZN(n4634) );
  INV_X1 U4546 ( .A(n3670), .ZN(n3673) );
  AND2_X1 U4547 ( .A1(a_13_), .A2(b_15_), .ZN(n3670) );
  INV_X1 U4548 ( .A(n3666), .ZN(n4632) );
  OR2_X1 U4549 ( .A1(n4635), .A2(n4636), .ZN(n3666) );
  AND2_X1 U4550 ( .A1(b_14_), .A2(n4637), .ZN(n4636) );
  OR2_X1 U4551 ( .A1(n4638), .A2(n3644), .ZN(n4637) );
  AND2_X1 U4552 ( .A1(a_14_), .A2(n3681), .ZN(n4638) );
  AND2_X1 U4553 ( .A1(b_13_), .A2(n4639), .ZN(n4635) );
  OR2_X1 U4554 ( .A1(n4640), .A2(n3647), .ZN(n4639) );
  AND2_X1 U4555 ( .A1(a_15_), .A2(n3645), .ZN(n4640) );
  OR2_X1 U4556 ( .A1(n4072), .A2(n3648), .ZN(n3697) );
  OR2_X1 U4557 ( .A1(n4641), .A2(n4642), .ZN(n3694) );
  AND2_X1 U4558 ( .A1(n4643), .A2(n4644), .ZN(n4642) );
  INV_X1 U4559 ( .A(n4645), .ZN(n4641) );
  OR2_X1 U4560 ( .A1(n4643), .A2(n4644), .ZN(n4645) );
  OR2_X1 U4561 ( .A1(n4646), .A2(n4647), .ZN(n4643) );
  AND2_X1 U4562 ( .A1(n4648), .A2(n4649), .ZN(n4647) );
  INV_X1 U4563 ( .A(n4650), .ZN(n4648) );
  AND2_X1 U4564 ( .A1(n4651), .A2(n4650), .ZN(n4646) );
  OR2_X1 U4565 ( .A1(n3735), .A2(n3648), .ZN(n3724) );
  OR2_X1 U4566 ( .A1(n4652), .A2(n4653), .ZN(n3718) );
  INV_X1 U4567 ( .A(n4654), .ZN(n4653) );
  OR2_X1 U4568 ( .A1(n4655), .A2(n4656), .ZN(n4654) );
  AND2_X1 U4569 ( .A1(n4656), .A2(n4655), .ZN(n4652) );
  AND2_X1 U4570 ( .A1(n4657), .A2(n4658), .ZN(n4655) );
  INV_X1 U4571 ( .A(n4659), .ZN(n4658) );
  AND2_X1 U4572 ( .A1(n4660), .A2(n4661), .ZN(n4659) );
  OR2_X1 U4573 ( .A1(n4661), .A2(n4660), .ZN(n4657) );
  INV_X1 U4574 ( .A(n4662), .ZN(n4660) );
  OR2_X1 U4575 ( .A1(n4059), .A2(n3648), .ZN(n3749) );
  OR2_X1 U4576 ( .A1(n4663), .A2(n4664), .ZN(n3746) );
  INV_X1 U4577 ( .A(n4665), .ZN(n4664) );
  OR2_X1 U4578 ( .A1(n4666), .A2(n4667), .ZN(n4665) );
  AND2_X1 U4579 ( .A1(n4667), .A2(n4666), .ZN(n4663) );
  AND2_X1 U4580 ( .A1(n4668), .A2(n4669), .ZN(n4666) );
  OR2_X1 U4581 ( .A1(n4670), .A2(n4671), .ZN(n4669) );
  INV_X1 U4582 ( .A(n4672), .ZN(n4671) );
  OR2_X1 U4583 ( .A1(n4672), .A2(n4673), .ZN(n4668) );
  INV_X1 U4584 ( .A(n4670), .ZN(n4673) );
  OR2_X1 U4585 ( .A1(n3786), .A2(n3648), .ZN(n3772) );
  OR2_X1 U4586 ( .A1(n4674), .A2(n4675), .ZN(n3769) );
  INV_X1 U4587 ( .A(n4676), .ZN(n4675) );
  OR2_X1 U4588 ( .A1(n4677), .A2(n4678), .ZN(n4676) );
  AND2_X1 U4589 ( .A1(n4678), .A2(n4677), .ZN(n4674) );
  AND2_X1 U4590 ( .A1(n4679), .A2(n4680), .ZN(n4677) );
  OR2_X1 U4591 ( .A1(n4681), .A2(n4682), .ZN(n4680) );
  INV_X1 U4592 ( .A(n4683), .ZN(n4679) );
  AND2_X1 U4593 ( .A1(n4682), .A2(n4681), .ZN(n4683) );
  INV_X1 U4594 ( .A(n4684), .ZN(n4682) );
  OR2_X1 U4595 ( .A1(n4053), .A2(n3648), .ZN(n3800) );
  OR2_X1 U4596 ( .A1(n4685), .A2(n4686), .ZN(n3797) );
  INV_X1 U4597 ( .A(n4687), .ZN(n4686) );
  OR2_X1 U4598 ( .A1(n4688), .A2(n4689), .ZN(n4687) );
  AND2_X1 U4599 ( .A1(n4689), .A2(n4688), .ZN(n4685) );
  AND2_X1 U4600 ( .A1(n4690), .A2(n4691), .ZN(n4688) );
  OR2_X1 U4601 ( .A1(n4692), .A2(n4693), .ZN(n4691) );
  INV_X1 U4602 ( .A(n4694), .ZN(n4693) );
  OR2_X1 U4603 ( .A1(n4694), .A2(n4695), .ZN(n4690) );
  INV_X1 U4604 ( .A(n4692), .ZN(n4695) );
  OR2_X1 U4605 ( .A1(n3837), .A2(n3648), .ZN(n3823) );
  OR2_X1 U4606 ( .A1(n4696), .A2(n4697), .ZN(n3820) );
  INV_X1 U4607 ( .A(n4698), .ZN(n4697) );
  OR2_X1 U4608 ( .A1(n4699), .A2(n4700), .ZN(n4698) );
  AND2_X1 U4609 ( .A1(n4700), .A2(n4699), .ZN(n4696) );
  AND2_X1 U4610 ( .A1(n4701), .A2(n4702), .ZN(n4699) );
  OR2_X1 U4611 ( .A1(n4703), .A2(n4704), .ZN(n4702) );
  INV_X1 U4612 ( .A(n4705), .ZN(n4704) );
  OR2_X1 U4613 ( .A1(n4705), .A2(n4706), .ZN(n4701) );
  INV_X1 U4614 ( .A(n4703), .ZN(n4706) );
  OR2_X1 U4615 ( .A1(n4047), .A2(n3648), .ZN(n3851) );
  OR2_X1 U4616 ( .A1(n4707), .A2(n4708), .ZN(n3848) );
  INV_X1 U4617 ( .A(n4709), .ZN(n4708) );
  OR2_X1 U4618 ( .A1(n4710), .A2(n4711), .ZN(n4709) );
  AND2_X1 U4619 ( .A1(n4711), .A2(n4710), .ZN(n4707) );
  AND2_X1 U4620 ( .A1(n4712), .A2(n4713), .ZN(n4710) );
  OR2_X1 U4621 ( .A1(n4714), .A2(n4715), .ZN(n4713) );
  INV_X1 U4622 ( .A(n4716), .ZN(n4715) );
  OR2_X1 U4623 ( .A1(n4716), .A2(n4717), .ZN(n4712) );
  INV_X1 U4624 ( .A(n4714), .ZN(n4717) );
  OR2_X1 U4625 ( .A1(n3888), .A2(n3648), .ZN(n3874) );
  OR2_X1 U4626 ( .A1(n4718), .A2(n4719), .ZN(n3871) );
  INV_X1 U4627 ( .A(n4720), .ZN(n4719) );
  OR2_X1 U4628 ( .A1(n4721), .A2(n4722), .ZN(n4720) );
  AND2_X1 U4629 ( .A1(n4722), .A2(n4721), .ZN(n4718) );
  AND2_X1 U4630 ( .A1(n4723), .A2(n4724), .ZN(n4721) );
  OR2_X1 U4631 ( .A1(n4725), .A2(n4726), .ZN(n4724) );
  INV_X1 U4632 ( .A(n4727), .ZN(n4726) );
  OR2_X1 U4633 ( .A1(n4727), .A2(n4728), .ZN(n4723) );
  INV_X1 U4634 ( .A(n4725), .ZN(n4728) );
  OR2_X1 U4635 ( .A1(n4041), .A2(n3648), .ZN(n3902) );
  OR2_X1 U4636 ( .A1(n4729), .A2(n4730), .ZN(n3899) );
  INV_X1 U4637 ( .A(n4731), .ZN(n4730) );
  OR2_X1 U4638 ( .A1(n4732), .A2(n4733), .ZN(n4731) );
  AND2_X1 U4639 ( .A1(n4733), .A2(n4732), .ZN(n4729) );
  AND2_X1 U4640 ( .A1(n4734), .A2(n4735), .ZN(n4732) );
  OR2_X1 U4641 ( .A1(n4736), .A2(n4737), .ZN(n4735) );
  INV_X1 U4642 ( .A(n4738), .ZN(n4737) );
  OR2_X1 U4643 ( .A1(n4738), .A2(n4739), .ZN(n4734) );
  INV_X1 U4644 ( .A(n4736), .ZN(n4739) );
  OR2_X1 U4645 ( .A1(n3951), .A2(n3648), .ZN(n3937) );
  OR2_X1 U4646 ( .A1(n4740), .A2(n4741), .ZN(n3934) );
  INV_X1 U4647 ( .A(n4742), .ZN(n4741) );
  OR2_X1 U4648 ( .A1(n4743), .A2(n4744), .ZN(n4742) );
  AND2_X1 U4649 ( .A1(n4744), .A2(n4743), .ZN(n4740) );
  AND2_X1 U4650 ( .A1(n4745), .A2(n4746), .ZN(n4743) );
  OR2_X1 U4651 ( .A1(n4747), .A2(n4748), .ZN(n4746) );
  INV_X1 U4652 ( .A(n4749), .ZN(n4748) );
  OR2_X1 U4653 ( .A1(n4749), .A2(n4750), .ZN(n4745) );
  INV_X1 U4654 ( .A(n4747), .ZN(n4750) );
  OR2_X1 U4655 ( .A1(n4035), .A2(n3648), .ZN(n3965) );
  OR2_X1 U4656 ( .A1(n4751), .A2(n4752), .ZN(n3962) );
  INV_X1 U4657 ( .A(n4753), .ZN(n4752) );
  OR2_X1 U4658 ( .A1(n4754), .A2(n4755), .ZN(n4753) );
  AND2_X1 U4659 ( .A1(n4755), .A2(n4754), .ZN(n4751) );
  AND2_X1 U4660 ( .A1(n4756), .A2(n4757), .ZN(n4754) );
  OR2_X1 U4661 ( .A1(n4758), .A2(n4759), .ZN(n4757) );
  INV_X1 U4662 ( .A(n4760), .ZN(n4759) );
  OR2_X1 U4663 ( .A1(n4760), .A2(n4761), .ZN(n4756) );
  INV_X1 U4664 ( .A(n4758), .ZN(n4761) );
  OR2_X1 U4665 ( .A1(n4002), .A2(n3648), .ZN(n3988) );
  INV_X1 U4666 ( .A(b_15_), .ZN(n3648) );
  OR2_X1 U4667 ( .A1(n4762), .A2(n4763), .ZN(n3985) );
  INV_X1 U4668 ( .A(n4764), .ZN(n4763) );
  OR2_X1 U4669 ( .A1(n4765), .A2(n4766), .ZN(n4764) );
  AND2_X1 U4670 ( .A1(n4766), .A2(n4765), .ZN(n4762) );
  AND2_X1 U4671 ( .A1(n4767), .A2(n4768), .ZN(n4765) );
  OR2_X1 U4672 ( .A1(n4769), .A2(n4770), .ZN(n4768) );
  INV_X1 U4673 ( .A(n4771), .ZN(n4770) );
  OR2_X1 U4674 ( .A1(n4771), .A2(n4772), .ZN(n4767) );
  INV_X1 U4675 ( .A(n4769), .ZN(n4772) );
  INV_X1 U4676 ( .A(n4019), .ZN(n4016) );
  AND2_X1 U4677 ( .A1(a_0_), .A2(b_15_), .ZN(n4019) );
  OR2_X1 U4678 ( .A1(n4773), .A2(n4774), .ZN(n4013) );
  INV_X1 U4679 ( .A(n4775), .ZN(n4774) );
  OR2_X1 U4680 ( .A1(n4776), .A2(n4539), .ZN(n4775) );
  AND2_X1 U4681 ( .A1(n4539), .A2(n4776), .ZN(n4773) );
  AND2_X1 U4682 ( .A1(n4777), .A2(n4778), .ZN(n4776) );
  OR2_X1 U4683 ( .A1(n4537), .A2(n4779), .ZN(n4778) );
  INV_X1 U4684 ( .A(n4538), .ZN(n4779) );
  OR2_X1 U4685 ( .A1(n4538), .A2(n4780), .ZN(n4777) );
  INV_X1 U4686 ( .A(n4537), .ZN(n4780) );
  OR2_X1 U4687 ( .A1(n4002), .A2(n3645), .ZN(n4537) );
  OR2_X1 U4688 ( .A1(n4781), .A2(n4782), .ZN(n4538) );
  AND2_X1 U4689 ( .A1(n4769), .A2(n4771), .ZN(n4782) );
  AND2_X1 U4690 ( .A1(n4766), .A2(n4783), .ZN(n4781) );
  OR2_X1 U4691 ( .A1(n4771), .A2(n4769), .ZN(n4783) );
  OR2_X1 U4692 ( .A1(n4035), .A2(n3645), .ZN(n4769) );
  OR2_X1 U4693 ( .A1(n4784), .A2(n4785), .ZN(n4771) );
  AND2_X1 U4694 ( .A1(n4758), .A2(n4760), .ZN(n4785) );
  AND2_X1 U4695 ( .A1(n4755), .A2(n4786), .ZN(n4784) );
  OR2_X1 U4696 ( .A1(n4760), .A2(n4758), .ZN(n4786) );
  OR2_X1 U4697 ( .A1(n3951), .A2(n3645), .ZN(n4758) );
  OR2_X1 U4698 ( .A1(n4787), .A2(n4788), .ZN(n4760) );
  AND2_X1 U4699 ( .A1(n4747), .A2(n4749), .ZN(n4788) );
  AND2_X1 U4700 ( .A1(n4744), .A2(n4789), .ZN(n4787) );
  OR2_X1 U4701 ( .A1(n4749), .A2(n4747), .ZN(n4789) );
  OR2_X1 U4702 ( .A1(n4041), .A2(n3645), .ZN(n4747) );
  OR2_X1 U4703 ( .A1(n4790), .A2(n4791), .ZN(n4749) );
  AND2_X1 U4704 ( .A1(n4736), .A2(n4738), .ZN(n4791) );
  AND2_X1 U4705 ( .A1(n4733), .A2(n4792), .ZN(n4790) );
  OR2_X1 U4706 ( .A1(n4738), .A2(n4736), .ZN(n4792) );
  OR2_X1 U4707 ( .A1(n3888), .A2(n3645), .ZN(n4736) );
  OR2_X1 U4708 ( .A1(n4793), .A2(n4794), .ZN(n4738) );
  AND2_X1 U4709 ( .A1(n4725), .A2(n4727), .ZN(n4794) );
  AND2_X1 U4710 ( .A1(n4722), .A2(n4795), .ZN(n4793) );
  OR2_X1 U4711 ( .A1(n4727), .A2(n4725), .ZN(n4795) );
  OR2_X1 U4712 ( .A1(n4047), .A2(n3645), .ZN(n4725) );
  OR2_X1 U4713 ( .A1(n4796), .A2(n4797), .ZN(n4727) );
  AND2_X1 U4714 ( .A1(n4714), .A2(n4716), .ZN(n4797) );
  AND2_X1 U4715 ( .A1(n4711), .A2(n4798), .ZN(n4796) );
  OR2_X1 U4716 ( .A1(n4716), .A2(n4714), .ZN(n4798) );
  OR2_X1 U4717 ( .A1(n3837), .A2(n3645), .ZN(n4714) );
  OR2_X1 U4718 ( .A1(n4799), .A2(n4800), .ZN(n4716) );
  AND2_X1 U4719 ( .A1(n4703), .A2(n4705), .ZN(n4800) );
  AND2_X1 U4720 ( .A1(n4700), .A2(n4801), .ZN(n4799) );
  OR2_X1 U4721 ( .A1(n4705), .A2(n4703), .ZN(n4801) );
  OR2_X1 U4722 ( .A1(n4053), .A2(n3645), .ZN(n4703) );
  OR2_X1 U4723 ( .A1(n4802), .A2(n4803), .ZN(n4705) );
  AND2_X1 U4724 ( .A1(n4692), .A2(n4694), .ZN(n4803) );
  AND2_X1 U4725 ( .A1(n4689), .A2(n4804), .ZN(n4802) );
  OR2_X1 U4726 ( .A1(n4694), .A2(n4692), .ZN(n4804) );
  OR2_X1 U4727 ( .A1(n3786), .A2(n3645), .ZN(n4692) );
  OR2_X1 U4728 ( .A1(n4805), .A2(n4806), .ZN(n4694) );
  AND2_X1 U4729 ( .A1(n4681), .A2(n4684), .ZN(n4806) );
  AND2_X1 U4730 ( .A1(n4678), .A2(n4807), .ZN(n4805) );
  OR2_X1 U4731 ( .A1(n4684), .A2(n4681), .ZN(n4807) );
  OR2_X1 U4732 ( .A1(n4059), .A2(n3645), .ZN(n4681) );
  OR2_X1 U4733 ( .A1(n4808), .A2(n4809), .ZN(n4684) );
  AND2_X1 U4734 ( .A1(n4670), .A2(n4672), .ZN(n4809) );
  AND2_X1 U4735 ( .A1(n4667), .A2(n4810), .ZN(n4808) );
  OR2_X1 U4736 ( .A1(n4672), .A2(n4670), .ZN(n4810) );
  OR2_X1 U4737 ( .A1(n3735), .A2(n3645), .ZN(n4670) );
  OR2_X1 U4738 ( .A1(n4811), .A2(n4812), .ZN(n4672) );
  AND2_X1 U4739 ( .A1(n4662), .A2(n4661), .ZN(n4812) );
  AND2_X1 U4740 ( .A1(n4656), .A2(n4813), .ZN(n4811) );
  OR2_X1 U4741 ( .A1(n4661), .A2(n4662), .ZN(n4813) );
  OR2_X1 U4742 ( .A1(n4072), .A2(n3645), .ZN(n4662) );
  OR2_X1 U4743 ( .A1(n4814), .A2(n4815), .ZN(n4661) );
  AND2_X1 U4744 ( .A1(n4644), .A2(n4650), .ZN(n4815) );
  AND2_X1 U4745 ( .A1(n4651), .A2(n4816), .ZN(n4814) );
  OR2_X1 U4746 ( .A1(n4650), .A2(n4644), .ZN(n4816) );
  OR2_X1 U4747 ( .A1(n3682), .A2(n3645), .ZN(n4644) );
  OR2_X1 U4748 ( .A1(n3645), .A2(n4817), .ZN(n4650) );
  INV_X1 U4749 ( .A(b_14_), .ZN(n3645) );
  INV_X1 U4750 ( .A(n4649), .ZN(n4651) );
  OR2_X1 U4751 ( .A1(n4818), .A2(n4819), .ZN(n4649) );
  AND2_X1 U4752 ( .A1(b_13_), .A2(n4820), .ZN(n4819) );
  OR2_X1 U4753 ( .A1(n4821), .A2(n3644), .ZN(n4820) );
  AND2_X1 U4754 ( .A1(a_14_), .A2(n4073), .ZN(n4821) );
  AND2_X1 U4755 ( .A1(b_12_), .A2(n4822), .ZN(n4818) );
  OR2_X1 U4756 ( .A1(n4823), .A2(n3647), .ZN(n4822) );
  AND2_X1 U4757 ( .A1(a_15_), .A2(n3681), .ZN(n4823) );
  OR2_X1 U4758 ( .A1(n4824), .A2(n4825), .ZN(n4656) );
  AND2_X1 U4759 ( .A1(n4826), .A2(n4067), .ZN(n4825) );
  AND2_X1 U4760 ( .A1(n4827), .A2(n3685), .ZN(n4824) );
  INV_X1 U4761 ( .A(n4067), .ZN(n3685) );
  INV_X1 U4762 ( .A(n4826), .ZN(n4827) );
  OR2_X1 U4763 ( .A1(n4828), .A2(n4829), .ZN(n4826) );
  AND2_X1 U4764 ( .A1(n4830), .A2(n4831), .ZN(n4829) );
  INV_X1 U4765 ( .A(n4832), .ZN(n4830) );
  AND2_X1 U4766 ( .A1(n4833), .A2(n4832), .ZN(n4828) );
  OR2_X1 U4767 ( .A1(n4834), .A2(n4835), .ZN(n4667) );
  INV_X1 U4768 ( .A(n4836), .ZN(n4835) );
  OR2_X1 U4769 ( .A1(n4837), .A2(n4838), .ZN(n4836) );
  AND2_X1 U4770 ( .A1(n4838), .A2(n4837), .ZN(n4834) );
  AND2_X1 U4771 ( .A1(n4839), .A2(n4840), .ZN(n4837) );
  OR2_X1 U4772 ( .A1(n4841), .A2(n4842), .ZN(n4840) );
  INV_X1 U4773 ( .A(n4843), .ZN(n4842) );
  OR2_X1 U4774 ( .A1(n4843), .A2(n4844), .ZN(n4839) );
  INV_X1 U4775 ( .A(n4841), .ZN(n4844) );
  OR2_X1 U4776 ( .A1(n4845), .A2(n4846), .ZN(n4678) );
  INV_X1 U4777 ( .A(n4847), .ZN(n4846) );
  OR2_X1 U4778 ( .A1(n4848), .A2(n4849), .ZN(n4847) );
  AND2_X1 U4779 ( .A1(n4849), .A2(n4848), .ZN(n4845) );
  AND2_X1 U4780 ( .A1(n4850), .A2(n4851), .ZN(n4848) );
  OR2_X1 U4781 ( .A1(n4852), .A2(n4853), .ZN(n4851) );
  INV_X1 U4782 ( .A(n4854), .ZN(n4853) );
  OR2_X1 U4783 ( .A1(n4854), .A2(n4855), .ZN(n4850) );
  INV_X1 U4784 ( .A(n4852), .ZN(n4855) );
  OR2_X1 U4785 ( .A1(n4856), .A2(n4857), .ZN(n4689) );
  INV_X1 U4786 ( .A(n4858), .ZN(n4857) );
  OR2_X1 U4787 ( .A1(n4859), .A2(n4860), .ZN(n4858) );
  AND2_X1 U4788 ( .A1(n4860), .A2(n4859), .ZN(n4856) );
  AND2_X1 U4789 ( .A1(n4861), .A2(n4862), .ZN(n4859) );
  OR2_X1 U4790 ( .A1(n4863), .A2(n4864), .ZN(n4862) );
  INV_X1 U4791 ( .A(n4865), .ZN(n4861) );
  AND2_X1 U4792 ( .A1(n4864), .A2(n4863), .ZN(n4865) );
  INV_X1 U4793 ( .A(n4866), .ZN(n4864) );
  OR2_X1 U4794 ( .A1(n4867), .A2(n4868), .ZN(n4700) );
  INV_X1 U4795 ( .A(n4869), .ZN(n4868) );
  OR2_X1 U4796 ( .A1(n4870), .A2(n4871), .ZN(n4869) );
  AND2_X1 U4797 ( .A1(n4871), .A2(n4870), .ZN(n4867) );
  AND2_X1 U4798 ( .A1(n4872), .A2(n4873), .ZN(n4870) );
  OR2_X1 U4799 ( .A1(n4874), .A2(n4875), .ZN(n4873) );
  INV_X1 U4800 ( .A(n4876), .ZN(n4875) );
  OR2_X1 U4801 ( .A1(n4876), .A2(n4877), .ZN(n4872) );
  INV_X1 U4802 ( .A(n4874), .ZN(n4877) );
  OR2_X1 U4803 ( .A1(n4878), .A2(n4879), .ZN(n4711) );
  INV_X1 U4804 ( .A(n4880), .ZN(n4879) );
  OR2_X1 U4805 ( .A1(n4881), .A2(n4882), .ZN(n4880) );
  AND2_X1 U4806 ( .A1(n4882), .A2(n4881), .ZN(n4878) );
  AND2_X1 U4807 ( .A1(n4883), .A2(n4884), .ZN(n4881) );
  OR2_X1 U4808 ( .A1(n4885), .A2(n4886), .ZN(n4884) );
  INV_X1 U4809 ( .A(n4887), .ZN(n4886) );
  OR2_X1 U4810 ( .A1(n4887), .A2(n4888), .ZN(n4883) );
  INV_X1 U4811 ( .A(n4885), .ZN(n4888) );
  OR2_X1 U4812 ( .A1(n4889), .A2(n4890), .ZN(n4722) );
  INV_X1 U4813 ( .A(n4891), .ZN(n4890) );
  OR2_X1 U4814 ( .A1(n4892), .A2(n4893), .ZN(n4891) );
  AND2_X1 U4815 ( .A1(n4893), .A2(n4892), .ZN(n4889) );
  AND2_X1 U4816 ( .A1(n4894), .A2(n4895), .ZN(n4892) );
  OR2_X1 U4817 ( .A1(n4896), .A2(n4897), .ZN(n4895) );
  INV_X1 U4818 ( .A(n4898), .ZN(n4897) );
  OR2_X1 U4819 ( .A1(n4898), .A2(n4899), .ZN(n4894) );
  INV_X1 U4820 ( .A(n4896), .ZN(n4899) );
  OR2_X1 U4821 ( .A1(n4900), .A2(n4901), .ZN(n4733) );
  INV_X1 U4822 ( .A(n4902), .ZN(n4901) );
  OR2_X1 U4823 ( .A1(n4903), .A2(n4904), .ZN(n4902) );
  AND2_X1 U4824 ( .A1(n4904), .A2(n4903), .ZN(n4900) );
  AND2_X1 U4825 ( .A1(n4905), .A2(n4906), .ZN(n4903) );
  OR2_X1 U4826 ( .A1(n4907), .A2(n4908), .ZN(n4906) );
  INV_X1 U4827 ( .A(n4909), .ZN(n4908) );
  OR2_X1 U4828 ( .A1(n4909), .A2(n4910), .ZN(n4905) );
  INV_X1 U4829 ( .A(n4907), .ZN(n4910) );
  OR2_X1 U4830 ( .A1(n4911), .A2(n4912), .ZN(n4744) );
  INV_X1 U4831 ( .A(n4913), .ZN(n4912) );
  OR2_X1 U4832 ( .A1(n4914), .A2(n4915), .ZN(n4913) );
  AND2_X1 U4833 ( .A1(n4915), .A2(n4914), .ZN(n4911) );
  AND2_X1 U4834 ( .A1(n4916), .A2(n4917), .ZN(n4914) );
  OR2_X1 U4835 ( .A1(n4918), .A2(n4919), .ZN(n4917) );
  INV_X1 U4836 ( .A(n4920), .ZN(n4919) );
  OR2_X1 U4837 ( .A1(n4920), .A2(n4921), .ZN(n4916) );
  INV_X1 U4838 ( .A(n4918), .ZN(n4921) );
  OR2_X1 U4839 ( .A1(n4922), .A2(n4923), .ZN(n4755) );
  INV_X1 U4840 ( .A(n4924), .ZN(n4923) );
  OR2_X1 U4841 ( .A1(n4925), .A2(n4926), .ZN(n4924) );
  AND2_X1 U4842 ( .A1(n4926), .A2(n4925), .ZN(n4922) );
  AND2_X1 U4843 ( .A1(n4927), .A2(n4928), .ZN(n4925) );
  OR2_X1 U4844 ( .A1(n4929), .A2(n4930), .ZN(n4928) );
  INV_X1 U4845 ( .A(n4931), .ZN(n4930) );
  OR2_X1 U4846 ( .A1(n4931), .A2(n4932), .ZN(n4927) );
  INV_X1 U4847 ( .A(n4929), .ZN(n4932) );
  OR2_X1 U4848 ( .A1(n4933), .A2(n4934), .ZN(n4766) );
  INV_X1 U4849 ( .A(n4935), .ZN(n4934) );
  OR2_X1 U4850 ( .A1(n4936), .A2(n4937), .ZN(n4935) );
  AND2_X1 U4851 ( .A1(n4937), .A2(n4936), .ZN(n4933) );
  AND2_X1 U4852 ( .A1(n4938), .A2(n4939), .ZN(n4936) );
  OR2_X1 U4853 ( .A1(n4940), .A2(n4941), .ZN(n4939) );
  INV_X1 U4854 ( .A(n4942), .ZN(n4941) );
  OR2_X1 U4855 ( .A1(n4942), .A2(n4943), .ZN(n4938) );
  INV_X1 U4856 ( .A(n4940), .ZN(n4943) );
  OR2_X1 U4857 ( .A1(n4944), .A2(n4945), .ZN(n4539) );
  INV_X1 U4858 ( .A(n4946), .ZN(n4945) );
  OR2_X1 U4859 ( .A1(n4947), .A2(n4567), .ZN(n4946) );
  AND2_X1 U4860 ( .A1(n4567), .A2(n4947), .ZN(n4944) );
  AND2_X1 U4861 ( .A1(n4948), .A2(n4949), .ZN(n4947) );
  OR2_X1 U4862 ( .A1(n4565), .A2(n4950), .ZN(n4949) );
  INV_X1 U4863 ( .A(n4566), .ZN(n4950) );
  OR2_X1 U4864 ( .A1(n4566), .A2(n4951), .ZN(n4948) );
  INV_X1 U4865 ( .A(n4565), .ZN(n4951) );
  OR2_X1 U4866 ( .A1(n4035), .A2(n3681), .ZN(n4565) );
  OR2_X1 U4867 ( .A1(n4952), .A2(n4953), .ZN(n4566) );
  AND2_X1 U4868 ( .A1(n4940), .A2(n4942), .ZN(n4953) );
  AND2_X1 U4869 ( .A1(n4937), .A2(n4954), .ZN(n4952) );
  OR2_X1 U4870 ( .A1(n4942), .A2(n4940), .ZN(n4954) );
  OR2_X1 U4871 ( .A1(n3951), .A2(n3681), .ZN(n4940) );
  OR2_X1 U4872 ( .A1(n4955), .A2(n4956), .ZN(n4942) );
  AND2_X1 U4873 ( .A1(n4929), .A2(n4931), .ZN(n4956) );
  AND2_X1 U4874 ( .A1(n4926), .A2(n4957), .ZN(n4955) );
  OR2_X1 U4875 ( .A1(n4931), .A2(n4929), .ZN(n4957) );
  OR2_X1 U4876 ( .A1(n4041), .A2(n3681), .ZN(n4929) );
  OR2_X1 U4877 ( .A1(n4958), .A2(n4959), .ZN(n4931) );
  AND2_X1 U4878 ( .A1(n4918), .A2(n4920), .ZN(n4959) );
  AND2_X1 U4879 ( .A1(n4915), .A2(n4960), .ZN(n4958) );
  OR2_X1 U4880 ( .A1(n4920), .A2(n4918), .ZN(n4960) );
  OR2_X1 U4881 ( .A1(n3888), .A2(n3681), .ZN(n4918) );
  OR2_X1 U4882 ( .A1(n4961), .A2(n4962), .ZN(n4920) );
  AND2_X1 U4883 ( .A1(n4907), .A2(n4909), .ZN(n4962) );
  AND2_X1 U4884 ( .A1(n4904), .A2(n4963), .ZN(n4961) );
  OR2_X1 U4885 ( .A1(n4909), .A2(n4907), .ZN(n4963) );
  OR2_X1 U4886 ( .A1(n4047), .A2(n3681), .ZN(n4907) );
  OR2_X1 U4887 ( .A1(n4964), .A2(n4965), .ZN(n4909) );
  AND2_X1 U4888 ( .A1(n4896), .A2(n4898), .ZN(n4965) );
  AND2_X1 U4889 ( .A1(n4893), .A2(n4966), .ZN(n4964) );
  OR2_X1 U4890 ( .A1(n4898), .A2(n4896), .ZN(n4966) );
  OR2_X1 U4891 ( .A1(n3837), .A2(n3681), .ZN(n4896) );
  OR2_X1 U4892 ( .A1(n4967), .A2(n4968), .ZN(n4898) );
  AND2_X1 U4893 ( .A1(n4885), .A2(n4887), .ZN(n4968) );
  AND2_X1 U4894 ( .A1(n4882), .A2(n4969), .ZN(n4967) );
  OR2_X1 U4895 ( .A1(n4887), .A2(n4885), .ZN(n4969) );
  OR2_X1 U4896 ( .A1(n4053), .A2(n3681), .ZN(n4885) );
  OR2_X1 U4897 ( .A1(n4970), .A2(n4971), .ZN(n4887) );
  AND2_X1 U4898 ( .A1(n4874), .A2(n4876), .ZN(n4971) );
  AND2_X1 U4899 ( .A1(n4871), .A2(n4972), .ZN(n4970) );
  OR2_X1 U4900 ( .A1(n4876), .A2(n4874), .ZN(n4972) );
  OR2_X1 U4901 ( .A1(n3786), .A2(n3681), .ZN(n4874) );
  OR2_X1 U4902 ( .A1(n4973), .A2(n4974), .ZN(n4876) );
  AND2_X1 U4903 ( .A1(n4863), .A2(n4866), .ZN(n4974) );
  AND2_X1 U4904 ( .A1(n4860), .A2(n4975), .ZN(n4973) );
  OR2_X1 U4905 ( .A1(n4866), .A2(n4863), .ZN(n4975) );
  OR2_X1 U4906 ( .A1(n4059), .A2(n3681), .ZN(n4863) );
  OR2_X1 U4907 ( .A1(n4976), .A2(n4977), .ZN(n4866) );
  AND2_X1 U4908 ( .A1(n4852), .A2(n4854), .ZN(n4977) );
  AND2_X1 U4909 ( .A1(n4849), .A2(n4978), .ZN(n4976) );
  OR2_X1 U4910 ( .A1(n4854), .A2(n4852), .ZN(n4978) );
  OR2_X1 U4911 ( .A1(n3735), .A2(n3681), .ZN(n4852) );
  OR2_X1 U4912 ( .A1(n4979), .A2(n4980), .ZN(n4854) );
  AND2_X1 U4913 ( .A1(n4841), .A2(n4843), .ZN(n4980) );
  AND2_X1 U4914 ( .A1(n4838), .A2(n4981), .ZN(n4979) );
  OR2_X1 U4915 ( .A1(n4843), .A2(n4841), .ZN(n4981) );
  OR2_X1 U4916 ( .A1(n4072), .A2(n3681), .ZN(n4841) );
  OR2_X1 U4917 ( .A1(n4982), .A2(n4983), .ZN(n4843) );
  AND2_X1 U4918 ( .A1(n4067), .A2(n4832), .ZN(n4983) );
  AND2_X1 U4919 ( .A1(n4833), .A2(n4984), .ZN(n4982) );
  OR2_X1 U4920 ( .A1(n4832), .A2(n4067), .ZN(n4984) );
  OR2_X1 U4921 ( .A1(n3682), .A2(n3681), .ZN(n4067) );
  OR2_X1 U4922 ( .A1(n4073), .A2(n4817), .ZN(n4832) );
  OR2_X1 U4923 ( .A1(n4070), .A2(n3681), .ZN(n4817) );
  INV_X1 U4924 ( .A(b_13_), .ZN(n3681) );
  INV_X1 U4925 ( .A(n4831), .ZN(n4833) );
  OR2_X1 U4926 ( .A1(n4985), .A2(n4986), .ZN(n4831) );
  AND2_X1 U4927 ( .A1(b_12_), .A2(n4987), .ZN(n4986) );
  OR2_X1 U4928 ( .A1(n4988), .A2(n3644), .ZN(n4987) );
  AND2_X1 U4929 ( .A1(a_14_), .A2(n3731), .ZN(n4988) );
  AND2_X1 U4930 ( .A1(b_11_), .A2(n4989), .ZN(n4985) );
  OR2_X1 U4931 ( .A1(n4990), .A2(n3647), .ZN(n4989) );
  AND2_X1 U4932 ( .A1(a_15_), .A2(n4073), .ZN(n4990) );
  OR2_X1 U4933 ( .A1(n4991), .A2(n4992), .ZN(n4838) );
  AND2_X1 U4934 ( .A1(n4993), .A2(n4994), .ZN(n4992) );
  INV_X1 U4935 ( .A(n4995), .ZN(n4991) );
  OR2_X1 U4936 ( .A1(n4993), .A2(n4994), .ZN(n4995) );
  OR2_X1 U4937 ( .A1(n4996), .A2(n4997), .ZN(n4993) );
  AND2_X1 U4938 ( .A1(n4998), .A2(n4999), .ZN(n4997) );
  INV_X1 U4939 ( .A(n5000), .ZN(n4998) );
  AND2_X1 U4940 ( .A1(n5001), .A2(n5000), .ZN(n4996) );
  OR2_X1 U4941 ( .A1(n5002), .A2(n5003), .ZN(n4849) );
  INV_X1 U4942 ( .A(n5004), .ZN(n5003) );
  OR2_X1 U4943 ( .A1(n5005), .A2(n5006), .ZN(n5004) );
  AND2_X1 U4944 ( .A1(n5006), .A2(n5005), .ZN(n5002) );
  AND2_X1 U4945 ( .A1(n5007), .A2(n5008), .ZN(n5005) );
  OR2_X1 U4946 ( .A1(n4065), .A2(n5009), .ZN(n5008) );
  INV_X1 U4947 ( .A(n5010), .ZN(n5009) );
  OR2_X1 U4948 ( .A1(n5010), .A2(n3709), .ZN(n5007) );
  INV_X1 U4949 ( .A(n4065), .ZN(n3709) );
  OR2_X1 U4950 ( .A1(n5011), .A2(n5012), .ZN(n4860) );
  INV_X1 U4951 ( .A(n5013), .ZN(n5012) );
  OR2_X1 U4952 ( .A1(n5014), .A2(n5015), .ZN(n5013) );
  AND2_X1 U4953 ( .A1(n5015), .A2(n5014), .ZN(n5011) );
  AND2_X1 U4954 ( .A1(n5016), .A2(n5017), .ZN(n5014) );
  OR2_X1 U4955 ( .A1(n5018), .A2(n5019), .ZN(n5017) );
  INV_X1 U4956 ( .A(n5020), .ZN(n5019) );
  OR2_X1 U4957 ( .A1(n5020), .A2(n5021), .ZN(n5016) );
  INV_X1 U4958 ( .A(n5018), .ZN(n5021) );
  OR2_X1 U4959 ( .A1(n5022), .A2(n5023), .ZN(n4871) );
  INV_X1 U4960 ( .A(n5024), .ZN(n5023) );
  OR2_X1 U4961 ( .A1(n5025), .A2(n5026), .ZN(n5024) );
  AND2_X1 U4962 ( .A1(n5026), .A2(n5025), .ZN(n5022) );
  AND2_X1 U4963 ( .A1(n5027), .A2(n5028), .ZN(n5025) );
  OR2_X1 U4964 ( .A1(n5029), .A2(n5030), .ZN(n5028) );
  INV_X1 U4965 ( .A(n5031), .ZN(n5027) );
  AND2_X1 U4966 ( .A1(n5030), .A2(n5029), .ZN(n5031) );
  INV_X1 U4967 ( .A(n5032), .ZN(n5030) );
  OR2_X1 U4968 ( .A1(n5033), .A2(n5034), .ZN(n4882) );
  INV_X1 U4969 ( .A(n5035), .ZN(n5034) );
  OR2_X1 U4970 ( .A1(n5036), .A2(n5037), .ZN(n5035) );
  AND2_X1 U4971 ( .A1(n5037), .A2(n5036), .ZN(n5033) );
  AND2_X1 U4972 ( .A1(n5038), .A2(n5039), .ZN(n5036) );
  OR2_X1 U4973 ( .A1(n5040), .A2(n5041), .ZN(n5039) );
  INV_X1 U4974 ( .A(n5042), .ZN(n5041) );
  OR2_X1 U4975 ( .A1(n5042), .A2(n5043), .ZN(n5038) );
  INV_X1 U4976 ( .A(n5040), .ZN(n5043) );
  OR2_X1 U4977 ( .A1(n5044), .A2(n5045), .ZN(n4893) );
  INV_X1 U4978 ( .A(n5046), .ZN(n5045) );
  OR2_X1 U4979 ( .A1(n5047), .A2(n5048), .ZN(n5046) );
  AND2_X1 U4980 ( .A1(n5048), .A2(n5047), .ZN(n5044) );
  AND2_X1 U4981 ( .A1(n5049), .A2(n5050), .ZN(n5047) );
  OR2_X1 U4982 ( .A1(n5051), .A2(n5052), .ZN(n5050) );
  INV_X1 U4983 ( .A(n5053), .ZN(n5052) );
  OR2_X1 U4984 ( .A1(n5053), .A2(n5054), .ZN(n5049) );
  INV_X1 U4985 ( .A(n5051), .ZN(n5054) );
  OR2_X1 U4986 ( .A1(n5055), .A2(n5056), .ZN(n4904) );
  INV_X1 U4987 ( .A(n5057), .ZN(n5056) );
  OR2_X1 U4988 ( .A1(n5058), .A2(n5059), .ZN(n5057) );
  AND2_X1 U4989 ( .A1(n5059), .A2(n5058), .ZN(n5055) );
  AND2_X1 U4990 ( .A1(n5060), .A2(n5061), .ZN(n5058) );
  OR2_X1 U4991 ( .A1(n5062), .A2(n5063), .ZN(n5061) );
  INV_X1 U4992 ( .A(n5064), .ZN(n5063) );
  OR2_X1 U4993 ( .A1(n5064), .A2(n5065), .ZN(n5060) );
  INV_X1 U4994 ( .A(n5062), .ZN(n5065) );
  OR2_X1 U4995 ( .A1(n5066), .A2(n5067), .ZN(n4915) );
  INV_X1 U4996 ( .A(n5068), .ZN(n5067) );
  OR2_X1 U4997 ( .A1(n5069), .A2(n5070), .ZN(n5068) );
  AND2_X1 U4998 ( .A1(n5070), .A2(n5069), .ZN(n5066) );
  AND2_X1 U4999 ( .A1(n5071), .A2(n5072), .ZN(n5069) );
  OR2_X1 U5000 ( .A1(n5073), .A2(n5074), .ZN(n5072) );
  INV_X1 U5001 ( .A(n5075), .ZN(n5074) );
  OR2_X1 U5002 ( .A1(n5075), .A2(n5076), .ZN(n5071) );
  INV_X1 U5003 ( .A(n5073), .ZN(n5076) );
  OR2_X1 U5004 ( .A1(n5077), .A2(n5078), .ZN(n4926) );
  INV_X1 U5005 ( .A(n5079), .ZN(n5078) );
  OR2_X1 U5006 ( .A1(n5080), .A2(n5081), .ZN(n5079) );
  AND2_X1 U5007 ( .A1(n5081), .A2(n5080), .ZN(n5077) );
  AND2_X1 U5008 ( .A1(n5082), .A2(n5083), .ZN(n5080) );
  OR2_X1 U5009 ( .A1(n5084), .A2(n5085), .ZN(n5083) );
  INV_X1 U5010 ( .A(n5086), .ZN(n5085) );
  OR2_X1 U5011 ( .A1(n5086), .A2(n5087), .ZN(n5082) );
  INV_X1 U5012 ( .A(n5084), .ZN(n5087) );
  OR2_X1 U5013 ( .A1(n5088), .A2(n5089), .ZN(n4937) );
  INV_X1 U5014 ( .A(n5090), .ZN(n5089) );
  OR2_X1 U5015 ( .A1(n5091), .A2(n5092), .ZN(n5090) );
  AND2_X1 U5016 ( .A1(n5092), .A2(n5091), .ZN(n5088) );
  AND2_X1 U5017 ( .A1(n5093), .A2(n5094), .ZN(n5091) );
  OR2_X1 U5018 ( .A1(n5095), .A2(n5096), .ZN(n5094) );
  INV_X1 U5019 ( .A(n5097), .ZN(n5096) );
  OR2_X1 U5020 ( .A1(n5097), .A2(n5098), .ZN(n5093) );
  INV_X1 U5021 ( .A(n5095), .ZN(n5098) );
  OR2_X1 U5022 ( .A1(n5099), .A2(n5100), .ZN(n4567) );
  INV_X1 U5023 ( .A(n5101), .ZN(n5100) );
  OR2_X1 U5024 ( .A1(n5102), .A2(n5103), .ZN(n5101) );
  AND2_X1 U5025 ( .A1(n5103), .A2(n5102), .ZN(n5099) );
  AND2_X1 U5026 ( .A1(n5104), .A2(n5105), .ZN(n5102) );
  OR2_X1 U5027 ( .A1(n5106), .A2(n5107), .ZN(n5105) );
  INV_X1 U5028 ( .A(n5108), .ZN(n5107) );
  OR2_X1 U5029 ( .A1(n5108), .A2(n5109), .ZN(n5104) );
  INV_X1 U5030 ( .A(n5106), .ZN(n5109) );
  AND2_X1 U5031 ( .A1(n5110), .A2(n4112), .ZN(n4108) );
  OR2_X1 U5032 ( .A1(n5111), .A2(n5112), .ZN(n4112) );
  INV_X1 U5033 ( .A(n5113), .ZN(n5110) );
  AND2_X1 U5034 ( .A1(n5111), .A2(n5112), .ZN(n5113) );
  OR2_X1 U5035 ( .A1(n5114), .A2(n5115), .ZN(n5112) );
  AND2_X1 U5036 ( .A1(n5116), .A2(n4514), .ZN(n5115) );
  AND2_X1 U5037 ( .A1(n4510), .A2(n5117), .ZN(n5114) );
  OR2_X1 U5038 ( .A1(n4514), .A2(n5116), .ZN(n5117) );
  INV_X1 U5039 ( .A(n4513), .ZN(n5116) );
  AND2_X1 U5040 ( .A1(a_0_), .A2(b_12_), .ZN(n4513) );
  OR2_X1 U5041 ( .A1(n5118), .A2(n5119), .ZN(n4514) );
  AND2_X1 U5042 ( .A1(n4587), .A2(n4589), .ZN(n5119) );
  AND2_X1 U5043 ( .A1(n4584), .A2(n5120), .ZN(n5118) );
  OR2_X1 U5044 ( .A1(n4589), .A2(n4587), .ZN(n5120) );
  OR2_X1 U5045 ( .A1(n4002), .A2(n4073), .ZN(n4587) );
  OR2_X1 U5046 ( .A1(n5121), .A2(n5122), .ZN(n4589) );
  AND2_X1 U5047 ( .A1(n4578), .A2(n4577), .ZN(n5122) );
  AND2_X1 U5048 ( .A1(n4573), .A2(n5123), .ZN(n5121) );
  OR2_X1 U5049 ( .A1(n4577), .A2(n4578), .ZN(n5123) );
  OR2_X1 U5050 ( .A1(n4035), .A2(n4073), .ZN(n4578) );
  OR2_X1 U5051 ( .A1(n5124), .A2(n5125), .ZN(n4577) );
  AND2_X1 U5052 ( .A1(n5106), .A2(n5108), .ZN(n5125) );
  AND2_X1 U5053 ( .A1(n5103), .A2(n5126), .ZN(n5124) );
  OR2_X1 U5054 ( .A1(n5108), .A2(n5106), .ZN(n5126) );
  OR2_X1 U5055 ( .A1(n3951), .A2(n4073), .ZN(n5106) );
  OR2_X1 U5056 ( .A1(n5127), .A2(n5128), .ZN(n5108) );
  AND2_X1 U5057 ( .A1(n5095), .A2(n5097), .ZN(n5128) );
  AND2_X1 U5058 ( .A1(n5092), .A2(n5129), .ZN(n5127) );
  OR2_X1 U5059 ( .A1(n5097), .A2(n5095), .ZN(n5129) );
  OR2_X1 U5060 ( .A1(n4041), .A2(n4073), .ZN(n5095) );
  OR2_X1 U5061 ( .A1(n5130), .A2(n5131), .ZN(n5097) );
  AND2_X1 U5062 ( .A1(n5084), .A2(n5086), .ZN(n5131) );
  AND2_X1 U5063 ( .A1(n5081), .A2(n5132), .ZN(n5130) );
  OR2_X1 U5064 ( .A1(n5086), .A2(n5084), .ZN(n5132) );
  OR2_X1 U5065 ( .A1(n3888), .A2(n4073), .ZN(n5084) );
  OR2_X1 U5066 ( .A1(n5133), .A2(n5134), .ZN(n5086) );
  AND2_X1 U5067 ( .A1(n5073), .A2(n5075), .ZN(n5134) );
  AND2_X1 U5068 ( .A1(n5070), .A2(n5135), .ZN(n5133) );
  OR2_X1 U5069 ( .A1(n5075), .A2(n5073), .ZN(n5135) );
  OR2_X1 U5070 ( .A1(n4047), .A2(n4073), .ZN(n5073) );
  OR2_X1 U5071 ( .A1(n5136), .A2(n5137), .ZN(n5075) );
  AND2_X1 U5072 ( .A1(n5062), .A2(n5064), .ZN(n5137) );
  AND2_X1 U5073 ( .A1(n5059), .A2(n5138), .ZN(n5136) );
  OR2_X1 U5074 ( .A1(n5064), .A2(n5062), .ZN(n5138) );
  OR2_X1 U5075 ( .A1(n3837), .A2(n4073), .ZN(n5062) );
  OR2_X1 U5076 ( .A1(n5139), .A2(n5140), .ZN(n5064) );
  AND2_X1 U5077 ( .A1(n5051), .A2(n5053), .ZN(n5140) );
  AND2_X1 U5078 ( .A1(n5048), .A2(n5141), .ZN(n5139) );
  OR2_X1 U5079 ( .A1(n5053), .A2(n5051), .ZN(n5141) );
  OR2_X1 U5080 ( .A1(n4053), .A2(n4073), .ZN(n5051) );
  OR2_X1 U5081 ( .A1(n5142), .A2(n5143), .ZN(n5053) );
  AND2_X1 U5082 ( .A1(n5040), .A2(n5042), .ZN(n5143) );
  AND2_X1 U5083 ( .A1(n5037), .A2(n5144), .ZN(n5142) );
  OR2_X1 U5084 ( .A1(n5042), .A2(n5040), .ZN(n5144) );
  OR2_X1 U5085 ( .A1(n3786), .A2(n4073), .ZN(n5040) );
  OR2_X1 U5086 ( .A1(n5145), .A2(n5146), .ZN(n5042) );
  AND2_X1 U5087 ( .A1(n5029), .A2(n5032), .ZN(n5146) );
  AND2_X1 U5088 ( .A1(n5026), .A2(n5147), .ZN(n5145) );
  OR2_X1 U5089 ( .A1(n5032), .A2(n5029), .ZN(n5147) );
  OR2_X1 U5090 ( .A1(n4059), .A2(n4073), .ZN(n5029) );
  OR2_X1 U5091 ( .A1(n5148), .A2(n5149), .ZN(n5032) );
  AND2_X1 U5092 ( .A1(n5018), .A2(n5020), .ZN(n5149) );
  AND2_X1 U5093 ( .A1(n5015), .A2(n5150), .ZN(n5148) );
  OR2_X1 U5094 ( .A1(n5020), .A2(n5018), .ZN(n5150) );
  OR2_X1 U5095 ( .A1(n3735), .A2(n4073), .ZN(n5018) );
  OR2_X1 U5096 ( .A1(n5151), .A2(n5152), .ZN(n5020) );
  AND2_X1 U5097 ( .A1(n4065), .A2(n5010), .ZN(n5152) );
  AND2_X1 U5098 ( .A1(n5006), .A2(n5153), .ZN(n5151) );
  OR2_X1 U5099 ( .A1(n5010), .A2(n4065), .ZN(n5153) );
  OR2_X1 U5100 ( .A1(n4072), .A2(n4073), .ZN(n4065) );
  OR2_X1 U5101 ( .A1(n5154), .A2(n5155), .ZN(n5010) );
  AND2_X1 U5102 ( .A1(n4994), .A2(n5000), .ZN(n5155) );
  AND2_X1 U5103 ( .A1(n5001), .A2(n5156), .ZN(n5154) );
  OR2_X1 U5104 ( .A1(n5000), .A2(n4994), .ZN(n5156) );
  OR2_X1 U5105 ( .A1(n3682), .A2(n4073), .ZN(n4994) );
  OR2_X1 U5106 ( .A1(n3731), .A2(n5157), .ZN(n5000) );
  OR2_X1 U5107 ( .A1(n4070), .A2(n4073), .ZN(n5157) );
  INV_X1 U5108 ( .A(b_12_), .ZN(n4073) );
  INV_X1 U5109 ( .A(n4999), .ZN(n5001) );
  OR2_X1 U5110 ( .A1(n5158), .A2(n5159), .ZN(n4999) );
  AND2_X1 U5111 ( .A1(b_11_), .A2(n5160), .ZN(n5159) );
  OR2_X1 U5112 ( .A1(n5161), .A2(n3644), .ZN(n5160) );
  AND2_X1 U5113 ( .A1(a_14_), .A2(n4060), .ZN(n5161) );
  AND2_X1 U5114 ( .A1(b_10_), .A2(n5162), .ZN(n5158) );
  OR2_X1 U5115 ( .A1(n5163), .A2(n3647), .ZN(n5162) );
  AND2_X1 U5116 ( .A1(a_15_), .A2(n3731), .ZN(n5163) );
  OR2_X1 U5117 ( .A1(n5164), .A2(n5165), .ZN(n5006) );
  AND2_X1 U5118 ( .A1(n5166), .A2(n5167), .ZN(n5165) );
  INV_X1 U5119 ( .A(n5168), .ZN(n5164) );
  OR2_X1 U5120 ( .A1(n5166), .A2(n5167), .ZN(n5168) );
  OR2_X1 U5121 ( .A1(n5169), .A2(n5170), .ZN(n5166) );
  AND2_X1 U5122 ( .A1(n5171), .A2(n5172), .ZN(n5170) );
  INV_X1 U5123 ( .A(n5173), .ZN(n5171) );
  AND2_X1 U5124 ( .A1(n5174), .A2(n5173), .ZN(n5169) );
  OR2_X1 U5125 ( .A1(n5175), .A2(n5176), .ZN(n5015) );
  INV_X1 U5126 ( .A(n5177), .ZN(n5176) );
  OR2_X1 U5127 ( .A1(n5178), .A2(n5179), .ZN(n5177) );
  AND2_X1 U5128 ( .A1(n5179), .A2(n5178), .ZN(n5175) );
  AND2_X1 U5129 ( .A1(n5180), .A2(n5181), .ZN(n5178) );
  OR2_X1 U5130 ( .A1(n5182), .A2(n5183), .ZN(n5181) );
  INV_X1 U5131 ( .A(n5184), .ZN(n5183) );
  OR2_X1 U5132 ( .A1(n5184), .A2(n5185), .ZN(n5180) );
  INV_X1 U5133 ( .A(n5182), .ZN(n5185) );
  OR2_X1 U5134 ( .A1(n5186), .A2(n5187), .ZN(n5026) );
  INV_X1 U5135 ( .A(n5188), .ZN(n5187) );
  OR2_X1 U5136 ( .A1(n5189), .A2(n5190), .ZN(n5188) );
  AND2_X1 U5137 ( .A1(n5190), .A2(n5189), .ZN(n5186) );
  AND2_X1 U5138 ( .A1(n5191), .A2(n5192), .ZN(n5189) );
  OR2_X1 U5139 ( .A1(n4064), .A2(n5193), .ZN(n5192) );
  INV_X1 U5140 ( .A(n5194), .ZN(n5193) );
  OR2_X1 U5141 ( .A1(n5194), .A2(n3738), .ZN(n5191) );
  INV_X1 U5142 ( .A(n4064), .ZN(n3738) );
  OR2_X1 U5143 ( .A1(n5195), .A2(n5196), .ZN(n5037) );
  INV_X1 U5144 ( .A(n5197), .ZN(n5196) );
  OR2_X1 U5145 ( .A1(n5198), .A2(n5199), .ZN(n5197) );
  AND2_X1 U5146 ( .A1(n5199), .A2(n5198), .ZN(n5195) );
  AND2_X1 U5147 ( .A1(n5200), .A2(n5201), .ZN(n5198) );
  OR2_X1 U5148 ( .A1(n5202), .A2(n5203), .ZN(n5201) );
  INV_X1 U5149 ( .A(n5204), .ZN(n5200) );
  AND2_X1 U5150 ( .A1(n5203), .A2(n5202), .ZN(n5204) );
  INV_X1 U5151 ( .A(n5205), .ZN(n5203) );
  OR2_X1 U5152 ( .A1(n5206), .A2(n5207), .ZN(n5048) );
  INV_X1 U5153 ( .A(n5208), .ZN(n5207) );
  OR2_X1 U5154 ( .A1(n5209), .A2(n5210), .ZN(n5208) );
  AND2_X1 U5155 ( .A1(n5210), .A2(n5209), .ZN(n5206) );
  AND2_X1 U5156 ( .A1(n5211), .A2(n5212), .ZN(n5209) );
  OR2_X1 U5157 ( .A1(n5213), .A2(n5214), .ZN(n5212) );
  INV_X1 U5158 ( .A(n5215), .ZN(n5214) );
  OR2_X1 U5159 ( .A1(n5215), .A2(n5216), .ZN(n5211) );
  INV_X1 U5160 ( .A(n5213), .ZN(n5216) );
  OR2_X1 U5161 ( .A1(n5217), .A2(n5218), .ZN(n5059) );
  INV_X1 U5162 ( .A(n5219), .ZN(n5218) );
  OR2_X1 U5163 ( .A1(n5220), .A2(n5221), .ZN(n5219) );
  AND2_X1 U5164 ( .A1(n5221), .A2(n5220), .ZN(n5217) );
  AND2_X1 U5165 ( .A1(n5222), .A2(n5223), .ZN(n5220) );
  OR2_X1 U5166 ( .A1(n5224), .A2(n5225), .ZN(n5223) );
  INV_X1 U5167 ( .A(n5226), .ZN(n5225) );
  OR2_X1 U5168 ( .A1(n5226), .A2(n5227), .ZN(n5222) );
  INV_X1 U5169 ( .A(n5224), .ZN(n5227) );
  OR2_X1 U5170 ( .A1(n5228), .A2(n5229), .ZN(n5070) );
  INV_X1 U5171 ( .A(n5230), .ZN(n5229) );
  OR2_X1 U5172 ( .A1(n5231), .A2(n5232), .ZN(n5230) );
  AND2_X1 U5173 ( .A1(n5232), .A2(n5231), .ZN(n5228) );
  AND2_X1 U5174 ( .A1(n5233), .A2(n5234), .ZN(n5231) );
  OR2_X1 U5175 ( .A1(n5235), .A2(n5236), .ZN(n5234) );
  INV_X1 U5176 ( .A(n5237), .ZN(n5236) );
  OR2_X1 U5177 ( .A1(n5237), .A2(n5238), .ZN(n5233) );
  INV_X1 U5178 ( .A(n5235), .ZN(n5238) );
  OR2_X1 U5179 ( .A1(n5239), .A2(n5240), .ZN(n5081) );
  INV_X1 U5180 ( .A(n5241), .ZN(n5240) );
  OR2_X1 U5181 ( .A1(n5242), .A2(n5243), .ZN(n5241) );
  AND2_X1 U5182 ( .A1(n5243), .A2(n5242), .ZN(n5239) );
  AND2_X1 U5183 ( .A1(n5244), .A2(n5245), .ZN(n5242) );
  OR2_X1 U5184 ( .A1(n5246), .A2(n5247), .ZN(n5245) );
  INV_X1 U5185 ( .A(n5248), .ZN(n5247) );
  OR2_X1 U5186 ( .A1(n5248), .A2(n5249), .ZN(n5244) );
  INV_X1 U5187 ( .A(n5246), .ZN(n5249) );
  OR2_X1 U5188 ( .A1(n5250), .A2(n5251), .ZN(n5092) );
  INV_X1 U5189 ( .A(n5252), .ZN(n5251) );
  OR2_X1 U5190 ( .A1(n5253), .A2(n5254), .ZN(n5252) );
  AND2_X1 U5191 ( .A1(n5254), .A2(n5253), .ZN(n5250) );
  AND2_X1 U5192 ( .A1(n5255), .A2(n5256), .ZN(n5253) );
  OR2_X1 U5193 ( .A1(n5257), .A2(n5258), .ZN(n5256) );
  INV_X1 U5194 ( .A(n5259), .ZN(n5258) );
  OR2_X1 U5195 ( .A1(n5259), .A2(n5260), .ZN(n5255) );
  INV_X1 U5196 ( .A(n5257), .ZN(n5260) );
  OR2_X1 U5197 ( .A1(n5261), .A2(n5262), .ZN(n5103) );
  INV_X1 U5198 ( .A(n5263), .ZN(n5262) );
  OR2_X1 U5199 ( .A1(n5264), .A2(n5265), .ZN(n5263) );
  AND2_X1 U5200 ( .A1(n5265), .A2(n5264), .ZN(n5261) );
  AND2_X1 U5201 ( .A1(n5266), .A2(n5267), .ZN(n5264) );
  OR2_X1 U5202 ( .A1(n5268), .A2(n5269), .ZN(n5267) );
  INV_X1 U5203 ( .A(n5270), .ZN(n5269) );
  OR2_X1 U5204 ( .A1(n5270), .A2(n5271), .ZN(n5266) );
  INV_X1 U5205 ( .A(n5268), .ZN(n5271) );
  AND2_X1 U5206 ( .A1(n5272), .A2(n5273), .ZN(n4573) );
  INV_X1 U5207 ( .A(n5274), .ZN(n5273) );
  AND2_X1 U5208 ( .A1(n5275), .A2(n5276), .ZN(n5274) );
  OR2_X1 U5209 ( .A1(n5276), .A2(n5275), .ZN(n5272) );
  OR2_X1 U5210 ( .A1(n5277), .A2(n5278), .ZN(n5275) );
  AND2_X1 U5211 ( .A1(n5279), .A2(n5280), .ZN(n5278) );
  INV_X1 U5212 ( .A(n5281), .ZN(n5279) );
  AND2_X1 U5213 ( .A1(n5282), .A2(n5281), .ZN(n5277) );
  INV_X1 U5214 ( .A(n5280), .ZN(n5282) );
  OR2_X1 U5215 ( .A1(n5283), .A2(n5284), .ZN(n4584) );
  INV_X1 U5216 ( .A(n5285), .ZN(n5284) );
  OR2_X1 U5217 ( .A1(n5286), .A2(n5287), .ZN(n5285) );
  AND2_X1 U5218 ( .A1(n5287), .A2(n5286), .ZN(n5283) );
  AND2_X1 U5219 ( .A1(n5288), .A2(n5289), .ZN(n5286) );
  OR2_X1 U5220 ( .A1(n5290), .A2(n5291), .ZN(n5289) );
  INV_X1 U5221 ( .A(n5292), .ZN(n5291) );
  OR2_X1 U5222 ( .A1(n5292), .A2(n5293), .ZN(n5288) );
  INV_X1 U5223 ( .A(n5290), .ZN(n5293) );
  AND2_X1 U5224 ( .A1(n5294), .A2(n5295), .ZN(n4510) );
  INV_X1 U5225 ( .A(n5296), .ZN(n5295) );
  AND2_X1 U5226 ( .A1(n5297), .A2(n5298), .ZN(n5296) );
  OR2_X1 U5227 ( .A1(n5298), .A2(n5297), .ZN(n5294) );
  OR2_X1 U5228 ( .A1(n5299), .A2(n5300), .ZN(n5297) );
  AND2_X1 U5229 ( .A1(n5301), .A2(n5302), .ZN(n5300) );
  INV_X1 U5230 ( .A(n5303), .ZN(n5301) );
  AND2_X1 U5231 ( .A1(n5304), .A2(n5303), .ZN(n5299) );
  INV_X1 U5232 ( .A(n5302), .ZN(n5304) );
  AND2_X1 U5233 ( .A1(n5305), .A2(n5306), .ZN(n5111) );
  INV_X1 U5234 ( .A(n5307), .ZN(n5306) );
  AND2_X1 U5235 ( .A1(n5308), .A2(n5309), .ZN(n5307) );
  OR2_X1 U5236 ( .A1(n5309), .A2(n5308), .ZN(n5305) );
  OR2_X1 U5237 ( .A1(n5310), .A2(n5311), .ZN(n5308) );
  AND2_X1 U5238 ( .A1(n5312), .A2(n5313), .ZN(n5311) );
  INV_X1 U5239 ( .A(n5314), .ZN(n5310) );
  OR2_X1 U5240 ( .A1(n5313), .A2(n5312), .ZN(n5314) );
  AND2_X1 U5241 ( .A1(n5315), .A2(n4124), .ZN(n4120) );
  OR2_X1 U5242 ( .A1(n5316), .A2(n5317), .ZN(n4124) );
  INV_X1 U5243 ( .A(n5318), .ZN(n5315) );
  AND2_X1 U5244 ( .A1(n5316), .A2(n5317), .ZN(n5318) );
  OR2_X1 U5245 ( .A1(n5319), .A2(n5320), .ZN(n5317) );
  AND2_X1 U5246 ( .A1(n5321), .A2(n5313), .ZN(n5320) );
  AND2_X1 U5247 ( .A1(n5309), .A2(n5322), .ZN(n5319) );
  OR2_X1 U5248 ( .A1(n5313), .A2(n5321), .ZN(n5322) );
  INV_X1 U5249 ( .A(n5312), .ZN(n5321) );
  AND2_X1 U5250 ( .A1(a_0_), .A2(b_11_), .ZN(n5312) );
  OR2_X1 U5251 ( .A1(n5323), .A2(n5324), .ZN(n5313) );
  AND2_X1 U5252 ( .A1(n5303), .A2(n5302), .ZN(n5324) );
  AND2_X1 U5253 ( .A1(n5298), .A2(n5325), .ZN(n5323) );
  OR2_X1 U5254 ( .A1(n5302), .A2(n5303), .ZN(n5325) );
  OR2_X1 U5255 ( .A1(n4002), .A2(n3731), .ZN(n5303) );
  OR2_X1 U5256 ( .A1(n5326), .A2(n5327), .ZN(n5302) );
  AND2_X1 U5257 ( .A1(n5290), .A2(n5292), .ZN(n5327) );
  AND2_X1 U5258 ( .A1(n5287), .A2(n5328), .ZN(n5326) );
  OR2_X1 U5259 ( .A1(n5292), .A2(n5290), .ZN(n5328) );
  OR2_X1 U5260 ( .A1(n4035), .A2(n3731), .ZN(n5290) );
  OR2_X1 U5261 ( .A1(n5329), .A2(n5330), .ZN(n5292) );
  AND2_X1 U5262 ( .A1(n5281), .A2(n5280), .ZN(n5330) );
  AND2_X1 U5263 ( .A1(n5276), .A2(n5331), .ZN(n5329) );
  OR2_X1 U5264 ( .A1(n5280), .A2(n5281), .ZN(n5331) );
  OR2_X1 U5265 ( .A1(n3951), .A2(n3731), .ZN(n5281) );
  OR2_X1 U5266 ( .A1(n5332), .A2(n5333), .ZN(n5280) );
  AND2_X1 U5267 ( .A1(n5268), .A2(n5270), .ZN(n5333) );
  AND2_X1 U5268 ( .A1(n5265), .A2(n5334), .ZN(n5332) );
  OR2_X1 U5269 ( .A1(n5270), .A2(n5268), .ZN(n5334) );
  OR2_X1 U5270 ( .A1(n4041), .A2(n3731), .ZN(n5268) );
  OR2_X1 U5271 ( .A1(n5335), .A2(n5336), .ZN(n5270) );
  AND2_X1 U5272 ( .A1(n5257), .A2(n5259), .ZN(n5336) );
  AND2_X1 U5273 ( .A1(n5254), .A2(n5337), .ZN(n5335) );
  OR2_X1 U5274 ( .A1(n5259), .A2(n5257), .ZN(n5337) );
  OR2_X1 U5275 ( .A1(n3888), .A2(n3731), .ZN(n5257) );
  OR2_X1 U5276 ( .A1(n5338), .A2(n5339), .ZN(n5259) );
  AND2_X1 U5277 ( .A1(n5246), .A2(n5248), .ZN(n5339) );
  AND2_X1 U5278 ( .A1(n5243), .A2(n5340), .ZN(n5338) );
  OR2_X1 U5279 ( .A1(n5248), .A2(n5246), .ZN(n5340) );
  OR2_X1 U5280 ( .A1(n4047), .A2(n3731), .ZN(n5246) );
  OR2_X1 U5281 ( .A1(n5341), .A2(n5342), .ZN(n5248) );
  AND2_X1 U5282 ( .A1(n5235), .A2(n5237), .ZN(n5342) );
  AND2_X1 U5283 ( .A1(n5232), .A2(n5343), .ZN(n5341) );
  OR2_X1 U5284 ( .A1(n5237), .A2(n5235), .ZN(n5343) );
  OR2_X1 U5285 ( .A1(n3837), .A2(n3731), .ZN(n5235) );
  OR2_X1 U5286 ( .A1(n5344), .A2(n5345), .ZN(n5237) );
  AND2_X1 U5287 ( .A1(n5224), .A2(n5226), .ZN(n5345) );
  AND2_X1 U5288 ( .A1(n5221), .A2(n5346), .ZN(n5344) );
  OR2_X1 U5289 ( .A1(n5226), .A2(n5224), .ZN(n5346) );
  OR2_X1 U5290 ( .A1(n4053), .A2(n3731), .ZN(n5224) );
  OR2_X1 U5291 ( .A1(n5347), .A2(n5348), .ZN(n5226) );
  AND2_X1 U5292 ( .A1(n5213), .A2(n5215), .ZN(n5348) );
  AND2_X1 U5293 ( .A1(n5210), .A2(n5349), .ZN(n5347) );
  OR2_X1 U5294 ( .A1(n5215), .A2(n5213), .ZN(n5349) );
  OR2_X1 U5295 ( .A1(n3786), .A2(n3731), .ZN(n5213) );
  OR2_X1 U5296 ( .A1(n5350), .A2(n5351), .ZN(n5215) );
  AND2_X1 U5297 ( .A1(n5202), .A2(n5205), .ZN(n5351) );
  AND2_X1 U5298 ( .A1(n5199), .A2(n5352), .ZN(n5350) );
  OR2_X1 U5299 ( .A1(n5205), .A2(n5202), .ZN(n5352) );
  OR2_X1 U5300 ( .A1(n4059), .A2(n3731), .ZN(n5202) );
  OR2_X1 U5301 ( .A1(n5353), .A2(n5354), .ZN(n5205) );
  AND2_X1 U5302 ( .A1(n4064), .A2(n5194), .ZN(n5354) );
  AND2_X1 U5303 ( .A1(n5190), .A2(n5355), .ZN(n5353) );
  OR2_X1 U5304 ( .A1(n5194), .A2(n4064), .ZN(n5355) );
  OR2_X1 U5305 ( .A1(n3735), .A2(n3731), .ZN(n4064) );
  OR2_X1 U5306 ( .A1(n5356), .A2(n5357), .ZN(n5194) );
  AND2_X1 U5307 ( .A1(n5182), .A2(n5184), .ZN(n5357) );
  AND2_X1 U5308 ( .A1(n5179), .A2(n5358), .ZN(n5356) );
  OR2_X1 U5309 ( .A1(n5184), .A2(n5182), .ZN(n5358) );
  OR2_X1 U5310 ( .A1(n4072), .A2(n3731), .ZN(n5182) );
  OR2_X1 U5311 ( .A1(n5359), .A2(n5360), .ZN(n5184) );
  AND2_X1 U5312 ( .A1(n5167), .A2(n5173), .ZN(n5360) );
  AND2_X1 U5313 ( .A1(n5174), .A2(n5361), .ZN(n5359) );
  OR2_X1 U5314 ( .A1(n5173), .A2(n5167), .ZN(n5361) );
  OR2_X1 U5315 ( .A1(n3682), .A2(n3731), .ZN(n5167) );
  OR2_X1 U5316 ( .A1(n3731), .A2(n5362), .ZN(n5173) );
  OR2_X1 U5317 ( .A1(n4070), .A2(n4060), .ZN(n5362) );
  INV_X1 U5318 ( .A(b_11_), .ZN(n3731) );
  INV_X1 U5319 ( .A(n5172), .ZN(n5174) );
  OR2_X1 U5320 ( .A1(n5363), .A2(n5364), .ZN(n5172) );
  AND2_X1 U5321 ( .A1(b_9_), .A2(n5365), .ZN(n5364) );
  OR2_X1 U5322 ( .A1(n5366), .A2(n3647), .ZN(n5365) );
  AND2_X1 U5323 ( .A1(a_15_), .A2(n4060), .ZN(n5366) );
  AND2_X1 U5324 ( .A1(b_10_), .A2(n5367), .ZN(n5363) );
  OR2_X1 U5325 ( .A1(n5368), .A2(n3644), .ZN(n5367) );
  AND2_X1 U5326 ( .A1(a_14_), .A2(n3782), .ZN(n5368) );
  OR2_X1 U5327 ( .A1(n5369), .A2(n5370), .ZN(n5179) );
  AND2_X1 U5328 ( .A1(n5371), .A2(n5372), .ZN(n5370) );
  INV_X1 U5329 ( .A(n5373), .ZN(n5369) );
  OR2_X1 U5330 ( .A1(n5371), .A2(n5372), .ZN(n5373) );
  OR2_X1 U5331 ( .A1(n5374), .A2(n5375), .ZN(n5371) );
  AND2_X1 U5332 ( .A1(n5376), .A2(n5377), .ZN(n5375) );
  INV_X1 U5333 ( .A(n5378), .ZN(n5376) );
  AND2_X1 U5334 ( .A1(n5379), .A2(n5378), .ZN(n5374) );
  OR2_X1 U5335 ( .A1(n5380), .A2(n5381), .ZN(n5190) );
  INV_X1 U5336 ( .A(n5382), .ZN(n5381) );
  OR2_X1 U5337 ( .A1(n5383), .A2(n5384), .ZN(n5382) );
  AND2_X1 U5338 ( .A1(n5384), .A2(n5383), .ZN(n5380) );
  AND2_X1 U5339 ( .A1(n5385), .A2(n5386), .ZN(n5383) );
  OR2_X1 U5340 ( .A1(n5387), .A2(n5388), .ZN(n5386) );
  INV_X1 U5341 ( .A(n5389), .ZN(n5388) );
  OR2_X1 U5342 ( .A1(n5389), .A2(n5390), .ZN(n5385) );
  INV_X1 U5343 ( .A(n5387), .ZN(n5390) );
  OR2_X1 U5344 ( .A1(n5391), .A2(n5392), .ZN(n5199) );
  INV_X1 U5345 ( .A(n5393), .ZN(n5392) );
  OR2_X1 U5346 ( .A1(n5394), .A2(n5395), .ZN(n5393) );
  AND2_X1 U5347 ( .A1(n5395), .A2(n5394), .ZN(n5391) );
  AND2_X1 U5348 ( .A1(n5396), .A2(n5397), .ZN(n5394) );
  OR2_X1 U5349 ( .A1(n5398), .A2(n5399), .ZN(n5397) );
  INV_X1 U5350 ( .A(n5400), .ZN(n5399) );
  OR2_X1 U5351 ( .A1(n5400), .A2(n5401), .ZN(n5396) );
  INV_X1 U5352 ( .A(n5398), .ZN(n5401) );
  OR2_X1 U5353 ( .A1(n5402), .A2(n5403), .ZN(n5210) );
  INV_X1 U5354 ( .A(n5404), .ZN(n5403) );
  OR2_X1 U5355 ( .A1(n5405), .A2(n5406), .ZN(n5404) );
  AND2_X1 U5356 ( .A1(n5406), .A2(n5405), .ZN(n5402) );
  AND2_X1 U5357 ( .A1(n5407), .A2(n5408), .ZN(n5405) );
  OR2_X1 U5358 ( .A1(n5409), .A2(n3761), .ZN(n5408) );
  OR2_X1 U5359 ( .A1(n4061), .A2(n5410), .ZN(n5407) );
  INV_X1 U5360 ( .A(n5409), .ZN(n5410) );
  OR2_X1 U5361 ( .A1(n5411), .A2(n5412), .ZN(n5221) );
  INV_X1 U5362 ( .A(n5413), .ZN(n5412) );
  OR2_X1 U5363 ( .A1(n5414), .A2(n5415), .ZN(n5413) );
  AND2_X1 U5364 ( .A1(n5415), .A2(n5414), .ZN(n5411) );
  AND2_X1 U5365 ( .A1(n5416), .A2(n5417), .ZN(n5414) );
  OR2_X1 U5366 ( .A1(n5418), .A2(n5419), .ZN(n5417) );
  INV_X1 U5367 ( .A(n5420), .ZN(n5419) );
  OR2_X1 U5368 ( .A1(n5420), .A2(n5421), .ZN(n5416) );
  INV_X1 U5369 ( .A(n5418), .ZN(n5421) );
  OR2_X1 U5370 ( .A1(n5422), .A2(n5423), .ZN(n5232) );
  INV_X1 U5371 ( .A(n5424), .ZN(n5423) );
  OR2_X1 U5372 ( .A1(n5425), .A2(n5426), .ZN(n5424) );
  AND2_X1 U5373 ( .A1(n5426), .A2(n5425), .ZN(n5422) );
  AND2_X1 U5374 ( .A1(n5427), .A2(n5428), .ZN(n5425) );
  OR2_X1 U5375 ( .A1(n5429), .A2(n5430), .ZN(n5428) );
  INV_X1 U5376 ( .A(n5431), .ZN(n5430) );
  OR2_X1 U5377 ( .A1(n5431), .A2(n5432), .ZN(n5427) );
  INV_X1 U5378 ( .A(n5429), .ZN(n5432) );
  OR2_X1 U5379 ( .A1(n5433), .A2(n5434), .ZN(n5243) );
  INV_X1 U5380 ( .A(n5435), .ZN(n5434) );
  OR2_X1 U5381 ( .A1(n5436), .A2(n5437), .ZN(n5435) );
  AND2_X1 U5382 ( .A1(n5437), .A2(n5436), .ZN(n5433) );
  AND2_X1 U5383 ( .A1(n5438), .A2(n5439), .ZN(n5436) );
  OR2_X1 U5384 ( .A1(n5440), .A2(n5441), .ZN(n5439) );
  INV_X1 U5385 ( .A(n5442), .ZN(n5441) );
  OR2_X1 U5386 ( .A1(n5442), .A2(n5443), .ZN(n5438) );
  INV_X1 U5387 ( .A(n5440), .ZN(n5443) );
  OR2_X1 U5388 ( .A1(n5444), .A2(n5445), .ZN(n5254) );
  INV_X1 U5389 ( .A(n5446), .ZN(n5445) );
  OR2_X1 U5390 ( .A1(n5447), .A2(n5448), .ZN(n5446) );
  AND2_X1 U5391 ( .A1(n5448), .A2(n5447), .ZN(n5444) );
  AND2_X1 U5392 ( .A1(n5449), .A2(n5450), .ZN(n5447) );
  OR2_X1 U5393 ( .A1(n5451), .A2(n5452), .ZN(n5450) );
  INV_X1 U5394 ( .A(n5453), .ZN(n5452) );
  OR2_X1 U5395 ( .A1(n5453), .A2(n5454), .ZN(n5449) );
  INV_X1 U5396 ( .A(n5451), .ZN(n5454) );
  OR2_X1 U5397 ( .A1(n5455), .A2(n5456), .ZN(n5265) );
  INV_X1 U5398 ( .A(n5457), .ZN(n5456) );
  OR2_X1 U5399 ( .A1(n5458), .A2(n5459), .ZN(n5457) );
  AND2_X1 U5400 ( .A1(n5459), .A2(n5458), .ZN(n5455) );
  AND2_X1 U5401 ( .A1(n5460), .A2(n5461), .ZN(n5458) );
  OR2_X1 U5402 ( .A1(n5462), .A2(n5463), .ZN(n5461) );
  INV_X1 U5403 ( .A(n5464), .ZN(n5463) );
  OR2_X1 U5404 ( .A1(n5464), .A2(n5465), .ZN(n5460) );
  INV_X1 U5405 ( .A(n5462), .ZN(n5465) );
  AND2_X1 U5406 ( .A1(n5466), .A2(n5467), .ZN(n5276) );
  INV_X1 U5407 ( .A(n5468), .ZN(n5467) );
  AND2_X1 U5408 ( .A1(n5469), .A2(n5470), .ZN(n5468) );
  OR2_X1 U5409 ( .A1(n5470), .A2(n5469), .ZN(n5466) );
  OR2_X1 U5410 ( .A1(n5471), .A2(n5472), .ZN(n5469) );
  AND2_X1 U5411 ( .A1(n5473), .A2(n5474), .ZN(n5472) );
  INV_X1 U5412 ( .A(n5475), .ZN(n5473) );
  AND2_X1 U5413 ( .A1(n5476), .A2(n5475), .ZN(n5471) );
  INV_X1 U5414 ( .A(n5474), .ZN(n5476) );
  OR2_X1 U5415 ( .A1(n5477), .A2(n5478), .ZN(n5287) );
  INV_X1 U5416 ( .A(n5479), .ZN(n5478) );
  OR2_X1 U5417 ( .A1(n5480), .A2(n5481), .ZN(n5479) );
  AND2_X1 U5418 ( .A1(n5481), .A2(n5480), .ZN(n5477) );
  AND2_X1 U5419 ( .A1(n5482), .A2(n5483), .ZN(n5480) );
  OR2_X1 U5420 ( .A1(n5484), .A2(n5485), .ZN(n5483) );
  INV_X1 U5421 ( .A(n5486), .ZN(n5485) );
  OR2_X1 U5422 ( .A1(n5486), .A2(n5487), .ZN(n5482) );
  INV_X1 U5423 ( .A(n5484), .ZN(n5487) );
  AND2_X1 U5424 ( .A1(n5488), .A2(n5489), .ZN(n5298) );
  INV_X1 U5425 ( .A(n5490), .ZN(n5489) );
  AND2_X1 U5426 ( .A1(n5491), .A2(n5492), .ZN(n5490) );
  OR2_X1 U5427 ( .A1(n5492), .A2(n5491), .ZN(n5488) );
  OR2_X1 U5428 ( .A1(n5493), .A2(n5494), .ZN(n5491) );
  AND2_X1 U5429 ( .A1(n5495), .A2(n5496), .ZN(n5494) );
  INV_X1 U5430 ( .A(n5497), .ZN(n5495) );
  AND2_X1 U5431 ( .A1(n5498), .A2(n5497), .ZN(n5493) );
  INV_X1 U5432 ( .A(n5496), .ZN(n5498) );
  AND2_X1 U5433 ( .A1(n5499), .A2(n5500), .ZN(n5309) );
  INV_X1 U5434 ( .A(n5501), .ZN(n5500) );
  AND2_X1 U5435 ( .A1(n5502), .A2(n5503), .ZN(n5501) );
  OR2_X1 U5436 ( .A1(n5503), .A2(n5502), .ZN(n5499) );
  OR2_X1 U5437 ( .A1(n5504), .A2(n5505), .ZN(n5502) );
  AND2_X1 U5438 ( .A1(n5506), .A2(n5507), .ZN(n5505) );
  INV_X1 U5439 ( .A(n5508), .ZN(n5506) );
  AND2_X1 U5440 ( .A1(n5509), .A2(n5508), .ZN(n5504) );
  INV_X1 U5441 ( .A(n5507), .ZN(n5509) );
  AND2_X1 U5442 ( .A1(n5510), .A2(n5511), .ZN(n5316) );
  INV_X1 U5443 ( .A(n5512), .ZN(n5511) );
  AND2_X1 U5444 ( .A1(n5513), .A2(n5514), .ZN(n5512) );
  OR2_X1 U5445 ( .A1(n5514), .A2(n5513), .ZN(n5510) );
  OR2_X1 U5446 ( .A1(n5515), .A2(n5516), .ZN(n5513) );
  AND2_X1 U5447 ( .A1(n5517), .A2(n5518), .ZN(n5516) );
  INV_X1 U5448 ( .A(n5519), .ZN(n5515) );
  OR2_X1 U5449 ( .A1(n5518), .A2(n5517), .ZN(n5519) );
  AND2_X1 U5450 ( .A1(n5520), .A2(n3541), .ZN(n4132) );
  OR2_X1 U5451 ( .A1(n5521), .A2(n5522), .ZN(n3541) );
  INV_X1 U5452 ( .A(n5523), .ZN(n5520) );
  AND2_X1 U5453 ( .A1(n5521), .A2(n5522), .ZN(n5523) );
  OR2_X1 U5454 ( .A1(n5524), .A2(n5525), .ZN(n5522) );
  AND2_X1 U5455 ( .A1(n5526), .A2(n5518), .ZN(n5525) );
  AND2_X1 U5456 ( .A1(n5514), .A2(n5527), .ZN(n5524) );
  OR2_X1 U5457 ( .A1(n5526), .A2(n5518), .ZN(n5527) );
  OR2_X1 U5458 ( .A1(n5528), .A2(n5529), .ZN(n5518) );
  AND2_X1 U5459 ( .A1(n5508), .A2(n5507), .ZN(n5529) );
  AND2_X1 U5460 ( .A1(n5503), .A2(n5530), .ZN(n5528) );
  OR2_X1 U5461 ( .A1(n5508), .A2(n5507), .ZN(n5530) );
  OR2_X1 U5462 ( .A1(n5531), .A2(n5532), .ZN(n5507) );
  AND2_X1 U5463 ( .A1(n5497), .A2(n5496), .ZN(n5532) );
  AND2_X1 U5464 ( .A1(n5492), .A2(n5533), .ZN(n5531) );
  OR2_X1 U5465 ( .A1(n5497), .A2(n5496), .ZN(n5533) );
  OR2_X1 U5466 ( .A1(n5534), .A2(n5535), .ZN(n5496) );
  AND2_X1 U5467 ( .A1(n5481), .A2(n5484), .ZN(n5535) );
  AND2_X1 U5468 ( .A1(n5536), .A2(n5486), .ZN(n5534) );
  OR2_X1 U5469 ( .A1(n5537), .A2(n5538), .ZN(n5486) );
  AND2_X1 U5470 ( .A1(n5475), .A2(n5474), .ZN(n5538) );
  AND2_X1 U5471 ( .A1(n5470), .A2(n5539), .ZN(n5537) );
  OR2_X1 U5472 ( .A1(n5475), .A2(n5474), .ZN(n5539) );
  OR2_X1 U5473 ( .A1(n5540), .A2(n5541), .ZN(n5474) );
  AND2_X1 U5474 ( .A1(n5459), .A2(n5462), .ZN(n5541) );
  AND2_X1 U5475 ( .A1(n5542), .A2(n5464), .ZN(n5540) );
  OR2_X1 U5476 ( .A1(n5543), .A2(n5544), .ZN(n5464) );
  AND2_X1 U5477 ( .A1(n5448), .A2(n5451), .ZN(n5544) );
  AND2_X1 U5478 ( .A1(n5545), .A2(n5453), .ZN(n5543) );
  OR2_X1 U5479 ( .A1(n5546), .A2(n5547), .ZN(n5453) );
  AND2_X1 U5480 ( .A1(n5437), .A2(n5440), .ZN(n5547) );
  AND2_X1 U5481 ( .A1(n5548), .A2(n5442), .ZN(n5546) );
  OR2_X1 U5482 ( .A1(n5549), .A2(n5550), .ZN(n5442) );
  AND2_X1 U5483 ( .A1(n5426), .A2(n5429), .ZN(n5550) );
  AND2_X1 U5484 ( .A1(n5551), .A2(n5431), .ZN(n5549) );
  OR2_X1 U5485 ( .A1(n5552), .A2(n5553), .ZN(n5431) );
  AND2_X1 U5486 ( .A1(n5415), .A2(n5418), .ZN(n5553) );
  AND2_X1 U5487 ( .A1(n5554), .A2(n5420), .ZN(n5552) );
  OR2_X1 U5488 ( .A1(n5555), .A2(n5556), .ZN(n5420) );
  AND2_X1 U5489 ( .A1(n5406), .A2(n4061), .ZN(n5556) );
  AND2_X1 U5490 ( .A1(n5557), .A2(n5409), .ZN(n5555) );
  OR2_X1 U5491 ( .A1(n5558), .A2(n5559), .ZN(n5409) );
  AND2_X1 U5492 ( .A1(n5395), .A2(n5398), .ZN(n5559) );
  AND2_X1 U5493 ( .A1(n5560), .A2(n5400), .ZN(n5558) );
  OR2_X1 U5494 ( .A1(n5561), .A2(n5562), .ZN(n5400) );
  AND2_X1 U5495 ( .A1(n5384), .A2(n5387), .ZN(n5562) );
  AND2_X1 U5496 ( .A1(n5563), .A2(n5389), .ZN(n5561) );
  OR2_X1 U5497 ( .A1(n5564), .A2(n5565), .ZN(n5389) );
  AND2_X1 U5498 ( .A1(n5372), .A2(n5378), .ZN(n5565) );
  AND2_X1 U5499 ( .A1(n5379), .A2(n5566), .ZN(n5564) );
  OR2_X1 U5500 ( .A1(n5372), .A2(n5378), .ZN(n5566) );
  OR2_X1 U5501 ( .A1(n4060), .A2(n5567), .ZN(n5378) );
  OR2_X1 U5502 ( .A1(n3782), .A2(n4070), .ZN(n5567) );
  OR2_X1 U5503 ( .A1(n4060), .A2(n3682), .ZN(n5372) );
  INV_X1 U5504 ( .A(n5377), .ZN(n5379) );
  OR2_X1 U5505 ( .A1(n5568), .A2(n5569), .ZN(n5377) );
  AND2_X1 U5506 ( .A1(b_9_), .A2(n5570), .ZN(n5569) );
  OR2_X1 U5507 ( .A1(n5571), .A2(n3644), .ZN(n5570) );
  AND2_X1 U5508 ( .A1(a_14_), .A2(n4054), .ZN(n5571) );
  AND2_X1 U5509 ( .A1(b_8_), .A2(n5572), .ZN(n5568) );
  OR2_X1 U5510 ( .A1(n5573), .A2(n3647), .ZN(n5572) );
  AND2_X1 U5511 ( .A1(a_15_), .A2(n3782), .ZN(n5573) );
  OR2_X1 U5512 ( .A1(n5384), .A2(n5387), .ZN(n5563) );
  OR2_X1 U5513 ( .A1(n4060), .A2(n4072), .ZN(n5387) );
  OR2_X1 U5514 ( .A1(n5574), .A2(n5575), .ZN(n5384) );
  AND2_X1 U5515 ( .A1(n5576), .A2(n5577), .ZN(n5575) );
  INV_X1 U5516 ( .A(n5578), .ZN(n5574) );
  OR2_X1 U5517 ( .A1(n5576), .A2(n5577), .ZN(n5578) );
  OR2_X1 U5518 ( .A1(n5579), .A2(n5580), .ZN(n5576) );
  AND2_X1 U5519 ( .A1(n5581), .A2(n5582), .ZN(n5580) );
  INV_X1 U5520 ( .A(n5583), .ZN(n5581) );
  AND2_X1 U5521 ( .A1(n5584), .A2(n5583), .ZN(n5579) );
  OR2_X1 U5522 ( .A1(n5395), .A2(n5398), .ZN(n5560) );
  OR2_X1 U5523 ( .A1(n4060), .A2(n3735), .ZN(n5398) );
  OR2_X1 U5524 ( .A1(n5585), .A2(n5586), .ZN(n5395) );
  INV_X1 U5525 ( .A(n5587), .ZN(n5586) );
  OR2_X1 U5526 ( .A1(n5588), .A2(n5589), .ZN(n5587) );
  AND2_X1 U5527 ( .A1(n5589), .A2(n5588), .ZN(n5585) );
  AND2_X1 U5528 ( .A1(n5590), .A2(n5591), .ZN(n5588) );
  OR2_X1 U5529 ( .A1(n5592), .A2(n5593), .ZN(n5591) );
  INV_X1 U5530 ( .A(n5594), .ZN(n5593) );
  OR2_X1 U5531 ( .A1(n5594), .A2(n5595), .ZN(n5590) );
  INV_X1 U5532 ( .A(n5592), .ZN(n5595) );
  OR2_X1 U5533 ( .A1(n5406), .A2(n4061), .ZN(n5557) );
  INV_X1 U5534 ( .A(n3761), .ZN(n4061) );
  AND2_X1 U5535 ( .A1(b_10_), .A2(a_10_), .ZN(n3761) );
  OR2_X1 U5536 ( .A1(n5596), .A2(n5597), .ZN(n5406) );
  INV_X1 U5537 ( .A(n5598), .ZN(n5597) );
  OR2_X1 U5538 ( .A1(n5599), .A2(n5600), .ZN(n5598) );
  AND2_X1 U5539 ( .A1(n5600), .A2(n5599), .ZN(n5596) );
  AND2_X1 U5540 ( .A1(n5601), .A2(n5602), .ZN(n5599) );
  OR2_X1 U5541 ( .A1(n5603), .A2(n5604), .ZN(n5602) );
  INV_X1 U5542 ( .A(n5605), .ZN(n5604) );
  OR2_X1 U5543 ( .A1(n5605), .A2(n5606), .ZN(n5601) );
  INV_X1 U5544 ( .A(n5603), .ZN(n5606) );
  OR2_X1 U5545 ( .A1(n5415), .A2(n5418), .ZN(n5554) );
  OR2_X1 U5546 ( .A1(n4060), .A2(n3786), .ZN(n5418) );
  OR2_X1 U5547 ( .A1(n5607), .A2(n5608), .ZN(n5415) );
  INV_X1 U5548 ( .A(n5609), .ZN(n5608) );
  OR2_X1 U5549 ( .A1(n5610), .A2(n5611), .ZN(n5609) );
  AND2_X1 U5550 ( .A1(n5611), .A2(n5610), .ZN(n5607) );
  AND2_X1 U5551 ( .A1(n5612), .A2(n5613), .ZN(n5610) );
  OR2_X1 U5552 ( .A1(n5614), .A2(n5615), .ZN(n5613) );
  INV_X1 U5553 ( .A(n5616), .ZN(n5612) );
  AND2_X1 U5554 ( .A1(n5615), .A2(n5614), .ZN(n5616) );
  INV_X1 U5555 ( .A(n5617), .ZN(n5615) );
  OR2_X1 U5556 ( .A1(n5426), .A2(n5429), .ZN(n5551) );
  OR2_X1 U5557 ( .A1(n4060), .A2(n4053), .ZN(n5429) );
  OR2_X1 U5558 ( .A1(n5618), .A2(n5619), .ZN(n5426) );
  INV_X1 U5559 ( .A(n5620), .ZN(n5619) );
  OR2_X1 U5560 ( .A1(n5621), .A2(n5622), .ZN(n5620) );
  AND2_X1 U5561 ( .A1(n5622), .A2(n5621), .ZN(n5618) );
  AND2_X1 U5562 ( .A1(n5623), .A2(n5624), .ZN(n5621) );
  OR2_X1 U5563 ( .A1(n4057), .A2(n5625), .ZN(n5624) );
  INV_X1 U5564 ( .A(n5626), .ZN(n5625) );
  OR2_X1 U5565 ( .A1(n5626), .A2(n3789), .ZN(n5623) );
  INV_X1 U5566 ( .A(n4057), .ZN(n3789) );
  OR2_X1 U5567 ( .A1(n5437), .A2(n5440), .ZN(n5548) );
  OR2_X1 U5568 ( .A1(n4060), .A2(n3837), .ZN(n5440) );
  OR2_X1 U5569 ( .A1(n5627), .A2(n5628), .ZN(n5437) );
  INV_X1 U5570 ( .A(n5629), .ZN(n5628) );
  OR2_X1 U5571 ( .A1(n5630), .A2(n5631), .ZN(n5629) );
  AND2_X1 U5572 ( .A1(n5631), .A2(n5630), .ZN(n5627) );
  AND2_X1 U5573 ( .A1(n5632), .A2(n5633), .ZN(n5630) );
  OR2_X1 U5574 ( .A1(n5634), .A2(n5635), .ZN(n5633) );
  INV_X1 U5575 ( .A(n5636), .ZN(n5635) );
  OR2_X1 U5576 ( .A1(n5636), .A2(n5637), .ZN(n5632) );
  INV_X1 U5577 ( .A(n5634), .ZN(n5637) );
  OR2_X1 U5578 ( .A1(n5448), .A2(n5451), .ZN(n5545) );
  OR2_X1 U5579 ( .A1(n4060), .A2(n4047), .ZN(n5451) );
  OR2_X1 U5580 ( .A1(n5638), .A2(n5639), .ZN(n5448) );
  INV_X1 U5581 ( .A(n5640), .ZN(n5639) );
  OR2_X1 U5582 ( .A1(n5641), .A2(n5642), .ZN(n5640) );
  AND2_X1 U5583 ( .A1(n5642), .A2(n5641), .ZN(n5638) );
  AND2_X1 U5584 ( .A1(n5643), .A2(n5644), .ZN(n5641) );
  OR2_X1 U5585 ( .A1(n5645), .A2(n5646), .ZN(n5644) );
  INV_X1 U5586 ( .A(n5647), .ZN(n5646) );
  OR2_X1 U5587 ( .A1(n5647), .A2(n5648), .ZN(n5643) );
  INV_X1 U5588 ( .A(n5645), .ZN(n5648) );
  OR2_X1 U5589 ( .A1(n5459), .A2(n5462), .ZN(n5542) );
  OR2_X1 U5590 ( .A1(n4060), .A2(n3888), .ZN(n5462) );
  OR2_X1 U5591 ( .A1(n5649), .A2(n5650), .ZN(n5459) );
  INV_X1 U5592 ( .A(n5651), .ZN(n5650) );
  OR2_X1 U5593 ( .A1(n5652), .A2(n5653), .ZN(n5651) );
  AND2_X1 U5594 ( .A1(n5653), .A2(n5652), .ZN(n5649) );
  AND2_X1 U5595 ( .A1(n5654), .A2(n5655), .ZN(n5652) );
  OR2_X1 U5596 ( .A1(n5656), .A2(n5657), .ZN(n5655) );
  INV_X1 U5597 ( .A(n5658), .ZN(n5657) );
  OR2_X1 U5598 ( .A1(n5658), .A2(n5659), .ZN(n5654) );
  INV_X1 U5599 ( .A(n5656), .ZN(n5659) );
  OR2_X1 U5600 ( .A1(n4060), .A2(n4041), .ZN(n5475) );
  AND2_X1 U5601 ( .A1(n5660), .A2(n5661), .ZN(n5470) );
  INV_X1 U5602 ( .A(n5662), .ZN(n5661) );
  AND2_X1 U5603 ( .A1(n5663), .A2(n5664), .ZN(n5662) );
  OR2_X1 U5604 ( .A1(n5664), .A2(n5663), .ZN(n5660) );
  OR2_X1 U5605 ( .A1(n5665), .A2(n5666), .ZN(n5663) );
  AND2_X1 U5606 ( .A1(n5667), .A2(n5668), .ZN(n5666) );
  INV_X1 U5607 ( .A(n5669), .ZN(n5667) );
  AND2_X1 U5608 ( .A1(n5670), .A2(n5669), .ZN(n5665) );
  INV_X1 U5609 ( .A(n5668), .ZN(n5670) );
  OR2_X1 U5610 ( .A1(n5481), .A2(n5484), .ZN(n5536) );
  OR2_X1 U5611 ( .A1(n4060), .A2(n3951), .ZN(n5484) );
  OR2_X1 U5612 ( .A1(n5671), .A2(n5672), .ZN(n5481) );
  INV_X1 U5613 ( .A(n5673), .ZN(n5672) );
  OR2_X1 U5614 ( .A1(n5674), .A2(n5675), .ZN(n5673) );
  AND2_X1 U5615 ( .A1(n5675), .A2(n5674), .ZN(n5671) );
  AND2_X1 U5616 ( .A1(n5676), .A2(n5677), .ZN(n5674) );
  OR2_X1 U5617 ( .A1(n5678), .A2(n5679), .ZN(n5677) );
  INV_X1 U5618 ( .A(n5680), .ZN(n5679) );
  OR2_X1 U5619 ( .A1(n5680), .A2(n5681), .ZN(n5676) );
  INV_X1 U5620 ( .A(n5678), .ZN(n5681) );
  OR2_X1 U5621 ( .A1(n4060), .A2(n4035), .ZN(n5497) );
  AND2_X1 U5622 ( .A1(n5682), .A2(n5683), .ZN(n5492) );
  INV_X1 U5623 ( .A(n5684), .ZN(n5683) );
  AND2_X1 U5624 ( .A1(n5685), .A2(n5686), .ZN(n5684) );
  OR2_X1 U5625 ( .A1(n5686), .A2(n5685), .ZN(n5682) );
  OR2_X1 U5626 ( .A1(n5687), .A2(n5688), .ZN(n5685) );
  AND2_X1 U5627 ( .A1(n5689), .A2(n5690), .ZN(n5688) );
  INV_X1 U5628 ( .A(n5691), .ZN(n5689) );
  AND2_X1 U5629 ( .A1(n5692), .A2(n5691), .ZN(n5687) );
  INV_X1 U5630 ( .A(n5690), .ZN(n5692) );
  OR2_X1 U5631 ( .A1(n4060), .A2(n4002), .ZN(n5508) );
  INV_X1 U5632 ( .A(b_10_), .ZN(n4060) );
  AND2_X1 U5633 ( .A1(n5693), .A2(n5694), .ZN(n5503) );
  INV_X1 U5634 ( .A(n5695), .ZN(n5694) );
  AND2_X1 U5635 ( .A1(n5696), .A2(n5697), .ZN(n5695) );
  OR2_X1 U5636 ( .A1(n5697), .A2(n5696), .ZN(n5693) );
  OR2_X1 U5637 ( .A1(n5698), .A2(n5699), .ZN(n5696) );
  AND2_X1 U5638 ( .A1(n5700), .A2(n5701), .ZN(n5699) );
  INV_X1 U5639 ( .A(n5702), .ZN(n5700) );
  AND2_X1 U5640 ( .A1(n5703), .A2(n5702), .ZN(n5698) );
  INV_X1 U5641 ( .A(n5701), .ZN(n5703) );
  INV_X1 U5642 ( .A(n5517), .ZN(n5526) );
  AND2_X1 U5643 ( .A1(b_10_), .A2(a_0_), .ZN(n5517) );
  AND2_X1 U5644 ( .A1(n5704), .A2(n5705), .ZN(n5514) );
  INV_X1 U5645 ( .A(n5706), .ZN(n5705) );
  AND2_X1 U5646 ( .A1(n5707), .A2(n5708), .ZN(n5706) );
  OR2_X1 U5647 ( .A1(n5708), .A2(n5707), .ZN(n5704) );
  OR2_X1 U5648 ( .A1(n5709), .A2(n5710), .ZN(n5707) );
  AND2_X1 U5649 ( .A1(n5711), .A2(n5712), .ZN(n5710) );
  INV_X1 U5650 ( .A(n5713), .ZN(n5711) );
  AND2_X1 U5651 ( .A1(n5714), .A2(n5713), .ZN(n5709) );
  INV_X1 U5652 ( .A(n5712), .ZN(n5714) );
  AND2_X1 U5653 ( .A1(n5715), .A2(n5716), .ZN(n5521) );
  INV_X1 U5654 ( .A(n5717), .ZN(n5716) );
  AND2_X1 U5655 ( .A1(n5718), .A2(n5719), .ZN(n5717) );
  OR2_X1 U5656 ( .A1(n5719), .A2(n5718), .ZN(n5715) );
  OR2_X1 U5657 ( .A1(n5720), .A2(n5721), .ZN(n5718) );
  AND2_X1 U5658 ( .A1(n5722), .A2(n5723), .ZN(n5721) );
  INV_X1 U5659 ( .A(n5724), .ZN(n5720) );
  OR2_X1 U5660 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  INV_X1 U5661 ( .A(n3557), .ZN(n3558) );
  OR2_X1 U5662 ( .A1(n4489), .A2(n4490), .ZN(n3557) );
  OR2_X1 U5663 ( .A1(n5725), .A2(n5726), .ZN(n4490) );
  AND2_X1 U5664 ( .A1(n5727), .A2(n5723), .ZN(n5726) );
  AND2_X1 U5665 ( .A1(n5719), .A2(n5728), .ZN(n5725) );
  OR2_X1 U5666 ( .A1(n5723), .A2(n5727), .ZN(n5728) );
  INV_X1 U5667 ( .A(n5722), .ZN(n5727) );
  AND2_X1 U5668 ( .A1(b_9_), .A2(a_0_), .ZN(n5722) );
  OR2_X1 U5669 ( .A1(n5729), .A2(n5730), .ZN(n5723) );
  AND2_X1 U5670 ( .A1(n5713), .A2(n5712), .ZN(n5730) );
  AND2_X1 U5671 ( .A1(n5708), .A2(n5731), .ZN(n5729) );
  OR2_X1 U5672 ( .A1(n5712), .A2(n5713), .ZN(n5731) );
  OR2_X1 U5673 ( .A1(n3782), .A2(n4002), .ZN(n5713) );
  OR2_X1 U5674 ( .A1(n5732), .A2(n5733), .ZN(n5712) );
  AND2_X1 U5675 ( .A1(n5702), .A2(n5701), .ZN(n5733) );
  AND2_X1 U5676 ( .A1(n5697), .A2(n5734), .ZN(n5732) );
  OR2_X1 U5677 ( .A1(n5701), .A2(n5702), .ZN(n5734) );
  OR2_X1 U5678 ( .A1(n3782), .A2(n4035), .ZN(n5702) );
  OR2_X1 U5679 ( .A1(n5735), .A2(n5736), .ZN(n5701) );
  AND2_X1 U5680 ( .A1(n5691), .A2(n5690), .ZN(n5736) );
  AND2_X1 U5681 ( .A1(n5686), .A2(n5737), .ZN(n5735) );
  OR2_X1 U5682 ( .A1(n5690), .A2(n5691), .ZN(n5737) );
  OR2_X1 U5683 ( .A1(n3782), .A2(n3951), .ZN(n5691) );
  OR2_X1 U5684 ( .A1(n5738), .A2(n5739), .ZN(n5690) );
  AND2_X1 U5685 ( .A1(n5675), .A2(n5678), .ZN(n5739) );
  AND2_X1 U5686 ( .A1(n5740), .A2(n5680), .ZN(n5738) );
  OR2_X1 U5687 ( .A1(n5741), .A2(n5742), .ZN(n5680) );
  AND2_X1 U5688 ( .A1(n5669), .A2(n5668), .ZN(n5742) );
  AND2_X1 U5689 ( .A1(n5664), .A2(n5743), .ZN(n5741) );
  OR2_X1 U5690 ( .A1(n5668), .A2(n5669), .ZN(n5743) );
  OR2_X1 U5691 ( .A1(n3782), .A2(n3888), .ZN(n5669) );
  OR2_X1 U5692 ( .A1(n5744), .A2(n5745), .ZN(n5668) );
  AND2_X1 U5693 ( .A1(n5653), .A2(n5656), .ZN(n5745) );
  AND2_X1 U5694 ( .A1(n5746), .A2(n5658), .ZN(n5744) );
  OR2_X1 U5695 ( .A1(n5747), .A2(n5748), .ZN(n5658) );
  AND2_X1 U5696 ( .A1(n5642), .A2(n5645), .ZN(n5748) );
  AND2_X1 U5697 ( .A1(n5749), .A2(n5647), .ZN(n5747) );
  OR2_X1 U5698 ( .A1(n5750), .A2(n5751), .ZN(n5647) );
  AND2_X1 U5699 ( .A1(n5631), .A2(n5634), .ZN(n5751) );
  AND2_X1 U5700 ( .A1(n5752), .A2(n5636), .ZN(n5750) );
  OR2_X1 U5701 ( .A1(n5753), .A2(n5754), .ZN(n5636) );
  AND2_X1 U5702 ( .A1(n5622), .A2(n4057), .ZN(n5754) );
  AND2_X1 U5703 ( .A1(n5755), .A2(n5626), .ZN(n5753) );
  OR2_X1 U5704 ( .A1(n5756), .A2(n5757), .ZN(n5626) );
  AND2_X1 U5705 ( .A1(n5611), .A2(n5614), .ZN(n5757) );
  AND2_X1 U5706 ( .A1(n5758), .A2(n5617), .ZN(n5756) );
  OR2_X1 U5707 ( .A1(n5759), .A2(n5760), .ZN(n5617) );
  AND2_X1 U5708 ( .A1(n5600), .A2(n5603), .ZN(n5760) );
  AND2_X1 U5709 ( .A1(n5761), .A2(n5605), .ZN(n5759) );
  OR2_X1 U5710 ( .A1(n5762), .A2(n5763), .ZN(n5605) );
  AND2_X1 U5711 ( .A1(n5589), .A2(n5592), .ZN(n5763) );
  AND2_X1 U5712 ( .A1(n5764), .A2(n5594), .ZN(n5762) );
  OR2_X1 U5713 ( .A1(n5765), .A2(n5766), .ZN(n5594) );
  AND2_X1 U5714 ( .A1(n5577), .A2(n5583), .ZN(n5766) );
  AND2_X1 U5715 ( .A1(n5584), .A2(n5767), .ZN(n5765) );
  OR2_X1 U5716 ( .A1(n5583), .A2(n5577), .ZN(n5767) );
  OR2_X1 U5717 ( .A1(n3782), .A2(n3682), .ZN(n5577) );
  OR2_X1 U5718 ( .A1(n4070), .A2(n5768), .ZN(n5583) );
  OR2_X1 U5719 ( .A1(n4054), .A2(n3782), .ZN(n5768) );
  INV_X1 U5720 ( .A(n5582), .ZN(n5584) );
  OR2_X1 U5721 ( .A1(n5769), .A2(n5770), .ZN(n5582) );
  AND2_X1 U5722 ( .A1(b_8_), .A2(n5771), .ZN(n5770) );
  OR2_X1 U5723 ( .A1(n5772), .A2(n3644), .ZN(n5771) );
  AND2_X1 U5724 ( .A1(a_14_), .A2(n3833), .ZN(n5772) );
  AND2_X1 U5725 ( .A1(b_7_), .A2(n5773), .ZN(n5769) );
  OR2_X1 U5726 ( .A1(n5774), .A2(n3647), .ZN(n5773) );
  AND2_X1 U5727 ( .A1(a_15_), .A2(n4054), .ZN(n5774) );
  OR2_X1 U5728 ( .A1(n5592), .A2(n5589), .ZN(n5764) );
  OR2_X1 U5729 ( .A1(n5775), .A2(n5776), .ZN(n5589) );
  AND2_X1 U5730 ( .A1(n5777), .A2(n5778), .ZN(n5776) );
  INV_X1 U5731 ( .A(n5779), .ZN(n5775) );
  OR2_X1 U5732 ( .A1(n5777), .A2(n5778), .ZN(n5779) );
  OR2_X1 U5733 ( .A1(n5780), .A2(n5781), .ZN(n5777) );
  AND2_X1 U5734 ( .A1(n5782), .A2(n5783), .ZN(n5781) );
  INV_X1 U5735 ( .A(n5784), .ZN(n5782) );
  AND2_X1 U5736 ( .A1(n5785), .A2(n5784), .ZN(n5780) );
  OR2_X1 U5737 ( .A1(n3782), .A2(n4072), .ZN(n5592) );
  OR2_X1 U5738 ( .A1(n5603), .A2(n5600), .ZN(n5761) );
  OR2_X1 U5739 ( .A1(n5786), .A2(n5787), .ZN(n5600) );
  INV_X1 U5740 ( .A(n5788), .ZN(n5787) );
  OR2_X1 U5741 ( .A1(n5789), .A2(n5790), .ZN(n5788) );
  AND2_X1 U5742 ( .A1(n5790), .A2(n5789), .ZN(n5786) );
  AND2_X1 U5743 ( .A1(n5791), .A2(n5792), .ZN(n5789) );
  OR2_X1 U5744 ( .A1(n5793), .A2(n5794), .ZN(n5792) );
  INV_X1 U5745 ( .A(n5795), .ZN(n5794) );
  OR2_X1 U5746 ( .A1(n5795), .A2(n5796), .ZN(n5791) );
  INV_X1 U5747 ( .A(n5793), .ZN(n5796) );
  OR2_X1 U5748 ( .A1(n3782), .A2(n3735), .ZN(n5603) );
  OR2_X1 U5749 ( .A1(n5614), .A2(n5611), .ZN(n5758) );
  OR2_X1 U5750 ( .A1(n5797), .A2(n5798), .ZN(n5611) );
  INV_X1 U5751 ( .A(n5799), .ZN(n5798) );
  OR2_X1 U5752 ( .A1(n5800), .A2(n5801), .ZN(n5799) );
  AND2_X1 U5753 ( .A1(n5801), .A2(n5800), .ZN(n5797) );
  AND2_X1 U5754 ( .A1(n5802), .A2(n5803), .ZN(n5800) );
  OR2_X1 U5755 ( .A1(n5804), .A2(n5805), .ZN(n5803) );
  INV_X1 U5756 ( .A(n5806), .ZN(n5805) );
  OR2_X1 U5757 ( .A1(n5806), .A2(n5807), .ZN(n5802) );
  INV_X1 U5758 ( .A(n5804), .ZN(n5807) );
  OR2_X1 U5759 ( .A1(n3782), .A2(n4059), .ZN(n5614) );
  OR2_X1 U5760 ( .A1(n4057), .A2(n5622), .ZN(n5755) );
  OR2_X1 U5761 ( .A1(n5808), .A2(n5809), .ZN(n5622) );
  INV_X1 U5762 ( .A(n5810), .ZN(n5809) );
  OR2_X1 U5763 ( .A1(n5811), .A2(n5812), .ZN(n5810) );
  AND2_X1 U5764 ( .A1(n5812), .A2(n5811), .ZN(n5808) );
  AND2_X1 U5765 ( .A1(n5813), .A2(n5814), .ZN(n5811) );
  OR2_X1 U5766 ( .A1(n5815), .A2(n5816), .ZN(n5814) );
  INV_X1 U5767 ( .A(n5817), .ZN(n5813) );
  AND2_X1 U5768 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  INV_X1 U5769 ( .A(n5818), .ZN(n5816) );
  OR2_X1 U5770 ( .A1(n3782), .A2(n3786), .ZN(n4057) );
  OR2_X1 U5771 ( .A1(n5634), .A2(n5631), .ZN(n5752) );
  OR2_X1 U5772 ( .A1(n5819), .A2(n5820), .ZN(n5631) );
  INV_X1 U5773 ( .A(n5821), .ZN(n5820) );
  OR2_X1 U5774 ( .A1(n5822), .A2(n5823), .ZN(n5821) );
  AND2_X1 U5775 ( .A1(n5823), .A2(n5822), .ZN(n5819) );
  AND2_X1 U5776 ( .A1(n5824), .A2(n5825), .ZN(n5822) );
  OR2_X1 U5777 ( .A1(n5826), .A2(n5827), .ZN(n5825) );
  INV_X1 U5778 ( .A(n5828), .ZN(n5827) );
  OR2_X1 U5779 ( .A1(n5828), .A2(n5829), .ZN(n5824) );
  INV_X1 U5780 ( .A(n5826), .ZN(n5829) );
  OR2_X1 U5781 ( .A1(n3782), .A2(n4053), .ZN(n5634) );
  OR2_X1 U5782 ( .A1(n5645), .A2(n5642), .ZN(n5749) );
  OR2_X1 U5783 ( .A1(n5830), .A2(n5831), .ZN(n5642) );
  INV_X1 U5784 ( .A(n5832), .ZN(n5831) );
  OR2_X1 U5785 ( .A1(n5833), .A2(n5834), .ZN(n5832) );
  AND2_X1 U5786 ( .A1(n5834), .A2(n5833), .ZN(n5830) );
  AND2_X1 U5787 ( .A1(n5835), .A2(n5836), .ZN(n5833) );
  OR2_X1 U5788 ( .A1(n5837), .A2(n5838), .ZN(n5836) );
  INV_X1 U5789 ( .A(n5839), .ZN(n5835) );
  AND2_X1 U5790 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  OR2_X1 U5791 ( .A1(n3782), .A2(n3837), .ZN(n5645) );
  OR2_X1 U5792 ( .A1(n5656), .A2(n5653), .ZN(n5746) );
  OR2_X1 U5793 ( .A1(n5840), .A2(n5841), .ZN(n5653) );
  INV_X1 U5794 ( .A(n5842), .ZN(n5841) );
  OR2_X1 U5795 ( .A1(n5843), .A2(n5844), .ZN(n5842) );
  AND2_X1 U5796 ( .A1(n5844), .A2(n5843), .ZN(n5840) );
  AND2_X1 U5797 ( .A1(n5845), .A2(n5846), .ZN(n5843) );
  OR2_X1 U5798 ( .A1(n5847), .A2(n5848), .ZN(n5846) );
  INV_X1 U5799 ( .A(n5849), .ZN(n5848) );
  OR2_X1 U5800 ( .A1(n5849), .A2(n5850), .ZN(n5845) );
  INV_X1 U5801 ( .A(n5847), .ZN(n5850) );
  OR2_X1 U5802 ( .A1(n3782), .A2(n4047), .ZN(n5656) );
  AND2_X1 U5803 ( .A1(n5851), .A2(n5852), .ZN(n5664) );
  INV_X1 U5804 ( .A(n5853), .ZN(n5852) );
  AND2_X1 U5805 ( .A1(n5854), .A2(n5855), .ZN(n5853) );
  OR2_X1 U5806 ( .A1(n5855), .A2(n5854), .ZN(n5851) );
  OR2_X1 U5807 ( .A1(n5856), .A2(n5857), .ZN(n5854) );
  AND2_X1 U5808 ( .A1(n5858), .A2(n5859), .ZN(n5857) );
  INV_X1 U5809 ( .A(n5860), .ZN(n5858) );
  AND2_X1 U5810 ( .A1(n5861), .A2(n5860), .ZN(n5856) );
  INV_X1 U5811 ( .A(n5859), .ZN(n5861) );
  OR2_X1 U5812 ( .A1(n5678), .A2(n5675), .ZN(n5740) );
  OR2_X1 U5813 ( .A1(n5862), .A2(n5863), .ZN(n5675) );
  INV_X1 U5814 ( .A(n5864), .ZN(n5863) );
  OR2_X1 U5815 ( .A1(n5865), .A2(n5866), .ZN(n5864) );
  AND2_X1 U5816 ( .A1(n5866), .A2(n5865), .ZN(n5862) );
  AND2_X1 U5817 ( .A1(n5867), .A2(n5868), .ZN(n5865) );
  OR2_X1 U5818 ( .A1(n5869), .A2(n5870), .ZN(n5868) );
  INV_X1 U5819 ( .A(n5871), .ZN(n5870) );
  OR2_X1 U5820 ( .A1(n5871), .A2(n5872), .ZN(n5867) );
  INV_X1 U5821 ( .A(n5869), .ZN(n5872) );
  OR2_X1 U5822 ( .A1(n3782), .A2(n4041), .ZN(n5678) );
  INV_X1 U5823 ( .A(b_9_), .ZN(n3782) );
  AND2_X1 U5824 ( .A1(n5873), .A2(n5874), .ZN(n5686) );
  INV_X1 U5825 ( .A(n5875), .ZN(n5874) );
  AND2_X1 U5826 ( .A1(n5876), .A2(n5877), .ZN(n5875) );
  OR2_X1 U5827 ( .A1(n5877), .A2(n5876), .ZN(n5873) );
  OR2_X1 U5828 ( .A1(n5878), .A2(n5879), .ZN(n5876) );
  AND2_X1 U5829 ( .A1(n5880), .A2(n5881), .ZN(n5879) );
  INV_X1 U5830 ( .A(n5882), .ZN(n5880) );
  AND2_X1 U5831 ( .A1(n5883), .A2(n5882), .ZN(n5878) );
  INV_X1 U5832 ( .A(n5881), .ZN(n5883) );
  AND2_X1 U5833 ( .A1(n5884), .A2(n5885), .ZN(n5697) );
  INV_X1 U5834 ( .A(n5886), .ZN(n5885) );
  AND2_X1 U5835 ( .A1(n5887), .A2(n5888), .ZN(n5886) );
  OR2_X1 U5836 ( .A1(n5888), .A2(n5887), .ZN(n5884) );
  OR2_X1 U5837 ( .A1(n5889), .A2(n5890), .ZN(n5887) );
  AND2_X1 U5838 ( .A1(n5891), .A2(n5892), .ZN(n5890) );
  INV_X1 U5839 ( .A(n5893), .ZN(n5891) );
  AND2_X1 U5840 ( .A1(n5894), .A2(n5893), .ZN(n5889) );
  INV_X1 U5841 ( .A(n5892), .ZN(n5894) );
  AND2_X1 U5842 ( .A1(n5895), .A2(n5896), .ZN(n5708) );
  INV_X1 U5843 ( .A(n5897), .ZN(n5896) );
  AND2_X1 U5844 ( .A1(n5898), .A2(n5899), .ZN(n5897) );
  OR2_X1 U5845 ( .A1(n5899), .A2(n5898), .ZN(n5895) );
  OR2_X1 U5846 ( .A1(n5900), .A2(n5901), .ZN(n5898) );
  AND2_X1 U5847 ( .A1(n5902), .A2(n5903), .ZN(n5901) );
  INV_X1 U5848 ( .A(n5904), .ZN(n5902) );
  AND2_X1 U5849 ( .A1(n5905), .A2(n5904), .ZN(n5900) );
  INV_X1 U5850 ( .A(n5903), .ZN(n5905) );
  AND2_X1 U5851 ( .A1(n5906), .A2(n5907), .ZN(n5719) );
  INV_X1 U5852 ( .A(n5908), .ZN(n5907) );
  AND2_X1 U5853 ( .A1(n5909), .A2(n5910), .ZN(n5908) );
  OR2_X1 U5854 ( .A1(n5910), .A2(n5909), .ZN(n5906) );
  OR2_X1 U5855 ( .A1(n5911), .A2(n5912), .ZN(n5909) );
  AND2_X1 U5856 ( .A1(n5913), .A2(n5914), .ZN(n5912) );
  INV_X1 U5857 ( .A(n5915), .ZN(n5913) );
  AND2_X1 U5858 ( .A1(n5916), .A2(n5915), .ZN(n5911) );
  INV_X1 U5859 ( .A(n5914), .ZN(n5916) );
  AND2_X1 U5860 ( .A1(n5917), .A2(n5918), .ZN(n4489) );
  OR2_X1 U5861 ( .A1(n5919), .A2(n4405), .ZN(n5918) );
  INV_X1 U5862 ( .A(n5920), .ZN(n5919) );
  OR2_X1 U5863 ( .A1(n5921), .A2(n5920), .ZN(n5917) );
  AND2_X1 U5864 ( .A1(n5922), .A2(n5923), .ZN(n5920) );
  OR2_X1 U5865 ( .A1(n4403), .A2(n5924), .ZN(n5923) );
  INV_X1 U5866 ( .A(n5925), .ZN(n5922) );
  AND2_X1 U5867 ( .A1(n5924), .A2(n4403), .ZN(n5925) );
  OR2_X1 U5868 ( .A1(n4054), .A2(n4028), .ZN(n4403) );
  INV_X1 U5869 ( .A(n4404), .ZN(n5924) );
  OR2_X1 U5870 ( .A1(n5926), .A2(n5927), .ZN(n4404) );
  AND2_X1 U5871 ( .A1(n5915), .A2(n5914), .ZN(n5927) );
  AND2_X1 U5872 ( .A1(n5910), .A2(n5928), .ZN(n5926) );
  OR2_X1 U5873 ( .A1(n5914), .A2(n5915), .ZN(n5928) );
  OR2_X1 U5874 ( .A1(n4054), .A2(n4002), .ZN(n5915) );
  OR2_X1 U5875 ( .A1(n5929), .A2(n5930), .ZN(n5914) );
  AND2_X1 U5876 ( .A1(n5904), .A2(n5903), .ZN(n5930) );
  AND2_X1 U5877 ( .A1(n5899), .A2(n5931), .ZN(n5929) );
  OR2_X1 U5878 ( .A1(n5903), .A2(n5904), .ZN(n5931) );
  OR2_X1 U5879 ( .A1(n4054), .A2(n4035), .ZN(n5904) );
  OR2_X1 U5880 ( .A1(n5932), .A2(n5933), .ZN(n5903) );
  AND2_X1 U5881 ( .A1(n5893), .A2(n5892), .ZN(n5933) );
  AND2_X1 U5882 ( .A1(n5888), .A2(n5934), .ZN(n5932) );
  OR2_X1 U5883 ( .A1(n5892), .A2(n5893), .ZN(n5934) );
  OR2_X1 U5884 ( .A1(n4054), .A2(n3951), .ZN(n5893) );
  OR2_X1 U5885 ( .A1(n5935), .A2(n5936), .ZN(n5892) );
  AND2_X1 U5886 ( .A1(n5882), .A2(n5881), .ZN(n5936) );
  AND2_X1 U5887 ( .A1(n5877), .A2(n5937), .ZN(n5935) );
  OR2_X1 U5888 ( .A1(n5881), .A2(n5882), .ZN(n5937) );
  OR2_X1 U5889 ( .A1(n4054), .A2(n4041), .ZN(n5882) );
  OR2_X1 U5890 ( .A1(n5938), .A2(n5939), .ZN(n5881) );
  AND2_X1 U5891 ( .A1(n5866), .A2(n5869), .ZN(n5939) );
  AND2_X1 U5892 ( .A1(n5940), .A2(n5871), .ZN(n5938) );
  OR2_X1 U5893 ( .A1(n5941), .A2(n5942), .ZN(n5871) );
  AND2_X1 U5894 ( .A1(n5860), .A2(n5859), .ZN(n5942) );
  AND2_X1 U5895 ( .A1(n5855), .A2(n5943), .ZN(n5941) );
  OR2_X1 U5896 ( .A1(n5859), .A2(n5860), .ZN(n5943) );
  OR2_X1 U5897 ( .A1(n4054), .A2(n4047), .ZN(n5860) );
  OR2_X1 U5898 ( .A1(n5944), .A2(n5945), .ZN(n5859) );
  AND2_X1 U5899 ( .A1(n5844), .A2(n5847), .ZN(n5945) );
  AND2_X1 U5900 ( .A1(n5946), .A2(n5849), .ZN(n5944) );
  OR2_X1 U5901 ( .A1(n5947), .A2(n5948), .ZN(n5849) );
  AND2_X1 U5902 ( .A1(n5834), .A2(n3811), .ZN(n5948) );
  AND2_X1 U5903 ( .A1(n5949), .A2(n5837), .ZN(n5947) );
  OR2_X1 U5904 ( .A1(n5950), .A2(n5951), .ZN(n5837) );
  AND2_X1 U5905 ( .A1(n5823), .A2(n5826), .ZN(n5951) );
  AND2_X1 U5906 ( .A1(n5952), .A2(n5828), .ZN(n5950) );
  OR2_X1 U5907 ( .A1(n5953), .A2(n5954), .ZN(n5828) );
  AND2_X1 U5908 ( .A1(n5812), .A2(n5815), .ZN(n5954) );
  AND2_X1 U5909 ( .A1(n5955), .A2(n5818), .ZN(n5953) );
  OR2_X1 U5910 ( .A1(n5956), .A2(n5957), .ZN(n5818) );
  AND2_X1 U5911 ( .A1(n5801), .A2(n5804), .ZN(n5957) );
  AND2_X1 U5912 ( .A1(n5958), .A2(n5806), .ZN(n5956) );
  OR2_X1 U5913 ( .A1(n5959), .A2(n5960), .ZN(n5806) );
  AND2_X1 U5914 ( .A1(n5790), .A2(n5793), .ZN(n5960) );
  AND2_X1 U5915 ( .A1(n5961), .A2(n5795), .ZN(n5959) );
  OR2_X1 U5916 ( .A1(n5962), .A2(n5963), .ZN(n5795) );
  AND2_X1 U5917 ( .A1(n5778), .A2(n5784), .ZN(n5963) );
  AND2_X1 U5918 ( .A1(n5785), .A2(n5964), .ZN(n5962) );
  OR2_X1 U5919 ( .A1(n5784), .A2(n5778), .ZN(n5964) );
  OR2_X1 U5920 ( .A1(n4054), .A2(n3682), .ZN(n5778) );
  OR2_X1 U5921 ( .A1(n3833), .A2(n5965), .ZN(n5784) );
  OR2_X1 U5922 ( .A1(n4054), .A2(n4070), .ZN(n5965) );
  INV_X1 U5923 ( .A(n5783), .ZN(n5785) );
  OR2_X1 U5924 ( .A1(n5966), .A2(n5967), .ZN(n5783) );
  AND2_X1 U5925 ( .A1(b_7_), .A2(n5968), .ZN(n5967) );
  OR2_X1 U5926 ( .A1(n5969), .A2(n3644), .ZN(n5968) );
  AND2_X1 U5927 ( .A1(a_14_), .A2(n4048), .ZN(n5969) );
  AND2_X1 U5928 ( .A1(b_6_), .A2(n5970), .ZN(n5966) );
  OR2_X1 U5929 ( .A1(n5971), .A2(n3647), .ZN(n5970) );
  AND2_X1 U5930 ( .A1(a_15_), .A2(n3833), .ZN(n5971) );
  OR2_X1 U5931 ( .A1(n5793), .A2(n5790), .ZN(n5961) );
  OR2_X1 U5932 ( .A1(n5972), .A2(n5973), .ZN(n5790) );
  AND2_X1 U5933 ( .A1(n5974), .A2(n5975), .ZN(n5973) );
  INV_X1 U5934 ( .A(n5976), .ZN(n5972) );
  OR2_X1 U5935 ( .A1(n5974), .A2(n5975), .ZN(n5976) );
  OR2_X1 U5936 ( .A1(n5977), .A2(n5978), .ZN(n5974) );
  AND2_X1 U5937 ( .A1(n5979), .A2(n5980), .ZN(n5978) );
  INV_X1 U5938 ( .A(n5981), .ZN(n5979) );
  AND2_X1 U5939 ( .A1(n5982), .A2(n5981), .ZN(n5977) );
  OR2_X1 U5940 ( .A1(n4054), .A2(n4072), .ZN(n5793) );
  OR2_X1 U5941 ( .A1(n5804), .A2(n5801), .ZN(n5958) );
  OR2_X1 U5942 ( .A1(n5983), .A2(n5984), .ZN(n5801) );
  INV_X1 U5943 ( .A(n5985), .ZN(n5984) );
  OR2_X1 U5944 ( .A1(n5986), .A2(n5987), .ZN(n5985) );
  AND2_X1 U5945 ( .A1(n5987), .A2(n5986), .ZN(n5983) );
  AND2_X1 U5946 ( .A1(n5988), .A2(n5989), .ZN(n5986) );
  OR2_X1 U5947 ( .A1(n5990), .A2(n5991), .ZN(n5989) );
  INV_X1 U5948 ( .A(n5992), .ZN(n5991) );
  OR2_X1 U5949 ( .A1(n5992), .A2(n5993), .ZN(n5988) );
  INV_X1 U5950 ( .A(n5990), .ZN(n5993) );
  OR2_X1 U5951 ( .A1(n4054), .A2(n3735), .ZN(n5804) );
  OR2_X1 U5952 ( .A1(n5815), .A2(n5812), .ZN(n5955) );
  OR2_X1 U5953 ( .A1(n5994), .A2(n5995), .ZN(n5812) );
  INV_X1 U5954 ( .A(n5996), .ZN(n5995) );
  OR2_X1 U5955 ( .A1(n5997), .A2(n5998), .ZN(n5996) );
  AND2_X1 U5956 ( .A1(n5998), .A2(n5997), .ZN(n5994) );
  AND2_X1 U5957 ( .A1(n5999), .A2(n6000), .ZN(n5997) );
  OR2_X1 U5958 ( .A1(n6001), .A2(n6002), .ZN(n6000) );
  INV_X1 U5959 ( .A(n6003), .ZN(n6002) );
  OR2_X1 U5960 ( .A1(n6003), .A2(n6004), .ZN(n5999) );
  INV_X1 U5961 ( .A(n6001), .ZN(n6004) );
  OR2_X1 U5962 ( .A1(n4054), .A2(n4059), .ZN(n5815) );
  OR2_X1 U5963 ( .A1(n5826), .A2(n5823), .ZN(n5952) );
  OR2_X1 U5964 ( .A1(n6005), .A2(n6006), .ZN(n5823) );
  INV_X1 U5965 ( .A(n6007), .ZN(n6006) );
  OR2_X1 U5966 ( .A1(n6008), .A2(n6009), .ZN(n6007) );
  AND2_X1 U5967 ( .A1(n6009), .A2(n6008), .ZN(n6005) );
  AND2_X1 U5968 ( .A1(n6010), .A2(n6011), .ZN(n6008) );
  OR2_X1 U5969 ( .A1(n6012), .A2(n6013), .ZN(n6011) );
  INV_X1 U5970 ( .A(n6014), .ZN(n6010) );
  AND2_X1 U5971 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  INV_X1 U5972 ( .A(n6015), .ZN(n6013) );
  OR2_X1 U5973 ( .A1(n4054), .A2(n3786), .ZN(n5826) );
  OR2_X1 U5974 ( .A1(n3811), .A2(n5834), .ZN(n5949) );
  OR2_X1 U5975 ( .A1(n6016), .A2(n6017), .ZN(n5834) );
  INV_X1 U5976 ( .A(n6018), .ZN(n6017) );
  OR2_X1 U5977 ( .A1(n6019), .A2(n6020), .ZN(n6018) );
  AND2_X1 U5978 ( .A1(n6020), .A2(n6019), .ZN(n6016) );
  AND2_X1 U5979 ( .A1(n6021), .A2(n6022), .ZN(n6019) );
  OR2_X1 U5980 ( .A1(n6023), .A2(n6024), .ZN(n6022) );
  INV_X1 U5981 ( .A(n6025), .ZN(n6024) );
  OR2_X1 U5982 ( .A1(n6025), .A2(n6026), .ZN(n6021) );
  INV_X1 U5983 ( .A(n6023), .ZN(n6026) );
  INV_X1 U5984 ( .A(n5838), .ZN(n3811) );
  AND2_X1 U5985 ( .A1(b_8_), .A2(a_8_), .ZN(n5838) );
  OR2_X1 U5986 ( .A1(n5847), .A2(n5844), .ZN(n5946) );
  OR2_X1 U5987 ( .A1(n6027), .A2(n6028), .ZN(n5844) );
  INV_X1 U5988 ( .A(n6029), .ZN(n6028) );
  OR2_X1 U5989 ( .A1(n6030), .A2(n6031), .ZN(n6029) );
  AND2_X1 U5990 ( .A1(n6031), .A2(n6030), .ZN(n6027) );
  AND2_X1 U5991 ( .A1(n6032), .A2(n6033), .ZN(n6030) );
  OR2_X1 U5992 ( .A1(n6034), .A2(n6035), .ZN(n6033) );
  INV_X1 U5993 ( .A(n6036), .ZN(n6035) );
  OR2_X1 U5994 ( .A1(n6036), .A2(n6037), .ZN(n6032) );
  INV_X1 U5995 ( .A(n6034), .ZN(n6037) );
  OR2_X1 U5996 ( .A1(n4054), .A2(n3837), .ZN(n5847) );
  AND2_X1 U5997 ( .A1(n6038), .A2(n6039), .ZN(n5855) );
  INV_X1 U5998 ( .A(n6040), .ZN(n6039) );
  AND2_X1 U5999 ( .A1(n6041), .A2(n6042), .ZN(n6040) );
  OR2_X1 U6000 ( .A1(n6042), .A2(n6041), .ZN(n6038) );
  OR2_X1 U6001 ( .A1(n6043), .A2(n6044), .ZN(n6041) );
  AND2_X1 U6002 ( .A1(n3840), .A2(n6045), .ZN(n6044) );
  INV_X1 U6003 ( .A(n4051), .ZN(n3840) );
  AND2_X1 U6004 ( .A1(n6046), .A2(n4051), .ZN(n6043) );
  INV_X1 U6005 ( .A(n6045), .ZN(n6046) );
  OR2_X1 U6006 ( .A1(n5869), .A2(n5866), .ZN(n5940) );
  OR2_X1 U6007 ( .A1(n6047), .A2(n6048), .ZN(n5866) );
  INV_X1 U6008 ( .A(n6049), .ZN(n6048) );
  OR2_X1 U6009 ( .A1(n6050), .A2(n6051), .ZN(n6049) );
  AND2_X1 U6010 ( .A1(n6051), .A2(n6050), .ZN(n6047) );
  AND2_X1 U6011 ( .A1(n6052), .A2(n6053), .ZN(n6050) );
  OR2_X1 U6012 ( .A1(n6054), .A2(n6055), .ZN(n6053) );
  INV_X1 U6013 ( .A(n6056), .ZN(n6055) );
  OR2_X1 U6014 ( .A1(n6056), .A2(n6057), .ZN(n6052) );
  INV_X1 U6015 ( .A(n6054), .ZN(n6057) );
  OR2_X1 U6016 ( .A1(n4054), .A2(n3888), .ZN(n5869) );
  INV_X1 U6017 ( .A(b_8_), .ZN(n4054) );
  AND2_X1 U6018 ( .A1(n6058), .A2(n6059), .ZN(n5877) );
  INV_X1 U6019 ( .A(n6060), .ZN(n6059) );
  AND2_X1 U6020 ( .A1(n6061), .A2(n6062), .ZN(n6060) );
  OR2_X1 U6021 ( .A1(n6062), .A2(n6061), .ZN(n6058) );
  OR2_X1 U6022 ( .A1(n6063), .A2(n6064), .ZN(n6061) );
  AND2_X1 U6023 ( .A1(n6065), .A2(n6066), .ZN(n6064) );
  INV_X1 U6024 ( .A(n6067), .ZN(n6065) );
  AND2_X1 U6025 ( .A1(n6068), .A2(n6067), .ZN(n6063) );
  INV_X1 U6026 ( .A(n6066), .ZN(n6068) );
  AND2_X1 U6027 ( .A1(n6069), .A2(n6070), .ZN(n5888) );
  INV_X1 U6028 ( .A(n6071), .ZN(n6070) );
  AND2_X1 U6029 ( .A1(n6072), .A2(n6073), .ZN(n6071) );
  OR2_X1 U6030 ( .A1(n6073), .A2(n6072), .ZN(n6069) );
  OR2_X1 U6031 ( .A1(n6074), .A2(n6075), .ZN(n6072) );
  AND2_X1 U6032 ( .A1(n6076), .A2(n6077), .ZN(n6075) );
  INV_X1 U6033 ( .A(n6078), .ZN(n6076) );
  AND2_X1 U6034 ( .A1(n6079), .A2(n6078), .ZN(n6074) );
  INV_X1 U6035 ( .A(n6077), .ZN(n6079) );
  AND2_X1 U6036 ( .A1(n6080), .A2(n6081), .ZN(n5899) );
  INV_X1 U6037 ( .A(n6082), .ZN(n6081) );
  AND2_X1 U6038 ( .A1(n6083), .A2(n6084), .ZN(n6082) );
  OR2_X1 U6039 ( .A1(n6084), .A2(n6083), .ZN(n6080) );
  OR2_X1 U6040 ( .A1(n6085), .A2(n6086), .ZN(n6083) );
  AND2_X1 U6041 ( .A1(n6087), .A2(n6088), .ZN(n6086) );
  INV_X1 U6042 ( .A(n6089), .ZN(n6087) );
  AND2_X1 U6043 ( .A1(n6090), .A2(n6089), .ZN(n6085) );
  INV_X1 U6044 ( .A(n6088), .ZN(n6090) );
  AND2_X1 U6045 ( .A1(n6091), .A2(n6092), .ZN(n5910) );
  INV_X1 U6046 ( .A(n6093), .ZN(n6092) );
  AND2_X1 U6047 ( .A1(n6094), .A2(n6095), .ZN(n6093) );
  OR2_X1 U6048 ( .A1(n6095), .A2(n6094), .ZN(n6091) );
  OR2_X1 U6049 ( .A1(n6096), .A2(n6097), .ZN(n6094) );
  AND2_X1 U6050 ( .A1(n6098), .A2(n6099), .ZN(n6097) );
  INV_X1 U6051 ( .A(n6100), .ZN(n6098) );
  AND2_X1 U6052 ( .A1(n6101), .A2(n6100), .ZN(n6096) );
  INV_X1 U6053 ( .A(n6099), .ZN(n6101) );
  INV_X1 U6054 ( .A(n4405), .ZN(n5921) );
  AND2_X1 U6055 ( .A1(n6102), .A2(n6103), .ZN(n4405) );
  INV_X1 U6056 ( .A(n6104), .ZN(n6103) );
  AND2_X1 U6057 ( .A1(n6105), .A2(n4418), .ZN(n6104) );
  OR2_X1 U6058 ( .A1(n4418), .A2(n6105), .ZN(n6102) );
  OR2_X1 U6059 ( .A1(n6106), .A2(n6107), .ZN(n6105) );
  AND2_X1 U6060 ( .A1(n6108), .A2(n4417), .ZN(n6107) );
  INV_X1 U6061 ( .A(n4416), .ZN(n6108) );
  AND2_X1 U6062 ( .A1(n6109), .A2(n4416), .ZN(n6106) );
  OR2_X1 U6063 ( .A1(n3833), .A2(n4002), .ZN(n4416) );
  INV_X1 U6064 ( .A(n4417), .ZN(n6109) );
  OR2_X1 U6065 ( .A1(n6110), .A2(n6111), .ZN(n4417) );
  AND2_X1 U6066 ( .A1(n6100), .A2(n6099), .ZN(n6111) );
  AND2_X1 U6067 ( .A1(n6095), .A2(n6112), .ZN(n6110) );
  OR2_X1 U6068 ( .A1(n6099), .A2(n6100), .ZN(n6112) );
  OR2_X1 U6069 ( .A1(n3833), .A2(n4035), .ZN(n6100) );
  OR2_X1 U6070 ( .A1(n6113), .A2(n6114), .ZN(n6099) );
  AND2_X1 U6071 ( .A1(n6089), .A2(n6088), .ZN(n6114) );
  AND2_X1 U6072 ( .A1(n6084), .A2(n6115), .ZN(n6113) );
  OR2_X1 U6073 ( .A1(n6088), .A2(n6089), .ZN(n6115) );
  OR2_X1 U6074 ( .A1(n3833), .A2(n3951), .ZN(n6089) );
  OR2_X1 U6075 ( .A1(n6116), .A2(n6117), .ZN(n6088) );
  AND2_X1 U6076 ( .A1(n6078), .A2(n6077), .ZN(n6117) );
  AND2_X1 U6077 ( .A1(n6073), .A2(n6118), .ZN(n6116) );
  OR2_X1 U6078 ( .A1(n6077), .A2(n6078), .ZN(n6118) );
  OR2_X1 U6079 ( .A1(n3833), .A2(n4041), .ZN(n6078) );
  OR2_X1 U6080 ( .A1(n6119), .A2(n6120), .ZN(n6077) );
  AND2_X1 U6081 ( .A1(n6067), .A2(n6066), .ZN(n6120) );
  AND2_X1 U6082 ( .A1(n6062), .A2(n6121), .ZN(n6119) );
  OR2_X1 U6083 ( .A1(n6066), .A2(n6067), .ZN(n6121) );
  OR2_X1 U6084 ( .A1(n3833), .A2(n3888), .ZN(n6067) );
  OR2_X1 U6085 ( .A1(n6122), .A2(n6123), .ZN(n6066) );
  AND2_X1 U6086 ( .A1(n6051), .A2(n6054), .ZN(n6123) );
  AND2_X1 U6087 ( .A1(n6124), .A2(n6056), .ZN(n6122) );
  OR2_X1 U6088 ( .A1(n6125), .A2(n6126), .ZN(n6056) );
  AND2_X1 U6089 ( .A1(n4051), .A2(n6045), .ZN(n6126) );
  AND2_X1 U6090 ( .A1(n6042), .A2(n6127), .ZN(n6125) );
  OR2_X1 U6091 ( .A1(n6045), .A2(n4051), .ZN(n6127) );
  OR2_X1 U6092 ( .A1(n3833), .A2(n3837), .ZN(n4051) );
  OR2_X1 U6093 ( .A1(n6128), .A2(n6129), .ZN(n6045) );
  AND2_X1 U6094 ( .A1(n6031), .A2(n6034), .ZN(n6129) );
  AND2_X1 U6095 ( .A1(n6130), .A2(n6036), .ZN(n6128) );
  OR2_X1 U6096 ( .A1(n6131), .A2(n6132), .ZN(n6036) );
  AND2_X1 U6097 ( .A1(n6020), .A2(n6023), .ZN(n6132) );
  AND2_X1 U6098 ( .A1(n6133), .A2(n6025), .ZN(n6131) );
  OR2_X1 U6099 ( .A1(n6134), .A2(n6135), .ZN(n6025) );
  AND2_X1 U6100 ( .A1(n6009), .A2(n6012), .ZN(n6135) );
  AND2_X1 U6101 ( .A1(n6136), .A2(n6015), .ZN(n6134) );
  OR2_X1 U6102 ( .A1(n6137), .A2(n6138), .ZN(n6015) );
  AND2_X1 U6103 ( .A1(n5998), .A2(n6001), .ZN(n6138) );
  AND2_X1 U6104 ( .A1(n6139), .A2(n6003), .ZN(n6137) );
  OR2_X1 U6105 ( .A1(n6140), .A2(n6141), .ZN(n6003) );
  AND2_X1 U6106 ( .A1(n5987), .A2(n5990), .ZN(n6141) );
  AND2_X1 U6107 ( .A1(n6142), .A2(n5992), .ZN(n6140) );
  OR2_X1 U6108 ( .A1(n6143), .A2(n6144), .ZN(n5992) );
  AND2_X1 U6109 ( .A1(n5975), .A2(n5981), .ZN(n6144) );
  AND2_X1 U6110 ( .A1(n5982), .A2(n6145), .ZN(n6143) );
  OR2_X1 U6111 ( .A1(n5981), .A2(n5975), .ZN(n6145) );
  OR2_X1 U6112 ( .A1(n3682), .A2(n3833), .ZN(n5975) );
  OR2_X1 U6113 ( .A1(n4048), .A2(n6146), .ZN(n5981) );
  OR2_X1 U6114 ( .A1(n4070), .A2(n3833), .ZN(n6146) );
  INV_X1 U6115 ( .A(n5980), .ZN(n5982) );
  OR2_X1 U6116 ( .A1(n6147), .A2(n6148), .ZN(n5980) );
  AND2_X1 U6117 ( .A1(b_6_), .A2(n6149), .ZN(n6148) );
  OR2_X1 U6118 ( .A1(n6150), .A2(n3644), .ZN(n6149) );
  AND2_X1 U6119 ( .A1(a_14_), .A2(n3884), .ZN(n6150) );
  AND2_X1 U6120 ( .A1(b_5_), .A2(n6151), .ZN(n6147) );
  OR2_X1 U6121 ( .A1(n6152), .A2(n3647), .ZN(n6151) );
  AND2_X1 U6122 ( .A1(a_15_), .A2(n4048), .ZN(n6152) );
  OR2_X1 U6123 ( .A1(n5990), .A2(n5987), .ZN(n6142) );
  OR2_X1 U6124 ( .A1(n6153), .A2(n6154), .ZN(n5987) );
  AND2_X1 U6125 ( .A1(n6155), .A2(n6156), .ZN(n6154) );
  INV_X1 U6126 ( .A(n6157), .ZN(n6153) );
  OR2_X1 U6127 ( .A1(n6155), .A2(n6156), .ZN(n6157) );
  OR2_X1 U6128 ( .A1(n6158), .A2(n6159), .ZN(n6155) );
  AND2_X1 U6129 ( .A1(n6160), .A2(n6161), .ZN(n6159) );
  INV_X1 U6130 ( .A(n6162), .ZN(n6160) );
  AND2_X1 U6131 ( .A1(n6163), .A2(n6162), .ZN(n6158) );
  OR2_X1 U6132 ( .A1(n4072), .A2(n3833), .ZN(n5990) );
  OR2_X1 U6133 ( .A1(n6001), .A2(n5998), .ZN(n6139) );
  OR2_X1 U6134 ( .A1(n6164), .A2(n6165), .ZN(n5998) );
  INV_X1 U6135 ( .A(n6166), .ZN(n6165) );
  OR2_X1 U6136 ( .A1(n6167), .A2(n6168), .ZN(n6166) );
  AND2_X1 U6137 ( .A1(n6168), .A2(n6167), .ZN(n6164) );
  AND2_X1 U6138 ( .A1(n6169), .A2(n6170), .ZN(n6167) );
  OR2_X1 U6139 ( .A1(n6171), .A2(n6172), .ZN(n6170) );
  INV_X1 U6140 ( .A(n6173), .ZN(n6172) );
  OR2_X1 U6141 ( .A1(n6173), .A2(n6174), .ZN(n6169) );
  INV_X1 U6142 ( .A(n6171), .ZN(n6174) );
  OR2_X1 U6143 ( .A1(n3833), .A2(n3735), .ZN(n6001) );
  OR2_X1 U6144 ( .A1(n6012), .A2(n6009), .ZN(n6136) );
  OR2_X1 U6145 ( .A1(n6175), .A2(n6176), .ZN(n6009) );
  INV_X1 U6146 ( .A(n6177), .ZN(n6176) );
  OR2_X1 U6147 ( .A1(n6178), .A2(n6179), .ZN(n6177) );
  AND2_X1 U6148 ( .A1(n6179), .A2(n6178), .ZN(n6175) );
  AND2_X1 U6149 ( .A1(n6180), .A2(n6181), .ZN(n6178) );
  OR2_X1 U6150 ( .A1(n6182), .A2(n6183), .ZN(n6181) );
  INV_X1 U6151 ( .A(n6184), .ZN(n6183) );
  OR2_X1 U6152 ( .A1(n6184), .A2(n6185), .ZN(n6180) );
  INV_X1 U6153 ( .A(n6182), .ZN(n6185) );
  OR2_X1 U6154 ( .A1(n3833), .A2(n4059), .ZN(n6012) );
  OR2_X1 U6155 ( .A1(n6023), .A2(n6020), .ZN(n6133) );
  OR2_X1 U6156 ( .A1(n6186), .A2(n6187), .ZN(n6020) );
  INV_X1 U6157 ( .A(n6188), .ZN(n6187) );
  OR2_X1 U6158 ( .A1(n6189), .A2(n6190), .ZN(n6188) );
  AND2_X1 U6159 ( .A1(n6190), .A2(n6189), .ZN(n6186) );
  AND2_X1 U6160 ( .A1(n6191), .A2(n6192), .ZN(n6189) );
  OR2_X1 U6161 ( .A1(n6193), .A2(n6194), .ZN(n6192) );
  INV_X1 U6162 ( .A(n6195), .ZN(n6191) );
  AND2_X1 U6163 ( .A1(n6194), .A2(n6193), .ZN(n6195) );
  INV_X1 U6164 ( .A(n6196), .ZN(n6194) );
  OR2_X1 U6165 ( .A1(n3833), .A2(n3786), .ZN(n6023) );
  OR2_X1 U6166 ( .A1(n6034), .A2(n6031), .ZN(n6130) );
  OR2_X1 U6167 ( .A1(n6197), .A2(n6198), .ZN(n6031) );
  INV_X1 U6168 ( .A(n6199), .ZN(n6198) );
  OR2_X1 U6169 ( .A1(n6200), .A2(n6201), .ZN(n6199) );
  AND2_X1 U6170 ( .A1(n6201), .A2(n6200), .ZN(n6197) );
  AND2_X1 U6171 ( .A1(n6202), .A2(n6203), .ZN(n6200) );
  OR2_X1 U6172 ( .A1(n6204), .A2(n6205), .ZN(n6203) );
  INV_X1 U6173 ( .A(n6206), .ZN(n6205) );
  OR2_X1 U6174 ( .A1(n6206), .A2(n6207), .ZN(n6202) );
  INV_X1 U6175 ( .A(n6204), .ZN(n6207) );
  OR2_X1 U6176 ( .A1(n3833), .A2(n4053), .ZN(n6034) );
  AND2_X1 U6177 ( .A1(n6208), .A2(n6209), .ZN(n6042) );
  INV_X1 U6178 ( .A(n6210), .ZN(n6209) );
  AND2_X1 U6179 ( .A1(n6211), .A2(n6212), .ZN(n6210) );
  OR2_X1 U6180 ( .A1(n6212), .A2(n6211), .ZN(n6208) );
  OR2_X1 U6181 ( .A1(n6213), .A2(n6214), .ZN(n6211) );
  AND2_X1 U6182 ( .A1(n6215), .A2(n6216), .ZN(n6214) );
  INV_X1 U6183 ( .A(n6217), .ZN(n6215) );
  AND2_X1 U6184 ( .A1(n6218), .A2(n6217), .ZN(n6213) );
  INV_X1 U6185 ( .A(n6216), .ZN(n6218) );
  OR2_X1 U6186 ( .A1(n6054), .A2(n6051), .ZN(n6124) );
  OR2_X1 U6187 ( .A1(n6219), .A2(n6220), .ZN(n6051) );
  INV_X1 U6188 ( .A(n6221), .ZN(n6220) );
  OR2_X1 U6189 ( .A1(n6222), .A2(n6223), .ZN(n6221) );
  AND2_X1 U6190 ( .A1(n6223), .A2(n6222), .ZN(n6219) );
  AND2_X1 U6191 ( .A1(n6224), .A2(n6225), .ZN(n6222) );
  OR2_X1 U6192 ( .A1(n6226), .A2(n6227), .ZN(n6225) );
  INV_X1 U6193 ( .A(n6228), .ZN(n6227) );
  OR2_X1 U6194 ( .A1(n6228), .A2(n6229), .ZN(n6224) );
  INV_X1 U6195 ( .A(n6226), .ZN(n6229) );
  OR2_X1 U6196 ( .A1(n3833), .A2(n4047), .ZN(n6054) );
  INV_X1 U6197 ( .A(b_7_), .ZN(n3833) );
  AND2_X1 U6198 ( .A1(n6230), .A2(n6231), .ZN(n6062) );
  INV_X1 U6199 ( .A(n6232), .ZN(n6231) );
  AND2_X1 U6200 ( .A1(n6233), .A2(n6234), .ZN(n6232) );
  OR2_X1 U6201 ( .A1(n6234), .A2(n6233), .ZN(n6230) );
  OR2_X1 U6202 ( .A1(n6235), .A2(n6236), .ZN(n6233) );
  AND2_X1 U6203 ( .A1(n6237), .A2(n6238), .ZN(n6236) );
  INV_X1 U6204 ( .A(n6239), .ZN(n6235) );
  OR2_X1 U6205 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  AND2_X1 U6206 ( .A1(n6240), .A2(n6241), .ZN(n6073) );
  INV_X1 U6207 ( .A(n6242), .ZN(n6241) );
  AND2_X1 U6208 ( .A1(n6243), .A2(n6244), .ZN(n6242) );
  OR2_X1 U6209 ( .A1(n6244), .A2(n6243), .ZN(n6240) );
  OR2_X1 U6210 ( .A1(n6245), .A2(n6246), .ZN(n6243) );
  AND2_X1 U6211 ( .A1(n6247), .A2(n6248), .ZN(n6246) );
  INV_X1 U6212 ( .A(n6249), .ZN(n6247) );
  AND2_X1 U6213 ( .A1(n6250), .A2(n6249), .ZN(n6245) );
  INV_X1 U6214 ( .A(n6248), .ZN(n6250) );
  AND2_X1 U6215 ( .A1(n6251), .A2(n6252), .ZN(n6084) );
  INV_X1 U6216 ( .A(n6253), .ZN(n6252) );
  AND2_X1 U6217 ( .A1(n6254), .A2(n6255), .ZN(n6253) );
  OR2_X1 U6218 ( .A1(n6255), .A2(n6254), .ZN(n6251) );
  OR2_X1 U6219 ( .A1(n6256), .A2(n6257), .ZN(n6254) );
  AND2_X1 U6220 ( .A1(n6258), .A2(n6259), .ZN(n6257) );
  INV_X1 U6221 ( .A(n6260), .ZN(n6258) );
  AND2_X1 U6222 ( .A1(n6261), .A2(n6260), .ZN(n6256) );
  INV_X1 U6223 ( .A(n6259), .ZN(n6261) );
  AND2_X1 U6224 ( .A1(n6262), .A2(n6263), .ZN(n6095) );
  INV_X1 U6225 ( .A(n6264), .ZN(n6263) );
  AND2_X1 U6226 ( .A1(n6265), .A2(n6266), .ZN(n6264) );
  OR2_X1 U6227 ( .A1(n6266), .A2(n6265), .ZN(n6262) );
  OR2_X1 U6228 ( .A1(n6267), .A2(n6268), .ZN(n6265) );
  AND2_X1 U6229 ( .A1(n6269), .A2(n6270), .ZN(n6268) );
  INV_X1 U6230 ( .A(n6271), .ZN(n6269) );
  AND2_X1 U6231 ( .A1(n6272), .A2(n6271), .ZN(n6267) );
  INV_X1 U6232 ( .A(n6270), .ZN(n6272) );
  AND2_X1 U6233 ( .A1(n6273), .A2(n6274), .ZN(n4418) );
  INV_X1 U6234 ( .A(n6275), .ZN(n6274) );
  AND2_X1 U6235 ( .A1(n6276), .A2(n4432), .ZN(n6275) );
  OR2_X1 U6236 ( .A1(n4432), .A2(n6276), .ZN(n6273) );
  OR2_X1 U6237 ( .A1(n6277), .A2(n6278), .ZN(n6276) );
  AND2_X1 U6238 ( .A1(n6279), .A2(n4431), .ZN(n6278) );
  INV_X1 U6239 ( .A(n4430), .ZN(n6279) );
  AND2_X1 U6240 ( .A1(n6280), .A2(n4430), .ZN(n6277) );
  OR2_X1 U6241 ( .A1(n4048), .A2(n4035), .ZN(n4430) );
  INV_X1 U6242 ( .A(n4431), .ZN(n6280) );
  OR2_X1 U6243 ( .A1(n6281), .A2(n6282), .ZN(n4431) );
  AND2_X1 U6244 ( .A1(n6271), .A2(n6270), .ZN(n6282) );
  AND2_X1 U6245 ( .A1(n6266), .A2(n6283), .ZN(n6281) );
  OR2_X1 U6246 ( .A1(n6270), .A2(n6271), .ZN(n6283) );
  OR2_X1 U6247 ( .A1(n4048), .A2(n3951), .ZN(n6271) );
  OR2_X1 U6248 ( .A1(n6284), .A2(n6285), .ZN(n6270) );
  AND2_X1 U6249 ( .A1(n6260), .A2(n6259), .ZN(n6285) );
  AND2_X1 U6250 ( .A1(n6255), .A2(n6286), .ZN(n6284) );
  OR2_X1 U6251 ( .A1(n6259), .A2(n6260), .ZN(n6286) );
  OR2_X1 U6252 ( .A1(n4048), .A2(n4041), .ZN(n6260) );
  OR2_X1 U6253 ( .A1(n6287), .A2(n6288), .ZN(n6259) );
  AND2_X1 U6254 ( .A1(n6249), .A2(n6248), .ZN(n6288) );
  AND2_X1 U6255 ( .A1(n6244), .A2(n6289), .ZN(n6287) );
  OR2_X1 U6256 ( .A1(n6248), .A2(n6249), .ZN(n6289) );
  OR2_X1 U6257 ( .A1(n4048), .A2(n3888), .ZN(n6249) );
  OR2_X1 U6258 ( .A1(n6290), .A2(n6291), .ZN(n6248) );
  AND2_X1 U6259 ( .A1(n3862), .A2(n6238), .ZN(n6291) );
  AND2_X1 U6260 ( .A1(n6234), .A2(n6292), .ZN(n6290) );
  OR2_X1 U6261 ( .A1(n6238), .A2(n3862), .ZN(n6292) );
  INV_X1 U6262 ( .A(n6237), .ZN(n3862) );
  AND2_X1 U6263 ( .A1(b_6_), .A2(a_6_), .ZN(n6237) );
  OR2_X1 U6264 ( .A1(n6293), .A2(n6294), .ZN(n6238) );
  AND2_X1 U6265 ( .A1(n6223), .A2(n6226), .ZN(n6294) );
  AND2_X1 U6266 ( .A1(n6295), .A2(n6228), .ZN(n6293) );
  OR2_X1 U6267 ( .A1(n6296), .A2(n6297), .ZN(n6228) );
  AND2_X1 U6268 ( .A1(n6217), .A2(n6216), .ZN(n6297) );
  AND2_X1 U6269 ( .A1(n6212), .A2(n6298), .ZN(n6296) );
  OR2_X1 U6270 ( .A1(n6216), .A2(n6217), .ZN(n6298) );
  OR2_X1 U6271 ( .A1(n4048), .A2(n4053), .ZN(n6217) );
  OR2_X1 U6272 ( .A1(n6299), .A2(n6300), .ZN(n6216) );
  AND2_X1 U6273 ( .A1(n6201), .A2(n6204), .ZN(n6300) );
  AND2_X1 U6274 ( .A1(n6301), .A2(n6206), .ZN(n6299) );
  OR2_X1 U6275 ( .A1(n6302), .A2(n6303), .ZN(n6206) );
  AND2_X1 U6276 ( .A1(n6190), .A2(n6193), .ZN(n6303) );
  AND2_X1 U6277 ( .A1(n6304), .A2(n6196), .ZN(n6302) );
  OR2_X1 U6278 ( .A1(n6305), .A2(n6306), .ZN(n6196) );
  AND2_X1 U6279 ( .A1(n6179), .A2(n6182), .ZN(n6306) );
  AND2_X1 U6280 ( .A1(n6307), .A2(n6184), .ZN(n6305) );
  OR2_X1 U6281 ( .A1(n6308), .A2(n6309), .ZN(n6184) );
  AND2_X1 U6282 ( .A1(n6168), .A2(n6171), .ZN(n6309) );
  AND2_X1 U6283 ( .A1(n6310), .A2(n6173), .ZN(n6308) );
  OR2_X1 U6284 ( .A1(n6311), .A2(n6312), .ZN(n6173) );
  AND2_X1 U6285 ( .A1(n6156), .A2(n6162), .ZN(n6312) );
  AND2_X1 U6286 ( .A1(n6163), .A2(n6313), .ZN(n6311) );
  OR2_X1 U6287 ( .A1(n6162), .A2(n6156), .ZN(n6313) );
  OR2_X1 U6288 ( .A1(n3682), .A2(n4048), .ZN(n6156) );
  OR2_X1 U6289 ( .A1(n3884), .A2(n6314), .ZN(n6162) );
  OR2_X1 U6290 ( .A1(n4070), .A2(n4048), .ZN(n6314) );
  INV_X1 U6291 ( .A(n6161), .ZN(n6163) );
  OR2_X1 U6292 ( .A1(n6315), .A2(n6316), .ZN(n6161) );
  AND2_X1 U6293 ( .A1(b_5_), .A2(n6317), .ZN(n6316) );
  OR2_X1 U6294 ( .A1(n6318), .A2(n3644), .ZN(n6317) );
  AND2_X1 U6295 ( .A1(a_14_), .A2(n4042), .ZN(n6318) );
  AND2_X1 U6296 ( .A1(b_4_), .A2(n6319), .ZN(n6315) );
  OR2_X1 U6297 ( .A1(n6320), .A2(n3647), .ZN(n6319) );
  AND2_X1 U6298 ( .A1(a_15_), .A2(n3884), .ZN(n6320) );
  OR2_X1 U6299 ( .A1(n6171), .A2(n6168), .ZN(n6310) );
  OR2_X1 U6300 ( .A1(n6321), .A2(n6322), .ZN(n6168) );
  AND2_X1 U6301 ( .A1(n6323), .A2(n6324), .ZN(n6322) );
  INV_X1 U6302 ( .A(n6325), .ZN(n6321) );
  OR2_X1 U6303 ( .A1(n6323), .A2(n6324), .ZN(n6325) );
  OR2_X1 U6304 ( .A1(n6326), .A2(n6327), .ZN(n6323) );
  AND2_X1 U6305 ( .A1(n6328), .A2(n6329), .ZN(n6327) );
  INV_X1 U6306 ( .A(n6330), .ZN(n6328) );
  AND2_X1 U6307 ( .A1(n6331), .A2(n6330), .ZN(n6326) );
  OR2_X1 U6308 ( .A1(n4072), .A2(n4048), .ZN(n6171) );
  OR2_X1 U6309 ( .A1(n6182), .A2(n6179), .ZN(n6307) );
  OR2_X1 U6310 ( .A1(n6332), .A2(n6333), .ZN(n6179) );
  INV_X1 U6311 ( .A(n6334), .ZN(n6333) );
  OR2_X1 U6312 ( .A1(n6335), .A2(n6336), .ZN(n6334) );
  AND2_X1 U6313 ( .A1(n6336), .A2(n6335), .ZN(n6332) );
  AND2_X1 U6314 ( .A1(n6337), .A2(n6338), .ZN(n6335) );
  OR2_X1 U6315 ( .A1(n6339), .A2(n6340), .ZN(n6338) );
  INV_X1 U6316 ( .A(n6341), .ZN(n6340) );
  OR2_X1 U6317 ( .A1(n6341), .A2(n6342), .ZN(n6337) );
  INV_X1 U6318 ( .A(n6339), .ZN(n6342) );
  OR2_X1 U6319 ( .A1(n3735), .A2(n4048), .ZN(n6182) );
  OR2_X1 U6320 ( .A1(n6193), .A2(n6190), .ZN(n6304) );
  OR2_X1 U6321 ( .A1(n6343), .A2(n6344), .ZN(n6190) );
  INV_X1 U6322 ( .A(n6345), .ZN(n6344) );
  OR2_X1 U6323 ( .A1(n6346), .A2(n6347), .ZN(n6345) );
  AND2_X1 U6324 ( .A1(n6347), .A2(n6346), .ZN(n6343) );
  AND2_X1 U6325 ( .A1(n6348), .A2(n6349), .ZN(n6346) );
  OR2_X1 U6326 ( .A1(n6350), .A2(n6351), .ZN(n6349) );
  INV_X1 U6327 ( .A(n6352), .ZN(n6351) );
  OR2_X1 U6328 ( .A1(n6352), .A2(n6353), .ZN(n6348) );
  INV_X1 U6329 ( .A(n6350), .ZN(n6353) );
  OR2_X1 U6330 ( .A1(n4048), .A2(n4059), .ZN(n6193) );
  OR2_X1 U6331 ( .A1(n6204), .A2(n6201), .ZN(n6301) );
  OR2_X1 U6332 ( .A1(n6354), .A2(n6355), .ZN(n6201) );
  INV_X1 U6333 ( .A(n6356), .ZN(n6355) );
  OR2_X1 U6334 ( .A1(n6357), .A2(n6358), .ZN(n6356) );
  AND2_X1 U6335 ( .A1(n6358), .A2(n6357), .ZN(n6354) );
  AND2_X1 U6336 ( .A1(n6359), .A2(n6360), .ZN(n6357) );
  OR2_X1 U6337 ( .A1(n6361), .A2(n6362), .ZN(n6360) );
  INV_X1 U6338 ( .A(n6363), .ZN(n6359) );
  AND2_X1 U6339 ( .A1(n6362), .A2(n6361), .ZN(n6363) );
  INV_X1 U6340 ( .A(n6364), .ZN(n6362) );
  OR2_X1 U6341 ( .A1(n4048), .A2(n3786), .ZN(n6204) );
  AND2_X1 U6342 ( .A1(n6365), .A2(n6366), .ZN(n6212) );
  INV_X1 U6343 ( .A(n6367), .ZN(n6366) );
  AND2_X1 U6344 ( .A1(n6368), .A2(n6369), .ZN(n6367) );
  OR2_X1 U6345 ( .A1(n6369), .A2(n6368), .ZN(n6365) );
  OR2_X1 U6346 ( .A1(n6370), .A2(n6371), .ZN(n6368) );
  AND2_X1 U6347 ( .A1(n6372), .A2(n6373), .ZN(n6371) );
  INV_X1 U6348 ( .A(n6374), .ZN(n6372) );
  AND2_X1 U6349 ( .A1(n6375), .A2(n6374), .ZN(n6370) );
  INV_X1 U6350 ( .A(n6373), .ZN(n6375) );
  OR2_X1 U6351 ( .A1(n6226), .A2(n6223), .ZN(n6295) );
  OR2_X1 U6352 ( .A1(n6376), .A2(n6377), .ZN(n6223) );
  INV_X1 U6353 ( .A(n6378), .ZN(n6377) );
  OR2_X1 U6354 ( .A1(n6379), .A2(n6380), .ZN(n6378) );
  AND2_X1 U6355 ( .A1(n6380), .A2(n6379), .ZN(n6376) );
  AND2_X1 U6356 ( .A1(n6381), .A2(n6382), .ZN(n6379) );
  OR2_X1 U6357 ( .A1(n6383), .A2(n6384), .ZN(n6382) );
  INV_X1 U6358 ( .A(n6385), .ZN(n6384) );
  OR2_X1 U6359 ( .A1(n6385), .A2(n6386), .ZN(n6381) );
  INV_X1 U6360 ( .A(n6383), .ZN(n6386) );
  OR2_X1 U6361 ( .A1(n4048), .A2(n3837), .ZN(n6226) );
  INV_X1 U6362 ( .A(b_6_), .ZN(n4048) );
  AND2_X1 U6363 ( .A1(n6387), .A2(n6388), .ZN(n6234) );
  INV_X1 U6364 ( .A(n6389), .ZN(n6388) );
  AND2_X1 U6365 ( .A1(n6390), .A2(n6391), .ZN(n6389) );
  OR2_X1 U6366 ( .A1(n6391), .A2(n6390), .ZN(n6387) );
  OR2_X1 U6367 ( .A1(n6392), .A2(n6393), .ZN(n6390) );
  AND2_X1 U6368 ( .A1(n6394), .A2(n6395), .ZN(n6393) );
  INV_X1 U6369 ( .A(n6396), .ZN(n6394) );
  AND2_X1 U6370 ( .A1(n6397), .A2(n6396), .ZN(n6392) );
  INV_X1 U6371 ( .A(n6395), .ZN(n6397) );
  AND2_X1 U6372 ( .A1(n6398), .A2(n6399), .ZN(n6244) );
  INV_X1 U6373 ( .A(n6400), .ZN(n6399) );
  AND2_X1 U6374 ( .A1(n6401), .A2(n6402), .ZN(n6400) );
  OR2_X1 U6375 ( .A1(n6402), .A2(n6401), .ZN(n6398) );
  OR2_X1 U6376 ( .A1(n6403), .A2(n6404), .ZN(n6401) );
  AND2_X1 U6377 ( .A1(n6405), .A2(n6406), .ZN(n6404) );
  INV_X1 U6378 ( .A(n6407), .ZN(n6405) );
  AND2_X1 U6379 ( .A1(n6408), .A2(n6407), .ZN(n6403) );
  INV_X1 U6380 ( .A(n6406), .ZN(n6408) );
  AND2_X1 U6381 ( .A1(n6409), .A2(n6410), .ZN(n6255) );
  INV_X1 U6382 ( .A(n6411), .ZN(n6410) );
  AND2_X1 U6383 ( .A1(n6412), .A2(n6413), .ZN(n6411) );
  OR2_X1 U6384 ( .A1(n6413), .A2(n6412), .ZN(n6409) );
  OR2_X1 U6385 ( .A1(n6414), .A2(n6415), .ZN(n6412) );
  AND2_X1 U6386 ( .A1(n3891), .A2(n6416), .ZN(n6415) );
  INV_X1 U6387 ( .A(n4045), .ZN(n3891) );
  AND2_X1 U6388 ( .A1(n6417), .A2(n4045), .ZN(n6414) );
  INV_X1 U6389 ( .A(n6416), .ZN(n6417) );
  AND2_X1 U6390 ( .A1(n6418), .A2(n6419), .ZN(n6266) );
  INV_X1 U6391 ( .A(n6420), .ZN(n6419) );
  AND2_X1 U6392 ( .A1(n6421), .A2(n6422), .ZN(n6420) );
  OR2_X1 U6393 ( .A1(n6422), .A2(n6421), .ZN(n6418) );
  OR2_X1 U6394 ( .A1(n6423), .A2(n6424), .ZN(n6421) );
  AND2_X1 U6395 ( .A1(n6425), .A2(n6426), .ZN(n6424) );
  INV_X1 U6396 ( .A(n6427), .ZN(n6425) );
  AND2_X1 U6397 ( .A1(n6428), .A2(n6427), .ZN(n6423) );
  INV_X1 U6398 ( .A(n6426), .ZN(n6428) );
  AND2_X1 U6399 ( .A1(n6429), .A2(n6430), .ZN(n4432) );
  INV_X1 U6400 ( .A(n6431), .ZN(n6430) );
  AND2_X1 U6401 ( .A1(n6432), .A2(n4446), .ZN(n6431) );
  OR2_X1 U6402 ( .A1(n4446), .A2(n6432), .ZN(n6429) );
  OR2_X1 U6403 ( .A1(n6433), .A2(n6434), .ZN(n6432) );
  AND2_X1 U6404 ( .A1(n6435), .A2(n4445), .ZN(n6434) );
  INV_X1 U6405 ( .A(n4444), .ZN(n6435) );
  AND2_X1 U6406 ( .A1(n6436), .A2(n4444), .ZN(n6433) );
  OR2_X1 U6407 ( .A1(n3884), .A2(n3951), .ZN(n4444) );
  INV_X1 U6408 ( .A(n4445), .ZN(n6436) );
  OR2_X1 U6409 ( .A1(n6437), .A2(n6438), .ZN(n4445) );
  AND2_X1 U6410 ( .A1(n6427), .A2(n6426), .ZN(n6438) );
  AND2_X1 U6411 ( .A1(n6422), .A2(n6439), .ZN(n6437) );
  OR2_X1 U6412 ( .A1(n6426), .A2(n6427), .ZN(n6439) );
  OR2_X1 U6413 ( .A1(n3884), .A2(n4041), .ZN(n6427) );
  OR2_X1 U6414 ( .A1(n6440), .A2(n6441), .ZN(n6426) );
  AND2_X1 U6415 ( .A1(n4045), .A2(n6416), .ZN(n6441) );
  AND2_X1 U6416 ( .A1(n6413), .A2(n6442), .ZN(n6440) );
  OR2_X1 U6417 ( .A1(n6416), .A2(n4045), .ZN(n6442) );
  OR2_X1 U6418 ( .A1(n3884), .A2(n3888), .ZN(n4045) );
  OR2_X1 U6419 ( .A1(n6443), .A2(n6444), .ZN(n6416) );
  AND2_X1 U6420 ( .A1(n6407), .A2(n6406), .ZN(n6444) );
  AND2_X1 U6421 ( .A1(n6402), .A2(n6445), .ZN(n6443) );
  OR2_X1 U6422 ( .A1(n6406), .A2(n6407), .ZN(n6445) );
  OR2_X1 U6423 ( .A1(n3884), .A2(n4047), .ZN(n6407) );
  OR2_X1 U6424 ( .A1(n6446), .A2(n6447), .ZN(n6406) );
  AND2_X1 U6425 ( .A1(n6396), .A2(n6395), .ZN(n6447) );
  AND2_X1 U6426 ( .A1(n6391), .A2(n6448), .ZN(n6446) );
  OR2_X1 U6427 ( .A1(n6395), .A2(n6396), .ZN(n6448) );
  OR2_X1 U6428 ( .A1(n3884), .A2(n3837), .ZN(n6396) );
  OR2_X1 U6429 ( .A1(n6449), .A2(n6450), .ZN(n6395) );
  AND2_X1 U6430 ( .A1(n6380), .A2(n6383), .ZN(n6450) );
  AND2_X1 U6431 ( .A1(n6451), .A2(n6385), .ZN(n6449) );
  OR2_X1 U6432 ( .A1(n6452), .A2(n6453), .ZN(n6385) );
  AND2_X1 U6433 ( .A1(n6374), .A2(n6373), .ZN(n6453) );
  AND2_X1 U6434 ( .A1(n6369), .A2(n6454), .ZN(n6452) );
  OR2_X1 U6435 ( .A1(n6373), .A2(n6374), .ZN(n6454) );
  OR2_X1 U6436 ( .A1(n3884), .A2(n3786), .ZN(n6374) );
  OR2_X1 U6437 ( .A1(n6455), .A2(n6456), .ZN(n6373) );
  AND2_X1 U6438 ( .A1(n6358), .A2(n6361), .ZN(n6456) );
  AND2_X1 U6439 ( .A1(n6457), .A2(n6364), .ZN(n6455) );
  OR2_X1 U6440 ( .A1(n6458), .A2(n6459), .ZN(n6364) );
  AND2_X1 U6441 ( .A1(n6347), .A2(n6350), .ZN(n6459) );
  AND2_X1 U6442 ( .A1(n6460), .A2(n6352), .ZN(n6458) );
  OR2_X1 U6443 ( .A1(n6461), .A2(n6462), .ZN(n6352) );
  AND2_X1 U6444 ( .A1(n6336), .A2(n6339), .ZN(n6462) );
  AND2_X1 U6445 ( .A1(n6463), .A2(n6341), .ZN(n6461) );
  OR2_X1 U6446 ( .A1(n6464), .A2(n6465), .ZN(n6341) );
  AND2_X1 U6447 ( .A1(n6324), .A2(n6330), .ZN(n6465) );
  AND2_X1 U6448 ( .A1(n6331), .A2(n6466), .ZN(n6464) );
  OR2_X1 U6449 ( .A1(n6330), .A2(n6324), .ZN(n6466) );
  OR2_X1 U6450 ( .A1(n3682), .A2(n3884), .ZN(n6324) );
  OR2_X1 U6451 ( .A1(n4042), .A2(n6467), .ZN(n6330) );
  OR2_X1 U6452 ( .A1(n4070), .A2(n3884), .ZN(n6467) );
  INV_X1 U6453 ( .A(n6329), .ZN(n6331) );
  OR2_X1 U6454 ( .A1(n6468), .A2(n6469), .ZN(n6329) );
  AND2_X1 U6455 ( .A1(b_4_), .A2(n6470), .ZN(n6469) );
  OR2_X1 U6456 ( .A1(n6471), .A2(n3644), .ZN(n6470) );
  AND2_X1 U6457 ( .A1(a_14_), .A2(n3947), .ZN(n6471) );
  AND2_X1 U6458 ( .A1(b_3_), .A2(n6472), .ZN(n6468) );
  OR2_X1 U6459 ( .A1(n6473), .A2(n3647), .ZN(n6472) );
  AND2_X1 U6460 ( .A1(a_15_), .A2(n4042), .ZN(n6473) );
  OR2_X1 U6461 ( .A1(n6339), .A2(n6336), .ZN(n6463) );
  OR2_X1 U6462 ( .A1(n6474), .A2(n6475), .ZN(n6336) );
  AND2_X1 U6463 ( .A1(n6476), .A2(n6477), .ZN(n6475) );
  INV_X1 U6464 ( .A(n6478), .ZN(n6474) );
  OR2_X1 U6465 ( .A1(n6476), .A2(n6477), .ZN(n6478) );
  OR2_X1 U6466 ( .A1(n6479), .A2(n6480), .ZN(n6476) );
  AND2_X1 U6467 ( .A1(n6481), .A2(n6482), .ZN(n6480) );
  INV_X1 U6468 ( .A(n6483), .ZN(n6481) );
  AND2_X1 U6469 ( .A1(n6484), .A2(n6483), .ZN(n6479) );
  OR2_X1 U6470 ( .A1(n4072), .A2(n3884), .ZN(n6339) );
  OR2_X1 U6471 ( .A1(n6350), .A2(n6347), .ZN(n6460) );
  OR2_X1 U6472 ( .A1(n6485), .A2(n6486), .ZN(n6347) );
  INV_X1 U6473 ( .A(n6487), .ZN(n6486) );
  OR2_X1 U6474 ( .A1(n6488), .A2(n6489), .ZN(n6487) );
  AND2_X1 U6475 ( .A1(n6489), .A2(n6488), .ZN(n6485) );
  AND2_X1 U6476 ( .A1(n6490), .A2(n6491), .ZN(n6488) );
  OR2_X1 U6477 ( .A1(n6492), .A2(n6493), .ZN(n6491) );
  INV_X1 U6478 ( .A(n6494), .ZN(n6493) );
  OR2_X1 U6479 ( .A1(n6494), .A2(n6495), .ZN(n6490) );
  INV_X1 U6480 ( .A(n6492), .ZN(n6495) );
  OR2_X1 U6481 ( .A1(n3735), .A2(n3884), .ZN(n6350) );
  OR2_X1 U6482 ( .A1(n6361), .A2(n6358), .ZN(n6457) );
  OR2_X1 U6483 ( .A1(n6496), .A2(n6497), .ZN(n6358) );
  INV_X1 U6484 ( .A(n6498), .ZN(n6497) );
  OR2_X1 U6485 ( .A1(n6499), .A2(n6500), .ZN(n6498) );
  AND2_X1 U6486 ( .A1(n6500), .A2(n6499), .ZN(n6496) );
  AND2_X1 U6487 ( .A1(n6501), .A2(n6502), .ZN(n6499) );
  OR2_X1 U6488 ( .A1(n6503), .A2(n6504), .ZN(n6502) );
  INV_X1 U6489 ( .A(n6505), .ZN(n6504) );
  OR2_X1 U6490 ( .A1(n6505), .A2(n6506), .ZN(n6501) );
  INV_X1 U6491 ( .A(n6503), .ZN(n6506) );
  OR2_X1 U6492 ( .A1(n4059), .A2(n3884), .ZN(n6361) );
  AND2_X1 U6493 ( .A1(n6507), .A2(n6508), .ZN(n6369) );
  INV_X1 U6494 ( .A(n6509), .ZN(n6508) );
  AND2_X1 U6495 ( .A1(n6510), .A2(n6511), .ZN(n6509) );
  OR2_X1 U6496 ( .A1(n6511), .A2(n6510), .ZN(n6507) );
  OR2_X1 U6497 ( .A1(n6512), .A2(n6513), .ZN(n6510) );
  AND2_X1 U6498 ( .A1(n6514), .A2(n6515), .ZN(n6513) );
  AND2_X1 U6499 ( .A1(n6516), .A2(n6517), .ZN(n6512) );
  INV_X1 U6500 ( .A(n6515), .ZN(n6516) );
  OR2_X1 U6501 ( .A1(n6383), .A2(n6380), .ZN(n6451) );
  OR2_X1 U6502 ( .A1(n6518), .A2(n6519), .ZN(n6380) );
  INV_X1 U6503 ( .A(n6520), .ZN(n6519) );
  OR2_X1 U6504 ( .A1(n6521), .A2(n6522), .ZN(n6520) );
  AND2_X1 U6505 ( .A1(n6522), .A2(n6521), .ZN(n6518) );
  AND2_X1 U6506 ( .A1(n6523), .A2(n6524), .ZN(n6521) );
  OR2_X1 U6507 ( .A1(n6525), .A2(n6526), .ZN(n6524) );
  INV_X1 U6508 ( .A(n6527), .ZN(n6526) );
  OR2_X1 U6509 ( .A1(n6527), .A2(n6528), .ZN(n6523) );
  INV_X1 U6510 ( .A(n6525), .ZN(n6528) );
  OR2_X1 U6511 ( .A1(n3884), .A2(n4053), .ZN(n6383) );
  INV_X1 U6512 ( .A(b_5_), .ZN(n3884) );
  AND2_X1 U6513 ( .A1(n6529), .A2(n6530), .ZN(n6391) );
  INV_X1 U6514 ( .A(n6531), .ZN(n6530) );
  AND2_X1 U6515 ( .A1(n6532), .A2(n6533), .ZN(n6531) );
  OR2_X1 U6516 ( .A1(n6533), .A2(n6532), .ZN(n6529) );
  OR2_X1 U6517 ( .A1(n6534), .A2(n6535), .ZN(n6532) );
  AND2_X1 U6518 ( .A1(n6536), .A2(n6537), .ZN(n6535) );
  INV_X1 U6519 ( .A(n6538), .ZN(n6536) );
  AND2_X1 U6520 ( .A1(n6539), .A2(n6538), .ZN(n6534) );
  INV_X1 U6521 ( .A(n6537), .ZN(n6539) );
  AND2_X1 U6522 ( .A1(n6540), .A2(n6541), .ZN(n6402) );
  INV_X1 U6523 ( .A(n6542), .ZN(n6541) );
  AND2_X1 U6524 ( .A1(n6543), .A2(n6544), .ZN(n6542) );
  OR2_X1 U6525 ( .A1(n6544), .A2(n6543), .ZN(n6540) );
  OR2_X1 U6526 ( .A1(n6545), .A2(n6546), .ZN(n6543) );
  AND2_X1 U6527 ( .A1(n6547), .A2(n6548), .ZN(n6546) );
  INV_X1 U6528 ( .A(n6549), .ZN(n6547) );
  AND2_X1 U6529 ( .A1(n6550), .A2(n6549), .ZN(n6545) );
  INV_X1 U6530 ( .A(n6548), .ZN(n6550) );
  AND2_X1 U6531 ( .A1(n6551), .A2(n6552), .ZN(n6413) );
  INV_X1 U6532 ( .A(n6553), .ZN(n6552) );
  AND2_X1 U6533 ( .A1(n6554), .A2(n6555), .ZN(n6553) );
  OR2_X1 U6534 ( .A1(n6555), .A2(n6554), .ZN(n6551) );
  OR2_X1 U6535 ( .A1(n6556), .A2(n6557), .ZN(n6554) );
  AND2_X1 U6536 ( .A1(n6558), .A2(n6559), .ZN(n6557) );
  INV_X1 U6537 ( .A(n6560), .ZN(n6558) );
  AND2_X1 U6538 ( .A1(n6561), .A2(n6560), .ZN(n6556) );
  INV_X1 U6539 ( .A(n6559), .ZN(n6561) );
  AND2_X1 U6540 ( .A1(n6562), .A2(n6563), .ZN(n6422) );
  INV_X1 U6541 ( .A(n6564), .ZN(n6563) );
  AND2_X1 U6542 ( .A1(n6565), .A2(n6566), .ZN(n6564) );
  OR2_X1 U6543 ( .A1(n6566), .A2(n6565), .ZN(n6562) );
  OR2_X1 U6544 ( .A1(n6567), .A2(n6568), .ZN(n6565) );
  AND2_X1 U6545 ( .A1(n6569), .A2(n6570), .ZN(n6568) );
  INV_X1 U6546 ( .A(n6571), .ZN(n6569) );
  AND2_X1 U6547 ( .A1(n6572), .A2(n6571), .ZN(n6567) );
  INV_X1 U6548 ( .A(n6570), .ZN(n6572) );
  AND2_X1 U6549 ( .A1(n6573), .A2(n6574), .ZN(n4446) );
  INV_X1 U6550 ( .A(n6575), .ZN(n6574) );
  AND2_X1 U6551 ( .A1(n6576), .A2(n4459), .ZN(n6575) );
  OR2_X1 U6552 ( .A1(n4459), .A2(n6576), .ZN(n6573) );
  OR2_X1 U6553 ( .A1(n6577), .A2(n6578), .ZN(n6576) );
  AND2_X1 U6554 ( .A1(n4461), .A2(n4458), .ZN(n6578) );
  INV_X1 U6555 ( .A(n6579), .ZN(n6577) );
  OR2_X1 U6556 ( .A1(n4458), .A2(n4461), .ZN(n6579) );
  AND2_X1 U6557 ( .A1(b_4_), .A2(a_4_), .ZN(n4461) );
  OR2_X1 U6558 ( .A1(n6580), .A2(n6581), .ZN(n4458) );
  AND2_X1 U6559 ( .A1(n6571), .A2(n6570), .ZN(n6581) );
  AND2_X1 U6560 ( .A1(n6566), .A2(n6582), .ZN(n6580) );
  OR2_X1 U6561 ( .A1(n6570), .A2(n6571), .ZN(n6582) );
  OR2_X1 U6562 ( .A1(n4042), .A2(n3888), .ZN(n6571) );
  OR2_X1 U6563 ( .A1(n6583), .A2(n6584), .ZN(n6570) );
  AND2_X1 U6564 ( .A1(n6560), .A2(n6559), .ZN(n6584) );
  AND2_X1 U6565 ( .A1(n6555), .A2(n6585), .ZN(n6583) );
  OR2_X1 U6566 ( .A1(n6559), .A2(n6560), .ZN(n6585) );
  OR2_X1 U6567 ( .A1(n4042), .A2(n4047), .ZN(n6560) );
  OR2_X1 U6568 ( .A1(n6586), .A2(n6587), .ZN(n6559) );
  AND2_X1 U6569 ( .A1(n6549), .A2(n6548), .ZN(n6587) );
  AND2_X1 U6570 ( .A1(n6544), .A2(n6588), .ZN(n6586) );
  OR2_X1 U6571 ( .A1(n6548), .A2(n6549), .ZN(n6588) );
  OR2_X1 U6572 ( .A1(n4042), .A2(n3837), .ZN(n6549) );
  OR2_X1 U6573 ( .A1(n6589), .A2(n6590), .ZN(n6548) );
  AND2_X1 U6574 ( .A1(n6538), .A2(n6537), .ZN(n6590) );
  AND2_X1 U6575 ( .A1(n6533), .A2(n6591), .ZN(n6589) );
  OR2_X1 U6576 ( .A1(n6537), .A2(n6538), .ZN(n6591) );
  OR2_X1 U6577 ( .A1(n4042), .A2(n4053), .ZN(n6538) );
  OR2_X1 U6578 ( .A1(n6592), .A2(n6593), .ZN(n6537) );
  AND2_X1 U6579 ( .A1(n6522), .A2(n6525), .ZN(n6593) );
  AND2_X1 U6580 ( .A1(n6594), .A2(n6527), .ZN(n6592) );
  OR2_X1 U6581 ( .A1(n6595), .A2(n6596), .ZN(n6527) );
  AND2_X1 U6582 ( .A1(n6517), .A2(n6515), .ZN(n6596) );
  AND2_X1 U6583 ( .A1(n6511), .A2(n6597), .ZN(n6595) );
  OR2_X1 U6584 ( .A1(n6515), .A2(n6517), .ZN(n6597) );
  INV_X1 U6585 ( .A(n6514), .ZN(n6517) );
  AND2_X1 U6586 ( .A1(a_10_), .A2(b_4_), .ZN(n6514) );
  OR2_X1 U6587 ( .A1(n6598), .A2(n6599), .ZN(n6515) );
  AND2_X1 U6588 ( .A1(n6500), .A2(n6503), .ZN(n6599) );
  AND2_X1 U6589 ( .A1(n6600), .A2(n6505), .ZN(n6598) );
  OR2_X1 U6590 ( .A1(n6601), .A2(n6602), .ZN(n6505) );
  AND2_X1 U6591 ( .A1(n6489), .A2(n6492), .ZN(n6602) );
  AND2_X1 U6592 ( .A1(n6603), .A2(n6494), .ZN(n6601) );
  OR2_X1 U6593 ( .A1(n6604), .A2(n6605), .ZN(n6494) );
  AND2_X1 U6594 ( .A1(n6477), .A2(n6483), .ZN(n6605) );
  AND2_X1 U6595 ( .A1(n6484), .A2(n6606), .ZN(n6604) );
  OR2_X1 U6596 ( .A1(n6483), .A2(n6477), .ZN(n6606) );
  OR2_X1 U6597 ( .A1(n3682), .A2(n4042), .ZN(n6477) );
  OR2_X1 U6598 ( .A1(n3947), .A2(n6607), .ZN(n6483) );
  OR2_X1 U6599 ( .A1(n4070), .A2(n4042), .ZN(n6607) );
  INV_X1 U6600 ( .A(n6482), .ZN(n6484) );
  OR2_X1 U6601 ( .A1(n6608), .A2(n6609), .ZN(n6482) );
  AND2_X1 U6602 ( .A1(b_3_), .A2(n6610), .ZN(n6609) );
  OR2_X1 U6603 ( .A1(n6611), .A2(n3644), .ZN(n6610) );
  AND2_X1 U6604 ( .A1(a_14_), .A2(n4036), .ZN(n6611) );
  AND2_X1 U6605 ( .A1(b_2_), .A2(n6612), .ZN(n6608) );
  OR2_X1 U6606 ( .A1(n6613), .A2(n3647), .ZN(n6612) );
  AND2_X1 U6607 ( .A1(a_15_), .A2(n3947), .ZN(n6613) );
  OR2_X1 U6608 ( .A1(n6492), .A2(n6489), .ZN(n6603) );
  OR2_X1 U6609 ( .A1(n6614), .A2(n6615), .ZN(n6489) );
  AND2_X1 U6610 ( .A1(n6616), .A2(n6617), .ZN(n6615) );
  INV_X1 U6611 ( .A(n6618), .ZN(n6614) );
  OR2_X1 U6612 ( .A1(n6616), .A2(n6617), .ZN(n6618) );
  OR2_X1 U6613 ( .A1(n6619), .A2(n6620), .ZN(n6616) );
  AND2_X1 U6614 ( .A1(n6621), .A2(n6622), .ZN(n6620) );
  INV_X1 U6615 ( .A(n6623), .ZN(n6621) );
  AND2_X1 U6616 ( .A1(n6624), .A2(n6623), .ZN(n6619) );
  OR2_X1 U6617 ( .A1(n4072), .A2(n4042), .ZN(n6492) );
  OR2_X1 U6618 ( .A1(n6503), .A2(n6500), .ZN(n6600) );
  OR2_X1 U6619 ( .A1(n6625), .A2(n6626), .ZN(n6500) );
  INV_X1 U6620 ( .A(n6627), .ZN(n6626) );
  OR2_X1 U6621 ( .A1(n6628), .A2(n6629), .ZN(n6627) );
  AND2_X1 U6622 ( .A1(n6629), .A2(n6628), .ZN(n6625) );
  AND2_X1 U6623 ( .A1(n6630), .A2(n6631), .ZN(n6628) );
  OR2_X1 U6624 ( .A1(n6632), .A2(n6633), .ZN(n6631) );
  INV_X1 U6625 ( .A(n6634), .ZN(n6633) );
  OR2_X1 U6626 ( .A1(n6634), .A2(n6635), .ZN(n6630) );
  INV_X1 U6627 ( .A(n6632), .ZN(n6635) );
  OR2_X1 U6628 ( .A1(n3735), .A2(n4042), .ZN(n6503) );
  AND2_X1 U6629 ( .A1(n6636), .A2(n6637), .ZN(n6511) );
  INV_X1 U6630 ( .A(n6638), .ZN(n6637) );
  AND2_X1 U6631 ( .A1(n6639), .A2(n6640), .ZN(n6638) );
  OR2_X1 U6632 ( .A1(n6640), .A2(n6639), .ZN(n6636) );
  OR2_X1 U6633 ( .A1(n6641), .A2(n6642), .ZN(n6639) );
  AND2_X1 U6634 ( .A1(n6643), .A2(n6644), .ZN(n6642) );
  INV_X1 U6635 ( .A(n6645), .ZN(n6643) );
  AND2_X1 U6636 ( .A1(n6646), .A2(n6645), .ZN(n6641) );
  INV_X1 U6637 ( .A(n6644), .ZN(n6646) );
  OR2_X1 U6638 ( .A1(n6525), .A2(n6522), .ZN(n6594) );
  OR2_X1 U6639 ( .A1(n6647), .A2(n6648), .ZN(n6522) );
  INV_X1 U6640 ( .A(n6649), .ZN(n6648) );
  OR2_X1 U6641 ( .A1(n6650), .A2(n6651), .ZN(n6649) );
  AND2_X1 U6642 ( .A1(n6651), .A2(n6650), .ZN(n6647) );
  AND2_X1 U6643 ( .A1(n6652), .A2(n6653), .ZN(n6650) );
  OR2_X1 U6644 ( .A1(n6654), .A2(n6655), .ZN(n6653) );
  INV_X1 U6645 ( .A(n6656), .ZN(n6652) );
  AND2_X1 U6646 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  INV_X1 U6647 ( .A(n6657), .ZN(n6655) );
  OR2_X1 U6648 ( .A1(n3786), .A2(n4042), .ZN(n6525) );
  INV_X1 U6649 ( .A(b_4_), .ZN(n4042) );
  AND2_X1 U6650 ( .A1(n6658), .A2(n6659), .ZN(n6533) );
  INV_X1 U6651 ( .A(n6660), .ZN(n6659) );
  AND2_X1 U6652 ( .A1(n6661), .A2(n6662), .ZN(n6660) );
  OR2_X1 U6653 ( .A1(n6662), .A2(n6661), .ZN(n6658) );
  OR2_X1 U6654 ( .A1(n6663), .A2(n6664), .ZN(n6661) );
  AND2_X1 U6655 ( .A1(n6665), .A2(n6666), .ZN(n6664) );
  INV_X1 U6656 ( .A(n6667), .ZN(n6665) );
  AND2_X1 U6657 ( .A1(n6668), .A2(n6667), .ZN(n6663) );
  INV_X1 U6658 ( .A(n6666), .ZN(n6668) );
  AND2_X1 U6659 ( .A1(n6669), .A2(n6670), .ZN(n6544) );
  INV_X1 U6660 ( .A(n6671), .ZN(n6670) );
  AND2_X1 U6661 ( .A1(n6672), .A2(n6673), .ZN(n6671) );
  OR2_X1 U6662 ( .A1(n6673), .A2(n6672), .ZN(n6669) );
  OR2_X1 U6663 ( .A1(n6674), .A2(n6675), .ZN(n6672) );
  AND2_X1 U6664 ( .A1(n6676), .A2(n6677), .ZN(n6675) );
  INV_X1 U6665 ( .A(n6678), .ZN(n6676) );
  AND2_X1 U6666 ( .A1(n6679), .A2(n6678), .ZN(n6674) );
  INV_X1 U6667 ( .A(n6677), .ZN(n6679) );
  AND2_X1 U6668 ( .A1(n6680), .A2(n6681), .ZN(n6555) );
  INV_X1 U6669 ( .A(n6682), .ZN(n6681) );
  AND2_X1 U6670 ( .A1(n6683), .A2(n6684), .ZN(n6682) );
  OR2_X1 U6671 ( .A1(n6684), .A2(n6683), .ZN(n6680) );
  OR2_X1 U6672 ( .A1(n6685), .A2(n6686), .ZN(n6683) );
  AND2_X1 U6673 ( .A1(n6687), .A2(n6688), .ZN(n6686) );
  INV_X1 U6674 ( .A(n6689), .ZN(n6687) );
  AND2_X1 U6675 ( .A1(n6690), .A2(n6689), .ZN(n6685) );
  INV_X1 U6676 ( .A(n6688), .ZN(n6690) );
  AND2_X1 U6677 ( .A1(n6691), .A2(n6692), .ZN(n6566) );
  INV_X1 U6678 ( .A(n6693), .ZN(n6692) );
  AND2_X1 U6679 ( .A1(n6694), .A2(n6695), .ZN(n6693) );
  OR2_X1 U6680 ( .A1(n6695), .A2(n6694), .ZN(n6691) );
  OR2_X1 U6681 ( .A1(n6696), .A2(n6697), .ZN(n6694) );
  AND2_X1 U6682 ( .A1(n6698), .A2(n6699), .ZN(n6697) );
  INV_X1 U6683 ( .A(n6700), .ZN(n6698) );
  AND2_X1 U6684 ( .A1(n6701), .A2(n6700), .ZN(n6696) );
  INV_X1 U6685 ( .A(n6699), .ZN(n6701) );
  AND2_X1 U6686 ( .A1(n6702), .A2(n6703), .ZN(n4459) );
  INV_X1 U6687 ( .A(n6704), .ZN(n6703) );
  AND2_X1 U6688 ( .A1(n6705), .A2(n4474), .ZN(n6704) );
  OR2_X1 U6689 ( .A1(n4474), .A2(n6705), .ZN(n6702) );
  OR2_X1 U6690 ( .A1(n6706), .A2(n6707), .ZN(n6705) );
  AND2_X1 U6691 ( .A1(n6708), .A2(n4473), .ZN(n6707) );
  INV_X1 U6692 ( .A(n4472), .ZN(n6708) );
  AND2_X1 U6693 ( .A1(n6709), .A2(n4472), .ZN(n6706) );
  OR2_X1 U6694 ( .A1(n3947), .A2(n3888), .ZN(n4472) );
  INV_X1 U6695 ( .A(n4473), .ZN(n6709) );
  OR2_X1 U6696 ( .A1(n6710), .A2(n6711), .ZN(n4473) );
  AND2_X1 U6697 ( .A1(n6700), .A2(n6699), .ZN(n6711) );
  AND2_X1 U6698 ( .A1(n6695), .A2(n6712), .ZN(n6710) );
  OR2_X1 U6699 ( .A1(n6699), .A2(n6700), .ZN(n6712) );
  OR2_X1 U6700 ( .A1(n3947), .A2(n4047), .ZN(n6700) );
  OR2_X1 U6701 ( .A1(n6713), .A2(n6714), .ZN(n6699) );
  AND2_X1 U6702 ( .A1(n6689), .A2(n6688), .ZN(n6714) );
  AND2_X1 U6703 ( .A1(n6684), .A2(n6715), .ZN(n6713) );
  OR2_X1 U6704 ( .A1(n6688), .A2(n6689), .ZN(n6715) );
  OR2_X1 U6705 ( .A1(n3947), .A2(n3837), .ZN(n6689) );
  OR2_X1 U6706 ( .A1(n6716), .A2(n6717), .ZN(n6688) );
  AND2_X1 U6707 ( .A1(n6678), .A2(n6677), .ZN(n6717) );
  AND2_X1 U6708 ( .A1(n6673), .A2(n6718), .ZN(n6716) );
  OR2_X1 U6709 ( .A1(n6677), .A2(n6678), .ZN(n6718) );
  OR2_X1 U6710 ( .A1(n4053), .A2(n3947), .ZN(n6678) );
  OR2_X1 U6711 ( .A1(n6719), .A2(n6720), .ZN(n6677) );
  AND2_X1 U6712 ( .A1(n6667), .A2(n6666), .ZN(n6720) );
  AND2_X1 U6713 ( .A1(n6662), .A2(n6721), .ZN(n6719) );
  OR2_X1 U6714 ( .A1(n6666), .A2(n6667), .ZN(n6721) );
  OR2_X1 U6715 ( .A1(n3786), .A2(n3947), .ZN(n6667) );
  OR2_X1 U6716 ( .A1(n6722), .A2(n6723), .ZN(n6666) );
  AND2_X1 U6717 ( .A1(n6651), .A2(n6654), .ZN(n6723) );
  AND2_X1 U6718 ( .A1(n6724), .A2(n6657), .ZN(n6722) );
  OR2_X1 U6719 ( .A1(n6725), .A2(n6726), .ZN(n6657) );
  AND2_X1 U6720 ( .A1(n6645), .A2(n6644), .ZN(n6726) );
  AND2_X1 U6721 ( .A1(n6640), .A2(n6727), .ZN(n6725) );
  OR2_X1 U6722 ( .A1(n6644), .A2(n6645), .ZN(n6727) );
  OR2_X1 U6723 ( .A1(n3735), .A2(n3947), .ZN(n6645) );
  OR2_X1 U6724 ( .A1(n6728), .A2(n6729), .ZN(n6644) );
  AND2_X1 U6725 ( .A1(n6629), .A2(n6632), .ZN(n6729) );
  AND2_X1 U6726 ( .A1(n6730), .A2(n6634), .ZN(n6728) );
  OR2_X1 U6727 ( .A1(n6731), .A2(n6732), .ZN(n6634) );
  AND2_X1 U6728 ( .A1(n6617), .A2(n6623), .ZN(n6732) );
  AND2_X1 U6729 ( .A1(n6624), .A2(n6733), .ZN(n6731) );
  OR2_X1 U6730 ( .A1(n6623), .A2(n6617), .ZN(n6733) );
  OR2_X1 U6731 ( .A1(n3682), .A2(n3947), .ZN(n6617) );
  OR2_X1 U6732 ( .A1(n4036), .A2(n6734), .ZN(n6623) );
  OR2_X1 U6733 ( .A1(n4070), .A2(n3947), .ZN(n6734) );
  INV_X1 U6734 ( .A(n6622), .ZN(n6624) );
  OR2_X1 U6735 ( .A1(n6735), .A2(n6736), .ZN(n6622) );
  AND2_X1 U6736 ( .A1(b_2_), .A2(n6737), .ZN(n6736) );
  OR2_X1 U6737 ( .A1(n6738), .A2(n3644), .ZN(n6737) );
  AND2_X1 U6738 ( .A1(a_14_), .A2(n3998), .ZN(n6738) );
  AND2_X1 U6739 ( .A1(b_1_), .A2(n6739), .ZN(n6735) );
  OR2_X1 U6740 ( .A1(n6740), .A2(n3647), .ZN(n6739) );
  AND2_X1 U6741 ( .A1(a_15_), .A2(n4036), .ZN(n6740) );
  OR2_X1 U6742 ( .A1(n6632), .A2(n6629), .ZN(n6730) );
  OR2_X1 U6743 ( .A1(n6741), .A2(n6742), .ZN(n6629) );
  AND2_X1 U6744 ( .A1(n6743), .A2(n6744), .ZN(n6742) );
  INV_X1 U6745 ( .A(n6745), .ZN(n6741) );
  OR2_X1 U6746 ( .A1(n6743), .A2(n6744), .ZN(n6745) );
  OR2_X1 U6747 ( .A1(n6746), .A2(n6747), .ZN(n6743) );
  AND2_X1 U6748 ( .A1(n6748), .A2(n6749), .ZN(n6747) );
  INV_X1 U6749 ( .A(n6750), .ZN(n6748) );
  AND2_X1 U6750 ( .A1(n6751), .A2(n6750), .ZN(n6746) );
  OR2_X1 U6751 ( .A1(n4072), .A2(n3947), .ZN(n6632) );
  AND2_X1 U6752 ( .A1(n6752), .A2(n6753), .ZN(n6640) );
  INV_X1 U6753 ( .A(n6754), .ZN(n6753) );
  AND2_X1 U6754 ( .A1(n6755), .A2(n6756), .ZN(n6754) );
  OR2_X1 U6755 ( .A1(n6756), .A2(n6755), .ZN(n6752) );
  OR2_X1 U6756 ( .A1(n6757), .A2(n6758), .ZN(n6755) );
  AND2_X1 U6757 ( .A1(n6759), .A2(n6760), .ZN(n6758) );
  INV_X1 U6758 ( .A(n6761), .ZN(n6759) );
  AND2_X1 U6759 ( .A1(n6762), .A2(n6761), .ZN(n6757) );
  INV_X1 U6760 ( .A(n6760), .ZN(n6762) );
  OR2_X1 U6761 ( .A1(n6654), .A2(n6651), .ZN(n6724) );
  OR2_X1 U6762 ( .A1(n6763), .A2(n6764), .ZN(n6651) );
  INV_X1 U6763 ( .A(n6765), .ZN(n6764) );
  OR2_X1 U6764 ( .A1(n6766), .A2(n6767), .ZN(n6765) );
  AND2_X1 U6765 ( .A1(n6767), .A2(n6766), .ZN(n6763) );
  AND2_X1 U6766 ( .A1(n6768), .A2(n6769), .ZN(n6766) );
  OR2_X1 U6767 ( .A1(n6770), .A2(n6771), .ZN(n6769) );
  INV_X1 U6768 ( .A(n6772), .ZN(n6771) );
  OR2_X1 U6769 ( .A1(n6772), .A2(n6773), .ZN(n6768) );
  INV_X1 U6770 ( .A(n6770), .ZN(n6773) );
  OR2_X1 U6771 ( .A1(n4059), .A2(n3947), .ZN(n6654) );
  INV_X1 U6772 ( .A(b_3_), .ZN(n3947) );
  AND2_X1 U6773 ( .A1(n6774), .A2(n6775), .ZN(n6662) );
  INV_X1 U6774 ( .A(n6776), .ZN(n6775) );
  AND2_X1 U6775 ( .A1(n6777), .A2(n6778), .ZN(n6776) );
  OR2_X1 U6776 ( .A1(n6778), .A2(n6777), .ZN(n6774) );
  OR2_X1 U6777 ( .A1(n6779), .A2(n6780), .ZN(n6777) );
  AND2_X1 U6778 ( .A1(n6781), .A2(n6782), .ZN(n6780) );
  AND2_X1 U6779 ( .A1(n6783), .A2(n6784), .ZN(n6779) );
  INV_X1 U6780 ( .A(n6782), .ZN(n6783) );
  AND2_X1 U6781 ( .A1(n6785), .A2(n6786), .ZN(n6673) );
  INV_X1 U6782 ( .A(n6787), .ZN(n6786) );
  AND2_X1 U6783 ( .A1(n6788), .A2(n6789), .ZN(n6787) );
  OR2_X1 U6784 ( .A1(n6789), .A2(n6788), .ZN(n6785) );
  OR2_X1 U6785 ( .A1(n6790), .A2(n6791), .ZN(n6788) );
  AND2_X1 U6786 ( .A1(n6792), .A2(n6793), .ZN(n6791) );
  INV_X1 U6787 ( .A(n6794), .ZN(n6792) );
  AND2_X1 U6788 ( .A1(n6795), .A2(n6794), .ZN(n6790) );
  INV_X1 U6789 ( .A(n6793), .ZN(n6795) );
  AND2_X1 U6790 ( .A1(n6796), .A2(n6797), .ZN(n6684) );
  INV_X1 U6791 ( .A(n6798), .ZN(n6797) );
  AND2_X1 U6792 ( .A1(n6799), .A2(n6800), .ZN(n6798) );
  OR2_X1 U6793 ( .A1(n6800), .A2(n6799), .ZN(n6796) );
  OR2_X1 U6794 ( .A1(n6801), .A2(n6802), .ZN(n6799) );
  AND2_X1 U6795 ( .A1(n6803), .A2(n6804), .ZN(n6802) );
  INV_X1 U6796 ( .A(n6805), .ZN(n6803) );
  AND2_X1 U6797 ( .A1(n6806), .A2(n6805), .ZN(n6801) );
  INV_X1 U6798 ( .A(n6804), .ZN(n6806) );
  AND2_X1 U6799 ( .A1(n6807), .A2(n6808), .ZN(n6695) );
  INV_X1 U6800 ( .A(n6809), .ZN(n6808) );
  AND2_X1 U6801 ( .A1(n6810), .A2(n6811), .ZN(n6809) );
  OR2_X1 U6802 ( .A1(n6811), .A2(n6810), .ZN(n6807) );
  OR2_X1 U6803 ( .A1(n6812), .A2(n6813), .ZN(n6810) );
  AND2_X1 U6804 ( .A1(n6814), .A2(n6815), .ZN(n6813) );
  INV_X1 U6805 ( .A(n6816), .ZN(n6814) );
  AND2_X1 U6806 ( .A1(n6817), .A2(n6816), .ZN(n6812) );
  INV_X1 U6807 ( .A(n6815), .ZN(n6817) );
  AND2_X1 U6808 ( .A1(n6818), .A2(n6819), .ZN(n4474) );
  INV_X1 U6809 ( .A(n6820), .ZN(n6819) );
  AND2_X1 U6810 ( .A1(n6821), .A2(n6822), .ZN(n6820) );
  OR2_X1 U6811 ( .A1(n6822), .A2(n6821), .ZN(n6818) );
  OR2_X1 U6812 ( .A1(n6823), .A2(n6824), .ZN(n6821) );
  AND2_X1 U6813 ( .A1(n6825), .A2(n6826), .ZN(n6824) );
  INV_X1 U6814 ( .A(n6827), .ZN(n6825) );
  AND2_X1 U6815 ( .A1(n6828), .A2(n6827), .ZN(n6823) );
  INV_X1 U6816 ( .A(n6826), .ZN(n6828) );
  AND2_X1 U6817 ( .A1(n3924), .A2(n3925), .ZN(n3926) );
  INV_X1 U6818 ( .A(n6829), .ZN(n3925) );
  OR2_X1 U6819 ( .A1(n4139), .A2(n4140), .ZN(n6829) );
  OR2_X1 U6820 ( .A1(n6830), .A2(n6831), .ZN(n4140) );
  AND2_X1 U6821 ( .A1(n4165), .A2(n4168), .ZN(n6831) );
  AND2_X1 U6822 ( .A1(n4160), .A2(n6832), .ZN(n6830) );
  OR2_X1 U6823 ( .A1(n4168), .A2(n4165), .ZN(n6832) );
  OR2_X1 U6824 ( .A1(n4036), .A2(n4028), .ZN(n4165) );
  OR2_X1 U6825 ( .A1(n6833), .A2(n6834), .ZN(n4168) );
  AND2_X1 U6826 ( .A1(n4200), .A2(n4199), .ZN(n6834) );
  AND2_X1 U6827 ( .A1(n4195), .A2(n6835), .ZN(n6833) );
  OR2_X1 U6828 ( .A1(n4199), .A2(n4200), .ZN(n6835) );
  OR2_X1 U6829 ( .A1(n4036), .A2(n4002), .ZN(n4200) );
  OR2_X1 U6830 ( .A1(n6836), .A2(n6837), .ZN(n4199) );
  AND2_X1 U6831 ( .A1(n3976), .A2(n4254), .ZN(n6837) );
  AND2_X1 U6832 ( .A1(n4250), .A2(n6838), .ZN(n6836) );
  OR2_X1 U6833 ( .A1(n4254), .A2(n3976), .ZN(n6838) );
  INV_X1 U6834 ( .A(n4253), .ZN(n3976) );
  AND2_X1 U6835 ( .A1(b_2_), .A2(a_2_), .ZN(n4253) );
  OR2_X1 U6836 ( .A1(n6839), .A2(n6840), .ZN(n4254) );
  AND2_X1 U6837 ( .A1(n4314), .A2(n4313), .ZN(n6840) );
  AND2_X1 U6838 ( .A1(n4309), .A2(n6841), .ZN(n6839) );
  OR2_X1 U6839 ( .A1(n4313), .A2(n4314), .ZN(n6841) );
  OR2_X1 U6840 ( .A1(n4036), .A2(n3951), .ZN(n4314) );
  OR2_X1 U6841 ( .A1(n6842), .A2(n6843), .ZN(n4313) );
  AND2_X1 U6842 ( .A1(n4396), .A2(n4395), .ZN(n6843) );
  AND2_X1 U6843 ( .A1(n4391), .A2(n6844), .ZN(n6842) );
  OR2_X1 U6844 ( .A1(n4395), .A2(n4396), .ZN(n6844) );
  OR2_X1 U6845 ( .A1(n4036), .A2(n4041), .ZN(n4396) );
  OR2_X1 U6846 ( .A1(n6845), .A2(n6846), .ZN(n4395) );
  AND2_X1 U6847 ( .A1(n4485), .A2(n4484), .ZN(n6846) );
  AND2_X1 U6848 ( .A1(n4480), .A2(n6847), .ZN(n6845) );
  OR2_X1 U6849 ( .A1(n4484), .A2(n4485), .ZN(n6847) );
  OR2_X1 U6850 ( .A1(n4036), .A2(n3888), .ZN(n4485) );
  OR2_X1 U6851 ( .A1(n6848), .A2(n6849), .ZN(n4484) );
  AND2_X1 U6852 ( .A1(n6827), .A2(n6826), .ZN(n6849) );
  AND2_X1 U6853 ( .A1(n6822), .A2(n6850), .ZN(n6848) );
  OR2_X1 U6854 ( .A1(n6826), .A2(n6827), .ZN(n6850) );
  OR2_X1 U6855 ( .A1(n4036), .A2(n4047), .ZN(n6827) );
  OR2_X1 U6856 ( .A1(n6851), .A2(n6852), .ZN(n6826) );
  AND2_X1 U6857 ( .A1(n6816), .A2(n6815), .ZN(n6852) );
  AND2_X1 U6858 ( .A1(n6811), .A2(n6853), .ZN(n6851) );
  OR2_X1 U6859 ( .A1(n6815), .A2(n6816), .ZN(n6853) );
  OR2_X1 U6860 ( .A1(n3837), .A2(n4036), .ZN(n6816) );
  OR2_X1 U6861 ( .A1(n6854), .A2(n6855), .ZN(n6815) );
  AND2_X1 U6862 ( .A1(n6805), .A2(n6804), .ZN(n6855) );
  AND2_X1 U6863 ( .A1(n6800), .A2(n6856), .ZN(n6854) );
  OR2_X1 U6864 ( .A1(n6804), .A2(n6805), .ZN(n6856) );
  OR2_X1 U6865 ( .A1(n4053), .A2(n4036), .ZN(n6805) );
  OR2_X1 U6866 ( .A1(n6857), .A2(n6858), .ZN(n6804) );
  AND2_X1 U6867 ( .A1(n6794), .A2(n6793), .ZN(n6858) );
  AND2_X1 U6868 ( .A1(n6789), .A2(n6859), .ZN(n6857) );
  OR2_X1 U6869 ( .A1(n6793), .A2(n6794), .ZN(n6859) );
  OR2_X1 U6870 ( .A1(n3786), .A2(n4036), .ZN(n6794) );
  OR2_X1 U6871 ( .A1(n6860), .A2(n6861), .ZN(n6793) );
  AND2_X1 U6872 ( .A1(n6784), .A2(n6782), .ZN(n6861) );
  AND2_X1 U6873 ( .A1(n6778), .A2(n6862), .ZN(n6860) );
  OR2_X1 U6874 ( .A1(n6782), .A2(n6784), .ZN(n6862) );
  INV_X1 U6875 ( .A(n6781), .ZN(n6784) );
  AND2_X1 U6876 ( .A1(a_10_), .A2(b_2_), .ZN(n6781) );
  OR2_X1 U6877 ( .A1(n6863), .A2(n6864), .ZN(n6782) );
  AND2_X1 U6878 ( .A1(n6767), .A2(n6770), .ZN(n6864) );
  AND2_X1 U6879 ( .A1(n6865), .A2(n6772), .ZN(n6863) );
  OR2_X1 U6880 ( .A1(n6866), .A2(n6867), .ZN(n6772) );
  AND2_X1 U6881 ( .A1(n6761), .A2(n6760), .ZN(n6867) );
  AND2_X1 U6882 ( .A1(n6756), .A2(n6868), .ZN(n6866) );
  OR2_X1 U6883 ( .A1(n6760), .A2(n6761), .ZN(n6868) );
  OR2_X1 U6884 ( .A1(n4072), .A2(n4036), .ZN(n6761) );
  OR2_X1 U6885 ( .A1(n6869), .A2(n6870), .ZN(n6760) );
  AND2_X1 U6886 ( .A1(n6744), .A2(n6750), .ZN(n6870) );
  AND2_X1 U6887 ( .A1(n6751), .A2(n6871), .ZN(n6869) );
  OR2_X1 U6888 ( .A1(n6750), .A2(n6744), .ZN(n6871) );
  OR2_X1 U6889 ( .A1(n3682), .A2(n4036), .ZN(n6744) );
  OR2_X1 U6890 ( .A1(n3998), .A2(n6872), .ZN(n6750) );
  OR2_X1 U6891 ( .A1(n4070), .A2(n4036), .ZN(n6872) );
  INV_X1 U6892 ( .A(n6749), .ZN(n6751) );
  OR2_X1 U6893 ( .A1(n6873), .A2(n6874), .ZN(n6749) );
  AND2_X1 U6894 ( .A1(b_1_), .A2(n6875), .ZN(n6874) );
  OR2_X1 U6895 ( .A1(n6876), .A2(n3644), .ZN(n6875) );
  AND2_X1 U6896 ( .A1(n3628), .A2(a_14_), .ZN(n3644) );
  AND2_X1 U6897 ( .A1(a_14_), .A2(n4029), .ZN(n6876) );
  AND2_X1 U6898 ( .A1(b_0_), .A2(n6877), .ZN(n6873) );
  OR2_X1 U6899 ( .A1(n6878), .A2(n3647), .ZN(n6877) );
  AND2_X1 U6900 ( .A1(n3639), .A2(a_15_), .ZN(n3647) );
  AND2_X1 U6901 ( .A1(a_15_), .A2(n3998), .ZN(n6878) );
  AND2_X1 U6902 ( .A1(n6879), .A2(n6880), .ZN(n6756) );
  INV_X1 U6903 ( .A(n6881), .ZN(n6880) );
  AND2_X1 U6904 ( .A1(n6882), .A2(n6883), .ZN(n6881) );
  OR2_X1 U6905 ( .A1(n6883), .A2(n6882), .ZN(n6879) );
  OR2_X1 U6906 ( .A1(n6884), .A2(n6885), .ZN(n6882) );
  AND2_X1 U6907 ( .A1(n6886), .A2(n6887), .ZN(n6885) );
  AND2_X1 U6908 ( .A1(b_0_), .A2(a_14_), .ZN(n6886) );
  AND2_X1 U6909 ( .A1(n6888), .A2(n6889), .ZN(n6884) );
  OR2_X1 U6910 ( .A1(n3639), .A2(n4029), .ZN(n6889) );
  INV_X1 U6911 ( .A(n6887), .ZN(n6888) );
  OR2_X1 U6912 ( .A1(n3682), .A2(n3998), .ZN(n6887) );
  OR2_X1 U6913 ( .A1(n6770), .A2(n6767), .ZN(n6865) );
  OR2_X1 U6914 ( .A1(n6890), .A2(n6891), .ZN(n6767) );
  AND2_X1 U6915 ( .A1(n6892), .A2(n6893), .ZN(n6891) );
  INV_X1 U6916 ( .A(n6894), .ZN(n6890) );
  OR2_X1 U6917 ( .A1(n6892), .A2(n6893), .ZN(n6894) );
  OR2_X1 U6918 ( .A1(n6895), .A2(n6896), .ZN(n6892) );
  AND2_X1 U6919 ( .A1(n6897), .A2(n6898), .ZN(n6896) );
  INV_X1 U6920 ( .A(n6899), .ZN(n6895) );
  OR2_X1 U6921 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  OR2_X1 U6922 ( .A1(n3735), .A2(n4036), .ZN(n6770) );
  INV_X1 U6923 ( .A(b_2_), .ZN(n4036) );
  AND2_X1 U6924 ( .A1(n6900), .A2(n6901), .ZN(n6778) );
  INV_X1 U6925 ( .A(n6902), .ZN(n6901) );
  AND2_X1 U6926 ( .A1(n6903), .A2(n6904), .ZN(n6902) );
  OR2_X1 U6927 ( .A1(n6903), .A2(n6904), .ZN(n6900) );
  OR2_X1 U6928 ( .A1(n6905), .A2(n6906), .ZN(n6903) );
  INV_X1 U6929 ( .A(n6907), .ZN(n6906) );
  OR2_X1 U6930 ( .A1(n6908), .A2(n6909), .ZN(n6907) );
  AND2_X1 U6931 ( .A1(n6909), .A2(n6908), .ZN(n6905) );
  AND2_X1 U6932 ( .A1(n6910), .A2(n6911), .ZN(n6789) );
  INV_X1 U6933 ( .A(n6912), .ZN(n6911) );
  AND2_X1 U6934 ( .A1(n6913), .A2(n6914), .ZN(n6912) );
  OR2_X1 U6935 ( .A1(n6913), .A2(n6914), .ZN(n6910) );
  OR2_X1 U6936 ( .A1(n6915), .A2(n6916), .ZN(n6913) );
  INV_X1 U6937 ( .A(n6917), .ZN(n6916) );
  OR2_X1 U6938 ( .A1(n6918), .A2(n6919), .ZN(n6917) );
  AND2_X1 U6939 ( .A1(n6919), .A2(n6918), .ZN(n6915) );
  AND2_X1 U6940 ( .A1(n6920), .A2(n6921), .ZN(n6800) );
  INV_X1 U6941 ( .A(n6922), .ZN(n6921) );
  AND2_X1 U6942 ( .A1(n6923), .A2(n6924), .ZN(n6922) );
  OR2_X1 U6943 ( .A1(n6923), .A2(n6924), .ZN(n6920) );
  OR2_X1 U6944 ( .A1(n6925), .A2(n6926), .ZN(n6923) );
  INV_X1 U6945 ( .A(n6927), .ZN(n6926) );
  OR2_X1 U6946 ( .A1(n6928), .A2(n6929), .ZN(n6927) );
  AND2_X1 U6947 ( .A1(n6929), .A2(n6928), .ZN(n6925) );
  AND2_X1 U6948 ( .A1(n6930), .A2(n6931), .ZN(n6811) );
  INV_X1 U6949 ( .A(n6932), .ZN(n6931) );
  AND2_X1 U6950 ( .A1(n6933), .A2(n6934), .ZN(n6932) );
  OR2_X1 U6951 ( .A1(n6933), .A2(n6934), .ZN(n6930) );
  OR2_X1 U6952 ( .A1(n6935), .A2(n6936), .ZN(n6933) );
  INV_X1 U6953 ( .A(n6937), .ZN(n6936) );
  OR2_X1 U6954 ( .A1(n6938), .A2(n6939), .ZN(n6937) );
  AND2_X1 U6955 ( .A1(n6939), .A2(n6938), .ZN(n6935) );
  AND2_X1 U6956 ( .A1(n6940), .A2(n6941), .ZN(n6822) );
  INV_X1 U6957 ( .A(n6942), .ZN(n6941) );
  AND2_X1 U6958 ( .A1(n6943), .A2(n6944), .ZN(n6942) );
  OR2_X1 U6959 ( .A1(n6943), .A2(n6944), .ZN(n6940) );
  OR2_X1 U6960 ( .A1(n6945), .A2(n6946), .ZN(n6943) );
  INV_X1 U6961 ( .A(n6947), .ZN(n6946) );
  OR2_X1 U6962 ( .A1(n6948), .A2(n6949), .ZN(n6947) );
  AND2_X1 U6963 ( .A1(n6949), .A2(n6948), .ZN(n6945) );
  AND2_X1 U6964 ( .A1(n6950), .A2(n6951), .ZN(n4480) );
  INV_X1 U6965 ( .A(n6952), .ZN(n6951) );
  AND2_X1 U6966 ( .A1(n6953), .A2(n6954), .ZN(n6952) );
  OR2_X1 U6967 ( .A1(n6953), .A2(n6954), .ZN(n6950) );
  OR2_X1 U6968 ( .A1(n6955), .A2(n6956), .ZN(n6953) );
  INV_X1 U6969 ( .A(n6957), .ZN(n6956) );
  OR2_X1 U6970 ( .A1(n6958), .A2(n6959), .ZN(n6957) );
  AND2_X1 U6971 ( .A1(n6959), .A2(n6958), .ZN(n6955) );
  AND2_X1 U6972 ( .A1(n6960), .A2(n6961), .ZN(n4391) );
  INV_X1 U6973 ( .A(n6962), .ZN(n6961) );
  AND2_X1 U6974 ( .A1(n6963), .A2(n6964), .ZN(n6962) );
  OR2_X1 U6975 ( .A1(n6963), .A2(n6964), .ZN(n6960) );
  OR2_X1 U6976 ( .A1(n6965), .A2(n6966), .ZN(n6963) );
  INV_X1 U6977 ( .A(n6967), .ZN(n6966) );
  OR2_X1 U6978 ( .A1(n6968), .A2(n6969), .ZN(n6967) );
  AND2_X1 U6979 ( .A1(n6969), .A2(n6968), .ZN(n6965) );
  AND2_X1 U6980 ( .A1(n6970), .A2(n6971), .ZN(n4309) );
  INV_X1 U6981 ( .A(n6972), .ZN(n6971) );
  AND2_X1 U6982 ( .A1(n6973), .A2(n6974), .ZN(n6972) );
  OR2_X1 U6983 ( .A1(n6973), .A2(n6974), .ZN(n6970) );
  OR2_X1 U6984 ( .A1(n6975), .A2(n6976), .ZN(n6973) );
  INV_X1 U6985 ( .A(n6977), .ZN(n6976) );
  OR2_X1 U6986 ( .A1(n6978), .A2(n6979), .ZN(n6977) );
  AND2_X1 U6987 ( .A1(n6979), .A2(n6978), .ZN(n6975) );
  AND2_X1 U6988 ( .A1(n6980), .A2(n6981), .ZN(n4250) );
  INV_X1 U6989 ( .A(n6982), .ZN(n6981) );
  AND2_X1 U6990 ( .A1(n6983), .A2(n6984), .ZN(n6982) );
  OR2_X1 U6991 ( .A1(n6983), .A2(n6984), .ZN(n6980) );
  OR2_X1 U6992 ( .A1(n6985), .A2(n6986), .ZN(n6983) );
  INV_X1 U6993 ( .A(n6987), .ZN(n6986) );
  OR2_X1 U6994 ( .A1(n6988), .A2(n6989), .ZN(n6987) );
  AND2_X1 U6995 ( .A1(n6989), .A2(n6988), .ZN(n6985) );
  AND2_X1 U6996 ( .A1(n6990), .A2(n6991), .ZN(n4195) );
  INV_X1 U6997 ( .A(n6992), .ZN(n6991) );
  AND2_X1 U6998 ( .A1(n6993), .A2(n6994), .ZN(n6992) );
  OR2_X1 U6999 ( .A1(n6993), .A2(n6994), .ZN(n6990) );
  OR2_X1 U7000 ( .A1(n6995), .A2(n6996), .ZN(n6993) );
  INV_X1 U7001 ( .A(n6997), .ZN(n6996) );
  OR2_X1 U7002 ( .A1(n6998), .A2(n6999), .ZN(n6997) );
  AND2_X1 U7003 ( .A1(n6999), .A2(n6998), .ZN(n6995) );
  INV_X1 U7004 ( .A(n4162), .ZN(n4160) );
  OR2_X1 U7005 ( .A1(n7000), .A2(n7001), .ZN(n4162) );
  AND2_X1 U7006 ( .A1(n7002), .A2(n7003), .ZN(n7001) );
  INV_X1 U7007 ( .A(n7004), .ZN(n7000) );
  OR2_X1 U7008 ( .A1(n7002), .A2(n7003), .ZN(n7004) );
  OR2_X1 U7009 ( .A1(n7005), .A2(n7006), .ZN(n7002) );
  AND2_X1 U7010 ( .A1(n7007), .A2(n4033), .ZN(n7006) );
  INV_X1 U7011 ( .A(n7008), .ZN(n7007) );
  AND2_X1 U7012 ( .A1(n4005), .A2(n7008), .ZN(n7005) );
  INV_X1 U7013 ( .A(n4033), .ZN(n4005) );
  AND2_X1 U7014 ( .A1(n7009), .A2(n7010), .ZN(n4139) );
  INV_X1 U7015 ( .A(n7011), .ZN(n7010) );
  AND2_X1 U7016 ( .A1(n7012), .A2(n7013), .ZN(n7011) );
  OR2_X1 U7017 ( .A1(n7012), .A2(n7013), .ZN(n7009) );
  OR2_X1 U7018 ( .A1(n7014), .A2(n7015), .ZN(n7012) );
  AND2_X1 U7019 ( .A1(n7016), .A2(n7017), .ZN(n7015) );
  INV_X1 U7020 ( .A(n7018), .ZN(n7014) );
  OR2_X1 U7021 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  INV_X1 U7022 ( .A(n7019), .ZN(n7016) );
  OR2_X1 U7023 ( .A1(n7020), .A2(n7021), .ZN(n3924) );
  INV_X1 U7024 ( .A(n7022), .ZN(n7021) );
  OR2_X1 U7025 ( .A1(n7023), .A2(n7024), .ZN(n7022) );
  AND2_X1 U7026 ( .A1(n7024), .A2(n7023), .ZN(n7020) );
  OR2_X1 U7027 ( .A1(n4029), .A2(n4028), .ZN(n7023) );
  AND2_X1 U7028 ( .A1(n7024), .A2(a_0_), .ZN(n4134) );
  INV_X1 U7029 ( .A(n7025), .ZN(n7024) );
  OR2_X1 U7030 ( .A1(n7026), .A2(n7027), .ZN(n7025) );
  AND2_X1 U7031 ( .A1(n7013), .A2(n7019), .ZN(n7027) );
  AND2_X1 U7032 ( .A1(n7028), .A2(n7017), .ZN(n7026) );
  OR2_X1 U7033 ( .A1(n3998), .A2(n4028), .ZN(n7017) );
  INV_X1 U7034 ( .A(a_0_), .ZN(n4028) );
  OR2_X1 U7035 ( .A1(n7019), .A2(n7013), .ZN(n7028) );
  OR2_X1 U7036 ( .A1(n4029), .A2(n4002), .ZN(n7013) );
  OR2_X1 U7037 ( .A1(n7029), .A2(n7030), .ZN(n7019) );
  AND2_X1 U7038 ( .A1(n7003), .A2(n7008), .ZN(n7030) );
  AND2_X1 U7039 ( .A1(n7031), .A2(n4033), .ZN(n7029) );
  OR2_X1 U7040 ( .A1(n3998), .A2(n4002), .ZN(n4033) );
  INV_X1 U7041 ( .A(a_1_), .ZN(n4002) );
  OR2_X1 U7042 ( .A1(n7008), .A2(n7003), .ZN(n7031) );
  OR2_X1 U7043 ( .A1(n4029), .A2(n4035), .ZN(n7003) );
  OR2_X1 U7044 ( .A1(n7032), .A2(n7033), .ZN(n7008) );
  AND2_X1 U7045 ( .A1(n6994), .A2(n6998), .ZN(n7033) );
  AND2_X1 U7046 ( .A1(n7034), .A2(n7035), .ZN(n7032) );
  INV_X1 U7047 ( .A(n6999), .ZN(n7035) );
  AND2_X1 U7048 ( .A1(b_0_), .A2(a_3_), .ZN(n6999) );
  OR2_X1 U7049 ( .A1(n6998), .A2(n6994), .ZN(n7034) );
  OR2_X1 U7050 ( .A1(n3998), .A2(n4035), .ZN(n6994) );
  INV_X1 U7051 ( .A(a_2_), .ZN(n4035) );
  OR2_X1 U7052 ( .A1(n7036), .A2(n7037), .ZN(n6998) );
  AND2_X1 U7053 ( .A1(n6984), .A2(n6988), .ZN(n7037) );
  AND2_X1 U7054 ( .A1(n7038), .A2(n7039), .ZN(n7036) );
  INV_X1 U7055 ( .A(n6989), .ZN(n7039) );
  AND2_X1 U7056 ( .A1(b_0_), .A2(a_4_), .ZN(n6989) );
  OR2_X1 U7057 ( .A1(n6988), .A2(n6984), .ZN(n7038) );
  OR2_X1 U7058 ( .A1(n3998), .A2(n3951), .ZN(n6984) );
  INV_X1 U7059 ( .A(a_3_), .ZN(n3951) );
  OR2_X1 U7060 ( .A1(n7040), .A2(n7041), .ZN(n6988) );
  AND2_X1 U7061 ( .A1(n6974), .A2(n6978), .ZN(n7041) );
  AND2_X1 U7062 ( .A1(n7042), .A2(n7043), .ZN(n7040) );
  INV_X1 U7063 ( .A(n6979), .ZN(n7043) );
  AND2_X1 U7064 ( .A1(a_5_), .A2(b_0_), .ZN(n6979) );
  OR2_X1 U7065 ( .A1(n6978), .A2(n6974), .ZN(n7042) );
  OR2_X1 U7066 ( .A1(n3998), .A2(n4041), .ZN(n6974) );
  INV_X1 U7067 ( .A(a_4_), .ZN(n4041) );
  OR2_X1 U7068 ( .A1(n7044), .A2(n7045), .ZN(n6978) );
  AND2_X1 U7069 ( .A1(n6964), .A2(n6968), .ZN(n7045) );
  AND2_X1 U7070 ( .A1(n7046), .A2(n7047), .ZN(n7044) );
  INV_X1 U7071 ( .A(n6969), .ZN(n7047) );
  AND2_X1 U7072 ( .A1(a_6_), .A2(b_0_), .ZN(n6969) );
  OR2_X1 U7073 ( .A1(n6968), .A2(n6964), .ZN(n7046) );
  OR2_X1 U7074 ( .A1(n3998), .A2(n3888), .ZN(n6964) );
  INV_X1 U7075 ( .A(a_5_), .ZN(n3888) );
  OR2_X1 U7076 ( .A1(n7048), .A2(n7049), .ZN(n6968) );
  AND2_X1 U7077 ( .A1(n6954), .A2(n6958), .ZN(n7049) );
  AND2_X1 U7078 ( .A1(n7050), .A2(n7051), .ZN(n7048) );
  INV_X1 U7079 ( .A(n6959), .ZN(n7051) );
  AND2_X1 U7080 ( .A1(a_7_), .A2(b_0_), .ZN(n6959) );
  OR2_X1 U7081 ( .A1(n6958), .A2(n6954), .ZN(n7050) );
  OR2_X1 U7082 ( .A1(n4047), .A2(n3998), .ZN(n6954) );
  INV_X1 U7083 ( .A(a_6_), .ZN(n4047) );
  OR2_X1 U7084 ( .A1(n7052), .A2(n7053), .ZN(n6958) );
  AND2_X1 U7085 ( .A1(n6944), .A2(n6948), .ZN(n7053) );
  AND2_X1 U7086 ( .A1(n7054), .A2(n7055), .ZN(n7052) );
  INV_X1 U7087 ( .A(n6949), .ZN(n7055) );
  AND2_X1 U7088 ( .A1(a_8_), .A2(b_0_), .ZN(n6949) );
  OR2_X1 U7089 ( .A1(n6948), .A2(n6944), .ZN(n7054) );
  OR2_X1 U7090 ( .A1(n3837), .A2(n3998), .ZN(n6944) );
  INV_X1 U7091 ( .A(a_7_), .ZN(n3837) );
  OR2_X1 U7092 ( .A1(n7056), .A2(n7057), .ZN(n6948) );
  AND2_X1 U7093 ( .A1(n6934), .A2(n6938), .ZN(n7057) );
  AND2_X1 U7094 ( .A1(n7058), .A2(n7059), .ZN(n7056) );
  INV_X1 U7095 ( .A(n6939), .ZN(n7059) );
  AND2_X1 U7096 ( .A1(a_9_), .A2(b_0_), .ZN(n6939) );
  OR2_X1 U7097 ( .A1(n6938), .A2(n6934), .ZN(n7058) );
  OR2_X1 U7098 ( .A1(n4053), .A2(n3998), .ZN(n6934) );
  INV_X1 U7099 ( .A(a_8_), .ZN(n4053) );
  OR2_X1 U7100 ( .A1(n7060), .A2(n7061), .ZN(n6938) );
  AND2_X1 U7101 ( .A1(n6924), .A2(n6928), .ZN(n7061) );
  AND2_X1 U7102 ( .A1(n7062), .A2(n7063), .ZN(n7060) );
  INV_X1 U7103 ( .A(n6929), .ZN(n7063) );
  AND2_X1 U7104 ( .A1(a_10_), .A2(b_0_), .ZN(n6929) );
  OR2_X1 U7105 ( .A1(n6928), .A2(n6924), .ZN(n7062) );
  OR2_X1 U7106 ( .A1(n3786), .A2(n3998), .ZN(n6924) );
  INV_X1 U7107 ( .A(a_9_), .ZN(n3786) );
  OR2_X1 U7108 ( .A1(n7064), .A2(n7065), .ZN(n6928) );
  AND2_X1 U7109 ( .A1(n6914), .A2(n6918), .ZN(n7065) );
  AND2_X1 U7110 ( .A1(n7066), .A2(n7067), .ZN(n7064) );
  INV_X1 U7111 ( .A(n6919), .ZN(n7067) );
  AND2_X1 U7112 ( .A1(a_11_), .A2(b_0_), .ZN(n6919) );
  OR2_X1 U7113 ( .A1(n6918), .A2(n6914), .ZN(n7066) );
  OR2_X1 U7114 ( .A1(n4059), .A2(n3998), .ZN(n6914) );
  INV_X1 U7115 ( .A(a_10_), .ZN(n4059) );
  OR2_X1 U7116 ( .A1(n7068), .A2(n7069), .ZN(n6918) );
  AND2_X1 U7117 ( .A1(n6904), .A2(n6908), .ZN(n7069) );
  AND2_X1 U7118 ( .A1(n7070), .A2(n7071), .ZN(n7068) );
  INV_X1 U7119 ( .A(n6909), .ZN(n7071) );
  AND2_X1 U7120 ( .A1(a_12_), .A2(b_0_), .ZN(n6909) );
  OR2_X1 U7121 ( .A1(n6908), .A2(n6904), .ZN(n7070) );
  OR2_X1 U7122 ( .A1(n3735), .A2(n3998), .ZN(n6904) );
  INV_X1 U7123 ( .A(a_11_), .ZN(n3735) );
  OR2_X1 U7124 ( .A1(n7072), .A2(n7073), .ZN(n6908) );
  AND2_X1 U7125 ( .A1(n6893), .A2(n6898), .ZN(n7073) );
  AND2_X1 U7126 ( .A1(n6897), .A2(n7074), .ZN(n7072) );
  OR2_X1 U7127 ( .A1(n6898), .A2(n6893), .ZN(n7074) );
  OR2_X1 U7128 ( .A1(n4072), .A2(n3998), .ZN(n6893) );
  INV_X1 U7129 ( .A(a_12_), .ZN(n4072) );
  AND2_X1 U7130 ( .A1(n7075), .A2(n6883), .ZN(n6897) );
  OR2_X1 U7131 ( .A1(n4029), .A2(n7076), .ZN(n6883) );
  OR2_X1 U7132 ( .A1(n4070), .A2(n3998), .ZN(n7076) );
  OR2_X1 U7133 ( .A1(n3628), .A2(n3639), .ZN(n4070) );
  INV_X1 U7134 ( .A(a_15_), .ZN(n3628) );
  OR2_X1 U7135 ( .A1(n7077), .A2(n6898), .ZN(n7075) );
  OR2_X1 U7136 ( .A1(n3682), .A2(n4029), .ZN(n6898) );
  INV_X1 U7137 ( .A(b_0_), .ZN(n4029) );
  INV_X1 U7138 ( .A(a_13_), .ZN(n3682) );
  OR2_X1 U7139 ( .A1(n3998), .A2(n3639), .ZN(n7077) );
  INV_X1 U7140 ( .A(a_14_), .ZN(n3639) );
  INV_X1 U7141 ( .A(b_1_), .ZN(n3998) );
endmodule

