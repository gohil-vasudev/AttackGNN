module s38417 ( CK, g1249, g16297, g16355, g16399, g16437, g16496, g1943, 
        g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g2637, 
        g27380, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, 
        g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, 
        g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, 
        g4450, g4590, g51, g5388, g5437, g5472, g5511, g5549, g5555, g5595, 
        g5612, g5629, g563, g5637, g5648, g5657, g5686, g5695, g5738, g5747, 
        g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, 
        g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, 
        g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, 
        g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, 
        g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, 
        g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, 
        g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, test_se, 
        test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, 
        test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, 
        test_si8, test_so8, test_si9, test_so9, test_si10, test_so10, 
        test_si11, test_so11, test_si12, test_so12, test_si13, test_so13, 
        test_si14, test_so14, test_si15, test_so15, test_si16, test_so16, 
        test_si17, test_so17, test_si18, test_so18, test_si19, test_so19, 
        test_si20, test_so20, test_si21, test_so21, test_si22, test_so22, 
        test_si23, test_so23, test_si24, test_so24, test_si25, test_so25, 
        test_si26, test_so26, test_si27, test_so27, test_si28, test_so28, 
        test_si29, test_so29, test_si30, test_so30, test_si31, test_so31, 
        test_si32, test_so32, test_si33, test_so33, test_si34, test_so34, 
        test_si35, test_so35, test_si36, test_so36, test_si37, test_so37, 
        test_si38, test_so38, test_si39, test_so39, test_si40, test_so40, 
        test_si41, test_so41, test_si42, test_so42, test_si43, test_so43, 
        test_si44, test_so44, test_si45, test_so45, test_si46, test_so46, 
        test_si47, test_so47, test_si48, test_so48, test_si49, test_so49, 
        test_si50, test_so50, test_si51, test_so51, test_si52, test_so52, 
        test_si53, test_so53, test_si54, test_so54, test_si55, test_so55, 
        test_si56, test_so56, test_si57, test_so57, test_si58, test_so58, 
        test_si59, test_so59, test_si60, test_so60, test_si61, test_so61, 
        test_si62, test_so62, test_si63, test_so63, test_si64, test_so64, 
        test_si65, test_so65, test_si66, test_so66, test_si67, test_so67, 
        test_si68, test_so68, test_si69, test_so69, test_si70, test_so70, 
        test_si71, test_so71, test_si72, test_so72, test_si73, test_so73, 
        test_si74, test_so74, test_si75, test_so75, test_si76, test_so76, 
        test_si77, test_so77, test_si78, test_so78, test_si79, test_so79, 
        test_si80, test_so80, test_si81, test_so81, test_si82, test_so82, 
        test_si83, test_so83, test_si84, test_so84, test_si85, test_so85, 
        test_si86, test_so86, test_si87, test_so87, test_si88, test_so88, 
        test_si89, test_so89, test_si90, test_so90, test_si91, test_so91, 
        test_si92, test_so92, test_si93, test_so93, test_si94, test_so94, 
        test_si95, test_so95, test_si96, test_so96, test_si97, test_so97, 
        test_si98, test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217,
         g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227,
         g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;
  output g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275,
         test_so1, test_so2, test_so3, test_so4, test_so5, test_so6, test_so7,
         test_so8, test_so9, test_so10, test_so11, test_so12, test_so13,
         test_so14, test_so15, test_so16, test_so17, test_so18, test_so19,
         test_so20, test_so21, test_so22, test_so23, test_so24, test_so25,
         test_so26, test_so27, test_so28, test_so29, test_so30, test_so31,
         test_so32, test_so33, test_so34, test_so35, test_so36, test_so37,
         test_so38, test_so39, test_so40, test_so41, test_so42, test_so43,
         test_so44, test_so45, test_so46, test_so47, test_so48, test_so49,
         test_so50, test_so51, test_so52, test_so53, test_so54, test_so55,
         test_so56, test_so57, test_so58, test_so59, test_so60, test_so61,
         test_so62, test_so63, test_so64, test_so65, test_so66, test_so67,
         test_so68, test_so69, test_so70, test_so71, test_so72, test_so73,
         test_so74, test_so75, test_so76, test_so77, test_so78, test_so79,
         test_so80, test_so81, test_so82, test_so83, test_so84, test_so85,
         test_so86, test_so87, test_so88, test_so89, test_so90, test_so91,
         test_so92, test_so93, test_so94, test_so95, test_so96, test_so97,
         test_so98, test_so99, test_so100;
  wire   test_so3, test_so4, test_so5, test_so23, test_so57, test_so63,
         test_so73, test_so99, test_so100, n2230, n2217, n2231, n2374, n2361,
         n2375, DFF_2_n1, n4264, n2445, n2446, n2440, n2426, n2670, n2671,
         n2669, n2685, n2686, n2684, n2718, n2719, n2717, g2124, n2981, g1430,
         n2984, g744, n2987, g56, n2990, n3741, n8104, g16802, n8103, g16823,
         n8102, g2950, n4423, g2883, n4330, g22026, g2888, g23358, g2896,
         n4431, g24473, g2892, g25201, g2903, n4305, g26037, g2900, n4291,
         g26798, g2908, n4355, n4273, g2912, n4482, g23357, g2917, n4479,
         g24476, g2924, n4349, g25199, g2920, n4280, n4281, n8099, n8098,
         DFF_18_n1, n4279, g2879, n4351, g2934, g2935, g2938, g2941, g2944,
         g2947, g2953, g2956, g2959, g2962, g2963, g2969, g2972, g2975, g2978,
         g2981, g2874, g18754, g1506, n4288, g18781, g1501, n4565, g18803,
         g1496, n4557, g18821, g1491, n4326, g18835, g1486, n4390, g18852,
         g1481, n4320, g18866, g1476, n4374, g18883, g1471, n4378, g21880,
         g2877, g19154, g813, n4289, g19163, g809, n4567, g19173, g805, n4559,
         g19184, g801, n4327, g20310, g797, n4391, g20343, g793, n4321, g20376,
         g789, n4375, g20417, g785, n4379, g21878, g2873, g19153, g125, n4290,
         g19162, g121, n4569, g19172, g117, n4561, g19144, g113, n4328, g19149,
         g109, n4392, g19157, g105, n4322, g19167, g101, n4376, g19178, g97,
         n4380, g20874, g2857, g18885, g2200, n4287, g18975, g2195, n4563,
         g18968, g2190, n4555, g18942, g2185, n4325, g18906, g2180, n4389,
         g18867, g2175, n4319, g18836, g2170, n4373, g18957, g2165, n4377,
         g21882, g2878, n4598, n4382, n4383, g3109, n4494, g18669, g18719,
         g3211, g18782, g3084, g17222, g3085, g17225, g3086, g17234, g3087,
         g17224, g3091, g17228, g3092, g17246, g3093, g17226, g3094, g17235,
         g3095, g17269, g3096, g25450, g3097, g25451, g3098, g25452, g3099,
         g28420, g3100, g28421, g28425, g3102, g29936, g3103, g29939, g3104,
         g29941, g3105, g30796, g3106, g30798, g3107, g30801, g3108, g17229,
         g3155, g17247, g3158, g17302, g3161, g17236, g3164, g17270, g3167,
         g17340, g3170, g17248, g3173, g17303, g3176, g17383, g17271, g3182,
         g17341, g3185, g17429, g3088, n8090, n8089, g3197, n8088, g3201,
         n4406, g3204, g3207, n4329, g3188, n4405, g3133, n8087, g3128, n8086,
         n8084, DFF_144_n1, g3124, n8083, DFF_146_n1, n8082, n8081, n8080,
         g3112, g3110, g3111, n8079, n8078, n8077, n8076, g3151, n4424, g3142,
         n4301, g185, n4384, n4318, n4512, g165, n4369, g22100, g130, g22122,
         g131, g22141, g129, g22123, g133, g22142, g134, g22161, g132, g22025,
         g142, g22027, g143, g22030, g141, g22028, g145, g22031, g146, g22037,
         g22032, g148, g22038, g149, g22047, g147, g22039, g151, g22048, g152,
         g22063, g150, g22049, g154, g22064, g155, g22079, g153, g22065, g157,
         g22080, g158, g22101, g156, g22081, g160, g22102, g161, g22124, g159,
         g22103, g22125, g164, g22143, g162, g25204, g169, g25206, g170,
         g25211, g168, g25207, g172, g25212, g173, g25218, g171, g25213, g175,
         g25219, g176, g25228, g174, g25220, g178, g25229, g179, g25239, g177,
         g30261, g186, g30267, g30275, g192, g30637, g231, g30640, g234,
         g30645, g237, g30668, g195, g30674, g198, g30680, g201, g30641, g240,
         g30646, g243, g30653, g246, g30276, g204, g30284, g207, g30292, g210,
         g30254, g249, g30257, g252, g30262, g30245, g213, g30246, g216,
         g30248, g219, g30258, g258, g30263, g261, g30268, g264, g30635, g222,
         g30636, g225, g30639, g228, g30661, g267, g30669, g270, g30675, g273,
         g25027, g92, g25932, g88, g26529, g83, g27120, g27594, g74, g28145,
         g70, g28634, g65, g29109, g61, g29353, g29579, g52, g180, g181, n4506,
         g309, n4388, g27253, g354, g27255, g343, g27258, g27256, g369, g27259,
         g358, g27265, g361, g27260, g384, g27266, g373, g27277, g376, g27267,
         g398, g27278, g388, g27293, g391, g28732, g408, g28735, g411, g28744,
         g414, g29194, g417, g29197, g420, g29201, g423, g28736, g28745, g428,
         g28754, g426, g26803, g429, g26804, g432, g26807, g435, g26805, g438,
         g26808, g441, g26812, g444, g27759, g448, g27760, g449, g27762, g447,
         g29606, g312, g29608, g313, g29611, g314, g30699, g315, g30700,
         g30702, g317, g30455, g318, g30468, g319, g30482, g320, g29167, g322,
         g29169, g323, g29172, g321, g26655, g403, g26659, g404, g26664, g402,
         g450, n8066, DFF_299_n1, g452, n8065, DFF_301_n1, g454, DFF_303_n1,
         g280, n8062, DFF_305_n1, g282, n8061, DFF_307_n1, g284, n8060,
         DFF_309_n1, g286, n8059, DFF_311_n1, g288, n8058, DFF_313_n1, g290,
         n8057, n4485, n4282, n8056, g21346, g305, n4278, n8055, DFF_328_n1,
         g349, g350, g351, g352, g353, g357, g364, g365, g366, g367, g368,
         g372, g379, g380, g381, g383, g387, g394, g395, g396, g397, g324,
         g337, n4298, n4372, g550, n4313, g21842, g554, g18678, g557, n4360,
         g18726, g513, g523, g524, g455, g564, g569, g458, g570, g571, g461,
         g572, g573, g465, g574, g565, g566, g567, g471, g568, g489, n4461,
         g485, n4466, g23067, g486, g23093, g487, g23117, g488, g23385, g23399,
         g24174, g24178, g477, g24207, g478, g24216, g479, g23092, g480,
         g23000, g484, g23022, g464, g24206, g24215, g24228, g528, g535, g542,
         g13149, g543, g544, g21851, g548, g13111, g549, g499, n4541, g13160,
         g558, g559, g27261, g576, g27268, g577, g27279, g575, g27269, g579,
         g27280, g27294, g578, g27281, g582, g27295, g583, g27311, g581,
         g27296, g585, g27312, g586, g27327, g584, g24491, g587, g24498, g590,
         g24507, g593, g24499, g596, g24508, g599, g24519, g602, g28345, g614,
         g28349, g617, g28353, g28342, g605, g28344, g608, g28348, g611,
         g26541, g490, g26545, g493, g26553, g496, g506, n4570, g22578, n4571,
         g525, n8047, n8046, n8045, n8044, n8043, g536, g537, g24059, g538,
         n4492, n8040, n4359, g629, n4295, g16654, g630, g20314, g659, n4429,
         g20682, g640, n4404, g23136, g633, n4478, g23324, g653, n4422, g24426,
         g646, n4414, g25185, g660, n4403, g26660, g672, n4413, g26776, g27672,
         g679, n4477, g28199, g686, n4396, g28668, g692, n4418, g20875, g699,
         g20879, g700, g20891, g698, g20880, g702, g20892, g703, g20901, g701,
         g20893, g705, g20902, g706, g20921, g704, g20903, g708, g20922, g709,
         g20944, g707, g20923, g20945, g712, g20966, g710, g20946, g714,
         g20967, g715, g20989, g713, g20968, g717, g20990, g718, g21009, g716,
         g20991, g720, g21010, g721, g21031, g719, g21011, g723, g21032, g724,
         g21051, g722, g20876, g726, g20881, g20894, g725, g20924, g729,
         g20947, g730, g20969, g728, g20948, g732, g20970, g733, g20992, g731,
         g25260, g735, g25262, g736, g25266, g734, g22218, g738, g22231, g739,
         g22242, g737, n4323, n4312, g22126, g818, g22145, g819, g22162, g817,
         g22146, g821, g22163, g822, g22177, g820, g22029, g830, g22033, g831,
         g22040, g829, g22034, g833, g22041, g834, g22054, g832, g22042, g836,
         g22055, g837, g22066, g835, g22056, g22067, g840, g22087, g838,
         g22068, g842, g22088, g843, g22104, g841, g22089, g845, g22105, g846,
         g22127, g844, g22106, g848, g22128, g849, g22147, g847, g22129, g851,
         g22148, g852, g22164, g850, g25209, g857, g25214, g25221, g856,
         g25215, g860, g25222, g861, g25230, g859, g25223, g863, g25231, g864,
         g25240, g862, g25232, g866, g25241, g867, g25248, g865, g30269, g873,
         g30277, g876, g30285, g879, g30643, g918, g30648, g921, g30654,
         g30676, g882, g30681, g885, g30687, g888, g30649, g927, g30655, g930,
         g30662, g933, g30286, g891, g30293, g894, g30298, g897, g30259, g936,
         g30264, g939, g30270, g942, g30247, g900, g30249, g903, g30251, g906,
         g30265, g30271, g948, g30278, g951, g30638, g909, g30642, g912,
         g30647, g915, g30670, g954, g30677, g957, g30682, g960, g25042, g780,
         g25935, g776, g26530, g771, g27123, g767, g27603, g762, g28146, g758,
         g28635, g753, g29110, g29354, g29580, g740, g868, g869, n4363, n4364,
         g1088, n4381, g996, n4387, g27257, g1041, g27262, g1030, g27270,
         g1033, g27263, g1056, g27271, g1045, g27282, g1048, g27272, g27283,
         g1060, g27297, g1063, g27284, g1085, g27298, g1075, g27313, g1078,
         g28738, g1095, g28746, g1098, g28758, g1101, g29198, g1104, g29204,
         g1107, g29209, g1110, g28747, g1114, g28759, g1115, g28767, g1113,
         g26806, g1116, g26809, g26813, g1122, g26810, g1125, g26814, g1128,
         g26818, g1131, g27761, g1135, g27763, g1136, g27765, g1134, g29609,
         g999, g29612, g1000, g29616, g1001, g30701, g1002, g30703, g1003,
         g30705, g1004, g30470, g1005, g30485, g1006, g30500, g29170, g1009,
         g29173, g1010, g29179, g1008, g26661, g1090, g26665, g1091, g26669,
         g1089, g1137, n8027, DFF_649_n1, g1139, n8026, DFF_651_n1, g1141,
         n8025, DFF_653_n1, g967, n8024, DFF_655_n1, g969, DFF_657_n1, g971,
         n8021, DFF_659_n1, g973, n8020, DFF_661_n1, g975, n8019, DFF_663_n1,
         g977, n8018, n4486, n4283, g986, n4432, g992, n4277, n8017, g1029,
         g1036, g1037, g1038, g1040, g1044, g1051, g1052, g1053, g1054, g1055,
         g1059, g1066, g1067, g1068, g1069, g1070, g1074, g1081, g1083, g1084,
         g1011, g1024, n4371, n4316, g1236, n4300, g21843, g1240, g18707,
         g1243, n4353, g18763, g1196, n4304, g1199, g1209, g1210, g1142, g1255,
         g1145, g1256, g1257, g1148, g1258, g1259, g1152, g1260, g1251, g1155,
         g1252, g1253, g1158, g1254, g1176, n4460, n4459, g1172, n4465, g23081,
         g1173, g23111, g23126, g1175, g23392, g23406, g24179, g24181, g1164,
         g24213, g1165, g24223, g1166, g23110, g1167, g23014, g1171, g23039,
         g1151, g24212, g24222, g24235, g1214, g1221, g13155, g1229, n4549,
         n4361, g13124, g1235, g1186, n4548, g13171, g1244, g1245, g27273,
         g1262, g27285, g1263, g27299, g1261, g27286, g1265, g27300, g1266,
         g27314, g1264, g27301, g1268, g27315, g1269, g27328, g27316, g1271,
         g27329, g1272, g27339, g1270, g24501, g1273, g24510, g1276, g24521,
         g1279, g24511, g1282, g24522, g1285, g24532, g1288, g28351, g1300,
         g28355, g1303, g28360, g1306, g28346, g1291, g28350, g1294, g28354,
         g1297, g26547, g26557, g1180, g26569, g1183, g1192, n4454, g22615,
         n8009, DFF_783_n1, DFF_792_n1, g1211, n8008, n8007, n8006, n8005,
         n8004, n8003, g1222, g1223, g24072, g1224, n4489, n4358, g1315, n4294,
         g16671, g1316, g20333, g1345, n4428, g20717, g1326, n4402, g21969,
         g1319, n4476, g23329, g1339, n4421, g24430, g1332, n4412, g25189,
         g1346, n4401, g26666, g1358, n4411, g26781, g1352, n4469, g27678,
         g1365, n4475, g27718, g1372, n4395, g28321, g1378, n4417, g20882,
         g20896, g1386, g20910, g1384, g20897, g1388, g20911, g1389, g20925,
         g1387, g20912, g1391, g20926, g1392, g20949, g1390, g20927, g1394,
         g20950, g1395, g20972, g1393, g20951, g1397, g20973, g1398, g20993,
         g1396, g20974, g1400, g20994, g21015, g1399, g20995, g1403, g21016,
         g1404, g21033, g1402, g21017, g1406, g21034, g1407, g21052, g1405,
         g21035, g1409, g21053, g1410, g21070, g1408, g20883, g1412, g20898,
         g1413, g20913, g1411, g20952, g1415, g20975, g1416, g20996, g20976,
         g1418, g20997, g1419, g21018, g1417, g25263, g1421, g25267, g1422,
         g25270, g1420, g22234, g1424, g22247, g1425, g22263, g1423, n4317,
         n4515, g1547, n4368, g22149, g1512, g22166, g1513, g22178, g1511,
         g22167, g22179, g1516, g22191, g1514, g22035, g1524, g22043, g1525,
         g22057, g1523, g22044, g1527, g22058, g1528, g22073, g1526, g22059,
         g1530, g22074, g1531, g22090, g1529, g22075, g1533, g22091, g1534,
         g22112, g1532, g22092, g1536, g22113, g22130, g1535, g22114, g1539,
         g22131, g1540, g22150, g1538, g22132, g1542, g22151, g1543, g22168,
         g1541, g22152, g1545, g22169, g1546, g22180, g1544, g25217, g1551,
         g25224, g1552, g25233, g1550, g25225, g1554, g25234, g1555, g25242,
         g25235, g1557, g25243, g1558, g25249, g1556, g25244, g1560, g25250,
         g1561, g25255, g1559, g30279, g1567, g30287, g1570, g30294, g1573,
         g30651, g1612, g30657, g1615, g30663, g1618, g30683, g1576, g30688,
         g1579, g30692, g1582, g30658, g30664, g1624, g30671, g1627, g30295,
         g1585, g30299, g1588, g30302, g1591, g30266, g1630, g30272, g1633,
         g30280, g1636, g30250, g1594, g30252, g1597, g30255, g1600, g30273,
         g1639, g30281, g1642, g30288, g1645, g30644, g1603, g30650, g30656,
         g1609, g30678, g1648, g30684, g1651, g30689, g1654, g25056, g1466,
         g25938, g1462, g26531, g1457, g27129, g1453, g27612, g1448, g28147,
         g1444, g28636, g1439, g29111, g1435, g29355, g29581, g1426, g1562,
         g1563, n4518, g1690, n4386, g27264, g1735, g27274, g1724, g27287,
         g1727, g27275, g1750, g27288, g1739, g27302, g1742, g27289, g1765,
         g27303, g1754, g27317, g1757, g27304, g1779, g27318, g27330, g1772,
         g28749, g1789, g28760, g1792, g28771, g1795, g29205, g1798, g29212,
         g1801, g29218, g1804, g28761, g1808, g28772, g1809, g28778, g1807,
         g26811, g1810, g26815, g1813, g26820, g1816, g26816, g1819, g26821,
         g1822, g26824, g27764, g1829, g27766, g1830, g27768, g1828, g29613,
         g1693, g29617, g1694, g29620, g1695, g30704, g1696, g30706, g1697,
         g30708, g1698, g30487, g1699, g30503, g1700, g30338, g1701, g29178,
         g1703, g29181, g1704, g29184, g1702, g26667, g26670, g1785, g26675,
         g1783, g1831, n7988, DFF_999_n1, g1833, n7987, DFF_1001_n1, g1835,
         n7986, DFF_1003_n1, g1661, n7985, DFF_1005_n1, g1663, n7984,
         DFF_1007_n1, g1665, n7983, DFF_1009_n1, g1667, DFF_1011_n1, g1669,
         n7980, DFF_1013_n1, g1671, n7979, n4484, n4284, g1680, n4488, g1686,
         n4276, n7978, g1723, g1730, g1731, g1732, g1733, g1734, g1738, g1745,
         g1747, g1748, g1749, g1753, g1760, g1761, g1762, g1763, g1764, g1768,
         g1775, g1776, g1777, g1778, g1705, g1718, n4296, n4315, g1930, n4366,
         g21845, g1934, g18743, g1937, g18794, g1890, n4297, g1893, g1903,
         g1904, g1836, g1944, g1949, g1950, g1951, g1842, g1953, g1846, g1954,
         g1945, g1849, g1946, g1947, g1852, g1948, g1870, n4458, n4457, g1866,
         n4464, g23097, g1867, g23124, g1868, g23137, g1869, g23400, g23413,
         g24182, g24208, g1858, g24219, g1859, g24231, g1860, g23123, g1861,
         g23030, g1865, g23058, g1845, g24218, g24230, g24243, g1908, g1915,
         g1922, g13164, g1923, DFF_1099_n1, n7971, DFF_1100_n1, g13135, g1929,
         g1880, n4545, g13182, g1938, g1939, g27290, g1956, g27305, g1957,
         g27319, g1955, g27306, g1959, g27320, g1960, g27331, g1958, g27321,
         g1962, g27332, g1963, g27340, g1961, g27333, g27341, g1966, g27346,
         g1964, g24513, g1967, g24524, g1970, g24534, g1973, g24525, g1976,
         g24535, g1979, g24545, g1982, g28357, g1994, g28362, g1997, g28366,
         g2000, g28352, g1985, g28356, g1988, g28361, g1991, g26559, g26573,
         g1874, g26592, g1877, g1886, n4493, g22651, n7968, DFF_1133_n1,
         DFF_1142_n1, g1905, n7967, n7966, n7965, n7964, n7963, n7962, g1916,
         g1917, g24083, n7960, n4357, g2009, n4293, g16692, g2010, g20353,
         g2039, n4427, g20752, g2020, n4400, g21972, g2013, n4474, g23339,
         g2033, n4420, g24434, g2026, n4410, g25194, g2040, n4399, g26671,
         g2052, n4409, g26789, g2046, n4468, g27682, g2059, n4473, g27722,
         g28325, g2072, n4416, g20899, g2079, g20915, g2080, g20934, g2078,
         g20916, g2082, g20935, g2083, g20953, g2081, g20936, g2085, g20954,
         g2086, g20977, g2084, g20955, g2088, g20978, g2089, g20999, g2087,
         g20979, g2091, g21000, g21019, g2090, g21001, g2094, g21020, g2095,
         g21039, g2093, g21021, g2097, g21040, g2098, g21054, g2096, g21041,
         g2100, g21055, g2101, g21071, g2099, g21056, g2103, g21072, g2104,
         g21080, g2102, g20900, g2106, g20917, g20937, g2105, g20980, g2109,
         g21002, g2110, g21022, g2108, g21003, g2112, g21023, g2113, g21042,
         g2111, g25268, g2115, g25271, g2116, g25279, g2114, g22249, g2118,
         g22267, g2119, g22280, g2117, n4324, g2241, n4367, g22170, g2206,
         g22182, g2207, g22192, g2205, g22183, g2209, g22193, g2210, g22200,
         g2208, g22045, g2218, g22060, g2219, g22076, g2217, g22061, g2221,
         g22077, g2222, g22097, g2220, g22078, g2224, g22098, g22115, g2223,
         g22099, g2227, g22116, g2228, g22138, g2226, g22117, g2230, g22139,
         g2231, g22153, g2229, g22140, g2233, g22154, g2234, g22171, g2232,
         g22155, g2236, g22172, g2237, g22184, g2235, g22173, g2239, g22185,
         g22194, g2238, g25227, g2245, g25236, g2246, g25245, g2244, g25237,
         g2248, g25246, g2249, g25251, g2247, g25247, g2251, g25252, g2252,
         g25256, g2250, g25253, g2254, g25257, g2255, g25259, g2253, g30289,
         g2261, g30296, g30300, g2267, g30660, g2306, g30666, g2309, g30672,
         g2312, g30690, g2270, g30693, g2273, g30695, g2276, g30667, g2315,
         g30673, g2318, g30679, g2321, g30301, g2279, g30303, g2282, g30304,
         g2285, g30274, g2324, g30282, g30290, g2330, g30253, g2288, g30256,
         g2291, g30260, g2294, g30283, g2333, g30291, g2336, g30297, g2339,
         g30652, g2297, g30659, g2300, g30665, g2303, g30686, g2342, g30691,
         g2345, g30694, g2348, g25067, g2160, g25940, g26532, g2151, g27131,
         g2147, g27621, g2142, g28148, g2138, g28637, g2133, g29112, g2129,
         g29357, g29582, g2120, g2256, g2257, n4516, g27276, g2429, g27291,
         g2418, g27307, g2421, g27292, g2444, g27308, g2433, g27322, g2436,
         g27309, g2459, g27323, g2448, g27334, g2451, g27324, g2473, g27335,
         g2463, g27342, g2466, g28763, g2483, g28773, g2486, g28782, g29213,
         g2492, g29221, g2495, g29226, g2498, g28774, g2502, g28783, g2503,
         g28788, g2501, g26817, g2504, g26822, g2507, g26825, g2510, g26823,
         g2513, g26826, g2516, g26827, g2519, g27767, g2523, g27769, g2524,
         g27771, g29618, g2387, g29621, g2388, g29623, g2389, g30707, g2390,
         g30709, g2391, g30566, g2392, g30505, g2393, g30341, g2394, g30356,
         g2395, g29182, g2397, g29185, g2398, g29187, g2396, g26672, g2478,
         g26676, g2479, g26025, g2525, n7946, DFF_1349_n1, g2527, n7945,
         DFF_1351_n1, g2529, n7944, DFF_1353_n1, g2355, n7943, DFF_1355_n1,
         g2357, n7942, DFF_1357_n1, g2359, n7941, DFF_1359_n1, g2361, n7940,
         DFF_1361_n1, n7938, DFF_1363_n1, g2365, n7937, n4483, n4285, g2374,
         n4487, g30055, g2380, n4275, n7936, DFF_1378_n1, g2417, g2424, g2425,
         g2426, g2427, g2428, g2432, g2439, g2441, g2442, g2443, g2447, g2454,
         g2455, g2456, g2457, g2458, g2462, g2469, g2470, g2471, g2472, g2412,
         n4314, n4370, g2624, n4299, g21847, g2628, g18780, g2631, n4352,
         g18820, g2584, n4303, g2587, g2597, g2598, g2530, g2638, g2643, g2533,
         g2645, g2536, g2646, g2647, g2540, g2648, g2639, g2543, g2640, g2641,
         g2546, g2642, g2564, n4456, n4455, g2560, n4463, g23114, g2561,
         g23133, g2562, g21970, g23407, g23418, g24209, g24214, g2552, g24226,
         g2553, g24238, g2554, g23132, g2555, g23047, g2559, g23076, g2539,
         g24225, g24237, g24250, g2602, g2609, g13175, g2617, n7930, g30072,
         n7929, g13143, g2623, g2574, n4543, g13194, g2632, g2633, g27310,
         g2650, g27325, g2651, g27336, g2649, g27326, g2653, g27337, g2654,
         g27343, g2652, g27338, g2656, g27344, g27347, g2655, g27345, g2659,
         g27348, g2660, g27354, g2658, g24527, g2661, g24537, g2664, g24547,
         g2667, g24538, g2670, g24548, g2673, g24557, g2676, g28364, g2688,
         g28368, g2691, g28371, g2694, g28358, g2679, g28363, g28367, g2685,
         g26575, g2565, g26596, g2568, g26616, g2571, g2580, g22687, n7926,
         g30061, g2599, n7925, n7924, n7923, n7922, n7921, n7920, g2611,
         g24092, g2612, n4490, n7918, n4356, g2703, n4292, g16718, g2704,
         g20375, g2733, n4426, g20789, g2714, n4398, g21974, g2707, n4472,
         g23348, g2727, n4419, g24438, g2720, n4408, g25197, g2734, n4397,
         g26677, g2746, n4407, g26795, g27243, g2753, n4471, g27724, g2760,
         n4393, g28328, g2766, n4415, g20918, g2773, g20939, g2774, g20962,
         g2772, g20940, g2776, g20963, g2777, g20981, g2775, g20964, g2779,
         g20982, g2780, g21004, g2778, g20983, g2782, g21005, g2783, g21025,
         g21006, g2785, g21026, g2786, g21043, g2784, g21027, g2788, g21044,
         g2789, g21060, g2787, g21045, g2791, g21061, g2792, g21073, g2790,
         g21062, g2794, g21074, g2795, g21081, g2793, g21075, g2797, g21082,
         g2798, g21094, g20919, g2800, g20941, g2801, g20965, g2799, g21007,
         g2803, g21028, g2804, g21046, g2802, g21029, g2806, g21047, g2807,
         g21063, g2805, g25272, g2809, g25280, g2810, g25288, g2808, g22269,
         g2812, g22284, g2813, g22299, g20877, n7913, g20884, n7912, n4263,
         n4269, g3043, n4268, g3044, n4267, g3045, n4266, g3046, n4265, g3047,
         n4272, g3048, n4271, g3049, n4270, g3050, n4259, g3051, n4236, g3052,
         n4239, g3053, n4237, n4234, g3056, n4233, g3057, n4238, g3058, n4235,
         g3059, n4240, g3060, n4232, g3061, n4245, g3062, n4248, g3063, n4246,
         g3064, n4243, g3065, n4242, g3066, n4247, g3067, n4244, g3068, n4249,
         g3069, n4241, n4254, g3071, n4257, g3072, n4255, g3073, n4252, g3074,
         n4251, g3075, n4256, g3076, n4253, g3077, n4258, g3078, n4250, g2997,
         g25265, g2993, g26048, n7909, g23330, g3006, g24445, g3002, g25191,
         g3013, g26031, g26786, g3024, n4262, g3018, n4481, g23359, g3028,
         n4350, g24446, g3036, n4480, g25202, g3032, n7907, DFF_1612_n1, g2987,
         n4365, g16824, g16844, g16853, g16860, g16803, g16835, g16851, g16857,
         g16866, g3083, n4261, N995, n4577, g16845, g16854, g16861, g16880,
         g18755, g18804, g18837, g18868, g18907, g2990, N690, n4578, n4260,
         n4309, n4308, n4307, n4306, n4524, n4525, n4511, n4509, n4499, n4520,
         n3683, n3887, n3686, n3890, n3692, n3896, n4513, n3897, n3424, n3427,
         n3433, n4529, n4530, n4522, n4523, n4521, n3171, n3159, n3163, n3893,
         n3689, n3430, n4527, n4528, n4526, n3167, n3894, n3888, n3891, n2302,
         n2289, n2303, n2275, n4066, n4065, n4606, n4618, n4640, n2489, n2542,
         n2617, n2279, n2207, n2381, n2309, n2237, n2459, n3936, n3260, n3252,
         n3254, n3293, n3334, n4102, n3374, n3038, n3070, n3102, n3130, n2800,
         n2798, n2616, n2594, n3940, n3705, n3933, n3939, n3700, n4058, n4123,
         n4101, n3938, n4182, n4073, n4057, n4122_Tj_Payload, n4122,
         n4160_Tj_Payload, n4149_Tj_Payload, n4149, n4161_Tj_Payload, Tj_OUT1,
         Tj_OUT2, Tj_OUT3, Tj_OUT4, Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7,
         Tj_OUT8, Tj_OUT5678, Tj_Trigger, n18, n29, n41, n97, n300, n323, n326,
         n330, n336, n339, n342, n375, n467, n470, n532, n534, n549, n578,
         n580, n608, n610, n631, n632, n633, n634, n680, n791, n879, n882,
         n885, n888, n962, n984, n1027, n1136, n1230, n1233, n1305, n1330,
         n1480, n1574, n1577, n1636, n1647, n1669, n1808, n9338, n9339, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9615, n9616,
         n9672, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9894, n9895, n9896, n9897, n9898,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10120,
         n10121, n10122, n10123, n10124, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, U4467_n1, U4904_n1, U4930_n1, U5128_n1, U5141_n1, U5749_n1,
         U5750_n1, U5751_n1, U5752_n1, U5753_n1, U5754_n1, U5755_n1, U5756_n1,
         U5757_n1, U5758_n1, U5759_n1, U5760_n1, U5761_n1, U5762_n1, U5763_n1,
         U5764_n1, U5882_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1, U6140_n1,
         U6460_n1, U6470_n1, U6562_n1, U6563_n1, U6718_n1, U7116_n1, U7118_n1,
         U7293_n1;
  assign g8251 = test_so3;
  assign g7519 = test_so4;
  assign g4450 = test_so5;
  assign g7909 = test_so23;
  assign g5612 = test_so57;
  assign g5695 = test_so63;
  assign g7084 = test_so73;
  assign g8270 = test_so99;
  assign g8258 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(g51), .SI(test_si1), .SE(n10227), .CLK(n10414), .Q(
        n8104), .QN(n18258) );
  SDFFX1 DFF_1_Q_reg ( .D(g16802), .SI(n8104), .SE(n10227), .CLK(n10414), .Q(
        n8103) );
  SDFFX1 DFF_2_Q_reg ( .D(g16823), .SI(n8103), .SE(n10227), .CLK(n10414), .Q(
        n8102), .QN(DFF_2_n1) );
  SDFFX1 DFF_3_Q_reg ( .D(n4264), .SI(n8102), .SE(n10227), .CLK(n10414), .Q(
        g2950), .QN(n4423) );
  SDFFX1 DFF_4_Q_reg ( .D(n18), .SI(g2950), .SE(n10228), .CLK(n10415), .Q(
        g2883), .QN(n4330) );
  SDFFX1 DFF_5_Q_reg ( .D(g22026), .SI(g2883), .SE(n10228), .CLK(n10415), .Q(
        g2888), .QN(n10152) );
  SDFFX1 DFF_6_Q_reg ( .D(g23358), .SI(g2888), .SE(n10233), .CLK(n10420), .Q(
        g2896), .QN(n4431) );
  SDFFX1 DFF_7_Q_reg ( .D(g24473), .SI(g2896), .SE(n10233), .CLK(n10420), .Q(
        g2892), .QN(n10173) );
  SDFFX1 DFF_8_Q_reg ( .D(g25201), .SI(g2892), .SE(n10233), .CLK(n10420), .Q(
        g2903), .QN(n4305) );
  SDFFX1 DFF_9_Q_reg ( .D(g26037), .SI(g2903), .SE(n10233), .CLK(n10420), .Q(
        g2900), .QN(n4291) );
  SDFFX1 DFF_10_Q_reg ( .D(g26798), .SI(g2900), .SE(n10233), .CLK(n10420), .Q(
        g2908), .QN(n4355) );
  SDFFX1 DFF_11_Q_reg ( .D(n4273), .SI(g2908), .SE(n10228), .CLK(n10415), .Q(
        g2912), .QN(n4482) );
  SDFFX1 DFF_12_Q_reg ( .D(g23357), .SI(g2912), .SE(n10228), .CLK(n10415), .Q(
        g2917), .QN(n4479) );
  SDFFX1 DFF_13_Q_reg ( .D(g24476), .SI(g2917), .SE(n10228), .CLK(n10415), .Q(
        g2924), .QN(n4349) );
  SDFFX1 DFF_14_Q_reg ( .D(g25199), .SI(g2924), .SE(n10228), .CLK(n10415), .Q(
        g2920), .QN(n9892) );
  SDFFX1 DFF_15_Q_reg ( .D(n4280), .SI(g2920), .SE(n10228), .CLK(n10415), .Q(
        test_so1) );
  SDFFX1 DFF_16_Q_reg ( .D(n4281), .SI(test_si2), .SE(n10225), .CLK(n10412), 
        .Q(n8099) );
  SDFFX1 DFF_17_Q_reg ( .D(g51), .SI(n8099), .SE(n10225), .CLK(n10412), .Q(
        g8021) );
  SDFFX1 DFF_18_Q_reg ( .D(g8021), .SI(g8021), .SE(n10225), .CLK(n10412), .Q(
        n8098), .QN(DFF_18_n1) );
  SDFFX1 DFF_19_Q_reg ( .D(n4279), .SI(n8098), .SE(n10225), .CLK(n10412), .Q(
        g2879), .QN(n4351) );
  SDFFX1 DFF_20_Q_reg ( .D(g3212), .SI(g2879), .SE(n10225), .CLK(n10412), .Q(
        g2934), .QN(n10148) );
  SDFFX1 DFF_21_Q_reg ( .D(g3228), .SI(g2934), .SE(n10225), .CLK(n10412), .Q(
        g2935), .QN(n10131) );
  SDFFX1 DFF_22_Q_reg ( .D(g3227), .SI(g2935), .SE(n10226), .CLK(n10413), .Q(
        g2938), .QN(n10132) );
  SDFFX1 DFF_23_Q_reg ( .D(g3226), .SI(g2938), .SE(n10226), .CLK(n10413), .Q(
        g2941), .QN(n10129) );
  SDFFX1 DFF_24_Q_reg ( .D(g3225), .SI(g2941), .SE(n10226), .CLK(n10413), .Q(
        g2944), .QN(n10135) );
  SDFFX1 DFF_25_Q_reg ( .D(g3224), .SI(g2944), .SE(n10226), .CLK(n10413), .Q(
        g2947), .QN(n10133) );
  SDFFX1 DFF_26_Q_reg ( .D(g3223), .SI(g2947), .SE(n10226), .CLK(n10413), .Q(
        g2953), .QN(n10134) );
  SDFFX1 DFF_27_Q_reg ( .D(g3222), .SI(g2953), .SE(n10226), .CLK(n10413), .Q(
        g2956), .QN(n10136) );
  SDFFX1 DFF_28_Q_reg ( .D(g3221), .SI(g2956), .SE(n10226), .CLK(n10413), .Q(
        g2959), .QN(n10130) );
  SDFFX1 DFF_29_Q_reg ( .D(g3232), .SI(g2959), .SE(n10226), .CLK(n10413), .Q(
        g2962), .QN(n10150) );
  SDFFX1 DFF_30_Q_reg ( .D(g3220), .SI(g2962), .SE(n10226), .CLK(n10413), .Q(
        g2963), .QN(n10139) );
  SDFFX1 DFF_31_Q_reg ( .D(g3219), .SI(g2963), .SE(n10226), .CLK(n10413), .Q(
        test_so2), .QN(n10198) );
  SDFFX1 DFF_32_Q_reg ( .D(g3218), .SI(test_si3), .SE(n10225), .CLK(n10412), 
        .Q(g2969), .QN(n10142) );
  SDFFX1 DFF_33_Q_reg ( .D(g3217), .SI(g2969), .SE(n10225), .CLK(n10412), .Q(
        g2972), .QN(n10140) );
  SDFFX1 DFF_34_Q_reg ( .D(g3216), .SI(g2972), .SE(n10225), .CLK(n10412), .Q(
        g2975), .QN(n10141) );
  SDFFX1 DFF_35_Q_reg ( .D(g3215), .SI(g2975), .SE(n10225), .CLK(n10412), .Q(
        g2978), .QN(n10137) );
  SDFFX1 DFF_36_Q_reg ( .D(g3214), .SI(g2978), .SE(n10225), .CLK(n10412), .Q(
        g2981), .QN(n10143) );
  SDFFX1 DFF_37_Q_reg ( .D(g3213), .SI(g2981), .SE(n10225), .CLK(n10412), .Q(
        g2874), .QN(n10138) );
  SDFFX1 DFF_38_Q_reg ( .D(g18754), .SI(g2874), .SE(n10226), .CLK(n10413), .Q(
        g1506), .QN(n4288) );
  SDFFX1 DFF_39_Q_reg ( .D(g18781), .SI(g1506), .SE(n10226), .CLK(n10413), .Q(
        g1501), .QN(n4565) );
  SDFFX1 DFF_40_Q_reg ( .D(g18803), .SI(g1501), .SE(n10227), .CLK(n10414), .Q(
        g1496), .QN(n4557) );
  SDFFX1 DFF_41_Q_reg ( .D(g18821), .SI(g1496), .SE(n10227), .CLK(n10414), .Q(
        g1491), .QN(n4326) );
  SDFFX1 DFF_42_Q_reg ( .D(g18835), .SI(g1491), .SE(n10227), .CLK(n10414), .Q(
        g1486), .QN(n4390) );
  SDFFX1 DFF_43_Q_reg ( .D(g18852), .SI(g1486), .SE(n10227), .CLK(n10414), .Q(
        g1481), .QN(n4320) );
  SDFFX1 DFF_44_Q_reg ( .D(g18866), .SI(g1481), .SE(n10227), .CLK(n10414), .Q(
        g1476), .QN(n4374) );
  SDFFX1 DFF_45_Q_reg ( .D(g18883), .SI(g1476), .SE(n10227), .CLK(n10414), .Q(
        g1471), .QN(n4378) );
  SDFFX1 DFF_46_Q_reg ( .D(g21880), .SI(g1471), .SE(n10238), .CLK(n10425), .Q(
        g2877) );
  SDFFX1 DFF_47_Q_reg ( .D(g19154), .SI(g2877), .SE(n10238), .CLK(n10425), .Q(
        test_so3) );
  SDFFX1 DFF_48_Q_reg ( .D(test_so3), .SI(test_si4), .SE(n10238), .CLK(n10425), 
        .Q(g813), .QN(n4289) );
  SDFFX1 DFF_49_Q_reg ( .D(g19163), .SI(g813), .SE(n10238), .CLK(n10425), .Q(
        g4090) );
  SDFFX1 DFF_50_Q_reg ( .D(g4090), .SI(g4090), .SE(n10238), .CLK(n10425), .Q(
        g809), .QN(n4567) );
  SDFFX1 DFF_51_Q_reg ( .D(g19173), .SI(g809), .SE(n10238), .CLK(n10425), .Q(
        g4323) );
  SDFFX1 DFF_52_Q_reg ( .D(g4323), .SI(g4323), .SE(n10239), .CLK(n10426), .Q(
        g805), .QN(n4559) );
  SDFFX1 DFF_53_Q_reg ( .D(g19184), .SI(g805), .SE(n10239), .CLK(n10426), .Q(
        g4590) );
  SDFFX1 DFF_54_Q_reg ( .D(g4590), .SI(g4590), .SE(n10239), .CLK(n10426), .Q(
        g801), .QN(n4327) );
  SDFFX1 DFF_55_Q_reg ( .D(g20310), .SI(g801), .SE(n10239), .CLK(n10426), .Q(
        g6225) );
  SDFFX1 DFF_56_Q_reg ( .D(g6225), .SI(g6225), .SE(n10239), .CLK(n10426), .Q(
        g797), .QN(n4391) );
  SDFFX1 DFF_57_Q_reg ( .D(g20343), .SI(g797), .SE(n10239), .CLK(n10426), .Q(
        g6442) );
  SDFFX1 DFF_58_Q_reg ( .D(g6442), .SI(g6442), .SE(n10239), .CLK(n10426), .Q(
        g793), .QN(n4321) );
  SDFFX1 DFF_59_Q_reg ( .D(g20376), .SI(g793), .SE(n10239), .CLK(n10426), .Q(
        g6895) );
  SDFFX1 DFF_60_Q_reg ( .D(g6895), .SI(g6895), .SE(n10239), .CLK(n10426), .Q(
        g789), .QN(n4375) );
  SDFFX1 DFF_61_Q_reg ( .D(g20417), .SI(g789), .SE(n10239), .CLK(n10426), .Q(
        g7334) );
  SDFFX1 DFF_62_Q_reg ( .D(g7334), .SI(g7334), .SE(n10239), .CLK(n10426), .Q(
        g785), .QN(n4379) );
  SDFFX1 DFF_63_Q_reg ( .D(g21878), .SI(g785), .SE(n10240), .CLK(n10427), .Q(
        test_so4) );
  SDFFX1 DFF_64_Q_reg ( .D(test_so4), .SI(test_si5), .SE(n10240), .CLK(n10427), 
        .Q(g2873) );
  SDFFX1 DFF_65_Q_reg ( .D(g19153), .SI(g2873), .SE(n10240), .CLK(n10427), .Q(
        g8249) );
  SDFFX1 DFF_66_Q_reg ( .D(g8249), .SI(g8249), .SE(n10240), .CLK(n10427), .Q(
        g125), .QN(n4290) );
  SDFFX1 DFF_67_Q_reg ( .D(g19162), .SI(g125), .SE(n10240), .CLK(n10427), .Q(
        g4088) );
  SDFFX1 DFF_68_Q_reg ( .D(g4088), .SI(g4088), .SE(n10241), .CLK(n10428), .Q(
        g121), .QN(n4569) );
  SDFFX1 DFF_69_Q_reg ( .D(g19172), .SI(g121), .SE(n10241), .CLK(n10428), .Q(
        g4321) );
  SDFFX1 DFF_70_Q_reg ( .D(g4321), .SI(g4321), .SE(n10241), .CLK(n10428), .Q(
        g117), .QN(n4561) );
  SDFFX1 DFF_71_Q_reg ( .D(g19144), .SI(g117), .SE(n10241), .CLK(n10428), .Q(
        g8023) );
  SDFFX1 DFF_72_Q_reg ( .D(g8023), .SI(g8023), .SE(n10241), .CLK(n10428), .Q(
        g113), .QN(n4328) );
  SDFFX1 DFF_73_Q_reg ( .D(g19149), .SI(g113), .SE(n10241), .CLK(n10428), .Q(
        g8175) );
  SDFFX1 DFF_74_Q_reg ( .D(g8175), .SI(g8175), .SE(n10241), .CLK(n10428), .Q(
        g109), .QN(n4392) );
  SDFFX1 DFF_75_Q_reg ( .D(g19157), .SI(g109), .SE(n10241), .CLK(n10428), .Q(
        g3993) );
  SDFFX1 DFF_76_Q_reg ( .D(g3993), .SI(g3993), .SE(n10241), .CLK(n10428), .Q(
        g105), .QN(n4322) );
  SDFFX1 DFF_77_Q_reg ( .D(g19167), .SI(g105), .SE(n10241), .CLK(n10428), .Q(
        g4200) );
  SDFFX1 DFF_78_Q_reg ( .D(g4200), .SI(g4200), .SE(n10241), .CLK(n10428), .Q(
        g101), .QN(n4376) );
  SDFFX1 DFF_79_Q_reg ( .D(g19178), .SI(g101), .SE(n10241), .CLK(n10428), .Q(
        test_so5) );
  SDFFX1 DFF_80_Q_reg ( .D(test_so5), .SI(test_si6), .SE(n10242), .CLK(n10429), 
        .Q(g97), .QN(n4380) );
  SDFFX1 DFF_81_Q_reg ( .D(g20874), .SI(g97), .SE(n10242), .CLK(n10429), .Q(
        g8096) );
  SDFFX1 DFF_82_Q_reg ( .D(g8096), .SI(g8096), .SE(n10242), .CLK(n10429), .Q(
        g2857) );
  SDFFX1 DFF_83_Q_reg ( .D(g18885), .SI(g2857), .SE(n10242), .CLK(n10429), .Q(
        g2200), .QN(n4287) );
  SDFFX1 DFF_84_Q_reg ( .D(g18975), .SI(g2200), .SE(n10242), .CLK(n10429), .Q(
        g2195), .QN(n4563) );
  SDFFX1 DFF_85_Q_reg ( .D(g18968), .SI(g2195), .SE(n10242), .CLK(n10429), .Q(
        g2190), .QN(n4555) );
  SDFFX1 DFF_86_Q_reg ( .D(g18942), .SI(g2190), .SE(n10242), .CLK(n10429), .Q(
        g2185), .QN(n4325) );
  SDFFX1 DFF_87_Q_reg ( .D(g18906), .SI(g2185), .SE(n10242), .CLK(n10429), .Q(
        g2180), .QN(n4389) );
  SDFFX1 DFF_88_Q_reg ( .D(g18867), .SI(g2180), .SE(n10242), .CLK(n10429), .Q(
        g2175), .QN(n4319) );
  SDFFX1 DFF_89_Q_reg ( .D(g18836), .SI(g2175), .SE(n10242), .CLK(n10429), .Q(
        g2170), .QN(n4373) );
  SDFFX1 DFF_90_Q_reg ( .D(g18957), .SI(g2170), .SE(n10242), .CLK(n10429), .Q(
        g2165), .QN(n4377) );
  SDFFX1 DFF_91_Q_reg ( .D(g21882), .SI(g2165), .SE(n10345), .CLK(n10532), .Q(
        g2878) );
  SDFFX1 DFF_92_Q_reg ( .D(n4598), .SI(g2878), .SE(n10350), .CLK(n10537), .Q(
        g8106), .QN(n4382) );
  SDFFX1 DFF_93_Q_reg ( .D(g8106), .SI(g8106), .SE(n10350), .CLK(n10537), .Q(
        g8030), .QN(n4383) );
  SDFFX1 DFF_94_Q_reg ( .D(g8030), .SI(g8030), .SE(n10350), .CLK(n10537), .Q(
        g3109), .QN(n4494) );
  SDFFX1 DFF_95_Q_reg ( .D(g18669), .SI(g3109), .SE(n10351), .CLK(n10538), .Q(
        test_so6) );
  SDFFX1 DFF_96_Q_reg ( .D(g18719), .SI(test_si7), .SE(n10350), .CLK(n10537), 
        .Q(g3211) );
  SDFFX1 DFF_97_Q_reg ( .D(g18782), .SI(g3211), .SE(n10350), .CLK(n10537), .Q(
        g3084) );
  SDFFX1 DFF_98_Q_reg ( .D(g17222), .SI(g3084), .SE(n10350), .CLK(n10537), .Q(
        g3085) );
  SDFFX1 DFF_99_Q_reg ( .D(g17225), .SI(g3085), .SE(n10350), .CLK(n10537), .Q(
        g3086) );
  SDFFX1 DFF_100_Q_reg ( .D(g17234), .SI(g3086), .SE(n10350), .CLK(n10537), 
        .Q(g3087) );
  SDFFX1 DFF_101_Q_reg ( .D(g17224), .SI(g3087), .SE(n10350), .CLK(n10537), 
        .Q(g3091) );
  SDFFX1 DFF_102_Q_reg ( .D(g17228), .SI(g3091), .SE(n10350), .CLK(n10537), 
        .Q(g3092) );
  SDFFX1 DFF_103_Q_reg ( .D(g17246), .SI(g3092), .SE(n10351), .CLK(n10538), 
        .Q(g3093) );
  SDFFX1 DFF_104_Q_reg ( .D(g17226), .SI(g3093), .SE(n10351), .CLK(n10538), 
        .Q(g3094) );
  SDFFX1 DFF_105_Q_reg ( .D(g17235), .SI(g3094), .SE(n10351), .CLK(n10538), 
        .Q(g3095) );
  SDFFX1 DFF_106_Q_reg ( .D(g17269), .SI(g3095), .SE(n10351), .CLK(n10538), 
        .Q(g3096) );
  SDFFX1 DFF_107_Q_reg ( .D(g25450), .SI(g3096), .SE(n10351), .CLK(n10538), 
        .Q(g3097) );
  SDFFX1 DFF_108_Q_reg ( .D(g25451), .SI(g3097), .SE(n10351), .CLK(n10538), 
        .Q(g3098) );
  SDFFX1 DFF_109_Q_reg ( .D(g25452), .SI(g3098), .SE(n10351), .CLK(n10538), 
        .Q(g3099) );
  SDFFX1 DFF_110_Q_reg ( .D(g28420), .SI(g3099), .SE(n10352), .CLK(n10539), 
        .Q(g3100) );
  SDFFX1 DFF_111_Q_reg ( .D(g28421), .SI(g3100), .SE(n10352), .CLK(n10539), 
        .Q(test_so7) );
  SDFFX1 DFF_112_Q_reg ( .D(g28425), .SI(test_si8), .SE(n10350), .CLK(n10537), 
        .Q(g3102) );
  SDFFX1 DFF_113_Q_reg ( .D(g29936), .SI(g3102), .SE(n10352), .CLK(n10539), 
        .Q(g3103) );
  SDFFX1 DFF_114_Q_reg ( .D(g29939), .SI(g3103), .SE(n10352), .CLK(n10539), 
        .Q(g3104) );
  SDFFX1 DFF_115_Q_reg ( .D(g29941), .SI(g3104), .SE(n10352), .CLK(n10539), 
        .Q(g3105) );
  SDFFX1 DFF_116_Q_reg ( .D(g30796), .SI(g3105), .SE(n10352), .CLK(n10539), 
        .Q(g3106) );
  SDFFX1 DFF_117_Q_reg ( .D(g30798), .SI(g3106), .SE(n10352), .CLK(n10539), 
        .Q(g3107) );
  SDFFX1 DFF_118_Q_reg ( .D(g30801), .SI(g3107), .SE(n10352), .CLK(n10539), 
        .Q(g3108) );
  SDFFX1 DFF_119_Q_reg ( .D(g17229), .SI(g3108), .SE(n10352), .CLK(n10539), 
        .Q(g3155) );
  SDFFX1 DFF_120_Q_reg ( .D(g17247), .SI(g3155), .SE(n10352), .CLK(n10539), 
        .Q(g3158) );
  SDFFX1 DFF_121_Q_reg ( .D(g17302), .SI(g3158), .SE(n10352), .CLK(n10539), 
        .Q(g3161) );
  SDFFX1 DFF_122_Q_reg ( .D(g17236), .SI(g3161), .SE(n10352), .CLK(n10539), 
        .Q(g3164) );
  SDFFX1 DFF_123_Q_reg ( .D(g17270), .SI(g3164), .SE(n10353), .CLK(n10540), 
        .Q(g3167) );
  SDFFX1 DFF_124_Q_reg ( .D(g17340), .SI(g3167), .SE(n10353), .CLK(n10540), 
        .Q(g3170) );
  SDFFX1 DFF_125_Q_reg ( .D(g17248), .SI(g3170), .SE(n10353), .CLK(n10540), 
        .Q(g3173) );
  SDFFX1 DFF_126_Q_reg ( .D(g17303), .SI(g3173), .SE(n10353), .CLK(n10540), 
        .Q(g3176) );
  SDFFX1 DFF_127_Q_reg ( .D(g17383), .SI(g3176), .SE(n10353), .CLK(n10540), 
        .Q(test_so8) );
  SDFFX1 DFF_128_Q_reg ( .D(g17271), .SI(test_si9), .SE(n10351), .CLK(n10538), 
        .Q(g3182) );
  SDFFX1 DFF_129_Q_reg ( .D(g17341), .SI(g3182), .SE(n10351), .CLK(n10538), 
        .Q(g3185) );
  SDFFX1 DFF_130_Q_reg ( .D(g17429), .SI(g3185), .SE(n10351), .CLK(n10538), 
        .Q(g3088) );
  SDFFX1 DFF_131_Q_reg ( .D(g24734), .SI(g3088), .SE(n10351), .CLK(n10538), 
        .Q(n8090) );
  SDFFX1 DFF_132_Q_reg ( .D(g25442), .SI(n8090), .SE(n10236), .CLK(n10423), 
        .Q(n8089) );
  SDFFX1 DFF_133_Q_reg ( .D(g25435), .SI(n8089), .SE(n10236), .CLK(n10423), 
        .Q(g3197) );
  SDFFX1 DFF_134_Q_reg ( .D(g25420), .SI(g3197), .SE(n10236), .CLK(n10423), 
        .Q(n8088) );
  SDFFX1 DFF_135_Q_reg ( .D(g26149), .SI(n8088), .SE(n10235), .CLK(n10422), 
        .Q(g3201), .QN(n4406) );
  SDFFX1 DFF_136_Q_reg ( .D(g26135), .SI(g3201), .SE(n10235), .CLK(n10422), 
        .Q(g3204) );
  SDFFX1 DFF_137_Q_reg ( .D(g26104), .SI(g3204), .SE(n10236), .CLK(n10423), 
        .Q(g3207), .QN(n4329) );
  SDFFX1 DFF_138_Q_reg ( .D(g27380), .SI(g3207), .SE(n10235), .CLK(n10422), 
        .Q(g3188), .QN(n4405) );
  SDFFX1 DFF_139_Q_reg ( .D(n97), .SI(g3188), .SE(n10235), .CLK(n10422), .Q(
        g3133), .QN(n9615) );
  SDFFX1 DFF_140_Q_reg ( .D(g26104), .SI(g3133), .SE(n10236), .CLK(n10423), 
        .Q(n8087) );
  SDFFX1 DFF_141_Q_reg ( .D(n300), .SI(n8087), .SE(n10236), .CLK(n10423), .Q(
        g3128), .QN(n9801) );
  SDFFX1 DFF_142_Q_reg ( .D(g26149), .SI(g3128), .SE(n10236), .CLK(n10423), 
        .Q(n8086) );
  SDFFX1 DFF_143_Q_reg ( .D(g25420), .SI(n8086), .SE(n10237), .CLK(n10424), 
        .Q(test_so9) );
  SDFFX1 DFF_144_Q_reg ( .D(n326), .SI(test_si10), .SE(n10236), .CLK(n10423), 
        .Q(n8084), .QN(DFF_144_n1) );
  SDFFX1 DFF_145_Q_reg ( .D(g25442), .SI(n8084), .SE(n10236), .CLK(n10423), 
        .Q(g3124) );
  SDFFX1 DFF_146_Q_reg ( .D(n330), .SI(g3124), .SE(n10236), .CLK(n10423), .Q(
        n8083), .QN(DFF_146_n1) );
  SDFFX1 DFF_147_Q_reg ( .D(g26104), .SI(n8083), .SE(n10236), .CLK(n10423), 
        .Q(n8082) );
  SDFFX1 DFF_148_Q_reg ( .D(g26135), .SI(n8082), .SE(n10236), .CLK(n10423), 
        .Q(n8081) );
  SDFFX1 DFF_149_Q_reg ( .D(g26149), .SI(n8081), .SE(n10237), .CLK(n10424), 
        .Q(n8080) );
  SDFFX1 DFF_150_Q_reg ( .D(g25420), .SI(n8080), .SE(n10237), .CLK(n10424), 
        .Q(g3112) );
  SDFFX1 DFF_151_Q_reg ( .D(g25435), .SI(g3112), .SE(n10237), .CLK(n10424), 
        .Q(g3110) );
  SDFFX1 DFF_152_Q_reg ( .D(g25442), .SI(g3110), .SE(n10237), .CLK(n10424), 
        .Q(g3111) );
  SDFFX1 DFF_153_Q_reg ( .D(g27380), .SI(g3111), .SE(n10237), .CLK(n10424), 
        .Q(n8079) );
  SDFFX1 DFF_154_Q_reg ( .D(g26104), .SI(n8079), .SE(n10237), .CLK(n10424), 
        .Q(n8078) );
  SDFFX1 DFF_155_Q_reg ( .D(g26135), .SI(n8078), .SE(n10237), .CLK(n10424), 
        .Q(n8077) );
  SDFFX1 DFF_156_Q_reg ( .D(g26149), .SI(n8077), .SE(n10237), .CLK(n10424), 
        .Q(n8076) );
  SDFFX1 DFF_157_Q_reg ( .D(g27380), .SI(n8076), .SE(n10237), .CLK(n10424), 
        .Q(g3151), .QN(n4424) );
  SDFFX1 DFF_158_Q_reg ( .D(g26104), .SI(g3151), .SE(n10237), .CLK(n10424), 
        .Q(g3142), .QN(n4301) );
  SDFFX1 DFF_159_Q_reg ( .D(g26135), .SI(g3142), .SE(n10237), .CLK(n10424), 
        .Q(test_so10), .QN(n10202) );
  SDFFX1 DFF_160_Q_reg ( .D(n97), .SI(test_si11), .SE(n10235), .CLK(n10422), 
        .Q(g185), .QN(n4384) );
  SDFFX1 DFF_161_Q_reg ( .D(g2950), .SI(g185), .SE(n10235), .CLK(n10422), .Q(
        g6231), .QN(n4318) );
  SDFFX1 DFF_162_Q_reg ( .D(g6231), .SI(g6231), .SE(n10235), .CLK(n10422), .Q(
        g6313), .QN(n4512) );
  SDFFX1 DFF_163_Q_reg ( .D(g6313), .SI(g6313), .SE(n10235), .CLK(n10422), .Q(
        g165), .QN(n4369) );
  SDFFX1 DFF_164_Q_reg ( .D(g22100), .SI(g165), .SE(n10264), .CLK(n10451), .Q(
        g130), .QN(n10112) );
  SDFFX1 DFF_165_Q_reg ( .D(g22122), .SI(g130), .SE(n10264), .CLK(n10451), .Q(
        g131), .QN(n10111) );
  SDFFX1 DFF_166_Q_reg ( .D(g22141), .SI(g131), .SE(n10264), .CLK(n10451), .Q(
        g129), .QN(n9738) );
  SDFFX1 DFF_167_Q_reg ( .D(g22123), .SI(g129), .SE(n10264), .CLK(n10451), .Q(
        g133), .QN(n10110) );
  SDFFX1 DFF_168_Q_reg ( .D(g22142), .SI(g133), .SE(n10264), .CLK(n10451), .Q(
        g134), .QN(n10109) );
  SDFFX1 DFF_169_Q_reg ( .D(g22161), .SI(g134), .SE(n10264), .CLK(n10451), .Q(
        g132), .QN(n9737) );
  SDFFX1 DFF_170_Q_reg ( .D(g22025), .SI(g132), .SE(n10264), .CLK(n10451), .Q(
        g142), .QN(n10108) );
  SDFFX1 DFF_171_Q_reg ( .D(g22027), .SI(g142), .SE(n10264), .CLK(n10451), .Q(
        g143), .QN(n10107) );
  SDFFX1 DFF_172_Q_reg ( .D(g22030), .SI(g143), .SE(n10264), .CLK(n10451), .Q(
        g141), .QN(n9736) );
  SDFFX1 DFF_173_Q_reg ( .D(g22028), .SI(g141), .SE(n10264), .CLK(n10451), .Q(
        g145), .QN(n10106) );
  SDFFX1 DFF_174_Q_reg ( .D(g22031), .SI(g145), .SE(n10265), .CLK(n10452), .Q(
        g146), .QN(n10105) );
  SDFFX1 DFF_175_Q_reg ( .D(g22037), .SI(g146), .SE(n10265), .CLK(n10452), .Q(
        test_so11), .QN(n10214) );
  SDFFX1 DFF_176_Q_reg ( .D(g22032), .SI(test_si12), .SE(n10263), .CLK(n10450), 
        .Q(g148), .QN(n10104) );
  SDFFX1 DFF_177_Q_reg ( .D(g22038), .SI(g148), .SE(n10263), .CLK(n10450), .Q(
        g149), .QN(n10103) );
  SDFFX1 DFF_178_Q_reg ( .D(g22047), .SI(g149), .SE(n10263), .CLK(n10450), .Q(
        g147), .QN(n9735) );
  SDFFX1 DFF_179_Q_reg ( .D(g22039), .SI(g147), .SE(n10263), .CLK(n10450), .Q(
        g151), .QN(n10102) );
  SDFFX1 DFF_180_Q_reg ( .D(g22048), .SI(g151), .SE(n10263), .CLK(n10450), .Q(
        g152), .QN(n10101) );
  SDFFX1 DFF_181_Q_reg ( .D(g22063), .SI(g152), .SE(n10263), .CLK(n10450), .Q(
        g150), .QN(n9734) );
  SDFFX1 DFF_182_Q_reg ( .D(g22049), .SI(g150), .SE(n10263), .CLK(n10450), .Q(
        g154), .QN(n10100) );
  SDFFX1 DFF_183_Q_reg ( .D(g22064), .SI(g154), .SE(n10263), .CLK(n10450), .Q(
        g155), .QN(n10099) );
  SDFFX1 DFF_184_Q_reg ( .D(g22079), .SI(g155), .SE(n10263), .CLK(n10450), .Q(
        g153), .QN(n9733) );
  SDFFX1 DFF_185_Q_reg ( .D(g22065), .SI(g153), .SE(n10259), .CLK(n10446), .Q(
        g157), .QN(n10098) );
  SDFFX1 DFF_186_Q_reg ( .D(g22080), .SI(g157), .SE(n10261), .CLK(n10448), .Q(
        g158), .QN(n10097) );
  SDFFX1 DFF_187_Q_reg ( .D(g22101), .SI(g158), .SE(n10261), .CLK(n10448), .Q(
        g156), .QN(n9732) );
  SDFFX1 DFF_188_Q_reg ( .D(g22081), .SI(g156), .SE(n10263), .CLK(n10450), .Q(
        g160), .QN(n9694) );
  SDFFX1 DFF_189_Q_reg ( .D(g22102), .SI(g160), .SE(n10263), .CLK(n10450), .Q(
        g161), .QN(n9693) );
  SDFFX1 DFF_190_Q_reg ( .D(g22124), .SI(g161), .SE(n10264), .CLK(n10451), .Q(
        g159), .QN(n9692) );
  SDFFX1 DFF_191_Q_reg ( .D(g22103), .SI(g159), .SE(n10264), .CLK(n10451), .Q(
        test_so12), .QN(n10213) );
  SDFFX1 DFF_192_Q_reg ( .D(g22125), .SI(test_si13), .SE(n10261), .CLK(n10448), 
        .Q(g164), .QN(n9731) );
  SDFFX1 DFF_193_Q_reg ( .D(g22143), .SI(g164), .SE(n10262), .CLK(n10449), .Q(
        g162), .QN(n9730) );
  SDFFX1 DFF_194_Q_reg ( .D(g25204), .SI(g162), .SE(n10262), .CLK(n10449), .Q(
        g169), .QN(n9800) );
  SDFFX1 DFF_195_Q_reg ( .D(g25206), .SI(g169), .SE(n10262), .CLK(n10449), .Q(
        g170), .QN(n9799) );
  SDFFX1 DFF_196_Q_reg ( .D(g25211), .SI(g170), .SE(n10262), .CLK(n10449), .Q(
        g168), .QN(n9798) );
  SDFFX1 DFF_197_Q_reg ( .D(g25207), .SI(g168), .SE(n10262), .CLK(n10449), .Q(
        g172), .QN(n9797) );
  SDFFX1 DFF_198_Q_reg ( .D(g25212), .SI(g172), .SE(n10262), .CLK(n10449), .Q(
        g173), .QN(n9796) );
  SDFFX1 DFF_199_Q_reg ( .D(g25218), .SI(g173), .SE(n10262), .CLK(n10449), .Q(
        g171), .QN(n9795) );
  SDFFX1 DFF_200_Q_reg ( .D(g25213), .SI(g171), .SE(n10262), .CLK(n10449), .Q(
        g175), .QN(n9794) );
  SDFFX1 DFF_201_Q_reg ( .D(g25219), .SI(g175), .SE(n10262), .CLK(n10449), .Q(
        g176), .QN(n9793) );
  SDFFX1 DFF_202_Q_reg ( .D(g25228), .SI(g176), .SE(n10262), .CLK(n10449), .Q(
        g174), .QN(n9792) );
  SDFFX1 DFF_203_Q_reg ( .D(g25220), .SI(g174), .SE(n10262), .CLK(n10449), .Q(
        g178) );
  SDFFX1 DFF_204_Q_reg ( .D(g25229), .SI(g178), .SE(n10262), .CLK(n10449), .Q(
        g179) );
  SDFFX1 DFF_205_Q_reg ( .D(g25239), .SI(g179), .SE(n10263), .CLK(n10450), .Q(
        g177) );
  SDFFX1 DFF_206_Q_reg ( .D(g30261), .SI(g177), .SE(n10269), .CLK(n10456), .Q(
        g186) );
  SDFFX1 DFF_207_Q_reg ( .D(g30267), .SI(g186), .SE(n10270), .CLK(n10457), .Q(
        test_so13) );
  SDFFX1 DFF_208_Q_reg ( .D(g30275), .SI(test_si14), .SE(n10270), .CLK(n10457), 
        .Q(g192) );
  SDFFX1 DFF_209_Q_reg ( .D(g30637), .SI(g192), .SE(n10270), .CLK(n10457), .Q(
        g231) );
  SDFFX1 DFF_210_Q_reg ( .D(g30640), .SI(g231), .SE(n10270), .CLK(n10457), .Q(
        g234) );
  SDFFX1 DFF_211_Q_reg ( .D(g30645), .SI(g234), .SE(n10270), .CLK(n10457), .Q(
        g237) );
  SDFFX1 DFF_212_Q_reg ( .D(g30668), .SI(g237), .SE(n10270), .CLK(n10457), .Q(
        g195) );
  SDFFX1 DFF_213_Q_reg ( .D(g30674), .SI(g195), .SE(n10270), .CLK(n10457), .Q(
        g198) );
  SDFFX1 DFF_214_Q_reg ( .D(g30680), .SI(g198), .SE(n10266), .CLK(n10453), .Q(
        g201) );
  SDFFX1 DFF_215_Q_reg ( .D(g30641), .SI(g201), .SE(n10266), .CLK(n10453), .Q(
        g240) );
  SDFFX1 DFF_216_Q_reg ( .D(g30646), .SI(g240), .SE(n10266), .CLK(n10453), .Q(
        g243) );
  SDFFX1 DFF_217_Q_reg ( .D(g30653), .SI(g243), .SE(n10265), .CLK(n10452), .Q(
        g246) );
  SDFFX1 DFF_218_Q_reg ( .D(g30276), .SI(g246), .SE(n10265), .CLK(n10452), .Q(
        g204) );
  SDFFX1 DFF_219_Q_reg ( .D(g30284), .SI(g204), .SE(n10265), .CLK(n10452), .Q(
        g207) );
  SDFFX1 DFF_220_Q_reg ( .D(g30292), .SI(g207), .SE(n10265), .CLK(n10452), .Q(
        g210) );
  SDFFX1 DFF_221_Q_reg ( .D(g30254), .SI(g210), .SE(n10265), .CLK(n10452), .Q(
        g249) );
  SDFFX1 DFF_222_Q_reg ( .D(g30257), .SI(g249), .SE(n10265), .CLK(n10452), .Q(
        g252) );
  SDFFX1 DFF_223_Q_reg ( .D(g30262), .SI(g252), .SE(n10265), .CLK(n10452), .Q(
        test_so14) );
  SDFFX1 DFF_224_Q_reg ( .D(g30245), .SI(test_si15), .SE(n10265), .CLK(n10452), 
        .Q(g213) );
  SDFFX1 DFF_225_Q_reg ( .D(g30246), .SI(g213), .SE(n10265), .CLK(n10452), .Q(
        g216) );
  SDFFX1 DFF_226_Q_reg ( .D(g30248), .SI(g216), .SE(n10265), .CLK(n10452), .Q(
        g219) );
  SDFFX1 DFF_227_Q_reg ( .D(g30258), .SI(g219), .SE(n10266), .CLK(n10453), .Q(
        g258) );
  SDFFX1 DFF_228_Q_reg ( .D(g30263), .SI(g258), .SE(n10266), .CLK(n10453), .Q(
        g261) );
  SDFFX1 DFF_229_Q_reg ( .D(g30268), .SI(g261), .SE(n10266), .CLK(n10453), .Q(
        g264) );
  SDFFX1 DFF_230_Q_reg ( .D(g30635), .SI(g264), .SE(n10266), .CLK(n10453), .Q(
        g222) );
  SDFFX1 DFF_231_Q_reg ( .D(g30636), .SI(g222), .SE(n10266), .CLK(n10453), .Q(
        g225) );
  SDFFX1 DFF_232_Q_reg ( .D(g30639), .SI(g225), .SE(n10266), .CLK(n10453), .Q(
        g228) );
  SDFFX1 DFF_233_Q_reg ( .D(g30661), .SI(g228), .SE(n10266), .CLK(n10453), .Q(
        g267) );
  SDFFX1 DFF_234_Q_reg ( .D(g30669), .SI(g267), .SE(n10266), .CLK(n10453), .Q(
        g270) );
  SDFFX1 DFF_235_Q_reg ( .D(g30675), .SI(g270), .SE(n10260), .CLK(n10447), .Q(
        g273) );
  SDFFX1 DFF_236_Q_reg ( .D(g25027), .SI(g273), .SE(n10260), .CLK(n10447), .Q(
        g92), .QN(n9891) );
  SDFFX1 DFF_237_Q_reg ( .D(g25932), .SI(g92), .SE(n10260), .CLK(n10447), .Q(
        g88), .QN(n10184) );
  SDFFX1 DFF_238_Q_reg ( .D(g26529), .SI(g88), .SE(n10260), .CLK(n10447), .Q(
        g83), .QN(n9890) );
  SDFFX1 DFF_239_Q_reg ( .D(g27120), .SI(g83), .SE(n10260), .CLK(n10447), .Q(
        test_so15), .QN(n10199) );
  SDFFX1 DFF_240_Q_reg ( .D(g27594), .SI(test_si16), .SE(n10260), .CLK(n10447), 
        .Q(g74), .QN(n9889) );
  SDFFX1 DFF_241_Q_reg ( .D(g28145), .SI(g74), .SE(n10260), .CLK(n10447), .Q(
        g70), .QN(n10167) );
  SDFFX1 DFF_242_Q_reg ( .D(g28634), .SI(g70), .SE(n10260), .CLK(n10447), .Q(
        g65), .QN(n9888) );
  SDFFX1 DFF_243_Q_reg ( .D(g29109), .SI(g65), .SE(n10260), .CLK(n10447), .Q(
        g61), .QN(n10176) );
  SDFFX1 DFF_244_Q_reg ( .D(g29353), .SI(g61), .SE(n10260), .CLK(n10447), .Q(
        g56), .QN(n9510) );
  SDFFX1 DFF_245_Q_reg ( .D(g29579), .SI(g56), .SE(n10260), .CLK(n10447), .Q(
        g52), .QN(n9356) );
  SDFFX1 DFF_246_Q_reg ( .D(n29), .SI(g52), .SE(n10261), .CLK(n10448), .Q(g180) );
  SDFFX1 DFF_247_Q_reg ( .D(g180), .SI(g180), .SE(n10261), .CLK(n10448), .Q(
        g5549) );
  SDFFX1 DFF_248_Q_reg ( .D(g5549), .SI(g5549), .SE(n10261), .CLK(n10448), .Q(
        g181), .QN(n10159) );
  SDFFX1 DFF_251_Q_reg ( .D(g6447), .SI(g6447), .SE(n10261), .CLK(n10448), .Q(
        n4640), .QN(n4506) );
  SDFFX1 DFF_252_Q_reg ( .D(g5549), .SI(n4640), .SE(n10261), .CLK(n10448), .Q(
        g309), .QN(n4388) );
  SDFFX1 DFF_253_Q_reg ( .D(g27253), .SI(g309), .SE(n10269), .CLK(n10456), .Q(
        g354), .QN(n9842) );
  SDFFX1 DFF_254_Q_reg ( .D(g27255), .SI(g354), .SE(n10269), .CLK(n10456), .Q(
        g343), .QN(n9841) );
  SDFFX1 DFF_255_Q_reg ( .D(g27258), .SI(g343), .SE(n10269), .CLK(n10456), .Q(
        test_so16), .QN(n10204) );
  SDFFX1 DFF_256_Q_reg ( .D(g27256), .SI(test_si17), .SE(n10269), .CLK(n10456), 
        .Q(g369), .QN(n9820) );
  SDFFX1 DFF_257_Q_reg ( .D(g27259), .SI(g369), .SE(n10269), .CLK(n10456), .Q(
        g358), .QN(n9819) );
  SDFFX1 DFF_258_Q_reg ( .D(g27265), .SI(g358), .SE(n10269), .CLK(n10456), .Q(
        g361), .QN(n9818) );
  SDFFX1 DFF_259_Q_reg ( .D(g27260), .SI(g361), .SE(n10269), .CLK(n10456), .Q(
        g384), .QN(n9564) );
  SDFFX1 DFF_260_Q_reg ( .D(g27266), .SI(g384), .SE(n10269), .CLK(n10456), .Q(
        g373), .QN(n9566) );
  SDFFX1 DFF_261_Q_reg ( .D(g27277), .SI(g373), .SE(n10269), .CLK(n10456), .Q(
        g376), .QN(n9565) );
  SDFFX1 DFF_262_Q_reg ( .D(g27267), .SI(g376), .SE(n10269), .CLK(n10456), .Q(
        g398), .QN(n9831) );
  SDFFX1 DFF_263_Q_reg ( .D(g27278), .SI(g398), .SE(n10269), .CLK(n10456), .Q(
        g388), .QN(n9830) );
  SDFFX1 DFF_264_Q_reg ( .D(g27293), .SI(g388), .SE(n10267), .CLK(n10454), .Q(
        g391), .QN(n9829) );
  SDFFX1 DFF_265_Q_reg ( .D(g28732), .SI(g391), .SE(n10267), .CLK(n10454), .Q(
        g408) );
  SDFFX1 DFF_266_Q_reg ( .D(g28735), .SI(g408), .SE(n10268), .CLK(n10455), .Q(
        g411) );
  SDFFX1 DFF_267_Q_reg ( .D(g28744), .SI(g411), .SE(n10268), .CLK(n10455), .Q(
        g414) );
  SDFFX1 DFF_268_Q_reg ( .D(g29194), .SI(g414), .SE(n10268), .CLK(n10455), .Q(
        g417) );
  SDFFX1 DFF_269_Q_reg ( .D(g29197), .SI(g417), .SE(n10268), .CLK(n10455), .Q(
        g420) );
  SDFFX1 DFF_270_Q_reg ( .D(g29201), .SI(g420), .SE(n10267), .CLK(n10454), .Q(
        g423) );
  SDFFX1 DFF_271_Q_reg ( .D(g28736), .SI(g423), .SE(n10267), .CLK(n10454), .Q(
        test_so17) );
  SDFFX1 DFF_272_Q_reg ( .D(g28745), .SI(test_si18), .SE(n10267), .CLK(n10454), 
        .Q(g428), .QN(n9874) );
  SDFFX1 DFF_273_Q_reg ( .D(g28754), .SI(g428), .SE(n10267), .CLK(n10454), .Q(
        g426), .QN(n9873) );
  SDFFX1 DFF_274_Q_reg ( .D(g26803), .SI(g426), .SE(n10267), .CLK(n10454), .Q(
        g429) );
  SDFFX1 DFF_275_Q_reg ( .D(g26804), .SI(g429), .SE(n10267), .CLK(n10454), .Q(
        g432) );
  SDFFX1 DFF_276_Q_reg ( .D(g26807), .SI(g432), .SE(n10267), .CLK(n10454), .Q(
        g435) );
  SDFFX1 DFF_277_Q_reg ( .D(g26805), .SI(g435), .SE(n10268), .CLK(n10455), .Q(
        g438) );
  SDFFX1 DFF_278_Q_reg ( .D(g26808), .SI(g438), .SE(n10268), .CLK(n10455), .Q(
        g441) );
  SDFFX1 DFF_279_Q_reg ( .D(g26812), .SI(g441), .SE(n10268), .CLK(n10455), .Q(
        g444) );
  SDFFX1 DFF_280_Q_reg ( .D(g27759), .SI(g444), .SE(n10268), .CLK(n10455), .Q(
        g448), .QN(n9872) );
  SDFFX1 DFF_281_Q_reg ( .D(g27760), .SI(g448), .SE(n10268), .CLK(n10455), .Q(
        g449), .QN(n9871) );
  SDFFX1 DFF_282_Q_reg ( .D(g27762), .SI(g449), .SE(n10267), .CLK(n10454), .Q(
        g447), .QN(n9870) );
  SDFFX1 DFF_283_Q_reg ( .D(g29606), .SI(g447), .SE(n10268), .CLK(n10455), .Q(
        g312), .QN(n9477) );
  SDFFX1 DFF_284_Q_reg ( .D(g29608), .SI(g312), .SE(n10268), .CLK(n10455), .Q(
        g313), .QN(n9476) );
  SDFFX1 DFF_285_Q_reg ( .D(g29611), .SI(g313), .SE(n10266), .CLK(n10453), .Q(
        g314), .QN(n9475) );
  SDFFX1 DFF_286_Q_reg ( .D(g30699), .SI(g314), .SE(n10267), .CLK(n10454), .Q(
        g315), .QN(n9474) );
  SDFFX1 DFF_287_Q_reg ( .D(g30700), .SI(g315), .SE(n10267), .CLK(n10454), .Q(
        test_so18), .QN(n10222) );
  SDFFX1 DFF_288_Q_reg ( .D(g30702), .SI(test_si19), .SE(n10259), .CLK(n10446), 
        .Q(g317), .QN(n9473) );
  SDFFX1 DFF_289_Q_reg ( .D(g30455), .SI(g317), .SE(n10261), .CLK(n10448), .Q(
        g318), .QN(n9472) );
  SDFFX1 DFF_290_Q_reg ( .D(g30468), .SI(g318), .SE(n10261), .CLK(n10448), .Q(
        g319), .QN(n9471) );
  SDFFX1 DFF_291_Q_reg ( .D(g30482), .SI(g319), .SE(n10260), .CLK(n10447), .Q(
        g320), .QN(n9470) );
  SDFFX1 DFF_292_Q_reg ( .D(g29167), .SI(g320), .SE(n10270), .CLK(n10457), .Q(
        g322) );
  SDFFX1 DFF_293_Q_reg ( .D(g29169), .SI(g322), .SE(n10270), .CLK(n10457), .Q(
        g323) );
  SDFFX1 DFF_294_Q_reg ( .D(g29172), .SI(g323), .SE(n10270), .CLK(n10457), .Q(
        g321) );
  SDFFX1 DFF_295_Q_reg ( .D(g26655), .SI(g321), .SE(n10270), .CLK(n10457), .Q(
        g403), .QN(n9869) );
  SDFFX1 DFF_296_Q_reg ( .D(g26659), .SI(g403), .SE(n10270), .CLK(n10457), .Q(
        g404), .QN(n9868) );
  SDFFX1 DFF_297_Q_reg ( .D(g26664), .SI(g404), .SE(n10271), .CLK(n10458), .Q(
        g402), .QN(n9867) );
  SDFFX1 DFF_298_Q_reg ( .D(n4290), .SI(g402), .SE(n10341), .CLK(n10528), .Q(
        g450) );
  SDFFX1 DFF_299_Q_reg ( .D(g450), .SI(g450), .SE(n10341), .CLK(n10528), .Q(
        n8066), .QN(DFF_299_n1) );
  SDFFX1 DFF_300_Q_reg ( .D(n4569), .SI(n8066), .SE(n10341), .CLK(n10528), .Q(
        g452) );
  SDFFX1 DFF_301_Q_reg ( .D(g452), .SI(g452), .SE(n10341), .CLK(n10528), .Q(
        n8065), .QN(DFF_301_n1) );
  SDFFX1 DFF_302_Q_reg ( .D(n4561), .SI(n8065), .SE(n10342), .CLK(n10529), .Q(
        g454) );
  SDFFX1 DFF_303_Q_reg ( .D(g454), .SI(g454), .SE(n10342), .CLK(n10529), .Q(
        test_so19), .QN(DFF_303_n1) );
  SDFFX1 DFF_304_Q_reg ( .D(n4328), .SI(test_si20), .SE(n10258), .CLK(n10445), 
        .Q(g280) );
  SDFFX1 DFF_305_Q_reg ( .D(g280), .SI(g280), .SE(n10258), .CLK(n10445), .Q(
        n8062), .QN(DFF_305_n1) );
  SDFFX1 DFF_306_Q_reg ( .D(n4392), .SI(n8062), .SE(n10258), .CLK(n10445), .Q(
        g282) );
  SDFFX1 DFF_307_Q_reg ( .D(g282), .SI(g282), .SE(n10258), .CLK(n10445), .Q(
        n8061), .QN(DFF_307_n1) );
  SDFFX1 DFF_308_Q_reg ( .D(n4322), .SI(n8061), .SE(n10259), .CLK(n10446), .Q(
        g284) );
  SDFFX1 DFF_309_Q_reg ( .D(g284), .SI(g284), .SE(n10259), .CLK(n10446), .Q(
        n8060), .QN(DFF_309_n1) );
  SDFFX1 DFF_310_Q_reg ( .D(n4376), .SI(n8060), .SE(n10259), .CLK(n10446), .Q(
        g286) );
  SDFFX1 DFF_311_Q_reg ( .D(g286), .SI(g286), .SE(n10259), .CLK(n10446), .Q(
        n8059), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(n4380), .SI(n8059), .SE(n10259), .CLK(n10446), .Q(
        g288) );
  SDFFX1 DFF_313_Q_reg ( .D(g288), .SI(g288), .SE(n10259), .CLK(n10446), .Q(
        n8058), .QN(DFF_313_n1) );
  SDFFX1 DFF_314_Q_reg ( .D(g2857), .SI(n8058), .SE(n10259), .CLK(n10446), .Q(
        g290) );
  SDFFX1 DFF_315_Q_reg ( .D(g290), .SI(g290), .SE(n10259), .CLK(n10446), .Q(
        n8057), .QN(n4485) );
  SDFFX1 DFF_316_Q_reg ( .D(n4282), .SI(n8057), .SE(n10268), .CLK(n10455), .Q(
        n8056), .QN(n18263) );
  SDFFX1 DFF_317_Q_reg ( .D(g21346), .SI(n8056), .SE(n10280), .CLK(n10467), 
        .Q(g305), .QN(n9616) );
  SDFFX1 DFF_328_Q_reg ( .D(n4278), .SI(g305), .SE(n10271), .CLK(n10458), .Q(
        n8055), .QN(DFF_328_n1) );
  SDFFX1 DFF_329_Q_reg ( .D(g354), .SI(n8055), .SE(n10271), .CLK(n10458), .Q(
        test_so20) );
  SDFFX1 DFF_330_Q_reg ( .D(test_so20), .SI(test_si21), .SE(n10271), .CLK(
        n10458), .Q(g349) );
  SDFFX1 DFF_331_Q_reg ( .D(g343), .SI(g349), .SE(n10271), .CLK(n10458), .Q(
        g350) );
  SDFFX1 DFF_332_Q_reg ( .D(g350), .SI(g350), .SE(n10271), .CLK(n10458), .Q(
        g351) );
  SDFFX1 DFF_333_Q_reg ( .D(test_so16), .SI(g351), .SE(n10271), .CLK(n10458), 
        .Q(g352) );
  SDFFX1 DFF_334_Q_reg ( .D(g352), .SI(g352), .SE(n10271), .CLK(n10458), .Q(
        g353) );
  SDFFX1 DFF_335_Q_reg ( .D(g369), .SI(g353), .SE(n10271), .CLK(n10458), .Q(
        g357) );
  SDFFX1 DFF_336_Q_reg ( .D(g357), .SI(g357), .SE(n10271), .CLK(n10458), .Q(
        g364) );
  SDFFX1 DFF_337_Q_reg ( .D(g358), .SI(g364), .SE(n10271), .CLK(n10458), .Q(
        g365) );
  SDFFX1 DFF_338_Q_reg ( .D(g365), .SI(g365), .SE(n10271), .CLK(n10458), .Q(
        g366) );
  SDFFX1 DFF_339_Q_reg ( .D(g361), .SI(g366), .SE(n10272), .CLK(n10459), .Q(
        g367) );
  SDFFX1 DFF_340_Q_reg ( .D(g367), .SI(g367), .SE(n10272), .CLK(n10459), .Q(
        g368) );
  SDFFX1 DFF_341_Q_reg ( .D(g384), .SI(g368), .SE(n10272), .CLK(n10459), .Q(
        g372) );
  SDFFX1 DFF_342_Q_reg ( .D(g372), .SI(g372), .SE(n10272), .CLK(n10459), .Q(
        g379) );
  SDFFX1 DFF_343_Q_reg ( .D(g373), .SI(g379), .SE(n10272), .CLK(n10459), .Q(
        g380) );
  SDFFX1 DFF_344_Q_reg ( .D(g380), .SI(g380), .SE(n10272), .CLK(n10459), .Q(
        g381) );
  SDFFX1 DFF_345_Q_reg ( .D(g376), .SI(g381), .SE(n10272), .CLK(n10459), .Q(
        test_so21) );
  SDFFX1 DFF_346_Q_reg ( .D(test_so21), .SI(test_si22), .SE(n10272), .CLK(
        n10459), .Q(g383) );
  SDFFX1 DFF_347_Q_reg ( .D(g398), .SI(g383), .SE(n10272), .CLK(n10459), .Q(
        g387) );
  SDFFX1 DFF_348_Q_reg ( .D(g387), .SI(g387), .SE(n10272), .CLK(n10459), .Q(
        g394) );
  SDFFX1 DFF_349_Q_reg ( .D(g388), .SI(g394), .SE(n10272), .CLK(n10459), .Q(
        g395) );
  SDFFX1 DFF_350_Q_reg ( .D(g395), .SI(g395), .SE(n10272), .CLK(n10459), .Q(
        g396) );
  SDFFX1 DFF_351_Q_reg ( .D(g391), .SI(g396), .SE(n10273), .CLK(n10460), .Q(
        g397) );
  SDFFX1 DFF_352_Q_reg ( .D(g397), .SI(g397), .SE(n10273), .CLK(n10460), .Q(
        g324) );
  SDFFX1 DFF_353_Q_reg ( .D(n4598), .SI(g324), .SE(n10273), .CLK(n10460), .Q(
        g5629) );
  SDFFX1 DFF_354_Q_reg ( .D(g5629), .SI(g5629), .SE(n10273), .CLK(n10460), .Q(
        g5648) );
  SDFFX1 DFF_355_Q_reg ( .D(g5648), .SI(g5648), .SE(n10273), .CLK(n10460), .Q(
        g337) );
  SDFFX1 DFF_356_Q_reg ( .D(n4598), .SI(g337), .SE(n10273), .CLK(n10460), .Q(
        g6485), .QN(n4298) );
  SDFFX1 DFF_357_Q_reg ( .D(g6485), .SI(g6485), .SE(n10273), .CLK(n10460), .Q(
        g6642), .QN(n4372) );
  SDFFX1 DFF_358_Q_reg ( .D(g6642), .SI(g6642), .SE(n10273), .CLK(n10460), .Q(
        g550), .QN(n4313) );
  SDFFX1 DFF_359_Q_reg ( .D(g21842), .SI(g550), .SE(n10273), .CLK(n10460), .Q(
        g554), .QN(n10123) );
  SDFFX1 DFF_360_Q_reg ( .D(g18678), .SI(g554), .SE(n10273), .CLK(n10460), .Q(
        g557), .QN(n4360) );
  SDFFX1 DFF_361_Q_reg ( .D(g18726), .SI(g557), .SE(n10273), .CLK(n10460), .Q(
        test_so22), .QN(n10200) );
  SDFFX1 DFF_362_Q_reg ( .D(n634), .SI(test_si23), .SE(n10273), .CLK(n10460), 
        .Q(g513) );
  SDFFX1 DFF_363_Q_reg ( .D(g513), .SI(g513), .SE(n10274), .CLK(n10461), .Q(
        g523) );
  SDFFX1 DFF_364_Q_reg ( .D(g523), .SI(g523), .SE(n10274), .CLK(n10461), .Q(
        g524) );
  SDFFX1 DFF_365_Q_reg ( .D(g455), .SI(g524), .SE(n10274), .CLK(n10461), .Q(
        g564) );
  SDFFX1 DFF_366_Q_reg ( .D(g564), .SI(g564), .SE(n10274), .CLK(n10461), .Q(
        g569) );
  SDFFX1 DFF_367_Q_reg ( .D(g458), .SI(g569), .SE(n10274), .CLK(n10461), .Q(
        g570) );
  SDFFX1 DFF_368_Q_reg ( .D(g570), .SI(g570), .SE(n10274), .CLK(n10461), .Q(
        g571) );
  SDFFX1 DFF_369_Q_reg ( .D(g461), .SI(g571), .SE(n10274), .CLK(n10461), .Q(
        g572) );
  SDFFX1 DFF_370_Q_reg ( .D(g572), .SI(g572), .SE(n10274), .CLK(n10461), .Q(
        g573) );
  SDFFX1 DFF_371_Q_reg ( .D(g465), .SI(g573), .SE(n10274), .CLK(n10461), .Q(
        g574) );
  SDFFX1 DFF_372_Q_reg ( .D(g574), .SI(g574), .SE(n10274), .CLK(n10461), .Q(
        g565) );
  SDFFX1 DFF_373_Q_reg ( .D(test_so24), .SI(g565), .SE(n10274), .CLK(n10461), 
        .Q(g566) );
  SDFFX1 DFF_374_Q_reg ( .D(g566), .SI(g566), .SE(n10274), .CLK(n10461), .Q(
        g567) );
  SDFFX1 DFF_375_Q_reg ( .D(g471), .SI(g567), .SE(n10275), .CLK(n10462), .Q(
        g568) );
  SDFFX1 DFF_376_Q_reg ( .D(g568), .SI(g568), .SE(n10275), .CLK(n10462), .Q(
        g489) );
  SDFFX1 DFF_377_Q_reg ( .D(g2950), .SI(g489), .SE(n10275), .CLK(n10462), .Q(
        test_so23), .QN(n10190) );
  SDFFX1 DFF_378_Q_reg ( .D(test_so23), .SI(test_si24), .SE(n10275), .CLK(
        n10462), .Q(g7956), .QN(n4461) );
  SDFFX1 DFF_379_Q_reg ( .D(g7956), .SI(g7956), .SE(n10275), .CLK(n10462), .Q(
        g485), .QN(n4466) );
  SDFFX1 DFF_380_Q_reg ( .D(g23067), .SI(g485), .SE(n10275), .CLK(n10462), .Q(
        g486) );
  SDFFX1 DFF_381_Q_reg ( .D(g23093), .SI(g486), .SE(n10275), .CLK(n10462), .Q(
        g487) );
  SDFFX1 DFF_382_Q_reg ( .D(g23117), .SI(g487), .SE(n10275), .CLK(n10462), .Q(
        g488) );
  SDFFX1 DFF_383_Q_reg ( .D(g23385), .SI(g488), .SE(n10275), .CLK(n10462), .Q(
        g455) );
  SDFFX1 DFF_384_Q_reg ( .D(g23399), .SI(g455), .SE(n10275), .CLK(n10462), .Q(
        g458) );
  SDFFX1 DFF_385_Q_reg ( .D(g24174), .SI(g458), .SE(n10275), .CLK(n10462), .Q(
        g461) );
  SDFFX1 DFF_386_Q_reg ( .D(g24178), .SI(g461), .SE(n10276), .CLK(n10463), .Q(
        g477) );
  SDFFX1 DFF_387_Q_reg ( .D(g24207), .SI(g477), .SE(n10276), .CLK(n10463), .Q(
        g478) );
  SDFFX1 DFF_388_Q_reg ( .D(g24216), .SI(g478), .SE(n10276), .CLK(n10463), .Q(
        g479) );
  SDFFX1 DFF_389_Q_reg ( .D(g23092), .SI(g479), .SE(n10276), .CLK(n10463), .Q(
        g480) );
  SDFFX1 DFF_390_Q_reg ( .D(g23000), .SI(g480), .SE(n10276), .CLK(n10463), .Q(
        g484) );
  SDFFX1 DFF_391_Q_reg ( .D(g23022), .SI(g484), .SE(n10276), .CLK(n10463), .Q(
        g464) );
  SDFFX1 DFF_392_Q_reg ( .D(g24206), .SI(g464), .SE(n10276), .CLK(n10463), .Q(
        g465) );
  SDFFX1 DFF_393_Q_reg ( .D(g24215), .SI(g465), .SE(n10276), .CLK(n10463), .Q(
        test_so24) );
  SDFFX1 DFF_394_Q_reg ( .D(g24228), .SI(test_si25), .SE(n10275), .CLK(n10462), 
        .Q(g471) );
  SDFFX1 DFF_395_Q_reg ( .D(n610), .SI(g471), .SE(n10276), .CLK(n10463), .Q(
        g528) );
  SDFFX1 DFF_396_Q_reg ( .D(g528), .SI(g528), .SE(n10276), .CLK(n10463), .Q(
        g535) );
  SDFFX1 DFF_397_Q_reg ( .D(g535), .SI(g535), .SE(n10276), .CLK(n10463), .Q(
        g542) );
  SDFFX1 DFF_398_Q_reg ( .D(g13149), .SI(g542), .SE(n10276), .CLK(n10463), .Q(
        g543) );
  SDFFX1 DFF_399_Q_reg ( .D(g543), .SI(g543), .SE(n10277), .CLK(n10464), .Q(
        g544) );
  SDFFX1 DFF_400_Q_reg ( .D(g21851), .SI(g544), .SE(n10277), .CLK(n10464), .Q(
        g548) );
  SDFFX1 DFF_401_Q_reg ( .D(g13111), .SI(g548), .SE(n10277), .CLK(n10464), .Q(
        g549) );
  SDFFX1 DFF_402_Q_reg ( .D(g549), .SI(g549), .SE(n10277), .CLK(n10464), .Q(
        g499), .QN(n4541) );
  SDFFX1 DFF_403_Q_reg ( .D(g13160), .SI(g499), .SE(n10277), .CLK(n10464), .Q(
        g558) );
  SDFFX1 DFF_404_Q_reg ( .D(g558), .SI(g558), .SE(n10277), .CLK(n10464), .Q(
        g559) );
  SDFFX1 DFF_405_Q_reg ( .D(g27261), .SI(g559), .SE(n10278), .CLK(n10465), .Q(
        g576), .QN(n9520) );
  SDFFX1 DFF_406_Q_reg ( .D(g27268), .SI(g576), .SE(n10278), .CLK(n10465), .Q(
        g577), .QN(n9522) );
  SDFFX1 DFF_407_Q_reg ( .D(g27279), .SI(g577), .SE(n10278), .CLK(n10465), .Q(
        g575), .QN(n9521) );
  SDFFX1 DFF_408_Q_reg ( .D(g27269), .SI(g575), .SE(n10278), .CLK(n10465), .Q(
        g579), .QN(n9532) );
  SDFFX1 DFF_409_Q_reg ( .D(g27280), .SI(g579), .SE(n10278), .CLK(n10465), .Q(
        test_so25) );
  SDFFX1 DFF_410_Q_reg ( .D(g27294), .SI(test_si26), .SE(n10277), .CLK(n10464), 
        .Q(g578), .QN(n9533) );
  SDFFX1 DFF_411_Q_reg ( .D(g27281), .SI(g578), .SE(n10277), .CLK(n10464), .Q(
        g582), .QN(n9364) );
  SDFFX1 DFF_412_Q_reg ( .D(g27295), .SI(g582), .SE(n10277), .CLK(n10464), .Q(
        g583), .QN(n9366) );
  SDFFX1 DFF_413_Q_reg ( .D(g27311), .SI(g583), .SE(n10277), .CLK(n10464), .Q(
        g581), .QN(n9365) );
  SDFFX1 DFF_414_Q_reg ( .D(g27296), .SI(g581), .SE(n10277), .CLK(n10464), .Q(
        g585), .QN(n9542) );
  SDFFX1 DFF_415_Q_reg ( .D(g27312), .SI(g585), .SE(n10278), .CLK(n10465), .Q(
        g586), .QN(n9544) );
  SDFFX1 DFF_416_Q_reg ( .D(g27327), .SI(g586), .SE(n10278), .CLK(n10465), .Q(
        g584), .QN(n9543) );
  SDFFX1 DFF_417_Q_reg ( .D(g24491), .SI(g584), .SE(n10278), .CLK(n10465), .Q(
        g587) );
  SDFFX1 DFF_418_Q_reg ( .D(g24498), .SI(g587), .SE(n10278), .CLK(n10465), .Q(
        g590) );
  SDFFX1 DFF_419_Q_reg ( .D(g24507), .SI(g590), .SE(n10278), .CLK(n10465), .Q(
        g593) );
  SDFFX1 DFF_420_Q_reg ( .D(g24499), .SI(g593), .SE(n10278), .CLK(n10465), .Q(
        g596) );
  SDFFX1 DFF_421_Q_reg ( .D(g24508), .SI(g596), .SE(n10278), .CLK(n10465), .Q(
        g599) );
  SDFFX1 DFF_422_Q_reg ( .D(g24519), .SI(g599), .SE(n10279), .CLK(n10466), .Q(
        g602) );
  SDFFX1 DFF_423_Q_reg ( .D(g28345), .SI(g602), .SE(n10279), .CLK(n10466), .Q(
        g614) );
  SDFFX1 DFF_424_Q_reg ( .D(g28349), .SI(g614), .SE(n10279), .CLK(n10466), .Q(
        g617) );
  SDFFX1 DFF_425_Q_reg ( .D(g28353), .SI(g617), .SE(n10277), .CLK(n10464), .Q(
        test_so26) );
  SDFFX1 DFF_426_Q_reg ( .D(g28342), .SI(test_si27), .SE(n10279), .CLK(n10466), 
        .Q(g605) );
  SDFFX1 DFF_427_Q_reg ( .D(g28344), .SI(g605), .SE(n10279), .CLK(n10466), .Q(
        g608) );
  SDFFX1 DFF_428_Q_reg ( .D(g28348), .SI(g608), .SE(n10279), .CLK(n10466), .Q(
        g611) );
  SDFFX1 DFF_429_Q_reg ( .D(g26541), .SI(g611), .SE(n10279), .CLK(n10466), .Q(
        g490) );
  SDFFX1 DFF_430_Q_reg ( .D(g26545), .SI(g490), .SE(n10279), .CLK(n10466), .Q(
        g493) );
  SDFFX1 DFF_431_Q_reg ( .D(g26553), .SI(g493), .SE(n10279), .CLK(n10466), .Q(
        g496) );
  SDFFX1 DFF_432_Q_reg ( .D(g499), .SI(g496), .SE(n10279), .CLK(n10466), .Q(
        g506), .QN(n4570) );
  SDFFX1 DFF_433_Q_reg ( .D(g22578), .SI(g506), .SE(n10279), .CLK(n10466), .Q(
        n4571) );
  SDFFX1 DFF_442_Q_reg ( .D(n633), .SI(n4571), .SE(n10279), .CLK(n10466), .Q(
        g16297) );
  SDFFX1 DFF_443_Q_reg ( .D(g16297), .SI(g16297), .SE(n10280), .CLK(n10467), 
        .Q(g525), .QN(n9898) );
  SDFFX1 DFF_444_Q_reg ( .D(DFF_299_n1), .SI(g525), .SE(n10342), .CLK(n10529), 
        .Q(n8047) );
  SDFFX1 DFF_445_Q_reg ( .D(DFF_301_n1), .SI(n8047), .SE(n10342), .CLK(n10529), 
        .Q(n8046) );
  SDFFX1 DFF_446_Q_reg ( .D(DFF_303_n1), .SI(n8046), .SE(n10342), .CLK(n10529), 
        .Q(n8045) );
  SDFFX1 DFF_447_Q_reg ( .D(DFF_305_n1), .SI(n8045), .SE(n10342), .CLK(n10529), 
        .Q(n8044) );
  SDFFX1 DFF_448_Q_reg ( .D(DFF_307_n1), .SI(n8044), .SE(n10343), .CLK(n10530), 
        .Q(n8043) );
  SDFFX1 DFF_449_Q_reg ( .D(DFF_309_n1), .SI(n8043), .SE(n10343), .CLK(n10530), 
        .Q(test_so27) );
  SDFFX1 DFF_450_Q_reg ( .D(DFF_311_n1), .SI(test_si28), .SE(n10259), .CLK(
        n10446), .Q(g536) );
  SDFFX1 DFF_451_Q_reg ( .D(DFF_313_n1), .SI(g536), .SE(n10259), .CLK(n10446), 
        .Q(g537) );
  SDFFX1 DFF_452_Q_reg ( .D(g24059), .SI(g537), .SE(n10280), .CLK(n10467), .Q(
        g538), .QN(n4492) );
  SDFFX1 DFF_453_Q_reg ( .D(n4485), .SI(g538), .SE(n10280), .CLK(n10467), .Q(
        n8040) );
  SDFFX1 DFF_455_Q_reg ( .D(g6677), .SI(g6677), .SE(n10280), .CLK(n10467), .Q(
        g6911), .QN(n4359) );
  SDFFX1 DFF_456_Q_reg ( .D(g6911), .SI(g6911), .SE(n10280), .CLK(n10467), .Q(
        g629), .QN(n4295) );
  SDFFX1 DFF_457_Q_reg ( .D(g16654), .SI(g629), .SE(n10280), .CLK(n10467), .Q(
        g630), .QN(n10153) );
  SDFFX1 DFF_458_Q_reg ( .D(g20314), .SI(g630), .SE(n10280), .CLK(n10467), .Q(
        g659), .QN(n4429) );
  SDFFX1 DFF_459_Q_reg ( .D(g20682), .SI(g659), .SE(n10280), .CLK(n10467), .Q(
        g640), .QN(n4404) );
  SDFFX1 DFF_460_Q_reg ( .D(g23136), .SI(g640), .SE(n10280), .CLK(n10467), .Q(
        g633), .QN(n4478) );
  SDFFX1 DFF_461_Q_reg ( .D(g23324), .SI(g633), .SE(n10280), .CLK(n10467), .Q(
        g653), .QN(n4422) );
  SDFFX1 DFF_462_Q_reg ( .D(g24426), .SI(g653), .SE(n10281), .CLK(n10468), .Q(
        g646), .QN(n4414) );
  SDFFX1 DFF_463_Q_reg ( .D(g25185), .SI(g646), .SE(n10281), .CLK(n10468), .Q(
        g660), .QN(n4403) );
  SDFFX1 DFF_464_Q_reg ( .D(g26660), .SI(g660), .SE(n10281), .CLK(n10468), .Q(
        g672), .QN(n4413) );
  SDFFX1 DFF_465_Q_reg ( .D(g26776), .SI(g672), .SE(n10281), .CLK(n10468), .Q(
        test_so28), .QN(n10193) );
  SDFFX1 DFF_466_Q_reg ( .D(g27672), .SI(test_si29), .SE(n10281), .CLK(n10468), 
        .Q(g679), .QN(n4477) );
  SDFFX1 DFF_467_Q_reg ( .D(g28199), .SI(g679), .SE(n10281), .CLK(n10468), .Q(
        g686), .QN(n4396) );
  SDFFX1 DFF_468_Q_reg ( .D(g28668), .SI(g686), .SE(n10281), .CLK(n10468), .Q(
        g692), .QN(n4418) );
  SDFFX1 DFF_469_Q_reg ( .D(g20875), .SI(g692), .SE(n10281), .CLK(n10468), .Q(
        g699), .QN(n10010) );
  SDFFX1 DFF_470_Q_reg ( .D(g20879), .SI(g699), .SE(n10281), .CLK(n10468), .Q(
        g700), .QN(n10009) );
  SDFFX1 DFF_471_Q_reg ( .D(g20891), .SI(g700), .SE(n10281), .CLK(n10468), .Q(
        g698), .QN(n10048) );
  SDFFX1 DFF_472_Q_reg ( .D(g20880), .SI(g698), .SE(n10281), .CLK(n10468), .Q(
        g702), .QN(n10008) );
  SDFFX1 DFF_473_Q_reg ( .D(g20892), .SI(g702), .SE(n10282), .CLK(n10469), .Q(
        g703), .QN(n10007) );
  SDFFX1 DFF_474_Q_reg ( .D(g20901), .SI(g703), .SE(n10282), .CLK(n10469), .Q(
        g701), .QN(n10047) );
  SDFFX1 DFF_475_Q_reg ( .D(g20893), .SI(g701), .SE(n10282), .CLK(n10469), .Q(
        g705), .QN(n10006) );
  SDFFX1 DFF_476_Q_reg ( .D(g20902), .SI(g705), .SE(n10282), .CLK(n10469), .Q(
        g706), .QN(n10005) );
  SDFFX1 DFF_477_Q_reg ( .D(g20921), .SI(g706), .SE(n10282), .CLK(n10469), .Q(
        g704), .QN(n10046) );
  SDFFX1 DFF_478_Q_reg ( .D(g20903), .SI(g704), .SE(n10283), .CLK(n10470), .Q(
        g708), .QN(n10004) );
  SDFFX1 DFF_479_Q_reg ( .D(g20922), .SI(g708), .SE(n10283), .CLK(n10470), .Q(
        g709), .QN(n10003) );
  SDFFX1 DFF_480_Q_reg ( .D(g20944), .SI(g709), .SE(n10283), .CLK(n10470), .Q(
        g707), .QN(n10045) );
  SDFFX1 DFF_481_Q_reg ( .D(g20923), .SI(g707), .SE(n10283), .CLK(n10470), .Q(
        test_so29) );
  SDFFX1 DFF_482_Q_reg ( .D(g20945), .SI(test_si30), .SE(n10281), .CLK(n10468), 
        .Q(g712), .QN(n10002) );
  SDFFX1 DFF_483_Q_reg ( .D(g20966), .SI(g712), .SE(n10283), .CLK(n10470), .Q(
        g710), .QN(n10044) );
  SDFFX1 DFF_484_Q_reg ( .D(g20946), .SI(g710), .SE(n10283), .CLK(n10470), .Q(
        g714), .QN(n10001) );
  SDFFX1 DFF_485_Q_reg ( .D(g20967), .SI(g714), .SE(n10283), .CLK(n10470), .Q(
        g715), .QN(n10000) );
  SDFFX1 DFF_486_Q_reg ( .D(g20989), .SI(g715), .SE(n10283), .CLK(n10470), .Q(
        g713), .QN(n10043) );
  SDFFX1 DFF_487_Q_reg ( .D(g20968), .SI(g713), .SE(n10283), .CLK(n10470), .Q(
        g717), .QN(n9999) );
  SDFFX1 DFF_488_Q_reg ( .D(g20990), .SI(g717), .SE(n10283), .CLK(n10470), .Q(
        g718), .QN(n9998) );
  SDFFX1 DFF_489_Q_reg ( .D(g21009), .SI(g718), .SE(n10283), .CLK(n10470), .Q(
        g716), .QN(n10042) );
  SDFFX1 DFF_490_Q_reg ( .D(g20991), .SI(g716), .SE(n10283), .CLK(n10470), .Q(
        g720), .QN(n9997) );
  SDFFX1 DFF_491_Q_reg ( .D(g21010), .SI(g720), .SE(n10284), .CLK(n10471), .Q(
        g721), .QN(n9996) );
  SDFFX1 DFF_492_Q_reg ( .D(g21031), .SI(g721), .SE(n10284), .CLK(n10471), .Q(
        g719), .QN(n10041) );
  SDFFX1 DFF_493_Q_reg ( .D(g21011), .SI(g719), .SE(n10284), .CLK(n10471), .Q(
        g723), .QN(n9995) );
  SDFFX1 DFF_494_Q_reg ( .D(g21032), .SI(g723), .SE(n10284), .CLK(n10471), .Q(
        g724), .QN(n9994) );
  SDFFX1 DFF_495_Q_reg ( .D(g21051), .SI(g724), .SE(n10284), .CLK(n10471), .Q(
        g722), .QN(n10040) );
  SDFFX1 DFF_496_Q_reg ( .D(g20876), .SI(g722), .SE(n10284), .CLK(n10471), .Q(
        g726), .QN(n9993) );
  SDFFX1 DFF_497_Q_reg ( .D(g20881), .SI(g726), .SE(n10284), .CLK(n10471), .Q(
        test_so30) );
  SDFFX1 DFF_498_Q_reg ( .D(g20894), .SI(test_si31), .SE(n10282), .CLK(n10469), 
        .Q(g725), .QN(n10039) );
  SDFFX1 DFF_499_Q_reg ( .D(g20924), .SI(g725), .SE(n10282), .CLK(n10469), .Q(
        g729), .QN(n9754) );
  SDFFX1 DFF_500_Q_reg ( .D(g20947), .SI(g729), .SE(n10282), .CLK(n10469), .Q(
        g730), .QN(n9746) );
  SDFFX1 DFF_501_Q_reg ( .D(g20969), .SI(g730), .SE(n10282), .CLK(n10469), .Q(
        g728), .QN(n9808) );
  SDFFX1 DFF_502_Q_reg ( .D(g20948), .SI(g728), .SE(n10282), .CLK(n10469), .Q(
        g732), .QN(n9753) );
  SDFFX1 DFF_503_Q_reg ( .D(g20970), .SI(g732), .SE(n10282), .CLK(n10469), .Q(
        g733), .QN(n9745) );
  SDFFX1 DFF_504_Q_reg ( .D(g20992), .SI(g733), .SE(n10282), .CLK(n10469), .Q(
        g731), .QN(n9807) );
  SDFFX1 DFF_505_Q_reg ( .D(g25260), .SI(g731), .SE(n10284), .CLK(n10471), .Q(
        g735) );
  SDFFX1 DFF_506_Q_reg ( .D(g25262), .SI(g735), .SE(n10284), .CLK(n10471), .Q(
        g736) );
  SDFFX1 DFF_507_Q_reg ( .D(g25266), .SI(g736), .SE(n10284), .CLK(n10471), .Q(
        g734) );
  SDFFX1 DFF_508_Q_reg ( .D(g22218), .SI(g734), .SE(n10284), .CLK(n10471), .Q(
        g738) );
  SDFFX1 DFF_509_Q_reg ( .D(g22231), .SI(g738), .SE(n10284), .CLK(n10471), .Q(
        g739) );
  SDFFX1 DFF_510_Q_reg ( .D(g22242), .SI(g739), .SE(n10285), .CLK(n10472), .Q(
        g737) );
  SDFFX1 DFF_511_Q_reg ( .D(g2950), .SI(g737), .SE(n10285), .CLK(n10472), .Q(
        g6368), .QN(n4323) );
  SDFFX1 DFF_512_Q_reg ( .D(g6368), .SI(g6368), .SE(n10285), .CLK(n10472), .Q(
        g6518), .QN(n4312) );
  SDFFX1 DFF_513_Q_reg ( .D(g6518), .SI(g6518), .SE(n10285), .CLK(n10472), .Q(
        test_so31), .QN(n10188) );
  SDFFX1 DFF_514_Q_reg ( .D(g22126), .SI(test_si32), .SE(n10286), .CLK(n10473), 
        .Q(g818), .QN(n10096) );
  SDFFX1 DFF_515_Q_reg ( .D(g22145), .SI(g818), .SE(n10289), .CLK(n10476), .Q(
        g819), .QN(n10095) );
  SDFFX1 DFF_516_Q_reg ( .D(g22162), .SI(g819), .SE(n10289), .CLK(n10476), .Q(
        g817), .QN(n9729) );
  SDFFX1 DFF_517_Q_reg ( .D(g22146), .SI(g817), .SE(n10286), .CLK(n10473), .Q(
        g821), .QN(n10094) );
  SDFFX1 DFF_518_Q_reg ( .D(g22163), .SI(g821), .SE(n10289), .CLK(n10476), .Q(
        g822), .QN(n10093) );
  SDFFX1 DFF_519_Q_reg ( .D(g22177), .SI(g822), .SE(n10289), .CLK(n10476), .Q(
        g820), .QN(n9728) );
  SDFFX1 DFF_520_Q_reg ( .D(g22029), .SI(g820), .SE(n10290), .CLK(n10477), .Q(
        g830), .QN(n10092) );
  SDFFX1 DFF_521_Q_reg ( .D(g22033), .SI(g830), .SE(n10290), .CLK(n10477), .Q(
        g831), .QN(n10091) );
  SDFFX1 DFF_522_Q_reg ( .D(g22040), .SI(g831), .SE(n10290), .CLK(n10477), .Q(
        g829), .QN(n9727) );
  SDFFX1 DFF_523_Q_reg ( .D(g22034), .SI(g829), .SE(n10290), .CLK(n10477), .Q(
        g833), .QN(n10090) );
  SDFFX1 DFF_524_Q_reg ( .D(g22041), .SI(g833), .SE(n10290), .CLK(n10477), .Q(
        g834), .QN(n10089) );
  SDFFX1 DFF_525_Q_reg ( .D(g22054), .SI(g834), .SE(n10290), .CLK(n10477), .Q(
        g832), .QN(n9726) );
  SDFFX1 DFF_526_Q_reg ( .D(g22042), .SI(g832), .SE(n10290), .CLK(n10477), .Q(
        g836), .QN(n10088) );
  SDFFX1 DFF_527_Q_reg ( .D(g22055), .SI(g836), .SE(n10290), .CLK(n10477), .Q(
        g837), .QN(n10087) );
  SDFFX1 DFF_528_Q_reg ( .D(g22066), .SI(g837), .SE(n10290), .CLK(n10477), .Q(
        g835), .QN(n9725) );
  SDFFX1 DFF_529_Q_reg ( .D(g22056), .SI(g835), .SE(n10290), .CLK(n10477), .Q(
        test_so32), .QN(n10212) );
  SDFFX1 DFF_530_Q_reg ( .D(g22067), .SI(test_si33), .SE(n10288), .CLK(n10475), 
        .Q(g840), .QN(n10086) );
  SDFFX1 DFF_531_Q_reg ( .D(g22087), .SI(g840), .SE(n10288), .CLK(n10475), .Q(
        g838), .QN(n9724) );
  SDFFX1 DFF_532_Q_reg ( .D(g22068), .SI(g838), .SE(n10288), .CLK(n10475), .Q(
        g842), .QN(n10085) );
  SDFFX1 DFF_533_Q_reg ( .D(g22088), .SI(g842), .SE(n10288), .CLK(n10475), .Q(
        g843), .QN(n10084) );
  SDFFX1 DFF_534_Q_reg ( .D(g22104), .SI(g843), .SE(n10288), .CLK(n10475), .Q(
        g841), .QN(n9723) );
  SDFFX1 DFF_535_Q_reg ( .D(g22089), .SI(g841), .SE(n10288), .CLK(n10475), .Q(
        g845), .QN(n10083) );
  SDFFX1 DFF_536_Q_reg ( .D(g22105), .SI(g845), .SE(n10288), .CLK(n10475), .Q(
        g846), .QN(n10082) );
  SDFFX1 DFF_537_Q_reg ( .D(g22127), .SI(g846), .SE(n10288), .CLK(n10475), .Q(
        g844), .QN(n9722) );
  SDFFX1 DFF_538_Q_reg ( .D(g22106), .SI(g844), .SE(n10289), .CLK(n10476), .Q(
        g848), .QN(n9721) );
  SDFFX1 DFF_539_Q_reg ( .D(g22128), .SI(g848), .SE(n10289), .CLK(n10476), .Q(
        g849), .QN(n9720) );
  SDFFX1 DFF_540_Q_reg ( .D(g22147), .SI(g849), .SE(n10289), .CLK(n10476), .Q(
        g847), .QN(n9719) );
  SDFFX1 DFF_541_Q_reg ( .D(g22129), .SI(g847), .SE(n10289), .CLK(n10476), .Q(
        g851), .QN(n9718) );
  SDFFX1 DFF_542_Q_reg ( .D(g22148), .SI(g851), .SE(n10289), .CLK(n10476), .Q(
        g852), .QN(n9717) );
  SDFFX1 DFF_543_Q_reg ( .D(g22164), .SI(g852), .SE(n10289), .CLK(n10476), .Q(
        g850), .QN(n9716) );
  SDFFX1 DFF_544_Q_reg ( .D(g25209), .SI(g850), .SE(n10289), .CLK(n10476), .Q(
        g857), .QN(n9788) );
  SDFFX1 DFF_545_Q_reg ( .D(g25214), .SI(g857), .SE(n10289), .CLK(n10476), .Q(
        test_so33), .QN(n10206) );
  SDFFX1 DFF_546_Q_reg ( .D(g25221), .SI(test_si34), .SE(n10285), .CLK(n10472), 
        .Q(g856), .QN(n9787) );
  SDFFX1 DFF_547_Q_reg ( .D(g25215), .SI(g856), .SE(n10285), .CLK(n10472), .Q(
        g860), .QN(n9786) );
  SDFFX1 DFF_548_Q_reg ( .D(g25222), .SI(g860), .SE(n10285), .CLK(n10472), .Q(
        g861), .QN(n9785) );
  SDFFX1 DFF_549_Q_reg ( .D(g25230), .SI(g861), .SE(n10285), .CLK(n10472), .Q(
        g859), .QN(n9784) );
  SDFFX1 DFF_550_Q_reg ( .D(g25223), .SI(g859), .SE(n10285), .CLK(n10472), .Q(
        g863), .QN(n9783) );
  SDFFX1 DFF_551_Q_reg ( .D(g25231), .SI(g863), .SE(n10285), .CLK(n10472), .Q(
        g864), .QN(n9782) );
  SDFFX1 DFF_552_Q_reg ( .D(g25240), .SI(g864), .SE(n10285), .CLK(n10472), .Q(
        g862), .QN(n9781) );
  SDFFX1 DFF_553_Q_reg ( .D(g25232), .SI(g862), .SE(n10285), .CLK(n10472), .Q(
        g866) );
  SDFFX1 DFF_554_Q_reg ( .D(g25241), .SI(g866), .SE(n10286), .CLK(n10473), .Q(
        g867) );
  SDFFX1 DFF_555_Q_reg ( .D(g25248), .SI(g867), .SE(n10286), .CLK(n10473), .Q(
        g865) );
  SDFFX1 DFF_556_Q_reg ( .D(g30269), .SI(g865), .SE(n10295), .CLK(n10482), .Q(
        g873) );
  SDFFX1 DFF_557_Q_reg ( .D(g30277), .SI(g873), .SE(n10295), .CLK(n10482), .Q(
        g876) );
  SDFFX1 DFF_558_Q_reg ( .D(g30285), .SI(g876), .SE(n10295), .CLK(n10482), .Q(
        g879) );
  SDFFX1 DFF_559_Q_reg ( .D(g30643), .SI(g879), .SE(n10295), .CLK(n10482), .Q(
        g918) );
  SDFFX1 DFF_560_Q_reg ( .D(g30648), .SI(g918), .SE(n10295), .CLK(n10482), .Q(
        g921) );
  SDFFX1 DFF_561_Q_reg ( .D(g30654), .SI(g921), .SE(n10296), .CLK(n10483), .Q(
        test_so34) );
  SDFFX1 DFF_562_Q_reg ( .D(g30676), .SI(test_si35), .SE(n10290), .CLK(n10477), 
        .Q(g882) );
  SDFFX1 DFF_563_Q_reg ( .D(g30681), .SI(g882), .SE(n10291), .CLK(n10478), .Q(
        g885) );
  SDFFX1 DFF_564_Q_reg ( .D(g30687), .SI(g885), .SE(n10291), .CLK(n10478), .Q(
        g888) );
  SDFFX1 DFF_565_Q_reg ( .D(g30649), .SI(g888), .SE(n10291), .CLK(n10478), .Q(
        g927) );
  SDFFX1 DFF_566_Q_reg ( .D(g30655), .SI(g927), .SE(n10291), .CLK(n10478), .Q(
        g930) );
  SDFFX1 DFF_567_Q_reg ( .D(g30662), .SI(g930), .SE(n10290), .CLK(n10477), .Q(
        g933) );
  SDFFX1 DFF_568_Q_reg ( .D(g30286), .SI(g933), .SE(n10291), .CLK(n10478), .Q(
        g891) );
  SDFFX1 DFF_569_Q_reg ( .D(g30293), .SI(g891), .SE(n10291), .CLK(n10478), .Q(
        g894) );
  SDFFX1 DFF_570_Q_reg ( .D(g30298), .SI(g894), .SE(n10291), .CLK(n10478), .Q(
        g897) );
  SDFFX1 DFF_571_Q_reg ( .D(g30259), .SI(g897), .SE(n10291), .CLK(n10478), .Q(
        g936) );
  SDFFX1 DFF_572_Q_reg ( .D(g30264), .SI(g936), .SE(n10291), .CLK(n10478), .Q(
        g939) );
  SDFFX1 DFF_573_Q_reg ( .D(g30270), .SI(g939), .SE(n10291), .CLK(n10478), .Q(
        g942) );
  SDFFX1 DFF_574_Q_reg ( .D(g30247), .SI(g942), .SE(n10291), .CLK(n10478), .Q(
        g900) );
  SDFFX1 DFF_575_Q_reg ( .D(g30249), .SI(g900), .SE(n10291), .CLK(n10478), .Q(
        g903) );
  SDFFX1 DFF_576_Q_reg ( .D(g30251), .SI(g903), .SE(n10292), .CLK(n10479), .Q(
        g906) );
  SDFFX1 DFF_577_Q_reg ( .D(g30265), .SI(g906), .SE(n10292), .CLK(n10479), .Q(
        test_so35) );
  SDFFX1 DFF_578_Q_reg ( .D(g30271), .SI(test_si36), .SE(n10292), .CLK(n10479), 
        .Q(g948) );
  SDFFX1 DFF_579_Q_reg ( .D(g30278), .SI(g948), .SE(n10292), .CLK(n10479), .Q(
        g951) );
  SDFFX1 DFF_580_Q_reg ( .D(g30638), .SI(g951), .SE(n10292), .CLK(n10479), .Q(
        g909) );
  SDFFX1 DFF_581_Q_reg ( .D(g30642), .SI(g909), .SE(n10292), .CLK(n10479), .Q(
        g912) );
  SDFFX1 DFF_582_Q_reg ( .D(g30647), .SI(g912), .SE(n10292), .CLK(n10479), .Q(
        g915) );
  SDFFX1 DFF_583_Q_reg ( .D(g30670), .SI(g915), .SE(n10292), .CLK(n10479), .Q(
        g954) );
  SDFFX1 DFF_584_Q_reg ( .D(g30677), .SI(g954), .SE(n10292), .CLK(n10479), .Q(
        g957) );
  SDFFX1 DFF_585_Q_reg ( .D(g30682), .SI(g957), .SE(n10286), .CLK(n10473), .Q(
        g960) );
  SDFFX1 DFF_586_Q_reg ( .D(g25042), .SI(g960), .SE(n10286), .CLK(n10473), .Q(
        g780), .QN(n9887) );
  SDFFX1 DFF_587_Q_reg ( .D(g25935), .SI(g780), .SE(n10286), .CLK(n10473), .Q(
        g776), .QN(n10172) );
  SDFFX1 DFF_588_Q_reg ( .D(g26530), .SI(g776), .SE(n10286), .CLK(n10473), .Q(
        g771), .QN(n9886) );
  SDFFX1 DFF_589_Q_reg ( .D(g27123), .SI(g771), .SE(n10286), .CLK(n10473), .Q(
        g767), .QN(n10171) );
  SDFFX1 DFF_590_Q_reg ( .D(g27603), .SI(g767), .SE(n10286), .CLK(n10473), .Q(
        g762), .QN(n9885) );
  SDFFX1 DFF_591_Q_reg ( .D(g28146), .SI(g762), .SE(n10287), .CLK(n10474), .Q(
        g758), .QN(n10170) );
  SDFFX1 DFF_592_Q_reg ( .D(g28635), .SI(g758), .SE(n10287), .CLK(n10474), .Q(
        g753), .QN(n9884) );
  SDFFX1 DFF_593_Q_reg ( .D(g29110), .SI(g753), .SE(n10287), .CLK(n10474), .Q(
        test_so36), .QN(n10195) );
  SDFFX1 DFF_594_Q_reg ( .D(g29354), .SI(test_si37), .SE(n10287), .CLK(n10474), 
        .Q(g744), .QN(n9509) );
  SDFFX1 DFF_595_Q_reg ( .D(g29580), .SI(g744), .SE(n10287), .CLK(n10474), .Q(
        g740), .QN(n9355) );
  SDFFX1 DFF_596_Q_reg ( .D(n29), .SI(g740), .SE(n10287), .CLK(n10474), .Q(
        g868) );
  SDFFX1 DFF_597_Q_reg ( .D(g868), .SI(g868), .SE(n10287), .CLK(n10474), .Q(
        g5595) );
  SDFFX1 DFF_598_Q_reg ( .D(g5595), .SI(g5595), .SE(n10287), .CLK(n10474), .Q(
        g869), .QN(n10160) );
  SDFFX1 DFF_599_Q_reg ( .D(g2950), .SI(g869), .SE(n10287), .CLK(n10474), .Q(
        g5472), .QN(n4363) );
  SDFFX1 DFF_600_Q_reg ( .D(g5472), .SI(g5472), .SE(n10287), .CLK(n10474), .Q(
        g6712), .QN(n4364) );
  SDFFX1 DFF_601_Q_reg ( .D(g6712), .SI(g6712), .SE(n10287), .CLK(n10474), .Q(
        g1088), .QN(n4381) );
  SDFFX1 DFF_602_Q_reg ( .D(g5595), .SI(g1088), .SE(n10287), .CLK(n10474), .Q(
        g996), .QN(n4387) );
  SDFFX1 DFF_603_Q_reg ( .D(g27257), .SI(g996), .SE(n10295), .CLK(n10482), .Q(
        g1041), .QN(n9840) );
  SDFFX1 DFF_604_Q_reg ( .D(g27262), .SI(g1041), .SE(n10295), .CLK(n10482), 
        .Q(g1030), .QN(n9839) );
  SDFFX1 DFF_605_Q_reg ( .D(g27270), .SI(g1030), .SE(n10295), .CLK(n10482), 
        .Q(g1033), .QN(n9838) );
  SDFFX1 DFF_606_Q_reg ( .D(g27263), .SI(g1033), .SE(n10295), .CLK(n10482), 
        .Q(g1056), .QN(n9817) );
  SDFFX1 DFF_607_Q_reg ( .D(g27271), .SI(g1056), .SE(n10295), .CLK(n10482), 
        .Q(g1045), .QN(n9816) );
  SDFFX1 DFF_608_Q_reg ( .D(g27282), .SI(g1045), .SE(n10294), .CLK(n10481), 
        .Q(g1048), .QN(n9815) );
  SDFFX1 DFF_609_Q_reg ( .D(g27272), .SI(g1048), .SE(n10294), .CLK(n10481), 
        .Q(test_so37), .QN(n10203) );
  SDFFX1 DFF_610_Q_reg ( .D(g27283), .SI(test_si38), .SE(n10294), .CLK(n10481), 
        .Q(g1060), .QN(n9562) );
  SDFFX1 DFF_611_Q_reg ( .D(g27297), .SI(g1060), .SE(n10294), .CLK(n10481), 
        .Q(g1063), .QN(n9563) );
  SDFFX1 DFF_612_Q_reg ( .D(g27284), .SI(g1063), .SE(n10295), .CLK(n10482), 
        .Q(g1085), .QN(n9828) );
  SDFFX1 DFF_613_Q_reg ( .D(g27298), .SI(g1085), .SE(n10295), .CLK(n10482), 
        .Q(g1075), .QN(n9827) );
  SDFFX1 DFF_614_Q_reg ( .D(g27313), .SI(g1075), .SE(n10292), .CLK(n10479), 
        .Q(g1078), .QN(n9826) );
  SDFFX1 DFF_615_Q_reg ( .D(g28738), .SI(g1078), .SE(n10292), .CLK(n10479), 
        .Q(g1095) );
  SDFFX1 DFF_616_Q_reg ( .D(g28746), .SI(g1095), .SE(n10294), .CLK(n10481), 
        .Q(g1098) );
  SDFFX1 DFF_617_Q_reg ( .D(g28758), .SI(g1098), .SE(n10294), .CLK(n10481), 
        .Q(g1101) );
  SDFFX1 DFF_618_Q_reg ( .D(g29198), .SI(g1101), .SE(n10294), .CLK(n10481), 
        .Q(g1104) );
  SDFFX1 DFF_619_Q_reg ( .D(g29204), .SI(g1104), .SE(n10294), .CLK(n10481), 
        .Q(g1107) );
  SDFFX1 DFF_620_Q_reg ( .D(g29209), .SI(g1107), .SE(n10293), .CLK(n10480), 
        .Q(g1110) );
  SDFFX1 DFF_621_Q_reg ( .D(g28747), .SI(g1110), .SE(n10293), .CLK(n10480), 
        .Q(g1114), .QN(n9866) );
  SDFFX1 DFF_622_Q_reg ( .D(g28759), .SI(g1114), .SE(n10293), .CLK(n10480), 
        .Q(g1115), .QN(n9851) );
  SDFFX1 DFF_623_Q_reg ( .D(g28767), .SI(g1115), .SE(n10293), .CLK(n10480), 
        .Q(g1113), .QN(n9865) );
  SDFFX1 DFF_624_Q_reg ( .D(g26806), .SI(g1113), .SE(n10293), .CLK(n10480), 
        .Q(g1116) );
  SDFFX1 DFF_625_Q_reg ( .D(g26809), .SI(g1116), .SE(n10293), .CLK(n10480), 
        .Q(test_so38) );
  SDFFX1 DFF_626_Q_reg ( .D(g26813), .SI(test_si39), .SE(n10293), .CLK(n10480), 
        .Q(g1122) );
  SDFFX1 DFF_627_Q_reg ( .D(g26810), .SI(g1122), .SE(n10293), .CLK(n10480), 
        .Q(g1125) );
  SDFFX1 DFF_628_Q_reg ( .D(g26814), .SI(g1125), .SE(n10293), .CLK(n10480), 
        .Q(g1128) );
  SDFFX1 DFF_629_Q_reg ( .D(g26818), .SI(g1128), .SE(n10294), .CLK(n10481), 
        .Q(g1131) );
  SDFFX1 DFF_630_Q_reg ( .D(g27761), .SI(g1131), .SE(n10294), .CLK(n10481), 
        .Q(g1135), .QN(n9864) );
  SDFFX1 DFF_631_Q_reg ( .D(g27763), .SI(g1135), .SE(n10294), .CLK(n10481), 
        .Q(g1136), .QN(n9850) );
  SDFFX1 DFF_632_Q_reg ( .D(g27765), .SI(g1136), .SE(n10293), .CLK(n10480), 
        .Q(g1134), .QN(n9863) );
  SDFFX1 DFF_633_Q_reg ( .D(g29609), .SI(g1134), .SE(n10293), .CLK(n10480), 
        .Q(g999), .QN(n9469) );
  SDFFX1 DFF_634_Q_reg ( .D(g29612), .SI(g999), .SE(n10293), .CLK(n10480), .Q(
        g1000), .QN(n9452) );
  SDFFX1 DFF_635_Q_reg ( .D(g29616), .SI(g1000), .SE(n10292), .CLK(n10479), 
        .Q(g1001), .QN(n9468) );
  SDFFX1 DFF_636_Q_reg ( .D(g30701), .SI(g1001), .SE(n10286), .CLK(n10473), 
        .Q(g1002), .QN(n9467) );
  SDFFX1 DFF_637_Q_reg ( .D(g30703), .SI(g1002), .SE(n10288), .CLK(n10475), 
        .Q(g1003), .QN(n9451) );
  SDFFX1 DFF_638_Q_reg ( .D(g30705), .SI(g1003), .SE(n10288), .CLK(n10475), 
        .Q(g1004), .QN(n9466) );
  SDFFX1 DFF_639_Q_reg ( .D(g30470), .SI(g1004), .SE(n10286), .CLK(n10473), 
        .Q(g1005), .QN(n9465) );
  SDFFX1 DFF_640_Q_reg ( .D(g30485), .SI(g1005), .SE(n10288), .CLK(n10475), 
        .Q(g1006), .QN(n9450) );
  SDFFX1 DFF_641_Q_reg ( .D(g30500), .SI(g1006), .SE(n10288), .CLK(n10475), 
        .Q(test_so39) );
  SDFFX1 DFF_642_Q_reg ( .D(g29170), .SI(test_si40), .SE(n10296), .CLK(n10483), 
        .Q(g1009) );
  SDFFX1 DFF_643_Q_reg ( .D(g29173), .SI(g1009), .SE(n10296), .CLK(n10483), 
        .Q(g1010) );
  SDFFX1 DFF_644_Q_reg ( .D(g29179), .SI(g1010), .SE(n10296), .CLK(n10483), 
        .Q(g1008) );
  SDFFX1 DFF_645_Q_reg ( .D(g26661), .SI(g1008), .SE(n10296), .CLK(n10483), 
        .Q(g1090), .QN(n9862) );
  SDFFX1 DFF_646_Q_reg ( .D(g26665), .SI(g1090), .SE(n10296), .CLK(n10483), 
        .Q(g1091), .QN(n9849) );
  SDFFX1 DFF_647_Q_reg ( .D(g26669), .SI(g1091), .SE(n10296), .CLK(n10483), 
        .Q(g1089), .QN(n9861) );
  SDFFX1 DFF_648_Q_reg ( .D(n4289), .SI(g1089), .SE(n10296), .CLK(n10483), .Q(
        g1137) );
  SDFFX1 DFF_649_Q_reg ( .D(g1137), .SI(g1137), .SE(n10296), .CLK(n10483), .Q(
        n8027), .QN(DFF_649_n1) );
  SDFFX1 DFF_650_Q_reg ( .D(n4567), .SI(n8027), .SE(n10296), .CLK(n10483), .Q(
        g1139) );
  SDFFX1 DFF_651_Q_reg ( .D(g1139), .SI(g1139), .SE(n10296), .CLK(n10483), .Q(
        n8026), .QN(DFF_651_n1) );
  SDFFX1 DFF_652_Q_reg ( .D(n4559), .SI(n8026), .SE(n10296), .CLK(n10483), .Q(
        g1141) );
  SDFFX1 DFF_653_Q_reg ( .D(g1141), .SI(g1141), .SE(n10297), .CLK(n10484), .Q(
        n8025), .QN(DFF_653_n1) );
  SDFFX1 DFF_654_Q_reg ( .D(n4327), .SI(n8025), .SE(n10297), .CLK(n10484), .Q(
        g967) );
  SDFFX1 DFF_655_Q_reg ( .D(g967), .SI(g967), .SE(n10297), .CLK(n10484), .Q(
        n8024), .QN(DFF_655_n1) );
  SDFFX1 DFF_656_Q_reg ( .D(n4391), .SI(n8024), .SE(n10297), .CLK(n10484), .Q(
        g969) );
  SDFFX1 DFF_657_Q_reg ( .D(g969), .SI(g969), .SE(n10297), .CLK(n10484), .Q(
        test_so40), .QN(DFF_657_n1) );
  SDFFX1 DFF_658_Q_reg ( .D(n4321), .SI(test_si41), .SE(n10239), .CLK(n10426), 
        .Q(g971) );
  SDFFX1 DFF_659_Q_reg ( .D(g971), .SI(g971), .SE(n10240), .CLK(n10427), .Q(
        n8021), .QN(DFF_659_n1) );
  SDFFX1 DFF_660_Q_reg ( .D(n4375), .SI(n8021), .SE(n10240), .CLK(n10427), .Q(
        g973) );
  SDFFX1 DFF_661_Q_reg ( .D(g973), .SI(g973), .SE(n10240), .CLK(n10427), .Q(
        n8020), .QN(DFF_661_n1) );
  SDFFX1 DFF_662_Q_reg ( .D(n4379), .SI(n8020), .SE(n10240), .CLK(n10427), .Q(
        g975) );
  SDFFX1 DFF_663_Q_reg ( .D(g975), .SI(g975), .SE(n10240), .CLK(n10427), .Q(
        n8019), .QN(DFF_663_n1) );
  SDFFX1 DFF_664_Q_reg ( .D(g2873), .SI(n8019), .SE(n10240), .CLK(n10427), .Q(
        g977) );
  SDFFX1 DFF_665_Q_reg ( .D(g977), .SI(g977), .SE(n10240), .CLK(n10427), .Q(
        n8018), .QN(n4486) );
  SDFFX1 DFF_666_Q_reg ( .D(n4283), .SI(n8018), .SE(n10294), .CLK(n10481), .Q(
        g986), .QN(n4432) );
  SDFFX1 DFF_667_Q_reg ( .D(n534), .SI(g986), .SE(n10297), .CLK(n10484), .Q(
        g992), .QN(n9894) );
  SDFFX1 DFF_678_Q_reg ( .D(n4277), .SI(g992), .SE(n10297), .CLK(n10484), .Q(
        n8017) );
  SDFFX1 DFF_679_Q_reg ( .D(g1041), .SI(n8017), .SE(n10297), .CLK(n10484), .Q(
        g1029) );
  SDFFX1 DFF_680_Q_reg ( .D(g1029), .SI(g1029), .SE(n10297), .CLK(n10484), .Q(
        g1036) );
  SDFFX1 DFF_681_Q_reg ( .D(g1030), .SI(g1036), .SE(n10297), .CLK(n10484), .Q(
        g1037) );
  SDFFX1 DFF_682_Q_reg ( .D(g1037), .SI(g1037), .SE(n10297), .CLK(n10484), .Q(
        g1038) );
  SDFFX1 DFF_683_Q_reg ( .D(g1033), .SI(g1038), .SE(n10297), .CLK(n10484), .Q(
        test_so41) );
  SDFFX1 DFF_684_Q_reg ( .D(test_so41), .SI(test_si42), .SE(n10298), .CLK(
        n10485), .Q(g1040) );
  SDFFX1 DFF_685_Q_reg ( .D(g1056), .SI(g1040), .SE(n10298), .CLK(n10485), .Q(
        g1044) );
  SDFFX1 DFF_686_Q_reg ( .D(g1044), .SI(g1044), .SE(n10298), .CLK(n10485), .Q(
        g1051) );
  SDFFX1 DFF_687_Q_reg ( .D(g1045), .SI(g1051), .SE(n10298), .CLK(n10485), .Q(
        g1052) );
  SDFFX1 DFF_688_Q_reg ( .D(g1052), .SI(g1052), .SE(n10298), .CLK(n10485), .Q(
        g1053) );
  SDFFX1 DFF_689_Q_reg ( .D(g1048), .SI(g1053), .SE(n10298), .CLK(n10485), .Q(
        g1054) );
  SDFFX1 DFF_690_Q_reg ( .D(g1054), .SI(g1054), .SE(n10298), .CLK(n10485), .Q(
        g1055) );
  SDFFX1 DFF_691_Q_reg ( .D(test_so37), .SI(g1055), .SE(n10298), .CLK(n10485), 
        .Q(g1059) );
  SDFFX1 DFF_692_Q_reg ( .D(g1059), .SI(g1059), .SE(n10298), .CLK(n10485), .Q(
        g1066) );
  SDFFX1 DFF_693_Q_reg ( .D(g1060), .SI(g1066), .SE(n10298), .CLK(n10485), .Q(
        g1067) );
  SDFFX1 DFF_694_Q_reg ( .D(g1067), .SI(g1067), .SE(n10298), .CLK(n10485), .Q(
        g1068) );
  SDFFX1 DFF_695_Q_reg ( .D(g1063), .SI(g1068), .SE(n10298), .CLK(n10485), .Q(
        g1069) );
  SDFFX1 DFF_696_Q_reg ( .D(g1069), .SI(g1069), .SE(n10299), .CLK(n10486), .Q(
        g1070) );
  SDFFX1 DFF_697_Q_reg ( .D(g1085), .SI(g1070), .SE(n10299), .CLK(n10486), .Q(
        g1074) );
  SDFFX1 DFF_698_Q_reg ( .D(g1074), .SI(g1074), .SE(n10299), .CLK(n10486), .Q(
        g1081) );
  SDFFX1 DFF_699_Q_reg ( .D(g1075), .SI(g1081), .SE(n10299), .CLK(n10486), .Q(
        test_so42) );
  SDFFX1 DFF_700_Q_reg ( .D(test_so42), .SI(test_si43), .SE(n10299), .CLK(
        n10486), .Q(g1083) );
  SDFFX1 DFF_701_Q_reg ( .D(g1078), .SI(g1083), .SE(n10299), .CLK(n10486), .Q(
        g1084) );
  SDFFX1 DFF_702_Q_reg ( .D(g1084), .SI(g1084), .SE(n10299), .CLK(n10486), .Q(
        g1011) );
  SDFFX1 DFF_703_Q_reg ( .D(n4598), .SI(g1011), .SE(n10299), .CLK(n10486), .Q(
        g5657) );
  SDFFX1 DFF_704_Q_reg ( .D(g5657), .SI(g5657), .SE(n10299), .CLK(n10486), .Q(
        g5686) );
  SDFFX1 DFF_705_Q_reg ( .D(g5686), .SI(g5686), .SE(n10299), .CLK(n10486), .Q(
        g1024) );
  SDFFX1 DFF_706_Q_reg ( .D(n4598), .SI(g1024), .SE(n10299), .CLK(n10486), .Q(
        g6750), .QN(n4371) );
  SDFFX1 DFF_707_Q_reg ( .D(g6750), .SI(g6750), .SE(n10299), .CLK(n10486), .Q(
        g6944), .QN(n4316) );
  SDFFX1 DFF_708_Q_reg ( .D(g6944), .SI(g6944), .SE(n10300), .CLK(n10487), .Q(
        g1236), .QN(n4300) );
  SDFFX1 DFF_709_Q_reg ( .D(g21843), .SI(g1236), .SE(n10300), .CLK(n10487), 
        .Q(g1240), .QN(n10122) );
  SDFFX1 DFF_710_Q_reg ( .D(g18707), .SI(g1240), .SE(n10300), .CLK(n10487), 
        .Q(g1243), .QN(n4353) );
  SDFFX1 DFF_711_Q_reg ( .D(g18763), .SI(g1243), .SE(n10300), .CLK(n10487), 
        .Q(g1196), .QN(n4304) );
  SDFFX1 DFF_712_Q_reg ( .D(n962), .SI(g1196), .SE(n10301), .CLK(n10488), .Q(
        g1199) );
  SDFFX1 DFF_713_Q_reg ( .D(g1199), .SI(g1199), .SE(n10301), .CLK(n10488), .Q(
        g1209) );
  SDFFX1 DFF_714_Q_reg ( .D(g1209), .SI(g1209), .SE(n10301), .CLK(n10488), .Q(
        g1210) );
  SDFFX1 DFF_715_Q_reg ( .D(g1142), .SI(g1210), .SE(n10301), .CLK(n10488), .Q(
        test_so43) );
  SDFFX1 DFF_716_Q_reg ( .D(test_so43), .SI(test_si44), .SE(n10301), .CLK(
        n10488), .Q(g1255) );
  SDFFX1 DFF_717_Q_reg ( .D(g1145), .SI(g1255), .SE(n10301), .CLK(n10488), .Q(
        g1256) );
  SDFFX1 DFF_718_Q_reg ( .D(g1256), .SI(g1256), .SE(n10301), .CLK(n10488), .Q(
        g1257) );
  SDFFX1 DFF_719_Q_reg ( .D(g1148), .SI(g1257), .SE(n10301), .CLK(n10488), .Q(
        g1258) );
  SDFFX1 DFF_720_Q_reg ( .D(g1258), .SI(g1258), .SE(n10302), .CLK(n10489), .Q(
        g1259) );
  SDFFX1 DFF_721_Q_reg ( .D(g1152), .SI(g1259), .SE(n10302), .CLK(n10489), .Q(
        g1260) );
  SDFFX1 DFF_722_Q_reg ( .D(g1260), .SI(g1260), .SE(n10302), .CLK(n10489), .Q(
        g1251) );
  SDFFX1 DFF_723_Q_reg ( .D(g1155), .SI(g1251), .SE(n10302), .CLK(n10489), .Q(
        g1252) );
  SDFFX1 DFF_724_Q_reg ( .D(g1252), .SI(g1252), .SE(n10302), .CLK(n10489), .Q(
        g1253) );
  SDFFX1 DFF_725_Q_reg ( .D(g1158), .SI(g1253), .SE(n10302), .CLK(n10489), .Q(
        g1254) );
  SDFFX1 DFF_726_Q_reg ( .D(g1254), .SI(g1254), .SE(n10302), .CLK(n10489), .Q(
        g1176) );
  SDFFX1 DFF_727_Q_reg ( .D(g2950), .SI(g1176), .SE(n10302), .CLK(n10489), .Q(
        g7961), .QN(n4460) );
  SDFFX1 DFF_728_Q_reg ( .D(g7961), .SI(g7961), .SE(n10302), .CLK(n10489), .Q(
        g8007), .QN(n4459) );
  SDFFX1 DFF_729_Q_reg ( .D(g8007), .SI(g8007), .SE(n10302), .CLK(n10489), .Q(
        g1172), .QN(n4465) );
  SDFFX1 DFF_730_Q_reg ( .D(g23081), .SI(g1172), .SE(n10304), .CLK(n10491), 
        .Q(g1173) );
  SDFFX1 DFF_731_Q_reg ( .D(g23111), .SI(g1173), .SE(n10304), .CLK(n10491), 
        .Q(test_so44) );
  SDFFX1 DFF_732_Q_reg ( .D(g23126), .SI(test_si45), .SE(n10302), .CLK(n10489), 
        .Q(g1175) );
  SDFFX1 DFF_733_Q_reg ( .D(g23392), .SI(g1175), .SE(n10302), .CLK(n10489), 
        .Q(g1142) );
  SDFFX1 DFF_734_Q_reg ( .D(g23406), .SI(g1142), .SE(n10303), .CLK(n10490), 
        .Q(g1145) );
  SDFFX1 DFF_735_Q_reg ( .D(g24179), .SI(g1145), .SE(n10303), .CLK(n10490), 
        .Q(g1148) );
  SDFFX1 DFF_736_Q_reg ( .D(g24181), .SI(g1148), .SE(n10303), .CLK(n10490), 
        .Q(g1164) );
  SDFFX1 DFF_737_Q_reg ( .D(g24213), .SI(g1164), .SE(n10303), .CLK(n10490), 
        .Q(g1165) );
  SDFFX1 DFF_738_Q_reg ( .D(g24223), .SI(g1165), .SE(n10303), .CLK(n10490), 
        .Q(g1166) );
  SDFFX1 DFF_739_Q_reg ( .D(g23110), .SI(g1166), .SE(n10303), .CLK(n10490), 
        .Q(g1167) );
  SDFFX1 DFF_740_Q_reg ( .D(g23014), .SI(g1167), .SE(n10303), .CLK(n10490), 
        .Q(g1171) );
  SDFFX1 DFF_741_Q_reg ( .D(g23039), .SI(g1171), .SE(n10303), .CLK(n10490), 
        .Q(g1151) );
  SDFFX1 DFF_742_Q_reg ( .D(g24212), .SI(g1151), .SE(n10303), .CLK(n10490), 
        .Q(g1152) );
  SDFFX1 DFF_743_Q_reg ( .D(g24222), .SI(g1152), .SE(n10303), .CLK(n10490), 
        .Q(g1155) );
  SDFFX1 DFF_744_Q_reg ( .D(g24235), .SI(g1155), .SE(n10303), .CLK(n10490), 
        .Q(g1158) );
  SDFFX1 DFF_745_Q_reg ( .D(n984), .SI(g1158), .SE(n10303), .CLK(n10490), .Q(
        g1214) );
  SDFFX1 DFF_746_Q_reg ( .D(g1214), .SI(g1214), .SE(n10304), .CLK(n10491), .Q(
        g1221) );
  SDFFX1 DFF_747_Q_reg ( .D(g1221), .SI(g1221), .SE(n10304), .CLK(n10491), .Q(
        test_so45) );
  SDFFX1 DFF_748_Q_reg ( .D(g13155), .SI(test_si46), .SE(n10304), .CLK(n10491), 
        .Q(g1229) );
  SDFFX1 DFF_749_Q_reg ( .D(g1229), .SI(g1229), .SE(n10304), .CLK(n10491), .Q(
        n4549), .QN(n9338) );
  SDFFX1 DFF_750_Q_reg ( .D(n578), .SI(n4549), .SE(n10304), .CLK(n10491), .Q(
        n4361), .QN(n9339) );
  SDFFX1 DFF_751_Q_reg ( .D(g13124), .SI(n4361), .SE(n10304), .CLK(n10491), 
        .Q(g1235) );
  SDFFX1 DFF_752_Q_reg ( .D(g1235), .SI(g1235), .SE(n10304), .CLK(n10491), .Q(
        g1186), .QN(n4548) );
  SDFFX1 DFF_753_Q_reg ( .D(g13171), .SI(g1186), .SE(n10304), .CLK(n10491), 
        .Q(g1244) );
  SDFFX1 DFF_754_Q_reg ( .D(g1244), .SI(g1244), .SE(n10304), .CLK(n10491), .Q(
        g1245) );
  SDFFX1 DFF_755_Q_reg ( .D(g27273), .SI(g1245), .SE(n10305), .CLK(n10492), 
        .Q(g1262), .QN(n9517) );
  SDFFX1 DFF_756_Q_reg ( .D(g27285), .SI(g1262), .SE(n10305), .CLK(n10492), 
        .Q(g1263), .QN(n9519) );
  SDFFX1 DFF_757_Q_reg ( .D(g27299), .SI(g1263), .SE(n10305), .CLK(n10492), 
        .Q(g1261), .QN(n9518) );
  SDFFX1 DFF_758_Q_reg ( .D(g27286), .SI(g1261), .SE(n10305), .CLK(n10492), 
        .Q(g1265), .QN(n9529) );
  SDFFX1 DFF_759_Q_reg ( .D(g27300), .SI(g1265), .SE(n10305), .CLK(n10492), 
        .Q(g1266), .QN(n9531) );
  SDFFX1 DFF_760_Q_reg ( .D(g27314), .SI(g1266), .SE(n10305), .CLK(n10492), 
        .Q(g1264), .QN(n9530) );
  SDFFX1 DFF_761_Q_reg ( .D(g27301), .SI(g1264), .SE(n10305), .CLK(n10492), 
        .Q(g1268), .QN(n9362) );
  SDFFX1 DFF_762_Q_reg ( .D(g27315), .SI(g1268), .SE(n10305), .CLK(n10492), 
        .Q(g1269), .QN(n9363) );
  SDFFX1 DFF_763_Q_reg ( .D(g27328), .SI(g1269), .SE(n10305), .CLK(n10492), 
        .Q(test_so46), .QN(n10207) );
  SDFFX1 DFF_764_Q_reg ( .D(g27316), .SI(test_si47), .SE(n10305), .CLK(n10492), 
        .Q(g1271), .QN(n9539) );
  SDFFX1 DFF_765_Q_reg ( .D(g27329), .SI(g1271), .SE(n10305), .CLK(n10492), 
        .Q(g1272), .QN(n9541) );
  SDFFX1 DFF_766_Q_reg ( .D(g27339), .SI(g1272), .SE(n10305), .CLK(n10492), 
        .Q(g1270), .QN(n9540) );
  SDFFX1 DFF_767_Q_reg ( .D(g24501), .SI(g1270), .SE(n10306), .CLK(n10493), 
        .Q(g1273) );
  SDFFX1 DFF_768_Q_reg ( .D(g24510), .SI(g1273), .SE(n10306), .CLK(n10493), 
        .Q(g1276) );
  SDFFX1 DFF_769_Q_reg ( .D(g24521), .SI(g1276), .SE(n10306), .CLK(n10493), 
        .Q(g1279) );
  SDFFX1 DFF_770_Q_reg ( .D(g24511), .SI(g1279), .SE(n10306), .CLK(n10493), 
        .Q(g1282) );
  SDFFX1 DFF_771_Q_reg ( .D(g24522), .SI(g1282), .SE(n10306), .CLK(n10493), 
        .Q(g1285) );
  SDFFX1 DFF_772_Q_reg ( .D(g24532), .SI(g1285), .SE(n10306), .CLK(n10493), 
        .Q(g1288) );
  SDFFX1 DFF_773_Q_reg ( .D(g28351), .SI(g1288), .SE(n10306), .CLK(n10493), 
        .Q(g1300) );
  SDFFX1 DFF_774_Q_reg ( .D(g28355), .SI(g1300), .SE(n10306), .CLK(n10493), 
        .Q(g1303) );
  SDFFX1 DFF_775_Q_reg ( .D(g28360), .SI(g1303), .SE(n10304), .CLK(n10491), 
        .Q(g1306) );
  SDFFX1 DFF_776_Q_reg ( .D(g28346), .SI(g1306), .SE(n10306), .CLK(n10493), 
        .Q(g1291) );
  SDFFX1 DFF_777_Q_reg ( .D(g28350), .SI(g1291), .SE(n10306), .CLK(n10493), 
        .Q(g1294) );
  SDFFX1 DFF_778_Q_reg ( .D(g28354), .SI(g1294), .SE(n10306), .CLK(n10493), 
        .Q(g1297) );
  SDFFX1 DFF_779_Q_reg ( .D(g26547), .SI(g1297), .SE(n10306), .CLK(n10493), 
        .Q(test_so47) );
  SDFFX1 DFF_780_Q_reg ( .D(g26557), .SI(test_si48), .SE(n10307), .CLK(n10494), 
        .Q(g1180) );
  SDFFX1 DFF_781_Q_reg ( .D(g26569), .SI(g1180), .SE(n10307), .CLK(n10494), 
        .Q(g1183) );
  SDFFX1 DFF_782_Q_reg ( .D(g1186), .SI(g1183), .SE(n10307), .CLK(n10494), .Q(
        g1192), .QN(n4454) );
  SDFFX1 DFF_783_Q_reg ( .D(g22615), .SI(g1192), .SE(n10307), .CLK(n10494), 
        .Q(n8009), .QN(DFF_783_n1) );
  SDFFX1 DFF_792_Q_reg ( .D(n632), .SI(n8009), .SE(n10307), .CLK(n10494), .Q(
        g16355), .QN(DFF_792_n1) );
  SDFFX1 DFF_793_Q_reg ( .D(g16355), .SI(g16355), .SE(n10307), .CLK(n10494), 
        .Q(g1211), .QN(n9897) );
  SDFFX1 DFF_794_Q_reg ( .D(DFF_649_n1), .SI(g1211), .SE(n10307), .CLK(n10494), 
        .Q(n8008) );
  SDFFX1 DFF_795_Q_reg ( .D(DFF_651_n1), .SI(n8008), .SE(n10307), .CLK(n10494), 
        .Q(n8007) );
  SDFFX1 DFF_796_Q_reg ( .D(DFF_653_n1), .SI(n8007), .SE(n10307), .CLK(n10494), 
        .Q(n8006) );
  SDFFX1 DFF_797_Q_reg ( .D(DFF_655_n1), .SI(n8006), .SE(n10308), .CLK(n10495), 
        .Q(n8005) );
  SDFFX1 DFF_798_Q_reg ( .D(DFF_657_n1), .SI(n8005), .SE(n10308), .CLK(n10495), 
        .Q(n8004) );
  SDFFX1 DFF_799_Q_reg ( .D(DFF_659_n1), .SI(n8004), .SE(n10308), .CLK(n10495), 
        .Q(n8003) );
  SDFFX1 DFF_800_Q_reg ( .D(DFF_661_n1), .SI(n8003), .SE(n10308), .CLK(n10495), 
        .Q(g1222) );
  SDFFX1 DFF_801_Q_reg ( .D(DFF_663_n1), .SI(g1222), .SE(n10308), .CLK(n10495), 
        .Q(g1223) );
  SDFFX1 DFF_802_Q_reg ( .D(g24072), .SI(g1223), .SE(n10308), .CLK(n10495), 
        .Q(g1224), .QN(n4489) );
  SDFFX1 DFF_803_Q_reg ( .D(n4486), .SI(g1224), .SE(n10308), .CLK(n10495), .Q(
        test_so48) );
  SDFFX1 DFF_805_Q_reg ( .D(g6979), .SI(g6979), .SE(n10224), .CLK(n10411), .Q(
        g7161), .QN(n4358) );
  SDFFX1 DFF_806_Q_reg ( .D(g7161), .SI(g7161), .SE(n10224), .CLK(n10411), .Q(
        g1315), .QN(n4294) );
  SDFFX1 DFF_807_Q_reg ( .D(g16671), .SI(g1315), .SE(n10300), .CLK(n10487), 
        .Q(g1316), .QN(n10154) );
  SDFFX1 DFF_808_Q_reg ( .D(g20333), .SI(g1316), .SE(n10300), .CLK(n10487), 
        .Q(g1345), .QN(n4428) );
  SDFFX1 DFF_809_Q_reg ( .D(g20717), .SI(g1345), .SE(n10300), .CLK(n10487), 
        .Q(g1326), .QN(n4402) );
  SDFFX1 DFF_810_Q_reg ( .D(g21969), .SI(g1326), .SE(n10300), .CLK(n10487), 
        .Q(g1319), .QN(n4476) );
  SDFFX1 DFF_811_Q_reg ( .D(g23329), .SI(g1319), .SE(n10300), .CLK(n10487), 
        .Q(g1339), .QN(n4421) );
  SDFFX1 DFF_812_Q_reg ( .D(g24430), .SI(g1339), .SE(n10300), .CLK(n10487), 
        .Q(g1332), .QN(n4412) );
  SDFFX1 DFF_813_Q_reg ( .D(g25189), .SI(g1332), .SE(n10300), .CLK(n10487), 
        .Q(g1346), .QN(n4401) );
  SDFFX1 DFF_814_Q_reg ( .D(g26666), .SI(g1346), .SE(n10300), .CLK(n10487), 
        .Q(g1358), .QN(n4411) );
  SDFFX1 DFF_815_Q_reg ( .D(g26781), .SI(g1358), .SE(n10301), .CLK(n10488), 
        .Q(g1352), .QN(n4469) );
  SDFFX1 DFF_816_Q_reg ( .D(g27678), .SI(g1352), .SE(n10301), .CLK(n10488), 
        .Q(g1365), .QN(n4475) );
  SDFFX1 DFF_817_Q_reg ( .D(g27718), .SI(g1365), .SE(n10301), .CLK(n10488), 
        .Q(g1372), .QN(n4395) );
  SDFFX1 DFF_818_Q_reg ( .D(g28321), .SI(g1372), .SE(n10301), .CLK(n10488), 
        .Q(g1378), .QN(n4417) );
  SDFFX1 DFF_819_Q_reg ( .D(g20882), .SI(g1378), .SE(n10308), .CLK(n10495), 
        .Q(test_so49), .QN(n10221) );
  SDFFX1 DFF_820_Q_reg ( .D(g20896), .SI(test_si50), .SE(n10308), .CLK(n10495), 
        .Q(g1386), .QN(n9992) );
  SDFFX1 DFF_821_Q_reg ( .D(g20910), .SI(g1386), .SE(n10308), .CLK(n10495), 
        .Q(g1384), .QN(n10038) );
  SDFFX1 DFF_822_Q_reg ( .D(g20897), .SI(g1384), .SE(n10308), .CLK(n10495), 
        .Q(g1388), .QN(n9991) );
  SDFFX1 DFF_823_Q_reg ( .D(g20911), .SI(g1388), .SE(n10308), .CLK(n10495), 
        .Q(g1389), .QN(n9990) );
  SDFFX1 DFF_824_Q_reg ( .D(g20925), .SI(g1389), .SE(n10309), .CLK(n10496), 
        .Q(g1387), .QN(n10037) );
  SDFFX1 DFF_825_Q_reg ( .D(g20912), .SI(g1387), .SE(n10309), .CLK(n10496), 
        .Q(g1391), .QN(n9989) );
  SDFFX1 DFF_826_Q_reg ( .D(g20926), .SI(g1391), .SE(n10309), .CLK(n10496), 
        .Q(g1392), .QN(n9988) );
  SDFFX1 DFF_827_Q_reg ( .D(g20949), .SI(g1392), .SE(n10309), .CLK(n10496), 
        .Q(g1390), .QN(n10036) );
  SDFFX1 DFF_828_Q_reg ( .D(g20927), .SI(g1390), .SE(n10309), .CLK(n10496), 
        .Q(g1394), .QN(n9987) );
  SDFFX1 DFF_829_Q_reg ( .D(g20950), .SI(g1394), .SE(n10309), .CLK(n10496), 
        .Q(g1395), .QN(n9986) );
  SDFFX1 DFF_830_Q_reg ( .D(g20972), .SI(g1395), .SE(n10309), .CLK(n10496), 
        .Q(g1393), .QN(n10035) );
  SDFFX1 DFF_831_Q_reg ( .D(g20951), .SI(g1393), .SE(n10309), .CLK(n10496), 
        .Q(g1397), .QN(n9985) );
  SDFFX1 DFF_832_Q_reg ( .D(g20973), .SI(g1397), .SE(n10309), .CLK(n10496), 
        .Q(g1398), .QN(n9984) );
  SDFFX1 DFF_833_Q_reg ( .D(g20993), .SI(g1398), .SE(n10309), .CLK(n10496), 
        .Q(g1396), .QN(n10034) );
  SDFFX1 DFF_834_Q_reg ( .D(g20974), .SI(g1396), .SE(n10309), .CLK(n10496), 
        .Q(g1400), .QN(n9983) );
  SDFFX1 DFF_835_Q_reg ( .D(g20994), .SI(g1400), .SE(n10309), .CLK(n10496), 
        .Q(test_so50) );
  SDFFX1 DFF_836_Q_reg ( .D(g21015), .SI(test_si51), .SE(n10310), .CLK(n10497), 
        .Q(g1399), .QN(n10033) );
  SDFFX1 DFF_837_Q_reg ( .D(g20995), .SI(g1399), .SE(n10310), .CLK(n10497), 
        .Q(g1403), .QN(n9982) );
  SDFFX1 DFF_838_Q_reg ( .D(g21016), .SI(g1403), .SE(n10310), .CLK(n10497), 
        .Q(g1404), .QN(n9981) );
  SDFFX1 DFF_839_Q_reg ( .D(g21033), .SI(g1404), .SE(n10310), .CLK(n10497), 
        .Q(g1402), .QN(n10032) );
  SDFFX1 DFF_840_Q_reg ( .D(g21017), .SI(g1402), .SE(n10310), .CLK(n10497), 
        .Q(g1406), .QN(n9980) );
  SDFFX1 DFF_841_Q_reg ( .D(g21034), .SI(g1406), .SE(n10310), .CLK(n10497), 
        .Q(g1407), .QN(n9979) );
  SDFFX1 DFF_842_Q_reg ( .D(g21052), .SI(g1407), .SE(n10310), .CLK(n10497), 
        .Q(g1405), .QN(n10031) );
  SDFFX1 DFF_843_Q_reg ( .D(g21035), .SI(g1405), .SE(n10310), .CLK(n10497), 
        .Q(g1409), .QN(n9978) );
  SDFFX1 DFF_844_Q_reg ( .D(g21053), .SI(g1409), .SE(n10310), .CLK(n10497), 
        .Q(g1410), .QN(n9977) );
  SDFFX1 DFF_845_Q_reg ( .D(g21070), .SI(g1410), .SE(n10310), .CLK(n10497), 
        .Q(g1408), .QN(n10030) );
  SDFFX1 DFF_846_Q_reg ( .D(g20883), .SI(g1408), .SE(n10310), .CLK(n10497), 
        .Q(g1412), .QN(n9976) );
  SDFFX1 DFF_847_Q_reg ( .D(g20898), .SI(g1412), .SE(n10310), .CLK(n10497), 
        .Q(g1413), .QN(n9975) );
  SDFFX1 DFF_848_Q_reg ( .D(g20913), .SI(g1413), .SE(n10311), .CLK(n10498), 
        .Q(g1411), .QN(n10029) );
  SDFFX1 DFF_849_Q_reg ( .D(g20952), .SI(g1411), .SE(n10311), .CLK(n10498), 
        .Q(g1415), .QN(n9752) );
  SDFFX1 DFF_850_Q_reg ( .D(g20975), .SI(g1415), .SE(n10311), .CLK(n10498), 
        .Q(g1416), .QN(n9744) );
  SDFFX1 DFF_851_Q_reg ( .D(g20996), .SI(g1416), .SE(n10311), .CLK(n10498), 
        .Q(test_so51), .QN(n10220) );
  SDFFX1 DFF_852_Q_reg ( .D(g20976), .SI(test_si52), .SE(n10307), .CLK(n10494), 
        .Q(g1418), .QN(n9751) );
  SDFFX1 DFF_853_Q_reg ( .D(g20997), .SI(g1418), .SE(n10307), .CLK(n10494), 
        .Q(g1419), .QN(n9743) );
  SDFFX1 DFF_854_Q_reg ( .D(g21018), .SI(g1419), .SE(n10307), .CLK(n10494), 
        .Q(g1417), .QN(n9806) );
  SDFFX1 DFF_855_Q_reg ( .D(g25263), .SI(g1417), .SE(n10311), .CLK(n10498), 
        .Q(g1421) );
  SDFFX1 DFF_856_Q_reg ( .D(g25267), .SI(g1421), .SE(n10311), .CLK(n10498), 
        .Q(g1422) );
  SDFFX1 DFF_857_Q_reg ( .D(g25270), .SI(g1422), .SE(n10311), .CLK(n10498), 
        .Q(g1420) );
  SDFFX1 DFF_858_Q_reg ( .D(g22234), .SI(g1420), .SE(n10311), .CLK(n10498), 
        .Q(g1424) );
  SDFFX1 DFF_859_Q_reg ( .D(g22247), .SI(g1424), .SE(n10311), .CLK(n10498), 
        .Q(g1425) );
  SDFFX1 DFF_860_Q_reg ( .D(g22263), .SI(g1425), .SE(n10311), .CLK(n10498), 
        .Q(g1423) );
  SDFFX1 DFF_861_Q_reg ( .D(g2950), .SI(g1423), .SE(n10311), .CLK(n10498), .Q(
        g6573), .QN(n4317) );
  SDFFX1 DFF_862_Q_reg ( .D(g6573), .SI(g6573), .SE(n10312), .CLK(n10499), .Q(
        g6782), .QN(n4515) );
  SDFFX1 DFF_863_Q_reg ( .D(g6782), .SI(g6782), .SE(n10312), .CLK(n10499), .Q(
        g1547), .QN(n4368) );
  SDFFX1 DFF_864_Q_reg ( .D(g22149), .SI(g1547), .SE(n10312), .CLK(n10499), 
        .Q(g1512), .QN(n10081) );
  SDFFX1 DFF_865_Q_reg ( .D(g22166), .SI(g1512), .SE(n10315), .CLK(n10502), 
        .Q(g1513), .QN(n10080) );
  SDFFX1 DFF_866_Q_reg ( .D(g22178), .SI(g1513), .SE(n10315), .CLK(n10502), 
        .Q(g1511), .QN(n9715) );
  SDFFX1 DFF_867_Q_reg ( .D(g22167), .SI(g1511), .SE(n10312), .CLK(n10499), 
        .Q(test_so52), .QN(n10209) );
  SDFFX1 DFF_868_Q_reg ( .D(g22179), .SI(test_si53), .SE(n10316), .CLK(n10503), 
        .Q(g1516), .QN(n10079) );
  SDFFX1 DFF_869_Q_reg ( .D(g22191), .SI(g1516), .SE(n10316), .CLK(n10503), 
        .Q(g1514), .QN(n9714) );
  SDFFX1 DFF_870_Q_reg ( .D(g22035), .SI(g1514), .SE(n10316), .CLK(n10503), 
        .Q(g1524), .QN(n10078) );
  SDFFX1 DFF_871_Q_reg ( .D(g22043), .SI(g1524), .SE(n10316), .CLK(n10503), 
        .Q(g1525), .QN(n10077) );
  SDFFX1 DFF_872_Q_reg ( .D(g22057), .SI(g1525), .SE(n10316), .CLK(n10503), 
        .Q(g1523), .QN(n9713) );
  SDFFX1 DFF_873_Q_reg ( .D(g22044), .SI(g1523), .SE(n10316), .CLK(n10503), 
        .Q(g1527), .QN(n10076) );
  SDFFX1 DFF_874_Q_reg ( .D(g22058), .SI(g1527), .SE(n10316), .CLK(n10503), 
        .Q(g1528), .QN(n10075) );
  SDFFX1 DFF_875_Q_reg ( .D(g22073), .SI(g1528), .SE(n10316), .CLK(n10503), 
        .Q(g1526), .QN(n9712) );
  SDFFX1 DFF_876_Q_reg ( .D(g22059), .SI(g1526), .SE(n10316), .CLK(n10503), 
        .Q(g1530), .QN(n10074) );
  SDFFX1 DFF_877_Q_reg ( .D(g22074), .SI(g1530), .SE(n10316), .CLK(n10503), 
        .Q(g1531), .QN(n10073) );
  SDFFX1 DFF_878_Q_reg ( .D(g22090), .SI(g1531), .SE(n10316), .CLK(n10503), 
        .Q(g1529), .QN(n9711) );
  SDFFX1 DFF_879_Q_reg ( .D(g22075), .SI(g1529), .SE(n10317), .CLK(n10504), 
        .Q(g1533), .QN(n10072) );
  SDFFX1 DFF_880_Q_reg ( .D(g22091), .SI(g1533), .SE(n10317), .CLK(n10504), 
        .Q(g1534), .QN(n10071) );
  SDFFX1 DFF_881_Q_reg ( .D(g22112), .SI(g1534), .SE(n10317), .CLK(n10504), 
        .Q(g1532), .QN(n9710) );
  SDFFX1 DFF_882_Q_reg ( .D(g22092), .SI(g1532), .SE(n10317), .CLK(n10504), 
        .Q(g1536), .QN(n10070) );
  SDFFX1 DFF_883_Q_reg ( .D(g22113), .SI(g1536), .SE(n10317), .CLK(n10504), 
        .Q(test_so53), .QN(n10210) );
  SDFFX1 DFF_884_Q_reg ( .D(g22130), .SI(test_si54), .SE(n10314), .CLK(n10501), 
        .Q(g1535), .QN(n9709) );
  SDFFX1 DFF_885_Q_reg ( .D(g22114), .SI(g1535), .SE(n10314), .CLK(n10501), 
        .Q(g1539), .QN(n10069) );
  SDFFX1 DFF_886_Q_reg ( .D(g22131), .SI(g1539), .SE(n10314), .CLK(n10501), 
        .Q(g1540), .QN(n10068) );
  SDFFX1 DFF_887_Q_reg ( .D(g22150), .SI(g1540), .SE(n10314), .CLK(n10501), 
        .Q(g1538), .QN(n9708) );
  SDFFX1 DFF_888_Q_reg ( .D(g22132), .SI(g1538), .SE(n10314), .CLK(n10501), 
        .Q(g1542), .QN(n9691) );
  SDFFX1 DFF_889_Q_reg ( .D(g22151), .SI(g1542), .SE(n10315), .CLK(n10502), 
        .Q(g1543), .QN(n9690) );
  SDFFX1 DFF_890_Q_reg ( .D(g22168), .SI(g1543), .SE(n10315), .CLK(n10502), 
        .Q(g1541), .QN(n9689) );
  SDFFX1 DFF_891_Q_reg ( .D(g22152), .SI(g1541), .SE(n10316), .CLK(n10503), 
        .Q(g1545), .QN(n9707) );
  SDFFX1 DFF_892_Q_reg ( .D(g22169), .SI(g1545), .SE(n10315), .CLK(n10502), 
        .Q(g1546), .QN(n9706) );
  SDFFX1 DFF_893_Q_reg ( .D(g22180), .SI(g1546), .SE(n10315), .CLK(n10502), 
        .Q(g1544), .QN(n9705) );
  SDFFX1 DFF_894_Q_reg ( .D(g25217), .SI(g1544), .SE(n10315), .CLK(n10502), 
        .Q(g1551), .QN(n9777) );
  SDFFX1 DFF_895_Q_reg ( .D(g25224), .SI(g1551), .SE(n10315), .CLK(n10502), 
        .Q(g1552), .QN(n9776) );
  SDFFX1 DFF_896_Q_reg ( .D(g25233), .SI(g1552), .SE(n10315), .CLK(n10502), 
        .Q(g1550), .QN(n9775) );
  SDFFX1 DFF_897_Q_reg ( .D(g25225), .SI(g1550), .SE(n10315), .CLK(n10502), 
        .Q(g1554), .QN(n9774) );
  SDFFX1 DFF_898_Q_reg ( .D(g25234), .SI(g1554), .SE(n10315), .CLK(n10502), 
        .Q(g1555), .QN(n9773) );
  SDFFX1 DFF_899_Q_reg ( .D(g25242), .SI(g1555), .SE(n10315), .CLK(n10502), 
        .Q(test_so54), .QN(n10223) );
  SDFFX1 DFF_900_Q_reg ( .D(g25235), .SI(test_si55), .SE(n10311), .CLK(n10498), 
        .Q(g1557), .QN(n9772) );
  SDFFX1 DFF_901_Q_reg ( .D(g25243), .SI(g1557), .SE(n10312), .CLK(n10499), 
        .Q(g1558), .QN(n9771) );
  SDFFX1 DFF_902_Q_reg ( .D(g25249), .SI(g1558), .SE(n10312), .CLK(n10499), 
        .Q(g1556), .QN(n9770) );
  SDFFX1 DFF_903_Q_reg ( .D(g25244), .SI(g1556), .SE(n10312), .CLK(n10499), 
        .Q(g1560) );
  SDFFX1 DFF_904_Q_reg ( .D(g25250), .SI(g1560), .SE(n10312), .CLK(n10499), 
        .Q(g1561) );
  SDFFX1 DFF_905_Q_reg ( .D(g25255), .SI(g1561), .SE(n10312), .CLK(n10499), 
        .Q(g1559) );
  SDFFX1 DFF_906_Q_reg ( .D(g30279), .SI(g1559), .SE(n10322), .CLK(n10509), 
        .Q(g1567) );
  SDFFX1 DFF_907_Q_reg ( .D(g30287), .SI(g1567), .SE(n10322), .CLK(n10509), 
        .Q(g1570) );
  SDFFX1 DFF_908_Q_reg ( .D(g30294), .SI(g1570), .SE(n10322), .CLK(n10509), 
        .Q(g1573) );
  SDFFX1 DFF_909_Q_reg ( .D(g30651), .SI(g1573), .SE(n10322), .CLK(n10509), 
        .Q(g1612) );
  SDFFX1 DFF_910_Q_reg ( .D(g30657), .SI(g1612), .SE(n10322), .CLK(n10509), 
        .Q(g1615) );
  SDFFX1 DFF_911_Q_reg ( .D(g30663), .SI(g1615), .SE(n10322), .CLK(n10509), 
        .Q(g1618) );
  SDFFX1 DFF_912_Q_reg ( .D(g30683), .SI(g1618), .SE(n10322), .CLK(n10509), 
        .Q(g1576) );
  SDFFX1 DFF_913_Q_reg ( .D(g30688), .SI(g1576), .SE(n10322), .CLK(n10509), 
        .Q(g1579) );
  SDFFX1 DFF_914_Q_reg ( .D(g30692), .SI(g1579), .SE(n10319), .CLK(n10506), 
        .Q(g1582) );
  SDFFX1 DFF_915_Q_reg ( .D(g30658), .SI(g1582), .SE(n10319), .CLK(n10506), 
        .Q(test_so55) );
  SDFFX1 DFF_916_Q_reg ( .D(g30664), .SI(test_si56), .SE(n10317), .CLK(n10504), 
        .Q(g1624) );
  SDFFX1 DFF_917_Q_reg ( .D(g30671), .SI(g1624), .SE(n10317), .CLK(n10504), 
        .Q(g1627) );
  SDFFX1 DFF_918_Q_reg ( .D(g30295), .SI(g1627), .SE(n10317), .CLK(n10504), 
        .Q(g1585) );
  SDFFX1 DFF_919_Q_reg ( .D(g30299), .SI(g1585), .SE(n10317), .CLK(n10504), 
        .Q(g1588) );
  SDFFX1 DFF_920_Q_reg ( .D(g30302), .SI(g1588), .SE(n10317), .CLK(n10504), 
        .Q(g1591) );
  SDFFX1 DFF_921_Q_reg ( .D(g30266), .SI(g1591), .SE(n10317), .CLK(n10504), 
        .Q(g1630) );
  SDFFX1 DFF_922_Q_reg ( .D(g30272), .SI(g1630), .SE(n10317), .CLK(n10504), 
        .Q(g1633) );
  SDFFX1 DFF_923_Q_reg ( .D(g30280), .SI(g1633), .SE(n10318), .CLK(n10505), 
        .Q(g1636) );
  SDFFX1 DFF_924_Q_reg ( .D(g30250), .SI(g1636), .SE(n10318), .CLK(n10505), 
        .Q(g1594) );
  SDFFX1 DFF_925_Q_reg ( .D(g30252), .SI(g1594), .SE(n10318), .CLK(n10505), 
        .Q(g1597) );
  SDFFX1 DFF_926_Q_reg ( .D(g30255), .SI(g1597), .SE(n10318), .CLK(n10505), 
        .Q(g1600) );
  SDFFX1 DFF_927_Q_reg ( .D(g30273), .SI(g1600), .SE(n10318), .CLK(n10505), 
        .Q(g1639) );
  SDFFX1 DFF_928_Q_reg ( .D(g30281), .SI(g1639), .SE(n10318), .CLK(n10505), 
        .Q(g1642) );
  SDFFX1 DFF_929_Q_reg ( .D(g30288), .SI(g1642), .SE(n10318), .CLK(n10505), 
        .Q(g1645) );
  SDFFX1 DFF_930_Q_reg ( .D(g30644), .SI(g1645), .SE(n10318), .CLK(n10505), 
        .Q(g1603) );
  SDFFX1 DFF_931_Q_reg ( .D(g30650), .SI(g1603), .SE(n10318), .CLK(n10505), 
        .Q(test_so56) );
  SDFFX1 DFF_932_Q_reg ( .D(g30656), .SI(test_si57), .SE(n10318), .CLK(n10505), 
        .Q(g1609) );
  SDFFX1 DFF_933_Q_reg ( .D(g30678), .SI(g1609), .SE(n10318), .CLK(n10505), 
        .Q(g1648) );
  SDFFX1 DFF_934_Q_reg ( .D(g30684), .SI(g1648), .SE(n10318), .CLK(n10505), 
        .Q(g1651) );
  SDFFX1 DFF_935_Q_reg ( .D(g30689), .SI(g1651), .SE(n10312), .CLK(n10499), 
        .Q(g1654) );
  SDFFX1 DFF_936_Q_reg ( .D(g25056), .SI(g1654), .SE(n10313), .CLK(n10500), 
        .Q(g1466), .QN(n9883) );
  SDFFX1 DFF_937_Q_reg ( .D(g25938), .SI(g1466), .SE(n10313), .CLK(n10500), 
        .Q(g1462), .QN(n10185) );
  SDFFX1 DFF_938_Q_reg ( .D(g26531), .SI(g1462), .SE(n10313), .CLK(n10500), 
        .Q(g1457), .QN(n9882) );
  SDFFX1 DFF_939_Q_reg ( .D(g27129), .SI(g1457), .SE(n10313), .CLK(n10500), 
        .Q(g1453), .QN(n10186) );
  SDFFX1 DFF_940_Q_reg ( .D(g27612), .SI(g1453), .SE(n10313), .CLK(n10500), 
        .Q(g1448), .QN(n9881) );
  SDFFX1 DFF_941_Q_reg ( .D(g28147), .SI(g1448), .SE(n10313), .CLK(n10500), 
        .Q(g1444), .QN(n10168) );
  SDFFX1 DFF_942_Q_reg ( .D(g28636), .SI(g1444), .SE(n10313), .CLK(n10500), 
        .Q(g1439), .QN(n9880) );
  SDFFX1 DFF_943_Q_reg ( .D(g29111), .SI(g1439), .SE(n10313), .CLK(n10500), 
        .Q(g1435), .QN(n10174) );
  SDFFX1 DFF_944_Q_reg ( .D(g29355), .SI(g1435), .SE(n10313), .CLK(n10500), 
        .Q(g1430), .QN(n9508) );
  SDFFX1 DFF_945_Q_reg ( .D(g29581), .SI(g1430), .SE(n10313), .CLK(n10500), 
        .Q(g1426), .QN(n9354) );
  SDFFX1 DFF_946_Q_reg ( .D(n29), .SI(g1426), .SE(n10313), .CLK(n10500), .Q(
        g1562) );
  SDFFX1 DFF_947_Q_reg ( .D(g1562), .SI(g1562), .SE(n10313), .CLK(n10500), .Q(
        test_so57) );
  SDFFX1 DFF_948_Q_reg ( .D(test_so57), .SI(test_si58), .SE(n10314), .CLK(
        n10501), .Q(g1563), .QN(n10161) );
  SDFFX1 DFF_949_Q_reg ( .D(g2950), .SI(g1563), .SE(n10314), .CLK(n10501), .Q(
        g5511), .QN(n4518) );
  SDFFX1 DFF_952_Q_reg ( .D(test_so57), .SI(n4618), .SE(n10314), .CLK(n10501), 
        .Q(g1690), .QN(n4386) );
  SDFFX1 DFF_953_Q_reg ( .D(g27264), .SI(g1690), .SE(n10321), .CLK(n10508), 
        .Q(g1735), .QN(n9837) );
  SDFFX1 DFF_954_Q_reg ( .D(g27274), .SI(g1735), .SE(n10321), .CLK(n10508), 
        .Q(g1724), .QN(n9836) );
  SDFFX1 DFF_955_Q_reg ( .D(g27287), .SI(g1724), .SE(n10321), .CLK(n10508), 
        .Q(g1727), .QN(n9835) );
  SDFFX1 DFF_956_Q_reg ( .D(g27275), .SI(g1727), .SE(n10321), .CLK(n10508), 
        .Q(g1750), .QN(n9814) );
  SDFFX1 DFF_957_Q_reg ( .D(g27288), .SI(g1750), .SE(n10321), .CLK(n10508), 
        .Q(g1739), .QN(n9813) );
  SDFFX1 DFF_958_Q_reg ( .D(g27302), .SI(g1739), .SE(n10321), .CLK(n10508), 
        .Q(g1742), .QN(n9812) );
  SDFFX1 DFF_959_Q_reg ( .D(g27289), .SI(g1742), .SE(n10321), .CLK(n10508), 
        .Q(g1765), .QN(n9559) );
  SDFFX1 DFF_960_Q_reg ( .D(g27303), .SI(g1765), .SE(n10321), .CLK(n10508), 
        .Q(g1754), .QN(n9561) );
  SDFFX1 DFF_961_Q_reg ( .D(g27317), .SI(g1754), .SE(n10321), .CLK(n10508), 
        .Q(g1757), .QN(n9560) );
  SDFFX1 DFF_962_Q_reg ( .D(g27304), .SI(g1757), .SE(n10322), .CLK(n10509), 
        .Q(g1779), .QN(n9825) );
  SDFFX1 DFF_963_Q_reg ( .D(g27318), .SI(g1779), .SE(n10322), .CLK(n10509), 
        .Q(test_so58) );
  SDFFX1 DFF_964_Q_reg ( .D(g27330), .SI(test_si59), .SE(n10319), .CLK(n10506), 
        .Q(g1772), .QN(n9824) );
  SDFFX1 DFF_965_Q_reg ( .D(g28749), .SI(g1772), .SE(n10319), .CLK(n10506), 
        .Q(g1789) );
  SDFFX1 DFF_966_Q_reg ( .D(g28760), .SI(g1789), .SE(n10320), .CLK(n10507), 
        .Q(g1792) );
  SDFFX1 DFF_967_Q_reg ( .D(g28771), .SI(g1792), .SE(n10320), .CLK(n10507), 
        .Q(g1795) );
  SDFFX1 DFF_968_Q_reg ( .D(g29205), .SI(g1795), .SE(n10321), .CLK(n10508), 
        .Q(g1798) );
  SDFFX1 DFF_969_Q_reg ( .D(g29212), .SI(g1798), .SE(n10321), .CLK(n10508), 
        .Q(g1801) );
  SDFFX1 DFF_970_Q_reg ( .D(g29218), .SI(g1801), .SE(n10319), .CLK(n10506), 
        .Q(g1804) );
  SDFFX1 DFF_971_Q_reg ( .D(g28761), .SI(g1804), .SE(n10319), .CLK(n10506), 
        .Q(g1808), .QN(n9860) );
  SDFFX1 DFF_972_Q_reg ( .D(g28772), .SI(g1808), .SE(n10319), .CLK(n10506), 
        .Q(g1809), .QN(n9848) );
  SDFFX1 DFF_973_Q_reg ( .D(g28778), .SI(g1809), .SE(n10319), .CLK(n10506), 
        .Q(g1807), .QN(n9859) );
  SDFFX1 DFF_974_Q_reg ( .D(g26811), .SI(g1807), .SE(n10319), .CLK(n10506), 
        .Q(g1810) );
  SDFFX1 DFF_975_Q_reg ( .D(g26815), .SI(g1810), .SE(n10320), .CLK(n10507), 
        .Q(g1813) );
  SDFFX1 DFF_976_Q_reg ( .D(g26820), .SI(g1813), .SE(n10320), .CLK(n10507), 
        .Q(g1816) );
  SDFFX1 DFF_977_Q_reg ( .D(g26816), .SI(g1816), .SE(n10320), .CLK(n10507), 
        .Q(g1819) );
  SDFFX1 DFF_978_Q_reg ( .D(g26821), .SI(g1819), .SE(n10320), .CLK(n10507), 
        .Q(g1822) );
  SDFFX1 DFF_979_Q_reg ( .D(g26824), .SI(g1822), .SE(n10320), .CLK(n10507), 
        .Q(test_so59) );
  SDFFX1 DFF_980_Q_reg ( .D(g27764), .SI(test_si60), .SE(n10320), .CLK(n10507), 
        .Q(g1829), .QN(n9858) );
  SDFFX1 DFF_981_Q_reg ( .D(g27766), .SI(g1829), .SE(n10320), .CLK(n10507), 
        .Q(g1830), .QN(n9847) );
  SDFFX1 DFF_982_Q_reg ( .D(g27768), .SI(g1830), .SE(n10320), .CLK(n10507), 
        .Q(g1828), .QN(n9857) );
  SDFFX1 DFF_983_Q_reg ( .D(g29613), .SI(g1828), .SE(n10320), .CLK(n10507), 
        .Q(g1693), .QN(n9464) );
  SDFFX1 DFF_984_Q_reg ( .D(g29617), .SI(g1693), .SE(n10320), .CLK(n10507), 
        .Q(g1694), .QN(n9449) );
  SDFFX1 DFF_985_Q_reg ( .D(g29620), .SI(g1694), .SE(n10319), .CLK(n10506), 
        .Q(g1695), .QN(n9463) );
  SDFFX1 DFF_986_Q_reg ( .D(g30704), .SI(g1695), .SE(n10319), .CLK(n10506), 
        .Q(g1696), .QN(n9462) );
  SDFFX1 DFF_987_Q_reg ( .D(g30706), .SI(g1696), .SE(n10319), .CLK(n10506), 
        .Q(g1697), .QN(n9448) );
  SDFFX1 DFF_988_Q_reg ( .D(g30708), .SI(g1697), .SE(n10312), .CLK(n10499), 
        .Q(g1698), .QN(n9461) );
  SDFFX1 DFF_989_Q_reg ( .D(g30487), .SI(g1698), .SE(n10314), .CLK(n10501), 
        .Q(g1699), .QN(n9460) );
  SDFFX1 DFF_990_Q_reg ( .D(g30503), .SI(g1699), .SE(n10312), .CLK(n10499), 
        .Q(g1700), .QN(n9447) );
  SDFFX1 DFF_991_Q_reg ( .D(g30338), .SI(g1700), .SE(n10314), .CLK(n10501), 
        .Q(g1701), .QN(n9459) );
  SDFFX1 DFF_992_Q_reg ( .D(g29178), .SI(g1701), .SE(n10322), .CLK(n10509), 
        .Q(g1703) );
  SDFFX1 DFF_993_Q_reg ( .D(g29181), .SI(g1703), .SE(n10322), .CLK(n10509), 
        .Q(g1704) );
  SDFFX1 DFF_994_Q_reg ( .D(g29184), .SI(g1704), .SE(n10323), .CLK(n10510), 
        .Q(g1702) );
  SDFFX1 DFF_995_Q_reg ( .D(g26667), .SI(g1702), .SE(n10323), .CLK(n10510), 
        .Q(test_so60), .QN(n10211) );
  SDFFX1 DFF_996_Q_reg ( .D(g26670), .SI(test_si61), .SE(n10323), .CLK(n10510), 
        .Q(g1785), .QN(n9846) );
  SDFFX1 DFF_997_Q_reg ( .D(g26675), .SI(g1785), .SE(n10323), .CLK(n10510), 
        .Q(g1783), .QN(n9856) );
  SDFFX1 DFF_998_Q_reg ( .D(n4288), .SI(g1783), .SE(n10323), .CLK(n10510), .Q(
        g1831) );
  SDFFX1 DFF_999_Q_reg ( .D(g1831), .SI(g1831), .SE(n10323), .CLK(n10510), .Q(
        n7988), .QN(DFF_999_n1) );
  SDFFX1 DFF_1000_Q_reg ( .D(n4565), .SI(n7988), .SE(n10323), .CLK(n10510), 
        .Q(g1833) );
  SDFFX1 DFF_1001_Q_reg ( .D(g1833), .SI(g1833), .SE(n10323), .CLK(n10510), 
        .Q(n7987), .QN(DFF_1001_n1) );
  SDFFX1 DFF_1002_Q_reg ( .D(n4557), .SI(n7987), .SE(n10323), .CLK(n10510), 
        .Q(g1835) );
  SDFFX1 DFF_1003_Q_reg ( .D(g1835), .SI(g1835), .SE(n10323), .CLK(n10510), 
        .Q(n7986), .QN(DFF_1003_n1) );
  SDFFX1 DFF_1004_Q_reg ( .D(n4326), .SI(n7986), .SE(n10323), .CLK(n10510), 
        .Q(g1661) );
  SDFFX1 DFF_1005_Q_reg ( .D(g1661), .SI(g1661), .SE(n10323), .CLK(n10510), 
        .Q(n7985), .QN(DFF_1005_n1) );
  SDFFX1 DFF_1006_Q_reg ( .D(n4390), .SI(n7985), .SE(n10324), .CLK(n10511), 
        .Q(g1663) );
  SDFFX1 DFF_1007_Q_reg ( .D(g1663), .SI(g1663), .SE(n10324), .CLK(n10511), 
        .Q(n7984), .QN(DFF_1007_n1) );
  SDFFX1 DFF_1008_Q_reg ( .D(n4320), .SI(n7984), .SE(n10324), .CLK(n10511), 
        .Q(g1665) );
  SDFFX1 DFF_1009_Q_reg ( .D(g1665), .SI(g1665), .SE(n10324), .CLK(n10511), 
        .Q(n7983), .QN(DFF_1009_n1) );
  SDFFX1 DFF_1010_Q_reg ( .D(n4374), .SI(n7983), .SE(n10324), .CLK(n10511), 
        .Q(g1667) );
  SDFFX1 DFF_1011_Q_reg ( .D(g1667), .SI(g1667), .SE(n10324), .CLK(n10511), 
        .Q(test_so61), .QN(DFF_1011_n1) );
  SDFFX1 DFF_1012_Q_reg ( .D(n4378), .SI(test_si62), .SE(n10227), .CLK(n10414), 
        .Q(g1669) );
  SDFFX1 DFF_1013_Q_reg ( .D(g1669), .SI(g1669), .SE(n10227), .CLK(n10414), 
        .Q(n7980), .QN(DFF_1013_n1) );
  SDFFX1 DFF_1014_Q_reg ( .D(g2877), .SI(n7980), .SE(n10238), .CLK(n10425), 
        .Q(g1671) );
  SDFFX1 DFF_1015_Q_reg ( .D(g1671), .SI(g1671), .SE(n10238), .CLK(n10425), 
        .Q(n7979), .QN(n4484) );
  SDFFX1 DFF_1016_Q_reg ( .D(n4284), .SI(n7979), .SE(n10321), .CLK(n10508), 
        .Q(g1680), .QN(n4488) );
  SDFFX1 DFF_1017_Q_reg ( .D(n532), .SI(g1680), .SE(n10337), .CLK(n10524), .Q(
        g1686) );
  SDFFX1 DFF_1028_Q_reg ( .D(n4276), .SI(g1686), .SE(n10324), .CLK(n10511), 
        .Q(n7978), .QN(n18261) );
  SDFFX1 DFF_1029_Q_reg ( .D(g1735), .SI(n7978), .SE(n10324), .CLK(n10511), 
        .Q(g1723) );
  SDFFX1 DFF_1030_Q_reg ( .D(g1723), .SI(g1723), .SE(n10324), .CLK(n10511), 
        .Q(g1730) );
  SDFFX1 DFF_1031_Q_reg ( .D(g1724), .SI(g1730), .SE(n10324), .CLK(n10511), 
        .Q(g1731) );
  SDFFX1 DFF_1032_Q_reg ( .D(g1731), .SI(g1731), .SE(n10324), .CLK(n10511), 
        .Q(g1732) );
  SDFFX1 DFF_1033_Q_reg ( .D(g1727), .SI(g1732), .SE(n10324), .CLK(n10511), 
        .Q(g1733) );
  SDFFX1 DFF_1034_Q_reg ( .D(g1733), .SI(g1733), .SE(n10325), .CLK(n10512), 
        .Q(g1734) );
  SDFFX1 DFF_1035_Q_reg ( .D(g1750), .SI(g1734), .SE(n10325), .CLK(n10512), 
        .Q(g1738) );
  SDFFX1 DFF_1036_Q_reg ( .D(g1738), .SI(g1738), .SE(n10325), .CLK(n10512), 
        .Q(g1745) );
  SDFFX1 DFF_1037_Q_reg ( .D(g1739), .SI(g1745), .SE(n10325), .CLK(n10512), 
        .Q(test_so62) );
  SDFFX1 DFF_1038_Q_reg ( .D(test_so62), .SI(test_si63), .SE(n10325), .CLK(
        n10512), .Q(g1747) );
  SDFFX1 DFF_1039_Q_reg ( .D(g1742), .SI(g1747), .SE(n10325), .CLK(n10512), 
        .Q(g1748) );
  SDFFX1 DFF_1040_Q_reg ( .D(g1748), .SI(g1748), .SE(n10325), .CLK(n10512), 
        .Q(g1749) );
  SDFFX1 DFF_1041_Q_reg ( .D(g1765), .SI(g1749), .SE(n10325), .CLK(n10512), 
        .Q(g1753) );
  SDFFX1 DFF_1042_Q_reg ( .D(g1753), .SI(g1753), .SE(n10325), .CLK(n10512), 
        .Q(g1760) );
  SDFFX1 DFF_1043_Q_reg ( .D(g1754), .SI(g1760), .SE(n10325), .CLK(n10512), 
        .Q(g1761) );
  SDFFX1 DFF_1044_Q_reg ( .D(g1761), .SI(g1761), .SE(n10325), .CLK(n10512), 
        .Q(g1762) );
  SDFFX1 DFF_1045_Q_reg ( .D(g1757), .SI(g1762), .SE(n10325), .CLK(n10512), 
        .Q(g1763) );
  SDFFX1 DFF_1046_Q_reg ( .D(g1763), .SI(g1763), .SE(n10326), .CLK(n10513), 
        .Q(g1764) );
  SDFFX1 DFF_1047_Q_reg ( .D(g1779), .SI(g1764), .SE(n10326), .CLK(n10513), 
        .Q(g1768) );
  SDFFX1 DFF_1048_Q_reg ( .D(g1768), .SI(g1768), .SE(n10326), .CLK(n10513), 
        .Q(g1775) );
  SDFFX1 DFF_1049_Q_reg ( .D(test_so58), .SI(g1775), .SE(n10326), .CLK(n10513), 
        .Q(g1776) );
  SDFFX1 DFF_1050_Q_reg ( .D(g1776), .SI(g1776), .SE(n10326), .CLK(n10513), 
        .Q(g1777) );
  SDFFX1 DFF_1051_Q_reg ( .D(g1772), .SI(g1777), .SE(n10326), .CLK(n10513), 
        .Q(g1778) );
  SDFFX1 DFF_1052_Q_reg ( .D(g1778), .SI(g1778), .SE(n10326), .CLK(n10513), 
        .Q(g1705) );
  SDFFX1 DFF_1053_Q_reg ( .D(n4598), .SI(g1705), .SE(n10326), .CLK(n10513), 
        .Q(test_so63) );
  SDFFX1 DFF_1054_Q_reg ( .D(test_so63), .SI(test_si64), .SE(n10326), .CLK(
        n10513), .Q(g5738) );
  SDFFX1 DFF_1055_Q_reg ( .D(g5738), .SI(g5738), .SE(n10326), .CLK(n10513), 
        .Q(g1718) );
  SDFFX1 DFF_1056_Q_reg ( .D(n4598), .SI(g1718), .SE(n10326), .CLK(n10513), 
        .Q(g7052), .QN(n4296) );
  SDFFX1 DFF_1057_Q_reg ( .D(g7052), .SI(g7052), .SE(n10326), .CLK(n10513), 
        .Q(g7194), .QN(n4315) );
  SDFFX1 DFF_1058_Q_reg ( .D(g7194), .SI(g7194), .SE(n10327), .CLK(n10514), 
        .Q(g1930), .QN(n4366) );
  SDFFX1 DFF_1059_Q_reg ( .D(g21845), .SI(g1930), .SE(n10327), .CLK(n10514), 
        .Q(g1934), .QN(n10121) );
  SDFFX1 DFF_1060_Q_reg ( .D(g18743), .SI(g1934), .SE(n10327), .CLK(n10514), 
        .Q(g1937) );
  SDFFX1 DFF_1061_Q_reg ( .D(g18794), .SI(g1937), .SE(n10327), .CLK(n10514), 
        .Q(g1890), .QN(n4297) );
  SDFFX1 DFF_1062_Q_reg ( .D(n1330), .SI(g1890), .SE(n10328), .CLK(n10515), 
        .Q(g1893) );
  SDFFX1 DFF_1063_Q_reg ( .D(g1893), .SI(g1893), .SE(n10328), .CLK(n10515), 
        .Q(g1903) );
  SDFFX1 DFF_1064_Q_reg ( .D(g1903), .SI(g1903), .SE(n10328), .CLK(n10515), 
        .Q(g1904) );
  SDFFX1 DFF_1065_Q_reg ( .D(g1836), .SI(g1904), .SE(n10328), .CLK(n10515), 
        .Q(g1944) );
  SDFFX1 DFF_1066_Q_reg ( .D(g1944), .SI(g1944), .SE(n10328), .CLK(n10515), 
        .Q(g1949) );
  SDFFX1 DFF_1067_Q_reg ( .D(test_so65), .SI(g1949), .SE(n10328), .CLK(n10515), 
        .Q(g1950) );
  SDFFX1 DFF_1068_Q_reg ( .D(g1950), .SI(g1950), .SE(n10328), .CLK(n10515), 
        .Q(g1951) );
  SDFFX1 DFF_1069_Q_reg ( .D(g1842), .SI(g1951), .SE(n10328), .CLK(n10515), 
        .Q(test_so64) );
  SDFFX1 DFF_1070_Q_reg ( .D(test_so64), .SI(test_si65), .SE(n10329), .CLK(
        n10516), .Q(g1953) );
  SDFFX1 DFF_1071_Q_reg ( .D(g1846), .SI(g1953), .SE(n10329), .CLK(n10516), 
        .Q(g1954) );
  SDFFX1 DFF_1072_Q_reg ( .D(g1954), .SI(g1954), .SE(n10329), .CLK(n10516), 
        .Q(g1945) );
  SDFFX1 DFF_1073_Q_reg ( .D(g1849), .SI(g1945), .SE(n10329), .CLK(n10516), 
        .Q(g1946) );
  SDFFX1 DFF_1074_Q_reg ( .D(g1946), .SI(g1946), .SE(n10329), .CLK(n10516), 
        .Q(g1947) );
  SDFFX1 DFF_1075_Q_reg ( .D(g1852), .SI(g1947), .SE(n10329), .CLK(n10516), 
        .Q(g1948) );
  SDFFX1 DFF_1076_Q_reg ( .D(g1948), .SI(g1948), .SE(n10329), .CLK(n10516), 
        .Q(g1870) );
  SDFFX1 DFF_1077_Q_reg ( .D(g2950), .SI(g1870), .SE(n10329), .CLK(n10516), 
        .Q(g8012), .QN(n4458) );
  SDFFX1 DFF_1078_Q_reg ( .D(g8012), .SI(g8012), .SE(n10329), .CLK(n10516), 
        .Q(g8082), .QN(n4457) );
  SDFFX1 DFF_1079_Q_reg ( .D(g8082), .SI(g8082), .SE(n10329), .CLK(n10516), 
        .Q(g1866), .QN(n4464) );
  SDFFX1 DFF_1080_Q_reg ( .D(g23097), .SI(g1866), .SE(n10330), .CLK(n10517), 
        .Q(g1867) );
  SDFFX1 DFF_1081_Q_reg ( .D(g23124), .SI(g1867), .SE(n10330), .CLK(n10517), 
        .Q(g1868) );
  SDFFX1 DFF_1082_Q_reg ( .D(g23137), .SI(g1868), .SE(n10330), .CLK(n10517), 
        .Q(g1869) );
  SDFFX1 DFF_1083_Q_reg ( .D(g23400), .SI(g1869), .SE(n10330), .CLK(n10517), 
        .Q(g1836) );
  SDFFX1 DFF_1084_Q_reg ( .D(g23413), .SI(g1836), .SE(n10331), .CLK(n10518), 
        .Q(test_so65) );
  SDFFX1 DFF_1085_Q_reg ( .D(g24182), .SI(test_si66), .SE(n10329), .CLK(n10516), .Q(g1842) );
  SDFFX1 DFF_1086_Q_reg ( .D(g24208), .SI(g1842), .SE(n10329), .CLK(n10516), 
        .Q(g1858) );
  SDFFX1 DFF_1087_Q_reg ( .D(g24219), .SI(g1858), .SE(n10330), .CLK(n10517), 
        .Q(g1859) );
  SDFFX1 DFF_1088_Q_reg ( .D(g24231), .SI(g1859), .SE(n10330), .CLK(n10517), 
        .Q(g1860) );
  SDFFX1 DFF_1089_Q_reg ( .D(g23123), .SI(g1860), .SE(n10330), .CLK(n10517), 
        .Q(g1861) );
  SDFFX1 DFF_1090_Q_reg ( .D(g23030), .SI(g1861), .SE(n10330), .CLK(n10517), 
        .Q(g1865) );
  SDFFX1 DFF_1091_Q_reg ( .D(g23058), .SI(g1865), .SE(n10330), .CLK(n10517), 
        .Q(g1845) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24218), .SI(g1845), .SE(n10330), .CLK(n10517), 
        .Q(g1846) );
  SDFFX1 DFF_1093_Q_reg ( .D(g24230), .SI(g1846), .SE(n10330), .CLK(n10517), 
        .Q(g1849) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24243), .SI(g1849), .SE(n10330), .CLK(n10517), 
        .Q(g1852) );
  SDFFX1 DFF_1095_Q_reg ( .D(n1305), .SI(g1852), .SE(n10331), .CLK(n10518), 
        .Q(g1908) );
  SDFFX1 DFF_1096_Q_reg ( .D(g1908), .SI(g1908), .SE(n10331), .CLK(n10518), 
        .Q(g1915) );
  SDFFX1 DFF_1097_Q_reg ( .D(g1915), .SI(g1915), .SE(n10331), .CLK(n10518), 
        .Q(g1922) );
  SDFFX1 DFF_1098_Q_reg ( .D(g13164), .SI(g1922), .SE(n10331), .CLK(n10518), 
        .Q(g1923) );
  SDFFX1 DFF_1099_Q_reg ( .D(g1923), .SI(g1923), .SE(n10331), .CLK(n10518), 
        .Q(test_so66), .QN(DFF_1099_n1) );
  SDFFX1 DFF_1100_Q_reg ( .D(n608), .SI(test_si67), .SE(n10333), .CLK(n10520), 
        .Q(n7971), .QN(DFF_1100_n1) );
  SDFFX1 DFF_1101_Q_reg ( .D(g13135), .SI(n7971), .SE(n10331), .CLK(n10518), 
        .Q(g1929) );
  SDFFX1 DFF_1102_Q_reg ( .D(g1929), .SI(g1929), .SE(n10331), .CLK(n10518), 
        .Q(g1880), .QN(n4545) );
  SDFFX1 DFF_1103_Q_reg ( .D(g13182), .SI(g1880), .SE(n10331), .CLK(n10518), 
        .Q(g1938) );
  SDFFX1 DFF_1104_Q_reg ( .D(g1938), .SI(g1938), .SE(n10331), .CLK(n10518), 
        .Q(g1939) );
  SDFFX1 DFF_1105_Q_reg ( .D(g27290), .SI(g1939), .SE(n10334), .CLK(n10521), 
        .Q(g1956), .QN(n9514) );
  SDFFX1 DFF_1106_Q_reg ( .D(g27305), .SI(g1956), .SE(n10334), .CLK(n10521), 
        .Q(g1957), .QN(n9516) );
  SDFFX1 DFF_1107_Q_reg ( .D(g27319), .SI(g1957), .SE(n10334), .CLK(n10521), 
        .Q(g1955), .QN(n9515) );
  SDFFX1 DFF_1108_Q_reg ( .D(g27306), .SI(g1955), .SE(n10334), .CLK(n10521), 
        .Q(g1959), .QN(n9526) );
  SDFFX1 DFF_1109_Q_reg ( .D(g27320), .SI(g1959), .SE(n10334), .CLK(n10521), 
        .Q(g1960), .QN(n9528) );
  SDFFX1 DFF_1110_Q_reg ( .D(g27331), .SI(g1960), .SE(n10334), .CLK(n10521), 
        .Q(g1958), .QN(n9527) );
  SDFFX1 DFF_1111_Q_reg ( .D(g27321), .SI(g1958), .SE(n10334), .CLK(n10521), 
        .Q(g1962), .QN(n9359) );
  SDFFX1 DFF_1112_Q_reg ( .D(g27332), .SI(g1962), .SE(n10334), .CLK(n10521), 
        .Q(g1963), .QN(n9361) );
  SDFFX1 DFF_1113_Q_reg ( .D(g27340), .SI(g1963), .SE(n10334), .CLK(n10521), 
        .Q(g1961), .QN(n9360) );
  SDFFX1 DFF_1114_Q_reg ( .D(g27333), .SI(g1961), .SE(n10334), .CLK(n10521), 
        .Q(test_so67), .QN(n10196) );
  SDFFX1 DFF_1115_Q_reg ( .D(g27341), .SI(test_si68), .SE(n10334), .CLK(n10521), .Q(g1966), .QN(n9538) );
  SDFFX1 DFF_1116_Q_reg ( .D(g27346), .SI(g1966), .SE(n10335), .CLK(n10522), 
        .Q(g1964), .QN(n9537) );
  SDFFX1 DFF_1117_Q_reg ( .D(g24513), .SI(g1964), .SE(n10335), .CLK(n10522), 
        .Q(g1967) );
  SDFFX1 DFF_1118_Q_reg ( .D(g24524), .SI(g1967), .SE(n10335), .CLK(n10522), 
        .Q(g1970) );
  SDFFX1 DFF_1119_Q_reg ( .D(g24534), .SI(g1970), .SE(n10335), .CLK(n10522), 
        .Q(g1973) );
  SDFFX1 DFF_1120_Q_reg ( .D(g24525), .SI(g1973), .SE(n10335), .CLK(n10522), 
        .Q(g1976) );
  SDFFX1 DFF_1121_Q_reg ( .D(g24535), .SI(g1976), .SE(n10335), .CLK(n10522), 
        .Q(g1979) );
  SDFFX1 DFF_1122_Q_reg ( .D(g24545), .SI(g1979), .SE(n10335), .CLK(n10522), 
        .Q(g1982) );
  SDFFX1 DFF_1123_Q_reg ( .D(g28357), .SI(g1982), .SE(n10335), .CLK(n10522), 
        .Q(g1994) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28362), .SI(g1994), .SE(n10335), .CLK(n10522), 
        .Q(g1997) );
  SDFFX1 DFF_1125_Q_reg ( .D(g28366), .SI(g1997), .SE(n10334), .CLK(n10521), 
        .Q(g2000) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28352), .SI(g2000), .SE(n10335), .CLK(n10522), 
        .Q(g1985) );
  SDFFX1 DFF_1127_Q_reg ( .D(g28356), .SI(g1985), .SE(n10335), .CLK(n10522), 
        .Q(g1988) );
  SDFFX1 DFF_1128_Q_reg ( .D(g28361), .SI(g1988), .SE(n10335), .CLK(n10522), 
        .Q(g1991) );
  SDFFX1 DFF_1129_Q_reg ( .D(g26559), .SI(g1991), .SE(n10336), .CLK(n10523), 
        .Q(test_so68) );
  SDFFX1 DFF_1130_Q_reg ( .D(g26573), .SI(test_si69), .SE(n10336), .CLK(n10523), .Q(g1874) );
  SDFFX1 DFF_1131_Q_reg ( .D(g26592), .SI(g1874), .SE(n10336), .CLK(n10523), 
        .Q(g1877) );
  SDFFX1 DFF_1132_Q_reg ( .D(g1880), .SI(g1877), .SE(n10336), .CLK(n10523), 
        .Q(g1886), .QN(n4493) );
  SDFFX1 DFF_1133_Q_reg ( .D(g22651), .SI(g1886), .SE(n10336), .CLK(n10523), 
        .Q(n7968), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(n631), .SI(n7968), .SE(n10336), .CLK(n10523), .Q(
        g16399), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(g16399), .SI(g16399), .SE(n10336), .CLK(n10523), 
        .Q(g1905), .QN(n9896) );
  SDFFX1 DFF_1144_Q_reg ( .D(DFF_999_n1), .SI(g1905), .SE(n10336), .CLK(n10523), .Q(n7967) );
  SDFFX1 DFF_1145_Q_reg ( .D(DFF_1001_n1), .SI(n7967), .SE(n10336), .CLK(
        n10523), .Q(n7966) );
  SDFFX1 DFF_1146_Q_reg ( .D(DFF_1003_n1), .SI(n7966), .SE(n10336), .CLK(
        n10523), .Q(n7965) );
  SDFFX1 DFF_1147_Q_reg ( .D(DFF_1005_n1), .SI(n7965), .SE(n10336), .CLK(
        n10523), .Q(n7964) );
  SDFFX1 DFF_1148_Q_reg ( .D(DFF_1007_n1), .SI(n7964), .SE(n10336), .CLK(
        n10523), .Q(n7963) );
  SDFFX1 DFF_1149_Q_reg ( .D(DFF_1009_n1), .SI(n7963), .SE(n10337), .CLK(
        n10524), .Q(n7962) );
  SDFFX1 DFF_1150_Q_reg ( .D(DFF_1011_n1), .SI(n7962), .SE(n10337), .CLK(
        n10524), .Q(g1916) );
  SDFFX1 DFF_1151_Q_reg ( .D(DFF_1013_n1), .SI(g1916), .SE(n10337), .CLK(
        n10524), .Q(g1917) );
  SDFFX1 DFF_1152_Q_reg ( .D(g24083), .SI(g1917), .SE(n10337), .CLK(n10524), 
        .Q(test_so69), .QN(n10201) );
  SDFFX1 DFF_1153_Q_reg ( .D(n4484), .SI(test_si70), .SE(n10238), .CLK(n10425), 
        .Q(n7960) );
  SDFFX1 DFF_1155_Q_reg ( .D(g7229), .SI(g7229), .SE(n10238), .CLK(n10425), 
        .Q(g7357), .QN(n4357) );
  SDFFX1 DFF_1156_Q_reg ( .D(g7357), .SI(g7357), .SE(n10238), .CLK(n10425), 
        .Q(g2009), .QN(n4293) );
  SDFFX1 DFF_1157_Q_reg ( .D(g16692), .SI(g2009), .SE(n10327), .CLK(n10514), 
        .Q(g2010), .QN(n10155) );
  SDFFX1 DFF_1158_Q_reg ( .D(g20353), .SI(g2010), .SE(n10327), .CLK(n10514), 
        .Q(g2039), .QN(n4427) );
  SDFFX1 DFF_1159_Q_reg ( .D(g20752), .SI(g2039), .SE(n10327), .CLK(n10514), 
        .Q(g2020), .QN(n4400) );
  SDFFX1 DFF_1160_Q_reg ( .D(g21972), .SI(g2020), .SE(n10327), .CLK(n10514), 
        .Q(g2013), .QN(n4474) );
  SDFFX1 DFF_1161_Q_reg ( .D(g23339), .SI(g2013), .SE(n10327), .CLK(n10514), 
        .Q(g2033), .QN(n4420) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24434), .SI(g2033), .SE(n10327), .CLK(n10514), 
        .Q(g2026), .QN(n4410) );
  SDFFX1 DFF_1163_Q_reg ( .D(g25194), .SI(g2026), .SE(n10327), .CLK(n10514), 
        .Q(g2040), .QN(n4399) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26671), .SI(g2040), .SE(n10327), .CLK(n10514), 
        .Q(g2052), .QN(n4409) );
  SDFFX1 DFF_1165_Q_reg ( .D(g26789), .SI(g2052), .SE(n10328), .CLK(n10515), 
        .Q(g2046), .QN(n4468) );
  SDFFX1 DFF_1166_Q_reg ( .D(g27682), .SI(g2046), .SE(n10328), .CLK(n10515), 
        .Q(g2059), .QN(n4473) );
  SDFFX1 DFF_1167_Q_reg ( .D(g27722), .SI(g2059), .SE(n10328), .CLK(n10515), 
        .Q(test_so70), .QN(n10194) );
  SDFFX1 DFF_1168_Q_reg ( .D(g28325), .SI(test_si71), .SE(n10328), .CLK(n10515), .Q(g2072), .QN(n4416) );
  SDFFX1 DFF_1169_Q_reg ( .D(g20899), .SI(g2072), .SE(n10337), .CLK(n10524), 
        .Q(g2079), .QN(n9974) );
  SDFFX1 DFF_1170_Q_reg ( .D(g20915), .SI(g2079), .SE(n10337), .CLK(n10524), 
        .Q(g2080), .QN(n9973) );
  SDFFX1 DFF_1171_Q_reg ( .D(g20934), .SI(g2080), .SE(n10337), .CLK(n10524), 
        .Q(g2078), .QN(n10028) );
  SDFFX1 DFF_1172_Q_reg ( .D(g20916), .SI(g2078), .SE(n10337), .CLK(n10524), 
        .Q(g2082), .QN(n9972) );
  SDFFX1 DFF_1173_Q_reg ( .D(g20935), .SI(g2082), .SE(n10337), .CLK(n10524), 
        .Q(g2083), .QN(n9971) );
  SDFFX1 DFF_1174_Q_reg ( .D(g20953), .SI(g2083), .SE(n10338), .CLK(n10525), 
        .Q(g2081), .QN(n10027) );
  SDFFX1 DFF_1175_Q_reg ( .D(g20936), .SI(g2081), .SE(n10338), .CLK(n10525), 
        .Q(g2085), .QN(n9970) );
  SDFFX1 DFF_1176_Q_reg ( .D(g20954), .SI(g2085), .SE(n10338), .CLK(n10525), 
        .Q(g2086), .QN(n9969) );
  SDFFX1 DFF_1177_Q_reg ( .D(g20977), .SI(g2086), .SE(n10338), .CLK(n10525), 
        .Q(g2084), .QN(n10026) );
  SDFFX1 DFF_1178_Q_reg ( .D(g20955), .SI(g2084), .SE(n10338), .CLK(n10525), 
        .Q(g2088), .QN(n9968) );
  SDFFX1 DFF_1179_Q_reg ( .D(g20978), .SI(g2088), .SE(n10338), .CLK(n10525), 
        .Q(g2089), .QN(n9967) );
  SDFFX1 DFF_1180_Q_reg ( .D(g20999), .SI(g2089), .SE(n10338), .CLK(n10525), 
        .Q(g2087), .QN(n10025) );
  SDFFX1 DFF_1181_Q_reg ( .D(g20979), .SI(g2087), .SE(n10339), .CLK(n10526), 
        .Q(g2091), .QN(n9966) );
  SDFFX1 DFF_1182_Q_reg ( .D(g21000), .SI(g2091), .SE(n10339), .CLK(n10526), 
        .Q(test_so71) );
  SDFFX1 DFF_1183_Q_reg ( .D(g21019), .SI(test_si72), .SE(n10339), .CLK(n10526), .Q(g2090), .QN(n10024) );
  SDFFX1 DFF_1184_Q_reg ( .D(g21001), .SI(g2090), .SE(n10339), .CLK(n10526), 
        .Q(g2094), .QN(n9965) );
  SDFFX1 DFF_1185_Q_reg ( .D(g21020), .SI(g2094), .SE(n10339), .CLK(n10526), 
        .Q(g2095), .QN(n9964) );
  SDFFX1 DFF_1186_Q_reg ( .D(g21039), .SI(g2095), .SE(n10339), .CLK(n10526), 
        .Q(g2093), .QN(n10023) );
  SDFFX1 DFF_1187_Q_reg ( .D(g21021), .SI(g2093), .SE(n10339), .CLK(n10526), 
        .Q(g2097), .QN(n9963) );
  SDFFX1 DFF_1188_Q_reg ( .D(g21040), .SI(g2097), .SE(n10339), .CLK(n10526), 
        .Q(g2098), .QN(n9962) );
  SDFFX1 DFF_1189_Q_reg ( .D(g21054), .SI(g2098), .SE(n10339), .CLK(n10526), 
        .Q(g2096), .QN(n10022) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21041), .SI(g2096), .SE(n10339), .CLK(n10526), 
        .Q(g2100), .QN(n9961) );
  SDFFX1 DFF_1191_Q_reg ( .D(g21055), .SI(g2100), .SE(n10339), .CLK(n10526), 
        .Q(g2101), .QN(n9960) );
  SDFFX1 DFF_1192_Q_reg ( .D(g21071), .SI(g2101), .SE(n10339), .CLK(n10526), 
        .Q(g2099), .QN(n10021) );
  SDFFX1 DFF_1193_Q_reg ( .D(g21056), .SI(g2099), .SE(n10340), .CLK(n10527), 
        .Q(g2103), .QN(n9959) );
  SDFFX1 DFF_1194_Q_reg ( .D(g21072), .SI(g2103), .SE(n10340), .CLK(n10527), 
        .Q(g2104), .QN(n9958) );
  SDFFX1 DFF_1195_Q_reg ( .D(g21080), .SI(g2104), .SE(n10340), .CLK(n10527), 
        .Q(g2102), .QN(n10020) );
  SDFFX1 DFF_1196_Q_reg ( .D(g20900), .SI(g2102), .SE(n10340), .CLK(n10527), 
        .Q(g2106), .QN(n9957) );
  SDFFX1 DFF_1197_Q_reg ( .D(g20917), .SI(g2106), .SE(n10340), .CLK(n10527), 
        .Q(test_so72) );
  SDFFX1 DFF_1198_Q_reg ( .D(g20937), .SI(test_si73), .SE(n10337), .CLK(n10524), .Q(g2105), .QN(n10019) );
  SDFFX1 DFF_1199_Q_reg ( .D(g20980), .SI(g2105), .SE(n10337), .CLK(n10524), 
        .Q(g2109), .QN(n9750) );
  SDFFX1 DFF_1200_Q_reg ( .D(g21002), .SI(g2109), .SE(n10338), .CLK(n10525), 
        .Q(g2110), .QN(n9742) );
  SDFFX1 DFF_1201_Q_reg ( .D(g21022), .SI(g2110), .SE(n10338), .CLK(n10525), 
        .Q(g2108), .QN(n9805) );
  SDFFX1 DFF_1202_Q_reg ( .D(g21003), .SI(g2108), .SE(n10338), .CLK(n10525), 
        .Q(g2112), .QN(n9749) );
  SDFFX1 DFF_1203_Q_reg ( .D(g21023), .SI(g2112), .SE(n10338), .CLK(n10525), 
        .Q(g2113), .QN(n9741) );
  SDFFX1 DFF_1204_Q_reg ( .D(g21042), .SI(g2113), .SE(n10338), .CLK(n10525), 
        .Q(g2111), .QN(n9804) );
  SDFFX1 DFF_1205_Q_reg ( .D(g25268), .SI(g2111), .SE(n10340), .CLK(n10527), 
        .Q(g2115) );
  SDFFX1 DFF_1206_Q_reg ( .D(g25271), .SI(g2115), .SE(n10340), .CLK(n10527), 
        .Q(g2116) );
  SDFFX1 DFF_1207_Q_reg ( .D(g25279), .SI(g2116), .SE(n10340), .CLK(n10527), 
        .Q(g2114) );
  SDFFX1 DFF_1208_Q_reg ( .D(g22249), .SI(g2114), .SE(n10340), .CLK(n10527), 
        .Q(g2118) );
  SDFFX1 DFF_1209_Q_reg ( .D(g22267), .SI(g2118), .SE(n10340), .CLK(n10527), 
        .Q(g2119) );
  SDFFX1 DFF_1210_Q_reg ( .D(g22280), .SI(g2119), .SE(n10233), .CLK(n10420), 
        .Q(g2117) );
  SDFFX1 DFF_1211_Q_reg ( .D(g2950), .SI(g2117), .SE(n10233), .CLK(n10420), 
        .Q(g6837), .QN(n4324) );
  SDFFX1 DFF_1212_Q_reg ( .D(g6837), .SI(g6837), .SE(n10233), .CLK(n10420), 
        .Q(test_so73), .QN(n10189) );
  SDFFX1 DFF_1213_Q_reg ( .D(test_so73), .SI(test_si74), .SE(n10233), .CLK(
        n10420), .Q(g2241), .QN(n4367) );
  SDFFX1 DFF_1214_Q_reg ( .D(g22170), .SI(g2241), .SE(n10242), .CLK(n10429), 
        .Q(g2206), .QN(n10067) );
  SDFFX1 DFF_1215_Q_reg ( .D(g22182), .SI(g2206), .SE(n10243), .CLK(n10430), 
        .Q(g2207), .QN(n10066) );
  SDFFX1 DFF_1216_Q_reg ( .D(g22192), .SI(g2207), .SE(n10243), .CLK(n10430), 
        .Q(g2205), .QN(n9704) );
  SDFFX1 DFF_1217_Q_reg ( .D(g22183), .SI(g2205), .SE(n10229), .CLK(n10416), 
        .Q(g2209), .QN(n10065) );
  SDFFX1 DFF_1218_Q_reg ( .D(g22193), .SI(g2209), .SE(n10243), .CLK(n10430), 
        .Q(g2210), .QN(n10064) );
  SDFFX1 DFF_1219_Q_reg ( .D(g22200), .SI(g2210), .SE(n10243), .CLK(n10430), 
        .Q(g2208), .QN(n9703) );
  SDFFX1 DFF_1220_Q_reg ( .D(g22045), .SI(g2208), .SE(n10243), .CLK(n10430), 
        .Q(g2218), .QN(n10063) );
  SDFFX1 DFF_1221_Q_reg ( .D(g22060), .SI(g2218), .SE(n10243), .CLK(n10430), 
        .Q(g2219), .QN(n10062) );
  SDFFX1 DFF_1222_Q_reg ( .D(g22076), .SI(g2219), .SE(n10243), .CLK(n10430), 
        .Q(g2217), .QN(n9702) );
  SDFFX1 DFF_1223_Q_reg ( .D(g22061), .SI(g2217), .SE(n10243), .CLK(n10430), 
        .Q(g2221), .QN(n10061) );
  SDFFX1 DFF_1224_Q_reg ( .D(g22077), .SI(g2221), .SE(n10243), .CLK(n10430), 
        .Q(g2222), .QN(n10060) );
  SDFFX1 DFF_1225_Q_reg ( .D(g22097), .SI(g2222), .SE(n10243), .CLK(n10430), 
        .Q(g2220), .QN(n9701) );
  SDFFX1 DFF_1226_Q_reg ( .D(g22078), .SI(g2220), .SE(n10243), .CLK(n10430), 
        .Q(g2224), .QN(n10059) );
  SDFFX1 DFF_1227_Q_reg ( .D(g22098), .SI(g2224), .SE(n10244), .CLK(n10431), 
        .Q(test_so74), .QN(n10216) );
  SDFFX1 DFF_1228_Q_reg ( .D(g22115), .SI(test_si75), .SE(n10243), .CLK(n10430), .Q(g2223), .QN(n9700) );
  SDFFX1 DFF_1229_Q_reg ( .D(g22099), .SI(g2223), .SE(n10244), .CLK(n10431), 
        .Q(g2227), .QN(n10058) );
  SDFFX1 DFF_1230_Q_reg ( .D(g22116), .SI(g2227), .SE(n10244), .CLK(n10431), 
        .Q(g2228), .QN(n10057) );
  SDFFX1 DFF_1231_Q_reg ( .D(g22138), .SI(g2228), .SE(n10244), .CLK(n10431), 
        .Q(g2226), .QN(n9699) );
  SDFFX1 DFF_1232_Q_reg ( .D(g22117), .SI(g2226), .SE(n10244), .CLK(n10431), 
        .Q(g2230), .QN(n10056) );
  SDFFX1 DFF_1233_Q_reg ( .D(g22139), .SI(g2230), .SE(n10244), .CLK(n10431), 
        .Q(g2231), .QN(n10055) );
  SDFFX1 DFF_1234_Q_reg ( .D(g22153), .SI(g2231), .SE(n10244), .CLK(n10431), 
        .Q(g2229), .QN(n9698) );
  SDFFX1 DFF_1235_Q_reg ( .D(g22140), .SI(g2229), .SE(n10245), .CLK(n10432), 
        .Q(g2233), .QN(n10054) );
  SDFFX1 DFF_1236_Q_reg ( .D(g22154), .SI(g2233), .SE(n10245), .CLK(n10432), 
        .Q(g2234), .QN(n10053) );
  SDFFX1 DFF_1237_Q_reg ( .D(g22171), .SI(g2234), .SE(n10245), .CLK(n10432), 
        .Q(g2232), .QN(n9697) );
  SDFFX1 DFF_1238_Q_reg ( .D(g22155), .SI(g2232), .SE(n10245), .CLK(n10432), 
        .Q(g2236), .QN(n9688) );
  SDFFX1 DFF_1239_Q_reg ( .D(g22172), .SI(g2236), .SE(n10246), .CLK(n10433), 
        .Q(g2237), .QN(n9687) );
  SDFFX1 DFF_1240_Q_reg ( .D(g22184), .SI(g2237), .SE(n10246), .CLK(n10433), 
        .Q(g2235), .QN(n9686) );
  SDFFX1 DFF_1241_Q_reg ( .D(g22173), .SI(g2235), .SE(n10246), .CLK(n10433), 
        .Q(g2239), .QN(n9696) );
  SDFFX1 DFF_1242_Q_reg ( .D(g22185), .SI(g2239), .SE(n10246), .CLK(n10433), 
        .Q(test_so75), .QN(n10215) );
  SDFFX1 DFF_1243_Q_reg ( .D(g22194), .SI(test_si76), .SE(n10245), .CLK(n10432), .Q(g2238), .QN(n9695) );
  SDFFX1 DFF_1244_Q_reg ( .D(g25227), .SI(g2238), .SE(n10245), .CLK(n10432), 
        .Q(g2245), .QN(n9766) );
  SDFFX1 DFF_1245_Q_reg ( .D(g25236), .SI(g2245), .SE(n10245), .CLK(n10432), 
        .Q(g2246), .QN(n9765) );
  SDFFX1 DFF_1246_Q_reg ( .D(g25245), .SI(g2246), .SE(n10244), .CLK(n10431), 
        .Q(g2244), .QN(n9764) );
  SDFFX1 DFF_1247_Q_reg ( .D(g25237), .SI(g2244), .SE(n10244), .CLK(n10431), 
        .Q(g2248), .QN(n9763) );
  SDFFX1 DFF_1248_Q_reg ( .D(g25246), .SI(g2248), .SE(n10244), .CLK(n10431), 
        .Q(g2249), .QN(n9762) );
  SDFFX1 DFF_1249_Q_reg ( .D(g25251), .SI(g2249), .SE(n10244), .CLK(n10431), 
        .Q(g2247), .QN(n9761) );
  SDFFX1 DFF_1250_Q_reg ( .D(g25247), .SI(g2247), .SE(n10244), .CLK(n10431), 
        .Q(g2251), .QN(n9760) );
  SDFFX1 DFF_1251_Q_reg ( .D(g25252), .SI(g2251), .SE(n10245), .CLK(n10432), 
        .Q(g2252), .QN(n9759) );
  SDFFX1 DFF_1252_Q_reg ( .D(g25256), .SI(g2252), .SE(n10245), .CLK(n10432), 
        .Q(g2250), .QN(n9758) );
  SDFFX1 DFF_1253_Q_reg ( .D(g25253), .SI(g2250), .SE(n10245), .CLK(n10432), 
        .Q(g2254) );
  SDFFX1 DFF_1254_Q_reg ( .D(g25257), .SI(g2254), .SE(n10245), .CLK(n10432), 
        .Q(g2255) );
  SDFFX1 DFF_1255_Q_reg ( .D(g25259), .SI(g2255), .SE(n10245), .CLK(n10432), 
        .Q(g2253) );
  SDFFX1 DFF_1256_Q_reg ( .D(g30289), .SI(g2253), .SE(n10256), .CLK(n10443), 
        .Q(g2261) );
  SDFFX1 DFF_1257_Q_reg ( .D(g30296), .SI(g2261), .SE(n10256), .CLK(n10443), 
        .Q(test_so76) );
  SDFFX1 DFF_1258_Q_reg ( .D(g30300), .SI(test_si77), .SE(n10256), .CLK(n10443), .Q(g2267) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30660), .SI(g2267), .SE(n10256), .CLK(n10443), 
        .Q(g2306) );
  SDFFX1 DFF_1260_Q_reg ( .D(g30666), .SI(g2306), .SE(n10256), .CLK(n10443), 
        .Q(g2309) );
  SDFFX1 DFF_1261_Q_reg ( .D(g30672), .SI(g2309), .SE(n10248), .CLK(n10435), 
        .Q(g2312) );
  SDFFX1 DFF_1262_Q_reg ( .D(g30690), .SI(g2312), .SE(n10248), .CLK(n10435), 
        .Q(g2270) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30693), .SI(g2270), .SE(n10248), .CLK(n10435), 
        .Q(g2273) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30695), .SI(g2273), .SE(n10246), .CLK(n10433), 
        .Q(g2276) );
  SDFFX1 DFF_1265_Q_reg ( .D(g30667), .SI(g2276), .SE(n10246), .CLK(n10433), 
        .Q(g2315) );
  SDFFX1 DFF_1266_Q_reg ( .D(g30673), .SI(g2315), .SE(n10247), .CLK(n10434), 
        .Q(g2318) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30679), .SI(g2318), .SE(n10247), .CLK(n10434), 
        .Q(g2321) );
  SDFFX1 DFF_1268_Q_reg ( .D(g30301), .SI(g2321), .SE(n10247), .CLK(n10434), 
        .Q(g2279) );
  SDFFX1 DFF_1269_Q_reg ( .D(g30303), .SI(g2279), .SE(n10247), .CLK(n10434), 
        .Q(g2282) );
  SDFFX1 DFF_1270_Q_reg ( .D(g30304), .SI(g2282), .SE(n10247), .CLK(n10434), 
        .Q(g2285) );
  SDFFX1 DFF_1271_Q_reg ( .D(g30274), .SI(g2285), .SE(n10247), .CLK(n10434), 
        .Q(g2324) );
  SDFFX1 DFF_1272_Q_reg ( .D(g30282), .SI(g2324), .SE(n10247), .CLK(n10434), 
        .Q(test_so77) );
  SDFFX1 DFF_1273_Q_reg ( .D(g30290), .SI(test_si78), .SE(n10247), .CLK(n10434), .Q(g2330) );
  SDFFX1 DFF_1274_Q_reg ( .D(g30253), .SI(g2330), .SE(n10247), .CLK(n10434), 
        .Q(g2288) );
  SDFFX1 DFF_1275_Q_reg ( .D(g30256), .SI(g2288), .SE(n10247), .CLK(n10434), 
        .Q(g2291) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30260), .SI(g2291), .SE(n10247), .CLK(n10434), 
        .Q(g2294) );
  SDFFX1 DFF_1277_Q_reg ( .D(g30283), .SI(g2294), .SE(n10247), .CLK(n10434), 
        .Q(g2333) );
  SDFFX1 DFF_1278_Q_reg ( .D(g30291), .SI(g2333), .SE(n10248), .CLK(n10435), 
        .Q(g2336) );
  SDFFX1 DFF_1279_Q_reg ( .D(g30297), .SI(g2336), .SE(n10246), .CLK(n10433), 
        .Q(g2339) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30652), .SI(g2339), .SE(n10246), .CLK(n10433), 
        .Q(g2297) );
  SDFFX1 DFF_1281_Q_reg ( .D(g30659), .SI(g2297), .SE(n10246), .CLK(n10433), 
        .Q(g2300) );
  SDFFX1 DFF_1282_Q_reg ( .D(g30665), .SI(g2300), .SE(n10246), .CLK(n10433), 
        .Q(g2303) );
  SDFFX1 DFF_1283_Q_reg ( .D(g30686), .SI(g2303), .SE(n10246), .CLK(n10433), 
        .Q(g2342) );
  SDFFX1 DFF_1284_Q_reg ( .D(g30691), .SI(g2342), .SE(n10246), .CLK(n10433), 
        .Q(g2345) );
  SDFFX1 DFF_1285_Q_reg ( .D(g30694), .SI(g2345), .SE(n10229), .CLK(n10416), 
        .Q(g2348) );
  SDFFX1 DFF_1286_Q_reg ( .D(g25067), .SI(g2348), .SE(n10233), .CLK(n10420), 
        .Q(g2160), .QN(n9879) );
  SDFFX1 DFF_1287_Q_reg ( .D(g25940), .SI(g2160), .SE(n10233), .CLK(n10420), 
        .Q(test_so78) );
  SDFFX1 DFF_1288_Q_reg ( .D(g26532), .SI(test_si79), .SE(n10233), .CLK(n10420), .Q(g2151), .QN(n9878) );
  SDFFX1 DFF_1289_Q_reg ( .D(g27131), .SI(g2151), .SE(n10234), .CLK(n10421), 
        .Q(g2147), .QN(n10187) );
  SDFFX1 DFF_1290_Q_reg ( .D(g27621), .SI(g2147), .SE(n10234), .CLK(n10421), 
        .Q(g2142), .QN(n9877) );
  SDFFX1 DFF_1291_Q_reg ( .D(g28148), .SI(g2142), .SE(n10234), .CLK(n10421), 
        .Q(g2138), .QN(n10169) );
  SDFFX1 DFF_1292_Q_reg ( .D(g28637), .SI(g2138), .SE(n10234), .CLK(n10421), 
        .Q(g2133), .QN(n9876) );
  SDFFX1 DFF_1293_Q_reg ( .D(g29112), .SI(g2133), .SE(n10234), .CLK(n10421), 
        .Q(g2129), .QN(n10175) );
  SDFFX1 DFF_1294_Q_reg ( .D(g29357), .SI(g2129), .SE(n10234), .CLK(n10421), 
        .Q(g2124), .QN(n9507) );
  SDFFX1 DFF_1295_Q_reg ( .D(g29582), .SI(g2124), .SE(n10234), .CLK(n10421), 
        .Q(g2120), .QN(n9353) );
  SDFFX1 DFF_1296_Q_reg ( .D(n29), .SI(g2120), .SE(n10228), .CLK(n10415), .Q(
        g2256) );
  SDFFX1 DFF_1297_Q_reg ( .D(g2256), .SI(g2256), .SE(n10228), .CLK(n10415), 
        .Q(g5637) );
  SDFFX1 DFF_1298_Q_reg ( .D(g5637), .SI(g5637), .SE(n10228), .CLK(n10415), 
        .Q(g2257), .QN(n10162) );
  SDFFX1 DFF_1299_Q_reg ( .D(g2950), .SI(g2257), .SE(n10228), .CLK(n10415), 
        .Q(g5555), .QN(n4516) );
  SDFFX1 DFF_1302_Q_reg ( .D(g5637), .SI(n4606), .SE(n10229), .CLK(n10416), 
        .Q(test_so79), .QN(n10191) );
  SDFFX1 DFF_1303_Q_reg ( .D(g27276), .SI(test_si80), .SE(n10253), .CLK(n10440), .Q(g2429), .QN(n9834) );
  SDFFX1 DFF_1304_Q_reg ( .D(g27291), .SI(g2429), .SE(n10254), .CLK(n10441), 
        .Q(g2418), .QN(n9833) );
  SDFFX1 DFF_1305_Q_reg ( .D(g27307), .SI(g2418), .SE(n10254), .CLK(n10441), 
        .Q(g2421), .QN(n9832) );
  SDFFX1 DFF_1306_Q_reg ( .D(g27292), .SI(g2421), .SE(n10254), .CLK(n10441), 
        .Q(g2444), .QN(n9811) );
  SDFFX1 DFF_1307_Q_reg ( .D(g27308), .SI(g2444), .SE(n10254), .CLK(n10441), 
        .Q(g2433), .QN(n9810) );
  SDFFX1 DFF_1308_Q_reg ( .D(g27322), .SI(g2433), .SE(n10253), .CLK(n10440), 
        .Q(g2436), .QN(n9809) );
  SDFFX1 DFF_1309_Q_reg ( .D(g27309), .SI(g2436), .SE(n10253), .CLK(n10440), 
        .Q(g2459), .QN(n9556) );
  SDFFX1 DFF_1310_Q_reg ( .D(g27323), .SI(g2459), .SE(n10253), .CLK(n10440), 
        .Q(g2448), .QN(n9558) );
  SDFFX1 DFF_1311_Q_reg ( .D(g27334), .SI(g2448), .SE(n10253), .CLK(n10440), 
        .Q(g2451), .QN(n9557) );
  SDFFX1 DFF_1312_Q_reg ( .D(g27324), .SI(g2451), .SE(n10255), .CLK(n10442), 
        .Q(g2473), .QN(n9823) );
  SDFFX1 DFF_1313_Q_reg ( .D(g27335), .SI(g2473), .SE(n10255), .CLK(n10442), 
        .Q(g2463), .QN(n9822) );
  SDFFX1 DFF_1314_Q_reg ( .D(g27342), .SI(g2463), .SE(n10248), .CLK(n10435), 
        .Q(g2466), .QN(n9821) );
  SDFFX1 DFF_1315_Q_reg ( .D(g28763), .SI(g2466), .SE(n10248), .CLK(n10435), 
        .Q(g2483) );
  SDFFX1 DFF_1316_Q_reg ( .D(g28773), .SI(g2483), .SE(n10253), .CLK(n10440), 
        .Q(g2486) );
  SDFFX1 DFF_1317_Q_reg ( .D(g28782), .SI(g2486), .SE(n10253), .CLK(n10440), 
        .Q(test_so80) );
  SDFFX1 DFF_1318_Q_reg ( .D(g29213), .SI(test_si81), .SE(n10248), .CLK(n10435), .Q(g2492) );
  SDFFX1 DFF_1319_Q_reg ( .D(g29221), .SI(g2492), .SE(n10248), .CLK(n10435), 
        .Q(g2495) );
  SDFFX1 DFF_1320_Q_reg ( .D(g29226), .SI(g2495), .SE(n10249), .CLK(n10436), 
        .Q(g2498) );
  SDFFX1 DFF_1321_Q_reg ( .D(g28774), .SI(g2498), .SE(n10252), .CLK(n10439), 
        .Q(g2502), .QN(n9855) );
  SDFFX1 DFF_1322_Q_reg ( .D(g28783), .SI(g2502), .SE(n10252), .CLK(n10439), 
        .Q(g2503), .QN(n9845) );
  SDFFX1 DFF_1323_Q_reg ( .D(g28788), .SI(g2503), .SE(n10252), .CLK(n10439), 
        .Q(g2501), .QN(n9854) );
  SDFFX1 DFF_1324_Q_reg ( .D(g26817), .SI(g2501), .SE(n10252), .CLK(n10439), 
        .Q(g2504) );
  SDFFX1 DFF_1325_Q_reg ( .D(g26822), .SI(g2504), .SE(n10252), .CLK(n10439), 
        .Q(g2507) );
  SDFFX1 DFF_1326_Q_reg ( .D(g26825), .SI(g2507), .SE(n10252), .CLK(n10439), 
        .Q(g2510) );
  SDFFX1 DFF_1327_Q_reg ( .D(g26823), .SI(g2510), .SE(n10252), .CLK(n10439), 
        .Q(g2513) );
  SDFFX1 DFF_1328_Q_reg ( .D(g26826), .SI(g2513), .SE(n10252), .CLK(n10439), 
        .Q(g2516) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26827), .SI(g2516), .SE(n10252), .CLK(n10439), 
        .Q(g2519) );
  SDFFX1 DFF_1330_Q_reg ( .D(g27767), .SI(g2519), .SE(n10253), .CLK(n10440), 
        .Q(g2523), .QN(n9853) );
  SDFFX1 DFF_1331_Q_reg ( .D(g27769), .SI(g2523), .SE(n10253), .CLK(n10440), 
        .Q(g2524), .QN(n9844) );
  SDFFX1 DFF_1332_Q_reg ( .D(g27771), .SI(g2524), .SE(n10252), .CLK(n10439), 
        .Q(test_so81), .QN(n10208) );
  SDFFX1 DFF_1333_Q_reg ( .D(g29618), .SI(test_si82), .SE(n10248), .CLK(n10435), .Q(g2387), .QN(n9458) );
  SDFFX1 DFF_1334_Q_reg ( .D(g29621), .SI(g2387), .SE(n10248), .CLK(n10435), 
        .Q(g2388), .QN(n9446) );
  SDFFX1 DFF_1335_Q_reg ( .D(g29623), .SI(g2388), .SE(n10248), .CLK(n10435), 
        .Q(g2389), .QN(n9457) );
  SDFFX1 DFF_1336_Q_reg ( .D(g30707), .SI(g2389), .SE(n10248), .CLK(n10435), 
        .Q(g2390), .QN(n9456) );
  SDFFX1 DFF_1337_Q_reg ( .D(g30709), .SI(g2390), .SE(n10229), .CLK(n10416), 
        .Q(g2391), .QN(n9445) );
  SDFFX1 DFF_1338_Q_reg ( .D(g30566), .SI(g2391), .SE(n10229), .CLK(n10416), 
        .Q(g2392), .QN(n9455) );
  SDFFX1 DFF_1339_Q_reg ( .D(g30505), .SI(g2392), .SE(n10229), .CLK(n10416), 
        .Q(g2393), .QN(n9454) );
  SDFFX1 DFF_1340_Q_reg ( .D(g30341), .SI(g2393), .SE(n10229), .CLK(n10416), 
        .Q(g2394), .QN(n9444) );
  SDFFX1 DFF_1341_Q_reg ( .D(g30356), .SI(g2394), .SE(n10229), .CLK(n10416), 
        .Q(g2395), .QN(n9453) );
  SDFFX1 DFF_1342_Q_reg ( .D(g29182), .SI(g2395), .SE(n10256), .CLK(n10443), 
        .Q(g2397) );
  SDFFX1 DFF_1343_Q_reg ( .D(g29185), .SI(g2397), .SE(n10256), .CLK(n10443), 
        .Q(g2398) );
  SDFFX1 DFF_1344_Q_reg ( .D(g29187), .SI(g2398), .SE(n10256), .CLK(n10443), 
        .Q(g2396) );
  SDFFX1 DFF_1345_Q_reg ( .D(g26672), .SI(g2396), .SE(n10257), .CLK(n10444), 
        .Q(g2478), .QN(n9852) );
  SDFFX1 DFF_1346_Q_reg ( .D(g26676), .SI(g2478), .SE(n10257), .CLK(n10444), 
        .Q(g2479), .QN(n9843) );
  SDFFX1 DFF_1347_Q_reg ( .D(g26025), .SI(g2479), .SE(n10257), .CLK(n10444), 
        .Q(test_so82), .QN(n10217) );
  SDFFX1 DFF_1348_Q_reg ( .D(n4287), .SI(test_si83), .SE(n10257), .CLK(n10444), 
        .Q(g2525) );
  SDFFX1 DFF_1349_Q_reg ( .D(g2525), .SI(g2525), .SE(n10257), .CLK(n10444), 
        .Q(n7946), .QN(DFF_1349_n1) );
  SDFFX1 DFF_1350_Q_reg ( .D(n4563), .SI(n7946), .SE(n10257), .CLK(n10444), 
        .Q(g2527) );
  SDFFX1 DFF_1351_Q_reg ( .D(g2527), .SI(g2527), .SE(n10257), .CLK(n10444), 
        .Q(n7945), .QN(DFF_1351_n1) );
  SDFFX1 DFF_1352_Q_reg ( .D(n4555), .SI(n7945), .SE(n10257), .CLK(n10444), 
        .Q(g2529) );
  SDFFX1 DFF_1353_Q_reg ( .D(g2529), .SI(g2529), .SE(n10257), .CLK(n10444), 
        .Q(n7944), .QN(DFF_1353_n1) );
  SDFFX1 DFF_1354_Q_reg ( .D(n4325), .SI(n7944), .SE(n10257), .CLK(n10444), 
        .Q(g2355) );
  SDFFX1 DFF_1355_Q_reg ( .D(g2355), .SI(g2355), .SE(n10257), .CLK(n10444), 
        .Q(n7943), .QN(DFF_1355_n1) );
  SDFFX1 DFF_1356_Q_reg ( .D(n4389), .SI(n7943), .SE(n10257), .CLK(n10444), 
        .Q(g2357) );
  SDFFX1 DFF_1357_Q_reg ( .D(g2357), .SI(g2357), .SE(n10258), .CLK(n10445), 
        .Q(n7942), .QN(DFF_1357_n1) );
  SDFFX1 DFF_1358_Q_reg ( .D(n4319), .SI(n7942), .SE(n10258), .CLK(n10445), 
        .Q(g2359) );
  SDFFX1 DFF_1359_Q_reg ( .D(g2359), .SI(g2359), .SE(n10258), .CLK(n10445), 
        .Q(n7941), .QN(DFF_1359_n1) );
  SDFFX1 DFF_1360_Q_reg ( .D(n4373), .SI(n7941), .SE(n10258), .CLK(n10445), 
        .Q(g2361) );
  SDFFX1 DFF_1361_Q_reg ( .D(g2361), .SI(g2361), .SE(n10258), .CLK(n10445), 
        .Q(n7940), .QN(DFF_1361_n1) );
  SDFFX1 DFF_1362_Q_reg ( .D(n4377), .SI(n7940), .SE(n10258), .CLK(n10445), 
        .Q(test_so83) );
  SDFFX1 DFF_1363_Q_reg ( .D(test_so83), .SI(test_si84), .SE(n10258), .CLK(
        n10445), .Q(n7938), .QN(DFF_1363_n1) );
  SDFFX1 DFF_1364_Q_reg ( .D(g2878), .SI(n7938), .SE(n10345), .CLK(n10532), 
        .Q(g2365) );
  SDFFX1 DFF_1365_Q_reg ( .D(g2365), .SI(g2365), .SE(n10345), .CLK(n10532), 
        .Q(n7937), .QN(n4483) );
  SDFFX1 DFF_1366_Q_reg ( .D(n4285), .SI(n7937), .SE(n10345), .CLK(n10532), 
        .Q(g2374), .QN(n4487) );
  SDFFX1 DFF_1367_Q_reg ( .D(g30055), .SI(g2374), .SE(n10229), .CLK(n10416), 
        .Q(g2380) );
  SDFFX1 DFF_1378_Q_reg ( .D(n4275), .SI(g2380), .SE(n10229), .CLK(n10416), 
        .Q(n7936), .QN(DFF_1378_n1) );
  SDFFX1 DFF_1379_Q_reg ( .D(g2429), .SI(n7936), .SE(n10253), .CLK(n10440), 
        .Q(g2417) );
  SDFFX1 DFF_1380_Q_reg ( .D(g2417), .SI(g2417), .SE(n10253), .CLK(n10440), 
        .Q(g2424) );
  SDFFX1 DFF_1381_Q_reg ( .D(g2418), .SI(g2424), .SE(n10254), .CLK(n10441), 
        .Q(g2425) );
  SDFFX1 DFF_1382_Q_reg ( .D(g2425), .SI(g2425), .SE(n10254), .CLK(n10441), 
        .Q(g2426) );
  SDFFX1 DFF_1383_Q_reg ( .D(g2421), .SI(g2426), .SE(n10254), .CLK(n10441), 
        .Q(g2427) );
  SDFFX1 DFF_1384_Q_reg ( .D(g2427), .SI(g2427), .SE(n10254), .CLK(n10441), 
        .Q(g2428) );
  SDFFX1 DFF_1385_Q_reg ( .D(g2444), .SI(g2428), .SE(n10254), .CLK(n10441), 
        .Q(g2432) );
  SDFFX1 DFF_1386_Q_reg ( .D(g2432), .SI(g2432), .SE(n10254), .CLK(n10441), 
        .Q(g2439) );
  SDFFX1 DFF_1387_Q_reg ( .D(g2433), .SI(g2439), .SE(n10254), .CLK(n10441), 
        .Q(test_so84) );
  SDFFX1 DFF_1388_Q_reg ( .D(test_so84), .SI(test_si85), .SE(n10254), .CLK(
        n10441), .Q(g2441) );
  SDFFX1 DFF_1389_Q_reg ( .D(g2436), .SI(g2441), .SE(n10255), .CLK(n10442), 
        .Q(g2442) );
  SDFFX1 DFF_1390_Q_reg ( .D(g2442), .SI(g2442), .SE(n10255), .CLK(n10442), 
        .Q(g2443) );
  SDFFX1 DFF_1391_Q_reg ( .D(g2459), .SI(g2443), .SE(n10255), .CLK(n10442), 
        .Q(g2447) );
  SDFFX1 DFF_1392_Q_reg ( .D(g2447), .SI(g2447), .SE(n10255), .CLK(n10442), 
        .Q(g2454) );
  SDFFX1 DFF_1393_Q_reg ( .D(g2448), .SI(g2454), .SE(n10255), .CLK(n10442), 
        .Q(g2455) );
  SDFFX1 DFF_1394_Q_reg ( .D(g2455), .SI(g2455), .SE(n10255), .CLK(n10442), 
        .Q(g2456) );
  SDFFX1 DFF_1395_Q_reg ( .D(g2451), .SI(g2456), .SE(n10255), .CLK(n10442), 
        .Q(g2457) );
  SDFFX1 DFF_1396_Q_reg ( .D(g2457), .SI(g2457), .SE(n10255), .CLK(n10442), 
        .Q(g2458) );
  SDFFX1 DFF_1397_Q_reg ( .D(g2473), .SI(g2458), .SE(n10255), .CLK(n10442), 
        .Q(g2462) );
  SDFFX1 DFF_1398_Q_reg ( .D(g2462), .SI(g2462), .SE(n10255), .CLK(n10442), 
        .Q(g2469) );
  SDFFX1 DFF_1399_Q_reg ( .D(g2463), .SI(g2469), .SE(n10256), .CLK(n10443), 
        .Q(g2470) );
  SDFFX1 DFF_1400_Q_reg ( .D(g2470), .SI(g2470), .SE(n10256), .CLK(n10443), 
        .Q(g2471) );
  SDFFX1 DFF_1401_Q_reg ( .D(g2466), .SI(g2471), .SE(n10256), .CLK(n10443), 
        .Q(g2472) );
  SDFFX1 DFF_1402_Q_reg ( .D(g2472), .SI(g2472), .SE(n10256), .CLK(n10443), 
        .Q(test_so85) );
  SDFFX1 DFF_1403_Q_reg ( .D(n4598), .SI(test_si86), .SE(n10224), .CLK(n10411), 
        .Q(g5747) );
  SDFFX1 DFF_1404_Q_reg ( .D(g5747), .SI(g5747), .SE(n10224), .CLK(n10411), 
        .Q(g5796) );
  SDFFX1 DFF_1405_Q_reg ( .D(g5796), .SI(g5796), .SE(n10224), .CLK(n10411), 
        .Q(g2412) );
  SDFFX1 DFF_1406_Q_reg ( .D(n4598), .SI(g2412), .SE(n10224), .CLK(n10411), 
        .Q(g7302), .QN(n4314) );
  SDFFX1 DFF_1407_Q_reg ( .D(g7302), .SI(g7302), .SE(n10224), .CLK(n10411), 
        .Q(g7390), .QN(n4370) );
  SDFFX1 DFF_1408_Q_reg ( .D(g7390), .SI(g7390), .SE(n10224), .CLK(n10411), 
        .Q(g2624), .QN(n4299) );
  SDFFX1 DFF_1409_Q_reg ( .D(g21847), .SI(g2624), .SE(n10232), .CLK(n10419), 
        .Q(g2628), .QN(n10120) );
  SDFFX1 DFF_1410_Q_reg ( .D(g18780), .SI(g2628), .SE(n10232), .CLK(n10419), 
        .Q(g2631), .QN(n4352) );
  SDFFX1 DFF_1411_Q_reg ( .D(g18820), .SI(g2631), .SE(n10232), .CLK(n10419), 
        .Q(g2584), .QN(n4303) );
  SDFFX1 DFF_1412_Q_reg ( .D(n1669), .SI(g2584), .SE(n10251), .CLK(n10438), 
        .Q(g2587) );
  SDFFX1 DFF_1413_Q_reg ( .D(g2587), .SI(g2587), .SE(n10251), .CLK(n10438), 
        .Q(g2597) );
  SDFFX1 DFF_1414_Q_reg ( .D(g2597), .SI(g2597), .SE(n10251), .CLK(n10438), 
        .Q(g2598) );
  SDFFX1 DFF_1415_Q_reg ( .D(g2530), .SI(g2598), .SE(n10250), .CLK(n10437), 
        .Q(g2638) );
  SDFFX1 DFF_1416_Q_reg ( .D(g2638), .SI(g2638), .SE(n10250), .CLK(n10437), 
        .Q(g2643) );
  SDFFX1 DFF_1417_Q_reg ( .D(g2533), .SI(g2643), .SE(n10251), .CLK(n10438), 
        .Q(test_so86) );
  SDFFX1 DFF_1418_Q_reg ( .D(test_so86), .SI(test_si87), .SE(n10251), .CLK(
        n10438), .Q(g2645) );
  SDFFX1 DFF_1419_Q_reg ( .D(g2536), .SI(g2645), .SE(n10251), .CLK(n10438), 
        .Q(g2646) );
  SDFFX1 DFF_1420_Q_reg ( .D(g2646), .SI(g2646), .SE(n10251), .CLK(n10438), 
        .Q(g2647) );
  SDFFX1 DFF_1421_Q_reg ( .D(g2540), .SI(g2647), .SE(n10249), .CLK(n10436), 
        .Q(g2648) );
  SDFFX1 DFF_1422_Q_reg ( .D(g2648), .SI(g2648), .SE(n10249), .CLK(n10436), 
        .Q(g2639) );
  SDFFX1 DFF_1423_Q_reg ( .D(g2543), .SI(g2639), .SE(n10249), .CLK(n10436), 
        .Q(g2640) );
  SDFFX1 DFF_1424_Q_reg ( .D(g2640), .SI(g2640), .SE(n10249), .CLK(n10436), 
        .Q(g2641) );
  SDFFX1 DFF_1425_Q_reg ( .D(g2546), .SI(g2641), .SE(n10249), .CLK(n10436), 
        .Q(g2642) );
  SDFFX1 DFF_1426_Q_reg ( .D(g2642), .SI(g2642), .SE(n10249), .CLK(n10436), 
        .Q(g2564) );
  SDFFX1 DFF_1427_Q_reg ( .D(g2950), .SI(g2564), .SE(n10249), .CLK(n10436), 
        .Q(g8087), .QN(n4456) );
  SDFFX1 DFF_1428_Q_reg ( .D(g8087), .SI(g8087), .SE(n10250), .CLK(n10437), 
        .Q(g8167), .QN(n4455) );
  SDFFX1 DFF_1429_Q_reg ( .D(g8167), .SI(g8167), .SE(n10250), .CLK(n10437), 
        .Q(g2560), .QN(n4463) );
  SDFFX1 DFF_1430_Q_reg ( .D(g23114), .SI(g2560), .SE(n10252), .CLK(n10439), 
        .Q(g2561) );
  SDFFX1 DFF_1431_Q_reg ( .D(g23133), .SI(g2561), .SE(n10252), .CLK(n10439), 
        .Q(g2562) );
  SDFFX1 DFF_1432_Q_reg ( .D(g21970), .SI(g2562), .SE(n10253), .CLK(n10440), 
        .Q(test_so87) );
  SDFFX1 DFF_1433_Q_reg ( .D(g23407), .SI(test_si88), .SE(n10250), .CLK(n10437), .Q(g2530) );
  SDFFX1 DFF_1434_Q_reg ( .D(g23418), .SI(g2530), .SE(n10250), .CLK(n10437), 
        .Q(g2533) );
  SDFFX1 DFF_1435_Q_reg ( .D(g24209), .SI(g2533), .SE(n10250), .CLK(n10437), 
        .Q(g2536) );
  SDFFX1 DFF_1436_Q_reg ( .D(g24214), .SI(g2536), .SE(n10251), .CLK(n10438), 
        .Q(g2552) );
  SDFFX1 DFF_1437_Q_reg ( .D(g24226), .SI(g2552), .SE(n10251), .CLK(n10438), 
        .Q(g2553) );
  SDFFX1 DFF_1438_Q_reg ( .D(g24238), .SI(g2553), .SE(n10251), .CLK(n10438), 
        .Q(g2554) );
  SDFFX1 DFF_1439_Q_reg ( .D(g23132), .SI(g2554), .SE(n10249), .CLK(n10436), 
        .Q(g2555) );
  SDFFX1 DFF_1440_Q_reg ( .D(g23047), .SI(g2555), .SE(n10249), .CLK(n10436), 
        .Q(g2559) );
  SDFFX1 DFF_1441_Q_reg ( .D(g23076), .SI(g2559), .SE(n10249), .CLK(n10436), 
        .Q(g2539) );
  SDFFX1 DFF_1442_Q_reg ( .D(g24225), .SI(g2539), .SE(n10249), .CLK(n10436), 
        .Q(g2540) );
  SDFFX1 DFF_1443_Q_reg ( .D(g24237), .SI(g2540), .SE(n10250), .CLK(n10437), 
        .Q(g2543) );
  SDFFX1 DFF_1444_Q_reg ( .D(g24250), .SI(g2543), .SE(n10250), .CLK(n10437), 
        .Q(g2546) );
  SDFFX1 DFF_1445_Q_reg ( .D(n1647), .SI(g2546), .SE(n10250), .CLK(n10437), 
        .Q(g2602) );
  SDFFX1 DFF_1446_Q_reg ( .D(g2602), .SI(g2602), .SE(n10250), .CLK(n10437), 
        .Q(g2609) );
  SDFFX1 DFF_1447_Q_reg ( .D(g2609), .SI(g2609), .SE(n10250), .CLK(n10437), 
        .Q(test_so88) );
  SDFFX1 DFF_1448_Q_reg ( .D(g13175), .SI(test_si89), .SE(n10251), .CLK(n10438), .Q(g2617) );
  SDFFX1 DFF_1449_Q_reg ( .D(g2617), .SI(g2617), .SE(n10251), .CLK(n10438), 
        .Q(n7930) );
  SDFFX1 DFF_1450_Q_reg ( .D(g30072), .SI(n7930), .SE(n10331), .CLK(n10518), 
        .Q(n7929) );
  SDFFX1 DFF_1451_Q_reg ( .D(g13143), .SI(n7929), .SE(n10331), .CLK(n10518), 
        .Q(g2623) );
  SDFFX1 DFF_1452_Q_reg ( .D(g2623), .SI(g2623), .SE(n10332), .CLK(n10519), 
        .Q(g2574), .QN(n4543) );
  SDFFX1 DFF_1453_Q_reg ( .D(g13194), .SI(g2574), .SE(n10332), .CLK(n10519), 
        .Q(g2632) );
  SDFFX1 DFF_1454_Q_reg ( .D(g2632), .SI(g2632), .SE(n10332), .CLK(n10519), 
        .Q(g2633) );
  SDFFX1 DFF_1455_Q_reg ( .D(g27310), .SI(g2633), .SE(n10332), .CLK(n10519), 
        .Q(g2650), .QN(n9511) );
  SDFFX1 DFF_1456_Q_reg ( .D(g27325), .SI(g2650), .SE(n10332), .CLK(n10519), 
        .Q(g2651), .QN(n9513) );
  SDFFX1 DFF_1457_Q_reg ( .D(g27336), .SI(g2651), .SE(n10332), .CLK(n10519), 
        .Q(g2649), .QN(n9512) );
  SDFFX1 DFF_1458_Q_reg ( .D(g27326), .SI(g2649), .SE(n10332), .CLK(n10519), 
        .Q(g2653), .QN(n9523) );
  SDFFX1 DFF_1459_Q_reg ( .D(g27337), .SI(g2653), .SE(n10333), .CLK(n10520), 
        .Q(g2654), .QN(n9525) );
  SDFFX1 DFF_1460_Q_reg ( .D(g27343), .SI(g2654), .SE(n10332), .CLK(n10519), 
        .Q(g2652), .QN(n9524) );
  SDFFX1 DFF_1461_Q_reg ( .D(g27338), .SI(g2652), .SE(n10332), .CLK(n10519), 
        .Q(g2656), .QN(n9357) );
  SDFFX1 DFF_1462_Q_reg ( .D(g27344), .SI(g2656), .SE(n10332), .CLK(n10519), 
        .Q(test_so89) );
  SDFFX1 DFF_1463_Q_reg ( .D(g27347), .SI(test_si90), .SE(n10332), .CLK(n10519), .Q(g2655), .QN(n9358) );
  SDFFX1 DFF_1464_Q_reg ( .D(g27345), .SI(g2655), .SE(n10232), .CLK(n10419), 
        .Q(g2659), .QN(n9534) );
  SDFFX1 DFF_1465_Q_reg ( .D(g27348), .SI(g2659), .SE(n10333), .CLK(n10520), 
        .Q(g2660), .QN(n9536) );
  SDFFX1 DFF_1466_Q_reg ( .D(g27354), .SI(g2660), .SE(n10333), .CLK(n10520), 
        .Q(g2658), .QN(n9535) );
  SDFFX1 DFF_1467_Q_reg ( .D(g24527), .SI(g2658), .SE(n10333), .CLK(n10520), 
        .Q(g2661) );
  SDFFX1 DFF_1468_Q_reg ( .D(g24537), .SI(g2661), .SE(n10333), .CLK(n10520), 
        .Q(g2664) );
  SDFFX1 DFF_1469_Q_reg ( .D(g24547), .SI(g2664), .SE(n10333), .CLK(n10520), 
        .Q(g2667) );
  SDFFX1 DFF_1470_Q_reg ( .D(g24538), .SI(g2667), .SE(n10333), .CLK(n10520), 
        .Q(g2670) );
  SDFFX1 DFF_1471_Q_reg ( .D(g24548), .SI(g2670), .SE(n10333), .CLK(n10520), 
        .Q(g2673) );
  SDFFX1 DFF_1472_Q_reg ( .D(g24557), .SI(g2673), .SE(n10333), .CLK(n10520), 
        .Q(g2676) );
  SDFFX1 DFF_1473_Q_reg ( .D(g28364), .SI(g2676), .SE(n10333), .CLK(n10520), 
        .Q(g2688) );
  SDFFX1 DFF_1474_Q_reg ( .D(g28368), .SI(g2688), .SE(n10333), .CLK(n10520), 
        .Q(g2691) );
  SDFFX1 DFF_1475_Q_reg ( .D(g28371), .SI(g2691), .SE(n10232), .CLK(n10419), 
        .Q(g2694) );
  SDFFX1 DFF_1476_Q_reg ( .D(g28358), .SI(g2694), .SE(n10232), .CLK(n10419), 
        .Q(g2679) );
  SDFFX1 DFF_1477_Q_reg ( .D(g28363), .SI(g2679), .SE(n10232), .CLK(n10419), 
        .Q(test_so90) );
  SDFFX1 DFF_1478_Q_reg ( .D(g28367), .SI(test_si91), .SE(n10232), .CLK(n10419), .Q(g2685) );
  SDFFX1 DFF_1479_Q_reg ( .D(g26575), .SI(g2685), .SE(n10232), .CLK(n10419), 
        .Q(g2565) );
  SDFFX1 DFF_1480_Q_reg ( .D(g26596), .SI(g2565), .SE(n10232), .CLK(n10419), 
        .Q(g2568) );
  SDFFX1 DFF_1481_Q_reg ( .D(g26616), .SI(g2568), .SE(n10232), .CLK(n10419), 
        .Q(g2571) );
  SDFFX1 DFF_1482_Q_reg ( .D(g2574), .SI(g2571), .SE(n10332), .CLK(n10519), 
        .Q(g2580), .QN(n9672) );
  SDFFX1 DFF_1483_Q_reg ( .D(g22687), .SI(g2580), .SE(n10353), .CLK(n10540), 
        .Q(n7926) );
  SDFFX1 DFF_1492_Q_reg ( .D(g30061), .SI(n7926), .SE(n10353), .CLK(n10540), 
        .Q(g16437) );
  SDFFX1 DFF_1493_Q_reg ( .D(g16437), .SI(g16437), .SE(n10353), .CLK(n10540), 
        .Q(g2599), .QN(n9895) );
  SDFFX1 DFF_1494_Q_reg ( .D(DFF_1349_n1), .SI(g2599), .SE(n10353), .CLK(
        n10540), .Q(n7925) );
  SDFFX1 DFF_1495_Q_reg ( .D(DFF_1351_n1), .SI(n7925), .SE(n10353), .CLK(
        n10540), .Q(n7924) );
  SDFFX1 DFF_1496_Q_reg ( .D(DFF_1353_n1), .SI(n7924), .SE(n10353), .CLK(
        n10540), .Q(n7923) );
  SDFFX1 DFF_1497_Q_reg ( .D(DFF_1355_n1), .SI(n7923), .SE(n10354), .CLK(
        n10541), .Q(n7922) );
  SDFFX1 DFF_1498_Q_reg ( .D(DFF_1357_n1), .SI(n7922), .SE(n10354), .CLK(
        n10541), .Q(n7921) );
  SDFFX1 DFF_1499_Q_reg ( .D(DFF_1359_n1), .SI(n7921), .SE(n10354), .CLK(
        n10541), .Q(n7920) );
  SDFFX1 DFF_1500_Q_reg ( .D(DFF_1361_n1), .SI(n7920), .SE(n10354), .CLK(
        n10541), .Q(test_so91) );
  SDFFX1 DFF_1501_Q_reg ( .D(DFF_1363_n1), .SI(test_si92), .SE(n10258), .CLK(
        n10445), .Q(g2611) );
  SDFFX1 DFF_1502_Q_reg ( .D(g24092), .SI(g2611), .SE(n10229), .CLK(n10416), 
        .Q(g2612), .QN(n4490) );
  SDFFX1 DFF_1503_Q_reg ( .D(n4483), .SI(g2612), .SE(n10345), .CLK(n10532), 
        .Q(n7918) );
  SDFFX1 DFF_1505_Q_reg ( .D(g7425), .SI(g7425), .SE(n10345), .CLK(n10532), 
        .Q(g7487), .QN(n4356) );
  SDFFX1 DFF_1506_Q_reg ( .D(g7487), .SI(g7487), .SE(n10345), .CLK(n10532), 
        .Q(g2703), .QN(n4292) );
  SDFFX1 DFF_1507_Q_reg ( .D(g16718), .SI(g2703), .SE(n10345), .CLK(n10532), 
        .Q(g2704), .QN(n10156) );
  SDFFX1 DFF_1508_Q_reg ( .D(g20375), .SI(g2704), .SE(n10345), .CLK(n10532), 
        .Q(g2733), .QN(n4426) );
  SDFFX1 DFF_1509_Q_reg ( .D(g20789), .SI(g2733), .SE(n10345), .CLK(n10532), 
        .Q(g2714), .QN(n4398) );
  SDFFX1 DFF_1510_Q_reg ( .D(g21974), .SI(g2714), .SE(n10346), .CLK(n10533), 
        .Q(g2707), .QN(n4472) );
  SDFFX1 DFF_1511_Q_reg ( .D(g23348), .SI(g2707), .SE(n10346), .CLK(n10533), 
        .Q(g2727), .QN(n4419) );
  SDFFX1 DFF_1512_Q_reg ( .D(g24438), .SI(g2727), .SE(n10346), .CLK(n10533), 
        .Q(g2720), .QN(n4408) );
  SDFFX1 DFF_1513_Q_reg ( .D(g25197), .SI(g2720), .SE(n10346), .CLK(n10533), 
        .Q(g2734), .QN(n4397) );
  SDFFX1 DFF_1514_Q_reg ( .D(g26677), .SI(g2734), .SE(n10346), .CLK(n10533), 
        .Q(g2746), .QN(n4407) );
  SDFFX1 DFF_1515_Q_reg ( .D(g26795), .SI(g2746), .SE(n10346), .CLK(n10533), 
        .Q(test_so92), .QN(n10192) );
  SDFFX1 DFF_1516_Q_reg ( .D(g27243), .SI(test_si93), .SE(n10346), .CLK(n10533), .Q(g2753), .QN(n4471) );
  SDFFX1 DFF_1517_Q_reg ( .D(g27724), .SI(g2753), .SE(n10346), .CLK(n10533), 
        .Q(g2760), .QN(n4393) );
  SDFFX1 DFF_1518_Q_reg ( .D(g28328), .SI(g2760), .SE(n10346), .CLK(n10533), 
        .Q(g2766), .QN(n4415) );
  SDFFX1 DFF_1519_Q_reg ( .D(g20918), .SI(g2766), .SE(n10347), .CLK(n10534), 
        .Q(g2773), .QN(n9956) );
  SDFFX1 DFF_1520_Q_reg ( .D(g20939), .SI(g2773), .SE(n10347), .CLK(n10534), 
        .Q(g2774), .QN(n9955) );
  SDFFX1 DFF_1521_Q_reg ( .D(g20962), .SI(g2774), .SE(n10347), .CLK(n10534), 
        .Q(g2772), .QN(n10018) );
  SDFFX1 DFF_1522_Q_reg ( .D(g20940), .SI(g2772), .SE(n10347), .CLK(n10534), 
        .Q(g2776), .QN(n9954) );
  SDFFX1 DFF_1523_Q_reg ( .D(g20963), .SI(g2776), .SE(n10348), .CLK(n10535), 
        .Q(g2777), .QN(n9953) );
  SDFFX1 DFF_1524_Q_reg ( .D(g20981), .SI(g2777), .SE(n10348), .CLK(n10535), 
        .Q(g2775), .QN(n10017) );
  SDFFX1 DFF_1525_Q_reg ( .D(g20964), .SI(g2775), .SE(n10348), .CLK(n10535), 
        .Q(g2779), .QN(n9952) );
  SDFFX1 DFF_1526_Q_reg ( .D(g20982), .SI(g2779), .SE(n10348), .CLK(n10535), 
        .Q(g2780), .QN(n9951) );
  SDFFX1 DFF_1527_Q_reg ( .D(g21004), .SI(g2780), .SE(n10348), .CLK(n10535), 
        .Q(g2778), .QN(n10016) );
  SDFFX1 DFF_1528_Q_reg ( .D(g20983), .SI(g2778), .SE(n10348), .CLK(n10535), 
        .Q(g2782), .QN(n9950) );
  SDFFX1 DFF_1529_Q_reg ( .D(g21005), .SI(g2782), .SE(n10348), .CLK(n10535), 
        .Q(g2783), .QN(n9949) );
  SDFFX1 DFF_1530_Q_reg ( .D(g21025), .SI(g2783), .SE(n10348), .CLK(n10535), 
        .Q(test_so93), .QN(n10219) );
  SDFFX1 DFF_1531_Q_reg ( .D(g21006), .SI(test_si94), .SE(n10348), .CLK(n10535), .Q(g2785), .QN(n9948) );
  SDFFX1 DFF_1532_Q_reg ( .D(g21026), .SI(g2785), .SE(n10348), .CLK(n10535), 
        .Q(g2786), .QN(n9947) );
  SDFFX1 DFF_1533_Q_reg ( .D(g21043), .SI(g2786), .SE(n10348), .CLK(n10535), 
        .Q(g2784), .QN(n10015) );
  SDFFX1 DFF_1534_Q_reg ( .D(g21027), .SI(g2784), .SE(n10348), .CLK(n10535), 
        .Q(g2788), .QN(n9946) );
  SDFFX1 DFF_1535_Q_reg ( .D(g21044), .SI(g2788), .SE(n10349), .CLK(n10536), 
        .Q(g2789), .QN(n9945) );
  SDFFX1 DFF_1536_Q_reg ( .D(g21060), .SI(g2789), .SE(n10349), .CLK(n10536), 
        .Q(g2787), .QN(n10014) );
  SDFFX1 DFF_1537_Q_reg ( .D(g21045), .SI(g2787), .SE(n10349), .CLK(n10536), 
        .Q(g2791), .QN(n9944) );
  SDFFX1 DFF_1538_Q_reg ( .D(g21061), .SI(g2791), .SE(n10349), .CLK(n10536), 
        .Q(g2792), .QN(n9943) );
  SDFFX1 DFF_1539_Q_reg ( .D(g21073), .SI(g2792), .SE(n10349), .CLK(n10536), 
        .Q(g2790), .QN(n10013) );
  SDFFX1 DFF_1540_Q_reg ( .D(g21062), .SI(g2790), .SE(n10349), .CLK(n10536), 
        .Q(g2794), .QN(n9942) );
  SDFFX1 DFF_1541_Q_reg ( .D(g21074), .SI(g2794), .SE(n10349), .CLK(n10536), 
        .Q(g2795), .QN(n9941) );
  SDFFX1 DFF_1542_Q_reg ( .D(g21081), .SI(g2795), .SE(n10349), .CLK(n10536), 
        .Q(g2793), .QN(n10012) );
  SDFFX1 DFF_1543_Q_reg ( .D(g21075), .SI(g2793), .SE(n10349), .CLK(n10536), 
        .Q(g2797), .QN(n9940) );
  SDFFX1 DFF_1544_Q_reg ( .D(g21082), .SI(g2797), .SE(n10349), .CLK(n10536), 
        .Q(g2798), .QN(n9939) );
  SDFFX1 DFF_1545_Q_reg ( .D(g21094), .SI(g2798), .SE(n10349), .CLK(n10536), 
        .Q(test_so94), .QN(n10218) );
  SDFFX1 DFF_1546_Q_reg ( .D(g20919), .SI(test_si95), .SE(n10347), .CLK(n10534), .Q(g2800), .QN(n9938) );
  SDFFX1 DFF_1547_Q_reg ( .D(g20941), .SI(g2800), .SE(n10347), .CLK(n10534), 
        .Q(g2801), .QN(n9937) );
  SDFFX1 DFF_1548_Q_reg ( .D(g20965), .SI(g2801), .SE(n10347), .CLK(n10534), 
        .Q(g2799), .QN(n10011) );
  SDFFX1 DFF_1549_Q_reg ( .D(g21007), .SI(g2799), .SE(n10347), .CLK(n10534), 
        .Q(g2803), .QN(n9748) );
  SDFFX1 DFF_1550_Q_reg ( .D(g21028), .SI(g2803), .SE(n10347), .CLK(n10534), 
        .Q(g2804), .QN(n9740) );
  SDFFX1 DFF_1551_Q_reg ( .D(g21046), .SI(g2804), .SE(n10347), .CLK(n10534), 
        .Q(g2802), .QN(n9803) );
  SDFFX1 DFF_1552_Q_reg ( .D(g21029), .SI(g2802), .SE(n10347), .CLK(n10534), 
        .Q(g2806), .QN(n9747) );
  SDFFX1 DFF_1553_Q_reg ( .D(g21047), .SI(g2806), .SE(n10347), .CLK(n10534), 
        .Q(g2807), .QN(n9739) );
  SDFFX1 DFF_1554_Q_reg ( .D(g21063), .SI(g2807), .SE(n10232), .CLK(n10419), 
        .Q(g2805), .QN(n9802) );
  SDFFX1 DFF_1555_Q_reg ( .D(g25272), .SI(g2805), .SE(n10349), .CLK(n10536), 
        .Q(g2809) );
  SDFFX1 DFF_1556_Q_reg ( .D(g25280), .SI(g2809), .SE(n10350), .CLK(n10537), 
        .Q(g2810) );
  SDFFX1 DFF_1557_Q_reg ( .D(g25288), .SI(g2810), .SE(n10230), .CLK(n10417), 
        .Q(g2808) );
  SDFFX1 DFF_1558_Q_reg ( .D(g22269), .SI(g2808), .SE(n10346), .CLK(n10533), 
        .Q(g2812) );
  SDFFX1 DFF_1559_Q_reg ( .D(g22284), .SI(g2812), .SE(n10346), .CLK(n10533), 
        .Q(g2813) );
  SDFFX1 DFF_1560_Q_reg ( .D(g22299), .SI(g2813), .SE(n10346), .CLK(n10533), 
        .Q(test_so95) );
  SDFFX1 DFF_1561_Q_reg ( .D(g20877), .SI(test_si96), .SE(n10224), .CLK(n10411), .Q(n7913) );
  SDFFX1 DFF_1562_Q_reg ( .D(g20884), .SI(n7913), .SE(n10224), .CLK(n10411), 
        .Q(n7912) );
  SDFFX1 DFF_1563_Q_reg ( .D(n4263), .SI(n7912), .SE(n10224), .CLK(n10411), 
        .Q(n4598), .QN(n10165) );
  SDFFX1 DFF_1564_Q_reg ( .D(n4269), .SI(n4598), .SE(n10342), .CLK(n10529), 
        .Q(g3043) );
  SDFFX1 DFF_1565_Q_reg ( .D(n4268), .SI(g3043), .SE(n10342), .CLK(n10529), 
        .Q(g3044) );
  SDFFX1 DFF_1566_Q_reg ( .D(n4267), .SI(g3044), .SE(n10342), .CLK(n10529), 
        .Q(g3045) );
  SDFFX1 DFF_1567_Q_reg ( .D(n4266), .SI(g3045), .SE(n10343), .CLK(n10530), 
        .Q(g3046) );
  SDFFX1 DFF_1568_Q_reg ( .D(n4265), .SI(g3046), .SE(n10343), .CLK(n10530), 
        .Q(g3047) );
  SDFFX1 DFF_1569_Q_reg ( .D(n4272), .SI(g3047), .SE(n10343), .CLK(n10530), 
        .Q(g3048) );
  SDFFX1 DFF_1570_Q_reg ( .D(n4271), .SI(g3048), .SE(n10343), .CLK(n10530), 
        .Q(g3049) );
  SDFFX1 DFF_1571_Q_reg ( .D(n4270), .SI(g3049), .SE(n10343), .CLK(n10530), 
        .Q(g3050) );
  SDFFX1 DFF_1572_Q_reg ( .D(n4259), .SI(g3050), .SE(n10344), .CLK(n10531), 
        .Q(g3051) );
  SDFFX1 DFF_1573_Q_reg ( .D(n4236), .SI(g3051), .SE(n10344), .CLK(n10531), 
        .Q(g3052) );
  SDFFX1 DFF_1574_Q_reg ( .D(n4239), .SI(g3052), .SE(n10344), .CLK(n10531), 
        .Q(g3053) );
  SDFFX1 DFF_1575_Q_reg ( .D(n4237), .SI(g3053), .SE(n10344), .CLK(n10531), 
        .Q(test_so96) );
  SDFFX1 DFF_1576_Q_reg ( .D(n4234), .SI(test_si97), .SE(n10340), .CLK(n10527), 
        .Q(g3056) );
  SDFFX1 DFF_1577_Q_reg ( .D(n4233), .SI(g3056), .SE(n10340), .CLK(n10527), 
        .Q(g3057) );
  SDFFX1 DFF_1578_Q_reg ( .D(n4238), .SI(g3057), .SE(n10341), .CLK(n10528), 
        .Q(g3058) );
  SDFFX1 DFF_1579_Q_reg ( .D(n4235), .SI(g3058), .SE(n10341), .CLK(n10528), 
        .Q(g3059) );
  SDFFX1 DFF_1580_Q_reg ( .D(n4240), .SI(g3059), .SE(n10341), .CLK(n10528), 
        .Q(g3060) );
  SDFFX1 DFF_1581_Q_reg ( .D(n4232), .SI(g3060), .SE(n10341), .CLK(n10528), 
        .Q(g3061) );
  SDFFX1 DFF_1582_Q_reg ( .D(n4245), .SI(g3061), .SE(n10341), .CLK(n10528), 
        .Q(g3062) );
  SDFFX1 DFF_1583_Q_reg ( .D(n4248), .SI(g3062), .SE(n10341), .CLK(n10528), 
        .Q(g3063) );
  SDFFX1 DFF_1584_Q_reg ( .D(n4246), .SI(g3063), .SE(n10341), .CLK(n10528), 
        .Q(g3064) );
  SDFFX1 DFF_1585_Q_reg ( .D(n4243), .SI(g3064), .SE(n10341), .CLK(n10528), 
        .Q(g3065) );
  SDFFX1 DFF_1586_Q_reg ( .D(n4242), .SI(g3065), .SE(n10234), .CLK(n10421), 
        .Q(g3066) );
  SDFFX1 DFF_1587_Q_reg ( .D(n4247), .SI(g3066), .SE(n10234), .CLK(n10421), 
        .Q(g3067) );
  SDFFX1 DFF_1588_Q_reg ( .D(n4244), .SI(g3067), .SE(n10234), .CLK(n10421), 
        .Q(g3068) );
  SDFFX1 DFF_1589_Q_reg ( .D(n4249), .SI(g3068), .SE(n10234), .CLK(n10421), 
        .Q(g3069) );
  SDFFX1 DFF_1590_Q_reg ( .D(n4241), .SI(g3069), .SE(n10234), .CLK(n10421), 
        .Q(test_so97) );
  SDFFX1 DFF_1591_Q_reg ( .D(n4254), .SI(test_si98), .SE(n10230), .CLK(n10417), 
        .Q(g3071) );
  SDFFX1 DFF_1592_Q_reg ( .D(n4257), .SI(g3071), .SE(n10230), .CLK(n10417), 
        .Q(g3072) );
  SDFFX1 DFF_1593_Q_reg ( .D(n4255), .SI(g3072), .SE(n10230), .CLK(n10417), 
        .Q(g3073) );
  SDFFX1 DFF_1594_Q_reg ( .D(n4252), .SI(g3073), .SE(n10230), .CLK(n10417), 
        .Q(g3074) );
  SDFFX1 DFF_1595_Q_reg ( .D(n4251), .SI(g3074), .SE(n10230), .CLK(n10417), 
        .Q(g3075) );
  SDFFX1 DFF_1596_Q_reg ( .D(n4256), .SI(g3075), .SE(n10230), .CLK(n10417), 
        .Q(g3076) );
  SDFFX1 DFF_1597_Q_reg ( .D(n4253), .SI(g3076), .SE(n10230), .CLK(n10417), 
        .Q(g3077) );
  SDFFX1 DFF_1598_Q_reg ( .D(n4258), .SI(g3077), .SE(n10230), .CLK(n10417), 
        .Q(g3078) );
  SDFFX1 DFF_1599_Q_reg ( .D(n4250), .SI(g3078), .SE(n10230), .CLK(n10417), 
        .Q(g2997) );
  SDFFX1 DFF_1600_Q_reg ( .D(g25265), .SI(g2997), .SE(n10230), .CLK(n10417), 
        .Q(g2993), .QN(n10166) );
  SDFFX1 DFF_1601_Q_reg ( .D(g26048), .SI(g2993), .SE(n10230), .CLK(n10417), 
        .Q(n7909), .QN(n18262) );
  SDFFX1 DFF_1602_Q_reg ( .D(g23330), .SI(n7909), .SE(n10231), .CLK(n10418), 
        .Q(g3006), .QN(n10164) );
  SDFFX1 DFF_1603_Q_reg ( .D(g24445), .SI(g3006), .SE(n10231), .CLK(n10418), 
        .Q(g3002), .QN(n9352) );
  SDFFX1 DFF_1604_Q_reg ( .D(g25191), .SI(g3002), .SE(n10231), .CLK(n10418), 
        .Q(g3013), .QN(n10163) );
  SDFFX1 DFF_1605_Q_reg ( .D(g26031), .SI(g3013), .SE(n10231), .CLK(n10418), 
        .Q(test_so98), .QN(n10197) );
  SDFFX1 DFF_1606_Q_reg ( .D(g26786), .SI(test_si99), .SE(n10231), .CLK(n10418), .Q(g3024), .QN(n9351) );
  SDFFX1 DFF_1607_Q_reg ( .D(n4262), .SI(g3024), .SE(n10231), .CLK(n10418), 
        .Q(g3018), .QN(n4481) );
  SDFFX1 DFF_1608_Q_reg ( .D(g23359), .SI(g3018), .SE(n10231), .CLK(n10418), 
        .Q(g3028), .QN(n4350) );
  SDFFX1 DFF_1609_Q_reg ( .D(g24446), .SI(g3028), .SE(n10231), .CLK(n10418), 
        .Q(g3036), .QN(n4480) );
  SDFFX1 DFF_1610_Q_reg ( .D(g25202), .SI(g3036), .SE(n10231), .CLK(n10418), 
        .Q(g3032), .QN(n10157) );
  SDFFX1 DFF_1611_Q_reg ( .D(g3234), .SI(g3032), .SE(n10231), .CLK(n10418), 
        .Q(g5388) );
  SDFFX1 DFF_1612_Q_reg ( .D(g5388), .SI(g5388), .SE(n10231), .CLK(n10418), 
        .Q(n7907), .QN(DFF_1612_n1) );
  SDFFX1 DFF_1613_Q_reg ( .D(g16496), .SI(n7907), .SE(n10231), .CLK(n10418), 
        .Q(g2987), .QN(n4365) );
  SDFFX1 DFF_1614_Q_reg ( .D(g16824), .SI(g2987), .SE(n10342), .CLK(n10529), 
        .Q(g8275), .QN(n10144) );
  SDFFX1 DFF_1615_Q_reg ( .D(g16844), .SI(g8275), .SE(n10342), .CLK(n10529), 
        .Q(g8274), .QN(n10146) );
  SDFFX1 DFF_1616_Q_reg ( .D(g16853), .SI(g8274), .SE(n10342), .CLK(n10529), 
        .Q(g8273), .QN(n18265) );
  SDFFX1 DFF_1617_Q_reg ( .D(g16860), .SI(g8273), .SE(n10343), .CLK(n10530), 
        .Q(g8272), .QN(n18259) );
  SDFFX1 DFF_1618_Q_reg ( .D(g16803), .SI(g8272), .SE(n10343), .CLK(n10530), 
        .Q(g8268), .QN(n18264) );
  SDFFX1 DFF_1619_Q_reg ( .D(g16835), .SI(g8268), .SE(n10343), .CLK(n10530), 
        .Q(g8269), .QN(n10147) );
  SDFFX1 DFF_1620_Q_reg ( .D(g16851), .SI(g8269), .SE(n10343), .CLK(n10530), 
        .Q(test_so99), .QN(n10205) );
  SDFFX1 DFF_1621_Q_reg ( .D(g16857), .SI(test_si100), .SE(n10343), .CLK(
        n10530), .Q(g8271) );
  SDFFX1 DFF_1622_Q_reg ( .D(g16866), .SI(g8271), .SE(n10235), .CLK(n10422), 
        .Q(g3083), .QN(n10149) );
  SDFFX1 DFF_1623_Q_reg ( .D(n4261), .SI(g3083), .SE(n10344), .CLK(n10531), 
        .Q(g8267) );
  SDFFX1 DFF_1624_Q_reg ( .D(N995), .SI(g8267), .SE(n10235), .CLK(n10422), .Q(
        n4577) );
  SDFFX1 DFF_1625_Q_reg ( .D(g16845), .SI(n4577), .SE(n10235), .CLK(n10422), 
        .Q(g8266), .QN(n18267) );
  SDFFX1 DFF_1626_Q_reg ( .D(g16854), .SI(g8266), .SE(n10344), .CLK(n10531), 
        .Q(g8265), .QN(n18260) );
  SDFFX1 DFF_1627_Q_reg ( .D(g16861), .SI(g8265), .SE(n10344), .CLK(n10531), 
        .Q(g8264), .QN(n10127) );
  SDFFX1 DFF_1628_Q_reg ( .D(g16880), .SI(g8264), .SE(n10344), .CLK(n10531), 
        .Q(g8262), .QN(n18266) );
  SDFFX1 DFF_1629_Q_reg ( .D(g18755), .SI(g8262), .SE(n10344), .CLK(n10531), 
        .Q(g8263), .QN(n10128) );
  SDFFX1 DFF_1630_Q_reg ( .D(g18804), .SI(g8263), .SE(n10344), .CLK(n10531), 
        .Q(g8260), .QN(n10124) );
  SDFFX1 DFF_1631_Q_reg ( .D(g18837), .SI(g8260), .SE(n10344), .CLK(n10531), 
        .Q(g8261) );
  SDFFX1 DFF_1632_Q_reg ( .D(g18868), .SI(g8261), .SE(n10344), .CLK(n10531), 
        .Q(g8259), .QN(n10126) );
  SDFFX1 DFF_1633_Q_reg ( .D(g18907), .SI(g8259), .SE(n10345), .CLK(n10532), 
        .Q(g2990), .QN(n10151) );
  SDFFX1 DFF_1634_Q_reg ( .D(N690), .SI(g2990), .SE(n10235), .CLK(n10422), .Q(
        n4578) );
  SDFFX1 DFF_1635_Q_reg ( .D(n4260), .SI(n4578), .SE(n10353), .CLK(n10540), 
        .Q(test_so100) );
  SDFFX1 DFF_454_Q_reg ( .D(n4598), .SI(n8040), .SE(n10280), .CLK(n10467), .Q(
        g6677), .QN(n4309) );
  SDFFX1 DFF_804_Q_reg ( .D(n4598), .SI(test_si49), .SE(n10224), .CLK(n10411), 
        .Q(g6979), .QN(n4308) );
  SDFFX1 DFF_1154_Q_reg ( .D(n4598), .SI(n7960), .SE(n10238), .CLK(n10425), 
        .Q(g7229), .QN(n4307) );
  SDFFX1 DFF_1504_Q_reg ( .D(n4598), .SI(n7918), .SE(n10345), .CLK(n10532), 
        .Q(g7425), .QN(n4306) );
  SDFFX1 DFF_1300_Q_reg ( .D(g5555), .SI(g5555), .SE(n10228), .CLK(n10415), 
        .Q(g7264), .QN(n4524) );
  SDFFX1 DFF_950_Q_reg ( .D(g5511), .SI(g5511), .SE(n10314), .CLK(n10501), .Q(
        g7014), .QN(n4525) );
  SDFFX1 DFF_951_Q_reg ( .D(g7014), .SI(g7014), .SE(n10314), .CLK(n10501), .Q(
        n4618), .QN(n4511) );
  SDFFX1 DFF_1301_Q_reg ( .D(g7264), .SI(g7264), .SE(n10229), .CLK(n10416), 
        .Q(n4606), .QN(n4509) );
  SDFFX1 DFF_250_Q_reg ( .D(g5437), .SI(g5437), .SE(n10261), .CLK(n10448), .Q(
        g6447), .QN(n4499) );
  SDFFX1 DFF_249_Q_reg ( .D(g2950), .SI(g181), .SE(n10261), .CLK(n10448), .Q(
        g5437), .QN(n4520) );
  NOR2X0 Trojan1 ( .IN1(n2459), .IN2(n2309), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(n2237), .IN2(n2279), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(n2381), .IN2(n2207), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(n2542), .IN2(n2489), .QN(Tj_OUT4) );
  AND4X1 Trojan1234 ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  OR2X1 Trojan5 ( .IN1(n3260), .IN2(n342), .Q(Tj_OUT5) );
  OR2X1 Trojan6 ( .IN1(n336), .IN2(n339), .Q(Tj_OUT6) );
  OR2X1 Trojan7 ( .IN1(n3374), .IN2(n3293), .Q(Tj_OUT7) );
  OR2X1 Trojan8 ( .IN1(n3334), .IN2(n41), .Q(Tj_OUT8) );
  AND4X1 Trojan5678 ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  AND2X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .Q(Tj_Trigger)
         );
  OR2X1 Trojan_Payload_1 ( .IN1(Tj_Trigger), .IN2(n4149), .Q(n4149_Tj_Payload)
         );
  OR2X1 Trojan_Payload_2 ( .IN1(Tj_Trigger), .IN2(n680), .Q(n4161_Tj_Payload)
         );
  OR2X1 Trojan_Payload_3 ( .IN1(Tj_Trigger), .IN2(n1027), .Q(n4160_Tj_Payload)
         );
  OR2X1 Trojan_Payload_4 ( .IN1(Tj_Trigger), .IN2(n4122), .Q(n4122_Tj_Payload)
         );
  NBUFFX2 U10085 ( .INP(n10398), .Z(n10224) );
  NBUFFX2 U10086 ( .INP(n10398), .Z(n10225) );
  NBUFFX2 U10087 ( .INP(n10396), .Z(n10231) );
  NBUFFX2 U10088 ( .INP(n10358), .Z(n10344) );
  NBUFFX2 U10089 ( .INP(n10396), .Z(n10230) );
  NBUFFX2 U10090 ( .INP(n10356), .Z(n10349) );
  NBUFFX2 U10091 ( .INP(n10357), .Z(n10348) );
  NBUFFX2 U10092 ( .INP(n10357), .Z(n10347) );
  NBUFFX2 U10093 ( .INP(n10357), .Z(n10346) );
  NBUFFX2 U10094 ( .INP(n10362), .Z(n10332) );
  NBUFFX2 U10095 ( .INP(n10389), .Z(n10250) );
  NBUFFX2 U10096 ( .INP(n10389), .Z(n10251) );
  NBUFFX2 U10097 ( .INP(n10395), .Z(n10232) );
  NBUFFX2 U10098 ( .INP(n10387), .Z(n10257) );
  NBUFFX2 U10099 ( .INP(n10389), .Z(n10252) );
  NBUFFX2 U10100 ( .INP(n10390), .Z(n10249) );
  NBUFFX2 U10101 ( .INP(n10388), .Z(n10255) );
  NBUFFX2 U10102 ( .INP(n10388), .Z(n10254) );
  NBUFFX2 U10103 ( .INP(n10388), .Z(n10253) );
  NBUFFX2 U10104 ( .INP(n10395), .Z(n10234) );
  NBUFFX2 U10105 ( .INP(n10390), .Z(n10247) );
  NBUFFX2 U10106 ( .INP(n10390), .Z(n10248) );
  NBUFFX2 U10107 ( .INP(n10387), .Z(n10256) );
  NBUFFX2 U10108 ( .INP(n10391), .Z(n10246) );
  NBUFFX2 U10109 ( .INP(n10391), .Z(n10245) );
  NBUFFX2 U10110 ( .INP(n10391), .Z(n10244) );
  NBUFFX2 U10111 ( .INP(n10396), .Z(n10229) );
  NBUFFX2 U10112 ( .INP(n10392), .Z(n10243) );
  NBUFFX2 U10113 ( .INP(n10359), .Z(n10340) );
  NBUFFX2 U10114 ( .INP(n10360), .Z(n10339) );
  NBUFFX2 U10115 ( .INP(n10360), .Z(n10338) );
  NBUFFX2 U10116 ( .INP(n10361), .Z(n10336) );
  NBUFFX2 U10117 ( .INP(n10361), .Z(n10335) );
  NBUFFX2 U10118 ( .INP(n10361), .Z(n10334) );
  NBUFFX2 U10119 ( .INP(n10362), .Z(n10333) );
  NBUFFX2 U10120 ( .INP(n10362), .Z(n10331) );
  NBUFFX2 U10121 ( .INP(n10363), .Z(n10330) );
  NBUFFX2 U10122 ( .INP(n10363), .Z(n10329) );
  NBUFFX2 U10123 ( .INP(n10363), .Z(n10328) );
  NBUFFX2 U10124 ( .INP(n10364), .Z(n10327) );
  NBUFFX2 U10125 ( .INP(n10364), .Z(n10326) );
  NBUFFX2 U10126 ( .INP(n10364), .Z(n10325) );
  NBUFFX2 U10127 ( .INP(n10360), .Z(n10337) );
  NBUFFX2 U10128 ( .INP(n10365), .Z(n10324) );
  NBUFFX2 U10129 ( .INP(n10365), .Z(n10323) );
  NBUFFX2 U10130 ( .INP(n10366), .Z(n10320) );
  NBUFFX2 U10131 ( .INP(n10366), .Z(n10321) );
  NBUFFX2 U10132 ( .INP(n10368), .Z(n10313) );
  NBUFFX2 U10133 ( .INP(n10367), .Z(n10318) );
  NBUFFX2 U10134 ( .INP(n10366), .Z(n10319) );
  NBUFFX2 U10135 ( .INP(n10365), .Z(n10322) );
  NBUFFX2 U10136 ( .INP(n10368), .Z(n10314) );
  NBUFFX2 U10137 ( .INP(n10367), .Z(n10317) );
  NBUFFX2 U10138 ( .INP(n10367), .Z(n10316) );
  NBUFFX2 U10139 ( .INP(n10368), .Z(n10315) );
  NBUFFX2 U10140 ( .INP(n10369), .Z(n10312) );
  NBUFFX2 U10141 ( .INP(n10369), .Z(n10311) );
  NBUFFX2 U10142 ( .INP(n10369), .Z(n10310) );
  NBUFFX2 U10143 ( .INP(n10370), .Z(n10309) );
  NBUFFX2 U10144 ( .INP(n10370), .Z(n10308) );
  NBUFFX2 U10145 ( .INP(n10370), .Z(n10307) );
  NBUFFX2 U10146 ( .INP(n10371), .Z(n10306) );
  NBUFFX2 U10147 ( .INP(n10371), .Z(n10305) );
  NBUFFX2 U10148 ( .INP(n10372), .Z(n10303) );
  NBUFFX2 U10149 ( .INP(n10371), .Z(n10304) );
  NBUFFX2 U10150 ( .INP(n10372), .Z(n10302) );
  NBUFFX2 U10151 ( .INP(n10372), .Z(n10301) );
  NBUFFX2 U10152 ( .INP(n10373), .Z(n10300) );
  NBUFFX2 U10153 ( .INP(n10373), .Z(n10299) );
  NBUFFX2 U10154 ( .INP(n10373), .Z(n10298) );
  NBUFFX2 U10155 ( .INP(n10374), .Z(n10297) );
  NBUFFX2 U10156 ( .INP(n10375), .Z(n10293) );
  NBUFFX2 U10157 ( .INP(n10375), .Z(n10294) );
  NBUFFX2 U10158 ( .INP(n10377), .Z(n10287) );
  NBUFFX2 U10159 ( .INP(n10375), .Z(n10292) );
  NBUFFX2 U10160 ( .INP(n10376), .Z(n10291) );
  NBUFFX2 U10161 ( .INP(n10374), .Z(n10296) );
  NBUFFX2 U10162 ( .INP(n10374), .Z(n10295) );
  NBUFFX2 U10163 ( .INP(n10377), .Z(n10288) );
  NBUFFX2 U10164 ( .INP(n10376), .Z(n10290) );
  NBUFFX2 U10165 ( .INP(n10376), .Z(n10289) );
  NBUFFX2 U10166 ( .INP(n10377), .Z(n10286) );
  NBUFFX2 U10167 ( .INP(n10378), .Z(n10285) );
  NBUFFX2 U10168 ( .INP(n10378), .Z(n10284) );
  NBUFFX2 U10169 ( .INP(n10378), .Z(n10283) );
  NBUFFX2 U10170 ( .INP(n10379), .Z(n10282) );
  NBUFFX2 U10171 ( .INP(n10379), .Z(n10281) );
  NBUFFX2 U10172 ( .INP(n10358), .Z(n10343) );
  NBUFFX2 U10173 ( .INP(n10380), .Z(n10279) );
  NBUFFX2 U10174 ( .INP(n10380), .Z(n10278) );
  NBUFFX2 U10175 ( .INP(n10380), .Z(n10277) );
  NBUFFX2 U10176 ( .INP(n10381), .Z(n10276) );
  NBUFFX2 U10177 ( .INP(n10381), .Z(n10275) );
  NBUFFX2 U10178 ( .INP(n10381), .Z(n10274) );
  NBUFFX2 U10179 ( .INP(n10382), .Z(n10273) );
  NBUFFX2 U10180 ( .INP(n10382), .Z(n10272) );
  NBUFFX2 U10181 ( .INP(n10379), .Z(n10280) );
  NBUFFX2 U10182 ( .INP(n10387), .Z(n10258) );
  NBUFFX2 U10183 ( .INP(n10359), .Z(n10342) );
  NBUFFX2 U10184 ( .INP(n10359), .Z(n10341) );
  NBUFFX2 U10185 ( .INP(n10382), .Z(n10271) );
  NBUFFX2 U10186 ( .INP(n10383), .Z(n10268) );
  NBUFFX2 U10187 ( .INP(n10384), .Z(n10267) );
  NBUFFX2 U10188 ( .INP(n10386), .Z(n10260) );
  NBUFFX2 U10189 ( .INP(n10384), .Z(n10266) );
  NBUFFX2 U10190 ( .INP(n10383), .Z(n10270) );
  NBUFFX2 U10191 ( .INP(n10383), .Z(n10269) );
  NBUFFX2 U10192 ( .INP(n10385), .Z(n10262) );
  NBUFFX2 U10193 ( .INP(n10386), .Z(n10261) );
  NBUFFX2 U10194 ( .INP(n10386), .Z(n10259) );
  NBUFFX2 U10195 ( .INP(n10385), .Z(n10263) );
  NBUFFX2 U10196 ( .INP(n10384), .Z(n10265) );
  NBUFFX2 U10197 ( .INP(n10385), .Z(n10264) );
  NBUFFX2 U10198 ( .INP(n10394), .Z(n10237) );
  NBUFFX2 U10199 ( .INP(n10394), .Z(n10235) );
  NBUFFX2 U10200 ( .INP(n10394), .Z(n10236) );
  NBUFFX2 U10201 ( .INP(n10355), .Z(n10353) );
  NBUFFX2 U10202 ( .INP(n10355), .Z(n10352) );
  NBUFFX2 U10203 ( .INP(n10356), .Z(n10351) );
  NBUFFX2 U10204 ( .INP(n10356), .Z(n10350) );
  NBUFFX2 U10205 ( .INP(n10358), .Z(n10345) );
  NBUFFX2 U10206 ( .INP(n10392), .Z(n10242) );
  NBUFFX2 U10207 ( .INP(n10392), .Z(n10241) );
  NBUFFX2 U10208 ( .INP(n10393), .Z(n10240) );
  NBUFFX2 U10209 ( .INP(n10393), .Z(n10239) );
  NBUFFX2 U10210 ( .INP(n10393), .Z(n10238) );
  NBUFFX2 U10211 ( .INP(n10397), .Z(n10226) );
  NBUFFX2 U10212 ( .INP(n10395), .Z(n10233) );
  NBUFFX2 U10213 ( .INP(n10397), .Z(n10228) );
  NBUFFX2 U10214 ( .INP(n10397), .Z(n10227) );
  NBUFFX2 U10215 ( .INP(n10585), .Z(n10411) );
  NBUFFX2 U10216 ( .INP(n10585), .Z(n10412) );
  NBUFFX2 U10217 ( .INP(n10583), .Z(n10418) );
  NBUFFX2 U10218 ( .INP(n10545), .Z(n10531) );
  NBUFFX2 U10219 ( .INP(n10583), .Z(n10417) );
  NBUFFX2 U10220 ( .INP(n10543), .Z(n10536) );
  NBUFFX2 U10221 ( .INP(n10544), .Z(n10535) );
  NBUFFX2 U10222 ( .INP(n10544), .Z(n10534) );
  NBUFFX2 U10223 ( .INP(n10544), .Z(n10533) );
  NBUFFX2 U10224 ( .INP(n10549), .Z(n10519) );
  NBUFFX2 U10225 ( .INP(n10576), .Z(n10437) );
  NBUFFX2 U10226 ( .INP(n10576), .Z(n10438) );
  NBUFFX2 U10227 ( .INP(n10582), .Z(n10419) );
  NBUFFX2 U10228 ( .INP(n10574), .Z(n10444) );
  NBUFFX2 U10229 ( .INP(n10576), .Z(n10439) );
  NBUFFX2 U10230 ( .INP(n10577), .Z(n10436) );
  NBUFFX2 U10231 ( .INP(n10575), .Z(n10442) );
  NBUFFX2 U10232 ( .INP(n10575), .Z(n10441) );
  NBUFFX2 U10233 ( .INP(n10575), .Z(n10440) );
  NBUFFX2 U10234 ( .INP(n10582), .Z(n10421) );
  NBUFFX2 U10235 ( .INP(n10577), .Z(n10434) );
  NBUFFX2 U10236 ( .INP(n10577), .Z(n10435) );
  NBUFFX2 U10237 ( .INP(n10574), .Z(n10443) );
  NBUFFX2 U10238 ( .INP(n10578), .Z(n10433) );
  NBUFFX2 U10239 ( .INP(n10578), .Z(n10432) );
  NBUFFX2 U10240 ( .INP(n10578), .Z(n10431) );
  NBUFFX2 U10241 ( .INP(n10583), .Z(n10416) );
  NBUFFX2 U10242 ( .INP(n10579), .Z(n10430) );
  NBUFFX2 U10243 ( .INP(n10546), .Z(n10527) );
  NBUFFX2 U10244 ( .INP(n10547), .Z(n10526) );
  NBUFFX2 U10245 ( .INP(n10547), .Z(n10525) );
  NBUFFX2 U10246 ( .INP(n10548), .Z(n10523) );
  NBUFFX2 U10247 ( .INP(n10548), .Z(n10522) );
  NBUFFX2 U10248 ( .INP(n10548), .Z(n10521) );
  NBUFFX2 U10249 ( .INP(n10549), .Z(n10520) );
  NBUFFX2 U10250 ( .INP(n10549), .Z(n10518) );
  NBUFFX2 U10251 ( .INP(n10550), .Z(n10517) );
  NBUFFX2 U10252 ( .INP(n10550), .Z(n10516) );
  NBUFFX2 U10253 ( .INP(n10550), .Z(n10515) );
  NBUFFX2 U10254 ( .INP(n10551), .Z(n10514) );
  NBUFFX2 U10255 ( .INP(n10551), .Z(n10513) );
  NBUFFX2 U10256 ( .INP(n10551), .Z(n10512) );
  NBUFFX2 U10257 ( .INP(n10547), .Z(n10524) );
  NBUFFX2 U10258 ( .INP(n10552), .Z(n10511) );
  NBUFFX2 U10259 ( .INP(n10552), .Z(n10510) );
  NBUFFX2 U10260 ( .INP(n10553), .Z(n10507) );
  NBUFFX2 U10261 ( .INP(n10553), .Z(n10508) );
  NBUFFX2 U10262 ( .INP(n10555), .Z(n10500) );
  NBUFFX2 U10263 ( .INP(n10554), .Z(n10505) );
  NBUFFX2 U10264 ( .INP(n10553), .Z(n10506) );
  NBUFFX2 U10265 ( .INP(n10552), .Z(n10509) );
  NBUFFX2 U10266 ( .INP(n10555), .Z(n10501) );
  NBUFFX2 U10267 ( .INP(n10554), .Z(n10504) );
  NBUFFX2 U10268 ( .INP(n10554), .Z(n10503) );
  NBUFFX2 U10269 ( .INP(n10555), .Z(n10502) );
  NBUFFX2 U10270 ( .INP(n10556), .Z(n10499) );
  NBUFFX2 U10271 ( .INP(n10556), .Z(n10498) );
  NBUFFX2 U10272 ( .INP(n10556), .Z(n10497) );
  NBUFFX2 U10273 ( .INP(n10557), .Z(n10496) );
  NBUFFX2 U10274 ( .INP(n10557), .Z(n10495) );
  NBUFFX2 U10275 ( .INP(n10557), .Z(n10494) );
  NBUFFX2 U10276 ( .INP(n10558), .Z(n10493) );
  NBUFFX2 U10277 ( .INP(n10558), .Z(n10492) );
  NBUFFX2 U10278 ( .INP(n10559), .Z(n10490) );
  NBUFFX2 U10279 ( .INP(n10558), .Z(n10491) );
  NBUFFX2 U10280 ( .INP(n10559), .Z(n10489) );
  NBUFFX2 U10281 ( .INP(n10559), .Z(n10488) );
  NBUFFX2 U10282 ( .INP(n10560), .Z(n10487) );
  NBUFFX2 U10283 ( .INP(n10560), .Z(n10486) );
  NBUFFX2 U10284 ( .INP(n10560), .Z(n10485) );
  NBUFFX2 U10285 ( .INP(n10561), .Z(n10484) );
  NBUFFX2 U10286 ( .INP(n10562), .Z(n10480) );
  NBUFFX2 U10287 ( .INP(n10562), .Z(n10481) );
  NBUFFX2 U10288 ( .INP(n10564), .Z(n10474) );
  NBUFFX2 U10289 ( .INP(n10562), .Z(n10479) );
  NBUFFX2 U10290 ( .INP(n10563), .Z(n10478) );
  NBUFFX2 U10291 ( .INP(n10561), .Z(n10483) );
  NBUFFX2 U10292 ( .INP(n10561), .Z(n10482) );
  NBUFFX2 U10293 ( .INP(n10564), .Z(n10475) );
  NBUFFX2 U10294 ( .INP(n10563), .Z(n10477) );
  NBUFFX2 U10295 ( .INP(n10563), .Z(n10476) );
  NBUFFX2 U10296 ( .INP(n10564), .Z(n10473) );
  NBUFFX2 U10297 ( .INP(n10565), .Z(n10472) );
  NBUFFX2 U10298 ( .INP(n10565), .Z(n10471) );
  NBUFFX2 U10299 ( .INP(n10565), .Z(n10470) );
  NBUFFX2 U10300 ( .INP(n10566), .Z(n10469) );
  NBUFFX2 U10301 ( .INP(n10566), .Z(n10468) );
  NBUFFX2 U10302 ( .INP(n10545), .Z(n10530) );
  NBUFFX2 U10303 ( .INP(n10567), .Z(n10466) );
  NBUFFX2 U10304 ( .INP(n10567), .Z(n10465) );
  NBUFFX2 U10305 ( .INP(n10567), .Z(n10464) );
  NBUFFX2 U10306 ( .INP(n10568), .Z(n10463) );
  NBUFFX2 U10307 ( .INP(n10568), .Z(n10462) );
  NBUFFX2 U10308 ( .INP(n10568), .Z(n10461) );
  NBUFFX2 U10309 ( .INP(n10569), .Z(n10460) );
  NBUFFX2 U10310 ( .INP(n10569), .Z(n10459) );
  NBUFFX2 U10311 ( .INP(n10566), .Z(n10467) );
  NBUFFX2 U10312 ( .INP(n10574), .Z(n10445) );
  NBUFFX2 U10313 ( .INP(n10546), .Z(n10529) );
  NBUFFX2 U10314 ( .INP(n10546), .Z(n10528) );
  NBUFFX2 U10315 ( .INP(n10569), .Z(n10458) );
  NBUFFX2 U10316 ( .INP(n10570), .Z(n10455) );
  NBUFFX2 U10317 ( .INP(n10571), .Z(n10454) );
  NBUFFX2 U10318 ( .INP(n10573), .Z(n10447) );
  NBUFFX2 U10319 ( .INP(n10571), .Z(n10453) );
  NBUFFX2 U10320 ( .INP(n10570), .Z(n10457) );
  NBUFFX2 U10321 ( .INP(n10570), .Z(n10456) );
  NBUFFX2 U10322 ( .INP(n10572), .Z(n10449) );
  NBUFFX2 U10323 ( .INP(n10573), .Z(n10448) );
  NBUFFX2 U10324 ( .INP(n10573), .Z(n10446) );
  NBUFFX2 U10325 ( .INP(n10572), .Z(n10450) );
  NBUFFX2 U10326 ( .INP(n10571), .Z(n10452) );
  NBUFFX2 U10327 ( .INP(n10572), .Z(n10451) );
  NBUFFX2 U10328 ( .INP(n10581), .Z(n10424) );
  NBUFFX2 U10329 ( .INP(n10581), .Z(n10422) );
  NBUFFX2 U10330 ( .INP(n10581), .Z(n10423) );
  NBUFFX2 U10331 ( .INP(n10542), .Z(n10540) );
  NBUFFX2 U10332 ( .INP(n10542), .Z(n10539) );
  NBUFFX2 U10333 ( .INP(n10543), .Z(n10538) );
  NBUFFX2 U10334 ( .INP(n10543), .Z(n10537) );
  NBUFFX2 U10335 ( .INP(n10545), .Z(n10532) );
  NBUFFX2 U10336 ( .INP(n10579), .Z(n10429) );
  NBUFFX2 U10337 ( .INP(n10579), .Z(n10428) );
  NBUFFX2 U10338 ( .INP(n10580), .Z(n10427) );
  NBUFFX2 U10339 ( .INP(n10580), .Z(n10426) );
  NBUFFX2 U10340 ( .INP(n10580), .Z(n10425) );
  NBUFFX2 U10341 ( .INP(n10584), .Z(n10413) );
  NBUFFX2 U10342 ( .INP(n10582), .Z(n10420) );
  NBUFFX2 U10343 ( .INP(n10584), .Z(n10415) );
  NBUFFX2 U10344 ( .INP(n10584), .Z(n10414) );
  NBUFFX2 U10345 ( .INP(n10355), .Z(n10354) );
  NBUFFX2 U10346 ( .INP(n10542), .Z(n10541) );
  NBUFFX2 U10347 ( .INP(n10594), .Z(n10544) );
  NBUFFX2 U10348 ( .INP(n10407), .Z(n10357) );
  NBUFFX2 U10349 ( .INP(n10594), .Z(n10542) );
  NBUFFX2 U10350 ( .INP(n10407), .Z(n10355) );
  NBUFFX2 U10351 ( .INP(n10594), .Z(n10543) );
  NBUFFX2 U10352 ( .INP(n10407), .Z(n10356) );
  NBUFFX2 U10353 ( .INP(n10594), .Z(n10545) );
  NBUFFX2 U10354 ( .INP(n10407), .Z(n10358) );
  NBUFFX2 U10355 ( .INP(n10587), .Z(n10576) );
  NBUFFX2 U10356 ( .INP(n10400), .Z(n10389) );
  NBUFFX2 U10357 ( .INP(n10588), .Z(n10575) );
  NBUFFX2 U10358 ( .INP(n10401), .Z(n10388) );
  NBUFFX2 U10359 ( .INP(n10587), .Z(n10577) );
  NBUFFX2 U10360 ( .INP(n10400), .Z(n10390) );
  NBUFFX2 U10361 ( .INP(n10587), .Z(n10578) );
  NBUFFX2 U10362 ( .INP(n10400), .Z(n10391) );
  NBUFFX2 U10363 ( .INP(n10586), .Z(n10583) );
  NBUFFX2 U10364 ( .INP(n10399), .Z(n10396) );
  NBUFFX2 U10365 ( .INP(n10593), .Z(n10548) );
  NBUFFX2 U10366 ( .INP(n10406), .Z(n10361) );
  NBUFFX2 U10367 ( .INP(n10593), .Z(n10549) );
  NBUFFX2 U10368 ( .INP(n10406), .Z(n10362) );
  NBUFFX2 U10369 ( .INP(n10593), .Z(n10550) );
  NBUFFX2 U10370 ( .INP(n10406), .Z(n10363) );
  NBUFFX2 U10371 ( .INP(n10592), .Z(n10551) );
  NBUFFX2 U10372 ( .INP(n10405), .Z(n10364) );
  NBUFFX2 U10373 ( .INP(n10593), .Z(n10547) );
  NBUFFX2 U10374 ( .INP(n10406), .Z(n10360) );
  NBUFFX2 U10375 ( .INP(n10592), .Z(n10553) );
  NBUFFX2 U10376 ( .INP(n10405), .Z(n10366) );
  NBUFFX2 U10377 ( .INP(n10592), .Z(n10552) );
  NBUFFX2 U10378 ( .INP(n10405), .Z(n10365) );
  NBUFFX2 U10379 ( .INP(n10592), .Z(n10554) );
  NBUFFX2 U10380 ( .INP(n10405), .Z(n10367) );
  NBUFFX2 U10381 ( .INP(n10592), .Z(n10555) );
  NBUFFX2 U10382 ( .INP(n10405), .Z(n10368) );
  NBUFFX2 U10383 ( .INP(n10591), .Z(n10556) );
  NBUFFX2 U10384 ( .INP(n10404), .Z(n10369) );
  NBUFFX2 U10385 ( .INP(n10591), .Z(n10557) );
  NBUFFX2 U10386 ( .INP(n10404), .Z(n10370) );
  NBUFFX2 U10387 ( .INP(n10591), .Z(n10558) );
  NBUFFX2 U10388 ( .INP(n10404), .Z(n10371) );
  NBUFFX2 U10389 ( .INP(n10591), .Z(n10559) );
  NBUFFX2 U10390 ( .INP(n10404), .Z(n10372) );
  NBUFFX2 U10391 ( .INP(n10591), .Z(n10560) );
  NBUFFX2 U10392 ( .INP(n10404), .Z(n10373) );
  NBUFFX2 U10393 ( .INP(n10590), .Z(n10562) );
  NBUFFX2 U10394 ( .INP(n10403), .Z(n10375) );
  NBUFFX2 U10395 ( .INP(n10590), .Z(n10561) );
  NBUFFX2 U10396 ( .INP(n10403), .Z(n10374) );
  NBUFFX2 U10397 ( .INP(n10590), .Z(n10563) );
  NBUFFX2 U10398 ( .INP(n10403), .Z(n10376) );
  NBUFFX2 U10399 ( .INP(n10590), .Z(n10564) );
  NBUFFX2 U10400 ( .INP(n10403), .Z(n10377) );
  NBUFFX2 U10401 ( .INP(n10590), .Z(n10565) );
  NBUFFX2 U10402 ( .INP(n10403), .Z(n10378) );
  NBUFFX2 U10403 ( .INP(n10589), .Z(n10567) );
  NBUFFX2 U10404 ( .INP(n10402), .Z(n10380) );
  NBUFFX2 U10405 ( .INP(n10589), .Z(n10568) );
  NBUFFX2 U10406 ( .INP(n10402), .Z(n10381) );
  NBUFFX2 U10407 ( .INP(n10589), .Z(n10566) );
  NBUFFX2 U10408 ( .INP(n10402), .Z(n10379) );
  NBUFFX2 U10409 ( .INP(n10588), .Z(n10574) );
  NBUFFX2 U10410 ( .INP(n10401), .Z(n10387) );
  NBUFFX2 U10411 ( .INP(n10593), .Z(n10546) );
  NBUFFX2 U10412 ( .INP(n10406), .Z(n10359) );
  NBUFFX2 U10413 ( .INP(n10589), .Z(n10569) );
  NBUFFX2 U10414 ( .INP(n10402), .Z(n10382) );
  NBUFFX2 U10415 ( .INP(n10589), .Z(n10570) );
  NBUFFX2 U10416 ( .INP(n10402), .Z(n10383) );
  NBUFFX2 U10417 ( .INP(n10588), .Z(n10573) );
  NBUFFX2 U10418 ( .INP(n10401), .Z(n10386) );
  NBUFFX2 U10419 ( .INP(n10588), .Z(n10571) );
  NBUFFX2 U10420 ( .INP(n10401), .Z(n10384) );
  NBUFFX2 U10421 ( .INP(n10588), .Z(n10572) );
  NBUFFX2 U10422 ( .INP(n10401), .Z(n10385) );
  NBUFFX2 U10423 ( .INP(n10586), .Z(n10581) );
  NBUFFX2 U10424 ( .INP(n10399), .Z(n10394) );
  NBUFFX2 U10425 ( .INP(n10587), .Z(n10579) );
  NBUFFX2 U10426 ( .INP(n10400), .Z(n10392) );
  NBUFFX2 U10427 ( .INP(n10587), .Z(n10580) );
  NBUFFX2 U10428 ( .INP(n10400), .Z(n10393) );
  NBUFFX2 U10429 ( .INP(n10586), .Z(n10582) );
  NBUFFX2 U10430 ( .INP(n10399), .Z(n10395) );
  NBUFFX2 U10431 ( .INP(n10586), .Z(n10584) );
  NBUFFX2 U10432 ( .INP(n10399), .Z(n10397) );
  NBUFFX2 U10433 ( .INP(n10586), .Z(n10585) );
  NBUFFX2 U10434 ( .INP(n10399), .Z(n10398) );
  NBUFFX2 U10435 ( .INP(n10410), .Z(n10399) );
  NBUFFX2 U10436 ( .INP(n10410), .Z(n10400) );
  NBUFFX2 U10437 ( .INP(n10410), .Z(n10401) );
  NBUFFX2 U10438 ( .INP(n10409), .Z(n10402) );
  NBUFFX2 U10439 ( .INP(n10409), .Z(n10403) );
  NBUFFX2 U10440 ( .INP(n10409), .Z(n10404) );
  NBUFFX2 U10441 ( .INP(n10408), .Z(n10405) );
  NBUFFX2 U10442 ( .INP(n10408), .Z(n10406) );
  NBUFFX2 U10443 ( .INP(n10408), .Z(n10407) );
  NBUFFX2 U10444 ( .INP(test_se), .Z(n10408) );
  NBUFFX2 U10445 ( .INP(test_se), .Z(n10409) );
  NBUFFX2 U10446 ( .INP(test_se), .Z(n10410) );
  NBUFFX2 U10447 ( .INP(n10597), .Z(n10586) );
  NBUFFX2 U10448 ( .INP(n10597), .Z(n10587) );
  NBUFFX2 U10449 ( .INP(n10597), .Z(n10588) );
  NBUFFX2 U10450 ( .INP(n10596), .Z(n10589) );
  NBUFFX2 U10451 ( .INP(n10596), .Z(n10590) );
  NBUFFX2 U10452 ( .INP(n10596), .Z(n10591) );
  NBUFFX2 U10453 ( .INP(n10595), .Z(n10592) );
  NBUFFX2 U10454 ( .INP(n10595), .Z(n10593) );
  NBUFFX2 U10455 ( .INP(n10595), .Z(n10594) );
  NBUFFX2 U10456 ( .INP(CK), .Z(n10595) );
  NBUFFX2 U10457 ( .INP(CK), .Z(n10596) );
  NBUFFX2 U10458 ( .INP(CK), .Z(n10597) );
  INVX0 U10459 ( .INP(n10598), .ZN(n984) );
  INVX0 U10460 ( .INP(g27380), .ZN(n97) );
  INVX0 U10461 ( .INP(n10599), .ZN(n962) );
  INVX0 U10462 ( .INP(n10600), .ZN(n791) );
  INVX0 U10463 ( .INP(n10601), .ZN(n634) );
  INVX0 U10464 ( .INP(n10602), .ZN(n632) );
  INVX0 U10465 ( .INP(n10603), .ZN(n610) );
  INVX0 U10466 ( .INP(n10604), .ZN(n4521) );
  AND2X1 U10467 ( .IN1(n3692), .IN2(test_so15), .Q(n10604) );
  OR2X1 U10468 ( .IN1(n10605), .IN2(n10606), .Q(n4281) );
  INVX0 U10469 ( .INP(n10607), .ZN(n10606) );
  OR2X1 U10470 ( .IN1(n10608), .IN2(n10150), .Q(n10607) );
  AND2X1 U10471 ( .IN1(n10150), .IN2(n10608), .Q(n10605) );
  AND2X1 U10472 ( .IN1(n10609), .IN2(n10610), .Q(n4280) );
  INVX0 U10473 ( .INP(n10611), .ZN(n10610) );
  AND2X1 U10474 ( .IN1(n10612), .IN2(n10148), .Q(n10611) );
  OR2X1 U10475 ( .IN1(n10148), .IN2(n10612), .Q(n10609) );
  OR2X1 U10476 ( .IN1(n10613), .IN2(n4351), .Q(n4279) );
  AND2X1 U10477 ( .IN1(DFF_18_n1), .IN2(g8021), .Q(n10613) );
  AND2X1 U10478 ( .IN1(n10614), .IN2(n10615), .Q(n4278) );
  OR2X1 U10479 ( .IN1(n10616), .IN2(n10617), .Q(n10615) );
  OR2X1 U10480 ( .IN1(n10618), .IN2(n10619), .Q(n10617) );
  OR2X1 U10481 ( .IN1(n10620), .IN2(n10621), .Q(n10619) );
  OR2X1 U10482 ( .IN1(n10622), .IN2(n10623), .Q(n10621) );
  OR2X1 U10483 ( .IN1(n10624), .IN2(n10625), .Q(n10623) );
  AND2X1 U10484 ( .IN1(n10626), .IN2(g88), .Q(n10625) );
  AND2X1 U10485 ( .IN1(n10184), .IN2(n10627), .Q(n10624) );
  OR2X1 U10486 ( .IN1(n10628), .IN2(n10629), .Q(n10622) );
  AND2X1 U10487 ( .IN1(n10630), .IN2(g70), .Q(n10629) );
  AND2X1 U10488 ( .IN1(n10167), .IN2(n10631), .Q(n10628) );
  OR2X1 U10489 ( .IN1(n10632), .IN2(n10633), .Q(n10620) );
  AND2X1 U10490 ( .IN1(n10634), .IN2(g61), .Q(n10633) );
  AND2X1 U10491 ( .IN1(n10176), .IN2(n10635), .Q(n10632) );
  OR2X1 U10492 ( .IN1(n10636), .IN2(n10637), .Q(n10618) );
  OR2X1 U10493 ( .IN1(n10638), .IN2(n10639), .Q(n10637) );
  OR2X1 U10494 ( .IN1(n10640), .IN2(n10641), .Q(n10639) );
  AND2X1 U10495 ( .IN1(n10642), .IN2(g65), .Q(n10641) );
  AND2X1 U10496 ( .IN1(n9888), .IN2(n10643), .Q(n10640) );
  OR2X1 U10497 ( .IN1(n10644), .IN2(n10645), .Q(n10638) );
  AND2X1 U10498 ( .IN1(n10646), .IN2(g52), .Q(n10645) );
  AND2X1 U10499 ( .IN1(n9356), .IN2(n10647), .Q(n10644) );
  OR2X1 U10500 ( .IN1(n10648), .IN2(n10649), .Q(n10636) );
  AND2X1 U10501 ( .IN1(n10650), .IN2(g56), .Q(n10649) );
  AND2X1 U10502 ( .IN1(n9510), .IN2(n10651), .Q(n10648) );
  OR2X1 U10503 ( .IN1(n10652), .IN2(n10653), .Q(n10616) );
  OR2X1 U10504 ( .IN1(n10654), .IN2(n10655), .Q(n10653) );
  OR2X1 U10505 ( .IN1(n10656), .IN2(n10657), .Q(n10655) );
  OR2X1 U10506 ( .IN1(n10658), .IN2(n10659), .Q(n10657) );
  AND2X1 U10507 ( .IN1(n4513), .IN2(g92), .Q(n10659) );
  AND2X1 U10508 ( .IN1(n9891), .IN2(n10660), .Q(n10658) );
  OR2X1 U10509 ( .IN1(n10661), .IN2(n10662), .Q(n10656) );
  AND2X1 U10510 ( .IN1(n10663), .IN2(g83), .Q(n10662) );
  AND2X1 U10511 ( .IN1(n9890), .IN2(n10664), .Q(n10661) );
  OR2X1 U10512 ( .IN1(n10665), .IN2(n10666), .Q(n10654) );
  AND2X1 U10513 ( .IN1(n10667), .IN2(g74), .Q(n10666) );
  AND2X1 U10514 ( .IN1(n9889), .IN2(n10668), .Q(n10665) );
  OR2X1 U10515 ( .IN1(n10669), .IN2(n10670), .Q(n10652) );
  OR2X1 U10516 ( .IN1(n10671), .IN2(n10672), .Q(n10670) );
  AND2X1 U10517 ( .IN1(n10673), .IN2(n10674), .Q(n10669) );
  OR2X1 U10518 ( .IN1(n10675), .IN2(n10199), .Q(n10674) );
  OR2X1 U10519 ( .IN1(test_so15), .IN2(n10676), .Q(n10673) );
  OR2X1 U10520 ( .IN1(n10677), .IN2(n10678), .Q(n10614) );
  AND2X1 U10521 ( .IN1(n10679), .IN2(n10680), .Q(n4277) );
  OR2X1 U10522 ( .IN1(n10681), .IN2(n10682), .Q(n10680) );
  OR2X1 U10523 ( .IN1(n10683), .IN2(n10684), .Q(n10682) );
  OR2X1 U10524 ( .IN1(n10685), .IN2(n10686), .Q(n10684) );
  OR2X1 U10525 ( .IN1(n10687), .IN2(n10688), .Q(n10686) );
  OR2X1 U10526 ( .IN1(n10689), .IN2(n10690), .Q(n10688) );
  AND2X1 U10527 ( .IN1(n10691), .IN2(g767), .Q(n10690) );
  AND2X1 U10528 ( .IN1(n10171), .IN2(n10692), .Q(n10689) );
  OR2X1 U10529 ( .IN1(n10693), .IN2(n10694), .Q(n10687) );
  AND2X1 U10530 ( .IN1(n10695), .IN2(g758), .Q(n10694) );
  AND2X1 U10531 ( .IN1(n10170), .IN2(n10696), .Q(n10693) );
  OR2X1 U10532 ( .IN1(n10697), .IN2(n10698), .Q(n10685) );
  AND2X1 U10533 ( .IN1(n10699), .IN2(g776), .Q(n10698) );
  AND2X1 U10534 ( .IN1(n10172), .IN2(n10700), .Q(n10697) );
  OR2X1 U10535 ( .IN1(n10701), .IN2(n10702), .Q(n10683) );
  OR2X1 U10536 ( .IN1(n10703), .IN2(n10704), .Q(n10702) );
  OR2X1 U10537 ( .IN1(n10705), .IN2(n10706), .Q(n10704) );
  AND2X1 U10538 ( .IN1(n10707), .IN2(g753), .Q(n10706) );
  AND2X1 U10539 ( .IN1(n9884), .IN2(n10708), .Q(n10705) );
  OR2X1 U10540 ( .IN1(n10709), .IN2(n10710), .Q(n10703) );
  AND2X1 U10541 ( .IN1(n10711), .IN2(g740), .Q(n10710) );
  AND2X1 U10542 ( .IN1(n9355), .IN2(n10712), .Q(n10709) );
  OR2X1 U10543 ( .IN1(n10713), .IN2(n10714), .Q(n10701) );
  AND2X1 U10544 ( .IN1(n10715), .IN2(g780), .Q(n10714) );
  AND2X1 U10545 ( .IN1(n9887), .IN2(n10716), .Q(n10713) );
  OR2X1 U10546 ( .IN1(n10717), .IN2(n10718), .Q(n10681) );
  OR2X1 U10547 ( .IN1(n10719), .IN2(n10720), .Q(n10718) );
  OR2X1 U10548 ( .IN1(n10721), .IN2(n10722), .Q(n10720) );
  OR2X1 U10549 ( .IN1(n10723), .IN2(n10724), .Q(n10722) );
  AND2X1 U10550 ( .IN1(n10725), .IN2(g762), .Q(n10724) );
  AND2X1 U10551 ( .IN1(n9885), .IN2(n10726), .Q(n10723) );
  OR2X1 U10552 ( .IN1(n10727), .IN2(n10728), .Q(n10721) );
  AND2X1 U10553 ( .IN1(n10729), .IN2(g744), .Q(n10728) );
  AND2X1 U10554 ( .IN1(n9509), .IN2(n10730), .Q(n10727) );
  OR2X1 U10555 ( .IN1(n10731), .IN2(n10732), .Q(n10719) );
  AND2X1 U10556 ( .IN1(n10733), .IN2(g771), .Q(n10732) );
  AND2X1 U10557 ( .IN1(n9886), .IN2(n10734), .Q(n10731) );
  OR2X1 U10558 ( .IN1(n10735), .IN2(n10736), .Q(n10717) );
  OR2X1 U10559 ( .IN1(n10737), .IN2(n10672), .Q(n10736) );
  AND2X1 U10560 ( .IN1(n10738), .IN2(n10739), .Q(n10735) );
  OR2X1 U10561 ( .IN1(n10740), .IN2(n10195), .Q(n10739) );
  OR2X1 U10562 ( .IN1(test_so36), .IN2(n10741), .Q(n10738) );
  OR2X1 U10563 ( .IN1(n2542), .IN2(n10742), .Q(n10679) );
  AND2X1 U10564 ( .IN1(n10743), .IN2(n10744), .Q(n4276) );
  OR2X1 U10565 ( .IN1(n10745), .IN2(n10746), .Q(n10744) );
  OR2X1 U10566 ( .IN1(n10747), .IN2(n10748), .Q(n10746) );
  OR2X1 U10567 ( .IN1(n10749), .IN2(n10750), .Q(n10748) );
  OR2X1 U10568 ( .IN1(n10751), .IN2(n10752), .Q(n10750) );
  OR2X1 U10569 ( .IN1(n10753), .IN2(n10754), .Q(n10752) );
  AND2X1 U10570 ( .IN1(n10755), .IN2(g1462), .Q(n10754) );
  AND2X1 U10571 ( .IN1(n10185), .IN2(n10756), .Q(n10753) );
  OR2X1 U10572 ( .IN1(n10757), .IN2(n10758), .Q(n10751) );
  AND2X1 U10573 ( .IN1(n10759), .IN2(g1444), .Q(n10758) );
  AND2X1 U10574 ( .IN1(n10168), .IN2(n10760), .Q(n10757) );
  OR2X1 U10575 ( .IN1(n10761), .IN2(n10762), .Q(n10749) );
  AND2X1 U10576 ( .IN1(n10763), .IN2(g1435), .Q(n10762) );
  AND2X1 U10577 ( .IN1(n10174), .IN2(n10764), .Q(n10761) );
  OR2X1 U10578 ( .IN1(n10765), .IN2(n10766), .Q(n10747) );
  OR2X1 U10579 ( .IN1(n10767), .IN2(n10768), .Q(n10766) );
  OR2X1 U10580 ( .IN1(n10769), .IN2(n10770), .Q(n10768) );
  AND2X1 U10581 ( .IN1(n10771), .IN2(g1466), .Q(n10770) );
  AND2X1 U10582 ( .IN1(n9883), .IN2(n10772), .Q(n10769) );
  OR2X1 U10583 ( .IN1(n10773), .IN2(n10774), .Q(n10767) );
  AND2X1 U10584 ( .IN1(n10775), .IN2(g1426), .Q(n10774) );
  AND2X1 U10585 ( .IN1(n9354), .IN2(n10776), .Q(n10773) );
  OR2X1 U10586 ( .IN1(n10777), .IN2(n10778), .Q(n10765) );
  AND2X1 U10587 ( .IN1(n10779), .IN2(g1453), .Q(n10778) );
  AND2X1 U10588 ( .IN1(n10186), .IN2(n10780), .Q(n10777) );
  OR2X1 U10589 ( .IN1(n10781), .IN2(n10782), .Q(n10745) );
  OR2X1 U10590 ( .IN1(n10783), .IN2(n10784), .Q(n10782) );
  OR2X1 U10591 ( .IN1(n10785), .IN2(n10786), .Q(n10784) );
  OR2X1 U10592 ( .IN1(n10787), .IN2(n10788), .Q(n10786) );
  AND2X1 U10593 ( .IN1(n10789), .IN2(g1457), .Q(n10788) );
  AND2X1 U10594 ( .IN1(n9882), .IN2(n10790), .Q(n10787) );
  OR2X1 U10595 ( .IN1(n10791), .IN2(n10792), .Q(n10785) );
  AND2X1 U10596 ( .IN1(n10793), .IN2(g1430), .Q(n10792) );
  AND2X1 U10597 ( .IN1(n9508), .IN2(n10794), .Q(n10791) );
  OR2X1 U10598 ( .IN1(n10795), .IN2(n10796), .Q(n10783) );
  AND2X1 U10599 ( .IN1(n10797), .IN2(g1439), .Q(n10796) );
  AND2X1 U10600 ( .IN1(n9880), .IN2(n10798), .Q(n10795) );
  OR2X1 U10601 ( .IN1(n10799), .IN2(n10800), .Q(n10781) );
  OR2X1 U10602 ( .IN1(n10801), .IN2(n10672), .Q(n10800) );
  OR2X1 U10603 ( .IN1(n10802), .IN2(n10803), .Q(n10799) );
  AND2X1 U10604 ( .IN1(n10804), .IN2(g1448), .Q(n10803) );
  AND2X1 U10605 ( .IN1(n9881), .IN2(n10805), .Q(n10802) );
  OR2X1 U10606 ( .IN1(n10806), .IN2(n10807), .Q(n10743) );
  AND2X1 U10607 ( .IN1(n10808), .IN2(n10809), .Q(n4275) );
  OR2X1 U10608 ( .IN1(n10810), .IN2(n10811), .Q(n10809) );
  OR2X1 U10609 ( .IN1(n10812), .IN2(n10813), .Q(n10811) );
  OR2X1 U10610 ( .IN1(n10814), .IN2(n10815), .Q(n10813) );
  OR2X1 U10611 ( .IN1(n10816), .IN2(n10817), .Q(n10815) );
  OR2X1 U10612 ( .IN1(n10818), .IN2(n10819), .Q(n10817) );
  AND2X1 U10613 ( .IN1(n10820), .IN2(g2120), .Q(n10819) );
  AND2X1 U10614 ( .IN1(n9353), .IN2(n10821), .Q(n10818) );
  OR2X1 U10615 ( .IN1(n10822), .IN2(n10823), .Q(n10816) );
  AND2X1 U10616 ( .IN1(n10824), .IN2(g2138), .Q(n10823) );
  AND2X1 U10617 ( .IN1(n10169), .IN2(n10825), .Q(n10822) );
  OR2X1 U10618 ( .IN1(n10826), .IN2(n10827), .Q(n10814) );
  AND2X1 U10619 ( .IN1(n10828), .IN2(g2129), .Q(n10827) );
  AND2X1 U10620 ( .IN1(n10175), .IN2(n10829), .Q(n10826) );
  OR2X1 U10621 ( .IN1(n10830), .IN2(n10831), .Q(n10812) );
  OR2X1 U10622 ( .IN1(n10832), .IN2(n10833), .Q(n10831) );
  OR2X1 U10623 ( .IN1(n10834), .IN2(n10835), .Q(n10833) );
  AND2X1 U10624 ( .IN1(n10836), .IN2(g2124), .Q(n10835) );
  AND2X1 U10625 ( .IN1(n9507), .IN2(n10837), .Q(n10834) );
  OR2X1 U10626 ( .IN1(n10838), .IN2(n10839), .Q(n10832) );
  AND2X1 U10627 ( .IN1(n10840), .IN2(g2147), .Q(n10839) );
  AND2X1 U10628 ( .IN1(n10187), .IN2(n10841), .Q(n10838) );
  OR2X1 U10629 ( .IN1(n10842), .IN2(n10843), .Q(n10830) );
  AND2X1 U10630 ( .IN1(n10844), .IN2(g2160), .Q(n10843) );
  AND2X1 U10631 ( .IN1(n9879), .IN2(n10845), .Q(n10842) );
  OR2X1 U10632 ( .IN1(n10846), .IN2(n10847), .Q(n10810) );
  OR2X1 U10633 ( .IN1(n10848), .IN2(n10849), .Q(n10847) );
  OR2X1 U10634 ( .IN1(n10850), .IN2(n10851), .Q(n10849) );
  OR2X1 U10635 ( .IN1(n10852), .IN2(n10853), .Q(n10851) );
  AND2X1 U10636 ( .IN1(n10854), .IN2(g2142), .Q(n10853) );
  AND2X1 U10637 ( .IN1(n9877), .IN2(n10855), .Q(n10852) );
  OR2X1 U10638 ( .IN1(n10856), .IN2(n10857), .Q(n10850) );
  AND2X1 U10639 ( .IN1(n10858), .IN2(g2133), .Q(n10857) );
  AND2X1 U10640 ( .IN1(n9876), .IN2(n10859), .Q(n10856) );
  OR2X1 U10641 ( .IN1(n10860), .IN2(n10861), .Q(n10848) );
  AND2X1 U10642 ( .IN1(n10862), .IN2(g2151), .Q(n10861) );
  AND2X1 U10643 ( .IN1(n9878), .IN2(n10863), .Q(n10860) );
  OR2X1 U10644 ( .IN1(n10864), .IN2(n10865), .Q(n10846) );
  OR2X1 U10645 ( .IN1(n10866), .IN2(n10672), .Q(n10865) );
  AND2X1 U10646 ( .IN1(n10867), .IN2(n10868), .Q(n10864) );
  INVX0 U10647 ( .INP(n10869), .ZN(n10868) );
  AND2X1 U10648 ( .IN1(n10870), .IN2(test_so78), .Q(n10869) );
  OR2X1 U10649 ( .IN1(test_so78), .IN2(n10870), .Q(n10867) );
  OR2X1 U10650 ( .IN1(n2489), .IN2(n10871), .Q(n10808) );
  INVX0 U10651 ( .INP(n10872), .ZN(n4273) );
  AND2X1 U10652 ( .IN1(n10873), .IN2(n10874), .Q(n10872) );
  OR2X1 U10653 ( .IN1(n10875), .IN2(n10876), .Q(n10873) );
  AND2X1 U10654 ( .IN1(n10877), .IN2(n4482), .Q(n10875) );
  OR2X1 U10655 ( .IN1(n10878), .IN2(n10879), .Q(n4272) );
  OR2X1 U10656 ( .IN1(n10880), .IN2(n10881), .Q(n10879) );
  AND2X1 U10657 ( .IN1(test_so27), .IN2(n10882), .Q(n10881) );
  AND2X1 U10658 ( .IN1(n10883), .IN2(n10884), .Q(n10880) );
  OR2X1 U10659 ( .IN1(n10885), .IN2(n10886), .Q(n4271) );
  OR2X1 U10660 ( .IN1(n10887), .IN2(n10888), .Q(n10886) );
  AND2X1 U10661 ( .IN1(n10882), .IN2(g536), .Q(n10888) );
  AND2X1 U10662 ( .IN1(n10883), .IN2(n10889), .Q(n10887) );
  AND2X1 U10663 ( .IN1(n2446), .IN2(n10890), .Q(n10885) );
  OR2X1 U10664 ( .IN1(n10891), .IN2(n10892), .Q(n4270) );
  OR2X1 U10665 ( .IN1(n10893), .IN2(n10894), .Q(n10892) );
  AND2X1 U10666 ( .IN1(n10882), .IN2(g537), .Q(n10894) );
  AND2X1 U10667 ( .IN1(n10883), .IN2(n10895), .Q(n10893) );
  AND2X1 U10668 ( .IN1(n2446), .IN2(n10896), .Q(n10891) );
  OR2X1 U10669 ( .IN1(n10897), .IN2(n10898), .Q(n4269) );
  OR2X1 U10670 ( .IN1(n10899), .IN2(n10900), .Q(n10898) );
  AND2X1 U10671 ( .IN1(n10882), .IN2(n8047), .Q(n10900) );
  AND2X1 U10672 ( .IN1(n10901), .IN2(n10902), .Q(n10899) );
  AND2X1 U10673 ( .IN1(n10903), .IN2(n10904), .Q(n10901) );
  OR2X1 U10674 ( .IN1(n10905), .IN2(n10906), .Q(n4268) );
  OR2X1 U10675 ( .IN1(n10907), .IN2(n10908), .Q(n10905) );
  AND2X1 U10676 ( .IN1(n10882), .IN2(n8046), .Q(n10908) );
  AND2X1 U10677 ( .IN1(n10909), .IN2(n10902), .Q(n10907) );
  AND2X1 U10678 ( .IN1(n10910), .IN2(n10904), .Q(n10909) );
  OR2X1 U10679 ( .IN1(n10911), .IN2(n10906), .Q(n4267) );
  OR2X1 U10680 ( .IN1(n10878), .IN2(n10912), .Q(n10906) );
  INVX0 U10681 ( .INP(n2440), .ZN(n10912) );
  OR2X1 U10682 ( .IN1(n10913), .IN2(n10914), .Q(n10911) );
  AND2X1 U10683 ( .IN1(n10882), .IN2(n8045), .Q(n10914) );
  AND2X1 U10684 ( .IN1(n10915), .IN2(n10902), .Q(n10913) );
  AND2X1 U10685 ( .IN1(n10916), .IN2(n10904), .Q(n10915) );
  OR2X1 U10686 ( .IN1(n10897), .IN2(n10917), .Q(n4266) );
  OR2X1 U10687 ( .IN1(n10918), .IN2(n10919), .Q(n10917) );
  AND2X1 U10688 ( .IN1(n10882), .IN2(n8044), .Q(n10919) );
  AND2X1 U10689 ( .IN1(n10920), .IN2(n10902), .Q(n10918) );
  AND2X1 U10690 ( .IN1(n10921), .IN2(n10904), .Q(n10920) );
  OR2X1 U10691 ( .IN1(n10922), .IN2(n10878), .Q(n10897) );
  AND2X1 U10692 ( .IN1(n2446), .IN2(n2445), .Q(n10922) );
  OR2X1 U10693 ( .IN1(n10878), .IN2(n10923), .Q(n4265) );
  OR2X1 U10694 ( .IN1(n10924), .IN2(n10925), .Q(n10923) );
  AND2X1 U10695 ( .IN1(n10882), .IN2(n8043), .Q(n10925) );
  AND2X1 U10696 ( .IN1(n10926), .IN2(n10902), .Q(n10882) );
  AND2X1 U10697 ( .IN1(n10883), .IN2(n10927), .Q(n10924) );
  AND2X1 U10698 ( .IN1(n10904), .IN2(n10902), .Q(n10883) );
  INVX0 U10699 ( .INP(n10928), .ZN(n10904) );
  INVX0 U10700 ( .INP(n2426), .ZN(n10878) );
  OR2X1 U10701 ( .IN1(g3234), .IN2(n7912), .Q(n4263) );
  OR2X1 U10702 ( .IN1(n10929), .IN2(n10930), .Q(n4262) );
  INVX0 U10703 ( .INP(n10931), .ZN(n10930) );
  AND2X1 U10704 ( .IN1(n10932), .IN2(n10933), .Q(n10929) );
  OR2X1 U10705 ( .IN1(n10934), .IN2(g3018), .Q(n10932) );
  AND2X1 U10706 ( .IN1(n10935), .IN2(n10936), .Q(n4261) );
  INVX0 U10707 ( .INP(n10937), .ZN(n10936) );
  AND2X1 U10708 ( .IN1(n10938), .IN2(n10939), .Q(n10937) );
  OR2X1 U10709 ( .IN1(n10939), .IN2(n10938), .Q(n10935) );
  OR2X1 U10710 ( .IN1(n10940), .IN2(n10941), .Q(n4260) );
  INVX0 U10711 ( .INP(n10942), .ZN(n10941) );
  OR2X1 U10712 ( .IN1(n10943), .IN2(n10939), .Q(n10942) );
  AND2X1 U10713 ( .IN1(n10939), .IN2(n10943), .Q(n10940) );
  AND2X1 U10714 ( .IN1(n8078), .IN2(n10944), .Q(n10939) );
  OR2X1 U10715 ( .IN1(n10945), .IN2(n10946), .Q(n4259) );
  OR2X1 U10716 ( .IN1(n10947), .IN2(n10948), .Q(n10946) );
  AND2X1 U10717 ( .IN1(n10949), .IN2(g557), .Q(n10948) );
  OR2X1 U10718 ( .IN1(n10950), .IN2(n10951), .Q(n10949) );
  INVX0 U10719 ( .INP(n10952), .ZN(n10951) );
  OR2X1 U10720 ( .IN1(n10896), .IN2(n10953), .Q(n10952) );
  AND2X1 U10721 ( .IN1(n10953), .IN2(n10896), .Q(n10950) );
  OR2X1 U10722 ( .IN1(n10954), .IN2(n10955), .Q(n10896) );
  OR2X1 U10723 ( .IN1(n10956), .IN2(n10957), .Q(n10954) );
  AND2X1 U10724 ( .IN1(n10958), .IN2(n10959), .Q(n10957) );
  AND2X1 U10725 ( .IN1(n10960), .IN2(n10961), .Q(n10956) );
  INVX0 U10726 ( .INP(n10890), .ZN(n10953) );
  OR2X1 U10727 ( .IN1(n10962), .IN2(n10963), .Q(n10890) );
  OR2X1 U10728 ( .IN1(n10964), .IN2(n10965), .Q(n10963) );
  AND2X1 U10729 ( .IN1(n10966), .IN2(n10967), .Q(n10965) );
  AND2X1 U10730 ( .IN1(n10968), .IN2(n10969), .Q(n10964) );
  AND2X1 U10731 ( .IN1(n10970), .IN2(n10971), .Q(n10947) );
  AND2X1 U10732 ( .IN1(n10972), .IN2(n10973), .Q(n10971) );
  OR2X1 U10733 ( .IN1(g3229), .IN2(n8040), .Q(n10973) );
  OR2X1 U10734 ( .IN1(n10974), .IN2(g538), .Q(n10972) );
  AND2X1 U10735 ( .IN1(n10928), .IN2(n10902), .Q(n10970) );
  INVX0 U10736 ( .INP(n10975), .ZN(n10902) );
  AND2X1 U10737 ( .IN1(n10926), .IN2(n549), .Q(n10928) );
  INVX0 U10738 ( .INP(n10976), .ZN(n549) );
  AND2X1 U10739 ( .IN1(test_so22), .IN2(n10977), .Q(n10945) );
  OR2X1 U10740 ( .IN1(n10978), .IN2(n10979), .Q(n10977) );
  INVX0 U10741 ( .INP(n10980), .ZN(n10979) );
  OR2X1 U10742 ( .IN1(n10981), .IN2(n10982), .Q(n10980) );
  AND2X1 U10743 ( .IN1(n10982), .IN2(n10981), .Q(n10978) );
  AND2X1 U10744 ( .IN1(n10983), .IN2(n10984), .Q(n10981) );
  INVX0 U10745 ( .INP(n10985), .ZN(n10984) );
  AND2X1 U10746 ( .IN1(n10986), .IN2(n10987), .Q(n10985) );
  OR2X1 U10747 ( .IN1(n10987), .IN2(n10986), .Q(n10983) );
  OR2X1 U10748 ( .IN1(n10988), .IN2(n10989), .Q(n10986) );
  AND2X1 U10749 ( .IN1(n10990), .IN2(n10921), .Q(n10989) );
  INVX0 U10750 ( .INP(n10991), .ZN(n10988) );
  OR2X1 U10751 ( .IN1(n10921), .IN2(n10990), .Q(n10991) );
  INVX0 U10752 ( .INP(n10927), .ZN(n10990) );
  OR2X1 U10753 ( .IN1(n10962), .IN2(n10992), .Q(n10927) );
  OR2X1 U10754 ( .IN1(n10993), .IN2(n10994), .Q(n10992) );
  AND2X1 U10755 ( .IN1(n10995), .IN2(n10967), .Q(n10994) );
  AND2X1 U10756 ( .IN1(n10968), .IN2(n10996), .Q(n10993) );
  OR2X1 U10757 ( .IN1(n10997), .IN2(n10998), .Q(n10921) );
  OR2X1 U10758 ( .IN1(n10999), .IN2(n11000), .Q(n10998) );
  AND2X1 U10759 ( .IN1(n10958), .IN2(n11001), .Q(n11000) );
  AND2X1 U10760 ( .IN1(n11002), .IN2(n10961), .Q(n10999) );
  AND2X1 U10761 ( .IN1(n11003), .IN2(n11004), .Q(n10987) );
  INVX0 U10762 ( .INP(n11005), .ZN(n11004) );
  AND2X1 U10763 ( .IN1(n11006), .IN2(n10910), .Q(n11005) );
  OR2X1 U10764 ( .IN1(n10910), .IN2(n11006), .Q(n11003) );
  INVX0 U10765 ( .INP(n10916), .ZN(n11006) );
  OR2X1 U10766 ( .IN1(n10997), .IN2(n11007), .Q(n10916) );
  OR2X1 U10767 ( .IN1(n11008), .IN2(n11009), .Q(n11007) );
  AND2X1 U10768 ( .IN1(n11010), .IN2(n10967), .Q(n11009) );
  AND2X1 U10769 ( .IN1(n10968), .IN2(n11011), .Q(n11008) );
  OR2X1 U10770 ( .IN1(n10997), .IN2(n11012), .Q(n10910) );
  OR2X1 U10771 ( .IN1(n11013), .IN2(n11014), .Q(n11012) );
  AND2X1 U10772 ( .IN1(n10958), .IN2(n11015), .Q(n11014) );
  AND2X1 U10773 ( .IN1(n11016), .IN2(n10961), .Q(n11013) );
  OR2X1 U10774 ( .IN1(n11017), .IN2(n11018), .Q(n10982) );
  INVX0 U10775 ( .INP(n11019), .ZN(n11018) );
  OR2X1 U10776 ( .IN1(n11020), .IN2(n11021), .Q(n11019) );
  AND2X1 U10777 ( .IN1(n11021), .IN2(n11020), .Q(n11017) );
  AND2X1 U10778 ( .IN1(n11022), .IN2(n11023), .Q(n11020) );
  INVX0 U10779 ( .INP(n11024), .ZN(n11023) );
  AND2X1 U10780 ( .IN1(n11025), .IN2(n10895), .Q(n11024) );
  OR2X1 U10781 ( .IN1(n10895), .IN2(n11025), .Q(n11022) );
  INVX0 U10782 ( .INP(n10903), .ZN(n11025) );
  OR2X1 U10783 ( .IN1(n10997), .IN2(n11026), .Q(n10903) );
  OR2X1 U10784 ( .IN1(n11027), .IN2(n11028), .Q(n11026) );
  AND2X1 U10785 ( .IN1(n11029), .IN2(n10967), .Q(n11028) );
  AND2X1 U10786 ( .IN1(n10968), .IN2(n11030), .Q(n11027) );
  OR2X1 U10787 ( .IN1(n10997), .IN2(n11031), .Q(n10895) );
  OR2X1 U10788 ( .IN1(n11032), .IN2(n11033), .Q(n11031) );
  AND2X1 U10789 ( .IN1(n10958), .IN2(n11034), .Q(n11033) );
  AND2X1 U10790 ( .IN1(n11035), .IN2(n10961), .Q(n11032) );
  OR2X1 U10791 ( .IN1(n11036), .IN2(n11037), .Q(n11021) );
  AND2X1 U10792 ( .IN1(n11038), .IN2(n10884), .Q(n11037) );
  INVX0 U10793 ( .INP(n10889), .ZN(n11038) );
  AND2X1 U10794 ( .IN1(n11039), .IN2(n10889), .Q(n11036) );
  OR2X1 U10795 ( .IN1(n10962), .IN2(n11040), .Q(n10889) );
  OR2X1 U10796 ( .IN1(n11041), .IN2(n11042), .Q(n11040) );
  AND2X1 U10797 ( .IN1(n11043), .IN2(n10967), .Q(n11042) );
  AND2X1 U10798 ( .IN1(n10968), .IN2(n11044), .Q(n11041) );
  AND2X1 U10799 ( .IN1(n11045), .IN2(n11046), .Q(n10968) );
  OR2X1 U10800 ( .IN1(n11047), .IN2(n10997), .Q(n10962) );
  INVX0 U10801 ( .INP(n11048), .ZN(n11047) );
  OR2X1 U10802 ( .IN1(n11045), .IN2(n11046), .Q(n11048) );
  INVX0 U10803 ( .INP(n10884), .ZN(n11039) );
  OR2X1 U10804 ( .IN1(n11049), .IN2(n10955), .Q(n10884) );
  OR2X1 U10805 ( .IN1(n11050), .IN2(n10997), .Q(n10955) );
  OR2X1 U10806 ( .IN1(n4541), .IN2(n10976), .Q(n10997) );
  OR2X1 U10807 ( .IN1(n11051), .IN2(n11052), .Q(n10976) );
  OR2X1 U10808 ( .IN1(g559), .IN2(g21851), .Q(n11052) );
  OR2X1 U10809 ( .IN1(g563), .IN2(n11053), .Q(n11051) );
  AND2X1 U10810 ( .IN1(n4541), .IN2(n11054), .Q(n11053) );
  INVX0 U10811 ( .INP(n2459), .ZN(n11050) );
  OR2X1 U10812 ( .IN1(n11055), .IN2(n11056), .Q(n11049) );
  AND2X1 U10813 ( .IN1(n10958), .IN2(n11057), .Q(n11056) );
  AND2X1 U10814 ( .IN1(n11045), .IN2(n11058), .Q(n10958) );
  AND2X1 U10815 ( .IN1(n11059), .IN2(n10961), .Q(n11055) );
  OR2X1 U10816 ( .IN1(n11060), .IN2(n11061), .Q(n4258) );
  OR2X1 U10817 ( .IN1(n11062), .IN2(n11063), .Q(n11061) );
  AND2X1 U10818 ( .IN1(n11064), .IN2(g2611), .Q(n11063) );
  AND2X1 U10819 ( .IN1(n11065), .IN2(n11066), .Q(n11062) );
  AND2X1 U10820 ( .IN1(n2361), .IN2(n11067), .Q(n11060) );
  OR2X1 U10821 ( .IN1(n11068), .IN2(n11069), .Q(n4257) );
  OR2X1 U10822 ( .IN1(n11070), .IN2(n11071), .Q(n11069) );
  AND2X1 U10823 ( .IN1(n11064), .IN2(n7924), .Q(n11070) );
  OR2X1 U10824 ( .IN1(n11072), .IN2(n11073), .Q(n11068) );
  AND2X1 U10825 ( .IN1(n11074), .IN2(n11075), .Q(n11073) );
  AND2X1 U10826 ( .IN1(n11076), .IN2(n11077), .Q(n11074) );
  OR2X1 U10827 ( .IN1(n11078), .IN2(n11079), .Q(n4256) );
  OR2X1 U10828 ( .IN1(n11072), .IN2(n11080), .Q(n11079) );
  AND2X1 U10829 ( .IN1(n11065), .IN2(n11081), .Q(n11080) );
  AND2X1 U10830 ( .IN1(n11064), .IN2(n7920), .Q(n11078) );
  OR2X1 U10831 ( .IN1(n11082), .IN2(n11083), .Q(n4255) );
  OR2X1 U10832 ( .IN1(n11084), .IN2(n11071), .Q(n11083) );
  INVX0 U10833 ( .INP(n2375), .ZN(n11071) );
  AND2X1 U10834 ( .IN1(n11064), .IN2(n7923), .Q(n11084) );
  OR2X1 U10835 ( .IN1(n11072), .IN2(n11085), .Q(n11082) );
  AND2X1 U10836 ( .IN1(n11086), .IN2(n11075), .Q(n11085) );
  AND2X1 U10837 ( .IN1(n11087), .IN2(n11077), .Q(n11086) );
  OR2X1 U10838 ( .IN1(n11088), .IN2(n11089), .Q(n4254) );
  OR2X1 U10839 ( .IN1(n11090), .IN2(n11091), .Q(n11089) );
  AND2X1 U10840 ( .IN1(n11064), .IN2(n7925), .Q(n11091) );
  AND2X1 U10841 ( .IN1(n11092), .IN2(n11075), .Q(n11090) );
  AND2X1 U10842 ( .IN1(n11093), .IN2(n11077), .Q(n11092) );
  OR2X1 U10843 ( .IN1(n11094), .IN2(n11095), .Q(n4253) );
  OR2X1 U10844 ( .IN1(n11096), .IN2(n11097), .Q(n11095) );
  AND2X1 U10845 ( .IN1(test_so91), .IN2(n11064), .Q(n11097) );
  AND2X1 U10846 ( .IN1(n11065), .IN2(n11098), .Q(n11096) );
  AND2X1 U10847 ( .IN1(n2361), .IN2(n11099), .Q(n11094) );
  OR2X1 U10848 ( .IN1(n11088), .IN2(n11100), .Q(n4252) );
  OR2X1 U10849 ( .IN1(n11101), .IN2(n11102), .Q(n11100) );
  AND2X1 U10850 ( .IN1(n11064), .IN2(n7922), .Q(n11102) );
  AND2X1 U10851 ( .IN1(n11103), .IN2(n11075), .Q(n11101) );
  AND2X1 U10852 ( .IN1(n11104), .IN2(n11077), .Q(n11103) );
  OR2X1 U10853 ( .IN1(n11072), .IN2(n11105), .Q(n11088) );
  AND2X1 U10854 ( .IN1(n2361), .IN2(n2374), .Q(n11105) );
  OR2X1 U10855 ( .IN1(n11106), .IN2(n11107), .Q(n4251) );
  OR2X1 U10856 ( .IN1(n11072), .IN2(n11108), .Q(n11107) );
  AND2X1 U10857 ( .IN1(n11065), .IN2(n11109), .Q(n11108) );
  AND2X1 U10858 ( .IN1(n11077), .IN2(n11075), .Q(n11065) );
  AND2X1 U10859 ( .IN1(n11110), .IN2(n2361), .Q(n11072) );
  AND2X1 U10860 ( .IN1(n11064), .IN2(n7921), .Q(n11106) );
  AND2X1 U10861 ( .IN1(n11111), .IN2(n11075), .Q(n11064) );
  OR2X1 U10862 ( .IN1(n11112), .IN2(n11113), .Q(n4250) );
  OR2X1 U10863 ( .IN1(n11114), .IN2(n11115), .Q(n11113) );
  AND2X1 U10864 ( .IN1(n11116), .IN2(g2584), .Q(n11115) );
  OR2X1 U10865 ( .IN1(n11117), .IN2(n11118), .Q(n11116) );
  INVX0 U10866 ( .INP(n11119), .ZN(n11118) );
  OR2X1 U10867 ( .IN1(n11120), .IN2(n11121), .Q(n11119) );
  AND2X1 U10868 ( .IN1(n11121), .IN2(n11120), .Q(n11117) );
  AND2X1 U10869 ( .IN1(n11122), .IN2(n11123), .Q(n11120) );
  INVX0 U10870 ( .INP(n11124), .ZN(n11123) );
  AND2X1 U10871 ( .IN1(n11125), .IN2(n11126), .Q(n11124) );
  OR2X1 U10872 ( .IN1(n11126), .IN2(n11125), .Q(n11122) );
  OR2X1 U10873 ( .IN1(n11127), .IN2(n11128), .Q(n11125) );
  AND2X1 U10874 ( .IN1(n11129), .IN2(n11104), .Q(n11128) );
  INVX0 U10875 ( .INP(n11130), .ZN(n11127) );
  OR2X1 U10876 ( .IN1(n11104), .IN2(n11129), .Q(n11130) );
  INVX0 U10877 ( .INP(n11109), .ZN(n11129) );
  OR2X1 U10878 ( .IN1(n11131), .IN2(n11132), .Q(n11109) );
  OR2X1 U10879 ( .IN1(n11133), .IN2(n11134), .Q(n11132) );
  AND2X1 U10880 ( .IN1(n11135), .IN2(n11136), .Q(n11134) );
  AND2X1 U10881 ( .IN1(n11137), .IN2(n11138), .Q(n11133) );
  OR2X1 U10882 ( .IN1(n11139), .IN2(n11140), .Q(n11104) );
  OR2X1 U10883 ( .IN1(n11141), .IN2(n11142), .Q(n11140) );
  AND2X1 U10884 ( .IN1(n11143), .IN2(n11144), .Q(n11142) );
  AND2X1 U10885 ( .IN1(n11145), .IN2(n11146), .Q(n11141) );
  AND2X1 U10886 ( .IN1(n11147), .IN2(n11148), .Q(n11126) );
  INVX0 U10887 ( .INP(n11149), .ZN(n11148) );
  AND2X1 U10888 ( .IN1(n11150), .IN2(n11093), .Q(n11149) );
  OR2X1 U10889 ( .IN1(n11093), .IN2(n11150), .Q(n11147) );
  INVX0 U10890 ( .INP(n11098), .ZN(n11150) );
  OR2X1 U10891 ( .IN1(n11131), .IN2(n11151), .Q(n11098) );
  OR2X1 U10892 ( .IN1(n11152), .IN2(n11153), .Q(n11151) );
  AND2X1 U10893 ( .IN1(n11154), .IN2(n11136), .Q(n11153) );
  AND2X1 U10894 ( .IN1(n11137), .IN2(n11155), .Q(n11152) );
  OR2X1 U10895 ( .IN1(n11139), .IN2(n11156), .Q(n11093) );
  OR2X1 U10896 ( .IN1(n11157), .IN2(n11158), .Q(n11156) );
  AND2X1 U10897 ( .IN1(n11159), .IN2(n11136), .Q(n11158) );
  AND2X1 U10898 ( .IN1(n11137), .IN2(n11160), .Q(n11157) );
  OR2X1 U10899 ( .IN1(n11161), .IN2(n11162), .Q(n11121) );
  INVX0 U10900 ( .INP(n11163), .ZN(n11162) );
  OR2X1 U10901 ( .IN1(n11164), .IN2(n11165), .Q(n11163) );
  AND2X1 U10902 ( .IN1(n11165), .IN2(n11164), .Q(n11161) );
  AND2X1 U10903 ( .IN1(n11166), .IN2(n11167), .Q(n11164) );
  INVX0 U10904 ( .INP(n11168), .ZN(n11167) );
  AND2X1 U10905 ( .IN1(n11169), .IN2(n11081), .Q(n11168) );
  OR2X1 U10906 ( .IN1(n11081), .IN2(n11169), .Q(n11166) );
  INVX0 U10907 ( .INP(n11087), .ZN(n11169) );
  OR2X1 U10908 ( .IN1(n11139), .IN2(n11170), .Q(n11087) );
  OR2X1 U10909 ( .IN1(n11171), .IN2(n11172), .Q(n11170) );
  AND2X1 U10910 ( .IN1(n11173), .IN2(n11136), .Q(n11172) );
  AND2X1 U10911 ( .IN1(n11137), .IN2(n11174), .Q(n11171) );
  OR2X1 U10912 ( .IN1(n11175), .IN2(n11176), .Q(n11081) );
  OR2X1 U10913 ( .IN1(n11177), .IN2(n11178), .Q(n11175) );
  AND2X1 U10914 ( .IN1(n11143), .IN2(n11179), .Q(n11178) );
  AND2X1 U10915 ( .IN1(n11180), .IN2(n11146), .Q(n11177) );
  OR2X1 U10916 ( .IN1(n11181), .IN2(n11182), .Q(n11165) );
  AND2X1 U10917 ( .IN1(n11183), .IN2(n11066), .Q(n11182) );
  INVX0 U10918 ( .INP(n11076), .ZN(n11183) );
  AND2X1 U10919 ( .IN1(n11184), .IN2(n11076), .Q(n11181) );
  OR2X1 U10920 ( .IN1(n11139), .IN2(n11185), .Q(n11076) );
  OR2X1 U10921 ( .IN1(n11186), .IN2(n11187), .Q(n11185) );
  AND2X1 U10922 ( .IN1(n11143), .IN2(n11188), .Q(n11187) );
  AND2X1 U10923 ( .IN1(n11189), .IN2(n11146), .Q(n11186) );
  INVX0 U10924 ( .INP(n11066), .ZN(n11184) );
  OR2X1 U10925 ( .IN1(n11139), .IN2(n11190), .Q(n11066) );
  OR2X1 U10926 ( .IN1(n11191), .IN2(n11192), .Q(n11190) );
  AND2X1 U10927 ( .IN1(n11143), .IN2(n11193), .Q(n11192) );
  AND2X1 U10928 ( .IN1(n11194), .IN2(n11146), .Q(n11191) );
  AND2X1 U10929 ( .IN1(n11195), .IN2(n11196), .Q(n11114) );
  AND2X1 U10930 ( .IN1(n11197), .IN2(n11198), .Q(n11196) );
  OR2X1 U10931 ( .IN1(g3229), .IN2(n7918), .Q(n11198) );
  OR2X1 U10932 ( .IN1(n10974), .IN2(g2612), .Q(n11197) );
  AND2X1 U10933 ( .IN1(n11199), .IN2(n11075), .Q(n11195) );
  INVX0 U10934 ( .INP(n11200), .ZN(n11075) );
  INVX0 U10935 ( .INP(n11077), .ZN(n11199) );
  OR2X1 U10936 ( .IN1(n11110), .IN2(n11201), .Q(n11077) );
  AND2X1 U10937 ( .IN1(n11202), .IN2(g2631), .Q(n11112) );
  OR2X1 U10938 ( .IN1(n11203), .IN2(n11204), .Q(n11202) );
  INVX0 U10939 ( .INP(n11205), .ZN(n11204) );
  OR2X1 U10940 ( .IN1(n11099), .IN2(n11206), .Q(n11205) );
  AND2X1 U10941 ( .IN1(n11206), .IN2(n11099), .Q(n11203) );
  OR2X1 U10942 ( .IN1(n11131), .IN2(n11207), .Q(n11099) );
  OR2X1 U10943 ( .IN1(n11208), .IN2(n11209), .Q(n11207) );
  AND2X1 U10944 ( .IN1(n11210), .IN2(n11136), .Q(n11209) );
  AND2X1 U10945 ( .IN1(n11137), .IN2(n11211), .Q(n11208) );
  AND2X1 U10946 ( .IN1(n11212), .IN2(n11213), .Q(n11137) );
  OR2X1 U10947 ( .IN1(n11214), .IN2(n11139), .Q(n11131) );
  INVX0 U10948 ( .INP(n11215), .ZN(n11214) );
  OR2X1 U10949 ( .IN1(n11212), .IN2(n11213), .Q(n11215) );
  INVX0 U10950 ( .INP(n11067), .ZN(n11206) );
  OR2X1 U10951 ( .IN1(n11216), .IN2(n11176), .Q(n11067) );
  OR2X1 U10952 ( .IN1(n11217), .IN2(n11139), .Q(n11176) );
  OR2X1 U10953 ( .IN1(n4543), .IN2(n11110), .Q(n11139) );
  OR2X1 U10954 ( .IN1(g2633), .IN2(n11218), .Q(n11110) );
  OR2X1 U10955 ( .IN1(g2637), .IN2(g30072), .Q(n11218) );
  INVX0 U10956 ( .INP(n2381), .ZN(n11217) );
  OR2X1 U10957 ( .IN1(n11219), .IN2(n11220), .Q(n11216) );
  AND2X1 U10958 ( .IN1(n11143), .IN2(n11221), .Q(n11220) );
  AND2X1 U10959 ( .IN1(n11212), .IN2(n11222), .Q(n11143) );
  AND2X1 U10960 ( .IN1(n11223), .IN2(n11146), .Q(n11219) );
  OR2X1 U10961 ( .IN1(n11224), .IN2(n11225), .Q(n4249) );
  OR2X1 U10962 ( .IN1(n11226), .IN2(n11227), .Q(n11225) );
  AND2X1 U10963 ( .IN1(n11228), .IN2(g1917), .Q(n11227) );
  AND2X1 U10964 ( .IN1(n11229), .IN2(n11230), .Q(n11226) );
  AND2X1 U10965 ( .IN1(n2289), .IN2(n11231), .Q(n11224) );
  OR2X1 U10966 ( .IN1(n11232), .IN2(n11233), .Q(n4248) );
  OR2X1 U10967 ( .IN1(n11234), .IN2(n11235), .Q(n11232) );
  AND2X1 U10968 ( .IN1(n11228), .IN2(n7966), .Q(n11235) );
  AND2X1 U10969 ( .IN1(n11236), .IN2(n11237), .Q(n11234) );
  AND2X1 U10970 ( .IN1(n11238), .IN2(n11239), .Q(n11236) );
  OR2X1 U10971 ( .IN1(n11240), .IN2(n11241), .Q(n4247) );
  OR2X1 U10972 ( .IN1(n11242), .IN2(n11243), .Q(n11241) );
  AND2X1 U10973 ( .IN1(n11228), .IN2(n7962), .Q(n11243) );
  AND2X1 U10974 ( .IN1(n11229), .IN2(n11244), .Q(n11242) );
  OR2X1 U10975 ( .IN1(n11245), .IN2(n11233), .Q(n4246) );
  OR2X1 U10976 ( .IN1(n11240), .IN2(n11246), .Q(n11233) );
  INVX0 U10977 ( .INP(n2303), .ZN(n11246) );
  OR2X1 U10978 ( .IN1(n11247), .IN2(n11248), .Q(n11245) );
  AND2X1 U10979 ( .IN1(n11228), .IN2(n7965), .Q(n11248) );
  AND2X1 U10980 ( .IN1(n11249), .IN2(n11237), .Q(n11247) );
  AND2X1 U10981 ( .IN1(n11250), .IN2(n11239), .Q(n11249) );
  OR2X1 U10982 ( .IN1(n11251), .IN2(n11252), .Q(n4245) );
  OR2X1 U10983 ( .IN1(n11253), .IN2(n11254), .Q(n11252) );
  AND2X1 U10984 ( .IN1(n11228), .IN2(n7967), .Q(n11254) );
  AND2X1 U10985 ( .IN1(n11255), .IN2(n11237), .Q(n11253) );
  AND2X1 U10986 ( .IN1(n11256), .IN2(n11239), .Q(n11255) );
  OR2X1 U10987 ( .IN1(n11257), .IN2(n11258), .Q(n4244) );
  OR2X1 U10988 ( .IN1(n11259), .IN2(n11260), .Q(n11258) );
  AND2X1 U10989 ( .IN1(n11228), .IN2(g1916), .Q(n11260) );
  AND2X1 U10990 ( .IN1(n11229), .IN2(n11261), .Q(n11259) );
  AND2X1 U10991 ( .IN1(n2289), .IN2(n11262), .Q(n11257) );
  OR2X1 U10992 ( .IN1(n11251), .IN2(n11263), .Q(n4243) );
  OR2X1 U10993 ( .IN1(n11264), .IN2(n11265), .Q(n11263) );
  AND2X1 U10994 ( .IN1(n11228), .IN2(n7964), .Q(n11265) );
  AND2X1 U10995 ( .IN1(n11266), .IN2(n11237), .Q(n11264) );
  AND2X1 U10996 ( .IN1(n11267), .IN2(n11239), .Q(n11266) );
  OR2X1 U10997 ( .IN1(n11268), .IN2(n11240), .Q(n11251) );
  AND2X1 U10998 ( .IN1(n2289), .IN2(n2302), .Q(n11268) );
  OR2X1 U10999 ( .IN1(n11240), .IN2(n11269), .Q(n4242) );
  OR2X1 U11000 ( .IN1(n11270), .IN2(n11271), .Q(n11269) );
  AND2X1 U11001 ( .IN1(n11228), .IN2(n7963), .Q(n11271) );
  AND2X1 U11002 ( .IN1(n11272), .IN2(n11237), .Q(n11228) );
  AND2X1 U11003 ( .IN1(n11229), .IN2(n11273), .Q(n11270) );
  AND2X1 U11004 ( .IN1(n11239), .IN2(n11237), .Q(n11229) );
  INVX0 U11005 ( .INP(n11274), .ZN(n11239) );
  INVX0 U11006 ( .INP(n2275), .ZN(n11240) );
  OR2X1 U11007 ( .IN1(n11275), .IN2(n11276), .Q(n4241) );
  OR2X1 U11008 ( .IN1(n11277), .IN2(n11278), .Q(n11276) );
  AND2X1 U11009 ( .IN1(n11279), .IN2(g1890), .Q(n11278) );
  OR2X1 U11010 ( .IN1(n11280), .IN2(n11281), .Q(n11279) );
  INVX0 U11011 ( .INP(n11282), .ZN(n11281) );
  OR2X1 U11012 ( .IN1(n11283), .IN2(n11284), .Q(n11282) );
  AND2X1 U11013 ( .IN1(n11284), .IN2(n11283), .Q(n11280) );
  AND2X1 U11014 ( .IN1(n11285), .IN2(n11286), .Q(n11283) );
  INVX0 U11015 ( .INP(n11287), .ZN(n11286) );
  AND2X1 U11016 ( .IN1(n11288), .IN2(n11289), .Q(n11287) );
  OR2X1 U11017 ( .IN1(n11289), .IN2(n11288), .Q(n11285) );
  OR2X1 U11018 ( .IN1(n11290), .IN2(n11291), .Q(n11288) );
  AND2X1 U11019 ( .IN1(n11292), .IN2(n11267), .Q(n11291) );
  INVX0 U11020 ( .INP(n11293), .ZN(n11290) );
  OR2X1 U11021 ( .IN1(n11267), .IN2(n11292), .Q(n11293) );
  INVX0 U11022 ( .INP(n11273), .ZN(n11292) );
  OR2X1 U11023 ( .IN1(n11294), .IN2(n11295), .Q(n11273) );
  OR2X1 U11024 ( .IN1(n11296), .IN2(n11297), .Q(n11295) );
  AND2X1 U11025 ( .IN1(n11298), .IN2(n11299), .Q(n11297) );
  AND2X1 U11026 ( .IN1(n11300), .IN2(n11301), .Q(n11296) );
  OR2X1 U11027 ( .IN1(n11302), .IN2(n11303), .Q(n11267) );
  OR2X1 U11028 ( .IN1(n11304), .IN2(n11305), .Q(n11303) );
  AND2X1 U11029 ( .IN1(n11306), .IN2(n11307), .Q(n11305) );
  AND2X1 U11030 ( .IN1(n11308), .IN2(n11309), .Q(n11304) );
  AND2X1 U11031 ( .IN1(n11310), .IN2(n11311), .Q(n11289) );
  INVX0 U11032 ( .INP(n11312), .ZN(n11311) );
  AND2X1 U11033 ( .IN1(n11313), .IN2(n11256), .Q(n11312) );
  OR2X1 U11034 ( .IN1(n11256), .IN2(n11313), .Q(n11310) );
  INVX0 U11035 ( .INP(n11261), .ZN(n11313) );
  OR2X1 U11036 ( .IN1(n11294), .IN2(n11314), .Q(n11261) );
  OR2X1 U11037 ( .IN1(n11315), .IN2(n11316), .Q(n11314) );
  AND2X1 U11038 ( .IN1(n11317), .IN2(n11299), .Q(n11316) );
  AND2X1 U11039 ( .IN1(n11300), .IN2(n11318), .Q(n11315) );
  OR2X1 U11040 ( .IN1(n11302), .IN2(n11319), .Q(n11256) );
  OR2X1 U11041 ( .IN1(n11320), .IN2(n11321), .Q(n11319) );
  AND2X1 U11042 ( .IN1(n11322), .IN2(n11299), .Q(n11321) );
  AND2X1 U11043 ( .IN1(n11300), .IN2(n11323), .Q(n11320) );
  OR2X1 U11044 ( .IN1(n11324), .IN2(n11325), .Q(n11284) );
  INVX0 U11045 ( .INP(n11326), .ZN(n11325) );
  OR2X1 U11046 ( .IN1(n11327), .IN2(n11328), .Q(n11326) );
  AND2X1 U11047 ( .IN1(n11328), .IN2(n11327), .Q(n11324) );
  AND2X1 U11048 ( .IN1(n11329), .IN2(n11330), .Q(n11327) );
  INVX0 U11049 ( .INP(n11331), .ZN(n11330) );
  AND2X1 U11050 ( .IN1(n11332), .IN2(n11244), .Q(n11331) );
  OR2X1 U11051 ( .IN1(n11244), .IN2(n11332), .Q(n11329) );
  INVX0 U11052 ( .INP(n11250), .ZN(n11332) );
  OR2X1 U11053 ( .IN1(n11302), .IN2(n11333), .Q(n11250) );
  OR2X1 U11054 ( .IN1(n11334), .IN2(n11335), .Q(n11333) );
  AND2X1 U11055 ( .IN1(n11336), .IN2(n11299), .Q(n11335) );
  AND2X1 U11056 ( .IN1(n11300), .IN2(n11337), .Q(n11334) );
  OR2X1 U11057 ( .IN1(n11338), .IN2(n11339), .Q(n11244) );
  OR2X1 U11058 ( .IN1(n11340), .IN2(n11341), .Q(n11338) );
  AND2X1 U11059 ( .IN1(n11306), .IN2(n11342), .Q(n11341) );
  AND2X1 U11060 ( .IN1(n11343), .IN2(n11309), .Q(n11340) );
  OR2X1 U11061 ( .IN1(n11344), .IN2(n11345), .Q(n11328) );
  AND2X1 U11062 ( .IN1(n11346), .IN2(n11230), .Q(n11345) );
  INVX0 U11063 ( .INP(n11238), .ZN(n11346) );
  AND2X1 U11064 ( .IN1(n11347), .IN2(n11238), .Q(n11344) );
  OR2X1 U11065 ( .IN1(n11302), .IN2(n11348), .Q(n11238) );
  OR2X1 U11066 ( .IN1(n11349), .IN2(n11350), .Q(n11348) );
  AND2X1 U11067 ( .IN1(n11306), .IN2(n11351), .Q(n11350) );
  AND2X1 U11068 ( .IN1(n11352), .IN2(n11309), .Q(n11349) );
  INVX0 U11069 ( .INP(n11230), .ZN(n11347) );
  OR2X1 U11070 ( .IN1(n11302), .IN2(n11353), .Q(n11230) );
  OR2X1 U11071 ( .IN1(n11354), .IN2(n11355), .Q(n11353) );
  AND2X1 U11072 ( .IN1(n11306), .IN2(n11356), .Q(n11355) );
  AND2X1 U11073 ( .IN1(n11357), .IN2(n11309), .Q(n11354) );
  AND2X1 U11074 ( .IN1(n11358), .IN2(n11359), .Q(n11277) );
  AND2X1 U11075 ( .IN1(n11360), .IN2(n11361), .Q(n11359) );
  OR2X1 U11076 ( .IN1(test_so69), .IN2(n10974), .Q(n11361) );
  OR2X1 U11077 ( .IN1(g3229), .IN2(n7960), .Q(n11360) );
  AND2X1 U11078 ( .IN1(n11274), .IN2(n11237), .Q(n11358) );
  INVX0 U11079 ( .INP(n11362), .ZN(n11237) );
  AND2X1 U11080 ( .IN1(n11272), .IN2(n580), .Q(n11274) );
  INVX0 U11081 ( .INP(n11363), .ZN(n580) );
  AND2X1 U11082 ( .IN1(n11364), .IN2(g1937), .Q(n11275) );
  OR2X1 U11083 ( .IN1(n11365), .IN2(n11366), .Q(n11364) );
  INVX0 U11084 ( .INP(n11367), .ZN(n11366) );
  OR2X1 U11085 ( .IN1(n11262), .IN2(n11368), .Q(n11367) );
  AND2X1 U11086 ( .IN1(n11368), .IN2(n11262), .Q(n11365) );
  OR2X1 U11087 ( .IN1(n11294), .IN2(n11369), .Q(n11262) );
  OR2X1 U11088 ( .IN1(n11370), .IN2(n11371), .Q(n11369) );
  AND2X1 U11089 ( .IN1(n11372), .IN2(n11299), .Q(n11371) );
  AND2X1 U11090 ( .IN1(n11300), .IN2(n11373), .Q(n11370) );
  AND2X1 U11091 ( .IN1(n11374), .IN2(n11375), .Q(n11300) );
  OR2X1 U11092 ( .IN1(n11376), .IN2(n11302), .Q(n11294) );
  INVX0 U11093 ( .INP(n2279), .ZN(n11376) );
  INVX0 U11094 ( .INP(n11231), .ZN(n11368) );
  OR2X1 U11095 ( .IN1(n11377), .IN2(n11339), .Q(n11231) );
  OR2X1 U11096 ( .IN1(n11378), .IN2(n11302), .Q(n11339) );
  OR2X1 U11097 ( .IN1(n4545), .IN2(n11363), .Q(n11302) );
  OR2X1 U11098 ( .IN1(g1939), .IN2(n11379), .Q(n11363) );
  OR2X1 U11099 ( .IN1(g1943), .IN2(n608), .Q(n11379) );
  INVX0 U11100 ( .INP(n2309), .ZN(n11378) );
  OR2X1 U11101 ( .IN1(n11380), .IN2(n11381), .Q(n11377) );
  AND2X1 U11102 ( .IN1(n11306), .IN2(n11382), .Q(n11381) );
  AND2X1 U11103 ( .IN1(n11374), .IN2(n11383), .Q(n11306) );
  AND2X1 U11104 ( .IN1(n11384), .IN2(n11309), .Q(n11380) );
  OR2X1 U11105 ( .IN1(n11385), .IN2(n11386), .Q(n4240) );
  OR2X1 U11106 ( .IN1(n11387), .IN2(n11388), .Q(n11386) );
  AND2X1 U11107 ( .IN1(n11389), .IN2(g1223), .Q(n11388) );
  AND2X1 U11108 ( .IN1(n11390), .IN2(n11391), .Q(n11387) );
  AND2X1 U11109 ( .IN1(n2217), .IN2(n11392), .Q(n11385) );
  OR2X1 U11110 ( .IN1(n11393), .IN2(n11394), .Q(n4239) );
  OR2X1 U11111 ( .IN1(n11395), .IN2(n11396), .Q(n11394) );
  AND2X1 U11112 ( .IN1(n11389), .IN2(n8007), .Q(n11395) );
  OR2X1 U11113 ( .IN1(n11397), .IN2(n11398), .Q(n11393) );
  AND2X1 U11114 ( .IN1(n11399), .IN2(n11400), .Q(n11398) );
  AND2X1 U11115 ( .IN1(n11401), .IN2(n11402), .Q(n11399) );
  OR2X1 U11116 ( .IN1(n11403), .IN2(n11404), .Q(n4238) );
  OR2X1 U11117 ( .IN1(n11397), .IN2(n11405), .Q(n11404) );
  AND2X1 U11118 ( .IN1(n11390), .IN2(n11406), .Q(n11405) );
  AND2X1 U11119 ( .IN1(n11389), .IN2(n8003), .Q(n11403) );
  OR2X1 U11120 ( .IN1(n11407), .IN2(n11408), .Q(n4237) );
  OR2X1 U11121 ( .IN1(n11409), .IN2(n11396), .Q(n11408) );
  INVX0 U11122 ( .INP(n2231), .ZN(n11396) );
  AND2X1 U11123 ( .IN1(n11389), .IN2(n8006), .Q(n11409) );
  OR2X1 U11124 ( .IN1(n11397), .IN2(n11410), .Q(n11407) );
  AND2X1 U11125 ( .IN1(n11411), .IN2(n11400), .Q(n11410) );
  AND2X1 U11126 ( .IN1(n11412), .IN2(n11402), .Q(n11411) );
  OR2X1 U11127 ( .IN1(n11413), .IN2(n11414), .Q(n4236) );
  OR2X1 U11128 ( .IN1(n11415), .IN2(n11416), .Q(n11414) );
  AND2X1 U11129 ( .IN1(n11389), .IN2(n8008), .Q(n11416) );
  AND2X1 U11130 ( .IN1(n11417), .IN2(n11400), .Q(n11415) );
  AND2X1 U11131 ( .IN1(n11418), .IN2(n11402), .Q(n11417) );
  OR2X1 U11132 ( .IN1(n11419), .IN2(n11420), .Q(n4235) );
  OR2X1 U11133 ( .IN1(n11421), .IN2(n11422), .Q(n11420) );
  AND2X1 U11134 ( .IN1(n11389), .IN2(g1222), .Q(n11422) );
  AND2X1 U11135 ( .IN1(n11390), .IN2(n11423), .Q(n11421) );
  AND2X1 U11136 ( .IN1(n2217), .IN2(n11424), .Q(n11419) );
  OR2X1 U11137 ( .IN1(n11413), .IN2(n11425), .Q(n4234) );
  OR2X1 U11138 ( .IN1(n11426), .IN2(n11427), .Q(n11425) );
  AND2X1 U11139 ( .IN1(n11389), .IN2(n8005), .Q(n11427) );
  AND2X1 U11140 ( .IN1(n11428), .IN2(n11400), .Q(n11426) );
  AND2X1 U11141 ( .IN1(n11429), .IN2(n11402), .Q(n11428) );
  OR2X1 U11142 ( .IN1(n11397), .IN2(n11430), .Q(n11413) );
  AND2X1 U11143 ( .IN1(n2217), .IN2(n2230), .Q(n11430) );
  OR2X1 U11144 ( .IN1(n11431), .IN2(n11432), .Q(n4233) );
  OR2X1 U11145 ( .IN1(n11397), .IN2(n11433), .Q(n11432) );
  AND2X1 U11146 ( .IN1(n11390), .IN2(n11434), .Q(n11433) );
  AND2X1 U11147 ( .IN1(n11402), .IN2(n11400), .Q(n11390) );
  AND2X1 U11148 ( .IN1(n11435), .IN2(n2217), .Q(n11397) );
  AND2X1 U11149 ( .IN1(n11389), .IN2(n8004), .Q(n11431) );
  AND2X1 U11150 ( .IN1(n11436), .IN2(n11400), .Q(n11389) );
  OR2X1 U11151 ( .IN1(n11437), .IN2(n11438), .Q(n4232) );
  OR2X1 U11152 ( .IN1(n11439), .IN2(n11440), .Q(n11438) );
  AND2X1 U11153 ( .IN1(n11441), .IN2(g1196), .Q(n11440) );
  OR2X1 U11154 ( .IN1(n11442), .IN2(n11443), .Q(n11441) );
  INVX0 U11155 ( .INP(n11444), .ZN(n11443) );
  OR2X1 U11156 ( .IN1(n11445), .IN2(n11446), .Q(n11444) );
  AND2X1 U11157 ( .IN1(n11446), .IN2(n11445), .Q(n11442) );
  AND2X1 U11158 ( .IN1(n11447), .IN2(n11448), .Q(n11445) );
  INVX0 U11159 ( .INP(n11449), .ZN(n11448) );
  AND2X1 U11160 ( .IN1(n11450), .IN2(n11451), .Q(n11449) );
  OR2X1 U11161 ( .IN1(n11451), .IN2(n11450), .Q(n11447) );
  OR2X1 U11162 ( .IN1(n11452), .IN2(n11453), .Q(n11450) );
  AND2X1 U11163 ( .IN1(n11454), .IN2(n11429), .Q(n11453) );
  INVX0 U11164 ( .INP(n11455), .ZN(n11452) );
  OR2X1 U11165 ( .IN1(n11429), .IN2(n11454), .Q(n11455) );
  INVX0 U11166 ( .INP(n11434), .ZN(n11454) );
  OR2X1 U11167 ( .IN1(n11456), .IN2(n11457), .Q(n11434) );
  OR2X1 U11168 ( .IN1(n11458), .IN2(n11459), .Q(n11457) );
  AND2X1 U11169 ( .IN1(n11460), .IN2(n11461), .Q(n11459) );
  AND2X1 U11170 ( .IN1(n11462), .IN2(n11463), .Q(n11458) );
  OR2X1 U11171 ( .IN1(n11464), .IN2(n11465), .Q(n11429) );
  OR2X1 U11172 ( .IN1(n11466), .IN2(n11467), .Q(n11465) );
  AND2X1 U11173 ( .IN1(n11468), .IN2(n11469), .Q(n11467) );
  AND2X1 U11174 ( .IN1(n11470), .IN2(n11471), .Q(n11466) );
  AND2X1 U11175 ( .IN1(n11472), .IN2(n11473), .Q(n11451) );
  INVX0 U11176 ( .INP(n11474), .ZN(n11473) );
  AND2X1 U11177 ( .IN1(n11475), .IN2(n11418), .Q(n11474) );
  OR2X1 U11178 ( .IN1(n11418), .IN2(n11475), .Q(n11472) );
  INVX0 U11179 ( .INP(n11423), .ZN(n11475) );
  OR2X1 U11180 ( .IN1(n11456), .IN2(n11476), .Q(n11423) );
  OR2X1 U11181 ( .IN1(n11477), .IN2(n11478), .Q(n11476) );
  AND2X1 U11182 ( .IN1(n11479), .IN2(n11461), .Q(n11478) );
  AND2X1 U11183 ( .IN1(n11462), .IN2(n11480), .Q(n11477) );
  OR2X1 U11184 ( .IN1(n11464), .IN2(n11481), .Q(n11418) );
  OR2X1 U11185 ( .IN1(n11482), .IN2(n11483), .Q(n11481) );
  AND2X1 U11186 ( .IN1(n11484), .IN2(n11461), .Q(n11483) );
  AND2X1 U11187 ( .IN1(n11462), .IN2(n11485), .Q(n11482) );
  OR2X1 U11188 ( .IN1(n11486), .IN2(n11487), .Q(n11446) );
  INVX0 U11189 ( .INP(n11488), .ZN(n11487) );
  OR2X1 U11190 ( .IN1(n11489), .IN2(n11490), .Q(n11488) );
  AND2X1 U11191 ( .IN1(n11490), .IN2(n11489), .Q(n11486) );
  AND2X1 U11192 ( .IN1(n11491), .IN2(n11492), .Q(n11489) );
  INVX0 U11193 ( .INP(n11493), .ZN(n11492) );
  AND2X1 U11194 ( .IN1(n11494), .IN2(n11406), .Q(n11493) );
  OR2X1 U11195 ( .IN1(n11406), .IN2(n11494), .Q(n11491) );
  INVX0 U11196 ( .INP(n11412), .ZN(n11494) );
  OR2X1 U11197 ( .IN1(n11464), .IN2(n11495), .Q(n11412) );
  OR2X1 U11198 ( .IN1(n11496), .IN2(n11497), .Q(n11495) );
  AND2X1 U11199 ( .IN1(n11498), .IN2(n11461), .Q(n11497) );
  AND2X1 U11200 ( .IN1(n11462), .IN2(n11499), .Q(n11496) );
  OR2X1 U11201 ( .IN1(n11500), .IN2(n11501), .Q(n11406) );
  OR2X1 U11202 ( .IN1(n11502), .IN2(n11503), .Q(n11500) );
  AND2X1 U11203 ( .IN1(n11468), .IN2(n11504), .Q(n11503) );
  AND2X1 U11204 ( .IN1(n11505), .IN2(n11471), .Q(n11502) );
  OR2X1 U11205 ( .IN1(n11506), .IN2(n11507), .Q(n11490) );
  AND2X1 U11206 ( .IN1(n11508), .IN2(n11391), .Q(n11507) );
  INVX0 U11207 ( .INP(n11401), .ZN(n11508) );
  AND2X1 U11208 ( .IN1(n11509), .IN2(n11401), .Q(n11506) );
  OR2X1 U11209 ( .IN1(n11464), .IN2(n11510), .Q(n11401) );
  OR2X1 U11210 ( .IN1(n11511), .IN2(n11512), .Q(n11510) );
  AND2X1 U11211 ( .IN1(n11468), .IN2(n11513), .Q(n11512) );
  AND2X1 U11212 ( .IN1(n11514), .IN2(n11471), .Q(n11511) );
  INVX0 U11213 ( .INP(n11391), .ZN(n11509) );
  OR2X1 U11214 ( .IN1(n11464), .IN2(n11515), .Q(n11391) );
  OR2X1 U11215 ( .IN1(n11516), .IN2(n11517), .Q(n11515) );
  AND2X1 U11216 ( .IN1(n11468), .IN2(n11518), .Q(n11517) );
  AND2X1 U11217 ( .IN1(n11519), .IN2(n11471), .Q(n11516) );
  AND2X1 U11218 ( .IN1(n11520), .IN2(n11521), .Q(n11439) );
  AND2X1 U11219 ( .IN1(n11522), .IN2(n11523), .Q(n11521) );
  OR2X1 U11220 ( .IN1(n10974), .IN2(g1224), .Q(n11523) );
  OR2X1 U11221 ( .IN1(test_so48), .IN2(g3229), .Q(n11522) );
  AND2X1 U11222 ( .IN1(n11524), .IN2(n11400), .Q(n11520) );
  INVX0 U11223 ( .INP(n11525), .ZN(n11400) );
  INVX0 U11224 ( .INP(n11402), .ZN(n11524) );
  OR2X1 U11225 ( .IN1(n11435), .IN2(n11526), .Q(n11402) );
  AND2X1 U11226 ( .IN1(n11527), .IN2(g1243), .Q(n11437) );
  OR2X1 U11227 ( .IN1(n11528), .IN2(n11529), .Q(n11527) );
  INVX0 U11228 ( .INP(n11530), .ZN(n11529) );
  OR2X1 U11229 ( .IN1(n11424), .IN2(n11531), .Q(n11530) );
  AND2X1 U11230 ( .IN1(n11531), .IN2(n11424), .Q(n11528) );
  OR2X1 U11231 ( .IN1(n11456), .IN2(n11532), .Q(n11424) );
  OR2X1 U11232 ( .IN1(n11533), .IN2(n11534), .Q(n11532) );
  AND2X1 U11233 ( .IN1(n11535), .IN2(n11461), .Q(n11534) );
  AND2X1 U11234 ( .IN1(n11462), .IN2(n11536), .Q(n11533) );
  AND2X1 U11235 ( .IN1(n11537), .IN2(n11538), .Q(n11462) );
  OR2X1 U11236 ( .IN1(n11539), .IN2(n11464), .Q(n11456) );
  INVX0 U11237 ( .INP(n2207), .ZN(n11539) );
  INVX0 U11238 ( .INP(n11392), .ZN(n11531) );
  OR2X1 U11239 ( .IN1(n11540), .IN2(n11501), .Q(n11392) );
  OR2X1 U11240 ( .IN1(n11541), .IN2(n11464), .Q(n11501) );
  OR2X1 U11241 ( .IN1(n4548), .IN2(n11435), .Q(n11464) );
  OR2X1 U11242 ( .IN1(g1245), .IN2(n11542), .Q(n11435) );
  OR2X1 U11243 ( .IN1(g1249), .IN2(n578), .Q(n11542) );
  INVX0 U11244 ( .INP(n2237), .ZN(n11541) );
  OR2X1 U11245 ( .IN1(n11543), .IN2(n11544), .Q(n11540) );
  AND2X1 U11246 ( .IN1(n11468), .IN2(n11545), .Q(n11544) );
  AND2X1 U11247 ( .IN1(n11537), .IN2(n11546), .Q(n11468) );
  AND2X1 U11248 ( .IN1(n11547), .IN2(n11471), .Q(n11543) );
  INVX0 U11249 ( .INP(n11548), .ZN(n375) );
  OR2X1 U11250 ( .IN1(n10184), .IN2(n11549), .Q(n4528) );
  INVX0 U11251 ( .INP(n3896), .ZN(n11549) );
  OR2X1 U11252 ( .IN1(n10185), .IN2(n11550), .Q(n4527) );
  INVX0 U11253 ( .INP(n3890), .ZN(n11550) );
  OR2X1 U11254 ( .IN1(n10186), .IN2(n11551), .Q(n4523) );
  INVX0 U11255 ( .INP(n3686), .ZN(n11551) );
  OR2X1 U11256 ( .IN1(n10187), .IN2(n11552), .Q(n4522) );
  INVX0 U11257 ( .INP(n3683), .ZN(n11552) );
  INVX0 U11258 ( .INP(g24734), .ZN(n330) );
  INVX0 U11259 ( .INP(g25435), .ZN(n326) );
  OR2X1 U11260 ( .IN1(n11553), .IN2(n11554), .Q(n3254) );
  AND2X1 U11261 ( .IN1(n11555), .IN2(n11556), .Q(n11554) );
  INVX0 U11262 ( .INP(n11557), .ZN(n11555) );
  INVX0 U11263 ( .INP(g26135), .ZN(n300) );
  INVX0 U11264 ( .INP(n11558), .ZN(n29) );
  OR2X1 U11265 ( .IN1(n11559), .IN2(n11560), .Q(n2800) );
  AND2X1 U11266 ( .IN1(n11561), .IN2(n11562), .Q(n11560) );
  AND2X1 U11267 ( .IN1(n11563), .IN2(n11564), .Q(n11561) );
  AND2X1 U11268 ( .IN1(n11565), .IN2(n11566), .Q(n11559) );
  INVX0 U11269 ( .INP(n11563), .ZN(n11565) );
  OR2X1 U11270 ( .IN1(n11567), .IN2(n11568), .Q(n11563) );
  OR2X1 U11271 ( .IN1(n11569), .IN2(n11570), .Q(n11568) );
  AND2X1 U11272 ( .IN1(n11571), .IN2(n11566), .Q(n11570) );
  OR2X1 U11273 ( .IN1(n11572), .IN2(n11573), .Q(n11567) );
  AND2X1 U11274 ( .IN1(n11574), .IN2(n11575), .Q(n11573) );
  AND2X1 U11275 ( .IN1(n11576), .IN2(n11577), .Q(n11574) );
  OR2X1 U11276 ( .IN1(n11578), .IN2(n11579), .Q(n11576) );
  AND2X1 U11277 ( .IN1(n11562), .IN2(n11580), .Q(n11578) );
  AND2X1 U11278 ( .IN1(n11581), .IN2(n11582), .Q(n11572) );
  OR2X1 U11279 ( .IN1(n4387), .IN2(n11583), .Q(n11582) );
  OR2X1 U11280 ( .IN1(n11584), .IN2(n11585), .Q(n2719) );
  AND2X1 U11281 ( .IN1(n11586), .IN2(n10651), .Q(n11585) );
  AND2X1 U11282 ( .IN1(n10650), .IN2(n11587), .Q(n11584) );
  OR2X1 U11283 ( .IN1(n11588), .IN2(n11589), .Q(n2686) );
  AND2X1 U11284 ( .IN1(n4530), .IN2(n10794), .Q(n11589) );
  AND2X1 U11285 ( .IN1(n10793), .IN2(n11590), .Q(n11588) );
  OR2X1 U11286 ( .IN1(n11591), .IN2(n11592), .Q(n2671) );
  AND2X1 U11287 ( .IN1(n4529), .IN2(n10837), .Q(n11592) );
  AND2X1 U11288 ( .IN1(n10836), .IN2(n11593), .Q(n11591) );
  OR2X1 U11289 ( .IN1(n11594), .IN2(n11595), .Q(n2616) );
  AND2X1 U11290 ( .IN1(n11596), .IN2(n11575), .Q(n11595) );
  INVX0 U11291 ( .INP(n11597), .ZN(n11596) );
  AND2X1 U11292 ( .IN1(n11581), .IN2(n11597), .Q(n11594) );
  OR2X1 U11293 ( .IN1(n11598), .IN2(n11599), .Q(n11597) );
  OR2X1 U11294 ( .IN1(n11600), .IN2(n11601), .Q(n11599) );
  AND2X1 U11295 ( .IN1(n11602), .IN2(n11581), .Q(n11601) );
  AND2X1 U11296 ( .IN1(n11603), .IN2(n11577), .Q(n11602) );
  AND2X1 U11297 ( .IN1(n11604), .IN2(n11605), .Q(n11603) );
  OR2X1 U11298 ( .IN1(n11562), .IN2(n11606), .Q(n11605) );
  OR2X1 U11299 ( .IN1(n11607), .IN2(n11566), .Q(n11604) );
  AND2X1 U11300 ( .IN1(n11608), .IN2(n11609), .Q(n11607) );
  AND2X1 U11301 ( .IN1(n11610), .IN2(n11564), .Q(n11609) );
  AND2X1 U11302 ( .IN1(n11611), .IN2(n11612), .Q(n11608) );
  OR2X1 U11303 ( .IN1(n11579), .IN2(n11580), .Q(n11612) );
  AND2X1 U11304 ( .IN1(n11613), .IN2(n11575), .Q(n11600) );
  OR2X1 U11305 ( .IN1(n11614), .IN2(n11579), .Q(n11613) );
  AND2X1 U11306 ( .IN1(n11615), .IN2(n11616), .Q(n11614) );
  INVX0 U11307 ( .INP(n11617), .ZN(n11616) );
  AND2X1 U11308 ( .IN1(n11618), .IN2(n11619), .Q(n11615) );
  INVX0 U11309 ( .INP(n11620), .ZN(n11619) );
  OR2X1 U11310 ( .IN1(n11566), .IN2(n11621), .Q(n11618) );
  OR2X1 U11311 ( .IN1(n11622), .IN2(n11623), .Q(n11621) );
  AND2X1 U11312 ( .IN1(n11569), .IN2(n11624), .Q(n11598) );
  OR2X1 U11313 ( .IN1(n11058), .IN2(n11045), .Q(n2459) );
  AND2X1 U11314 ( .IN1(n10975), .IN2(n10926), .Q(n2446) );
  INVX0 U11315 ( .INP(n11625), .ZN(n10926) );
  OR2X1 U11316 ( .IN1(n11626), .IN2(test_so22), .Q(n11625) );
  AND2X1 U11317 ( .IN1(n4360), .IN2(n9898), .Q(n11626) );
  OR2X1 U11318 ( .IN1(n11627), .IN2(g557), .Q(n10975) );
  AND2X1 U11319 ( .IN1(n9898), .IN2(n10200), .Q(n11627) );
  OR2X1 U11320 ( .IN1(n11628), .IN2(n4541), .Q(n2445) );
  AND2X1 U11321 ( .IN1(n11629), .IN2(n11630), .Q(n11628) );
  AND2X1 U11322 ( .IN1(n11631), .IN2(n11045), .Q(n11630) );
  OR2X1 U11323 ( .IN1(n11632), .IN2(n11633), .Q(n11045) );
  OR2X1 U11324 ( .IN1(n11634), .IN2(n11635), .Q(n11633) );
  OR2X1 U11325 ( .IN1(n11030), .IN2(n11636), .Q(n11635) );
  OR2X1 U11326 ( .IN1(n11001), .IN2(n11034), .Q(n11636) );
  OR2X1 U11327 ( .IN1(n11011), .IN2(n11637), .Q(n11634) );
  OR2X1 U11328 ( .IN1(n11638), .IN2(n11015), .Q(n11637) );
  AND2X1 U11329 ( .IN1(n11639), .IN2(n11640), .Q(n11638) );
  OR2X1 U11330 ( .IN1(n4295), .IN2(g737), .Q(n11640) );
  AND2X1 U11331 ( .IN1(n11641), .IN2(n11642), .Q(n11639) );
  OR2X1 U11332 ( .IN1(n4359), .IN2(g739), .Q(n11642) );
  OR2X1 U11333 ( .IN1(n4309), .IN2(g738), .Q(n11641) );
  OR2X1 U11334 ( .IN1(n11643), .IN2(n11644), .Q(n11632) );
  OR2X1 U11335 ( .IN1(n11645), .IN2(n11646), .Q(n11644) );
  OR2X1 U11336 ( .IN1(n10966), .IN2(n10960), .Q(n11646) );
  INVX0 U11337 ( .INP(n10959), .ZN(n10960) );
  INVX0 U11338 ( .INP(n10969), .ZN(n10966) );
  INVX0 U11339 ( .INP(n11647), .ZN(n11645) );
  OR2X1 U11340 ( .IN1(n10995), .IN2(n11648), .Q(n11643) );
  OR2X1 U11341 ( .IN1(n11059), .IN2(n11043), .Q(n11648) );
  OR2X1 U11342 ( .IN1(n4359), .IN2(g736), .Q(n11631) );
  AND2X1 U11343 ( .IN1(n11649), .IN2(n11650), .Q(n11629) );
  OR2X1 U11344 ( .IN1(n4309), .IN2(g735), .Q(n11650) );
  OR2X1 U11345 ( .IN1(n4295), .IN2(g734), .Q(n11649) );
  OR2X1 U11346 ( .IN1(n11222), .IN2(n11212), .Q(n2381) );
  OR2X1 U11347 ( .IN1(n11651), .IN2(n4543), .Q(n2374) );
  AND2X1 U11348 ( .IN1(n11652), .IN2(n11653), .Q(n11651) );
  AND2X1 U11349 ( .IN1(n11654), .IN2(n11212), .Q(n11653) );
  OR2X1 U11350 ( .IN1(n11655), .IN2(n11656), .Q(n11212) );
  OR2X1 U11351 ( .IN1(n11657), .IN2(n11658), .Q(n11656) );
  OR2X1 U11352 ( .IN1(n11193), .IN2(n11659), .Q(n11658) );
  OR2X1 U11353 ( .IN1(n11144), .IN2(n11160), .Q(n11659) );
  OR2X1 U11354 ( .IN1(n11174), .IN2(n11660), .Q(n11657) );
  OR2X1 U11355 ( .IN1(n11661), .IN2(n11188), .Q(n11660) );
  AND2X1 U11356 ( .IN1(n11662), .IN2(n11663), .Q(n11661) );
  OR2X1 U11357 ( .IN1(n4292), .IN2(test_so95), .Q(n11663) );
  AND2X1 U11358 ( .IN1(n11664), .IN2(n11665), .Q(n11662) );
  OR2X1 U11359 ( .IN1(n4356), .IN2(g2813), .Q(n11665) );
  OR2X1 U11360 ( .IN1(n4306), .IN2(g2812), .Q(n11664) );
  OR2X1 U11361 ( .IN1(n11666), .IN2(n11667), .Q(n11655) );
  OR2X1 U11362 ( .IN1(n11668), .IN2(n11669), .Q(n11667) );
  OR2X1 U11363 ( .IN1(n11210), .IN2(n11223), .Q(n11669) );
  INVX0 U11364 ( .INP(n11221), .ZN(n11223) );
  INVX0 U11365 ( .INP(n11211), .ZN(n11210) );
  INVX0 U11366 ( .INP(n11670), .ZN(n11668) );
  OR2X1 U11367 ( .IN1(n11135), .IN2(n11671), .Q(n11666) );
  OR2X1 U11368 ( .IN1(n11180), .IN2(n11154), .Q(n11671) );
  OR2X1 U11369 ( .IN1(n4356), .IN2(g2810), .Q(n11654) );
  AND2X1 U11370 ( .IN1(n11672), .IN2(n11673), .Q(n11652) );
  OR2X1 U11371 ( .IN1(n4306), .IN2(g2809), .Q(n11673) );
  OR2X1 U11372 ( .IN1(n4292), .IN2(g2808), .Q(n11672) );
  AND2X1 U11373 ( .IN1(n11200), .IN2(n11111), .Q(n2361) );
  INVX0 U11374 ( .INP(n11201), .ZN(n11111) );
  OR2X1 U11375 ( .IN1(n11674), .IN2(g2584), .Q(n11201) );
  AND2X1 U11376 ( .IN1(n4352), .IN2(n9895), .Q(n11674) );
  OR2X1 U11377 ( .IN1(n11675), .IN2(g2631), .Q(n11200) );
  AND2X1 U11378 ( .IN1(n9895), .IN2(n4303), .Q(n11675) );
  OR2X1 U11379 ( .IN1(n11383), .IN2(n11374), .Q(n2309) );
  OR2X1 U11380 ( .IN1(n11676), .IN2(n4545), .Q(n2302) );
  AND2X1 U11381 ( .IN1(n11677), .IN2(n11678), .Q(n11676) );
  AND2X1 U11382 ( .IN1(n11679), .IN2(n11374), .Q(n11678) );
  OR2X1 U11383 ( .IN1(n4357), .IN2(g2116), .Q(n11679) );
  AND2X1 U11384 ( .IN1(n11680), .IN2(n11681), .Q(n11677) );
  OR2X1 U11385 ( .IN1(n4307), .IN2(g2115), .Q(n11681) );
  OR2X1 U11386 ( .IN1(n4293), .IN2(g2114), .Q(n11680) );
  AND2X1 U11387 ( .IN1(n11362), .IN2(n11272), .Q(n2289) );
  AND2X1 U11388 ( .IN1(n11682), .IN2(n4297), .Q(n11272) );
  OR2X1 U11389 ( .IN1(g1905), .IN2(g1937), .Q(n11682) );
  OR2X1 U11390 ( .IN1(n11683), .IN2(g1937), .Q(n11362) );
  AND2X1 U11391 ( .IN1(n4297), .IN2(n9896), .Q(n11683) );
  OR2X1 U11392 ( .IN1(n11375), .IN2(n11374), .Q(n2279) );
  OR2X1 U11393 ( .IN1(n11684), .IN2(n11685), .Q(n11374) );
  OR2X1 U11394 ( .IN1(n11686), .IN2(n11687), .Q(n11685) );
  OR2X1 U11395 ( .IN1(n11356), .IN2(n11688), .Q(n11687) );
  OR2X1 U11396 ( .IN1(n11323), .IN2(n11307), .Q(n11688) );
  OR2X1 U11397 ( .IN1(n11351), .IN2(n11689), .Q(n11686) );
  OR2X1 U11398 ( .IN1(n11690), .IN2(n11337), .Q(n11689) );
  AND2X1 U11399 ( .IN1(n11691), .IN2(n11692), .Q(n11690) );
  OR2X1 U11400 ( .IN1(n4293), .IN2(g2117), .Q(n11692) );
  AND2X1 U11401 ( .IN1(n11693), .IN2(n11694), .Q(n11691) );
  OR2X1 U11402 ( .IN1(n4357), .IN2(g2119), .Q(n11694) );
  OR2X1 U11403 ( .IN1(n4307), .IN2(g2118), .Q(n11693) );
  OR2X1 U11404 ( .IN1(n11695), .IN2(n11696), .Q(n11684) );
  OR2X1 U11405 ( .IN1(n11697), .IN2(n11698), .Q(n11696) );
  OR2X1 U11406 ( .IN1(n11372), .IN2(n11384), .Q(n11698) );
  INVX0 U11407 ( .INP(n11699), .ZN(n11697) );
  OR2X1 U11408 ( .IN1(n11298), .IN2(n11700), .Q(n11695) );
  OR2X1 U11409 ( .IN1(n11343), .IN2(n11317), .Q(n11700) );
  OR2X1 U11410 ( .IN1(n11546), .IN2(n11537), .Q(n2237) );
  OR2X1 U11411 ( .IN1(n11701), .IN2(n4548), .Q(n2230) );
  AND2X1 U11412 ( .IN1(n11702), .IN2(n11703), .Q(n11701) );
  AND2X1 U11413 ( .IN1(n11704), .IN2(n11537), .Q(n11703) );
  OR2X1 U11414 ( .IN1(n4358), .IN2(g1422), .Q(n11704) );
  AND2X1 U11415 ( .IN1(n11705), .IN2(n11706), .Q(n11702) );
  OR2X1 U11416 ( .IN1(n4308), .IN2(g1421), .Q(n11706) );
  OR2X1 U11417 ( .IN1(n4294), .IN2(g1420), .Q(n11705) );
  AND2X1 U11418 ( .IN1(n11525), .IN2(n11436), .Q(n2217) );
  INVX0 U11419 ( .INP(n11526), .ZN(n11436) );
  OR2X1 U11420 ( .IN1(n11707), .IN2(g1196), .Q(n11526) );
  AND2X1 U11421 ( .IN1(n4353), .IN2(n9897), .Q(n11707) );
  OR2X1 U11422 ( .IN1(n11708), .IN2(g1243), .Q(n11525) );
  AND2X1 U11423 ( .IN1(n9897), .IN2(n4304), .Q(n11708) );
  OR2X1 U11424 ( .IN1(n11538), .IN2(n11537), .Q(n2207) );
  OR2X1 U11425 ( .IN1(n11709), .IN2(n11710), .Q(n11537) );
  OR2X1 U11426 ( .IN1(n11711), .IN2(n11712), .Q(n11710) );
  OR2X1 U11427 ( .IN1(n11518), .IN2(n11713), .Q(n11712) );
  OR2X1 U11428 ( .IN1(n11485), .IN2(n11469), .Q(n11713) );
  OR2X1 U11429 ( .IN1(n11513), .IN2(n11714), .Q(n11711) );
  OR2X1 U11430 ( .IN1(n11715), .IN2(n11499), .Q(n11714) );
  AND2X1 U11431 ( .IN1(n11716), .IN2(n11717), .Q(n11715) );
  OR2X1 U11432 ( .IN1(n4294), .IN2(g1423), .Q(n11717) );
  AND2X1 U11433 ( .IN1(n11718), .IN2(n11719), .Q(n11716) );
  OR2X1 U11434 ( .IN1(n4358), .IN2(g1425), .Q(n11719) );
  OR2X1 U11435 ( .IN1(n4308), .IN2(g1424), .Q(n11718) );
  OR2X1 U11436 ( .IN1(n11720), .IN2(n11721), .Q(n11709) );
  OR2X1 U11437 ( .IN1(n11722), .IN2(n11723), .Q(n11721) );
  OR2X1 U11438 ( .IN1(n11547), .IN2(n11535), .Q(n11723) );
  INVX0 U11439 ( .INP(n11724), .ZN(n11722) );
  OR2X1 U11440 ( .IN1(n11460), .IN2(n11725), .Q(n11720) );
  OR2X1 U11441 ( .IN1(n11505), .IN2(n11479), .Q(n11725) );
  OR2X1 U11442 ( .IN1(n11726), .IN2(n11727), .Q(n18) );
  OR2X1 U11443 ( .IN1(n11728), .IN2(n11729), .Q(n11727) );
  AND2X1 U11444 ( .IN1(n4330), .IN2(g2950), .Q(n11729) );
  AND2X1 U11445 ( .IN1(n4423), .IN2(g2883), .Q(n11728) );
  INVX0 U11446 ( .INP(n11730), .ZN(n11726) );
  INVX0 U11447 ( .INP(n11731), .ZN(n1669) );
  INVX0 U11448 ( .INP(n11732), .ZN(n1647) );
  INVX0 U11449 ( .INP(n11733), .ZN(n4526) );
  AND2X1 U11450 ( .IN1(test_so78), .IN2(n3887), .Q(n11733) );
  INVX0 U11451 ( .INP(n11734), .ZN(n1480) );
  INVX0 U11452 ( .INP(n11735), .ZN(n1330) );
  INVX0 U11453 ( .INP(n11736), .ZN(n1305) );
  INVX0 U11454 ( .INP(n11737), .ZN(n1136) );
  OR2X1 U11455 ( .IN1(n11738), .IN2(n11739), .Q(g30801) );
  AND2X1 U11456 ( .IN1(g30072), .IN2(g3109), .Q(n11739) );
  AND2X1 U11457 ( .IN1(n4494), .IN2(g3108), .Q(n11738) );
  OR2X1 U11458 ( .IN1(n11740), .IN2(n11741), .Q(g30798) );
  AND2X1 U11459 ( .IN1(g30072), .IN2(g8030), .Q(n11741) );
  AND2X1 U11460 ( .IN1(n4383), .IN2(g3107), .Q(n11740) );
  OR2X1 U11461 ( .IN1(n11742), .IN2(n11743), .Q(g30796) );
  AND2X1 U11462 ( .IN1(g30072), .IN2(g8106), .Q(n11743) );
  AND2X1 U11463 ( .IN1(n4382), .IN2(g3106), .Q(n11742) );
  OR2X1 U11464 ( .IN1(n11744), .IN2(n11745), .Q(g30709) );
  AND2X1 U11465 ( .IN1(n4524), .IN2(g2391), .Q(n11745) );
  AND2X1 U11466 ( .IN1(n11746), .IN2(g7264), .Q(n11744) );
  OR2X1 U11467 ( .IN1(n11747), .IN2(n11748), .Q(g30708) );
  AND2X1 U11468 ( .IN1(n4511), .IN2(g1698), .Q(n11748) );
  AND2X1 U11469 ( .IN1(n11749), .IN2(n4618), .Q(n11747) );
  OR2X1 U11470 ( .IN1(n11750), .IN2(n11751), .Q(g30707) );
  AND2X1 U11471 ( .IN1(n4516), .IN2(g2390), .Q(n11751) );
  AND2X1 U11472 ( .IN1(n11746), .IN2(g5555), .Q(n11750) );
  OR2X1 U11473 ( .IN1(n11752), .IN2(n11753), .Q(g30706) );
  AND2X1 U11474 ( .IN1(n4525), .IN2(g1697), .Q(n11753) );
  AND2X1 U11475 ( .IN1(n11749), .IN2(g7014), .Q(n11752) );
  OR2X1 U11476 ( .IN1(n11754), .IN2(n11755), .Q(g30705) );
  AND2X1 U11477 ( .IN1(n2594), .IN2(g1088), .Q(n11755) );
  AND2X1 U11478 ( .IN1(n4381), .IN2(g1004), .Q(n11754) );
  OR2X1 U11479 ( .IN1(n11756), .IN2(n11757), .Q(g30704) );
  AND2X1 U11480 ( .IN1(n4518), .IN2(g1696), .Q(n11757) );
  AND2X1 U11481 ( .IN1(n11749), .IN2(g5511), .Q(n11756) );
  AND2X1 U11482 ( .IN1(n11758), .IN2(n11759), .Q(n11749) );
  OR2X1 U11483 ( .IN1(n11760), .IN2(n11761), .Q(n11759) );
  AND2X1 U11484 ( .IN1(n11762), .IN2(n11763), .Q(n11761) );
  AND2X1 U11485 ( .IN1(n11764), .IN2(n11765), .Q(n11760) );
  INVX0 U11486 ( .INP(n11762), .ZN(n11765) );
  OR2X1 U11487 ( .IN1(n11766), .IN2(n11767), .Q(n11762) );
  OR2X1 U11488 ( .IN1(n11768), .IN2(n11769), .Q(n11767) );
  AND2X1 U11489 ( .IN1(n11770), .IN2(n11763), .Q(n11769) );
  AND2X1 U11490 ( .IN1(n11771), .IN2(n11772), .Q(n11770) );
  AND2X1 U11491 ( .IN1(n11773), .IN2(n11774), .Q(n11771) );
  OR2X1 U11492 ( .IN1(n11775), .IN2(n11776), .Q(n11774) );
  OR2X1 U11493 ( .IN1(n11777), .IN2(n11778), .Q(n11773) );
  AND2X1 U11494 ( .IN1(n11779), .IN2(n11780), .Q(n11777) );
  AND2X1 U11495 ( .IN1(n11781), .IN2(n11782), .Q(n11780) );
  AND2X1 U11496 ( .IN1(n11783), .IN2(n11784), .Q(n11779) );
  OR2X1 U11497 ( .IN1(n11785), .IN2(n11786), .Q(n11784) );
  AND2X1 U11498 ( .IN1(n11787), .IN2(n11764), .Q(n11768) );
  OR2X1 U11499 ( .IN1(n11788), .IN2(n11785), .Q(n11787) );
  AND2X1 U11500 ( .IN1(n11789), .IN2(n11790), .Q(n11788) );
  INVX0 U11501 ( .INP(n11791), .ZN(n11790) );
  AND2X1 U11502 ( .IN1(n11792), .IN2(n11793), .Q(n11789) );
  INVX0 U11503 ( .INP(n11794), .ZN(n11793) );
  OR2X1 U11504 ( .IN1(n11778), .IN2(n11795), .Q(n11792) );
  OR2X1 U11505 ( .IN1(n11796), .IN2(n11797), .Q(n11795) );
  AND2X1 U11506 ( .IN1(n11798), .IN2(n11799), .Q(n11766) );
  OR2X1 U11507 ( .IN1(n11800), .IN2(n11801), .Q(g30703) );
  AND2X1 U11508 ( .IN1(n2594), .IN2(g6712), .Q(n11801) );
  AND2X1 U11509 ( .IN1(n4364), .IN2(g1003), .Q(n11800) );
  OR2X1 U11510 ( .IN1(n11802), .IN2(n11803), .Q(g30702) );
  AND2X1 U11511 ( .IN1(n4506), .IN2(g317), .Q(n11803) );
  AND2X1 U11512 ( .IN1(n11804), .IN2(n4640), .Q(n11802) );
  OR2X1 U11513 ( .IN1(n11805), .IN2(n11806), .Q(g30701) );
  AND2X1 U11514 ( .IN1(n2594), .IN2(g5472), .Q(n11806) );
  AND2X1 U11515 ( .IN1(n4363), .IN2(g1002), .Q(n11805) );
  OR2X1 U11516 ( .IN1(n11807), .IN2(n11808), .Q(g30700) );
  AND2X1 U11517 ( .IN1(test_so18), .IN2(n4499), .Q(n11808) );
  AND2X1 U11518 ( .IN1(n11804), .IN2(g6447), .Q(n11807) );
  OR2X1 U11519 ( .IN1(n11809), .IN2(n11810), .Q(g30699) );
  AND2X1 U11520 ( .IN1(n4520), .IN2(g315), .Q(n11810) );
  AND2X1 U11521 ( .IN1(n11804), .IN2(g5437), .Q(n11809) );
  AND2X1 U11522 ( .IN1(n11811), .IN2(n11812), .Q(n11804) );
  OR2X1 U11523 ( .IN1(n11813), .IN2(n11814), .Q(n11812) );
  AND2X1 U11524 ( .IN1(n11815), .IN2(n11816), .Q(n11814) );
  AND2X1 U11525 ( .IN1(n11817), .IN2(n11818), .Q(n11813) );
  INVX0 U11526 ( .INP(n11815), .ZN(n11818) );
  OR2X1 U11527 ( .IN1(n11819), .IN2(n11820), .Q(n11815) );
  OR2X1 U11528 ( .IN1(n11821), .IN2(n11822), .Q(n11820) );
  AND2X1 U11529 ( .IN1(n11823), .IN2(n11816), .Q(n11822) );
  AND2X1 U11530 ( .IN1(n11824), .IN2(n11825), .Q(n11823) );
  AND2X1 U11531 ( .IN1(n11826), .IN2(n11827), .Q(n11824) );
  OR2X1 U11532 ( .IN1(n11828), .IN2(n11829), .Q(n11827) );
  OR2X1 U11533 ( .IN1(n11830), .IN2(n11831), .Q(n11826) );
  AND2X1 U11534 ( .IN1(n11832), .IN2(n11833), .Q(n11830) );
  AND2X1 U11535 ( .IN1(n11834), .IN2(n11835), .Q(n11833) );
  AND2X1 U11536 ( .IN1(n11836), .IN2(n11837), .Q(n11832) );
  OR2X1 U11537 ( .IN1(n11838), .IN2(n11839), .Q(n11837) );
  AND2X1 U11538 ( .IN1(n11840), .IN2(n11817), .Q(n11821) );
  OR2X1 U11539 ( .IN1(n11841), .IN2(n11838), .Q(n11840) );
  AND2X1 U11540 ( .IN1(n11842), .IN2(n11843), .Q(n11841) );
  INVX0 U11541 ( .INP(n11844), .ZN(n11843) );
  AND2X1 U11542 ( .IN1(n11845), .IN2(n11846), .Q(n11842) );
  INVX0 U11543 ( .INP(n11847), .ZN(n11846) );
  OR2X1 U11544 ( .IN1(n11831), .IN2(n11848), .Q(n11845) );
  OR2X1 U11545 ( .IN1(n11849), .IN2(n11850), .Q(n11848) );
  AND2X1 U11546 ( .IN1(n11851), .IN2(n11852), .Q(n11819) );
  OR2X1 U11547 ( .IN1(n11853), .IN2(n11854), .Q(g30695) );
  AND2X1 U11548 ( .IN1(n11855), .IN2(g2241), .Q(n11854) );
  AND2X1 U11549 ( .IN1(n4367), .IN2(g2276), .Q(n11853) );
  OR2X1 U11550 ( .IN1(n11856), .IN2(n11857), .Q(g30694) );
  AND2X1 U11551 ( .IN1(n11858), .IN2(g2241), .Q(n11857) );
  AND2X1 U11552 ( .IN1(n4367), .IN2(g2348), .Q(n11856) );
  OR2X1 U11553 ( .IN1(n11859), .IN2(n11860), .Q(g30693) );
  AND2X1 U11554 ( .IN1(test_so73), .IN2(n11855), .Q(n11860) );
  AND2X1 U11555 ( .IN1(g2273), .IN2(n10189), .Q(n11859) );
  OR2X1 U11556 ( .IN1(n11861), .IN2(n11862), .Q(g30692) );
  AND2X1 U11557 ( .IN1(n11863), .IN2(g1547), .Q(n11862) );
  AND2X1 U11558 ( .IN1(n4368), .IN2(g1582), .Q(n11861) );
  OR2X1 U11559 ( .IN1(n11864), .IN2(n11865), .Q(g30691) );
  AND2X1 U11560 ( .IN1(n11858), .IN2(test_so73), .Q(n11865) );
  AND2X1 U11561 ( .IN1(g2345), .IN2(n10189), .Q(n11864) );
  OR2X1 U11562 ( .IN1(n11866), .IN2(n11867), .Q(g30690) );
  AND2X1 U11563 ( .IN1(n11855), .IN2(g6837), .Q(n11867) );
  OR2X1 U11564 ( .IN1(n11868), .IN2(n11869), .Q(n11855) );
  OR2X1 U11565 ( .IN1(n11870), .IN2(n11871), .Q(n11869) );
  AND2X1 U11566 ( .IN1(n11872), .IN2(g2175), .Q(n11871) );
  AND2X1 U11567 ( .IN1(n11873), .IN2(n11874), .Q(n11870) );
  AND2X1 U11568 ( .IN1(n11875), .IN2(n11876), .Q(n11873) );
  OR2X1 U11569 ( .IN1(n11877), .IN2(n10863), .Q(n11876) );
  INVX0 U11570 ( .INP(n11878), .ZN(n11877) );
  OR2X1 U11571 ( .IN1(n10862), .IN2(n11878), .Q(n11875) );
  AND2X1 U11572 ( .IN1(n4324), .IN2(g2270), .Q(n11866) );
  OR2X1 U11573 ( .IN1(n11879), .IN2(n11880), .Q(g30689) );
  AND2X1 U11574 ( .IN1(n11881), .IN2(g1547), .Q(n11880) );
  AND2X1 U11575 ( .IN1(n4368), .IN2(g1654), .Q(n11879) );
  OR2X1 U11576 ( .IN1(n11882), .IN2(n11883), .Q(g30688) );
  AND2X1 U11577 ( .IN1(n11863), .IN2(g6782), .Q(n11883) );
  AND2X1 U11578 ( .IN1(n4515), .IN2(g1579), .Q(n11882) );
  OR2X1 U11579 ( .IN1(n11884), .IN2(n11885), .Q(g30687) );
  AND2X1 U11580 ( .IN1(test_so31), .IN2(n11886), .Q(n11885) );
  AND2X1 U11581 ( .IN1(g888), .IN2(n10188), .Q(n11884) );
  OR2X1 U11582 ( .IN1(n11887), .IN2(n11888), .Q(g30686) );
  AND2X1 U11583 ( .IN1(n11858), .IN2(g6837), .Q(n11888) );
  INVX0 U11584 ( .INP(n11889), .ZN(n11858) );
  OR2X1 U11585 ( .IN1(n11890), .IN2(n11891), .Q(n11889) );
  OR2X1 U11586 ( .IN1(n11892), .IN2(n11893), .Q(n11891) );
  AND2X1 U11587 ( .IN1(n11894), .IN2(n11874), .Q(n11893) );
  AND2X1 U11588 ( .IN1(n11895), .IN2(n11896), .Q(n11894) );
  OR2X1 U11589 ( .IN1(n10820), .IN2(n11897), .Q(n11896) );
  INVX0 U11590 ( .INP(n2669), .ZN(n11897) );
  OR2X1 U11591 ( .IN1(n2669), .IN2(n10821), .Q(n11895) );
  AND2X1 U11592 ( .IN1(n11872), .IN2(n11898), .Q(n11890) );
  AND2X1 U11593 ( .IN1(n4324), .IN2(g2342), .Q(n11887) );
  OR2X1 U11594 ( .IN1(n11899), .IN2(n11900), .Q(g30684) );
  AND2X1 U11595 ( .IN1(n11881), .IN2(g6782), .Q(n11900) );
  AND2X1 U11596 ( .IN1(n4515), .IN2(g1651), .Q(n11899) );
  OR2X1 U11597 ( .IN1(n11901), .IN2(n11902), .Q(g30683) );
  AND2X1 U11598 ( .IN1(n11863), .IN2(g6573), .Q(n11902) );
  OR2X1 U11599 ( .IN1(n11903), .IN2(n11904), .Q(n11863) );
  OR2X1 U11600 ( .IN1(n11905), .IN2(n11906), .Q(n11904) );
  AND2X1 U11601 ( .IN1(n11907), .IN2(g1481), .Q(n11906) );
  AND2X1 U11602 ( .IN1(n11908), .IN2(n11909), .Q(n11905) );
  AND2X1 U11603 ( .IN1(n11910), .IN2(n11911), .Q(n11908) );
  OR2X1 U11604 ( .IN1(n11912), .IN2(n10790), .Q(n11911) );
  INVX0 U11605 ( .INP(n11913), .ZN(n11912) );
  OR2X1 U11606 ( .IN1(n10789), .IN2(n11913), .Q(n11910) );
  AND2X1 U11607 ( .IN1(n4317), .IN2(g1576), .Q(n11901) );
  OR2X1 U11608 ( .IN1(n11914), .IN2(n11915), .Q(g30682) );
  AND2X1 U11609 ( .IN1(n11916), .IN2(test_so31), .Q(n11915) );
  AND2X1 U11610 ( .IN1(g960), .IN2(n10188), .Q(n11914) );
  OR2X1 U11611 ( .IN1(n11917), .IN2(n11918), .Q(g30681) );
  AND2X1 U11612 ( .IN1(n11886), .IN2(g6518), .Q(n11918) );
  AND2X1 U11613 ( .IN1(n4312), .IN2(g885), .Q(n11917) );
  OR2X1 U11614 ( .IN1(n11919), .IN2(n11920), .Q(g30680) );
  AND2X1 U11615 ( .IN1(n11921), .IN2(g165), .Q(n11920) );
  AND2X1 U11616 ( .IN1(n4369), .IN2(g201), .Q(n11919) );
  OR2X1 U11617 ( .IN1(n11922), .IN2(n11923), .Q(g30679) );
  AND2X1 U11618 ( .IN1(n11924), .IN2(g2241), .Q(n11923) );
  AND2X1 U11619 ( .IN1(n4367), .IN2(g2321), .Q(n11922) );
  OR2X1 U11620 ( .IN1(n11925), .IN2(n11926), .Q(g30678) );
  AND2X1 U11621 ( .IN1(n11881), .IN2(g6573), .Q(n11926) );
  INVX0 U11622 ( .INP(n11927), .ZN(n11881) );
  OR2X1 U11623 ( .IN1(n11928), .IN2(n11929), .Q(n11927) );
  OR2X1 U11624 ( .IN1(n11930), .IN2(n11931), .Q(n11929) );
  AND2X1 U11625 ( .IN1(n11932), .IN2(n11909), .Q(n11931) );
  AND2X1 U11626 ( .IN1(n11933), .IN2(n11934), .Q(n11932) );
  OR2X1 U11627 ( .IN1(n10775), .IN2(n11935), .Q(n11934) );
  INVX0 U11628 ( .INP(n2684), .ZN(n11935) );
  OR2X1 U11629 ( .IN1(n2684), .IN2(n10776), .Q(n11933) );
  AND2X1 U11630 ( .IN1(n11907), .IN2(n11936), .Q(n11928) );
  AND2X1 U11631 ( .IN1(n4317), .IN2(g1648), .Q(n11925) );
  OR2X1 U11632 ( .IN1(n11937), .IN2(n11938), .Q(g30677) );
  AND2X1 U11633 ( .IN1(n11916), .IN2(g6518), .Q(n11938) );
  AND2X1 U11634 ( .IN1(n4312), .IN2(g957), .Q(n11937) );
  OR2X1 U11635 ( .IN1(n11939), .IN2(n11940), .Q(g30676) );
  AND2X1 U11636 ( .IN1(n11886), .IN2(g6368), .Q(n11940) );
  OR2X1 U11637 ( .IN1(n11941), .IN2(n11942), .Q(n11886) );
  OR2X1 U11638 ( .IN1(n11943), .IN2(n11944), .Q(n11942) );
  AND2X1 U11639 ( .IN1(n11945), .IN2(n11946), .Q(n11944) );
  AND2X1 U11640 ( .IN1(n11947), .IN2(n11948), .Q(n11945) );
  OR2X1 U11641 ( .IN1(n11949), .IN2(n10734), .Q(n11948) );
  INVX0 U11642 ( .INP(n11950), .ZN(n11949) );
  OR2X1 U11643 ( .IN1(n10733), .IN2(n11950), .Q(n11947) );
  AND2X1 U11644 ( .IN1(n11951), .IN2(g793), .Q(n11941) );
  AND2X1 U11645 ( .IN1(n4323), .IN2(g882), .Q(n11939) );
  OR2X1 U11646 ( .IN1(n11952), .IN2(n11953), .Q(g30675) );
  AND2X1 U11647 ( .IN1(n11954), .IN2(g165), .Q(n11953) );
  AND2X1 U11648 ( .IN1(n4369), .IN2(g273), .Q(n11952) );
  OR2X1 U11649 ( .IN1(n11955), .IN2(n11956), .Q(g30674) );
  AND2X1 U11650 ( .IN1(n11921), .IN2(g6313), .Q(n11956) );
  AND2X1 U11651 ( .IN1(n4512), .IN2(g198), .Q(n11955) );
  OR2X1 U11652 ( .IN1(n11957), .IN2(n11958), .Q(g30673) );
  AND2X1 U11653 ( .IN1(n11924), .IN2(test_so73), .Q(n11958) );
  AND2X1 U11654 ( .IN1(g2318), .IN2(n10189), .Q(n11957) );
  OR2X1 U11655 ( .IN1(n11959), .IN2(n11960), .Q(g30672) );
  AND2X1 U11656 ( .IN1(n11961), .IN2(g2241), .Q(n11960) );
  AND2X1 U11657 ( .IN1(n4367), .IN2(g2312), .Q(n11959) );
  OR2X1 U11658 ( .IN1(n11962), .IN2(n11963), .Q(g30671) );
  AND2X1 U11659 ( .IN1(n11964), .IN2(g1547), .Q(n11963) );
  AND2X1 U11660 ( .IN1(n4368), .IN2(g1627), .Q(n11962) );
  OR2X1 U11661 ( .IN1(n11965), .IN2(n11966), .Q(g30670) );
  AND2X1 U11662 ( .IN1(n11916), .IN2(g6368), .Q(n11966) );
  INVX0 U11663 ( .INP(n11967), .ZN(n11916) );
  OR2X1 U11664 ( .IN1(n11968), .IN2(n11969), .Q(n11967) );
  OR2X1 U11665 ( .IN1(n11970), .IN2(n11971), .Q(n11969) );
  AND2X1 U11666 ( .IN1(n11946), .IN2(n11972), .Q(n11971) );
  OR2X1 U11667 ( .IN1(n11973), .IN2(n11974), .Q(n11972) );
  AND2X1 U11668 ( .IN1(n11975), .IN2(n10712), .Q(n11974) );
  INVX0 U11669 ( .INP(n11976), .ZN(n11975) );
  AND2X1 U11670 ( .IN1(n10711), .IN2(n11976), .Q(n11973) );
  OR2X1 U11671 ( .IN1(n11977), .IN2(n11978), .Q(n11976) );
  AND2X1 U11672 ( .IN1(n11979), .IN2(n11980), .Q(n11977) );
  OR2X1 U11673 ( .IN1(n11981), .IN2(n10730), .Q(n11980) );
  OR2X1 U11674 ( .IN1(n10729), .IN2(n11982), .Q(n11979) );
  AND2X1 U11675 ( .IN1(n11951), .IN2(n11983), .Q(n11968) );
  AND2X1 U11676 ( .IN1(n4323), .IN2(g954), .Q(n11965) );
  OR2X1 U11677 ( .IN1(n11984), .IN2(n11985), .Q(g30669) );
  AND2X1 U11678 ( .IN1(n11954), .IN2(g6313), .Q(n11985) );
  AND2X1 U11679 ( .IN1(n4512), .IN2(g270), .Q(n11984) );
  OR2X1 U11680 ( .IN1(n11986), .IN2(n11987), .Q(g30668) );
  AND2X1 U11681 ( .IN1(n11921), .IN2(g6231), .Q(n11987) );
  OR2X1 U11682 ( .IN1(n11988), .IN2(n11989), .Q(n11921) );
  OR2X1 U11683 ( .IN1(n11990), .IN2(n11991), .Q(n11989) );
  AND2X1 U11684 ( .IN1(n11992), .IN2(n11993), .Q(n11991) );
  AND2X1 U11685 ( .IN1(n11994), .IN2(n11995), .Q(n11992) );
  OR2X1 U11686 ( .IN1(n11996), .IN2(n10664), .Q(n11995) );
  INVX0 U11687 ( .INP(n11997), .ZN(n11996) );
  OR2X1 U11688 ( .IN1(n10663), .IN2(n11997), .Q(n11994) );
  AND2X1 U11689 ( .IN1(n11998), .IN2(g105), .Q(n11988) );
  AND2X1 U11690 ( .IN1(n4318), .IN2(g195), .Q(n11986) );
  OR2X1 U11691 ( .IN1(n11999), .IN2(n12000), .Q(g30667) );
  AND2X1 U11692 ( .IN1(n11924), .IN2(g6837), .Q(n12000) );
  INVX0 U11693 ( .INP(n12001), .ZN(n11924) );
  OR2X1 U11694 ( .IN1(n12002), .IN2(n12003), .Q(n12001) );
  OR2X1 U11695 ( .IN1(n11892), .IN2(n12004), .Q(n12003) );
  AND2X1 U11696 ( .IN1(n11874), .IN2(n12005), .Q(n12004) );
  OR2X1 U11697 ( .IN1(n12006), .IN2(n12007), .Q(n12005) );
  AND2X1 U11698 ( .IN1(n12008), .IN2(n10841), .Q(n12007) );
  INVX0 U11699 ( .INP(n12009), .ZN(n12008) );
  AND2X1 U11700 ( .IN1(n10840), .IN2(n12009), .Q(n12006) );
  OR2X1 U11701 ( .IN1(n12010), .IN2(n12011), .Q(n12009) );
  AND2X1 U11702 ( .IN1(n4529), .IN2(n10862), .Q(n12010) );
  AND2X1 U11703 ( .IN1(n11872), .IN2(n4389), .Q(n12002) );
  AND2X1 U11704 ( .IN1(n4324), .IN2(g2315), .Q(n11999) );
  OR2X1 U11705 ( .IN1(n12012), .IN2(n12013), .Q(g30666) );
  AND2X1 U11706 ( .IN1(n11961), .IN2(test_so73), .Q(n12013) );
  AND2X1 U11707 ( .IN1(g2309), .IN2(n10189), .Q(n12012) );
  OR2X1 U11708 ( .IN1(n12014), .IN2(n12015), .Q(g30665) );
  AND2X1 U11709 ( .IN1(n12016), .IN2(g2241), .Q(n12015) );
  AND2X1 U11710 ( .IN1(n4367), .IN2(g2303), .Q(n12014) );
  OR2X1 U11711 ( .IN1(n12017), .IN2(n12018), .Q(g30664) );
  AND2X1 U11712 ( .IN1(n11964), .IN2(g6782), .Q(n12018) );
  AND2X1 U11713 ( .IN1(n4515), .IN2(g1624), .Q(n12017) );
  OR2X1 U11714 ( .IN1(n12019), .IN2(n12020), .Q(g30663) );
  AND2X1 U11715 ( .IN1(n12021), .IN2(g1547), .Q(n12020) );
  AND2X1 U11716 ( .IN1(n4368), .IN2(g1618), .Q(n12019) );
  OR2X1 U11717 ( .IN1(n12022), .IN2(n12023), .Q(g30662) );
  AND2X1 U11718 ( .IN1(n12024), .IN2(test_so31), .Q(n12023) );
  AND2X1 U11719 ( .IN1(g933), .IN2(n10188), .Q(n12022) );
  OR2X1 U11720 ( .IN1(n12025), .IN2(n12026), .Q(g30661) );
  AND2X1 U11721 ( .IN1(n11954), .IN2(g6231), .Q(n12026) );
  INVX0 U11722 ( .INP(n12027), .ZN(n11954) );
  OR2X1 U11723 ( .IN1(n12028), .IN2(n12029), .Q(n12027) );
  OR2X1 U11724 ( .IN1(n12030), .IN2(n12031), .Q(n12029) );
  AND2X1 U11725 ( .IN1(n12032), .IN2(n11993), .Q(n12031) );
  AND2X1 U11726 ( .IN1(n12033), .IN2(n12034), .Q(n12032) );
  OR2X1 U11727 ( .IN1(n10646), .IN2(n12035), .Q(n12034) );
  INVX0 U11728 ( .INP(n2717), .ZN(n12035) );
  OR2X1 U11729 ( .IN1(n2717), .IN2(n10647), .Q(n12033) );
  AND2X1 U11730 ( .IN1(n11998), .IN2(n12036), .Q(n12028) );
  AND2X1 U11731 ( .IN1(n4318), .IN2(g267), .Q(n12025) );
  OR2X1 U11732 ( .IN1(n12037), .IN2(n12038), .Q(g30660) );
  AND2X1 U11733 ( .IN1(n11961), .IN2(g6837), .Q(n12038) );
  INVX0 U11734 ( .INP(n12039), .ZN(n11961) );
  OR2X1 U11735 ( .IN1(n12040), .IN2(n12041), .Q(n12039) );
  OR2X1 U11736 ( .IN1(n11892), .IN2(n12042), .Q(n12041) );
  AND2X1 U11737 ( .IN1(n11874), .IN2(n12043), .Q(n12042) );
  OR2X1 U11738 ( .IN1(n12044), .IN2(n12045), .Q(n12043) );
  AND2X1 U11739 ( .IN1(n12046), .IN2(n10870), .Q(n12045) );
  INVX0 U11740 ( .INP(n12047), .ZN(n12046) );
  AND2X1 U11741 ( .IN1(n12048), .IN2(n12047), .Q(n12044) );
  AND2X1 U11742 ( .IN1(n4529), .IN2(n12049), .Q(n11892) );
  AND2X1 U11743 ( .IN1(n11872), .IN2(n4373), .Q(n12040) );
  AND2X1 U11744 ( .IN1(n4324), .IN2(g2306), .Q(n12037) );
  OR2X1 U11745 ( .IN1(n12050), .IN2(n12051), .Q(g30659) );
  AND2X1 U11746 ( .IN1(test_so73), .IN2(n12016), .Q(n12051) );
  AND2X1 U11747 ( .IN1(g2300), .IN2(n10189), .Q(n12050) );
  OR2X1 U11748 ( .IN1(n12052), .IN2(n12053), .Q(g30658) );
  AND2X1 U11749 ( .IN1(test_so55), .IN2(n4317), .Q(n12053) );
  AND2X1 U11750 ( .IN1(n11964), .IN2(g6573), .Q(n12052) );
  INVX0 U11751 ( .INP(n12054), .ZN(n11964) );
  OR2X1 U11752 ( .IN1(n12055), .IN2(n12056), .Q(n12054) );
  OR2X1 U11753 ( .IN1(n11930), .IN2(n12057), .Q(n12056) );
  AND2X1 U11754 ( .IN1(n11909), .IN2(n12058), .Q(n12057) );
  OR2X1 U11755 ( .IN1(n12059), .IN2(n12060), .Q(n12058) );
  AND2X1 U11756 ( .IN1(n12061), .IN2(n10780), .Q(n12060) );
  INVX0 U11757 ( .INP(n12062), .ZN(n12061) );
  AND2X1 U11758 ( .IN1(n10779), .IN2(n12062), .Q(n12059) );
  OR2X1 U11759 ( .IN1(n12063), .IN2(n12064), .Q(n12062) );
  AND2X1 U11760 ( .IN1(n4530), .IN2(n10789), .Q(n12063) );
  AND2X1 U11761 ( .IN1(n11907), .IN2(n4390), .Q(n12055) );
  OR2X1 U11762 ( .IN1(n12065), .IN2(n12066), .Q(g30657) );
  AND2X1 U11763 ( .IN1(n12021), .IN2(g6782), .Q(n12066) );
  AND2X1 U11764 ( .IN1(n4515), .IN2(g1615), .Q(n12065) );
  OR2X1 U11765 ( .IN1(n12067), .IN2(n12068), .Q(g30656) );
  AND2X1 U11766 ( .IN1(n12069), .IN2(g1547), .Q(n12068) );
  AND2X1 U11767 ( .IN1(n4368), .IN2(g1609), .Q(n12067) );
  OR2X1 U11768 ( .IN1(n12070), .IN2(n12071), .Q(g30655) );
  AND2X1 U11769 ( .IN1(n12024), .IN2(g6518), .Q(n12071) );
  AND2X1 U11770 ( .IN1(n4312), .IN2(g930), .Q(n12070) );
  OR2X1 U11771 ( .IN1(n12072), .IN2(n12073), .Q(g30654) );
  AND2X1 U11772 ( .IN1(n12074), .IN2(test_so31), .Q(n12073) );
  AND2X1 U11773 ( .IN1(test_so34), .IN2(n10188), .Q(n12072) );
  OR2X1 U11774 ( .IN1(n12075), .IN2(n12076), .Q(g30653) );
  AND2X1 U11775 ( .IN1(n12077), .IN2(g165), .Q(n12076) );
  AND2X1 U11776 ( .IN1(n4369), .IN2(g246), .Q(n12075) );
  OR2X1 U11777 ( .IN1(n12078), .IN2(n12079), .Q(g30652) );
  AND2X1 U11778 ( .IN1(n12016), .IN2(g6837), .Q(n12079) );
  OR2X1 U11779 ( .IN1(n11868), .IN2(n12080), .Q(n12016) );
  OR2X1 U11780 ( .IN1(n12081), .IN2(n12082), .Q(n12080) );
  AND2X1 U11781 ( .IN1(n11872), .IN2(n12083), .Q(n12082) );
  AND2X1 U11782 ( .IN1(n12084), .IN2(n11874), .Q(n12081) );
  AND2X1 U11783 ( .IN1(n12085), .IN2(n12086), .Q(n12084) );
  OR2X1 U11784 ( .IN1(n12087), .IN2(n10837), .Q(n12086) );
  INVX0 U11785 ( .INP(n2670), .ZN(n12087) );
  OR2X1 U11786 ( .IN1(n2670), .IN2(n10836), .Q(n12085) );
  OR2X1 U11787 ( .IN1(n12088), .IN2(n12089), .Q(n2670) );
  AND2X1 U11788 ( .IN1(n12090), .IN2(n12091), .Q(n12088) );
  OR2X1 U11789 ( .IN1(n4529), .IN2(n10829), .Q(n12091) );
  OR2X1 U11790 ( .IN1(n10828), .IN2(n11593), .Q(n12090) );
  AND2X1 U11791 ( .IN1(n12049), .IN2(n12092), .Q(n11868) );
  AND2X1 U11792 ( .IN1(n4324), .IN2(g2297), .Q(n12078) );
  OR2X1 U11793 ( .IN1(n12093), .IN2(n12094), .Q(g30651) );
  AND2X1 U11794 ( .IN1(n12021), .IN2(g6573), .Q(n12094) );
  INVX0 U11795 ( .INP(n12095), .ZN(n12021) );
  OR2X1 U11796 ( .IN1(n12096), .IN2(n12097), .Q(n12095) );
  OR2X1 U11797 ( .IN1(n11930), .IN2(n12098), .Q(n12097) );
  AND2X1 U11798 ( .IN1(n11909), .IN2(n12099), .Q(n12098) );
  OR2X1 U11799 ( .IN1(n12100), .IN2(n12101), .Q(n12099) );
  AND2X1 U11800 ( .IN1(n12102), .IN2(n10756), .Q(n12101) );
  INVX0 U11801 ( .INP(n12103), .ZN(n12102) );
  AND2X1 U11802 ( .IN1(n10755), .IN2(n12103), .Q(n12100) );
  AND2X1 U11803 ( .IN1(n4530), .IN2(n12104), .Q(n11930) );
  AND2X1 U11804 ( .IN1(n11907), .IN2(n4374), .Q(n12096) );
  AND2X1 U11805 ( .IN1(n4317), .IN2(g1612), .Q(n12093) );
  OR2X1 U11806 ( .IN1(n12105), .IN2(n12106), .Q(g30650) );
  AND2X1 U11807 ( .IN1(n12069), .IN2(g6782), .Q(n12106) );
  AND2X1 U11808 ( .IN1(test_so56), .IN2(n4515), .Q(n12105) );
  OR2X1 U11809 ( .IN1(n12107), .IN2(n12108), .Q(g30649) );
  AND2X1 U11810 ( .IN1(n12024), .IN2(g6368), .Q(n12108) );
  INVX0 U11811 ( .INP(n12109), .ZN(n12024) );
  OR2X1 U11812 ( .IN1(n12110), .IN2(n12111), .Q(n12109) );
  OR2X1 U11813 ( .IN1(n11970), .IN2(n12112), .Q(n12111) );
  AND2X1 U11814 ( .IN1(n11946), .IN2(n12113), .Q(n12112) );
  OR2X1 U11815 ( .IN1(n12114), .IN2(n12115), .Q(n12113) );
  AND2X1 U11816 ( .IN1(n12116), .IN2(n10692), .Q(n12115) );
  INVX0 U11817 ( .INP(n12117), .ZN(n12116) );
  AND2X1 U11818 ( .IN1(n10691), .IN2(n12117), .Q(n12114) );
  OR2X1 U11819 ( .IN1(n12118), .IN2(n12119), .Q(n12117) );
  AND2X1 U11820 ( .IN1(n11981), .IN2(n10733), .Q(n12118) );
  AND2X1 U11821 ( .IN1(n11951), .IN2(n4391), .Q(n12110) );
  AND2X1 U11822 ( .IN1(n4323), .IN2(g927), .Q(n12107) );
  OR2X1 U11823 ( .IN1(n12120), .IN2(n12121), .Q(g30648) );
  AND2X1 U11824 ( .IN1(n12074), .IN2(g6518), .Q(n12121) );
  AND2X1 U11825 ( .IN1(n4312), .IN2(g921), .Q(n12120) );
  OR2X1 U11826 ( .IN1(n12122), .IN2(n12123), .Q(g30647) );
  AND2X1 U11827 ( .IN1(test_so31), .IN2(n12124), .Q(n12123) );
  AND2X1 U11828 ( .IN1(g915), .IN2(n10188), .Q(n12122) );
  OR2X1 U11829 ( .IN1(n12125), .IN2(n12126), .Q(g30646) );
  AND2X1 U11830 ( .IN1(n12077), .IN2(g6313), .Q(n12126) );
  AND2X1 U11831 ( .IN1(n4512), .IN2(g243), .Q(n12125) );
  OR2X1 U11832 ( .IN1(n12127), .IN2(n12128), .Q(g30645) );
  AND2X1 U11833 ( .IN1(n12129), .IN2(g165), .Q(n12128) );
  AND2X1 U11834 ( .IN1(n4369), .IN2(g237), .Q(n12127) );
  OR2X1 U11835 ( .IN1(n12130), .IN2(n12131), .Q(g30644) );
  AND2X1 U11836 ( .IN1(n12069), .IN2(g6573), .Q(n12131) );
  OR2X1 U11837 ( .IN1(n11903), .IN2(n12132), .Q(n12069) );
  OR2X1 U11838 ( .IN1(n12133), .IN2(n12134), .Q(n12132) );
  AND2X1 U11839 ( .IN1(n11907), .IN2(n12135), .Q(n12134) );
  AND2X1 U11840 ( .IN1(n12136), .IN2(n11909), .Q(n12133) );
  AND2X1 U11841 ( .IN1(n12137), .IN2(n12138), .Q(n12136) );
  OR2X1 U11842 ( .IN1(n12139), .IN2(n10794), .Q(n12138) );
  INVX0 U11843 ( .INP(n2685), .ZN(n12139) );
  OR2X1 U11844 ( .IN1(n2685), .IN2(n10793), .Q(n12137) );
  OR2X1 U11845 ( .IN1(n12140), .IN2(n12141), .Q(n2685) );
  AND2X1 U11846 ( .IN1(n12142), .IN2(n12143), .Q(n12140) );
  OR2X1 U11847 ( .IN1(n4530), .IN2(n10764), .Q(n12143) );
  OR2X1 U11848 ( .IN1(n10763), .IN2(n11590), .Q(n12142) );
  AND2X1 U11849 ( .IN1(n12104), .IN2(n12144), .Q(n11903) );
  AND2X1 U11850 ( .IN1(n4317), .IN2(g1603), .Q(n12130) );
  OR2X1 U11851 ( .IN1(n12145), .IN2(n12146), .Q(g30643) );
  AND2X1 U11852 ( .IN1(n12074), .IN2(g6368), .Q(n12146) );
  INVX0 U11853 ( .INP(n12147), .ZN(n12074) );
  OR2X1 U11854 ( .IN1(n12148), .IN2(n12149), .Q(n12147) );
  OR2X1 U11855 ( .IN1(n11970), .IN2(n12150), .Q(n12149) );
  AND2X1 U11856 ( .IN1(n11946), .IN2(n12151), .Q(n12150) );
  OR2X1 U11857 ( .IN1(n12152), .IN2(n12153), .Q(n12151) );
  AND2X1 U11858 ( .IN1(n12154), .IN2(n10700), .Q(n12153) );
  INVX0 U11859 ( .INP(n12155), .ZN(n12154) );
  AND2X1 U11860 ( .IN1(n10699), .IN2(n12155), .Q(n12152) );
  AND2X1 U11861 ( .IN1(n11981), .IN2(n12156), .Q(n11970) );
  AND2X1 U11862 ( .IN1(n11951), .IN2(n4375), .Q(n12148) );
  AND2X1 U11863 ( .IN1(n4323), .IN2(g918), .Q(n12145) );
  OR2X1 U11864 ( .IN1(n12157), .IN2(n12158), .Q(g30642) );
  AND2X1 U11865 ( .IN1(n12124), .IN2(g6518), .Q(n12158) );
  AND2X1 U11866 ( .IN1(n4312), .IN2(g912), .Q(n12157) );
  OR2X1 U11867 ( .IN1(n12159), .IN2(n12160), .Q(g30641) );
  AND2X1 U11868 ( .IN1(n12077), .IN2(g6231), .Q(n12160) );
  INVX0 U11869 ( .INP(n12161), .ZN(n12077) );
  OR2X1 U11870 ( .IN1(n12162), .IN2(n12163), .Q(n12161) );
  OR2X1 U11871 ( .IN1(n12030), .IN2(n12164), .Q(n12163) );
  AND2X1 U11872 ( .IN1(n11993), .IN2(n12165), .Q(n12164) );
  OR2X1 U11873 ( .IN1(n12166), .IN2(n12167), .Q(n12165) );
  AND2X1 U11874 ( .IN1(n12168), .IN2(n10676), .Q(n12167) );
  INVX0 U11875 ( .INP(n12169), .ZN(n12168) );
  AND2X1 U11876 ( .IN1(n10675), .IN2(n12169), .Q(n12166) );
  OR2X1 U11877 ( .IN1(n12170), .IN2(n12171), .Q(n12169) );
  AND2X1 U11878 ( .IN1(n11586), .IN2(n10663), .Q(n12170) );
  AND2X1 U11879 ( .IN1(n11998), .IN2(n4392), .Q(n12162) );
  AND2X1 U11880 ( .IN1(n4318), .IN2(g240), .Q(n12159) );
  OR2X1 U11881 ( .IN1(n12172), .IN2(n12173), .Q(g30640) );
  AND2X1 U11882 ( .IN1(n12129), .IN2(g6313), .Q(n12173) );
  AND2X1 U11883 ( .IN1(n4512), .IN2(g234), .Q(n12172) );
  OR2X1 U11884 ( .IN1(n12174), .IN2(n12175), .Q(g30639) );
  AND2X1 U11885 ( .IN1(n12176), .IN2(g165), .Q(n12175) );
  AND2X1 U11886 ( .IN1(n4369), .IN2(g228), .Q(n12174) );
  OR2X1 U11887 ( .IN1(n12177), .IN2(n12178), .Q(g30638) );
  AND2X1 U11888 ( .IN1(n12124), .IN2(g6368), .Q(n12178) );
  OR2X1 U11889 ( .IN1(n12179), .IN2(n12180), .Q(n12124) );
  OR2X1 U11890 ( .IN1(n11943), .IN2(n12181), .Q(n12180) );
  AND2X1 U11891 ( .IN1(n12182), .IN2(n11946), .Q(n12181) );
  AND2X1 U11892 ( .IN1(n12183), .IN2(n12184), .Q(n12182) );
  OR2X1 U11893 ( .IN1(n12185), .IN2(n10730), .Q(n12184) );
  INVX0 U11894 ( .INP(n11978), .ZN(n12185) );
  OR2X1 U11895 ( .IN1(n10729), .IN2(n11978), .Q(n12183) );
  OR2X1 U11896 ( .IN1(n12186), .IN2(n12187), .Q(n11978) );
  OR2X1 U11897 ( .IN1(n12188), .IN2(n12189), .Q(n12187) );
  AND2X1 U11898 ( .IN1(n11981), .IN2(n10740), .Q(n12189) );
  AND2X1 U11899 ( .IN1(n10707), .IN2(n10741), .Q(n12188) );
  AND2X1 U11900 ( .IN1(n11982), .IN2(n12156), .Q(n11943) );
  AND2X1 U11901 ( .IN1(n11951), .IN2(n12190), .Q(n12179) );
  AND2X1 U11902 ( .IN1(n4323), .IN2(g909), .Q(n12177) );
  OR2X1 U11903 ( .IN1(n12191), .IN2(n12192), .Q(g30637) );
  AND2X1 U11904 ( .IN1(n12129), .IN2(g6231), .Q(n12192) );
  INVX0 U11905 ( .INP(n12193), .ZN(n12129) );
  OR2X1 U11906 ( .IN1(n12194), .IN2(n12195), .Q(n12193) );
  OR2X1 U11907 ( .IN1(n12030), .IN2(n12196), .Q(n12195) );
  AND2X1 U11908 ( .IN1(n11993), .IN2(n12197), .Q(n12196) );
  OR2X1 U11909 ( .IN1(n12198), .IN2(n12199), .Q(n12197) );
  AND2X1 U11910 ( .IN1(n12200), .IN2(n10627), .Q(n12199) );
  INVX0 U11911 ( .INP(n12201), .ZN(n12200) );
  AND2X1 U11912 ( .IN1(n10626), .IN2(n12201), .Q(n12198) );
  AND2X1 U11913 ( .IN1(n11586), .IN2(n12202), .Q(n12030) );
  AND2X1 U11914 ( .IN1(n11998), .IN2(n4376), .Q(n12194) );
  AND2X1 U11915 ( .IN1(n4318), .IN2(g231), .Q(n12191) );
  OR2X1 U11916 ( .IN1(n12203), .IN2(n12204), .Q(g30636) );
  AND2X1 U11917 ( .IN1(n12176), .IN2(g6313), .Q(n12204) );
  AND2X1 U11918 ( .IN1(n4512), .IN2(g225), .Q(n12203) );
  OR2X1 U11919 ( .IN1(n12205), .IN2(n12206), .Q(g30635) );
  AND2X1 U11920 ( .IN1(n12176), .IN2(g6231), .Q(n12206) );
  OR2X1 U11921 ( .IN1(n12207), .IN2(n12208), .Q(n12176) );
  OR2X1 U11922 ( .IN1(n11990), .IN2(n12209), .Q(n12208) );
  AND2X1 U11923 ( .IN1(n12210), .IN2(n11993), .Q(n12209) );
  AND2X1 U11924 ( .IN1(n12211), .IN2(n12212), .Q(n12210) );
  OR2X1 U11925 ( .IN1(n12213), .IN2(n10651), .Q(n12212) );
  INVX0 U11926 ( .INP(n2718), .ZN(n12213) );
  OR2X1 U11927 ( .IN1(n2718), .IN2(n10650), .Q(n12211) );
  OR2X1 U11928 ( .IN1(n12214), .IN2(n12215), .Q(n2718) );
  AND2X1 U11929 ( .IN1(n12216), .IN2(n12217), .Q(n12214) );
  OR2X1 U11930 ( .IN1(n11586), .IN2(n10635), .Q(n12217) );
  OR2X1 U11931 ( .IN1(n10634), .IN2(n11587), .Q(n12216) );
  AND2X1 U11932 ( .IN1(n11587), .IN2(n12202), .Q(n11990) );
  AND2X1 U11933 ( .IN1(n11998), .IN2(n12218), .Q(n12207) );
  AND2X1 U11934 ( .IN1(n4318), .IN2(g222), .Q(n12205) );
  OR2X1 U11935 ( .IN1(n12219), .IN2(n12220), .Q(g30566) );
  AND2X1 U11936 ( .IN1(n4509), .IN2(g2392), .Q(n12220) );
  AND2X1 U11937 ( .IN1(n11746), .IN2(n4606), .Q(n12219) );
  AND2X1 U11938 ( .IN1(n12221), .IN2(n12222), .Q(n11746) );
  OR2X1 U11939 ( .IN1(n12223), .IN2(n12224), .Q(n12222) );
  AND2X1 U11940 ( .IN1(n12225), .IN2(n12226), .Q(n12224) );
  AND2X1 U11941 ( .IN1(n12227), .IN2(n12228), .Q(n12223) );
  INVX0 U11942 ( .INP(n12225), .ZN(n12228) );
  OR2X1 U11943 ( .IN1(n12229), .IN2(n12230), .Q(n12225) );
  OR2X1 U11944 ( .IN1(n12231), .IN2(n12232), .Q(n12230) );
  AND2X1 U11945 ( .IN1(n12233), .IN2(n12226), .Q(n12232) );
  AND2X1 U11946 ( .IN1(n12234), .IN2(n12235), .Q(n12233) );
  AND2X1 U11947 ( .IN1(n12236), .IN2(n12237), .Q(n12234) );
  OR2X1 U11948 ( .IN1(n12238), .IN2(n12239), .Q(n12237) );
  OR2X1 U11949 ( .IN1(n12240), .IN2(n12241), .Q(n12236) );
  AND2X1 U11950 ( .IN1(n12242), .IN2(n12243), .Q(n12240) );
  AND2X1 U11951 ( .IN1(n12244), .IN2(n12245), .Q(n12243) );
  AND2X1 U11952 ( .IN1(n12246), .IN2(n12247), .Q(n12242) );
  OR2X1 U11953 ( .IN1(n12248), .IN2(n12249), .Q(n12247) );
  AND2X1 U11954 ( .IN1(n12250), .IN2(n12227), .Q(n12231) );
  OR2X1 U11955 ( .IN1(n12251), .IN2(n12248), .Q(n12250) );
  AND2X1 U11956 ( .IN1(n12252), .IN2(n12253), .Q(n12251) );
  INVX0 U11957 ( .INP(n12254), .ZN(n12253) );
  AND2X1 U11958 ( .IN1(n12255), .IN2(n12256), .Q(n12252) );
  INVX0 U11959 ( .INP(n12257), .ZN(n12256) );
  OR2X1 U11960 ( .IN1(n12241), .IN2(n12258), .Q(n12255) );
  OR2X1 U11961 ( .IN1(n12259), .IN2(n12260), .Q(n12258) );
  AND2X1 U11962 ( .IN1(n12261), .IN2(n12262), .Q(n12229) );
  OR2X1 U11963 ( .IN1(n12263), .IN2(n12264), .Q(g30505) );
  AND2X1 U11964 ( .IN1(n4516), .IN2(g2393), .Q(n12264) );
  AND2X1 U11965 ( .IN1(n12265), .IN2(g5555), .Q(n12263) );
  OR2X1 U11966 ( .IN1(n12266), .IN2(n12267), .Q(g30503) );
  AND2X1 U11967 ( .IN1(n4525), .IN2(g1700), .Q(n12267) );
  AND2X1 U11968 ( .IN1(n12268), .IN2(g7014), .Q(n12266) );
  OR2X1 U11969 ( .IN1(n12269), .IN2(n12270), .Q(g30500) );
  AND2X1 U11970 ( .IN1(test_so39), .IN2(n4381), .Q(n12270) );
  AND2X1 U11971 ( .IN1(n2798), .IN2(g1088), .Q(n12269) );
  OR2X1 U11972 ( .IN1(n12271), .IN2(n12272), .Q(g30487) );
  AND2X1 U11973 ( .IN1(n4518), .IN2(g1699), .Q(n12272) );
  AND2X1 U11974 ( .IN1(n12268), .IN2(g5511), .Q(n12271) );
  OR2X1 U11975 ( .IN1(n12273), .IN2(n12274), .Q(g30485) );
  AND2X1 U11976 ( .IN1(n2798), .IN2(g6712), .Q(n12274) );
  AND2X1 U11977 ( .IN1(n4364), .IN2(g1006), .Q(n12273) );
  OR2X1 U11978 ( .IN1(n12275), .IN2(n12276), .Q(g30482) );
  AND2X1 U11979 ( .IN1(n4506), .IN2(g320), .Q(n12276) );
  AND2X1 U11980 ( .IN1(n12277), .IN2(n4640), .Q(n12275) );
  OR2X1 U11981 ( .IN1(n12278), .IN2(n12279), .Q(g30470) );
  AND2X1 U11982 ( .IN1(n2798), .IN2(g5472), .Q(n12279) );
  AND2X1 U11983 ( .IN1(n4363), .IN2(g1005), .Q(n12278) );
  OR2X1 U11984 ( .IN1(n12280), .IN2(n12281), .Q(g30468) );
  AND2X1 U11985 ( .IN1(n4499), .IN2(g319), .Q(n12281) );
  AND2X1 U11986 ( .IN1(n12277), .IN2(g6447), .Q(n12280) );
  OR2X1 U11987 ( .IN1(n12282), .IN2(n12283), .Q(g30455) );
  AND2X1 U11988 ( .IN1(n4520), .IN2(g318), .Q(n12283) );
  AND2X1 U11989 ( .IN1(n12277), .IN2(g5437), .Q(n12282) );
  AND2X1 U11990 ( .IN1(n11811), .IN2(n12284), .Q(n12277) );
  AND2X1 U11991 ( .IN1(n12285), .IN2(n12286), .Q(n12284) );
  INVX0 U11992 ( .INP(n12287), .ZN(n12286) );
  AND2X1 U11993 ( .IN1(n12288), .IN2(n12289), .Q(n12287) );
  OR2X1 U11994 ( .IN1(n11851), .IN2(n11831), .Q(n12288) );
  OR2X1 U11995 ( .IN1(n12289), .IN2(n11831), .Q(n12285) );
  OR2X1 U11996 ( .IN1(n12290), .IN2(n12291), .Q(n12289) );
  OR2X1 U11997 ( .IN1(n11851), .IN2(n12292), .Q(n12291) );
  AND2X1 U11998 ( .IN1(n12293), .IN2(n11831), .Q(n12292) );
  OR2X1 U11999 ( .IN1(n12294), .IN2(n12295), .Q(n12290) );
  AND2X1 U12000 ( .IN1(n12296), .IN2(n11817), .Q(n12295) );
  AND2X1 U12001 ( .IN1(n12297), .IN2(n11825), .Q(n12296) );
  OR2X1 U12002 ( .IN1(n12298), .IN2(n11838), .Q(n12297) );
  AND2X1 U12003 ( .IN1(n11828), .IN2(n11839), .Q(n12298) );
  AND2X1 U12004 ( .IN1(n11816), .IN2(n12299), .Q(n12294) );
  OR2X1 U12005 ( .IN1(n4388), .IN2(n12300), .Q(n12299) );
  OR2X1 U12006 ( .IN1(n12301), .IN2(n12302), .Q(g30356) );
  AND2X1 U12007 ( .IN1(n4509), .IN2(g2395), .Q(n12302) );
  AND2X1 U12008 ( .IN1(n12265), .IN2(n4606), .Q(n12301) );
  OR2X1 U12009 ( .IN1(n12303), .IN2(n12304), .Q(g30341) );
  AND2X1 U12010 ( .IN1(n4524), .IN2(g2394), .Q(n12304) );
  AND2X1 U12011 ( .IN1(n12265), .IN2(g7264), .Q(n12303) );
  AND2X1 U12012 ( .IN1(n12221), .IN2(n12305), .Q(n12265) );
  AND2X1 U12013 ( .IN1(n12306), .IN2(n12307), .Q(n12305) );
  INVX0 U12014 ( .INP(n12308), .ZN(n12307) );
  AND2X1 U12015 ( .IN1(n12309), .IN2(n12310), .Q(n12308) );
  OR2X1 U12016 ( .IN1(n12261), .IN2(n12241), .Q(n12309) );
  OR2X1 U12017 ( .IN1(n12310), .IN2(n12241), .Q(n12306) );
  OR2X1 U12018 ( .IN1(n12311), .IN2(n12312), .Q(n12310) );
  OR2X1 U12019 ( .IN1(n12261), .IN2(n12313), .Q(n12312) );
  AND2X1 U12020 ( .IN1(n12314), .IN2(n12241), .Q(n12313) );
  OR2X1 U12021 ( .IN1(n12315), .IN2(n12316), .Q(n12311) );
  AND2X1 U12022 ( .IN1(n12317), .IN2(n12227), .Q(n12316) );
  AND2X1 U12023 ( .IN1(n12318), .IN2(n12235), .Q(n12317) );
  OR2X1 U12024 ( .IN1(n12319), .IN2(n12248), .Q(n12318) );
  AND2X1 U12025 ( .IN1(n12238), .IN2(n12249), .Q(n12319) );
  AND2X1 U12026 ( .IN1(n12226), .IN2(n12320), .Q(n12315) );
  OR2X1 U12027 ( .IN1(n12321), .IN2(n10191), .Q(n12320) );
  OR2X1 U12028 ( .IN1(n12322), .IN2(n12323), .Q(g30338) );
  AND2X1 U12029 ( .IN1(n4511), .IN2(g1701), .Q(n12323) );
  AND2X1 U12030 ( .IN1(n12268), .IN2(n4618), .Q(n12322) );
  AND2X1 U12031 ( .IN1(n11758), .IN2(n12324), .Q(n12268) );
  AND2X1 U12032 ( .IN1(n12325), .IN2(n12326), .Q(n12324) );
  INVX0 U12033 ( .INP(n12327), .ZN(n12326) );
  AND2X1 U12034 ( .IN1(n12328), .IN2(n12329), .Q(n12327) );
  OR2X1 U12035 ( .IN1(n11798), .IN2(n11778), .Q(n12328) );
  OR2X1 U12036 ( .IN1(n12329), .IN2(n11778), .Q(n12325) );
  OR2X1 U12037 ( .IN1(n12330), .IN2(n12331), .Q(n12329) );
  OR2X1 U12038 ( .IN1(n11798), .IN2(n12332), .Q(n12331) );
  AND2X1 U12039 ( .IN1(n12333), .IN2(n11778), .Q(n12332) );
  OR2X1 U12040 ( .IN1(n12334), .IN2(n12335), .Q(n12330) );
  AND2X1 U12041 ( .IN1(n12336), .IN2(n11764), .Q(n12335) );
  AND2X1 U12042 ( .IN1(n12337), .IN2(n11772), .Q(n12336) );
  OR2X1 U12043 ( .IN1(n12338), .IN2(n11785), .Q(n12337) );
  AND2X1 U12044 ( .IN1(n11775), .IN2(n11786), .Q(n12338) );
  AND2X1 U12045 ( .IN1(n11763), .IN2(n12339), .Q(n12334) );
  OR2X1 U12046 ( .IN1(n4386), .IN2(n12340), .Q(n12339) );
  OR2X1 U12047 ( .IN1(n12341), .IN2(n12342), .Q(g30304) );
  AND2X1 U12048 ( .IN1(n12343), .IN2(g2241), .Q(n12342) );
  AND2X1 U12049 ( .IN1(n4367), .IN2(g2285), .Q(n12341) );
  OR2X1 U12050 ( .IN1(n12344), .IN2(n12345), .Q(g30303) );
  AND2X1 U12051 ( .IN1(test_so73), .IN2(n12343), .Q(n12345) );
  AND2X1 U12052 ( .IN1(g2282), .IN2(n10189), .Q(n12344) );
  OR2X1 U12053 ( .IN1(n12346), .IN2(n12347), .Q(g30302) );
  AND2X1 U12054 ( .IN1(n12348), .IN2(g1547), .Q(n12347) );
  AND2X1 U12055 ( .IN1(n4368), .IN2(g1591), .Q(n12346) );
  OR2X1 U12056 ( .IN1(n12349), .IN2(n12350), .Q(g30301) );
  AND2X1 U12057 ( .IN1(n12343), .IN2(g6837), .Q(n12350) );
  OR2X1 U12058 ( .IN1(n12351), .IN2(n12352), .Q(n12343) );
  AND2X1 U12059 ( .IN1(n11872), .IN2(g2185), .Q(n12352) );
  AND2X1 U12060 ( .IN1(n12353), .IN2(n11874), .Q(n12351) );
  AND2X1 U12061 ( .IN1(n12354), .IN2(n12355), .Q(n12353) );
  OR2X1 U12062 ( .IN1(n12356), .IN2(n10855), .Q(n12355) );
  OR2X1 U12063 ( .IN1(n10854), .IN2(n12357), .Q(n12354) );
  AND2X1 U12064 ( .IN1(n4324), .IN2(g2279), .Q(n12349) );
  OR2X1 U12065 ( .IN1(n12358), .IN2(n12359), .Q(g30300) );
  AND2X1 U12066 ( .IN1(n12360), .IN2(g2241), .Q(n12359) );
  AND2X1 U12067 ( .IN1(n4367), .IN2(g2267), .Q(n12358) );
  OR2X1 U12068 ( .IN1(n12361), .IN2(n12362), .Q(g30299) );
  AND2X1 U12069 ( .IN1(n12348), .IN2(g6782), .Q(n12362) );
  AND2X1 U12070 ( .IN1(n4515), .IN2(g1588), .Q(n12361) );
  OR2X1 U12071 ( .IN1(n12363), .IN2(n12364), .Q(g30298) );
  AND2X1 U12072 ( .IN1(test_so31), .IN2(n12365), .Q(n12364) );
  AND2X1 U12073 ( .IN1(g897), .IN2(n10188), .Q(n12363) );
  OR2X1 U12074 ( .IN1(n12366), .IN2(n12367), .Q(g30297) );
  AND2X1 U12075 ( .IN1(n12368), .IN2(g2241), .Q(n12367) );
  AND2X1 U12076 ( .IN1(n4367), .IN2(g2339), .Q(n12366) );
  OR2X1 U12077 ( .IN1(n12369), .IN2(n12370), .Q(g30296) );
  AND2X1 U12078 ( .IN1(test_so73), .IN2(n12360), .Q(n12370) );
  AND2X1 U12079 ( .IN1(test_so76), .IN2(n10189), .Q(n12369) );
  OR2X1 U12080 ( .IN1(n12371), .IN2(n12372), .Q(g30295) );
  AND2X1 U12081 ( .IN1(n12348), .IN2(g6573), .Q(n12372) );
  OR2X1 U12082 ( .IN1(n12373), .IN2(n12374), .Q(n12348) );
  AND2X1 U12083 ( .IN1(n11907), .IN2(g1491), .Q(n12374) );
  AND2X1 U12084 ( .IN1(n12375), .IN2(n11909), .Q(n12373) );
  AND2X1 U12085 ( .IN1(n12376), .IN2(n12377), .Q(n12375) );
  OR2X1 U12086 ( .IN1(n12378), .IN2(n10805), .Q(n12377) );
  OR2X1 U12087 ( .IN1(n10804), .IN2(n12379), .Q(n12376) );
  AND2X1 U12088 ( .IN1(n4317), .IN2(g1585), .Q(n12371) );
  OR2X1 U12089 ( .IN1(n12380), .IN2(n12381), .Q(g30294) );
  AND2X1 U12090 ( .IN1(n12382), .IN2(g1547), .Q(n12381) );
  AND2X1 U12091 ( .IN1(n4368), .IN2(g1573), .Q(n12380) );
  OR2X1 U12092 ( .IN1(n12383), .IN2(n12384), .Q(g30293) );
  AND2X1 U12093 ( .IN1(n12365), .IN2(g6518), .Q(n12384) );
  AND2X1 U12094 ( .IN1(n4312), .IN2(g894), .Q(n12383) );
  OR2X1 U12095 ( .IN1(n12385), .IN2(n12386), .Q(g30292) );
  AND2X1 U12096 ( .IN1(n12387), .IN2(g165), .Q(n12386) );
  AND2X1 U12097 ( .IN1(n4369), .IN2(g210), .Q(n12385) );
  OR2X1 U12098 ( .IN1(n12388), .IN2(n12389), .Q(g30291) );
  AND2X1 U12099 ( .IN1(test_so73), .IN2(n12368), .Q(n12389) );
  AND2X1 U12100 ( .IN1(g2336), .IN2(n10189), .Q(n12388) );
  OR2X1 U12101 ( .IN1(n12390), .IN2(n12391), .Q(g30290) );
  AND2X1 U12102 ( .IN1(n12392), .IN2(g2241), .Q(n12391) );
  AND2X1 U12103 ( .IN1(n4367), .IN2(g2330), .Q(n12390) );
  OR2X1 U12104 ( .IN1(n12393), .IN2(n12394), .Q(g30289) );
  AND2X1 U12105 ( .IN1(n12360), .IN2(g6837), .Q(n12394) );
  OR2X1 U12106 ( .IN1(n12395), .IN2(n12396), .Q(n12360) );
  AND2X1 U12107 ( .IN1(n11872), .IN2(g2165), .Q(n12396) );
  AND2X1 U12108 ( .IN1(n11874), .IN2(n12397), .Q(n12395) );
  OR2X1 U12109 ( .IN1(n12398), .IN2(n12399), .Q(n12397) );
  AND2X1 U12110 ( .IN1(n12400), .IN2(n10845), .Q(n12399) );
  AND2X1 U12111 ( .IN1(n10844), .IN2(n12401), .Q(n12398) );
  INVX0 U12112 ( .INP(n12400), .ZN(n12401) );
  AND2X1 U12113 ( .IN1(n4324), .IN2(g2261), .Q(n12393) );
  OR2X1 U12114 ( .IN1(n12402), .IN2(n12403), .Q(g30288) );
  AND2X1 U12115 ( .IN1(n12404), .IN2(g1547), .Q(n12403) );
  AND2X1 U12116 ( .IN1(n4368), .IN2(g1645), .Q(n12402) );
  OR2X1 U12117 ( .IN1(n12405), .IN2(n12406), .Q(g30287) );
  AND2X1 U12118 ( .IN1(n12382), .IN2(g6782), .Q(n12406) );
  AND2X1 U12119 ( .IN1(n4515), .IN2(g1570), .Q(n12405) );
  OR2X1 U12120 ( .IN1(n12407), .IN2(n12408), .Q(g30286) );
  AND2X1 U12121 ( .IN1(n12365), .IN2(g6368), .Q(n12408) );
  OR2X1 U12122 ( .IN1(n12409), .IN2(n12410), .Q(n12365) );
  AND2X1 U12123 ( .IN1(n11951), .IN2(g801), .Q(n12410) );
  AND2X1 U12124 ( .IN1(n12411), .IN2(n11946), .Q(n12409) );
  AND2X1 U12125 ( .IN1(n12412), .IN2(n12413), .Q(n12411) );
  OR2X1 U12126 ( .IN1(n12414), .IN2(n10726), .Q(n12413) );
  OR2X1 U12127 ( .IN1(n10725), .IN2(n12415), .Q(n12412) );
  AND2X1 U12128 ( .IN1(n4323), .IN2(g891), .Q(n12407) );
  OR2X1 U12129 ( .IN1(n12416), .IN2(n12417), .Q(g30285) );
  AND2X1 U12130 ( .IN1(test_so31), .IN2(n12418), .Q(n12417) );
  AND2X1 U12131 ( .IN1(g879), .IN2(n10188), .Q(n12416) );
  OR2X1 U12132 ( .IN1(n12419), .IN2(n12420), .Q(g30284) );
  AND2X1 U12133 ( .IN1(n12387), .IN2(g6313), .Q(n12420) );
  AND2X1 U12134 ( .IN1(n4512), .IN2(g207), .Q(n12419) );
  OR2X1 U12135 ( .IN1(n12421), .IN2(n12422), .Q(g30283) );
  AND2X1 U12136 ( .IN1(n12368), .IN2(g6837), .Q(n12422) );
  OR2X1 U12137 ( .IN1(n12423), .IN2(n12424), .Q(n12368) );
  AND2X1 U12138 ( .IN1(n11872), .IN2(g2200), .Q(n12424) );
  AND2X1 U12139 ( .IN1(n12425), .IN2(n12426), .Q(n12423) );
  AND2X1 U12140 ( .IN1(n12427), .IN2(n12428), .Q(n12426) );
  OR2X1 U12141 ( .IN1(n12429), .IN2(n10829), .Q(n12428) );
  INVX0 U12142 ( .INP(n12089), .ZN(n12429) );
  OR2X1 U12143 ( .IN1(n10828), .IN2(n12089), .Q(n12427) );
  OR2X1 U12144 ( .IN1(n12430), .IN2(n12431), .Q(n12089) );
  AND2X1 U12145 ( .IN1(n12432), .IN2(n12433), .Q(n12430) );
  OR2X1 U12146 ( .IN1(n4529), .IN2(n10859), .Q(n12433) );
  OR2X1 U12147 ( .IN1(n10858), .IN2(n11593), .Q(n12432) );
  AND2X1 U12148 ( .IN1(n4324), .IN2(g2333), .Q(n12421) );
  OR2X1 U12149 ( .IN1(n12434), .IN2(n12435), .Q(g30282) );
  AND2X1 U12150 ( .IN1(test_so73), .IN2(n12392), .Q(n12435) );
  AND2X1 U12151 ( .IN1(test_so77), .IN2(n10189), .Q(n12434) );
  OR2X1 U12152 ( .IN1(n12436), .IN2(n12437), .Q(g30281) );
  AND2X1 U12153 ( .IN1(n12404), .IN2(g6782), .Q(n12437) );
  AND2X1 U12154 ( .IN1(n4515), .IN2(g1642), .Q(n12436) );
  OR2X1 U12155 ( .IN1(n12438), .IN2(n12439), .Q(g30280) );
  AND2X1 U12156 ( .IN1(n12440), .IN2(g1547), .Q(n12439) );
  AND2X1 U12157 ( .IN1(n4368), .IN2(g1636), .Q(n12438) );
  OR2X1 U12158 ( .IN1(n12441), .IN2(n12442), .Q(g30279) );
  AND2X1 U12159 ( .IN1(n12382), .IN2(g6573), .Q(n12442) );
  OR2X1 U12160 ( .IN1(n12443), .IN2(n12444), .Q(n12382) );
  AND2X1 U12161 ( .IN1(n11907), .IN2(g1471), .Q(n12444) );
  AND2X1 U12162 ( .IN1(n11909), .IN2(n12445), .Q(n12443) );
  OR2X1 U12163 ( .IN1(n12446), .IN2(n12447), .Q(n12445) );
  AND2X1 U12164 ( .IN1(n12448), .IN2(n10772), .Q(n12447) );
  AND2X1 U12165 ( .IN1(n10771), .IN2(n12449), .Q(n12446) );
  INVX0 U12166 ( .INP(n12448), .ZN(n12449) );
  AND2X1 U12167 ( .IN1(n4317), .IN2(g1567), .Q(n12441) );
  OR2X1 U12168 ( .IN1(n12450), .IN2(n12451), .Q(g30278) );
  AND2X1 U12169 ( .IN1(test_so31), .IN2(n12452), .Q(n12451) );
  AND2X1 U12170 ( .IN1(g951), .IN2(n10188), .Q(n12450) );
  OR2X1 U12171 ( .IN1(n12453), .IN2(n12454), .Q(g30277) );
  AND2X1 U12172 ( .IN1(n12418), .IN2(g6518), .Q(n12454) );
  AND2X1 U12173 ( .IN1(n4312), .IN2(g876), .Q(n12453) );
  OR2X1 U12174 ( .IN1(n12455), .IN2(n12456), .Q(g30276) );
  AND2X1 U12175 ( .IN1(n12387), .IN2(g6231), .Q(n12456) );
  OR2X1 U12176 ( .IN1(n12457), .IN2(n12458), .Q(n12387) );
  AND2X1 U12177 ( .IN1(n11998), .IN2(g113), .Q(n12458) );
  AND2X1 U12178 ( .IN1(n12459), .IN2(n11993), .Q(n12457) );
  AND2X1 U12179 ( .IN1(n12460), .IN2(n12461), .Q(n12459) );
  OR2X1 U12180 ( .IN1(n12462), .IN2(n10668), .Q(n12461) );
  OR2X1 U12181 ( .IN1(n10667), .IN2(n12463), .Q(n12460) );
  AND2X1 U12182 ( .IN1(n4318), .IN2(g204), .Q(n12455) );
  OR2X1 U12183 ( .IN1(n12464), .IN2(n12465), .Q(g30275) );
  AND2X1 U12184 ( .IN1(n12466), .IN2(g165), .Q(n12465) );
  AND2X1 U12185 ( .IN1(n4369), .IN2(g192), .Q(n12464) );
  OR2X1 U12186 ( .IN1(n12467), .IN2(n12468), .Q(g30274) );
  AND2X1 U12187 ( .IN1(n12392), .IN2(g6837), .Q(n12468) );
  OR2X1 U12188 ( .IN1(n12469), .IN2(n12470), .Q(n12392) );
  AND2X1 U12189 ( .IN1(n11872), .IN2(g2190), .Q(n12470) );
  AND2X1 U12190 ( .IN1(n12425), .IN2(n12471), .Q(n12469) );
  AND2X1 U12191 ( .IN1(n12472), .IN2(n12473), .Q(n12471) );
  OR2X1 U12192 ( .IN1(n12474), .IN2(n10825), .Q(n12473) );
  AND2X1 U12193 ( .IN1(n12356), .IN2(n12475), .Q(n12474) );
  OR2X1 U12194 ( .IN1(n12476), .IN2(n12477), .Q(n12475) );
  AND2X1 U12195 ( .IN1(n4529), .IN2(n10855), .Q(n12477) );
  AND2X1 U12196 ( .IN1(n10854), .IN2(n11593), .Q(n12476) );
  INVX0 U12197 ( .INP(n12357), .ZN(n12356) );
  OR2X1 U12198 ( .IN1(n10824), .IN2(n12478), .Q(n12472) );
  OR2X1 U12199 ( .IN1(n12479), .IN2(n12480), .Q(n12478) );
  AND2X1 U12200 ( .IN1(n4529), .IN2(n10854), .Q(n12479) );
  AND2X1 U12201 ( .IN1(n11874), .IN2(n12481), .Q(n12425) );
  INVX0 U12202 ( .INP(n12049), .ZN(n12481) );
  AND2X1 U12203 ( .IN1(n4324), .IN2(g2324), .Q(n12467) );
  OR2X1 U12204 ( .IN1(n12482), .IN2(n12483), .Q(g30273) );
  AND2X1 U12205 ( .IN1(n12404), .IN2(g6573), .Q(n12483) );
  OR2X1 U12206 ( .IN1(n12484), .IN2(n12485), .Q(n12404) );
  AND2X1 U12207 ( .IN1(n11907), .IN2(g1506), .Q(n12485) );
  AND2X1 U12208 ( .IN1(n12486), .IN2(n12487), .Q(n12484) );
  AND2X1 U12209 ( .IN1(n12488), .IN2(n12489), .Q(n12487) );
  OR2X1 U12210 ( .IN1(n12490), .IN2(n10764), .Q(n12489) );
  INVX0 U12211 ( .INP(n12141), .ZN(n12490) );
  OR2X1 U12212 ( .IN1(n10763), .IN2(n12141), .Q(n12488) );
  OR2X1 U12213 ( .IN1(n12491), .IN2(n12492), .Q(n12141) );
  AND2X1 U12214 ( .IN1(n12493), .IN2(n12494), .Q(n12491) );
  OR2X1 U12215 ( .IN1(n4530), .IN2(n10798), .Q(n12494) );
  OR2X1 U12216 ( .IN1(n10797), .IN2(n11590), .Q(n12493) );
  AND2X1 U12217 ( .IN1(n4317), .IN2(g1639), .Q(n12482) );
  OR2X1 U12218 ( .IN1(n12495), .IN2(n12496), .Q(g30272) );
  AND2X1 U12219 ( .IN1(n12440), .IN2(g6782), .Q(n12496) );
  AND2X1 U12220 ( .IN1(n4515), .IN2(g1633), .Q(n12495) );
  OR2X1 U12221 ( .IN1(n12497), .IN2(n12498), .Q(g30271) );
  AND2X1 U12222 ( .IN1(n12452), .IN2(g6518), .Q(n12498) );
  AND2X1 U12223 ( .IN1(n4312), .IN2(g948), .Q(n12497) );
  OR2X1 U12224 ( .IN1(n12499), .IN2(n12500), .Q(g30270) );
  AND2X1 U12225 ( .IN1(test_so31), .IN2(n12501), .Q(n12500) );
  AND2X1 U12226 ( .IN1(g942), .IN2(n10188), .Q(n12499) );
  OR2X1 U12227 ( .IN1(n12502), .IN2(n12503), .Q(g30269) );
  AND2X1 U12228 ( .IN1(n12418), .IN2(g6368), .Q(n12503) );
  OR2X1 U12229 ( .IN1(n12504), .IN2(n12505), .Q(n12418) );
  AND2X1 U12230 ( .IN1(n11951), .IN2(g785), .Q(n12505) );
  AND2X1 U12231 ( .IN1(n11946), .IN2(n12506), .Q(n12504) );
  OR2X1 U12232 ( .IN1(n12507), .IN2(n12508), .Q(n12506) );
  AND2X1 U12233 ( .IN1(n12509), .IN2(n10716), .Q(n12508) );
  AND2X1 U12234 ( .IN1(n10715), .IN2(n12510), .Q(n12507) );
  INVX0 U12235 ( .INP(n12509), .ZN(n12510) );
  AND2X1 U12236 ( .IN1(n4323), .IN2(g873), .Q(n12502) );
  OR2X1 U12237 ( .IN1(n12511), .IN2(n12512), .Q(g30268) );
  AND2X1 U12238 ( .IN1(n12513), .IN2(g165), .Q(n12512) );
  AND2X1 U12239 ( .IN1(n4369), .IN2(g264), .Q(n12511) );
  OR2X1 U12240 ( .IN1(n12514), .IN2(n12515), .Q(g30267) );
  AND2X1 U12241 ( .IN1(n12466), .IN2(g6313), .Q(n12515) );
  AND2X1 U12242 ( .IN1(test_so13), .IN2(n4512), .Q(n12514) );
  OR2X1 U12243 ( .IN1(n12516), .IN2(n12517), .Q(g30266) );
  AND2X1 U12244 ( .IN1(n12440), .IN2(g6573), .Q(n12517) );
  OR2X1 U12245 ( .IN1(n12518), .IN2(n12519), .Q(n12440) );
  AND2X1 U12246 ( .IN1(n11907), .IN2(g1496), .Q(n12519) );
  AND2X1 U12247 ( .IN1(n12486), .IN2(n12520), .Q(n12518) );
  AND2X1 U12248 ( .IN1(n12521), .IN2(n12522), .Q(n12520) );
  OR2X1 U12249 ( .IN1(n12523), .IN2(n10760), .Q(n12522) );
  AND2X1 U12250 ( .IN1(n12378), .IN2(n12524), .Q(n12523) );
  OR2X1 U12251 ( .IN1(n12525), .IN2(n12526), .Q(n12524) );
  AND2X1 U12252 ( .IN1(n4530), .IN2(n10805), .Q(n12526) );
  AND2X1 U12253 ( .IN1(n10804), .IN2(n11590), .Q(n12525) );
  INVX0 U12254 ( .INP(n12379), .ZN(n12378) );
  OR2X1 U12255 ( .IN1(n10759), .IN2(n12527), .Q(n12521) );
  OR2X1 U12256 ( .IN1(n12528), .IN2(n12529), .Q(n12527) );
  AND2X1 U12257 ( .IN1(n4530), .IN2(n10804), .Q(n12528) );
  AND2X1 U12258 ( .IN1(n11909), .IN2(n12530), .Q(n12486) );
  INVX0 U12259 ( .INP(n12104), .ZN(n12530) );
  AND2X1 U12260 ( .IN1(n4317), .IN2(g1630), .Q(n12516) );
  OR2X1 U12261 ( .IN1(n12531), .IN2(n12532), .Q(g30265) );
  AND2X1 U12262 ( .IN1(n12452), .IN2(g6368), .Q(n12532) );
  OR2X1 U12263 ( .IN1(n12533), .IN2(n12534), .Q(n12452) );
  AND2X1 U12264 ( .IN1(n11951), .IN2(g813), .Q(n12534) );
  AND2X1 U12265 ( .IN1(n12535), .IN2(n11946), .Q(n12533) );
  AND2X1 U12266 ( .IN1(n12536), .IN2(n12537), .Q(n12535) );
  OR2X1 U12267 ( .IN1(n12538), .IN2(n10741), .Q(n12537) );
  AND2X1 U12268 ( .IN1(n12539), .IN2(n12540), .Q(n12538) );
  OR2X1 U12269 ( .IN1(n12541), .IN2(n12542), .Q(n12540) );
  AND2X1 U12270 ( .IN1(n11981), .IN2(n10708), .Q(n12542) );
  AND2X1 U12271 ( .IN1(n10707), .IN2(n11982), .Q(n12541) );
  OR2X1 U12272 ( .IN1(n10740), .IN2(n12543), .Q(n12536) );
  OR2X1 U12273 ( .IN1(n12544), .IN2(n12186), .Q(n12543) );
  OR2X1 U12274 ( .IN1(n12545), .IN2(n12546), .Q(n12186) );
  AND2X1 U12275 ( .IN1(n11982), .IN2(n10708), .Q(n12545) );
  AND2X1 U12276 ( .IN1(n11981), .IN2(n10707), .Q(n12544) );
  AND2X1 U12277 ( .IN1(test_so35), .IN2(n4323), .Q(n12531) );
  OR2X1 U12278 ( .IN1(n12547), .IN2(n12548), .Q(g30264) );
  AND2X1 U12279 ( .IN1(n12501), .IN2(g6518), .Q(n12548) );
  AND2X1 U12280 ( .IN1(n4312), .IN2(g939), .Q(n12547) );
  OR2X1 U12281 ( .IN1(n12549), .IN2(n12550), .Q(g30263) );
  AND2X1 U12282 ( .IN1(n12513), .IN2(g6313), .Q(n12550) );
  AND2X1 U12283 ( .IN1(n4512), .IN2(g261), .Q(n12549) );
  OR2X1 U12284 ( .IN1(n12551), .IN2(n12552), .Q(g30262) );
  AND2X1 U12285 ( .IN1(n12553), .IN2(g165), .Q(n12552) );
  AND2X1 U12286 ( .IN1(n4369), .IN2(test_so14), .Q(n12551) );
  OR2X1 U12287 ( .IN1(n12554), .IN2(n12555), .Q(g30261) );
  AND2X1 U12288 ( .IN1(n12466), .IN2(g6231), .Q(n12555) );
  OR2X1 U12289 ( .IN1(n12556), .IN2(n12557), .Q(n12466) );
  AND2X1 U12290 ( .IN1(n11998), .IN2(g97), .Q(n12557) );
  AND2X1 U12291 ( .IN1(n11993), .IN2(n12558), .Q(n12556) );
  OR2X1 U12292 ( .IN1(n12559), .IN2(n12560), .Q(n12558) );
  AND2X1 U12293 ( .IN1(n4513), .IN2(n12561), .Q(n12560) );
  INVX0 U12294 ( .INP(n12562), .ZN(n12561) );
  AND2X1 U12295 ( .IN1(n12562), .IN2(n10660), .Q(n12559) );
  AND2X1 U12296 ( .IN1(n4318), .IN2(g186), .Q(n12554) );
  OR2X1 U12297 ( .IN1(n12563), .IN2(n12564), .Q(g30260) );
  AND2X1 U12298 ( .IN1(n12565), .IN2(g2241), .Q(n12564) );
  AND2X1 U12299 ( .IN1(n4367), .IN2(g2294), .Q(n12563) );
  OR2X1 U12300 ( .IN1(n12566), .IN2(n12567), .Q(g30259) );
  AND2X1 U12301 ( .IN1(n12501), .IN2(g6368), .Q(n12567) );
  OR2X1 U12302 ( .IN1(n12568), .IN2(n12569), .Q(n12501) );
  AND2X1 U12303 ( .IN1(n11951), .IN2(g805), .Q(n12569) );
  AND2X1 U12304 ( .IN1(n12570), .IN2(n11946), .Q(n12568) );
  AND2X1 U12305 ( .IN1(n12571), .IN2(n12572), .Q(n12570) );
  OR2X1 U12306 ( .IN1(n12573), .IN2(n10696), .Q(n12572) );
  AND2X1 U12307 ( .IN1(n12414), .IN2(n12574), .Q(n12573) );
  OR2X1 U12308 ( .IN1(n12575), .IN2(n12576), .Q(n12574) );
  AND2X1 U12309 ( .IN1(n11981), .IN2(n10726), .Q(n12576) );
  AND2X1 U12310 ( .IN1(n10725), .IN2(n11982), .Q(n12575) );
  INVX0 U12311 ( .INP(n12415), .ZN(n12414) );
  OR2X1 U12312 ( .IN1(n10695), .IN2(n12577), .Q(n12571) );
  OR2X1 U12313 ( .IN1(n12578), .IN2(n12579), .Q(n12577) );
  AND2X1 U12314 ( .IN1(n11981), .IN2(n10725), .Q(n12578) );
  AND2X1 U12315 ( .IN1(n4323), .IN2(g936), .Q(n12566) );
  OR2X1 U12316 ( .IN1(n12580), .IN2(n12581), .Q(g30258) );
  AND2X1 U12317 ( .IN1(n12513), .IN2(g6231), .Q(n12581) );
  OR2X1 U12318 ( .IN1(n12582), .IN2(n12583), .Q(n12513) );
  AND2X1 U12319 ( .IN1(n11998), .IN2(g125), .Q(n12583) );
  AND2X1 U12320 ( .IN1(n12584), .IN2(n11993), .Q(n12582) );
  AND2X1 U12321 ( .IN1(n12585), .IN2(n12586), .Q(n12584) );
  OR2X1 U12322 ( .IN1(n12587), .IN2(n10635), .Q(n12586) );
  INVX0 U12323 ( .INP(n12215), .ZN(n12587) );
  OR2X1 U12324 ( .IN1(n10634), .IN2(n12215), .Q(n12585) );
  OR2X1 U12325 ( .IN1(n12588), .IN2(n12589), .Q(n12215) );
  AND2X1 U12326 ( .IN1(n12590), .IN2(n12591), .Q(n12588) );
  OR2X1 U12327 ( .IN1(n11586), .IN2(n10643), .Q(n12591) );
  OR2X1 U12328 ( .IN1(n10642), .IN2(n11587), .Q(n12590) );
  AND2X1 U12329 ( .IN1(n4318), .IN2(g258), .Q(n12580) );
  OR2X1 U12330 ( .IN1(n12592), .IN2(n12593), .Q(g30257) );
  AND2X1 U12331 ( .IN1(n12553), .IN2(g6313), .Q(n12593) );
  AND2X1 U12332 ( .IN1(n4512), .IN2(g252), .Q(n12592) );
  OR2X1 U12333 ( .IN1(n12594), .IN2(n12595), .Q(g30256) );
  AND2X1 U12334 ( .IN1(test_so73), .IN2(n12565), .Q(n12595) );
  AND2X1 U12335 ( .IN1(g2291), .IN2(n10189), .Q(n12594) );
  OR2X1 U12336 ( .IN1(n12596), .IN2(n12597), .Q(g30255) );
  AND2X1 U12337 ( .IN1(n12598), .IN2(g1547), .Q(n12597) );
  AND2X1 U12338 ( .IN1(n4368), .IN2(g1600), .Q(n12596) );
  OR2X1 U12339 ( .IN1(n12599), .IN2(n12600), .Q(g30254) );
  AND2X1 U12340 ( .IN1(n12553), .IN2(g6231), .Q(n12600) );
  OR2X1 U12341 ( .IN1(n12601), .IN2(n12602), .Q(n12553) );
  AND2X1 U12342 ( .IN1(n11998), .IN2(g117), .Q(n12602) );
  AND2X1 U12343 ( .IN1(n12603), .IN2(n11993), .Q(n12601) );
  AND2X1 U12344 ( .IN1(n12604), .IN2(n12605), .Q(n12603) );
  OR2X1 U12345 ( .IN1(n12606), .IN2(n10631), .Q(n12605) );
  AND2X1 U12346 ( .IN1(n12462), .IN2(n12607), .Q(n12606) );
  OR2X1 U12347 ( .IN1(n12608), .IN2(n12609), .Q(n12607) );
  AND2X1 U12348 ( .IN1(n11586), .IN2(n10668), .Q(n12609) );
  AND2X1 U12349 ( .IN1(n10667), .IN2(n11587), .Q(n12608) );
  INVX0 U12350 ( .INP(n12463), .ZN(n12462) );
  OR2X1 U12351 ( .IN1(n10630), .IN2(n12610), .Q(n12604) );
  OR2X1 U12352 ( .IN1(n12611), .IN2(n12612), .Q(n12610) );
  AND2X1 U12353 ( .IN1(n11586), .IN2(n10667), .Q(n12611) );
  AND2X1 U12354 ( .IN1(n4318), .IN2(g249), .Q(n12599) );
  OR2X1 U12355 ( .IN1(n12613), .IN2(n12614), .Q(g30253) );
  AND2X1 U12356 ( .IN1(n12565), .IN2(g6837), .Q(n12614) );
  OR2X1 U12357 ( .IN1(n12615), .IN2(n12616), .Q(n12565) );
  AND2X1 U12358 ( .IN1(n11872), .IN2(g2195), .Q(n12616) );
  INVX0 U12359 ( .INP(n12617), .ZN(n11872) );
  OR2X1 U12360 ( .IN1(n11874), .IN2(n12049), .Q(n12617) );
  AND2X1 U12361 ( .IN1(n12618), .IN2(n12619), .Q(n12049) );
  INVX0 U12362 ( .INP(n12620), .ZN(n12619) );
  OR2X1 U12363 ( .IN1(n12400), .IN2(n12621), .Q(n12620) );
  AND2X1 U12364 ( .IN1(n12622), .IN2(n2489), .Q(n12621) );
  AND2X1 U12365 ( .IN1(n12623), .IN2(n11874), .Q(n12615) );
  AND2X1 U12366 ( .IN1(n12624), .IN2(n12618), .Q(n11874) );
  AND2X1 U12367 ( .IN1(n12625), .IN2(n12626), .Q(n12618) );
  AND2X1 U12368 ( .IN1(n12221), .IN2(n12627), .Q(n12626) );
  OR2X1 U12369 ( .IN1(n12628), .IN2(n12261), .Q(n12627) );
  AND2X1 U12370 ( .IN1(n12629), .IN2(n12235), .Q(n12628) );
  OR2X1 U12371 ( .IN1(n12246), .IN2(n12227), .Q(n12629) );
  OR2X1 U12372 ( .IN1(n12239), .IN2(n12630), .Q(n12246) );
  OR2X1 U12373 ( .IN1(n12631), .IN2(n12239), .Q(n12625) );
  OR2X1 U12374 ( .IN1(n12632), .IN2(n12633), .Q(n12239) );
  AND2X1 U12375 ( .IN1(n12634), .IN2(n12635), .Q(n12632) );
  OR2X1 U12376 ( .IN1(n4524), .IN2(g2398), .Q(n12635) );
  AND2X1 U12377 ( .IN1(n12636), .IN2(n12637), .Q(n12634) );
  OR2X1 U12378 ( .IN1(n4516), .IN2(g2397), .Q(n12637) );
  OR2X1 U12379 ( .IN1(n4509), .IN2(g2396), .Q(n12636) );
  OR2X1 U12380 ( .IN1(n12638), .IN2(n12400), .Q(n12624) );
  AND2X1 U12381 ( .IN1(n12639), .IN2(n12622), .Q(n12638) );
  OR2X1 U12382 ( .IN1(n12640), .IN2(n12641), .Q(n12622) );
  OR2X1 U12383 ( .IN1(n12092), .IN2(n12642), .Q(n12641) );
  OR2X1 U12384 ( .IN1(n10862), .IN2(n12643), .Q(n12642) );
  INVX0 U12385 ( .INP(n4529), .ZN(n12092) );
  OR2X1 U12386 ( .IN1(n12644), .IN2(n12645), .Q(n12640) );
  OR2X1 U12387 ( .IN1(n10840), .IN2(n10836), .Q(n12645) );
  OR2X1 U12388 ( .IN1(n12048), .IN2(n10820), .Q(n12644) );
  OR2X1 U12389 ( .IN1(n2489), .IN2(n4529), .Q(n12639) );
  OR2X1 U12390 ( .IN1(n12646), .IN2(n12647), .Q(n2489) );
  OR2X1 U12391 ( .IN1(n12643), .IN2(n12648), .Q(n12647) );
  OR2X1 U12392 ( .IN1(n10837), .IN2(n10821), .Q(n12648) );
  OR2X1 U12393 ( .IN1(n12649), .IN2(n12650), .Q(n12643) );
  OR2X1 U12394 ( .IN1(n10825), .IN2(n10829), .Q(n12650) );
  OR2X1 U12395 ( .IN1(n10845), .IN2(n12651), .Q(n12649) );
  OR2X1 U12396 ( .IN1(n10859), .IN2(n10855), .Q(n12651) );
  OR2X1 U12397 ( .IN1(n10841), .IN2(n12652), .Q(n12646) );
  OR2X1 U12398 ( .IN1(n10870), .IN2(n10863), .Q(n12652) );
  AND2X1 U12399 ( .IN1(n12653), .IN2(n12654), .Q(n12623) );
  OR2X1 U12400 ( .IN1(n12655), .IN2(n10859), .Q(n12654) );
  INVX0 U12401 ( .INP(n12431), .ZN(n12655) );
  OR2X1 U12402 ( .IN1(n10858), .IN2(n12431), .Q(n12653) );
  OR2X1 U12403 ( .IN1(n12480), .IN2(n12656), .Q(n12431) );
  OR2X1 U12404 ( .IN1(n12657), .IN2(n12658), .Q(n12656) );
  AND2X1 U12405 ( .IN1(n4529), .IN2(n10824), .Q(n12658) );
  AND2X1 U12406 ( .IN1(n10854), .IN2(n10825), .Q(n12657) );
  OR2X1 U12407 ( .IN1(n12659), .IN2(n12357), .Q(n12480) );
  OR2X1 U12408 ( .IN1(n12011), .IN2(n12660), .Q(n12357) );
  OR2X1 U12409 ( .IN1(n12661), .IN2(n12662), .Q(n12660) );
  AND2X1 U12410 ( .IN1(n4529), .IN2(n10840), .Q(n12662) );
  AND2X1 U12411 ( .IN1(n10862), .IN2(n10841), .Q(n12661) );
  OR2X1 U12412 ( .IN1(n12663), .IN2(n11878), .Q(n12011) );
  OR2X1 U12413 ( .IN1(n12664), .IN2(n12047), .Q(n11878) );
  OR2X1 U12414 ( .IN1(n12400), .IN2(n12665), .Q(n12047) );
  AND2X1 U12415 ( .IN1(n12666), .IN2(n12667), .Q(n12665) );
  OR2X1 U12416 ( .IN1(n4529), .IN2(n10845), .Q(n12667) );
  OR2X1 U12417 ( .IN1(n10844), .IN2(n11593), .Q(n12666) );
  AND2X1 U12418 ( .IN1(n11593), .IN2(n10871), .Q(n12400) );
  AND2X1 U12419 ( .IN1(n12668), .IN2(n12669), .Q(n12664) );
  OR2X1 U12420 ( .IN1(n4529), .IN2(n10870), .Q(n12669) );
  OR2X1 U12421 ( .IN1(n12048), .IN2(n11593), .Q(n12668) );
  AND2X1 U12422 ( .IN1(n11593), .IN2(n10863), .Q(n12663) );
  AND2X1 U12423 ( .IN1(n11593), .IN2(n10855), .Q(n12659) );
  AND2X1 U12424 ( .IN1(n4324), .IN2(g2288), .Q(n12613) );
  OR2X1 U12425 ( .IN1(n12670), .IN2(n12671), .Q(g30252) );
  AND2X1 U12426 ( .IN1(n12598), .IN2(g6782), .Q(n12671) );
  AND2X1 U12427 ( .IN1(n4515), .IN2(g1597), .Q(n12670) );
  OR2X1 U12428 ( .IN1(n12672), .IN2(n12673), .Q(g30251) );
  AND2X1 U12429 ( .IN1(test_so31), .IN2(n12674), .Q(n12673) );
  AND2X1 U12430 ( .IN1(g906), .IN2(n10188), .Q(n12672) );
  OR2X1 U12431 ( .IN1(n12675), .IN2(n12676), .Q(g30250) );
  AND2X1 U12432 ( .IN1(n12598), .IN2(g6573), .Q(n12676) );
  OR2X1 U12433 ( .IN1(n12677), .IN2(n12678), .Q(n12598) );
  AND2X1 U12434 ( .IN1(n11907), .IN2(g1501), .Q(n12678) );
  INVX0 U12435 ( .INP(n12679), .ZN(n11907) );
  OR2X1 U12436 ( .IN1(n11909), .IN2(n12104), .Q(n12679) );
  AND2X1 U12437 ( .IN1(n12680), .IN2(n12681), .Q(n12104) );
  INVX0 U12438 ( .INP(n12682), .ZN(n12681) );
  OR2X1 U12439 ( .IN1(n12448), .IN2(n12683), .Q(n12682) );
  AND2X1 U12440 ( .IN1(n12684), .IN2(n10806), .Q(n12683) );
  AND2X1 U12441 ( .IN1(n12685), .IN2(n11909), .Q(n12677) );
  AND2X1 U12442 ( .IN1(n12686), .IN2(n12680), .Q(n11909) );
  AND2X1 U12443 ( .IN1(n12687), .IN2(n12688), .Q(n12680) );
  AND2X1 U12444 ( .IN1(n11758), .IN2(n12689), .Q(n12688) );
  OR2X1 U12445 ( .IN1(n12690), .IN2(n11798), .Q(n12689) );
  AND2X1 U12446 ( .IN1(n12691), .IN2(n11772), .Q(n12690) );
  OR2X1 U12447 ( .IN1(n11783), .IN2(n11764), .Q(n12691) );
  OR2X1 U12448 ( .IN1(n11776), .IN2(n12692), .Q(n11783) );
  OR2X1 U12449 ( .IN1(n12693), .IN2(n11776), .Q(n12687) );
  OR2X1 U12450 ( .IN1(n12694), .IN2(n12695), .Q(n11776) );
  AND2X1 U12451 ( .IN1(n12696), .IN2(n12697), .Q(n12694) );
  OR2X1 U12452 ( .IN1(n4525), .IN2(g1704), .Q(n12697) );
  AND2X1 U12453 ( .IN1(n12698), .IN2(n12699), .Q(n12696) );
  OR2X1 U12454 ( .IN1(n4518), .IN2(g1703), .Q(n12699) );
  OR2X1 U12455 ( .IN1(n4511), .IN2(g1702), .Q(n12698) );
  OR2X1 U12456 ( .IN1(n12700), .IN2(n12448), .Q(n12686) );
  AND2X1 U12457 ( .IN1(n12701), .IN2(n12684), .Q(n12700) );
  OR2X1 U12458 ( .IN1(n12702), .IN2(n12703), .Q(n12684) );
  OR2X1 U12459 ( .IN1(n12144), .IN2(n12704), .Q(n12703) );
  OR2X1 U12460 ( .IN1(n10789), .IN2(n12705), .Q(n12704) );
  INVX0 U12461 ( .INP(n4530), .ZN(n12144) );
  OR2X1 U12462 ( .IN1(n12706), .IN2(n12707), .Q(n12702) );
  OR2X1 U12463 ( .IN1(n10779), .IN2(n10793), .Q(n12707) );
  OR2X1 U12464 ( .IN1(n10755), .IN2(n10775), .Q(n12706) );
  OR2X1 U12465 ( .IN1(n10806), .IN2(n4530), .Q(n12701) );
  OR2X1 U12466 ( .IN1(n12708), .IN2(n12709), .Q(n10806) );
  OR2X1 U12467 ( .IN1(n12705), .IN2(n12710), .Q(n12709) );
  OR2X1 U12468 ( .IN1(n10780), .IN2(n10756), .Q(n12710) );
  OR2X1 U12469 ( .IN1(n12711), .IN2(n12712), .Q(n12705) );
  OR2X1 U12470 ( .IN1(n10760), .IN2(n10764), .Q(n12712) );
  OR2X1 U12471 ( .IN1(n10772), .IN2(n12713), .Q(n12711) );
  OR2X1 U12472 ( .IN1(n10805), .IN2(n10798), .Q(n12713) );
  OR2X1 U12473 ( .IN1(n10776), .IN2(n12714), .Q(n12708) );
  OR2X1 U12474 ( .IN1(n10794), .IN2(n10790), .Q(n12714) );
  AND2X1 U12475 ( .IN1(n12715), .IN2(n12716), .Q(n12685) );
  OR2X1 U12476 ( .IN1(n12717), .IN2(n10798), .Q(n12716) );
  INVX0 U12477 ( .INP(n12492), .ZN(n12717) );
  OR2X1 U12478 ( .IN1(n10797), .IN2(n12492), .Q(n12715) );
  OR2X1 U12479 ( .IN1(n12529), .IN2(n12718), .Q(n12492) );
  OR2X1 U12480 ( .IN1(n12719), .IN2(n12720), .Q(n12718) );
  AND2X1 U12481 ( .IN1(n4530), .IN2(n10759), .Q(n12720) );
  AND2X1 U12482 ( .IN1(n10804), .IN2(n10760), .Q(n12719) );
  OR2X1 U12483 ( .IN1(n12721), .IN2(n12379), .Q(n12529) );
  OR2X1 U12484 ( .IN1(n12064), .IN2(n12722), .Q(n12379) );
  OR2X1 U12485 ( .IN1(n12723), .IN2(n12724), .Q(n12722) );
  AND2X1 U12486 ( .IN1(n4530), .IN2(n10779), .Q(n12724) );
  AND2X1 U12487 ( .IN1(n10789), .IN2(n10780), .Q(n12723) );
  OR2X1 U12488 ( .IN1(n12725), .IN2(n11913), .Q(n12064) );
  OR2X1 U12489 ( .IN1(n12726), .IN2(n12103), .Q(n11913) );
  OR2X1 U12490 ( .IN1(n12448), .IN2(n12727), .Q(n12103) );
  AND2X1 U12491 ( .IN1(n12728), .IN2(n12729), .Q(n12727) );
  OR2X1 U12492 ( .IN1(n4530), .IN2(n10772), .Q(n12729) );
  OR2X1 U12493 ( .IN1(n10771), .IN2(n11590), .Q(n12728) );
  AND2X1 U12494 ( .IN1(n11590), .IN2(n10807), .Q(n12448) );
  AND2X1 U12495 ( .IN1(n12730), .IN2(n12731), .Q(n12726) );
  OR2X1 U12496 ( .IN1(n4530), .IN2(n10756), .Q(n12731) );
  OR2X1 U12497 ( .IN1(n10755), .IN2(n11590), .Q(n12730) );
  AND2X1 U12498 ( .IN1(n11590), .IN2(n10790), .Q(n12725) );
  AND2X1 U12499 ( .IN1(n11590), .IN2(n10805), .Q(n12721) );
  AND2X1 U12500 ( .IN1(n4317), .IN2(g1594), .Q(n12675) );
  OR2X1 U12501 ( .IN1(n12732), .IN2(n12733), .Q(g30249) );
  AND2X1 U12502 ( .IN1(n12674), .IN2(g6518), .Q(n12733) );
  AND2X1 U12503 ( .IN1(n4312), .IN2(g903), .Q(n12732) );
  OR2X1 U12504 ( .IN1(n12734), .IN2(n12735), .Q(g30248) );
  AND2X1 U12505 ( .IN1(n12736), .IN2(g165), .Q(n12735) );
  AND2X1 U12506 ( .IN1(n4369), .IN2(g219), .Q(n12734) );
  OR2X1 U12507 ( .IN1(n12737), .IN2(n12738), .Q(g30247) );
  AND2X1 U12508 ( .IN1(n12674), .IN2(g6368), .Q(n12738) );
  OR2X1 U12509 ( .IN1(n12739), .IN2(n12740), .Q(n12674) );
  AND2X1 U12510 ( .IN1(n11951), .IN2(g809), .Q(n12740) );
  INVX0 U12511 ( .INP(n12741), .ZN(n11951) );
  OR2X1 U12512 ( .IN1(n12156), .IN2(n11946), .Q(n12741) );
  AND2X1 U12513 ( .IN1(n12742), .IN2(n12743), .Q(n12156) );
  INVX0 U12514 ( .INP(n12744), .ZN(n12742) );
  AND2X1 U12515 ( .IN1(n12745), .IN2(n11946), .Q(n12739) );
  AND2X1 U12516 ( .IN1(n12746), .IN2(n12743), .Q(n11946) );
  AND2X1 U12517 ( .IN1(n12747), .IN2(n12748), .Q(n12743) );
  AND2X1 U12518 ( .IN1(n12749), .IN2(n12750), .Q(n12748) );
  OR2X1 U12519 ( .IN1(n12751), .IN2(n11569), .Q(n12750) );
  AND2X1 U12520 ( .IN1(n12752), .IN2(n11577), .Q(n12751) );
  OR2X1 U12521 ( .IN1(n11611), .IN2(n11575), .Q(n12752) );
  OR2X1 U12522 ( .IN1(n12753), .IN2(n11606), .Q(n11611) );
  OR2X1 U12523 ( .IN1(n12754), .IN2(n11606), .Q(n12747) );
  OR2X1 U12524 ( .IN1(n12755), .IN2(n12756), .Q(n11606) );
  AND2X1 U12525 ( .IN1(n12757), .IN2(n12758), .Q(n12755) );
  OR2X1 U12526 ( .IN1(n4364), .IN2(g1010), .Q(n12758) );
  AND2X1 U12527 ( .IN1(n12759), .IN2(n12760), .Q(n12757) );
  OR2X1 U12528 ( .IN1(n4363), .IN2(g1009), .Q(n12760) );
  OR2X1 U12529 ( .IN1(n4381), .IN2(g1008), .Q(n12759) );
  OR2X1 U12530 ( .IN1(n12744), .IN2(n12761), .Q(n12746) );
  AND2X1 U12531 ( .IN1(n12762), .IN2(n11981), .Q(n12761) );
  OR2X1 U12532 ( .IN1(n12763), .IN2(n12509), .Q(n12744) );
  AND2X1 U12533 ( .IN1(n12762), .IN2(n2542), .Q(n12763) );
  OR2X1 U12534 ( .IN1(n12764), .IN2(n12765), .Q(n2542) );
  OR2X1 U12535 ( .IN1(n12766), .IN2(n12767), .Q(n12765) );
  OR2X1 U12536 ( .IN1(n10692), .IN2(n10700), .Q(n12767) );
  OR2X1 U12537 ( .IN1(n10712), .IN2(n12768), .Q(n12764) );
  OR2X1 U12538 ( .IN1(n10730), .IN2(n10734), .Q(n12768) );
  OR2X1 U12539 ( .IN1(n12769), .IN2(n12770), .Q(n12762) );
  OR2X1 U12540 ( .IN1(n11982), .IN2(n12771), .Q(n12770) );
  OR2X1 U12541 ( .IN1(n10733), .IN2(n12766), .Q(n12771) );
  OR2X1 U12542 ( .IN1(n12772), .IN2(n12773), .Q(n12766) );
  OR2X1 U12543 ( .IN1(n10716), .IN2(n10696), .Q(n12773) );
  OR2X1 U12544 ( .IN1(n10708), .IN2(n12774), .Q(n12772) );
  OR2X1 U12545 ( .IN1(n10741), .IN2(n10726), .Q(n12774) );
  OR2X1 U12546 ( .IN1(n12775), .IN2(n12776), .Q(n12769) );
  OR2X1 U12547 ( .IN1(n10711), .IN2(n10729), .Q(n12776) );
  OR2X1 U12548 ( .IN1(n10699), .IN2(n10691), .Q(n12775) );
  AND2X1 U12549 ( .IN1(n12777), .IN2(n12778), .Q(n12745) );
  OR2X1 U12550 ( .IN1(n12539), .IN2(n10708), .Q(n12778) );
  INVX0 U12551 ( .INP(n12546), .ZN(n12539) );
  OR2X1 U12552 ( .IN1(n10707), .IN2(n12546), .Q(n12777) );
  OR2X1 U12553 ( .IN1(n12579), .IN2(n12779), .Q(n12546) );
  OR2X1 U12554 ( .IN1(n12780), .IN2(n12781), .Q(n12779) );
  AND2X1 U12555 ( .IN1(n11981), .IN2(n10695), .Q(n12781) );
  AND2X1 U12556 ( .IN1(n10725), .IN2(n10696), .Q(n12780) );
  OR2X1 U12557 ( .IN1(n12782), .IN2(n12415), .Q(n12579) );
  OR2X1 U12558 ( .IN1(n12119), .IN2(n12783), .Q(n12415) );
  OR2X1 U12559 ( .IN1(n12784), .IN2(n12785), .Q(n12783) );
  AND2X1 U12560 ( .IN1(n11981), .IN2(n10691), .Q(n12785) );
  INVX0 U12561 ( .INP(n10692), .ZN(n10691) );
  AND2X1 U12562 ( .IN1(n10733), .IN2(n10692), .Q(n12784) );
  OR2X1 U12563 ( .IN1(n12786), .IN2(n11950), .Q(n12119) );
  OR2X1 U12564 ( .IN1(n12787), .IN2(n12155), .Q(n11950) );
  OR2X1 U12565 ( .IN1(n12509), .IN2(n12788), .Q(n12155) );
  AND2X1 U12566 ( .IN1(n12789), .IN2(n12790), .Q(n12788) );
  OR2X1 U12567 ( .IN1(n11981), .IN2(n10716), .Q(n12790) );
  OR2X1 U12568 ( .IN1(n10715), .IN2(n11982), .Q(n12789) );
  AND2X1 U12569 ( .IN1(n11982), .IN2(n10742), .Q(n12509) );
  AND2X1 U12570 ( .IN1(n12791), .IN2(n12792), .Q(n12787) );
  OR2X1 U12571 ( .IN1(n11981), .IN2(n10700), .Q(n12792) );
  OR2X1 U12572 ( .IN1(n10699), .IN2(n11982), .Q(n12791) );
  INVX0 U12573 ( .INP(n10700), .ZN(n10699) );
  AND2X1 U12574 ( .IN1(n11982), .IN2(n10734), .Q(n12786) );
  AND2X1 U12575 ( .IN1(n11982), .IN2(n10726), .Q(n12782) );
  AND2X1 U12576 ( .IN1(n4323), .IN2(g900), .Q(n12737) );
  OR2X1 U12577 ( .IN1(n12793), .IN2(n12794), .Q(g30246) );
  AND2X1 U12578 ( .IN1(n12736), .IN2(g6313), .Q(n12794) );
  AND2X1 U12579 ( .IN1(n4512), .IN2(g216), .Q(n12793) );
  OR2X1 U12580 ( .IN1(n12795), .IN2(n12796), .Q(g30245) );
  AND2X1 U12581 ( .IN1(n12736), .IN2(g6231), .Q(n12796) );
  OR2X1 U12582 ( .IN1(n12797), .IN2(n12798), .Q(n12736) );
  AND2X1 U12583 ( .IN1(n11998), .IN2(g121), .Q(n12798) );
  INVX0 U12584 ( .INP(n12799), .ZN(n11998) );
  OR2X1 U12585 ( .IN1(n12202), .IN2(n11993), .Q(n12799) );
  AND2X1 U12586 ( .IN1(n12800), .IN2(n12801), .Q(n12202) );
  INVX0 U12587 ( .INP(n12802), .ZN(n12800) );
  AND2X1 U12588 ( .IN1(n12803), .IN2(n11993), .Q(n12797) );
  AND2X1 U12589 ( .IN1(n12804), .IN2(n12801), .Q(n11993) );
  AND2X1 U12590 ( .IN1(n12805), .IN2(n12806), .Q(n12801) );
  AND2X1 U12591 ( .IN1(n11811), .IN2(n12807), .Q(n12806) );
  OR2X1 U12592 ( .IN1(n12808), .IN2(n11851), .Q(n12807) );
  AND2X1 U12593 ( .IN1(n12809), .IN2(n11825), .Q(n12808) );
  OR2X1 U12594 ( .IN1(n11836), .IN2(n11817), .Q(n12809) );
  OR2X1 U12595 ( .IN1(n11829), .IN2(n12810), .Q(n11836) );
  OR2X1 U12596 ( .IN1(n12811), .IN2(n11829), .Q(n12805) );
  OR2X1 U12597 ( .IN1(n12812), .IN2(n12813), .Q(n11829) );
  AND2X1 U12598 ( .IN1(n12814), .IN2(n12815), .Q(n12812) );
  OR2X1 U12599 ( .IN1(n4499), .IN2(g323), .Q(n12815) );
  AND2X1 U12600 ( .IN1(n12816), .IN2(n12817), .Q(n12814) );
  OR2X1 U12601 ( .IN1(n4520), .IN2(g322), .Q(n12817) );
  OR2X1 U12602 ( .IN1(n4506), .IN2(g321), .Q(n12816) );
  OR2X1 U12603 ( .IN1(n12802), .IN2(n12818), .Q(n12804) );
  AND2X1 U12604 ( .IN1(n12819), .IN2(n11586), .Q(n12818) );
  OR2X1 U12605 ( .IN1(n12820), .IN2(n12562), .Q(n12802) );
  AND2X1 U12606 ( .IN1(n12819), .IN2(n10677), .Q(n12820) );
  OR2X1 U12607 ( .IN1(n12821), .IN2(n12822), .Q(n10677) );
  OR2X1 U12608 ( .IN1(n12823), .IN2(n12824), .Q(n12822) );
  OR2X1 U12609 ( .IN1(n10651), .IN2(n10627), .Q(n12824) );
  OR2X1 U12610 ( .IN1(n10647), .IN2(n12825), .Q(n12821) );
  OR2X1 U12611 ( .IN1(n10676), .IN2(n10664), .Q(n12825) );
  OR2X1 U12612 ( .IN1(n12826), .IN2(n12827), .Q(n12819) );
  OR2X1 U12613 ( .IN1(n11587), .IN2(n12828), .Q(n12827) );
  OR2X1 U12614 ( .IN1(n10663), .IN2(n12823), .Q(n12828) );
  OR2X1 U12615 ( .IN1(n12829), .IN2(n12830), .Q(n12823) );
  OR2X1 U12616 ( .IN1(n10635), .IN2(n12831), .Q(n12830) );
  OR2X1 U12617 ( .IN1(n10631), .IN2(n12832), .Q(n12829) );
  OR2X1 U12618 ( .IN1(n10668), .IN2(n10643), .Q(n12832) );
  OR2X1 U12619 ( .IN1(n12833), .IN2(n12834), .Q(n12826) );
  OR2X1 U12620 ( .IN1(n10675), .IN2(n10650), .Q(n12834) );
  OR2X1 U12621 ( .IN1(n10626), .IN2(n10646), .Q(n12833) );
  AND2X1 U12622 ( .IN1(n12835), .IN2(n12836), .Q(n12803) );
  OR2X1 U12623 ( .IN1(n12837), .IN2(n10643), .Q(n12836) );
  INVX0 U12624 ( .INP(n12589), .ZN(n12837) );
  OR2X1 U12625 ( .IN1(n10642), .IN2(n12589), .Q(n12835) );
  OR2X1 U12626 ( .IN1(n12612), .IN2(n12838), .Q(n12589) );
  OR2X1 U12627 ( .IN1(n12839), .IN2(n12840), .Q(n12838) );
  AND2X1 U12628 ( .IN1(n11586), .IN2(n10630), .Q(n12840) );
  AND2X1 U12629 ( .IN1(n10667), .IN2(n10631), .Q(n12839) );
  OR2X1 U12630 ( .IN1(n12841), .IN2(n12463), .Q(n12612) );
  OR2X1 U12631 ( .IN1(n12171), .IN2(n12842), .Q(n12463) );
  OR2X1 U12632 ( .IN1(n12843), .IN2(n12844), .Q(n12842) );
  AND2X1 U12633 ( .IN1(n11586), .IN2(n10675), .Q(n12844) );
  AND2X1 U12634 ( .IN1(n10663), .IN2(n10676), .Q(n12843) );
  OR2X1 U12635 ( .IN1(n12845), .IN2(n11997), .Q(n12171) );
  OR2X1 U12636 ( .IN1(n12846), .IN2(n12201), .Q(n11997) );
  OR2X1 U12637 ( .IN1(n12562), .IN2(n12847), .Q(n12201) );
  AND2X1 U12638 ( .IN1(n12848), .IN2(n12849), .Q(n12847) );
  OR2X1 U12639 ( .IN1(n11586), .IN2(n10660), .Q(n12849) );
  OR2X1 U12640 ( .IN1(n4513), .IN2(n11587), .Q(n12848) );
  INVX0 U12641 ( .INP(n10660), .ZN(n4513) );
  OR2X1 U12642 ( .IN1(n12850), .IN2(n12851), .Q(n10660) );
  OR2X1 U12643 ( .IN1(n12852), .IN2(n12853), .Q(n12851) );
  AND2X1 U12644 ( .IN1(g186), .IN2(g6231), .Q(n12853) );
  AND2X1 U12645 ( .IN1(g192), .IN2(g165), .Q(n12852) );
  AND2X1 U12646 ( .IN1(test_so13), .IN2(g6313), .Q(n12850) );
  AND2X1 U12647 ( .IN1(n10678), .IN2(n11587), .Q(n12562) );
  AND2X1 U12648 ( .IN1(n12854), .IN2(n12855), .Q(n12846) );
  OR2X1 U12649 ( .IN1(n11586), .IN2(n10627), .Q(n12855) );
  OR2X1 U12650 ( .IN1(n10626), .IN2(n11587), .Q(n12854) );
  AND2X1 U12651 ( .IN1(n11587), .IN2(n10664), .Q(n12845) );
  AND2X1 U12652 ( .IN1(n11587), .IN2(n10668), .Q(n12841) );
  AND2X1 U12653 ( .IN1(n4318), .IN2(g213), .Q(n12795) );
  OR2X1 U12654 ( .IN1(n12856), .IN2(n12857), .Q(g30072) );
  AND2X1 U12655 ( .IN1(n4543), .IN2(n12858), .Q(n12857) );
  OR2X1 U12656 ( .IN1(n12859), .IN2(n12860), .Q(n12858) );
  AND2X1 U12657 ( .IN1(n12861), .IN2(n7929), .Q(n12860) );
  INVX0 U12658 ( .INP(g7302), .ZN(n12861) );
  AND2X1 U12659 ( .IN1(n608), .IN2(n12862), .Q(n12859) );
  AND2X1 U12660 ( .IN1(g2574), .IN2(n7930), .Q(n12856) );
  OR2X1 U12661 ( .IN1(n12863), .IN2(n12864), .Q(g30061) );
  AND2X1 U12662 ( .IN1(n9672), .IN2(n12865), .Q(n12864) );
  OR2X1 U12663 ( .IN1(n12866), .IN2(n12867), .Q(n12865) );
  AND2X1 U12664 ( .IN1(n631), .IN2(g7390), .Q(n12867) );
  INVX0 U12665 ( .INP(n12868), .ZN(n631) );
  OR2X1 U12666 ( .IN1(n12869), .IN2(n12870), .Q(n12868) );
  AND2X1 U12667 ( .IN1(n4493), .IN2(n12871), .Q(n12870) );
  OR2X1 U12668 ( .IN1(n12872), .IN2(n12873), .Q(n12871) );
  AND2X1 U12669 ( .IN1(n10602), .IN2(g7194), .Q(n12873) );
  OR2X1 U12670 ( .IN1(n12874), .IN2(n12875), .Q(n10602) );
  AND2X1 U12671 ( .IN1(n4454), .IN2(n12876), .Q(n12875) );
  OR2X1 U12672 ( .IN1(n12877), .IN2(n12878), .Q(n12876) );
  AND2X1 U12673 ( .IN1(n12879), .IN2(g6944), .Q(n12878) );
  INVX0 U12674 ( .INP(n633), .ZN(n12879) );
  OR2X1 U12675 ( .IN1(n12880), .IN2(n12881), .Q(n633) );
  AND2X1 U12676 ( .IN1(n4570), .IN2(n12882), .Q(n12881) );
  OR2X1 U12677 ( .IN1(g6642), .IN2(g16297), .Q(n12882) );
  AND2X1 U12678 ( .IN1(g506), .IN2(n4571), .Q(n12880) );
  AND2X1 U12679 ( .IN1(n4316), .IN2(DFF_792_n1), .Q(n12877) );
  AND2X1 U12680 ( .IN1(g1192), .IN2(DFF_783_n1), .Q(n12874) );
  AND2X1 U12681 ( .IN1(n4315), .IN2(DFF_1142_n1), .Q(n12872) );
  AND2X1 U12682 ( .IN1(g1886), .IN2(DFF_1133_n1), .Q(n12869) );
  AND2X1 U12683 ( .IN1(n4370), .IN2(g16437), .Q(n12866) );
  AND2X1 U12684 ( .IN1(g2580), .IN2(n7926), .Q(n12863) );
  OR2X1 U12685 ( .IN1(n12883), .IN2(n12884), .Q(g30055) );
  AND2X1 U12686 ( .IN1(n12885), .IN2(g2374), .Q(n12884) );
  OR2X1 U12687 ( .IN1(n12886), .IN2(n12887), .Q(n12885) );
  AND2X1 U12688 ( .IN1(n4524), .IN2(g2380), .Q(n12887) );
  AND2X1 U12689 ( .IN1(g7264), .IN2(n532), .Q(n12886) );
  OR2X1 U12690 ( .IN1(n12888), .IN2(n12889), .Q(n532) );
  AND2X1 U12691 ( .IN1(n12890), .IN2(g1680), .Q(n12889) );
  OR2X1 U12692 ( .IN1(n12891), .IN2(n12892), .Q(n12890) );
  AND2X1 U12693 ( .IN1(n4525), .IN2(g1686), .Q(n12892) );
  AND2X1 U12694 ( .IN1(g7014), .IN2(n534), .Q(n12891) );
  INVX0 U12695 ( .INP(n12893), .ZN(n534) );
  OR2X1 U12696 ( .IN1(n12894), .IN2(n12895), .Q(n12893) );
  AND2X1 U12697 ( .IN1(n12896), .IN2(g986), .Q(n12895) );
  OR2X1 U12698 ( .IN1(n12897), .IN2(n12898), .Q(n12896) );
  AND2X1 U12699 ( .IN1(n12899), .IN2(g6712), .Q(n12898) );
  INVX0 U12700 ( .INP(g21346), .ZN(n12899) );
  AND2X1 U12701 ( .IN1(n4364), .IN2(n9894), .Q(n12897) );
  AND2X1 U12702 ( .IN1(n4432), .IN2(n8017), .Q(n12894) );
  AND2X1 U12703 ( .IN1(n18261), .IN2(n4488), .Q(n12888) );
  AND2X1 U12704 ( .IN1(n4487), .IN2(DFF_1378_n1), .Q(n12883) );
  OR2X1 U12705 ( .IN1(n12900), .IN2(n12901), .Q(g29941) );
  AND2X1 U12706 ( .IN1(n608), .IN2(g3109), .Q(n12901) );
  AND2X1 U12707 ( .IN1(n4494), .IN2(g3105), .Q(n12900) );
  OR2X1 U12708 ( .IN1(n12902), .IN2(n12903), .Q(g29939) );
  AND2X1 U12709 ( .IN1(n608), .IN2(g8030), .Q(n12903) );
  AND2X1 U12710 ( .IN1(n4383), .IN2(g3104), .Q(n12902) );
  OR2X1 U12711 ( .IN1(n12904), .IN2(n12905), .Q(g29936) );
  AND2X1 U12712 ( .IN1(n608), .IN2(g8106), .Q(n12905) );
  INVX0 U12713 ( .INP(n12906), .ZN(n608) );
  OR2X1 U12714 ( .IN1(n12907), .IN2(n12908), .Q(n12906) );
  AND2X1 U12715 ( .IN1(n12909), .IN2(n4545), .Q(n12908) );
  AND2X1 U12716 ( .IN1(n12910), .IN2(n12911), .Q(n12909) );
  OR2X1 U12717 ( .IN1(n4296), .IN2(n12912), .Q(n12911) );
  OR2X1 U12718 ( .IN1(g7052), .IN2(DFF_1100_n1), .Q(n12910) );
  AND2X1 U12719 ( .IN1(g1880), .IN2(DFF_1099_n1), .Q(n12907) );
  AND2X1 U12720 ( .IN1(n4382), .IN2(g3103), .Q(n12904) );
  OR2X1 U12721 ( .IN1(n12913), .IN2(n12914), .Q(g29623) );
  AND2X1 U12722 ( .IN1(n4509), .IN2(g2389), .Q(n12914) );
  AND2X1 U12723 ( .IN1(n12915), .IN2(n4606), .Q(n12913) );
  OR2X1 U12724 ( .IN1(n12916), .IN2(n12917), .Q(g29621) );
  AND2X1 U12725 ( .IN1(n4524), .IN2(g2388), .Q(n12917) );
  AND2X1 U12726 ( .IN1(n12915), .IN2(g7264), .Q(n12916) );
  OR2X1 U12727 ( .IN1(n12918), .IN2(n12919), .Q(g29620) );
  AND2X1 U12728 ( .IN1(n4511), .IN2(g1695), .Q(n12919) );
  AND2X1 U12729 ( .IN1(n12920), .IN2(n4618), .Q(n12918) );
  OR2X1 U12730 ( .IN1(n12921), .IN2(n12922), .Q(g29618) );
  AND2X1 U12731 ( .IN1(n4516), .IN2(g2387), .Q(n12922) );
  AND2X1 U12732 ( .IN1(n12915), .IN2(g5555), .Q(n12921) );
  AND2X1 U12733 ( .IN1(n12923), .IN2(n12221), .Q(n12915) );
  OR2X1 U12734 ( .IN1(n12924), .IN2(n12633), .Q(n12221) );
  INVX0 U12735 ( .INP(n12925), .ZN(n12924) );
  OR2X1 U12736 ( .IN1(n12926), .IN2(n4529), .Q(n12923) );
  INVX0 U12737 ( .INP(n11593), .ZN(n4529) );
  OR2X1 U12738 ( .IN1(n12241), .IN2(n12927), .Q(n11593) );
  OR2X1 U12739 ( .IN1(n12226), .IN2(n12245), .Q(n12927) );
  INVX0 U12740 ( .INP(n12227), .ZN(n12226) );
  AND2X1 U12741 ( .IN1(n12631), .IN2(n12928), .Q(n12926) );
  AND2X1 U12742 ( .IN1(n12630), .IN2(n12245), .Q(n12928) );
  OR2X1 U12743 ( .IN1(n12929), .IN2(n12930), .Q(g29617) );
  AND2X1 U12744 ( .IN1(n4525), .IN2(g1694), .Q(n12930) );
  AND2X1 U12745 ( .IN1(n12920), .IN2(g7014), .Q(n12929) );
  OR2X1 U12746 ( .IN1(n12931), .IN2(n12932), .Q(g29616) );
  AND2X1 U12747 ( .IN1(n12933), .IN2(g1088), .Q(n12932) );
  AND2X1 U12748 ( .IN1(n4381), .IN2(g1001), .Q(n12931) );
  OR2X1 U12749 ( .IN1(n12934), .IN2(n12935), .Q(g29613) );
  AND2X1 U12750 ( .IN1(n4518), .IN2(g1693), .Q(n12935) );
  AND2X1 U12751 ( .IN1(n12920), .IN2(g5511), .Q(n12934) );
  AND2X1 U12752 ( .IN1(n12936), .IN2(n11758), .Q(n12920) );
  OR2X1 U12753 ( .IN1(n12937), .IN2(n12695), .Q(n11758) );
  INVX0 U12754 ( .INP(n12938), .ZN(n12937) );
  OR2X1 U12755 ( .IN1(n12939), .IN2(n4530), .Q(n12936) );
  INVX0 U12756 ( .INP(n11590), .ZN(n4530) );
  OR2X1 U12757 ( .IN1(n11778), .IN2(n12940), .Q(n11590) );
  OR2X1 U12758 ( .IN1(n11763), .IN2(n11782), .Q(n12940) );
  INVX0 U12759 ( .INP(n11764), .ZN(n11763) );
  AND2X1 U12760 ( .IN1(n12693), .IN2(n12941), .Q(n12939) );
  AND2X1 U12761 ( .IN1(n12692), .IN2(n11782), .Q(n12941) );
  OR2X1 U12762 ( .IN1(n12942), .IN2(n12943), .Q(g29612) );
  AND2X1 U12763 ( .IN1(n12933), .IN2(g6712), .Q(n12943) );
  AND2X1 U12764 ( .IN1(n4364), .IN2(g1000), .Q(n12942) );
  OR2X1 U12765 ( .IN1(n12944), .IN2(n12945), .Q(g29611) );
  AND2X1 U12766 ( .IN1(n4506), .IN2(g314), .Q(n12945) );
  AND2X1 U12767 ( .IN1(n12946), .IN2(n4640), .Q(n12944) );
  OR2X1 U12768 ( .IN1(n12947), .IN2(n12948), .Q(g29609) );
  AND2X1 U12769 ( .IN1(n12933), .IN2(g5472), .Q(n12948) );
  AND2X1 U12770 ( .IN1(n12949), .IN2(n12749), .Q(n12933) );
  INVX0 U12771 ( .INP(n2617), .ZN(n12749) );
  AND2X1 U12772 ( .IN1(n12950), .IN2(n12951), .Q(n2617) );
  INVX0 U12773 ( .INP(n12756), .ZN(n12951) );
  OR2X1 U12774 ( .IN1(n12952), .IN2(n11981), .Q(n12949) );
  INVX0 U12775 ( .INP(n11982), .ZN(n11981) );
  OR2X1 U12776 ( .IN1(n11566), .IN2(n12953), .Q(n11982) );
  OR2X1 U12777 ( .IN1(n11581), .IN2(n11564), .Q(n12953) );
  INVX0 U12778 ( .INP(n11575), .ZN(n11581) );
  AND2X1 U12779 ( .IN1(n12754), .IN2(n12954), .Q(n12952) );
  AND2X1 U12780 ( .IN1(n12753), .IN2(n11564), .Q(n12954) );
  AND2X1 U12781 ( .IN1(n4363), .IN2(g999), .Q(n12947) );
  OR2X1 U12782 ( .IN1(n12955), .IN2(n12956), .Q(g29608) );
  AND2X1 U12783 ( .IN1(n4499), .IN2(g313), .Q(n12956) );
  AND2X1 U12784 ( .IN1(n12946), .IN2(g6447), .Q(n12955) );
  OR2X1 U12785 ( .IN1(n12957), .IN2(n12958), .Q(g29606) );
  AND2X1 U12786 ( .IN1(n4520), .IN2(g312), .Q(n12958) );
  AND2X1 U12787 ( .IN1(n12946), .IN2(g5437), .Q(n12957) );
  AND2X1 U12788 ( .IN1(n12959), .IN2(n11811), .Q(n12946) );
  OR2X1 U12789 ( .IN1(n12960), .IN2(n12813), .Q(n11811) );
  INVX0 U12790 ( .INP(n12961), .ZN(n12960) );
  OR2X1 U12791 ( .IN1(n12962), .IN2(n11586), .Q(n12959) );
  INVX0 U12792 ( .INP(n11587), .ZN(n11586) );
  OR2X1 U12793 ( .IN1(n11831), .IN2(n12963), .Q(n11587) );
  OR2X1 U12794 ( .IN1(n11816), .IN2(n11835), .Q(n12963) );
  INVX0 U12795 ( .INP(n11817), .ZN(n11816) );
  AND2X1 U12796 ( .IN1(n12811), .IN2(n12964), .Q(n12962) );
  AND2X1 U12797 ( .IN1(n12810), .IN2(n11835), .Q(n12964) );
  AND2X1 U12798 ( .IN1(n12965), .IN2(n12966), .Q(g29582) );
  OR2X1 U12799 ( .IN1(n12967), .IN2(n12968), .Q(n12965) );
  AND2X1 U12800 ( .IN1(n2981), .IN2(g2120), .Q(n12968) );
  AND2X1 U12801 ( .IN1(n9353), .IN2(n12969), .Q(n12967) );
  INVX0 U12802 ( .INP(n2981), .ZN(n12969) );
  AND2X1 U12803 ( .IN1(n12970), .IN2(n12971), .Q(g29581) );
  OR2X1 U12804 ( .IN1(n12972), .IN2(n12973), .Q(n12970) );
  AND2X1 U12805 ( .IN1(n2984), .IN2(g1426), .Q(n12973) );
  AND2X1 U12806 ( .IN1(n9354), .IN2(n12974), .Q(n12972) );
  INVX0 U12807 ( .INP(n2984), .ZN(n12974) );
  AND2X1 U12808 ( .IN1(n12975), .IN2(n12976), .Q(g29580) );
  OR2X1 U12809 ( .IN1(n12977), .IN2(n12978), .Q(n12975) );
  AND2X1 U12810 ( .IN1(n2987), .IN2(g740), .Q(n12978) );
  AND2X1 U12811 ( .IN1(n9355), .IN2(n12979), .Q(n12977) );
  INVX0 U12812 ( .INP(n2987), .ZN(n12979) );
  AND2X1 U12813 ( .IN1(n12980), .IN2(n12981), .Q(g29579) );
  OR2X1 U12814 ( .IN1(n12982), .IN2(n12983), .Q(n12980) );
  AND2X1 U12815 ( .IN1(n2990), .IN2(g52), .Q(n12983) );
  AND2X1 U12816 ( .IN1(n9356), .IN2(n12984), .Q(n12982) );
  INVX0 U12817 ( .INP(n2990), .ZN(n12984) );
  AND2X1 U12818 ( .IN1(n12985), .IN2(n12966), .Q(g29357) );
  AND2X1 U12819 ( .IN1(n12986), .IN2(n12987), .Q(n12985) );
  INVX0 U12820 ( .INP(n12988), .ZN(n12987) );
  AND2X1 U12821 ( .IN1(n1577), .IN2(n9507), .Q(n12988) );
  OR2X1 U12822 ( .IN1(n9507), .IN2(n1577), .Q(n12986) );
  AND2X1 U12823 ( .IN1(n12989), .IN2(n12971), .Q(g29355) );
  AND2X1 U12824 ( .IN1(n12990), .IN2(n12991), .Q(n12989) );
  INVX0 U12825 ( .INP(n12992), .ZN(n12991) );
  AND2X1 U12826 ( .IN1(n1233), .IN2(n9508), .Q(n12992) );
  OR2X1 U12827 ( .IN1(n9508), .IN2(n1233), .Q(n12990) );
  AND2X1 U12828 ( .IN1(n12993), .IN2(n12976), .Q(g29354) );
  AND2X1 U12829 ( .IN1(n12994), .IN2(n12995), .Q(n12993) );
  INVX0 U12830 ( .INP(n12996), .ZN(n12995) );
  AND2X1 U12831 ( .IN1(n888), .IN2(n9509), .Q(n12996) );
  OR2X1 U12832 ( .IN1(n9509), .IN2(n888), .Q(n12994) );
  OR2X1 U12833 ( .IN1(n12997), .IN2(n10195), .Q(n888) );
  AND2X1 U12834 ( .IN1(n12998), .IN2(n12981), .Q(g29353) );
  AND2X1 U12835 ( .IN1(n12999), .IN2(n13000), .Q(n12998) );
  INVX0 U12836 ( .INP(n13001), .ZN(n13000) );
  AND2X1 U12837 ( .IN1(n470), .IN2(n9510), .Q(n13001) );
  OR2X1 U12838 ( .IN1(n9510), .IN2(n470), .Q(n12999) );
  OR2X1 U12839 ( .IN1(n13002), .IN2(n13003), .Q(g29226) );
  AND2X1 U12840 ( .IN1(n4509), .IN2(g2498), .Q(n13003) );
  AND2X1 U12841 ( .IN1(n13004), .IN2(n4606), .Q(n13002) );
  OR2X1 U12842 ( .IN1(n13005), .IN2(n13006), .Q(g29221) );
  AND2X1 U12843 ( .IN1(n4524), .IN2(g2495), .Q(n13006) );
  AND2X1 U12844 ( .IN1(n13004), .IN2(g7264), .Q(n13005) );
  OR2X1 U12845 ( .IN1(n13007), .IN2(n13008), .Q(g29218) );
  AND2X1 U12846 ( .IN1(n4511), .IN2(g1804), .Q(n13008) );
  AND2X1 U12847 ( .IN1(n13009), .IN2(n4618), .Q(n13007) );
  OR2X1 U12848 ( .IN1(n13010), .IN2(n13011), .Q(g29213) );
  AND2X1 U12849 ( .IN1(n4516), .IN2(g2492), .Q(n13011) );
  AND2X1 U12850 ( .IN1(n13004), .IN2(g5555), .Q(n13010) );
  AND2X1 U12851 ( .IN1(n13012), .IN2(n13013), .Q(n13004) );
  OR2X1 U12852 ( .IN1(n13014), .IN2(n4285), .Q(n13013) );
  INVX0 U12853 ( .INP(n13015), .ZN(n13014) );
  OR2X1 U12854 ( .IN1(n13015), .IN2(n13016), .Q(n13012) );
  OR2X1 U12855 ( .IN1(n10191), .IN2(n13017), .Q(n13015) );
  OR2X1 U12856 ( .IN1(n13018), .IN2(n13019), .Q(n13017) );
  AND2X1 U12857 ( .IN1(n13020), .IN2(n13016), .Q(n13019) );
  OR2X1 U12858 ( .IN1(n13021), .IN2(n13022), .Q(n13020) );
  AND2X1 U12859 ( .IN1(n12235), .IN2(n13023), .Q(n13021) );
  OR2X1 U12860 ( .IN1(n13024), .IN2(n13025), .Q(n13023) );
  AND2X1 U12861 ( .IN1(n13026), .IN2(n4285), .Q(n13018) );
  OR2X1 U12862 ( .IN1(n13025), .IN2(n13027), .Q(n13026) );
  OR2X1 U12863 ( .IN1(n13024), .IN2(n13028), .Q(n13027) );
  OR2X1 U12864 ( .IN1(n13029), .IN2(n13030), .Q(g29212) );
  AND2X1 U12865 ( .IN1(n4525), .IN2(g1801), .Q(n13030) );
  AND2X1 U12866 ( .IN1(n13009), .IN2(g7014), .Q(n13029) );
  OR2X1 U12867 ( .IN1(n13031), .IN2(n13032), .Q(g29209) );
  AND2X1 U12868 ( .IN1(n13033), .IN2(g1088), .Q(n13032) );
  AND2X1 U12869 ( .IN1(n4381), .IN2(g1110), .Q(n13031) );
  OR2X1 U12870 ( .IN1(n13034), .IN2(n13035), .Q(g29205) );
  AND2X1 U12871 ( .IN1(n4518), .IN2(g1798), .Q(n13035) );
  AND2X1 U12872 ( .IN1(n13009), .IN2(g5511), .Q(n13034) );
  AND2X1 U12873 ( .IN1(n13036), .IN2(n13037), .Q(n13009) );
  OR2X1 U12874 ( .IN1(n13038), .IN2(n4284), .Q(n13037) );
  INVX0 U12875 ( .INP(n13039), .ZN(n13038) );
  OR2X1 U12876 ( .IN1(n13039), .IN2(n13040), .Q(n13036) );
  OR2X1 U12877 ( .IN1(n4386), .IN2(n13041), .Q(n13039) );
  OR2X1 U12878 ( .IN1(n13042), .IN2(n13043), .Q(n13041) );
  AND2X1 U12879 ( .IN1(n13044), .IN2(n13040), .Q(n13043) );
  OR2X1 U12880 ( .IN1(n13045), .IN2(n13046), .Q(n13044) );
  AND2X1 U12881 ( .IN1(n11772), .IN2(n13047), .Q(n13045) );
  OR2X1 U12882 ( .IN1(n13048), .IN2(n13049), .Q(n13047) );
  AND2X1 U12883 ( .IN1(n13050), .IN2(n4284), .Q(n13042) );
  OR2X1 U12884 ( .IN1(n13049), .IN2(n13051), .Q(n13050) );
  OR2X1 U12885 ( .IN1(n13048), .IN2(n13052), .Q(n13051) );
  OR2X1 U12886 ( .IN1(n13053), .IN2(n13054), .Q(g29204) );
  AND2X1 U12887 ( .IN1(n13033), .IN2(g6712), .Q(n13054) );
  AND2X1 U12888 ( .IN1(n4364), .IN2(g1107), .Q(n13053) );
  OR2X1 U12889 ( .IN1(n13055), .IN2(n13056), .Q(g29201) );
  AND2X1 U12890 ( .IN1(n4506), .IN2(g423), .Q(n13056) );
  AND2X1 U12891 ( .IN1(n13057), .IN2(n4640), .Q(n13055) );
  OR2X1 U12892 ( .IN1(n13058), .IN2(n13059), .Q(g29198) );
  AND2X1 U12893 ( .IN1(n13033), .IN2(g5472), .Q(n13059) );
  AND2X1 U12894 ( .IN1(n13060), .IN2(n13061), .Q(n13033) );
  OR2X1 U12895 ( .IN1(n13062), .IN2(n4283), .Q(n13061) );
  INVX0 U12896 ( .INP(n13063), .ZN(n13062) );
  OR2X1 U12897 ( .IN1(n13063), .IN2(n13064), .Q(n13060) );
  OR2X1 U12898 ( .IN1(n4387), .IN2(n13065), .Q(n13063) );
  OR2X1 U12899 ( .IN1(n13066), .IN2(n13067), .Q(n13065) );
  AND2X1 U12900 ( .IN1(n13068), .IN2(n13064), .Q(n13067) );
  OR2X1 U12901 ( .IN1(n13069), .IN2(n13070), .Q(n13068) );
  AND2X1 U12902 ( .IN1(n11577), .IN2(n13071), .Q(n13069) );
  OR2X1 U12903 ( .IN1(n13072), .IN2(n13073), .Q(n13071) );
  AND2X1 U12904 ( .IN1(n13074), .IN2(n4283), .Q(n13066) );
  OR2X1 U12905 ( .IN1(n13073), .IN2(n13075), .Q(n13074) );
  OR2X1 U12906 ( .IN1(n13072), .IN2(n13076), .Q(n13075) );
  AND2X1 U12907 ( .IN1(n4363), .IN2(g1104), .Q(n13058) );
  OR2X1 U12908 ( .IN1(n13077), .IN2(n13078), .Q(g29197) );
  AND2X1 U12909 ( .IN1(n4499), .IN2(g420), .Q(n13078) );
  AND2X1 U12910 ( .IN1(n13057), .IN2(g6447), .Q(n13077) );
  OR2X1 U12911 ( .IN1(n13079), .IN2(n13080), .Q(g29194) );
  AND2X1 U12912 ( .IN1(n4520), .IN2(g417), .Q(n13080) );
  AND2X1 U12913 ( .IN1(n13057), .IN2(g5437), .Q(n13079) );
  AND2X1 U12914 ( .IN1(n13081), .IN2(n13082), .Q(n13057) );
  OR2X1 U12915 ( .IN1(n13083), .IN2(n4282), .Q(n13082) );
  INVX0 U12916 ( .INP(n13084), .ZN(n13083) );
  OR2X1 U12917 ( .IN1(n13084), .IN2(n13085), .Q(n13081) );
  OR2X1 U12918 ( .IN1(n4388), .IN2(n13086), .Q(n13084) );
  OR2X1 U12919 ( .IN1(n13087), .IN2(n13088), .Q(n13086) );
  AND2X1 U12920 ( .IN1(n13089), .IN2(n13085), .Q(n13088) );
  OR2X1 U12921 ( .IN1(n13090), .IN2(n13091), .Q(n13089) );
  AND2X1 U12922 ( .IN1(n11825), .IN2(n13092), .Q(n13090) );
  OR2X1 U12923 ( .IN1(n13093), .IN2(n13094), .Q(n13092) );
  AND2X1 U12924 ( .IN1(n13095), .IN2(n4282), .Q(n13087) );
  OR2X1 U12925 ( .IN1(n13094), .IN2(n13096), .Q(n13095) );
  OR2X1 U12926 ( .IN1(n13093), .IN2(n13097), .Q(n13096) );
  OR2X1 U12927 ( .IN1(n13098), .IN2(n13099), .Q(g29187) );
  AND2X1 U12928 ( .IN1(n13100), .IN2(n13101), .Q(n13099) );
  AND2X1 U12929 ( .IN1(n13102), .IN2(g2396), .Q(n13098) );
  OR2X1 U12930 ( .IN1(n4509), .IN2(n13103), .Q(n13102) );
  OR2X1 U12931 ( .IN1(n13104), .IN2(n13105), .Q(g29185) );
  AND2X1 U12932 ( .IN1(n13100), .IN2(n13106), .Q(n13105) );
  AND2X1 U12933 ( .IN1(n13107), .IN2(g2398), .Q(n13104) );
  OR2X1 U12934 ( .IN1(n4524), .IN2(n13103), .Q(n13107) );
  OR2X1 U12935 ( .IN1(n13108), .IN2(n13109), .Q(g29184) );
  AND2X1 U12936 ( .IN1(n13110), .IN2(n13111), .Q(n13109) );
  AND2X1 U12937 ( .IN1(n13112), .IN2(g1702), .Q(n13108) );
  OR2X1 U12938 ( .IN1(n4511), .IN2(n13113), .Q(n13112) );
  OR2X1 U12939 ( .IN1(n13114), .IN2(n13115), .Q(g29182) );
  AND2X1 U12940 ( .IN1(n13100), .IN2(n13116), .Q(n13115) );
  AND2X1 U12941 ( .IN1(n13103), .IN2(n13117), .Q(n13100) );
  INVX0 U12942 ( .INP(n13118), .ZN(n13117) );
  OR2X1 U12943 ( .IN1(n13119), .IN2(n13120), .Q(n13118) );
  AND2X1 U12944 ( .IN1(n12314), .IN2(n12631), .Q(n13120) );
  AND2X1 U12945 ( .IN1(n13121), .IN2(g2397), .Q(n13114) );
  OR2X1 U12946 ( .IN1(n4516), .IN2(n13103), .Q(n13121) );
  OR2X1 U12947 ( .IN1(n12633), .IN2(n13122), .Q(n13103) );
  OR2X1 U12948 ( .IN1(n13119), .IN2(n13123), .Q(n13122) );
  AND2X1 U12949 ( .IN1(n13124), .IN2(n12631), .Q(n13123) );
  OR2X1 U12950 ( .IN1(n12314), .IN2(n13125), .Q(n13124) );
  OR2X1 U12951 ( .IN1(n12261), .IN2(n12321), .Q(n13125) );
  OR2X1 U12952 ( .IN1(n12241), .IN2(n12630), .Q(n12321) );
  OR2X1 U12953 ( .IN1(n12259), .IN2(n13126), .Q(n12630) );
  AND2X1 U12954 ( .IN1(n3038), .IN2(n13127), .Q(n13126) );
  OR2X1 U12955 ( .IN1(n12257), .IN2(n12254), .Q(n13127) );
  OR2X1 U12956 ( .IN1(n13128), .IN2(n13129), .Q(n12254) );
  AND2X1 U12957 ( .IN1(n13130), .IN2(n13131), .Q(n13129) );
  AND2X1 U12958 ( .IN1(n13132), .IN2(n13133), .Q(n13130) );
  OR2X1 U12959 ( .IN1(n13134), .IN2(n13135), .Q(n13133) );
  OR2X1 U12960 ( .IN1(n13136), .IN2(n13137), .Q(n13132) );
  AND2X1 U12961 ( .IN1(n13138), .IN2(n13135), .Q(n13128) );
  AND2X1 U12962 ( .IN1(n13139), .IN2(n13140), .Q(n13138) );
  OR2X1 U12963 ( .IN1(n13131), .IN2(n13137), .Q(n13140) );
  AND2X1 U12964 ( .IN1(n13136), .IN2(n13141), .Q(n12257) );
  AND2X1 U12965 ( .IN1(n13142), .IN2(n13143), .Q(n13141) );
  OR2X1 U12966 ( .IN1(n13131), .IN2(n13134), .Q(n13142) );
  INVX0 U12967 ( .INP(n12244), .ZN(n12259) );
  OR2X1 U12968 ( .IN1(n13144), .IN2(n12248), .Q(n12244) );
  AND2X1 U12969 ( .IN1(n13145), .IN2(n13146), .Q(n13144) );
  OR2X1 U12970 ( .IN1(n13147), .IN2(n13148), .Q(n13146) );
  OR2X1 U12971 ( .IN1(n13149), .IN2(n13150), .Q(n13148) );
  AND2X1 U12972 ( .IN1(n13151), .IN2(n13152), .Q(n13150) );
  AND2X1 U12973 ( .IN1(n13153), .IN2(n13154), .Q(n13149) );
  AND2X1 U12974 ( .IN1(n13155), .IN2(n13156), .Q(n13145) );
  OR2X1 U12975 ( .IN1(n13153), .IN2(n13157), .Q(n13156) );
  OR2X1 U12976 ( .IN1(n13158), .IN2(n13159), .Q(n13157) );
  AND2X1 U12977 ( .IN1(n13147), .IN2(n13151), .Q(n13159) );
  AND2X1 U12978 ( .IN1(n13154), .IN2(n13152), .Q(n13158) );
  OR2X1 U12979 ( .IN1(n13152), .IN2(n13160), .Q(n13155) );
  OR2X1 U12980 ( .IN1(n13161), .IN2(n13162), .Q(n13160) );
  AND2X1 U12981 ( .IN1(n13153), .IN2(n13151), .Q(n13162) );
  INVX0 U12982 ( .INP(n13163), .ZN(n13151) );
  INVX0 U12983 ( .INP(n13164), .ZN(n13153) );
  AND2X1 U12984 ( .IN1(n13147), .IN2(n13154), .Q(n13161) );
  INVX0 U12985 ( .INP(n13165), .ZN(n13154) );
  INVX0 U12986 ( .INP(n13166), .ZN(n13147) );
  INVX0 U12987 ( .INP(n13167), .ZN(n13152) );
  OR2X1 U12988 ( .IN1(n12260), .IN2(n12248), .Q(n12314) );
  INVX0 U12989 ( .INP(n12249), .ZN(n12260) );
  OR2X1 U12990 ( .IN1(n13168), .IN2(n13169), .Q(n12249) );
  OR2X1 U12991 ( .IN1(n13170), .IN2(n13143), .Q(n13169) );
  OR2X1 U12992 ( .IN1(n13135), .IN2(n13137), .Q(n13143) );
  OR2X1 U12993 ( .IN1(n13171), .IN2(n13172), .Q(n13137) );
  AND2X1 U12994 ( .IN1(n10858), .IN2(g2195), .Q(n13172) );
  INVX0 U12995 ( .INP(n10859), .ZN(n10858) );
  AND2X1 U12996 ( .IN1(n4563), .IN2(n10859), .Q(n13171) );
  OR2X1 U12997 ( .IN1(n13173), .IN2(n13174), .Q(n10859) );
  OR2X1 U12998 ( .IN1(n13175), .IN2(n13176), .Q(n13174) );
  AND2X1 U12999 ( .IN1(g2241), .IN2(g2294), .Q(n13176) );
  AND2X1 U13000 ( .IN1(g6837), .IN2(g2288), .Q(n13175) );
  AND2X1 U13001 ( .IN1(test_so73), .IN2(g2291), .Q(n13173) );
  OR2X1 U13002 ( .IN1(n13177), .IN2(n13178), .Q(n13135) );
  AND2X1 U13003 ( .IN1(n13179), .IN2(n10837), .Q(n13178) );
  AND2X1 U13004 ( .IN1(n10836), .IN2(n12083), .Q(n13177) );
  INVX0 U13005 ( .INP(n10837), .ZN(n10836) );
  OR2X1 U13006 ( .IN1(n13180), .IN2(n13181), .Q(n10837) );
  OR2X1 U13007 ( .IN1(n13182), .IN2(n13183), .Q(n13181) );
  AND2X1 U13008 ( .IN1(g2241), .IN2(g2303), .Q(n13183) );
  AND2X1 U13009 ( .IN1(g6837), .IN2(g2297), .Q(n13182) );
  AND2X1 U13010 ( .IN1(test_so73), .IN2(g2300), .Q(n13180) );
  OR2X1 U13011 ( .IN1(n13131), .IN2(n13139), .Q(n13170) );
  OR2X1 U13012 ( .IN1(n13134), .IN2(n13136), .Q(n13139) );
  OR2X1 U13013 ( .IN1(n13184), .IN2(n13185), .Q(n13136) );
  AND2X1 U13014 ( .IN1(n10844), .IN2(g2165), .Q(n13185) );
  INVX0 U13015 ( .INP(n10845), .ZN(n10844) );
  AND2X1 U13016 ( .IN1(n4377), .IN2(n10845), .Q(n13184) );
  OR2X1 U13017 ( .IN1(n13186), .IN2(n13187), .Q(n10845) );
  OR2X1 U13018 ( .IN1(n13188), .IN2(n13189), .Q(n13187) );
  AND2X1 U13019 ( .IN1(g2261), .IN2(g6837), .Q(n13189) );
  AND2X1 U13020 ( .IN1(g2267), .IN2(g2241), .Q(n13188) );
  AND2X1 U13021 ( .IN1(test_so76), .IN2(test_so73), .Q(n13186) );
  OR2X1 U13022 ( .IN1(n13190), .IN2(n13191), .Q(n13134) );
  AND2X1 U13023 ( .IN1(n10862), .IN2(g2175), .Q(n13191) );
  INVX0 U13024 ( .INP(n10863), .ZN(n10862) );
  AND2X1 U13025 ( .IN1(n4319), .IN2(n10863), .Q(n13190) );
  OR2X1 U13026 ( .IN1(n13192), .IN2(n13193), .Q(n10863) );
  OR2X1 U13027 ( .IN1(n13194), .IN2(n13195), .Q(n13193) );
  AND2X1 U13028 ( .IN1(g2241), .IN2(g2276), .Q(n13195) );
  AND2X1 U13029 ( .IN1(g6837), .IN2(g2270), .Q(n13194) );
  AND2X1 U13030 ( .IN1(test_so73), .IN2(g2273), .Q(n13192) );
  OR2X1 U13031 ( .IN1(n13196), .IN2(n13197), .Q(n13131) );
  AND2X1 U13032 ( .IN1(n10854), .IN2(g2185), .Q(n13197) );
  INVX0 U13033 ( .INP(n10855), .ZN(n10854) );
  AND2X1 U13034 ( .IN1(n4325), .IN2(n10855), .Q(n13196) );
  OR2X1 U13035 ( .IN1(n13198), .IN2(n13199), .Q(n10855) );
  OR2X1 U13036 ( .IN1(n13200), .IN2(n13201), .Q(n13199) );
  AND2X1 U13037 ( .IN1(g2241), .IN2(g2285), .Q(n13201) );
  AND2X1 U13038 ( .IN1(g6837), .IN2(g2279), .Q(n13200) );
  AND2X1 U13039 ( .IN1(test_so73), .IN2(g2282), .Q(n13198) );
  OR2X1 U13040 ( .IN1(n13202), .IN2(n13203), .Q(n13168) );
  OR2X1 U13041 ( .IN1(n13166), .IN2(n13164), .Q(n13203) );
  OR2X1 U13042 ( .IN1(n13204), .IN2(n13205), .Q(n13164) );
  AND2X1 U13043 ( .IN1(n11898), .IN2(n10821), .Q(n13205) );
  AND2X1 U13044 ( .IN1(n10820), .IN2(n13206), .Q(n13204) );
  INVX0 U13045 ( .INP(n10821), .ZN(n10820) );
  OR2X1 U13046 ( .IN1(n13207), .IN2(n13208), .Q(n10821) );
  OR2X1 U13047 ( .IN1(n13209), .IN2(n13210), .Q(n13208) );
  AND2X1 U13048 ( .IN1(g2241), .IN2(g2348), .Q(n13210) );
  AND2X1 U13049 ( .IN1(g6837), .IN2(g2342), .Q(n13209) );
  AND2X1 U13050 ( .IN1(test_so73), .IN2(g2345), .Q(n13207) );
  OR2X1 U13051 ( .IN1(n13211), .IN2(n13212), .Q(n13166) );
  AND2X1 U13052 ( .IN1(n10824), .IN2(g2190), .Q(n13212) );
  INVX0 U13053 ( .INP(n10825), .ZN(n10824) );
  AND2X1 U13054 ( .IN1(n4555), .IN2(n10825), .Q(n13211) );
  OR2X1 U13055 ( .IN1(n13213), .IN2(n13214), .Q(n10825) );
  OR2X1 U13056 ( .IN1(n13215), .IN2(n13216), .Q(n13214) );
  AND2X1 U13057 ( .IN1(g2241), .IN2(g2330), .Q(n13216) );
  AND2X1 U13058 ( .IN1(g6837), .IN2(g2324), .Q(n13215) );
  AND2X1 U13059 ( .IN1(test_so77), .IN2(test_so73), .Q(n13213) );
  OR2X1 U13060 ( .IN1(n13163), .IN2(n13217), .Q(n13202) );
  OR2X1 U13061 ( .IN1(n13167), .IN2(n13165), .Q(n13217) );
  OR2X1 U13062 ( .IN1(n13218), .IN2(n13219), .Q(n13165) );
  AND2X1 U13063 ( .IN1(n10840), .IN2(g2180), .Q(n13219) );
  INVX0 U13064 ( .INP(n10841), .ZN(n10840) );
  AND2X1 U13065 ( .IN1(n4389), .IN2(n10841), .Q(n13218) );
  OR2X1 U13066 ( .IN1(n13220), .IN2(n13221), .Q(n10841) );
  OR2X1 U13067 ( .IN1(n13222), .IN2(n13223), .Q(n13221) );
  AND2X1 U13068 ( .IN1(g2241), .IN2(g2321), .Q(n13223) );
  AND2X1 U13069 ( .IN1(g6837), .IN2(g2315), .Q(n13222) );
  AND2X1 U13070 ( .IN1(test_so73), .IN2(g2318), .Q(n13220) );
  OR2X1 U13071 ( .IN1(n13224), .IN2(n13225), .Q(n13167) );
  AND2X1 U13072 ( .IN1(n12048), .IN2(g2170), .Q(n13225) );
  INVX0 U13073 ( .INP(n10870), .ZN(n12048) );
  AND2X1 U13074 ( .IN1(n4373), .IN2(n10870), .Q(n13224) );
  OR2X1 U13075 ( .IN1(n13226), .IN2(n13227), .Q(n10870) );
  OR2X1 U13076 ( .IN1(n13228), .IN2(n13229), .Q(n13227) );
  AND2X1 U13077 ( .IN1(g2241), .IN2(g2312), .Q(n13229) );
  AND2X1 U13078 ( .IN1(g6837), .IN2(g2306), .Q(n13228) );
  AND2X1 U13079 ( .IN1(test_so73), .IN2(g2309), .Q(n13226) );
  OR2X1 U13080 ( .IN1(n13230), .IN2(n13231), .Q(n13163) );
  AND2X1 U13081 ( .IN1(n10828), .IN2(g2200), .Q(n13231) );
  INVX0 U13082 ( .INP(n10829), .ZN(n10828) );
  AND2X1 U13083 ( .IN1(n4287), .IN2(n10829), .Q(n13230) );
  OR2X1 U13084 ( .IN1(n13232), .IN2(n13233), .Q(n10829) );
  OR2X1 U13085 ( .IN1(n13234), .IN2(n13235), .Q(n13233) );
  AND2X1 U13086 ( .IN1(g2241), .IN2(g2339), .Q(n13235) );
  AND2X1 U13087 ( .IN1(g6837), .IN2(g2333), .Q(n13234) );
  AND2X1 U13088 ( .IN1(test_so73), .IN2(g2336), .Q(n13232) );
  AND2X1 U13089 ( .IN1(n13236), .IN2(n10191), .Q(n13119) );
  OR2X1 U13090 ( .IN1(n13237), .IN2(n13238), .Q(g29181) );
  AND2X1 U13091 ( .IN1(n13110), .IN2(n13239), .Q(n13238) );
  AND2X1 U13092 ( .IN1(n13240), .IN2(g1704), .Q(n13237) );
  OR2X1 U13093 ( .IN1(n4525), .IN2(n13113), .Q(n13240) );
  OR2X1 U13094 ( .IN1(n13241), .IN2(n13242), .Q(g29179) );
  AND2X1 U13095 ( .IN1(n13243), .IN2(g1088), .Q(n13242) );
  AND2X1 U13096 ( .IN1(n13244), .IN2(g1008), .Q(n13241) );
  OR2X1 U13097 ( .IN1(n4381), .IN2(n13245), .Q(n13244) );
  OR2X1 U13098 ( .IN1(n13246), .IN2(n13247), .Q(g29178) );
  AND2X1 U13099 ( .IN1(n13110), .IN2(n13248), .Q(n13247) );
  AND2X1 U13100 ( .IN1(n13113), .IN2(n13249), .Q(n13110) );
  INVX0 U13101 ( .INP(n13250), .ZN(n13249) );
  OR2X1 U13102 ( .IN1(n13251), .IN2(n13252), .Q(n13250) );
  AND2X1 U13103 ( .IN1(n12333), .IN2(n12693), .Q(n13252) );
  AND2X1 U13104 ( .IN1(n13253), .IN2(g1703), .Q(n13246) );
  OR2X1 U13105 ( .IN1(n4518), .IN2(n13113), .Q(n13253) );
  OR2X1 U13106 ( .IN1(n12695), .IN2(n13254), .Q(n13113) );
  OR2X1 U13107 ( .IN1(n13251), .IN2(n13255), .Q(n13254) );
  AND2X1 U13108 ( .IN1(n13256), .IN2(n12693), .Q(n13255) );
  OR2X1 U13109 ( .IN1(n12333), .IN2(n13257), .Q(n13256) );
  OR2X1 U13110 ( .IN1(n11798), .IN2(n12340), .Q(n13257) );
  OR2X1 U13111 ( .IN1(n11778), .IN2(n12692), .Q(n12340) );
  OR2X1 U13112 ( .IN1(n11796), .IN2(n13258), .Q(n12692) );
  AND2X1 U13113 ( .IN1(n3070), .IN2(n13259), .Q(n13258) );
  OR2X1 U13114 ( .IN1(n11794), .IN2(n11791), .Q(n13259) );
  OR2X1 U13115 ( .IN1(n13260), .IN2(n13261), .Q(n11791) );
  AND2X1 U13116 ( .IN1(n13262), .IN2(n13263), .Q(n13261) );
  AND2X1 U13117 ( .IN1(n13264), .IN2(n13265), .Q(n13262) );
  OR2X1 U13118 ( .IN1(n13266), .IN2(n13267), .Q(n13265) );
  OR2X1 U13119 ( .IN1(n13268), .IN2(n13269), .Q(n13264) );
  AND2X1 U13120 ( .IN1(n13270), .IN2(n13267), .Q(n13260) );
  AND2X1 U13121 ( .IN1(n13271), .IN2(n13272), .Q(n13270) );
  OR2X1 U13122 ( .IN1(n13263), .IN2(n13269), .Q(n13272) );
  AND2X1 U13123 ( .IN1(n13268), .IN2(n13273), .Q(n11794) );
  AND2X1 U13124 ( .IN1(n13274), .IN2(n13275), .Q(n13273) );
  OR2X1 U13125 ( .IN1(n13263), .IN2(n13266), .Q(n13274) );
  INVX0 U13126 ( .INP(n11781), .ZN(n11796) );
  OR2X1 U13127 ( .IN1(n13276), .IN2(n11785), .Q(n11781) );
  AND2X1 U13128 ( .IN1(n13277), .IN2(n13278), .Q(n13276) );
  OR2X1 U13129 ( .IN1(n13279), .IN2(n13280), .Q(n13278) );
  OR2X1 U13130 ( .IN1(n13281), .IN2(n13282), .Q(n13280) );
  AND2X1 U13131 ( .IN1(n13283), .IN2(n13284), .Q(n13282) );
  AND2X1 U13132 ( .IN1(n13285), .IN2(n13286), .Q(n13281) );
  AND2X1 U13133 ( .IN1(n13287), .IN2(n13288), .Q(n13277) );
  OR2X1 U13134 ( .IN1(n13285), .IN2(n13289), .Q(n13288) );
  OR2X1 U13135 ( .IN1(n13290), .IN2(n13291), .Q(n13289) );
  AND2X1 U13136 ( .IN1(n13279), .IN2(n13283), .Q(n13291) );
  AND2X1 U13137 ( .IN1(n13286), .IN2(n13284), .Q(n13290) );
  OR2X1 U13138 ( .IN1(n13284), .IN2(n13292), .Q(n13287) );
  OR2X1 U13139 ( .IN1(n13293), .IN2(n13294), .Q(n13292) );
  AND2X1 U13140 ( .IN1(n13285), .IN2(n13283), .Q(n13294) );
  INVX0 U13141 ( .INP(n13295), .ZN(n13283) );
  INVX0 U13142 ( .INP(n13296), .ZN(n13285) );
  AND2X1 U13143 ( .IN1(n13279), .IN2(n13286), .Q(n13293) );
  INVX0 U13144 ( .INP(n13297), .ZN(n13286) );
  INVX0 U13145 ( .INP(n13298), .ZN(n13279) );
  INVX0 U13146 ( .INP(n13299), .ZN(n13284) );
  OR2X1 U13147 ( .IN1(n11797), .IN2(n11785), .Q(n12333) );
  INVX0 U13148 ( .INP(n11786), .ZN(n11797) );
  OR2X1 U13149 ( .IN1(n13300), .IN2(n13301), .Q(n11786) );
  OR2X1 U13150 ( .IN1(n13302), .IN2(n13275), .Q(n13301) );
  OR2X1 U13151 ( .IN1(n13267), .IN2(n13269), .Q(n13275) );
  OR2X1 U13152 ( .IN1(n13303), .IN2(n13304), .Q(n13269) );
  AND2X1 U13153 ( .IN1(n10797), .IN2(g1501), .Q(n13304) );
  INVX0 U13154 ( .INP(n10798), .ZN(n10797) );
  AND2X1 U13155 ( .IN1(n4565), .IN2(n10798), .Q(n13303) );
  OR2X1 U13156 ( .IN1(n13305), .IN2(n13306), .Q(n10798) );
  OR2X1 U13157 ( .IN1(n13307), .IN2(n13308), .Q(n13306) );
  AND2X1 U13158 ( .IN1(g1547), .IN2(g1600), .Q(n13308) );
  AND2X1 U13159 ( .IN1(g6573), .IN2(g1594), .Q(n13307) );
  AND2X1 U13160 ( .IN1(g6782), .IN2(g1597), .Q(n13305) );
  OR2X1 U13161 ( .IN1(n13309), .IN2(n13310), .Q(n13267) );
  AND2X1 U13162 ( .IN1(n13311), .IN2(n10794), .Q(n13310) );
  AND2X1 U13163 ( .IN1(n10793), .IN2(n12135), .Q(n13309) );
  INVX0 U13164 ( .INP(n10794), .ZN(n10793) );
  OR2X1 U13165 ( .IN1(n13312), .IN2(n13313), .Q(n10794) );
  OR2X1 U13166 ( .IN1(n13314), .IN2(n13315), .Q(n13313) );
  AND2X1 U13167 ( .IN1(g1547), .IN2(g1609), .Q(n13315) );
  AND2X1 U13168 ( .IN1(g6573), .IN2(g1603), .Q(n13314) );
  AND2X1 U13169 ( .IN1(test_so56), .IN2(g6782), .Q(n13312) );
  OR2X1 U13170 ( .IN1(n13263), .IN2(n13271), .Q(n13302) );
  OR2X1 U13171 ( .IN1(n13266), .IN2(n13268), .Q(n13271) );
  OR2X1 U13172 ( .IN1(n13316), .IN2(n13317), .Q(n13268) );
  AND2X1 U13173 ( .IN1(n10771), .IN2(g1471), .Q(n13317) );
  INVX0 U13174 ( .INP(n10772), .ZN(n10771) );
  AND2X1 U13175 ( .IN1(n4378), .IN2(n10772), .Q(n13316) );
  OR2X1 U13176 ( .IN1(n13318), .IN2(n13319), .Q(n10772) );
  OR2X1 U13177 ( .IN1(n13320), .IN2(n13321), .Q(n13319) );
  AND2X1 U13178 ( .IN1(g1570), .IN2(g6782), .Q(n13321) );
  AND2X1 U13179 ( .IN1(g1573), .IN2(g1547), .Q(n13320) );
  AND2X1 U13180 ( .IN1(g1567), .IN2(g6573), .Q(n13318) );
  OR2X1 U13181 ( .IN1(n13322), .IN2(n13323), .Q(n13266) );
  AND2X1 U13182 ( .IN1(n10789), .IN2(g1481), .Q(n13323) );
  INVX0 U13183 ( .INP(n10790), .ZN(n10789) );
  AND2X1 U13184 ( .IN1(n4320), .IN2(n10790), .Q(n13322) );
  OR2X1 U13185 ( .IN1(n13324), .IN2(n13325), .Q(n10790) );
  OR2X1 U13186 ( .IN1(n13326), .IN2(n13327), .Q(n13325) );
  AND2X1 U13187 ( .IN1(g1547), .IN2(g1582), .Q(n13327) );
  AND2X1 U13188 ( .IN1(g6573), .IN2(g1576), .Q(n13326) );
  AND2X1 U13189 ( .IN1(g6782), .IN2(g1579), .Q(n13324) );
  OR2X1 U13190 ( .IN1(n13328), .IN2(n13329), .Q(n13263) );
  AND2X1 U13191 ( .IN1(n10804), .IN2(g1491), .Q(n13329) );
  INVX0 U13192 ( .INP(n10805), .ZN(n10804) );
  AND2X1 U13193 ( .IN1(n4326), .IN2(n10805), .Q(n13328) );
  OR2X1 U13194 ( .IN1(n13330), .IN2(n13331), .Q(n10805) );
  OR2X1 U13195 ( .IN1(n13332), .IN2(n13333), .Q(n13331) );
  AND2X1 U13196 ( .IN1(g1547), .IN2(g1591), .Q(n13333) );
  AND2X1 U13197 ( .IN1(g6573), .IN2(g1585), .Q(n13332) );
  AND2X1 U13198 ( .IN1(g6782), .IN2(g1588), .Q(n13330) );
  OR2X1 U13199 ( .IN1(n13334), .IN2(n13335), .Q(n13300) );
  OR2X1 U13200 ( .IN1(n13298), .IN2(n13296), .Q(n13335) );
  OR2X1 U13201 ( .IN1(n13336), .IN2(n13337), .Q(n13296) );
  AND2X1 U13202 ( .IN1(n11936), .IN2(n10776), .Q(n13337) );
  AND2X1 U13203 ( .IN1(n10775), .IN2(n13338), .Q(n13336) );
  INVX0 U13204 ( .INP(n10776), .ZN(n10775) );
  OR2X1 U13205 ( .IN1(n13339), .IN2(n13340), .Q(n10776) );
  OR2X1 U13206 ( .IN1(n13341), .IN2(n13342), .Q(n13340) );
  AND2X1 U13207 ( .IN1(g1547), .IN2(g1654), .Q(n13342) );
  AND2X1 U13208 ( .IN1(g6573), .IN2(g1648), .Q(n13341) );
  AND2X1 U13209 ( .IN1(g6782), .IN2(g1651), .Q(n13339) );
  OR2X1 U13210 ( .IN1(n13343), .IN2(n13344), .Q(n13298) );
  AND2X1 U13211 ( .IN1(n10759), .IN2(g1496), .Q(n13344) );
  INVX0 U13212 ( .INP(n10760), .ZN(n10759) );
  AND2X1 U13213 ( .IN1(n4557), .IN2(n10760), .Q(n13343) );
  OR2X1 U13214 ( .IN1(n13345), .IN2(n13346), .Q(n10760) );
  OR2X1 U13215 ( .IN1(n13347), .IN2(n13348), .Q(n13346) );
  AND2X1 U13216 ( .IN1(g1547), .IN2(g1636), .Q(n13348) );
  AND2X1 U13217 ( .IN1(g6573), .IN2(g1630), .Q(n13347) );
  AND2X1 U13218 ( .IN1(g6782), .IN2(g1633), .Q(n13345) );
  OR2X1 U13219 ( .IN1(n13295), .IN2(n13349), .Q(n13334) );
  OR2X1 U13220 ( .IN1(n13299), .IN2(n13297), .Q(n13349) );
  OR2X1 U13221 ( .IN1(n13350), .IN2(n13351), .Q(n13297) );
  AND2X1 U13222 ( .IN1(n10779), .IN2(g1486), .Q(n13351) );
  INVX0 U13223 ( .INP(n10780), .ZN(n10779) );
  AND2X1 U13224 ( .IN1(n4390), .IN2(n10780), .Q(n13350) );
  OR2X1 U13225 ( .IN1(n13352), .IN2(n13353), .Q(n10780) );
  OR2X1 U13226 ( .IN1(n13354), .IN2(n13355), .Q(n13353) );
  AND2X1 U13227 ( .IN1(g1547), .IN2(g1627), .Q(n13355) );
  AND2X1 U13228 ( .IN1(test_so55), .IN2(g6573), .Q(n13354) );
  AND2X1 U13229 ( .IN1(g6782), .IN2(g1624), .Q(n13352) );
  OR2X1 U13230 ( .IN1(n13356), .IN2(n13357), .Q(n13299) );
  AND2X1 U13231 ( .IN1(n10755), .IN2(g1476), .Q(n13357) );
  INVX0 U13232 ( .INP(n10756), .ZN(n10755) );
  AND2X1 U13233 ( .IN1(n4374), .IN2(n10756), .Q(n13356) );
  OR2X1 U13234 ( .IN1(n13358), .IN2(n13359), .Q(n10756) );
  OR2X1 U13235 ( .IN1(n13360), .IN2(n13361), .Q(n13359) );
  AND2X1 U13236 ( .IN1(g1547), .IN2(g1618), .Q(n13361) );
  AND2X1 U13237 ( .IN1(g6573), .IN2(g1612), .Q(n13360) );
  AND2X1 U13238 ( .IN1(g6782), .IN2(g1615), .Q(n13358) );
  OR2X1 U13239 ( .IN1(n13362), .IN2(n13363), .Q(n13295) );
  AND2X1 U13240 ( .IN1(n10763), .IN2(g1506), .Q(n13363) );
  INVX0 U13241 ( .INP(n10764), .ZN(n10763) );
  AND2X1 U13242 ( .IN1(n4288), .IN2(n10764), .Q(n13362) );
  OR2X1 U13243 ( .IN1(n13364), .IN2(n13365), .Q(n10764) );
  OR2X1 U13244 ( .IN1(n13366), .IN2(n13367), .Q(n13365) );
  AND2X1 U13245 ( .IN1(g1547), .IN2(g1645), .Q(n13367) );
  AND2X1 U13246 ( .IN1(g6573), .IN2(g1639), .Q(n13366) );
  AND2X1 U13247 ( .IN1(g6782), .IN2(g1642), .Q(n13364) );
  AND2X1 U13248 ( .IN1(n4386), .IN2(n13368), .Q(n13251) );
  OR2X1 U13249 ( .IN1(n13369), .IN2(n13370), .Q(g29173) );
  AND2X1 U13250 ( .IN1(n13243), .IN2(g6712), .Q(n13370) );
  AND2X1 U13251 ( .IN1(n13371), .IN2(g1010), .Q(n13369) );
  OR2X1 U13252 ( .IN1(n4364), .IN2(n13245), .Q(n13371) );
  OR2X1 U13253 ( .IN1(n13372), .IN2(n13373), .Q(g29172) );
  AND2X1 U13254 ( .IN1(n13374), .IN2(n13375), .Q(n13373) );
  AND2X1 U13255 ( .IN1(n13376), .IN2(g321), .Q(n13372) );
  OR2X1 U13256 ( .IN1(n4506), .IN2(n13377), .Q(n13376) );
  OR2X1 U13257 ( .IN1(n13378), .IN2(n13379), .Q(g29170) );
  AND2X1 U13258 ( .IN1(n13243), .IN2(g5472), .Q(n13379) );
  AND2X1 U13259 ( .IN1(n13245), .IN2(n13380), .Q(n13243) );
  INVX0 U13260 ( .INP(n13381), .ZN(n13380) );
  OR2X1 U13261 ( .IN1(n13382), .IN2(n13383), .Q(n13381) );
  AND2X1 U13262 ( .IN1(n12754), .IN2(n11571), .Q(n13383) );
  AND2X1 U13263 ( .IN1(n13384), .IN2(g1009), .Q(n13378) );
  OR2X1 U13264 ( .IN1(n4363), .IN2(n13245), .Q(n13384) );
  OR2X1 U13265 ( .IN1(n12756), .IN2(n13385), .Q(n13245) );
  OR2X1 U13266 ( .IN1(n13382), .IN2(n13386), .Q(n13385) );
  AND2X1 U13267 ( .IN1(n13387), .IN2(n12754), .Q(n13386) );
  OR2X1 U13268 ( .IN1(n11571), .IN2(n13388), .Q(n13387) );
  OR2X1 U13269 ( .IN1(n11569), .IN2(n11583), .Q(n13388) );
  OR2X1 U13270 ( .IN1(n11566), .IN2(n12753), .Q(n11583) );
  OR2X1 U13271 ( .IN1(n11623), .IN2(n13389), .Q(n12753) );
  AND2X1 U13272 ( .IN1(n3102), .IN2(n13390), .Q(n13389) );
  OR2X1 U13273 ( .IN1(n11620), .IN2(n11617), .Q(n13390) );
  OR2X1 U13274 ( .IN1(n13391), .IN2(n13392), .Q(n11617) );
  AND2X1 U13275 ( .IN1(n13393), .IN2(n13394), .Q(n13392) );
  AND2X1 U13276 ( .IN1(n13395), .IN2(n13396), .Q(n13393) );
  OR2X1 U13277 ( .IN1(n13397), .IN2(n13398), .Q(n13396) );
  OR2X1 U13278 ( .IN1(n13399), .IN2(n13400), .Q(n13395) );
  AND2X1 U13279 ( .IN1(n13401), .IN2(n13398), .Q(n13391) );
  AND2X1 U13280 ( .IN1(n13402), .IN2(n13403), .Q(n13401) );
  OR2X1 U13281 ( .IN1(n13394), .IN2(n13400), .Q(n13403) );
  AND2X1 U13282 ( .IN1(n13399), .IN2(n13404), .Q(n11620) );
  AND2X1 U13283 ( .IN1(n13405), .IN2(n13406), .Q(n13404) );
  OR2X1 U13284 ( .IN1(n13394), .IN2(n13397), .Q(n13405) );
  INVX0 U13285 ( .INP(n11610), .ZN(n11623) );
  OR2X1 U13286 ( .IN1(n13407), .IN2(n11579), .Q(n11610) );
  AND2X1 U13287 ( .IN1(n13408), .IN2(n13409), .Q(n13407) );
  OR2X1 U13288 ( .IN1(n13410), .IN2(n13411), .Q(n13409) );
  OR2X1 U13289 ( .IN1(n13412), .IN2(n13413), .Q(n13411) );
  AND2X1 U13290 ( .IN1(n13414), .IN2(n13415), .Q(n13412) );
  AND2X1 U13291 ( .IN1(n13416), .IN2(n13417), .Q(n13408) );
  OR2X1 U13292 ( .IN1(n13414), .IN2(n13418), .Q(n13417) );
  OR2X1 U13293 ( .IN1(n13419), .IN2(n13420), .Q(n13418) );
  AND2X1 U13294 ( .IN1(n13410), .IN2(n13421), .Q(n13420) );
  AND2X1 U13295 ( .IN1(n13415), .IN2(n13422), .Q(n13419) );
  OR2X1 U13296 ( .IN1(n13422), .IN2(n13423), .Q(n13416) );
  OR2X1 U13297 ( .IN1(n13424), .IN2(n13425), .Q(n13423) );
  AND2X1 U13298 ( .IN1(n13410), .IN2(n13415), .Q(n13425) );
  INVX0 U13299 ( .INP(n13426), .ZN(n13410) );
  AND2X1 U13300 ( .IN1(n13414), .IN2(n13421), .Q(n13424) );
  INVX0 U13301 ( .INP(n13427), .ZN(n13414) );
  OR2X1 U13302 ( .IN1(n11622), .IN2(n11579), .Q(n11571) );
  INVX0 U13303 ( .INP(n11580), .ZN(n11622) );
  OR2X1 U13304 ( .IN1(n13428), .IN2(n13429), .Q(n11580) );
  OR2X1 U13305 ( .IN1(n13430), .IN2(n13431), .Q(n13429) );
  OR2X1 U13306 ( .IN1(n13427), .IN2(n13426), .Q(n13431) );
  OR2X1 U13307 ( .IN1(n13432), .IN2(n13433), .Q(n13426) );
  AND2X1 U13308 ( .IN1(n10695), .IN2(g805), .Q(n13433) );
  INVX0 U13309 ( .INP(n10696), .ZN(n10695) );
  AND2X1 U13310 ( .IN1(n4559), .IN2(n10696), .Q(n13432) );
  OR2X1 U13311 ( .IN1(n13434), .IN2(n13435), .Q(n10696) );
  OR2X1 U13312 ( .IN1(n13436), .IN2(n13437), .Q(n13435) );
  AND2X1 U13313 ( .IN1(g6368), .IN2(g936), .Q(n13437) );
  AND2X1 U13314 ( .IN1(g6518), .IN2(g939), .Q(n13436) );
  AND2X1 U13315 ( .IN1(test_so31), .IN2(g942), .Q(n13434) );
  OR2X1 U13316 ( .IN1(n13438), .IN2(n13439), .Q(n13427) );
  AND2X1 U13317 ( .IN1(n11983), .IN2(n10712), .Q(n13439) );
  AND2X1 U13318 ( .IN1(n10711), .IN2(n13440), .Q(n13438) );
  INVX0 U13319 ( .INP(n10712), .ZN(n10711) );
  OR2X1 U13320 ( .IN1(n13441), .IN2(n13442), .Q(n10712) );
  OR2X1 U13321 ( .IN1(n13443), .IN2(n13444), .Q(n13442) );
  AND2X1 U13322 ( .IN1(g6368), .IN2(g954), .Q(n13444) );
  AND2X1 U13323 ( .IN1(g6518), .IN2(g957), .Q(n13443) );
  AND2X1 U13324 ( .IN1(test_so31), .IN2(g960), .Q(n13441) );
  INVX0 U13325 ( .INP(n13445), .ZN(n13430) );
  AND2X1 U13326 ( .IN1(n13415), .IN2(n13413), .Q(n13445) );
  AND2X1 U13327 ( .IN1(n13422), .IN2(n13421), .Q(n13413) );
  INVX0 U13328 ( .INP(n13446), .ZN(n13421) );
  OR2X1 U13329 ( .IN1(n13447), .IN2(n13448), .Q(n13446) );
  AND2X1 U13330 ( .IN1(n10740), .IN2(g813), .Q(n13448) );
  INVX0 U13331 ( .INP(n10741), .ZN(n10740) );
  AND2X1 U13332 ( .IN1(n4289), .IN2(n10741), .Q(n13447) );
  OR2X1 U13333 ( .IN1(n13449), .IN2(n13450), .Q(n10741) );
  OR2X1 U13334 ( .IN1(n13451), .IN2(n13452), .Q(n13450) );
  AND2X1 U13335 ( .IN1(test_so35), .IN2(g6368), .Q(n13452) );
  AND2X1 U13336 ( .IN1(g6518), .IN2(g948), .Q(n13451) );
  AND2X1 U13337 ( .IN1(test_so31), .IN2(g951), .Q(n13449) );
  AND2X1 U13338 ( .IN1(n13453), .IN2(n13454), .Q(n13422) );
  OR2X1 U13339 ( .IN1(n10700), .IN2(n4375), .Q(n13454) );
  INVX0 U13340 ( .INP(n13455), .ZN(n13453) );
  AND2X1 U13341 ( .IN1(n4375), .IN2(n10700), .Q(n13455) );
  OR2X1 U13342 ( .IN1(n13456), .IN2(n13457), .Q(n10700) );
  OR2X1 U13343 ( .IN1(n13458), .IN2(n13459), .Q(n13457) );
  AND2X1 U13344 ( .IN1(g6368), .IN2(g918), .Q(n13459) );
  AND2X1 U13345 ( .IN1(g6518), .IN2(g921), .Q(n13458) );
  AND2X1 U13346 ( .IN1(test_so34), .IN2(test_so31), .Q(n13456) );
  AND2X1 U13347 ( .IN1(n13460), .IN2(n13461), .Q(n13415) );
  OR2X1 U13348 ( .IN1(n10692), .IN2(n4391), .Q(n13461) );
  INVX0 U13349 ( .INP(n13462), .ZN(n13460) );
  AND2X1 U13350 ( .IN1(n4391), .IN2(n10692), .Q(n13462) );
  OR2X1 U13351 ( .IN1(n13463), .IN2(n13464), .Q(n10692) );
  OR2X1 U13352 ( .IN1(n13465), .IN2(n13466), .Q(n13464) );
  AND2X1 U13353 ( .IN1(g6368), .IN2(g927), .Q(n13466) );
  AND2X1 U13354 ( .IN1(g6518), .IN2(g930), .Q(n13465) );
  AND2X1 U13355 ( .IN1(test_so31), .IN2(g933), .Q(n13463) );
  OR2X1 U13356 ( .IN1(n13467), .IN2(n13406), .Q(n13428) );
  OR2X1 U13357 ( .IN1(n13400), .IN2(n13398), .Q(n13406) );
  OR2X1 U13358 ( .IN1(n13468), .IN2(n13469), .Q(n13398) );
  AND2X1 U13359 ( .IN1(n13470), .IN2(n10730), .Q(n13469) );
  AND2X1 U13360 ( .IN1(n10729), .IN2(n12190), .Q(n13468) );
  INVX0 U13361 ( .INP(n10730), .ZN(n10729) );
  OR2X1 U13362 ( .IN1(n13471), .IN2(n13472), .Q(n10730) );
  OR2X1 U13363 ( .IN1(n13473), .IN2(n13474), .Q(n13472) );
  AND2X1 U13364 ( .IN1(g6368), .IN2(g909), .Q(n13474) );
  AND2X1 U13365 ( .IN1(g6518), .IN2(g912), .Q(n13473) );
  AND2X1 U13366 ( .IN1(test_so31), .IN2(g915), .Q(n13471) );
  OR2X1 U13367 ( .IN1(n13475), .IN2(n13476), .Q(n13400) );
  AND2X1 U13368 ( .IN1(n10707), .IN2(g809), .Q(n13476) );
  INVX0 U13369 ( .INP(n10708), .ZN(n10707) );
  AND2X1 U13370 ( .IN1(n4567), .IN2(n10708), .Q(n13475) );
  OR2X1 U13371 ( .IN1(n13477), .IN2(n13478), .Q(n10708) );
  OR2X1 U13372 ( .IN1(n13479), .IN2(n13480), .Q(n13478) );
  AND2X1 U13373 ( .IN1(g6368), .IN2(g900), .Q(n13480) );
  AND2X1 U13374 ( .IN1(g6518), .IN2(g903), .Q(n13479) );
  AND2X1 U13375 ( .IN1(test_so31), .IN2(g906), .Q(n13477) );
  OR2X1 U13376 ( .IN1(n13394), .IN2(n13402), .Q(n13467) );
  OR2X1 U13377 ( .IN1(n13397), .IN2(n13399), .Q(n13402) );
  OR2X1 U13378 ( .IN1(n13481), .IN2(n13482), .Q(n13399) );
  AND2X1 U13379 ( .IN1(n10715), .IN2(g785), .Q(n13482) );
  INVX0 U13380 ( .INP(n10716), .ZN(n10715) );
  AND2X1 U13381 ( .IN1(n4379), .IN2(n10716), .Q(n13481) );
  OR2X1 U13382 ( .IN1(n13483), .IN2(n13484), .Q(n10716) );
  OR2X1 U13383 ( .IN1(n13485), .IN2(n13486), .Q(n13484) );
  AND2X1 U13384 ( .IN1(g6368), .IN2(g873), .Q(n13486) );
  AND2X1 U13385 ( .IN1(g6518), .IN2(g876), .Q(n13485) );
  AND2X1 U13386 ( .IN1(test_so31), .IN2(g879), .Q(n13483) );
  OR2X1 U13387 ( .IN1(n13487), .IN2(n13488), .Q(n13397) );
  AND2X1 U13388 ( .IN1(n10733), .IN2(g793), .Q(n13488) );
  INVX0 U13389 ( .INP(n10734), .ZN(n10733) );
  AND2X1 U13390 ( .IN1(n4321), .IN2(n10734), .Q(n13487) );
  OR2X1 U13391 ( .IN1(n13489), .IN2(n13490), .Q(n10734) );
  OR2X1 U13392 ( .IN1(n13491), .IN2(n13492), .Q(n13490) );
  AND2X1 U13393 ( .IN1(g6368), .IN2(g882), .Q(n13492) );
  AND2X1 U13394 ( .IN1(g6518), .IN2(g885), .Q(n13491) );
  AND2X1 U13395 ( .IN1(test_so31), .IN2(g888), .Q(n13489) );
  OR2X1 U13396 ( .IN1(n13493), .IN2(n13494), .Q(n13394) );
  AND2X1 U13397 ( .IN1(n10725), .IN2(g801), .Q(n13494) );
  INVX0 U13398 ( .INP(n10726), .ZN(n10725) );
  AND2X1 U13399 ( .IN1(n4327), .IN2(n10726), .Q(n13493) );
  OR2X1 U13400 ( .IN1(n13495), .IN2(n13496), .Q(n10726) );
  OR2X1 U13401 ( .IN1(n13497), .IN2(n13498), .Q(n13496) );
  AND2X1 U13402 ( .IN1(g6368), .IN2(g891), .Q(n13498) );
  AND2X1 U13403 ( .IN1(g6518), .IN2(g894), .Q(n13497) );
  AND2X1 U13404 ( .IN1(test_so31), .IN2(g897), .Q(n13495) );
  AND2X1 U13405 ( .IN1(n4387), .IN2(n13499), .Q(n13382) );
  OR2X1 U13406 ( .IN1(n13500), .IN2(n13501), .Q(g29169) );
  AND2X1 U13407 ( .IN1(n13374), .IN2(n13502), .Q(n13501) );
  AND2X1 U13408 ( .IN1(n13503), .IN2(g323), .Q(n13500) );
  OR2X1 U13409 ( .IN1(n4499), .IN2(n13377), .Q(n13503) );
  OR2X1 U13410 ( .IN1(n13504), .IN2(n13505), .Q(g29167) );
  AND2X1 U13411 ( .IN1(n13374), .IN2(n13506), .Q(n13505) );
  AND2X1 U13412 ( .IN1(n13377), .IN2(n13507), .Q(n13374) );
  INVX0 U13413 ( .INP(n13508), .ZN(n13507) );
  OR2X1 U13414 ( .IN1(n13509), .IN2(n13510), .Q(n13508) );
  AND2X1 U13415 ( .IN1(n12293), .IN2(n12811), .Q(n13510) );
  AND2X1 U13416 ( .IN1(n13511), .IN2(g322), .Q(n13504) );
  OR2X1 U13417 ( .IN1(n4520), .IN2(n13377), .Q(n13511) );
  OR2X1 U13418 ( .IN1(n12813), .IN2(n13512), .Q(n13377) );
  OR2X1 U13419 ( .IN1(n13509), .IN2(n13513), .Q(n13512) );
  AND2X1 U13420 ( .IN1(n13514), .IN2(n12811), .Q(n13513) );
  OR2X1 U13421 ( .IN1(n12293), .IN2(n13515), .Q(n13514) );
  OR2X1 U13422 ( .IN1(n11851), .IN2(n12300), .Q(n13515) );
  OR2X1 U13423 ( .IN1(n11831), .IN2(n12810), .Q(n12300) );
  OR2X1 U13424 ( .IN1(n11849), .IN2(n13516), .Q(n12810) );
  AND2X1 U13425 ( .IN1(n3130), .IN2(n13517), .Q(n13516) );
  OR2X1 U13426 ( .IN1(n11847), .IN2(n11844), .Q(n13517) );
  OR2X1 U13427 ( .IN1(n13518), .IN2(n13519), .Q(n11844) );
  AND2X1 U13428 ( .IN1(n13520), .IN2(n13521), .Q(n13519) );
  AND2X1 U13429 ( .IN1(n13522), .IN2(n13523), .Q(n13520) );
  OR2X1 U13430 ( .IN1(n13524), .IN2(n13525), .Q(n13523) );
  OR2X1 U13431 ( .IN1(n13526), .IN2(n13527), .Q(n13522) );
  AND2X1 U13432 ( .IN1(n13528), .IN2(n13525), .Q(n13518) );
  AND2X1 U13433 ( .IN1(n13529), .IN2(n13530), .Q(n13528) );
  OR2X1 U13434 ( .IN1(n13521), .IN2(n13527), .Q(n13530) );
  AND2X1 U13435 ( .IN1(n13526), .IN2(n13531), .Q(n11847) );
  AND2X1 U13436 ( .IN1(n13532), .IN2(n13533), .Q(n13531) );
  OR2X1 U13437 ( .IN1(n13521), .IN2(n13524), .Q(n13532) );
  INVX0 U13438 ( .INP(n11834), .ZN(n11849) );
  OR2X1 U13439 ( .IN1(n13534), .IN2(n11838), .Q(n11834) );
  AND2X1 U13440 ( .IN1(n13535), .IN2(n13536), .Q(n13534) );
  OR2X1 U13441 ( .IN1(n13537), .IN2(n13538), .Q(n13536) );
  OR2X1 U13442 ( .IN1(n13539), .IN2(n13540), .Q(n13538) );
  AND2X1 U13443 ( .IN1(n13541), .IN2(n13542), .Q(n13540) );
  AND2X1 U13444 ( .IN1(n13543), .IN2(n13544), .Q(n13539) );
  AND2X1 U13445 ( .IN1(n13545), .IN2(n13546), .Q(n13535) );
  OR2X1 U13446 ( .IN1(n13543), .IN2(n13547), .Q(n13546) );
  OR2X1 U13447 ( .IN1(n13548), .IN2(n13549), .Q(n13547) );
  AND2X1 U13448 ( .IN1(n13537), .IN2(n13541), .Q(n13549) );
  OR2X1 U13449 ( .IN1(n13542), .IN2(n13550), .Q(n13545) );
  OR2X1 U13450 ( .IN1(n13551), .IN2(n13552), .Q(n13550) );
  AND2X1 U13451 ( .IN1(n13543), .IN2(n13541), .Q(n13552) );
  INVX0 U13452 ( .INP(n13553), .ZN(n13541) );
  INVX0 U13453 ( .INP(n13554), .ZN(n13543) );
  AND2X1 U13454 ( .IN1(n13537), .IN2(n13544), .Q(n13551) );
  INVX0 U13455 ( .INP(n13555), .ZN(n13537) );
  OR2X1 U13456 ( .IN1(n11850), .IN2(n11838), .Q(n12293) );
  INVX0 U13457 ( .INP(n11839), .ZN(n11850) );
  OR2X1 U13458 ( .IN1(n13556), .IN2(n13557), .Q(n11839) );
  OR2X1 U13459 ( .IN1(n13558), .IN2(n13533), .Q(n13557) );
  OR2X1 U13460 ( .IN1(n13525), .IN2(n13527), .Q(n13533) );
  OR2X1 U13461 ( .IN1(n13559), .IN2(n13560), .Q(n13527) );
  AND2X1 U13462 ( .IN1(n10642), .IN2(g121), .Q(n13560) );
  INVX0 U13463 ( .INP(n10643), .ZN(n10642) );
  AND2X1 U13464 ( .IN1(n4569), .IN2(n10643), .Q(n13559) );
  OR2X1 U13465 ( .IN1(n13561), .IN2(n13562), .Q(n10643) );
  OR2X1 U13466 ( .IN1(n13563), .IN2(n13564), .Q(n13562) );
  AND2X1 U13467 ( .IN1(g165), .IN2(g219), .Q(n13564) );
  AND2X1 U13468 ( .IN1(g6231), .IN2(g213), .Q(n13563) );
  AND2X1 U13469 ( .IN1(g6313), .IN2(g216), .Q(n13561) );
  OR2X1 U13470 ( .IN1(n13565), .IN2(n13566), .Q(n13525) );
  AND2X1 U13471 ( .IN1(n13567), .IN2(n10651), .Q(n13566) );
  AND2X1 U13472 ( .IN1(n10650), .IN2(n12218), .Q(n13565) );
  INVX0 U13473 ( .INP(n10651), .ZN(n10650) );
  OR2X1 U13474 ( .IN1(n13568), .IN2(n13569), .Q(n10651) );
  OR2X1 U13475 ( .IN1(n13570), .IN2(n13571), .Q(n13569) );
  AND2X1 U13476 ( .IN1(g165), .IN2(g228), .Q(n13571) );
  AND2X1 U13477 ( .IN1(g6231), .IN2(g222), .Q(n13570) );
  AND2X1 U13478 ( .IN1(g6313), .IN2(g225), .Q(n13568) );
  OR2X1 U13479 ( .IN1(n13521), .IN2(n13529), .Q(n13558) );
  OR2X1 U13480 ( .IN1(n13524), .IN2(n13526), .Q(n13529) );
  OR2X1 U13481 ( .IN1(n13572), .IN2(n13573), .Q(n13526) );
  AND2X1 U13482 ( .IN1(n4380), .IN2(n12831), .Q(n13573) );
  INVX0 U13483 ( .INP(n4513), .ZN(n12831) );
  AND2X1 U13484 ( .IN1(n4513), .IN2(g97), .Q(n13572) );
  OR2X1 U13485 ( .IN1(n13574), .IN2(n13575), .Q(n13524) );
  AND2X1 U13486 ( .IN1(n10663), .IN2(g105), .Q(n13575) );
  INVX0 U13487 ( .INP(n10664), .ZN(n10663) );
  AND2X1 U13488 ( .IN1(n4322), .IN2(n10664), .Q(n13574) );
  OR2X1 U13489 ( .IN1(n13576), .IN2(n13577), .Q(n10664) );
  OR2X1 U13490 ( .IN1(n13578), .IN2(n13579), .Q(n13577) );
  AND2X1 U13491 ( .IN1(g165), .IN2(g201), .Q(n13579) );
  AND2X1 U13492 ( .IN1(g6231), .IN2(g195), .Q(n13578) );
  AND2X1 U13493 ( .IN1(g6313), .IN2(g198), .Q(n13576) );
  OR2X1 U13494 ( .IN1(n13580), .IN2(n13581), .Q(n13521) );
  AND2X1 U13495 ( .IN1(n10667), .IN2(g113), .Q(n13581) );
  INVX0 U13496 ( .INP(n10668), .ZN(n10667) );
  AND2X1 U13497 ( .IN1(n4328), .IN2(n10668), .Q(n13580) );
  OR2X1 U13498 ( .IN1(n13582), .IN2(n13583), .Q(n10668) );
  OR2X1 U13499 ( .IN1(n13584), .IN2(n13585), .Q(n13583) );
  AND2X1 U13500 ( .IN1(g165), .IN2(g210), .Q(n13585) );
  AND2X1 U13501 ( .IN1(g6231), .IN2(g204), .Q(n13584) );
  AND2X1 U13502 ( .IN1(g6313), .IN2(g207), .Q(n13582) );
  OR2X1 U13503 ( .IN1(n13586), .IN2(n13587), .Q(n13556) );
  OR2X1 U13504 ( .IN1(n13555), .IN2(n13554), .Q(n13587) );
  OR2X1 U13505 ( .IN1(n13588), .IN2(n13589), .Q(n13554) );
  AND2X1 U13506 ( .IN1(n12036), .IN2(n10647), .Q(n13589) );
  AND2X1 U13507 ( .IN1(n10646), .IN2(n13590), .Q(n13588) );
  INVX0 U13508 ( .INP(n10647), .ZN(n10646) );
  OR2X1 U13509 ( .IN1(n13591), .IN2(n13592), .Q(n10647) );
  OR2X1 U13510 ( .IN1(n13593), .IN2(n13594), .Q(n13592) );
  AND2X1 U13511 ( .IN1(g165), .IN2(g273), .Q(n13594) );
  AND2X1 U13512 ( .IN1(g6231), .IN2(g267), .Q(n13593) );
  AND2X1 U13513 ( .IN1(g6313), .IN2(g270), .Q(n13591) );
  OR2X1 U13514 ( .IN1(n13595), .IN2(n13596), .Q(n13555) );
  AND2X1 U13515 ( .IN1(n10630), .IN2(g117), .Q(n13596) );
  INVX0 U13516 ( .INP(n10631), .ZN(n10630) );
  AND2X1 U13517 ( .IN1(n4561), .IN2(n10631), .Q(n13595) );
  OR2X1 U13518 ( .IN1(n13597), .IN2(n13598), .Q(n10631) );
  OR2X1 U13519 ( .IN1(n13599), .IN2(n13600), .Q(n13598) );
  AND2X1 U13520 ( .IN1(test_so14), .IN2(g165), .Q(n13600) );
  AND2X1 U13521 ( .IN1(g6231), .IN2(g249), .Q(n13599) );
  AND2X1 U13522 ( .IN1(g6313), .IN2(g252), .Q(n13597) );
  OR2X1 U13523 ( .IN1(n13553), .IN2(n13601), .Q(n13586) );
  INVX0 U13524 ( .INP(n13548), .ZN(n13601) );
  AND2X1 U13525 ( .IN1(n13542), .IN2(n13544), .Q(n13548) );
  AND2X1 U13526 ( .IN1(n13602), .IN2(n13603), .Q(n13544) );
  OR2X1 U13527 ( .IN1(n10676), .IN2(n4392), .Q(n13603) );
  OR2X1 U13528 ( .IN1(g109), .IN2(n10675), .Q(n13602) );
  INVX0 U13529 ( .INP(n10676), .ZN(n10675) );
  OR2X1 U13530 ( .IN1(n13604), .IN2(n13605), .Q(n10676) );
  OR2X1 U13531 ( .IN1(n13606), .IN2(n13607), .Q(n13605) );
  AND2X1 U13532 ( .IN1(g165), .IN2(g246), .Q(n13607) );
  AND2X1 U13533 ( .IN1(g6231), .IN2(g240), .Q(n13606) );
  AND2X1 U13534 ( .IN1(g6313), .IN2(g243), .Q(n13604) );
  AND2X1 U13535 ( .IN1(n13608), .IN2(n13609), .Q(n13542) );
  OR2X1 U13536 ( .IN1(n10627), .IN2(n4376), .Q(n13609) );
  OR2X1 U13537 ( .IN1(g101), .IN2(n10626), .Q(n13608) );
  INVX0 U13538 ( .INP(n10627), .ZN(n10626) );
  OR2X1 U13539 ( .IN1(n13610), .IN2(n13611), .Q(n10627) );
  OR2X1 U13540 ( .IN1(n13612), .IN2(n13613), .Q(n13611) );
  AND2X1 U13541 ( .IN1(g165), .IN2(g237), .Q(n13613) );
  AND2X1 U13542 ( .IN1(g6231), .IN2(g231), .Q(n13612) );
  AND2X1 U13543 ( .IN1(g6313), .IN2(g234), .Q(n13610) );
  OR2X1 U13544 ( .IN1(n13614), .IN2(n13615), .Q(n13553) );
  AND2X1 U13545 ( .IN1(n10634), .IN2(g125), .Q(n13615) );
  INVX0 U13546 ( .INP(n10635), .ZN(n10634) );
  AND2X1 U13547 ( .IN1(n4290), .IN2(n10635), .Q(n13614) );
  OR2X1 U13548 ( .IN1(n13616), .IN2(n13617), .Q(n10635) );
  OR2X1 U13549 ( .IN1(n13618), .IN2(n13619), .Q(n13617) );
  AND2X1 U13550 ( .IN1(g165), .IN2(g264), .Q(n13619) );
  AND2X1 U13551 ( .IN1(g6231), .IN2(g258), .Q(n13618) );
  AND2X1 U13552 ( .IN1(g6313), .IN2(g261), .Q(n13616) );
  AND2X1 U13553 ( .IN1(n4388), .IN2(n13620), .Q(n13509) );
  AND2X1 U13554 ( .IN1(n13621), .IN2(n12966), .Q(g29112) );
  AND2X1 U13555 ( .IN1(n13622), .IN2(n1577), .Q(n13621) );
  OR2X1 U13556 ( .IN1(n10175), .IN2(n13623), .Q(n1577) );
  INVX0 U13557 ( .INP(n3159), .ZN(n13623) );
  OR2X1 U13558 ( .IN1(n3159), .IN2(g2129), .Q(n13622) );
  AND2X1 U13559 ( .IN1(n13624), .IN2(n12971), .Q(g29111) );
  AND2X1 U13560 ( .IN1(n13625), .IN2(n1233), .Q(n13624) );
  OR2X1 U13561 ( .IN1(n10174), .IN2(n13626), .Q(n1233) );
  INVX0 U13562 ( .INP(n3163), .ZN(n13626) );
  OR2X1 U13563 ( .IN1(n3163), .IN2(g1435), .Q(n13625) );
  AND2X1 U13564 ( .IN1(n13627), .IN2(n12976), .Q(g29110) );
  OR2X1 U13565 ( .IN1(n13628), .IN2(n13629), .Q(n13627) );
  AND2X1 U13566 ( .IN1(n3167), .IN2(n10195), .Q(n13629) );
  AND2X1 U13567 ( .IN1(test_so36), .IN2(n12997), .Q(n13628) );
  INVX0 U13568 ( .INP(n3167), .ZN(n12997) );
  AND2X1 U13569 ( .IN1(n13630), .IN2(n12981), .Q(g29109) );
  AND2X1 U13570 ( .IN1(n13631), .IN2(n470), .Q(n13630) );
  OR2X1 U13571 ( .IN1(n10176), .IN2(n13632), .Q(n470) );
  INVX0 U13572 ( .INP(n3171), .ZN(n13632) );
  OR2X1 U13573 ( .IN1(n3171), .IN2(g61), .Q(n13631) );
  OR2X1 U13574 ( .IN1(n13633), .IN2(n13634), .Q(g28788) );
  AND2X1 U13575 ( .IN1(n13635), .IN2(n13101), .Q(n13634) );
  AND2X1 U13576 ( .IN1(n13636), .IN2(g2501), .Q(n13633) );
  OR2X1 U13577 ( .IN1(n4509), .IN2(n13637), .Q(n13636) );
  OR2X1 U13578 ( .IN1(n13638), .IN2(n13639), .Q(g28783) );
  AND2X1 U13579 ( .IN1(n13635), .IN2(n13106), .Q(n13639) );
  AND2X1 U13580 ( .IN1(n13640), .IN2(g2503), .Q(n13638) );
  OR2X1 U13581 ( .IN1(n4524), .IN2(n13637), .Q(n13640) );
  OR2X1 U13582 ( .IN1(n13641), .IN2(n13642), .Q(g28782) );
  AND2X1 U13583 ( .IN1(test_so80), .IN2(n4509), .Q(n13642) );
  AND2X1 U13584 ( .IN1(n4606), .IN2(n13643), .Q(n13641) );
  OR2X1 U13585 ( .IN1(n13644), .IN2(n13645), .Q(g28778) );
  AND2X1 U13586 ( .IN1(n13646), .IN2(n13111), .Q(n13645) );
  AND2X1 U13587 ( .IN1(n13647), .IN2(g1807), .Q(n13644) );
  OR2X1 U13588 ( .IN1(n4511), .IN2(n13648), .Q(n13647) );
  OR2X1 U13589 ( .IN1(n13649), .IN2(n13650), .Q(g28774) );
  AND2X1 U13590 ( .IN1(n13635), .IN2(n13116), .Q(n13650) );
  AND2X1 U13591 ( .IN1(n13651), .IN2(g2502), .Q(n13649) );
  OR2X1 U13592 ( .IN1(n4516), .IN2(n13637), .Q(n13651) );
  OR2X1 U13593 ( .IN1(n13652), .IN2(n13653), .Q(n13637) );
  OR2X1 U13594 ( .IN1(n13654), .IN2(n10191), .Q(n13653) );
  INVX0 U13595 ( .INP(n13655), .ZN(n13654) );
  OR2X1 U13596 ( .IN1(n13656), .IN2(n13657), .Q(g28773) );
  AND2X1 U13597 ( .IN1(n4524), .IN2(g2486), .Q(n13657) );
  AND2X1 U13598 ( .IN1(g7264), .IN2(n13643), .Q(n13656) );
  OR2X1 U13599 ( .IN1(n13658), .IN2(n13659), .Q(g28772) );
  AND2X1 U13600 ( .IN1(n13646), .IN2(n13239), .Q(n13659) );
  AND2X1 U13601 ( .IN1(n13660), .IN2(g1809), .Q(n13658) );
  OR2X1 U13602 ( .IN1(n4525), .IN2(n13648), .Q(n13660) );
  OR2X1 U13603 ( .IN1(n13661), .IN2(n13662), .Q(g28771) );
  AND2X1 U13604 ( .IN1(n4511), .IN2(g1795), .Q(n13662) );
  AND2X1 U13605 ( .IN1(n4618), .IN2(n13663), .Q(n13661) );
  OR2X1 U13606 ( .IN1(n13664), .IN2(n13665), .Q(g28767) );
  AND2X1 U13607 ( .IN1(n13666), .IN2(g1088), .Q(n13665) );
  AND2X1 U13608 ( .IN1(n13667), .IN2(g1113), .Q(n13664) );
  OR2X1 U13609 ( .IN1(n4381), .IN2(n13668), .Q(n13667) );
  OR2X1 U13610 ( .IN1(n13669), .IN2(n13670), .Q(g28763) );
  AND2X1 U13611 ( .IN1(n4516), .IN2(g2483), .Q(n13670) );
  AND2X1 U13612 ( .IN1(g5555), .IN2(n13643), .Q(n13669) );
  OR2X1 U13613 ( .IN1(n13671), .IN2(n13635), .Q(n13643) );
  AND2X1 U13614 ( .IN1(n13024), .IN2(n13672), .Q(n13635) );
  AND2X1 U13615 ( .IN1(n13655), .IN2(test_so79), .Q(n13672) );
  INVX0 U13616 ( .INP(n13673), .ZN(n13024) );
  AND2X1 U13617 ( .IN1(n13674), .IN2(n13673), .Q(n13671) );
  OR2X1 U13618 ( .IN1(n13675), .IN2(n13676), .Q(n13673) );
  OR2X1 U13619 ( .IN1(n13677), .IN2(n13678), .Q(n13676) );
  AND2X1 U13620 ( .IN1(g7264), .IN2(g2486), .Q(n13678) );
  AND2X1 U13621 ( .IN1(test_so80), .IN2(n4606), .Q(n13677) );
  AND2X1 U13622 ( .IN1(g5555), .IN2(g2483), .Q(n13675) );
  OR2X1 U13623 ( .IN1(n13679), .IN2(n10191), .Q(n13674) );
  AND2X1 U13624 ( .IN1(n13025), .IN2(n13655), .Q(n13679) );
  OR2X1 U13625 ( .IN1(n13680), .IN2(n13681), .Q(n13655) );
  AND2X1 U13626 ( .IN1(n13682), .IN2(n13016), .Q(n13681) );
  AND2X1 U13627 ( .IN1(n13028), .IN2(n12235), .Q(n13682) );
  OR2X1 U13628 ( .IN1(n10162), .IN2(n11734), .Q(n12235) );
  OR2X1 U13629 ( .IN1(n13683), .IN2(n13684), .Q(n11734) );
  OR2X1 U13630 ( .IN1(n13685), .IN2(n13686), .Q(n13684) );
  AND2X1 U13631 ( .IN1(n9764), .IN2(g2241), .Q(n13686) );
  AND2X1 U13632 ( .IN1(n9766), .IN2(g6837), .Q(n13685) );
  AND2X1 U13633 ( .IN1(n9765), .IN2(test_so73), .Q(n13683) );
  INVX0 U13634 ( .INP(n13022), .ZN(n13028) );
  AND2X1 U13635 ( .IN1(n13022), .IN2(n4285), .Q(n13680) );
  OR2X1 U13636 ( .IN1(n13687), .IN2(n13688), .Q(n13022) );
  OR2X1 U13637 ( .IN1(n13179), .IN2(n11898), .Q(n13688) );
  INVX0 U13638 ( .INP(n13652), .ZN(n13025) );
  OR2X1 U13639 ( .IN1(n13689), .IN2(n13690), .Q(n13652) );
  OR2X1 U13640 ( .IN1(n13691), .IN2(n13692), .Q(n13690) );
  AND2X1 U13641 ( .IN1(n9855), .IN2(n13116), .Q(n13692) );
  AND2X1 U13642 ( .IN1(n9854), .IN2(n13101), .Q(n13691) );
  AND2X1 U13643 ( .IN1(n9845), .IN2(n13106), .Q(n13689) );
  OR2X1 U13644 ( .IN1(n13693), .IN2(n13694), .Q(g28761) );
  AND2X1 U13645 ( .IN1(n13646), .IN2(n13248), .Q(n13694) );
  AND2X1 U13646 ( .IN1(n13695), .IN2(g1808), .Q(n13693) );
  OR2X1 U13647 ( .IN1(n4518), .IN2(n13648), .Q(n13695) );
  OR2X1 U13648 ( .IN1(n13696), .IN2(n13697), .Q(n13648) );
  OR2X1 U13649 ( .IN1(n4386), .IN2(n13698), .Q(n13697) );
  INVX0 U13650 ( .INP(n13699), .ZN(n13698) );
  OR2X1 U13651 ( .IN1(n13700), .IN2(n13701), .Q(g28760) );
  AND2X1 U13652 ( .IN1(n4525), .IN2(g1792), .Q(n13701) );
  AND2X1 U13653 ( .IN1(g7014), .IN2(n13663), .Q(n13700) );
  OR2X1 U13654 ( .IN1(n13702), .IN2(n13703), .Q(g28759) );
  AND2X1 U13655 ( .IN1(n13666), .IN2(g6712), .Q(n13703) );
  AND2X1 U13656 ( .IN1(n13704), .IN2(g1115), .Q(n13702) );
  OR2X1 U13657 ( .IN1(n4364), .IN2(n13668), .Q(n13704) );
  OR2X1 U13658 ( .IN1(n13705), .IN2(n13706), .Q(g28758) );
  AND2X1 U13659 ( .IN1(n13707), .IN2(g1088), .Q(n13706) );
  AND2X1 U13660 ( .IN1(n4381), .IN2(g1101), .Q(n13705) );
  OR2X1 U13661 ( .IN1(n13708), .IN2(n13709), .Q(g28754) );
  AND2X1 U13662 ( .IN1(n13710), .IN2(n13375), .Q(n13709) );
  AND2X1 U13663 ( .IN1(n13711), .IN2(g426), .Q(n13708) );
  OR2X1 U13664 ( .IN1(n4506), .IN2(n13712), .Q(n13711) );
  OR2X1 U13665 ( .IN1(n13713), .IN2(n13714), .Q(g28749) );
  AND2X1 U13666 ( .IN1(n4518), .IN2(g1789), .Q(n13714) );
  AND2X1 U13667 ( .IN1(g5511), .IN2(n13663), .Q(n13713) );
  OR2X1 U13668 ( .IN1(n13715), .IN2(n13646), .Q(n13663) );
  AND2X1 U13669 ( .IN1(n13048), .IN2(n13716), .Q(n13646) );
  AND2X1 U13670 ( .IN1(g1690), .IN2(n13699), .Q(n13716) );
  INVX0 U13671 ( .INP(n13717), .ZN(n13048) );
  AND2X1 U13672 ( .IN1(n13718), .IN2(n13717), .Q(n13715) );
  OR2X1 U13673 ( .IN1(n13719), .IN2(n13720), .Q(n13717) );
  OR2X1 U13674 ( .IN1(n13721), .IN2(n13722), .Q(n13720) );
  AND2X1 U13675 ( .IN1(g7014), .IN2(g1792), .Q(n13722) );
  AND2X1 U13676 ( .IN1(n4618), .IN2(g1795), .Q(n13721) );
  AND2X1 U13677 ( .IN1(g5511), .IN2(g1789), .Q(n13719) );
  OR2X1 U13678 ( .IN1(n13723), .IN2(n4386), .Q(n13718) );
  AND2X1 U13679 ( .IN1(n13049), .IN2(n13699), .Q(n13723) );
  OR2X1 U13680 ( .IN1(n13724), .IN2(n13725), .Q(n13699) );
  AND2X1 U13681 ( .IN1(n13726), .IN2(n13040), .Q(n13725) );
  AND2X1 U13682 ( .IN1(n13052), .IN2(n11772), .Q(n13726) );
  OR2X1 U13683 ( .IN1(n10161), .IN2(n11737), .Q(n11772) );
  OR2X1 U13684 ( .IN1(n13727), .IN2(n13728), .Q(n11737) );
  OR2X1 U13685 ( .IN1(n13729), .IN2(n13730), .Q(n13728) );
  AND2X1 U13686 ( .IN1(n9775), .IN2(g1547), .Q(n13730) );
  AND2X1 U13687 ( .IN1(n9777), .IN2(g6573), .Q(n13729) );
  AND2X1 U13688 ( .IN1(n9776), .IN2(g6782), .Q(n13727) );
  INVX0 U13689 ( .INP(n13046), .ZN(n13052) );
  AND2X1 U13690 ( .IN1(n13046), .IN2(n4284), .Q(n13724) );
  OR2X1 U13691 ( .IN1(n13731), .IN2(n13732), .Q(n13046) );
  OR2X1 U13692 ( .IN1(n13311), .IN2(n11936), .Q(n13732) );
  INVX0 U13693 ( .INP(n13696), .ZN(n13049) );
  OR2X1 U13694 ( .IN1(n13733), .IN2(n13734), .Q(n13696) );
  OR2X1 U13695 ( .IN1(n13735), .IN2(n13736), .Q(n13734) );
  AND2X1 U13696 ( .IN1(n9860), .IN2(n13248), .Q(n13736) );
  AND2X1 U13697 ( .IN1(n9859), .IN2(n13111), .Q(n13735) );
  AND2X1 U13698 ( .IN1(n9848), .IN2(n13239), .Q(n13733) );
  OR2X1 U13699 ( .IN1(n13737), .IN2(n13738), .Q(g28747) );
  AND2X1 U13700 ( .IN1(n13666), .IN2(g5472), .Q(n13738) );
  AND2X1 U13701 ( .IN1(n13739), .IN2(g1114), .Q(n13737) );
  OR2X1 U13702 ( .IN1(n4363), .IN2(n13668), .Q(n13739) );
  OR2X1 U13703 ( .IN1(n13740), .IN2(n13741), .Q(n13668) );
  OR2X1 U13704 ( .IN1(n4387), .IN2(n13742), .Q(n13741) );
  INVX0 U13705 ( .INP(n13743), .ZN(n13742) );
  OR2X1 U13706 ( .IN1(n13744), .IN2(n13745), .Q(g28746) );
  AND2X1 U13707 ( .IN1(n13707), .IN2(g6712), .Q(n13745) );
  AND2X1 U13708 ( .IN1(n4364), .IN2(g1098), .Q(n13744) );
  OR2X1 U13709 ( .IN1(n13746), .IN2(n13747), .Q(g28745) );
  AND2X1 U13710 ( .IN1(n13710), .IN2(n13502), .Q(n13747) );
  AND2X1 U13711 ( .IN1(n13748), .IN2(g428), .Q(n13746) );
  OR2X1 U13712 ( .IN1(n4499), .IN2(n13712), .Q(n13748) );
  OR2X1 U13713 ( .IN1(n13749), .IN2(n13750), .Q(g28744) );
  AND2X1 U13714 ( .IN1(n4506), .IN2(g414), .Q(n13750) );
  AND2X1 U13715 ( .IN1(n4640), .IN2(n13751), .Q(n13749) );
  OR2X1 U13716 ( .IN1(n13752), .IN2(n13753), .Q(g28738) );
  AND2X1 U13717 ( .IN1(n13707), .IN2(g5472), .Q(n13753) );
  OR2X1 U13718 ( .IN1(n13754), .IN2(n13666), .Q(n13707) );
  AND2X1 U13719 ( .IN1(n13072), .IN2(n13755), .Q(n13666) );
  AND2X1 U13720 ( .IN1(g996), .IN2(n13743), .Q(n13755) );
  INVX0 U13721 ( .INP(n13756), .ZN(n13072) );
  AND2X1 U13722 ( .IN1(n13757), .IN2(n13756), .Q(n13754) );
  OR2X1 U13723 ( .IN1(n13758), .IN2(n13759), .Q(n13756) );
  OR2X1 U13724 ( .IN1(n13760), .IN2(n13761), .Q(n13759) );
  AND2X1 U13725 ( .IN1(g6712), .IN2(g1098), .Q(n13761) );
  AND2X1 U13726 ( .IN1(g5472), .IN2(g1095), .Q(n13760) );
  AND2X1 U13727 ( .IN1(g1088), .IN2(g1101), .Q(n13758) );
  OR2X1 U13728 ( .IN1(n13762), .IN2(n4387), .Q(n13757) );
  AND2X1 U13729 ( .IN1(n13073), .IN2(n13743), .Q(n13762) );
  OR2X1 U13730 ( .IN1(n13763), .IN2(n13764), .Q(n13743) );
  AND2X1 U13731 ( .IN1(n13765), .IN2(n13064), .Q(n13764) );
  AND2X1 U13732 ( .IN1(n13076), .IN2(n11577), .Q(n13765) );
  OR2X1 U13733 ( .IN1(n10160), .IN2(n10600), .Q(n11577) );
  OR2X1 U13734 ( .IN1(n13766), .IN2(n13767), .Q(n10600) );
  OR2X1 U13735 ( .IN1(n13768), .IN2(n13769), .Q(n13767) );
  AND2X1 U13736 ( .IN1(n9788), .IN2(g6368), .Q(n13769) );
  AND2X1 U13737 ( .IN1(g6518), .IN2(n10206), .Q(n13768) );
  AND2X1 U13738 ( .IN1(test_so31), .IN2(n9787), .Q(n13766) );
  INVX0 U13739 ( .INP(n13070), .ZN(n13076) );
  AND2X1 U13740 ( .IN1(n13070), .IN2(n4283), .Q(n13763) );
  OR2X1 U13741 ( .IN1(n13770), .IN2(n13771), .Q(n13070) );
  OR2X1 U13742 ( .IN1(n11983), .IN2(n13470), .Q(n13771) );
  INVX0 U13743 ( .INP(n13740), .ZN(n13073) );
  OR2X1 U13744 ( .IN1(n13772), .IN2(n13773), .Q(n13740) );
  OR2X1 U13745 ( .IN1(n13774), .IN2(n13775), .Q(n13773) );
  AND2X1 U13746 ( .IN1(n9851), .IN2(g6712), .Q(n13775) );
  AND2X1 U13747 ( .IN1(n9866), .IN2(g5472), .Q(n13774) );
  AND2X1 U13748 ( .IN1(n9865), .IN2(g1088), .Q(n13772) );
  AND2X1 U13749 ( .IN1(n4363), .IN2(g1095), .Q(n13752) );
  OR2X1 U13750 ( .IN1(n13776), .IN2(n13777), .Q(g28736) );
  AND2X1 U13751 ( .IN1(n13710), .IN2(n13506), .Q(n13777) );
  AND2X1 U13752 ( .IN1(test_so17), .IN2(n13778), .Q(n13776) );
  OR2X1 U13753 ( .IN1(n4520), .IN2(n13712), .Q(n13778) );
  INVX0 U13754 ( .INP(n13779), .ZN(n13712) );
  AND2X1 U13755 ( .IN1(n13094), .IN2(n13780), .Q(n13779) );
  OR2X1 U13756 ( .IN1(n13781), .IN2(n13782), .Q(g28735) );
  AND2X1 U13757 ( .IN1(n4499), .IN2(g411), .Q(n13782) );
  AND2X1 U13758 ( .IN1(g6447), .IN2(n13751), .Q(n13781) );
  OR2X1 U13759 ( .IN1(n13783), .IN2(n13784), .Q(g28732) );
  AND2X1 U13760 ( .IN1(n4520), .IN2(g408), .Q(n13784) );
  AND2X1 U13761 ( .IN1(g5437), .IN2(n13751), .Q(n13783) );
  OR2X1 U13762 ( .IN1(n13785), .IN2(n13710), .Q(n13751) );
  AND2X1 U13763 ( .IN1(n13093), .IN2(n13780), .Q(n13710) );
  AND2X1 U13764 ( .IN1(g309), .IN2(n13786), .Q(n13780) );
  INVX0 U13765 ( .INP(n13787), .ZN(n13093) );
  AND2X1 U13766 ( .IN1(n13788), .IN2(n13787), .Q(n13785) );
  OR2X1 U13767 ( .IN1(n13789), .IN2(n13790), .Q(n13787) );
  OR2X1 U13768 ( .IN1(n13791), .IN2(n13792), .Q(n13790) );
  AND2X1 U13769 ( .IN1(g6447), .IN2(g411), .Q(n13792) );
  AND2X1 U13770 ( .IN1(n4640), .IN2(g414), .Q(n13791) );
  AND2X1 U13771 ( .IN1(g5437), .IN2(g408), .Q(n13789) );
  OR2X1 U13772 ( .IN1(n13793), .IN2(n4388), .Q(n13788) );
  AND2X1 U13773 ( .IN1(n13094), .IN2(n13786), .Q(n13793) );
  OR2X1 U13774 ( .IN1(n13794), .IN2(n13795), .Q(n13786) );
  AND2X1 U13775 ( .IN1(n13796), .IN2(n13085), .Q(n13795) );
  AND2X1 U13776 ( .IN1(n13097), .IN2(n11825), .Q(n13796) );
  OR2X1 U13777 ( .IN1(n10159), .IN2(n11548), .Q(n11825) );
  OR2X1 U13778 ( .IN1(n13797), .IN2(n13798), .Q(n11548) );
  OR2X1 U13779 ( .IN1(n13799), .IN2(n13800), .Q(n13798) );
  AND2X1 U13780 ( .IN1(n9798), .IN2(g165), .Q(n13800) );
  AND2X1 U13781 ( .IN1(n9800), .IN2(g6231), .Q(n13799) );
  AND2X1 U13782 ( .IN1(n9799), .IN2(g6313), .Q(n13797) );
  INVX0 U13783 ( .INP(n13091), .ZN(n13097) );
  AND2X1 U13784 ( .IN1(n13091), .IN2(n4282), .Q(n13794) );
  OR2X1 U13785 ( .IN1(n13801), .IN2(n13802), .Q(n13091) );
  OR2X1 U13786 ( .IN1(n13567), .IN2(n12036), .Q(n13802) );
  AND2X1 U13787 ( .IN1(n13803), .IN2(n13804), .Q(n13094) );
  INVX0 U13788 ( .INP(n13805), .ZN(n13804) );
  OR2X1 U13789 ( .IN1(n13806), .IN2(n13807), .Q(n13805) );
  AND2X1 U13790 ( .IN1(n9873), .IN2(n13375), .Q(n13807) );
  AND2X1 U13791 ( .IN1(n9874), .IN2(n13502), .Q(n13806) );
  OR2X1 U13792 ( .IN1(n4520), .IN2(test_so17), .Q(n13803) );
  AND2X1 U13793 ( .IN1(n13808), .IN2(n13809), .Q(g28668) );
  AND2X1 U13794 ( .IN1(n13810), .IN2(n13811), .Q(n13808) );
  INVX0 U13795 ( .INP(n13812), .ZN(n13811) );
  AND2X1 U13796 ( .IN1(n13813), .IN2(n4418), .Q(n13812) );
  OR2X1 U13797 ( .IN1(n4418), .IN2(n13813), .Q(n13810) );
  AND2X1 U13798 ( .IN1(n13814), .IN2(n12966), .Q(g28637) );
  AND2X1 U13799 ( .IN1(n13815), .IN2(n13816), .Q(n13814) );
  INVX0 U13800 ( .INP(n13817), .ZN(n13816) );
  AND2X1 U13801 ( .IN1(n1574), .IN2(n9876), .Q(n13817) );
  OR2X1 U13802 ( .IN1(n9876), .IN2(n1574), .Q(n13815) );
  AND2X1 U13803 ( .IN1(n13818), .IN2(n12971), .Q(g28636) );
  AND2X1 U13804 ( .IN1(n13819), .IN2(n13820), .Q(n13818) );
  INVX0 U13805 ( .INP(n13821), .ZN(n13820) );
  AND2X1 U13806 ( .IN1(n1230), .IN2(n9880), .Q(n13821) );
  OR2X1 U13807 ( .IN1(n9880), .IN2(n1230), .Q(n13819) );
  AND2X1 U13808 ( .IN1(n13822), .IN2(n12976), .Q(g28635) );
  AND2X1 U13809 ( .IN1(n13823), .IN2(n13824), .Q(n13822) );
  INVX0 U13810 ( .INP(n13825), .ZN(n13824) );
  AND2X1 U13811 ( .IN1(n885), .IN2(n9884), .Q(n13825) );
  OR2X1 U13812 ( .IN1(n9884), .IN2(n885), .Q(n13823) );
  AND2X1 U13813 ( .IN1(n13826), .IN2(n12981), .Q(g28634) );
  AND2X1 U13814 ( .IN1(n13827), .IN2(n13828), .Q(n13826) );
  INVX0 U13815 ( .INP(n13829), .ZN(n13828) );
  AND2X1 U13816 ( .IN1(n467), .IN2(n9888), .Q(n13829) );
  OR2X1 U13817 ( .IN1(n9888), .IN2(n467), .Q(n13827) );
  OR2X1 U13818 ( .IN1(n13830), .IN2(n13831), .Q(g28425) );
  AND2X1 U13819 ( .IN1(n578), .IN2(g3109), .Q(n13831) );
  AND2X1 U13820 ( .IN1(n4494), .IN2(g3102), .Q(n13830) );
  OR2X1 U13821 ( .IN1(n13832), .IN2(n13833), .Q(g28421) );
  AND2X1 U13822 ( .IN1(n578), .IN2(g8030), .Q(n13833) );
  AND2X1 U13823 ( .IN1(n4383), .IN2(test_so7), .Q(n13832) );
  OR2X1 U13824 ( .IN1(n13834), .IN2(n13835), .Q(g28420) );
  AND2X1 U13825 ( .IN1(n578), .IN2(g8106), .Q(n13835) );
  INVX0 U13826 ( .INP(n12912), .ZN(n578) );
  OR2X1 U13827 ( .IN1(n13836), .IN2(n13837), .Q(n12912) );
  AND2X1 U13828 ( .IN1(n13838), .IN2(n4548), .Q(n13837) );
  AND2X1 U13829 ( .IN1(n13839), .IN2(n13840), .Q(n13838) );
  INVX0 U13830 ( .INP(n13841), .ZN(n13840) );
  AND2X1 U13831 ( .IN1(g21851), .IN2(g6750), .Q(n13841) );
  OR2X1 U13832 ( .IN1(n9339), .IN2(n13842), .Q(n13839) );
  AND2X1 U13833 ( .IN1(n9338), .IN2(g1186), .Q(n13836) );
  AND2X1 U13834 ( .IN1(n4382), .IN2(g3100), .Q(n13834) );
  OR2X1 U13835 ( .IN1(n13843), .IN2(n13844), .Q(g28371) );
  AND2X1 U13836 ( .IN1(n13845), .IN2(g2624), .Q(n13844) );
  AND2X1 U13837 ( .IN1(n4299), .IN2(g2694), .Q(n13843) );
  OR2X1 U13838 ( .IN1(n13846), .IN2(n13847), .Q(g28368) );
  AND2X1 U13839 ( .IN1(n13845), .IN2(g7390), .Q(n13847) );
  AND2X1 U13840 ( .IN1(n4370), .IN2(g2691), .Q(n13846) );
  OR2X1 U13841 ( .IN1(n13848), .IN2(n13849), .Q(g28367) );
  AND2X1 U13842 ( .IN1(n13850), .IN2(g2624), .Q(n13849) );
  AND2X1 U13843 ( .IN1(n4299), .IN2(g2685), .Q(n13848) );
  OR2X1 U13844 ( .IN1(n13851), .IN2(n13852), .Q(g28366) );
  AND2X1 U13845 ( .IN1(n13853), .IN2(g1930), .Q(n13852) );
  AND2X1 U13846 ( .IN1(n4366), .IN2(g2000), .Q(n13851) );
  OR2X1 U13847 ( .IN1(n13854), .IN2(n13855), .Q(g28364) );
  AND2X1 U13848 ( .IN1(n13845), .IN2(n12862), .Q(n13855) );
  OR2X1 U13849 ( .IN1(n13856), .IN2(n13857), .Q(n13845) );
  AND2X1 U13850 ( .IN1(n11146), .IN2(n13858), .Q(n13857) );
  AND2X1 U13851 ( .IN1(n3252), .IN2(n13859), .Q(n13856) );
  AND2X1 U13852 ( .IN1(n4314), .IN2(g2688), .Q(n13854) );
  OR2X1 U13853 ( .IN1(n13860), .IN2(n13861), .Q(g28363) );
  AND2X1 U13854 ( .IN1(n13850), .IN2(g7390), .Q(n13861) );
  AND2X1 U13855 ( .IN1(n4370), .IN2(test_so90), .Q(n13860) );
  OR2X1 U13856 ( .IN1(n13862), .IN2(n13863), .Q(g28362) );
  AND2X1 U13857 ( .IN1(n13853), .IN2(g7194), .Q(n13863) );
  AND2X1 U13858 ( .IN1(n4315), .IN2(g1997), .Q(n13862) );
  OR2X1 U13859 ( .IN1(n13864), .IN2(n13865), .Q(g28361) );
  AND2X1 U13860 ( .IN1(n13866), .IN2(g1930), .Q(n13865) );
  AND2X1 U13861 ( .IN1(n4366), .IN2(g1991), .Q(n13864) );
  OR2X1 U13862 ( .IN1(n13867), .IN2(n13868), .Q(g28360) );
  AND2X1 U13863 ( .IN1(n13869), .IN2(g1236), .Q(n13868) );
  AND2X1 U13864 ( .IN1(n4300), .IN2(g1306), .Q(n13867) );
  OR2X1 U13865 ( .IN1(n13870), .IN2(n13871), .Q(g28358) );
  AND2X1 U13866 ( .IN1(n4314), .IN2(g2679), .Q(n13871) );
  AND2X1 U13867 ( .IN1(g7302), .IN2(n13850), .Q(n13870) );
  OR2X1 U13868 ( .IN1(n13872), .IN2(n13873), .Q(n13850) );
  AND2X1 U13869 ( .IN1(n11136), .IN2(n13858), .Q(n13873) );
  AND2X1 U13870 ( .IN1(n3260), .IN2(n11556), .Q(n13872) );
  INVX0 U13871 ( .INP(n13874), .ZN(n11556) );
  OR2X1 U13872 ( .IN1(n13875), .IN2(n13876), .Q(n13874) );
  OR2X1 U13873 ( .IN1(n13877), .IN2(n13878), .Q(n13876) );
  AND2X1 U13874 ( .IN1(n13879), .IN2(n13880), .Q(n13878) );
  AND2X1 U13875 ( .IN1(n13881), .IN2(n13882), .Q(n13879) );
  OR2X1 U13876 ( .IN1(n13883), .IN2(n13884), .Q(n13881) );
  AND2X1 U13877 ( .IN1(n13885), .IN2(n13886), .Q(n13883) );
  OR2X1 U13878 ( .IN1(n13887), .IN2(n13888), .Q(n13886) );
  AND2X1 U13879 ( .IN1(n13889), .IN2(n13890), .Q(n13877) );
  OR2X1 U13880 ( .IN1(n13891), .IN2(n13892), .Q(n13890) );
  AND2X1 U13881 ( .IN1(n13893), .IN2(n13894), .Q(n13892) );
  OR2X1 U13882 ( .IN1(n13895), .IN2(n13885), .Q(n13893) );
  AND2X1 U13883 ( .IN1(n13896), .IN2(n13897), .Q(n13895) );
  AND2X1 U13884 ( .IN1(n13898), .IN2(n13899), .Q(n13891) );
  AND2X1 U13885 ( .IN1(n13887), .IN2(n13888), .Q(n13899) );
  AND2X1 U13886 ( .IN1(n13885), .IN2(n13900), .Q(n13898) );
  OR2X1 U13887 ( .IN1(n13901), .IN2(n13902), .Q(n13875) );
  AND2X1 U13888 ( .IN1(n13903), .IN2(n13897), .Q(n13902) );
  AND2X1 U13889 ( .IN1(n13904), .IN2(n13905), .Q(n13903) );
  OR2X1 U13890 ( .IN1(n13906), .IN2(n13907), .Q(n13905) );
  AND2X1 U13891 ( .IN1(n13908), .IN2(n13909), .Q(n13906) );
  AND2X1 U13892 ( .IN1(n13910), .IN2(n13911), .Q(n13901) );
  OR2X1 U13893 ( .IN1(n13912), .IN2(n13913), .Q(n13911) );
  AND2X1 U13894 ( .IN1(n13914), .IN2(n13908), .Q(n13913) );
  OR2X1 U13895 ( .IN1(n13915), .IN2(n13916), .Q(n13908) );
  AND2X1 U13896 ( .IN1(n13917), .IN2(n13880), .Q(n13915) );
  AND2X1 U13897 ( .IN1(n13918), .IN2(n13907), .Q(n13912) );
  OR2X1 U13898 ( .IN1(n13919), .IN2(n13920), .Q(n13907) );
  AND2X1 U13899 ( .IN1(n13916), .IN2(n13880), .Q(n13920) );
  AND2X1 U13900 ( .IN1(n13900), .IN2(n13889), .Q(n13919) );
  INVX0 U13901 ( .INP(n13921), .ZN(n3260) );
  OR2X1 U13902 ( .IN1(n13858), .IN2(n13922), .Q(n13921) );
  OR2X1 U13903 ( .IN1(n11553), .IN2(n13923), .Q(n13922) );
  AND2X1 U13904 ( .IN1(n1636), .IN2(n13924), .Q(n13923) );
  INVX0 U13905 ( .INP(n13925), .ZN(n13924) );
  INVX0 U13906 ( .INP(n13926), .ZN(n1636) );
  OR2X1 U13907 ( .IN1(n13927), .IN2(n13928), .Q(n13926) );
  OR2X1 U13908 ( .IN1(n13929), .IN2(n13930), .Q(n13928) );
  AND2X1 U13909 ( .IN1(n13931), .IN2(n13880), .Q(n13930) );
  OR2X1 U13910 ( .IN1(n13932), .IN2(n13933), .Q(n13931) );
  AND2X1 U13911 ( .IN1(n13910), .IN2(n13934), .Q(n13933) );
  OR2X1 U13912 ( .IN1(n13935), .IN2(n13936), .Q(n13934) );
  OR2X1 U13913 ( .IN1(n13937), .IN2(n13938), .Q(n13936) );
  AND2X1 U13914 ( .IN1(n13884), .IN2(n13900), .Q(n13938) );
  AND2X1 U13915 ( .IN1(n13887), .IN2(n13939), .Q(n13884) );
  AND2X1 U13916 ( .IN1(n13888), .IN2(n13896), .Q(n13939) );
  AND2X1 U13917 ( .IN1(n13940), .IN2(n13885), .Q(n13937) );
  AND2X1 U13918 ( .IN1(n13904), .IN2(n13916), .Q(n13935) );
  AND2X1 U13919 ( .IN1(n13918), .IN2(n13894), .Q(n13932) );
  AND2X1 U13920 ( .IN1(n13941), .IN2(n13904), .Q(n13929) );
  INVX0 U13921 ( .INP(n13888), .ZN(n13904) );
  AND2X1 U13922 ( .IN1(n13942), .IN2(n13882), .Q(n13941) );
  OR2X1 U13923 ( .IN1(n13943), .IN2(n13944), .Q(n13942) );
  AND2X1 U13924 ( .IN1(n13910), .IN2(n13909), .Q(n13944) );
  AND2X1 U13925 ( .IN1(n13889), .IN2(n13887), .Q(n13943) );
  AND2X1 U13926 ( .IN1(n13945), .IN2(n13897), .Q(n13927) );
  OR2X1 U13927 ( .IN1(n13946), .IN2(n13947), .Q(n13945) );
  AND2X1 U13928 ( .IN1(n13889), .IN2(n13948), .Q(n13947) );
  OR2X1 U13929 ( .IN1(n13949), .IN2(n13950), .Q(n13948) );
  OR2X1 U13930 ( .IN1(n13951), .IN2(n13952), .Q(n13950) );
  AND2X1 U13931 ( .IN1(n13940), .IN2(n13918), .Q(n13952) );
  AND2X1 U13932 ( .IN1(n13888), .IN2(n13909), .Q(n13918) );
  AND2X1 U13933 ( .IN1(n13953), .IN2(n13896), .Q(n13951) );
  AND2X1 U13934 ( .IN1(n13916), .IN2(n13888), .Q(n13953) );
  OR2X1 U13935 ( .IN1(n13954), .IN2(n13955), .Q(n13888) );
  OR2X1 U13936 ( .IN1(n13956), .IN2(n13957), .Q(n13955) );
  AND2X1 U13937 ( .IN1(g2412), .IN2(g2443), .Q(n13957) );
  AND2X1 U13938 ( .IN1(g5747), .IN2(g2439), .Q(n13956) );
  AND2X1 U13939 ( .IN1(g5796), .IN2(g2441), .Q(n13954) );
  AND2X1 U13940 ( .IN1(n13885), .IN2(n13882), .Q(n13949) );
  INVX0 U13941 ( .INP(n13909), .ZN(n13885) );
  OR2X1 U13942 ( .IN1(n13958), .IN2(n13959), .Q(n13909) );
  OR2X1 U13943 ( .IN1(n13960), .IN2(n13961), .Q(n13959) );
  AND2X1 U13944 ( .IN1(g2412), .IN2(g2458), .Q(n13961) );
  AND2X1 U13945 ( .IN1(g5747), .IN2(g2454), .Q(n13960) );
  AND2X1 U13946 ( .IN1(g5796), .IN2(g2456), .Q(n13958) );
  INVX0 U13947 ( .INP(n13880), .ZN(n13889) );
  OR2X1 U13948 ( .IN1(n13962), .IN2(n13963), .Q(n13880) );
  OR2X1 U13949 ( .IN1(n13964), .IN2(n13965), .Q(n13963) );
  AND2X1 U13950 ( .IN1(g2412), .IN2(g2428), .Q(n13965) );
  AND2X1 U13951 ( .IN1(g5747), .IN2(g2424), .Q(n13964) );
  AND2X1 U13952 ( .IN1(g5796), .IN2(g2426), .Q(n13962) );
  AND2X1 U13953 ( .IN1(n13966), .IN2(n13914), .Q(n13946) );
  INVX0 U13954 ( .INP(n13896), .ZN(n13914) );
  OR2X1 U13955 ( .IN1(n13967), .IN2(n13968), .Q(n13896) );
  OR2X1 U13956 ( .IN1(n13969), .IN2(n13970), .Q(n13968) );
  AND2X1 U13957 ( .IN1(test_so85), .IN2(g2412), .Q(n13970) );
  AND2X1 U13958 ( .IN1(g5747), .IN2(g2469), .Q(n13969) );
  AND2X1 U13959 ( .IN1(g5796), .IN2(g2471), .Q(n13967) );
  AND2X1 U13960 ( .IN1(n13900), .IN2(n13887), .Q(n13966) );
  AND2X1 U13961 ( .IN1(n11557), .IN2(n13925), .Q(n11553) );
  OR2X1 U13962 ( .IN1(n13971), .IN2(n13972), .Q(g28357) );
  AND2X1 U13963 ( .IN1(n13853), .IN2(n13973), .Q(n13972) );
  OR2X1 U13964 ( .IN1(n13974), .IN2(n13975), .Q(n13853) );
  AND2X1 U13965 ( .IN1(n11309), .IN2(n13858), .Q(n13975) );
  AND2X1 U13966 ( .IN1(n3293), .IN2(n13976), .Q(n13974) );
  INVX0 U13967 ( .INP(n13977), .ZN(n3293) );
  OR2X1 U13968 ( .IN1(n13858), .IN2(n13978), .Q(n13977) );
  OR2X1 U13969 ( .IN1(n13979), .IN2(n13980), .Q(n13978) );
  AND2X1 U13970 ( .IN1(n13981), .IN2(n13982), .Q(n13980) );
  INVX0 U13971 ( .INP(n13983), .ZN(n13981) );
  AND2X1 U13972 ( .IN1(n4296), .IN2(g1994), .Q(n13971) );
  OR2X1 U13973 ( .IN1(n13984), .IN2(n13985), .Q(g28356) );
  AND2X1 U13974 ( .IN1(n13866), .IN2(g7194), .Q(n13985) );
  AND2X1 U13975 ( .IN1(n4315), .IN2(g1988), .Q(n13984) );
  OR2X1 U13976 ( .IN1(n13986), .IN2(n13987), .Q(g28355) );
  AND2X1 U13977 ( .IN1(n13869), .IN2(g6944), .Q(n13987) );
  AND2X1 U13978 ( .IN1(n4316), .IN2(g1303), .Q(n13986) );
  OR2X1 U13979 ( .IN1(n13988), .IN2(n13989), .Q(g28354) );
  AND2X1 U13980 ( .IN1(n13990), .IN2(g1236), .Q(n13989) );
  AND2X1 U13981 ( .IN1(n4300), .IN2(g1297), .Q(n13988) );
  OR2X1 U13982 ( .IN1(n13991), .IN2(n13992), .Q(g28353) );
  AND2X1 U13983 ( .IN1(n13993), .IN2(g550), .Q(n13992) );
  AND2X1 U13984 ( .IN1(n4313), .IN2(test_so26), .Q(n13991) );
  OR2X1 U13985 ( .IN1(n13994), .IN2(n13995), .Q(g28352) );
  AND2X1 U13986 ( .IN1(n4296), .IN2(g1985), .Q(n13995) );
  AND2X1 U13987 ( .IN1(g7052), .IN2(n13866), .Q(n13994) );
  OR2X1 U13988 ( .IN1(n13996), .IN2(n13997), .Q(n13866) );
  AND2X1 U13989 ( .IN1(n11299), .IN2(n13858), .Q(n13997) );
  AND2X1 U13990 ( .IN1(n342), .IN2(n13982), .Q(n13996) );
  INVX0 U13991 ( .INP(n13998), .ZN(n13982) );
  OR2X1 U13992 ( .IN1(n13999), .IN2(n14000), .Q(n13998) );
  OR2X1 U13993 ( .IN1(n14001), .IN2(n14002), .Q(n14000) );
  AND2X1 U13994 ( .IN1(n14003), .IN2(n14004), .Q(n14002) );
  AND2X1 U13995 ( .IN1(n14005), .IN2(n14006), .Q(n14003) );
  OR2X1 U13996 ( .IN1(n14007), .IN2(n14008), .Q(n14005) );
  AND2X1 U13997 ( .IN1(n14009), .IN2(n14010), .Q(n14007) );
  OR2X1 U13998 ( .IN1(n14011), .IN2(n14012), .Q(n14010) );
  AND2X1 U13999 ( .IN1(n14013), .IN2(n14014), .Q(n14001) );
  OR2X1 U14000 ( .IN1(n14015), .IN2(n14016), .Q(n14014) );
  AND2X1 U14001 ( .IN1(n14017), .IN2(n14018), .Q(n14016) );
  OR2X1 U14002 ( .IN1(n14019), .IN2(n14009), .Q(n14017) );
  AND2X1 U14003 ( .IN1(n14020), .IN2(n14021), .Q(n14019) );
  AND2X1 U14004 ( .IN1(n14022), .IN2(n14023), .Q(n14015) );
  AND2X1 U14005 ( .IN1(n14011), .IN2(n14012), .Q(n14023) );
  AND2X1 U14006 ( .IN1(n14009), .IN2(n14024), .Q(n14022) );
  OR2X1 U14007 ( .IN1(n14025), .IN2(n14026), .Q(n13999) );
  AND2X1 U14008 ( .IN1(n14027), .IN2(n14021), .Q(n14026) );
  AND2X1 U14009 ( .IN1(n14028), .IN2(n14029), .Q(n14027) );
  OR2X1 U14010 ( .IN1(n14030), .IN2(n14031), .Q(n14029) );
  AND2X1 U14011 ( .IN1(n14032), .IN2(n14033), .Q(n14030) );
  AND2X1 U14012 ( .IN1(n14034), .IN2(n14035), .Q(n14025) );
  OR2X1 U14013 ( .IN1(n14036), .IN2(n14037), .Q(n14035) );
  AND2X1 U14014 ( .IN1(n14038), .IN2(n14032), .Q(n14037) );
  OR2X1 U14015 ( .IN1(n14039), .IN2(n14040), .Q(n14032) );
  AND2X1 U14016 ( .IN1(n14041), .IN2(n14004), .Q(n14039) );
  AND2X1 U14017 ( .IN1(n14042), .IN2(n14031), .Q(n14036) );
  OR2X1 U14018 ( .IN1(n14043), .IN2(n14044), .Q(n14031) );
  AND2X1 U14019 ( .IN1(n14040), .IN2(n14004), .Q(n14044) );
  AND2X1 U14020 ( .IN1(n14024), .IN2(n14013), .Q(n14043) );
  INVX0 U14021 ( .INP(n14045), .ZN(n342) );
  OR2X1 U14022 ( .IN1(n13858), .IN2(n14046), .Q(n14045) );
  OR2X1 U14023 ( .IN1(n13979), .IN2(n14047), .Q(n14046) );
  AND2X1 U14024 ( .IN1(n14048), .IN2(n13976), .Q(n14047) );
  INVX0 U14025 ( .INP(n14049), .ZN(n13976) );
  OR2X1 U14026 ( .IN1(n14050), .IN2(n14051), .Q(n14049) );
  OR2X1 U14027 ( .IN1(n14052), .IN2(n14053), .Q(n14051) );
  AND2X1 U14028 ( .IN1(n14054), .IN2(n14004), .Q(n14053) );
  OR2X1 U14029 ( .IN1(n14055), .IN2(n14056), .Q(n14054) );
  AND2X1 U14030 ( .IN1(n14034), .IN2(n14057), .Q(n14056) );
  OR2X1 U14031 ( .IN1(n14058), .IN2(n14059), .Q(n14057) );
  OR2X1 U14032 ( .IN1(n14060), .IN2(n14061), .Q(n14059) );
  AND2X1 U14033 ( .IN1(n14008), .IN2(n14024), .Q(n14061) );
  AND2X1 U14034 ( .IN1(n14011), .IN2(n14062), .Q(n14008) );
  AND2X1 U14035 ( .IN1(n14012), .IN2(n14020), .Q(n14062) );
  AND2X1 U14036 ( .IN1(n14063), .IN2(n14009), .Q(n14060) );
  AND2X1 U14037 ( .IN1(n14028), .IN2(n14040), .Q(n14058) );
  AND2X1 U14038 ( .IN1(n14042), .IN2(n14018), .Q(n14055) );
  AND2X1 U14039 ( .IN1(n14064), .IN2(n14028), .Q(n14052) );
  INVX0 U14040 ( .INP(n14012), .ZN(n14028) );
  AND2X1 U14041 ( .IN1(n14065), .IN2(n14006), .Q(n14064) );
  OR2X1 U14042 ( .IN1(n14066), .IN2(n14067), .Q(n14065) );
  AND2X1 U14043 ( .IN1(n14034), .IN2(n14033), .Q(n14067) );
  AND2X1 U14044 ( .IN1(n14013), .IN2(n14011), .Q(n14066) );
  AND2X1 U14045 ( .IN1(n14068), .IN2(n14021), .Q(n14050) );
  OR2X1 U14046 ( .IN1(n14069), .IN2(n14070), .Q(n14068) );
  AND2X1 U14047 ( .IN1(n14013), .IN2(n14071), .Q(n14070) );
  OR2X1 U14048 ( .IN1(n14072), .IN2(n14073), .Q(n14071) );
  OR2X1 U14049 ( .IN1(n14074), .IN2(n14075), .Q(n14073) );
  AND2X1 U14050 ( .IN1(n14063), .IN2(n14042), .Q(n14075) );
  AND2X1 U14051 ( .IN1(n14012), .IN2(n14033), .Q(n14042) );
  AND2X1 U14052 ( .IN1(n14076), .IN2(n14020), .Q(n14074) );
  AND2X1 U14053 ( .IN1(n14040), .IN2(n14012), .Q(n14076) );
  OR2X1 U14054 ( .IN1(n14077), .IN2(n14078), .Q(n14012) );
  OR2X1 U14055 ( .IN1(n14079), .IN2(n14080), .Q(n14078) );
  AND2X1 U14056 ( .IN1(g5738), .IN2(g1747), .Q(n14080) );
  AND2X1 U14057 ( .IN1(g1718), .IN2(g1749), .Q(n14079) );
  AND2X1 U14058 ( .IN1(test_so63), .IN2(g1745), .Q(n14077) );
  AND2X1 U14059 ( .IN1(n14009), .IN2(n14006), .Q(n14072) );
  INVX0 U14060 ( .INP(n14033), .ZN(n14009) );
  OR2X1 U14061 ( .IN1(n14081), .IN2(n14082), .Q(n14033) );
  OR2X1 U14062 ( .IN1(n14083), .IN2(n14084), .Q(n14082) );
  AND2X1 U14063 ( .IN1(g5738), .IN2(g1762), .Q(n14084) );
  AND2X1 U14064 ( .IN1(g1718), .IN2(g1764), .Q(n14083) );
  AND2X1 U14065 ( .IN1(test_so63), .IN2(g1760), .Q(n14081) );
  INVX0 U14066 ( .INP(n14004), .ZN(n14013) );
  OR2X1 U14067 ( .IN1(n14085), .IN2(n14086), .Q(n14004) );
  OR2X1 U14068 ( .IN1(n14087), .IN2(n14088), .Q(n14086) );
  AND2X1 U14069 ( .IN1(g5738), .IN2(g1732), .Q(n14088) );
  AND2X1 U14070 ( .IN1(g1718), .IN2(g1734), .Q(n14087) );
  AND2X1 U14071 ( .IN1(test_so63), .IN2(g1730), .Q(n14085) );
  AND2X1 U14072 ( .IN1(n14089), .IN2(n14038), .Q(n14069) );
  INVX0 U14073 ( .INP(n14020), .ZN(n14038) );
  OR2X1 U14074 ( .IN1(n14090), .IN2(n14091), .Q(n14020) );
  OR2X1 U14075 ( .IN1(n14092), .IN2(n14093), .Q(n14091) );
  AND2X1 U14076 ( .IN1(g5738), .IN2(g1777), .Q(n14093) );
  AND2X1 U14077 ( .IN1(g1718), .IN2(g1705), .Q(n14092) );
  AND2X1 U14078 ( .IN1(test_so63), .IN2(g1775), .Q(n14090) );
  AND2X1 U14079 ( .IN1(n14024), .IN2(n14011), .Q(n14089) );
  INVX0 U14080 ( .INP(n14094), .ZN(n14048) );
  AND2X1 U14081 ( .IN1(n13983), .IN2(n14094), .Q(n13979) );
  OR2X1 U14082 ( .IN1(n14095), .IN2(n14096), .Q(g28351) );
  AND2X1 U14083 ( .IN1(n13869), .IN2(n13842), .Q(n14096) );
  OR2X1 U14084 ( .IN1(n14097), .IN2(n14098), .Q(n13869) );
  AND2X1 U14085 ( .IN1(n11471), .IN2(n13858), .Q(n14098) );
  AND2X1 U14086 ( .IN1(n3334), .IN2(n14099), .Q(n14097) );
  INVX0 U14087 ( .INP(n14100), .ZN(n3334) );
  OR2X1 U14088 ( .IN1(n13858), .IN2(n14101), .Q(n14100) );
  OR2X1 U14089 ( .IN1(n14102), .IN2(n14103), .Q(n14101) );
  AND2X1 U14090 ( .IN1(n14104), .IN2(n14105), .Q(n14103) );
  INVX0 U14091 ( .INP(n14106), .ZN(n14104) );
  AND2X1 U14092 ( .IN1(n4371), .IN2(g1300), .Q(n14095) );
  OR2X1 U14093 ( .IN1(n14107), .IN2(n14108), .Q(g28350) );
  AND2X1 U14094 ( .IN1(n13990), .IN2(g6944), .Q(n14108) );
  AND2X1 U14095 ( .IN1(n4316), .IN2(g1294), .Q(n14107) );
  OR2X1 U14096 ( .IN1(n14109), .IN2(n14110), .Q(g28349) );
  AND2X1 U14097 ( .IN1(n13993), .IN2(g6642), .Q(n14110) );
  AND2X1 U14098 ( .IN1(n4372), .IN2(g617), .Q(n14109) );
  OR2X1 U14099 ( .IN1(n14111), .IN2(n14112), .Q(g28348) );
  AND2X1 U14100 ( .IN1(n14113), .IN2(g550), .Q(n14112) );
  AND2X1 U14101 ( .IN1(n4313), .IN2(g611), .Q(n14111) );
  OR2X1 U14102 ( .IN1(n14114), .IN2(n14115), .Q(g28346) );
  AND2X1 U14103 ( .IN1(n4371), .IN2(g1291), .Q(n14115) );
  AND2X1 U14104 ( .IN1(g6750), .IN2(n13990), .Q(n14114) );
  OR2X1 U14105 ( .IN1(n14116), .IN2(n14117), .Q(n13990) );
  AND2X1 U14106 ( .IN1(n11461), .IN2(n13858), .Q(n14117) );
  AND2X1 U14107 ( .IN1(n339), .IN2(n14105), .Q(n14116) );
  INVX0 U14108 ( .INP(n14118), .ZN(n14105) );
  OR2X1 U14109 ( .IN1(n14119), .IN2(n14120), .Q(n14118) );
  OR2X1 U14110 ( .IN1(n14121), .IN2(n14122), .Q(n14120) );
  AND2X1 U14111 ( .IN1(n14123), .IN2(n14124), .Q(n14122) );
  AND2X1 U14112 ( .IN1(n14125), .IN2(n14126), .Q(n14123) );
  OR2X1 U14113 ( .IN1(n14127), .IN2(n14128), .Q(n14125) );
  AND2X1 U14114 ( .IN1(n14129), .IN2(n14130), .Q(n14127) );
  OR2X1 U14115 ( .IN1(n14131), .IN2(n14132), .Q(n14130) );
  AND2X1 U14116 ( .IN1(n14133), .IN2(n14134), .Q(n14121) );
  OR2X1 U14117 ( .IN1(n14135), .IN2(n14136), .Q(n14134) );
  AND2X1 U14118 ( .IN1(n14137), .IN2(n14138), .Q(n14136) );
  OR2X1 U14119 ( .IN1(n14139), .IN2(n14129), .Q(n14137) );
  AND2X1 U14120 ( .IN1(n14140), .IN2(n14141), .Q(n14139) );
  AND2X1 U14121 ( .IN1(n14142), .IN2(n14143), .Q(n14135) );
  AND2X1 U14122 ( .IN1(n14131), .IN2(n14132), .Q(n14143) );
  AND2X1 U14123 ( .IN1(n14129), .IN2(n14144), .Q(n14142) );
  OR2X1 U14124 ( .IN1(n14145), .IN2(n14146), .Q(n14119) );
  AND2X1 U14125 ( .IN1(n14147), .IN2(n14141), .Q(n14146) );
  AND2X1 U14126 ( .IN1(n14148), .IN2(n14149), .Q(n14147) );
  OR2X1 U14127 ( .IN1(n14150), .IN2(n14151), .Q(n14149) );
  AND2X1 U14128 ( .IN1(n14152), .IN2(n14153), .Q(n14150) );
  AND2X1 U14129 ( .IN1(n14154), .IN2(n14155), .Q(n14145) );
  OR2X1 U14130 ( .IN1(n14156), .IN2(n14157), .Q(n14155) );
  AND2X1 U14131 ( .IN1(n14158), .IN2(n14152), .Q(n14157) );
  OR2X1 U14132 ( .IN1(n14159), .IN2(n14160), .Q(n14152) );
  AND2X1 U14133 ( .IN1(n14161), .IN2(n14124), .Q(n14159) );
  AND2X1 U14134 ( .IN1(n14162), .IN2(n14151), .Q(n14156) );
  OR2X1 U14135 ( .IN1(n14163), .IN2(n14164), .Q(n14151) );
  AND2X1 U14136 ( .IN1(n14160), .IN2(n14124), .Q(n14164) );
  AND2X1 U14137 ( .IN1(n14144), .IN2(n14133), .Q(n14163) );
  INVX0 U14138 ( .INP(n14165), .ZN(n339) );
  OR2X1 U14139 ( .IN1(n13858), .IN2(n14166), .Q(n14165) );
  OR2X1 U14140 ( .IN1(n14102), .IN2(n14167), .Q(n14166) );
  AND2X1 U14141 ( .IN1(n14168), .IN2(n14099), .Q(n14167) );
  INVX0 U14142 ( .INP(n14169), .ZN(n14099) );
  OR2X1 U14143 ( .IN1(n14170), .IN2(n14171), .Q(n14169) );
  OR2X1 U14144 ( .IN1(n14172), .IN2(n14173), .Q(n14171) );
  AND2X1 U14145 ( .IN1(n14174), .IN2(n14124), .Q(n14173) );
  OR2X1 U14146 ( .IN1(n14175), .IN2(n14176), .Q(n14174) );
  AND2X1 U14147 ( .IN1(n14154), .IN2(n14177), .Q(n14176) );
  OR2X1 U14148 ( .IN1(n14178), .IN2(n14179), .Q(n14177) );
  OR2X1 U14149 ( .IN1(n14180), .IN2(n14181), .Q(n14179) );
  AND2X1 U14150 ( .IN1(n14128), .IN2(n14144), .Q(n14181) );
  AND2X1 U14151 ( .IN1(n14131), .IN2(n14182), .Q(n14128) );
  AND2X1 U14152 ( .IN1(n14132), .IN2(n14140), .Q(n14182) );
  AND2X1 U14153 ( .IN1(n14183), .IN2(n14129), .Q(n14180) );
  AND2X1 U14154 ( .IN1(n14148), .IN2(n14160), .Q(n14178) );
  AND2X1 U14155 ( .IN1(n14162), .IN2(n14138), .Q(n14175) );
  AND2X1 U14156 ( .IN1(n14184), .IN2(n14148), .Q(n14172) );
  INVX0 U14157 ( .INP(n14132), .ZN(n14148) );
  AND2X1 U14158 ( .IN1(n14185), .IN2(n14126), .Q(n14184) );
  OR2X1 U14159 ( .IN1(n14186), .IN2(n14187), .Q(n14185) );
  AND2X1 U14160 ( .IN1(n14154), .IN2(n14153), .Q(n14187) );
  AND2X1 U14161 ( .IN1(n14133), .IN2(n14131), .Q(n14186) );
  AND2X1 U14162 ( .IN1(n14188), .IN2(n14141), .Q(n14170) );
  OR2X1 U14163 ( .IN1(n14189), .IN2(n14190), .Q(n14188) );
  AND2X1 U14164 ( .IN1(n14133), .IN2(n14191), .Q(n14190) );
  OR2X1 U14165 ( .IN1(n14192), .IN2(n14193), .Q(n14191) );
  OR2X1 U14166 ( .IN1(n14194), .IN2(n14195), .Q(n14193) );
  AND2X1 U14167 ( .IN1(n14183), .IN2(n14162), .Q(n14195) );
  AND2X1 U14168 ( .IN1(n14132), .IN2(n14153), .Q(n14162) );
  AND2X1 U14169 ( .IN1(n14196), .IN2(n14140), .Q(n14194) );
  AND2X1 U14170 ( .IN1(n14160), .IN2(n14132), .Q(n14196) );
  OR2X1 U14171 ( .IN1(n14197), .IN2(n14198), .Q(n14132) );
  OR2X1 U14172 ( .IN1(n14199), .IN2(n14200), .Q(n14198) );
  AND2X1 U14173 ( .IN1(g1024), .IN2(g1055), .Q(n14200) );
  AND2X1 U14174 ( .IN1(g5657), .IN2(g1051), .Q(n14199) );
  AND2X1 U14175 ( .IN1(g5686), .IN2(g1053), .Q(n14197) );
  AND2X1 U14176 ( .IN1(n14129), .IN2(n14126), .Q(n14192) );
  INVX0 U14177 ( .INP(n14153), .ZN(n14129) );
  OR2X1 U14178 ( .IN1(n14201), .IN2(n14202), .Q(n14153) );
  OR2X1 U14179 ( .IN1(n14203), .IN2(n14204), .Q(n14202) );
  AND2X1 U14180 ( .IN1(g1024), .IN2(g1070), .Q(n14204) );
  AND2X1 U14181 ( .IN1(g5657), .IN2(g1066), .Q(n14203) );
  AND2X1 U14182 ( .IN1(g5686), .IN2(g1068), .Q(n14201) );
  INVX0 U14183 ( .INP(n14124), .ZN(n14133) );
  OR2X1 U14184 ( .IN1(n14205), .IN2(n14206), .Q(n14124) );
  OR2X1 U14185 ( .IN1(n14207), .IN2(n14208), .Q(n14206) );
  AND2X1 U14186 ( .IN1(g1024), .IN2(g1040), .Q(n14208) );
  AND2X1 U14187 ( .IN1(g5657), .IN2(g1036), .Q(n14207) );
  AND2X1 U14188 ( .IN1(g5686), .IN2(g1038), .Q(n14205) );
  AND2X1 U14189 ( .IN1(n14209), .IN2(n14158), .Q(n14189) );
  INVX0 U14190 ( .INP(n14140), .ZN(n14158) );
  OR2X1 U14191 ( .IN1(n14210), .IN2(n14211), .Q(n14140) );
  OR2X1 U14192 ( .IN1(n14212), .IN2(n14213), .Q(n14211) );
  AND2X1 U14193 ( .IN1(g1024), .IN2(g1011), .Q(n14213) );
  AND2X1 U14194 ( .IN1(g5657), .IN2(g1081), .Q(n14212) );
  AND2X1 U14195 ( .IN1(g5686), .IN2(g1083), .Q(n14210) );
  AND2X1 U14196 ( .IN1(n14144), .IN2(n14131), .Q(n14209) );
  INVX0 U14197 ( .INP(n14214), .ZN(n14168) );
  AND2X1 U14198 ( .IN1(n14106), .IN2(n14214), .Q(n14102) );
  OR2X1 U14199 ( .IN1(n14215), .IN2(n14216), .Q(g28345) );
  AND2X1 U14200 ( .IN1(n13993), .IN2(n11054), .Q(n14216) );
  OR2X1 U14201 ( .IN1(n14217), .IN2(n14218), .Q(n13993) );
  AND2X1 U14202 ( .IN1(n10961), .IN2(n13858), .Q(n14218) );
  AND2X1 U14203 ( .IN1(n3374), .IN2(n14219), .Q(n14217) );
  INVX0 U14204 ( .INP(n14220), .ZN(n3374) );
  OR2X1 U14205 ( .IN1(n13858), .IN2(n14221), .Q(n14220) );
  OR2X1 U14206 ( .IN1(n14222), .IN2(n14223), .Q(n14221) );
  AND2X1 U14207 ( .IN1(n14224), .IN2(n14225), .Q(n14223) );
  INVX0 U14208 ( .INP(n14226), .ZN(n14224) );
  AND2X1 U14209 ( .IN1(n4298), .IN2(g614), .Q(n14215) );
  OR2X1 U14210 ( .IN1(n14227), .IN2(n14228), .Q(g28344) );
  AND2X1 U14211 ( .IN1(n14113), .IN2(g6642), .Q(n14228) );
  AND2X1 U14212 ( .IN1(n4372), .IN2(g608), .Q(n14227) );
  OR2X1 U14213 ( .IN1(n14229), .IN2(n14230), .Q(g28342) );
  AND2X1 U14214 ( .IN1(n4298), .IN2(g605), .Q(n14230) );
  AND2X1 U14215 ( .IN1(g6485), .IN2(n14113), .Q(n14229) );
  OR2X1 U14216 ( .IN1(n14231), .IN2(n14232), .Q(n14113) );
  AND2X1 U14217 ( .IN1(n10967), .IN2(n13858), .Q(n14232) );
  AND2X1 U14218 ( .IN1(n336), .IN2(n14225), .Q(n14231) );
  INVX0 U14219 ( .INP(n14233), .ZN(n14225) );
  OR2X1 U14220 ( .IN1(n14234), .IN2(n14235), .Q(n14233) );
  OR2X1 U14221 ( .IN1(n14236), .IN2(n14237), .Q(n14235) );
  AND2X1 U14222 ( .IN1(n14238), .IN2(n14239), .Q(n14237) );
  AND2X1 U14223 ( .IN1(n14240), .IN2(n14241), .Q(n14238) );
  OR2X1 U14224 ( .IN1(n14242), .IN2(n14243), .Q(n14240) );
  AND2X1 U14225 ( .IN1(n14244), .IN2(n14245), .Q(n14242) );
  OR2X1 U14226 ( .IN1(n14246), .IN2(n14247), .Q(n14245) );
  AND2X1 U14227 ( .IN1(n14248), .IN2(n14249), .Q(n14236) );
  OR2X1 U14228 ( .IN1(n14250), .IN2(n14251), .Q(n14249) );
  AND2X1 U14229 ( .IN1(n14252), .IN2(n14253), .Q(n14251) );
  OR2X1 U14230 ( .IN1(n14254), .IN2(n14244), .Q(n14252) );
  AND2X1 U14231 ( .IN1(n14255), .IN2(n14256), .Q(n14254) );
  AND2X1 U14232 ( .IN1(n14257), .IN2(n14258), .Q(n14250) );
  AND2X1 U14233 ( .IN1(n14246), .IN2(n14247), .Q(n14258) );
  AND2X1 U14234 ( .IN1(n14244), .IN2(n14259), .Q(n14257) );
  OR2X1 U14235 ( .IN1(n14260), .IN2(n14261), .Q(n14234) );
  AND2X1 U14236 ( .IN1(n14262), .IN2(n14256), .Q(n14261) );
  AND2X1 U14237 ( .IN1(n14263), .IN2(n14264), .Q(n14262) );
  OR2X1 U14238 ( .IN1(n14265), .IN2(n14266), .Q(n14264) );
  AND2X1 U14239 ( .IN1(n14267), .IN2(n14268), .Q(n14265) );
  AND2X1 U14240 ( .IN1(n14269), .IN2(n14270), .Q(n14260) );
  OR2X1 U14241 ( .IN1(n14271), .IN2(n14272), .Q(n14270) );
  AND2X1 U14242 ( .IN1(n14273), .IN2(n14267), .Q(n14272) );
  OR2X1 U14243 ( .IN1(n14274), .IN2(n14275), .Q(n14267) );
  AND2X1 U14244 ( .IN1(n14276), .IN2(n14239), .Q(n14274) );
  AND2X1 U14245 ( .IN1(n14277), .IN2(n14266), .Q(n14271) );
  OR2X1 U14246 ( .IN1(n14278), .IN2(n14279), .Q(n14266) );
  AND2X1 U14247 ( .IN1(n14275), .IN2(n14239), .Q(n14279) );
  AND2X1 U14248 ( .IN1(n14259), .IN2(n14248), .Q(n14278) );
  INVX0 U14249 ( .INP(n14280), .ZN(n336) );
  OR2X1 U14250 ( .IN1(n13858), .IN2(n14281), .Q(n14280) );
  OR2X1 U14251 ( .IN1(n14222), .IN2(n14282), .Q(n14281) );
  AND2X1 U14252 ( .IN1(n14283), .IN2(n14219), .Q(n14282) );
  INVX0 U14253 ( .INP(n14284), .ZN(n14219) );
  OR2X1 U14254 ( .IN1(n14285), .IN2(n14286), .Q(n14284) );
  OR2X1 U14255 ( .IN1(n14287), .IN2(n14288), .Q(n14286) );
  AND2X1 U14256 ( .IN1(n14289), .IN2(n14239), .Q(n14288) );
  OR2X1 U14257 ( .IN1(n14290), .IN2(n14291), .Q(n14289) );
  AND2X1 U14258 ( .IN1(n14269), .IN2(n14292), .Q(n14291) );
  OR2X1 U14259 ( .IN1(n14293), .IN2(n14294), .Q(n14292) );
  OR2X1 U14260 ( .IN1(n14295), .IN2(n14296), .Q(n14294) );
  AND2X1 U14261 ( .IN1(n14243), .IN2(n14259), .Q(n14296) );
  AND2X1 U14262 ( .IN1(n14246), .IN2(n14297), .Q(n14243) );
  AND2X1 U14263 ( .IN1(n14247), .IN2(n14255), .Q(n14297) );
  AND2X1 U14264 ( .IN1(n14298), .IN2(n14244), .Q(n14295) );
  AND2X1 U14265 ( .IN1(n14263), .IN2(n14275), .Q(n14293) );
  AND2X1 U14266 ( .IN1(n14277), .IN2(n14253), .Q(n14290) );
  AND2X1 U14267 ( .IN1(n14299), .IN2(n14263), .Q(n14287) );
  INVX0 U14268 ( .INP(n14247), .ZN(n14263) );
  AND2X1 U14269 ( .IN1(n14300), .IN2(n14241), .Q(n14299) );
  OR2X1 U14270 ( .IN1(n14301), .IN2(n14302), .Q(n14300) );
  AND2X1 U14271 ( .IN1(n14269), .IN2(n14268), .Q(n14302) );
  AND2X1 U14272 ( .IN1(n14248), .IN2(n14246), .Q(n14301) );
  AND2X1 U14273 ( .IN1(n14303), .IN2(n14256), .Q(n14285) );
  OR2X1 U14274 ( .IN1(n14304), .IN2(n14305), .Q(n14303) );
  AND2X1 U14275 ( .IN1(n14248), .IN2(n14306), .Q(n14305) );
  OR2X1 U14276 ( .IN1(n14307), .IN2(n14308), .Q(n14306) );
  OR2X1 U14277 ( .IN1(n14309), .IN2(n14310), .Q(n14308) );
  AND2X1 U14278 ( .IN1(n14298), .IN2(n14277), .Q(n14310) );
  AND2X1 U14279 ( .IN1(n14247), .IN2(n14268), .Q(n14277) );
  AND2X1 U14280 ( .IN1(n14311), .IN2(n14255), .Q(n14309) );
  AND2X1 U14281 ( .IN1(n14275), .IN2(n14247), .Q(n14311) );
  OR2X1 U14282 ( .IN1(n14312), .IN2(n14313), .Q(n14247) );
  OR2X1 U14283 ( .IN1(n14314), .IN2(n14315), .Q(n14313) );
  AND2X1 U14284 ( .IN1(g337), .IN2(g368), .Q(n14315) );
  AND2X1 U14285 ( .IN1(g5629), .IN2(g364), .Q(n14314) );
  AND2X1 U14286 ( .IN1(g5648), .IN2(g366), .Q(n14312) );
  AND2X1 U14287 ( .IN1(n14244), .IN2(n14241), .Q(n14307) );
  INVX0 U14288 ( .INP(n14268), .ZN(n14244) );
  OR2X1 U14289 ( .IN1(n14316), .IN2(n14317), .Q(n14268) );
  OR2X1 U14290 ( .IN1(n14318), .IN2(n14319), .Q(n14317) );
  AND2X1 U14291 ( .IN1(g337), .IN2(g383), .Q(n14319) );
  AND2X1 U14292 ( .IN1(g5629), .IN2(g379), .Q(n14318) );
  AND2X1 U14293 ( .IN1(g5648), .IN2(g381), .Q(n14316) );
  INVX0 U14294 ( .INP(n14239), .ZN(n14248) );
  OR2X1 U14295 ( .IN1(n14320), .IN2(n14321), .Q(n14239) );
  OR2X1 U14296 ( .IN1(n14322), .IN2(n14323), .Q(n14321) );
  AND2X1 U14297 ( .IN1(g337), .IN2(g353), .Q(n14323) );
  AND2X1 U14298 ( .IN1(g5629), .IN2(g349), .Q(n14322) );
  AND2X1 U14299 ( .IN1(g5648), .IN2(g351), .Q(n14320) );
  AND2X1 U14300 ( .IN1(n14324), .IN2(n14273), .Q(n14304) );
  INVX0 U14301 ( .INP(n14255), .ZN(n14273) );
  OR2X1 U14302 ( .IN1(n14325), .IN2(n14326), .Q(n14255) );
  OR2X1 U14303 ( .IN1(n14327), .IN2(n14328), .Q(n14326) );
  AND2X1 U14304 ( .IN1(g337), .IN2(g324), .Q(n14328) );
  AND2X1 U14305 ( .IN1(g5629), .IN2(g394), .Q(n14327) );
  AND2X1 U14306 ( .IN1(g5648), .IN2(g396), .Q(n14325) );
  AND2X1 U14307 ( .IN1(n14259), .IN2(n14246), .Q(n14324) );
  INVX0 U14308 ( .INP(n14329), .ZN(n14283) );
  AND2X1 U14309 ( .IN1(n14226), .IN2(n14329), .Q(n14222) );
  AND2X1 U14310 ( .IN1(n14330), .IN2(n14331), .Q(g28328) );
  AND2X1 U14311 ( .IN1(n14332), .IN2(n14333), .Q(n14330) );
  INVX0 U14312 ( .INP(n14334), .ZN(n14333) );
  AND2X1 U14313 ( .IN1(n14335), .IN2(n4415), .Q(n14334) );
  OR2X1 U14314 ( .IN1(n4415), .IN2(n14335), .Q(n14332) );
  AND2X1 U14315 ( .IN1(n14336), .IN2(n14337), .Q(g28325) );
  AND2X1 U14316 ( .IN1(n14338), .IN2(n14339), .Q(n14336) );
  OR2X1 U14317 ( .IN1(n14340), .IN2(g2072), .Q(n14339) );
  AND2X1 U14318 ( .IN1(test_so70), .IN2(n14341), .Q(n14340) );
  OR2X1 U14319 ( .IN1(n4416), .IN2(n14342), .Q(n14338) );
  OR2X1 U14320 ( .IN1(n14343), .IN2(n10194), .Q(n14342) );
  AND2X1 U14321 ( .IN1(n14344), .IN2(n14345), .Q(g28321) );
  AND2X1 U14322 ( .IN1(n14346), .IN2(n14347), .Q(n14344) );
  OR2X1 U14323 ( .IN1(n14348), .IN2(g1378), .Q(n14347) );
  AND2X1 U14324 ( .IN1(n14349), .IN2(g1372), .Q(n14348) );
  OR2X1 U14325 ( .IN1(n4417), .IN2(n14350), .Q(n14346) );
  AND2X1 U14326 ( .IN1(n14351), .IN2(n13809), .Q(g28199) );
  AND2X1 U14327 ( .IN1(n13813), .IN2(n14352), .Q(n14351) );
  INVX0 U14328 ( .INP(n14353), .ZN(n14352) );
  AND2X1 U14329 ( .IN1(n14354), .IN2(n4396), .Q(n14353) );
  OR2X1 U14330 ( .IN1(n4396), .IN2(n14354), .Q(n13813) );
  AND2X1 U14331 ( .IN1(n14355), .IN2(n12966), .Q(g28148) );
  AND2X1 U14332 ( .IN1(n14356), .IN2(n1574), .Q(n14355) );
  OR2X1 U14333 ( .IN1(n10169), .IN2(n14357), .Q(n1574) );
  INVX0 U14334 ( .INP(n3424), .ZN(n14357) );
  OR2X1 U14335 ( .IN1(n3424), .IN2(g2138), .Q(n14356) );
  AND2X1 U14336 ( .IN1(n14358), .IN2(n12971), .Q(g28147) );
  AND2X1 U14337 ( .IN1(n14359), .IN2(n1230), .Q(n14358) );
  OR2X1 U14338 ( .IN1(n10168), .IN2(n14360), .Q(n1230) );
  INVX0 U14339 ( .INP(n3427), .ZN(n14360) );
  OR2X1 U14340 ( .IN1(n3427), .IN2(g1444), .Q(n14359) );
  AND2X1 U14341 ( .IN1(n14361), .IN2(n12976), .Q(g28146) );
  AND2X1 U14342 ( .IN1(n14362), .IN2(n885), .Q(n14361) );
  OR2X1 U14343 ( .IN1(n10170), .IN2(n14363), .Q(n885) );
  INVX0 U14344 ( .INP(n3430), .ZN(n14363) );
  OR2X1 U14345 ( .IN1(n3430), .IN2(g758), .Q(n14362) );
  AND2X1 U14346 ( .IN1(n14364), .IN2(n12981), .Q(g28145) );
  AND2X1 U14347 ( .IN1(n14365), .IN2(n467), .Q(n14364) );
  OR2X1 U14348 ( .IN1(n10167), .IN2(n14366), .Q(n467) );
  INVX0 U14349 ( .INP(n3433), .ZN(n14366) );
  OR2X1 U14350 ( .IN1(n3433), .IN2(g70), .Q(n14365) );
  OR2X1 U14351 ( .IN1(n14367), .IN2(n14368), .Q(g27771) );
  AND2X1 U14352 ( .IN1(n14369), .IN2(n13101), .Q(n14368) );
  AND2X1 U14353 ( .IN1(test_so81), .IN2(n14370), .Q(n14367) );
  OR2X1 U14354 ( .IN1(n4509), .IN2(n14371), .Q(n14370) );
  OR2X1 U14355 ( .IN1(n14372), .IN2(n14373), .Q(g27769) );
  AND2X1 U14356 ( .IN1(n14369), .IN2(n13106), .Q(n14373) );
  AND2X1 U14357 ( .IN1(n14374), .IN2(g2524), .Q(n14372) );
  OR2X1 U14358 ( .IN1(n4524), .IN2(n14371), .Q(n14374) );
  OR2X1 U14359 ( .IN1(n14375), .IN2(n14376), .Q(g27768) );
  AND2X1 U14360 ( .IN1(n14377), .IN2(n13111), .Q(n14376) );
  AND2X1 U14361 ( .IN1(n14378), .IN2(g1828), .Q(n14375) );
  OR2X1 U14362 ( .IN1(n4511), .IN2(n14379), .Q(n14378) );
  OR2X1 U14363 ( .IN1(n14380), .IN2(n14381), .Q(g27767) );
  AND2X1 U14364 ( .IN1(n14369), .IN2(n13116), .Q(n14381) );
  INVX0 U14365 ( .INP(n14382), .ZN(n14369) );
  OR2X1 U14366 ( .IN1(n10191), .IN2(n14383), .Q(n14382) );
  OR2X1 U14367 ( .IN1(n14384), .IN2(n14385), .Q(n14383) );
  AND2X1 U14368 ( .IN1(n14386), .IN2(n14387), .Q(n14385) );
  AND2X1 U14369 ( .IN1(n14388), .IN2(n14389), .Q(n14384) );
  AND2X1 U14370 ( .IN1(n14390), .IN2(g2523), .Q(n14380) );
  OR2X1 U14371 ( .IN1(n4516), .IN2(n14371), .Q(n14390) );
  OR2X1 U14372 ( .IN1(n14391), .IN2(n14392), .Q(n14371) );
  OR2X1 U14373 ( .IN1(n14393), .IN2(n14394), .Q(g27766) );
  AND2X1 U14374 ( .IN1(n14377), .IN2(n13239), .Q(n14394) );
  AND2X1 U14375 ( .IN1(n14395), .IN2(g1830), .Q(n14393) );
  OR2X1 U14376 ( .IN1(n4525), .IN2(n14379), .Q(n14395) );
  OR2X1 U14377 ( .IN1(n14396), .IN2(n14397), .Q(g27765) );
  AND2X1 U14378 ( .IN1(n14398), .IN2(g1088), .Q(n14397) );
  AND2X1 U14379 ( .IN1(n14399), .IN2(g1134), .Q(n14396) );
  OR2X1 U14380 ( .IN1(n4381), .IN2(n14400), .Q(n14399) );
  OR2X1 U14381 ( .IN1(n14401), .IN2(n14402), .Q(g27764) );
  AND2X1 U14382 ( .IN1(n14377), .IN2(n13248), .Q(n14402) );
  INVX0 U14383 ( .INP(n14403), .ZN(n14377) );
  OR2X1 U14384 ( .IN1(n4386), .IN2(n14404), .Q(n14403) );
  OR2X1 U14385 ( .IN1(n14405), .IN2(n14406), .Q(n14404) );
  AND2X1 U14386 ( .IN1(n14407), .IN2(n14408), .Q(n14406) );
  AND2X1 U14387 ( .IN1(n14409), .IN2(n14410), .Q(n14405) );
  AND2X1 U14388 ( .IN1(n14411), .IN2(g1829), .Q(n14401) );
  OR2X1 U14389 ( .IN1(n4518), .IN2(n14379), .Q(n14411) );
  OR2X1 U14390 ( .IN1(n14412), .IN2(n14413), .Q(n14379) );
  OR2X1 U14391 ( .IN1(n14414), .IN2(n14415), .Q(g27763) );
  AND2X1 U14392 ( .IN1(n14398), .IN2(g6712), .Q(n14415) );
  AND2X1 U14393 ( .IN1(n14416), .IN2(g1136), .Q(n14414) );
  OR2X1 U14394 ( .IN1(n4364), .IN2(n14400), .Q(n14416) );
  OR2X1 U14395 ( .IN1(n14417), .IN2(n14418), .Q(g27762) );
  AND2X1 U14396 ( .IN1(n14419), .IN2(n13375), .Q(n14418) );
  AND2X1 U14397 ( .IN1(n14420), .IN2(g447), .Q(n14417) );
  OR2X1 U14398 ( .IN1(n4506), .IN2(n14421), .Q(n14420) );
  OR2X1 U14399 ( .IN1(n14422), .IN2(n14423), .Q(g27761) );
  AND2X1 U14400 ( .IN1(n14398), .IN2(g5472), .Q(n14423) );
  INVX0 U14401 ( .INP(n14424), .ZN(n14398) );
  OR2X1 U14402 ( .IN1(n4387), .IN2(n14425), .Q(n14424) );
  OR2X1 U14403 ( .IN1(n14426), .IN2(n14427), .Q(n14425) );
  AND2X1 U14404 ( .IN1(n14428), .IN2(n14429), .Q(n14427) );
  AND2X1 U14405 ( .IN1(n14430), .IN2(n14431), .Q(n14426) );
  AND2X1 U14406 ( .IN1(n14432), .IN2(g1135), .Q(n14422) );
  OR2X1 U14407 ( .IN1(n4363), .IN2(n14400), .Q(n14432) );
  OR2X1 U14408 ( .IN1(n14433), .IN2(n14434), .Q(n14400) );
  OR2X1 U14409 ( .IN1(n14435), .IN2(n14436), .Q(g27760) );
  AND2X1 U14410 ( .IN1(n14419), .IN2(n13502), .Q(n14436) );
  AND2X1 U14411 ( .IN1(n14437), .IN2(g449), .Q(n14435) );
  OR2X1 U14412 ( .IN1(n4499), .IN2(n14421), .Q(n14437) );
  OR2X1 U14413 ( .IN1(n14438), .IN2(n14439), .Q(g27759) );
  AND2X1 U14414 ( .IN1(n14419), .IN2(n13506), .Q(n14439) );
  INVX0 U14415 ( .INP(n14440), .ZN(n14419) );
  OR2X1 U14416 ( .IN1(n4388), .IN2(n14441), .Q(n14440) );
  OR2X1 U14417 ( .IN1(n14442), .IN2(n14443), .Q(n14441) );
  AND2X1 U14418 ( .IN1(n14444), .IN2(n14445), .Q(n14443) );
  AND2X1 U14419 ( .IN1(n14446), .IN2(n14447), .Q(n14442) );
  AND2X1 U14420 ( .IN1(n14448), .IN2(g448), .Q(n14438) );
  OR2X1 U14421 ( .IN1(n4520), .IN2(n14421), .Q(n14448) );
  OR2X1 U14422 ( .IN1(n14449), .IN2(n14450), .Q(n14421) );
  AND2X1 U14423 ( .IN1(n14451), .IN2(n14331), .Q(g27724) );
  AND2X1 U14424 ( .IN1(n14335), .IN2(n14452), .Q(n14451) );
  INVX0 U14425 ( .INP(n14453), .ZN(n14452) );
  AND2X1 U14426 ( .IN1(n14454), .IN2(n4393), .Q(n14453) );
  OR2X1 U14427 ( .IN1(n4393), .IN2(n14454), .Q(n14335) );
  AND2X1 U14428 ( .IN1(n14455), .IN2(n14337), .Q(g27722) );
  OR2X1 U14429 ( .IN1(n14456), .IN2(n14457), .Q(n14455) );
  AND2X1 U14430 ( .IN1(n14341), .IN2(n10194), .Q(n14457) );
  INVX0 U14431 ( .INP(n14343), .ZN(n14341) );
  AND2X1 U14432 ( .IN1(test_so70), .IN2(n14343), .Q(n14456) );
  AND2X1 U14433 ( .IN1(n14458), .IN2(n14345), .Q(g27718) );
  AND2X1 U14434 ( .IN1(n14350), .IN2(n14459), .Q(n14458) );
  OR2X1 U14435 ( .IN1(n14349), .IN2(g1372), .Q(n14459) );
  INVX0 U14436 ( .INP(n14460), .ZN(n14349) );
  OR2X1 U14437 ( .IN1(n4395), .IN2(n14460), .Q(n14350) );
  AND2X1 U14438 ( .IN1(n14461), .IN2(n14462), .Q(g27682) );
  OR2X1 U14439 ( .IN1(n14463), .IN2(g2059), .Q(n14462) );
  AND2X1 U14440 ( .IN1(n14464), .IN2(g2046), .Q(n14463) );
  AND2X1 U14441 ( .IN1(n14337), .IN2(n14343), .Q(n14461) );
  OR2X1 U14442 ( .IN1(n14465), .IN2(n14466), .Q(n14343) );
  OR2X1 U14443 ( .IN1(n4473), .IN2(n4468), .Q(n14466) );
  AND2X1 U14444 ( .IN1(n14467), .IN2(n14468), .Q(g27678) );
  OR2X1 U14445 ( .IN1(n14469), .IN2(g1365), .Q(n14468) );
  AND2X1 U14446 ( .IN1(n14470), .IN2(g1352), .Q(n14469) );
  AND2X1 U14447 ( .IN1(n14345), .IN2(n14460), .Q(n14467) );
  OR2X1 U14448 ( .IN1(n14471), .IN2(n14472), .Q(n14460) );
  OR2X1 U14449 ( .IN1(n4475), .IN2(n4469), .Q(n14472) );
  AND2X1 U14450 ( .IN1(n14473), .IN2(n14474), .Q(g27672) );
  OR2X1 U14451 ( .IN1(n14475), .IN2(g679), .Q(n14474) );
  AND2X1 U14452 ( .IN1(test_so28), .IN2(n14476), .Q(n14475) );
  AND2X1 U14453 ( .IN1(n14354), .IN2(n13809), .Q(n14473) );
  OR2X1 U14454 ( .IN1(n10193), .IN2(n14477), .Q(n14354) );
  OR2X1 U14455 ( .IN1(n4477), .IN2(n14478), .Q(n14477) );
  AND2X1 U14456 ( .IN1(n14479), .IN2(n12966), .Q(g27621) );
  OR2X1 U14457 ( .IN1(n14480), .IN2(n14481), .Q(n14479) );
  AND2X1 U14458 ( .IN1(n4522), .IN2(g2142), .Q(n14481) );
  AND2X1 U14459 ( .IN1(n9877), .IN2(n14482), .Q(n14480) );
  INVX0 U14460 ( .INP(n4522), .ZN(n14482) );
  AND2X1 U14461 ( .IN1(n14483), .IN2(n12971), .Q(g27612) );
  OR2X1 U14462 ( .IN1(n14484), .IN2(n14485), .Q(n14483) );
  AND2X1 U14463 ( .IN1(n4523), .IN2(g1448), .Q(n14485) );
  AND2X1 U14464 ( .IN1(n9881), .IN2(n14486), .Q(n14484) );
  INVX0 U14465 ( .INP(n4523), .ZN(n14486) );
  AND2X1 U14466 ( .IN1(n14487), .IN2(n12976), .Q(g27603) );
  AND2X1 U14467 ( .IN1(n14488), .IN2(n14489), .Q(n14487) );
  INVX0 U14468 ( .INP(n14490), .ZN(n14489) );
  AND2X1 U14469 ( .IN1(n882), .IN2(n9885), .Q(n14490) );
  OR2X1 U14470 ( .IN1(n9885), .IN2(n882), .Q(n14488) );
  AND2X1 U14471 ( .IN1(n14491), .IN2(n12981), .Q(g27594) );
  OR2X1 U14472 ( .IN1(n14492), .IN2(n14493), .Q(n14491) );
  AND2X1 U14473 ( .IN1(n4521), .IN2(g74), .Q(n14493) );
  AND2X1 U14474 ( .IN1(n9889), .IN2(n14494), .Q(n14492) );
  INVX0 U14475 ( .INP(n4521), .ZN(n14494) );
  OR2X1 U14476 ( .IN1(n14495), .IN2(n14496), .Q(g27380) );
  OR2X1 U14477 ( .IN1(n14497), .IN2(n14498), .Q(n14496) );
  OR2X1 U14478 ( .IN1(n14499), .IN2(n14500), .Q(n14498) );
  AND2X1 U14479 ( .IN1(n9615), .IN2(n14501), .Q(n14500) );
  AND2X1 U14480 ( .IN1(n14502), .IN2(n8079), .Q(n14499) );
  OR2X1 U14481 ( .IN1(n14503), .IN2(n14504), .Q(n14495) );
  OR2X1 U14482 ( .IN1(n14505), .IN2(n14506), .Q(n14504) );
  AND2X1 U14483 ( .IN1(n14507), .IN2(g3151), .Q(n14506) );
  AND2X1 U14484 ( .IN1(n14508), .IN2(n14509), .Q(n14505) );
  OR2X1 U14485 ( .IN1(n14510), .IN2(n3705), .Q(n14509) );
  AND2X1 U14486 ( .IN1(n4384), .IN2(n14511), .Q(n14510) );
  OR2X1 U14487 ( .IN1(n14512), .IN2(n14513), .Q(n14503) );
  AND2X1 U14488 ( .IN1(n14514), .IN2(n14515), .Q(n14513) );
  INVX0 U14489 ( .INP(n14516), .ZN(n14515) );
  OR2X1 U14490 ( .IN1(n14517), .IN2(n14518), .Q(n14516) );
  AND2X1 U14491 ( .IN1(n8081), .IN2(n14519), .Q(n14518) );
  AND2X1 U14492 ( .IN1(n8082), .IN2(n14520), .Q(n14517) );
  AND2X1 U14493 ( .IN1(n14521), .IN2(n14522), .Q(n14514) );
  OR2X1 U14494 ( .IN1(n14523), .IN2(n14524), .Q(g27354) );
  AND2X1 U14495 ( .IN1(n14525), .IN2(n14526), .Q(n14524) );
  INVX0 U14496 ( .INP(n14527), .ZN(n14523) );
  OR2X1 U14497 ( .IN1(n14525), .IN2(n9535), .Q(n14527) );
  OR2X1 U14498 ( .IN1(n14528), .IN2(n14529), .Q(g27348) );
  AND2X1 U14499 ( .IN1(n14530), .IN2(n14526), .Q(n14529) );
  AND2X1 U14500 ( .IN1(n14531), .IN2(g2660), .Q(n14528) );
  OR2X1 U14501 ( .IN1(n14532), .IN2(n14533), .Q(g27347) );
  AND2X1 U14502 ( .IN1(n14525), .IN2(n14534), .Q(n14533) );
  INVX0 U14503 ( .INP(n14535), .ZN(n14532) );
  OR2X1 U14504 ( .IN1(n14525), .IN2(n9358), .Q(n14535) );
  OR2X1 U14505 ( .IN1(n14536), .IN2(n14537), .Q(g27346) );
  AND2X1 U14506 ( .IN1(n14538), .IN2(n14539), .Q(n14537) );
  INVX0 U14507 ( .INP(n14540), .ZN(n14536) );
  OR2X1 U14508 ( .IN1(n14538), .IN2(n9537), .Q(n14540) );
  OR2X1 U14509 ( .IN1(n14541), .IN2(n14542), .Q(g27345) );
  AND2X1 U14510 ( .IN1(n14543), .IN2(n14526), .Q(n14542) );
  OR2X1 U14511 ( .IN1(n14544), .IN2(n14545), .Q(n14526) );
  OR2X1 U14512 ( .IN1(n13916), .IN2(n13882), .Q(n14545) );
  INVX0 U14513 ( .INP(n14546), .ZN(n14541) );
  OR2X1 U14514 ( .IN1(n14543), .IN2(n9534), .Q(n14546) );
  OR2X1 U14515 ( .IN1(n14547), .IN2(n14548), .Q(g27344) );
  AND2X1 U14516 ( .IN1(n14530), .IN2(n14534), .Q(n14548) );
  AND2X1 U14517 ( .IN1(test_so89), .IN2(n14531), .Q(n14547) );
  OR2X1 U14518 ( .IN1(n14549), .IN2(n14550), .Q(g27343) );
  AND2X1 U14519 ( .IN1(n14551), .IN2(n14525), .Q(n14550) );
  INVX0 U14520 ( .INP(n14552), .ZN(n14549) );
  OR2X1 U14521 ( .IN1(n14525), .IN2(n9524), .Q(n14552) );
  OR2X1 U14522 ( .IN1(n14553), .IN2(n14554), .Q(g27342) );
  AND2X1 U14523 ( .IN1(n14555), .IN2(n14556), .Q(n14554) );
  INVX0 U14524 ( .INP(n14557), .ZN(n14553) );
  OR2X1 U14525 ( .IN1(n14555), .IN2(n9821), .Q(n14557) );
  OR2X1 U14526 ( .IN1(n14558), .IN2(n14559), .Q(g27341) );
  AND2X1 U14527 ( .IN1(n14560), .IN2(n14539), .Q(n14559) );
  INVX0 U14528 ( .INP(n14561), .ZN(n14558) );
  OR2X1 U14529 ( .IN1(n14560), .IN2(n9538), .Q(n14561) );
  OR2X1 U14530 ( .IN1(n14562), .IN2(n14563), .Q(g27340) );
  AND2X1 U14531 ( .IN1(n14538), .IN2(n14564), .Q(n14563) );
  INVX0 U14532 ( .INP(n14565), .ZN(n14562) );
  OR2X1 U14533 ( .IN1(n14538), .IN2(n9360), .Q(n14565) );
  OR2X1 U14534 ( .IN1(n14566), .IN2(n14567), .Q(g27339) );
  AND2X1 U14535 ( .IN1(n14568), .IN2(n14569), .Q(n14567) );
  AND2X1 U14536 ( .IN1(n14570), .IN2(g1270), .Q(n14566) );
  OR2X1 U14537 ( .IN1(n14571), .IN2(n14572), .Q(g27338) );
  AND2X1 U14538 ( .IN1(n14543), .IN2(n14534), .Q(n14572) );
  AND2X1 U14539 ( .IN1(n14573), .IN2(n14574), .Q(n14534) );
  OR2X1 U14540 ( .IN1(n14544), .IN2(n13900), .Q(n14574) );
  OR2X1 U14541 ( .IN1(n14575), .IN2(n14576), .Q(n14573) );
  INVX0 U14542 ( .INP(n13940), .ZN(n14576) );
  AND2X1 U14543 ( .IN1(n13917), .IN2(n13900), .Q(n13940) );
  INVX0 U14544 ( .INP(n14577), .ZN(n14571) );
  OR2X1 U14545 ( .IN1(n14543), .IN2(n9357), .Q(n14577) );
  OR2X1 U14546 ( .IN1(n14578), .IN2(n14579), .Q(g27337) );
  AND2X1 U14547 ( .IN1(n14551), .IN2(n14530), .Q(n14579) );
  AND2X1 U14548 ( .IN1(n14531), .IN2(g2654), .Q(n14578) );
  OR2X1 U14549 ( .IN1(n14580), .IN2(n14581), .Q(g27336) );
  AND2X1 U14550 ( .IN1(n14582), .IN2(n14525), .Q(n14581) );
  INVX0 U14551 ( .INP(n14583), .ZN(n14580) );
  OR2X1 U14552 ( .IN1(n14525), .IN2(n9512), .Q(n14583) );
  AND2X1 U14553 ( .IN1(g2624), .IN2(g22687), .Q(n14525) );
  OR2X1 U14554 ( .IN1(n14584), .IN2(n14585), .Q(g27335) );
  AND2X1 U14555 ( .IN1(n14586), .IN2(n14556), .Q(n14585) );
  INVX0 U14556 ( .INP(n14587), .ZN(n14584) );
  OR2X1 U14557 ( .IN1(n14586), .IN2(n9822), .Q(n14587) );
  OR2X1 U14558 ( .IN1(n14588), .IN2(n14589), .Q(g27334) );
  AND2X1 U14559 ( .IN1(n14555), .IN2(n14590), .Q(n14589) );
  INVX0 U14560 ( .INP(n14591), .ZN(n14588) );
  OR2X1 U14561 ( .IN1(n14555), .IN2(n9557), .Q(n14591) );
  OR2X1 U14562 ( .IN1(n14592), .IN2(n14593), .Q(g27333) );
  AND2X1 U14563 ( .IN1(n14594), .IN2(n14539), .Q(n14593) );
  OR2X1 U14564 ( .IN1(n14595), .IN2(n14596), .Q(n14539) );
  OR2X1 U14565 ( .IN1(n14040), .IN2(n14006), .Q(n14596) );
  INVX0 U14566 ( .INP(n14597), .ZN(n14592) );
  OR2X1 U14567 ( .IN1(n10196), .IN2(n14594), .Q(n14597) );
  OR2X1 U14568 ( .IN1(n14598), .IN2(n14599), .Q(g27332) );
  AND2X1 U14569 ( .IN1(n14560), .IN2(n14564), .Q(n14599) );
  INVX0 U14570 ( .INP(n14600), .ZN(n14598) );
  OR2X1 U14571 ( .IN1(n14560), .IN2(n9361), .Q(n14600) );
  OR2X1 U14572 ( .IN1(n14601), .IN2(n14602), .Q(g27331) );
  AND2X1 U14573 ( .IN1(n14603), .IN2(n14538), .Q(n14602) );
  INVX0 U14574 ( .INP(n14604), .ZN(n14601) );
  OR2X1 U14575 ( .IN1(n14538), .IN2(n9527), .Q(n14604) );
  OR2X1 U14576 ( .IN1(n14605), .IN2(n14606), .Q(g27330) );
  AND2X1 U14577 ( .IN1(n14607), .IN2(n14608), .Q(n14606) );
  INVX0 U14578 ( .INP(n14609), .ZN(n14605) );
  OR2X1 U14579 ( .IN1(n14607), .IN2(n9824), .Q(n14609) );
  OR2X1 U14580 ( .IN1(n14610), .IN2(n14611), .Q(g27329) );
  AND2X1 U14581 ( .IN1(n14612), .IN2(n14569), .Q(n14611) );
  INVX0 U14582 ( .INP(n14613), .ZN(n14610) );
  OR2X1 U14583 ( .IN1(n14612), .IN2(n9541), .Q(n14613) );
  OR2X1 U14584 ( .IN1(n14614), .IN2(n14615), .Q(g27328) );
  AND2X1 U14585 ( .IN1(n14568), .IN2(n14616), .Q(n14615) );
  AND2X1 U14586 ( .IN1(test_so46), .IN2(n14570), .Q(n14614) );
  OR2X1 U14587 ( .IN1(n14617), .IN2(n14618), .Q(g27327) );
  AND2X1 U14588 ( .IN1(n14619), .IN2(n14620), .Q(n14618) );
  INVX0 U14589 ( .INP(n14621), .ZN(n14617) );
  OR2X1 U14590 ( .IN1(n14619), .IN2(n9543), .Q(n14621) );
  OR2X1 U14591 ( .IN1(n14622), .IN2(n14623), .Q(g27326) );
  AND2X1 U14592 ( .IN1(n14551), .IN2(n14543), .Q(n14623) );
  AND2X1 U14593 ( .IN1(n14624), .IN2(n14625), .Q(n14551) );
  OR2X1 U14594 ( .IN1(n14575), .IN2(n13887), .Q(n14624) );
  INVX0 U14595 ( .INP(n13916), .ZN(n13887) );
  INVX0 U14596 ( .INP(n14544), .ZN(n14575) );
  OR2X1 U14597 ( .IN1(n14626), .IN2(n14627), .Q(n14544) );
  AND2X1 U14598 ( .IN1(n13910), .IN2(n10974), .Q(n14627) );
  INVX0 U14599 ( .INP(n13897), .ZN(n13910) );
  AND2X1 U14600 ( .IN1(g3229), .IN2(n13897), .Q(n14626) );
  INVX0 U14601 ( .INP(n14628), .ZN(n14622) );
  OR2X1 U14602 ( .IN1(n14543), .IN2(n9523), .Q(n14628) );
  OR2X1 U14603 ( .IN1(n14629), .IN2(n14630), .Q(g27325) );
  AND2X1 U14604 ( .IN1(n14582), .IN2(n14530), .Q(n14630) );
  AND2X1 U14605 ( .IN1(n14531), .IN2(g2651), .Q(n14629) );
  INVX0 U14606 ( .INP(n14530), .ZN(n14531) );
  AND2X1 U14607 ( .IN1(g7390), .IN2(g22687), .Q(n14530) );
  OR2X1 U14608 ( .IN1(n14631), .IN2(n14632), .Q(g27324) );
  AND2X1 U14609 ( .IN1(n14633), .IN2(n14556), .Q(n14632) );
  OR2X1 U14610 ( .IN1(n14634), .IN2(n14635), .Q(n14556) );
  OR2X1 U14611 ( .IN1(n14636), .IN2(n14637), .Q(n14635) );
  INVX0 U14612 ( .INP(n14638), .ZN(n14631) );
  OR2X1 U14613 ( .IN1(n14633), .IN2(n9823), .Q(n14638) );
  OR2X1 U14614 ( .IN1(n14639), .IN2(n14640), .Q(g27323) );
  AND2X1 U14615 ( .IN1(n14586), .IN2(n14590), .Q(n14640) );
  INVX0 U14616 ( .INP(n14641), .ZN(n14639) );
  OR2X1 U14617 ( .IN1(n14586), .IN2(n9558), .Q(n14641) );
  OR2X1 U14618 ( .IN1(n14642), .IN2(n14643), .Q(g27322) );
  AND2X1 U14619 ( .IN1(n14644), .IN2(n14555), .Q(n14643) );
  INVX0 U14620 ( .INP(n14645), .ZN(n14642) );
  OR2X1 U14621 ( .IN1(n14555), .IN2(n9809), .Q(n14645) );
  OR2X1 U14622 ( .IN1(n14646), .IN2(n14647), .Q(g27321) );
  AND2X1 U14623 ( .IN1(n14594), .IN2(n14564), .Q(n14647) );
  AND2X1 U14624 ( .IN1(n14648), .IN2(n14649), .Q(n14564) );
  OR2X1 U14625 ( .IN1(n14595), .IN2(n14024), .Q(n14649) );
  OR2X1 U14626 ( .IN1(n14650), .IN2(n14651), .Q(n14648) );
  INVX0 U14627 ( .INP(n14063), .ZN(n14651) );
  AND2X1 U14628 ( .IN1(n14041), .IN2(n14024), .Q(n14063) );
  INVX0 U14629 ( .INP(n14652), .ZN(n14646) );
  OR2X1 U14630 ( .IN1(n14594), .IN2(n9359), .Q(n14652) );
  OR2X1 U14631 ( .IN1(n14653), .IN2(n14654), .Q(g27320) );
  AND2X1 U14632 ( .IN1(n14603), .IN2(n14560), .Q(n14654) );
  INVX0 U14633 ( .INP(n14655), .ZN(n14653) );
  OR2X1 U14634 ( .IN1(n14560), .IN2(n9528), .Q(n14655) );
  OR2X1 U14635 ( .IN1(n14656), .IN2(n14657), .Q(g27319) );
  AND2X1 U14636 ( .IN1(n14658), .IN2(n14538), .Q(n14657) );
  INVX0 U14637 ( .INP(n14659), .ZN(n14656) );
  OR2X1 U14638 ( .IN1(n14538), .IN2(n9515), .Q(n14659) );
  AND2X1 U14639 ( .IN1(g1930), .IN2(g22651), .Q(n14538) );
  OR2X1 U14640 ( .IN1(n14660), .IN2(n14661), .Q(g27318) );
  AND2X1 U14641 ( .IN1(n14662), .IN2(n14608), .Q(n14661) );
  AND2X1 U14642 ( .IN1(test_so58), .IN2(n14663), .Q(n14660) );
  OR2X1 U14643 ( .IN1(n14664), .IN2(n14665), .Q(g27317) );
  AND2X1 U14644 ( .IN1(n14607), .IN2(n14666), .Q(n14665) );
  INVX0 U14645 ( .INP(n14667), .ZN(n14664) );
  OR2X1 U14646 ( .IN1(n14607), .IN2(n9560), .Q(n14667) );
  OR2X1 U14647 ( .IN1(n14668), .IN2(n14669), .Q(g27316) );
  AND2X1 U14648 ( .IN1(n14670), .IN2(n14569), .Q(n14669) );
  OR2X1 U14649 ( .IN1(n14671), .IN2(n14672), .Q(n14569) );
  OR2X1 U14650 ( .IN1(n14160), .IN2(n14126), .Q(n14672) );
  INVX0 U14651 ( .INP(n14673), .ZN(n14668) );
  OR2X1 U14652 ( .IN1(n14670), .IN2(n9539), .Q(n14673) );
  OR2X1 U14653 ( .IN1(n14674), .IN2(n14675), .Q(g27315) );
  AND2X1 U14654 ( .IN1(n14612), .IN2(n14616), .Q(n14675) );
  INVX0 U14655 ( .INP(n14676), .ZN(n14674) );
  OR2X1 U14656 ( .IN1(n14612), .IN2(n9363), .Q(n14676) );
  OR2X1 U14657 ( .IN1(n14677), .IN2(n14678), .Q(g27314) );
  AND2X1 U14658 ( .IN1(n14679), .IN2(n14568), .Q(n14678) );
  AND2X1 U14659 ( .IN1(n14570), .IN2(g1264), .Q(n14677) );
  OR2X1 U14660 ( .IN1(n14680), .IN2(n14681), .Q(g27313) );
  AND2X1 U14661 ( .IN1(n14682), .IN2(n14683), .Q(n14681) );
  INVX0 U14662 ( .INP(n14684), .ZN(n14680) );
  OR2X1 U14663 ( .IN1(n14682), .IN2(n9826), .Q(n14684) );
  OR2X1 U14664 ( .IN1(n14685), .IN2(n14686), .Q(g27312) );
  AND2X1 U14665 ( .IN1(n14687), .IN2(n14620), .Q(n14686) );
  AND2X1 U14666 ( .IN1(n14688), .IN2(g586), .Q(n14685) );
  OR2X1 U14667 ( .IN1(n14689), .IN2(n14690), .Q(g27311) );
  AND2X1 U14668 ( .IN1(n14619), .IN2(n14691), .Q(n14690) );
  INVX0 U14669 ( .INP(n14692), .ZN(n14689) );
  OR2X1 U14670 ( .IN1(n14619), .IN2(n9365), .Q(n14692) );
  OR2X1 U14671 ( .IN1(n14693), .IN2(n14694), .Q(g27310) );
  AND2X1 U14672 ( .IN1(n14582), .IN2(n14543), .Q(n14694) );
  INVX0 U14673 ( .INP(n14695), .ZN(n14582) );
  OR2X1 U14674 ( .IN1(n14696), .IN2(n14697), .Q(n14695) );
  OR2X1 U14675 ( .IN1(n14698), .IN2(n14699), .Q(n14697) );
  AND2X1 U14676 ( .IN1(n14700), .IN2(n14625), .Q(n14699) );
  AND2X1 U14677 ( .IN1(n13917), .IN2(n13897), .Q(n14700) );
  OR2X1 U14678 ( .IN1(n14701), .IN2(n14702), .Q(n13897) );
  OR2X1 U14679 ( .IN1(n14703), .IN2(n14704), .Q(n14702) );
  AND2X1 U14680 ( .IN1(n9511), .IN2(n12862), .Q(n14704) );
  AND2X1 U14681 ( .IN1(n9512), .IN2(g2624), .Q(n14703) );
  AND2X1 U14682 ( .IN1(n9513), .IN2(g7390), .Q(n14701) );
  INVX0 U14683 ( .INP(n13894), .ZN(n13917) );
  AND2X1 U14684 ( .IN1(n14705), .IN2(n10974), .Q(n14698) );
  INVX0 U14685 ( .INP(n14625), .ZN(n14705) );
  OR2X1 U14686 ( .IN1(n13900), .IN2(n13916), .Q(n14625) );
  OR2X1 U14687 ( .IN1(n14706), .IN2(n14707), .Q(n13916) );
  OR2X1 U14688 ( .IN1(n14708), .IN2(n14709), .Q(n14707) );
  AND2X1 U14689 ( .IN1(n9357), .IN2(n12862), .Q(n14709) );
  AND2X1 U14690 ( .IN1(n9358), .IN2(g2624), .Q(n14708) );
  INVX0 U14691 ( .INP(n14710), .ZN(n14706) );
  OR2X1 U14692 ( .IN1(n4370), .IN2(test_so89), .Q(n14710) );
  INVX0 U14693 ( .INP(n13882), .ZN(n13900) );
  OR2X1 U14694 ( .IN1(n14711), .IN2(n14712), .Q(n13882) );
  OR2X1 U14695 ( .IN1(n14713), .IN2(n14714), .Q(n14712) );
  AND2X1 U14696 ( .IN1(n9523), .IN2(n12862), .Q(n14714) );
  AND2X1 U14697 ( .IN1(n9524), .IN2(g2624), .Q(n14713) );
  AND2X1 U14698 ( .IN1(n9525), .IN2(g7390), .Q(n14711) );
  AND2X1 U14699 ( .IN1(g3229), .IN2(n13894), .Q(n14696) );
  OR2X1 U14700 ( .IN1(n14715), .IN2(n14716), .Q(n13894) );
  OR2X1 U14701 ( .IN1(n14717), .IN2(n14718), .Q(n14716) );
  AND2X1 U14702 ( .IN1(n9534), .IN2(n12862), .Q(n14718) );
  AND2X1 U14703 ( .IN1(n9535), .IN2(g2624), .Q(n14717) );
  AND2X1 U14704 ( .IN1(n9536), .IN2(g7390), .Q(n14715) );
  INVX0 U14705 ( .INP(n14719), .ZN(n14693) );
  OR2X1 U14706 ( .IN1(n14543), .IN2(n9511), .Q(n14719) );
  AND2X1 U14707 ( .IN1(g22687), .IN2(g7302), .Q(n14543) );
  OR2X1 U14708 ( .IN1(n14720), .IN2(n14721), .Q(g27309) );
  AND2X1 U14709 ( .IN1(n14633), .IN2(n14590), .Q(n14721) );
  AND2X1 U14710 ( .IN1(n14722), .IN2(n14723), .Q(n14590) );
  OR2X1 U14711 ( .IN1(n14724), .IN2(n14634), .Q(n14723) );
  OR2X1 U14712 ( .IN1(n14725), .IN2(n14726), .Q(n14724) );
  OR2X1 U14713 ( .IN1(n14637), .IN2(n14727), .Q(n14722) );
  INVX0 U14714 ( .INP(n14728), .ZN(n14720) );
  OR2X1 U14715 ( .IN1(n14633), .IN2(n9556), .Q(n14728) );
  OR2X1 U14716 ( .IN1(n14729), .IN2(n14730), .Q(g27308) );
  AND2X1 U14717 ( .IN1(n14644), .IN2(n14586), .Q(n14730) );
  INVX0 U14718 ( .INP(n14731), .ZN(n14729) );
  OR2X1 U14719 ( .IN1(n14586), .IN2(n9810), .Q(n14731) );
  OR2X1 U14720 ( .IN1(n14732), .IN2(n14733), .Q(g27307) );
  AND2X1 U14721 ( .IN1(n14734), .IN2(n14555), .Q(n14733) );
  INVX0 U14722 ( .INP(n14735), .ZN(n14732) );
  OR2X1 U14723 ( .IN1(n14555), .IN2(n9832), .Q(n14735) );
  AND2X1 U14724 ( .IN1(n13101), .IN2(n14736), .Q(n14555) );
  OR2X1 U14725 ( .IN1(n14737), .IN2(n14738), .Q(g27306) );
  AND2X1 U14726 ( .IN1(n14603), .IN2(n14594), .Q(n14738) );
  AND2X1 U14727 ( .IN1(n14739), .IN2(n14740), .Q(n14603) );
  OR2X1 U14728 ( .IN1(n14650), .IN2(n14011), .Q(n14739) );
  INVX0 U14729 ( .INP(n14040), .ZN(n14011) );
  INVX0 U14730 ( .INP(n14595), .ZN(n14650) );
  OR2X1 U14731 ( .IN1(n14741), .IN2(n14742), .Q(n14595) );
  AND2X1 U14732 ( .IN1(n14034), .IN2(n10974), .Q(n14742) );
  INVX0 U14733 ( .INP(n14021), .ZN(n14034) );
  AND2X1 U14734 ( .IN1(g3229), .IN2(n14021), .Q(n14741) );
  INVX0 U14735 ( .INP(n14743), .ZN(n14737) );
  OR2X1 U14736 ( .IN1(n14594), .IN2(n9526), .Q(n14743) );
  OR2X1 U14737 ( .IN1(n14744), .IN2(n14745), .Q(g27305) );
  AND2X1 U14738 ( .IN1(n14658), .IN2(n14560), .Q(n14745) );
  INVX0 U14739 ( .INP(n14746), .ZN(n14744) );
  OR2X1 U14740 ( .IN1(n14560), .IN2(n9516), .Q(n14746) );
  AND2X1 U14741 ( .IN1(g7194), .IN2(g22651), .Q(n14560) );
  OR2X1 U14742 ( .IN1(n14747), .IN2(n14748), .Q(g27304) );
  AND2X1 U14743 ( .IN1(n14749), .IN2(n14608), .Q(n14748) );
  OR2X1 U14744 ( .IN1(n14750), .IN2(n14751), .Q(n14608) );
  OR2X1 U14745 ( .IN1(n14752), .IN2(n14753), .Q(n14751) );
  INVX0 U14746 ( .INP(n14754), .ZN(n14747) );
  OR2X1 U14747 ( .IN1(n14749), .IN2(n9825), .Q(n14754) );
  OR2X1 U14748 ( .IN1(n14755), .IN2(n14756), .Q(g27303) );
  AND2X1 U14749 ( .IN1(n14662), .IN2(n14666), .Q(n14756) );
  AND2X1 U14750 ( .IN1(n14663), .IN2(g1754), .Q(n14755) );
  OR2X1 U14751 ( .IN1(n14757), .IN2(n14758), .Q(g27302) );
  AND2X1 U14752 ( .IN1(n14759), .IN2(n14607), .Q(n14758) );
  INVX0 U14753 ( .INP(n14760), .ZN(n14757) );
  OR2X1 U14754 ( .IN1(n14607), .IN2(n9812), .Q(n14760) );
  OR2X1 U14755 ( .IN1(n14761), .IN2(n14762), .Q(g27301) );
  AND2X1 U14756 ( .IN1(n14670), .IN2(n14616), .Q(n14762) );
  AND2X1 U14757 ( .IN1(n14763), .IN2(n14764), .Q(n14616) );
  OR2X1 U14758 ( .IN1(n14671), .IN2(n14144), .Q(n14764) );
  OR2X1 U14759 ( .IN1(n14765), .IN2(n14766), .Q(n14763) );
  INVX0 U14760 ( .INP(n14183), .ZN(n14766) );
  AND2X1 U14761 ( .IN1(n14161), .IN2(n14144), .Q(n14183) );
  INVX0 U14762 ( .INP(n14767), .ZN(n14761) );
  OR2X1 U14763 ( .IN1(n14670), .IN2(n9362), .Q(n14767) );
  OR2X1 U14764 ( .IN1(n14768), .IN2(n14769), .Q(g27300) );
  AND2X1 U14765 ( .IN1(n14679), .IN2(n14612), .Q(n14769) );
  INVX0 U14766 ( .INP(n14770), .ZN(n14768) );
  OR2X1 U14767 ( .IN1(n14612), .IN2(n9531), .Q(n14770) );
  OR2X1 U14768 ( .IN1(n14771), .IN2(n14772), .Q(g27299) );
  AND2X1 U14769 ( .IN1(n14773), .IN2(n14568), .Q(n14772) );
  AND2X1 U14770 ( .IN1(n14570), .IN2(g1261), .Q(n14771) );
  INVX0 U14771 ( .INP(n14568), .ZN(n14570) );
  AND2X1 U14772 ( .IN1(g1236), .IN2(g22615), .Q(n14568) );
  OR2X1 U14773 ( .IN1(n14774), .IN2(n14775), .Q(g27298) );
  AND2X1 U14774 ( .IN1(n14776), .IN2(n14683), .Q(n14775) );
  INVX0 U14775 ( .INP(n14777), .ZN(n14774) );
  OR2X1 U14776 ( .IN1(n14776), .IN2(n9827), .Q(n14777) );
  OR2X1 U14777 ( .IN1(n14778), .IN2(n14779), .Q(g27297) );
  AND2X1 U14778 ( .IN1(n14682), .IN2(n14780), .Q(n14779) );
  INVX0 U14779 ( .INP(n14781), .ZN(n14778) );
  OR2X1 U14780 ( .IN1(n14682), .IN2(n9563), .Q(n14781) );
  OR2X1 U14781 ( .IN1(n14782), .IN2(n14783), .Q(g27296) );
  AND2X1 U14782 ( .IN1(n14784), .IN2(n14620), .Q(n14783) );
  OR2X1 U14783 ( .IN1(n14785), .IN2(n14786), .Q(n14620) );
  OR2X1 U14784 ( .IN1(n14275), .IN2(n14241), .Q(n14786) );
  INVX0 U14785 ( .INP(n14787), .ZN(n14782) );
  OR2X1 U14786 ( .IN1(n14784), .IN2(n9542), .Q(n14787) );
  OR2X1 U14787 ( .IN1(n14788), .IN2(n14789), .Q(g27295) );
  AND2X1 U14788 ( .IN1(n14687), .IN2(n14691), .Q(n14789) );
  AND2X1 U14789 ( .IN1(n14688), .IN2(g583), .Q(n14788) );
  OR2X1 U14790 ( .IN1(n14790), .IN2(n14791), .Q(g27294) );
  AND2X1 U14791 ( .IN1(n14792), .IN2(n14619), .Q(n14791) );
  INVX0 U14792 ( .INP(n14793), .ZN(n14790) );
  OR2X1 U14793 ( .IN1(n14619), .IN2(n9533), .Q(n14793) );
  OR2X1 U14794 ( .IN1(n14794), .IN2(n14795), .Q(g27293) );
  AND2X1 U14795 ( .IN1(n14796), .IN2(n14797), .Q(n14795) );
  AND2X1 U14796 ( .IN1(n14798), .IN2(g391), .Q(n14794) );
  OR2X1 U14797 ( .IN1(n14799), .IN2(n14800), .Q(g27292) );
  AND2X1 U14798 ( .IN1(n14644), .IN2(n14633), .Q(n14800) );
  AND2X1 U14799 ( .IN1(n14801), .IN2(n14802), .Q(n14644) );
  OR2X1 U14800 ( .IN1(n14726), .IN2(n14803), .Q(n14801) );
  INVX0 U14801 ( .INP(n14636), .ZN(n14803) );
  INVX0 U14802 ( .INP(n14637), .ZN(n14726) );
  OR2X1 U14803 ( .IN1(n14804), .IN2(n14805), .Q(n14637) );
  AND2X1 U14804 ( .IN1(n14806), .IN2(n10974), .Q(n14805) );
  INVX0 U14805 ( .INP(n14807), .ZN(n14806) );
  AND2X1 U14806 ( .IN1(g3229), .IN2(n14807), .Q(n14804) );
  INVX0 U14807 ( .INP(n14808), .ZN(n14799) );
  OR2X1 U14808 ( .IN1(n14633), .IN2(n9811), .Q(n14808) );
  OR2X1 U14809 ( .IN1(n14809), .IN2(n14810), .Q(g27291) );
  AND2X1 U14810 ( .IN1(n14734), .IN2(n14586), .Q(n14810) );
  INVX0 U14811 ( .INP(n14811), .ZN(n14809) );
  OR2X1 U14812 ( .IN1(n14586), .IN2(n9833), .Q(n14811) );
  AND2X1 U14813 ( .IN1(g7264), .IN2(n14736), .Q(n14586) );
  OR2X1 U14814 ( .IN1(n14812), .IN2(n14813), .Q(g27290) );
  AND2X1 U14815 ( .IN1(n14658), .IN2(n14594), .Q(n14813) );
  INVX0 U14816 ( .INP(n14814), .ZN(n14658) );
  OR2X1 U14817 ( .IN1(n14815), .IN2(n14816), .Q(n14814) );
  OR2X1 U14818 ( .IN1(n14817), .IN2(n14818), .Q(n14816) );
  AND2X1 U14819 ( .IN1(n14819), .IN2(n14740), .Q(n14818) );
  AND2X1 U14820 ( .IN1(n14041), .IN2(n14021), .Q(n14819) );
  OR2X1 U14821 ( .IN1(n14820), .IN2(n14821), .Q(n14021) );
  OR2X1 U14822 ( .IN1(n14822), .IN2(n14823), .Q(n14821) );
  AND2X1 U14823 ( .IN1(n9516), .IN2(g7194), .Q(n14823) );
  AND2X1 U14824 ( .IN1(n9514), .IN2(n13973), .Q(n14822) );
  AND2X1 U14825 ( .IN1(n9515), .IN2(g1930), .Q(n14820) );
  INVX0 U14826 ( .INP(n14018), .ZN(n14041) );
  AND2X1 U14827 ( .IN1(n14824), .IN2(n10974), .Q(n14817) );
  INVX0 U14828 ( .INP(n14740), .ZN(n14824) );
  OR2X1 U14829 ( .IN1(n14024), .IN2(n14040), .Q(n14740) );
  OR2X1 U14830 ( .IN1(n14825), .IN2(n14826), .Q(n14040) );
  OR2X1 U14831 ( .IN1(n14827), .IN2(n14828), .Q(n14826) );
  AND2X1 U14832 ( .IN1(n9361), .IN2(g7194), .Q(n14828) );
  AND2X1 U14833 ( .IN1(n9359), .IN2(n13973), .Q(n14827) );
  AND2X1 U14834 ( .IN1(n9360), .IN2(g1930), .Q(n14825) );
  INVX0 U14835 ( .INP(n14006), .ZN(n14024) );
  OR2X1 U14836 ( .IN1(n14829), .IN2(n14830), .Q(n14006) );
  OR2X1 U14837 ( .IN1(n14831), .IN2(n14832), .Q(n14830) );
  AND2X1 U14838 ( .IN1(n9528), .IN2(g7194), .Q(n14832) );
  AND2X1 U14839 ( .IN1(n9526), .IN2(n13973), .Q(n14831) );
  AND2X1 U14840 ( .IN1(n9527), .IN2(g1930), .Q(n14829) );
  AND2X1 U14841 ( .IN1(g3229), .IN2(n14018), .Q(n14815) );
  OR2X1 U14842 ( .IN1(n14833), .IN2(n14834), .Q(n14018) );
  OR2X1 U14843 ( .IN1(n14835), .IN2(n14836), .Q(n14834) );
  AND2X1 U14844 ( .IN1(n9538), .IN2(g7194), .Q(n14836) );
  AND2X1 U14845 ( .IN1(n13973), .IN2(n10196), .Q(n14835) );
  AND2X1 U14846 ( .IN1(n9537), .IN2(g1930), .Q(n14833) );
  INVX0 U14847 ( .INP(n14837), .ZN(n14812) );
  OR2X1 U14848 ( .IN1(n14594), .IN2(n9514), .Q(n14837) );
  AND2X1 U14849 ( .IN1(g22651), .IN2(g7052), .Q(n14594) );
  OR2X1 U14850 ( .IN1(n14838), .IN2(n14839), .Q(g27289) );
  AND2X1 U14851 ( .IN1(n14749), .IN2(n14666), .Q(n14839) );
  AND2X1 U14852 ( .IN1(n14840), .IN2(n14841), .Q(n14666) );
  INVX0 U14853 ( .INP(n14842), .ZN(n14841) );
  AND2X1 U14854 ( .IN1(n14843), .IN2(n14844), .Q(n14842) );
  AND2X1 U14855 ( .IN1(n14845), .IN2(n14753), .Q(n14843) );
  OR2X1 U14856 ( .IN1(n14753), .IN2(n14844), .Q(n14840) );
  INVX0 U14857 ( .INP(n14846), .ZN(n14838) );
  OR2X1 U14858 ( .IN1(n14749), .IN2(n9559), .Q(n14846) );
  OR2X1 U14859 ( .IN1(n14847), .IN2(n14848), .Q(g27288) );
  AND2X1 U14860 ( .IN1(n14759), .IN2(n14662), .Q(n14848) );
  AND2X1 U14861 ( .IN1(n14663), .IN2(g1739), .Q(n14847) );
  OR2X1 U14862 ( .IN1(n14849), .IN2(n14850), .Q(g27287) );
  AND2X1 U14863 ( .IN1(n14851), .IN2(n14607), .Q(n14850) );
  INVX0 U14864 ( .INP(n14852), .ZN(n14849) );
  OR2X1 U14865 ( .IN1(n14607), .IN2(n9835), .Q(n14852) );
  AND2X1 U14866 ( .IN1(n13111), .IN2(n14853), .Q(n14607) );
  OR2X1 U14867 ( .IN1(n14854), .IN2(n14855), .Q(g27286) );
  AND2X1 U14868 ( .IN1(n14679), .IN2(n14670), .Q(n14855) );
  AND2X1 U14869 ( .IN1(n14856), .IN2(n14857), .Q(n14679) );
  OR2X1 U14870 ( .IN1(n14765), .IN2(n14131), .Q(n14856) );
  INVX0 U14871 ( .INP(n14160), .ZN(n14131) );
  INVX0 U14872 ( .INP(n14671), .ZN(n14765) );
  OR2X1 U14873 ( .IN1(n14858), .IN2(n14859), .Q(n14671) );
  AND2X1 U14874 ( .IN1(n14154), .IN2(n10974), .Q(n14859) );
  INVX0 U14875 ( .INP(n14141), .ZN(n14154) );
  AND2X1 U14876 ( .IN1(g3229), .IN2(n14141), .Q(n14858) );
  INVX0 U14877 ( .INP(n14860), .ZN(n14854) );
  OR2X1 U14878 ( .IN1(n14670), .IN2(n9529), .Q(n14860) );
  OR2X1 U14879 ( .IN1(n14861), .IN2(n14862), .Q(g27285) );
  AND2X1 U14880 ( .IN1(n14773), .IN2(n14612), .Q(n14862) );
  INVX0 U14881 ( .INP(n14863), .ZN(n14861) );
  OR2X1 U14882 ( .IN1(n14612), .IN2(n9519), .Q(n14863) );
  AND2X1 U14883 ( .IN1(g6944), .IN2(g22615), .Q(n14612) );
  OR2X1 U14884 ( .IN1(n14864), .IN2(n14865), .Q(g27284) );
  AND2X1 U14885 ( .IN1(n14866), .IN2(n14683), .Q(n14865) );
  OR2X1 U14886 ( .IN1(n14867), .IN2(n14868), .Q(n14683) );
  OR2X1 U14887 ( .IN1(n14869), .IN2(n14870), .Q(n14868) );
  AND2X1 U14888 ( .IN1(n14871), .IN2(g1085), .Q(n14864) );
  OR2X1 U14889 ( .IN1(n14872), .IN2(n14873), .Q(g27283) );
  AND2X1 U14890 ( .IN1(n14776), .IN2(n14780), .Q(n14873) );
  INVX0 U14891 ( .INP(n14874), .ZN(n14872) );
  OR2X1 U14892 ( .IN1(n14776), .IN2(n9562), .Q(n14874) );
  OR2X1 U14893 ( .IN1(n14875), .IN2(n14876), .Q(g27282) );
  AND2X1 U14894 ( .IN1(n14877), .IN2(n14682), .Q(n14876) );
  INVX0 U14895 ( .INP(n14878), .ZN(n14875) );
  OR2X1 U14896 ( .IN1(n14682), .IN2(n9815), .Q(n14878) );
  OR2X1 U14897 ( .IN1(n14879), .IN2(n14880), .Q(g27281) );
  AND2X1 U14898 ( .IN1(n14784), .IN2(n14691), .Q(n14880) );
  AND2X1 U14899 ( .IN1(n14881), .IN2(n14882), .Q(n14691) );
  OR2X1 U14900 ( .IN1(n14785), .IN2(n14259), .Q(n14882) );
  OR2X1 U14901 ( .IN1(n14883), .IN2(n14884), .Q(n14881) );
  INVX0 U14902 ( .INP(n14298), .ZN(n14884) );
  AND2X1 U14903 ( .IN1(n14276), .IN2(n14259), .Q(n14298) );
  INVX0 U14904 ( .INP(n14885), .ZN(n14879) );
  OR2X1 U14905 ( .IN1(n14784), .IN2(n9364), .Q(n14885) );
  OR2X1 U14906 ( .IN1(n14886), .IN2(n14887), .Q(g27280) );
  AND2X1 U14907 ( .IN1(n14792), .IN2(n14687), .Q(n14887) );
  AND2X1 U14908 ( .IN1(test_so25), .IN2(n14688), .Q(n14886) );
  OR2X1 U14909 ( .IN1(n14888), .IN2(n14889), .Q(g27279) );
  AND2X1 U14910 ( .IN1(n14890), .IN2(n14619), .Q(n14889) );
  INVX0 U14911 ( .INP(n14891), .ZN(n14888) );
  OR2X1 U14912 ( .IN1(n14619), .IN2(n9521), .Q(n14891) );
  AND2X1 U14913 ( .IN1(g550), .IN2(g22578), .Q(n14619) );
  OR2X1 U14914 ( .IN1(n14892), .IN2(n14893), .Q(g27278) );
  AND2X1 U14915 ( .IN1(n14894), .IN2(n14797), .Q(n14893) );
  INVX0 U14916 ( .INP(n14895), .ZN(n14892) );
  OR2X1 U14917 ( .IN1(n14894), .IN2(n9830), .Q(n14895) );
  OR2X1 U14918 ( .IN1(n14896), .IN2(n14897), .Q(g27277) );
  AND2X1 U14919 ( .IN1(n14796), .IN2(n14898), .Q(n14897) );
  AND2X1 U14920 ( .IN1(n14798), .IN2(g376), .Q(n14896) );
  OR2X1 U14921 ( .IN1(n14899), .IN2(n14900), .Q(g27276) );
  AND2X1 U14922 ( .IN1(n14734), .IN2(n14633), .Q(n14900) );
  INVX0 U14923 ( .INP(n14901), .ZN(n14734) );
  OR2X1 U14924 ( .IN1(n14902), .IN2(n14903), .Q(n14901) );
  OR2X1 U14925 ( .IN1(n14904), .IN2(n14905), .Q(n14903) );
  AND2X1 U14926 ( .IN1(n14906), .IN2(n14802), .Q(n14905) );
  AND2X1 U14927 ( .IN1(n14907), .IN2(n14807), .Q(n14906) );
  OR2X1 U14928 ( .IN1(n14908), .IN2(n14909), .Q(n14807) );
  OR2X1 U14929 ( .IN1(n14910), .IN2(n14911), .Q(n14909) );
  AND2X1 U14930 ( .IN1(n9834), .IN2(n13116), .Q(n14911) );
  AND2X1 U14931 ( .IN1(n9832), .IN2(n13101), .Q(n14910) );
  AND2X1 U14932 ( .IN1(n9833), .IN2(n13106), .Q(n14908) );
  INVX0 U14933 ( .INP(n14725), .ZN(n14907) );
  INVX0 U14934 ( .INP(n14912), .ZN(n14904) );
  OR2X1 U14935 ( .IN1(n14802), .IN2(g3229), .Q(n14912) );
  OR2X1 U14936 ( .IN1(n14727), .IN2(n14636), .Q(n14802) );
  OR2X1 U14937 ( .IN1(n14913), .IN2(n14914), .Q(n14636) );
  OR2X1 U14938 ( .IN1(n14915), .IN2(n14916), .Q(n14914) );
  AND2X1 U14939 ( .IN1(n9556), .IN2(n13116), .Q(n14916) );
  AND2X1 U14940 ( .IN1(n9557), .IN2(n13101), .Q(n14915) );
  AND2X1 U14941 ( .IN1(n9558), .IN2(n13106), .Q(n14913) );
  INVX0 U14942 ( .INP(n14634), .ZN(n14727) );
  OR2X1 U14943 ( .IN1(n14917), .IN2(n14918), .Q(n14634) );
  OR2X1 U14944 ( .IN1(n14919), .IN2(n14920), .Q(n14918) );
  AND2X1 U14945 ( .IN1(n9811), .IN2(n13116), .Q(n14920) );
  AND2X1 U14946 ( .IN1(n9809), .IN2(n13101), .Q(n14919) );
  AND2X1 U14947 ( .IN1(n9810), .IN2(n13106), .Q(n14917) );
  AND2X1 U14948 ( .IN1(g3229), .IN2(n14725), .Q(n14902) );
  OR2X1 U14949 ( .IN1(n14921), .IN2(n14922), .Q(n14725) );
  OR2X1 U14950 ( .IN1(n14923), .IN2(n14924), .Q(n14922) );
  AND2X1 U14951 ( .IN1(n9823), .IN2(n13116), .Q(n14924) );
  AND2X1 U14952 ( .IN1(n9821), .IN2(n13101), .Q(n14923) );
  AND2X1 U14953 ( .IN1(n9822), .IN2(n13106), .Q(n14921) );
  INVX0 U14954 ( .INP(n14925), .ZN(n14899) );
  OR2X1 U14955 ( .IN1(n14633), .IN2(n9834), .Q(n14925) );
  AND2X1 U14956 ( .IN1(g5555), .IN2(n14736), .Q(n14633) );
  INVX0 U14957 ( .INP(n14926), .ZN(n14736) );
  OR2X1 U14958 ( .IN1(n14927), .IN2(n10866), .Q(n14926) );
  AND2X1 U14959 ( .IN1(n10672), .IN2(n10871), .Q(n14927) );
  OR2X1 U14960 ( .IN1(n14928), .IN2(n14929), .Q(g27275) );
  AND2X1 U14961 ( .IN1(n14759), .IN2(n14749), .Q(n14929) );
  AND2X1 U14962 ( .IN1(n14930), .IN2(n14931), .Q(n14759) );
  INVX0 U14963 ( .INP(n14932), .ZN(n14930) );
  AND2X1 U14964 ( .IN1(n14753), .IN2(n14752), .Q(n14932) );
  OR2X1 U14965 ( .IN1(n14933), .IN2(n14934), .Q(n14753) );
  AND2X1 U14966 ( .IN1(n14935), .IN2(n10974), .Q(n14934) );
  INVX0 U14967 ( .INP(n14936), .ZN(n14935) );
  AND2X1 U14968 ( .IN1(g3229), .IN2(n14936), .Q(n14933) );
  INVX0 U14969 ( .INP(n14937), .ZN(n14928) );
  OR2X1 U14970 ( .IN1(n14749), .IN2(n9814), .Q(n14937) );
  OR2X1 U14971 ( .IN1(n14938), .IN2(n14939), .Q(g27274) );
  AND2X1 U14972 ( .IN1(n14851), .IN2(n14662), .Q(n14939) );
  AND2X1 U14973 ( .IN1(n14663), .IN2(g1724), .Q(n14938) );
  INVX0 U14974 ( .INP(n14662), .ZN(n14663) );
  AND2X1 U14975 ( .IN1(g7014), .IN2(n14853), .Q(n14662) );
  OR2X1 U14976 ( .IN1(n14940), .IN2(n14941), .Q(g27273) );
  AND2X1 U14977 ( .IN1(n14773), .IN2(n14670), .Q(n14941) );
  INVX0 U14978 ( .INP(n14942), .ZN(n14773) );
  OR2X1 U14979 ( .IN1(n14943), .IN2(n14944), .Q(n14942) );
  OR2X1 U14980 ( .IN1(n14945), .IN2(n14946), .Q(n14944) );
  AND2X1 U14981 ( .IN1(n14947), .IN2(n14857), .Q(n14946) );
  AND2X1 U14982 ( .IN1(n14161), .IN2(n14141), .Q(n14947) );
  OR2X1 U14983 ( .IN1(n14948), .IN2(n14949), .Q(n14141) );
  OR2X1 U14984 ( .IN1(n14950), .IN2(n14951), .Q(n14949) );
  AND2X1 U14985 ( .IN1(n9519), .IN2(g6944), .Q(n14951) );
  AND2X1 U14986 ( .IN1(n9518), .IN2(g1236), .Q(n14950) );
  AND2X1 U14987 ( .IN1(n9517), .IN2(n13842), .Q(n14948) );
  INVX0 U14988 ( .INP(n14138), .ZN(n14161) );
  AND2X1 U14989 ( .IN1(n14952), .IN2(n10974), .Q(n14945) );
  INVX0 U14990 ( .INP(n14857), .ZN(n14952) );
  OR2X1 U14991 ( .IN1(n14144), .IN2(n14160), .Q(n14857) );
  OR2X1 U14992 ( .IN1(n14953), .IN2(n14954), .Q(n14160) );
  OR2X1 U14993 ( .IN1(n14955), .IN2(n14956), .Q(n14954) );
  AND2X1 U14994 ( .IN1(n9363), .IN2(g6944), .Q(n14956) );
  AND2X1 U14995 ( .IN1(g1236), .IN2(n10207), .Q(n14955) );
  AND2X1 U14996 ( .IN1(n9362), .IN2(n13842), .Q(n14953) );
  INVX0 U14997 ( .INP(n14126), .ZN(n14144) );
  OR2X1 U14998 ( .IN1(n14957), .IN2(n14958), .Q(n14126) );
  OR2X1 U14999 ( .IN1(n14959), .IN2(n14960), .Q(n14958) );
  AND2X1 U15000 ( .IN1(n9531), .IN2(g6944), .Q(n14960) );
  AND2X1 U15001 ( .IN1(n9530), .IN2(g1236), .Q(n14959) );
  AND2X1 U15002 ( .IN1(n9529), .IN2(n13842), .Q(n14957) );
  AND2X1 U15003 ( .IN1(g3229), .IN2(n14138), .Q(n14943) );
  OR2X1 U15004 ( .IN1(n14961), .IN2(n14962), .Q(n14138) );
  OR2X1 U15005 ( .IN1(n14963), .IN2(n14964), .Q(n14962) );
  AND2X1 U15006 ( .IN1(n9541), .IN2(g6944), .Q(n14964) );
  AND2X1 U15007 ( .IN1(n9540), .IN2(g1236), .Q(n14963) );
  AND2X1 U15008 ( .IN1(n9539), .IN2(n13842), .Q(n14961) );
  INVX0 U15009 ( .INP(n14965), .ZN(n14940) );
  OR2X1 U15010 ( .IN1(n14670), .IN2(n9517), .Q(n14965) );
  AND2X1 U15011 ( .IN1(g22615), .IN2(g6750), .Q(n14670) );
  OR2X1 U15012 ( .IN1(n14966), .IN2(n14967), .Q(g27272) );
  AND2X1 U15013 ( .IN1(n14866), .IN2(n14780), .Q(n14967) );
  AND2X1 U15014 ( .IN1(n14968), .IN2(n14969), .Q(n14780) );
  OR2X1 U15015 ( .IN1(n14970), .IN2(n14867), .Q(n14969) );
  OR2X1 U15016 ( .IN1(n14971), .IN2(n14972), .Q(n14970) );
  OR2X1 U15017 ( .IN1(n14870), .IN2(n14973), .Q(n14968) );
  AND2X1 U15018 ( .IN1(test_so37), .IN2(n14871), .Q(n14966) );
  OR2X1 U15019 ( .IN1(n14974), .IN2(n14975), .Q(g27271) );
  AND2X1 U15020 ( .IN1(n14877), .IN2(n14776), .Q(n14975) );
  INVX0 U15021 ( .INP(n14976), .ZN(n14974) );
  OR2X1 U15022 ( .IN1(n14776), .IN2(n9816), .Q(n14976) );
  OR2X1 U15023 ( .IN1(n14977), .IN2(n14978), .Q(g27270) );
  AND2X1 U15024 ( .IN1(n14979), .IN2(n14682), .Q(n14978) );
  INVX0 U15025 ( .INP(n14980), .ZN(n14977) );
  OR2X1 U15026 ( .IN1(n14682), .IN2(n9838), .Q(n14980) );
  AND2X1 U15027 ( .IN1(g1088), .IN2(n14981), .Q(n14682) );
  OR2X1 U15028 ( .IN1(n14982), .IN2(n14983), .Q(g27269) );
  AND2X1 U15029 ( .IN1(n14792), .IN2(n14784), .Q(n14983) );
  AND2X1 U15030 ( .IN1(n14984), .IN2(n14985), .Q(n14792) );
  OR2X1 U15031 ( .IN1(n14883), .IN2(n14246), .Q(n14984) );
  INVX0 U15032 ( .INP(n14275), .ZN(n14246) );
  INVX0 U15033 ( .INP(n14785), .ZN(n14883) );
  OR2X1 U15034 ( .IN1(n14986), .IN2(n14987), .Q(n14785) );
  AND2X1 U15035 ( .IN1(n14269), .IN2(n10974), .Q(n14987) );
  INVX0 U15036 ( .INP(n14256), .ZN(n14269) );
  AND2X1 U15037 ( .IN1(g3229), .IN2(n14256), .Q(n14986) );
  INVX0 U15038 ( .INP(n14988), .ZN(n14982) );
  OR2X1 U15039 ( .IN1(n14784), .IN2(n9532), .Q(n14988) );
  OR2X1 U15040 ( .IN1(n14989), .IN2(n14990), .Q(g27268) );
  AND2X1 U15041 ( .IN1(n14890), .IN2(n14687), .Q(n14990) );
  AND2X1 U15042 ( .IN1(n14688), .IN2(g577), .Q(n14989) );
  INVX0 U15043 ( .INP(n14687), .ZN(n14688) );
  AND2X1 U15044 ( .IN1(g6642), .IN2(g22578), .Q(n14687) );
  OR2X1 U15045 ( .IN1(n14991), .IN2(n14992), .Q(g27267) );
  AND2X1 U15046 ( .IN1(n14993), .IN2(n14797), .Q(n14992) );
  OR2X1 U15047 ( .IN1(n14994), .IN2(n14995), .Q(n14797) );
  OR2X1 U15048 ( .IN1(n14996), .IN2(n14997), .Q(n14995) );
  INVX0 U15049 ( .INP(n14998), .ZN(n14991) );
  OR2X1 U15050 ( .IN1(n14993), .IN2(n9831), .Q(n14998) );
  OR2X1 U15051 ( .IN1(n14999), .IN2(n15000), .Q(g27266) );
  AND2X1 U15052 ( .IN1(n14894), .IN2(n14898), .Q(n15000) );
  INVX0 U15053 ( .INP(n15001), .ZN(n14999) );
  OR2X1 U15054 ( .IN1(n14894), .IN2(n9566), .Q(n15001) );
  OR2X1 U15055 ( .IN1(n15002), .IN2(n15003), .Q(g27265) );
  AND2X1 U15056 ( .IN1(n15004), .IN2(n14796), .Q(n15003) );
  AND2X1 U15057 ( .IN1(n14798), .IN2(g361), .Q(n15002) );
  OR2X1 U15058 ( .IN1(n15005), .IN2(n15006), .Q(g27264) );
  AND2X1 U15059 ( .IN1(n14851), .IN2(n14749), .Q(n15006) );
  AND2X1 U15060 ( .IN1(n15007), .IN2(n15008), .Q(n14851) );
  AND2X1 U15061 ( .IN1(n15009), .IN2(n15010), .Q(n15008) );
  INVX0 U15062 ( .INP(n15011), .ZN(n15010) );
  AND2X1 U15063 ( .IN1(n15012), .IN2(n14931), .Q(n15011) );
  AND2X1 U15064 ( .IN1(n14845), .IN2(n14936), .Q(n15012) );
  OR2X1 U15065 ( .IN1(n15013), .IN2(n15014), .Q(n14936) );
  OR2X1 U15066 ( .IN1(n15015), .IN2(n15016), .Q(n15014) );
  AND2X1 U15067 ( .IN1(n9837), .IN2(n13248), .Q(n15016) );
  AND2X1 U15068 ( .IN1(n9835), .IN2(n13111), .Q(n15015) );
  AND2X1 U15069 ( .IN1(n9836), .IN2(n13239), .Q(n15013) );
  OR2X1 U15070 ( .IN1(n14931), .IN2(g3229), .Q(n15009) );
  OR2X1 U15071 ( .IN1(n14844), .IN2(n14752), .Q(n14931) );
  OR2X1 U15072 ( .IN1(n15017), .IN2(n15018), .Q(n14752) );
  OR2X1 U15073 ( .IN1(n15019), .IN2(n15020), .Q(n15018) );
  AND2X1 U15074 ( .IN1(n9559), .IN2(n13248), .Q(n15020) );
  AND2X1 U15075 ( .IN1(n9560), .IN2(n13111), .Q(n15019) );
  AND2X1 U15076 ( .IN1(n9561), .IN2(n13239), .Q(n15017) );
  INVX0 U15077 ( .INP(n14750), .ZN(n14844) );
  OR2X1 U15078 ( .IN1(n15021), .IN2(n15022), .Q(n14750) );
  OR2X1 U15079 ( .IN1(n15023), .IN2(n15024), .Q(n15022) );
  AND2X1 U15080 ( .IN1(n9814), .IN2(n13248), .Q(n15024) );
  AND2X1 U15081 ( .IN1(n9812), .IN2(n13111), .Q(n15023) );
  AND2X1 U15082 ( .IN1(n9813), .IN2(n13239), .Q(n15021) );
  OR2X1 U15083 ( .IN1(n10974), .IN2(n14845), .Q(n15007) );
  AND2X1 U15084 ( .IN1(n15025), .IN2(n15026), .Q(n14845) );
  INVX0 U15085 ( .INP(n15027), .ZN(n15026) );
  OR2X1 U15086 ( .IN1(n15028), .IN2(n15029), .Q(n15027) );
  AND2X1 U15087 ( .IN1(n9825), .IN2(n13248), .Q(n15029) );
  AND2X1 U15088 ( .IN1(n9824), .IN2(n13111), .Q(n15028) );
  OR2X1 U15089 ( .IN1(n4525), .IN2(test_so58), .Q(n15025) );
  INVX0 U15090 ( .INP(n15030), .ZN(n15005) );
  OR2X1 U15091 ( .IN1(n14749), .IN2(n9837), .Q(n15030) );
  AND2X1 U15092 ( .IN1(g5511), .IN2(n14853), .Q(n14749) );
  INVX0 U15093 ( .INP(n15031), .ZN(n14853) );
  OR2X1 U15094 ( .IN1(n15032), .IN2(n10801), .Q(n15031) );
  AND2X1 U15095 ( .IN1(n10672), .IN2(n10807), .Q(n15032) );
  OR2X1 U15096 ( .IN1(n15033), .IN2(n15034), .Q(g27263) );
  AND2X1 U15097 ( .IN1(n14877), .IN2(n14866), .Q(n15034) );
  AND2X1 U15098 ( .IN1(n15035), .IN2(n15036), .Q(n14877) );
  OR2X1 U15099 ( .IN1(n14972), .IN2(n15037), .Q(n15035) );
  INVX0 U15100 ( .INP(n14869), .ZN(n15037) );
  INVX0 U15101 ( .INP(n14870), .ZN(n14972) );
  OR2X1 U15102 ( .IN1(n15038), .IN2(n15039), .Q(n14870) );
  AND2X1 U15103 ( .IN1(n15040), .IN2(n10974), .Q(n15039) );
  INVX0 U15104 ( .INP(n15041), .ZN(n15040) );
  AND2X1 U15105 ( .IN1(g3229), .IN2(n15041), .Q(n15038) );
  AND2X1 U15106 ( .IN1(n14871), .IN2(g1056), .Q(n15033) );
  OR2X1 U15107 ( .IN1(n15042), .IN2(n15043), .Q(g27262) );
  AND2X1 U15108 ( .IN1(n14979), .IN2(n14776), .Q(n15043) );
  INVX0 U15109 ( .INP(n15044), .ZN(n15042) );
  OR2X1 U15110 ( .IN1(n14776), .IN2(n9839), .Q(n15044) );
  AND2X1 U15111 ( .IN1(g6712), .IN2(n14981), .Q(n14776) );
  OR2X1 U15112 ( .IN1(n15045), .IN2(n15046), .Q(g27261) );
  AND2X1 U15113 ( .IN1(n14890), .IN2(n14784), .Q(n15046) );
  INVX0 U15114 ( .INP(n15047), .ZN(n14890) );
  OR2X1 U15115 ( .IN1(n15048), .IN2(n15049), .Q(n15047) );
  OR2X1 U15116 ( .IN1(n15050), .IN2(n15051), .Q(n15049) );
  AND2X1 U15117 ( .IN1(n15052), .IN2(n14985), .Q(n15051) );
  AND2X1 U15118 ( .IN1(n14276), .IN2(n14256), .Q(n15052) );
  OR2X1 U15119 ( .IN1(n15053), .IN2(n15054), .Q(n14256) );
  OR2X1 U15120 ( .IN1(n15055), .IN2(n15056), .Q(n15054) );
  AND2X1 U15121 ( .IN1(n9521), .IN2(g550), .Q(n15056) );
  AND2X1 U15122 ( .IN1(n9520), .IN2(n11054), .Q(n15055) );
  AND2X1 U15123 ( .IN1(n9522), .IN2(g6642), .Q(n15053) );
  INVX0 U15124 ( .INP(n14253), .ZN(n14276) );
  AND2X1 U15125 ( .IN1(n15057), .IN2(n10974), .Q(n15050) );
  INVX0 U15126 ( .INP(n14985), .ZN(n15057) );
  OR2X1 U15127 ( .IN1(n14259), .IN2(n14275), .Q(n14985) );
  OR2X1 U15128 ( .IN1(n15058), .IN2(n15059), .Q(n14275) );
  OR2X1 U15129 ( .IN1(n15060), .IN2(n15061), .Q(n15059) );
  AND2X1 U15130 ( .IN1(n9365), .IN2(g550), .Q(n15061) );
  AND2X1 U15131 ( .IN1(n9364), .IN2(n11054), .Q(n15060) );
  AND2X1 U15132 ( .IN1(n9366), .IN2(g6642), .Q(n15058) );
  INVX0 U15133 ( .INP(n14241), .ZN(n14259) );
  OR2X1 U15134 ( .IN1(n15062), .IN2(n15063), .Q(n14241) );
  OR2X1 U15135 ( .IN1(n15064), .IN2(n15065), .Q(n15063) );
  AND2X1 U15136 ( .IN1(n9533), .IN2(g550), .Q(n15065) );
  AND2X1 U15137 ( .IN1(n9532), .IN2(n11054), .Q(n15064) );
  INVX0 U15138 ( .INP(n15066), .ZN(n15062) );
  OR2X1 U15139 ( .IN1(n4372), .IN2(test_so25), .Q(n15066) );
  AND2X1 U15140 ( .IN1(g3229), .IN2(n14253), .Q(n15048) );
  OR2X1 U15141 ( .IN1(n15067), .IN2(n15068), .Q(n14253) );
  OR2X1 U15142 ( .IN1(n15069), .IN2(n15070), .Q(n15068) );
  AND2X1 U15143 ( .IN1(n9543), .IN2(g550), .Q(n15070) );
  AND2X1 U15144 ( .IN1(n9542), .IN2(n11054), .Q(n15069) );
  AND2X1 U15145 ( .IN1(n9544), .IN2(g6642), .Q(n15067) );
  INVX0 U15146 ( .INP(n15071), .ZN(n15045) );
  OR2X1 U15147 ( .IN1(n14784), .IN2(n9520), .Q(n15071) );
  AND2X1 U15148 ( .IN1(g22578), .IN2(g6485), .Q(n14784) );
  OR2X1 U15149 ( .IN1(n15072), .IN2(n15073), .Q(g27260) );
  AND2X1 U15150 ( .IN1(n14993), .IN2(n14898), .Q(n15073) );
  AND2X1 U15151 ( .IN1(n15074), .IN2(n15075), .Q(n14898) );
  OR2X1 U15152 ( .IN1(n15076), .IN2(n14994), .Q(n15075) );
  OR2X1 U15153 ( .IN1(n15077), .IN2(n15078), .Q(n15076) );
  OR2X1 U15154 ( .IN1(n14997), .IN2(n15079), .Q(n15074) );
  INVX0 U15155 ( .INP(n15080), .ZN(n15072) );
  OR2X1 U15156 ( .IN1(n14993), .IN2(n9564), .Q(n15080) );
  OR2X1 U15157 ( .IN1(n15081), .IN2(n15082), .Q(g27259) );
  AND2X1 U15158 ( .IN1(n15004), .IN2(n14894), .Q(n15082) );
  INVX0 U15159 ( .INP(n15083), .ZN(n15081) );
  OR2X1 U15160 ( .IN1(n14894), .IN2(n9819), .Q(n15083) );
  OR2X1 U15161 ( .IN1(n15084), .IN2(n15085), .Q(g27258) );
  AND2X1 U15162 ( .IN1(n15086), .IN2(n14796), .Q(n15085) );
  AND2X1 U15163 ( .IN1(test_so16), .IN2(n14798), .Q(n15084) );
  INVX0 U15164 ( .INP(n14796), .ZN(n14798) );
  AND2X1 U15165 ( .IN1(n13375), .IN2(n15087), .Q(n14796) );
  OR2X1 U15166 ( .IN1(n15088), .IN2(n15089), .Q(g27257) );
  AND2X1 U15167 ( .IN1(n14979), .IN2(n14866), .Q(n15089) );
  INVX0 U15168 ( .INP(n15090), .ZN(n14979) );
  OR2X1 U15169 ( .IN1(n15091), .IN2(n15092), .Q(n15090) );
  OR2X1 U15170 ( .IN1(n15093), .IN2(n15094), .Q(n15092) );
  AND2X1 U15171 ( .IN1(n15095), .IN2(n15036), .Q(n15094) );
  AND2X1 U15172 ( .IN1(n15096), .IN2(n15041), .Q(n15095) );
  OR2X1 U15173 ( .IN1(n15097), .IN2(n15098), .Q(n15041) );
  OR2X1 U15174 ( .IN1(n15099), .IN2(n15100), .Q(n15098) );
  AND2X1 U15175 ( .IN1(n9839), .IN2(g6712), .Q(n15100) );
  AND2X1 U15176 ( .IN1(n9840), .IN2(g5472), .Q(n15099) );
  AND2X1 U15177 ( .IN1(n9838), .IN2(g1088), .Q(n15097) );
  INVX0 U15178 ( .INP(n14971), .ZN(n15096) );
  INVX0 U15179 ( .INP(n15101), .ZN(n15093) );
  OR2X1 U15180 ( .IN1(n15036), .IN2(g3229), .Q(n15101) );
  OR2X1 U15181 ( .IN1(n14973), .IN2(n14869), .Q(n15036) );
  OR2X1 U15182 ( .IN1(n15102), .IN2(n15103), .Q(n14869) );
  OR2X1 U15183 ( .IN1(n15104), .IN2(n15105), .Q(n15103) );
  AND2X1 U15184 ( .IN1(n9562), .IN2(g6712), .Q(n15105) );
  AND2X1 U15185 ( .IN1(g5472), .IN2(n10203), .Q(n15104) );
  AND2X1 U15186 ( .IN1(n9563), .IN2(g1088), .Q(n15102) );
  INVX0 U15187 ( .INP(n14867), .ZN(n14973) );
  OR2X1 U15188 ( .IN1(n15106), .IN2(n15107), .Q(n14867) );
  OR2X1 U15189 ( .IN1(n15108), .IN2(n15109), .Q(n15107) );
  AND2X1 U15190 ( .IN1(n9816), .IN2(g6712), .Q(n15109) );
  AND2X1 U15191 ( .IN1(n9817), .IN2(g5472), .Q(n15108) );
  AND2X1 U15192 ( .IN1(n9815), .IN2(g1088), .Q(n15106) );
  AND2X1 U15193 ( .IN1(g3229), .IN2(n14971), .Q(n15091) );
  OR2X1 U15194 ( .IN1(n15110), .IN2(n15111), .Q(n14971) );
  OR2X1 U15195 ( .IN1(n15112), .IN2(n15113), .Q(n15111) );
  AND2X1 U15196 ( .IN1(n9827), .IN2(g6712), .Q(n15113) );
  AND2X1 U15197 ( .IN1(n9828), .IN2(g5472), .Q(n15112) );
  AND2X1 U15198 ( .IN1(n9826), .IN2(g1088), .Q(n15110) );
  AND2X1 U15199 ( .IN1(n14871), .IN2(g1041), .Q(n15088) );
  INVX0 U15200 ( .INP(n14866), .ZN(n14871) );
  AND2X1 U15201 ( .IN1(g5472), .IN2(n14981), .Q(n14866) );
  INVX0 U15202 ( .INP(n15114), .ZN(n14981) );
  OR2X1 U15203 ( .IN1(n15115), .IN2(n10737), .Q(n15114) );
  AND2X1 U15204 ( .IN1(n10672), .IN2(n10742), .Q(n15115) );
  OR2X1 U15205 ( .IN1(n15116), .IN2(n15117), .Q(g27256) );
  AND2X1 U15206 ( .IN1(n15004), .IN2(n14993), .Q(n15117) );
  AND2X1 U15207 ( .IN1(n15118), .IN2(n15119), .Q(n15004) );
  OR2X1 U15208 ( .IN1(n15078), .IN2(n15120), .Q(n15118) );
  INVX0 U15209 ( .INP(n14996), .ZN(n15120) );
  INVX0 U15210 ( .INP(n14997), .ZN(n15078) );
  OR2X1 U15211 ( .IN1(n15121), .IN2(n15122), .Q(n14997) );
  AND2X1 U15212 ( .IN1(n15123), .IN2(n10974), .Q(n15122) );
  INVX0 U15213 ( .INP(n15124), .ZN(n15123) );
  AND2X1 U15214 ( .IN1(g3229), .IN2(n15124), .Q(n15121) );
  INVX0 U15215 ( .INP(n15125), .ZN(n15116) );
  OR2X1 U15216 ( .IN1(n14993), .IN2(n9820), .Q(n15125) );
  OR2X1 U15217 ( .IN1(n15126), .IN2(n15127), .Q(g27255) );
  AND2X1 U15218 ( .IN1(n15086), .IN2(n14894), .Q(n15127) );
  INVX0 U15219 ( .INP(n15128), .ZN(n15126) );
  OR2X1 U15220 ( .IN1(n14894), .IN2(n9841), .Q(n15128) );
  AND2X1 U15221 ( .IN1(g6447), .IN2(n15087), .Q(n14894) );
  OR2X1 U15222 ( .IN1(n15129), .IN2(n15130), .Q(g27253) );
  AND2X1 U15223 ( .IN1(n15086), .IN2(n14993), .Q(n15130) );
  INVX0 U15224 ( .INP(n15131), .ZN(n15086) );
  OR2X1 U15225 ( .IN1(n15132), .IN2(n15133), .Q(n15131) );
  OR2X1 U15226 ( .IN1(n15134), .IN2(n15135), .Q(n15133) );
  AND2X1 U15227 ( .IN1(n15136), .IN2(n15119), .Q(n15135) );
  AND2X1 U15228 ( .IN1(n15137), .IN2(n15124), .Q(n15136) );
  OR2X1 U15229 ( .IN1(n15138), .IN2(n15139), .Q(n15124) );
  OR2X1 U15230 ( .IN1(n15140), .IN2(n15141), .Q(n15139) );
  AND2X1 U15231 ( .IN1(n13375), .IN2(n10204), .Q(n15141) );
  AND2X1 U15232 ( .IN1(n9841), .IN2(n13502), .Q(n15140) );
  AND2X1 U15233 ( .IN1(n9842), .IN2(n13506), .Q(n15138) );
  INVX0 U15234 ( .INP(n15077), .ZN(n15137) );
  INVX0 U15235 ( .INP(n15142), .ZN(n15134) );
  OR2X1 U15236 ( .IN1(n15119), .IN2(g3229), .Q(n15142) );
  OR2X1 U15237 ( .IN1(n15079), .IN2(n14996), .Q(n15119) );
  OR2X1 U15238 ( .IN1(n15143), .IN2(n15144), .Q(n14996) );
  OR2X1 U15239 ( .IN1(n15145), .IN2(n15146), .Q(n15144) );
  AND2X1 U15240 ( .IN1(n9565), .IN2(n13375), .Q(n15146) );
  AND2X1 U15241 ( .IN1(n9566), .IN2(n13502), .Q(n15145) );
  AND2X1 U15242 ( .IN1(n9564), .IN2(n13506), .Q(n15143) );
  INVX0 U15243 ( .INP(n14994), .ZN(n15079) );
  OR2X1 U15244 ( .IN1(n15147), .IN2(n15148), .Q(n14994) );
  OR2X1 U15245 ( .IN1(n15149), .IN2(n15150), .Q(n15148) );
  AND2X1 U15246 ( .IN1(n9818), .IN2(n13375), .Q(n15150) );
  AND2X1 U15247 ( .IN1(n9819), .IN2(n13502), .Q(n15149) );
  AND2X1 U15248 ( .IN1(n9820), .IN2(n13506), .Q(n15147) );
  AND2X1 U15249 ( .IN1(g3229), .IN2(n15077), .Q(n15132) );
  OR2X1 U15250 ( .IN1(n15151), .IN2(n15152), .Q(n15077) );
  OR2X1 U15251 ( .IN1(n15153), .IN2(n15154), .Q(n15152) );
  AND2X1 U15252 ( .IN1(n9829), .IN2(n13375), .Q(n15154) );
  AND2X1 U15253 ( .IN1(n9830), .IN2(n13502), .Q(n15153) );
  AND2X1 U15254 ( .IN1(n9831), .IN2(n13506), .Q(n15151) );
  INVX0 U15255 ( .INP(n15155), .ZN(n15129) );
  OR2X1 U15256 ( .IN1(n14993), .IN2(n9842), .Q(n15155) );
  AND2X1 U15257 ( .IN1(g5437), .IN2(n15087), .Q(n14993) );
  INVX0 U15258 ( .INP(n15156), .ZN(n15087) );
  OR2X1 U15259 ( .IN1(n15157), .IN2(n10671), .Q(n15156) );
  AND2X1 U15260 ( .IN1(n10672), .IN2(n10678), .Q(n15157) );
  AND2X1 U15261 ( .IN1(n15158), .IN2(n15159), .Q(g27243) );
  OR2X1 U15262 ( .IN1(n15160), .IN2(g2753), .Q(n15159) );
  AND2X1 U15263 ( .IN1(test_so92), .IN2(n15161), .Q(n15160) );
  AND2X1 U15264 ( .IN1(n14454), .IN2(n14331), .Q(n15158) );
  OR2X1 U15265 ( .IN1(n10192), .IN2(n15162), .Q(n14454) );
  OR2X1 U15266 ( .IN1(n4471), .IN2(n15163), .Q(n15162) );
  AND2X1 U15267 ( .IN1(n15164), .IN2(n4522), .Q(g27131) );
  AND2X1 U15268 ( .IN1(n15165), .IN2(n12966), .Q(n15164) );
  OR2X1 U15269 ( .IN1(n3683), .IN2(g2147), .Q(n15165) );
  AND2X1 U15270 ( .IN1(n15166), .IN2(n4523), .Q(g27129) );
  AND2X1 U15271 ( .IN1(n15167), .IN2(n12971), .Q(n15166) );
  OR2X1 U15272 ( .IN1(n3686), .IN2(g1453), .Q(n15167) );
  AND2X1 U15273 ( .IN1(n15168), .IN2(n12976), .Q(g27123) );
  AND2X1 U15274 ( .IN1(n15169), .IN2(n882), .Q(n15168) );
  OR2X1 U15275 ( .IN1(n10171), .IN2(n15170), .Q(n882) );
  INVX0 U15276 ( .INP(n3689), .ZN(n15170) );
  OR2X1 U15277 ( .IN1(n3689), .IN2(g767), .Q(n15169) );
  AND2X1 U15278 ( .IN1(n15171), .IN2(n4521), .Q(g27120) );
  AND2X1 U15279 ( .IN1(n15172), .IN2(n12981), .Q(n15171) );
  OR2X1 U15280 ( .IN1(n3692), .IN2(test_so15), .Q(n15172) );
  OR2X1 U15281 ( .IN1(n15173), .IN2(n15174), .Q(g26827) );
  AND2X1 U15282 ( .IN1(n4509), .IN2(g2519), .Q(n15174) );
  AND2X1 U15283 ( .IN1(n15175), .IN2(n4606), .Q(n15173) );
  OR2X1 U15284 ( .IN1(n15176), .IN2(n15177), .Q(g26826) );
  AND2X1 U15285 ( .IN1(n4524), .IN2(g2516), .Q(n15177) );
  AND2X1 U15286 ( .IN1(n15175), .IN2(g7264), .Q(n15176) );
  OR2X1 U15287 ( .IN1(n15178), .IN2(n15179), .Q(g26825) );
  AND2X1 U15288 ( .IN1(n4509), .IN2(g2510), .Q(n15179) );
  AND2X1 U15289 ( .IN1(n4606), .IN2(n15180), .Q(n15178) );
  OR2X1 U15290 ( .IN1(n15181), .IN2(n15182), .Q(g26824) );
  AND2X1 U15291 ( .IN1(test_so59), .IN2(n4511), .Q(n15182) );
  AND2X1 U15292 ( .IN1(n15183), .IN2(n4618), .Q(n15181) );
  OR2X1 U15293 ( .IN1(n15184), .IN2(n15185), .Q(g26823) );
  AND2X1 U15294 ( .IN1(n4516), .IN2(g2513), .Q(n15185) );
  AND2X1 U15295 ( .IN1(n15175), .IN2(g5555), .Q(n15184) );
  AND2X1 U15296 ( .IN1(n15186), .IN2(n15187), .Q(n15175) );
  OR2X1 U15297 ( .IN1(n15188), .IN2(n15189), .Q(n15187) );
  OR2X1 U15298 ( .IN1(n14392), .IN2(n15190), .Q(n15188) );
  INVX0 U15299 ( .INP(n14391), .ZN(n15190) );
  OR2X1 U15300 ( .IN1(n15191), .IN2(n15192), .Q(n15186) );
  AND2X1 U15301 ( .IN1(n14391), .IN2(n15193), .Q(n15192) );
  INVX0 U15302 ( .INP(n14392), .ZN(n15193) );
  OR2X1 U15303 ( .IN1(n10191), .IN2(n15194), .Q(n14392) );
  OR2X1 U15304 ( .IN1(n15195), .IN2(n15196), .Q(n15194) );
  AND2X1 U15305 ( .IN1(n14388), .IN2(n14386), .Q(n15196) );
  OR2X1 U15306 ( .IN1(n15189), .IN2(n15197), .Q(n14386) );
  INVX0 U15307 ( .INP(n15191), .ZN(n15189) );
  INVX0 U15308 ( .INP(n14387), .ZN(n14388) );
  AND2X1 U15309 ( .IN1(n14389), .IN2(n14387), .Q(n15195) );
  OR2X1 U15310 ( .IN1(n15198), .IN2(n15191), .Q(n14389) );
  OR2X1 U15311 ( .IN1(n15199), .IN2(n15200), .Q(n14391) );
  OR2X1 U15312 ( .IN1(n15201), .IN2(n15202), .Q(n15200) );
  AND2X1 U15313 ( .IN1(n9853), .IN2(n13116), .Q(n15202) );
  AND2X1 U15314 ( .IN1(n13101), .IN2(n10208), .Q(n15201) );
  AND2X1 U15315 ( .IN1(n9844), .IN2(n13106), .Q(n15199) );
  OR2X1 U15316 ( .IN1(n15203), .IN2(n15204), .Q(g26822) );
  AND2X1 U15317 ( .IN1(n4524), .IN2(g2507), .Q(n15204) );
  AND2X1 U15318 ( .IN1(g7264), .IN2(n15180), .Q(n15203) );
  OR2X1 U15319 ( .IN1(n15205), .IN2(n15206), .Q(g26821) );
  AND2X1 U15320 ( .IN1(n4525), .IN2(g1822), .Q(n15206) );
  AND2X1 U15321 ( .IN1(n15183), .IN2(g7014), .Q(n15205) );
  OR2X1 U15322 ( .IN1(n15207), .IN2(n15208), .Q(g26820) );
  AND2X1 U15323 ( .IN1(n4511), .IN2(g1816), .Q(n15208) );
  AND2X1 U15324 ( .IN1(n4618), .IN2(n15209), .Q(n15207) );
  OR2X1 U15325 ( .IN1(n15210), .IN2(n15211), .Q(g26818) );
  AND2X1 U15326 ( .IN1(n15212), .IN2(g1088), .Q(n15211) );
  AND2X1 U15327 ( .IN1(n4381), .IN2(g1131), .Q(n15210) );
  OR2X1 U15328 ( .IN1(n15213), .IN2(n15214), .Q(g26817) );
  AND2X1 U15329 ( .IN1(n4516), .IN2(g2504), .Q(n15214) );
  AND2X1 U15330 ( .IN1(g5555), .IN2(n15180), .Q(n15213) );
  OR2X1 U15331 ( .IN1(n15215), .IN2(n15216), .Q(n15180) );
  AND2X1 U15332 ( .IN1(n14387), .IN2(n10191), .Q(n15216) );
  OR2X1 U15333 ( .IN1(n15217), .IN2(n15218), .Q(n14387) );
  OR2X1 U15334 ( .IN1(n15219), .IN2(n15220), .Q(n15218) );
  AND2X1 U15335 ( .IN1(g7264), .IN2(g2507), .Q(n15220) );
  AND2X1 U15336 ( .IN1(n4606), .IN2(g2510), .Q(n15219) );
  AND2X1 U15337 ( .IN1(g5555), .IN2(g2504), .Q(n15217) );
  AND2X1 U15338 ( .IN1(n15197), .IN2(test_so79), .Q(n15215) );
  INVX0 U15339 ( .INP(n15198), .ZN(n15197) );
  OR2X1 U15340 ( .IN1(n15221), .IN2(n13687), .Q(n15198) );
  AND2X1 U15341 ( .IN1(n15222), .IN2(n15223), .Q(n15221) );
  OR2X1 U15342 ( .IN1(n4324), .IN2(g2254), .Q(n15223) );
  AND2X1 U15343 ( .IN1(n15224), .IN2(n15225), .Q(n15222) );
  OR2X1 U15344 ( .IN1(n10189), .IN2(g2255), .Q(n15225) );
  OR2X1 U15345 ( .IN1(n4367), .IN2(g2253), .Q(n15224) );
  OR2X1 U15346 ( .IN1(n15226), .IN2(n15227), .Q(g26816) );
  AND2X1 U15347 ( .IN1(n4518), .IN2(g1819), .Q(n15227) );
  AND2X1 U15348 ( .IN1(n15183), .IN2(g5511), .Q(n15226) );
  AND2X1 U15349 ( .IN1(n15228), .IN2(n15229), .Q(n15183) );
  OR2X1 U15350 ( .IN1(n15230), .IN2(n15231), .Q(n15229) );
  OR2X1 U15351 ( .IN1(n14413), .IN2(n15232), .Q(n15230) );
  INVX0 U15352 ( .INP(n14412), .ZN(n15232) );
  OR2X1 U15353 ( .IN1(n15233), .IN2(n15234), .Q(n15228) );
  AND2X1 U15354 ( .IN1(n14412), .IN2(n15235), .Q(n15234) );
  INVX0 U15355 ( .INP(n14413), .ZN(n15235) );
  OR2X1 U15356 ( .IN1(n4386), .IN2(n15236), .Q(n14413) );
  OR2X1 U15357 ( .IN1(n15237), .IN2(n15238), .Q(n15236) );
  AND2X1 U15358 ( .IN1(n14409), .IN2(n14407), .Q(n15238) );
  OR2X1 U15359 ( .IN1(n15231), .IN2(n15239), .Q(n14407) );
  INVX0 U15360 ( .INP(n15233), .ZN(n15231) );
  INVX0 U15361 ( .INP(n14408), .ZN(n14409) );
  AND2X1 U15362 ( .IN1(n14410), .IN2(n14408), .Q(n15237) );
  OR2X1 U15363 ( .IN1(n15240), .IN2(n15233), .Q(n14410) );
  OR2X1 U15364 ( .IN1(n15241), .IN2(n15242), .Q(n14412) );
  OR2X1 U15365 ( .IN1(n15243), .IN2(n15244), .Q(n15242) );
  AND2X1 U15366 ( .IN1(n9858), .IN2(n13248), .Q(n15244) );
  AND2X1 U15367 ( .IN1(n9857), .IN2(n13111), .Q(n15243) );
  AND2X1 U15368 ( .IN1(n9847), .IN2(n13239), .Q(n15241) );
  OR2X1 U15369 ( .IN1(n15245), .IN2(n15246), .Q(g26815) );
  AND2X1 U15370 ( .IN1(n4525), .IN2(g1813), .Q(n15246) );
  AND2X1 U15371 ( .IN1(g7014), .IN2(n15209), .Q(n15245) );
  OR2X1 U15372 ( .IN1(n15247), .IN2(n15248), .Q(g26814) );
  AND2X1 U15373 ( .IN1(n15212), .IN2(g6712), .Q(n15248) );
  AND2X1 U15374 ( .IN1(n4364), .IN2(g1128), .Q(n15247) );
  OR2X1 U15375 ( .IN1(n15249), .IN2(n15250), .Q(g26813) );
  AND2X1 U15376 ( .IN1(n15251), .IN2(g1088), .Q(n15250) );
  AND2X1 U15377 ( .IN1(n4381), .IN2(g1122), .Q(n15249) );
  OR2X1 U15378 ( .IN1(n15252), .IN2(n15253), .Q(g26812) );
  AND2X1 U15379 ( .IN1(n4506), .IN2(g444), .Q(n15253) );
  AND2X1 U15380 ( .IN1(n15254), .IN2(n4640), .Q(n15252) );
  OR2X1 U15381 ( .IN1(n15255), .IN2(n15256), .Q(g26811) );
  AND2X1 U15382 ( .IN1(n4518), .IN2(g1810), .Q(n15256) );
  AND2X1 U15383 ( .IN1(g5511), .IN2(n15209), .Q(n15255) );
  OR2X1 U15384 ( .IN1(n15257), .IN2(n15258), .Q(n15209) );
  AND2X1 U15385 ( .IN1(n4386), .IN2(n14408), .Q(n15258) );
  OR2X1 U15386 ( .IN1(n15259), .IN2(n15260), .Q(n14408) );
  OR2X1 U15387 ( .IN1(n15261), .IN2(n15262), .Q(n15260) );
  AND2X1 U15388 ( .IN1(g7014), .IN2(g1813), .Q(n15262) );
  AND2X1 U15389 ( .IN1(n4618), .IN2(g1816), .Q(n15261) );
  AND2X1 U15390 ( .IN1(g5511), .IN2(g1810), .Q(n15259) );
  AND2X1 U15391 ( .IN1(n15239), .IN2(g1690), .Q(n15257) );
  INVX0 U15392 ( .INP(n15240), .ZN(n15239) );
  OR2X1 U15393 ( .IN1(n15263), .IN2(n13731), .Q(n15240) );
  AND2X1 U15394 ( .IN1(n15264), .IN2(n15265), .Q(n15263) );
  OR2X1 U15395 ( .IN1(n4317), .IN2(g1560), .Q(n15265) );
  AND2X1 U15396 ( .IN1(n15266), .IN2(n15267), .Q(n15264) );
  OR2X1 U15397 ( .IN1(n4515), .IN2(g1561), .Q(n15267) );
  OR2X1 U15398 ( .IN1(n4368), .IN2(g1559), .Q(n15266) );
  OR2X1 U15399 ( .IN1(n15268), .IN2(n15269), .Q(g26810) );
  AND2X1 U15400 ( .IN1(n15212), .IN2(g5472), .Q(n15269) );
  AND2X1 U15401 ( .IN1(n15270), .IN2(n15271), .Q(n15212) );
  OR2X1 U15402 ( .IN1(n15272), .IN2(n15273), .Q(n15271) );
  OR2X1 U15403 ( .IN1(n14434), .IN2(n15274), .Q(n15272) );
  INVX0 U15404 ( .INP(n14433), .ZN(n15274) );
  OR2X1 U15405 ( .IN1(n15275), .IN2(n15276), .Q(n15270) );
  AND2X1 U15406 ( .IN1(n14433), .IN2(n15277), .Q(n15276) );
  INVX0 U15407 ( .INP(n14434), .ZN(n15277) );
  OR2X1 U15408 ( .IN1(n4387), .IN2(n15278), .Q(n14434) );
  OR2X1 U15409 ( .IN1(n15279), .IN2(n15280), .Q(n15278) );
  AND2X1 U15410 ( .IN1(n14430), .IN2(n14428), .Q(n15280) );
  OR2X1 U15411 ( .IN1(n15273), .IN2(n15281), .Q(n14428) );
  INVX0 U15412 ( .INP(n15275), .ZN(n15273) );
  INVX0 U15413 ( .INP(n14429), .ZN(n14430) );
  AND2X1 U15414 ( .IN1(n14431), .IN2(n14429), .Q(n15279) );
  OR2X1 U15415 ( .IN1(n15282), .IN2(n15275), .Q(n14431) );
  OR2X1 U15416 ( .IN1(n15283), .IN2(n15284), .Q(n14433) );
  OR2X1 U15417 ( .IN1(n15285), .IN2(n15286), .Q(n15284) );
  AND2X1 U15418 ( .IN1(n9850), .IN2(g6712), .Q(n15286) );
  AND2X1 U15419 ( .IN1(n9864), .IN2(g5472), .Q(n15285) );
  AND2X1 U15420 ( .IN1(n9863), .IN2(g1088), .Q(n15283) );
  AND2X1 U15421 ( .IN1(n4363), .IN2(g1125), .Q(n15268) );
  OR2X1 U15422 ( .IN1(n15287), .IN2(n15288), .Q(g26809) );
  AND2X1 U15423 ( .IN1(n4364), .IN2(test_so38), .Q(n15288) );
  AND2X1 U15424 ( .IN1(n15251), .IN2(g6712), .Q(n15287) );
  OR2X1 U15425 ( .IN1(n15289), .IN2(n15290), .Q(g26808) );
  AND2X1 U15426 ( .IN1(n4499), .IN2(g441), .Q(n15290) );
  AND2X1 U15427 ( .IN1(n15254), .IN2(g6447), .Q(n15289) );
  OR2X1 U15428 ( .IN1(n15291), .IN2(n15292), .Q(g26807) );
  AND2X1 U15429 ( .IN1(n4506), .IN2(g435), .Q(n15292) );
  AND2X1 U15430 ( .IN1(n4640), .IN2(n15293), .Q(n15291) );
  OR2X1 U15431 ( .IN1(n15294), .IN2(n15295), .Q(g26806) );
  AND2X1 U15432 ( .IN1(n15251), .IN2(g5472), .Q(n15295) );
  OR2X1 U15433 ( .IN1(n15296), .IN2(n15297), .Q(n15251) );
  AND2X1 U15434 ( .IN1(n4387), .IN2(n14429), .Q(n15297) );
  OR2X1 U15435 ( .IN1(n15298), .IN2(n15299), .Q(n14429) );
  OR2X1 U15436 ( .IN1(n15300), .IN2(n15301), .Q(n15299) );
  AND2X1 U15437 ( .IN1(test_so38), .IN2(g6712), .Q(n15301) );
  AND2X1 U15438 ( .IN1(g5472), .IN2(g1116), .Q(n15300) );
  AND2X1 U15439 ( .IN1(g1088), .IN2(g1122), .Q(n15298) );
  AND2X1 U15440 ( .IN1(n15281), .IN2(g996), .Q(n15296) );
  INVX0 U15441 ( .INP(n15282), .ZN(n15281) );
  OR2X1 U15442 ( .IN1(n15302), .IN2(n13770), .Q(n15282) );
  AND2X1 U15443 ( .IN1(n15303), .IN2(n15304), .Q(n15302) );
  OR2X1 U15444 ( .IN1(n4312), .IN2(g867), .Q(n15304) );
  AND2X1 U15445 ( .IN1(n15305), .IN2(n15306), .Q(n15303) );
  OR2X1 U15446 ( .IN1(n10188), .IN2(g865), .Q(n15306) );
  OR2X1 U15447 ( .IN1(n4323), .IN2(g866), .Q(n15305) );
  AND2X1 U15448 ( .IN1(n4363), .IN2(g1116), .Q(n15294) );
  OR2X1 U15449 ( .IN1(n15307), .IN2(n15308), .Q(g26805) );
  AND2X1 U15450 ( .IN1(n4520), .IN2(g438), .Q(n15308) );
  AND2X1 U15451 ( .IN1(n15254), .IN2(g5437), .Q(n15307) );
  AND2X1 U15452 ( .IN1(n15309), .IN2(n15310), .Q(n15254) );
  OR2X1 U15453 ( .IN1(n15311), .IN2(n15312), .Q(n15310) );
  OR2X1 U15454 ( .IN1(n14450), .IN2(n15313), .Q(n15311) );
  INVX0 U15455 ( .INP(n14449), .ZN(n15313) );
  OR2X1 U15456 ( .IN1(n15314), .IN2(n15315), .Q(n15309) );
  AND2X1 U15457 ( .IN1(n14449), .IN2(n15316), .Q(n15315) );
  INVX0 U15458 ( .INP(n14450), .ZN(n15316) );
  OR2X1 U15459 ( .IN1(n4388), .IN2(n15317), .Q(n14450) );
  OR2X1 U15460 ( .IN1(n15318), .IN2(n15319), .Q(n15317) );
  AND2X1 U15461 ( .IN1(n14446), .IN2(n14444), .Q(n15319) );
  OR2X1 U15462 ( .IN1(n15312), .IN2(n15320), .Q(n14444) );
  INVX0 U15463 ( .INP(n15314), .ZN(n15312) );
  INVX0 U15464 ( .INP(n14445), .ZN(n14446) );
  AND2X1 U15465 ( .IN1(n14447), .IN2(n14445), .Q(n15318) );
  OR2X1 U15466 ( .IN1(n15321), .IN2(n15314), .Q(n14447) );
  OR2X1 U15467 ( .IN1(n15322), .IN2(n15323), .Q(n14449) );
  OR2X1 U15468 ( .IN1(n15324), .IN2(n15325), .Q(n15323) );
  AND2X1 U15469 ( .IN1(n9870), .IN2(n13375), .Q(n15325) );
  AND2X1 U15470 ( .IN1(n9871), .IN2(n13502), .Q(n15324) );
  AND2X1 U15471 ( .IN1(n9872), .IN2(n13506), .Q(n15322) );
  OR2X1 U15472 ( .IN1(n15326), .IN2(n15327), .Q(g26804) );
  AND2X1 U15473 ( .IN1(n4499), .IN2(g432), .Q(n15327) );
  AND2X1 U15474 ( .IN1(g6447), .IN2(n15293), .Q(n15326) );
  OR2X1 U15475 ( .IN1(n15328), .IN2(n15329), .Q(g26803) );
  AND2X1 U15476 ( .IN1(n4520), .IN2(g429), .Q(n15329) );
  AND2X1 U15477 ( .IN1(g5437), .IN2(n15293), .Q(n15328) );
  OR2X1 U15478 ( .IN1(n15330), .IN2(n15331), .Q(n15293) );
  AND2X1 U15479 ( .IN1(n4388), .IN2(n14445), .Q(n15331) );
  OR2X1 U15480 ( .IN1(n15332), .IN2(n15333), .Q(n14445) );
  OR2X1 U15481 ( .IN1(n15334), .IN2(n15335), .Q(n15333) );
  AND2X1 U15482 ( .IN1(g6447), .IN2(g432), .Q(n15335) );
  AND2X1 U15483 ( .IN1(n4640), .IN2(g435), .Q(n15334) );
  AND2X1 U15484 ( .IN1(g5437), .IN2(g429), .Q(n15332) );
  AND2X1 U15485 ( .IN1(n15320), .IN2(g309), .Q(n15330) );
  INVX0 U15486 ( .INP(n15321), .ZN(n15320) );
  OR2X1 U15487 ( .IN1(n15336), .IN2(n13801), .Q(n15321) );
  AND2X1 U15488 ( .IN1(n15337), .IN2(n15338), .Q(n15336) );
  OR2X1 U15489 ( .IN1(n4318), .IN2(g178), .Q(n15338) );
  AND2X1 U15490 ( .IN1(n15339), .IN2(n15340), .Q(n15337) );
  OR2X1 U15491 ( .IN1(n4512), .IN2(g179), .Q(n15340) );
  OR2X1 U15492 ( .IN1(n4369), .IN2(g177), .Q(n15339) );
  AND2X1 U15493 ( .IN1(n15341), .IN2(n11730), .Q(g26798) );
  AND2X1 U15494 ( .IN1(n15342), .IN2(n15343), .Q(n15341) );
  INVX0 U15495 ( .INP(n15344), .ZN(n15343) );
  AND2X1 U15496 ( .IN1(n15345), .IN2(n4355), .Q(n15344) );
  OR2X1 U15497 ( .IN1(n4355), .IN2(n15345), .Q(n15342) );
  AND2X1 U15498 ( .IN1(n15346), .IN2(n14331), .Q(g26795) );
  OR2X1 U15499 ( .IN1(n15347), .IN2(n15348), .Q(n15346) );
  AND2X1 U15500 ( .IN1(n15161), .IN2(n10192), .Q(n15348) );
  INVX0 U15501 ( .INP(n15163), .ZN(n15161) );
  AND2X1 U15502 ( .IN1(test_so92), .IN2(n15163), .Q(n15347) );
  AND2X1 U15503 ( .IN1(n15349), .IN2(n14337), .Q(g26789) );
  AND2X1 U15504 ( .IN1(n15350), .IN2(n15351), .Q(n15349) );
  OR2X1 U15505 ( .IN1(n14464), .IN2(g2046), .Q(n15351) );
  INVX0 U15506 ( .INP(n14465), .ZN(n14464) );
  OR2X1 U15507 ( .IN1(n4468), .IN2(n14465), .Q(n15350) );
  AND2X1 U15508 ( .IN1(n15352), .IN2(n15353), .Q(g26786) );
  OR2X1 U15509 ( .IN1(n15354), .IN2(n15355), .Q(n15353) );
  INVX0 U15510 ( .INP(n15356), .ZN(n15355) );
  OR2X1 U15511 ( .IN1(n15357), .IN2(n9351), .Q(n15356) );
  AND2X1 U15512 ( .IN1(n9351), .IN2(n15357), .Q(n15354) );
  INVX0 U15513 ( .INP(n3741), .ZN(n15357) );
  AND2X1 U15514 ( .IN1(n15358), .IN2(n14345), .Q(g26781) );
  AND2X1 U15515 ( .IN1(n15359), .IN2(n15360), .Q(n15358) );
  OR2X1 U15516 ( .IN1(n14470), .IN2(g1352), .Q(n15360) );
  INVX0 U15517 ( .INP(n14471), .ZN(n14470) );
  OR2X1 U15518 ( .IN1(n4469), .IN2(n14471), .Q(n15359) );
  AND2X1 U15519 ( .IN1(n15361), .IN2(n13809), .Q(g26776) );
  OR2X1 U15520 ( .IN1(n15362), .IN2(n15363), .Q(n15361) );
  AND2X1 U15521 ( .IN1(n14476), .IN2(n10193), .Q(n15363) );
  INVX0 U15522 ( .INP(n14478), .ZN(n14476) );
  AND2X1 U15523 ( .IN1(test_so28), .IN2(n14478), .Q(n15362) );
  AND2X1 U15524 ( .IN1(n15364), .IN2(n15365), .Q(g26677) );
  OR2X1 U15525 ( .IN1(n15366), .IN2(g2746), .Q(n15365) );
  AND2X1 U15526 ( .IN1(n15367), .IN2(g2734), .Q(n15366) );
  AND2X1 U15527 ( .IN1(n14331), .IN2(n15163), .Q(n15364) );
  OR2X1 U15528 ( .IN1(n15368), .IN2(n15369), .Q(n15163) );
  OR2X1 U15529 ( .IN1(n4407), .IN2(n4397), .Q(n15369) );
  OR2X1 U15530 ( .IN1(n15370), .IN2(n15371), .Q(g26676) );
  AND2X1 U15531 ( .IN1(n15372), .IN2(n13106), .Q(n15371) );
  AND2X1 U15532 ( .IN1(n15373), .IN2(g2479), .Q(n15370) );
  OR2X1 U15533 ( .IN1(n4524), .IN2(n15374), .Q(n15373) );
  OR2X1 U15534 ( .IN1(n15375), .IN2(n15376), .Q(g26675) );
  AND2X1 U15535 ( .IN1(n15377), .IN2(n13111), .Q(n15376) );
  AND2X1 U15536 ( .IN1(n15378), .IN2(g1783), .Q(n15375) );
  OR2X1 U15537 ( .IN1(n4511), .IN2(n15379), .Q(n15378) );
  OR2X1 U15538 ( .IN1(n15380), .IN2(n15381), .Q(g26672) );
  AND2X1 U15539 ( .IN1(n15372), .IN2(n13116), .Q(n15381) );
  AND2X1 U15540 ( .IN1(n15382), .IN2(g2478), .Q(n15380) );
  OR2X1 U15541 ( .IN1(n4516), .IN2(n15374), .Q(n15382) );
  AND2X1 U15542 ( .IN1(n15383), .IN2(n15384), .Q(g26671) );
  OR2X1 U15543 ( .IN1(n15385), .IN2(g2052), .Q(n15384) );
  AND2X1 U15544 ( .IN1(n15386), .IN2(g2040), .Q(n15385) );
  AND2X1 U15545 ( .IN1(n14465), .IN2(n14337), .Q(n15383) );
  OR2X1 U15546 ( .IN1(n15387), .IN2(n15388), .Q(n14465) );
  OR2X1 U15547 ( .IN1(n4409), .IN2(n4399), .Q(n15388) );
  OR2X1 U15548 ( .IN1(n15389), .IN2(n15390), .Q(g26670) );
  AND2X1 U15549 ( .IN1(n15377), .IN2(n13239), .Q(n15390) );
  AND2X1 U15550 ( .IN1(n15391), .IN2(g1785), .Q(n15389) );
  OR2X1 U15551 ( .IN1(n4525), .IN2(n15379), .Q(n15391) );
  OR2X1 U15552 ( .IN1(n15392), .IN2(n15393), .Q(g26669) );
  AND2X1 U15553 ( .IN1(n15394), .IN2(g1088), .Q(n15393) );
  AND2X1 U15554 ( .IN1(n15395), .IN2(g1089), .Q(n15392) );
  OR2X1 U15555 ( .IN1(n4381), .IN2(n15396), .Q(n15395) );
  OR2X1 U15556 ( .IN1(n15397), .IN2(n15398), .Q(g26667) );
  AND2X1 U15557 ( .IN1(n15377), .IN2(n13248), .Q(n15398) );
  AND2X1 U15558 ( .IN1(g1690), .IN2(n15379), .Q(n15377) );
  AND2X1 U15559 ( .IN1(test_so60), .IN2(n15399), .Q(n15397) );
  OR2X1 U15560 ( .IN1(n4518), .IN2(n15379), .Q(n15399) );
  OR2X1 U15561 ( .IN1(n12938), .IN2(n15400), .Q(n15379) );
  OR2X1 U15562 ( .IN1(n4386), .IN2(n12695), .Q(n15400) );
  OR2X1 U15563 ( .IN1(n15401), .IN2(n15402), .Q(n12695) );
  OR2X1 U15564 ( .IN1(n15403), .IN2(n15404), .Q(n15402) );
  OR2X1 U15565 ( .IN1(n15405), .IN2(n15406), .Q(n15404) );
  OR2X1 U15566 ( .IN1(n15407), .IN2(n15408), .Q(n15406) );
  AND2X1 U15567 ( .IN1(n15409), .IN2(n12135), .Q(n15408) );
  INVX0 U15568 ( .INP(n15410), .ZN(n15409) );
  AND2X1 U15569 ( .IN1(n13311), .IN2(n15410), .Q(n15407) );
  OR2X1 U15570 ( .IN1(n15411), .IN2(n15412), .Q(n15410) );
  OR2X1 U15571 ( .IN1(n15413), .IN2(n15414), .Q(n15412) );
  AND2X1 U15572 ( .IN1(n9689), .IN2(g1547), .Q(n15414) );
  AND2X1 U15573 ( .IN1(n9691), .IN2(g6573), .Q(n15413) );
  AND2X1 U15574 ( .IN1(n9690), .IN2(g6782), .Q(n15411) );
  OR2X1 U15575 ( .IN1(n15415), .IN2(n15416), .Q(n15405) );
  AND2X1 U15576 ( .IN1(n15417), .IN2(g1481), .Q(n15416) );
  INVX0 U15577 ( .INP(n15418), .ZN(n15417) );
  AND2X1 U15578 ( .IN1(n4320), .IN2(n15418), .Q(n15415) );
  OR2X1 U15579 ( .IN1(n15419), .IN2(n15420), .Q(n15418) );
  OR2X1 U15580 ( .IN1(n15421), .IN2(n15422), .Q(n15420) );
  AND2X1 U15581 ( .IN1(n10078), .IN2(g6573), .Q(n15422) );
  AND2X1 U15582 ( .IN1(n10077), .IN2(g6782), .Q(n15421) );
  AND2X1 U15583 ( .IN1(n9713), .IN2(g1547), .Q(n15419) );
  OR2X1 U15584 ( .IN1(n15423), .IN2(n15424), .Q(n15403) );
  OR2X1 U15585 ( .IN1(n15425), .IN2(n15426), .Q(n15424) );
  OR2X1 U15586 ( .IN1(n15427), .IN2(n15428), .Q(n15426) );
  AND2X1 U15587 ( .IN1(n15429), .IN2(g1471), .Q(n15428) );
  INVX0 U15588 ( .INP(n15430), .ZN(n15429) );
  AND2X1 U15589 ( .IN1(n4378), .IN2(n15430), .Q(n15427) );
  OR2X1 U15590 ( .IN1(n15431), .IN2(n15432), .Q(n15430) );
  OR2X1 U15591 ( .IN1(n15433), .IN2(n15434), .Q(n15432) );
  AND2X1 U15592 ( .IN1(n10081), .IN2(g6573), .Q(n15434) );
  AND2X1 U15593 ( .IN1(n10080), .IN2(g6782), .Q(n15433) );
  AND2X1 U15594 ( .IN1(n9715), .IN2(g1547), .Q(n15431) );
  OR2X1 U15595 ( .IN1(n15435), .IN2(n15436), .Q(n15425) );
  AND2X1 U15596 ( .IN1(n15437), .IN2(g1476), .Q(n15436) );
  INVX0 U15597 ( .INP(n15438), .ZN(n15437) );
  AND2X1 U15598 ( .IN1(n4374), .IN2(n15438), .Q(n15435) );
  OR2X1 U15599 ( .IN1(n15439), .IN2(n15440), .Q(n15438) );
  OR2X1 U15600 ( .IN1(n15441), .IN2(n15442), .Q(n15440) );
  AND2X1 U15601 ( .IN1(g6573), .IN2(n10209), .Q(n15442) );
  AND2X1 U15602 ( .IN1(n10079), .IN2(g6782), .Q(n15441) );
  AND2X1 U15603 ( .IN1(n9714), .IN2(g1547), .Q(n15439) );
  OR2X1 U15604 ( .IN1(n15443), .IN2(n15444), .Q(n15423) );
  AND2X1 U15605 ( .IN1(n15445), .IN2(n13338), .Q(n15444) );
  INVX0 U15606 ( .INP(n15446), .ZN(n15445) );
  AND2X1 U15607 ( .IN1(n11936), .IN2(n15446), .Q(n15443) );
  OR2X1 U15608 ( .IN1(n15447), .IN2(n15448), .Q(n15446) );
  OR2X1 U15609 ( .IN1(n15449), .IN2(n15450), .Q(n15448) );
  AND2X1 U15610 ( .IN1(n9705), .IN2(g1547), .Q(n15450) );
  AND2X1 U15611 ( .IN1(n9707), .IN2(g6573), .Q(n15449) );
  AND2X1 U15612 ( .IN1(n9706), .IN2(g6782), .Q(n15447) );
  OR2X1 U15613 ( .IN1(n15451), .IN2(n15452), .Q(n15401) );
  OR2X1 U15614 ( .IN1(n15453), .IN2(n15454), .Q(n15452) );
  OR2X1 U15615 ( .IN1(n15455), .IN2(n15456), .Q(n15454) );
  OR2X1 U15616 ( .IN1(n15457), .IN2(n15458), .Q(n15456) );
  AND2X1 U15617 ( .IN1(n15459), .IN2(g1501), .Q(n15458) );
  INVX0 U15618 ( .INP(n15460), .ZN(n15459) );
  AND2X1 U15619 ( .IN1(n4565), .IN2(n15460), .Q(n15457) );
  OR2X1 U15620 ( .IN1(n15461), .IN2(n15462), .Q(n15460) );
  OR2X1 U15621 ( .IN1(n15463), .IN2(n15464), .Q(n15462) );
  AND2X1 U15622 ( .IN1(n9709), .IN2(g1547), .Q(n15464) );
  AND2X1 U15623 ( .IN1(n10070), .IN2(g6573), .Q(n15463) );
  AND2X1 U15624 ( .IN1(g6782), .IN2(n10210), .Q(n15461) );
  OR2X1 U15625 ( .IN1(n15465), .IN2(n15466), .Q(n15455) );
  AND2X1 U15626 ( .IN1(n15467), .IN2(g1496), .Q(n15466) );
  INVX0 U15627 ( .INP(n15468), .ZN(n15467) );
  AND2X1 U15628 ( .IN1(n4557), .IN2(n15468), .Q(n15465) );
  OR2X1 U15629 ( .IN1(n15469), .IN2(n15470), .Q(n15468) );
  OR2X1 U15630 ( .IN1(n15471), .IN2(n15472), .Q(n15470) );
  AND2X1 U15631 ( .IN1(n10072), .IN2(g6573), .Q(n15472) );
  AND2X1 U15632 ( .IN1(n10071), .IN2(g6782), .Q(n15471) );
  AND2X1 U15633 ( .IN1(n9710), .IN2(g1547), .Q(n15469) );
  OR2X1 U15634 ( .IN1(n15473), .IN2(n15474), .Q(n15453) );
  AND2X1 U15635 ( .IN1(n15475), .IN2(g1486), .Q(n15474) );
  INVX0 U15636 ( .INP(n15476), .ZN(n15475) );
  AND2X1 U15637 ( .IN1(n4390), .IN2(n15476), .Q(n15473) );
  OR2X1 U15638 ( .IN1(n15477), .IN2(n15478), .Q(n15476) );
  OR2X1 U15639 ( .IN1(n15479), .IN2(n15480), .Q(n15478) );
  AND2X1 U15640 ( .IN1(n10076), .IN2(g6573), .Q(n15480) );
  AND2X1 U15641 ( .IN1(n10075), .IN2(g6782), .Q(n15479) );
  AND2X1 U15642 ( .IN1(n9712), .IN2(g1547), .Q(n15477) );
  OR2X1 U15643 ( .IN1(n15481), .IN2(n15482), .Q(n15451) );
  OR2X1 U15644 ( .IN1(n11785), .IN2(n15483), .Q(n15482) );
  OR2X1 U15645 ( .IN1(n15484), .IN2(n15485), .Q(n15483) );
  AND2X1 U15646 ( .IN1(n15486), .IN2(g1506), .Q(n15485) );
  INVX0 U15647 ( .INP(n15487), .ZN(n15486) );
  AND2X1 U15648 ( .IN1(n4288), .IN2(n15487), .Q(n15484) );
  OR2X1 U15649 ( .IN1(n15488), .IN2(n15489), .Q(n15487) );
  OR2X1 U15650 ( .IN1(n15490), .IN2(n15491), .Q(n15489) );
  AND2X1 U15651 ( .IN1(n10069), .IN2(g6573), .Q(n15491) );
  AND2X1 U15652 ( .IN1(n10068), .IN2(g6782), .Q(n15490) );
  AND2X1 U15653 ( .IN1(n9708), .IN2(g1547), .Q(n15488) );
  INVX0 U15654 ( .INP(n3070), .ZN(n11785) );
  OR2X1 U15655 ( .IN1(n15492), .IN2(n15493), .Q(n15481) );
  AND2X1 U15656 ( .IN1(n15494), .IN2(g1491), .Q(n15493) );
  INVX0 U15657 ( .INP(n15495), .ZN(n15494) );
  AND2X1 U15658 ( .IN1(n4326), .IN2(n15495), .Q(n15492) );
  OR2X1 U15659 ( .IN1(n15496), .IN2(n15497), .Q(n15495) );
  OR2X1 U15660 ( .IN1(n15498), .IN2(n15499), .Q(n15497) );
  AND2X1 U15661 ( .IN1(n10074), .IN2(g6573), .Q(n15499) );
  AND2X1 U15662 ( .IN1(n10073), .IN2(g6782), .Q(n15498) );
  AND2X1 U15663 ( .IN1(n9711), .IN2(g1547), .Q(n15496) );
  OR2X1 U15664 ( .IN1(n15500), .IN2(n15501), .Q(n12938) );
  OR2X1 U15665 ( .IN1(n15502), .IN2(n15503), .Q(n15501) );
  AND2X1 U15666 ( .IN1(n13248), .IN2(n10211), .Q(n15503) );
  AND2X1 U15667 ( .IN1(n9856), .IN2(n13111), .Q(n15502) );
  AND2X1 U15668 ( .IN1(n9846), .IN2(n13239), .Q(n15500) );
  AND2X1 U15669 ( .IN1(n15504), .IN2(n15505), .Q(g26666) );
  OR2X1 U15670 ( .IN1(n15506), .IN2(g1358), .Q(n15505) );
  AND2X1 U15671 ( .IN1(n15507), .IN2(g1346), .Q(n15506) );
  AND2X1 U15672 ( .IN1(n14471), .IN2(n14345), .Q(n15504) );
  OR2X1 U15673 ( .IN1(n15508), .IN2(n15509), .Q(n14471) );
  OR2X1 U15674 ( .IN1(n4411), .IN2(n4401), .Q(n15509) );
  OR2X1 U15675 ( .IN1(n15510), .IN2(n15511), .Q(g26665) );
  AND2X1 U15676 ( .IN1(n15394), .IN2(g6712), .Q(n15511) );
  AND2X1 U15677 ( .IN1(n15512), .IN2(g1091), .Q(n15510) );
  OR2X1 U15678 ( .IN1(n4364), .IN2(n15396), .Q(n15512) );
  OR2X1 U15679 ( .IN1(n15513), .IN2(n15514), .Q(g26664) );
  AND2X1 U15680 ( .IN1(n15515), .IN2(n13375), .Q(n15514) );
  AND2X1 U15681 ( .IN1(n15516), .IN2(g402), .Q(n15513) );
  OR2X1 U15682 ( .IN1(n4506), .IN2(n15517), .Q(n15516) );
  OR2X1 U15683 ( .IN1(n15518), .IN2(n15519), .Q(g26661) );
  AND2X1 U15684 ( .IN1(n15394), .IN2(g5472), .Q(n15519) );
  AND2X1 U15685 ( .IN1(g996), .IN2(n15396), .Q(n15394) );
  AND2X1 U15686 ( .IN1(n15520), .IN2(g1090), .Q(n15518) );
  OR2X1 U15687 ( .IN1(n4363), .IN2(n15396), .Q(n15520) );
  OR2X1 U15688 ( .IN1(n12950), .IN2(n15521), .Q(n15396) );
  OR2X1 U15689 ( .IN1(n4387), .IN2(n12756), .Q(n15521) );
  OR2X1 U15690 ( .IN1(n15522), .IN2(n15523), .Q(n12756) );
  OR2X1 U15691 ( .IN1(n15524), .IN2(n15525), .Q(n15523) );
  OR2X1 U15692 ( .IN1(n15526), .IN2(n15527), .Q(n15525) );
  OR2X1 U15693 ( .IN1(n15528), .IN2(n15529), .Q(n15527) );
  AND2X1 U15694 ( .IN1(n15530), .IN2(n12190), .Q(n15529) );
  INVX0 U15695 ( .INP(n15531), .ZN(n15530) );
  AND2X1 U15696 ( .IN1(n13470), .IN2(n15531), .Q(n15528) );
  OR2X1 U15697 ( .IN1(n15532), .IN2(n15533), .Q(n15531) );
  OR2X1 U15698 ( .IN1(n15534), .IN2(n15535), .Q(n15533) );
  AND2X1 U15699 ( .IN1(n9721), .IN2(g6368), .Q(n15535) );
  AND2X1 U15700 ( .IN1(n9720), .IN2(g6518), .Q(n15534) );
  AND2X1 U15701 ( .IN1(n9719), .IN2(test_so31), .Q(n15532) );
  OR2X1 U15702 ( .IN1(n15536), .IN2(n15537), .Q(n15526) );
  AND2X1 U15703 ( .IN1(n15538), .IN2(n13440), .Q(n15537) );
  INVX0 U15704 ( .INP(n15539), .ZN(n15538) );
  AND2X1 U15705 ( .IN1(n11983), .IN2(n15539), .Q(n15536) );
  OR2X1 U15706 ( .IN1(n15540), .IN2(n15541), .Q(n15539) );
  OR2X1 U15707 ( .IN1(n15542), .IN2(n15543), .Q(n15541) );
  AND2X1 U15708 ( .IN1(n9718), .IN2(g6368), .Q(n15543) );
  AND2X1 U15709 ( .IN1(n9717), .IN2(g6518), .Q(n15542) );
  AND2X1 U15710 ( .IN1(n9716), .IN2(test_so31), .Q(n15540) );
  OR2X1 U15711 ( .IN1(n15544), .IN2(n15545), .Q(n15524) );
  OR2X1 U15712 ( .IN1(n15546), .IN2(n15547), .Q(n15545) );
  OR2X1 U15713 ( .IN1(n15548), .IN2(n15549), .Q(n15547) );
  AND2X1 U15714 ( .IN1(n15550), .IN2(g793), .Q(n15549) );
  INVX0 U15715 ( .INP(n15551), .ZN(n15550) );
  AND2X1 U15716 ( .IN1(n4321), .IN2(n15551), .Q(n15548) );
  OR2X1 U15717 ( .IN1(n15552), .IN2(n15553), .Q(n15551) );
  OR2X1 U15718 ( .IN1(n15554), .IN2(n15555), .Q(n15553) );
  AND2X1 U15719 ( .IN1(n10092), .IN2(g6368), .Q(n15555) );
  AND2X1 U15720 ( .IN1(n10091), .IN2(g6518), .Q(n15554) );
  AND2X1 U15721 ( .IN1(n9727), .IN2(test_so31), .Q(n15552) );
  OR2X1 U15722 ( .IN1(n15556), .IN2(n15557), .Q(n15546) );
  AND2X1 U15723 ( .IN1(n15558), .IN2(g785), .Q(n15557) );
  INVX0 U15724 ( .INP(n15559), .ZN(n15558) );
  AND2X1 U15725 ( .IN1(n4379), .IN2(n15559), .Q(n15556) );
  OR2X1 U15726 ( .IN1(n15560), .IN2(n15561), .Q(n15559) );
  OR2X1 U15727 ( .IN1(n15562), .IN2(n15563), .Q(n15561) );
  AND2X1 U15728 ( .IN1(n10096), .IN2(g6368), .Q(n15563) );
  AND2X1 U15729 ( .IN1(n10095), .IN2(g6518), .Q(n15562) );
  AND2X1 U15730 ( .IN1(n9729), .IN2(test_so31), .Q(n15560) );
  OR2X1 U15731 ( .IN1(n15564), .IN2(n15565), .Q(n15544) );
  INVX0 U15732 ( .INP(n15566), .ZN(n15565) );
  OR2X1 U15733 ( .IN1(n15567), .IN2(n4375), .Q(n15566) );
  AND2X1 U15734 ( .IN1(n4375), .IN2(n15567), .Q(n15564) );
  OR2X1 U15735 ( .IN1(n15568), .IN2(n15569), .Q(n15567) );
  OR2X1 U15736 ( .IN1(n15570), .IN2(n15571), .Q(n15569) );
  AND2X1 U15737 ( .IN1(n10094), .IN2(g6368), .Q(n15571) );
  AND2X1 U15738 ( .IN1(n10093), .IN2(g6518), .Q(n15570) );
  AND2X1 U15739 ( .IN1(n9728), .IN2(test_so31), .Q(n15568) );
  OR2X1 U15740 ( .IN1(n15572), .IN2(n15573), .Q(n15522) );
  OR2X1 U15741 ( .IN1(n15574), .IN2(n15575), .Q(n15573) );
  OR2X1 U15742 ( .IN1(n15576), .IN2(n15577), .Q(n15575) );
  OR2X1 U15743 ( .IN1(n15578), .IN2(n15579), .Q(n15577) );
  AND2X1 U15744 ( .IN1(n15580), .IN2(g809), .Q(n15579) );
  INVX0 U15745 ( .INP(n15581), .ZN(n15580) );
  AND2X1 U15746 ( .IN1(n4567), .IN2(n15581), .Q(n15578) );
  OR2X1 U15747 ( .IN1(n15582), .IN2(n15583), .Q(n15581) );
  OR2X1 U15748 ( .IN1(n15584), .IN2(n15585), .Q(n15583) );
  AND2X1 U15749 ( .IN1(n10085), .IN2(g6368), .Q(n15585) );
  AND2X1 U15750 ( .IN1(n10084), .IN2(g6518), .Q(n15584) );
  AND2X1 U15751 ( .IN1(n9723), .IN2(test_so31), .Q(n15582) );
  OR2X1 U15752 ( .IN1(n15586), .IN2(n15587), .Q(n15576) );
  AND2X1 U15753 ( .IN1(n15588), .IN2(g805), .Q(n15587) );
  INVX0 U15754 ( .INP(n15589), .ZN(n15588) );
  AND2X1 U15755 ( .IN1(n4559), .IN2(n15589), .Q(n15586) );
  OR2X1 U15756 ( .IN1(n15590), .IN2(n15591), .Q(n15589) );
  OR2X1 U15757 ( .IN1(n15592), .IN2(n15593), .Q(n15591) );
  AND2X1 U15758 ( .IN1(g6368), .IN2(n10212), .Q(n15593) );
  AND2X1 U15759 ( .IN1(n10086), .IN2(g6518), .Q(n15592) );
  AND2X1 U15760 ( .IN1(n9724), .IN2(test_so31), .Q(n15590) );
  OR2X1 U15761 ( .IN1(n15594), .IN2(n15595), .Q(n15574) );
  INVX0 U15762 ( .INP(n15596), .ZN(n15595) );
  OR2X1 U15763 ( .IN1(n15597), .IN2(n4391), .Q(n15596) );
  AND2X1 U15764 ( .IN1(n4391), .IN2(n15597), .Q(n15594) );
  OR2X1 U15765 ( .IN1(n15598), .IN2(n15599), .Q(n15597) );
  OR2X1 U15766 ( .IN1(n15600), .IN2(n15601), .Q(n15599) );
  AND2X1 U15767 ( .IN1(n10090), .IN2(g6368), .Q(n15601) );
  AND2X1 U15768 ( .IN1(n10089), .IN2(g6518), .Q(n15600) );
  AND2X1 U15769 ( .IN1(n9726), .IN2(test_so31), .Q(n15598) );
  OR2X1 U15770 ( .IN1(n15602), .IN2(n15603), .Q(n15572) );
  OR2X1 U15771 ( .IN1(n11579), .IN2(n15604), .Q(n15603) );
  OR2X1 U15772 ( .IN1(n15605), .IN2(n15606), .Q(n15604) );
  AND2X1 U15773 ( .IN1(n15607), .IN2(g813), .Q(n15606) );
  INVX0 U15774 ( .INP(n15608), .ZN(n15607) );
  AND2X1 U15775 ( .IN1(n4289), .IN2(n15608), .Q(n15605) );
  OR2X1 U15776 ( .IN1(n15609), .IN2(n15610), .Q(n15608) );
  OR2X1 U15777 ( .IN1(n15611), .IN2(n15612), .Q(n15610) );
  AND2X1 U15778 ( .IN1(n10083), .IN2(g6368), .Q(n15612) );
  AND2X1 U15779 ( .IN1(n10082), .IN2(g6518), .Q(n15611) );
  AND2X1 U15780 ( .IN1(n9722), .IN2(test_so31), .Q(n15609) );
  INVX0 U15781 ( .INP(n3102), .ZN(n11579) );
  OR2X1 U15782 ( .IN1(n15613), .IN2(n15614), .Q(n15602) );
  AND2X1 U15783 ( .IN1(n15615), .IN2(g801), .Q(n15614) );
  INVX0 U15784 ( .INP(n15616), .ZN(n15615) );
  AND2X1 U15785 ( .IN1(n4327), .IN2(n15616), .Q(n15613) );
  OR2X1 U15786 ( .IN1(n15617), .IN2(n15618), .Q(n15616) );
  OR2X1 U15787 ( .IN1(n15619), .IN2(n15620), .Q(n15618) );
  AND2X1 U15788 ( .IN1(n10088), .IN2(g6368), .Q(n15620) );
  AND2X1 U15789 ( .IN1(n10087), .IN2(g6518), .Q(n15619) );
  AND2X1 U15790 ( .IN1(n9725), .IN2(test_so31), .Q(n15617) );
  OR2X1 U15791 ( .IN1(n15621), .IN2(n15622), .Q(n12950) );
  OR2X1 U15792 ( .IN1(n15623), .IN2(n15624), .Q(n15622) );
  AND2X1 U15793 ( .IN1(n9849), .IN2(g6712), .Q(n15624) );
  AND2X1 U15794 ( .IN1(n9862), .IN2(g5472), .Q(n15623) );
  AND2X1 U15795 ( .IN1(n9861), .IN2(g1088), .Q(n15621) );
  AND2X1 U15796 ( .IN1(n15625), .IN2(n15626), .Q(g26660) );
  OR2X1 U15797 ( .IN1(n15627), .IN2(g672), .Q(n15626) );
  AND2X1 U15798 ( .IN1(n15628), .IN2(g660), .Q(n15627) );
  AND2X1 U15799 ( .IN1(n13809), .IN2(n14478), .Q(n15625) );
  OR2X1 U15800 ( .IN1(n15629), .IN2(n15630), .Q(n14478) );
  OR2X1 U15801 ( .IN1(n4413), .IN2(n4403), .Q(n15630) );
  OR2X1 U15802 ( .IN1(n15631), .IN2(n15632), .Q(g26659) );
  AND2X1 U15803 ( .IN1(n15515), .IN2(n13502), .Q(n15632) );
  AND2X1 U15804 ( .IN1(n15633), .IN2(g404), .Q(n15631) );
  OR2X1 U15805 ( .IN1(n4499), .IN2(n15517), .Q(n15633) );
  OR2X1 U15806 ( .IN1(n15634), .IN2(n15635), .Q(g26655) );
  AND2X1 U15807 ( .IN1(n15515), .IN2(n13506), .Q(n15635) );
  AND2X1 U15808 ( .IN1(g309), .IN2(n15517), .Q(n15515) );
  AND2X1 U15809 ( .IN1(n15636), .IN2(g403), .Q(n15634) );
  OR2X1 U15810 ( .IN1(n4520), .IN2(n15517), .Q(n15636) );
  OR2X1 U15811 ( .IN1(n12961), .IN2(n15637), .Q(n15517) );
  OR2X1 U15812 ( .IN1(n4388), .IN2(n12813), .Q(n15637) );
  OR2X1 U15813 ( .IN1(n15638), .IN2(n15639), .Q(n12813) );
  OR2X1 U15814 ( .IN1(n15640), .IN2(n15641), .Q(n15639) );
  OR2X1 U15815 ( .IN1(n15642), .IN2(n15643), .Q(n15641) );
  OR2X1 U15816 ( .IN1(n15644), .IN2(n15645), .Q(n15643) );
  AND2X1 U15817 ( .IN1(n15646), .IN2(n12218), .Q(n15645) );
  INVX0 U15818 ( .INP(n15647), .ZN(n15646) );
  AND2X1 U15819 ( .IN1(n13567), .IN2(n15647), .Q(n15644) );
  OR2X1 U15820 ( .IN1(n15648), .IN2(n15649), .Q(n15647) );
  OR2X1 U15821 ( .IN1(n15650), .IN2(n15651), .Q(n15649) );
  AND2X1 U15822 ( .IN1(n9692), .IN2(g165), .Q(n15651) );
  AND2X1 U15823 ( .IN1(n9694), .IN2(g6231), .Q(n15650) );
  AND2X1 U15824 ( .IN1(n9693), .IN2(g6313), .Q(n15648) );
  OR2X1 U15825 ( .IN1(n15652), .IN2(n15653), .Q(n15642) );
  AND2X1 U15826 ( .IN1(n15654), .IN2(g105), .Q(n15653) );
  INVX0 U15827 ( .INP(n15655), .ZN(n15654) );
  AND2X1 U15828 ( .IN1(n4322), .IN2(n15655), .Q(n15652) );
  OR2X1 U15829 ( .IN1(n15656), .IN2(n15657), .Q(n15655) );
  OR2X1 U15830 ( .IN1(n15658), .IN2(n15659), .Q(n15657) );
  AND2X1 U15831 ( .IN1(n10108), .IN2(g6231), .Q(n15659) );
  AND2X1 U15832 ( .IN1(n10107), .IN2(g6313), .Q(n15658) );
  AND2X1 U15833 ( .IN1(n9736), .IN2(g165), .Q(n15656) );
  OR2X1 U15834 ( .IN1(n15660), .IN2(n15661), .Q(n15640) );
  OR2X1 U15835 ( .IN1(n15662), .IN2(n15663), .Q(n15661) );
  OR2X1 U15836 ( .IN1(n15664), .IN2(n15665), .Q(n15663) );
  AND2X1 U15837 ( .IN1(n15666), .IN2(g97), .Q(n15665) );
  INVX0 U15838 ( .INP(n15667), .ZN(n15666) );
  AND2X1 U15839 ( .IN1(n4380), .IN2(n15667), .Q(n15664) );
  OR2X1 U15840 ( .IN1(n15668), .IN2(n15669), .Q(n15667) );
  OR2X1 U15841 ( .IN1(n15670), .IN2(n15671), .Q(n15669) );
  AND2X1 U15842 ( .IN1(n10112), .IN2(g6231), .Q(n15671) );
  AND2X1 U15843 ( .IN1(n10111), .IN2(g6313), .Q(n15670) );
  AND2X1 U15844 ( .IN1(n9738), .IN2(g165), .Q(n15668) );
  OR2X1 U15845 ( .IN1(n15672), .IN2(n15673), .Q(n15662) );
  INVX0 U15846 ( .INP(n15674), .ZN(n15673) );
  OR2X1 U15847 ( .IN1(n15675), .IN2(n4376), .Q(n15674) );
  AND2X1 U15848 ( .IN1(n4376), .IN2(n15675), .Q(n15672) );
  OR2X1 U15849 ( .IN1(n15676), .IN2(n15677), .Q(n15675) );
  OR2X1 U15850 ( .IN1(n15678), .IN2(n15679), .Q(n15677) );
  AND2X1 U15851 ( .IN1(n10110), .IN2(g6231), .Q(n15679) );
  AND2X1 U15852 ( .IN1(n10109), .IN2(g6313), .Q(n15678) );
  AND2X1 U15853 ( .IN1(n9737), .IN2(g165), .Q(n15676) );
  OR2X1 U15854 ( .IN1(n15680), .IN2(n15681), .Q(n15660) );
  AND2X1 U15855 ( .IN1(n15682), .IN2(n13590), .Q(n15681) );
  INVX0 U15856 ( .INP(n15683), .ZN(n15682) );
  AND2X1 U15857 ( .IN1(n12036), .IN2(n15683), .Q(n15680) );
  OR2X1 U15858 ( .IN1(n15684), .IN2(n15685), .Q(n15683) );
  OR2X1 U15859 ( .IN1(n15686), .IN2(n15687), .Q(n15685) );
  AND2X1 U15860 ( .IN1(n9730), .IN2(g165), .Q(n15687) );
  AND2X1 U15861 ( .IN1(g6231), .IN2(n10213), .Q(n15686) );
  AND2X1 U15862 ( .IN1(n9731), .IN2(g6313), .Q(n15684) );
  OR2X1 U15863 ( .IN1(n15688), .IN2(n15689), .Q(n15638) );
  OR2X1 U15864 ( .IN1(n15690), .IN2(n15691), .Q(n15689) );
  OR2X1 U15865 ( .IN1(n15692), .IN2(n15693), .Q(n15691) );
  OR2X1 U15866 ( .IN1(n15694), .IN2(n15695), .Q(n15693) );
  AND2X1 U15867 ( .IN1(n15696), .IN2(g121), .Q(n15695) );
  INVX0 U15868 ( .INP(n15697), .ZN(n15696) );
  AND2X1 U15869 ( .IN1(n4569), .IN2(n15697), .Q(n15694) );
  OR2X1 U15870 ( .IN1(n15698), .IN2(n15699), .Q(n15697) );
  OR2X1 U15871 ( .IN1(n15700), .IN2(n15701), .Q(n15699) );
  AND2X1 U15872 ( .IN1(n10100), .IN2(g6231), .Q(n15701) );
  AND2X1 U15873 ( .IN1(n10099), .IN2(g6313), .Q(n15700) );
  AND2X1 U15874 ( .IN1(n9733), .IN2(g165), .Q(n15698) );
  OR2X1 U15875 ( .IN1(n15702), .IN2(n15703), .Q(n15692) );
  AND2X1 U15876 ( .IN1(n15704), .IN2(g117), .Q(n15703) );
  INVX0 U15877 ( .INP(n15705), .ZN(n15704) );
  AND2X1 U15878 ( .IN1(n4561), .IN2(n15705), .Q(n15702) );
  OR2X1 U15879 ( .IN1(n15706), .IN2(n15707), .Q(n15705) );
  OR2X1 U15880 ( .IN1(n15708), .IN2(n15709), .Q(n15707) );
  AND2X1 U15881 ( .IN1(n10102), .IN2(g6231), .Q(n15709) );
  AND2X1 U15882 ( .IN1(n10101), .IN2(g6313), .Q(n15708) );
  AND2X1 U15883 ( .IN1(n9734), .IN2(g165), .Q(n15706) );
  OR2X1 U15884 ( .IN1(n15710), .IN2(n15711), .Q(n15690) );
  AND2X1 U15885 ( .IN1(n15712), .IN2(g109), .Q(n15711) );
  INVX0 U15886 ( .INP(n15713), .ZN(n15712) );
  AND2X1 U15887 ( .IN1(n4392), .IN2(n15713), .Q(n15710) );
  OR2X1 U15888 ( .IN1(n15714), .IN2(n15715), .Q(n15713) );
  OR2X1 U15889 ( .IN1(n15716), .IN2(n15717), .Q(n15715) );
  AND2X1 U15890 ( .IN1(n10106), .IN2(g6231), .Q(n15717) );
  AND2X1 U15891 ( .IN1(n10105), .IN2(g6313), .Q(n15716) );
  AND2X1 U15892 ( .IN1(g165), .IN2(n10214), .Q(n15714) );
  OR2X1 U15893 ( .IN1(n15718), .IN2(n15719), .Q(n15688) );
  OR2X1 U15894 ( .IN1(n11838), .IN2(n15720), .Q(n15719) );
  OR2X1 U15895 ( .IN1(n15721), .IN2(n15722), .Q(n15720) );
  AND2X1 U15896 ( .IN1(n15723), .IN2(g125), .Q(n15722) );
  INVX0 U15897 ( .INP(n15724), .ZN(n15723) );
  AND2X1 U15898 ( .IN1(n4290), .IN2(n15724), .Q(n15721) );
  OR2X1 U15899 ( .IN1(n15725), .IN2(n15726), .Q(n15724) );
  OR2X1 U15900 ( .IN1(n15727), .IN2(n15728), .Q(n15726) );
  AND2X1 U15901 ( .IN1(n10098), .IN2(g6231), .Q(n15728) );
  AND2X1 U15902 ( .IN1(n10097), .IN2(g6313), .Q(n15727) );
  AND2X1 U15903 ( .IN1(n9732), .IN2(g165), .Q(n15725) );
  INVX0 U15904 ( .INP(n3130), .ZN(n11838) );
  OR2X1 U15905 ( .IN1(n15729), .IN2(n15730), .Q(n15718) );
  AND2X1 U15906 ( .IN1(n15731), .IN2(g113), .Q(n15730) );
  INVX0 U15907 ( .INP(n15732), .ZN(n15731) );
  AND2X1 U15908 ( .IN1(n4328), .IN2(n15732), .Q(n15729) );
  OR2X1 U15909 ( .IN1(n15733), .IN2(n15734), .Q(n15732) );
  OR2X1 U15910 ( .IN1(n15735), .IN2(n15736), .Q(n15734) );
  AND2X1 U15911 ( .IN1(n10104), .IN2(g6231), .Q(n15736) );
  AND2X1 U15912 ( .IN1(n10103), .IN2(g6313), .Q(n15735) );
  AND2X1 U15913 ( .IN1(n9735), .IN2(g165), .Q(n15733) );
  OR2X1 U15914 ( .IN1(n15737), .IN2(n15738), .Q(n12961) );
  OR2X1 U15915 ( .IN1(n15739), .IN2(n15740), .Q(n15738) );
  AND2X1 U15916 ( .IN1(n9867), .IN2(n13375), .Q(n15740) );
  AND2X1 U15917 ( .IN1(n9868), .IN2(n13502), .Q(n15739) );
  AND2X1 U15918 ( .IN1(n9869), .IN2(n13506), .Q(n15737) );
  OR2X1 U15919 ( .IN1(n15741), .IN2(n15742), .Q(g26616) );
  AND2X1 U15920 ( .IN1(n15743), .IN2(g2624), .Q(n15742) );
  AND2X1 U15921 ( .IN1(n4299), .IN2(g2571), .Q(n15741) );
  OR2X1 U15922 ( .IN1(n15744), .IN2(n15745), .Q(g26596) );
  AND2X1 U15923 ( .IN1(n15743), .IN2(g7390), .Q(n15745) );
  AND2X1 U15924 ( .IN1(n4370), .IN2(g2568), .Q(n15744) );
  OR2X1 U15925 ( .IN1(n15746), .IN2(n15747), .Q(g26592) );
  AND2X1 U15926 ( .IN1(n15748), .IN2(g1930), .Q(n15747) );
  AND2X1 U15927 ( .IN1(n4366), .IN2(g1877), .Q(n15746) );
  OR2X1 U15928 ( .IN1(n15749), .IN2(n15750), .Q(g26575) );
  AND2X1 U15929 ( .IN1(n15743), .IN2(n12862), .Q(n15750) );
  AND2X1 U15930 ( .IN1(n15751), .IN2(n15752), .Q(n15743) );
  AND2X1 U15931 ( .IN1(g2584), .IN2(n11222), .Q(n15752) );
  AND2X1 U15932 ( .IN1(n4314), .IN2(g2565), .Q(n15749) );
  OR2X1 U15933 ( .IN1(n15753), .IN2(n15754), .Q(g26573) );
  AND2X1 U15934 ( .IN1(n15748), .IN2(g7194), .Q(n15754) );
  AND2X1 U15935 ( .IN1(n4315), .IN2(g1874), .Q(n15753) );
  OR2X1 U15936 ( .IN1(n15755), .IN2(n15756), .Q(g26569) );
  AND2X1 U15937 ( .IN1(n15757), .IN2(g1236), .Q(n15756) );
  AND2X1 U15938 ( .IN1(n4300), .IN2(g1183), .Q(n15755) );
  OR2X1 U15939 ( .IN1(n15758), .IN2(n15759), .Q(g26559) );
  AND2X1 U15940 ( .IN1(test_so68), .IN2(n4296), .Q(n15759) );
  AND2X1 U15941 ( .IN1(n15748), .IN2(n13973), .Q(n15758) );
  AND2X1 U15942 ( .IN1(n15760), .IN2(n15761), .Q(n15748) );
  AND2X1 U15943 ( .IN1(g1890), .IN2(n11383), .Q(n15761) );
  OR2X1 U15944 ( .IN1(n15762), .IN2(n15763), .Q(g26557) );
  AND2X1 U15945 ( .IN1(n15757), .IN2(g6944), .Q(n15763) );
  AND2X1 U15946 ( .IN1(n4316), .IN2(g1180), .Q(n15762) );
  OR2X1 U15947 ( .IN1(n15764), .IN2(n15765), .Q(g26553) );
  AND2X1 U15948 ( .IN1(n15766), .IN2(g550), .Q(n15765) );
  AND2X1 U15949 ( .IN1(n4313), .IN2(g496), .Q(n15764) );
  OR2X1 U15950 ( .IN1(n15767), .IN2(n15768), .Q(g26547) );
  AND2X1 U15951 ( .IN1(test_so47), .IN2(n4371), .Q(n15768) );
  AND2X1 U15952 ( .IN1(n15757), .IN2(n13842), .Q(n15767) );
  AND2X1 U15953 ( .IN1(n15769), .IN2(n15770), .Q(n15757) );
  AND2X1 U15954 ( .IN1(g1196), .IN2(n11546), .Q(n15770) );
  OR2X1 U15955 ( .IN1(n15771), .IN2(n15772), .Q(g26545) );
  AND2X1 U15956 ( .IN1(n15766), .IN2(g6642), .Q(n15772) );
  AND2X1 U15957 ( .IN1(n4372), .IN2(g493), .Q(n15771) );
  OR2X1 U15958 ( .IN1(n15773), .IN2(n15774), .Q(g26541) );
  AND2X1 U15959 ( .IN1(n15766), .IN2(n11054), .Q(n15774) );
  AND2X1 U15960 ( .IN1(n15775), .IN2(n15776), .Q(n15766) );
  AND2X1 U15961 ( .IN1(n11058), .IN2(test_so22), .Q(n15776) );
  AND2X1 U15962 ( .IN1(n4298), .IN2(g490), .Q(n15773) );
  AND2X1 U15963 ( .IN1(n15777), .IN2(n12966), .Q(g26532) );
  OR2X1 U15964 ( .IN1(n15778), .IN2(n15779), .Q(n15777) );
  AND2X1 U15965 ( .IN1(n4526), .IN2(g2151), .Q(n15779) );
  AND2X1 U15966 ( .IN1(n9878), .IN2(n15780), .Q(n15778) );
  INVX0 U15967 ( .INP(n4526), .ZN(n15780) );
  AND2X1 U15968 ( .IN1(n15781), .IN2(n12971), .Q(g26531) );
  OR2X1 U15969 ( .IN1(n15782), .IN2(n15783), .Q(n15781) );
  AND2X1 U15970 ( .IN1(n4527), .IN2(g1457), .Q(n15783) );
  AND2X1 U15971 ( .IN1(n9882), .IN2(n15784), .Q(n15782) );
  INVX0 U15972 ( .INP(n4527), .ZN(n15784) );
  AND2X1 U15973 ( .IN1(n15785), .IN2(n12976), .Q(g26530) );
  AND2X1 U15974 ( .IN1(n15786), .IN2(n15787), .Q(n15785) );
  INVX0 U15975 ( .INP(n15788), .ZN(n15787) );
  AND2X1 U15976 ( .IN1(n879), .IN2(n9886), .Q(n15788) );
  OR2X1 U15977 ( .IN1(n9886), .IN2(n879), .Q(n15786) );
  AND2X1 U15978 ( .IN1(n15789), .IN2(n12981), .Q(g26529) );
  OR2X1 U15979 ( .IN1(n15790), .IN2(n15791), .Q(n15789) );
  AND2X1 U15980 ( .IN1(n4528), .IN2(g83), .Q(n15791) );
  AND2X1 U15981 ( .IN1(n9890), .IN2(n15792), .Q(n15790) );
  INVX0 U15982 ( .INP(n4528), .ZN(n15792) );
  OR2X1 U15983 ( .IN1(n15793), .IN2(n15794), .Q(g26149) );
  OR2X1 U15984 ( .IN1(n15795), .IN2(n15796), .Q(n15794) );
  OR2X1 U15985 ( .IN1(n15797), .IN2(n14497), .Q(n15796) );
  AND2X1 U15986 ( .IN1(n14501), .IN2(n8086), .Q(n15797) );
  OR2X1 U15987 ( .IN1(n15798), .IN2(n15799), .Q(n15795) );
  OR2X1 U15988 ( .IN1(n15800), .IN2(n15801), .Q(n15799) );
  AND2X1 U15989 ( .IN1(n15802), .IN2(g3170), .Q(n15801) );
  AND2X1 U15990 ( .IN1(n15803), .IN2(g3173), .Q(n15800) );
  AND2X1 U15991 ( .IN1(n15804), .IN2(n8080), .Q(n15798) );
  OR2X1 U15992 ( .IN1(n15805), .IN2(n15806), .Q(n15793) );
  OR2X1 U15993 ( .IN1(n15807), .IN2(n15808), .Q(n15806) );
  OR2X1 U15994 ( .IN1(n15809), .IN2(n15810), .Q(n15808) );
  AND2X1 U15995 ( .IN1(n15811), .IN2(g3176), .Q(n15810) );
  AND2X1 U15996 ( .IN1(n14502), .IN2(n8076), .Q(n15809) );
  AND2X1 U15997 ( .IN1(n15812), .IN2(g3161), .Q(n15807) );
  OR2X1 U15998 ( .IN1(n15813), .IN2(n15814), .Q(n15805) );
  OR2X1 U15999 ( .IN1(n15815), .IN2(n15816), .Q(n15814) );
  AND2X1 U16000 ( .IN1(n3939), .IN2(n15817), .Q(n15816) );
  OR2X1 U16001 ( .IN1(n15818), .IN2(n15819), .Q(n15817) );
  OR2X1 U16002 ( .IN1(n15820), .IN2(n15821), .Q(n15819) );
  AND2X1 U16003 ( .IN1(n15822), .IN2(g3155), .Q(n15821) );
  AND2X1 U16004 ( .IN1(test_so8), .IN2(n14522), .Q(n15820) );
  AND2X1 U16005 ( .IN1(n3940), .IN2(g3185), .Q(n15818) );
  AND2X1 U16006 ( .IN1(n15823), .IN2(g3167), .Q(n15815) );
  AND2X1 U16007 ( .IN1(n3936), .IN2(n15824), .Q(n15813) );
  OR2X1 U16008 ( .IN1(n15825), .IN2(n15826), .Q(n15824) );
  OR2X1 U16009 ( .IN1(n15827), .IN2(n15828), .Q(n15826) );
  AND2X1 U16010 ( .IN1(n14508), .IN2(g3182), .Q(n15828) );
  AND2X1 U16011 ( .IN1(n15829), .IN2(g3158), .Q(n15827) );
  OR2X1 U16012 ( .IN1(n15830), .IN2(n15831), .Q(n15825) );
  AND2X1 U16013 ( .IN1(n15832), .IN2(g3164), .Q(n15831) );
  AND2X1 U16014 ( .IN1(n15833), .IN2(g3088), .Q(n15830) );
  OR2X1 U16015 ( .IN1(n15834), .IN2(n15835), .Q(g26135) );
  OR2X1 U16016 ( .IN1(n15836), .IN2(n15837), .Q(n15835) );
  OR2X1 U16017 ( .IN1(n14497), .IN2(n15838), .Q(n15837) );
  OR2X1 U16018 ( .IN1(n15839), .IN2(n15840), .Q(n15838) );
  AND2X1 U16019 ( .IN1(n9801), .IN2(n14501), .Q(n15840) );
  AND2X1 U16020 ( .IN1(n15804), .IN2(n8081), .Q(n15839) );
  OR2X1 U16021 ( .IN1(n15841), .IN2(n15842), .Q(n15836) );
  OR2X1 U16022 ( .IN1(n15843), .IN2(n15844), .Q(n15842) );
  AND2X1 U16023 ( .IN1(n15803), .IN2(g3103), .Q(n15844) );
  AND2X1 U16024 ( .IN1(n15812), .IN2(g3099), .Q(n15843) );
  AND2X1 U16025 ( .IN1(n15802), .IN2(g3102), .Q(n15841) );
  OR2X1 U16026 ( .IN1(n15845), .IN2(n15846), .Q(n15834) );
  OR2X1 U16027 ( .IN1(n15847), .IN2(n15848), .Q(n15846) );
  OR2X1 U16028 ( .IN1(n15849), .IN2(n15850), .Q(n15848) );
  AND2X1 U16029 ( .IN1(n14502), .IN2(n8077), .Q(n15850) );
  AND2X1 U16030 ( .IN1(n3936), .IN2(n15851), .Q(n15849) );
  OR2X1 U16031 ( .IN1(n15852), .IN2(n15853), .Q(n15851) );
  OR2X1 U16032 ( .IN1(n15854), .IN2(n15855), .Q(n15853) );
  AND2X1 U16033 ( .IN1(n14508), .IN2(g3106), .Q(n15855) );
  AND2X1 U16034 ( .IN1(n15829), .IN2(g3098), .Q(n15854) );
  OR2X1 U16035 ( .IN1(n15856), .IN2(n15857), .Q(n15852) );
  AND2X1 U16036 ( .IN1(n15832), .IN2(g3100), .Q(n15857) );
  AND2X1 U16037 ( .IN1(n15833), .IN2(g3108), .Q(n15856) );
  AND2X1 U16038 ( .IN1(n15811), .IN2(g3104), .Q(n15847) );
  OR2X1 U16039 ( .IN1(n15858), .IN2(n15859), .Q(n15845) );
  OR2X1 U16040 ( .IN1(n15860), .IN2(n15861), .Q(n15859) );
  AND2X1 U16041 ( .IN1(n3939), .IN2(n15862), .Q(n15861) );
  OR2X1 U16042 ( .IN1(n15863), .IN2(n15864), .Q(n15862) );
  OR2X1 U16043 ( .IN1(n15865), .IN2(n15866), .Q(n15864) );
  AND2X1 U16044 ( .IN1(n15822), .IN2(g3097), .Q(n15866) );
  AND2X1 U16045 ( .IN1(n14522), .IN2(g3105), .Q(n15865) );
  AND2X1 U16046 ( .IN1(n3940), .IN2(g3107), .Q(n15863) );
  AND2X1 U16047 ( .IN1(test_so10), .IN2(n14507), .Q(n15860) );
  OR2X1 U16048 ( .IN1(n15867), .IN2(n15868), .Q(n15858) );
  AND2X1 U16049 ( .IN1(n14512), .IN2(n14519), .Q(n15868) );
  AND2X1 U16050 ( .IN1(test_so7), .IN2(n15823), .Q(n15867) );
  OR2X1 U16051 ( .IN1(n15869), .IN2(n15870), .Q(g26104) );
  OR2X1 U16052 ( .IN1(n15871), .IN2(n15872), .Q(n15870) );
  OR2X1 U16053 ( .IN1(n14497), .IN2(n15873), .Q(n15872) );
  OR2X1 U16054 ( .IN1(n15874), .IN2(n15875), .Q(n15873) );
  AND2X1 U16055 ( .IN1(n14501), .IN2(n8087), .Q(n15875) );
  AND2X1 U16056 ( .IN1(n15804), .IN2(n8082), .Q(n15874) );
  OR2X1 U16057 ( .IN1(n15876), .IN2(n15877), .Q(n15871) );
  OR2X1 U16058 ( .IN1(n15878), .IN2(n15879), .Q(n15877) );
  AND2X1 U16059 ( .IN1(n15803), .IN2(g3091), .Q(n15879) );
  AND2X1 U16060 ( .IN1(n3933), .IN2(n15880), .Q(n15803) );
  AND2X1 U16061 ( .IN1(n4406), .IN2(n14521), .Q(n15880) );
  AND2X1 U16062 ( .IN1(n15812), .IN2(g3084), .Q(n15878) );
  AND2X1 U16063 ( .IN1(n3933), .IN2(n15881), .Q(n15812) );
  AND2X1 U16064 ( .IN1(n4406), .IN2(n3939), .Q(n15881) );
  AND2X1 U16065 ( .IN1(g3207), .IN2(n4405), .Q(n3933) );
  AND2X1 U16066 ( .IN1(n15802), .IN2(g3087), .Q(n15876) );
  AND2X1 U16067 ( .IN1(n15829), .IN2(n14511), .Q(n15802) );
  OR2X1 U16068 ( .IN1(n15882), .IN2(n15883), .Q(n15869) );
  OR2X1 U16069 ( .IN1(n15884), .IN2(n15885), .Q(n15883) );
  OR2X1 U16070 ( .IN1(n15886), .IN2(n15887), .Q(n15885) );
  AND2X1 U16071 ( .IN1(n14502), .IN2(n8078), .Q(n15887) );
  AND2X1 U16072 ( .IN1(n14522), .IN2(n15888), .Q(n14502) );
  AND2X1 U16073 ( .IN1(n3936), .IN2(n15889), .Q(n15886) );
  OR2X1 U16074 ( .IN1(n15890), .IN2(n15891), .Q(n15889) );
  OR2X1 U16075 ( .IN1(n15892), .IN2(n15893), .Q(n15891) );
  AND2X1 U16076 ( .IN1(n14508), .IN2(g3094), .Q(n15893) );
  AND2X1 U16077 ( .IN1(n15829), .IN2(g3211), .Q(n15892) );
  OR2X1 U16078 ( .IN1(n15894), .IN2(n15895), .Q(n15890) );
  AND2X1 U16079 ( .IN1(n15832), .IN2(g3085), .Q(n15895) );
  AND2X1 U16080 ( .IN1(n15833), .IN2(g3096), .Q(n15894) );
  AND2X1 U16081 ( .IN1(g3201), .IN2(g3207), .Q(n15833) );
  AND2X1 U16082 ( .IN1(n15811), .IN2(g3092), .Q(n15884) );
  AND2X1 U16083 ( .IN1(n14511), .IN2(n15832), .Q(n15811) );
  AND2X1 U16084 ( .IN1(g3207), .IN2(n4406), .Q(n15832) );
  AND2X1 U16085 ( .IN1(g3188), .IN2(n14521), .Q(n14511) );
  OR2X1 U16086 ( .IN1(n15896), .IN2(n15897), .Q(n15882) );
  OR2X1 U16087 ( .IN1(n15898), .IN2(n15899), .Q(n15897) );
  AND2X1 U16088 ( .IN1(n3939), .IN2(n15900), .Q(n15899) );
  OR2X1 U16089 ( .IN1(n15901), .IN2(n15902), .Q(n15900) );
  OR2X1 U16090 ( .IN1(n15903), .IN2(n15904), .Q(n15902) );
  AND2X1 U16091 ( .IN1(test_so6), .IN2(n15822), .Q(n15904) );
  AND2X1 U16092 ( .IN1(n14522), .IN2(g3093), .Q(n15903) );
  AND2X1 U16093 ( .IN1(n4405), .IN2(n14508), .Q(n14522) );
  AND2X1 U16094 ( .IN1(g3201), .IN2(n4329), .Q(n14508) );
  AND2X1 U16095 ( .IN1(n3940), .IN2(g3095), .Q(n15901) );
  AND2X1 U16096 ( .IN1(n14507), .IN2(g3142), .Q(n15898) );
  AND2X1 U16097 ( .IN1(n15888), .IN2(n3940), .Q(n14507) );
  OR2X1 U16098 ( .IN1(n15905), .IN2(n15906), .Q(n15896) );
  AND2X1 U16099 ( .IN1(n14512), .IN2(n14520), .Q(n15906) );
  AND2X1 U16100 ( .IN1(n15822), .IN2(n3705), .Q(n14512) );
  AND2X1 U16101 ( .IN1(n15823), .IN2(g3086), .Q(n15905) );
  AND2X1 U16102 ( .IN1(n15822), .IN2(n14521), .Q(n15823) );
  AND2X1 U16103 ( .IN1(g3204), .IN2(n3938), .Q(n14521) );
  AND2X1 U16104 ( .IN1(g3197), .IN2(n323), .Q(n3938) );
  INVX0 U16105 ( .INP(n15907), .ZN(n323) );
  OR2X1 U16106 ( .IN1(n8088), .IN2(n15908), .Q(n15907) );
  OR2X1 U16107 ( .IN1(n8090), .IN2(n8089), .Q(n15908) );
  AND2X1 U16108 ( .IN1(n15909), .IN2(n15910), .Q(g26048) );
  OR2X1 U16109 ( .IN1(n15911), .IN2(n15912), .Q(n15909) );
  AND2X1 U16110 ( .IN1(n15913), .IN2(n15914), .Q(n15911) );
  OR2X1 U16111 ( .IN1(n15915), .IN2(n7909), .Q(n15914) );
  OR2X1 U16112 ( .IN1(n18262), .IN2(n15916), .Q(n15913) );
  AND2X1 U16113 ( .IN1(n15917), .IN2(n11730), .Q(g26037) );
  AND2X1 U16114 ( .IN1(n15918), .IN2(n15345), .Q(n15917) );
  OR2X1 U16115 ( .IN1(n4291), .IN2(n15919), .Q(n15345) );
  OR2X1 U16116 ( .IN1(n15920), .IN2(g2900), .Q(n15918) );
  INVX0 U16117 ( .INP(n15919), .ZN(n15920) );
  AND2X1 U16118 ( .IN1(n15352), .IN2(n15921), .Q(g26031) );
  OR2X1 U16119 ( .IN1(n15922), .IN2(n15923), .Q(n15921) );
  AND2X1 U16120 ( .IN1(n15924), .IN2(n10197), .Q(n15923) );
  AND2X1 U16121 ( .IN1(test_so98), .IN2(n1808), .Q(n15922) );
  OR2X1 U16122 ( .IN1(n15925), .IN2(n15926), .Q(g26025) );
  AND2X1 U16123 ( .IN1(n15372), .IN2(n13101), .Q(n15926) );
  AND2X1 U16124 ( .IN1(n15374), .IN2(test_so79), .Q(n15372) );
  AND2X1 U16125 ( .IN1(test_so82), .IN2(n15927), .Q(n15925) );
  OR2X1 U16126 ( .IN1(n4509), .IN2(n15374), .Q(n15927) );
  OR2X1 U16127 ( .IN1(n12925), .IN2(n15928), .Q(n15374) );
  OR2X1 U16128 ( .IN1(n12633), .IN2(n10191), .Q(n15928) );
  OR2X1 U16129 ( .IN1(n15929), .IN2(n15930), .Q(n12633) );
  OR2X1 U16130 ( .IN1(n15931), .IN2(n15932), .Q(n15930) );
  OR2X1 U16131 ( .IN1(n15933), .IN2(n15934), .Q(n15932) );
  OR2X1 U16132 ( .IN1(n15935), .IN2(n15936), .Q(n15934) );
  AND2X1 U16133 ( .IN1(n15937), .IN2(n12083), .Q(n15936) );
  INVX0 U16134 ( .INP(n15938), .ZN(n15937) );
  AND2X1 U16135 ( .IN1(n13179), .IN2(n15938), .Q(n15935) );
  OR2X1 U16136 ( .IN1(n15939), .IN2(n15940), .Q(n15938) );
  OR2X1 U16137 ( .IN1(n15941), .IN2(n15942), .Q(n15940) );
  AND2X1 U16138 ( .IN1(n9686), .IN2(g2241), .Q(n15942) );
  AND2X1 U16139 ( .IN1(n9688), .IN2(g6837), .Q(n15941) );
  AND2X1 U16140 ( .IN1(n9687), .IN2(test_so73), .Q(n15939) );
  OR2X1 U16141 ( .IN1(n15943), .IN2(n15944), .Q(n15933) );
  AND2X1 U16142 ( .IN1(n15945), .IN2(g2175), .Q(n15944) );
  INVX0 U16143 ( .INP(n15946), .ZN(n15945) );
  AND2X1 U16144 ( .IN1(n4319), .IN2(n15946), .Q(n15943) );
  OR2X1 U16145 ( .IN1(n15947), .IN2(n15948), .Q(n15946) );
  OR2X1 U16146 ( .IN1(n15949), .IN2(n15950), .Q(n15948) );
  AND2X1 U16147 ( .IN1(n10063), .IN2(g6837), .Q(n15950) );
  AND2X1 U16148 ( .IN1(n10062), .IN2(test_so73), .Q(n15949) );
  AND2X1 U16149 ( .IN1(n9702), .IN2(g2241), .Q(n15947) );
  OR2X1 U16150 ( .IN1(n15951), .IN2(n15952), .Q(n15931) );
  OR2X1 U16151 ( .IN1(n15953), .IN2(n15954), .Q(n15952) );
  OR2X1 U16152 ( .IN1(n15955), .IN2(n15956), .Q(n15954) );
  AND2X1 U16153 ( .IN1(n15957), .IN2(g2165), .Q(n15956) );
  INVX0 U16154 ( .INP(n15958), .ZN(n15957) );
  AND2X1 U16155 ( .IN1(n4377), .IN2(n15958), .Q(n15955) );
  OR2X1 U16156 ( .IN1(n15959), .IN2(n15960), .Q(n15958) );
  OR2X1 U16157 ( .IN1(n15961), .IN2(n15962), .Q(n15960) );
  AND2X1 U16158 ( .IN1(n10067), .IN2(g6837), .Q(n15962) );
  AND2X1 U16159 ( .IN1(n10066), .IN2(test_so73), .Q(n15961) );
  AND2X1 U16160 ( .IN1(n9704), .IN2(g2241), .Q(n15959) );
  OR2X1 U16161 ( .IN1(n15963), .IN2(n15964), .Q(n15953) );
  AND2X1 U16162 ( .IN1(n15965), .IN2(g2170), .Q(n15964) );
  INVX0 U16163 ( .INP(n15966), .ZN(n15965) );
  AND2X1 U16164 ( .IN1(n4373), .IN2(n15966), .Q(n15963) );
  OR2X1 U16165 ( .IN1(n15967), .IN2(n15968), .Q(n15966) );
  OR2X1 U16166 ( .IN1(n15969), .IN2(n15970), .Q(n15968) );
  AND2X1 U16167 ( .IN1(n10065), .IN2(g6837), .Q(n15970) );
  AND2X1 U16168 ( .IN1(n10064), .IN2(test_so73), .Q(n15969) );
  AND2X1 U16169 ( .IN1(n9703), .IN2(g2241), .Q(n15967) );
  OR2X1 U16170 ( .IN1(n15971), .IN2(n15972), .Q(n15951) );
  AND2X1 U16171 ( .IN1(n15973), .IN2(n13206), .Q(n15972) );
  INVX0 U16172 ( .INP(n15974), .ZN(n15973) );
  AND2X1 U16173 ( .IN1(n11898), .IN2(n15974), .Q(n15971) );
  OR2X1 U16174 ( .IN1(n15975), .IN2(n15976), .Q(n15974) );
  OR2X1 U16175 ( .IN1(n15977), .IN2(n15978), .Q(n15976) );
  AND2X1 U16176 ( .IN1(n9695), .IN2(g2241), .Q(n15978) );
  AND2X1 U16177 ( .IN1(n9696), .IN2(g6837), .Q(n15977) );
  AND2X1 U16178 ( .IN1(test_so73), .IN2(n10215), .Q(n15975) );
  OR2X1 U16179 ( .IN1(n15979), .IN2(n15980), .Q(n15929) );
  OR2X1 U16180 ( .IN1(n15981), .IN2(n15982), .Q(n15980) );
  OR2X1 U16181 ( .IN1(n15983), .IN2(n15984), .Q(n15982) );
  OR2X1 U16182 ( .IN1(n15985), .IN2(n15986), .Q(n15984) );
  AND2X1 U16183 ( .IN1(n15987), .IN2(g2195), .Q(n15986) );
  INVX0 U16184 ( .INP(n15988), .ZN(n15987) );
  AND2X1 U16185 ( .IN1(n4563), .IN2(n15988), .Q(n15985) );
  OR2X1 U16186 ( .IN1(n15989), .IN2(n15990), .Q(n15988) );
  OR2X1 U16187 ( .IN1(n15991), .IN2(n15992), .Q(n15990) );
  AND2X1 U16188 ( .IN1(n10056), .IN2(g6837), .Q(n15992) );
  AND2X1 U16189 ( .IN1(n10055), .IN2(test_so73), .Q(n15991) );
  AND2X1 U16190 ( .IN1(n9698), .IN2(g2241), .Q(n15989) );
  OR2X1 U16191 ( .IN1(n15993), .IN2(n15994), .Q(n15983) );
  AND2X1 U16192 ( .IN1(n15995), .IN2(g2190), .Q(n15994) );
  INVX0 U16193 ( .INP(n15996), .ZN(n15995) );
  AND2X1 U16194 ( .IN1(n4555), .IN2(n15996), .Q(n15993) );
  OR2X1 U16195 ( .IN1(n15997), .IN2(n15998), .Q(n15996) );
  OR2X1 U16196 ( .IN1(n15999), .IN2(n16000), .Q(n15998) );
  AND2X1 U16197 ( .IN1(n10058), .IN2(g6837), .Q(n16000) );
  AND2X1 U16198 ( .IN1(n10057), .IN2(test_so73), .Q(n15999) );
  AND2X1 U16199 ( .IN1(n9699), .IN2(g2241), .Q(n15997) );
  OR2X1 U16200 ( .IN1(n16001), .IN2(n16002), .Q(n15981) );
  AND2X1 U16201 ( .IN1(n16003), .IN2(g2180), .Q(n16002) );
  INVX0 U16202 ( .INP(n16004), .ZN(n16003) );
  AND2X1 U16203 ( .IN1(n4389), .IN2(n16004), .Q(n16001) );
  OR2X1 U16204 ( .IN1(n16005), .IN2(n16006), .Q(n16004) );
  OR2X1 U16205 ( .IN1(n16007), .IN2(n16008), .Q(n16006) );
  AND2X1 U16206 ( .IN1(n10061), .IN2(g6837), .Q(n16008) );
  AND2X1 U16207 ( .IN1(n10060), .IN2(test_so73), .Q(n16007) );
  AND2X1 U16208 ( .IN1(n9701), .IN2(g2241), .Q(n16005) );
  OR2X1 U16209 ( .IN1(n16009), .IN2(n16010), .Q(n15979) );
  OR2X1 U16210 ( .IN1(n12248), .IN2(n16011), .Q(n16010) );
  OR2X1 U16211 ( .IN1(n16012), .IN2(n16013), .Q(n16011) );
  AND2X1 U16212 ( .IN1(n16014), .IN2(g2200), .Q(n16013) );
  INVX0 U16213 ( .INP(n16015), .ZN(n16014) );
  AND2X1 U16214 ( .IN1(n4287), .IN2(n16015), .Q(n16012) );
  OR2X1 U16215 ( .IN1(n16016), .IN2(n16017), .Q(n16015) );
  OR2X1 U16216 ( .IN1(n16018), .IN2(n16019), .Q(n16017) );
  AND2X1 U16217 ( .IN1(n10054), .IN2(g6837), .Q(n16019) );
  AND2X1 U16218 ( .IN1(n10053), .IN2(test_so73), .Q(n16018) );
  AND2X1 U16219 ( .IN1(n9697), .IN2(g2241), .Q(n16016) );
  INVX0 U16220 ( .INP(n3038), .ZN(n12248) );
  OR2X1 U16221 ( .IN1(n16020), .IN2(n16021), .Q(n16009) );
  AND2X1 U16222 ( .IN1(n16022), .IN2(g2185), .Q(n16021) );
  INVX0 U16223 ( .INP(n16023), .ZN(n16022) );
  AND2X1 U16224 ( .IN1(n4325), .IN2(n16023), .Q(n16020) );
  OR2X1 U16225 ( .IN1(n16024), .IN2(n16025), .Q(n16023) );
  OR2X1 U16226 ( .IN1(n16026), .IN2(n16027), .Q(n16025) );
  AND2X1 U16227 ( .IN1(n9700), .IN2(g2241), .Q(n16027) );
  AND2X1 U16228 ( .IN1(n10059), .IN2(g6837), .Q(n16026) );
  AND2X1 U16229 ( .IN1(test_so73), .IN2(n10216), .Q(n16024) );
  OR2X1 U16230 ( .IN1(n16028), .IN2(n16029), .Q(n12925) );
  OR2X1 U16231 ( .IN1(n16030), .IN2(n16031), .Q(n16029) );
  AND2X1 U16232 ( .IN1(n9852), .IN2(n13116), .Q(n16031) );
  AND2X1 U16233 ( .IN1(n13101), .IN2(n10217), .Q(n16030) );
  AND2X1 U16234 ( .IN1(n9843), .IN2(n13106), .Q(n16028) );
  AND2X1 U16235 ( .IN1(n16032), .IN2(n4526), .Q(g25940) );
  AND2X1 U16236 ( .IN1(n16033), .IN2(n12966), .Q(n16032) );
  OR2X1 U16237 ( .IN1(n3887), .IN2(test_so78), .Q(n16033) );
  AND2X1 U16238 ( .IN1(n16034), .IN2(n4527), .Q(g25938) );
  AND2X1 U16239 ( .IN1(n16035), .IN2(n12971), .Q(n16034) );
  OR2X1 U16240 ( .IN1(n3890), .IN2(g1462), .Q(n16035) );
  AND2X1 U16241 ( .IN1(n16036), .IN2(n12976), .Q(g25935) );
  AND2X1 U16242 ( .IN1(n16037), .IN2(n879), .Q(n16036) );
  OR2X1 U16243 ( .IN1(n10172), .IN2(n16038), .Q(n879) );
  INVX0 U16244 ( .INP(n3893), .ZN(n16038) );
  OR2X1 U16245 ( .IN1(n3893), .IN2(g776), .Q(n16037) );
  AND2X1 U16246 ( .IN1(n16039), .IN2(n4528), .Q(g25932) );
  AND2X1 U16247 ( .IN1(n16040), .IN2(n12981), .Q(n16039) );
  OR2X1 U16248 ( .IN1(n3896), .IN2(g88), .Q(n16040) );
  OR2X1 U16249 ( .IN1(n16041), .IN2(n16042), .Q(g25489) );
  AND2X1 U16250 ( .IN1(n16043), .IN2(test_so10), .Q(n16042) );
  AND2X1 U16251 ( .IN1(n16044), .IN2(g3142), .Q(n16043) );
  AND2X1 U16252 ( .IN1(g3151), .IN2(g3097), .Q(n16044) );
  AND2X1 U16253 ( .IN1(n16045), .IN2(n10202), .Q(n16041) );
  OR2X1 U16254 ( .IN1(n16046), .IN2(n16047), .Q(n16045) );
  AND2X1 U16255 ( .IN1(n4301), .IN2(n14520), .Q(n16047) );
  OR2X1 U16256 ( .IN1(test_so1), .IN2(n8099), .Q(n14520) );
  AND2X1 U16257 ( .IN1(n4424), .IN2(n16048), .Q(n16046) );
  OR2X1 U16258 ( .IN1(n4301), .IN2(n14519), .Q(n16048) );
  OR2X1 U16259 ( .IN1(n4577), .IN2(n4578), .Q(n14519) );
  OR2X1 U16260 ( .IN1(n16049), .IN2(n16050), .Q(g25452) );
  AND2X1 U16261 ( .IN1(g21851), .IN2(g3109), .Q(n16050) );
  AND2X1 U16262 ( .IN1(n4494), .IN2(g3099), .Q(n16049) );
  OR2X1 U16263 ( .IN1(n16051), .IN2(n16052), .Q(g25451) );
  AND2X1 U16264 ( .IN1(g21851), .IN2(g8030), .Q(n16052) );
  AND2X1 U16265 ( .IN1(n4383), .IN2(g3098), .Q(n16051) );
  OR2X1 U16266 ( .IN1(n16053), .IN2(n16054), .Q(g25450) );
  AND2X1 U16267 ( .IN1(g21851), .IN2(g8106), .Q(n16054) );
  AND2X1 U16268 ( .IN1(n4382), .IN2(g3097), .Q(n16053) );
  OR2X1 U16269 ( .IN1(n14497), .IN2(n16055), .Q(g25442) );
  OR2X1 U16270 ( .IN1(n16056), .IN2(n16057), .Q(n16055) );
  AND2X1 U16271 ( .IN1(n14501), .IN2(g3124), .Q(n16057) );
  AND2X1 U16272 ( .IN1(n15804), .IN2(g3111), .Q(n16056) );
  OR2X1 U16273 ( .IN1(n14497), .IN2(n16058), .Q(g25435) );
  OR2X1 U16274 ( .IN1(n16059), .IN2(n16060), .Q(n16058) );
  AND2X1 U16275 ( .IN1(n14501), .IN2(DFF_144_n1), .Q(n16060) );
  AND2X1 U16276 ( .IN1(n15804), .IN2(g3110), .Q(n16059) );
  OR2X1 U16277 ( .IN1(n14497), .IN2(n16061), .Q(g25420) );
  OR2X1 U16278 ( .IN1(n16062), .IN2(n16063), .Q(n16061) );
  AND2X1 U16279 ( .IN1(test_so9), .IN2(n14501), .Q(n16063) );
  AND2X1 U16280 ( .IN1(n15804), .IN2(g3112), .Q(n16062) );
  AND2X1 U16281 ( .IN1(n15822), .IN2(n15888), .Q(n15804) );
  AND2X1 U16282 ( .IN1(g3204), .IN2(n4073), .Q(n15888) );
  AND2X1 U16283 ( .IN1(n15829), .IN2(n4405), .Q(n15822) );
  AND2X1 U16284 ( .IN1(n4329), .IN2(n4406), .Q(n15829) );
  OR2X1 U16285 ( .IN1(n16064), .IN2(n16065), .Q(g25288) );
  AND2X1 U16286 ( .IN1(n16066), .IN2(n16067), .Q(n16065) );
  AND2X1 U16287 ( .IN1(n16068), .IN2(g2808), .Q(n16064) );
  OR2X1 U16288 ( .IN1(n16069), .IN2(n16070), .Q(g25280) );
  AND2X1 U16289 ( .IN1(n16071), .IN2(g2810), .Q(n16070) );
  AND2X1 U16290 ( .IN1(n16072), .IN2(n16066), .Q(n16069) );
  OR2X1 U16291 ( .IN1(n16073), .IN2(n16074), .Q(g25279) );
  AND2X1 U16292 ( .IN1(n16075), .IN2(n4149), .Q(n16074) );
  AND2X1 U16293 ( .IN1(n16076), .IN2(g2114), .Q(n16073) );
  OR2X1 U16294 ( .IN1(n16077), .IN2(n16078), .Q(g25272) );
  AND2X1 U16295 ( .IN1(n16079), .IN2(g2809), .Q(n16078) );
  AND2X1 U16296 ( .IN1(n16080), .IN2(n16066), .Q(n16077) );
  INVX0 U16297 ( .INP(n16081), .ZN(n16066) );
  OR2X1 U16298 ( .IN1(n16082), .IN2(n16083), .Q(n16081) );
  OR2X1 U16299 ( .IN1(n16084), .IN2(n11670), .Q(n16083) );
  OR2X1 U16300 ( .IN1(n16085), .IN2(n16086), .Q(n11670) );
  OR2X1 U16301 ( .IN1(n16087), .IN2(n16088), .Q(n16086) );
  AND2X1 U16302 ( .IN1(n9747), .IN2(g7425), .Q(n16088) );
  AND2X1 U16303 ( .IN1(n9802), .IN2(g2703), .Q(n16087) );
  AND2X1 U16304 ( .IN1(n9739), .IN2(g7487), .Q(n16085) );
  AND2X1 U16305 ( .IN1(n9740), .IN2(g7487), .Q(n16084) );
  OR2X1 U16306 ( .IN1(n16089), .IN2(n16090), .Q(n16082) );
  OR2X1 U16307 ( .IN1(n16091), .IN2(n16092), .Q(n16090) );
  AND2X1 U16308 ( .IN1(n9803), .IN2(g2703), .Q(n16092) );
  AND2X1 U16309 ( .IN1(n16093), .IN2(n16094), .Q(n16091) );
  AND2X1 U16310 ( .IN1(n16095), .IN2(n16096), .Q(n16094) );
  AND2X1 U16311 ( .IN1(n16097), .IN2(n16098), .Q(n16096) );
  AND2X1 U16312 ( .IN1(n16099), .IN2(n16100), .Q(n16098) );
  OR2X1 U16313 ( .IN1(n11154), .IN2(g2707), .Q(n16100) );
  INVX0 U16314 ( .INP(n11155), .ZN(n11154) );
  OR2X1 U16315 ( .IN1(n4472), .IN2(n11155), .Q(n16099) );
  OR2X1 U16316 ( .IN1(n16101), .IN2(n16102), .Q(n11155) );
  OR2X1 U16317 ( .IN1(n16103), .IN2(n16104), .Q(n16102) );
  AND2X1 U16318 ( .IN1(n9954), .IN2(g7425), .Q(n16104) );
  AND2X1 U16319 ( .IN1(n10017), .IN2(g2703), .Q(n16103) );
  AND2X1 U16320 ( .IN1(n9953), .IN2(g7487), .Q(n16101) );
  AND2X1 U16321 ( .IN1(n16105), .IN2(n16106), .Q(n16097) );
  OR2X1 U16322 ( .IN1(n16107), .IN2(n16108), .Q(n16106) );
  AND2X1 U16323 ( .IN1(n11189), .IN2(n10192), .Q(n16108) );
  INVX0 U16324 ( .INP(n11188), .ZN(n11189) );
  AND2X1 U16325 ( .IN1(test_so92), .IN2(n11188), .Q(n16107) );
  OR2X1 U16326 ( .IN1(n16109), .IN2(n16110), .Q(n11188) );
  OR2X1 U16327 ( .IN1(n16111), .IN2(n16112), .Q(n16110) );
  AND2X1 U16328 ( .IN1(n9944), .IN2(g7425), .Q(n16112) );
  AND2X1 U16329 ( .IN1(n10013), .IN2(g2703), .Q(n16111) );
  AND2X1 U16330 ( .IN1(n9943), .IN2(g7487), .Q(n16109) );
  AND2X1 U16331 ( .IN1(n16113), .IN2(n16114), .Q(n16105) );
  OR2X1 U16332 ( .IN1(n11194), .IN2(g2714), .Q(n16114) );
  INVX0 U16333 ( .INP(n11193), .ZN(n11194) );
  OR2X1 U16334 ( .IN1(n4398), .IN2(n11193), .Q(n16113) );
  OR2X1 U16335 ( .IN1(n16115), .IN2(n16116), .Q(n11193) );
  OR2X1 U16336 ( .IN1(n16117), .IN2(n16118), .Q(n16116) );
  AND2X1 U16337 ( .IN1(n9956), .IN2(g7425), .Q(n16118) );
  AND2X1 U16338 ( .IN1(n10018), .IN2(g2703), .Q(n16117) );
  AND2X1 U16339 ( .IN1(n9955), .IN2(g7487), .Q(n16115) );
  AND2X1 U16340 ( .IN1(n16119), .IN2(n16120), .Q(n16095) );
  AND2X1 U16341 ( .IN1(n16121), .IN2(n16122), .Q(n16120) );
  OR2X1 U16342 ( .IN1(n11145), .IN2(g2734), .Q(n16122) );
  INVX0 U16343 ( .INP(n11144), .ZN(n11145) );
  OR2X1 U16344 ( .IN1(n4397), .IN2(n11144), .Q(n16121) );
  OR2X1 U16345 ( .IN1(n16123), .IN2(n16124), .Q(n11144) );
  OR2X1 U16346 ( .IN1(n16125), .IN2(n16126), .Q(n16124) );
  AND2X1 U16347 ( .IN1(n9948), .IN2(g7425), .Q(n16126) );
  AND2X1 U16348 ( .IN1(n10015), .IN2(g2703), .Q(n16125) );
  AND2X1 U16349 ( .IN1(n9947), .IN2(g7487), .Q(n16123) );
  AND2X1 U16350 ( .IN1(n16127), .IN2(n16128), .Q(n16119) );
  OR2X1 U16351 ( .IN1(n11173), .IN2(g2746), .Q(n16128) );
  INVX0 U16352 ( .INP(n11174), .ZN(n11173) );
  OR2X1 U16353 ( .IN1(n4407), .IN2(n11174), .Q(n16127) );
  OR2X1 U16354 ( .IN1(n16129), .IN2(n16130), .Q(n11174) );
  OR2X1 U16355 ( .IN1(n16131), .IN2(n16132), .Q(n16130) );
  AND2X1 U16356 ( .IN1(n9946), .IN2(g7425), .Q(n16132) );
  AND2X1 U16357 ( .IN1(n10014), .IN2(g2703), .Q(n16131) );
  AND2X1 U16358 ( .IN1(n9945), .IN2(g7487), .Q(n16129) );
  AND2X1 U16359 ( .IN1(n16133), .IN2(n16134), .Q(n16093) );
  AND2X1 U16360 ( .IN1(n16135), .IN2(n16136), .Q(n16134) );
  AND2X1 U16361 ( .IN1(n16137), .IN2(n16138), .Q(n16136) );
  OR2X1 U16362 ( .IN1(n11159), .IN2(g2753), .Q(n16138) );
  INVX0 U16363 ( .INP(n11160), .ZN(n11159) );
  OR2X1 U16364 ( .IN1(n4471), .IN2(n11160), .Q(n16137) );
  OR2X1 U16365 ( .IN1(n16139), .IN2(n16140), .Q(n11160) );
  OR2X1 U16366 ( .IN1(n16141), .IN2(n16142), .Q(n16140) );
  AND2X1 U16367 ( .IN1(n9942), .IN2(g7425), .Q(n16142) );
  AND2X1 U16368 ( .IN1(n10012), .IN2(g2703), .Q(n16141) );
  AND2X1 U16369 ( .IN1(n9941), .IN2(g7487), .Q(n16139) );
  AND2X1 U16370 ( .IN1(n16143), .IN2(n16144), .Q(n16135) );
  AND2X1 U16371 ( .IN1(n16145), .IN2(n16146), .Q(n16144) );
  INVX0 U16372 ( .INP(n16147), .ZN(n16146) );
  AND2X1 U16373 ( .IN1(n11211), .IN2(n4415), .Q(n16147) );
  OR2X1 U16374 ( .IN1(n4415), .IN2(n11211), .Q(n16145) );
  OR2X1 U16375 ( .IN1(n16148), .IN2(n16149), .Q(n11211) );
  OR2X1 U16376 ( .IN1(n16150), .IN2(n16151), .Q(n16149) );
  AND2X1 U16377 ( .IN1(n9938), .IN2(g7425), .Q(n16151) );
  AND2X1 U16378 ( .IN1(n10011), .IN2(g2703), .Q(n16150) );
  AND2X1 U16379 ( .IN1(n9937), .IN2(g7487), .Q(n16148) );
  AND2X1 U16380 ( .IN1(n16152), .IN2(n16153), .Q(n16143) );
  INVX0 U16381 ( .INP(n16154), .ZN(n16153) );
  AND2X1 U16382 ( .IN1(n11221), .IN2(n4393), .Q(n16154) );
  OR2X1 U16383 ( .IN1(n4393), .IN2(n11221), .Q(n16152) );
  OR2X1 U16384 ( .IN1(n16155), .IN2(n16156), .Q(n11221) );
  OR2X1 U16385 ( .IN1(n16157), .IN2(n16158), .Q(n16156) );
  AND2X1 U16386 ( .IN1(n9940), .IN2(g7425), .Q(n16158) );
  AND2X1 U16387 ( .IN1(g2703), .IN2(n10218), .Q(n16157) );
  AND2X1 U16388 ( .IN1(n9939), .IN2(g7487), .Q(n16155) );
  AND2X1 U16389 ( .IN1(n16159), .IN2(n16160), .Q(n16133) );
  AND2X1 U16390 ( .IN1(n16161), .IN2(n16162), .Q(n16160) );
  OR2X1 U16391 ( .IN1(n11135), .IN2(g2720), .Q(n16162) );
  INVX0 U16392 ( .INP(n11138), .ZN(n11135) );
  OR2X1 U16393 ( .IN1(n4408), .IN2(n11138), .Q(n16161) );
  OR2X1 U16394 ( .IN1(n16163), .IN2(n16164), .Q(n11138) );
  OR2X1 U16395 ( .IN1(n16165), .IN2(n16166), .Q(n16164) );
  AND2X1 U16396 ( .IN1(n9950), .IN2(g7425), .Q(n16166) );
  AND2X1 U16397 ( .IN1(g2703), .IN2(n10219), .Q(n16165) );
  AND2X1 U16398 ( .IN1(n9949), .IN2(g7487), .Q(n16163) );
  AND2X1 U16399 ( .IN1(n16167), .IN2(n16168), .Q(n16159) );
  OR2X1 U16400 ( .IN1(n11180), .IN2(g2727), .Q(n16168) );
  INVX0 U16401 ( .INP(n11179), .ZN(n11180) );
  OR2X1 U16402 ( .IN1(n4419), .IN2(n11179), .Q(n16167) );
  OR2X1 U16403 ( .IN1(n16169), .IN2(n16170), .Q(n11179) );
  OR2X1 U16404 ( .IN1(n16171), .IN2(n16172), .Q(n16170) );
  AND2X1 U16405 ( .IN1(n9952), .IN2(g7425), .Q(n16172) );
  AND2X1 U16406 ( .IN1(n10016), .IN2(g2703), .Q(n16171) );
  AND2X1 U16407 ( .IN1(n9951), .IN2(g7487), .Q(n16169) );
  AND2X1 U16408 ( .IN1(n9748), .IN2(g7425), .Q(n16089) );
  OR2X1 U16409 ( .IN1(n16173), .IN2(n16174), .Q(g25271) );
  AND2X1 U16410 ( .IN1(n16175), .IN2(n16075), .Q(n16174) );
  AND2X1 U16411 ( .IN1(n16176), .IN2(g2116), .Q(n16173) );
  OR2X1 U16412 ( .IN1(n16177), .IN2(n16178), .Q(g25270) );
  AND2X1 U16413 ( .IN1(n16179), .IN2(n16180), .Q(n16178) );
  AND2X1 U16414 ( .IN1(n16181), .IN2(g1420), .Q(n16177) );
  OR2X1 U16415 ( .IN1(n16182), .IN2(n16183), .Q(g25268) );
  AND2X1 U16416 ( .IN1(n16184), .IN2(n16075), .Q(n16183) );
  INVX0 U16417 ( .INP(n16185), .ZN(n16075) );
  OR2X1 U16418 ( .IN1(n16186), .IN2(n16187), .Q(n16185) );
  OR2X1 U16419 ( .IN1(n16188), .IN2(n11699), .Q(n16187) );
  OR2X1 U16420 ( .IN1(n16189), .IN2(n16190), .Q(n11699) );
  OR2X1 U16421 ( .IN1(n16191), .IN2(n16192), .Q(n16190) );
  AND2X1 U16422 ( .IN1(n9749), .IN2(g7229), .Q(n16192) );
  AND2X1 U16423 ( .IN1(n9804), .IN2(g2009), .Q(n16191) );
  AND2X1 U16424 ( .IN1(n9741), .IN2(g7357), .Q(n16189) );
  AND2X1 U16425 ( .IN1(n9742), .IN2(g7357), .Q(n16188) );
  OR2X1 U16426 ( .IN1(n16193), .IN2(n16194), .Q(n16186) );
  OR2X1 U16427 ( .IN1(n16195), .IN2(n16196), .Q(n16194) );
  AND2X1 U16428 ( .IN1(n9805), .IN2(g2009), .Q(n16196) );
  AND2X1 U16429 ( .IN1(n16197), .IN2(n16198), .Q(n16195) );
  AND2X1 U16430 ( .IN1(n16199), .IN2(n16200), .Q(n16198) );
  AND2X1 U16431 ( .IN1(n16201), .IN2(n16202), .Q(n16200) );
  AND2X1 U16432 ( .IN1(n16203), .IN2(n16204), .Q(n16202) );
  OR2X1 U16433 ( .IN1(n11317), .IN2(g2013), .Q(n16204) );
  INVX0 U16434 ( .INP(n11318), .ZN(n11317) );
  OR2X1 U16435 ( .IN1(n4474), .IN2(n11318), .Q(n16203) );
  OR2X1 U16436 ( .IN1(n16205), .IN2(n16206), .Q(n11318) );
  OR2X1 U16437 ( .IN1(n16207), .IN2(n16208), .Q(n16206) );
  AND2X1 U16438 ( .IN1(n9972), .IN2(g7229), .Q(n16208) );
  AND2X1 U16439 ( .IN1(n10027), .IN2(g2009), .Q(n16207) );
  AND2X1 U16440 ( .IN1(n9971), .IN2(g7357), .Q(n16205) );
  AND2X1 U16441 ( .IN1(n16209), .IN2(n16210), .Q(n16201) );
  OR2X1 U16442 ( .IN1(n16211), .IN2(n16212), .Q(n16210) );
  AND2X1 U16443 ( .IN1(n11384), .IN2(n10194), .Q(n16212) );
  INVX0 U16444 ( .INP(n11382), .ZN(n11384) );
  AND2X1 U16445 ( .IN1(test_so70), .IN2(n11382), .Q(n16211) );
  OR2X1 U16446 ( .IN1(n16213), .IN2(n16214), .Q(n11382) );
  OR2X1 U16447 ( .IN1(n16215), .IN2(n16216), .Q(n16214) );
  AND2X1 U16448 ( .IN1(n9959), .IN2(g7229), .Q(n16216) );
  AND2X1 U16449 ( .IN1(n10020), .IN2(g2009), .Q(n16215) );
  AND2X1 U16450 ( .IN1(n9958), .IN2(g7357), .Q(n16213) );
  AND2X1 U16451 ( .IN1(n16217), .IN2(n16218), .Q(n16209) );
  OR2X1 U16452 ( .IN1(n11322), .IN2(g2059), .Q(n16218) );
  INVX0 U16453 ( .INP(n11323), .ZN(n11322) );
  OR2X1 U16454 ( .IN1(n4473), .IN2(n11323), .Q(n16217) );
  OR2X1 U16455 ( .IN1(n16219), .IN2(n16220), .Q(n11323) );
  OR2X1 U16456 ( .IN1(n16221), .IN2(n16222), .Q(n16220) );
  AND2X1 U16457 ( .IN1(n9961), .IN2(g7229), .Q(n16222) );
  AND2X1 U16458 ( .IN1(n10021), .IN2(g2009), .Q(n16221) );
  AND2X1 U16459 ( .IN1(n9960), .IN2(g7357), .Q(n16219) );
  AND2X1 U16460 ( .IN1(n16223), .IN2(n16224), .Q(n16199) );
  AND2X1 U16461 ( .IN1(n16225), .IN2(n16226), .Q(n16224) );
  OR2X1 U16462 ( .IN1(n11352), .IN2(g2046), .Q(n16226) );
  INVX0 U16463 ( .INP(n11351), .ZN(n11352) );
  OR2X1 U16464 ( .IN1(n4468), .IN2(n11351), .Q(n16225) );
  OR2X1 U16465 ( .IN1(n16227), .IN2(n16228), .Q(n11351) );
  OR2X1 U16466 ( .IN1(n16229), .IN2(n16230), .Q(n16228) );
  AND2X1 U16467 ( .IN1(n9963), .IN2(g7229), .Q(n16230) );
  AND2X1 U16468 ( .IN1(n10022), .IN2(g2009), .Q(n16229) );
  AND2X1 U16469 ( .IN1(n9962), .IN2(g7357), .Q(n16227) );
  AND2X1 U16470 ( .IN1(n16231), .IN2(n16232), .Q(n16223) );
  OR2X1 U16471 ( .IN1(n11298), .IN2(g2026), .Q(n16232) );
  INVX0 U16472 ( .INP(n11301), .ZN(n11298) );
  OR2X1 U16473 ( .IN1(n4410), .IN2(n11301), .Q(n16231) );
  OR2X1 U16474 ( .IN1(n16233), .IN2(n16234), .Q(n11301) );
  OR2X1 U16475 ( .IN1(n16235), .IN2(n16236), .Q(n16234) );
  AND2X1 U16476 ( .IN1(n9968), .IN2(g7229), .Q(n16236) );
  AND2X1 U16477 ( .IN1(n10025), .IN2(g2009), .Q(n16235) );
  AND2X1 U16478 ( .IN1(n9967), .IN2(g7357), .Q(n16233) );
  AND2X1 U16479 ( .IN1(n16237), .IN2(n16238), .Q(n16197) );
  AND2X1 U16480 ( .IN1(n16239), .IN2(n16240), .Q(n16238) );
  AND2X1 U16481 ( .IN1(n16241), .IN2(n16242), .Q(n16240) );
  OR2X1 U16482 ( .IN1(n11308), .IN2(g2040), .Q(n16242) );
  INVX0 U16483 ( .INP(n11307), .ZN(n11308) );
  OR2X1 U16484 ( .IN1(n4399), .IN2(n11307), .Q(n16241) );
  OR2X1 U16485 ( .IN1(n16243), .IN2(n16244), .Q(n11307) );
  OR2X1 U16486 ( .IN1(n16245), .IN2(n16246), .Q(n16244) );
  AND2X1 U16487 ( .IN1(n9966), .IN2(g7229), .Q(n16246) );
  AND2X1 U16488 ( .IN1(n10024), .IN2(g2009), .Q(n16245) );
  INVX0 U16489 ( .INP(n16247), .ZN(n16243) );
  OR2X1 U16490 ( .IN1(n4357), .IN2(test_so71), .Q(n16247) );
  AND2X1 U16491 ( .IN1(n16248), .IN2(n16249), .Q(n16239) );
  AND2X1 U16492 ( .IN1(n16250), .IN2(n16251), .Q(n16249) );
  OR2X1 U16493 ( .IN1(n11372), .IN2(g2072), .Q(n16251) );
  INVX0 U16494 ( .INP(n11373), .ZN(n11372) );
  OR2X1 U16495 ( .IN1(n4416), .IN2(n11373), .Q(n16250) );
  OR2X1 U16496 ( .IN1(n16252), .IN2(n16253), .Q(n11373) );
  OR2X1 U16497 ( .IN1(n16254), .IN2(n16255), .Q(n16253) );
  AND2X1 U16498 ( .IN1(n9957), .IN2(g7229), .Q(n16255) );
  AND2X1 U16499 ( .IN1(n10019), .IN2(g2009), .Q(n16254) );
  INVX0 U16500 ( .INP(n16256), .ZN(n16252) );
  OR2X1 U16501 ( .IN1(n4357), .IN2(test_so72), .Q(n16256) );
  AND2X1 U16502 ( .IN1(n16257), .IN2(n16258), .Q(n16248) );
  OR2X1 U16503 ( .IN1(n11336), .IN2(g2052), .Q(n16258) );
  INVX0 U16504 ( .INP(n11337), .ZN(n11336) );
  OR2X1 U16505 ( .IN1(n4409), .IN2(n11337), .Q(n16257) );
  OR2X1 U16506 ( .IN1(n16259), .IN2(n16260), .Q(n11337) );
  OR2X1 U16507 ( .IN1(n16261), .IN2(n16262), .Q(n16260) );
  AND2X1 U16508 ( .IN1(n9965), .IN2(g7229), .Q(n16262) );
  AND2X1 U16509 ( .IN1(n10023), .IN2(g2009), .Q(n16261) );
  AND2X1 U16510 ( .IN1(n9964), .IN2(g7357), .Q(n16259) );
  AND2X1 U16511 ( .IN1(n16263), .IN2(n16264), .Q(n16237) );
  AND2X1 U16512 ( .IN1(n16265), .IN2(n16266), .Q(n16264) );
  OR2X1 U16513 ( .IN1(n11357), .IN2(g2020), .Q(n16266) );
  INVX0 U16514 ( .INP(n11356), .ZN(n11357) );
  OR2X1 U16515 ( .IN1(n4400), .IN2(n11356), .Q(n16265) );
  OR2X1 U16516 ( .IN1(n16267), .IN2(n16268), .Q(n11356) );
  OR2X1 U16517 ( .IN1(n16269), .IN2(n16270), .Q(n16268) );
  AND2X1 U16518 ( .IN1(n9974), .IN2(g7229), .Q(n16270) );
  AND2X1 U16519 ( .IN1(n10028), .IN2(g2009), .Q(n16269) );
  AND2X1 U16520 ( .IN1(n9973), .IN2(g7357), .Q(n16267) );
  AND2X1 U16521 ( .IN1(n16271), .IN2(n16272), .Q(n16263) );
  OR2X1 U16522 ( .IN1(n11343), .IN2(g2033), .Q(n16272) );
  INVX0 U16523 ( .INP(n11342), .ZN(n11343) );
  OR2X1 U16524 ( .IN1(n4420), .IN2(n11342), .Q(n16271) );
  OR2X1 U16525 ( .IN1(n16273), .IN2(n16274), .Q(n11342) );
  OR2X1 U16526 ( .IN1(n16275), .IN2(n16276), .Q(n16274) );
  AND2X1 U16527 ( .IN1(n9970), .IN2(g7229), .Q(n16276) );
  AND2X1 U16528 ( .IN1(n10026), .IN2(g2009), .Q(n16275) );
  AND2X1 U16529 ( .IN1(n9969), .IN2(g7357), .Q(n16273) );
  AND2X1 U16530 ( .IN1(n9750), .IN2(g7229), .Q(n16193) );
  AND2X1 U16531 ( .IN1(n16277), .IN2(g2115), .Q(n16182) );
  OR2X1 U16532 ( .IN1(n16278), .IN2(n16279), .Q(g25267) );
  AND2X1 U16533 ( .IN1(n1027), .IN2(n16179), .Q(n16279) );
  AND2X1 U16534 ( .IN1(n16280), .IN2(g1422), .Q(n16278) );
  OR2X1 U16535 ( .IN1(n16281), .IN2(n16282), .Q(g25266) );
  AND2X1 U16536 ( .IN1(n16283), .IN2(n680), .Q(n16282) );
  AND2X1 U16537 ( .IN1(n16284), .IN2(g734), .Q(n16281) );
  OR2X1 U16538 ( .IN1(n16285), .IN2(n16286), .Q(g25265) );
  INVX0 U16539 ( .INP(n15910), .ZN(n16286) );
  OR2X1 U16540 ( .IN1(n15352), .IN2(g3234), .Q(n15910) );
  AND2X1 U16541 ( .IN1(n15352), .IN2(n16287), .Q(n16285) );
  OR2X1 U16542 ( .IN1(n16288), .IN2(n16289), .Q(n16287) );
  AND2X1 U16543 ( .IN1(n10165), .IN2(g2993), .Q(n16289) );
  AND2X1 U16544 ( .IN1(n10166), .IN2(n4598), .Q(n16288) );
  OR2X1 U16545 ( .IN1(n16290), .IN2(n16291), .Q(g25263) );
  AND2X1 U16546 ( .IN1(n16292), .IN2(g1421), .Q(n16291) );
  AND2X1 U16547 ( .IN1(n16293), .IN2(n16179), .Q(n16290) );
  INVX0 U16548 ( .INP(n16294), .ZN(n16179) );
  OR2X1 U16549 ( .IN1(n16295), .IN2(n16296), .Q(n16294) );
  OR2X1 U16550 ( .IN1(n16297), .IN2(n11724), .Q(n16296) );
  OR2X1 U16551 ( .IN1(n16298), .IN2(n16299), .Q(n11724) );
  OR2X1 U16552 ( .IN1(n16300), .IN2(n16301), .Q(n16299) );
  AND2X1 U16553 ( .IN1(n9751), .IN2(g6979), .Q(n16301) );
  AND2X1 U16554 ( .IN1(n9806), .IN2(g1315), .Q(n16300) );
  AND2X1 U16555 ( .IN1(n9743), .IN2(g7161), .Q(n16298) );
  AND2X1 U16556 ( .IN1(n9744), .IN2(g7161), .Q(n16297) );
  OR2X1 U16557 ( .IN1(n16302), .IN2(n16303), .Q(n16295) );
  OR2X1 U16558 ( .IN1(n16304), .IN2(n16305), .Q(n16303) );
  AND2X1 U16559 ( .IN1(g1315), .IN2(n10220), .Q(n16305) );
  AND2X1 U16560 ( .IN1(n16306), .IN2(n16307), .Q(n16304) );
  AND2X1 U16561 ( .IN1(n16308), .IN2(n16309), .Q(n16307) );
  AND2X1 U16562 ( .IN1(n16310), .IN2(n16311), .Q(n16309) );
  AND2X1 U16563 ( .IN1(n16312), .IN2(n16313), .Q(n16311) );
  OR2X1 U16564 ( .IN1(n11484), .IN2(g1365), .Q(n16313) );
  INVX0 U16565 ( .INP(n11485), .ZN(n11484) );
  OR2X1 U16566 ( .IN1(n4475), .IN2(n11485), .Q(n16312) );
  OR2X1 U16567 ( .IN1(n16314), .IN2(n16315), .Q(n11485) );
  OR2X1 U16568 ( .IN1(n16316), .IN2(n16317), .Q(n16315) );
  AND2X1 U16569 ( .IN1(n9980), .IN2(g6979), .Q(n16317) );
  AND2X1 U16570 ( .IN1(n10031), .IN2(g1315), .Q(n16316) );
  AND2X1 U16571 ( .IN1(n9979), .IN2(g7161), .Q(n16314) );
  AND2X1 U16572 ( .IN1(n16318), .IN2(n16319), .Q(n16310) );
  AND2X1 U16573 ( .IN1(n16320), .IN2(n16321), .Q(n16319) );
  OR2X1 U16574 ( .IN1(n11514), .IN2(g1352), .Q(n16321) );
  INVX0 U16575 ( .INP(n11513), .ZN(n11514) );
  OR2X1 U16576 ( .IN1(n4469), .IN2(n11513), .Q(n16320) );
  OR2X1 U16577 ( .IN1(n16322), .IN2(n16323), .Q(n11513) );
  OR2X1 U16578 ( .IN1(n16324), .IN2(n16325), .Q(n16323) );
  AND2X1 U16579 ( .IN1(n9982), .IN2(g6979), .Q(n16325) );
  AND2X1 U16580 ( .IN1(n10032), .IN2(g1315), .Q(n16324) );
  AND2X1 U16581 ( .IN1(n9981), .IN2(g7161), .Q(n16322) );
  AND2X1 U16582 ( .IN1(n16326), .IN2(n16327), .Q(n16318) );
  OR2X1 U16583 ( .IN1(n11479), .IN2(g1319), .Q(n16327) );
  INVX0 U16584 ( .INP(n11480), .ZN(n11479) );
  OR2X1 U16585 ( .IN1(n4476), .IN2(n11480), .Q(n16326) );
  OR2X1 U16586 ( .IN1(n16328), .IN2(n16329), .Q(n11480) );
  OR2X1 U16587 ( .IN1(n16330), .IN2(n16331), .Q(n16329) );
  AND2X1 U16588 ( .IN1(n9991), .IN2(g6979), .Q(n16331) );
  AND2X1 U16589 ( .IN1(n10037), .IN2(g1315), .Q(n16330) );
  AND2X1 U16590 ( .IN1(n9990), .IN2(g7161), .Q(n16328) );
  AND2X1 U16591 ( .IN1(n16332), .IN2(n16333), .Q(n16308) );
  AND2X1 U16592 ( .IN1(n16334), .IN2(n16335), .Q(n16333) );
  OR2X1 U16593 ( .IN1(n11460), .IN2(g1332), .Q(n16335) );
  INVX0 U16594 ( .INP(n11463), .ZN(n11460) );
  OR2X1 U16595 ( .IN1(n4412), .IN2(n11463), .Q(n16334) );
  OR2X1 U16596 ( .IN1(n16336), .IN2(n16337), .Q(n11463) );
  OR2X1 U16597 ( .IN1(n16338), .IN2(n16339), .Q(n16337) );
  AND2X1 U16598 ( .IN1(n9987), .IN2(g6979), .Q(n16339) );
  AND2X1 U16599 ( .IN1(n10035), .IN2(g1315), .Q(n16338) );
  AND2X1 U16600 ( .IN1(n9986), .IN2(g7161), .Q(n16336) );
  AND2X1 U16601 ( .IN1(n16340), .IN2(n16341), .Q(n16332) );
  OR2X1 U16602 ( .IN1(n11535), .IN2(g1378), .Q(n16341) );
  INVX0 U16603 ( .INP(n11536), .ZN(n11535) );
  OR2X1 U16604 ( .IN1(n4417), .IN2(n11536), .Q(n16340) );
  OR2X1 U16605 ( .IN1(n16342), .IN2(n16343), .Q(n11536) );
  OR2X1 U16606 ( .IN1(n16344), .IN2(n16345), .Q(n16343) );
  AND2X1 U16607 ( .IN1(n9976), .IN2(g6979), .Q(n16345) );
  AND2X1 U16608 ( .IN1(n10029), .IN2(g1315), .Q(n16344) );
  AND2X1 U16609 ( .IN1(n9975), .IN2(g7161), .Q(n16342) );
  AND2X1 U16610 ( .IN1(n16346), .IN2(n16347), .Q(n16306) );
  AND2X1 U16611 ( .IN1(n16348), .IN2(n16349), .Q(n16347) );
  AND2X1 U16612 ( .IN1(n16350), .IN2(n16351), .Q(n16349) );
  OR2X1 U16613 ( .IN1(n11470), .IN2(g1346), .Q(n16351) );
  INVX0 U16614 ( .INP(n11469), .ZN(n11470) );
  OR2X1 U16615 ( .IN1(n4401), .IN2(n11469), .Q(n16350) );
  OR2X1 U16616 ( .IN1(n16352), .IN2(n16353), .Q(n11469) );
  OR2X1 U16617 ( .IN1(n16354), .IN2(n16355), .Q(n16353) );
  AND2X1 U16618 ( .IN1(n9985), .IN2(g6979), .Q(n16355) );
  AND2X1 U16619 ( .IN1(n10034), .IN2(g1315), .Q(n16354) );
  AND2X1 U16620 ( .IN1(n9984), .IN2(g7161), .Q(n16352) );
  AND2X1 U16621 ( .IN1(n16356), .IN2(n16357), .Q(n16348) );
  AND2X1 U16622 ( .IN1(n16358), .IN2(n16359), .Q(n16357) );
  OR2X1 U16623 ( .IN1(n11547), .IN2(g1372), .Q(n16359) );
  INVX0 U16624 ( .INP(n11545), .ZN(n11547) );
  OR2X1 U16625 ( .IN1(n4395), .IN2(n11545), .Q(n16358) );
  OR2X1 U16626 ( .IN1(n16360), .IN2(n16361), .Q(n11545) );
  OR2X1 U16627 ( .IN1(n16362), .IN2(n16363), .Q(n16361) );
  AND2X1 U16628 ( .IN1(n9978), .IN2(g6979), .Q(n16363) );
  AND2X1 U16629 ( .IN1(n10030), .IN2(g1315), .Q(n16362) );
  AND2X1 U16630 ( .IN1(n9977), .IN2(g7161), .Q(n16360) );
  AND2X1 U16631 ( .IN1(n16364), .IN2(n16365), .Q(n16356) );
  OR2X1 U16632 ( .IN1(n11498), .IN2(g1358), .Q(n16365) );
  INVX0 U16633 ( .INP(n11499), .ZN(n11498) );
  OR2X1 U16634 ( .IN1(n4411), .IN2(n11499), .Q(n16364) );
  OR2X1 U16635 ( .IN1(n16366), .IN2(n16367), .Q(n11499) );
  OR2X1 U16636 ( .IN1(n16368), .IN2(n16369), .Q(n16367) );
  AND2X1 U16637 ( .IN1(n9983), .IN2(g6979), .Q(n16369) );
  AND2X1 U16638 ( .IN1(n10033), .IN2(g1315), .Q(n16368) );
  INVX0 U16639 ( .INP(n16370), .ZN(n16366) );
  OR2X1 U16640 ( .IN1(n4358), .IN2(test_so50), .Q(n16370) );
  AND2X1 U16641 ( .IN1(n16371), .IN2(n16372), .Q(n16346) );
  AND2X1 U16642 ( .IN1(n16373), .IN2(n16374), .Q(n16372) );
  OR2X1 U16643 ( .IN1(n11519), .IN2(g1326), .Q(n16374) );
  INVX0 U16644 ( .INP(n11518), .ZN(n11519) );
  OR2X1 U16645 ( .IN1(n4402), .IN2(n11518), .Q(n16373) );
  OR2X1 U16646 ( .IN1(n16375), .IN2(n16376), .Q(n11518) );
  OR2X1 U16647 ( .IN1(n16377), .IN2(n16378), .Q(n16376) );
  AND2X1 U16648 ( .IN1(g6979), .IN2(n10221), .Q(n16378) );
  AND2X1 U16649 ( .IN1(n10038), .IN2(g1315), .Q(n16377) );
  AND2X1 U16650 ( .IN1(n9992), .IN2(g7161), .Q(n16375) );
  AND2X1 U16651 ( .IN1(n16379), .IN2(n16380), .Q(n16371) );
  OR2X1 U16652 ( .IN1(n11505), .IN2(g1339), .Q(n16380) );
  INVX0 U16653 ( .INP(n11504), .ZN(n11505) );
  OR2X1 U16654 ( .IN1(n4421), .IN2(n11504), .Q(n16379) );
  OR2X1 U16655 ( .IN1(n16381), .IN2(n16382), .Q(n11504) );
  OR2X1 U16656 ( .IN1(n16383), .IN2(n16384), .Q(n16382) );
  AND2X1 U16657 ( .IN1(n9989), .IN2(g6979), .Q(n16384) );
  AND2X1 U16658 ( .IN1(n10036), .IN2(g1315), .Q(n16383) );
  AND2X1 U16659 ( .IN1(n9988), .IN2(g7161), .Q(n16381) );
  AND2X1 U16660 ( .IN1(n9752), .IN2(g6979), .Q(n16302) );
  OR2X1 U16661 ( .IN1(n16385), .IN2(n16386), .Q(g25262) );
  AND2X1 U16662 ( .IN1(n16387), .IN2(g736), .Q(n16386) );
  AND2X1 U16663 ( .IN1(n16388), .IN2(n16283), .Q(n16385) );
  OR2X1 U16664 ( .IN1(n16389), .IN2(n16390), .Q(g25260) );
  AND2X1 U16665 ( .IN1(n16391), .IN2(g735), .Q(n16390) );
  AND2X1 U16666 ( .IN1(n16392), .IN2(n16283), .Q(n16389) );
  INVX0 U16667 ( .INP(n16393), .ZN(n16283) );
  OR2X1 U16668 ( .IN1(n16394), .IN2(n16395), .Q(n16393) );
  OR2X1 U16669 ( .IN1(n16396), .IN2(n11647), .Q(n16395) );
  OR2X1 U16670 ( .IN1(n16397), .IN2(n16398), .Q(n11647) );
  OR2X1 U16671 ( .IN1(n16399), .IN2(n16400), .Q(n16398) );
  AND2X1 U16672 ( .IN1(n9753), .IN2(g6677), .Q(n16400) );
  AND2X1 U16673 ( .IN1(n9807), .IN2(g629), .Q(n16399) );
  AND2X1 U16674 ( .IN1(n9745), .IN2(g6911), .Q(n16397) );
  AND2X1 U16675 ( .IN1(n9746), .IN2(g6911), .Q(n16396) );
  OR2X1 U16676 ( .IN1(n16401), .IN2(n16402), .Q(n16394) );
  OR2X1 U16677 ( .IN1(n16403), .IN2(n16404), .Q(n16402) );
  AND2X1 U16678 ( .IN1(n9808), .IN2(g629), .Q(n16404) );
  AND2X1 U16679 ( .IN1(n16405), .IN2(n16406), .Q(n16403) );
  AND2X1 U16680 ( .IN1(n16407), .IN2(n16408), .Q(n16406) );
  AND2X1 U16681 ( .IN1(n16409), .IN2(n16410), .Q(n16408) );
  AND2X1 U16682 ( .IN1(n16411), .IN2(n16412), .Q(n16410) );
  OR2X1 U16683 ( .IN1(n11043), .IN2(g633), .Q(n16412) );
  INVX0 U16684 ( .INP(n11044), .ZN(n11043) );
  OR2X1 U16685 ( .IN1(n4478), .IN2(n11044), .Q(n16411) );
  OR2X1 U16686 ( .IN1(n16413), .IN2(n16414), .Q(n11044) );
  OR2X1 U16687 ( .IN1(n16415), .IN2(n16416), .Q(n16414) );
  AND2X1 U16688 ( .IN1(n10008), .IN2(g6677), .Q(n16416) );
  AND2X1 U16689 ( .IN1(n10007), .IN2(g6911), .Q(n16415) );
  AND2X1 U16690 ( .IN1(n10047), .IN2(g629), .Q(n16413) );
  AND2X1 U16691 ( .IN1(n16417), .IN2(n16418), .Q(n16409) );
  OR2X1 U16692 ( .IN1(n16419), .IN2(n16420), .Q(n16418) );
  AND2X1 U16693 ( .IN1(n11016), .IN2(n10193), .Q(n16420) );
  INVX0 U16694 ( .INP(n11015), .ZN(n11016) );
  AND2X1 U16695 ( .IN1(test_so28), .IN2(n11015), .Q(n16419) );
  OR2X1 U16696 ( .IN1(n16421), .IN2(n16422), .Q(n11015) );
  OR2X1 U16697 ( .IN1(n16423), .IN2(n16424), .Q(n16422) );
  AND2X1 U16698 ( .IN1(n9999), .IN2(g6677), .Q(n16424) );
  AND2X1 U16699 ( .IN1(n10042), .IN2(g629), .Q(n16423) );
  AND2X1 U16700 ( .IN1(n9998), .IN2(g6911), .Q(n16421) );
  AND2X1 U16701 ( .IN1(n16425), .IN2(n16426), .Q(n16417) );
  OR2X1 U16702 ( .IN1(n11035), .IN2(g640), .Q(n16426) );
  INVX0 U16703 ( .INP(n11034), .ZN(n11035) );
  OR2X1 U16704 ( .IN1(n4404), .IN2(n11034), .Q(n16425) );
  OR2X1 U16705 ( .IN1(n16427), .IN2(n16428), .Q(n11034) );
  OR2X1 U16706 ( .IN1(n16429), .IN2(n16430), .Q(n16428) );
  AND2X1 U16707 ( .IN1(n10010), .IN2(g6677), .Q(n16430) );
  AND2X1 U16708 ( .IN1(n10009), .IN2(g6911), .Q(n16429) );
  AND2X1 U16709 ( .IN1(n10048), .IN2(g629), .Q(n16427) );
  AND2X1 U16710 ( .IN1(n16431), .IN2(n16432), .Q(n16407) );
  AND2X1 U16711 ( .IN1(n16433), .IN2(n16434), .Q(n16432) );
  OR2X1 U16712 ( .IN1(n11002), .IN2(g660), .Q(n16434) );
  INVX0 U16713 ( .INP(n11001), .ZN(n11002) );
  OR2X1 U16714 ( .IN1(n4403), .IN2(n11001), .Q(n16433) );
  OR2X1 U16715 ( .IN1(n16435), .IN2(n16436), .Q(n11001) );
  OR2X1 U16716 ( .IN1(n16437), .IN2(n16438), .Q(n16436) );
  AND2X1 U16717 ( .IN1(n10044), .IN2(g629), .Q(n16438) );
  AND2X1 U16718 ( .IN1(n10002), .IN2(g6911), .Q(n16437) );
  INVX0 U16719 ( .INP(n16439), .ZN(n16435) );
  OR2X1 U16720 ( .IN1(n4309), .IN2(test_so29), .Q(n16439) );
  AND2X1 U16721 ( .IN1(n16440), .IN2(n16441), .Q(n16431) );
  OR2X1 U16722 ( .IN1(n11010), .IN2(g672), .Q(n16441) );
  INVX0 U16723 ( .INP(n11011), .ZN(n11010) );
  OR2X1 U16724 ( .IN1(n4413), .IN2(n11011), .Q(n16440) );
  OR2X1 U16725 ( .IN1(n16442), .IN2(n16443), .Q(n11011) );
  OR2X1 U16726 ( .IN1(n16444), .IN2(n16445), .Q(n16443) );
  AND2X1 U16727 ( .IN1(n10001), .IN2(g6677), .Q(n16445) );
  AND2X1 U16728 ( .IN1(n10000), .IN2(g6911), .Q(n16444) );
  AND2X1 U16729 ( .IN1(n10043), .IN2(g629), .Q(n16442) );
  AND2X1 U16730 ( .IN1(n16446), .IN2(n16447), .Q(n16405) );
  AND2X1 U16731 ( .IN1(n16448), .IN2(n16449), .Q(n16447) );
  AND2X1 U16732 ( .IN1(n16450), .IN2(n16451), .Q(n16449) );
  OR2X1 U16733 ( .IN1(n11029), .IN2(g679), .Q(n16451) );
  INVX0 U16734 ( .INP(n11030), .ZN(n11029) );
  OR2X1 U16735 ( .IN1(n4477), .IN2(n11030), .Q(n16450) );
  OR2X1 U16736 ( .IN1(n16452), .IN2(n16453), .Q(n11030) );
  OR2X1 U16737 ( .IN1(n16454), .IN2(n16455), .Q(n16453) );
  AND2X1 U16738 ( .IN1(n9997), .IN2(g6677), .Q(n16455) );
  AND2X1 U16739 ( .IN1(n10041), .IN2(g629), .Q(n16454) );
  AND2X1 U16740 ( .IN1(n9996), .IN2(g6911), .Q(n16452) );
  AND2X1 U16741 ( .IN1(n16456), .IN2(n16457), .Q(n16448) );
  AND2X1 U16742 ( .IN1(n16458), .IN2(n16459), .Q(n16457) );
  INVX0 U16743 ( .INP(n16460), .ZN(n16459) );
  AND2X1 U16744 ( .IN1(n10969), .IN2(n4418), .Q(n16460) );
  OR2X1 U16745 ( .IN1(n4418), .IN2(n10969), .Q(n16458) );
  OR2X1 U16746 ( .IN1(n16461), .IN2(n16462), .Q(n10969) );
  OR2X1 U16747 ( .IN1(n16463), .IN2(n16464), .Q(n16462) );
  AND2X1 U16748 ( .IN1(n9993), .IN2(g6677), .Q(n16464) );
  AND2X1 U16749 ( .IN1(n10039), .IN2(g629), .Q(n16463) );
  INVX0 U16750 ( .INP(n16465), .ZN(n16461) );
  OR2X1 U16751 ( .IN1(n4359), .IN2(test_so30), .Q(n16465) );
  AND2X1 U16752 ( .IN1(n16466), .IN2(n16467), .Q(n16456) );
  INVX0 U16753 ( .INP(n16468), .ZN(n16467) );
  AND2X1 U16754 ( .IN1(n10959), .IN2(n4396), .Q(n16468) );
  OR2X1 U16755 ( .IN1(n4396), .IN2(n10959), .Q(n16466) );
  OR2X1 U16756 ( .IN1(n16469), .IN2(n16470), .Q(n10959) );
  OR2X1 U16757 ( .IN1(n16471), .IN2(n16472), .Q(n16470) );
  AND2X1 U16758 ( .IN1(n9995), .IN2(g6677), .Q(n16472) );
  AND2X1 U16759 ( .IN1(n10040), .IN2(g629), .Q(n16471) );
  AND2X1 U16760 ( .IN1(n9994), .IN2(g6911), .Q(n16469) );
  AND2X1 U16761 ( .IN1(n16473), .IN2(n16474), .Q(n16446) );
  AND2X1 U16762 ( .IN1(n16475), .IN2(n16476), .Q(n16474) );
  OR2X1 U16763 ( .IN1(n10995), .IN2(g646), .Q(n16476) );
  INVX0 U16764 ( .INP(n10996), .ZN(n10995) );
  OR2X1 U16765 ( .IN1(n4414), .IN2(n10996), .Q(n16475) );
  OR2X1 U16766 ( .IN1(n16477), .IN2(n16478), .Q(n10996) );
  OR2X1 U16767 ( .IN1(n16479), .IN2(n16480), .Q(n16478) );
  AND2X1 U16768 ( .IN1(n10004), .IN2(g6677), .Q(n16480) );
  AND2X1 U16769 ( .IN1(n10003), .IN2(g6911), .Q(n16479) );
  AND2X1 U16770 ( .IN1(n10045), .IN2(g629), .Q(n16477) );
  AND2X1 U16771 ( .IN1(n16481), .IN2(n16482), .Q(n16473) );
  OR2X1 U16772 ( .IN1(n11059), .IN2(g653), .Q(n16482) );
  INVX0 U16773 ( .INP(n11057), .ZN(n11059) );
  OR2X1 U16774 ( .IN1(n4422), .IN2(n11057), .Q(n16481) );
  OR2X1 U16775 ( .IN1(n16483), .IN2(n16484), .Q(n11057) );
  OR2X1 U16776 ( .IN1(n16485), .IN2(n16486), .Q(n16484) );
  AND2X1 U16777 ( .IN1(n10006), .IN2(g6677), .Q(n16486) );
  AND2X1 U16778 ( .IN1(n10005), .IN2(g6911), .Q(n16485) );
  AND2X1 U16779 ( .IN1(n10046), .IN2(g629), .Q(n16483) );
  AND2X1 U16780 ( .IN1(n9754), .IN2(g6677), .Q(n16401) );
  OR2X1 U16781 ( .IN1(n16487), .IN2(n16488), .Q(g25259) );
  AND2X1 U16782 ( .IN1(n16489), .IN2(g2253), .Q(n16488) );
  AND2X1 U16783 ( .IN1(n16490), .IN2(n13687), .Q(n16487) );
  OR2X1 U16784 ( .IN1(n16491), .IN2(n16492), .Q(g25257) );
  AND2X1 U16785 ( .IN1(n41), .IN2(n13687), .Q(n16492) );
  AND2X1 U16786 ( .IN1(n16493), .IN2(g2255), .Q(n16491) );
  OR2X1 U16787 ( .IN1(n16494), .IN2(n16495), .Q(g25256) );
  AND2X1 U16788 ( .IN1(n16489), .IN2(g2250), .Q(n16495) );
  AND2X1 U16789 ( .IN1(n16490), .IN2(n4377), .Q(n16494) );
  OR2X1 U16790 ( .IN1(n16496), .IN2(n16497), .Q(g25255) );
  AND2X1 U16791 ( .IN1(n16498), .IN2(g1559), .Q(n16497) );
  AND2X1 U16792 ( .IN1(n16499), .IN2(n13731), .Q(n16496) );
  OR2X1 U16793 ( .IN1(n16500), .IN2(n16501), .Q(g25253) );
  AND2X1 U16794 ( .IN1(n16502), .IN2(g2254), .Q(n16501) );
  AND2X1 U16795 ( .IN1(n16503), .IN2(n13687), .Q(n16500) );
  OR2X1 U16796 ( .IN1(n16504), .IN2(n16505), .Q(n13687) );
  OR2X1 U16797 ( .IN1(n16506), .IN2(n16507), .Q(n16505) );
  OR2X1 U16798 ( .IN1(n4319), .IN2(n4287), .Q(n16507) );
  OR2X1 U16799 ( .IN1(n4373), .IN2(n4325), .Q(n16506) );
  OR2X1 U16800 ( .IN1(n16508), .IN2(n16509), .Q(n16504) );
  OR2X1 U16801 ( .IN1(n4389), .IN2(n4377), .Q(n16509) );
  OR2X1 U16802 ( .IN1(n4563), .IN2(n4555), .Q(n16508) );
  OR2X1 U16803 ( .IN1(n16510), .IN2(n16511), .Q(g25252) );
  AND2X1 U16804 ( .IN1(n16493), .IN2(g2252), .Q(n16511) );
  AND2X1 U16805 ( .IN1(n41), .IN2(n4377), .Q(n16510) );
  OR2X1 U16806 ( .IN1(n16512), .IN2(n16513), .Q(g25251) );
  AND2X1 U16807 ( .IN1(n16489), .IN2(g2247), .Q(n16513) );
  AND2X1 U16808 ( .IN1(n16490), .IN2(n4373), .Q(n16512) );
  OR2X1 U16809 ( .IN1(n16514), .IN2(n16515), .Q(g25250) );
  AND2X1 U16810 ( .IN1(n16516), .IN2(g1561), .Q(n16515) );
  AND2X1 U16811 ( .IN1(n16517), .IN2(n13731), .Q(n16514) );
  OR2X1 U16812 ( .IN1(n16518), .IN2(n16519), .Q(g25249) );
  AND2X1 U16813 ( .IN1(n16498), .IN2(g1556), .Q(n16519) );
  AND2X1 U16814 ( .IN1(n16499), .IN2(n4378), .Q(n16518) );
  OR2X1 U16815 ( .IN1(n16520), .IN2(n16521), .Q(g25248) );
  AND2X1 U16816 ( .IN1(n16522), .IN2(g865), .Q(n16521) );
  AND2X1 U16817 ( .IN1(n16523), .IN2(n13770), .Q(n16520) );
  OR2X1 U16818 ( .IN1(n16524), .IN2(n16525), .Q(g25247) );
  AND2X1 U16819 ( .IN1(n16502), .IN2(g2251), .Q(n16525) );
  AND2X1 U16820 ( .IN1(n16503), .IN2(n4377), .Q(n16524) );
  OR2X1 U16821 ( .IN1(n16526), .IN2(n16527), .Q(g25246) );
  AND2X1 U16822 ( .IN1(n16493), .IN2(g2249), .Q(n16527) );
  AND2X1 U16823 ( .IN1(n41), .IN2(n4373), .Q(n16526) );
  OR2X1 U16824 ( .IN1(n16528), .IN2(n16529), .Q(g25245) );
  AND2X1 U16825 ( .IN1(n16530), .IN2(n16490), .Q(n16529) );
  INVX0 U16826 ( .INP(n16489), .ZN(n16490) );
  AND2X1 U16827 ( .IN1(n16489), .IN2(g2244), .Q(n16528) );
  OR2X1 U16828 ( .IN1(n4367), .IN2(n11558), .Q(n16489) );
  OR2X1 U16829 ( .IN1(n16531), .IN2(n16532), .Q(g25244) );
  AND2X1 U16830 ( .IN1(n16533), .IN2(g1560), .Q(n16532) );
  AND2X1 U16831 ( .IN1(n16534), .IN2(n13731), .Q(n16531) );
  OR2X1 U16832 ( .IN1(n16535), .IN2(n16536), .Q(n13731) );
  OR2X1 U16833 ( .IN1(n16537), .IN2(n16538), .Q(n16536) );
  OR2X1 U16834 ( .IN1(n4320), .IN2(n4288), .Q(n16538) );
  OR2X1 U16835 ( .IN1(n4374), .IN2(n4326), .Q(n16537) );
  OR2X1 U16836 ( .IN1(n16539), .IN2(n16540), .Q(n16535) );
  OR2X1 U16837 ( .IN1(n4390), .IN2(n4378), .Q(n16540) );
  OR2X1 U16838 ( .IN1(n4565), .IN2(n4557), .Q(n16539) );
  OR2X1 U16839 ( .IN1(n16541), .IN2(n16542), .Q(g25243) );
  AND2X1 U16840 ( .IN1(n16516), .IN2(g1558), .Q(n16542) );
  AND2X1 U16841 ( .IN1(n16517), .IN2(n4378), .Q(n16541) );
  OR2X1 U16842 ( .IN1(n16543), .IN2(n16544), .Q(g25242) );
  AND2X1 U16843 ( .IN1(n16499), .IN2(n4374), .Q(n16544) );
  AND2X1 U16844 ( .IN1(test_so54), .IN2(n16498), .Q(n16543) );
  OR2X1 U16845 ( .IN1(n16545), .IN2(n16546), .Q(g25241) );
  AND2X1 U16846 ( .IN1(n16547), .IN2(g867), .Q(n16546) );
  AND2X1 U16847 ( .IN1(n16548), .IN2(n13770), .Q(n16545) );
  OR2X1 U16848 ( .IN1(n16549), .IN2(n16550), .Q(g25240) );
  AND2X1 U16849 ( .IN1(n16522), .IN2(g862), .Q(n16550) );
  AND2X1 U16850 ( .IN1(n16523), .IN2(n4379), .Q(n16549) );
  OR2X1 U16851 ( .IN1(n16551), .IN2(n16552), .Q(g25239) );
  AND2X1 U16852 ( .IN1(n16553), .IN2(g177), .Q(n16552) );
  AND2X1 U16853 ( .IN1(n16554), .IN2(n13801), .Q(n16551) );
  OR2X1 U16854 ( .IN1(n16555), .IN2(n16556), .Q(g25237) );
  AND2X1 U16855 ( .IN1(n16502), .IN2(g2248), .Q(n16556) );
  AND2X1 U16856 ( .IN1(n16503), .IN2(n4373), .Q(n16555) );
  OR2X1 U16857 ( .IN1(n16557), .IN2(n16558), .Q(g25236) );
  AND2X1 U16858 ( .IN1(n16530), .IN2(n41), .Q(n16558) );
  INVX0 U16859 ( .INP(n16493), .ZN(n41) );
  AND2X1 U16860 ( .IN1(n16493), .IN2(g2246), .Q(n16557) );
  OR2X1 U16861 ( .IN1(n10189), .IN2(n11558), .Q(n16493) );
  OR2X1 U16862 ( .IN1(n16559), .IN2(n16560), .Q(g25235) );
  AND2X1 U16863 ( .IN1(n16533), .IN2(g1557), .Q(n16560) );
  AND2X1 U16864 ( .IN1(n16534), .IN2(n4378), .Q(n16559) );
  OR2X1 U16865 ( .IN1(n16561), .IN2(n16562), .Q(g25234) );
  AND2X1 U16866 ( .IN1(n16516), .IN2(g1555), .Q(n16562) );
  AND2X1 U16867 ( .IN1(n16517), .IN2(n4374), .Q(n16561) );
  OR2X1 U16868 ( .IN1(n16563), .IN2(n16564), .Q(g25233) );
  AND2X1 U16869 ( .IN1(n16565), .IN2(n16499), .Q(n16564) );
  INVX0 U16870 ( .INP(n16498), .ZN(n16499) );
  AND2X1 U16871 ( .IN1(n16498), .IN2(g1550), .Q(n16563) );
  OR2X1 U16872 ( .IN1(n4368), .IN2(n11558), .Q(n16498) );
  OR2X1 U16873 ( .IN1(n16566), .IN2(n16567), .Q(g25232) );
  AND2X1 U16874 ( .IN1(n16568), .IN2(g866), .Q(n16567) );
  AND2X1 U16875 ( .IN1(n16569), .IN2(n13770), .Q(n16566) );
  OR2X1 U16876 ( .IN1(n16570), .IN2(n16571), .Q(n13770) );
  OR2X1 U16877 ( .IN1(n16572), .IN2(n16573), .Q(n16571) );
  OR2X1 U16878 ( .IN1(n4321), .IN2(n4289), .Q(n16573) );
  OR2X1 U16879 ( .IN1(n4375), .IN2(n4327), .Q(n16572) );
  OR2X1 U16880 ( .IN1(n16574), .IN2(n16575), .Q(n16570) );
  OR2X1 U16881 ( .IN1(n4391), .IN2(n4379), .Q(n16575) );
  OR2X1 U16882 ( .IN1(n4567), .IN2(n4559), .Q(n16574) );
  OR2X1 U16883 ( .IN1(n16576), .IN2(n16577), .Q(g25231) );
  AND2X1 U16884 ( .IN1(n16547), .IN2(g864), .Q(n16577) );
  AND2X1 U16885 ( .IN1(n16548), .IN2(n4379), .Q(n16576) );
  OR2X1 U16886 ( .IN1(n16578), .IN2(n16579), .Q(g25230) );
  AND2X1 U16887 ( .IN1(n16522), .IN2(g859), .Q(n16579) );
  AND2X1 U16888 ( .IN1(n16523), .IN2(n4375), .Q(n16578) );
  OR2X1 U16889 ( .IN1(n16580), .IN2(n16581), .Q(g25229) );
  AND2X1 U16890 ( .IN1(n16582), .IN2(g179), .Q(n16581) );
  AND2X1 U16891 ( .IN1(n16583), .IN2(n13801), .Q(n16580) );
  OR2X1 U16892 ( .IN1(n16584), .IN2(n16585), .Q(g25228) );
  AND2X1 U16893 ( .IN1(n16553), .IN2(g174), .Q(n16585) );
  AND2X1 U16894 ( .IN1(n16554), .IN2(n4380), .Q(n16584) );
  OR2X1 U16895 ( .IN1(n16586), .IN2(n16587), .Q(g25227) );
  AND2X1 U16896 ( .IN1(n16530), .IN2(n16503), .Q(n16587) );
  INVX0 U16897 ( .INP(n16502), .ZN(n16503) );
  INVX0 U16898 ( .INP(n16588), .ZN(n16530) );
  OR2X1 U16899 ( .IN1(n16589), .IN2(n16590), .Q(n16588) );
  OR2X1 U16900 ( .IN1(g2190), .IN2(g2195), .Q(n16590) );
  OR2X1 U16901 ( .IN1(n4325), .IN2(n4287), .Q(n16589) );
  AND2X1 U16902 ( .IN1(n16502), .IN2(g2245), .Q(n16586) );
  OR2X1 U16903 ( .IN1(n4324), .IN2(n11558), .Q(n16502) );
  OR2X1 U16904 ( .IN1(n16591), .IN2(n16592), .Q(g25225) );
  AND2X1 U16905 ( .IN1(n16533), .IN2(g1554), .Q(n16592) );
  AND2X1 U16906 ( .IN1(n16534), .IN2(n4374), .Q(n16591) );
  OR2X1 U16907 ( .IN1(n16593), .IN2(n16594), .Q(g25224) );
  AND2X1 U16908 ( .IN1(n16565), .IN2(n16517), .Q(n16594) );
  INVX0 U16909 ( .INP(n16516), .ZN(n16517) );
  AND2X1 U16910 ( .IN1(n16516), .IN2(g1552), .Q(n16593) );
  OR2X1 U16911 ( .IN1(n4515), .IN2(n11558), .Q(n16516) );
  OR2X1 U16912 ( .IN1(n16595), .IN2(n16596), .Q(g25223) );
  AND2X1 U16913 ( .IN1(n16568), .IN2(g863), .Q(n16596) );
  AND2X1 U16914 ( .IN1(n16569), .IN2(n4379), .Q(n16595) );
  OR2X1 U16915 ( .IN1(n16597), .IN2(n16598), .Q(g25222) );
  AND2X1 U16916 ( .IN1(n16547), .IN2(g861), .Q(n16598) );
  AND2X1 U16917 ( .IN1(n16548), .IN2(n4375), .Q(n16597) );
  OR2X1 U16918 ( .IN1(n16599), .IN2(n16600), .Q(g25221) );
  AND2X1 U16919 ( .IN1(n16601), .IN2(n16523), .Q(n16600) );
  INVX0 U16920 ( .INP(n16522), .ZN(n16523) );
  AND2X1 U16921 ( .IN1(n16522), .IN2(g856), .Q(n16599) );
  OR2X1 U16922 ( .IN1(n10188), .IN2(n11558), .Q(n16522) );
  OR2X1 U16923 ( .IN1(n16602), .IN2(n16603), .Q(g25220) );
  AND2X1 U16924 ( .IN1(n16604), .IN2(g178), .Q(n16603) );
  AND2X1 U16925 ( .IN1(n16605), .IN2(n13801), .Q(n16602) );
  OR2X1 U16926 ( .IN1(n16606), .IN2(n16607), .Q(n13801) );
  OR2X1 U16927 ( .IN1(n16608), .IN2(n16609), .Q(n16607) );
  OR2X1 U16928 ( .IN1(n4322), .IN2(n4290), .Q(n16609) );
  OR2X1 U16929 ( .IN1(n4376), .IN2(n4328), .Q(n16608) );
  OR2X1 U16930 ( .IN1(n16610), .IN2(n16611), .Q(n16606) );
  OR2X1 U16931 ( .IN1(n4392), .IN2(n4380), .Q(n16611) );
  OR2X1 U16932 ( .IN1(n4569), .IN2(n4561), .Q(n16610) );
  OR2X1 U16933 ( .IN1(n16612), .IN2(n16613), .Q(g25219) );
  AND2X1 U16934 ( .IN1(n16582), .IN2(g176), .Q(n16613) );
  AND2X1 U16935 ( .IN1(n16583), .IN2(n4380), .Q(n16612) );
  OR2X1 U16936 ( .IN1(n16614), .IN2(n16615), .Q(g25218) );
  AND2X1 U16937 ( .IN1(n16553), .IN2(g171), .Q(n16615) );
  AND2X1 U16938 ( .IN1(n16554), .IN2(n4376), .Q(n16614) );
  OR2X1 U16939 ( .IN1(n16616), .IN2(n16617), .Q(g25217) );
  AND2X1 U16940 ( .IN1(n16565), .IN2(n16534), .Q(n16617) );
  INVX0 U16941 ( .INP(n16533), .ZN(n16534) );
  INVX0 U16942 ( .INP(n16618), .ZN(n16565) );
  OR2X1 U16943 ( .IN1(n16619), .IN2(n16620), .Q(n16618) );
  OR2X1 U16944 ( .IN1(g1496), .IN2(g1501), .Q(n16620) );
  OR2X1 U16945 ( .IN1(n4326), .IN2(n4288), .Q(n16619) );
  AND2X1 U16946 ( .IN1(n16533), .IN2(g1551), .Q(n16616) );
  OR2X1 U16947 ( .IN1(n4317), .IN2(n11558), .Q(n16533) );
  OR2X1 U16948 ( .IN1(n16621), .IN2(n16622), .Q(g25215) );
  AND2X1 U16949 ( .IN1(n16568), .IN2(g860), .Q(n16622) );
  AND2X1 U16950 ( .IN1(n16569), .IN2(n4375), .Q(n16621) );
  OR2X1 U16951 ( .IN1(n16623), .IN2(n16624), .Q(g25214) );
  AND2X1 U16952 ( .IN1(n16601), .IN2(n16548), .Q(n16624) );
  INVX0 U16953 ( .INP(n16547), .ZN(n16548) );
  AND2X1 U16954 ( .IN1(test_so33), .IN2(n16547), .Q(n16623) );
  OR2X1 U16955 ( .IN1(n4312), .IN2(n11558), .Q(n16547) );
  OR2X1 U16956 ( .IN1(n16625), .IN2(n16626), .Q(g25213) );
  AND2X1 U16957 ( .IN1(n16604), .IN2(g175), .Q(n16626) );
  AND2X1 U16958 ( .IN1(n16605), .IN2(n4380), .Q(n16625) );
  OR2X1 U16959 ( .IN1(n16627), .IN2(n16628), .Q(g25212) );
  AND2X1 U16960 ( .IN1(n16582), .IN2(g173), .Q(n16628) );
  AND2X1 U16961 ( .IN1(n16583), .IN2(n4376), .Q(n16627) );
  OR2X1 U16962 ( .IN1(n16629), .IN2(n16630), .Q(g25211) );
  AND2X1 U16963 ( .IN1(n16631), .IN2(n16554), .Q(n16630) );
  INVX0 U16964 ( .INP(n16553), .ZN(n16554) );
  AND2X1 U16965 ( .IN1(n16553), .IN2(g168), .Q(n16629) );
  OR2X1 U16966 ( .IN1(n4369), .IN2(n11558), .Q(n16553) );
  OR2X1 U16967 ( .IN1(n16632), .IN2(n16633), .Q(g25209) );
  AND2X1 U16968 ( .IN1(n16601), .IN2(n16569), .Q(n16633) );
  INVX0 U16969 ( .INP(n16568), .ZN(n16569) );
  INVX0 U16970 ( .INP(n16634), .ZN(n16601) );
  OR2X1 U16971 ( .IN1(n16635), .IN2(n16636), .Q(n16634) );
  OR2X1 U16972 ( .IN1(g805), .IN2(g809), .Q(n16636) );
  OR2X1 U16973 ( .IN1(n4327), .IN2(n4289), .Q(n16635) );
  AND2X1 U16974 ( .IN1(n16568), .IN2(g857), .Q(n16632) );
  OR2X1 U16975 ( .IN1(n4323), .IN2(n11558), .Q(n16568) );
  OR2X1 U16976 ( .IN1(n16637), .IN2(n16638), .Q(g25207) );
  AND2X1 U16977 ( .IN1(n16604), .IN2(g172), .Q(n16638) );
  AND2X1 U16978 ( .IN1(n16605), .IN2(n4376), .Q(n16637) );
  OR2X1 U16979 ( .IN1(n16639), .IN2(n16640), .Q(g25206) );
  AND2X1 U16980 ( .IN1(n16631), .IN2(n16583), .Q(n16640) );
  INVX0 U16981 ( .INP(n16582), .ZN(n16583) );
  AND2X1 U16982 ( .IN1(n16582), .IN2(g170), .Q(n16639) );
  OR2X1 U16983 ( .IN1(n4512), .IN2(n11558), .Q(n16582) );
  OR2X1 U16984 ( .IN1(n16641), .IN2(n16642), .Q(g25204) );
  AND2X1 U16985 ( .IN1(n16631), .IN2(n16605), .Q(n16642) );
  INVX0 U16986 ( .INP(n16604), .ZN(n16605) );
  INVX0 U16987 ( .INP(n16643), .ZN(n16631) );
  OR2X1 U16988 ( .IN1(n16644), .IN2(n16645), .Q(n16643) );
  OR2X1 U16989 ( .IN1(g117), .IN2(g121), .Q(n16645) );
  OR2X1 U16990 ( .IN1(n4328), .IN2(n4290), .Q(n16644) );
  AND2X1 U16991 ( .IN1(n16604), .IN2(g169), .Q(n16641) );
  OR2X1 U16992 ( .IN1(n4318), .IN2(n11558), .Q(n16604) );
  OR2X1 U16993 ( .IN1(n16646), .IN2(n16647), .Q(n11558) );
  OR2X1 U16994 ( .IN1(g2920), .IN2(n16648), .Q(n16647) );
  OR2X1 U16995 ( .IN1(n16649), .IN2(g2888), .Q(n16648) );
  OR2X1 U16996 ( .IN1(n16650), .IN2(n16651), .Q(n16646) );
  OR2X1 U16997 ( .IN1(g2912), .IN2(g2917), .Q(n16651) );
  OR2X1 U16998 ( .IN1(n4349), .IN2(n4330), .Q(n16650) );
  AND2X1 U16999 ( .IN1(n16652), .IN2(n10931), .Q(g25202) );
  AND2X1 U17000 ( .IN1(n16653), .IN2(n16654), .Q(n16652) );
  INVX0 U17001 ( .INP(n16655), .ZN(n16654) );
  AND2X1 U17002 ( .IN1(n16656), .IN2(n10157), .Q(n16655) );
  OR2X1 U17003 ( .IN1(n10157), .IN2(n16656), .Q(n16653) );
  AND2X1 U17004 ( .IN1(n16657), .IN2(n11730), .Q(g25201) );
  AND2X1 U17005 ( .IN1(n15919), .IN2(n16658), .Q(n16657) );
  INVX0 U17006 ( .INP(n4057), .ZN(n16658) );
  OR2X1 U17007 ( .IN1(n4305), .IN2(n4058), .Q(n15919) );
  AND2X1 U17008 ( .IN1(n16659), .IN2(n10874), .Q(g25199) );
  AND2X1 U17009 ( .IN1(n16660), .IN2(n16661), .Q(n16659) );
  OR2X1 U17010 ( .IN1(n16662), .IN2(g2920), .Q(n16661) );
  INVX0 U17011 ( .INP(n16663), .ZN(n16662) );
  OR2X1 U17012 ( .IN1(n9892), .IN2(n16663), .Q(n16660) );
  AND2X1 U17013 ( .IN1(n16664), .IN2(n14331), .Q(g25197) );
  AND2X1 U17014 ( .IN1(n16665), .IN2(n16666), .Q(n16664) );
  OR2X1 U17015 ( .IN1(n15367), .IN2(g2734), .Q(n16666) );
  INVX0 U17016 ( .INP(n15368), .ZN(n15367) );
  OR2X1 U17017 ( .IN1(n4397), .IN2(n15368), .Q(n16665) );
  AND2X1 U17018 ( .IN1(n16667), .IN2(n14337), .Q(g25194) );
  AND2X1 U17019 ( .IN1(n16668), .IN2(n16669), .Q(n16667) );
  OR2X1 U17020 ( .IN1(n15386), .IN2(g2040), .Q(n16669) );
  INVX0 U17021 ( .INP(n15387), .ZN(n15386) );
  OR2X1 U17022 ( .IN1(n4399), .IN2(n15387), .Q(n16668) );
  AND2X1 U17023 ( .IN1(n16670), .IN2(n15352), .Q(g25191) );
  AND2X1 U17024 ( .IN1(n16671), .IN2(n1808), .Q(n16670) );
  INVX0 U17025 ( .INP(n15924), .ZN(n1808) );
  AND2X1 U17026 ( .IN1(g3013), .IN2(n4065), .Q(n15924) );
  OR2X1 U17027 ( .IN1(n4065), .IN2(g3013), .Q(n16671) );
  AND2X1 U17028 ( .IN1(n16672), .IN2(n14345), .Q(g25189) );
  AND2X1 U17029 ( .IN1(n16673), .IN2(n16674), .Q(n16672) );
  OR2X1 U17030 ( .IN1(n15507), .IN2(g1346), .Q(n16674) );
  INVX0 U17031 ( .INP(n15508), .ZN(n15507) );
  OR2X1 U17032 ( .IN1(n4401), .IN2(n15508), .Q(n16673) );
  AND2X1 U17033 ( .IN1(n16675), .IN2(n13809), .Q(g25185) );
  AND2X1 U17034 ( .IN1(n16676), .IN2(n16677), .Q(n16675) );
  OR2X1 U17035 ( .IN1(n15628), .IN2(g660), .Q(n16677) );
  INVX0 U17036 ( .INP(n15629), .ZN(n15628) );
  OR2X1 U17037 ( .IN1(n4403), .IN2(n15629), .Q(n16676) );
  AND2X1 U17038 ( .IN1(n16678), .IN2(n12966), .Q(g25067) );
  OR2X1 U17039 ( .IN1(n16649), .IN2(n16679), .Q(n12966) );
  AND2X1 U17040 ( .IN1(n16680), .IN2(n16681), .Q(n16678) );
  OR2X1 U17041 ( .IN1(n16682), .IN2(g2160), .Q(n16681) );
  INVX0 U17042 ( .INP(n3888), .ZN(n16682) );
  OR2X1 U17043 ( .IN1(n9879), .IN2(n3888), .Q(n16680) );
  OR2X1 U17044 ( .IN1(n10672), .IN2(n4367), .Q(n3888) );
  AND2X1 U17045 ( .IN1(n16683), .IN2(n12971), .Q(g25056) );
  OR2X1 U17046 ( .IN1(n16649), .IN2(n16684), .Q(n12971) );
  AND2X1 U17047 ( .IN1(n16685), .IN2(n16686), .Q(n16683) );
  OR2X1 U17048 ( .IN1(n16687), .IN2(g1466), .Q(n16686) );
  INVX0 U17049 ( .INP(n3891), .ZN(n16687) );
  OR2X1 U17050 ( .IN1(n9883), .IN2(n3891), .Q(n16685) );
  OR2X1 U17051 ( .IN1(n10672), .IN2(n4368), .Q(n3891) );
  AND2X1 U17052 ( .IN1(n16688), .IN2(n12976), .Q(g25042) );
  OR2X1 U17053 ( .IN1(n16649), .IN2(n16689), .Q(n12976) );
  AND2X1 U17054 ( .IN1(n16690), .IN2(n16691), .Q(n16688) );
  OR2X1 U17055 ( .IN1(n16692), .IN2(g780), .Q(n16691) );
  INVX0 U17056 ( .INP(n3894), .ZN(n16692) );
  OR2X1 U17057 ( .IN1(n9887), .IN2(n3894), .Q(n16690) );
  OR2X1 U17058 ( .IN1(n10672), .IN2(n10188), .Q(n3894) );
  AND2X1 U17059 ( .IN1(n16693), .IN2(n12981), .Q(g25027) );
  OR2X1 U17060 ( .IN1(n16649), .IN2(n16694), .Q(n12981) );
  INVX0 U17061 ( .INP(n10672), .ZN(n16649) );
  AND2X1 U17062 ( .IN1(n16695), .IN2(n16696), .Q(n16693) );
  OR2X1 U17063 ( .IN1(n16697), .IN2(g92), .Q(n16696) );
  INVX0 U17064 ( .INP(n3897), .ZN(n16697) );
  OR2X1 U17065 ( .IN1(n9891), .IN2(n3897), .Q(n16695) );
  OR2X1 U17066 ( .IN1(n10672), .IN2(n4369), .Q(n3897) );
  AND2X1 U17067 ( .IN1(n16698), .IN2(n16699), .Q(n10672) );
  AND2X1 U17068 ( .IN1(n4355), .IN2(n4431), .Q(n16699) );
  AND2X1 U17069 ( .IN1(n4305), .IN2(n16700), .Q(n16698) );
  AND2X1 U17070 ( .IN1(n10173), .IN2(n4291), .Q(n16700) );
  OR2X1 U17071 ( .IN1(n16701), .IN2(n14497), .Q(g24734) );
  INVX0 U17072 ( .INP(n3700), .ZN(n14497) );
  AND2X1 U17073 ( .IN1(n14501), .IN2(DFF_146_n1), .Q(n16701) );
  AND2X1 U17074 ( .IN1(n3705), .IN2(n3940), .Q(n14501) );
  OR2X1 U17075 ( .IN1(n16702), .IN2(n16703), .Q(g24557) );
  AND2X1 U17076 ( .IN1(n4299), .IN2(g2676), .Q(n16703) );
  AND2X1 U17077 ( .IN1(n16704), .IN2(n11557), .Q(n16702) );
  OR2X1 U17078 ( .IN1(n16705), .IN2(n16706), .Q(g24548) );
  AND2X1 U17079 ( .IN1(n16707), .IN2(g7390), .Q(n16706) );
  AND2X1 U17080 ( .IN1(n4370), .IN2(g2673), .Q(n16705) );
  OR2X1 U17081 ( .IN1(n16708), .IN2(n16709), .Q(g24547) );
  AND2X1 U17082 ( .IN1(n4299), .IN2(g2667), .Q(n16709) );
  AND2X1 U17083 ( .IN1(n16704), .IN2(n13925), .Q(n16708) );
  OR2X1 U17084 ( .IN1(n16710), .IN2(n16711), .Q(g24545) );
  AND2X1 U17085 ( .IN1(n4366), .IN2(g1982), .Q(n16711) );
  AND2X1 U17086 ( .IN1(n16712), .IN2(n13983), .Q(n16710) );
  OR2X1 U17087 ( .IN1(n16713), .IN2(n16714), .Q(g24538) );
  AND2X1 U17088 ( .IN1(n4314), .IN2(g2670), .Q(n16714) );
  AND2X1 U17089 ( .IN1(n16707), .IN2(g7302), .Q(n16713) );
  AND2X1 U17090 ( .IN1(n11557), .IN2(n13858), .Q(n16707) );
  OR2X1 U17091 ( .IN1(n16715), .IN2(n16716), .Q(n11557) );
  OR2X1 U17092 ( .IN1(n16717), .IN2(n16718), .Q(n16716) );
  AND2X1 U17093 ( .IN1(g7390), .IN2(g2673), .Q(n16718) );
  AND2X1 U17094 ( .IN1(n12862), .IN2(g2670), .Q(n16717) );
  OR2X1 U17095 ( .IN1(n16719), .IN2(n16720), .Q(n16715) );
  AND2X1 U17096 ( .IN1(g2624), .IN2(g2676), .Q(n16720) );
  AND2X1 U17097 ( .IN1(n16721), .IN2(test_so88), .Q(n16719) );
  AND2X1 U17098 ( .IN1(n11732), .IN2(g185), .Q(n16721) );
  OR2X1 U17099 ( .IN1(n16722), .IN2(n16723), .Q(n11732) );
  OR2X1 U17100 ( .IN1(n16724), .IN2(n16725), .Q(n16723) );
  AND2X1 U17101 ( .IN1(n12862), .IN2(g2639), .Q(n16725) );
  AND2X1 U17102 ( .IN1(g2624), .IN2(g2564), .Q(n16724) );
  AND2X1 U17103 ( .IN1(g7390), .IN2(g2641), .Q(n16722) );
  OR2X1 U17104 ( .IN1(n16726), .IN2(n16727), .Q(g24537) );
  AND2X1 U17105 ( .IN1(n16728), .IN2(g7390), .Q(n16727) );
  AND2X1 U17106 ( .IN1(n4370), .IN2(g2664), .Q(n16726) );
  OR2X1 U17107 ( .IN1(n16729), .IN2(n16730), .Q(g24535) );
  AND2X1 U17108 ( .IN1(n16731), .IN2(g7194), .Q(n16730) );
  AND2X1 U17109 ( .IN1(n4315), .IN2(g1979), .Q(n16729) );
  OR2X1 U17110 ( .IN1(n16732), .IN2(n16733), .Q(g24534) );
  AND2X1 U17111 ( .IN1(n4366), .IN2(g1973), .Q(n16733) );
  AND2X1 U17112 ( .IN1(n16712), .IN2(n14094), .Q(n16732) );
  OR2X1 U17113 ( .IN1(n16734), .IN2(n16735), .Q(g24532) );
  AND2X1 U17114 ( .IN1(n4300), .IN2(g1288), .Q(n16735) );
  AND2X1 U17115 ( .IN1(n16736), .IN2(n14106), .Q(n16734) );
  OR2X1 U17116 ( .IN1(n16737), .IN2(n16738), .Q(g24527) );
  AND2X1 U17117 ( .IN1(n16728), .IN2(n12862), .Q(n16738) );
  AND2X1 U17118 ( .IN1(n13925), .IN2(n13858), .Q(n16728) );
  OR2X1 U17119 ( .IN1(n16739), .IN2(n16740), .Q(n13925) );
  OR2X1 U17120 ( .IN1(n16741), .IN2(n16742), .Q(n16740) );
  AND2X1 U17121 ( .IN1(g7390), .IN2(g2664), .Q(n16742) );
  AND2X1 U17122 ( .IN1(g2624), .IN2(g2667), .Q(n16741) );
  OR2X1 U17123 ( .IN1(n16743), .IN2(n16744), .Q(n16739) );
  AND2X1 U17124 ( .IN1(g7302), .IN2(g2661), .Q(n16744) );
  AND2X1 U17125 ( .IN1(n16745), .IN2(n11731), .Q(n16743) );
  OR2X1 U17126 ( .IN1(n16746), .IN2(n16747), .Q(n11731) );
  OR2X1 U17127 ( .IN1(n16748), .IN2(n16749), .Q(n16747) );
  AND2X1 U17128 ( .IN1(g2624), .IN2(g2647), .Q(n16749) );
  AND2X1 U17129 ( .IN1(g7302), .IN2(g2643), .Q(n16748) );
  AND2X1 U17130 ( .IN1(g7390), .IN2(g2645), .Q(n16746) );
  AND2X1 U17131 ( .IN1(g185), .IN2(g2598), .Q(n16745) );
  AND2X1 U17132 ( .IN1(n4314), .IN2(g2661), .Q(n16737) );
  OR2X1 U17133 ( .IN1(n16750), .IN2(n16751), .Q(g24525) );
  AND2X1 U17134 ( .IN1(n4296), .IN2(g1976), .Q(n16751) );
  AND2X1 U17135 ( .IN1(n16731), .IN2(g7052), .Q(n16750) );
  AND2X1 U17136 ( .IN1(n13983), .IN2(n13858), .Q(n16731) );
  OR2X1 U17137 ( .IN1(n16752), .IN2(n16753), .Q(n13983) );
  OR2X1 U17138 ( .IN1(n16754), .IN2(n16755), .Q(n16753) );
  AND2X1 U17139 ( .IN1(g1930), .IN2(g1982), .Q(n16755) );
  AND2X1 U17140 ( .IN1(g7194), .IN2(g1979), .Q(n16754) );
  OR2X1 U17141 ( .IN1(n16756), .IN2(n16757), .Q(n16752) );
  AND2X1 U17142 ( .IN1(n13973), .IN2(g1976), .Q(n16757) );
  AND2X1 U17143 ( .IN1(n16758), .IN2(n11736), .Q(n16756) );
  OR2X1 U17144 ( .IN1(n16759), .IN2(n16760), .Q(n11736) );
  OR2X1 U17145 ( .IN1(n16761), .IN2(n16762), .Q(n16760) );
  AND2X1 U17146 ( .IN1(g7194), .IN2(g1947), .Q(n16762) );
  AND2X1 U17147 ( .IN1(n13973), .IN2(g1945), .Q(n16761) );
  AND2X1 U17148 ( .IN1(g1930), .IN2(g1870), .Q(n16759) );
  AND2X1 U17149 ( .IN1(g185), .IN2(g1922), .Q(n16758) );
  OR2X1 U17150 ( .IN1(n16763), .IN2(n16764), .Q(g24524) );
  AND2X1 U17151 ( .IN1(n16765), .IN2(g7194), .Q(n16764) );
  AND2X1 U17152 ( .IN1(n4315), .IN2(g1970), .Q(n16763) );
  OR2X1 U17153 ( .IN1(n16766), .IN2(n16767), .Q(g24522) );
  AND2X1 U17154 ( .IN1(n16768), .IN2(g6944), .Q(n16767) );
  AND2X1 U17155 ( .IN1(n4316), .IN2(g1285), .Q(n16766) );
  OR2X1 U17156 ( .IN1(n16769), .IN2(n16770), .Q(g24521) );
  AND2X1 U17157 ( .IN1(n4300), .IN2(g1279), .Q(n16770) );
  AND2X1 U17158 ( .IN1(n16736), .IN2(n14214), .Q(n16769) );
  OR2X1 U17159 ( .IN1(n16771), .IN2(n16772), .Q(g24519) );
  AND2X1 U17160 ( .IN1(n4313), .IN2(g602), .Q(n16772) );
  AND2X1 U17161 ( .IN1(n16773), .IN2(n14226), .Q(n16771) );
  OR2X1 U17162 ( .IN1(n16774), .IN2(n16775), .Q(g24513) );
  AND2X1 U17163 ( .IN1(n16765), .IN2(n13973), .Q(n16775) );
  AND2X1 U17164 ( .IN1(n14094), .IN2(n13858), .Q(n16765) );
  OR2X1 U17165 ( .IN1(n16776), .IN2(n16777), .Q(n14094) );
  OR2X1 U17166 ( .IN1(n16778), .IN2(n16779), .Q(n16777) );
  AND2X1 U17167 ( .IN1(g1930), .IN2(g1973), .Q(n16779) );
  AND2X1 U17168 ( .IN1(g7194), .IN2(g1970), .Q(n16778) );
  OR2X1 U17169 ( .IN1(n16780), .IN2(n16781), .Q(n16776) );
  AND2X1 U17170 ( .IN1(g7052), .IN2(g1967), .Q(n16781) );
  AND2X1 U17171 ( .IN1(n16782), .IN2(n11735), .Q(n16780) );
  OR2X1 U17172 ( .IN1(n16783), .IN2(n16784), .Q(n11735) );
  OR2X1 U17173 ( .IN1(n16785), .IN2(n16786), .Q(n16784) );
  AND2X1 U17174 ( .IN1(g7194), .IN2(g1951), .Q(n16786) );
  AND2X1 U17175 ( .IN1(g7052), .IN2(g1949), .Q(n16785) );
  AND2X1 U17176 ( .IN1(g1930), .IN2(g1953), .Q(n16783) );
  AND2X1 U17177 ( .IN1(g185), .IN2(g1904), .Q(n16782) );
  AND2X1 U17178 ( .IN1(n4296), .IN2(g1967), .Q(n16774) );
  OR2X1 U17179 ( .IN1(n16787), .IN2(n16788), .Q(g24511) );
  AND2X1 U17180 ( .IN1(n4371), .IN2(g1282), .Q(n16788) );
  AND2X1 U17181 ( .IN1(n16768), .IN2(g6750), .Q(n16787) );
  AND2X1 U17182 ( .IN1(n14106), .IN2(n13858), .Q(n16768) );
  OR2X1 U17183 ( .IN1(n16789), .IN2(n16790), .Q(n14106) );
  OR2X1 U17184 ( .IN1(n16791), .IN2(n16792), .Q(n16790) );
  AND2X1 U17185 ( .IN1(n13842), .IN2(g1282), .Q(n16792) );
  AND2X1 U17186 ( .IN1(g6944), .IN2(g1285), .Q(n16791) );
  OR2X1 U17187 ( .IN1(n16793), .IN2(n16794), .Q(n16789) );
  AND2X1 U17188 ( .IN1(g1236), .IN2(g1288), .Q(n16794) );
  AND2X1 U17189 ( .IN1(n16795), .IN2(test_so45), .Q(n16793) );
  AND2X1 U17190 ( .IN1(n10598), .IN2(g185), .Q(n16795) );
  OR2X1 U17191 ( .IN1(n16796), .IN2(n16797), .Q(n10598) );
  OR2X1 U17192 ( .IN1(n16798), .IN2(n16799), .Q(n16797) );
  AND2X1 U17193 ( .IN1(g1236), .IN2(g1176), .Q(n16799) );
  AND2X1 U17194 ( .IN1(g6750), .IN2(g1251), .Q(n16798) );
  AND2X1 U17195 ( .IN1(g6944), .IN2(g1253), .Q(n16796) );
  OR2X1 U17196 ( .IN1(n16800), .IN2(n16801), .Q(g24510) );
  AND2X1 U17197 ( .IN1(n16802), .IN2(g6944), .Q(n16801) );
  AND2X1 U17198 ( .IN1(n4316), .IN2(g1276), .Q(n16800) );
  OR2X1 U17199 ( .IN1(n16803), .IN2(n16804), .Q(g24508) );
  AND2X1 U17200 ( .IN1(n16805), .IN2(g6642), .Q(n16804) );
  AND2X1 U17201 ( .IN1(n4372), .IN2(g599), .Q(n16803) );
  OR2X1 U17202 ( .IN1(n16806), .IN2(n16807), .Q(g24507) );
  AND2X1 U17203 ( .IN1(n4313), .IN2(g593), .Q(n16807) );
  AND2X1 U17204 ( .IN1(n16773), .IN2(n14329), .Q(n16806) );
  OR2X1 U17205 ( .IN1(n16808), .IN2(n16809), .Q(g24501) );
  AND2X1 U17206 ( .IN1(n16802), .IN2(n13842), .Q(n16809) );
  AND2X1 U17207 ( .IN1(n14214), .IN2(n13858), .Q(n16802) );
  OR2X1 U17208 ( .IN1(n16810), .IN2(n16811), .Q(n14214) );
  OR2X1 U17209 ( .IN1(n16812), .IN2(n16813), .Q(n16811) );
  AND2X1 U17210 ( .IN1(g6944), .IN2(g1276), .Q(n16813) );
  AND2X1 U17211 ( .IN1(g1236), .IN2(g1279), .Q(n16812) );
  OR2X1 U17212 ( .IN1(n16814), .IN2(n16815), .Q(n16810) );
  AND2X1 U17213 ( .IN1(g6750), .IN2(g1273), .Q(n16815) );
  AND2X1 U17214 ( .IN1(n16816), .IN2(n10599), .Q(n16814) );
  OR2X1 U17215 ( .IN1(n16817), .IN2(n16818), .Q(n10599) );
  OR2X1 U17216 ( .IN1(n16819), .IN2(n16820), .Q(n16818) );
  AND2X1 U17217 ( .IN1(g6944), .IN2(g1257), .Q(n16820) );
  AND2X1 U17218 ( .IN1(g1236), .IN2(g1259), .Q(n16819) );
  AND2X1 U17219 ( .IN1(n13842), .IN2(g1255), .Q(n16817) );
  AND2X1 U17220 ( .IN1(g185), .IN2(g1210), .Q(n16816) );
  AND2X1 U17221 ( .IN1(n4371), .IN2(g1273), .Q(n16808) );
  OR2X1 U17222 ( .IN1(n16821), .IN2(n16822), .Q(g24499) );
  AND2X1 U17223 ( .IN1(n4298), .IN2(g596), .Q(n16822) );
  AND2X1 U17224 ( .IN1(n16805), .IN2(g6485), .Q(n16821) );
  AND2X1 U17225 ( .IN1(n14226), .IN2(n13858), .Q(n16805) );
  OR2X1 U17226 ( .IN1(n16823), .IN2(n16824), .Q(n14226) );
  OR2X1 U17227 ( .IN1(n16825), .IN2(n16826), .Q(n16824) );
  AND2X1 U17228 ( .IN1(g6642), .IN2(g599), .Q(n16826) );
  AND2X1 U17229 ( .IN1(g550), .IN2(g602), .Q(n16825) );
  OR2X1 U17230 ( .IN1(n16827), .IN2(n16828), .Q(n16823) );
  AND2X1 U17231 ( .IN1(g6485), .IN2(g596), .Q(n16828) );
  AND2X1 U17232 ( .IN1(n16829), .IN2(n10603), .Q(n16827) );
  OR2X1 U17233 ( .IN1(n16830), .IN2(n16831), .Q(n10603) );
  OR2X1 U17234 ( .IN1(n16832), .IN2(n16833), .Q(n16831) );
  AND2X1 U17235 ( .IN1(g550), .IN2(g489), .Q(n16833) );
  AND2X1 U17236 ( .IN1(n11054), .IN2(g565), .Q(n16832) );
  AND2X1 U17237 ( .IN1(g6642), .IN2(g567), .Q(n16830) );
  AND2X1 U17238 ( .IN1(g185), .IN2(g542), .Q(n16829) );
  OR2X1 U17239 ( .IN1(n16834), .IN2(n16835), .Q(g24498) );
  AND2X1 U17240 ( .IN1(n16836), .IN2(g6642), .Q(n16835) );
  AND2X1 U17241 ( .IN1(n4372), .IN2(g590), .Q(n16834) );
  OR2X1 U17242 ( .IN1(n16837), .IN2(n16838), .Q(g24491) );
  AND2X1 U17243 ( .IN1(n16836), .IN2(n11054), .Q(n16838) );
  AND2X1 U17244 ( .IN1(n14329), .IN2(n13858), .Q(n16836) );
  OR2X1 U17245 ( .IN1(n16839), .IN2(n16840), .Q(n14329) );
  OR2X1 U17246 ( .IN1(n16841), .IN2(n16842), .Q(n16840) );
  AND2X1 U17247 ( .IN1(g6642), .IN2(g590), .Q(n16842) );
  AND2X1 U17248 ( .IN1(g550), .IN2(g593), .Q(n16841) );
  OR2X1 U17249 ( .IN1(n16843), .IN2(n16844), .Q(n16839) );
  AND2X1 U17250 ( .IN1(n11054), .IN2(g587), .Q(n16844) );
  AND2X1 U17251 ( .IN1(n16845), .IN2(n10601), .Q(n16843) );
  OR2X1 U17252 ( .IN1(n16846), .IN2(n16847), .Q(n10601) );
  OR2X1 U17253 ( .IN1(n16848), .IN2(n16849), .Q(n16847) );
  AND2X1 U17254 ( .IN1(g550), .IN2(g573), .Q(n16849) );
  AND2X1 U17255 ( .IN1(g6485), .IN2(g569), .Q(n16848) );
  AND2X1 U17256 ( .IN1(g6642), .IN2(g571), .Q(n16846) );
  AND2X1 U17257 ( .IN1(g185), .IN2(g524), .Q(n16845) );
  AND2X1 U17258 ( .IN1(n4298), .IN2(g587), .Q(n16837) );
  AND2X1 U17259 ( .IN1(n16850), .IN2(n16851), .Q(g24476) );
  OR2X1 U17260 ( .IN1(n16852), .IN2(g2924), .Q(n16851) );
  AND2X1 U17261 ( .IN1(n10876), .IN2(g2917), .Q(n16852) );
  AND2X1 U17262 ( .IN1(n16663), .IN2(n10874), .Q(n16850) );
  OR2X1 U17263 ( .IN1(n16853), .IN2(n16854), .Q(n16663) );
  OR2X1 U17264 ( .IN1(n4479), .IN2(n4349), .Q(n16854) );
  AND2X1 U17265 ( .IN1(n16855), .IN2(n11730), .Q(g24473) );
  AND2X1 U17266 ( .IN1(n16856), .IN2(n4058), .Q(n16855) );
  OR2X1 U17267 ( .IN1(n10173), .IN2(n16857), .Q(n4058) );
  INVX0 U17268 ( .INP(n16858), .ZN(n16856) );
  AND2X1 U17269 ( .IN1(n16857), .IN2(n10173), .Q(n16858) );
  AND2X1 U17270 ( .IN1(n16859), .IN2(n16656), .Q(g24446) );
  OR2X1 U17271 ( .IN1(n4480), .IN2(n4102), .Q(n16656) );
  AND2X1 U17272 ( .IN1(n10931), .IN2(n16860), .Q(n16859) );
  INVX0 U17273 ( .INP(n4101), .ZN(n16860) );
  AND2X1 U17274 ( .IN1(n16861), .IN2(n15352), .Q(g24445) );
  AND2X1 U17275 ( .IN1(n16862), .IN2(n16863), .Q(n16861) );
  INVX0 U17276 ( .INP(n16864), .ZN(n16863) );
  AND2X1 U17277 ( .IN1(n4066), .IN2(n9352), .Q(n16864) );
  OR2X1 U17278 ( .IN1(n9352), .IN2(n4066), .Q(n16862) );
  AND2X1 U17279 ( .IN1(n16865), .IN2(n16866), .Q(g24438) );
  OR2X1 U17280 ( .IN1(n16867), .IN2(g2720), .Q(n16866) );
  AND2X1 U17281 ( .IN1(n16868), .IN2(g2727), .Q(n16867) );
  AND2X1 U17282 ( .IN1(n15368), .IN2(n14331), .Q(n16865) );
  OR2X1 U17283 ( .IN1(n16869), .IN2(n16870), .Q(n15368) );
  OR2X1 U17284 ( .IN1(n4419), .IN2(n4408), .Q(n16870) );
  AND2X1 U17285 ( .IN1(n16871), .IN2(n16872), .Q(g24434) );
  OR2X1 U17286 ( .IN1(n16873), .IN2(g2026), .Q(n16872) );
  AND2X1 U17287 ( .IN1(n16874), .IN2(g2033), .Q(n16873) );
  AND2X1 U17288 ( .IN1(n15387), .IN2(n14337), .Q(n16871) );
  OR2X1 U17289 ( .IN1(n16875), .IN2(n16876), .Q(n15387) );
  OR2X1 U17290 ( .IN1(n4420), .IN2(n4410), .Q(n16876) );
  AND2X1 U17291 ( .IN1(n16877), .IN2(n16878), .Q(g24430) );
  OR2X1 U17292 ( .IN1(n16879), .IN2(g1332), .Q(n16878) );
  AND2X1 U17293 ( .IN1(n16880), .IN2(g1339), .Q(n16879) );
  AND2X1 U17294 ( .IN1(n15508), .IN2(n14345), .Q(n16877) );
  OR2X1 U17295 ( .IN1(n16881), .IN2(n16882), .Q(n15508) );
  OR2X1 U17296 ( .IN1(n4421), .IN2(n4412), .Q(n16882) );
  AND2X1 U17297 ( .IN1(n16883), .IN2(n16884), .Q(g24426) );
  OR2X1 U17298 ( .IN1(n16885), .IN2(g646), .Q(n16884) );
  AND2X1 U17299 ( .IN1(n16886), .IN2(g653), .Q(n16885) );
  AND2X1 U17300 ( .IN1(n15629), .IN2(n13809), .Q(n16883) );
  OR2X1 U17301 ( .IN1(n16887), .IN2(n16888), .Q(n15629) );
  OR2X1 U17302 ( .IN1(n4422), .IN2(n4414), .Q(n16888) );
  OR2X1 U17303 ( .IN1(n16889), .IN2(n16890), .Q(g24250) );
  AND2X1 U17304 ( .IN1(n16891), .IN2(g2560), .Q(n16890) );
  AND2X1 U17305 ( .IN1(n4463), .IN2(g2546), .Q(n16889) );
  OR2X1 U17306 ( .IN1(n16892), .IN2(n16893), .Q(g24243) );
  AND2X1 U17307 ( .IN1(n16894), .IN2(g1866), .Q(n16893) );
  AND2X1 U17308 ( .IN1(n4464), .IN2(g1852), .Q(n16892) );
  OR2X1 U17309 ( .IN1(n16895), .IN2(n16896), .Q(g24238) );
  AND2X1 U17310 ( .IN1(n13236), .IN2(g2560), .Q(n16896) );
  AND2X1 U17311 ( .IN1(n4463), .IN2(g2554), .Q(n16895) );
  OR2X1 U17312 ( .IN1(n16897), .IN2(n16898), .Q(g24237) );
  AND2X1 U17313 ( .IN1(n16891), .IN2(g8167), .Q(n16898) );
  AND2X1 U17314 ( .IN1(n4455), .IN2(g2543), .Q(n16897) );
  OR2X1 U17315 ( .IN1(n16899), .IN2(n16900), .Q(g24235) );
  AND2X1 U17316 ( .IN1(n16901), .IN2(g1172), .Q(n16900) );
  AND2X1 U17317 ( .IN1(n4465), .IN2(g1158), .Q(n16899) );
  OR2X1 U17318 ( .IN1(n16902), .IN2(n16903), .Q(g24231) );
  AND2X1 U17319 ( .IN1(n13368), .IN2(g1866), .Q(n16903) );
  AND2X1 U17320 ( .IN1(n4464), .IN2(g1860), .Q(n16902) );
  OR2X1 U17321 ( .IN1(n16904), .IN2(n16905), .Q(g24230) );
  AND2X1 U17322 ( .IN1(n16894), .IN2(g8082), .Q(n16905) );
  AND2X1 U17323 ( .IN1(n4457), .IN2(g1849), .Q(n16904) );
  OR2X1 U17324 ( .IN1(n16906), .IN2(n16907), .Q(g24228) );
  AND2X1 U17325 ( .IN1(n16908), .IN2(g485), .Q(n16907) );
  AND2X1 U17326 ( .IN1(n4466), .IN2(g471), .Q(n16906) );
  OR2X1 U17327 ( .IN1(n16909), .IN2(n16910), .Q(g24226) );
  AND2X1 U17328 ( .IN1(n13236), .IN2(g8167), .Q(n16910) );
  AND2X1 U17329 ( .IN1(n4455), .IN2(g2553), .Q(n16909) );
  OR2X1 U17330 ( .IN1(n16911), .IN2(n16912), .Q(g24225) );
  AND2X1 U17331 ( .IN1(n16891), .IN2(g8087), .Q(n16912) );
  INVX0 U17332 ( .INP(n10871), .ZN(n16891) );
  OR2X1 U17333 ( .IN1(n12245), .IN2(n12262), .Q(n10871) );
  OR2X1 U17334 ( .IN1(n12241), .IN2(n12227), .Q(n12262) );
  AND2X1 U17335 ( .IN1(n4456), .IN2(g2540), .Q(n16911) );
  OR2X1 U17336 ( .IN1(n16913), .IN2(n16914), .Q(g24223) );
  AND2X1 U17337 ( .IN1(n13499), .IN2(g1172), .Q(n16914) );
  AND2X1 U17338 ( .IN1(n4465), .IN2(g1166), .Q(n16913) );
  OR2X1 U17339 ( .IN1(n16915), .IN2(n16916), .Q(g24222) );
  AND2X1 U17340 ( .IN1(n16901), .IN2(g8007), .Q(n16916) );
  AND2X1 U17341 ( .IN1(n4459), .IN2(g1155), .Q(n16915) );
  OR2X1 U17342 ( .IN1(n16917), .IN2(n16918), .Q(g24219) );
  AND2X1 U17343 ( .IN1(n13368), .IN2(g8082), .Q(n16918) );
  AND2X1 U17344 ( .IN1(n4457), .IN2(g1859), .Q(n16917) );
  OR2X1 U17345 ( .IN1(n16919), .IN2(n16920), .Q(g24218) );
  AND2X1 U17346 ( .IN1(n16894), .IN2(g8012), .Q(n16920) );
  INVX0 U17347 ( .INP(n10807), .ZN(n16894) );
  OR2X1 U17348 ( .IN1(n11782), .IN2(n11799), .Q(n10807) );
  OR2X1 U17349 ( .IN1(n11778), .IN2(n11764), .Q(n11799) );
  AND2X1 U17350 ( .IN1(n4458), .IN2(g1846), .Q(n16919) );
  OR2X1 U17351 ( .IN1(n16921), .IN2(n16922), .Q(g24216) );
  AND2X1 U17352 ( .IN1(n13620), .IN2(g485), .Q(n16922) );
  AND2X1 U17353 ( .IN1(n4466), .IN2(g479), .Q(n16921) );
  OR2X1 U17354 ( .IN1(n16923), .IN2(n16924), .Q(g24215) );
  AND2X1 U17355 ( .IN1(test_so24), .IN2(n4461), .Q(n16924) );
  AND2X1 U17356 ( .IN1(n16908), .IN2(g7956), .Q(n16923) );
  OR2X1 U17357 ( .IN1(n16925), .IN2(n16926), .Q(g24214) );
  AND2X1 U17358 ( .IN1(n13236), .IN2(g8087), .Q(n16926) );
  INVX0 U17359 ( .INP(n12631), .ZN(n13236) );
  OR2X1 U17360 ( .IN1(n12227), .IN2(n16927), .Q(n12631) );
  OR2X1 U17361 ( .IN1(n12261), .IN2(n12238), .Q(n16927) );
  INVX0 U17362 ( .INP(n12241), .ZN(n12238) );
  AND2X1 U17363 ( .IN1(n4456), .IN2(g2552), .Q(n16925) );
  OR2X1 U17364 ( .IN1(n16928), .IN2(n16929), .Q(g24213) );
  AND2X1 U17365 ( .IN1(n13499), .IN2(g8007), .Q(n16929) );
  AND2X1 U17366 ( .IN1(n4459), .IN2(g1165), .Q(n16928) );
  OR2X1 U17367 ( .IN1(n16930), .IN2(n16931), .Q(g24212) );
  AND2X1 U17368 ( .IN1(n16901), .IN2(g7961), .Q(n16931) );
  INVX0 U17369 ( .INP(n10742), .ZN(n16901) );
  OR2X1 U17370 ( .IN1(n11564), .IN2(n11624), .Q(n10742) );
  OR2X1 U17371 ( .IN1(n11566), .IN2(n11575), .Q(n11624) );
  AND2X1 U17372 ( .IN1(n4460), .IN2(g1152), .Q(n16930) );
  OR2X1 U17373 ( .IN1(n16932), .IN2(n16933), .Q(g24209) );
  AND2X1 U17374 ( .IN1(n10866), .IN2(g2560), .Q(n16933) );
  AND2X1 U17375 ( .IN1(n4463), .IN2(g2536), .Q(n16932) );
  OR2X1 U17376 ( .IN1(n16934), .IN2(n16935), .Q(g24208) );
  AND2X1 U17377 ( .IN1(n13368), .IN2(g8012), .Q(n16935) );
  INVX0 U17378 ( .INP(n12693), .ZN(n13368) );
  OR2X1 U17379 ( .IN1(n11764), .IN2(n16936), .Q(n12693) );
  OR2X1 U17380 ( .IN1(n11798), .IN2(n11775), .Q(n16936) );
  INVX0 U17381 ( .INP(n11778), .ZN(n11775) );
  AND2X1 U17382 ( .IN1(n4458), .IN2(g1858), .Q(n16934) );
  OR2X1 U17383 ( .IN1(n16937), .IN2(n16938), .Q(g24207) );
  AND2X1 U17384 ( .IN1(n13620), .IN2(g7956), .Q(n16938) );
  AND2X1 U17385 ( .IN1(n4461), .IN2(g478), .Q(n16937) );
  OR2X1 U17386 ( .IN1(n16939), .IN2(n16940), .Q(g24206) );
  AND2X1 U17387 ( .IN1(test_so23), .IN2(n16908), .Q(n16940) );
  INVX0 U17388 ( .INP(n10678), .ZN(n16908) );
  OR2X1 U17389 ( .IN1(n11835), .IN2(n11852), .Q(n10678) );
  OR2X1 U17390 ( .IN1(n11831), .IN2(n11817), .Q(n11852) );
  AND2X1 U17391 ( .IN1(g465), .IN2(n10190), .Q(n16939) );
  OR2X1 U17392 ( .IN1(n16941), .IN2(n16942), .Q(g24182) );
  AND2X1 U17393 ( .IN1(n10801), .IN2(g1866), .Q(n16942) );
  AND2X1 U17394 ( .IN1(n4464), .IN2(g1842), .Q(n16941) );
  OR2X1 U17395 ( .IN1(n16943), .IN2(n16944), .Q(g24181) );
  AND2X1 U17396 ( .IN1(n13499), .IN2(g7961), .Q(n16944) );
  INVX0 U17397 ( .INP(n12754), .ZN(n13499) );
  OR2X1 U17398 ( .IN1(n11575), .IN2(n16945), .Q(n12754) );
  OR2X1 U17399 ( .IN1(n11569), .IN2(n11562), .Q(n16945) );
  INVX0 U17400 ( .INP(n11566), .ZN(n11562) );
  AND2X1 U17401 ( .IN1(n4460), .IN2(g1164), .Q(n16943) );
  OR2X1 U17402 ( .IN1(n16946), .IN2(n16947), .Q(g24179) );
  AND2X1 U17403 ( .IN1(n10737), .IN2(g1172), .Q(n16947) );
  AND2X1 U17404 ( .IN1(n4465), .IN2(g1148), .Q(n16946) );
  OR2X1 U17405 ( .IN1(n16948), .IN2(n16949), .Q(g24178) );
  AND2X1 U17406 ( .IN1(test_so23), .IN2(n13620), .Q(n16949) );
  INVX0 U17407 ( .INP(n12811), .ZN(n13620) );
  OR2X1 U17408 ( .IN1(n11817), .IN2(n16950), .Q(n12811) );
  OR2X1 U17409 ( .IN1(n11851), .IN2(n11828), .Q(n16950) );
  INVX0 U17410 ( .INP(n11831), .ZN(n11828) );
  AND2X1 U17411 ( .IN1(g477), .IN2(n10190), .Q(n16948) );
  OR2X1 U17412 ( .IN1(n16951), .IN2(n16952), .Q(g24174) );
  AND2X1 U17413 ( .IN1(n10671), .IN2(g485), .Q(n16952) );
  AND2X1 U17414 ( .IN1(n4466), .IN2(g461), .Q(n16951) );
  OR2X1 U17415 ( .IN1(n16953), .IN2(n16954), .Q(g24092) );
  AND2X1 U17416 ( .IN1(n10974), .IN2(g2380), .Q(n16954) );
  AND2X1 U17417 ( .IN1(g3229), .IN2(n4483), .Q(n16953) );
  OR2X1 U17418 ( .IN1(n16955), .IN2(n16956), .Q(g24083) );
  AND2X1 U17419 ( .IN1(n10974), .IN2(g1686), .Q(n16956) );
  AND2X1 U17420 ( .IN1(g3229), .IN2(n4484), .Q(n16955) );
  OR2X1 U17421 ( .IN1(n16957), .IN2(n16958), .Q(g24072) );
  AND2X1 U17422 ( .IN1(n10974), .IN2(g992), .Q(n16958) );
  AND2X1 U17423 ( .IN1(g3229), .IN2(n4486), .Q(n16957) );
  OR2X1 U17424 ( .IN1(n16959), .IN2(n16960), .Q(g24059) );
  AND2X1 U17425 ( .IN1(n10974), .IN2(g305), .Q(n16960) );
  INVX0 U17426 ( .INP(g3229), .ZN(n10974) );
  AND2X1 U17427 ( .IN1(g3229), .IN2(n4485), .Q(n16959) );
  OR2X1 U17428 ( .IN1(n16961), .IN2(n16962), .Q(g23418) );
  AND2X1 U17429 ( .IN1(n10866), .IN2(g8167), .Q(n16962) );
  AND2X1 U17430 ( .IN1(n4455), .IN2(g2533), .Q(n16961) );
  OR2X1 U17431 ( .IN1(n16963), .IN2(n16964), .Q(g23413) );
  AND2X1 U17432 ( .IN1(test_so65), .IN2(n4457), .Q(n16964) );
  AND2X1 U17433 ( .IN1(n10801), .IN2(g8082), .Q(n16963) );
  OR2X1 U17434 ( .IN1(n16965), .IN2(n16966), .Q(g23407) );
  AND2X1 U17435 ( .IN1(n10866), .IN2(g8087), .Q(n16966) );
  AND2X1 U17436 ( .IN1(n12261), .IN2(n16967), .Q(n10866) );
  AND2X1 U17437 ( .IN1(n12227), .IN2(n12241), .Q(n16967) );
  OR2X1 U17438 ( .IN1(n16968), .IN2(n16969), .Q(n12241) );
  OR2X1 U17439 ( .IN1(n16970), .IN2(n16971), .Q(n16969) );
  AND2X1 U17440 ( .IN1(n9454), .IN2(n13116), .Q(n16971) );
  AND2X1 U17441 ( .IN1(n9453), .IN2(n13101), .Q(n16970) );
  AND2X1 U17442 ( .IN1(n9444), .IN2(n13106), .Q(n16968) );
  OR2X1 U17443 ( .IN1(n16972), .IN2(n16973), .Q(n12227) );
  OR2X1 U17444 ( .IN1(n16974), .IN2(n16975), .Q(n16973) );
  AND2X1 U17445 ( .IN1(n9456), .IN2(n13116), .Q(n16975) );
  AND2X1 U17446 ( .IN1(n9455), .IN2(n13101), .Q(n16974) );
  AND2X1 U17447 ( .IN1(n9445), .IN2(n13106), .Q(n16972) );
  INVX0 U17448 ( .INP(n12245), .ZN(n12261) );
  OR2X1 U17449 ( .IN1(n16976), .IN2(n16977), .Q(n12245) );
  OR2X1 U17450 ( .IN1(n16978), .IN2(n16979), .Q(n16977) );
  AND2X1 U17451 ( .IN1(n9458), .IN2(n13116), .Q(n16979) );
  INVX0 U17452 ( .INP(n4516), .ZN(n13116) );
  AND2X1 U17453 ( .IN1(n9457), .IN2(n13101), .Q(n16978) );
  INVX0 U17454 ( .INP(n4509), .ZN(n13101) );
  AND2X1 U17455 ( .IN1(n9446), .IN2(n13106), .Q(n16976) );
  INVX0 U17456 ( .INP(n4524), .ZN(n13106) );
  AND2X1 U17457 ( .IN1(n4456), .IN2(g2530), .Q(n16965) );
  OR2X1 U17458 ( .IN1(n16980), .IN2(n16981), .Q(g23406) );
  AND2X1 U17459 ( .IN1(n10737), .IN2(g8007), .Q(n16981) );
  AND2X1 U17460 ( .IN1(n4459), .IN2(g1145), .Q(n16980) );
  OR2X1 U17461 ( .IN1(n16982), .IN2(n16983), .Q(g23400) );
  AND2X1 U17462 ( .IN1(n10801), .IN2(g8012), .Q(n16983) );
  AND2X1 U17463 ( .IN1(n11798), .IN2(n16984), .Q(n10801) );
  AND2X1 U17464 ( .IN1(n11764), .IN2(n11778), .Q(n16984) );
  OR2X1 U17465 ( .IN1(n16985), .IN2(n16986), .Q(n11778) );
  OR2X1 U17466 ( .IN1(n16987), .IN2(n16988), .Q(n16986) );
  AND2X1 U17467 ( .IN1(n9460), .IN2(n13248), .Q(n16988) );
  AND2X1 U17468 ( .IN1(n9459), .IN2(n13111), .Q(n16987) );
  AND2X1 U17469 ( .IN1(n9447), .IN2(n13239), .Q(n16985) );
  OR2X1 U17470 ( .IN1(n16989), .IN2(n16990), .Q(n11764) );
  OR2X1 U17471 ( .IN1(n16991), .IN2(n16992), .Q(n16990) );
  AND2X1 U17472 ( .IN1(n9462), .IN2(n13248), .Q(n16992) );
  AND2X1 U17473 ( .IN1(n9461), .IN2(n13111), .Q(n16991) );
  AND2X1 U17474 ( .IN1(n9448), .IN2(n13239), .Q(n16989) );
  INVX0 U17475 ( .INP(n11782), .ZN(n11798) );
  OR2X1 U17476 ( .IN1(n16993), .IN2(n16994), .Q(n11782) );
  OR2X1 U17477 ( .IN1(n16995), .IN2(n16996), .Q(n16994) );
  AND2X1 U17478 ( .IN1(n9464), .IN2(n13248), .Q(n16996) );
  INVX0 U17479 ( .INP(n4518), .ZN(n13248) );
  AND2X1 U17480 ( .IN1(n9463), .IN2(n13111), .Q(n16995) );
  INVX0 U17481 ( .INP(n4511), .ZN(n13111) );
  AND2X1 U17482 ( .IN1(n9449), .IN2(n13239), .Q(n16993) );
  INVX0 U17483 ( .INP(n4525), .ZN(n13239) );
  AND2X1 U17484 ( .IN1(n4458), .IN2(g1836), .Q(n16982) );
  OR2X1 U17485 ( .IN1(n16997), .IN2(n16998), .Q(g23399) );
  AND2X1 U17486 ( .IN1(n10671), .IN2(g7956), .Q(n16998) );
  AND2X1 U17487 ( .IN1(n4461), .IN2(g458), .Q(n16997) );
  OR2X1 U17488 ( .IN1(n16999), .IN2(n17000), .Q(g23392) );
  AND2X1 U17489 ( .IN1(n10737), .IN2(g7961), .Q(n17000) );
  AND2X1 U17490 ( .IN1(n11569), .IN2(n17001), .Q(n10737) );
  AND2X1 U17491 ( .IN1(n11575), .IN2(n11566), .Q(n17001) );
  OR2X1 U17492 ( .IN1(n17002), .IN2(n17003), .Q(n11566) );
  OR2X1 U17493 ( .IN1(n17004), .IN2(n17005), .Q(n17003) );
  AND2X1 U17494 ( .IN1(n9450), .IN2(g6712), .Q(n17005) );
  AND2X1 U17495 ( .IN1(n9465), .IN2(g5472), .Q(n17004) );
  INVX0 U17496 ( .INP(n17006), .ZN(n17002) );
  OR2X1 U17497 ( .IN1(n4381), .IN2(test_so39), .Q(n17006) );
  OR2X1 U17498 ( .IN1(n17007), .IN2(n17008), .Q(n11575) );
  OR2X1 U17499 ( .IN1(n17009), .IN2(n17010), .Q(n17008) );
  AND2X1 U17500 ( .IN1(n9451), .IN2(g6712), .Q(n17010) );
  AND2X1 U17501 ( .IN1(n9467), .IN2(g5472), .Q(n17009) );
  AND2X1 U17502 ( .IN1(n9466), .IN2(g1088), .Q(n17007) );
  INVX0 U17503 ( .INP(n11564), .ZN(n11569) );
  OR2X1 U17504 ( .IN1(n17011), .IN2(n17012), .Q(n11564) );
  OR2X1 U17505 ( .IN1(n17013), .IN2(n17014), .Q(n17012) );
  AND2X1 U17506 ( .IN1(n9452), .IN2(g6712), .Q(n17014) );
  AND2X1 U17507 ( .IN1(n9469), .IN2(g5472), .Q(n17013) );
  AND2X1 U17508 ( .IN1(n9468), .IN2(g1088), .Q(n17011) );
  AND2X1 U17509 ( .IN1(n4460), .IN2(g1142), .Q(n16999) );
  OR2X1 U17510 ( .IN1(n17015), .IN2(n17016), .Q(g23385) );
  AND2X1 U17511 ( .IN1(n10671), .IN2(test_so23), .Q(n17016) );
  AND2X1 U17512 ( .IN1(n11851), .IN2(n17017), .Q(n10671) );
  AND2X1 U17513 ( .IN1(n11817), .IN2(n11831), .Q(n17017) );
  OR2X1 U17514 ( .IN1(n17018), .IN2(n17019), .Q(n11831) );
  OR2X1 U17515 ( .IN1(n17020), .IN2(n17021), .Q(n17019) );
  AND2X1 U17516 ( .IN1(n9470), .IN2(n13375), .Q(n17021) );
  AND2X1 U17517 ( .IN1(n9471), .IN2(n13502), .Q(n17020) );
  AND2X1 U17518 ( .IN1(n9472), .IN2(n13506), .Q(n17018) );
  OR2X1 U17519 ( .IN1(n17022), .IN2(n17023), .Q(n11817) );
  OR2X1 U17520 ( .IN1(n17024), .IN2(n17025), .Q(n17023) );
  AND2X1 U17521 ( .IN1(n9473), .IN2(n13375), .Q(n17025) );
  AND2X1 U17522 ( .IN1(n13502), .IN2(n10222), .Q(n17024) );
  AND2X1 U17523 ( .IN1(n9474), .IN2(n13506), .Q(n17022) );
  INVX0 U17524 ( .INP(n11835), .ZN(n11851) );
  OR2X1 U17525 ( .IN1(n17026), .IN2(n17027), .Q(n11835) );
  OR2X1 U17526 ( .IN1(n17028), .IN2(n17029), .Q(n17027) );
  AND2X1 U17527 ( .IN1(n9475), .IN2(n13375), .Q(n17029) );
  INVX0 U17528 ( .INP(n4506), .ZN(n13375) );
  AND2X1 U17529 ( .IN1(n9476), .IN2(n13502), .Q(n17028) );
  INVX0 U17530 ( .INP(n4499), .ZN(n13502) );
  AND2X1 U17531 ( .IN1(n9477), .IN2(n13506), .Q(n17026) );
  INVX0 U17532 ( .INP(n4520), .ZN(n13506) );
  AND2X1 U17533 ( .IN1(g455), .IN2(n10190), .Q(n17015) );
  AND2X1 U17534 ( .IN1(n17030), .IN2(n10931), .Q(g23359) );
  OR2X1 U17535 ( .IN1(n17031), .IN2(n15352), .Q(n10931) );
  AND2X1 U17536 ( .IN1(n17032), .IN2(n17033), .Q(n17031) );
  OR2X1 U17537 ( .IN1(n17034), .IN2(n17035), .Q(n17032) );
  INVX0 U17538 ( .INP(n17036), .ZN(n17035) );
  AND2X1 U17539 ( .IN1(n4350), .IN2(n4480), .Q(n17036) );
  OR2X1 U17540 ( .IN1(n4481), .IN2(n10157), .Q(n17034) );
  AND2X1 U17541 ( .IN1(n4102), .IN2(n17037), .Q(n17030) );
  INVX0 U17542 ( .INP(n17038), .ZN(n17037) );
  AND2X1 U17543 ( .IN1(n10933), .IN2(n4350), .Q(n17038) );
  OR2X1 U17544 ( .IN1(n4350), .IN2(n10933), .Q(n4102) );
  OR2X1 U17545 ( .IN1(n17039), .IN2(n17040), .Q(n10933) );
  OR2X1 U17546 ( .IN1(n4481), .IN2(n10165), .Q(n17040) );
  AND2X1 U17547 ( .IN1(n17041), .IN2(n11730), .Q(g23358) );
  AND2X1 U17548 ( .IN1(n16857), .IN2(n17042), .Q(n17041) );
  INVX0 U17549 ( .INP(n4122_Tj_Payload), .ZN(n17042) );
  OR2X1 U17550 ( .IN1(n4431), .IN2(n4123), .Q(n16857) );
  AND2X1 U17551 ( .IN1(n17043), .IN2(n10874), .Q(g23357) );
  OR2X1 U17552 ( .IN1(n17044), .IN2(n11730), .Q(n10874) );
  AND2X1 U17553 ( .IN1(n18258), .IN2(n17045), .Q(n17044) );
  OR2X1 U17554 ( .IN1(n17046), .IN2(n17047), .Q(n17045) );
  OR2X1 U17555 ( .IN1(g2924), .IN2(g2917), .Q(n17047) );
  OR2X1 U17556 ( .IN1(n9892), .IN2(n4482), .Q(n17046) );
  AND2X1 U17557 ( .IN1(n17048), .IN2(n17049), .Q(n17043) );
  OR2X1 U17558 ( .IN1(n10876), .IN2(g2917), .Q(n17049) );
  INVX0 U17559 ( .INP(n16853), .ZN(n10876) );
  OR2X1 U17560 ( .IN1(n4479), .IN2(n16853), .Q(n17048) );
  OR2X1 U17561 ( .IN1(n4482), .IN2(n10877), .Q(n16853) );
  AND2X1 U17562 ( .IN1(n17050), .IN2(n14331), .Q(g23348) );
  AND2X1 U17563 ( .IN1(n17051), .IN2(n17052), .Q(n17050) );
  OR2X1 U17564 ( .IN1(n16868), .IN2(g2727), .Q(n17052) );
  INVX0 U17565 ( .INP(n16869), .ZN(n16868) );
  OR2X1 U17566 ( .IN1(n4419), .IN2(n16869), .Q(n17051) );
  AND2X1 U17567 ( .IN1(n17053), .IN2(n14337), .Q(g23339) );
  AND2X1 U17568 ( .IN1(n17054), .IN2(n17055), .Q(n17053) );
  OR2X1 U17569 ( .IN1(n16874), .IN2(g2033), .Q(n17055) );
  INVX0 U17570 ( .INP(n16875), .ZN(n16874) );
  OR2X1 U17571 ( .IN1(n4420), .IN2(n16875), .Q(n17054) );
  AND2X1 U17572 ( .IN1(n17056), .IN2(n15352), .Q(g23330) );
  INVX0 U17573 ( .INP(n15912), .ZN(n15352) );
  OR2X1 U17574 ( .IN1(n10934), .IN2(g3234), .Q(n15912) );
  AND2X1 U17575 ( .IN1(n17057), .IN2(n4598), .Q(n10934) );
  AND2X1 U17576 ( .IN1(n17058), .IN2(n4066), .Q(n17056) );
  OR2X1 U17577 ( .IN1(n15916), .IN2(n17059), .Q(n4066) );
  OR2X1 U17578 ( .IN1(n18262), .IN2(n10164), .Q(n17059) );
  OR2X1 U17579 ( .IN1(n17060), .IN2(g3006), .Q(n17058) );
  AND2X1 U17580 ( .IN1(n15915), .IN2(n7909), .Q(n17060) );
  INVX0 U17581 ( .INP(n15916), .ZN(n15915) );
  OR2X1 U17582 ( .IN1(n10165), .IN2(n10166), .Q(n15916) );
  AND2X1 U17583 ( .IN1(n17061), .IN2(n14345), .Q(g23329) );
  AND2X1 U17584 ( .IN1(n17062), .IN2(n17063), .Q(n17061) );
  OR2X1 U17585 ( .IN1(n16880), .IN2(g1339), .Q(n17063) );
  INVX0 U17586 ( .INP(n16881), .ZN(n16880) );
  OR2X1 U17587 ( .IN1(n4421), .IN2(n16881), .Q(n17062) );
  AND2X1 U17588 ( .IN1(n17064), .IN2(n13809), .Q(g23324) );
  AND2X1 U17589 ( .IN1(n17065), .IN2(n17066), .Q(n17064) );
  OR2X1 U17590 ( .IN1(n16886), .IN2(g653), .Q(n17066) );
  INVX0 U17591 ( .INP(n16887), .ZN(n16886) );
  OR2X1 U17592 ( .IN1(n4422), .IN2(n16887), .Q(n17065) );
  OR2X1 U17593 ( .IN1(n17067), .IN2(n17068), .Q(g23137) );
  AND2X1 U17594 ( .IN1(n15233), .IN2(g1866), .Q(n17068) );
  AND2X1 U17595 ( .IN1(n4464), .IN2(g1869), .Q(n17067) );
  AND2X1 U17596 ( .IN1(n17069), .IN2(n17070), .Q(g23136) );
  OR2X1 U17597 ( .IN1(n17071), .IN2(g633), .Q(n17070) );
  INVX0 U17598 ( .INP(n17072), .ZN(n17071) );
  AND2X1 U17599 ( .IN1(n16887), .IN2(n13809), .Q(n17069) );
  OR2X1 U17600 ( .IN1(n4478), .IN2(n17072), .Q(n16887) );
  OR2X1 U17601 ( .IN1(n17073), .IN2(n17074), .Q(g23133) );
  AND2X1 U17602 ( .IN1(n15191), .IN2(g8167), .Q(n17074) );
  AND2X1 U17603 ( .IN1(n4455), .IN2(g2562), .Q(n17073) );
  OR2X1 U17604 ( .IN1(n17075), .IN2(n17076), .Q(g23132) );
  AND2X1 U17605 ( .IN1(n13016), .IN2(g8087), .Q(n17076) );
  AND2X1 U17606 ( .IN1(n4456), .IN2(g2555), .Q(n17075) );
  OR2X1 U17607 ( .IN1(n17077), .IN2(n17078), .Q(g23126) );
  AND2X1 U17608 ( .IN1(n15275), .IN2(g1172), .Q(n17078) );
  AND2X1 U17609 ( .IN1(n4465), .IN2(g1175), .Q(n17077) );
  OR2X1 U17610 ( .IN1(n17079), .IN2(n17080), .Q(g23124) );
  AND2X1 U17611 ( .IN1(n15233), .IN2(g8082), .Q(n17080) );
  AND2X1 U17612 ( .IN1(n4457), .IN2(g1868), .Q(n17079) );
  OR2X1 U17613 ( .IN1(n17081), .IN2(n17082), .Q(g23123) );
  AND2X1 U17614 ( .IN1(n13040), .IN2(g8012), .Q(n17082) );
  AND2X1 U17615 ( .IN1(n4458), .IN2(g1861), .Q(n17081) );
  OR2X1 U17616 ( .IN1(n17083), .IN2(n17084), .Q(g23117) );
  AND2X1 U17617 ( .IN1(n15314), .IN2(g485), .Q(n17084) );
  AND2X1 U17618 ( .IN1(n4466), .IN2(g488), .Q(n17083) );
  OR2X1 U17619 ( .IN1(n17085), .IN2(n17086), .Q(g23114) );
  AND2X1 U17620 ( .IN1(n15191), .IN2(g8087), .Q(n17086) );
  AND2X1 U17621 ( .IN1(n4456), .IN2(g2561), .Q(n17085) );
  OR2X1 U17622 ( .IN1(n17087), .IN2(n17088), .Q(g23111) );
  AND2X1 U17623 ( .IN1(n15275), .IN2(g8007), .Q(n17088) );
  AND2X1 U17624 ( .IN1(test_so44), .IN2(n4459), .Q(n17087) );
  OR2X1 U17625 ( .IN1(n17089), .IN2(n17090), .Q(g23110) );
  AND2X1 U17626 ( .IN1(n13064), .IN2(g7961), .Q(n17090) );
  AND2X1 U17627 ( .IN1(n4460), .IN2(g1167), .Q(n17089) );
  OR2X1 U17628 ( .IN1(n17091), .IN2(n17092), .Q(g23097) );
  AND2X1 U17629 ( .IN1(n15233), .IN2(g8012), .Q(n17092) );
  OR2X1 U17630 ( .IN1(n17093), .IN2(n17094), .Q(n15233) );
  OR2X1 U17631 ( .IN1(n17095), .IN2(n17096), .Q(n17094) );
  AND2X1 U17632 ( .IN1(g7014), .IN2(g1822), .Q(n17096) );
  AND2X1 U17633 ( .IN1(test_so59), .IN2(n4618), .Q(n17095) );
  AND2X1 U17634 ( .IN1(g5511), .IN2(g1819), .Q(n17093) );
  AND2X1 U17635 ( .IN1(n4458), .IN2(g1867), .Q(n17091) );
  OR2X1 U17636 ( .IN1(n17097), .IN2(n17098), .Q(g23093) );
  AND2X1 U17637 ( .IN1(n15314), .IN2(g7956), .Q(n17098) );
  AND2X1 U17638 ( .IN1(n4461), .IN2(g487), .Q(n17097) );
  OR2X1 U17639 ( .IN1(n17099), .IN2(n17100), .Q(g23092) );
  AND2X1 U17640 ( .IN1(test_so23), .IN2(n13085), .Q(n17100) );
  AND2X1 U17641 ( .IN1(g480), .IN2(n10190), .Q(n17099) );
  OR2X1 U17642 ( .IN1(n17101), .IN2(n17102), .Q(g23081) );
  AND2X1 U17643 ( .IN1(n15275), .IN2(g7961), .Q(n17102) );
  OR2X1 U17644 ( .IN1(n17103), .IN2(n17104), .Q(n15275) );
  OR2X1 U17645 ( .IN1(n17105), .IN2(n17106), .Q(n17104) );
  AND2X1 U17646 ( .IN1(g6712), .IN2(g1128), .Q(n17106) );
  AND2X1 U17647 ( .IN1(g5472), .IN2(g1125), .Q(n17105) );
  AND2X1 U17648 ( .IN1(g1088), .IN2(g1131), .Q(n17103) );
  AND2X1 U17649 ( .IN1(n4460), .IN2(g1173), .Q(n17101) );
  OR2X1 U17650 ( .IN1(n17107), .IN2(n17108), .Q(g23076) );
  AND2X1 U17651 ( .IN1(n13016), .IN2(g2560), .Q(n17108) );
  AND2X1 U17652 ( .IN1(n4463), .IN2(g2539), .Q(n17107) );
  OR2X1 U17653 ( .IN1(n17109), .IN2(n17110), .Q(g23067) );
  AND2X1 U17654 ( .IN1(test_so23), .IN2(n15314), .Q(n17110) );
  OR2X1 U17655 ( .IN1(n17111), .IN2(n17112), .Q(n15314) );
  OR2X1 U17656 ( .IN1(n17113), .IN2(n17114), .Q(n17112) );
  AND2X1 U17657 ( .IN1(g6447), .IN2(g441), .Q(n17114) );
  AND2X1 U17658 ( .IN1(n4640), .IN2(g444), .Q(n17113) );
  AND2X1 U17659 ( .IN1(g5437), .IN2(g438), .Q(n17111) );
  AND2X1 U17660 ( .IN1(g486), .IN2(n10190), .Q(n17109) );
  OR2X1 U17661 ( .IN1(n17115), .IN2(n17116), .Q(g23058) );
  AND2X1 U17662 ( .IN1(n13040), .IN2(g1866), .Q(n17116) );
  AND2X1 U17663 ( .IN1(n4464), .IN2(g1845), .Q(n17115) );
  OR2X1 U17664 ( .IN1(n17117), .IN2(n17118), .Q(g23047) );
  AND2X1 U17665 ( .IN1(n13016), .IN2(g8167), .Q(n17118) );
  INVX0 U17666 ( .INP(n4285), .ZN(n13016) );
  OR2X1 U17667 ( .IN1(n17119), .IN2(n17120), .Q(n4285) );
  OR2X1 U17668 ( .IN1(n17121), .IN2(n17122), .Q(n17120) );
  AND2X1 U17669 ( .IN1(g7264), .IN2(g2495), .Q(n17122) );
  AND2X1 U17670 ( .IN1(n4606), .IN2(g2498), .Q(n17121) );
  AND2X1 U17671 ( .IN1(g5555), .IN2(g2492), .Q(n17119) );
  AND2X1 U17672 ( .IN1(n4455), .IN2(g2559), .Q(n17117) );
  OR2X1 U17673 ( .IN1(n17123), .IN2(n17124), .Q(g23039) );
  AND2X1 U17674 ( .IN1(n13064), .IN2(g1172), .Q(n17124) );
  AND2X1 U17675 ( .IN1(n4465), .IN2(g1151), .Q(n17123) );
  OR2X1 U17676 ( .IN1(n17125), .IN2(n17126), .Q(g23030) );
  AND2X1 U17677 ( .IN1(n13040), .IN2(g8082), .Q(n17126) );
  INVX0 U17678 ( .INP(n4284), .ZN(n13040) );
  OR2X1 U17679 ( .IN1(n17127), .IN2(n17128), .Q(n4284) );
  OR2X1 U17680 ( .IN1(n17129), .IN2(n17130), .Q(n17128) );
  AND2X1 U17681 ( .IN1(g7014), .IN2(g1801), .Q(n17130) );
  AND2X1 U17682 ( .IN1(n4618), .IN2(g1804), .Q(n17129) );
  AND2X1 U17683 ( .IN1(g5511), .IN2(g1798), .Q(n17127) );
  AND2X1 U17684 ( .IN1(n4457), .IN2(g1865), .Q(n17125) );
  OR2X1 U17685 ( .IN1(n17131), .IN2(n17132), .Q(g23022) );
  AND2X1 U17686 ( .IN1(n13085), .IN2(g485), .Q(n17132) );
  AND2X1 U17687 ( .IN1(n4466), .IN2(g464), .Q(n17131) );
  OR2X1 U17688 ( .IN1(n17133), .IN2(n17134), .Q(g23014) );
  AND2X1 U17689 ( .IN1(n13064), .IN2(g8007), .Q(n17134) );
  INVX0 U17690 ( .INP(n4283), .ZN(n13064) );
  OR2X1 U17691 ( .IN1(n17135), .IN2(n17136), .Q(n4283) );
  OR2X1 U17692 ( .IN1(n17137), .IN2(n17138), .Q(n17136) );
  AND2X1 U17693 ( .IN1(g6712), .IN2(g1107), .Q(n17138) );
  AND2X1 U17694 ( .IN1(g5472), .IN2(g1104), .Q(n17137) );
  AND2X1 U17695 ( .IN1(g1088), .IN2(g1110), .Q(n17135) );
  AND2X1 U17696 ( .IN1(n4459), .IN2(g1171), .Q(n17133) );
  OR2X1 U17697 ( .IN1(n17139), .IN2(n17140), .Q(g23000) );
  AND2X1 U17698 ( .IN1(n13085), .IN2(g7956), .Q(n17140) );
  INVX0 U17699 ( .INP(n4282), .ZN(n13085) );
  OR2X1 U17700 ( .IN1(n17141), .IN2(n17142), .Q(n4282) );
  OR2X1 U17701 ( .IN1(n17143), .IN2(n17144), .Q(n17142) );
  AND2X1 U17702 ( .IN1(g6447), .IN2(g420), .Q(n17144) );
  AND2X1 U17703 ( .IN1(n4640), .IN2(g423), .Q(n17143) );
  AND2X1 U17704 ( .IN1(g5437), .IN2(g417), .Q(n17141) );
  AND2X1 U17705 ( .IN1(n4461), .IN2(g484), .Q(n17139) );
  OR2X1 U17706 ( .IN1(n17145), .IN2(n17146), .Q(g22687) );
  AND2X1 U17707 ( .IN1(n17147), .IN2(n17148), .Q(n17146) );
  OR2X1 U17708 ( .IN1(n15751), .IN2(n11213), .Q(n17147) );
  AND2X1 U17709 ( .IN1(n17149), .IN2(n15751), .Q(n17145) );
  INVX0 U17710 ( .INP(n17150), .ZN(n15751) );
  OR2X1 U17711 ( .IN1(n17151), .IN2(n17152), .Q(n17150) );
  OR2X1 U17712 ( .IN1(n17153), .IN2(n17154), .Q(n17152) );
  AND2X1 U17713 ( .IN1(n12862), .IN2(g2565), .Q(n17154) );
  AND2X1 U17714 ( .IN1(g2624), .IN2(g2571), .Q(n17153) );
  AND2X1 U17715 ( .IN1(g7390), .IN2(g2568), .Q(n17151) );
  AND2X1 U17716 ( .IN1(n11146), .IN2(g2584), .Q(n17149) );
  OR2X1 U17717 ( .IN1(n17155), .IN2(n17156), .Q(g22651) );
  AND2X1 U17718 ( .IN1(n17157), .IN2(n17148), .Q(n17156) );
  OR2X1 U17719 ( .IN1(n15760), .IN2(n11375), .Q(n17157) );
  AND2X1 U17720 ( .IN1(n17158), .IN2(n15760), .Q(n17155) );
  INVX0 U17721 ( .INP(n17159), .ZN(n15760) );
  OR2X1 U17722 ( .IN1(n17160), .IN2(n17161), .Q(n17159) );
  OR2X1 U17723 ( .IN1(n17162), .IN2(n17163), .Q(n17161) );
  AND2X1 U17724 ( .IN1(g7194), .IN2(g1874), .Q(n17163) );
  AND2X1 U17725 ( .IN1(test_so68), .IN2(n13973), .Q(n17162) );
  AND2X1 U17726 ( .IN1(g1930), .IN2(g1877), .Q(n17160) );
  AND2X1 U17727 ( .IN1(n11309), .IN2(g1890), .Q(n17158) );
  OR2X1 U17728 ( .IN1(n17164), .IN2(n17165), .Q(g22615) );
  AND2X1 U17729 ( .IN1(n17166), .IN2(n17148), .Q(n17165) );
  OR2X1 U17730 ( .IN1(n15769), .IN2(n11538), .Q(n17166) );
  AND2X1 U17731 ( .IN1(n17167), .IN2(n15769), .Q(n17164) );
  INVX0 U17732 ( .INP(n17168), .ZN(n15769) );
  OR2X1 U17733 ( .IN1(n17169), .IN2(n17170), .Q(n17168) );
  OR2X1 U17734 ( .IN1(n17171), .IN2(n17172), .Q(n17170) );
  AND2X1 U17735 ( .IN1(g6944), .IN2(g1180), .Q(n17172) );
  AND2X1 U17736 ( .IN1(g1236), .IN2(g1183), .Q(n17171) );
  AND2X1 U17737 ( .IN1(test_so47), .IN2(n13842), .Q(n17169) );
  AND2X1 U17738 ( .IN1(n11471), .IN2(g1196), .Q(n17167) );
  OR2X1 U17739 ( .IN1(n17173), .IN2(n17174), .Q(g22578) );
  AND2X1 U17740 ( .IN1(n17175), .IN2(n17148), .Q(n17174) );
  INVX0 U17741 ( .INP(n17176), .ZN(n17148) );
  OR2X1 U17742 ( .IN1(n15775), .IN2(n11046), .Q(n17175) );
  AND2X1 U17743 ( .IN1(n17177), .IN2(n15775), .Q(n17173) );
  INVX0 U17744 ( .INP(n17178), .ZN(n15775) );
  OR2X1 U17745 ( .IN1(n17179), .IN2(n17180), .Q(n17178) );
  OR2X1 U17746 ( .IN1(n17181), .IN2(n17182), .Q(n17180) );
  AND2X1 U17747 ( .IN1(g550), .IN2(g496), .Q(n17182) );
  AND2X1 U17748 ( .IN1(g6485), .IN2(g490), .Q(n17181) );
  AND2X1 U17749 ( .IN1(g6642), .IN2(g493), .Q(n17179) );
  AND2X1 U17750 ( .IN1(test_so22), .IN2(n10961), .Q(n17177) );
  AND2X1 U17751 ( .IN1(n17183), .IN2(n17184), .Q(g22299) );
  OR2X1 U17752 ( .IN1(n16067), .IN2(test_so95), .Q(n17183) );
  AND2X1 U17753 ( .IN1(n17185), .IN2(n14331), .Q(g22284) );
  OR2X1 U17754 ( .IN1(n16072), .IN2(g2813), .Q(n17185) );
  AND2X1 U17755 ( .IN1(n17186), .IN2(n17187), .Q(g22280) );
  OR2X1 U17756 ( .IN1(n4149_Tj_Payload), .IN2(g2117), .Q(n17186) );
  AND2X1 U17757 ( .IN1(n17188), .IN2(n17189), .Q(g22269) );
  OR2X1 U17758 ( .IN1(n16080), .IN2(g2812), .Q(n17188) );
  AND2X1 U17759 ( .IN1(n17190), .IN2(n14337), .Q(g22267) );
  OR2X1 U17760 ( .IN1(n16175), .IN2(g2119), .Q(n17190) );
  AND2X1 U17761 ( .IN1(n17191), .IN2(n17192), .Q(g22263) );
  OR2X1 U17762 ( .IN1(n16180), .IN2(g1423), .Q(n17191) );
  AND2X1 U17763 ( .IN1(n17193), .IN2(n17194), .Q(g22249) );
  OR2X1 U17764 ( .IN1(n16184), .IN2(g2118), .Q(n17193) );
  AND2X1 U17765 ( .IN1(n17195), .IN2(n14345), .Q(g22247) );
  OR2X1 U17766 ( .IN1(n4160_Tj_Payload), .IN2(g1425), .Q(n17195) );
  AND2X1 U17767 ( .IN1(n17196), .IN2(n17197), .Q(g22242) );
  OR2X1 U17768 ( .IN1(n4161_Tj_Payload), .IN2(g737), .Q(n17196) );
  AND2X1 U17769 ( .IN1(n17198), .IN2(n17199), .Q(g22234) );
  OR2X1 U17770 ( .IN1(n16293), .IN2(g1424), .Q(n17198) );
  AND2X1 U17771 ( .IN1(n17200), .IN2(n13809), .Q(g22231) );
  OR2X1 U17772 ( .IN1(n16388), .IN2(g739), .Q(n17200) );
  AND2X1 U17773 ( .IN1(n17201), .IN2(n17202), .Q(g22218) );
  OR2X1 U17774 ( .IN1(n16392), .IN2(g738), .Q(n17201) );
  OR2X1 U17775 ( .IN1(n17203), .IN2(n17204), .Q(g22200) );
  AND2X1 U17776 ( .IN1(n16679), .IN2(g2208), .Q(n17204) );
  AND2X1 U17777 ( .IN1(n17205), .IN2(n4373), .Q(n17203) );
  OR2X1 U17778 ( .IN1(n17206), .IN2(n17207), .Q(g22194) );
  AND2X1 U17779 ( .IN1(n16679), .IN2(g2238), .Q(n17207) );
  AND2X1 U17780 ( .IN1(n17205), .IN2(n11898), .Q(n17206) );
  OR2X1 U17781 ( .IN1(n17208), .IN2(n17209), .Q(g22193) );
  AND2X1 U17782 ( .IN1(n17210), .IN2(g2210), .Q(n17209) );
  AND2X1 U17783 ( .IN1(n17211), .IN2(n4373), .Q(n17208) );
  OR2X1 U17784 ( .IN1(n17212), .IN2(n17213), .Q(g22192) );
  AND2X1 U17785 ( .IN1(n16679), .IN2(g2205), .Q(n17213) );
  AND2X1 U17786 ( .IN1(n17205), .IN2(n4377), .Q(n17212) );
  OR2X1 U17787 ( .IN1(n17214), .IN2(n17215), .Q(g22191) );
  AND2X1 U17788 ( .IN1(n16684), .IN2(g1514), .Q(n17215) );
  AND2X1 U17789 ( .IN1(n17216), .IN2(n4374), .Q(n17214) );
  OR2X1 U17790 ( .IN1(n17217), .IN2(n17218), .Q(g22185) );
  AND2X1 U17791 ( .IN1(n17211), .IN2(n11898), .Q(n17218) );
  AND2X1 U17792 ( .IN1(test_so75), .IN2(n17210), .Q(n17217) );
  OR2X1 U17793 ( .IN1(n17219), .IN2(n17220), .Q(g22184) );
  AND2X1 U17794 ( .IN1(n16679), .IN2(g2235), .Q(n17220) );
  AND2X1 U17795 ( .IN1(n13179), .IN2(n17205), .Q(n17219) );
  OR2X1 U17796 ( .IN1(n17221), .IN2(n17222), .Q(g22183) );
  AND2X1 U17797 ( .IN1(n17223), .IN2(g2209), .Q(n17222) );
  AND2X1 U17798 ( .IN1(n17224), .IN2(n4373), .Q(n17221) );
  OR2X1 U17799 ( .IN1(n17225), .IN2(n17226), .Q(g22182) );
  AND2X1 U17800 ( .IN1(n17210), .IN2(g2207), .Q(n17226) );
  AND2X1 U17801 ( .IN1(n17211), .IN2(n4377), .Q(n17225) );
  OR2X1 U17802 ( .IN1(n17227), .IN2(n17228), .Q(g22180) );
  AND2X1 U17803 ( .IN1(n16684), .IN2(g1544), .Q(n17228) );
  AND2X1 U17804 ( .IN1(n17216), .IN2(n11936), .Q(n17227) );
  OR2X1 U17805 ( .IN1(n17229), .IN2(n17230), .Q(g22179) );
  AND2X1 U17806 ( .IN1(n17231), .IN2(g1516), .Q(n17230) );
  AND2X1 U17807 ( .IN1(n17232), .IN2(n4374), .Q(n17229) );
  OR2X1 U17808 ( .IN1(n17233), .IN2(n17234), .Q(g22178) );
  AND2X1 U17809 ( .IN1(n16684), .IN2(g1511), .Q(n17234) );
  AND2X1 U17810 ( .IN1(n17216), .IN2(n4378), .Q(n17233) );
  OR2X1 U17811 ( .IN1(n17235), .IN2(n17236), .Q(g22177) );
  AND2X1 U17812 ( .IN1(n16689), .IN2(g820), .Q(n17236) );
  AND2X1 U17813 ( .IN1(n17237), .IN2(n4375), .Q(n17235) );
  OR2X1 U17814 ( .IN1(n17238), .IN2(n17239), .Q(g22173) );
  AND2X1 U17815 ( .IN1(n17223), .IN2(g2239), .Q(n17239) );
  AND2X1 U17816 ( .IN1(n17224), .IN2(n11898), .Q(n17238) );
  INVX0 U17817 ( .INP(n13206), .ZN(n11898) );
  OR2X1 U17818 ( .IN1(n17240), .IN2(n17241), .Q(n13206) );
  OR2X1 U17819 ( .IN1(n17242), .IN2(n17243), .Q(n17241) );
  AND2X1 U17820 ( .IN1(n9761), .IN2(g2241), .Q(n17243) );
  AND2X1 U17821 ( .IN1(n9763), .IN2(g6837), .Q(n17242) );
  AND2X1 U17822 ( .IN1(n9762), .IN2(test_so73), .Q(n17240) );
  OR2X1 U17823 ( .IN1(n17244), .IN2(n17245), .Q(g22172) );
  AND2X1 U17824 ( .IN1(n17210), .IN2(g2237), .Q(n17245) );
  AND2X1 U17825 ( .IN1(n17211), .IN2(n13179), .Q(n17244) );
  OR2X1 U17826 ( .IN1(n17246), .IN2(n17247), .Q(g22171) );
  AND2X1 U17827 ( .IN1(n16679), .IN2(g2232), .Q(n17247) );
  AND2X1 U17828 ( .IN1(n17205), .IN2(n4287), .Q(n17246) );
  OR2X1 U17829 ( .IN1(n17248), .IN2(n17249), .Q(g22170) );
  AND2X1 U17830 ( .IN1(n17223), .IN2(g2206), .Q(n17249) );
  AND2X1 U17831 ( .IN1(n17224), .IN2(n4377), .Q(n17248) );
  OR2X1 U17832 ( .IN1(n17250), .IN2(n17251), .Q(g22169) );
  AND2X1 U17833 ( .IN1(n17231), .IN2(g1546), .Q(n17251) );
  AND2X1 U17834 ( .IN1(n17232), .IN2(n11936), .Q(n17250) );
  OR2X1 U17835 ( .IN1(n17252), .IN2(n17253), .Q(g22168) );
  AND2X1 U17836 ( .IN1(n16684), .IN2(g1541), .Q(n17253) );
  AND2X1 U17837 ( .IN1(n13311), .IN2(n17216), .Q(n17252) );
  OR2X1 U17838 ( .IN1(n17254), .IN2(n17255), .Q(g22167) );
  AND2X1 U17839 ( .IN1(n17256), .IN2(n4374), .Q(n17255) );
  AND2X1 U17840 ( .IN1(test_so52), .IN2(n17257), .Q(n17254) );
  OR2X1 U17841 ( .IN1(n17258), .IN2(n17259), .Q(g22166) );
  AND2X1 U17842 ( .IN1(n17231), .IN2(g1513), .Q(n17259) );
  AND2X1 U17843 ( .IN1(n17232), .IN2(n4378), .Q(n17258) );
  OR2X1 U17844 ( .IN1(n17260), .IN2(n17261), .Q(g22164) );
  AND2X1 U17845 ( .IN1(n16689), .IN2(g850), .Q(n17261) );
  AND2X1 U17846 ( .IN1(n17237), .IN2(n11983), .Q(n17260) );
  OR2X1 U17847 ( .IN1(n17262), .IN2(n17263), .Q(g22163) );
  AND2X1 U17848 ( .IN1(n17264), .IN2(g822), .Q(n17263) );
  AND2X1 U17849 ( .IN1(n17265), .IN2(n4375), .Q(n17262) );
  OR2X1 U17850 ( .IN1(n17266), .IN2(n17267), .Q(g22162) );
  AND2X1 U17851 ( .IN1(n16689), .IN2(g817), .Q(n17267) );
  AND2X1 U17852 ( .IN1(n4379), .IN2(n17237), .Q(n17266) );
  OR2X1 U17853 ( .IN1(n17268), .IN2(n17269), .Q(g22161) );
  AND2X1 U17854 ( .IN1(n16694), .IN2(g132), .Q(n17269) );
  AND2X1 U17855 ( .IN1(n17270), .IN2(n4376), .Q(n17268) );
  OR2X1 U17856 ( .IN1(n17271), .IN2(n17272), .Q(g22155) );
  AND2X1 U17857 ( .IN1(n17223), .IN2(g2236), .Q(n17272) );
  AND2X1 U17858 ( .IN1(n17224), .IN2(n13179), .Q(n17271) );
  INVX0 U17859 ( .INP(n12083), .ZN(n13179) );
  OR2X1 U17860 ( .IN1(n17273), .IN2(n17274), .Q(n12083) );
  OR2X1 U17861 ( .IN1(n17275), .IN2(n17276), .Q(n17274) );
  AND2X1 U17862 ( .IN1(n9758), .IN2(g2241), .Q(n17276) );
  AND2X1 U17863 ( .IN1(n9760), .IN2(g6837), .Q(n17275) );
  AND2X1 U17864 ( .IN1(n9759), .IN2(test_so73), .Q(n17273) );
  OR2X1 U17865 ( .IN1(n17277), .IN2(n17278), .Q(g22154) );
  AND2X1 U17866 ( .IN1(n17210), .IN2(g2234), .Q(n17278) );
  AND2X1 U17867 ( .IN1(n17211), .IN2(n4287), .Q(n17277) );
  OR2X1 U17868 ( .IN1(n17279), .IN2(n17280), .Q(g22153) );
  AND2X1 U17869 ( .IN1(n16679), .IN2(g2229), .Q(n17280) );
  AND2X1 U17870 ( .IN1(n17205), .IN2(n4563), .Q(n17279) );
  OR2X1 U17871 ( .IN1(n17281), .IN2(n17282), .Q(g22152) );
  AND2X1 U17872 ( .IN1(n17257), .IN2(g1545), .Q(n17282) );
  AND2X1 U17873 ( .IN1(n17256), .IN2(n11936), .Q(n17281) );
  INVX0 U17874 ( .INP(n13338), .ZN(n11936) );
  OR2X1 U17875 ( .IN1(n17283), .IN2(n17284), .Q(n13338) );
  OR2X1 U17876 ( .IN1(n17285), .IN2(n17286), .Q(n17284) );
  AND2X1 U17877 ( .IN1(g1547), .IN2(n10223), .Q(n17286) );
  AND2X1 U17878 ( .IN1(n9774), .IN2(g6573), .Q(n17285) );
  AND2X1 U17879 ( .IN1(n9773), .IN2(g6782), .Q(n17283) );
  OR2X1 U17880 ( .IN1(n17287), .IN2(n17288), .Q(g22151) );
  AND2X1 U17881 ( .IN1(n17231), .IN2(g1543), .Q(n17288) );
  AND2X1 U17882 ( .IN1(n17232), .IN2(n13311), .Q(n17287) );
  OR2X1 U17883 ( .IN1(n17289), .IN2(n17290), .Q(g22150) );
  AND2X1 U17884 ( .IN1(n16684), .IN2(g1538), .Q(n17290) );
  AND2X1 U17885 ( .IN1(n17216), .IN2(n4288), .Q(n17289) );
  OR2X1 U17886 ( .IN1(n17291), .IN2(n17292), .Q(g22149) );
  AND2X1 U17887 ( .IN1(n17257), .IN2(g1512), .Q(n17292) );
  AND2X1 U17888 ( .IN1(n17256), .IN2(n4378), .Q(n17291) );
  OR2X1 U17889 ( .IN1(n17293), .IN2(n17294), .Q(g22148) );
  AND2X1 U17890 ( .IN1(n17264), .IN2(g852), .Q(n17294) );
  AND2X1 U17891 ( .IN1(n17265), .IN2(n11983), .Q(n17293) );
  OR2X1 U17892 ( .IN1(n17295), .IN2(n17296), .Q(g22147) );
  AND2X1 U17893 ( .IN1(n16689), .IN2(g847), .Q(n17296) );
  AND2X1 U17894 ( .IN1(n13470), .IN2(n17237), .Q(n17295) );
  OR2X1 U17895 ( .IN1(n17297), .IN2(n17298), .Q(g22146) );
  AND2X1 U17896 ( .IN1(n17299), .IN2(g821), .Q(n17298) );
  AND2X1 U17897 ( .IN1(n17300), .IN2(n4375), .Q(n17297) );
  OR2X1 U17898 ( .IN1(n17301), .IN2(n17302), .Q(g22145) );
  AND2X1 U17899 ( .IN1(n17264), .IN2(g819), .Q(n17302) );
  AND2X1 U17900 ( .IN1(n17265), .IN2(n4379), .Q(n17301) );
  OR2X1 U17901 ( .IN1(n17303), .IN2(n17304), .Q(g22143) );
  AND2X1 U17902 ( .IN1(n16694), .IN2(g162), .Q(n17304) );
  AND2X1 U17903 ( .IN1(n17270), .IN2(n12036), .Q(n17303) );
  OR2X1 U17904 ( .IN1(n17305), .IN2(n17306), .Q(g22142) );
  AND2X1 U17905 ( .IN1(n17307), .IN2(g134), .Q(n17306) );
  AND2X1 U17906 ( .IN1(n17308), .IN2(n4376), .Q(n17305) );
  OR2X1 U17907 ( .IN1(n17309), .IN2(n17310), .Q(g22141) );
  AND2X1 U17908 ( .IN1(n16694), .IN2(g129), .Q(n17310) );
  AND2X1 U17909 ( .IN1(n4380), .IN2(n17270), .Q(n17309) );
  OR2X1 U17910 ( .IN1(n17311), .IN2(n17312), .Q(g22140) );
  AND2X1 U17911 ( .IN1(n17223), .IN2(g2233), .Q(n17312) );
  AND2X1 U17912 ( .IN1(n17224), .IN2(n4287), .Q(n17311) );
  OR2X1 U17913 ( .IN1(n17313), .IN2(n17314), .Q(g22139) );
  AND2X1 U17914 ( .IN1(n17210), .IN2(g2231), .Q(n17314) );
  AND2X1 U17915 ( .IN1(n17211), .IN2(n4563), .Q(n17313) );
  OR2X1 U17916 ( .IN1(n17315), .IN2(n17316), .Q(g22138) );
  AND2X1 U17917 ( .IN1(n16679), .IN2(g2226), .Q(n17316) );
  AND2X1 U17918 ( .IN1(n17205), .IN2(n4555), .Q(n17315) );
  OR2X1 U17919 ( .IN1(n17317), .IN2(n17318), .Q(g22132) );
  AND2X1 U17920 ( .IN1(n17257), .IN2(g1542), .Q(n17318) );
  AND2X1 U17921 ( .IN1(n17256), .IN2(n13311), .Q(n17317) );
  INVX0 U17922 ( .INP(n12135), .ZN(n13311) );
  OR2X1 U17923 ( .IN1(n17319), .IN2(n17320), .Q(n12135) );
  OR2X1 U17924 ( .IN1(n17321), .IN2(n17322), .Q(n17320) );
  AND2X1 U17925 ( .IN1(n9770), .IN2(g1547), .Q(n17322) );
  AND2X1 U17926 ( .IN1(n9772), .IN2(g6573), .Q(n17321) );
  AND2X1 U17927 ( .IN1(n9771), .IN2(g6782), .Q(n17319) );
  OR2X1 U17928 ( .IN1(n17323), .IN2(n17324), .Q(g22131) );
  AND2X1 U17929 ( .IN1(n17231), .IN2(g1540), .Q(n17324) );
  AND2X1 U17930 ( .IN1(n17232), .IN2(n4288), .Q(n17323) );
  OR2X1 U17931 ( .IN1(n17325), .IN2(n17326), .Q(g22130) );
  AND2X1 U17932 ( .IN1(n16684), .IN2(g1535), .Q(n17326) );
  AND2X1 U17933 ( .IN1(n17216), .IN2(n4565), .Q(n17325) );
  OR2X1 U17934 ( .IN1(n17327), .IN2(n17328), .Q(g22129) );
  AND2X1 U17935 ( .IN1(n17299), .IN2(g851), .Q(n17328) );
  AND2X1 U17936 ( .IN1(n17300), .IN2(n11983), .Q(n17327) );
  INVX0 U17937 ( .INP(n13440), .ZN(n11983) );
  OR2X1 U17938 ( .IN1(n17329), .IN2(n17330), .Q(n13440) );
  OR2X1 U17939 ( .IN1(n17331), .IN2(n17332), .Q(n17330) );
  AND2X1 U17940 ( .IN1(n9786), .IN2(g6368), .Q(n17332) );
  AND2X1 U17941 ( .IN1(n9785), .IN2(g6518), .Q(n17331) );
  AND2X1 U17942 ( .IN1(n9784), .IN2(test_so31), .Q(n17329) );
  OR2X1 U17943 ( .IN1(n17333), .IN2(n17334), .Q(g22128) );
  AND2X1 U17944 ( .IN1(n17264), .IN2(g849), .Q(n17334) );
  AND2X1 U17945 ( .IN1(n17265), .IN2(n13470), .Q(n17333) );
  OR2X1 U17946 ( .IN1(n17335), .IN2(n17336), .Q(g22127) );
  AND2X1 U17947 ( .IN1(n16689), .IN2(g844), .Q(n17336) );
  AND2X1 U17948 ( .IN1(n4289), .IN2(n17237), .Q(n17335) );
  OR2X1 U17949 ( .IN1(n17337), .IN2(n17338), .Q(g22126) );
  AND2X1 U17950 ( .IN1(n17299), .IN2(g818), .Q(n17338) );
  AND2X1 U17951 ( .IN1(n17300), .IN2(n4379), .Q(n17337) );
  OR2X1 U17952 ( .IN1(n17339), .IN2(n17340), .Q(g22125) );
  AND2X1 U17953 ( .IN1(n17307), .IN2(g164), .Q(n17340) );
  AND2X1 U17954 ( .IN1(n17308), .IN2(n12036), .Q(n17339) );
  OR2X1 U17955 ( .IN1(n17341), .IN2(n17342), .Q(g22124) );
  AND2X1 U17956 ( .IN1(n16694), .IN2(g159), .Q(n17342) );
  AND2X1 U17957 ( .IN1(n13567), .IN2(n17270), .Q(n17341) );
  OR2X1 U17958 ( .IN1(n17343), .IN2(n17344), .Q(g22123) );
  AND2X1 U17959 ( .IN1(n17345), .IN2(g133), .Q(n17344) );
  AND2X1 U17960 ( .IN1(n17346), .IN2(n4376), .Q(n17343) );
  OR2X1 U17961 ( .IN1(n17347), .IN2(n17348), .Q(g22122) );
  AND2X1 U17962 ( .IN1(n17307), .IN2(g131), .Q(n17348) );
  AND2X1 U17963 ( .IN1(n17308), .IN2(n4380), .Q(n17347) );
  OR2X1 U17964 ( .IN1(n17349), .IN2(n17350), .Q(g22117) );
  AND2X1 U17965 ( .IN1(n17223), .IN2(g2230), .Q(n17350) );
  AND2X1 U17966 ( .IN1(n17224), .IN2(n4563), .Q(n17349) );
  OR2X1 U17967 ( .IN1(n17351), .IN2(n17352), .Q(g22116) );
  AND2X1 U17968 ( .IN1(n17210), .IN2(g2228), .Q(n17352) );
  AND2X1 U17969 ( .IN1(n17211), .IN2(n4555), .Q(n17351) );
  OR2X1 U17970 ( .IN1(n17353), .IN2(n17354), .Q(g22115) );
  AND2X1 U17971 ( .IN1(n16679), .IN2(g2223), .Q(n17354) );
  AND2X1 U17972 ( .IN1(n17205), .IN2(n4325), .Q(n17353) );
  OR2X1 U17973 ( .IN1(n17355), .IN2(n17356), .Q(g22114) );
  AND2X1 U17974 ( .IN1(n17257), .IN2(g1539), .Q(n17356) );
  AND2X1 U17975 ( .IN1(n17256), .IN2(n4288), .Q(n17355) );
  OR2X1 U17976 ( .IN1(n17357), .IN2(n17358), .Q(g22113) );
  AND2X1 U17977 ( .IN1(n17232), .IN2(n4565), .Q(n17358) );
  AND2X1 U17978 ( .IN1(test_so53), .IN2(n17231), .Q(n17357) );
  OR2X1 U17979 ( .IN1(n17359), .IN2(n17360), .Q(g22112) );
  AND2X1 U17980 ( .IN1(n16684), .IN2(g1532), .Q(n17360) );
  AND2X1 U17981 ( .IN1(n17216), .IN2(n4557), .Q(n17359) );
  OR2X1 U17982 ( .IN1(n17361), .IN2(n17362), .Q(g22106) );
  AND2X1 U17983 ( .IN1(n17299), .IN2(g848), .Q(n17362) );
  AND2X1 U17984 ( .IN1(n17300), .IN2(n13470), .Q(n17361) );
  INVX0 U17985 ( .INP(n12190), .ZN(n13470) );
  OR2X1 U17986 ( .IN1(n17363), .IN2(n17364), .Q(n12190) );
  OR2X1 U17987 ( .IN1(n17365), .IN2(n17366), .Q(n17364) );
  AND2X1 U17988 ( .IN1(n9783), .IN2(g6368), .Q(n17366) );
  AND2X1 U17989 ( .IN1(n9782), .IN2(g6518), .Q(n17365) );
  AND2X1 U17990 ( .IN1(n9781), .IN2(test_so31), .Q(n17363) );
  OR2X1 U17991 ( .IN1(n17367), .IN2(n17368), .Q(g22105) );
  AND2X1 U17992 ( .IN1(n17264), .IN2(g846), .Q(n17368) );
  AND2X1 U17993 ( .IN1(n17265), .IN2(n4289), .Q(n17367) );
  OR2X1 U17994 ( .IN1(n17369), .IN2(n17370), .Q(g22104) );
  AND2X1 U17995 ( .IN1(n16689), .IN2(g841), .Q(n17370) );
  AND2X1 U17996 ( .IN1(n17237), .IN2(n4567), .Q(n17369) );
  OR2X1 U17997 ( .IN1(n17371), .IN2(n17372), .Q(g22103) );
  AND2X1 U17998 ( .IN1(n17346), .IN2(n12036), .Q(n17372) );
  INVX0 U17999 ( .INP(n13590), .ZN(n12036) );
  OR2X1 U18000 ( .IN1(n17373), .IN2(n17374), .Q(n13590) );
  OR2X1 U18001 ( .IN1(n17375), .IN2(n17376), .Q(n17374) );
  AND2X1 U18002 ( .IN1(n9795), .IN2(g165), .Q(n17376) );
  AND2X1 U18003 ( .IN1(n9797), .IN2(g6231), .Q(n17375) );
  AND2X1 U18004 ( .IN1(n9796), .IN2(g6313), .Q(n17373) );
  AND2X1 U18005 ( .IN1(test_so12), .IN2(n17345), .Q(n17371) );
  OR2X1 U18006 ( .IN1(n17377), .IN2(n17378), .Q(g22102) );
  AND2X1 U18007 ( .IN1(n17307), .IN2(g161), .Q(n17378) );
  AND2X1 U18008 ( .IN1(n17308), .IN2(n13567), .Q(n17377) );
  OR2X1 U18009 ( .IN1(n17379), .IN2(n17380), .Q(g22101) );
  AND2X1 U18010 ( .IN1(n16694), .IN2(g156), .Q(n17380) );
  AND2X1 U18011 ( .IN1(n4290), .IN2(n17270), .Q(n17379) );
  OR2X1 U18012 ( .IN1(n17381), .IN2(n17382), .Q(g22100) );
  AND2X1 U18013 ( .IN1(n17345), .IN2(g130), .Q(n17382) );
  AND2X1 U18014 ( .IN1(n17346), .IN2(n4380), .Q(n17381) );
  OR2X1 U18015 ( .IN1(n17383), .IN2(n17384), .Q(g22099) );
  AND2X1 U18016 ( .IN1(n17223), .IN2(g2227), .Q(n17384) );
  AND2X1 U18017 ( .IN1(n17224), .IN2(n4555), .Q(n17383) );
  OR2X1 U18018 ( .IN1(n17385), .IN2(n17386), .Q(g22098) );
  AND2X1 U18019 ( .IN1(n17211), .IN2(n4325), .Q(n17386) );
  AND2X1 U18020 ( .IN1(test_so74), .IN2(n17210), .Q(n17385) );
  OR2X1 U18021 ( .IN1(n17387), .IN2(n17388), .Q(g22097) );
  AND2X1 U18022 ( .IN1(n16679), .IN2(g2220), .Q(n17388) );
  AND2X1 U18023 ( .IN1(n17205), .IN2(n4389), .Q(n17387) );
  OR2X1 U18024 ( .IN1(n17389), .IN2(n17390), .Q(g22092) );
  AND2X1 U18025 ( .IN1(n17257), .IN2(g1536), .Q(n17390) );
  AND2X1 U18026 ( .IN1(n17256), .IN2(n4565), .Q(n17389) );
  OR2X1 U18027 ( .IN1(n17391), .IN2(n17392), .Q(g22091) );
  AND2X1 U18028 ( .IN1(n17231), .IN2(g1534), .Q(n17392) );
  AND2X1 U18029 ( .IN1(n17232), .IN2(n4557), .Q(n17391) );
  OR2X1 U18030 ( .IN1(n17393), .IN2(n17394), .Q(g22090) );
  AND2X1 U18031 ( .IN1(n16684), .IN2(g1529), .Q(n17394) );
  AND2X1 U18032 ( .IN1(n17216), .IN2(n4326), .Q(n17393) );
  OR2X1 U18033 ( .IN1(n17395), .IN2(n17396), .Q(g22089) );
  AND2X1 U18034 ( .IN1(n17299), .IN2(g845), .Q(n17396) );
  AND2X1 U18035 ( .IN1(n17300), .IN2(n4289), .Q(n17395) );
  OR2X1 U18036 ( .IN1(n17397), .IN2(n17398), .Q(g22088) );
  AND2X1 U18037 ( .IN1(n17264), .IN2(g843), .Q(n17398) );
  AND2X1 U18038 ( .IN1(n17265), .IN2(n4567), .Q(n17397) );
  OR2X1 U18039 ( .IN1(n17399), .IN2(n17400), .Q(g22087) );
  AND2X1 U18040 ( .IN1(n16689), .IN2(g838), .Q(n17400) );
  AND2X1 U18041 ( .IN1(n17237), .IN2(n4559), .Q(n17399) );
  OR2X1 U18042 ( .IN1(n17401), .IN2(n17402), .Q(g22081) );
  AND2X1 U18043 ( .IN1(n17345), .IN2(g160), .Q(n17402) );
  AND2X1 U18044 ( .IN1(n17346), .IN2(n13567), .Q(n17401) );
  INVX0 U18045 ( .INP(n12218), .ZN(n13567) );
  OR2X1 U18046 ( .IN1(n17403), .IN2(n17404), .Q(n12218) );
  OR2X1 U18047 ( .IN1(n17405), .IN2(n17406), .Q(n17404) );
  AND2X1 U18048 ( .IN1(n9792), .IN2(g165), .Q(n17406) );
  AND2X1 U18049 ( .IN1(n9794), .IN2(g6231), .Q(n17405) );
  AND2X1 U18050 ( .IN1(n9793), .IN2(g6313), .Q(n17403) );
  OR2X1 U18051 ( .IN1(n17407), .IN2(n17408), .Q(g22080) );
  AND2X1 U18052 ( .IN1(n17307), .IN2(g158), .Q(n17408) );
  AND2X1 U18053 ( .IN1(n17308), .IN2(n4290), .Q(n17407) );
  OR2X1 U18054 ( .IN1(n17409), .IN2(n17410), .Q(g22079) );
  AND2X1 U18055 ( .IN1(n16694), .IN2(g153), .Q(n17410) );
  AND2X1 U18056 ( .IN1(n17270), .IN2(n4569), .Q(n17409) );
  OR2X1 U18057 ( .IN1(n17411), .IN2(n17412), .Q(g22078) );
  AND2X1 U18058 ( .IN1(n17223), .IN2(g2224), .Q(n17412) );
  AND2X1 U18059 ( .IN1(n17224), .IN2(n4325), .Q(n17411) );
  OR2X1 U18060 ( .IN1(n17413), .IN2(n17414), .Q(g22077) );
  AND2X1 U18061 ( .IN1(n17210), .IN2(g2222), .Q(n17414) );
  AND2X1 U18062 ( .IN1(n17211), .IN2(n4389), .Q(n17413) );
  OR2X1 U18063 ( .IN1(n17415), .IN2(n17416), .Q(g22076) );
  AND2X1 U18064 ( .IN1(n16679), .IN2(g2217), .Q(n17416) );
  AND2X1 U18065 ( .IN1(n17205), .IN2(n4319), .Q(n17415) );
  INVX0 U18066 ( .INP(n16679), .ZN(n17205) );
  OR2X1 U18067 ( .IN1(n10162), .IN2(n4367), .Q(n16679) );
  OR2X1 U18068 ( .IN1(n17417), .IN2(n17418), .Q(g22075) );
  AND2X1 U18069 ( .IN1(n17257), .IN2(g1533), .Q(n17418) );
  AND2X1 U18070 ( .IN1(n17256), .IN2(n4557), .Q(n17417) );
  OR2X1 U18071 ( .IN1(n17419), .IN2(n17420), .Q(g22074) );
  AND2X1 U18072 ( .IN1(n17231), .IN2(g1531), .Q(n17420) );
  AND2X1 U18073 ( .IN1(n17232), .IN2(n4326), .Q(n17419) );
  OR2X1 U18074 ( .IN1(n17421), .IN2(n17422), .Q(g22073) );
  AND2X1 U18075 ( .IN1(n16684), .IN2(g1526), .Q(n17422) );
  AND2X1 U18076 ( .IN1(n17216), .IN2(n4390), .Q(n17421) );
  OR2X1 U18077 ( .IN1(n17423), .IN2(n17424), .Q(g22068) );
  AND2X1 U18078 ( .IN1(n17299), .IN2(g842), .Q(n17424) );
  AND2X1 U18079 ( .IN1(n17300), .IN2(n4567), .Q(n17423) );
  OR2X1 U18080 ( .IN1(n17425), .IN2(n17426), .Q(g22067) );
  AND2X1 U18081 ( .IN1(n17264), .IN2(g840), .Q(n17426) );
  AND2X1 U18082 ( .IN1(n17265), .IN2(n4559), .Q(n17425) );
  OR2X1 U18083 ( .IN1(n17427), .IN2(n17428), .Q(g22066) );
  AND2X1 U18084 ( .IN1(n16689), .IN2(g835), .Q(n17428) );
  AND2X1 U18085 ( .IN1(n4327), .IN2(n17237), .Q(n17427) );
  OR2X1 U18086 ( .IN1(n17429), .IN2(n17430), .Q(g22065) );
  AND2X1 U18087 ( .IN1(n17345), .IN2(g157), .Q(n17430) );
  AND2X1 U18088 ( .IN1(n17346), .IN2(n4290), .Q(n17429) );
  OR2X1 U18089 ( .IN1(n17431), .IN2(n17432), .Q(g22064) );
  AND2X1 U18090 ( .IN1(n17307), .IN2(g155), .Q(n17432) );
  AND2X1 U18091 ( .IN1(n17308), .IN2(n4569), .Q(n17431) );
  OR2X1 U18092 ( .IN1(n17433), .IN2(n17434), .Q(g22063) );
  AND2X1 U18093 ( .IN1(n16694), .IN2(g150), .Q(n17434) );
  AND2X1 U18094 ( .IN1(n17270), .IN2(n4561), .Q(n17433) );
  OR2X1 U18095 ( .IN1(n17435), .IN2(n17436), .Q(g22061) );
  AND2X1 U18096 ( .IN1(n17223), .IN2(g2221), .Q(n17436) );
  AND2X1 U18097 ( .IN1(n17224), .IN2(n4389), .Q(n17435) );
  OR2X1 U18098 ( .IN1(n17437), .IN2(n17438), .Q(g22060) );
  AND2X1 U18099 ( .IN1(n17210), .IN2(g2219), .Q(n17438) );
  AND2X1 U18100 ( .IN1(n17211), .IN2(n4319), .Q(n17437) );
  INVX0 U18101 ( .INP(n17210), .ZN(n17211) );
  OR2X1 U18102 ( .IN1(n10162), .IN2(n10189), .Q(n17210) );
  OR2X1 U18103 ( .IN1(n17439), .IN2(n17440), .Q(g22059) );
  AND2X1 U18104 ( .IN1(n17257), .IN2(g1530), .Q(n17440) );
  AND2X1 U18105 ( .IN1(n17256), .IN2(n4326), .Q(n17439) );
  OR2X1 U18106 ( .IN1(n17441), .IN2(n17442), .Q(g22058) );
  AND2X1 U18107 ( .IN1(n17231), .IN2(g1528), .Q(n17442) );
  AND2X1 U18108 ( .IN1(n17232), .IN2(n4390), .Q(n17441) );
  OR2X1 U18109 ( .IN1(n17443), .IN2(n17444), .Q(g22057) );
  AND2X1 U18110 ( .IN1(n16684), .IN2(g1523), .Q(n17444) );
  AND2X1 U18111 ( .IN1(n17216), .IN2(n4320), .Q(n17443) );
  INVX0 U18112 ( .INP(n16684), .ZN(n17216) );
  OR2X1 U18113 ( .IN1(n10161), .IN2(n4368), .Q(n16684) );
  OR2X1 U18114 ( .IN1(n17445), .IN2(n17446), .Q(g22056) );
  AND2X1 U18115 ( .IN1(n17300), .IN2(n4559), .Q(n17446) );
  AND2X1 U18116 ( .IN1(test_so32), .IN2(n17299), .Q(n17445) );
  OR2X1 U18117 ( .IN1(n17447), .IN2(n17448), .Q(g22055) );
  AND2X1 U18118 ( .IN1(n17264), .IN2(g837), .Q(n17448) );
  AND2X1 U18119 ( .IN1(n17265), .IN2(n4327), .Q(n17447) );
  OR2X1 U18120 ( .IN1(n17449), .IN2(n17450), .Q(g22054) );
  AND2X1 U18121 ( .IN1(n16689), .IN2(g832), .Q(n17450) );
  AND2X1 U18122 ( .IN1(n17237), .IN2(n4391), .Q(n17449) );
  OR2X1 U18123 ( .IN1(n17451), .IN2(n17452), .Q(g22049) );
  AND2X1 U18124 ( .IN1(n17345), .IN2(g154), .Q(n17452) );
  AND2X1 U18125 ( .IN1(n17346), .IN2(n4569), .Q(n17451) );
  OR2X1 U18126 ( .IN1(n17453), .IN2(n17454), .Q(g22048) );
  AND2X1 U18127 ( .IN1(n17307), .IN2(g152), .Q(n17454) );
  AND2X1 U18128 ( .IN1(n17308), .IN2(n4561), .Q(n17453) );
  OR2X1 U18129 ( .IN1(n17455), .IN2(n17456), .Q(g22047) );
  AND2X1 U18130 ( .IN1(n16694), .IN2(g147), .Q(n17456) );
  AND2X1 U18131 ( .IN1(n4328), .IN2(n17270), .Q(n17455) );
  OR2X1 U18132 ( .IN1(n17457), .IN2(n17458), .Q(g22045) );
  AND2X1 U18133 ( .IN1(n17223), .IN2(g2218), .Q(n17458) );
  AND2X1 U18134 ( .IN1(n17224), .IN2(n4319), .Q(n17457) );
  INVX0 U18135 ( .INP(n17223), .ZN(n17224) );
  OR2X1 U18136 ( .IN1(n10162), .IN2(n4324), .Q(n17223) );
  OR2X1 U18137 ( .IN1(n17459), .IN2(n17460), .Q(g22044) );
  AND2X1 U18138 ( .IN1(n17257), .IN2(g1527), .Q(n17460) );
  AND2X1 U18139 ( .IN1(n17256), .IN2(n4390), .Q(n17459) );
  OR2X1 U18140 ( .IN1(n17461), .IN2(n17462), .Q(g22043) );
  AND2X1 U18141 ( .IN1(n17231), .IN2(g1525), .Q(n17462) );
  AND2X1 U18142 ( .IN1(n17232), .IN2(n4320), .Q(n17461) );
  INVX0 U18143 ( .INP(n17231), .ZN(n17232) );
  OR2X1 U18144 ( .IN1(n10161), .IN2(n4515), .Q(n17231) );
  OR2X1 U18145 ( .IN1(n17463), .IN2(n17464), .Q(g22042) );
  AND2X1 U18146 ( .IN1(n17299), .IN2(g836), .Q(n17464) );
  AND2X1 U18147 ( .IN1(n17300), .IN2(n4327), .Q(n17463) );
  OR2X1 U18148 ( .IN1(n17465), .IN2(n17466), .Q(g22041) );
  AND2X1 U18149 ( .IN1(n17264), .IN2(g834), .Q(n17466) );
  AND2X1 U18150 ( .IN1(n17265), .IN2(n4391), .Q(n17465) );
  OR2X1 U18151 ( .IN1(n17467), .IN2(n17468), .Q(g22040) );
  AND2X1 U18152 ( .IN1(n16689), .IN2(g829), .Q(n17468) );
  AND2X1 U18153 ( .IN1(n4321), .IN2(n17237), .Q(n17467) );
  INVX0 U18154 ( .INP(n16689), .ZN(n17237) );
  OR2X1 U18155 ( .IN1(n10160), .IN2(n10188), .Q(n16689) );
  OR2X1 U18156 ( .IN1(n17469), .IN2(n17470), .Q(g22039) );
  AND2X1 U18157 ( .IN1(n17345), .IN2(g151), .Q(n17470) );
  AND2X1 U18158 ( .IN1(n17346), .IN2(n4561), .Q(n17469) );
  OR2X1 U18159 ( .IN1(n17471), .IN2(n17472), .Q(g22038) );
  AND2X1 U18160 ( .IN1(n17307), .IN2(g149), .Q(n17472) );
  AND2X1 U18161 ( .IN1(n17308), .IN2(n4328), .Q(n17471) );
  OR2X1 U18162 ( .IN1(n17473), .IN2(n17474), .Q(g22037) );
  AND2X1 U18163 ( .IN1(n17270), .IN2(n4392), .Q(n17474) );
  AND2X1 U18164 ( .IN1(test_so11), .IN2(n16694), .Q(n17473) );
  OR2X1 U18165 ( .IN1(n17475), .IN2(n17476), .Q(g22035) );
  AND2X1 U18166 ( .IN1(n17257), .IN2(g1524), .Q(n17476) );
  AND2X1 U18167 ( .IN1(n17256), .IN2(n4320), .Q(n17475) );
  INVX0 U18168 ( .INP(n17257), .ZN(n17256) );
  OR2X1 U18169 ( .IN1(n10161), .IN2(n4317), .Q(n17257) );
  OR2X1 U18170 ( .IN1(n17477), .IN2(n17478), .Q(g22034) );
  AND2X1 U18171 ( .IN1(n17299), .IN2(g833), .Q(n17478) );
  AND2X1 U18172 ( .IN1(n17300), .IN2(n4391), .Q(n17477) );
  OR2X1 U18173 ( .IN1(n17479), .IN2(n17480), .Q(g22033) );
  AND2X1 U18174 ( .IN1(n17264), .IN2(g831), .Q(n17480) );
  AND2X1 U18175 ( .IN1(n17265), .IN2(n4321), .Q(n17479) );
  INVX0 U18176 ( .INP(n17264), .ZN(n17265) );
  OR2X1 U18177 ( .IN1(n10160), .IN2(n4312), .Q(n17264) );
  OR2X1 U18178 ( .IN1(n17481), .IN2(n17482), .Q(g22032) );
  AND2X1 U18179 ( .IN1(n17345), .IN2(g148), .Q(n17482) );
  AND2X1 U18180 ( .IN1(n17346), .IN2(n4328), .Q(n17481) );
  OR2X1 U18181 ( .IN1(n17483), .IN2(n17484), .Q(g22031) );
  AND2X1 U18182 ( .IN1(n17307), .IN2(g146), .Q(n17484) );
  AND2X1 U18183 ( .IN1(n17308), .IN2(n4392), .Q(n17483) );
  OR2X1 U18184 ( .IN1(n17485), .IN2(n17486), .Q(g22030) );
  AND2X1 U18185 ( .IN1(n16694), .IN2(g141), .Q(n17486) );
  AND2X1 U18186 ( .IN1(n4322), .IN2(n17270), .Q(n17485) );
  INVX0 U18187 ( .INP(n16694), .ZN(n17270) );
  OR2X1 U18188 ( .IN1(n10159), .IN2(n4369), .Q(n16694) );
  OR2X1 U18189 ( .IN1(n17487), .IN2(n17488), .Q(g22029) );
  AND2X1 U18190 ( .IN1(n17299), .IN2(g830), .Q(n17488) );
  AND2X1 U18191 ( .IN1(n17300), .IN2(n4321), .Q(n17487) );
  INVX0 U18192 ( .INP(n17299), .ZN(n17300) );
  OR2X1 U18193 ( .IN1(n10160), .IN2(n4323), .Q(n17299) );
  OR2X1 U18194 ( .IN1(n17489), .IN2(n17490), .Q(g22028) );
  AND2X1 U18195 ( .IN1(n17345), .IN2(g145), .Q(n17490) );
  AND2X1 U18196 ( .IN1(n17346), .IN2(n4392), .Q(n17489) );
  OR2X1 U18197 ( .IN1(n17491), .IN2(n17492), .Q(g22027) );
  AND2X1 U18198 ( .IN1(n17307), .IN2(g143), .Q(n17492) );
  AND2X1 U18199 ( .IN1(n17308), .IN2(n4322), .Q(n17491) );
  INVX0 U18200 ( .INP(n17307), .ZN(n17308) );
  OR2X1 U18201 ( .IN1(n10159), .IN2(n4512), .Q(n17307) );
  AND2X1 U18202 ( .IN1(n17493), .IN2(n11730), .Q(g22026) );
  AND2X1 U18203 ( .IN1(n10877), .IN2(n18258), .Q(n11730) );
  OR2X1 U18204 ( .IN1(n17494), .IN2(n17495), .Q(n10877) );
  OR2X1 U18205 ( .IN1(n17496), .IN2(g2883), .Q(n17495) );
  INVX0 U18206 ( .INP(n17497), .ZN(n17496) );
  AND2X1 U18207 ( .IN1(n4182), .IN2(n4431), .Q(n17497) );
  OR2X1 U18208 ( .IN1(n17498), .IN2(n17499), .Q(n17494) );
  OR2X1 U18209 ( .IN1(n10152), .IN2(g2900), .Q(n17499) );
  OR2X1 U18210 ( .IN1(n4423), .IN2(n4355), .Q(n17498) );
  AND2X1 U18211 ( .IN1(n17500), .IN2(n4123), .Q(n17493) );
  OR2X1 U18212 ( .IN1(n10152), .IN2(n17501), .Q(n4123) );
  OR2X1 U18213 ( .IN1(n4423), .IN2(n4330), .Q(n17501) );
  OR2X1 U18214 ( .IN1(n17502), .IN2(g2888), .Q(n17500) );
  AND2X1 U18215 ( .IN1(g2883), .IN2(g2950), .Q(n17502) );
  OR2X1 U18216 ( .IN1(n17503), .IN2(n17504), .Q(g22025) );
  AND2X1 U18217 ( .IN1(n17345), .IN2(g142), .Q(n17504) );
  AND2X1 U18218 ( .IN1(n17346), .IN2(n4322), .Q(n17503) );
  INVX0 U18219 ( .INP(n17345), .ZN(n17346) );
  OR2X1 U18220 ( .IN1(n10159), .IN2(n4318), .Q(n17345) );
  AND2X1 U18221 ( .IN1(n17505), .IN2(n17506), .Q(g21974) );
  OR2X1 U18222 ( .IN1(n17507), .IN2(g2707), .Q(n17506) );
  INVX0 U18223 ( .INP(n17508), .ZN(n17507) );
  AND2X1 U18224 ( .IN1(n16869), .IN2(n14331), .Q(n17505) );
  OR2X1 U18225 ( .IN1(n4472), .IN2(n17508), .Q(n16869) );
  AND2X1 U18226 ( .IN1(n17509), .IN2(n17510), .Q(g21972) );
  OR2X1 U18227 ( .IN1(n17511), .IN2(g2013), .Q(n17510) );
  INVX0 U18228 ( .INP(n17512), .ZN(n17511) );
  AND2X1 U18229 ( .IN1(n16875), .IN2(n14337), .Q(n17509) );
  OR2X1 U18230 ( .IN1(n4474), .IN2(n17512), .Q(n16875) );
  OR2X1 U18231 ( .IN1(n17513), .IN2(n17514), .Q(g21970) );
  AND2X1 U18232 ( .IN1(n15191), .IN2(g2560), .Q(n17514) );
  OR2X1 U18233 ( .IN1(n17515), .IN2(n17516), .Q(n15191) );
  OR2X1 U18234 ( .IN1(n17517), .IN2(n17518), .Q(n17516) );
  AND2X1 U18235 ( .IN1(g7264), .IN2(g2516), .Q(n17518) );
  AND2X1 U18236 ( .IN1(n4606), .IN2(g2519), .Q(n17517) );
  AND2X1 U18237 ( .IN1(g5555), .IN2(g2513), .Q(n17515) );
  AND2X1 U18238 ( .IN1(test_so87), .IN2(n4463), .Q(n17513) );
  AND2X1 U18239 ( .IN1(n17519), .IN2(n17520), .Q(g21969) );
  OR2X1 U18240 ( .IN1(n17521), .IN2(g1319), .Q(n17520) );
  INVX0 U18241 ( .INP(n17522), .ZN(n17521) );
  AND2X1 U18242 ( .IN1(n16881), .IN2(n14345), .Q(n17519) );
  OR2X1 U18243 ( .IN1(n4476), .IN2(n17522), .Q(n16881) );
  OR2X1 U18244 ( .IN1(n17523), .IN2(n17524), .Q(g21882) );
  AND2X1 U18245 ( .IN1(n17525), .IN2(g2879), .Q(n17524) );
  AND2X1 U18246 ( .IN1(n4351), .IN2(g2878), .Q(n17523) );
  OR2X1 U18247 ( .IN1(n17526), .IN2(n17527), .Q(g21880) );
  AND2X1 U18248 ( .IN1(n17528), .IN2(g2879), .Q(n17527) );
  AND2X1 U18249 ( .IN1(n4351), .IN2(g2877), .Q(n17526) );
  OR2X1 U18250 ( .IN1(n17529), .IN2(n17530), .Q(g21878) );
  AND2X1 U18251 ( .IN1(n4351), .IN2(n17525), .Q(n17530) );
  OR2X1 U18252 ( .IN1(n17531), .IN2(n17532), .Q(n17525) );
  INVX0 U18253 ( .INP(n17533), .ZN(n17532) );
  OR2X1 U18254 ( .IN1(n10608), .IN2(n17534), .Q(n17533) );
  AND2X1 U18255 ( .IN1(n17534), .IN2(n10608), .Q(n17531) );
  AND2X1 U18256 ( .IN1(n17535), .IN2(n17536), .Q(n10608) );
  INVX0 U18257 ( .INP(n17537), .ZN(n17536) );
  AND2X1 U18258 ( .IN1(n17538), .IN2(n17539), .Q(n17537) );
  OR2X1 U18259 ( .IN1(n17539), .IN2(n17538), .Q(n17535) );
  OR2X1 U18260 ( .IN1(n17540), .IN2(n17541), .Q(n17538) );
  AND2X1 U18261 ( .IN1(n17542), .IN2(n17543), .Q(n17541) );
  INVX0 U18262 ( .INP(n17544), .ZN(n17540) );
  OR2X1 U18263 ( .IN1(n17543), .IN2(n17542), .Q(n17544) );
  OR2X1 U18264 ( .IN1(n17545), .IN2(n17546), .Q(n17542) );
  AND2X1 U18265 ( .IN1(n10137), .IN2(g2874), .Q(n17546) );
  AND2X1 U18266 ( .IN1(n10138), .IN2(g2978), .Q(n17545) );
  INVX0 U18267 ( .INP(n17547), .ZN(n17543) );
  OR2X1 U18268 ( .IN1(n17548), .IN2(n17549), .Q(n17547) );
  AND2X1 U18269 ( .IN1(n10139), .IN2(g2972), .Q(n17549) );
  AND2X1 U18270 ( .IN1(n10140), .IN2(g2963), .Q(n17548) );
  AND2X1 U18271 ( .IN1(n17550), .IN2(n17551), .Q(n17539) );
  INVX0 U18272 ( .INP(n17552), .ZN(n17551) );
  AND2X1 U18273 ( .IN1(n17553), .IN2(n17554), .Q(n17552) );
  OR2X1 U18274 ( .IN1(n17554), .IN2(n17553), .Q(n17550) );
  OR2X1 U18275 ( .IN1(n17555), .IN2(n17556), .Q(n17553) );
  AND2X1 U18276 ( .IN1(n10141), .IN2(g2969), .Q(n17556) );
  AND2X1 U18277 ( .IN1(n10142), .IN2(g2975), .Q(n17555) );
  AND2X1 U18278 ( .IN1(n17557), .IN2(n17558), .Q(n17554) );
  OR2X1 U18279 ( .IN1(g2981), .IN2(test_so2), .Q(n17558) );
  OR2X1 U18280 ( .IN1(n10198), .IN2(n10143), .Q(n17557) );
  AND2X1 U18281 ( .IN1(test_so4), .IN2(g2879), .Q(n17529) );
  OR2X1 U18282 ( .IN1(n17559), .IN2(n17560), .Q(g21851) );
  AND2X1 U18283 ( .IN1(n17561), .IN2(n4541), .Q(n17560) );
  AND2X1 U18284 ( .IN1(n4298), .IN2(g548), .Q(n17561) );
  AND2X1 U18285 ( .IN1(g499), .IN2(g544), .Q(n17559) );
  OR2X1 U18286 ( .IN1(n17562), .IN2(n16704), .Q(g21847) );
  AND2X1 U18287 ( .IN1(g2624), .IN2(n13858), .Q(n16704) );
  AND2X1 U18288 ( .IN1(n4299), .IN2(g2628), .Q(n17562) );
  OR2X1 U18289 ( .IN1(n17563), .IN2(n16712), .Q(g21845) );
  AND2X1 U18290 ( .IN1(g1930), .IN2(n13858), .Q(n16712) );
  AND2X1 U18291 ( .IN1(n4366), .IN2(g1934), .Q(n17563) );
  OR2X1 U18292 ( .IN1(n17564), .IN2(n16736), .Q(g21843) );
  AND2X1 U18293 ( .IN1(g1236), .IN2(n13858), .Q(n16736) );
  AND2X1 U18294 ( .IN1(n4300), .IN2(g1240), .Q(n17564) );
  OR2X1 U18295 ( .IN1(n17565), .IN2(n16773), .Q(g21842) );
  AND2X1 U18296 ( .IN1(g550), .IN2(n13858), .Q(n16773) );
  INVX0 U18297 ( .INP(n13859), .ZN(n13858) );
  AND2X1 U18298 ( .IN1(n17566), .IN2(n17567), .Q(n13859) );
  AND2X1 U18299 ( .IN1(n4480), .IN2(n10157), .Q(n17567) );
  AND2X1 U18300 ( .IN1(n17057), .IN2(n17568), .Q(n17566) );
  INVX0 U18301 ( .INP(n17569), .ZN(n17568) );
  OR2X1 U18302 ( .IN1(n4481), .IN2(n4350), .Q(n17569) );
  INVX0 U18303 ( .INP(n17039), .ZN(n17057) );
  OR2X1 U18304 ( .IN1(n17570), .IN2(n17571), .Q(n17039) );
  OR2X1 U18305 ( .IN1(g2993), .IN2(n17572), .Q(n17571) );
  OR2X1 U18306 ( .IN1(n10163), .IN2(g3006), .Q(n17572) );
  OR2X1 U18307 ( .IN1(n17573), .IN2(n17574), .Q(n17570) );
  OR2X1 U18308 ( .IN1(n9352), .IN2(n9351), .Q(n17574) );
  OR2X1 U18309 ( .IN1(test_so98), .IN2(n18262), .Q(n17573) );
  AND2X1 U18310 ( .IN1(n4313), .IN2(g554), .Q(n17565) );
  OR2X1 U18311 ( .IN1(n17575), .IN2(n17576), .Q(g21346) );
  INVX0 U18312 ( .INP(n17577), .ZN(n17576) );
  OR2X1 U18313 ( .IN1(n17578), .IN2(n18263), .Q(n17577) );
  OR2X1 U18314 ( .IN1(g6447), .IN2(n9616), .Q(n17578) );
  AND2X1 U18315 ( .IN1(n18263), .IN2(DFF_328_n1), .Q(n17575) );
  OR2X1 U18316 ( .IN1(n17579), .IN2(n17580), .Q(g21094) );
  AND2X1 U18317 ( .IN1(n16067), .IN2(n4393), .Q(n17580) );
  AND2X1 U18318 ( .IN1(test_so94), .IN2(n16068), .Q(n17579) );
  OR2X1 U18319 ( .IN1(n17581), .IN2(n17582), .Q(g21082) );
  AND2X1 U18320 ( .IN1(n16071), .IN2(g2798), .Q(n17582) );
  AND2X1 U18321 ( .IN1(n16072), .IN2(n4393), .Q(n17581) );
  OR2X1 U18322 ( .IN1(n17583), .IN2(n17584), .Q(g21081) );
  AND2X1 U18323 ( .IN1(n16068), .IN2(g2793), .Q(n17584) );
  AND2X1 U18324 ( .IN1(n16067), .IN2(n4471), .Q(n17583) );
  OR2X1 U18325 ( .IN1(n17585), .IN2(n17586), .Q(g21080) );
  AND2X1 U18326 ( .IN1(n16076), .IN2(g2102), .Q(n17586) );
  AND2X1 U18327 ( .IN1(n4149), .IN2(n10194), .Q(n17585) );
  OR2X1 U18328 ( .IN1(n17587), .IN2(n17588), .Q(g21075) );
  AND2X1 U18329 ( .IN1(n16079), .IN2(g2797), .Q(n17588) );
  AND2X1 U18330 ( .IN1(n16080), .IN2(n4393), .Q(n17587) );
  OR2X1 U18331 ( .IN1(n17589), .IN2(n17590), .Q(g21074) );
  AND2X1 U18332 ( .IN1(n16071), .IN2(g2795), .Q(n17590) );
  AND2X1 U18333 ( .IN1(n16072), .IN2(n4471), .Q(n17589) );
  OR2X1 U18334 ( .IN1(n17591), .IN2(n17592), .Q(g21073) );
  AND2X1 U18335 ( .IN1(n16068), .IN2(g2790), .Q(n17592) );
  AND2X1 U18336 ( .IN1(n16067), .IN2(n10192), .Q(n17591) );
  OR2X1 U18337 ( .IN1(n17593), .IN2(n17594), .Q(g21072) );
  AND2X1 U18338 ( .IN1(n16176), .IN2(g2104), .Q(n17594) );
  AND2X1 U18339 ( .IN1(n16175), .IN2(n10194), .Q(n17593) );
  OR2X1 U18340 ( .IN1(n17595), .IN2(n17596), .Q(g21071) );
  AND2X1 U18341 ( .IN1(n16076), .IN2(g2099), .Q(n17596) );
  AND2X1 U18342 ( .IN1(n4149), .IN2(n4473), .Q(n17595) );
  OR2X1 U18343 ( .IN1(n17597), .IN2(n17598), .Q(g21070) );
  AND2X1 U18344 ( .IN1(n16181), .IN2(g1408), .Q(n17598) );
  AND2X1 U18345 ( .IN1(n16180), .IN2(n4395), .Q(n17597) );
  OR2X1 U18346 ( .IN1(n17599), .IN2(n17600), .Q(g21063) );
  AND2X1 U18347 ( .IN1(n17184), .IN2(g2805), .Q(n17600) );
  AND2X1 U18348 ( .IN1(n17601), .IN2(n11213), .Q(n17599) );
  OR2X1 U18349 ( .IN1(n17602), .IN2(n17603), .Q(g21062) );
  AND2X1 U18350 ( .IN1(n16079), .IN2(g2794), .Q(n17603) );
  AND2X1 U18351 ( .IN1(n16080), .IN2(n4471), .Q(n17602) );
  OR2X1 U18352 ( .IN1(n17604), .IN2(n17605), .Q(g21061) );
  AND2X1 U18353 ( .IN1(n16071), .IN2(g2792), .Q(n17605) );
  AND2X1 U18354 ( .IN1(n16072), .IN2(n10192), .Q(n17604) );
  OR2X1 U18355 ( .IN1(n17606), .IN2(n17607), .Q(g21060) );
  AND2X1 U18356 ( .IN1(n16068), .IN2(g2787), .Q(n17607) );
  AND2X1 U18357 ( .IN1(n16067), .IN2(n4407), .Q(n17606) );
  OR2X1 U18358 ( .IN1(n17608), .IN2(n17609), .Q(g21056) );
  AND2X1 U18359 ( .IN1(n16277), .IN2(g2103), .Q(n17609) );
  AND2X1 U18360 ( .IN1(n16184), .IN2(n10194), .Q(n17608) );
  OR2X1 U18361 ( .IN1(n17610), .IN2(n17611), .Q(g21055) );
  AND2X1 U18362 ( .IN1(n16176), .IN2(g2101), .Q(n17611) );
  AND2X1 U18363 ( .IN1(n16175), .IN2(n4473), .Q(n17610) );
  OR2X1 U18364 ( .IN1(n17612), .IN2(n17613), .Q(g21054) );
  AND2X1 U18365 ( .IN1(n16076), .IN2(g2096), .Q(n17613) );
  AND2X1 U18366 ( .IN1(n4149), .IN2(n4468), .Q(n17612) );
  OR2X1 U18367 ( .IN1(n17614), .IN2(n17615), .Q(g21053) );
  AND2X1 U18368 ( .IN1(n16280), .IN2(g1410), .Q(n17615) );
  AND2X1 U18369 ( .IN1(n1027), .IN2(n4395), .Q(n17614) );
  OR2X1 U18370 ( .IN1(n17616), .IN2(n17617), .Q(g21052) );
  AND2X1 U18371 ( .IN1(n16181), .IN2(g1405), .Q(n17617) );
  AND2X1 U18372 ( .IN1(n16180), .IN2(n4475), .Q(n17616) );
  OR2X1 U18373 ( .IN1(n17618), .IN2(n17619), .Q(g21051) );
  AND2X1 U18374 ( .IN1(n16284), .IN2(g722), .Q(n17619) );
  AND2X1 U18375 ( .IN1(n680), .IN2(n4396), .Q(n17618) );
  OR2X1 U18376 ( .IN1(n17620), .IN2(n17621), .Q(g21047) );
  AND2X1 U18377 ( .IN1(n14331), .IN2(g2807), .Q(n17621) );
  AND2X1 U18378 ( .IN1(n17622), .IN2(n11213), .Q(n17620) );
  OR2X1 U18379 ( .IN1(n17623), .IN2(n17624), .Q(g21046) );
  AND2X1 U18380 ( .IN1(n17184), .IN2(g2802), .Q(n17624) );
  AND2X1 U18381 ( .IN1(n17601), .IN2(n11222), .Q(n17623) );
  INVX0 U18382 ( .INP(n17184), .ZN(n17601) );
  OR2X1 U18383 ( .IN1(n10156), .IN2(n4292), .Q(n17184) );
  OR2X1 U18384 ( .IN1(n17625), .IN2(n17626), .Q(g21045) );
  AND2X1 U18385 ( .IN1(n16079), .IN2(g2791), .Q(n17626) );
  AND2X1 U18386 ( .IN1(n16080), .IN2(n10192), .Q(n17625) );
  OR2X1 U18387 ( .IN1(n17627), .IN2(n17628), .Q(g21044) );
  AND2X1 U18388 ( .IN1(n16071), .IN2(g2789), .Q(n17628) );
  AND2X1 U18389 ( .IN1(n16072), .IN2(n4407), .Q(n17627) );
  OR2X1 U18390 ( .IN1(n17629), .IN2(n17630), .Q(g21043) );
  AND2X1 U18391 ( .IN1(n16068), .IN2(g2784), .Q(n17630) );
  AND2X1 U18392 ( .IN1(n16067), .IN2(n4397), .Q(n17629) );
  OR2X1 U18393 ( .IN1(n17631), .IN2(n17632), .Q(g21042) );
  AND2X1 U18394 ( .IN1(n17187), .IN2(g2111), .Q(n17632) );
  AND2X1 U18395 ( .IN1(n17633), .IN2(n11375), .Q(n17631) );
  OR2X1 U18396 ( .IN1(n17634), .IN2(n17635), .Q(g21041) );
  AND2X1 U18397 ( .IN1(n16277), .IN2(g2100), .Q(n17635) );
  AND2X1 U18398 ( .IN1(n16184), .IN2(n4473), .Q(n17634) );
  OR2X1 U18399 ( .IN1(n17636), .IN2(n17637), .Q(g21040) );
  AND2X1 U18400 ( .IN1(n16176), .IN2(g2098), .Q(n17637) );
  AND2X1 U18401 ( .IN1(n16175), .IN2(n4468), .Q(n17636) );
  OR2X1 U18402 ( .IN1(n17638), .IN2(n17639), .Q(g21039) );
  AND2X1 U18403 ( .IN1(n16076), .IN2(g2093), .Q(n17639) );
  AND2X1 U18404 ( .IN1(n4149), .IN2(n4409), .Q(n17638) );
  OR2X1 U18405 ( .IN1(n17640), .IN2(n17641), .Q(g21035) );
  AND2X1 U18406 ( .IN1(n16292), .IN2(g1409), .Q(n17641) );
  AND2X1 U18407 ( .IN1(n16293), .IN2(n4395), .Q(n17640) );
  OR2X1 U18408 ( .IN1(n17642), .IN2(n17643), .Q(g21034) );
  AND2X1 U18409 ( .IN1(n16280), .IN2(g1407), .Q(n17643) );
  AND2X1 U18410 ( .IN1(n1027), .IN2(n4475), .Q(n17642) );
  OR2X1 U18411 ( .IN1(n17644), .IN2(n17645), .Q(g21033) );
  AND2X1 U18412 ( .IN1(n16181), .IN2(g1402), .Q(n17645) );
  AND2X1 U18413 ( .IN1(n16180), .IN2(n4469), .Q(n17644) );
  OR2X1 U18414 ( .IN1(n17646), .IN2(n17647), .Q(g21032) );
  AND2X1 U18415 ( .IN1(n16387), .IN2(g724), .Q(n17647) );
  AND2X1 U18416 ( .IN1(n16388), .IN2(n4396), .Q(n17646) );
  OR2X1 U18417 ( .IN1(n17648), .IN2(n17649), .Q(g21031) );
  AND2X1 U18418 ( .IN1(n16284), .IN2(g719), .Q(n17649) );
  AND2X1 U18419 ( .IN1(n680), .IN2(n4477), .Q(n17648) );
  OR2X1 U18420 ( .IN1(n17650), .IN2(n17651), .Q(g21029) );
  AND2X1 U18421 ( .IN1(n17189), .IN2(g2806), .Q(n17651) );
  AND2X1 U18422 ( .IN1(n17652), .IN2(n11213), .Q(n17650) );
  INVX0 U18423 ( .INP(n11136), .ZN(n11213) );
  OR2X1 U18424 ( .IN1(n17653), .IN2(n17654), .Q(n11136) );
  OR2X1 U18425 ( .IN1(n17655), .IN2(n17656), .Q(n17654) );
  AND2X1 U18426 ( .IN1(g2624), .IN2(g2685), .Q(n17656) );
  AND2X1 U18427 ( .IN1(g7302), .IN2(g2679), .Q(n17655) );
  AND2X1 U18428 ( .IN1(test_so90), .IN2(g7390), .Q(n17653) );
  OR2X1 U18429 ( .IN1(n17657), .IN2(n17658), .Q(g21028) );
  AND2X1 U18430 ( .IN1(n14331), .IN2(g2804), .Q(n17658) );
  AND2X1 U18431 ( .IN1(n17622), .IN2(n11222), .Q(n17657) );
  INVX0 U18432 ( .INP(n14331), .ZN(n17622) );
  OR2X1 U18433 ( .IN1(n17659), .IN2(n17660), .Q(g21027) );
  AND2X1 U18434 ( .IN1(n16079), .IN2(g2788), .Q(n17660) );
  AND2X1 U18435 ( .IN1(n16080), .IN2(n4407), .Q(n17659) );
  OR2X1 U18436 ( .IN1(n17661), .IN2(n17662), .Q(g21026) );
  AND2X1 U18437 ( .IN1(n16071), .IN2(g2786), .Q(n17662) );
  AND2X1 U18438 ( .IN1(n16072), .IN2(n4397), .Q(n17661) );
  OR2X1 U18439 ( .IN1(n17663), .IN2(n17664), .Q(g21025) );
  AND2X1 U18440 ( .IN1(n16067), .IN2(n4408), .Q(n17664) );
  AND2X1 U18441 ( .IN1(test_so93), .IN2(n16068), .Q(n17663) );
  OR2X1 U18442 ( .IN1(n17665), .IN2(n17666), .Q(g21023) );
  AND2X1 U18443 ( .IN1(n14337), .IN2(g2113), .Q(n17666) );
  AND2X1 U18444 ( .IN1(n17667), .IN2(n11375), .Q(n17665) );
  OR2X1 U18445 ( .IN1(n17668), .IN2(n17669), .Q(g21022) );
  AND2X1 U18446 ( .IN1(n17187), .IN2(g2108), .Q(n17669) );
  AND2X1 U18447 ( .IN1(n17633), .IN2(n11383), .Q(n17668) );
  INVX0 U18448 ( .INP(n17187), .ZN(n17633) );
  OR2X1 U18449 ( .IN1(n10155), .IN2(n4293), .Q(n17187) );
  OR2X1 U18450 ( .IN1(n17670), .IN2(n17671), .Q(g21021) );
  AND2X1 U18451 ( .IN1(n16277), .IN2(g2097), .Q(n17671) );
  AND2X1 U18452 ( .IN1(n16184), .IN2(n4468), .Q(n17670) );
  OR2X1 U18453 ( .IN1(n17672), .IN2(n17673), .Q(g21020) );
  AND2X1 U18454 ( .IN1(n16176), .IN2(g2095), .Q(n17673) );
  AND2X1 U18455 ( .IN1(n16175), .IN2(n4409), .Q(n17672) );
  OR2X1 U18456 ( .IN1(n17674), .IN2(n17675), .Q(g21019) );
  AND2X1 U18457 ( .IN1(n16076), .IN2(g2090), .Q(n17675) );
  AND2X1 U18458 ( .IN1(n4149), .IN2(n4399), .Q(n17674) );
  OR2X1 U18459 ( .IN1(n17676), .IN2(n17677), .Q(g21018) );
  AND2X1 U18460 ( .IN1(n17192), .IN2(g1417), .Q(n17677) );
  AND2X1 U18461 ( .IN1(n17678), .IN2(n11538), .Q(n17676) );
  OR2X1 U18462 ( .IN1(n17679), .IN2(n17680), .Q(g21017) );
  AND2X1 U18463 ( .IN1(n16292), .IN2(g1406), .Q(n17680) );
  AND2X1 U18464 ( .IN1(n16293), .IN2(n4475), .Q(n17679) );
  OR2X1 U18465 ( .IN1(n17681), .IN2(n17682), .Q(g21016) );
  AND2X1 U18466 ( .IN1(n16280), .IN2(g1404), .Q(n17682) );
  AND2X1 U18467 ( .IN1(n1027), .IN2(n4469), .Q(n17681) );
  OR2X1 U18468 ( .IN1(n17683), .IN2(n17684), .Q(g21015) );
  AND2X1 U18469 ( .IN1(n16181), .IN2(g1399), .Q(n17684) );
  AND2X1 U18470 ( .IN1(n16180), .IN2(n4411), .Q(n17683) );
  OR2X1 U18471 ( .IN1(n17685), .IN2(n17686), .Q(g21011) );
  AND2X1 U18472 ( .IN1(n16391), .IN2(g723), .Q(n17686) );
  AND2X1 U18473 ( .IN1(n16392), .IN2(n4396), .Q(n17685) );
  OR2X1 U18474 ( .IN1(n17687), .IN2(n17688), .Q(g21010) );
  AND2X1 U18475 ( .IN1(n16387), .IN2(g721), .Q(n17688) );
  AND2X1 U18476 ( .IN1(n16388), .IN2(n4477), .Q(n17687) );
  OR2X1 U18477 ( .IN1(n17689), .IN2(n17690), .Q(g21009) );
  AND2X1 U18478 ( .IN1(n16284), .IN2(g716), .Q(n17690) );
  AND2X1 U18479 ( .IN1(n680), .IN2(n10193), .Q(n17689) );
  OR2X1 U18480 ( .IN1(n17691), .IN2(n17692), .Q(g21007) );
  AND2X1 U18481 ( .IN1(n17189), .IN2(g2803), .Q(n17692) );
  AND2X1 U18482 ( .IN1(n17652), .IN2(n11222), .Q(n17691) );
  INVX0 U18483 ( .INP(n11146), .ZN(n11222) );
  OR2X1 U18484 ( .IN1(n17693), .IN2(n17694), .Q(n11146) );
  OR2X1 U18485 ( .IN1(n17695), .IN2(n17696), .Q(n17694) );
  AND2X1 U18486 ( .IN1(n12862), .IN2(g2688), .Q(n17696) );
  INVX0 U18487 ( .INP(n4314), .ZN(n12862) );
  AND2X1 U18488 ( .IN1(g2624), .IN2(g2694), .Q(n17695) );
  AND2X1 U18489 ( .IN1(g7390), .IN2(g2691), .Q(n17693) );
  INVX0 U18490 ( .INP(n17189), .ZN(n17652) );
  OR2X1 U18491 ( .IN1(n10156), .IN2(n4306), .Q(n17189) );
  OR2X1 U18492 ( .IN1(n17697), .IN2(n17698), .Q(g21006) );
  AND2X1 U18493 ( .IN1(n16079), .IN2(g2785), .Q(n17698) );
  AND2X1 U18494 ( .IN1(n16080), .IN2(n4397), .Q(n17697) );
  OR2X1 U18495 ( .IN1(n17699), .IN2(n17700), .Q(g21005) );
  AND2X1 U18496 ( .IN1(n16071), .IN2(g2783), .Q(n17700) );
  AND2X1 U18497 ( .IN1(n16072), .IN2(n4408), .Q(n17699) );
  OR2X1 U18498 ( .IN1(n17701), .IN2(n17702), .Q(g21004) );
  AND2X1 U18499 ( .IN1(n16068), .IN2(g2778), .Q(n17702) );
  AND2X1 U18500 ( .IN1(n16067), .IN2(n4419), .Q(n17701) );
  OR2X1 U18501 ( .IN1(n17703), .IN2(n17704), .Q(g21003) );
  AND2X1 U18502 ( .IN1(n17194), .IN2(g2112), .Q(n17704) );
  AND2X1 U18503 ( .IN1(n17705), .IN2(n11375), .Q(n17703) );
  INVX0 U18504 ( .INP(n11299), .ZN(n11375) );
  OR2X1 U18505 ( .IN1(n17706), .IN2(n17707), .Q(n11299) );
  OR2X1 U18506 ( .IN1(n17708), .IN2(n17709), .Q(n17707) );
  AND2X1 U18507 ( .IN1(g7194), .IN2(g1988), .Q(n17709) );
  AND2X1 U18508 ( .IN1(g7052), .IN2(g1985), .Q(n17708) );
  AND2X1 U18509 ( .IN1(g1930), .IN2(g1991), .Q(n17706) );
  OR2X1 U18510 ( .IN1(n17710), .IN2(n17711), .Q(g21002) );
  AND2X1 U18511 ( .IN1(n14337), .IN2(g2110), .Q(n17711) );
  AND2X1 U18512 ( .IN1(n17667), .IN2(n11383), .Q(n17710) );
  INVX0 U18513 ( .INP(n14337), .ZN(n17667) );
  OR2X1 U18514 ( .IN1(n17712), .IN2(n17713), .Q(g21001) );
  AND2X1 U18515 ( .IN1(n16277), .IN2(g2094), .Q(n17713) );
  AND2X1 U18516 ( .IN1(n16184), .IN2(n4409), .Q(n17712) );
  OR2X1 U18517 ( .IN1(n17714), .IN2(n17715), .Q(g21000) );
  AND2X1 U18518 ( .IN1(n16175), .IN2(n4399), .Q(n17715) );
  AND2X1 U18519 ( .IN1(test_so71), .IN2(n16176), .Q(n17714) );
  OR2X1 U18520 ( .IN1(n17716), .IN2(n17717), .Q(g20999) );
  AND2X1 U18521 ( .IN1(n16076), .IN2(g2087), .Q(n17717) );
  AND2X1 U18522 ( .IN1(n4149), .IN2(n4410), .Q(n17716) );
  OR2X1 U18523 ( .IN1(n17718), .IN2(n17719), .Q(g20997) );
  AND2X1 U18524 ( .IN1(n14345), .IN2(g1419), .Q(n17719) );
  AND2X1 U18525 ( .IN1(n17720), .IN2(n11538), .Q(n17718) );
  OR2X1 U18526 ( .IN1(n17721), .IN2(n17722), .Q(g20996) );
  AND2X1 U18527 ( .IN1(n17678), .IN2(n11546), .Q(n17722) );
  INVX0 U18528 ( .INP(n17192), .ZN(n17678) );
  AND2X1 U18529 ( .IN1(test_so51), .IN2(n17192), .Q(n17721) );
  OR2X1 U18530 ( .IN1(n10154), .IN2(n4294), .Q(n17192) );
  OR2X1 U18531 ( .IN1(n17723), .IN2(n17724), .Q(g20995) );
  AND2X1 U18532 ( .IN1(n16292), .IN2(g1403), .Q(n17724) );
  AND2X1 U18533 ( .IN1(n16293), .IN2(n4469), .Q(n17723) );
  OR2X1 U18534 ( .IN1(n17725), .IN2(n17726), .Q(g20994) );
  AND2X1 U18535 ( .IN1(n1027), .IN2(n4411), .Q(n17726) );
  AND2X1 U18536 ( .IN1(test_so50), .IN2(n16280), .Q(n17725) );
  OR2X1 U18537 ( .IN1(n17727), .IN2(n17728), .Q(g20993) );
  AND2X1 U18538 ( .IN1(n16181), .IN2(g1396), .Q(n17728) );
  AND2X1 U18539 ( .IN1(n16180), .IN2(n4401), .Q(n17727) );
  OR2X1 U18540 ( .IN1(n17729), .IN2(n17730), .Q(g20992) );
  AND2X1 U18541 ( .IN1(n17197), .IN2(g731), .Q(n17730) );
  AND2X1 U18542 ( .IN1(n17731), .IN2(n11046), .Q(n17729) );
  OR2X1 U18543 ( .IN1(n17732), .IN2(n17733), .Q(g20991) );
  AND2X1 U18544 ( .IN1(n16391), .IN2(g720), .Q(n17733) );
  AND2X1 U18545 ( .IN1(n16392), .IN2(n4477), .Q(n17732) );
  OR2X1 U18546 ( .IN1(n17734), .IN2(n17735), .Q(g20990) );
  AND2X1 U18547 ( .IN1(n16387), .IN2(g718), .Q(n17735) );
  AND2X1 U18548 ( .IN1(n16388), .IN2(n10193), .Q(n17734) );
  OR2X1 U18549 ( .IN1(n17736), .IN2(n17737), .Q(g20989) );
  AND2X1 U18550 ( .IN1(n16284), .IN2(g713), .Q(n17737) );
  AND2X1 U18551 ( .IN1(n680), .IN2(n4413), .Q(n17736) );
  OR2X1 U18552 ( .IN1(n17738), .IN2(n17739), .Q(g20983) );
  AND2X1 U18553 ( .IN1(n16079), .IN2(g2782), .Q(n17739) );
  AND2X1 U18554 ( .IN1(n16080), .IN2(n4408), .Q(n17738) );
  OR2X1 U18555 ( .IN1(n17740), .IN2(n17741), .Q(g20982) );
  AND2X1 U18556 ( .IN1(n16071), .IN2(g2780), .Q(n17741) );
  AND2X1 U18557 ( .IN1(n16072), .IN2(n4419), .Q(n17740) );
  OR2X1 U18558 ( .IN1(n17742), .IN2(n17743), .Q(g20981) );
  AND2X1 U18559 ( .IN1(n16068), .IN2(g2775), .Q(n17743) );
  AND2X1 U18560 ( .IN1(n16067), .IN2(n4472), .Q(n17742) );
  OR2X1 U18561 ( .IN1(n17744), .IN2(n17745), .Q(g20980) );
  AND2X1 U18562 ( .IN1(n17194), .IN2(g2109), .Q(n17745) );
  AND2X1 U18563 ( .IN1(n17705), .IN2(n11383), .Q(n17744) );
  INVX0 U18564 ( .INP(n11309), .ZN(n11383) );
  OR2X1 U18565 ( .IN1(n17746), .IN2(n17747), .Q(n11309) );
  OR2X1 U18566 ( .IN1(n17748), .IN2(n17749), .Q(n17747) );
  AND2X1 U18567 ( .IN1(g7194), .IN2(g1997), .Q(n17749) );
  AND2X1 U18568 ( .IN1(n13973), .IN2(g1994), .Q(n17748) );
  INVX0 U18569 ( .INP(n4296), .ZN(n13973) );
  AND2X1 U18570 ( .IN1(g1930), .IN2(g2000), .Q(n17746) );
  INVX0 U18571 ( .INP(n17194), .ZN(n17705) );
  OR2X1 U18572 ( .IN1(n10155), .IN2(n4307), .Q(n17194) );
  OR2X1 U18573 ( .IN1(n17750), .IN2(n17751), .Q(g20979) );
  AND2X1 U18574 ( .IN1(n16277), .IN2(g2091), .Q(n17751) );
  AND2X1 U18575 ( .IN1(n16184), .IN2(n4399), .Q(n17750) );
  OR2X1 U18576 ( .IN1(n17752), .IN2(n17753), .Q(g20978) );
  AND2X1 U18577 ( .IN1(n16176), .IN2(g2089), .Q(n17753) );
  AND2X1 U18578 ( .IN1(n16175), .IN2(n4410), .Q(n17752) );
  OR2X1 U18579 ( .IN1(n17754), .IN2(n17755), .Q(g20977) );
  AND2X1 U18580 ( .IN1(n16076), .IN2(g2084), .Q(n17755) );
  AND2X1 U18581 ( .IN1(n4149), .IN2(n4420), .Q(n17754) );
  OR2X1 U18582 ( .IN1(n17756), .IN2(n17757), .Q(g20976) );
  AND2X1 U18583 ( .IN1(n17199), .IN2(g1418), .Q(n17757) );
  AND2X1 U18584 ( .IN1(n17758), .IN2(n11538), .Q(n17756) );
  INVX0 U18585 ( .INP(n11461), .ZN(n11538) );
  OR2X1 U18586 ( .IN1(n17759), .IN2(n17760), .Q(n11461) );
  OR2X1 U18587 ( .IN1(n17761), .IN2(n17762), .Q(n17760) );
  AND2X1 U18588 ( .IN1(g1236), .IN2(g1297), .Q(n17762) );
  AND2X1 U18589 ( .IN1(g6750), .IN2(g1291), .Q(n17761) );
  AND2X1 U18590 ( .IN1(g6944), .IN2(g1294), .Q(n17759) );
  OR2X1 U18591 ( .IN1(n17763), .IN2(n17764), .Q(g20975) );
  AND2X1 U18592 ( .IN1(n14345), .IN2(g1416), .Q(n17764) );
  AND2X1 U18593 ( .IN1(n17720), .IN2(n11546), .Q(n17763) );
  INVX0 U18594 ( .INP(n14345), .ZN(n17720) );
  OR2X1 U18595 ( .IN1(n17765), .IN2(n17766), .Q(g20974) );
  AND2X1 U18596 ( .IN1(n16292), .IN2(g1400), .Q(n17766) );
  AND2X1 U18597 ( .IN1(n16293), .IN2(n4411), .Q(n17765) );
  OR2X1 U18598 ( .IN1(n17767), .IN2(n17768), .Q(g20973) );
  AND2X1 U18599 ( .IN1(n16280), .IN2(g1398), .Q(n17768) );
  AND2X1 U18600 ( .IN1(n1027), .IN2(n4401), .Q(n17767) );
  OR2X1 U18601 ( .IN1(n17769), .IN2(n17770), .Q(g20972) );
  AND2X1 U18602 ( .IN1(n16181), .IN2(g1393), .Q(n17770) );
  AND2X1 U18603 ( .IN1(n16180), .IN2(n4412), .Q(n17769) );
  OR2X1 U18604 ( .IN1(n17771), .IN2(n17772), .Q(g20970) );
  AND2X1 U18605 ( .IN1(n13809), .IN2(g733), .Q(n17772) );
  AND2X1 U18606 ( .IN1(n17773), .IN2(n11046), .Q(n17771) );
  OR2X1 U18607 ( .IN1(n17774), .IN2(n17775), .Q(g20969) );
  AND2X1 U18608 ( .IN1(n17197), .IN2(g728), .Q(n17775) );
  AND2X1 U18609 ( .IN1(n17731), .IN2(n11058), .Q(n17774) );
  INVX0 U18610 ( .INP(n17197), .ZN(n17731) );
  OR2X1 U18611 ( .IN1(n10153), .IN2(n4295), .Q(n17197) );
  OR2X1 U18612 ( .IN1(n17776), .IN2(n17777), .Q(g20968) );
  AND2X1 U18613 ( .IN1(n16391), .IN2(g717), .Q(n17777) );
  AND2X1 U18614 ( .IN1(n16392), .IN2(n10193), .Q(n17776) );
  OR2X1 U18615 ( .IN1(n17778), .IN2(n17779), .Q(g20967) );
  AND2X1 U18616 ( .IN1(n16387), .IN2(g715), .Q(n17779) );
  AND2X1 U18617 ( .IN1(n16388), .IN2(n4413), .Q(n17778) );
  OR2X1 U18618 ( .IN1(n17780), .IN2(n17781), .Q(g20966) );
  AND2X1 U18619 ( .IN1(n16284), .IN2(g710), .Q(n17781) );
  AND2X1 U18620 ( .IN1(n680), .IN2(n4403), .Q(n17780) );
  OR2X1 U18621 ( .IN1(n17782), .IN2(n17783), .Q(g20965) );
  AND2X1 U18622 ( .IN1(n16068), .IN2(g2799), .Q(n17783) );
  AND2X1 U18623 ( .IN1(n16067), .IN2(n4415), .Q(n17782) );
  OR2X1 U18624 ( .IN1(n17784), .IN2(n17785), .Q(g20964) );
  AND2X1 U18625 ( .IN1(n16079), .IN2(g2779), .Q(n17785) );
  AND2X1 U18626 ( .IN1(n16080), .IN2(n4419), .Q(n17784) );
  OR2X1 U18627 ( .IN1(n17786), .IN2(n17787), .Q(g20963) );
  AND2X1 U18628 ( .IN1(n16071), .IN2(g2777), .Q(n17787) );
  AND2X1 U18629 ( .IN1(n16072), .IN2(n4472), .Q(n17786) );
  OR2X1 U18630 ( .IN1(n17788), .IN2(n17789), .Q(g20962) );
  AND2X1 U18631 ( .IN1(n16068), .IN2(g2772), .Q(n17789) );
  AND2X1 U18632 ( .IN1(n16067), .IN2(n4398), .Q(n17788) );
  INVX0 U18633 ( .INP(n16068), .ZN(n16067) );
  OR2X1 U18634 ( .IN1(n4292), .IN2(n17790), .Q(n16068) );
  OR2X1 U18635 ( .IN1(n17791), .IN2(n17792), .Q(g20955) );
  AND2X1 U18636 ( .IN1(n16277), .IN2(g2088), .Q(n17792) );
  AND2X1 U18637 ( .IN1(n16184), .IN2(n4410), .Q(n17791) );
  OR2X1 U18638 ( .IN1(n17793), .IN2(n17794), .Q(g20954) );
  AND2X1 U18639 ( .IN1(n16176), .IN2(g2086), .Q(n17794) );
  AND2X1 U18640 ( .IN1(n16175), .IN2(n4420), .Q(n17793) );
  OR2X1 U18641 ( .IN1(n17795), .IN2(n17796), .Q(g20953) );
  AND2X1 U18642 ( .IN1(n16076), .IN2(g2081), .Q(n17796) );
  AND2X1 U18643 ( .IN1(n4149), .IN2(n4474), .Q(n17795) );
  OR2X1 U18644 ( .IN1(n17797), .IN2(n17798), .Q(g20952) );
  AND2X1 U18645 ( .IN1(n17199), .IN2(g1415), .Q(n17798) );
  AND2X1 U18646 ( .IN1(n17758), .IN2(n11546), .Q(n17797) );
  INVX0 U18647 ( .INP(n11471), .ZN(n11546) );
  OR2X1 U18648 ( .IN1(n17799), .IN2(n17800), .Q(n11471) );
  OR2X1 U18649 ( .IN1(n17801), .IN2(n17802), .Q(n17800) );
  AND2X1 U18650 ( .IN1(g6944), .IN2(g1303), .Q(n17802) );
  AND2X1 U18651 ( .IN1(g1236), .IN2(g1306), .Q(n17801) );
  AND2X1 U18652 ( .IN1(n13842), .IN2(g1300), .Q(n17799) );
  INVX0 U18653 ( .INP(n4371), .ZN(n13842) );
  INVX0 U18654 ( .INP(n17199), .ZN(n17758) );
  OR2X1 U18655 ( .IN1(n10154), .IN2(n4308), .Q(n17199) );
  OR2X1 U18656 ( .IN1(n17803), .IN2(n17804), .Q(g20951) );
  AND2X1 U18657 ( .IN1(n16292), .IN2(g1397), .Q(n17804) );
  AND2X1 U18658 ( .IN1(n16293), .IN2(n4401), .Q(n17803) );
  OR2X1 U18659 ( .IN1(n17805), .IN2(n17806), .Q(g20950) );
  AND2X1 U18660 ( .IN1(n16280), .IN2(g1395), .Q(n17806) );
  AND2X1 U18661 ( .IN1(n1027), .IN2(n4412), .Q(n17805) );
  OR2X1 U18662 ( .IN1(n17807), .IN2(n17808), .Q(g20949) );
  AND2X1 U18663 ( .IN1(n16181), .IN2(g1390), .Q(n17808) );
  AND2X1 U18664 ( .IN1(n16180), .IN2(n4421), .Q(n17807) );
  OR2X1 U18665 ( .IN1(n17809), .IN2(n17810), .Q(g20948) );
  AND2X1 U18666 ( .IN1(n17202), .IN2(g732), .Q(n17810) );
  AND2X1 U18667 ( .IN1(n17811), .IN2(n11046), .Q(n17809) );
  INVX0 U18668 ( .INP(n10967), .ZN(n11046) );
  OR2X1 U18669 ( .IN1(n17812), .IN2(n17813), .Q(n10967) );
  OR2X1 U18670 ( .IN1(n17814), .IN2(n17815), .Q(n17813) );
  AND2X1 U18671 ( .IN1(g550), .IN2(g611), .Q(n17815) );
  AND2X1 U18672 ( .IN1(n11054), .IN2(g605), .Q(n17814) );
  INVX0 U18673 ( .INP(n4298), .ZN(n11054) );
  AND2X1 U18674 ( .IN1(g6642), .IN2(g608), .Q(n17812) );
  OR2X1 U18675 ( .IN1(n17816), .IN2(n17817), .Q(g20947) );
  AND2X1 U18676 ( .IN1(n13809), .IN2(g730), .Q(n17817) );
  AND2X1 U18677 ( .IN1(n17773), .IN2(n11058), .Q(n17816) );
  INVX0 U18678 ( .INP(n13809), .ZN(n17773) );
  OR2X1 U18679 ( .IN1(n17818), .IN2(n17819), .Q(g20946) );
  AND2X1 U18680 ( .IN1(n16391), .IN2(g714), .Q(n17819) );
  AND2X1 U18681 ( .IN1(n16392), .IN2(n4413), .Q(n17818) );
  OR2X1 U18682 ( .IN1(n17820), .IN2(n17821), .Q(g20945) );
  AND2X1 U18683 ( .IN1(n16387), .IN2(g712), .Q(n17821) );
  AND2X1 U18684 ( .IN1(n16388), .IN2(n4403), .Q(n17820) );
  OR2X1 U18685 ( .IN1(n17822), .IN2(n17823), .Q(g20944) );
  AND2X1 U18686 ( .IN1(n16284), .IN2(g707), .Q(n17823) );
  AND2X1 U18687 ( .IN1(n680), .IN2(n4414), .Q(n17822) );
  OR2X1 U18688 ( .IN1(n17824), .IN2(n17825), .Q(g20941) );
  AND2X1 U18689 ( .IN1(n16071), .IN2(g2801), .Q(n17825) );
  AND2X1 U18690 ( .IN1(n16072), .IN2(n4415), .Q(n17824) );
  OR2X1 U18691 ( .IN1(n17826), .IN2(n17827), .Q(g20940) );
  AND2X1 U18692 ( .IN1(n16079), .IN2(g2776), .Q(n17827) );
  AND2X1 U18693 ( .IN1(n16080), .IN2(n4472), .Q(n17826) );
  OR2X1 U18694 ( .IN1(n17828), .IN2(n17829), .Q(g20939) );
  AND2X1 U18695 ( .IN1(n16071), .IN2(g2774), .Q(n17829) );
  AND2X1 U18696 ( .IN1(n16072), .IN2(n4398), .Q(n17828) );
  INVX0 U18697 ( .INP(n16071), .ZN(n16072) );
  OR2X1 U18698 ( .IN1(n4356), .IN2(n17790), .Q(n16071) );
  OR2X1 U18699 ( .IN1(n17830), .IN2(n17831), .Q(g20937) );
  AND2X1 U18700 ( .IN1(n16076), .IN2(g2105), .Q(n17831) );
  AND2X1 U18701 ( .IN1(n4149), .IN2(n4416), .Q(n17830) );
  OR2X1 U18702 ( .IN1(n17832), .IN2(n17833), .Q(g20936) );
  AND2X1 U18703 ( .IN1(n16277), .IN2(g2085), .Q(n17833) );
  AND2X1 U18704 ( .IN1(n16184), .IN2(n4420), .Q(n17832) );
  OR2X1 U18705 ( .IN1(n17834), .IN2(n17835), .Q(g20935) );
  AND2X1 U18706 ( .IN1(n16176), .IN2(g2083), .Q(n17835) );
  AND2X1 U18707 ( .IN1(n16175), .IN2(n4474), .Q(n17834) );
  OR2X1 U18708 ( .IN1(n17836), .IN2(n17837), .Q(g20934) );
  AND2X1 U18709 ( .IN1(n16076), .IN2(g2078), .Q(n17837) );
  AND2X1 U18710 ( .IN1(n4149), .IN2(n4400), .Q(n17836) );
  INVX0 U18711 ( .INP(n16076), .ZN(n4149) );
  OR2X1 U18712 ( .IN1(n4293), .IN2(n17838), .Q(n16076) );
  OR2X1 U18713 ( .IN1(n17839), .IN2(n17840), .Q(g20927) );
  AND2X1 U18714 ( .IN1(n16292), .IN2(g1394), .Q(n17840) );
  AND2X1 U18715 ( .IN1(n16293), .IN2(n4412), .Q(n17839) );
  OR2X1 U18716 ( .IN1(n17841), .IN2(n17842), .Q(g20926) );
  AND2X1 U18717 ( .IN1(n16280), .IN2(g1392), .Q(n17842) );
  AND2X1 U18718 ( .IN1(n1027), .IN2(n4421), .Q(n17841) );
  OR2X1 U18719 ( .IN1(n17843), .IN2(n17844), .Q(g20925) );
  AND2X1 U18720 ( .IN1(n16181), .IN2(g1387), .Q(n17844) );
  AND2X1 U18721 ( .IN1(n16180), .IN2(n4476), .Q(n17843) );
  OR2X1 U18722 ( .IN1(n17845), .IN2(n17846), .Q(g20924) );
  AND2X1 U18723 ( .IN1(n17202), .IN2(g729), .Q(n17846) );
  AND2X1 U18724 ( .IN1(n17811), .IN2(n11058), .Q(n17845) );
  INVX0 U18725 ( .INP(n10961), .ZN(n11058) );
  OR2X1 U18726 ( .IN1(n17847), .IN2(n17848), .Q(n10961) );
  OR2X1 U18727 ( .IN1(n17849), .IN2(n17850), .Q(n17848) );
  AND2X1 U18728 ( .IN1(test_so26), .IN2(g550), .Q(n17850) );
  AND2X1 U18729 ( .IN1(g6485), .IN2(g614), .Q(n17849) );
  AND2X1 U18730 ( .IN1(g6642), .IN2(g617), .Q(n17847) );
  INVX0 U18731 ( .INP(n17202), .ZN(n17811) );
  OR2X1 U18732 ( .IN1(n10153), .IN2(n4309), .Q(n17202) );
  OR2X1 U18733 ( .IN1(n17851), .IN2(n17852), .Q(g20923) );
  AND2X1 U18734 ( .IN1(n16392), .IN2(n4403), .Q(n17852) );
  AND2X1 U18735 ( .IN1(test_so29), .IN2(n16391), .Q(n17851) );
  OR2X1 U18736 ( .IN1(n17853), .IN2(n17854), .Q(g20922) );
  AND2X1 U18737 ( .IN1(n16387), .IN2(g709), .Q(n17854) );
  AND2X1 U18738 ( .IN1(n16388), .IN2(n4414), .Q(n17853) );
  OR2X1 U18739 ( .IN1(n17855), .IN2(n17856), .Q(g20921) );
  AND2X1 U18740 ( .IN1(n16284), .IN2(g704), .Q(n17856) );
  AND2X1 U18741 ( .IN1(n680), .IN2(n4422), .Q(n17855) );
  OR2X1 U18742 ( .IN1(n17857), .IN2(n17858), .Q(g20919) );
  AND2X1 U18743 ( .IN1(n16079), .IN2(g2800), .Q(n17858) );
  AND2X1 U18744 ( .IN1(n16080), .IN2(n4415), .Q(n17857) );
  OR2X1 U18745 ( .IN1(n17859), .IN2(n17860), .Q(g20918) );
  AND2X1 U18746 ( .IN1(n16079), .IN2(g2773), .Q(n17860) );
  AND2X1 U18747 ( .IN1(n16080), .IN2(n4398), .Q(n17859) );
  INVX0 U18748 ( .INP(n16079), .ZN(n16080) );
  OR2X1 U18749 ( .IN1(n4306), .IN2(n17790), .Q(n16079) );
  OR2X1 U18750 ( .IN1(g2733), .IN2(n17861), .Q(n17790) );
  OR2X1 U18751 ( .IN1(n9895), .IN2(n4490), .Q(n17861) );
  OR2X1 U18752 ( .IN1(n17862), .IN2(n17863), .Q(g20917) );
  AND2X1 U18753 ( .IN1(n16175), .IN2(n4416), .Q(n17863) );
  AND2X1 U18754 ( .IN1(test_so72), .IN2(n16176), .Q(n17862) );
  OR2X1 U18755 ( .IN1(n17864), .IN2(n17865), .Q(g20916) );
  AND2X1 U18756 ( .IN1(n16277), .IN2(g2082), .Q(n17865) );
  AND2X1 U18757 ( .IN1(n16184), .IN2(n4474), .Q(n17864) );
  OR2X1 U18758 ( .IN1(n17866), .IN2(n17867), .Q(g20915) );
  AND2X1 U18759 ( .IN1(n16176), .IN2(g2080), .Q(n17867) );
  AND2X1 U18760 ( .IN1(n16175), .IN2(n4400), .Q(n17866) );
  INVX0 U18761 ( .INP(n16176), .ZN(n16175) );
  OR2X1 U18762 ( .IN1(n4357), .IN2(n17838), .Q(n16176) );
  OR2X1 U18763 ( .IN1(n17868), .IN2(n17869), .Q(g20913) );
  AND2X1 U18764 ( .IN1(n16181), .IN2(g1411), .Q(n17869) );
  AND2X1 U18765 ( .IN1(n16180), .IN2(n4417), .Q(n17868) );
  OR2X1 U18766 ( .IN1(n17870), .IN2(n17871), .Q(g20912) );
  AND2X1 U18767 ( .IN1(n16292), .IN2(g1391), .Q(n17871) );
  AND2X1 U18768 ( .IN1(n16293), .IN2(n4421), .Q(n17870) );
  OR2X1 U18769 ( .IN1(n17872), .IN2(n17873), .Q(g20911) );
  AND2X1 U18770 ( .IN1(n16280), .IN2(g1389), .Q(n17873) );
  AND2X1 U18771 ( .IN1(n1027), .IN2(n4476), .Q(n17872) );
  OR2X1 U18772 ( .IN1(n17874), .IN2(n17875), .Q(g20910) );
  AND2X1 U18773 ( .IN1(n16181), .IN2(g1384), .Q(n17875) );
  AND2X1 U18774 ( .IN1(n16180), .IN2(n4402), .Q(n17874) );
  INVX0 U18775 ( .INP(n16181), .ZN(n16180) );
  OR2X1 U18776 ( .IN1(n4294), .IN2(n17876), .Q(n16181) );
  OR2X1 U18777 ( .IN1(n17877), .IN2(n17878), .Q(g20903) );
  AND2X1 U18778 ( .IN1(n16391), .IN2(g708), .Q(n17878) );
  AND2X1 U18779 ( .IN1(n16392), .IN2(n4414), .Q(n17877) );
  OR2X1 U18780 ( .IN1(n17879), .IN2(n17880), .Q(g20902) );
  AND2X1 U18781 ( .IN1(n16387), .IN2(g706), .Q(n17880) );
  AND2X1 U18782 ( .IN1(n16388), .IN2(n4422), .Q(n17879) );
  OR2X1 U18783 ( .IN1(n17881), .IN2(n17882), .Q(g20901) );
  AND2X1 U18784 ( .IN1(n16284), .IN2(g701), .Q(n17882) );
  AND2X1 U18785 ( .IN1(n680), .IN2(n4478), .Q(n17881) );
  OR2X1 U18786 ( .IN1(n17883), .IN2(n17884), .Q(g20900) );
  AND2X1 U18787 ( .IN1(n16277), .IN2(g2106), .Q(n17884) );
  AND2X1 U18788 ( .IN1(n16184), .IN2(n4416), .Q(n17883) );
  OR2X1 U18789 ( .IN1(n17885), .IN2(n17886), .Q(g20899) );
  AND2X1 U18790 ( .IN1(n16277), .IN2(g2079), .Q(n17886) );
  AND2X1 U18791 ( .IN1(n16184), .IN2(n4400), .Q(n17885) );
  INVX0 U18792 ( .INP(n16277), .ZN(n16184) );
  OR2X1 U18793 ( .IN1(n4307), .IN2(n17838), .Q(n16277) );
  OR2X1 U18794 ( .IN1(n10201), .IN2(n17887), .Q(n17838) );
  OR2X1 U18795 ( .IN1(n9896), .IN2(g2039), .Q(n17887) );
  OR2X1 U18796 ( .IN1(n17888), .IN2(n17889), .Q(g20898) );
  AND2X1 U18797 ( .IN1(n16280), .IN2(g1413), .Q(n17889) );
  AND2X1 U18798 ( .IN1(n1027), .IN2(n4417), .Q(n17888) );
  OR2X1 U18799 ( .IN1(n17890), .IN2(n17891), .Q(g20897) );
  AND2X1 U18800 ( .IN1(n16292), .IN2(g1388), .Q(n17891) );
  AND2X1 U18801 ( .IN1(n16293), .IN2(n4476), .Q(n17890) );
  OR2X1 U18802 ( .IN1(n17892), .IN2(n17893), .Q(g20896) );
  AND2X1 U18803 ( .IN1(n16280), .IN2(g1386), .Q(n17893) );
  AND2X1 U18804 ( .IN1(n1027), .IN2(n4402), .Q(n17892) );
  INVX0 U18805 ( .INP(n16280), .ZN(n1027) );
  OR2X1 U18806 ( .IN1(n4358), .IN2(n17876), .Q(n16280) );
  OR2X1 U18807 ( .IN1(n17894), .IN2(n17895), .Q(g20894) );
  AND2X1 U18808 ( .IN1(n16284), .IN2(g725), .Q(n17895) );
  AND2X1 U18809 ( .IN1(n680), .IN2(n4418), .Q(n17894) );
  OR2X1 U18810 ( .IN1(n17896), .IN2(n17897), .Q(g20893) );
  AND2X1 U18811 ( .IN1(n16391), .IN2(g705), .Q(n17897) );
  AND2X1 U18812 ( .IN1(n16392), .IN2(n4422), .Q(n17896) );
  OR2X1 U18813 ( .IN1(n17898), .IN2(n17899), .Q(g20892) );
  AND2X1 U18814 ( .IN1(n16387), .IN2(g703), .Q(n17899) );
  AND2X1 U18815 ( .IN1(n16388), .IN2(n4478), .Q(n17898) );
  OR2X1 U18816 ( .IN1(n17900), .IN2(n17901), .Q(g20891) );
  AND2X1 U18817 ( .IN1(n16284), .IN2(g698), .Q(n17901) );
  AND2X1 U18818 ( .IN1(n680), .IN2(n4404), .Q(n17900) );
  INVX0 U18819 ( .INP(n16284), .ZN(n680) );
  OR2X1 U18820 ( .IN1(n4295), .IN2(n17902), .Q(n16284) );
  AND2X1 U18821 ( .IN1(n17033), .IN2(n7913), .Q(g20884) );
  INVX0 U18822 ( .INP(g3234), .ZN(n17033) );
  OR2X1 U18823 ( .IN1(n17903), .IN2(n17904), .Q(g20883) );
  AND2X1 U18824 ( .IN1(n16292), .IN2(g1412), .Q(n17904) );
  AND2X1 U18825 ( .IN1(n16293), .IN2(n4417), .Q(n17903) );
  OR2X1 U18826 ( .IN1(n17905), .IN2(n17906), .Q(g20882) );
  AND2X1 U18827 ( .IN1(n16293), .IN2(n4402), .Q(n17906) );
  INVX0 U18828 ( .INP(n16292), .ZN(n16293) );
  AND2X1 U18829 ( .IN1(test_so49), .IN2(n16292), .Q(n17905) );
  OR2X1 U18830 ( .IN1(n4308), .IN2(n17876), .Q(n16292) );
  OR2X1 U18831 ( .IN1(g1345), .IN2(n17907), .Q(n17876) );
  OR2X1 U18832 ( .IN1(n9897), .IN2(n4489), .Q(n17907) );
  OR2X1 U18833 ( .IN1(n17908), .IN2(n17909), .Q(g20881) );
  AND2X1 U18834 ( .IN1(n16388), .IN2(n4418), .Q(n17909) );
  AND2X1 U18835 ( .IN1(test_so30), .IN2(n16387), .Q(n17908) );
  OR2X1 U18836 ( .IN1(n17910), .IN2(n17911), .Q(g20880) );
  AND2X1 U18837 ( .IN1(n16391), .IN2(g702), .Q(n17911) );
  AND2X1 U18838 ( .IN1(n16392), .IN2(n4478), .Q(n17910) );
  OR2X1 U18839 ( .IN1(n17912), .IN2(n17913), .Q(g20879) );
  AND2X1 U18840 ( .IN1(n16387), .IN2(g700), .Q(n17913) );
  AND2X1 U18841 ( .IN1(n16388), .IN2(n4404), .Q(n17912) );
  INVX0 U18842 ( .INP(n16387), .ZN(n16388) );
  OR2X1 U18843 ( .IN1(n4359), .IN2(n17902), .Q(n16387) );
  OR2X1 U18844 ( .IN1(n17914), .IN2(n17915), .Q(g20876) );
  AND2X1 U18845 ( .IN1(n16391), .IN2(g726), .Q(n17915) );
  AND2X1 U18846 ( .IN1(n16392), .IN2(n4418), .Q(n17914) );
  OR2X1 U18847 ( .IN1(n17916), .IN2(n17917), .Q(g20875) );
  AND2X1 U18848 ( .IN1(n16391), .IN2(g699), .Q(n17917) );
  AND2X1 U18849 ( .IN1(n16392), .IN2(n4404), .Q(n17916) );
  INVX0 U18850 ( .INP(n16391), .ZN(n16392) );
  OR2X1 U18851 ( .IN1(n4309), .IN2(n17902), .Q(n16391) );
  OR2X1 U18852 ( .IN1(g659), .IN2(n17918), .Q(n17902) );
  OR2X1 U18853 ( .IN1(n9898), .IN2(n4492), .Q(n17918) );
  OR2X1 U18854 ( .IN1(n17919), .IN2(n17920), .Q(g20874) );
  AND2X1 U18855 ( .IN1(n4351), .IN2(n17528), .Q(n17920) );
  AND2X1 U18856 ( .IN1(n17921), .IN2(n17922), .Q(n17528) );
  OR2X1 U18857 ( .IN1(n10612), .IN2(n17534), .Q(n17922) );
  INVX0 U18858 ( .INP(n17923), .ZN(n17921) );
  AND2X1 U18859 ( .IN1(n17534), .IN2(n10612), .Q(n17923) );
  AND2X1 U18860 ( .IN1(n17924), .IN2(n17925), .Q(n10612) );
  INVX0 U18861 ( .INP(n17926), .ZN(n17925) );
  AND2X1 U18862 ( .IN1(n17927), .IN2(n17928), .Q(n17926) );
  OR2X1 U18863 ( .IN1(n17928), .IN2(n17927), .Q(n17924) );
  OR2X1 U18864 ( .IN1(n17929), .IN2(n17930), .Q(n17927) );
  AND2X1 U18865 ( .IN1(n17931), .IN2(n17932), .Q(n17930) );
  INVX0 U18866 ( .INP(n17933), .ZN(n17929) );
  OR2X1 U18867 ( .IN1(n17932), .IN2(n17931), .Q(n17933) );
  OR2X1 U18868 ( .IN1(n17934), .IN2(n17935), .Q(n17931) );
  AND2X1 U18869 ( .IN1(n10129), .IN2(g2959), .Q(n17935) );
  AND2X1 U18870 ( .IN1(n10130), .IN2(g2941), .Q(n17934) );
  INVX0 U18871 ( .INP(n17936), .ZN(n17932) );
  OR2X1 U18872 ( .IN1(n17937), .IN2(n17938), .Q(n17936) );
  AND2X1 U18873 ( .IN1(n10131), .IN2(g2938), .Q(n17938) );
  AND2X1 U18874 ( .IN1(n10132), .IN2(g2935), .Q(n17937) );
  AND2X1 U18875 ( .IN1(n17939), .IN2(n17940), .Q(n17928) );
  INVX0 U18876 ( .INP(n17941), .ZN(n17940) );
  AND2X1 U18877 ( .IN1(n17942), .IN2(n17943), .Q(n17941) );
  OR2X1 U18878 ( .IN1(n17943), .IN2(n17942), .Q(n17939) );
  OR2X1 U18879 ( .IN1(n17944), .IN2(n17945), .Q(n17942) );
  AND2X1 U18880 ( .IN1(n10133), .IN2(g2953), .Q(n17945) );
  AND2X1 U18881 ( .IN1(n10134), .IN2(g2947), .Q(n17944) );
  INVX0 U18882 ( .INP(n17946), .ZN(n17943) );
  OR2X1 U18883 ( .IN1(n17947), .IN2(n17948), .Q(n17946) );
  AND2X1 U18884 ( .IN1(n10135), .IN2(g2956), .Q(n17948) );
  AND2X1 U18885 ( .IN1(n10136), .IN2(g2944), .Q(n17947) );
  AND2X1 U18886 ( .IN1(n10944), .IN2(n8079), .Q(n17534) );
  INVX0 U18887 ( .INP(g3231), .ZN(n10944) );
  AND2X1 U18888 ( .IN1(g2879), .IN2(g8096), .Q(n17919) );
  AND2X1 U18889 ( .IN1(n17949), .IN2(n17950), .Q(g20789) );
  OR2X1 U18890 ( .IN1(n17951), .IN2(g2714), .Q(n17950) );
  AND2X1 U18891 ( .IN1(n4426), .IN2(g2703), .Q(n17951) );
  AND2X1 U18892 ( .IN1(n17508), .IN2(n14331), .Q(n17949) );
  OR2X1 U18893 ( .IN1(n10156), .IN2(n4356), .Q(n14331) );
  OR2X1 U18894 ( .IN1(g2733), .IN2(n17952), .Q(n17508) );
  OR2X1 U18895 ( .IN1(n4398), .IN2(n4292), .Q(n17952) );
  AND2X1 U18896 ( .IN1(n17953), .IN2(n17954), .Q(g20752) );
  OR2X1 U18897 ( .IN1(n17955), .IN2(g2020), .Q(n17954) );
  AND2X1 U18898 ( .IN1(n4427), .IN2(g2009), .Q(n17955) );
  AND2X1 U18899 ( .IN1(n17512), .IN2(n14337), .Q(n17953) );
  OR2X1 U18900 ( .IN1(n10155), .IN2(n4357), .Q(n14337) );
  OR2X1 U18901 ( .IN1(g2039), .IN2(n17956), .Q(n17512) );
  OR2X1 U18902 ( .IN1(n4400), .IN2(n4293), .Q(n17956) );
  AND2X1 U18903 ( .IN1(n17957), .IN2(n17958), .Q(g20717) );
  OR2X1 U18904 ( .IN1(n17959), .IN2(g1326), .Q(n17958) );
  AND2X1 U18905 ( .IN1(n4428), .IN2(g1315), .Q(n17959) );
  AND2X1 U18906 ( .IN1(n17522), .IN2(n14345), .Q(n17957) );
  OR2X1 U18907 ( .IN1(n10154), .IN2(n4358), .Q(n14345) );
  OR2X1 U18908 ( .IN1(g1345), .IN2(n17960), .Q(n17522) );
  OR2X1 U18909 ( .IN1(n4402), .IN2(n4294), .Q(n17960) );
  AND2X1 U18910 ( .IN1(n17961), .IN2(n17962), .Q(g20682) );
  OR2X1 U18911 ( .IN1(n17963), .IN2(g640), .Q(n17962) );
  AND2X1 U18912 ( .IN1(n4429), .IN2(g629), .Q(n17963) );
  AND2X1 U18913 ( .IN1(n17072), .IN2(n13809), .Q(n17961) );
  OR2X1 U18914 ( .IN1(n10153), .IN2(n4359), .Q(n13809) );
  OR2X1 U18915 ( .IN1(g659), .IN2(n17964), .Q(n17072) );
  OR2X1 U18916 ( .IN1(n4404), .IN2(n4295), .Q(n17964) );
  OR2X1 U18917 ( .IN1(n17965), .IN2(n17966), .Q(g20417) );
  AND2X1 U18918 ( .IN1(n4351), .IN2(g2963), .Q(n17966) );
  AND2X1 U18919 ( .IN1(g2879), .IN2(g7334), .Q(n17965) );
  OR2X1 U18920 ( .IN1(n17967), .IN2(n17968), .Q(g20376) );
  AND2X1 U18921 ( .IN1(g2879), .IN2(g6895), .Q(n17968) );
  AND2X1 U18922 ( .IN1(n4351), .IN2(test_so2), .Q(n17967) );
  OR2X1 U18923 ( .IN1(n17969), .IN2(n17970), .Q(g20375) );
  AND2X1 U18924 ( .IN1(n17176), .IN2(g2703), .Q(n17970) );
  AND2X1 U18925 ( .IN1(n4292), .IN2(g2733), .Q(n17969) );
  OR2X1 U18926 ( .IN1(n17971), .IN2(n17972), .Q(g20353) );
  AND2X1 U18927 ( .IN1(n17176), .IN2(g2009), .Q(n17972) );
  AND2X1 U18928 ( .IN1(n4293), .IN2(g2039), .Q(n17971) );
  OR2X1 U18929 ( .IN1(n17973), .IN2(n17974), .Q(g20343) );
  AND2X1 U18930 ( .IN1(n4351), .IN2(g2969), .Q(n17974) );
  AND2X1 U18931 ( .IN1(g2879), .IN2(g6442), .Q(n17973) );
  OR2X1 U18932 ( .IN1(n17975), .IN2(n17976), .Q(g20333) );
  AND2X1 U18933 ( .IN1(n17176), .IN2(g1315), .Q(n17976) );
  AND2X1 U18934 ( .IN1(n4294), .IN2(g1345), .Q(n17975) );
  OR2X1 U18935 ( .IN1(n17977), .IN2(n17978), .Q(g20314) );
  AND2X1 U18936 ( .IN1(n17176), .IN2(g629), .Q(n17978) );
  AND2X1 U18937 ( .IN1(n17979), .IN2(n17980), .Q(n17176) );
  AND2X1 U18938 ( .IN1(n9351), .IN2(n9352), .Q(n17980) );
  AND2X1 U18939 ( .IN1(n10163), .IN2(n17981), .Q(n17979) );
  AND2X1 U18940 ( .IN1(n10197), .IN2(n10164), .Q(n17981) );
  AND2X1 U18941 ( .IN1(n4295), .IN2(g659), .Q(n17977) );
  OR2X1 U18942 ( .IN1(n17982), .IN2(n17983), .Q(g20310) );
  AND2X1 U18943 ( .IN1(n4351), .IN2(g2972), .Q(n17983) );
  AND2X1 U18944 ( .IN1(g2879), .IN2(g6225), .Q(n17982) );
  OR2X1 U18945 ( .IN1(n17984), .IN2(n17985), .Q(g19184) );
  AND2X1 U18946 ( .IN1(n4351), .IN2(g2975), .Q(n17985) );
  AND2X1 U18947 ( .IN1(g2879), .IN2(g4590), .Q(n17984) );
  OR2X1 U18948 ( .IN1(n17986), .IN2(n17987), .Q(g19178) );
  AND2X1 U18949 ( .IN1(n4351), .IN2(g2935), .Q(n17987) );
  AND2X1 U18950 ( .IN1(test_so5), .IN2(g2879), .Q(n17986) );
  OR2X1 U18951 ( .IN1(n17988), .IN2(n17989), .Q(g19173) );
  AND2X1 U18952 ( .IN1(n4351), .IN2(g2978), .Q(n17989) );
  AND2X1 U18953 ( .IN1(g2879), .IN2(g4323), .Q(n17988) );
  OR2X1 U18954 ( .IN1(n17990), .IN2(n17991), .Q(g19172) );
  AND2X1 U18955 ( .IN1(n4351), .IN2(g2953), .Q(n17991) );
  AND2X1 U18956 ( .IN1(g2879), .IN2(g4321), .Q(n17990) );
  OR2X1 U18957 ( .IN1(n17992), .IN2(n17993), .Q(g19167) );
  AND2X1 U18958 ( .IN1(n4351), .IN2(g2938), .Q(n17993) );
  AND2X1 U18959 ( .IN1(g2879), .IN2(g4200), .Q(n17992) );
  OR2X1 U18960 ( .IN1(n17994), .IN2(n17995), .Q(g19163) );
  AND2X1 U18961 ( .IN1(n4351), .IN2(g2981), .Q(n17995) );
  AND2X1 U18962 ( .IN1(g2879), .IN2(g4090), .Q(n17994) );
  OR2X1 U18963 ( .IN1(n17996), .IN2(n17997), .Q(g19162) );
  AND2X1 U18964 ( .IN1(n4351), .IN2(g2956), .Q(n17997) );
  AND2X1 U18965 ( .IN1(g2879), .IN2(g4088), .Q(n17996) );
  OR2X1 U18966 ( .IN1(n17998), .IN2(n17999), .Q(g19157) );
  AND2X1 U18967 ( .IN1(n4351), .IN2(g2941), .Q(n17999) );
  AND2X1 U18968 ( .IN1(g2879), .IN2(g3993), .Q(n17998) );
  OR2X1 U18969 ( .IN1(n18000), .IN2(n18001), .Q(g19154) );
  AND2X1 U18970 ( .IN1(n4351), .IN2(g2874), .Q(n18001) );
  AND2X1 U18971 ( .IN1(test_so3), .IN2(g2879), .Q(n18000) );
  OR2X1 U18972 ( .IN1(n18002), .IN2(n18003), .Q(g19153) );
  AND2X1 U18973 ( .IN1(n4351), .IN2(g2959), .Q(n18003) );
  AND2X1 U18974 ( .IN1(g2879), .IN2(g8249), .Q(n18002) );
  OR2X1 U18975 ( .IN1(n18004), .IN2(n18005), .Q(g19149) );
  AND2X1 U18976 ( .IN1(n4351), .IN2(g2944), .Q(n18005) );
  AND2X1 U18977 ( .IN1(g2879), .IN2(g8175), .Q(n18004) );
  OR2X1 U18978 ( .IN1(n18006), .IN2(n18007), .Q(g19144) );
  AND2X1 U18979 ( .IN1(n4351), .IN2(g2947), .Q(n18007) );
  AND2X1 U18980 ( .IN1(g2879), .IN2(g8023), .Q(n18006) );
  OR2X1 U18981 ( .IN1(n18008), .IN2(n18009), .Q(g18975) );
  AND2X1 U18982 ( .IN1(g2981), .IN2(g2879), .Q(n18009) );
  AND2X1 U18983 ( .IN1(n4351), .IN2(g2195), .Q(n18008) );
  OR2X1 U18984 ( .IN1(n18010), .IN2(n18011), .Q(g18968) );
  AND2X1 U18985 ( .IN1(g2978), .IN2(g2879), .Q(n18011) );
  AND2X1 U18986 ( .IN1(n4351), .IN2(g2190), .Q(n18010) );
  OR2X1 U18987 ( .IN1(n18012), .IN2(n18013), .Q(g18957) );
  AND2X1 U18988 ( .IN1(g2963), .IN2(g2879), .Q(n18013) );
  AND2X1 U18989 ( .IN1(n4351), .IN2(g2165), .Q(n18012) );
  OR2X1 U18990 ( .IN1(n18014), .IN2(n18015), .Q(g18942) );
  AND2X1 U18991 ( .IN1(g2975), .IN2(g2879), .Q(n18015) );
  AND2X1 U18992 ( .IN1(n4351), .IN2(g2185), .Q(n18014) );
  OR2X1 U18993 ( .IN1(n18016), .IN2(n18017), .Q(g18907) );
  AND2X1 U18994 ( .IN1(g2987), .IN2(g2997), .Q(n18017) );
  AND2X1 U18995 ( .IN1(n4365), .IN2(g3061), .Q(n18016) );
  OR2X1 U18996 ( .IN1(n18018), .IN2(n18019), .Q(g18906) );
  AND2X1 U18997 ( .IN1(g2972), .IN2(g2879), .Q(n18019) );
  AND2X1 U18998 ( .IN1(n4351), .IN2(g2180), .Q(n18018) );
  OR2X1 U18999 ( .IN1(n18020), .IN2(n18021), .Q(g18885) );
  AND2X1 U19000 ( .IN1(g2874), .IN2(g2879), .Q(n18021) );
  AND2X1 U19001 ( .IN1(n4351), .IN2(g2200), .Q(n18020) );
  OR2X1 U19002 ( .IN1(n18022), .IN2(n18023), .Q(g18883) );
  AND2X1 U19003 ( .IN1(g2935), .IN2(g2879), .Q(n18023) );
  AND2X1 U19004 ( .IN1(n4351), .IN2(g1471), .Q(n18022) );
  OR2X1 U19005 ( .IN1(n18024), .IN2(n18025), .Q(g18868) );
  AND2X1 U19006 ( .IN1(g2987), .IN2(g3078), .Q(n18025) );
  AND2X1 U19007 ( .IN1(n4365), .IN2(g3060), .Q(n18024) );
  OR2X1 U19008 ( .IN1(n18026), .IN2(n18027), .Q(g18867) );
  AND2X1 U19009 ( .IN1(g2969), .IN2(g2879), .Q(n18027) );
  AND2X1 U19010 ( .IN1(n4351), .IN2(g2175), .Q(n18026) );
  OR2X1 U19011 ( .IN1(n18028), .IN2(n18029), .Q(g18866) );
  AND2X1 U19012 ( .IN1(g2938), .IN2(g2879), .Q(n18029) );
  AND2X1 U19013 ( .IN1(n4351), .IN2(g1476), .Q(n18028) );
  OR2X1 U19014 ( .IN1(n18030), .IN2(n18031), .Q(g18852) );
  AND2X1 U19015 ( .IN1(g2941), .IN2(g2879), .Q(n18031) );
  AND2X1 U19016 ( .IN1(n4351), .IN2(g1481), .Q(n18030) );
  OR2X1 U19017 ( .IN1(n18032), .IN2(n18033), .Q(g18837) );
  AND2X1 U19018 ( .IN1(g2987), .IN2(g3077), .Q(n18033) );
  AND2X1 U19019 ( .IN1(n4365), .IN2(g3059), .Q(n18032) );
  OR2X1 U19020 ( .IN1(n18034), .IN2(n18035), .Q(g18836) );
  AND2X1 U19021 ( .IN1(test_so2), .IN2(g2879), .Q(n18035) );
  AND2X1 U19022 ( .IN1(n4351), .IN2(g2170), .Q(n18034) );
  OR2X1 U19023 ( .IN1(n18036), .IN2(n18037), .Q(g18835) );
  AND2X1 U19024 ( .IN1(g2944), .IN2(g2879), .Q(n18037) );
  AND2X1 U19025 ( .IN1(n4351), .IN2(g1486), .Q(n18036) );
  OR2X1 U19026 ( .IN1(n18038), .IN2(n18039), .Q(g18821) );
  AND2X1 U19027 ( .IN1(g2947), .IN2(g2879), .Q(n18039) );
  AND2X1 U19028 ( .IN1(n4351), .IN2(g1491), .Q(n18038) );
  OR2X1 U19029 ( .IN1(n18040), .IN2(n18041), .Q(g18820) );
  AND2X1 U19030 ( .IN1(g2624), .IN2(g2631), .Q(n18041) );
  AND2X1 U19031 ( .IN1(n4299), .IN2(g2584), .Q(n18040) );
  OR2X1 U19032 ( .IN1(n18042), .IN2(n18043), .Q(g18804) );
  AND2X1 U19033 ( .IN1(g2987), .IN2(g3076), .Q(n18043) );
  AND2X1 U19034 ( .IN1(n4365), .IN2(g3058), .Q(n18042) );
  OR2X1 U19035 ( .IN1(n18044), .IN2(n18045), .Q(g18803) );
  AND2X1 U19036 ( .IN1(g2953), .IN2(g2879), .Q(n18045) );
  AND2X1 U19037 ( .IN1(n4351), .IN2(g1496), .Q(n18044) );
  OR2X1 U19038 ( .IN1(n18046), .IN2(n18047), .Q(g18794) );
  AND2X1 U19039 ( .IN1(n4366), .IN2(g1890), .Q(n18047) );
  AND2X1 U19040 ( .IN1(g1937), .IN2(g1930), .Q(n18046) );
  OR2X1 U19041 ( .IN1(n18048), .IN2(n18049), .Q(g18782) );
  AND2X1 U19042 ( .IN1(n4494), .IN2(g3084), .Q(n18049) );
  AND2X1 U19043 ( .IN1(g3109), .IN2(g559), .Q(n18048) );
  OR2X1 U19044 ( .IN1(n18050), .IN2(n18051), .Q(g18781) );
  AND2X1 U19045 ( .IN1(g2956), .IN2(g2879), .Q(n18051) );
  AND2X1 U19046 ( .IN1(n4351), .IN2(g1501), .Q(n18050) );
  OR2X1 U19047 ( .IN1(n18052), .IN2(n18053), .Q(g18780) );
  AND2X1 U19048 ( .IN1(n10120), .IN2(g2624), .Q(n18053) );
  AND2X1 U19049 ( .IN1(n4299), .IN2(g2631), .Q(n18052) );
  OR2X1 U19050 ( .IN1(n18054), .IN2(n18055), .Q(g18763) );
  AND2X1 U19051 ( .IN1(g1236), .IN2(g1243), .Q(n18055) );
  AND2X1 U19052 ( .IN1(n4300), .IN2(g1196), .Q(n18054) );
  OR2X1 U19053 ( .IN1(n18056), .IN2(n18057), .Q(g18755) );
  AND2X1 U19054 ( .IN1(g2987), .IN2(g3075), .Q(n18057) );
  AND2X1 U19055 ( .IN1(n4365), .IN2(g3057), .Q(n18056) );
  OR2X1 U19056 ( .IN1(n18058), .IN2(n18059), .Q(g18754) );
  AND2X1 U19057 ( .IN1(g2959), .IN2(g2879), .Q(n18059) );
  AND2X1 U19058 ( .IN1(n4351), .IN2(g1506), .Q(n18058) );
  OR2X1 U19059 ( .IN1(n18060), .IN2(n18061), .Q(g18743) );
  AND2X1 U19060 ( .IN1(n10121), .IN2(g1930), .Q(n18061) );
  AND2X1 U19061 ( .IN1(n4366), .IN2(g1937), .Q(n18060) );
  OR2X1 U19062 ( .IN1(n18062), .IN2(n18063), .Q(g18726) );
  AND2X1 U19063 ( .IN1(g550), .IN2(g557), .Q(n18063) );
  AND2X1 U19064 ( .IN1(n4313), .IN2(test_so22), .Q(n18062) );
  OR2X1 U19065 ( .IN1(n18064), .IN2(n18065), .Q(g18719) );
  AND2X1 U19066 ( .IN1(g8030), .IN2(g559), .Q(n18065) );
  AND2X1 U19067 ( .IN1(n4383), .IN2(g3211), .Q(n18064) );
  OR2X1 U19068 ( .IN1(n18066), .IN2(n18067), .Q(g18707) );
  AND2X1 U19069 ( .IN1(n10122), .IN2(g1236), .Q(n18067) );
  AND2X1 U19070 ( .IN1(n4300), .IN2(g1243), .Q(n18066) );
  OR2X1 U19071 ( .IN1(n18068), .IN2(n18069), .Q(g18678) );
  AND2X1 U19072 ( .IN1(n10123), .IN2(g550), .Q(n18069) );
  AND2X1 U19073 ( .IN1(n4313), .IN2(g557), .Q(n18068) );
  OR2X1 U19074 ( .IN1(n18070), .IN2(n18071), .Q(g18669) );
  AND2X1 U19075 ( .IN1(g8106), .IN2(g559), .Q(n18071) );
  AND2X1 U19076 ( .IN1(n4382), .IN2(test_so6), .Q(n18070) );
  OR2X1 U19077 ( .IN1(n18072), .IN2(n18073), .Q(g17429) );
  AND2X1 U19078 ( .IN1(n4494), .IN2(g3088), .Q(n18073) );
  AND2X1 U19079 ( .IN1(g3109), .IN2(g2574), .Q(n18072) );
  OR2X1 U19080 ( .IN1(n18074), .IN2(n18075), .Q(g17383) );
  AND2X1 U19081 ( .IN1(g3109), .IN2(g1880), .Q(n18075) );
  AND2X1 U19082 ( .IN1(n4494), .IN2(test_so8), .Q(n18074) );
  OR2X1 U19083 ( .IN1(n18076), .IN2(n18077), .Q(g17341) );
  AND2X1 U19084 ( .IN1(g8030), .IN2(g2574), .Q(n18077) );
  AND2X1 U19085 ( .IN1(n4383), .IN2(g3185), .Q(n18076) );
  OR2X1 U19086 ( .IN1(n18078), .IN2(n18079), .Q(g17340) );
  AND2X1 U19087 ( .IN1(n4494), .IN2(g3170), .Q(n18079) );
  AND2X1 U19088 ( .IN1(g3109), .IN2(g1186), .Q(n18078) );
  OR2X1 U19089 ( .IN1(n18080), .IN2(n18081), .Q(g17303) );
  AND2X1 U19090 ( .IN1(g8030), .IN2(g1880), .Q(n18081) );
  AND2X1 U19091 ( .IN1(n4383), .IN2(g3176), .Q(n18080) );
  OR2X1 U19092 ( .IN1(n18082), .IN2(n18083), .Q(g17302) );
  AND2X1 U19093 ( .IN1(n4494), .IN2(g3161), .Q(n18083) );
  AND2X1 U19094 ( .IN1(g3109), .IN2(g499), .Q(n18082) );
  OR2X1 U19095 ( .IN1(n18084), .IN2(n18085), .Q(g17271) );
  AND2X1 U19096 ( .IN1(g8106), .IN2(g2574), .Q(n18085) );
  AND2X1 U19097 ( .IN1(n4382), .IN2(g3182), .Q(n18084) );
  OR2X1 U19098 ( .IN1(n18086), .IN2(n18087), .Q(g17270) );
  AND2X1 U19099 ( .IN1(n4383), .IN2(g3167), .Q(n18087) );
  AND2X1 U19100 ( .IN1(g8030), .IN2(g1186), .Q(n18086) );
  OR2X1 U19101 ( .IN1(n18088), .IN2(n18089), .Q(g17269) );
  AND2X1 U19102 ( .IN1(n4494), .IN2(g3096), .Q(n18089) );
  AND2X1 U19103 ( .IN1(g3109), .IN2(g2633), .Q(n18088) );
  OR2X1 U19104 ( .IN1(n18090), .IN2(n18091), .Q(g17248) );
  AND2X1 U19105 ( .IN1(n4382), .IN2(g3173), .Q(n18091) );
  AND2X1 U19106 ( .IN1(g8106), .IN2(g1880), .Q(n18090) );
  OR2X1 U19107 ( .IN1(n18092), .IN2(n18093), .Q(g17247) );
  AND2X1 U19108 ( .IN1(g8030), .IN2(g499), .Q(n18093) );
  AND2X1 U19109 ( .IN1(n4383), .IN2(g3158), .Q(n18092) );
  OR2X1 U19110 ( .IN1(n18094), .IN2(n18095), .Q(g17246) );
  AND2X1 U19111 ( .IN1(n4494), .IN2(g3093), .Q(n18095) );
  AND2X1 U19112 ( .IN1(g3109), .IN2(g1939), .Q(n18094) );
  OR2X1 U19113 ( .IN1(n18096), .IN2(n18097), .Q(g17236) );
  AND2X1 U19114 ( .IN1(n4382), .IN2(g3164), .Q(n18097) );
  AND2X1 U19115 ( .IN1(g8106), .IN2(g1186), .Q(n18096) );
  OR2X1 U19116 ( .IN1(n18098), .IN2(n18099), .Q(g17235) );
  AND2X1 U19117 ( .IN1(g8030), .IN2(g2633), .Q(n18099) );
  AND2X1 U19118 ( .IN1(n4383), .IN2(g3095), .Q(n18098) );
  OR2X1 U19119 ( .IN1(n18100), .IN2(n18101), .Q(g17234) );
  AND2X1 U19120 ( .IN1(n4494), .IN2(g3087), .Q(n18101) );
  AND2X1 U19121 ( .IN1(g3109), .IN2(g1245), .Q(n18100) );
  OR2X1 U19122 ( .IN1(n18102), .IN2(n18103), .Q(g17229) );
  AND2X1 U19123 ( .IN1(g8106), .IN2(g499), .Q(n18103) );
  AND2X1 U19124 ( .IN1(n4382), .IN2(g3155), .Q(n18102) );
  OR2X1 U19125 ( .IN1(n18104), .IN2(n18105), .Q(g17228) );
  AND2X1 U19126 ( .IN1(g8030), .IN2(g1939), .Q(n18105) );
  AND2X1 U19127 ( .IN1(n4383), .IN2(g3092), .Q(n18104) );
  OR2X1 U19128 ( .IN1(n18106), .IN2(n18107), .Q(g17226) );
  AND2X1 U19129 ( .IN1(g8106), .IN2(g2633), .Q(n18107) );
  AND2X1 U19130 ( .IN1(n4382), .IN2(g3094), .Q(n18106) );
  OR2X1 U19131 ( .IN1(n18108), .IN2(n18109), .Q(g17225) );
  AND2X1 U19132 ( .IN1(n4383), .IN2(g3086), .Q(n18109) );
  AND2X1 U19133 ( .IN1(g8030), .IN2(g1245), .Q(n18108) );
  OR2X1 U19134 ( .IN1(n18110), .IN2(n18111), .Q(g17224) );
  AND2X1 U19135 ( .IN1(g8106), .IN2(g1939), .Q(n18111) );
  AND2X1 U19136 ( .IN1(n4382), .IN2(g3091), .Q(n18110) );
  OR2X1 U19137 ( .IN1(n18112), .IN2(n18113), .Q(g17222) );
  AND2X1 U19138 ( .IN1(n4382), .IN2(g3085), .Q(n18113) );
  AND2X1 U19139 ( .IN1(g8106), .IN2(g1245), .Q(n18112) );
  OR2X1 U19140 ( .IN1(n18114), .IN2(n18115), .Q(g16880) );
  AND2X1 U19141 ( .IN1(g2987), .IN2(g3074), .Q(n18115) );
  AND2X1 U19142 ( .IN1(n4365), .IN2(g3056), .Q(n18114) );
  OR2X1 U19143 ( .IN1(n18116), .IN2(n18117), .Q(g16866) );
  AND2X1 U19144 ( .IN1(test_so97), .IN2(g2987), .Q(n18117) );
  AND2X1 U19145 ( .IN1(n4365), .IN2(g3051), .Q(n18116) );
  OR2X1 U19146 ( .IN1(n18118), .IN2(n18119), .Q(g16861) );
  AND2X1 U19147 ( .IN1(g2987), .IN2(g3073), .Q(n18119) );
  AND2X1 U19148 ( .IN1(test_so96), .IN2(n4365), .Q(n18118) );
  OR2X1 U19149 ( .IN1(n18120), .IN2(n18121), .Q(g16860) );
  AND2X1 U19150 ( .IN1(g2987), .IN2(g3065), .Q(n18121) );
  AND2X1 U19151 ( .IN1(n4365), .IN2(g3046), .Q(n18120) );
  OR2X1 U19152 ( .IN1(n18122), .IN2(n18123), .Q(g16857) );
  AND2X1 U19153 ( .IN1(g2987), .IN2(g3069), .Q(n18123) );
  AND2X1 U19154 ( .IN1(n4365), .IN2(g3050), .Q(n18122) );
  OR2X1 U19155 ( .IN1(n18124), .IN2(n18125), .Q(g16854) );
  AND2X1 U19156 ( .IN1(g2987), .IN2(g3072), .Q(n18125) );
  AND2X1 U19157 ( .IN1(n4365), .IN2(g3053), .Q(n18124) );
  OR2X1 U19158 ( .IN1(n18126), .IN2(n18127), .Q(g16853) );
  AND2X1 U19159 ( .IN1(g2987), .IN2(g3064), .Q(n18127) );
  AND2X1 U19160 ( .IN1(n4365), .IN2(g3045), .Q(n18126) );
  OR2X1 U19161 ( .IN1(n18128), .IN2(n18129), .Q(g16851) );
  AND2X1 U19162 ( .IN1(g2987), .IN2(g3068), .Q(n18129) );
  AND2X1 U19163 ( .IN1(n4365), .IN2(g3049), .Q(n18128) );
  OR2X1 U19164 ( .IN1(n18130), .IN2(n18131), .Q(g16845) );
  AND2X1 U19165 ( .IN1(g2987), .IN2(g3071), .Q(n18131) );
  AND2X1 U19166 ( .IN1(n4365), .IN2(g3052), .Q(n18130) );
  OR2X1 U19167 ( .IN1(n18132), .IN2(n18133), .Q(g16844) );
  AND2X1 U19168 ( .IN1(g2987), .IN2(g3063), .Q(n18133) );
  AND2X1 U19169 ( .IN1(n4365), .IN2(g3044), .Q(n18132) );
  OR2X1 U19170 ( .IN1(n18134), .IN2(n18135), .Q(g16835) );
  AND2X1 U19171 ( .IN1(g2987), .IN2(g3067), .Q(n18135) );
  AND2X1 U19172 ( .IN1(n4365), .IN2(g3048), .Q(n18134) );
  OR2X1 U19173 ( .IN1(n18136), .IN2(n18137), .Q(g16824) );
  AND2X1 U19174 ( .IN1(g2987), .IN2(g3062), .Q(n18137) );
  AND2X1 U19175 ( .IN1(n4365), .IN2(g3043), .Q(n18136) );
  AND2X1 U19176 ( .IN1(n18138), .IN2(n8103), .Q(g16823) );
  OR2X1 U19177 ( .IN1(n18139), .IN2(n18140), .Q(g16803) );
  AND2X1 U19178 ( .IN1(g2987), .IN2(g3066), .Q(n18140) );
  AND2X1 U19179 ( .IN1(n4365), .IN2(g3047), .Q(n18139) );
  AND2X1 U19180 ( .IN1(n18138), .IN2(g2950), .Q(g16802) );
  INVX0 U19181 ( .INP(g51), .ZN(n18138) );
  OR2X1 U19182 ( .IN1(n18141), .IN2(n18142), .Q(g16718) );
  INVX0 U19183 ( .INP(n18143), .ZN(n18142) );
  OR2X1 U19184 ( .IN1(g2703), .IN2(n10156), .Q(n18143) );
  AND2X1 U19185 ( .IN1(g2703), .IN2(g2584), .Q(n18141) );
  OR2X1 U19186 ( .IN1(n18144), .IN2(n18145), .Q(g16692) );
  INVX0 U19187 ( .INP(n18146), .ZN(n18145) );
  OR2X1 U19188 ( .IN1(g2009), .IN2(n10155), .Q(n18146) );
  AND2X1 U19189 ( .IN1(g2009), .IN2(g1890), .Q(n18144) );
  OR2X1 U19190 ( .IN1(n18147), .IN2(n18148), .Q(g16671) );
  INVX0 U19191 ( .INP(n18149), .ZN(n18148) );
  OR2X1 U19192 ( .IN1(g1315), .IN2(n10154), .Q(n18149) );
  AND2X1 U19193 ( .IN1(g1315), .IN2(g1196), .Q(n18147) );
  OR2X1 U19194 ( .IN1(n18150), .IN2(n18151), .Q(g16654) );
  INVX0 U19195 ( .INP(n18152), .ZN(n18151) );
  OR2X1 U19196 ( .IN1(g629), .IN2(n10153), .Q(n18152) );
  AND2X1 U19197 ( .IN1(test_so22), .IN2(g629), .Q(n18150) );
  OR2X1 U19198 ( .IN1(n4365), .IN2(n18153), .Q(g16496) );
  AND2X1 U19199 ( .IN1(DFF_1612_n1), .IN2(g5388), .Q(n18153) );
  AND2X1 U19200 ( .IN1(n18154), .IN2(n18155), .Q(g13194) );
  OR2X1 U19201 ( .IN1(n4370), .IN2(g2561), .Q(n18155) );
  AND2X1 U19202 ( .IN1(n18156), .IN2(n18157), .Q(n18154) );
  OR2X1 U19203 ( .IN1(n4299), .IN2(g2562), .Q(n18157) );
  OR2X1 U19204 ( .IN1(n4314), .IN2(test_so87), .Q(n18156) );
  AND2X1 U19205 ( .IN1(n18158), .IN2(n18159), .Q(g13182) );
  OR2X1 U19206 ( .IN1(n4315), .IN2(g1867), .Q(n18159) );
  AND2X1 U19207 ( .IN1(n18160), .IN2(n18161), .Q(n18158) );
  OR2X1 U19208 ( .IN1(n4366), .IN2(g1868), .Q(n18161) );
  OR2X1 U19209 ( .IN1(n4296), .IN2(g1869), .Q(n18160) );
  AND2X1 U19210 ( .IN1(n18162), .IN2(n18163), .Q(g13175) );
  OR2X1 U19211 ( .IN1(n4370), .IN2(g2552), .Q(n18163) );
  AND2X1 U19212 ( .IN1(n18164), .IN2(n18165), .Q(n18162) );
  OR2X1 U19213 ( .IN1(n4299), .IN2(g2553), .Q(n18165) );
  OR2X1 U19214 ( .IN1(n4314), .IN2(g2554), .Q(n18164) );
  AND2X1 U19215 ( .IN1(n18166), .IN2(n18167), .Q(g13171) );
  OR2X1 U19216 ( .IN1(n4316), .IN2(g1173), .Q(n18167) );
  AND2X1 U19217 ( .IN1(n18168), .IN2(n18169), .Q(n18166) );
  OR2X1 U19218 ( .IN1(n4371), .IN2(g1175), .Q(n18169) );
  OR2X1 U19219 ( .IN1(n4300), .IN2(test_so44), .Q(n18168) );
  AND2X1 U19220 ( .IN1(n18170), .IN2(n18171), .Q(g13164) );
  OR2X1 U19221 ( .IN1(n4315), .IN2(g1858), .Q(n18171) );
  AND2X1 U19222 ( .IN1(n18172), .IN2(n18173), .Q(n18170) );
  OR2X1 U19223 ( .IN1(n4366), .IN2(g1859), .Q(n18173) );
  OR2X1 U19224 ( .IN1(n4296), .IN2(g1860), .Q(n18172) );
  AND2X1 U19225 ( .IN1(n18174), .IN2(n18175), .Q(g13160) );
  OR2X1 U19226 ( .IN1(n4372), .IN2(g486), .Q(n18175) );
  AND2X1 U19227 ( .IN1(n18176), .IN2(n18177), .Q(n18174) );
  OR2X1 U19228 ( .IN1(n4313), .IN2(g487), .Q(n18177) );
  OR2X1 U19229 ( .IN1(n4298), .IN2(g488), .Q(n18176) );
  AND2X1 U19230 ( .IN1(n18178), .IN2(n18179), .Q(g13155) );
  OR2X1 U19231 ( .IN1(n4316), .IN2(g1164), .Q(n18179) );
  AND2X1 U19232 ( .IN1(n18180), .IN2(n18181), .Q(n18178) );
  OR2X1 U19233 ( .IN1(n4300), .IN2(g1165), .Q(n18181) );
  OR2X1 U19234 ( .IN1(n4371), .IN2(g1166), .Q(n18180) );
  AND2X1 U19235 ( .IN1(n18182), .IN2(n18183), .Q(g13149) );
  OR2X1 U19236 ( .IN1(n4372), .IN2(g477), .Q(n18183) );
  AND2X1 U19237 ( .IN1(n18184), .IN2(n18185), .Q(n18182) );
  OR2X1 U19238 ( .IN1(n4313), .IN2(g478), .Q(n18185) );
  OR2X1 U19239 ( .IN1(n4298), .IN2(g479), .Q(n18184) );
  AND2X1 U19240 ( .IN1(n18186), .IN2(n18187), .Q(g13143) );
  OR2X1 U19241 ( .IN1(n4370), .IN2(g2555), .Q(n18187) );
  AND2X1 U19242 ( .IN1(n18188), .IN2(n18189), .Q(n18186) );
  OR2X1 U19243 ( .IN1(n4299), .IN2(g2559), .Q(n18189) );
  OR2X1 U19244 ( .IN1(n4314), .IN2(g2539), .Q(n18188) );
  AND2X1 U19245 ( .IN1(n18190), .IN2(n18191), .Q(g13135) );
  OR2X1 U19246 ( .IN1(n4315), .IN2(g1861), .Q(n18191) );
  AND2X1 U19247 ( .IN1(n18192), .IN2(n18193), .Q(n18190) );
  OR2X1 U19248 ( .IN1(n4366), .IN2(g1865), .Q(n18193) );
  OR2X1 U19249 ( .IN1(n4296), .IN2(g1845), .Q(n18192) );
  AND2X1 U19250 ( .IN1(n18194), .IN2(n18195), .Q(g13124) );
  OR2X1 U19251 ( .IN1(n4316), .IN2(g1167), .Q(n18195) );
  AND2X1 U19252 ( .IN1(n18196), .IN2(n18197), .Q(n18194) );
  OR2X1 U19253 ( .IN1(n4300), .IN2(g1171), .Q(n18197) );
  OR2X1 U19254 ( .IN1(n4371), .IN2(g1151), .Q(n18196) );
  AND2X1 U19255 ( .IN1(n18198), .IN2(n18199), .Q(g13111) );
  OR2X1 U19256 ( .IN1(n4372), .IN2(g480), .Q(n18199) );
  AND2X1 U19257 ( .IN1(n18200), .IN2(n18201), .Q(n18198) );
  OR2X1 U19258 ( .IN1(n4313), .IN2(g484), .Q(n18201) );
  OR2X1 U19259 ( .IN1(n4298), .IN2(g464), .Q(n18200) );
  OR2X1 U19260 ( .IN1(n18202), .IN2(n18203), .Q(N995) );
  INVX0 U19261 ( .INP(n18204), .ZN(n18203) );
  OR2X1 U19262 ( .IN1(n10938), .IN2(n10149), .Q(n18204) );
  AND2X1 U19263 ( .IN1(n10149), .IN2(n10938), .Q(n18202) );
  AND2X1 U19264 ( .IN1(n18205), .IN2(n18206), .Q(n10938) );
  INVX0 U19265 ( .INP(n18207), .ZN(n18206) );
  AND2X1 U19266 ( .IN1(n18208), .IN2(n18209), .Q(n18207) );
  OR2X1 U19267 ( .IN1(n18209), .IN2(n18208), .Q(n18205) );
  OR2X1 U19268 ( .IN1(n18210), .IN2(n18211), .Q(n18208) );
  INVX0 U19269 ( .INP(n18212), .ZN(n18211) );
  OR2X1 U19270 ( .IN1(n18213), .IN2(n18214), .Q(n18212) );
  AND2X1 U19271 ( .IN1(n18214), .IN2(n18213), .Q(n18210) );
  AND2X1 U19272 ( .IN1(n18215), .IN2(n18216), .Q(n18213) );
  INVX0 U19273 ( .INP(n18217), .ZN(n18216) );
  AND2X1 U19274 ( .IN1(n10144), .IN2(g8271), .Q(n18217) );
  OR2X1 U19275 ( .IN1(g8271), .IN2(n10144), .Q(n18215) );
  OR2X1 U19276 ( .IN1(n18218), .IN2(n18219), .Q(n18214) );
  AND2X1 U19277 ( .IN1(n10146), .IN2(g8269), .Q(n18219) );
  AND2X1 U19278 ( .IN1(n10147), .IN2(g8274), .Q(n18218) );
  AND2X1 U19279 ( .IN1(n18220), .IN2(n18221), .Q(n18209) );
  INVX0 U19280 ( .INP(n18222), .ZN(n18221) );
  AND2X1 U19281 ( .IN1(n18223), .IN2(n18224), .Q(n18222) );
  OR2X1 U19282 ( .IN1(n18224), .IN2(n18223), .Q(n18220) );
  OR2X1 U19283 ( .IN1(n18225), .IN2(n18226), .Q(n18223) );
  AND2X1 U19284 ( .IN1(n18265), .IN2(g8268), .Q(n18226) );
  AND2X1 U19285 ( .IN1(n18264), .IN2(g8273), .Q(n18225) );
  INVX0 U19286 ( .INP(n18227), .ZN(n18224) );
  OR2X1 U19287 ( .IN1(n18228), .IN2(n18229), .Q(n18227) );
  AND2X1 U19288 ( .IN1(n18259), .IN2(n10205), .Q(n18229) );
  AND2X1 U19289 ( .IN1(test_so99), .IN2(g8272), .Q(n18228) );
  AND2X1 U19290 ( .IN1(n18230), .IN2(n18231), .Q(N690) );
  INVX0 U19291 ( .INP(n18232), .ZN(n18231) );
  AND2X1 U19292 ( .IN1(n10943), .IN2(n10151), .Q(n18232) );
  OR2X1 U19293 ( .IN1(n10151), .IN2(n10943), .Q(n18230) );
  AND2X1 U19294 ( .IN1(n18233), .IN2(n18234), .Q(n10943) );
  INVX0 U19295 ( .INP(n18235), .ZN(n18234) );
  AND2X1 U19296 ( .IN1(n18236), .IN2(n18237), .Q(n18235) );
  OR2X1 U19297 ( .IN1(n18237), .IN2(n18236), .Q(n18233) );
  OR2X1 U19298 ( .IN1(n18238), .IN2(n18239), .Q(n18236) );
  INVX0 U19299 ( .INP(n18240), .ZN(n18239) );
  OR2X1 U19300 ( .IN1(n18241), .IN2(n18242), .Q(n18240) );
  AND2X1 U19301 ( .IN1(n18242), .IN2(n18241), .Q(n18238) );
  AND2X1 U19302 ( .IN1(n18243), .IN2(n18244), .Q(n18241) );
  INVX0 U19303 ( .INP(n18245), .ZN(n18244) );
  AND2X1 U19304 ( .IN1(n10124), .IN2(g8261), .Q(n18245) );
  OR2X1 U19305 ( .IN1(g8261), .IN2(n10124), .Q(n18243) );
  OR2X1 U19306 ( .IN1(n18246), .IN2(n18247), .Q(n18242) );
  AND2X1 U19307 ( .IN1(n10126), .IN2(g8264), .Q(n18247) );
  AND2X1 U19308 ( .IN1(n10127), .IN2(g8259), .Q(n18246) );
  AND2X1 U19309 ( .IN1(n18248), .IN2(n18249), .Q(n18237) );
  INVX0 U19310 ( .INP(n18250), .ZN(n18249) );
  AND2X1 U19311 ( .IN1(n18251), .IN2(n18252), .Q(n18250) );
  OR2X1 U19312 ( .IN1(n18252), .IN2(n18251), .Q(n18248) );
  OR2X1 U19313 ( .IN1(n18253), .IN2(n18254), .Q(n18251) );
  AND2X1 U19314 ( .IN1(n10128), .IN2(g8266), .Q(n18254) );
  AND2X1 U19315 ( .IN1(n18267), .IN2(g8263), .Q(n18253) );
  INVX0 U19316 ( .INP(n18255), .ZN(n18252) );
  OR2X1 U19317 ( .IN1(n18256), .IN2(n18257), .Q(n18255) );
  AND2X1 U19318 ( .IN1(n18266), .IN2(g8265), .Q(n18257) );
  AND2X1 U19319 ( .IN1(n18260), .IN2(g8262), .Q(n18256) );
  OR2X1 U3772_U1 ( .IN1(n2230), .IN2(n2217), .Q(n2231) );
  OR2X1 U3776_U1 ( .IN1(n2374), .IN2(n2361), .Q(n2375) );
  OR2X1 U3777_U1 ( .IN1(g51), .IN2(DFF_2_n1), .Q(n4264) );
  OR2X1 U3778_U1 ( .IN1(n2445), .IN2(n2446), .Q(n2440) );
  OR2X1 U3779_U1 ( .IN1(n549), .IN2(n2446), .Q(n2426) );
  OR2X1 U3780_U1 ( .IN1(n2670), .IN2(n2671), .Q(n2669) );
  OR2X1 U3781_U1 ( .IN1(n2685), .IN2(n2686), .Q(n2684) );
  OR2X1 U3782_U1 ( .IN1(n2718), .IN2(n2719), .Q(n2717) );
  OR2X1 U3783_U1 ( .IN1(n1577), .IN2(g2124), .Q(n2981) );
  OR2X1 U3784_U1 ( .IN1(n1233), .IN2(g1430), .Q(n2984) );
  OR2X1 U3785_U1 ( .IN1(n888), .IN2(g744), .Q(n2987) );
  OR2X1 U3786_U1 ( .IN1(n470), .IN2(g56), .Q(n2990) );
  OR2X1 U3787_U1 ( .IN1(n1808), .IN2(test_so98), .Q(n3741) );
  OR2X1 U3901_U1 ( .IN1(n2302), .IN2(n2289), .Q(n2303) );
  OR2X1 U3902_U1 ( .IN1(n580), .IN2(n2289), .Q(n2275) );
  INVX0 U4467_U2 ( .INP(n3254), .ZN(U4467_n1) );
  AND2X1 U4467_U1 ( .IN1(n1636), .IN2(U4467_n1), .Q(n3252) );
  INVX0 U4904_U2 ( .INP(n2617), .ZN(U4904_n1) );
  AND2X1 U4904_U1 ( .IN1(n2800), .IN2(U4904_n1), .Q(n2798) );
  INVX0 U4930_U2 ( .INP(n2617), .ZN(U4930_n1) );
  AND2X1 U4930_U1 ( .IN1(n2616), .IN2(U4930_n1), .Q(n2594) );
  INVX0 U5128_U2 ( .INP(n4406), .ZN(U5128_n1) );
  AND2X1 U5128_U1 ( .IN1(n3933), .IN2(U5128_n1), .Q(n3940) );
  INVX0 U5141_U2 ( .INP(n4405), .ZN(U5141_n1) );
  AND2X1 U5141_U1 ( .IN1(n3939), .IN2(U5141_n1), .Q(n3936) );
  INVX0 U5749_U2 ( .INP(n1574), .ZN(U5749_n1) );
  AND2X1 U5749_U1 ( .IN1(g2133), .IN2(U5749_n1), .Q(n3159) );
  INVX0 U5750_U2 ( .INP(n1230), .ZN(U5750_n1) );
  AND2X1 U5750_U1 ( .IN1(g1439), .IN2(U5750_n1), .Q(n3163) );
  INVX0 U5751_U2 ( .INP(n885), .ZN(U5751_n1) );
  AND2X1 U5751_U1 ( .IN1(g753), .IN2(U5751_n1), .Q(n3167) );
  INVX0 U5752_U2 ( .INP(n467), .ZN(U5752_n1) );
  AND2X1 U5752_U1 ( .IN1(g65), .IN2(U5752_n1), .Q(n3171) );
  INVX0 U5753_U2 ( .INP(n4522), .ZN(U5753_n1) );
  AND2X1 U5753_U1 ( .IN1(g2142), .IN2(U5753_n1), .Q(n3424) );
  INVX0 U5754_U2 ( .INP(n4526), .ZN(U5754_n1) );
  AND2X1 U5754_U1 ( .IN1(g2151), .IN2(U5754_n1), .Q(n3683) );
  INVX0 U5755_U2 ( .INP(n3888), .ZN(U5755_n1) );
  AND2X1 U5755_U1 ( .IN1(g2160), .IN2(U5755_n1), .Q(n3887) );
  INVX0 U5756_U2 ( .INP(n4523), .ZN(U5756_n1) );
  AND2X1 U5756_U1 ( .IN1(g1448), .IN2(U5756_n1), .Q(n3427) );
  INVX0 U5757_U2 ( .INP(n4527), .ZN(U5757_n1) );
  AND2X1 U5757_U1 ( .IN1(g1457), .IN2(U5757_n1), .Q(n3686) );
  INVX0 U5758_U2 ( .INP(n3891), .ZN(U5758_n1) );
  AND2X1 U5758_U1 ( .IN1(g1466), .IN2(U5758_n1), .Q(n3890) );
  INVX0 U5759_U2 ( .INP(n882), .ZN(U5759_n1) );
  AND2X1 U5759_U1 ( .IN1(g762), .IN2(U5759_n1), .Q(n3430) );
  INVX0 U5760_U2 ( .INP(n879), .ZN(U5760_n1) );
  AND2X1 U5760_U1 ( .IN1(g771), .IN2(U5760_n1), .Q(n3689) );
  INVX0 U5761_U2 ( .INP(n3894), .ZN(U5761_n1) );
  AND2X1 U5761_U1 ( .IN1(g780), .IN2(U5761_n1), .Q(n3893) );
  INVX0 U5762_U2 ( .INP(n4521), .ZN(U5762_n1) );
  AND2X1 U5762_U1 ( .IN1(g74), .IN2(U5762_n1), .Q(n3433) );
  INVX0 U5763_U2 ( .INP(n4528), .ZN(U5763_n1) );
  AND2X1 U5763_U1 ( .IN1(g83), .IN2(U5763_n1), .Q(n3692) );
  INVX0 U5764_U2 ( .INP(n3897), .ZN(U5764_n1) );
  AND2X1 U5764_U1 ( .IN1(g92), .IN2(U5764_n1), .Q(n3896) );
  INVX0 U5882_U2 ( .INP(g3036), .ZN(U5882_n1) );
  AND2X1 U5882_U1 ( .IN1(n4102), .IN2(U5882_n1), .Q(n4101) );
  INVX0 U5939_U2 ( .INP(n1480), .ZN(U5939_n1) );
  AND2X1 U5939_U1 ( .IN1(g2257), .IN2(U5939_n1), .Q(n3038) );
  INVX0 U5940_U2 ( .INP(n1136), .ZN(U5940_n1) );
  AND2X1 U5940_U1 ( .IN1(g1563), .IN2(U5940_n1), .Q(n3070) );
  INVX0 U5941_U2 ( .INP(n791), .ZN(U5941_n1) );
  AND2X1 U5941_U1 ( .IN1(g869), .IN2(U5941_n1), .Q(n3102) );
  INVX0 U5942_U2 ( .INP(n375), .ZN(U5942_n1) );
  AND2X1 U5942_U1 ( .IN1(g181), .IN2(U5942_n1), .Q(n3130) );
  INVX0 U6140_U2 ( .INP(n4066), .ZN(U6140_n1) );
  AND2X1 U6140_U1 ( .IN1(g3002), .IN2(U6140_n1), .Q(n4065) );
  INVX0 U6460_U2 ( .INP(g3230), .ZN(U6460_n1) );
  AND2X1 U6460_U1 ( .IN1(g3233), .IN2(U6460_n1), .Q(n3700) );
  INVX0 U6470_U2 ( .INP(n4305), .ZN(U6470_n1) );
  AND2X1 U6470_U1 ( .IN1(g2892), .IN2(U6470_n1), .Q(n4182) );
  INVX0 U6562_U2 ( .INP(g3204), .ZN(U6562_n1) );
  AND2X1 U6562_U1 ( .IN1(n3938), .IN2(U6562_n1), .Q(n3939) );
  INVX0 U6563_U2 ( .INP(g3204), .ZN(U6563_n1) );
  AND2X1 U6563_U1 ( .IN1(n4073), .IN2(U6563_n1), .Q(n3705) );
  INVX0 U6718_U2 ( .INP(g3197), .ZN(U6718_n1) );
  AND2X1 U6718_U1 ( .IN1(n323), .IN2(U6718_n1), .Q(n4073) );
  INVX0 U7116_U2 ( .INP(g2903), .ZN(U7116_n1) );
  AND2X1 U7116_U1 ( .IN1(n4058), .IN2(U7116_n1), .Q(n4057) );
  INVX0 U7118_U2 ( .INP(g2896), .ZN(U7118_n1) );
  AND2X1 U7118_U1 ( .IN1(n4123), .IN2(U7118_n1), .Q(n4122) );
  INVX0 U7293_U2 ( .INP(g3234), .ZN(U7293_n1) );
  AND2X1 U7293_U1 ( .IN1(n4598), .IN2(U7293_n1), .Q(g20877) );
endmodule

