module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n288_, new_n421_, new_n620_, new_n368_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n240_, new_n526_, new_n442_, new_n642_, new_n211_, new_n552_, new_n342_, new_n462_, new_n603_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n248_, new_n350_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n227_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n598_, new_n570_, new_n143_, new_n520_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n605_, new_n182_, new_n407_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n255_, new_n533_, new_n569_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n412_, new_n327_, new_n594_, new_n561_, new_n495_, new_n196_, new_n574_, new_n319_, new_n640_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n138_, keyIn_0_6 );
xnor g001 ( new_n139_, N73, N77 );
xnor g002 ( new_n140_, new_n139_, new_n138_ );
xnor g003 ( new_n141_, N65, N69 );
xnor g004 ( new_n142_, new_n141_, keyIn_0_5 );
xnor g005 ( new_n143_, new_n140_, new_n142_ );
xnor g006 ( new_n144_, N81, N85 );
xnor g007 ( new_n145_, N89, N93 );
xnor g008 ( new_n146_, new_n144_, new_n145_ );
xnor g009 ( new_n147_, new_n143_, new_n146_ );
nand g010 ( new_n148_, N129, N137 );
not g011 ( new_n149_, new_n148_ );
nand g012 ( new_n150_, new_n147_, new_n149_ );
nand g013 ( new_n151_, new_n143_, new_n146_ );
not g014 ( new_n152_, new_n143_ );
not g015 ( new_n153_, new_n146_ );
nand g016 ( new_n154_, new_n152_, new_n153_ );
nand g017 ( new_n155_, new_n154_, new_n151_, new_n148_ );
nand g018 ( new_n156_, new_n150_, new_n155_ );
xnor g019 ( new_n157_, N1, N17 );
xnor g020 ( new_n158_, N33, N49 );
xnor g021 ( new_n159_, new_n157_, new_n158_ );
not g022 ( new_n160_, new_n159_ );
nand g023 ( new_n161_, new_n156_, new_n160_ );
nand g024 ( new_n162_, new_n150_, new_n155_, new_n159_ );
nand g025 ( new_n163_, new_n161_, new_n162_ );
not g026 ( new_n164_, keyIn_0_23 );
not g027 ( new_n165_, keyIn_0_19 );
xnor g028 ( new_n166_, N121, N125 );
xnor g029 ( new_n167_, new_n166_, keyIn_0_7 );
xor g030 ( new_n168_, N113, N117 );
xnor g031 ( new_n169_, new_n167_, new_n168_ );
xnor g032 ( new_n170_, new_n169_, new_n165_ );
nand g033 ( new_n171_, new_n170_, new_n153_ );
xnor g034 ( new_n172_, new_n169_, keyIn_0_19 );
nand g035 ( new_n173_, new_n172_, new_n146_ );
nand g036 ( new_n174_, new_n171_, new_n173_ );
nand g037 ( new_n175_, N132, N137 );
xnor g038 ( new_n176_, new_n175_, keyIn_0_9 );
not g039 ( new_n177_, new_n176_ );
nand g040 ( new_n178_, new_n174_, new_n177_ );
nand g041 ( new_n179_, new_n171_, new_n173_, new_n176_ );
nand g042 ( new_n180_, new_n178_, new_n179_ );
nand g043 ( new_n181_, new_n180_, new_n164_ );
nand g044 ( new_n182_, new_n178_, keyIn_0_23, new_n179_ );
nand g045 ( new_n183_, new_n181_, new_n182_ );
xnor g046 ( new_n184_, N13, N29 );
xnor g047 ( new_n185_, new_n184_, keyIn_0_14 );
xnor g048 ( new_n186_, N45, N61 );
xnor g049 ( new_n187_, new_n185_, new_n186_ );
not g050 ( new_n188_, new_n187_ );
nand g051 ( new_n189_, new_n183_, new_n188_ );
nand g052 ( new_n190_, new_n181_, new_n182_, new_n187_ );
nand g053 ( new_n191_, new_n189_, new_n190_ );
xnor g054 ( new_n192_, N105, N109 );
xnor g055 ( new_n193_, N97, N101 );
xnor g056 ( new_n194_, new_n192_, new_n193_ );
xnor g057 ( new_n195_, new_n194_, keyIn_0_18 );
nand g058 ( new_n196_, new_n170_, new_n195_ );
not g059 ( new_n197_, new_n195_ );
nand g060 ( new_n198_, new_n172_, new_n197_ );
nand g061 ( new_n199_, new_n196_, new_n198_ );
nand g062 ( new_n200_, new_n199_, keyIn_0_22 );
not g063 ( new_n201_, keyIn_0_22 );
nand g064 ( new_n202_, new_n196_, new_n198_, new_n201_ );
nand g065 ( new_n203_, new_n200_, new_n202_ );
nand g066 ( new_n204_, N130, N137 );
xor g067 ( new_n205_, new_n204_, keyIn_0_8 );
not g068 ( new_n206_, new_n205_ );
nand g069 ( new_n207_, new_n203_, new_n206_ );
nand g070 ( new_n208_, new_n200_, new_n202_, new_n205_ );
nand g071 ( new_n209_, new_n207_, new_n208_ );
xor g072 ( new_n210_, N37, N53 );
xnor g073 ( new_n211_, new_n210_, keyIn_0_13 );
xnor g074 ( new_n212_, N5, N21 );
xnor g075 ( new_n213_, new_n212_, keyIn_0_12 );
xor g076 ( new_n214_, new_n211_, new_n213_ );
not g077 ( new_n215_, new_n214_ );
nand g078 ( new_n216_, new_n209_, new_n215_ );
nand g079 ( new_n217_, new_n207_, new_n208_, new_n214_ );
nand g080 ( new_n218_, new_n216_, new_n217_ );
not g081 ( new_n219_, keyIn_0_26 );
nand g082 ( new_n220_, new_n143_, new_n195_ );
nand g083 ( new_n221_, new_n152_, new_n197_ );
nand g084 ( new_n222_, new_n221_, new_n220_ );
nand g085 ( new_n223_, N131, N137 );
not g086 ( new_n224_, new_n223_ );
nand g087 ( new_n225_, new_n222_, new_n224_ );
nand g088 ( new_n226_, new_n221_, new_n220_, new_n223_ );
nand g089 ( new_n227_, new_n225_, new_n226_ );
xnor g090 ( new_n228_, N9, N25 );
xnor g091 ( new_n229_, N41, N57 );
xor g092 ( new_n230_, new_n228_, new_n229_ );
not g093 ( new_n231_, new_n230_ );
nand g094 ( new_n232_, new_n227_, new_n231_ );
nand g095 ( new_n233_, new_n225_, new_n226_, new_n230_ );
nand g096 ( new_n234_, new_n232_, new_n233_ );
nand g097 ( new_n235_, new_n234_, keyIn_0_24 );
not g098 ( new_n236_, keyIn_0_24 );
nand g099 ( new_n237_, new_n232_, new_n236_, new_n233_ );
nand g100 ( new_n238_, new_n235_, new_n237_ );
nand g101 ( new_n239_, new_n238_, new_n219_ );
nand g102 ( new_n240_, new_n235_, keyIn_0_26, new_n237_ );
nand g103 ( new_n241_, new_n239_, new_n240_ );
nand g104 ( new_n242_, new_n241_, new_n191_, new_n218_, new_n163_ );
nand g105 ( new_n243_, new_n242_, keyIn_0_36 );
not g106 ( new_n244_, keyIn_0_36 );
and g107 ( new_n245_, new_n218_, new_n163_ );
nand g108 ( new_n246_, new_n245_, new_n244_, new_n191_, new_n241_ );
not g109 ( new_n247_, new_n163_ );
nand g110 ( new_n248_, new_n216_, new_n247_, new_n217_, new_n238_ );
not g111 ( new_n249_, keyIn_0_25 );
xnor g112 ( new_n250_, new_n163_, new_n249_ );
nor g113 ( new_n251_, new_n250_, new_n238_ );
nand g114 ( new_n252_, new_n218_, new_n251_ );
nand g115 ( new_n253_, new_n252_, new_n248_ );
nand g116 ( new_n254_, new_n253_, new_n191_ );
not g117 ( new_n255_, new_n191_ );
nand g118 ( new_n256_, new_n255_, new_n247_, new_n218_, new_n238_ );
nand g119 ( new_n257_, new_n246_, new_n254_, new_n243_, new_n256_ );
nand g120 ( new_n258_, N33, N37 );
not g121 ( new_n259_, N33 );
not g122 ( new_n260_, N37 );
nand g123 ( new_n261_, new_n259_, new_n260_ );
nand g124 ( new_n262_, new_n261_, new_n258_ );
nand g125 ( new_n263_, new_n262_, keyIn_0_2 );
not g126 ( new_n264_, keyIn_0_2 );
nand g127 ( new_n265_, new_n261_, new_n264_, new_n258_ );
nand g128 ( new_n266_, new_n263_, new_n265_ );
xnor g129 ( new_n267_, N41, N45 );
nand g130 ( new_n268_, new_n267_, keyIn_0_3 );
not g131 ( new_n269_, keyIn_0_3 );
nand g132 ( new_n270_, N41, N45 );
not g133 ( new_n271_, N41 );
not g134 ( new_n272_, N45 );
nand g135 ( new_n273_, new_n271_, new_n272_ );
nand g136 ( new_n274_, new_n273_, new_n269_, new_n270_ );
nand g137 ( new_n275_, new_n268_, new_n274_ );
nand g138 ( new_n276_, new_n266_, new_n275_ );
nand g139 ( new_n277_, new_n263_, new_n268_, new_n265_, new_n274_ );
nand g140 ( new_n278_, new_n276_, new_n277_ );
nand g141 ( new_n279_, new_n278_, keyIn_0_17 );
not g142 ( new_n280_, keyIn_0_17 );
nand g143 ( new_n281_, new_n276_, new_n280_, new_n277_ );
nand g144 ( new_n282_, new_n279_, new_n281_ );
nand g145 ( new_n283_, N1, N5 );
not g146 ( new_n284_, N1 );
not g147 ( new_n285_, N5 );
nand g148 ( new_n286_, new_n284_, new_n285_ );
nand g149 ( new_n287_, new_n286_, new_n283_ );
xnor g150 ( new_n288_, N9, N13 );
nand g151 ( new_n289_, new_n287_, new_n288_ );
nand g152 ( new_n290_, N9, N13 );
or g153 ( new_n291_, N9, N13 );
nand g154 ( new_n292_, new_n291_, new_n286_, new_n283_, new_n290_ );
nand g155 ( new_n293_, new_n289_, new_n292_ );
nand g156 ( new_n294_, new_n293_, keyIn_0_16 );
not g157 ( new_n295_, keyIn_0_16 );
nand g158 ( new_n296_, new_n289_, new_n295_, new_n292_ );
nand g159 ( new_n297_, new_n294_, new_n296_ );
nand g160 ( new_n298_, new_n282_, new_n297_ );
nand g161 ( new_n299_, new_n279_, new_n281_, new_n294_, new_n296_ );
nand g162 ( new_n300_, new_n298_, new_n299_ );
nand g163 ( new_n301_, new_n300_, keyIn_0_21 );
not g164 ( new_n302_, keyIn_0_21 );
nand g165 ( new_n303_, new_n298_, new_n302_, new_n299_ );
nand g166 ( new_n304_, new_n301_, new_n303_ );
nand g167 ( new_n305_, N135, N137 );
xnor g168 ( new_n306_, new_n305_, keyIn_0_10 );
not g169 ( new_n307_, new_n306_ );
nand g170 ( new_n308_, new_n304_, new_n307_ );
nand g171 ( new_n309_, new_n301_, new_n303_, new_n306_ );
nand g172 ( new_n310_, new_n308_, new_n309_ );
xor g173 ( new_n311_, N73, N89 );
xnor g174 ( new_n312_, N105, N121 );
xnor g175 ( new_n313_, new_n311_, new_n312_ );
xor g176 ( new_n314_, new_n313_, keyIn_0_20 );
not g177 ( new_n315_, new_n314_ );
nand g178 ( new_n316_, new_n310_, new_n315_ );
nand g179 ( new_n317_, new_n308_, new_n309_, new_n314_ );
nand g180 ( new_n318_, new_n316_, new_n317_ );
nand g181 ( new_n319_, N57, N61 );
or g182 ( new_n320_, N57, N61 );
nand g183 ( new_n321_, new_n320_, new_n319_ );
nand g184 ( new_n322_, new_n321_, keyIn_0_4 );
not g185 ( new_n323_, keyIn_0_4 );
nand g186 ( new_n324_, new_n320_, new_n323_, new_n319_ );
nand g187 ( new_n325_, new_n322_, new_n324_ );
xor g188 ( new_n326_, N49, N53 );
not g189 ( new_n327_, new_n326_ );
nand g190 ( new_n328_, new_n325_, new_n327_ );
nand g191 ( new_n329_, new_n322_, new_n324_, new_n326_ );
nand g192 ( new_n330_, new_n328_, new_n329_ );
nand g193 ( new_n331_, new_n282_, new_n330_ );
nand g194 ( new_n332_, new_n279_, new_n281_, new_n328_, new_n329_ );
nand g195 ( new_n333_, new_n331_, new_n332_ );
nand g196 ( new_n334_, N134, N137 );
not g197 ( new_n335_, new_n334_ );
nand g198 ( new_n336_, new_n333_, new_n335_ );
nand g199 ( new_n337_, new_n331_, new_n332_, new_n334_ );
nand g200 ( new_n338_, new_n336_, new_n337_ );
xnor g201 ( new_n339_, N69, N85 );
xnor g202 ( new_n340_, N101, N117 );
xnor g203 ( new_n341_, new_n339_, new_n340_ );
not g204 ( new_n342_, new_n341_ );
nand g205 ( new_n343_, new_n338_, new_n342_ );
nand g206 ( new_n344_, new_n336_, new_n337_, new_n341_ );
and g207 ( new_n345_, new_n343_, new_n344_ );
not g208 ( new_n346_, N21 );
nand g209 ( new_n347_, new_n346_, N17 );
not g210 ( new_n348_, N17 );
nand g211 ( new_n349_, new_n348_, N21 );
nand g212 ( new_n350_, new_n347_, new_n349_ );
nand g213 ( new_n351_, new_n350_, keyIn_0_0 );
not g214 ( new_n352_, keyIn_0_0 );
nand g215 ( new_n353_, new_n347_, new_n349_, new_n352_ );
nand g216 ( new_n354_, new_n351_, new_n353_ );
not g217 ( new_n355_, N29 );
nand g218 ( new_n356_, new_n355_, N25 );
not g219 ( new_n357_, N25 );
nand g220 ( new_n358_, new_n357_, N29 );
nand g221 ( new_n359_, new_n356_, new_n358_ );
nand g222 ( new_n360_, new_n359_, keyIn_0_1 );
not g223 ( new_n361_, keyIn_0_1 );
nand g224 ( new_n362_, new_n356_, new_n358_, new_n361_ );
nand g225 ( new_n363_, new_n360_, new_n362_ );
nand g226 ( new_n364_, new_n354_, new_n363_ );
nand g227 ( new_n365_, new_n351_, new_n360_, new_n353_, new_n362_ );
nand g228 ( new_n366_, new_n364_, new_n365_ );
nand g229 ( new_n367_, new_n366_, new_n297_ );
nand g230 ( new_n368_, new_n364_, new_n294_, new_n296_, new_n365_ );
nand g231 ( new_n369_, new_n367_, new_n368_ );
nand g232 ( new_n370_, new_n369_, N133, N137 );
nand g233 ( new_n371_, N133, N137 );
nand g234 ( new_n372_, new_n367_, new_n368_, new_n371_ );
nand g235 ( new_n373_, new_n370_, new_n372_ );
xnor g236 ( new_n374_, N97, N113 );
xnor g237 ( new_n375_, new_n374_, keyIn_0_15 );
xnor g238 ( new_n376_, N65, N81 );
xnor g239 ( new_n377_, new_n375_, new_n376_ );
not g240 ( new_n378_, new_n377_ );
nand g241 ( new_n379_, new_n373_, new_n378_ );
nand g242 ( new_n380_, new_n370_, new_n372_, new_n377_ );
nand g243 ( new_n381_, new_n379_, new_n380_ );
not g244 ( new_n382_, new_n381_ );
nor g245 ( new_n383_, new_n345_, new_n382_ );
nand g246 ( new_n384_, new_n366_, new_n330_ );
nand g247 ( new_n385_, new_n364_, new_n328_, new_n329_, new_n365_ );
nand g248 ( new_n386_, new_n384_, new_n385_ );
nand g249 ( new_n387_, N136, N137 );
xor g250 ( new_n388_, new_n387_, keyIn_0_11 );
not g251 ( new_n389_, new_n388_ );
nand g252 ( new_n390_, new_n386_, new_n389_ );
nand g253 ( new_n391_, new_n384_, new_n385_, new_n388_ );
nand g254 ( new_n392_, new_n390_, new_n391_ );
xnor g255 ( new_n393_, N77, N93 );
xnor g256 ( new_n394_, N109, N125 );
xnor g257 ( new_n395_, new_n393_, new_n394_ );
not g258 ( new_n396_, new_n395_ );
nand g259 ( new_n397_, new_n392_, new_n396_ );
nand g260 ( new_n398_, new_n390_, new_n391_, new_n395_ );
and g261 ( new_n399_, new_n397_, new_n398_ );
and g262 ( new_n400_, new_n257_, new_n318_, new_n383_, new_n399_ );
nand g263 ( new_n401_, new_n400_, keyIn_0_41, new_n163_ );
not g264 ( new_n402_, keyIn_0_41 );
nand g265 ( new_n403_, new_n400_, new_n163_ );
nand g266 ( new_n404_, new_n403_, new_n402_ );
nand g267 ( new_n405_, new_n404_, new_n401_ );
xnor g268 ( N724, new_n405_, N1 );
not g269 ( new_n407_, new_n218_ );
nand g270 ( new_n408_, new_n400_, keyIn_0_42, new_n407_ );
not g271 ( new_n409_, keyIn_0_42 );
nand g272 ( new_n410_, new_n400_, new_n407_ );
nand g273 ( new_n411_, new_n410_, new_n409_ );
nand g274 ( new_n412_, new_n411_, new_n408_ );
xnor g275 ( N725, new_n412_, new_n285_ );
not g276 ( new_n414_, new_n238_ );
nand g277 ( new_n415_, new_n400_, new_n414_ );
xnor g278 ( N726, new_n415_, N9 );
nand g279 ( new_n417_, new_n400_, new_n255_ );
xnor g280 ( N727, new_n417_, N13 );
not g281 ( new_n419_, new_n318_ );
nand g282 ( new_n420_, new_n397_, new_n398_ );
and g283 ( new_n421_, new_n257_, new_n419_, new_n383_, new_n420_ );
nand g284 ( new_n422_, new_n421_, N17, new_n163_ );
nand g285 ( new_n423_, new_n421_, new_n163_ );
nand g286 ( new_n424_, new_n423_, new_n348_ );
nand g287 ( new_n425_, new_n424_, new_n422_ );
xor g288 ( N728, new_n425_, keyIn_0_54 );
nand g289 ( new_n427_, new_n421_, N21, new_n407_ );
nand g290 ( new_n428_, new_n421_, new_n407_ );
nand g291 ( new_n429_, new_n428_, new_n346_ );
nand g292 ( new_n430_, new_n429_, new_n427_ );
xor g293 ( N729, new_n430_, keyIn_0_55 );
nand g294 ( new_n432_, new_n421_, new_n414_ );
xnor g295 ( N730, new_n432_, N25 );
nand g296 ( new_n434_, new_n421_, keyIn_0_43, new_n255_ );
not g297 ( new_n435_, keyIn_0_43 );
nand g298 ( new_n436_, new_n421_, new_n255_ );
nand g299 ( new_n437_, new_n436_, new_n435_ );
nand g300 ( new_n438_, new_n437_, new_n434_ );
xnor g301 ( N731, new_n438_, N29 );
nand g302 ( new_n440_, new_n345_, new_n382_ );
nor g303 ( new_n441_, new_n440_, new_n420_ );
and g304 ( new_n442_, new_n257_, new_n318_, new_n441_ );
nand g305 ( new_n443_, new_n442_, N33, new_n163_ );
nand g306 ( new_n444_, new_n442_, new_n163_ );
nand g307 ( new_n445_, new_n444_, new_n259_ );
nand g308 ( new_n446_, new_n445_, new_n443_ );
xor g309 ( N732, new_n446_, keyIn_0_56 );
nand g310 ( new_n448_, new_n442_, N37, new_n407_ );
nand g311 ( new_n449_, new_n442_, new_n407_ );
nand g312 ( new_n450_, new_n449_, new_n260_ );
nand g313 ( new_n451_, new_n450_, new_n448_ );
xnor g314 ( N733, new_n451_, keyIn_0_57 );
nand g315 ( new_n453_, new_n442_, keyIn_0_44, new_n414_ );
and g316 ( new_n454_, new_n442_, new_n414_ );
or g317 ( new_n455_, new_n454_, keyIn_0_44 );
nand g318 ( new_n456_, new_n455_, new_n453_ );
nand g319 ( new_n457_, new_n456_, N41 );
nand g320 ( new_n458_, new_n455_, new_n271_, new_n453_ );
nand g321 ( N734, new_n457_, new_n458_ );
nand g322 ( new_n460_, new_n442_, keyIn_0_45, new_n255_ );
not g323 ( new_n461_, keyIn_0_45 );
nand g324 ( new_n462_, new_n257_, new_n255_, new_n318_, new_n441_ );
nand g325 ( new_n463_, new_n462_, new_n461_ );
nand g326 ( new_n464_, new_n460_, new_n463_ );
nand g327 ( new_n465_, new_n464_, N45 );
nand g328 ( new_n466_, new_n460_, new_n272_, new_n463_ );
nand g329 ( new_n467_, new_n465_, new_n466_ );
nand g330 ( new_n468_, new_n467_, keyIn_0_58 );
not g331 ( new_n469_, keyIn_0_58 );
nand g332 ( new_n470_, new_n465_, new_n469_, new_n466_ );
nand g333 ( N735, new_n468_, new_n470_ );
not g334 ( new_n472_, N49 );
nor g335 ( new_n473_, new_n419_, keyIn_0_27 );
and g336 ( new_n474_, new_n419_, keyIn_0_27 );
nor g337 ( new_n475_, new_n474_, new_n473_, new_n440_ );
nand g338 ( new_n476_, new_n257_, keyIn_0_39, new_n420_, new_n475_ );
not g339 ( new_n477_, keyIn_0_39 );
nand g340 ( new_n478_, new_n257_, new_n420_, new_n475_ );
nand g341 ( new_n479_, new_n478_, new_n477_ );
nand g342 ( new_n480_, new_n479_, new_n476_ );
nand g343 ( new_n481_, new_n480_, new_n472_, new_n163_ );
nand g344 ( new_n482_, new_n480_, new_n163_ );
nand g345 ( new_n483_, new_n482_, N49 );
nand g346 ( new_n484_, new_n483_, new_n481_ );
nand g347 ( new_n485_, new_n484_, keyIn_0_59 );
not g348 ( new_n486_, keyIn_0_59 );
nand g349 ( new_n487_, new_n483_, new_n486_, new_n481_ );
nand g350 ( N736, new_n485_, new_n487_ );
not g351 ( new_n489_, keyIn_0_46 );
nand g352 ( new_n490_, new_n480_, new_n489_, new_n407_ );
nand g353 ( new_n491_, new_n480_, new_n407_ );
nand g354 ( new_n492_, new_n491_, keyIn_0_46 );
nand g355 ( new_n493_, new_n492_, new_n490_ );
nand g356 ( new_n494_, new_n493_, N53 );
not g357 ( new_n495_, N53 );
nand g358 ( new_n496_, new_n492_, new_n495_, new_n490_ );
nand g359 ( N737, new_n494_, new_n496_ );
nand g360 ( new_n498_, new_n480_, new_n414_ );
xnor g361 ( N738, new_n498_, N57 );
nand g362 ( new_n500_, new_n480_, new_n255_ );
xnor g363 ( N739, new_n500_, N61 );
not g364 ( new_n502_, keyIn_0_40 );
not g365 ( new_n503_, keyIn_0_31 );
nand g366 ( new_n504_, new_n316_, new_n503_, new_n317_ );
nand g367 ( new_n505_, new_n318_, keyIn_0_31 );
nand g368 ( new_n506_, new_n505_, new_n441_, new_n504_ );
nand g369 ( new_n507_, new_n506_, keyIn_0_37 );
not g370 ( new_n508_, keyIn_0_37 );
nand g371 ( new_n509_, new_n505_, new_n441_, new_n508_, new_n504_ );
not g372 ( new_n510_, keyIn_0_32 );
nand g373 ( new_n511_, new_n316_, new_n510_, new_n317_ );
nand g374 ( new_n512_, new_n318_, keyIn_0_32 );
nand g375 ( new_n513_, new_n343_, new_n344_ );
or g376 ( new_n514_, new_n399_, keyIn_0_33 );
nand g377 ( new_n515_, new_n399_, keyIn_0_33 );
and g378 ( new_n516_, new_n513_, new_n514_, new_n381_, new_n515_ );
nand g379 ( new_n517_, new_n512_, new_n511_, new_n516_ );
not g380 ( new_n518_, keyIn_0_28 );
nand g381 ( new_n519_, new_n343_, new_n518_, new_n344_ );
nand g382 ( new_n520_, new_n513_, keyIn_0_28 );
nor g383 ( new_n521_, new_n399_, new_n381_ );
nand g384 ( new_n522_, new_n520_, new_n519_, new_n521_ );
or g385 ( new_n523_, new_n522_, new_n318_ );
nand g386 ( new_n524_, new_n381_, keyIn_0_29 );
not g387 ( new_n525_, keyIn_0_29 );
nand g388 ( new_n526_, new_n379_, new_n525_, new_n380_ );
nand g389 ( new_n527_, new_n420_, keyIn_0_30 );
not g390 ( new_n528_, keyIn_0_30 );
nand g391 ( new_n529_, new_n397_, new_n528_, new_n398_ );
nand g392 ( new_n530_, new_n524_, new_n527_, new_n526_, new_n529_ );
nor g393 ( new_n531_, new_n530_, new_n345_ );
nand g394 ( new_n532_, new_n531_, new_n318_ );
and g395 ( new_n533_, new_n517_, new_n523_, new_n532_ );
nand g396 ( new_n534_, new_n533_, keyIn_0_38, new_n507_, new_n509_ );
not g397 ( new_n535_, keyIn_0_38 );
nor g398 ( new_n536_, new_n522_, new_n318_ );
and g399 ( new_n537_, new_n531_, new_n318_ );
nor g400 ( new_n538_, new_n537_, new_n536_ );
nand g401 ( new_n539_, new_n507_, new_n509_, new_n538_, new_n517_ );
nand g402 ( new_n540_, new_n539_, new_n535_ );
nand g403 ( new_n541_, new_n540_, new_n534_ );
and g404 ( new_n542_, new_n245_, new_n191_, new_n414_ );
nand g405 ( new_n543_, new_n541_, new_n502_, new_n542_ );
nand g406 ( new_n544_, new_n541_, new_n542_ );
nand g407 ( new_n545_, new_n544_, keyIn_0_40 );
nand g408 ( new_n546_, new_n545_, new_n543_ );
nand g409 ( new_n547_, new_n546_, keyIn_0_47, new_n381_ );
not g410 ( new_n548_, keyIn_0_47 );
nand g411 ( new_n549_, new_n546_, new_n381_ );
nand g412 ( new_n550_, new_n549_, new_n548_ );
nand g413 ( new_n551_, new_n550_, new_n547_ );
nand g414 ( new_n552_, new_n551_, N65 );
not g415 ( new_n553_, N65 );
nand g416 ( new_n554_, new_n550_, new_n553_, new_n547_ );
nand g417 ( N740, new_n552_, new_n554_ );
nand g418 ( new_n556_, new_n546_, keyIn_0_48, new_n345_ );
not g419 ( new_n557_, keyIn_0_48 );
nand g420 ( new_n558_, new_n546_, new_n345_ );
nand g421 ( new_n559_, new_n558_, new_n557_ );
nand g422 ( new_n560_, new_n559_, new_n556_ );
nand g423 ( new_n561_, new_n560_, N69 );
not g424 ( new_n562_, N69 );
nand g425 ( new_n563_, new_n559_, new_n562_, new_n556_ );
nand g426 ( N741, new_n561_, new_n563_ );
nand g427 ( new_n565_, new_n546_, new_n318_ );
xnor g428 ( N742, new_n565_, N73 );
not g429 ( new_n567_, N77 );
nand g430 ( new_n568_, new_n546_, new_n567_, new_n420_ );
nand g431 ( new_n569_, new_n546_, new_n420_ );
nand g432 ( new_n570_, new_n569_, N77 );
nand g433 ( new_n571_, new_n570_, new_n568_ );
nand g434 ( new_n572_, new_n571_, keyIn_0_60 );
not g435 ( new_n573_, keyIn_0_60 );
nand g436 ( new_n574_, new_n570_, new_n573_, new_n568_ );
nand g437 ( N743, new_n572_, new_n574_ );
xnor g438 ( new_n576_, new_n218_, keyIn_0_34 );
nor g439 ( new_n577_, new_n191_, new_n247_, new_n414_ );
nand g440 ( new_n578_, new_n541_, new_n576_, new_n577_ );
not g441 ( new_n579_, new_n578_ );
nand g442 ( new_n580_, new_n579_, new_n381_ );
xnor g443 ( N744, new_n580_, N81 );
nand g444 ( new_n582_, new_n579_, new_n345_ );
or g445 ( new_n583_, new_n582_, keyIn_0_49 );
nand g446 ( new_n584_, new_n582_, keyIn_0_49 );
nand g447 ( new_n585_, new_n583_, new_n584_ );
nand g448 ( new_n586_, new_n585_, N85 );
not g449 ( new_n587_, N85 );
nand g450 ( new_n588_, new_n583_, new_n587_, new_n584_ );
nand g451 ( N745, new_n586_, new_n588_ );
nand g452 ( new_n590_, new_n579_, new_n318_ );
or g453 ( new_n591_, new_n590_, N89 );
nand g454 ( new_n592_, new_n590_, N89 );
nand g455 ( new_n593_, new_n591_, new_n592_ );
nand g456 ( new_n594_, new_n593_, keyIn_0_61 );
not g457 ( new_n595_, keyIn_0_61 );
nand g458 ( new_n596_, new_n591_, new_n595_, new_n592_ );
nand g459 ( N746, new_n594_, new_n596_ );
nand g460 ( new_n598_, new_n579_, new_n420_ );
xnor g461 ( N747, new_n598_, N93 );
xor g462 ( new_n600_, new_n163_, keyIn_0_35 );
nor g463 ( new_n601_, new_n255_, new_n218_, new_n238_, new_n600_ );
and g464 ( new_n602_, new_n541_, new_n601_ );
nand g465 ( new_n603_, new_n602_, new_n381_ );
xnor g466 ( N748, new_n603_, N97 );
nand g467 ( new_n605_, new_n602_, new_n345_ );
xnor g468 ( new_n606_, new_n605_, keyIn_0_50 );
xnor g469 ( N749, new_n606_, N101 );
nand g470 ( new_n608_, new_n602_, new_n318_ );
xnor g471 ( N750, new_n608_, N105 );
nand g472 ( new_n610_, new_n602_, new_n420_ );
xnor g473 ( N751, new_n610_, N109 );
nor g474 ( new_n612_, new_n248_, new_n191_ );
and g475 ( new_n613_, new_n541_, new_n612_ );
nand g476 ( new_n614_, new_n613_, new_n381_ );
xnor g477 ( N752, new_n614_, N113 );
not g478 ( new_n616_, keyIn_0_51 );
nand g479 ( new_n617_, new_n613_, new_n345_ );
xnor g480 ( new_n618_, new_n617_, new_n616_ );
xnor g481 ( N753, new_n618_, N117 );
not g482 ( new_n620_, keyIn_0_62 );
nand g483 ( new_n621_, new_n613_, keyIn_0_52, new_n318_ );
not g484 ( new_n622_, keyIn_0_52 );
nand g485 ( new_n623_, new_n541_, new_n318_, new_n612_ );
nand g486 ( new_n624_, new_n623_, new_n622_ );
nand g487 ( new_n625_, new_n621_, new_n624_ );
nand g488 ( new_n626_, new_n625_, N121 );
not g489 ( new_n627_, N121 );
nand g490 ( new_n628_, new_n621_, new_n627_, new_n624_ );
nand g491 ( new_n629_, new_n626_, new_n628_ );
nand g492 ( new_n630_, new_n629_, new_n620_ );
nand g493 ( new_n631_, new_n626_, keyIn_0_62, new_n628_ );
nand g494 ( N754, new_n630_, new_n631_ );
not g495 ( new_n633_, keyIn_0_63 );
nand g496 ( new_n634_, new_n541_, new_n420_, new_n612_ );
xnor g497 ( new_n635_, new_n634_, keyIn_0_53 );
nand g498 ( new_n636_, new_n635_, N125 );
not g499 ( new_n637_, N125 );
or g500 ( new_n638_, new_n634_, keyIn_0_53 );
nand g501 ( new_n639_, new_n634_, keyIn_0_53 );
nand g502 ( new_n640_, new_n638_, new_n637_, new_n639_ );
nand g503 ( new_n641_, new_n636_, new_n640_ );
nand g504 ( new_n642_, new_n641_, new_n633_ );
nand g505 ( new_n643_, new_n636_, keyIn_0_63, new_n640_ );
nand g506 ( N755, new_n642_, new_n643_ );
endmodule