module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n318_, new_n155_, new_n163_, new_n236_, new_n238_, new_n148_, new_n321_, new_n92_, new_n79_, new_n122_, new_n324_, new_n250_, new_n113_, new_n111_, new_n288_, new_n158_, new_n97_, new_n252_, new_n202_, new_n262_, new_n296_, new_n160_, new_n308_, new_n271_, new_n274_, new_n100_, new_n242_, new_n232_, new_n218_, new_n115_, new_n258_, new_n76_, new_n190_, new_n307_, new_n176_, new_n305_, new_n156_, new_n223_, new_n283_, new_n306_, new_n291_, new_n261_, new_n241_, new_n309_, new_n186_, new_n213_, new_n134_, new_n197_, new_n205_, new_n82_, new_n141_, new_n323_, new_n259_, new_n206_, new_n109_, new_n254_, new_n227_, new_n222_, new_n85_, new_n265_, new_n246_, new_n170_, new_n328_, new_n266_, new_n278_, new_n304_, new_n173_, new_n220_, new_n268_, new_n217_, new_n101_, new_n269_, new_n194_, new_n214_, new_n116_, new_n129_, new_n138_, new_n142_, new_n299_, new_n144_, new_n275_, new_n114_, new_n188_, new_n139_, new_n240_, new_n314_, new_n118_, new_n165_, new_n123_, new_n127_, new_n211_, new_n126_, new_n327_, new_n216_, new_n177_, new_n77_, new_n196_, new_n280_, new_n264_, new_n319_, new_n235_, new_n273_, new_n224_, new_n301_, new_n169_, new_n270_, new_n317_, new_n210_, new_n102_, new_n143_, new_n207_, new_n125_, new_n145_, new_n267_, new_n287_, new_n253_, new_n140_, new_n247_, new_n90_, new_n237_, new_n330_, new_n234_, new_n149_, new_n294_, new_n187_, new_n260_, new_n86_, new_n311_, new_n251_, new_n189_, new_n300_, new_n84_, new_n292_, new_n195_, new_n106_, new_n263_, new_n215_, new_n152_, new_n157_, new_n107_, new_n93_, new_n182_, new_n153_, new_n81_, new_n320_, new_n244_, new_n172_, new_n133_, new_n277_, new_n257_, new_n245_, new_n212_, new_n89_, new_n151_, new_n286_, new_n193_, new_n231_, new_n313_, new_n78_, new_n239_, new_n272_, new_n91_, new_n282_, new_n198_, new_n201_, new_n128_, new_n192_, new_n199_, new_n146_, new_n88_, new_n208_, new_n98_, new_n159_, new_n83_, new_n110_, new_n228_, new_n315_, new_n302_, new_n322_, new_n191_, new_n124_, new_n95_, new_n289_, new_n326_, new_n179_, new_n225_, new_n164_, new_n230_, new_n175_, new_n226_, new_n281_, new_n104_, new_n185_, new_n87_, new_n103_, new_n112_, new_n171_, new_n248_, new_n117_, new_n121_, new_n167_, new_n221_, new_n243_, new_n200_, new_n298_, new_n184_, new_n99_, new_n131_, new_n154_, new_n255_, new_n329_, new_n249_, new_n136_, new_n233_, new_n284_, new_n119_, new_n293_, new_n96_, new_n178_, new_n168_, new_n174_, new_n297_, new_n279_, new_n150_, new_n295_, new_n120_, new_n132_, new_n166_, new_n108_, new_n137_, new_n162_, new_n183_, new_n303_, new_n105_, new_n161_, new_n147_, new_n285_, new_n80_, new_n229_, new_n209_, new_n290_, new_n203_, new_n94_, new_n204_, new_n325_, new_n181_, new_n135_, new_n180_, new_n276_;

not g000 ( new_n76_, keyIn_0_18 );
or g001 ( new_n77_, keyIn_0_8, N102 );
and g002 ( new_n78_, keyIn_0_8, N102 );
not g003 ( new_n79_, new_n78_ );
and g004 ( new_n80_, new_n79_, N108, new_n77_ );
xnor g005 ( new_n81_, new_n80_, keyIn_0_17 );
not g006 ( new_n82_, keyIn_0_16 );
xnor g007 ( new_n83_, keyIn_0_7, N89 );
and g008 ( new_n84_, new_n83_, N95 );
xnor g009 ( new_n85_, new_n84_, new_n82_ );
not g010 ( new_n86_, N24 );
or g011 ( new_n87_, new_n86_, keyIn_0_2 );
not g012 ( new_n88_, keyIn_0_2 );
or g013 ( new_n89_, new_n88_, N24 );
and g014 ( new_n90_, new_n87_, new_n89_, N30 );
xnor g015 ( new_n91_, new_n90_, keyIn_0_11 );
and g016 ( new_n92_, new_n91_, new_n85_, new_n81_ );
not g017 ( new_n93_, keyIn_0_10 );
not g018 ( new_n94_, N17 );
xnor g019 ( new_n95_, keyIn_0_1, N11 );
or g020 ( new_n96_, new_n95_, new_n94_ );
xnor g021 ( new_n97_, new_n96_, new_n93_ );
not g022 ( new_n98_, N63 );
or g023 ( new_n99_, new_n98_, keyIn_0_5 );
not g024 ( new_n100_, keyIn_0_5 );
or g025 ( new_n101_, new_n100_, N63 );
and g026 ( new_n102_, new_n99_, new_n101_, N69 );
xnor g027 ( new_n103_, new_n102_, keyIn_0_14 );
and g028 ( new_n104_, new_n97_, new_n103_ );
xnor g029 ( new_n105_, keyIn_0_4, N50 );
and g030 ( new_n106_, new_n105_, N56 );
xnor g031 ( new_n107_, new_n106_, keyIn_0_13 );
not g032 ( new_n108_, keyIn_0_15 );
or g033 ( new_n109_, keyIn_0_6, N76 );
and g034 ( new_n110_, keyIn_0_6, N76 );
not g035 ( new_n111_, new_n110_ );
and g036 ( new_n112_, new_n111_, N82, new_n109_ );
xnor g037 ( new_n113_, new_n112_, new_n108_ );
and g038 ( new_n114_, new_n107_, new_n113_ );
xor g039 ( new_n115_, keyIn_0_0, N1 );
and g040 ( new_n116_, new_n115_, N4 );
or g041 ( new_n117_, new_n116_, keyIn_0_9 );
not g042 ( new_n118_, keyIn_0_9 );
not g043 ( new_n119_, N4 );
xnor g044 ( new_n120_, keyIn_0_0, N1 );
or g045 ( new_n121_, new_n120_, new_n118_, new_n119_ );
not g046 ( new_n122_, keyIn_0_12 );
xnor g047 ( new_n123_, keyIn_0_3, N37 );
and g048 ( new_n124_, new_n123_, N43 );
or g049 ( new_n125_, new_n124_, new_n122_ );
and g050 ( new_n126_, new_n123_, new_n122_, N43 );
not g051 ( new_n127_, new_n126_ );
and g052 ( new_n128_, new_n117_, new_n121_, new_n125_, new_n127_ );
and g053 ( new_n129_, new_n92_, new_n104_, new_n128_, new_n114_ );
xnor g054 ( N223, new_n129_, new_n76_ );
not g055 ( new_n131_, N56 );
not g056 ( new_n132_, keyIn_0_24 );
xnor g057 ( new_n133_, N223, keyIn_0_19 );
or g058 ( new_n134_, new_n133_, new_n107_ );
not g059 ( new_n135_, new_n107_ );
not g060 ( new_n136_, keyIn_0_19 );
and g061 ( new_n137_, N223, new_n136_ );
xnor g062 ( new_n138_, new_n129_, keyIn_0_18 );
and g063 ( new_n139_, new_n138_, keyIn_0_19 );
or g064 ( new_n140_, new_n137_, new_n139_, new_n135_ );
and g065 ( new_n141_, new_n134_, new_n132_, new_n140_ );
xnor g066 ( new_n142_, new_n133_, new_n107_ );
and g067 ( new_n143_, new_n142_, keyIn_0_24 );
or g068 ( new_n144_, new_n143_, new_n141_, new_n131_, N60 );
not g069 ( new_n145_, N43 );
not g070 ( new_n146_, keyIn_0_23 );
and g071 ( new_n147_, new_n125_, new_n127_ );
or g072 ( new_n148_, new_n133_, new_n147_ );
not g073 ( new_n149_, new_n147_ );
or g074 ( new_n150_, new_n137_, new_n139_, new_n149_ );
and g075 ( new_n151_, new_n148_, new_n146_, new_n150_ );
xnor g076 ( new_n152_, new_n133_, new_n147_ );
and g077 ( new_n153_, new_n152_, keyIn_0_23 );
or g078 ( new_n154_, new_n153_, new_n151_, new_n145_, N47 );
not g079 ( new_n155_, N69 );
or g080 ( new_n156_, new_n133_, new_n103_ );
not g081 ( new_n157_, new_n103_ );
or g082 ( new_n158_, new_n137_, new_n139_, new_n157_ );
and g083 ( new_n159_, new_n156_, keyIn_0_25, new_n158_ );
not g084 ( new_n160_, keyIn_0_25 );
xnor g085 ( new_n161_, new_n133_, new_n103_ );
and g086 ( new_n162_, new_n161_, new_n160_ );
or g087 ( new_n163_, new_n162_, new_n159_, new_n155_, N73 );
and g088 ( new_n164_, new_n144_, new_n154_, new_n163_ );
not g089 ( new_n165_, N108 );
not g090 ( new_n166_, keyIn_0_28 );
not g091 ( new_n167_, new_n81_ );
or g092 ( new_n168_, new_n137_, new_n139_, new_n167_ );
or g093 ( new_n169_, new_n133_, new_n81_ );
and g094 ( new_n170_, new_n169_, new_n166_, new_n168_ );
xnor g095 ( new_n171_, new_n133_, new_n81_ );
and g096 ( new_n172_, new_n171_, keyIn_0_28 );
or g097 ( new_n173_, new_n172_, new_n170_, new_n165_, N112 );
not g098 ( new_n174_, new_n85_ );
xnor g099 ( new_n175_, new_n133_, new_n174_ );
xnor g100 ( new_n176_, new_n175_, keyIn_0_27 );
not g101 ( new_n177_, N95 );
or g102 ( new_n178_, new_n177_, N99 );
or g103 ( new_n179_, new_n176_, new_n178_ );
and g104 ( new_n180_, new_n179_, new_n173_ );
not g105 ( new_n181_, N82 );
not g106 ( new_n182_, new_n113_ );
or g107 ( new_n183_, new_n137_, new_n139_, new_n182_ );
or g108 ( new_n184_, new_n133_, new_n113_ );
and g109 ( new_n185_, new_n184_, keyIn_0_26, new_n183_ );
not g110 ( new_n186_, keyIn_0_26 );
xnor g111 ( new_n187_, new_n133_, new_n113_ );
and g112 ( new_n188_, new_n187_, new_n186_ );
or g113 ( new_n189_, new_n188_, new_n185_, new_n181_, N86 );
not g114 ( new_n190_, N30 );
not g115 ( new_n191_, keyIn_0_22 );
not g116 ( new_n192_, new_n91_ );
or g117 ( new_n193_, new_n137_, new_n139_, new_n192_ );
or g118 ( new_n194_, new_n133_, new_n91_ );
and g119 ( new_n195_, new_n194_, new_n191_, new_n193_ );
xnor g120 ( new_n196_, new_n133_, new_n91_ );
and g121 ( new_n197_, new_n196_, keyIn_0_22 );
or g122 ( new_n198_, new_n197_, new_n195_, new_n190_, N34 );
and g123 ( new_n199_, new_n189_, new_n198_ );
and g124 ( new_n200_, new_n117_, new_n121_ );
not g125 ( new_n201_, new_n200_ );
or g126 ( new_n202_, new_n137_, new_n139_, new_n201_ );
or g127 ( new_n203_, new_n133_, new_n200_ );
and g128 ( new_n204_, new_n203_, keyIn_0_20, new_n202_ );
not g129 ( new_n205_, keyIn_0_20 );
xnor g130 ( new_n206_, new_n133_, new_n200_ );
and g131 ( new_n207_, new_n206_, new_n205_ );
or g132 ( new_n208_, new_n207_, new_n204_, new_n119_, N8 );
not g133 ( new_n209_, keyIn_0_21 );
not g134 ( new_n210_, new_n97_ );
or g135 ( new_n211_, new_n137_, new_n139_, new_n210_ );
or g136 ( new_n212_, new_n133_, new_n97_ );
and g137 ( new_n213_, new_n212_, new_n209_, new_n211_ );
xnor g138 ( new_n214_, new_n133_, new_n97_ );
and g139 ( new_n215_, new_n214_, keyIn_0_21 );
or g140 ( new_n216_, new_n215_, new_n213_, new_n94_, N21 );
and g141 ( new_n217_, new_n208_, new_n216_ );
and g142 ( new_n218_, new_n164_, new_n180_, new_n199_, new_n217_ );
xnor g143 ( N329, new_n218_, keyIn_0_29 );
not g144 ( new_n220_, keyIn_0_30 );
xnor g145 ( new_n221_, N329, new_n208_ );
or g146 ( new_n222_, new_n207_, new_n204_, new_n119_, N14 );
or g147 ( new_n223_, new_n221_, new_n222_ );
xnor g148 ( new_n224_, N329, new_n173_ );
or g149 ( new_n225_, new_n172_, new_n170_, new_n165_, N115 );
or g150 ( new_n226_, new_n224_, new_n225_ );
xnor g151 ( new_n227_, N329, new_n189_ );
or g152 ( new_n228_, new_n188_, new_n185_, new_n181_, N92 );
or g153 ( new_n229_, new_n227_, new_n228_ );
and g154 ( new_n230_, new_n223_, new_n226_, new_n229_ );
or g155 ( new_n231_, new_n162_, new_n155_, new_n159_ );
xnor g156 ( new_n232_, N329, new_n163_ );
or g157 ( new_n233_, new_n232_, N79, new_n231_ );
xnor g158 ( new_n234_, N329, new_n179_ );
or g159 ( new_n235_, new_n176_, new_n177_, N105 );
or g160 ( new_n236_, new_n234_, new_n235_ );
and g161 ( new_n237_, new_n233_, new_n236_ );
xnor g162 ( new_n238_, N329, new_n154_ );
or g163 ( new_n239_, new_n153_, new_n151_, new_n145_, N53 );
or g164 ( new_n240_, new_n238_, new_n239_ );
not g165 ( new_n241_, new_n144_ );
or g166 ( new_n242_, N329, new_n241_ );
or g167 ( new_n243_, new_n144_, keyIn_0_29 );
and g168 ( new_n244_, new_n242_, new_n243_ );
or g169 ( new_n245_, new_n143_, new_n141_, new_n131_, N66 );
or g170 ( new_n246_, new_n244_, new_n245_ );
and g171 ( new_n247_, new_n246_, new_n240_ );
xnor g172 ( new_n248_, N329, new_n198_ );
or g173 ( new_n249_, new_n197_, new_n195_, new_n190_, N40 );
or g174 ( new_n250_, new_n248_, new_n249_ );
xnor g175 ( new_n251_, N329, new_n216_ );
or g176 ( new_n252_, new_n215_, new_n213_, new_n94_, N27 );
or g177 ( new_n253_, new_n251_, new_n252_ );
and g178 ( new_n254_, new_n250_, new_n253_ );
and g179 ( new_n255_, new_n247_, new_n230_, new_n237_, new_n254_ );
xnor g180 ( N370, new_n255_, new_n220_ );
and g181 ( new_n257_, N370, N27 );
and g182 ( new_n258_, N329, N21 );
and g183 ( new_n259_, N223, N11 );
or g184 ( new_n260_, new_n258_, new_n94_, new_n259_ );
or g185 ( new_n261_, new_n257_, new_n260_ );
and g186 ( new_n262_, N370, N40 );
and g187 ( new_n263_, N329, N34 );
and g188 ( new_n264_, N223, N24 );
or g189 ( new_n265_, new_n263_, new_n190_, new_n264_ );
or g190 ( new_n266_, new_n262_, new_n265_ );
and g191 ( new_n267_, new_n261_, new_n266_ );
and g192 ( new_n268_, N370, N66 );
and g193 ( new_n269_, N329, N60 );
and g194 ( new_n270_, N223, N50 );
or g195 ( new_n271_, new_n269_, new_n131_, new_n270_ );
or g196 ( new_n272_, new_n268_, new_n271_ );
and g197 ( new_n273_, N370, N53 );
and g198 ( new_n274_, N329, N47 );
and g199 ( new_n275_, N223, N37 );
or g200 ( new_n276_, new_n274_, new_n145_, new_n275_ );
or g201 ( new_n277_, new_n273_, new_n276_ );
and g202 ( new_n278_, new_n272_, new_n277_ );
and g203 ( new_n279_, N370, N79 );
and g204 ( new_n280_, N329, N73 );
and g205 ( new_n281_, N223, N63 );
or g206 ( new_n282_, new_n280_, new_n155_, new_n281_ );
or g207 ( new_n283_, new_n279_, new_n282_ );
and g208 ( new_n284_, N370, N92 );
and g209 ( new_n285_, N329, N86 );
and g210 ( new_n286_, N223, N76 );
or g211 ( new_n287_, new_n285_, new_n181_, new_n286_ );
or g212 ( new_n288_, new_n284_, new_n287_ );
and g213 ( new_n289_, N370, N115 );
and g214 ( new_n290_, N329, N112 );
and g215 ( new_n291_, N223, N102 );
or g216 ( new_n292_, new_n290_, new_n165_, new_n291_ );
or g217 ( new_n293_, new_n289_, new_n292_ );
and g218 ( new_n294_, N370, N105 );
and g219 ( new_n295_, N329, N99 );
and g220 ( new_n296_, N223, N89 );
or g221 ( new_n297_, new_n295_, new_n177_, new_n296_ );
or g222 ( new_n298_, new_n294_, new_n297_ );
and g223 ( new_n299_, new_n283_, new_n288_, new_n293_, new_n298_ );
and g224 ( new_n300_, new_n299_, keyIn_0_31, new_n267_, new_n278_ );
not g225 ( new_n301_, new_n300_ );
and g226 ( new_n302_, new_n283_, new_n288_ );
and g227 ( new_n303_, new_n293_, new_n298_ );
and g228 ( new_n304_, new_n267_, new_n278_, new_n302_, new_n303_ );
or g229 ( new_n305_, new_n304_, keyIn_0_31 );
and g230 ( new_n306_, N370, N14 );
and g231 ( new_n307_, N329, N8 );
and g232 ( new_n308_, N223, N1 );
or g233 ( new_n309_, new_n306_, new_n119_, new_n307_, new_n308_ );
and g234 ( N421, new_n305_, new_n301_, new_n309_ );
and g235 ( new_n311_, new_n267_, new_n278_ );
not g236 ( N430, new_n311_ );
not g237 ( new_n313_, new_n267_ );
not g238 ( new_n314_, new_n302_ );
and g239 ( new_n315_, new_n314_, new_n278_ );
or g240 ( N431, new_n315_, new_n313_ );
not g241 ( new_n317_, new_n261_ );
not g242 ( new_n318_, new_n277_ );
not g243 ( new_n319_, N79 );
xnor g244 ( new_n320_, new_n255_, keyIn_0_30 );
or g245 ( new_n321_, new_n320_, new_n319_ );
not g246 ( new_n322_, new_n282_ );
and g247 ( new_n323_, new_n272_, new_n321_, new_n322_ );
not g248 ( new_n324_, N105 );
or g249 ( new_n325_, new_n320_, new_n324_ );
not g250 ( new_n326_, new_n297_ );
and g251 ( new_n327_, new_n325_, new_n326_ );
and g252 ( new_n328_, new_n288_, new_n327_ );
or g253 ( new_n329_, new_n323_, new_n328_, new_n318_ );
and g254 ( new_n330_, new_n329_, new_n266_ );
or g255 ( N432, new_n330_, new_n317_ );
endmodule