module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n155_, new_n384_, new_n410_, new_n445_, new_n236_, new_n238_, new_n479_, new_n543_, new_n250_, new_n113_, new_n501_, new_n288_, new_n371_, new_n509_, new_n421_, new_n202_, new_n296_, new_n308_, new_n368_, new_n232_, new_n258_, new_n439_, new_n176_, new_n283_, new_n223_, new_n390_, new_n156_, new_n306_, new_n366_, new_n291_, new_n261_, new_n241_, new_n309_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n323_, new_n401_, new_n389_, new_n259_, new_n362_, new_n514_, new_n227_, new_n416_, new_n222_, new_n456_, new_n170_, new_n246_, new_n571_, new_n400_, new_n328_, new_n266_, new_n367_, new_n173_, new_n220_, new_n130_, new_n505_, new_n419_, new_n471_, new_n268_, new_n374_, new_n577_, new_n534_, new_n376_, new_n380_, new_n214_, new_n451_, new_n489_, new_n424_, new_n138_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n240_, new_n413_, new_n526_, new_n352_, new_n442_, new_n575_, new_n485_, new_n525_, new_n211_, new_n123_, new_n127_, new_n342_, new_n562_, new_n126_, new_n462_, new_n564_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n500_, new_n273_, new_n224_, new_n270_, new_n570_, new_n317_, new_n344_, new_n143_, new_n520_, new_n287_, new_n125_, new_n145_, new_n253_, new_n504_, new_n403_, new_n475_, new_n237_, new_n427_, new_n234_, new_n532_, new_n149_, new_n472_, new_n557_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n106_, new_n411_, new_n215_, new_n152_, new_n157_, new_n107_, new_n182_, new_n407_, new_n153_, new_n480_, new_n133_, new_n257_, new_n212_, new_n151_, new_n513_, new_n364_, new_n449_, new_n580_, new_n484_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n272_, new_n282_, new_n239_, new_n583_, new_n522_, new_n588_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n110_, new_n315_, new_n302_, new_n191_, new_n124_, new_n326_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n387_, new_n544_, new_n476_, new_n589_, new_n112_, new_n248_, new_n350_, new_n117_, new_n121_, new_n415_, new_n167_, new_n537_, new_n221_, new_n385_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n478_, new_n461_, new_n459_, new_n555_, new_n174_, new_n297_, new_n361_, new_n468_, new_n150_, new_n354_, new_n392_, new_n444_, new_n518_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n340_, new_n147_, new_n510_, new_n285_, new_n502_, new_n351_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n517_, new_n325_, new_n417_, new_n180_, new_n530_, new_n332_, new_n318_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n531_, new_n111_, new_n158_, new_n252_, new_n585_, new_n491_, new_n549_, new_n466_, new_n262_, new_n160_, new_n312_, new_n271_, new_n535_, new_n274_, new_n372_, new_n242_, new_n527_, new_n218_, new_n497_, new_n115_, new_n307_, new_n190_, new_n305_, new_n420_, new_n568_, new_n408_, new_n470_, new_n423_, new_n205_, new_n492_, new_n496_, new_n213_, new_n141_, new_n134_, new_n433_, new_n435_, new_n206_, new_n109_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n265_, new_n506_, new_n370_, new_n256_, new_n584_, new_n452_, new_n278_, new_n304_, new_n381_, new_n523_, new_n388_, new_n550_, new_n217_, new_n269_, new_n508_, new_n512_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n129_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n412_, new_n165_, new_n441_, new_n327_, new_n216_, new_n495_, new_n431_, new_n196_, new_n280_, new_n574_, new_n426_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n338_, new_n207_, new_n267_, new_n336_, new_n140_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n587_, new_n465_, new_n195_, new_n567_, new_n263_, new_n334_, new_n331_, new_n576_, new_n341_, new_n378_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n488_, new_n277_, new_n245_, new_n402_, new_n474_, new_n579_, new_n467_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n560_, new_n346_, new_n396_, new_n198_, new_n438_, new_n128_, new_n358_, new_n208_, new_n348_, new_n159_, new_n322_, new_n228_, new_n545_, new_n289_, new_n528_, new_n179_, new_n572_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n185_, new_n399_, new_n373_, new_n171_, new_n559_, new_n540_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n233_, new_n136_, new_n284_, new_n119_, new_n293_, new_n391_, new_n178_, new_n437_, new_n551_, new_n168_, new_n279_, new_n455_, new_n295_, new_n359_, new_n132_, new_n120_, new_n521_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n406_, new_n356_, new_n333_, new_n229_, new_n290_, new_n464_, new_n204_, new_n369_, new_n181_, new_n135_, new_n448_, new_n276_, new_n405_;

not g000 ( new_n106_, keyIn_0_20 );
not g001 ( new_n107_, N85 );
nand g002 ( new_n108_, new_n107_, N81 );
not g003 ( new_n109_, N81 );
nand g004 ( new_n110_, new_n109_, N85 );
nand g005 ( new_n111_, new_n108_, new_n110_ );
xnor g006 ( new_n112_, N89, N93 );
nand g007 ( new_n113_, new_n111_, new_n112_ );
xnor g008 ( new_n114_, N81, N85 );
not g009 ( new_n115_, N93 );
nand g010 ( new_n116_, new_n115_, N89 );
not g011 ( new_n117_, N89 );
nand g012 ( new_n118_, new_n117_, N93 );
nand g013 ( new_n119_, new_n116_, new_n118_ );
nand g014 ( new_n120_, new_n119_, new_n114_ );
nand g015 ( new_n121_, new_n113_, new_n120_ );
nand g016 ( new_n122_, new_n121_, keyIn_0_5 );
not g017 ( new_n123_, keyIn_0_5 );
nand g018 ( new_n124_, new_n113_, new_n120_, new_n123_ );
nand g019 ( new_n125_, new_n122_, new_n124_ );
not g020 ( new_n126_, keyIn_0_4 );
not g021 ( new_n127_, N77 );
nand g022 ( new_n128_, new_n127_, N73 );
not g023 ( new_n129_, N73 );
nand g024 ( new_n130_, new_n129_, N77 );
not g025 ( new_n131_, N65 );
not g026 ( new_n132_, N69 );
nand g027 ( new_n133_, new_n131_, new_n132_ );
nand g028 ( new_n134_, N65, N69 );
nand g029 ( new_n135_, new_n133_, new_n128_, new_n130_, new_n134_ );
nand g030 ( new_n136_, new_n128_, new_n130_ );
xnor g031 ( new_n137_, N65, N69 );
nand g032 ( new_n138_, new_n136_, new_n137_ );
nand g033 ( new_n139_, new_n138_, new_n135_ );
nand g034 ( new_n140_, new_n139_, new_n126_ );
nand g035 ( new_n141_, new_n138_, keyIn_0_4, new_n135_ );
nand g036 ( new_n142_, new_n125_, new_n140_, new_n141_ );
nand g037 ( new_n143_, new_n140_, new_n141_ );
nand g038 ( new_n144_, new_n143_, new_n122_, new_n124_ );
nand g039 ( new_n145_, new_n142_, new_n144_ );
nand g040 ( new_n146_, new_n145_, new_n106_ );
nand g041 ( new_n147_, new_n142_, new_n144_, keyIn_0_20 );
nand g042 ( new_n148_, new_n146_, new_n147_ );
nand g043 ( new_n149_, N129, N137 );
not g044 ( new_n150_, new_n149_ );
nand g045 ( new_n151_, new_n148_, new_n150_ );
nand g046 ( new_n152_, new_n146_, new_n147_, new_n149_ );
nand g047 ( new_n153_, new_n151_, new_n152_ );
nand g048 ( new_n154_, new_n153_, keyIn_0_24 );
not g049 ( new_n155_, keyIn_0_24 );
nand g050 ( new_n156_, new_n151_, new_n155_, new_n152_ );
nand g051 ( new_n157_, new_n154_, new_n156_ );
xor g052 ( new_n158_, N1, N17 );
xnor g053 ( new_n159_, N33, N49 );
xnor g054 ( new_n160_, new_n158_, new_n159_ );
xor g055 ( new_n161_, new_n160_, keyIn_0_8 );
nand g056 ( new_n162_, new_n157_, new_n161_ );
not g057 ( new_n163_, new_n161_ );
nand g058 ( new_n164_, new_n154_, new_n156_, new_n163_ );
nand g059 ( new_n165_, new_n162_, new_n164_ );
not g060 ( new_n166_, keyIn_0_25 );
not g061 ( new_n167_, keyIn_0_21 );
not g062 ( new_n168_, N101 );
nand g063 ( new_n169_, new_n168_, N97 );
not g064 ( new_n170_, N97 );
nand g065 ( new_n171_, new_n170_, N101 );
not g066 ( new_n172_, N109 );
nand g067 ( new_n173_, new_n172_, N105 );
not g068 ( new_n174_, N105 );
nand g069 ( new_n175_, new_n174_, N109 );
nand g070 ( new_n176_, new_n169_, new_n171_, new_n173_, new_n175_ );
nand g071 ( new_n177_, new_n169_, new_n171_ );
nand g072 ( new_n178_, new_n173_, new_n175_ );
nand g073 ( new_n179_, new_n177_, new_n178_ );
nand g074 ( new_n180_, new_n179_, new_n176_, keyIn_0_6 );
not g075 ( new_n181_, keyIn_0_6 );
nand g076 ( new_n182_, new_n179_, new_n176_ );
nand g077 ( new_n183_, new_n182_, new_n181_ );
not g078 ( new_n184_, keyIn_0_7 );
not g079 ( new_n185_, N117 );
nand g080 ( new_n186_, new_n185_, N113 );
not g081 ( new_n187_, N113 );
nand g082 ( new_n188_, new_n187_, N117 );
nand g083 ( new_n189_, new_n186_, new_n188_ );
xnor g084 ( new_n190_, N121, N125 );
nand g085 ( new_n191_, new_n189_, new_n190_ );
xnor g086 ( new_n192_, N113, N117 );
not g087 ( new_n193_, N125 );
nand g088 ( new_n194_, new_n193_, N121 );
not g089 ( new_n195_, N121 );
nand g090 ( new_n196_, new_n195_, N125 );
nand g091 ( new_n197_, new_n194_, new_n196_ );
nand g092 ( new_n198_, new_n197_, new_n192_ );
nand g093 ( new_n199_, new_n191_, new_n198_ );
nand g094 ( new_n200_, new_n199_, new_n184_ );
nand g095 ( new_n201_, new_n191_, new_n198_, keyIn_0_7 );
nand g096 ( new_n202_, new_n200_, new_n183_, new_n180_, new_n201_ );
nand g097 ( new_n203_, new_n183_, new_n180_ );
nand g098 ( new_n204_, new_n200_, new_n201_ );
nand g099 ( new_n205_, new_n204_, new_n203_ );
nand g100 ( new_n206_, new_n205_, new_n167_, new_n202_ );
nand g101 ( new_n207_, new_n205_, new_n202_ );
nand g102 ( new_n208_, new_n207_, keyIn_0_21 );
nand g103 ( new_n209_, new_n208_, new_n206_ );
nand g104 ( new_n210_, N130, N137 );
nand g105 ( new_n211_, new_n209_, new_n210_ );
nand g106 ( new_n212_, new_n208_, N130, N137, new_n206_ );
nand g107 ( new_n213_, new_n211_, new_n212_ );
nand g108 ( new_n214_, new_n213_, new_n166_ );
nand g109 ( new_n215_, new_n211_, keyIn_0_25, new_n212_ );
nand g110 ( new_n216_, new_n214_, new_n215_ );
xor g111 ( new_n217_, N5, N21 );
xnor g112 ( new_n218_, N37, N53 );
xnor g113 ( new_n219_, new_n217_, new_n218_ );
xnor g114 ( new_n220_, new_n219_, keyIn_0_9 );
not g115 ( new_n221_, new_n220_ );
nand g116 ( new_n222_, new_n216_, new_n221_ );
nand g117 ( new_n223_, new_n214_, new_n215_, new_n220_ );
nand g118 ( new_n224_, new_n222_, new_n223_ );
nand g119 ( new_n225_, new_n183_, new_n140_, new_n141_, new_n180_ );
nand g120 ( new_n226_, new_n203_, new_n143_ );
nand g121 ( new_n227_, new_n226_, keyIn_0_22, new_n225_ );
not g122 ( new_n228_, keyIn_0_22 );
nand g123 ( new_n229_, new_n226_, new_n225_ );
nand g124 ( new_n230_, new_n229_, new_n228_ );
nand g125 ( new_n231_, new_n230_, new_n227_ );
nand g126 ( new_n232_, N131, N137 );
not g127 ( new_n233_, new_n232_ );
nand g128 ( new_n234_, new_n231_, new_n233_ );
nand g129 ( new_n235_, new_n230_, new_n227_, new_n232_ );
nand g130 ( new_n236_, new_n234_, new_n235_ );
nand g131 ( new_n237_, new_n236_, keyIn_0_26 );
not g132 ( new_n238_, keyIn_0_26 );
nand g133 ( new_n239_, new_n234_, new_n238_, new_n235_ );
nand g134 ( new_n240_, new_n237_, new_n239_ );
xor g135 ( new_n241_, N9, N25 );
xnor g136 ( new_n242_, N41, N57 );
xnor g137 ( new_n243_, new_n241_, new_n242_ );
xor g138 ( new_n244_, new_n243_, keyIn_0_10 );
xnor g139 ( new_n245_, new_n240_, new_n244_ );
not g140 ( new_n246_, keyIn_0_27 );
nand g141 ( new_n247_, new_n125_, new_n200_, new_n201_ );
nand g142 ( new_n248_, new_n204_, new_n122_, new_n124_ );
nand g143 ( new_n249_, new_n247_, new_n248_ );
nand g144 ( new_n250_, new_n249_, keyIn_0_23 );
not g145 ( new_n251_, keyIn_0_23 );
nand g146 ( new_n252_, new_n247_, new_n248_, new_n251_ );
nand g147 ( new_n253_, new_n250_, N132, N137, new_n252_ );
nand g148 ( new_n254_, new_n250_, new_n252_ );
nand g149 ( new_n255_, N132, N137 );
nand g150 ( new_n256_, new_n254_, new_n255_ );
nand g151 ( new_n257_, new_n256_, new_n253_ );
nand g152 ( new_n258_, new_n257_, new_n246_ );
nand g153 ( new_n259_, new_n256_, keyIn_0_27, new_n253_ );
nand g154 ( new_n260_, new_n258_, new_n259_ );
xor g155 ( new_n261_, N13, N29 );
xnor g156 ( new_n262_, N45, N61 );
xnor g157 ( new_n263_, new_n261_, new_n262_ );
xnor g158 ( new_n264_, new_n263_, keyIn_0_11 );
xnor g159 ( new_n265_, new_n260_, new_n264_ );
nand g160 ( new_n266_, new_n265_, new_n165_, new_n224_, new_n245_ );
not g161 ( new_n267_, new_n266_ );
not g162 ( new_n268_, N53 );
nand g163 ( new_n269_, new_n268_, N49 );
not g164 ( new_n270_, N49 );
nand g165 ( new_n271_, new_n270_, N53 );
not g166 ( new_n272_, N61 );
nand g167 ( new_n273_, new_n272_, N57 );
not g168 ( new_n274_, N57 );
nand g169 ( new_n275_, new_n274_, N61 );
nand g170 ( new_n276_, new_n269_, new_n271_, new_n273_, new_n275_ );
nand g171 ( new_n277_, new_n269_, new_n271_ );
nand g172 ( new_n278_, new_n273_, new_n275_ );
nand g173 ( new_n279_, new_n277_, new_n278_ );
nand g174 ( new_n280_, new_n279_, new_n276_, keyIn_0_3 );
not g175 ( new_n281_, keyIn_0_3 );
nand g176 ( new_n282_, new_n279_, new_n276_ );
nand g177 ( new_n283_, new_n282_, new_n281_ );
nand g178 ( new_n284_, new_n283_, new_n280_ );
not g179 ( new_n285_, N21 );
nand g180 ( new_n286_, new_n285_, N17 );
not g181 ( new_n287_, N17 );
nand g182 ( new_n288_, new_n287_, N21 );
nand g183 ( new_n289_, new_n286_, new_n288_ );
not g184 ( new_n290_, N29 );
nand g185 ( new_n291_, new_n290_, N25 );
not g186 ( new_n292_, N25 );
nand g187 ( new_n293_, new_n292_, N29 );
nand g188 ( new_n294_, new_n289_, new_n291_, new_n293_ );
xnor g189 ( new_n295_, N17, N21 );
nand g190 ( new_n296_, new_n291_, new_n293_ );
nand g191 ( new_n297_, new_n296_, new_n295_ );
nand g192 ( new_n298_, new_n294_, new_n297_, keyIn_0_1 );
not g193 ( new_n299_, keyIn_0_1 );
nand g194 ( new_n300_, new_n294_, new_n297_ );
nand g195 ( new_n301_, new_n300_, new_n299_ );
nand g196 ( new_n302_, new_n284_, new_n298_, new_n301_ );
nand g197 ( new_n303_, new_n301_, new_n298_ );
nand g198 ( new_n304_, new_n303_, new_n280_, new_n283_ );
nand g199 ( new_n305_, new_n304_, new_n302_ );
nand g200 ( new_n306_, new_n305_, keyIn_0_19 );
not g201 ( new_n307_, keyIn_0_19 );
nand g202 ( new_n308_, new_n304_, new_n302_, new_n307_ );
nand g203 ( new_n309_, new_n306_, N136, N137, new_n308_ );
nand g204 ( new_n310_, new_n306_, new_n308_ );
nand g205 ( new_n311_, N136, N137 );
nand g206 ( new_n312_, new_n310_, new_n311_ );
nand g207 ( new_n313_, new_n312_, new_n309_ );
nand g208 ( new_n314_, new_n313_, keyIn_0_31 );
not g209 ( new_n315_, keyIn_0_31 );
nand g210 ( new_n316_, new_n312_, new_n315_, new_n309_ );
xor g211 ( new_n317_, N77, N93 );
xnor g212 ( new_n318_, N109, N125 );
xnor g213 ( new_n319_, new_n317_, new_n318_ );
xor g214 ( new_n320_, new_n319_, keyIn_0_15 );
nand g215 ( new_n321_, new_n314_, new_n316_, new_n320_ );
nand g216 ( new_n322_, new_n314_, new_n316_ );
not g217 ( new_n323_, new_n320_ );
nand g218 ( new_n324_, new_n322_, new_n323_ );
nand g219 ( new_n325_, new_n324_, new_n321_ );
not g220 ( new_n326_, keyIn_0_0 );
not g221 ( new_n327_, N5 );
nand g222 ( new_n328_, new_n327_, N1 );
not g223 ( new_n329_, N1 );
nand g224 ( new_n330_, new_n329_, N5 );
not g225 ( new_n331_, N13 );
nand g226 ( new_n332_, new_n331_, N9 );
not g227 ( new_n333_, N9 );
nand g228 ( new_n334_, new_n333_, N13 );
nand g229 ( new_n335_, new_n328_, new_n330_, new_n332_, new_n334_ );
nand g230 ( new_n336_, new_n328_, new_n330_ );
nand g231 ( new_n337_, new_n332_, new_n334_ );
nand g232 ( new_n338_, new_n336_, new_n337_ );
nand g233 ( new_n339_, new_n338_, new_n335_, new_n326_ );
nand g234 ( new_n340_, new_n338_, new_n335_ );
nand g235 ( new_n341_, new_n340_, keyIn_0_0 );
nand g236 ( new_n342_, new_n341_, new_n339_ );
not g237 ( new_n343_, keyIn_0_2 );
not g238 ( new_n344_, N45 );
nand g239 ( new_n345_, new_n344_, N41 );
not g240 ( new_n346_, N41 );
nand g241 ( new_n347_, new_n346_, N45 );
not g242 ( new_n348_, N33 );
not g243 ( new_n349_, N37 );
nand g244 ( new_n350_, new_n348_, new_n349_ );
nand g245 ( new_n351_, N33, N37 );
nand g246 ( new_n352_, new_n350_, new_n345_, new_n347_, new_n351_ );
nand g247 ( new_n353_, new_n345_, new_n347_ );
xnor g248 ( new_n354_, N33, N37 );
nand g249 ( new_n355_, new_n353_, new_n354_ );
nand g250 ( new_n356_, new_n355_, new_n352_ );
nand g251 ( new_n357_, new_n356_, new_n343_ );
nand g252 ( new_n358_, new_n355_, keyIn_0_2, new_n352_ );
nand g253 ( new_n359_, new_n342_, new_n357_, new_n358_ );
nand g254 ( new_n360_, new_n357_, new_n358_ );
nand g255 ( new_n361_, new_n360_, new_n339_, new_n341_ );
nand g256 ( new_n362_, new_n359_, new_n361_ );
nand g257 ( new_n363_, new_n362_, keyIn_0_18 );
not g258 ( new_n364_, keyIn_0_18 );
nand g259 ( new_n365_, new_n359_, new_n361_, new_n364_ );
nand g260 ( new_n366_, new_n363_, new_n365_ );
nand g261 ( new_n367_, N135, N137 );
not g262 ( new_n368_, new_n367_ );
nand g263 ( new_n369_, new_n366_, new_n368_ );
nand g264 ( new_n370_, new_n363_, new_n365_, new_n367_ );
nand g265 ( new_n371_, new_n369_, new_n370_ );
nand g266 ( new_n372_, new_n371_, keyIn_0_30 );
not g267 ( new_n373_, keyIn_0_30 );
nand g268 ( new_n374_, new_n369_, new_n373_, new_n370_ );
nand g269 ( new_n375_, new_n372_, new_n374_ );
xor g270 ( new_n376_, N73, N89 );
xnor g271 ( new_n377_, N105, N121 );
xnor g272 ( new_n378_, new_n376_, new_n377_ );
xor g273 ( new_n379_, new_n378_, keyIn_0_14 );
not g274 ( new_n380_, new_n379_ );
xnor g275 ( new_n381_, new_n375_, new_n380_ );
nand g276 ( new_n382_, new_n301_, new_n341_, new_n298_, new_n339_ );
nand g277 ( new_n383_, new_n303_, new_n342_ );
nand g278 ( new_n384_, new_n383_, keyIn_0_16, new_n382_ );
not g279 ( new_n385_, keyIn_0_16 );
nand g280 ( new_n386_, new_n383_, new_n382_ );
nand g281 ( new_n387_, new_n386_, new_n385_ );
nand g282 ( new_n388_, new_n387_, new_n384_ );
nand g283 ( new_n389_, N133, N137 );
not g284 ( new_n390_, new_n389_ );
nand g285 ( new_n391_, new_n388_, new_n390_ );
nand g286 ( new_n392_, new_n387_, new_n384_, new_n389_ );
nand g287 ( new_n393_, new_n391_, new_n392_ );
nand g288 ( new_n394_, new_n393_, keyIn_0_28 );
not g289 ( new_n395_, keyIn_0_28 );
nand g290 ( new_n396_, new_n391_, new_n395_, new_n392_ );
nand g291 ( new_n397_, new_n394_, new_n396_ );
xor g292 ( new_n398_, N65, N81 );
xnor g293 ( new_n399_, N97, N113 );
xnor g294 ( new_n400_, new_n398_, new_n399_ );
xnor g295 ( new_n401_, new_n400_, keyIn_0_12 );
not g296 ( new_n402_, new_n401_ );
nand g297 ( new_n403_, new_n397_, new_n402_ );
nand g298 ( new_n404_, new_n394_, new_n396_, new_n401_ );
nand g299 ( new_n405_, new_n403_, new_n404_ );
not g300 ( new_n406_, keyIn_0_17 );
nand g301 ( new_n407_, new_n283_, new_n357_, new_n280_, new_n358_ );
nand g302 ( new_n408_, new_n284_, new_n360_ );
nand g303 ( new_n409_, new_n408_, new_n406_, new_n407_ );
nand g304 ( new_n410_, new_n408_, new_n407_ );
nand g305 ( new_n411_, new_n410_, keyIn_0_17 );
nand g306 ( new_n412_, new_n411_, new_n409_ );
nand g307 ( new_n413_, N134, N137 );
nand g308 ( new_n414_, new_n412_, new_n413_ );
nand g309 ( new_n415_, new_n411_, N134, N137, new_n409_ );
nand g310 ( new_n416_, new_n414_, new_n415_ );
nand g311 ( new_n417_, new_n416_, keyIn_0_29 );
not g312 ( new_n418_, keyIn_0_29 );
nand g313 ( new_n419_, new_n414_, new_n418_, new_n415_ );
nand g314 ( new_n420_, new_n417_, new_n419_ );
xor g315 ( new_n421_, N69, N85 );
xnor g316 ( new_n422_, N101, N117 );
xnor g317 ( new_n423_, new_n421_, new_n422_ );
xnor g318 ( new_n424_, new_n423_, keyIn_0_13 );
not g319 ( new_n425_, new_n424_ );
nand g320 ( new_n426_, new_n420_, new_n425_ );
nand g321 ( new_n427_, new_n417_, new_n419_, new_n424_ );
nand g322 ( new_n428_, new_n426_, new_n427_ );
nand g323 ( new_n429_, new_n405_, new_n428_ );
nor g324 ( new_n430_, new_n429_, new_n381_, new_n325_ );
nand g325 ( new_n431_, new_n267_, new_n430_ );
nand g326 ( new_n432_, new_n431_, N1 );
nand g327 ( new_n433_, new_n267_, new_n329_, new_n430_ );
nand g328 ( N724, new_n432_, new_n433_ );
not g329 ( new_n435_, new_n244_ );
nand g330 ( new_n436_, new_n240_, new_n435_ );
nand g331 ( new_n437_, new_n237_, new_n239_, new_n244_ );
nand g332 ( new_n438_, new_n436_, new_n437_ );
not g333 ( new_n439_, new_n264_ );
nand g334 ( new_n440_, new_n260_, new_n439_ );
nand g335 ( new_n441_, new_n258_, new_n259_, new_n264_ );
nand g336 ( new_n442_, new_n440_, new_n441_ );
nor g337 ( new_n443_, new_n165_, new_n442_, new_n224_, new_n438_ );
nand g338 ( new_n444_, new_n443_, new_n430_ );
nand g339 ( new_n445_, new_n444_, N5 );
nand g340 ( new_n446_, new_n443_, new_n327_, new_n430_ );
nand g341 ( N725, new_n445_, new_n446_ );
xnor g342 ( new_n448_, new_n157_, new_n163_ );
nand g343 ( new_n449_, new_n265_, new_n448_, new_n224_, new_n438_ );
not g344 ( new_n450_, new_n449_ );
nand g345 ( new_n451_, new_n450_, new_n430_ );
nand g346 ( new_n452_, new_n451_, N9 );
nand g347 ( new_n453_, new_n450_, new_n333_, new_n430_ );
nand g348 ( N726, new_n452_, new_n453_ );
nand g349 ( new_n455_, new_n448_, new_n245_, new_n224_, new_n442_ );
not g350 ( new_n456_, new_n455_ );
nand g351 ( new_n457_, new_n456_, new_n430_ );
nand g352 ( new_n458_, new_n457_, N13 );
nand g353 ( new_n459_, new_n456_, new_n430_, new_n331_ );
nand g354 ( N727, new_n458_, new_n459_ );
xnor g355 ( new_n461_, new_n322_, new_n320_ );
nand g356 ( new_n462_, new_n375_, new_n379_ );
nand g357 ( new_n463_, new_n372_, new_n374_, new_n380_ );
nand g358 ( new_n464_, new_n462_, new_n463_ );
nor g359 ( new_n465_, new_n429_, new_n461_, new_n464_ );
nand g360 ( new_n466_, new_n267_, new_n465_ );
nand g361 ( new_n467_, new_n466_, N17 );
nand g362 ( new_n468_, new_n267_, new_n465_, new_n287_ );
nand g363 ( N728, new_n467_, new_n468_ );
nand g364 ( new_n470_, new_n443_, new_n465_ );
nand g365 ( new_n471_, new_n470_, N21 );
nand g366 ( new_n472_, new_n443_, new_n465_, new_n285_ );
nand g367 ( N729, new_n471_, new_n472_ );
nand g368 ( new_n474_, new_n450_, new_n465_ );
nand g369 ( new_n475_, new_n474_, N25 );
nand g370 ( new_n476_, new_n450_, new_n292_, new_n465_ );
nand g371 ( N730, new_n475_, new_n476_ );
nand g372 ( new_n478_, new_n456_, new_n465_ );
nand g373 ( new_n479_, new_n478_, N29 );
nand g374 ( new_n480_, new_n456_, new_n465_, new_n290_ );
nand g375 ( N731, new_n479_, new_n480_ );
nor g376 ( new_n482_, new_n381_, new_n325_, new_n405_, new_n428_ );
nand g377 ( new_n483_, new_n267_, new_n482_ );
nand g378 ( new_n484_, new_n483_, N33 );
nand g379 ( new_n485_, new_n267_, new_n482_, new_n348_ );
nand g380 ( N732, new_n484_, new_n485_ );
nand g381 ( new_n487_, new_n443_, new_n482_ );
nand g382 ( new_n488_, new_n487_, N37 );
nand g383 ( new_n489_, new_n443_, new_n482_, new_n349_ );
nand g384 ( N733, new_n488_, new_n489_ );
nand g385 ( new_n491_, new_n450_, new_n482_ );
nand g386 ( new_n492_, new_n491_, N41 );
nand g387 ( new_n493_, new_n450_, new_n482_, new_n346_ );
nand g388 ( N734, new_n492_, new_n493_ );
nand g389 ( new_n495_, new_n482_, new_n456_ );
nand g390 ( new_n496_, new_n495_, N45 );
nand g391 ( new_n497_, new_n482_, new_n456_, new_n344_ );
nand g392 ( N735, new_n496_, new_n497_ );
nor g393 ( new_n499_, new_n461_, new_n464_, new_n405_, new_n428_ );
nand g394 ( new_n500_, new_n267_, new_n499_ );
nand g395 ( new_n501_, new_n500_, N49 );
nand g396 ( new_n502_, new_n267_, new_n499_, new_n270_ );
nand g397 ( N736, new_n501_, new_n502_ );
nand g398 ( new_n504_, new_n443_, new_n499_ );
nand g399 ( new_n505_, new_n504_, N53 );
nand g400 ( new_n506_, new_n443_, new_n499_, new_n268_ );
nand g401 ( N737, new_n505_, new_n506_ );
nand g402 ( new_n508_, new_n450_, new_n499_ );
nand g403 ( new_n509_, new_n508_, N57 );
nand g404 ( new_n510_, new_n450_, new_n499_, new_n274_ );
nand g405 ( N738, new_n509_, new_n510_ );
nand g406 ( new_n512_, new_n499_, new_n456_ );
nand g407 ( new_n513_, new_n512_, N61 );
nand g408 ( new_n514_, new_n499_, new_n456_, new_n272_ );
nand g409 ( N739, new_n513_, new_n514_ );
nand g410 ( new_n516_, new_n461_, new_n381_, new_n405_, new_n428_ );
not g411 ( new_n517_, new_n516_ );
nand g412 ( new_n518_, new_n165_, new_n224_ );
nand g413 ( new_n519_, new_n438_, new_n440_, new_n441_ );
nor g414 ( new_n520_, new_n518_, new_n519_ );
nand g415 ( new_n521_, new_n517_, new_n520_ );
nand g416 ( new_n522_, new_n521_, N65 );
nand g417 ( new_n523_, new_n517_, new_n131_, new_n520_ );
nand g418 ( N740, new_n522_, new_n523_ );
nor g419 ( new_n525_, new_n325_, new_n464_, new_n405_, new_n428_ );
nand g420 ( new_n526_, new_n525_, new_n520_ );
nand g421 ( new_n527_, new_n526_, N69 );
nand g422 ( new_n528_, new_n525_, new_n520_, new_n132_ );
nand g423 ( N741, new_n527_, new_n528_ );
xnor g424 ( new_n530_, new_n397_, new_n401_ );
nand g425 ( new_n531_, new_n461_, new_n530_, new_n464_, new_n428_ );
not g426 ( new_n532_, new_n531_ );
nand g427 ( new_n533_, new_n532_, new_n520_ );
nand g428 ( new_n534_, new_n533_, N73 );
nand g429 ( new_n535_, new_n532_, new_n129_, new_n520_ );
nand g430 ( N742, new_n534_, new_n535_ );
nand g431 ( new_n537_, new_n381_, new_n530_, new_n325_, new_n428_ );
not g432 ( new_n538_, new_n537_ );
nand g433 ( new_n539_, new_n538_, new_n520_ );
nand g434 ( new_n540_, new_n539_, N77 );
nand g435 ( new_n541_, new_n538_, new_n520_, new_n127_ );
nand g436 ( N743, new_n540_, new_n541_ );
nand g437 ( new_n543_, new_n245_, new_n442_, new_n165_, new_n224_ );
not g438 ( new_n544_, new_n543_ );
nand g439 ( new_n545_, new_n517_, new_n544_ );
nand g440 ( new_n546_, new_n545_, N81 );
nand g441 ( new_n547_, new_n517_, new_n109_, new_n544_ );
nand g442 ( N744, new_n546_, new_n547_ );
nand g443 ( new_n549_, new_n525_, new_n544_ );
nand g444 ( new_n550_, new_n549_, N85 );
nand g445 ( new_n551_, new_n525_, new_n107_, new_n544_ );
nand g446 ( N745, new_n550_, new_n551_ );
nor g447 ( new_n553_, new_n531_, new_n543_ );
xnor g448 ( N746, new_n553_, new_n117_ );
nor g449 ( new_n555_, new_n537_, new_n543_ );
xnor g450 ( N747, new_n555_, new_n115_ );
nor g451 ( new_n557_, new_n519_, new_n165_, new_n224_ );
nand g452 ( new_n558_, new_n517_, new_n557_ );
nand g453 ( new_n559_, new_n558_, N97 );
nand g454 ( new_n560_, new_n517_, new_n170_, new_n557_ );
nand g455 ( N748, new_n559_, new_n560_ );
nand g456 ( new_n562_, new_n525_, new_n557_ );
nand g457 ( new_n563_, new_n562_, N101 );
nand g458 ( new_n564_, new_n525_, new_n557_, new_n168_ );
nand g459 ( N749, new_n563_, new_n564_ );
nand g460 ( new_n566_, new_n532_, new_n557_ );
nand g461 ( new_n567_, new_n566_, N105 );
nand g462 ( new_n568_, new_n532_, new_n174_, new_n557_ );
nand g463 ( N750, new_n567_, new_n568_ );
nand g464 ( new_n570_, new_n538_, new_n557_ );
nand g465 ( new_n571_, new_n570_, N109 );
nand g466 ( new_n572_, new_n538_, new_n557_, new_n172_ );
nand g467 ( N751, new_n571_, new_n572_ );
nor g468 ( new_n574_, new_n265_, new_n165_, new_n224_, new_n438_ );
nand g469 ( new_n575_, new_n517_, new_n574_ );
nand g470 ( new_n576_, new_n575_, N113 );
nand g471 ( new_n577_, new_n517_, new_n574_, new_n187_ );
nand g472 ( N752, new_n576_, new_n577_ );
nand g473 ( new_n579_, new_n525_, new_n574_ );
nand g474 ( new_n580_, new_n579_, N117 );
nand g475 ( new_n581_, new_n525_, new_n574_, new_n185_ );
nand g476 ( N753, new_n580_, new_n581_ );
nand g477 ( new_n583_, new_n532_, new_n574_ );
nand g478 ( new_n584_, new_n583_, N121 );
nand g479 ( new_n585_, new_n532_, new_n574_, new_n195_ );
nand g480 ( N754, new_n584_, new_n585_ );
nand g481 ( new_n587_, new_n574_, new_n538_ );
nand g482 ( new_n588_, new_n587_, N125 );
nand g483 ( new_n589_, new_n574_, new_n538_, new_n193_ );
nand g484 ( N755, new_n588_, new_n589_ );
endmodule