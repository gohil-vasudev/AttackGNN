module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n170_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n257_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n326_, new_n554_, new_n648_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n297_, new_n361_, new_n565_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n578_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n407_, new_n666_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n662_, new_n531_, new_n593_, new_n252_, new_n585_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n269_, new_n512_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n697_, new_n373_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n151_, N75 );
nand g001 ( new_n152_, N29, N42 );
nor g002 ( N388, new_n152_, new_n151_ );
not g003 ( new_n154_, N29 );
not g004 ( new_n155_, N36 );
nor g005 ( new_n156_, new_n154_, new_n155_ );
and g006 ( N389, new_n156_, N80 );
nand g007 ( new_n158_, new_n156_, N42 );
not g008 ( N390, new_n158_ );
and g009 ( N391, N85, N86 );
not g010 ( new_n161_, N13 );
nand g011 ( new_n162_, N1, N8 );
nor g012 ( new_n163_, new_n162_, new_n161_ );
and g013 ( N418, new_n163_, N17 );
nand g014 ( new_n165_, N1, N26 );
nand g015 ( new_n166_, N13, N17 );
nor g016 ( new_n167_, new_n165_, new_n166_ );
nand g017 ( N419, new_n158_, new_n167_ );
not g018 ( new_n169_, N59 );
nor g019 ( new_n170_, new_n169_, new_n151_ );
nand g020 ( N420, new_n170_, N80 );
nor g021 ( new_n172_, new_n155_, new_n169_ );
nand g022 ( N421, new_n172_, N80 );
nand g023 ( N422, new_n172_, N42 );
not g024 ( new_n175_, N90 );
nor g025 ( new_n176_, N87, N88 );
nor g026 ( N423, new_n176_, new_n175_ );
nand g027 ( N446, N390, new_n167_ );
not g028 ( new_n179_, keyIn_0_0 );
not g029 ( new_n180_, N51 );
nor g030 ( new_n181_, new_n165_, new_n180_ );
xnor g031 ( N447, new_n181_, new_n179_ );
nand g032 ( new_n183_, new_n163_, N55 );
nand g033 ( new_n184_, N29, N68 );
nor g034 ( N448, new_n183_, new_n184_ );
and g035 ( new_n186_, N59, N68 );
nand g036 ( new_n187_, new_n186_, N74 );
nor g037 ( N449, new_n183_, new_n187_ );
not g038 ( new_n189_, N89 );
nor g039 ( N450, new_n176_, new_n189_ );
not g040 ( new_n191_, N135 );
xnor g041 ( new_n192_, N111, N116 );
xnor g042 ( new_n193_, N121, N126 );
xnor g043 ( new_n194_, new_n192_, new_n193_ );
nand g044 ( new_n195_, new_n194_, new_n191_ );
xor g045 ( new_n196_, new_n195_, keyIn_0_21 );
nor g046 ( new_n197_, new_n194_, new_n191_ );
nor g047 ( new_n198_, new_n196_, new_n197_ );
xnor g048 ( new_n199_, N91, N96 );
xnor g049 ( new_n200_, N101, N106 );
xor g050 ( new_n201_, new_n199_, new_n200_ );
xnor g051 ( new_n202_, new_n201_, N130 );
xnor g052 ( N767, new_n198_, new_n202_ );
nand g053 ( new_n204_, N183, N189 );
xnor g054 ( new_n205_, new_n204_, keyIn_0_6 );
not g055 ( new_n206_, N183 );
not g056 ( new_n207_, N189 );
nand g057 ( new_n208_, new_n206_, new_n207_ );
nand g058 ( new_n209_, new_n205_, new_n208_ );
xnor g059 ( new_n210_, N195, N201 );
xnor g060 ( new_n211_, new_n209_, new_n210_ );
xnor g061 ( new_n212_, new_n211_, N207 );
xor g062 ( new_n213_, N159, N165 );
xnor g063 ( new_n214_, N171, N177 );
xnor g064 ( new_n215_, new_n213_, new_n214_ );
xnor g065 ( new_n216_, new_n215_, N130 );
xnor g066 ( N768, new_n212_, new_n216_ );
not g067 ( new_n218_, N261 );
not g068 ( new_n219_, N201 );
not g069 ( new_n220_, keyIn_0_15 );
nand g070 ( new_n221_, new_n181_, keyIn_0_0 );
and g071 ( new_n222_, N1, N26 );
nand g072 ( new_n223_, new_n222_, N51 );
nand g073 ( new_n224_, new_n223_, new_n179_ );
nand g074 ( new_n225_, new_n224_, new_n221_ );
nand g075 ( new_n226_, new_n225_, keyIn_0_8 );
not g076 ( new_n227_, keyIn_0_8 );
nand g077 ( new_n228_, N447, new_n227_ );
nand g078 ( new_n229_, new_n228_, new_n226_ );
xnor g079 ( new_n230_, new_n229_, keyIn_0_12 );
nor g080 ( new_n231_, N17, N42 );
xor g081 ( new_n232_, new_n231_, keyIn_0_4 );
nand g082 ( new_n233_, N17, N42 );
xnor g083 ( new_n234_, new_n233_, keyIn_0_5 );
nand g084 ( new_n235_, new_n232_, new_n234_ );
nor g085 ( new_n236_, new_n235_, keyIn_0_11 );
not g086 ( new_n237_, new_n236_ );
nand g087 ( new_n238_, new_n235_, keyIn_0_11 );
nand g088 ( new_n239_, N59, N156 );
not g089 ( new_n240_, new_n239_ );
and g090 ( new_n241_, new_n238_, new_n240_ );
nand g091 ( new_n242_, new_n241_, new_n237_ );
nor g092 ( new_n243_, new_n230_, new_n242_ );
nand g093 ( new_n244_, new_n243_, new_n220_ );
xnor g094 ( new_n245_, new_n225_, new_n227_ );
nand g095 ( new_n246_, new_n245_, keyIn_0_12 );
not g096 ( new_n247_, keyIn_0_12 );
nand g097 ( new_n248_, new_n229_, new_n247_ );
nand g098 ( new_n249_, new_n246_, new_n248_ );
nand g099 ( new_n250_, new_n238_, new_n240_ );
nor g100 ( new_n251_, new_n250_, new_n236_ );
nand g101 ( new_n252_, new_n249_, new_n251_ );
nand g102 ( new_n253_, new_n252_, keyIn_0_15 );
nand g103 ( new_n254_, new_n244_, new_n253_ );
nand g104 ( new_n255_, N42, N59 );
nor g105 ( new_n256_, new_n255_, new_n151_ );
xor g106 ( new_n257_, new_n256_, keyIn_0_2 );
xnor g107 ( new_n258_, new_n257_, keyIn_0_10 );
nand g108 ( new_n259_, N17, N51 );
nor g109 ( new_n260_, new_n162_, new_n259_ );
xor g110 ( new_n261_, new_n260_, keyIn_0_1 );
xnor g111 ( new_n262_, new_n261_, keyIn_0_9 );
nand g112 ( new_n263_, new_n262_, new_n258_ );
xor g113 ( new_n264_, new_n263_, keyIn_0_13 );
nand g114 ( new_n265_, new_n254_, new_n264_ );
nand g115 ( new_n266_, new_n265_, keyIn_0_17 );
not g116 ( new_n267_, keyIn_0_17 );
xnor g117 ( new_n268_, new_n252_, new_n220_ );
xnor g118 ( new_n269_, new_n263_, keyIn_0_13 );
nor g119 ( new_n270_, new_n268_, new_n269_ );
nand g120 ( new_n271_, new_n270_, new_n267_ );
nand g121 ( new_n272_, new_n271_, new_n266_ );
nand g122 ( new_n273_, new_n272_, N126 );
not g123 ( new_n274_, keyIn_0_18 );
not g124 ( new_n275_, keyIn_0_16 );
not g125 ( new_n276_, N17 );
xnor g126 ( new_n277_, new_n239_, keyIn_0_3 );
nor g127 ( new_n278_, new_n277_, new_n276_ );
nand g128 ( new_n279_, new_n249_, new_n278_ );
nor g129 ( new_n280_, new_n279_, new_n275_ );
nand g130 ( new_n281_, new_n279_, new_n275_ );
nand g131 ( new_n282_, new_n281_, N1 );
nor g132 ( new_n283_, new_n282_, new_n280_ );
xnor g133 ( new_n284_, new_n283_, new_n274_ );
nand g134 ( new_n285_, new_n284_, N153 );
nand g135 ( new_n286_, new_n273_, new_n285_ );
xnor g136 ( new_n287_, new_n286_, keyIn_0_27 );
nor g137 ( new_n288_, new_n154_, new_n151_ );
nand g138 ( new_n289_, new_n288_, N80 );
nor g139 ( new_n290_, new_n230_, new_n289_ );
nand g140 ( new_n291_, new_n290_, N55 );
xnor g141 ( new_n292_, new_n291_, keyIn_0_14 );
nor g142 ( new_n293_, new_n292_, N268 );
not g143 ( new_n294_, new_n293_ );
nand g144 ( new_n295_, new_n287_, new_n294_ );
xor g145 ( new_n296_, new_n295_, keyIn_0_30 );
nand g146 ( new_n297_, new_n296_, new_n219_ );
xnor g147 ( new_n298_, new_n297_, keyIn_0_35 );
nor g148 ( new_n299_, new_n296_, new_n219_ );
not g149 ( new_n300_, new_n299_ );
nand g150 ( new_n301_, new_n298_, new_n300_ );
nand g151 ( new_n302_, new_n301_, new_n218_ );
not g152 ( new_n303_, N219 );
nor g153 ( new_n304_, new_n301_, new_n218_ );
nor g154 ( new_n305_, new_n304_, new_n303_ );
nand g155 ( new_n306_, new_n305_, new_n302_ );
not g156 ( new_n307_, N228 );
nor g157 ( new_n308_, new_n301_, new_n307_ );
nand g158 ( new_n309_, new_n299_, N237 );
not g159 ( new_n310_, N246 );
nor g160 ( new_n311_, new_n296_, new_n310_ );
and g161 ( new_n312_, N42, N72 );
and g162 ( new_n313_, new_n312_, N73 );
nand g163 ( new_n314_, new_n313_, new_n186_ );
nor g164 ( new_n315_, new_n314_, new_n183_ );
nand g165 ( new_n316_, new_n315_, N201 );
nand g166 ( new_n317_, N121, N210 );
xnor g167 ( new_n318_, new_n317_, keyIn_0_7 );
nand g168 ( new_n319_, N255, N267 );
and g169 ( new_n320_, new_n318_, new_n319_ );
nand g170 ( new_n321_, new_n316_, new_n320_ );
nor g171 ( new_n322_, new_n311_, new_n321_ );
nand g172 ( new_n323_, new_n322_, new_n309_ );
nor g173 ( new_n324_, new_n308_, new_n323_ );
nand g174 ( N850, new_n306_, new_n324_ );
not g175 ( new_n326_, keyIn_0_42 );
not g176 ( new_n327_, keyIn_0_40 );
not g177 ( new_n328_, keyIn_0_28 );
not g178 ( new_n329_, keyIn_0_22 );
nand g179 ( new_n330_, new_n284_, N146 );
xnor g180 ( new_n331_, new_n330_, new_n329_ );
not g181 ( new_n332_, keyIn_0_23 );
nand g182 ( new_n333_, new_n272_, N116 );
nand g183 ( new_n334_, new_n333_, new_n332_ );
not g184 ( new_n335_, N116 );
xnor g185 ( new_n336_, new_n265_, new_n267_ );
nor g186 ( new_n337_, new_n336_, new_n335_ );
nand g187 ( new_n338_, new_n337_, keyIn_0_23 );
nand g188 ( new_n339_, new_n338_, new_n334_ );
nor g189 ( new_n340_, new_n331_, new_n339_ );
nand g190 ( new_n341_, new_n340_, keyIn_0_25 );
not g191 ( new_n342_, keyIn_0_25 );
xnor g192 ( new_n343_, new_n330_, keyIn_0_22 );
xnor g193 ( new_n344_, new_n333_, keyIn_0_23 );
nand g194 ( new_n345_, new_n343_, new_n344_ );
nand g195 ( new_n346_, new_n345_, new_n342_ );
nand g196 ( new_n347_, new_n341_, new_n346_ );
xnor g197 ( new_n348_, new_n293_, keyIn_0_20 );
nand g198 ( new_n349_, new_n347_, new_n348_ );
xnor g199 ( new_n350_, new_n349_, new_n328_ );
nor g200 ( new_n351_, new_n350_, N189 );
nand g201 ( new_n352_, new_n351_, keyIn_0_32 );
not g202 ( new_n353_, keyIn_0_32 );
xnor g203 ( new_n354_, new_n349_, keyIn_0_28 );
nand g204 ( new_n355_, new_n354_, new_n207_ );
nand g205 ( new_n356_, new_n355_, new_n353_ );
nand g206 ( new_n357_, new_n352_, new_n356_ );
not g207 ( new_n358_, new_n357_ );
not g208 ( new_n359_, N195 );
not g209 ( new_n360_, keyIn_0_24 );
nand g210 ( new_n361_, new_n272_, N121 );
nor g211 ( new_n362_, new_n361_, new_n360_ );
nand g212 ( new_n363_, new_n361_, new_n360_ );
nand g213 ( new_n364_, new_n284_, N149 );
nand g214 ( new_n365_, new_n363_, new_n364_ );
or g215 ( new_n366_, new_n365_, new_n362_ );
nor g216 ( new_n367_, new_n366_, keyIn_0_26 );
nand g217 ( new_n368_, new_n366_, keyIn_0_26 );
nand g218 ( new_n369_, new_n368_, new_n294_ );
nor g219 ( new_n370_, new_n369_, new_n367_ );
nand g220 ( new_n371_, new_n370_, keyIn_0_29 );
not g221 ( new_n372_, keyIn_0_29 );
not g222 ( new_n373_, new_n367_ );
not g223 ( new_n374_, keyIn_0_26 );
nor g224 ( new_n375_, new_n365_, new_n362_ );
nor g225 ( new_n376_, new_n375_, new_n374_ );
nor g226 ( new_n377_, new_n376_, new_n293_ );
nand g227 ( new_n378_, new_n373_, new_n377_ );
nand g228 ( new_n379_, new_n378_, new_n372_ );
nand g229 ( new_n380_, new_n371_, new_n379_ );
nor g230 ( new_n381_, new_n380_, new_n359_ );
xnor g231 ( new_n382_, new_n381_, keyIn_0_33 );
xnor g232 ( new_n383_, new_n382_, keyIn_0_37 );
nor g233 ( new_n384_, new_n383_, new_n358_ );
xnor g234 ( new_n385_, new_n384_, new_n327_ );
not g235 ( new_n386_, keyIn_0_34 );
nand g236 ( new_n387_, new_n380_, new_n359_ );
xnor g237 ( new_n388_, new_n387_, new_n386_ );
nand g238 ( new_n389_, new_n357_, new_n388_ );
nor g239 ( new_n390_, new_n389_, new_n300_ );
xnor g240 ( new_n391_, new_n390_, keyIn_0_41 );
not g241 ( new_n392_, keyIn_0_36 );
nand g242 ( new_n393_, new_n350_, N189 );
nand g243 ( new_n394_, new_n393_, keyIn_0_31 );
not g244 ( new_n395_, keyIn_0_31 );
nor g245 ( new_n396_, new_n354_, new_n207_ );
nand g246 ( new_n397_, new_n396_, new_n395_ );
nand g247 ( new_n398_, new_n397_, new_n394_ );
nand g248 ( new_n399_, new_n398_, new_n392_ );
xnor g249 ( new_n400_, new_n393_, new_n395_ );
nand g250 ( new_n401_, new_n400_, keyIn_0_36 );
nand g251 ( new_n402_, new_n401_, new_n399_ );
nand g252 ( new_n403_, new_n402_, keyIn_0_39 );
not g253 ( new_n404_, keyIn_0_39 );
xnor g254 ( new_n405_, new_n398_, keyIn_0_36 );
nand g255 ( new_n406_, new_n405_, new_n404_ );
nand g256 ( new_n407_, new_n406_, new_n403_ );
nand g257 ( new_n408_, new_n298_, N261 );
nor g258 ( new_n409_, new_n389_, new_n408_ );
xnor g259 ( new_n410_, new_n409_, keyIn_0_38 );
nand g260 ( new_n411_, new_n410_, new_n407_ );
nor g261 ( new_n412_, new_n411_, new_n391_ );
nand g262 ( new_n413_, new_n412_, new_n385_ );
xnor g263 ( new_n414_, new_n413_, new_n326_ );
nand g264 ( new_n415_, new_n284_, N143 );
xor g265 ( new_n416_, new_n293_, keyIn_0_19 );
not g266 ( new_n417_, N111 );
nor g267 ( new_n418_, new_n336_, new_n417_ );
nor g268 ( new_n419_, new_n416_, new_n418_ );
and g269 ( new_n420_, new_n419_, new_n415_ );
nand g270 ( new_n421_, new_n420_, new_n206_ );
not g271 ( new_n422_, new_n421_ );
nor g272 ( new_n423_, new_n414_, new_n422_ );
nor g273 ( new_n424_, new_n420_, new_n206_ );
not g274 ( new_n425_, new_n424_ );
nand g275 ( new_n426_, new_n423_, new_n425_ );
nand g276 ( new_n427_, new_n425_, new_n421_ );
nand g277 ( new_n428_, new_n414_, new_n427_ );
and g278 ( new_n429_, new_n428_, N219 );
nand g279 ( new_n430_, new_n429_, new_n426_ );
nor g280 ( new_n431_, new_n427_, new_n307_ );
nand g281 ( new_n432_, new_n424_, N237 );
nor g282 ( new_n433_, new_n420_, new_n310_ );
nand g283 ( new_n434_, new_n315_, N183 );
nand g284 ( new_n435_, N106, N210 );
nand g285 ( new_n436_, new_n434_, new_n435_ );
nor g286 ( new_n437_, new_n433_, new_n436_ );
nand g287 ( new_n438_, new_n437_, new_n432_ );
nor g288 ( new_n439_, new_n431_, new_n438_ );
nand g289 ( N863, new_n430_, new_n439_ );
not g290 ( new_n441_, new_n408_ );
nor g291 ( new_n442_, new_n441_, new_n299_ );
not g292 ( new_n443_, new_n442_ );
nand g293 ( new_n444_, new_n443_, new_n388_ );
nand g294 ( new_n445_, new_n444_, new_n383_ );
nor g295 ( new_n446_, new_n358_, new_n398_ );
nor g296 ( new_n447_, new_n445_, new_n446_ );
nand g297 ( new_n448_, new_n445_, new_n446_ );
nand g298 ( new_n449_, new_n448_, N219 );
nor g299 ( new_n450_, new_n449_, new_n447_ );
and g300 ( new_n451_, N111, N210 );
nor g301 ( new_n452_, new_n450_, new_n451_ );
xnor g302 ( new_n453_, new_n452_, keyIn_0_50 );
not g303 ( new_n454_, N237 );
nor g304 ( new_n455_, new_n402_, new_n454_ );
nand g305 ( new_n456_, new_n446_, N228 );
nor g306 ( new_n457_, new_n354_, new_n310_ );
nand g307 ( new_n458_, new_n315_, N189 );
nand g308 ( new_n459_, N255, N259 );
nand g309 ( new_n460_, new_n458_, new_n459_ );
nor g310 ( new_n461_, new_n457_, new_n460_ );
nand g311 ( new_n462_, new_n456_, new_n461_ );
nor g312 ( new_n463_, new_n462_, new_n455_ );
nand g313 ( N864, new_n453_, new_n463_ );
nand g314 ( new_n465_, new_n382_, new_n388_ );
nand g315 ( new_n466_, new_n442_, new_n465_ );
nor g316 ( new_n467_, new_n442_, new_n465_ );
nor g317 ( new_n468_, new_n467_, new_n303_ );
nand g318 ( new_n469_, new_n468_, new_n466_ );
nor g319 ( new_n470_, new_n383_, new_n454_ );
or g320 ( new_n471_, new_n465_, new_n307_ );
nor g321 ( new_n472_, new_n380_, new_n310_ );
nand g322 ( new_n473_, new_n315_, N195 );
nand g323 ( new_n474_, N116, N210 );
nand g324 ( new_n475_, N255, N260 );
and g325 ( new_n476_, new_n474_, new_n475_ );
nand g326 ( new_n477_, new_n473_, new_n476_ );
nor g327 ( new_n478_, new_n472_, new_n477_ );
nand g328 ( new_n479_, new_n471_, new_n478_ );
nor g329 ( new_n480_, new_n470_, new_n479_ );
nand g330 ( N865, new_n480_, new_n469_ );
not g331 ( new_n482_, keyIn_0_48 );
not g332 ( new_n483_, keyIn_0_43 );
nand g333 ( new_n484_, new_n423_, new_n483_ );
xnor g334 ( new_n485_, new_n384_, keyIn_0_40 );
not g335 ( new_n486_, new_n391_ );
xnor g336 ( new_n487_, new_n402_, new_n404_ );
not g337 ( new_n488_, keyIn_0_38 );
nand g338 ( new_n489_, new_n409_, new_n488_ );
and g339 ( new_n490_, new_n357_, new_n388_ );
nand g340 ( new_n491_, new_n490_, new_n441_ );
nand g341 ( new_n492_, new_n491_, keyIn_0_38 );
nand g342 ( new_n493_, new_n492_, new_n489_ );
nor g343 ( new_n494_, new_n487_, new_n493_ );
nand g344 ( new_n495_, new_n494_, new_n486_ );
nor g345 ( new_n496_, new_n495_, new_n485_ );
nand g346 ( new_n497_, new_n496_, new_n326_ );
nand g347 ( new_n498_, new_n413_, keyIn_0_42 );
nand g348 ( new_n499_, new_n497_, new_n498_ );
nand g349 ( new_n500_, new_n499_, new_n421_ );
nand g350 ( new_n501_, new_n500_, keyIn_0_43 );
nand g351 ( new_n502_, new_n484_, new_n501_ );
nand g352 ( new_n503_, new_n502_, new_n425_ );
xnor g353 ( new_n504_, new_n503_, keyIn_0_44 );
nand g354 ( new_n505_, new_n272_, N96 );
not g355 ( new_n506_, N146 );
not g356 ( new_n507_, N55 );
nor g357 ( new_n508_, new_n277_, new_n507_ );
nand g358 ( new_n509_, new_n249_, new_n508_ );
nor g359 ( new_n510_, new_n509_, new_n506_ );
nor g360 ( new_n511_, new_n276_, N268 );
nand g361 ( new_n512_, new_n290_, new_n511_ );
nand g362 ( new_n513_, N51, N138 );
nand g363 ( new_n514_, new_n512_, new_n513_ );
nor g364 ( new_n515_, new_n514_, new_n510_ );
nand g365 ( new_n516_, new_n505_, new_n515_ );
nor g366 ( new_n517_, new_n516_, N165 );
nand g367 ( new_n518_, new_n272_, N101 );
not g368 ( new_n519_, N149 );
nor g369 ( new_n520_, new_n509_, new_n519_ );
nand g370 ( new_n521_, N17, N138 );
nand g371 ( new_n522_, new_n512_, new_n521_ );
nor g372 ( new_n523_, new_n522_, new_n520_ );
nand g373 ( new_n524_, new_n518_, new_n523_ );
nor g374 ( new_n525_, new_n524_, N171 );
nor g375 ( new_n526_, new_n517_, new_n525_ );
not g376 ( new_n527_, new_n526_ );
nand g377 ( new_n528_, new_n272_, N106 );
not g378 ( new_n529_, N153 );
nor g379 ( new_n530_, new_n509_, new_n529_ );
nand g380 ( new_n531_, N138, N152 );
nand g381 ( new_n532_, new_n512_, new_n531_ );
nor g382 ( new_n533_, new_n532_, new_n530_ );
nand g383 ( new_n534_, new_n528_, new_n533_ );
nor g384 ( new_n535_, new_n534_, N177 );
nor g385 ( new_n536_, new_n527_, new_n535_ );
nand g386 ( new_n537_, new_n504_, new_n536_ );
nor g387 ( new_n538_, new_n537_, keyIn_0_47 );
nand g388 ( new_n539_, new_n537_, keyIn_0_47 );
nand g389 ( new_n540_, new_n534_, N177 );
nor g390 ( new_n541_, new_n527_, new_n540_ );
nand g391 ( new_n542_, new_n524_, N171 );
nor g392 ( new_n543_, new_n517_, new_n542_ );
nand g393 ( new_n544_, new_n516_, N165 );
not g394 ( new_n545_, new_n544_ );
nor g395 ( new_n546_, new_n543_, new_n545_ );
not g396 ( new_n547_, new_n546_ );
nor g397 ( new_n548_, new_n541_, new_n547_ );
nand g398 ( new_n549_, new_n539_, new_n548_ );
nor g399 ( new_n550_, new_n549_, new_n538_ );
xnor g400 ( new_n551_, new_n550_, new_n482_ );
nand g401 ( new_n552_, new_n272_, N91 );
not g402 ( new_n553_, N143 );
nor g403 ( new_n554_, new_n509_, new_n553_ );
nand g404 ( new_n555_, N8, N138 );
nand g405 ( new_n556_, new_n512_, new_n555_ );
nor g406 ( new_n557_, new_n556_, new_n554_ );
nand g407 ( new_n558_, new_n552_, new_n557_ );
nor g408 ( new_n559_, new_n558_, N159 );
or g409 ( new_n560_, new_n551_, new_n559_ );
nand g410 ( new_n561_, new_n558_, N159 );
nand g411 ( N866, new_n560_, new_n561_ );
not g412 ( new_n563_, keyIn_0_49 );
not g413 ( new_n564_, keyIn_0_44 );
nand g414 ( new_n565_, new_n503_, new_n564_ );
xnor g415 ( new_n566_, new_n500_, new_n483_ );
nor g416 ( new_n567_, new_n566_, new_n424_ );
nand g417 ( new_n568_, new_n567_, keyIn_0_44 );
nand g418 ( new_n569_, new_n568_, new_n565_ );
not g419 ( new_n570_, new_n535_ );
nand g420 ( new_n571_, new_n570_, new_n540_ );
nor g421 ( new_n572_, new_n569_, new_n571_ );
xnor g422 ( new_n573_, new_n572_, keyIn_0_46 );
nand g423 ( new_n574_, new_n569_, new_n571_ );
xor g424 ( new_n575_, new_n574_, keyIn_0_45 );
nand g425 ( new_n576_, new_n575_, new_n573_ );
nor g426 ( new_n577_, new_n576_, new_n563_ );
nand g427 ( new_n578_, new_n576_, new_n563_ );
nand g428 ( new_n579_, new_n578_, N219 );
nor g429 ( new_n580_, new_n579_, new_n577_ );
xor g430 ( new_n581_, new_n580_, keyIn_0_53 );
nand g431 ( new_n582_, N101, N210 );
nand g432 ( new_n583_, new_n581_, new_n582_ );
xnor g433 ( new_n584_, new_n583_, keyIn_0_55 );
nor g434 ( new_n585_, new_n571_, new_n307_ );
nor g435 ( new_n586_, new_n540_, new_n454_ );
nand g436 ( new_n587_, new_n534_, N246 );
nand g437 ( new_n588_, new_n315_, N177 );
nand g438 ( new_n589_, new_n587_, new_n588_ );
or g439 ( new_n590_, new_n586_, new_n589_ );
nor g440 ( new_n591_, new_n585_, new_n590_ );
nand g441 ( new_n592_, new_n584_, new_n591_ );
xnor g442 ( new_n593_, new_n592_, keyIn_0_57 );
xnor g443 ( new_n594_, new_n593_, keyIn_0_59 );
xnor g444 ( N874, new_n594_, keyIn_0_61 );
not g445 ( new_n596_, keyIn_0_62 );
not g446 ( new_n597_, keyIn_0_56 );
not g447 ( new_n598_, new_n538_ );
not g448 ( new_n599_, keyIn_0_47 );
not g449 ( new_n600_, new_n536_ );
nor g450 ( new_n601_, new_n569_, new_n600_ );
nor g451 ( new_n602_, new_n601_, new_n599_ );
not g452 ( new_n603_, new_n548_ );
nor g453 ( new_n604_, new_n602_, new_n603_ );
nand g454 ( new_n605_, new_n604_, new_n598_ );
nand g455 ( new_n606_, new_n605_, new_n482_ );
nand g456 ( new_n607_, new_n550_, keyIn_0_48 );
nand g457 ( new_n608_, new_n606_, new_n607_ );
not g458 ( new_n609_, new_n561_ );
nor g459 ( new_n610_, new_n609_, new_n559_ );
nand g460 ( new_n611_, new_n608_, new_n610_ );
nand g461 ( new_n612_, new_n611_, keyIn_0_52 );
not g462 ( new_n613_, keyIn_0_52 );
and g463 ( new_n614_, new_n608_, new_n610_ );
nand g464 ( new_n615_, new_n614_, new_n613_ );
nand g465 ( new_n616_, new_n615_, new_n612_ );
not g466 ( new_n617_, new_n610_ );
nand g467 ( new_n618_, new_n551_, new_n617_ );
nand g468 ( new_n619_, new_n618_, keyIn_0_51 );
not g469 ( new_n620_, keyIn_0_51 );
nor g470 ( new_n621_, new_n608_, new_n610_ );
nand g471 ( new_n622_, new_n621_, new_n620_ );
nand g472 ( new_n623_, new_n619_, new_n622_ );
nor g473 ( new_n624_, new_n616_, new_n623_ );
nand g474 ( new_n625_, new_n624_, keyIn_0_54 );
not g475 ( new_n626_, keyIn_0_54 );
xnor g476 ( new_n627_, new_n611_, new_n613_ );
and g477 ( new_n628_, new_n619_, new_n622_ );
nand g478 ( new_n629_, new_n628_, new_n627_ );
nand g479 ( new_n630_, new_n629_, new_n626_ );
nand g480 ( new_n631_, new_n630_, new_n625_ );
and g481 ( new_n632_, new_n631_, N219 );
nand g482 ( new_n633_, new_n632_, new_n597_ );
nand g483 ( new_n634_, new_n631_, N219 );
nand g484 ( new_n635_, new_n634_, keyIn_0_56 );
nand g485 ( new_n636_, new_n633_, new_n635_ );
nand g486 ( new_n637_, N210, N268 );
nand g487 ( new_n638_, new_n636_, new_n637_ );
nor g488 ( new_n639_, new_n638_, keyIn_0_58 );
not g489 ( new_n640_, new_n639_ );
nand g490 ( new_n641_, new_n638_, keyIn_0_58 );
nor g491 ( new_n642_, new_n617_, new_n307_ );
nand g492 ( new_n643_, new_n609_, N237 );
nand g493 ( new_n644_, new_n558_, N246 );
nand g494 ( new_n645_, new_n315_, N159 );
and g495 ( new_n646_, new_n644_, new_n645_ );
nand g496 ( new_n647_, new_n643_, new_n646_ );
nor g497 ( new_n648_, new_n642_, new_n647_ );
and g498 ( new_n649_, new_n641_, new_n648_ );
nand g499 ( new_n650_, new_n649_, new_n640_ );
nand g500 ( new_n651_, new_n650_, keyIn_0_60 );
not g501 ( new_n652_, keyIn_0_60 );
nand g502 ( new_n653_, new_n641_, new_n648_ );
nor g503 ( new_n654_, new_n653_, new_n639_ );
nand g504 ( new_n655_, new_n654_, new_n652_ );
nand g505 ( new_n656_, new_n651_, new_n655_ );
nand g506 ( new_n657_, new_n656_, new_n596_ );
xnor g507 ( new_n658_, new_n654_, keyIn_0_60 );
nand g508 ( new_n659_, new_n658_, keyIn_0_62 );
nand g509 ( new_n660_, new_n659_, new_n657_ );
nand g510 ( new_n661_, new_n660_, keyIn_0_63 );
not g511 ( new_n662_, keyIn_0_63 );
xnor g512 ( new_n663_, new_n656_, keyIn_0_62 );
nand g513 ( new_n664_, new_n663_, new_n662_ );
nand g514 ( N878, new_n664_, new_n661_ );
not g515 ( new_n666_, new_n525_ );
nand g516 ( new_n667_, new_n504_, new_n570_ );
nand g517 ( new_n668_, new_n667_, new_n540_ );
nand g518 ( new_n669_, new_n668_, new_n666_ );
nand g519 ( new_n670_, new_n669_, new_n542_ );
nor g520 ( new_n671_, new_n545_, new_n517_ );
nand g521 ( new_n672_, new_n670_, new_n671_ );
nor g522 ( new_n673_, new_n670_, new_n671_ );
nor g523 ( new_n674_, new_n673_, new_n303_ );
nand g524 ( new_n675_, new_n674_, new_n672_ );
and g525 ( new_n676_, new_n671_, N228 );
nand g526 ( new_n677_, new_n545_, N237 );
and g527 ( new_n678_, new_n516_, N246 );
nand g528 ( new_n679_, new_n315_, N165 );
nand g529 ( new_n680_, N91, N210 );
nand g530 ( new_n681_, new_n679_, new_n680_ );
nor g531 ( new_n682_, new_n678_, new_n681_ );
nand g532 ( new_n683_, new_n682_, new_n677_ );
nor g533 ( new_n684_, new_n676_, new_n683_ );
nand g534 ( N879, new_n675_, new_n684_ );
not g535 ( new_n686_, new_n542_ );
nor g536 ( new_n687_, new_n686_, new_n525_ );
nand g537 ( new_n688_, new_n668_, new_n687_ );
nor g538 ( new_n689_, new_n668_, new_n687_ );
nor g539 ( new_n690_, new_n689_, new_n303_ );
nand g540 ( new_n691_, new_n690_, new_n688_ );
and g541 ( new_n692_, new_n687_, N228 );
nand g542 ( new_n693_, new_n686_, N237 );
and g543 ( new_n694_, new_n524_, N246 );
nand g544 ( new_n695_, new_n315_, N171 );
nand g545 ( new_n696_, N96, N210 );
nand g546 ( new_n697_, new_n695_, new_n696_ );
nor g547 ( new_n698_, new_n694_, new_n697_ );
nand g548 ( new_n699_, new_n698_, new_n693_ );
nor g549 ( new_n700_, new_n692_, new_n699_ );
nand g550 ( N880, new_n691_, new_n700_ );
endmodule