module add_mul_combine_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_mul_0_, 
        Result_mul_1_, Result_mul_2_, Result_mul_3_, Result_mul_4_, 
        Result_mul_5_, Result_mul_6_, Result_mul_7_, Result_mul_8_, 
        Result_mul_9_, Result_mul_10_, Result_mul_11_, Result_mul_12_, 
        Result_mul_13_, Result_mul_14_, Result_mul_15_, Result_add_0_, 
        Result_add_1_, Result_add_2_, Result_add_3_, Result_add_4_, 
        Result_add_5_, Result_add_6_, Result_add_7_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_;
  wire   n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858;

  XNOR2_X1 U445 ( .A(n421), .B(n422), .ZN(Result_mul_9_) );
  XOR2_X1 U446 ( .A(n423), .B(n424), .Z(n422) );
  XNOR2_X1 U447 ( .A(n425), .B(n426), .ZN(Result_mul_8_) );
  XOR2_X1 U448 ( .A(n427), .B(n428), .Z(n426) );
  XOR2_X1 U449 ( .A(n429), .B(n430), .Z(Result_mul_7_) );
  AND2_X1 U450 ( .A1(n431), .A2(n432), .ZN(Result_mul_6_) );
  OR2_X1 U451 ( .A1(n433), .A2(n434), .ZN(n431) );
  XOR2_X1 U452 ( .A(n435), .B(n436), .Z(n434) );
  INV_X1 U453 ( .A(n437), .ZN(n433) );
  OR2_X1 U454 ( .A1(n429), .A2(n430), .ZN(n437) );
  XNOR2_X1 U455 ( .A(n438), .B(n439), .ZN(Result_mul_5_) );
  OR2_X1 U456 ( .A1(n440), .A2(n441), .ZN(n438) );
  XOR2_X1 U457 ( .A(n442), .B(n443), .Z(Result_mul_4_) );
  XOR2_X1 U458 ( .A(n444), .B(n445), .Z(Result_mul_3_) );
  AND2_X1 U459 ( .A1(n446), .A2(n447), .ZN(n445) );
  OR2_X1 U460 ( .A1(n448), .A2(n449), .ZN(n447) );
  AND2_X1 U461 ( .A1(n450), .A2(n451), .ZN(n449) );
  INV_X1 U462 ( .A(n452), .ZN(n446) );
  XOR2_X1 U463 ( .A(n453), .B(n454), .Z(Result_mul_2_) );
  XOR2_X1 U464 ( .A(n455), .B(n456), .Z(Result_mul_1_) );
  AND2_X1 U465 ( .A1(n457), .A2(n458), .ZN(n456) );
  OR2_X1 U466 ( .A1(n459), .A2(n460), .ZN(n458) );
  AND2_X1 U467 ( .A1(n461), .A2(n462), .ZN(n459) );
  INV_X1 U468 ( .A(n463), .ZN(n457) );
  XNOR2_X1 U469 ( .A(n464), .B(n465), .ZN(Result_mul_14_) );
  AND2_X1 U470 ( .A1(b_7_), .A2(a_6_), .ZN(n465) );
  XNOR2_X1 U471 ( .A(n466), .B(n467), .ZN(Result_mul_13_) );
  XOR2_X1 U472 ( .A(n468), .B(n469), .Z(n467) );
  XNOR2_X1 U473 ( .A(n470), .B(n471), .ZN(Result_mul_12_) );
  XOR2_X1 U474 ( .A(n472), .B(n473), .Z(n471) );
  XNOR2_X1 U475 ( .A(n474), .B(n475), .ZN(Result_mul_11_) );
  XOR2_X1 U476 ( .A(n476), .B(n477), .Z(n475) );
  XNOR2_X1 U477 ( .A(n478), .B(n479), .ZN(Result_mul_10_) );
  XOR2_X1 U478 ( .A(n480), .B(n481), .Z(n479) );
  OR3_X1 U479 ( .A1(n463), .A2(n482), .A3(n483), .ZN(Result_mul_0_) );
  AND2_X1 U480 ( .A1(n484), .A2(a_0_), .ZN(n483) );
  AND2_X1 U481 ( .A1(n455), .A2(n460), .ZN(n482) );
  AND2_X1 U482 ( .A1(n453), .A2(n454), .ZN(n455) );
  XOR2_X1 U483 ( .A(n462), .B(n461), .Z(n454) );
  OR2_X1 U484 ( .A1(n485), .A2(n486), .ZN(n453) );
  INV_X1 U485 ( .A(n487), .ZN(n486) );
  OR2_X1 U486 ( .A1(n488), .A2(n452), .ZN(n485) );
  AND3_X1 U487 ( .A1(n451), .A2(n450), .A3(n448), .ZN(n452) );
  AND2_X1 U488 ( .A1(n444), .A2(n448), .ZN(n488) );
  AND2_X1 U489 ( .A1(n489), .A2(n487), .ZN(n448) );
  OR2_X1 U490 ( .A1(n490), .A2(n491), .ZN(n487) );
  INV_X1 U491 ( .A(n492), .ZN(n489) );
  AND2_X1 U492 ( .A1(n490), .A2(n491), .ZN(n492) );
  OR2_X1 U493 ( .A1(n493), .A2(n494), .ZN(n491) );
  AND2_X1 U494 ( .A1(n495), .A2(n496), .ZN(n494) );
  AND2_X1 U495 ( .A1(n497), .A2(n498), .ZN(n493) );
  OR2_X1 U496 ( .A1(n496), .A2(n495), .ZN(n498) );
  XOR2_X1 U497 ( .A(n499), .B(n500), .Z(n490) );
  XOR2_X1 U498 ( .A(n501), .B(n502), .Z(n500) );
  AND2_X1 U499 ( .A1(n442), .A2(n443), .ZN(n444) );
  XOR2_X1 U500 ( .A(n451), .B(n450), .Z(n443) );
  INV_X1 U501 ( .A(n503), .ZN(n450) );
  OR2_X1 U502 ( .A1(n504), .A2(n505), .ZN(n503) );
  AND2_X1 U503 ( .A1(n506), .A2(n507), .ZN(n505) );
  AND2_X1 U504 ( .A1(n508), .A2(n509), .ZN(n504) );
  OR2_X1 U505 ( .A1(n507), .A2(n506), .ZN(n509) );
  XOR2_X1 U506 ( .A(n510), .B(n497), .Z(n451) );
  XOR2_X1 U507 ( .A(n511), .B(n512), .Z(n497) );
  XOR2_X1 U508 ( .A(n513), .B(n514), .Z(n512) );
  XNOR2_X1 U509 ( .A(n496), .B(n495), .ZN(n510) );
  OR2_X1 U510 ( .A1(n515), .A2(n516), .ZN(n495) );
  AND2_X1 U511 ( .A1(n517), .A2(n518), .ZN(n516) );
  AND2_X1 U512 ( .A1(n519), .A2(n520), .ZN(n515) );
  OR2_X1 U513 ( .A1(n518), .A2(n517), .ZN(n520) );
  OR2_X1 U514 ( .A1(n521), .A2(n522), .ZN(n496) );
  OR2_X1 U515 ( .A1(n523), .A2(n524), .ZN(n442) );
  OR2_X1 U516 ( .A1(n525), .A2(n526), .ZN(n523) );
  AND2_X1 U517 ( .A1(n440), .A2(n527), .ZN(n526) );
  AND2_X1 U518 ( .A1(n441), .A2(n527), .ZN(n525) );
  INV_X1 U519 ( .A(n439), .ZN(n527) );
  OR2_X1 U520 ( .A1(n528), .A2(n524), .ZN(n439) );
  INV_X1 U521 ( .A(n529), .ZN(n524) );
  OR2_X1 U522 ( .A1(n530), .A2(n531), .ZN(n529) );
  AND2_X1 U523 ( .A1(n530), .A2(n531), .ZN(n528) );
  OR2_X1 U524 ( .A1(n532), .A2(n533), .ZN(n531) );
  AND2_X1 U525 ( .A1(n534), .A2(n535), .ZN(n533) );
  AND2_X1 U526 ( .A1(n536), .A2(n537), .ZN(n532) );
  OR2_X1 U527 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U528 ( .A(n508), .B(n538), .Z(n530) );
  XOR2_X1 U529 ( .A(n507), .B(n506), .Z(n538) );
  OR2_X1 U530 ( .A1(n539), .A2(n522), .ZN(n506) );
  OR2_X1 U531 ( .A1(n540), .A2(n541), .ZN(n507) );
  AND2_X1 U532 ( .A1(n542), .A2(n543), .ZN(n541) );
  AND2_X1 U533 ( .A1(n544), .A2(n545), .ZN(n540) );
  OR2_X1 U534 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U535 ( .A(n546), .B(n519), .ZN(n508) );
  XNOR2_X1 U536 ( .A(n547), .B(n548), .ZN(n519) );
  XNOR2_X1 U537 ( .A(n549), .B(n550), .ZN(n547) );
  XNOR2_X1 U538 ( .A(n518), .B(n517), .ZN(n546) );
  OR2_X1 U539 ( .A1(n551), .A2(n552), .ZN(n517) );
  AND2_X1 U540 ( .A1(n553), .A2(n554), .ZN(n552) );
  AND2_X1 U541 ( .A1(n555), .A2(n556), .ZN(n551) );
  OR2_X1 U542 ( .A1(n554), .A2(n553), .ZN(n556) );
  OR2_X1 U543 ( .A1(n521), .A2(n557), .ZN(n518) );
  INV_X1 U544 ( .A(n432), .ZN(n441) );
  OR4_X1 U545 ( .A1(n430), .A2(n429), .A3(n440), .A4(n558), .ZN(n432) );
  AND2_X1 U546 ( .A1(n435), .A2(n436), .ZN(n558) );
  INV_X1 U547 ( .A(n559), .ZN(n440) );
  OR2_X1 U548 ( .A1(n435), .A2(n436), .ZN(n559) );
  OR2_X1 U549 ( .A1(n560), .A2(n561), .ZN(n436) );
  AND2_X1 U550 ( .A1(n562), .A2(n563), .ZN(n561) );
  AND2_X1 U551 ( .A1(n564), .A2(n565), .ZN(n560) );
  OR2_X1 U552 ( .A1(n563), .A2(n562), .ZN(n565) );
  XOR2_X1 U553 ( .A(n534), .B(n566), .Z(n435) );
  XOR2_X1 U554 ( .A(n537), .B(n535), .Z(n566) );
  OR2_X1 U555 ( .A1(n567), .A2(n522), .ZN(n535) );
  OR2_X1 U556 ( .A1(n568), .A2(n569), .ZN(n537) );
  AND2_X1 U557 ( .A1(n570), .A2(n571), .ZN(n569) );
  AND2_X1 U558 ( .A1(n572), .A2(n573), .ZN(n568) );
  OR2_X1 U559 ( .A1(n571), .A2(n570), .ZN(n573) );
  XOR2_X1 U560 ( .A(n542), .B(n574), .Z(n534) );
  XOR2_X1 U561 ( .A(n545), .B(n543), .Z(n574) );
  OR2_X1 U562 ( .A1(n539), .A2(n557), .ZN(n543) );
  OR2_X1 U563 ( .A1(n575), .A2(n576), .ZN(n545) );
  AND2_X1 U564 ( .A1(n577), .A2(n578), .ZN(n576) );
  AND2_X1 U565 ( .A1(n579), .A2(n580), .ZN(n575) );
  OR2_X1 U566 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U567 ( .A(n581), .B(n555), .ZN(n542) );
  XNOR2_X1 U568 ( .A(n582), .B(n583), .ZN(n555) );
  XNOR2_X1 U569 ( .A(n584), .B(n585), .ZN(n582) );
  XNOR2_X1 U570 ( .A(n554), .B(n553), .ZN(n581) );
  OR2_X1 U571 ( .A1(n586), .A2(n587), .ZN(n553) );
  AND2_X1 U572 ( .A1(n588), .A2(n589), .ZN(n587) );
  AND2_X1 U573 ( .A1(n590), .A2(n591), .ZN(n586) );
  OR2_X1 U574 ( .A1(n588), .A2(n589), .ZN(n590) );
  OR2_X1 U575 ( .A1(n521), .A2(n592), .ZN(n554) );
  OR2_X1 U576 ( .A1(n593), .A2(n594), .ZN(n429) );
  AND2_X1 U577 ( .A1(n428), .A2(n427), .ZN(n594) );
  AND2_X1 U578 ( .A1(n425), .A2(n595), .ZN(n593) );
  OR2_X1 U579 ( .A1(n427), .A2(n428), .ZN(n595) );
  OR2_X1 U580 ( .A1(n596), .A2(n522), .ZN(n428) );
  OR2_X1 U581 ( .A1(n597), .A2(n598), .ZN(n427) );
  AND2_X1 U582 ( .A1(n424), .A2(n423), .ZN(n598) );
  AND2_X1 U583 ( .A1(n421), .A2(n599), .ZN(n597) );
  OR2_X1 U584 ( .A1(n423), .A2(n424), .ZN(n599) );
  OR2_X1 U585 ( .A1(n596), .A2(n557), .ZN(n424) );
  OR2_X1 U586 ( .A1(n600), .A2(n601), .ZN(n423) );
  AND2_X1 U587 ( .A1(n481), .A2(n480), .ZN(n601) );
  AND2_X1 U588 ( .A1(n478), .A2(n602), .ZN(n600) );
  OR2_X1 U589 ( .A1(n481), .A2(n480), .ZN(n602) );
  OR2_X1 U590 ( .A1(n603), .A2(n604), .ZN(n480) );
  AND2_X1 U591 ( .A1(n477), .A2(n476), .ZN(n604) );
  AND2_X1 U592 ( .A1(n474), .A2(n605), .ZN(n603) );
  OR2_X1 U593 ( .A1(n477), .A2(n476), .ZN(n605) );
  OR2_X1 U594 ( .A1(n606), .A2(n607), .ZN(n476) );
  AND2_X1 U595 ( .A1(n473), .A2(n472), .ZN(n607) );
  AND2_X1 U596 ( .A1(n470), .A2(n608), .ZN(n606) );
  OR2_X1 U597 ( .A1(n473), .A2(n472), .ZN(n608) );
  OR2_X1 U598 ( .A1(n609), .A2(n610), .ZN(n472) );
  AND2_X1 U599 ( .A1(n469), .A2(n468), .ZN(n610) );
  AND2_X1 U600 ( .A1(n466), .A2(n611), .ZN(n609) );
  OR2_X1 U601 ( .A1(n469), .A2(n468), .ZN(n611) );
  INV_X1 U602 ( .A(n612), .ZN(n468) );
  OR2_X1 U603 ( .A1(n613), .A2(n596), .ZN(n469) );
  XOR2_X1 U604 ( .A(n614), .B(n615), .Z(n466) );
  OR2_X1 U605 ( .A1(n616), .A2(n596), .ZN(n473) );
  XOR2_X1 U606 ( .A(n617), .B(n618), .Z(n470) );
  XOR2_X1 U607 ( .A(n619), .B(n620), .Z(n618) );
  OR2_X1 U608 ( .A1(n621), .A2(n596), .ZN(n477) );
  XOR2_X1 U609 ( .A(n622), .B(n623), .Z(n474) );
  XOR2_X1 U610 ( .A(n624), .B(n625), .Z(n623) );
  OR2_X1 U611 ( .A1(n592), .A2(n596), .ZN(n481) );
  XOR2_X1 U612 ( .A(n626), .B(n627), .Z(n478) );
  XOR2_X1 U613 ( .A(n628), .B(n629), .Z(n627) );
  XOR2_X1 U614 ( .A(n630), .B(n631), .Z(n421) );
  XOR2_X1 U615 ( .A(n632), .B(n633), .Z(n631) );
  XOR2_X1 U616 ( .A(n634), .B(n635), .Z(n425) );
  XOR2_X1 U617 ( .A(n636), .B(n637), .Z(n635) );
  XOR2_X1 U618 ( .A(n564), .B(n638), .Z(n430) );
  XOR2_X1 U619 ( .A(n563), .B(n562), .Z(n638) );
  OR2_X1 U620 ( .A1(n639), .A2(n522), .ZN(n562) );
  OR2_X1 U621 ( .A1(n640), .A2(n641), .ZN(n563) );
  AND2_X1 U622 ( .A1(n637), .A2(n636), .ZN(n641) );
  AND2_X1 U623 ( .A1(n634), .A2(n642), .ZN(n640) );
  OR2_X1 U624 ( .A1(n636), .A2(n637), .ZN(n642) );
  OR2_X1 U625 ( .A1(n639), .A2(n557), .ZN(n637) );
  OR2_X1 U626 ( .A1(n643), .A2(n644), .ZN(n636) );
  AND2_X1 U627 ( .A1(n633), .A2(n632), .ZN(n644) );
  AND2_X1 U628 ( .A1(n630), .A2(n645), .ZN(n643) );
  OR2_X1 U629 ( .A1(n632), .A2(n633), .ZN(n645) );
  OR2_X1 U630 ( .A1(n639), .A2(n592), .ZN(n633) );
  OR2_X1 U631 ( .A1(n646), .A2(n647), .ZN(n632) );
  AND2_X1 U632 ( .A1(n629), .A2(n628), .ZN(n647) );
  AND2_X1 U633 ( .A1(n626), .A2(n648), .ZN(n646) );
  OR2_X1 U634 ( .A1(n629), .A2(n628), .ZN(n648) );
  OR2_X1 U635 ( .A1(n649), .A2(n650), .ZN(n628) );
  AND2_X1 U636 ( .A1(n625), .A2(n624), .ZN(n650) );
  AND2_X1 U637 ( .A1(n622), .A2(n651), .ZN(n649) );
  OR2_X1 U638 ( .A1(n625), .A2(n624), .ZN(n651) );
  OR2_X1 U639 ( .A1(n652), .A2(n653), .ZN(n624) );
  AND2_X1 U640 ( .A1(n620), .A2(n619), .ZN(n653) );
  AND2_X1 U641 ( .A1(n617), .A2(n654), .ZN(n652) );
  OR2_X1 U642 ( .A1(n620), .A2(n619), .ZN(n654) );
  OR2_X1 U643 ( .A1(n464), .A2(n655), .ZN(n619) );
  OR2_X1 U644 ( .A1(n656), .A2(n639), .ZN(n464) );
  OR2_X1 U645 ( .A1(n613), .A2(n639), .ZN(n620) );
  XNOR2_X1 U646 ( .A(n657), .B(n655), .ZN(n617) );
  OR2_X1 U647 ( .A1(n658), .A2(n567), .ZN(n655) );
  OR2_X1 U648 ( .A1(n656), .A2(n539), .ZN(n657) );
  OR2_X1 U649 ( .A1(n616), .A2(n639), .ZN(n625) );
  XNOR2_X1 U650 ( .A(n659), .B(n660), .ZN(n622) );
  XOR2_X1 U651 ( .A(n661), .B(n662), .Z(n659) );
  OR2_X1 U652 ( .A1(n621), .A2(n639), .ZN(n629) );
  XOR2_X1 U653 ( .A(n663), .B(n664), .Z(n626) );
  XOR2_X1 U654 ( .A(n665), .B(n666), .Z(n664) );
  XOR2_X1 U655 ( .A(n667), .B(n668), .Z(n630) );
  XOR2_X1 U656 ( .A(n669), .B(n670), .Z(n668) );
  XOR2_X1 U657 ( .A(n671), .B(n672), .Z(n634) );
  XOR2_X1 U658 ( .A(n673), .B(n674), .Z(n672) );
  XOR2_X1 U659 ( .A(n572), .B(n675), .Z(n564) );
  XOR2_X1 U660 ( .A(n571), .B(n570), .Z(n675) );
  OR2_X1 U661 ( .A1(n567), .A2(n557), .ZN(n570) );
  OR2_X1 U662 ( .A1(n676), .A2(n677), .ZN(n571) );
  AND2_X1 U663 ( .A1(n674), .A2(n673), .ZN(n677) );
  AND2_X1 U664 ( .A1(n671), .A2(n678), .ZN(n676) );
  OR2_X1 U665 ( .A1(n673), .A2(n674), .ZN(n678) );
  OR2_X1 U666 ( .A1(n567), .A2(n592), .ZN(n674) );
  OR2_X1 U667 ( .A1(n679), .A2(n680), .ZN(n673) );
  AND2_X1 U668 ( .A1(n670), .A2(n669), .ZN(n680) );
  AND2_X1 U669 ( .A1(n667), .A2(n681), .ZN(n679) );
  OR2_X1 U670 ( .A1(n669), .A2(n670), .ZN(n681) );
  OR2_X1 U671 ( .A1(n567), .A2(n621), .ZN(n670) );
  OR2_X1 U672 ( .A1(n682), .A2(n683), .ZN(n669) );
  AND2_X1 U673 ( .A1(n666), .A2(n665), .ZN(n683) );
  AND2_X1 U674 ( .A1(n663), .A2(n684), .ZN(n682) );
  OR2_X1 U675 ( .A1(n666), .A2(n665), .ZN(n684) );
  OR2_X1 U676 ( .A1(n685), .A2(n686), .ZN(n665) );
  AND2_X1 U677 ( .A1(n660), .A2(n661), .ZN(n686) );
  AND2_X1 U678 ( .A1(n687), .A2(n688), .ZN(n685) );
  OR2_X1 U679 ( .A1(n660), .A2(n661), .ZN(n687) );
  OR2_X1 U680 ( .A1(n689), .A2(n690), .ZN(n661) );
  AND2_X1 U681 ( .A1(n691), .A2(n692), .ZN(n689) );
  OR2_X1 U682 ( .A1(n691), .A2(n614), .ZN(n660) );
  OR2_X1 U683 ( .A1(n656), .A2(n567), .ZN(n614) );
  OR2_X1 U684 ( .A1(n616), .A2(n567), .ZN(n666) );
  XNOR2_X1 U685 ( .A(n693), .B(n694), .ZN(n663) );
  XOR2_X1 U686 ( .A(n695), .B(n690), .Z(n693) );
  INV_X1 U687 ( .A(n696), .ZN(n690) );
  XNOR2_X1 U688 ( .A(n697), .B(n698), .ZN(n667) );
  XNOR2_X1 U689 ( .A(n699), .B(n700), .ZN(n697) );
  XOR2_X1 U690 ( .A(n701), .B(n702), .Z(n671) );
  XOR2_X1 U691 ( .A(n703), .B(n704), .Z(n702) );
  XOR2_X1 U692 ( .A(n579), .B(n705), .Z(n572) );
  XOR2_X1 U693 ( .A(n578), .B(n577), .Z(n705) );
  OR2_X1 U694 ( .A1(n539), .A2(n592), .ZN(n577) );
  OR2_X1 U695 ( .A1(n706), .A2(n707), .ZN(n578) );
  AND2_X1 U696 ( .A1(n704), .A2(n703), .ZN(n707) );
  AND2_X1 U697 ( .A1(n701), .A2(n708), .ZN(n706) );
  OR2_X1 U698 ( .A1(n703), .A2(n704), .ZN(n708) );
  OR2_X1 U699 ( .A1(n539), .A2(n621), .ZN(n704) );
  OR2_X1 U700 ( .A1(n709), .A2(n710), .ZN(n703) );
  AND2_X1 U701 ( .A1(n698), .A2(n700), .ZN(n710) );
  AND2_X1 U702 ( .A1(n711), .A2(n699), .ZN(n709) );
  OR2_X1 U703 ( .A1(n698), .A2(n700), .ZN(n711) );
  OR2_X1 U704 ( .A1(n712), .A2(n713), .ZN(n700) );
  AND2_X1 U705 ( .A1(n694), .A2(n696), .ZN(n713) );
  AND2_X1 U706 ( .A1(n714), .A2(n695), .ZN(n712) );
  OR2_X1 U707 ( .A1(n715), .A2(n716), .ZN(n695) );
  INV_X1 U708 ( .A(n717), .ZN(n716) );
  AND2_X1 U709 ( .A1(n718), .A2(n719), .ZN(n715) );
  OR2_X1 U710 ( .A1(n720), .A2(n656), .ZN(n719) );
  OR2_X1 U711 ( .A1(n658), .A2(n521), .ZN(n718) );
  OR2_X1 U712 ( .A1(n694), .A2(n696), .ZN(n714) );
  OR2_X1 U713 ( .A1(n692), .A2(n691), .ZN(n696) );
  OR2_X1 U714 ( .A1(n658), .A2(n539), .ZN(n691) );
  OR2_X1 U715 ( .A1(n613), .A2(n539), .ZN(n694) );
  XNOR2_X1 U716 ( .A(n721), .B(n717), .ZN(n698) );
  XNOR2_X1 U717 ( .A(n722), .B(n723), .ZN(n721) );
  XNOR2_X1 U718 ( .A(n724), .B(n725), .ZN(n701) );
  XNOR2_X1 U719 ( .A(n726), .B(n727), .ZN(n724) );
  XNOR2_X1 U720 ( .A(n728), .B(n588), .ZN(n579) );
  XNOR2_X1 U721 ( .A(n729), .B(n730), .ZN(n588) );
  XNOR2_X1 U722 ( .A(n731), .B(n732), .ZN(n729) );
  XOR2_X1 U723 ( .A(n733), .B(n589), .Z(n728) );
  OR2_X1 U724 ( .A1(n734), .A2(n735), .ZN(n589) );
  AND2_X1 U725 ( .A1(n727), .A2(n726), .ZN(n735) );
  AND2_X1 U726 ( .A1(n725), .A2(n736), .ZN(n734) );
  OR2_X1 U727 ( .A1(n726), .A2(n727), .ZN(n736) );
  OR2_X1 U728 ( .A1(n737), .A2(n738), .ZN(n727) );
  AND2_X1 U729 ( .A1(n717), .A2(n723), .ZN(n738) );
  AND2_X1 U730 ( .A1(n739), .A2(n722), .ZN(n737) );
  OR2_X1 U731 ( .A1(n740), .A2(n741), .ZN(n722) );
  AND2_X1 U732 ( .A1(n742), .A2(n743), .ZN(n740) );
  OR2_X1 U733 ( .A1(n723), .A2(n717), .ZN(n739) );
  OR2_X1 U734 ( .A1(n692), .A2(n743), .ZN(n717) );
  OR2_X1 U735 ( .A1(n656), .A2(n521), .ZN(n692) );
  OR2_X1 U736 ( .A1(n521), .A2(n613), .ZN(n723) );
  OR2_X1 U737 ( .A1(n521), .A2(n616), .ZN(n726) );
  XNOR2_X1 U738 ( .A(n744), .B(n745), .ZN(n725) );
  XOR2_X1 U739 ( .A(n746), .B(n741), .Z(n744) );
  INV_X1 U740 ( .A(n747), .ZN(n741) );
  AND3_X1 U741 ( .A1(n462), .A2(n460), .A3(n461), .ZN(n463) );
  INV_X1 U742 ( .A(n748), .ZN(n461) );
  OR2_X1 U743 ( .A1(n749), .A2(n750), .ZN(n748) );
  AND2_X1 U744 ( .A1(n502), .A2(n501), .ZN(n750) );
  AND2_X1 U745 ( .A1(n499), .A2(n751), .ZN(n749) );
  OR2_X1 U746 ( .A1(n501), .A2(n502), .ZN(n751) );
  OR2_X1 U747 ( .A1(n720), .A2(n522), .ZN(n502) );
  OR2_X1 U748 ( .A1(n752), .A2(n753), .ZN(n501) );
  AND2_X1 U749 ( .A1(n514), .A2(n513), .ZN(n753) );
  AND2_X1 U750 ( .A1(n511), .A2(n754), .ZN(n752) );
  OR2_X1 U751 ( .A1(n513), .A2(n514), .ZN(n754) );
  OR2_X1 U752 ( .A1(n720), .A2(n557), .ZN(n514) );
  OR2_X1 U753 ( .A1(n755), .A2(n756), .ZN(n513) );
  AND2_X1 U754 ( .A1(n548), .A2(n550), .ZN(n756) );
  AND2_X1 U755 ( .A1(n757), .A2(n549), .ZN(n755) );
  OR2_X1 U756 ( .A1(n548), .A2(n550), .ZN(n757) );
  OR2_X1 U757 ( .A1(n758), .A2(n759), .ZN(n550) );
  AND2_X1 U758 ( .A1(n584), .A2(n585), .ZN(n759) );
  AND2_X1 U759 ( .A1(n583), .A2(n760), .ZN(n758) );
  OR2_X1 U760 ( .A1(n585), .A2(n584), .ZN(n760) );
  OR2_X1 U761 ( .A1(n761), .A2(n762), .ZN(n584) );
  AND2_X1 U762 ( .A1(n732), .A2(n731), .ZN(n762) );
  AND2_X1 U763 ( .A1(n730), .A2(n763), .ZN(n761) );
  OR2_X1 U764 ( .A1(n731), .A2(n732), .ZN(n763) );
  OR2_X1 U765 ( .A1(n720), .A2(n616), .ZN(n732) );
  OR2_X1 U766 ( .A1(n764), .A2(n765), .ZN(n731) );
  AND2_X1 U767 ( .A1(n745), .A2(n747), .ZN(n765) );
  AND2_X1 U768 ( .A1(n766), .A2(n746), .ZN(n764) );
  OR2_X1 U769 ( .A1(n767), .A2(n768), .ZN(n746) );
  AND2_X1 U770 ( .A1(n769), .A2(n770), .ZN(n767) );
  OR2_X1 U771 ( .A1(n656), .A2(n771), .ZN(n769) );
  OR2_X1 U772 ( .A1(n747), .A2(n745), .ZN(n766) );
  OR2_X1 U773 ( .A1(n720), .A2(n613), .ZN(n745) );
  OR2_X1 U774 ( .A1(n743), .A2(n742), .ZN(n747) );
  OR2_X1 U775 ( .A1(n656), .A2(n772), .ZN(n742) );
  OR2_X1 U776 ( .A1(n658), .A2(n720), .ZN(n743) );
  XOR2_X1 U777 ( .A(n773), .B(n768), .Z(n730) );
  INV_X1 U778 ( .A(n774), .ZN(n768) );
  OR2_X1 U779 ( .A1(n775), .A2(n776), .ZN(n773) );
  INV_X1 U780 ( .A(n777), .ZN(n776) );
  AND2_X1 U781 ( .A1(n778), .A2(n779), .ZN(n775) );
  OR2_X1 U782 ( .A1(n658), .A2(n771), .ZN(n778) );
  OR2_X1 U783 ( .A1(n720), .A2(n621), .ZN(n585) );
  XOR2_X1 U784 ( .A(n780), .B(n781), .Z(n583) );
  XOR2_X1 U785 ( .A(n782), .B(n783), .Z(n780) );
  XOR2_X1 U786 ( .A(n784), .B(n785), .Z(n548) );
  XOR2_X1 U787 ( .A(n786), .B(n787), .Z(n785) );
  XOR2_X1 U788 ( .A(n788), .B(n789), .Z(n511) );
  XOR2_X1 U789 ( .A(n790), .B(n791), .Z(n789) );
  XOR2_X1 U790 ( .A(n792), .B(n793), .Z(n499) );
  XOR2_X1 U791 ( .A(n794), .B(n795), .Z(n793) );
  XNOR2_X1 U792 ( .A(n796), .B(n484), .ZN(n460) );
  INV_X1 U793 ( .A(n797), .ZN(n484) );
  OR2_X1 U794 ( .A1(n798), .A2(n799), .ZN(n797) );
  AND2_X1 U795 ( .A1(n800), .A2(n801), .ZN(n799) );
  AND2_X1 U796 ( .A1(n802), .A2(n803), .ZN(n798) );
  OR2_X1 U797 ( .A1(n801), .A2(n800), .ZN(n802) );
  OR2_X1 U798 ( .A1(n771), .A2(n522), .ZN(n796) );
  XNOR2_X1 U799 ( .A(n800), .B(n804), .ZN(n462) );
  XOR2_X1 U800 ( .A(n801), .B(n803), .Z(n804) );
  OR2_X1 U801 ( .A1(n772), .A2(n522), .ZN(n803) );
  OR2_X1 U802 ( .A1(n805), .A2(n806), .ZN(n801) );
  AND2_X1 U803 ( .A1(n792), .A2(n794), .ZN(n806) );
  AND2_X1 U804 ( .A1(n807), .A2(n795), .ZN(n805) );
  OR2_X1 U805 ( .A1(n794), .A2(n792), .ZN(n807) );
  OR2_X1 U806 ( .A1(n592), .A2(n771), .ZN(n792) );
  OR2_X1 U807 ( .A1(n808), .A2(n809), .ZN(n794) );
  AND2_X1 U808 ( .A1(n788), .A2(n790), .ZN(n809) );
  AND2_X1 U809 ( .A1(n810), .A2(n791), .ZN(n808) );
  OR2_X1 U810 ( .A1(n621), .A2(n771), .ZN(n791) );
  OR2_X1 U811 ( .A1(n790), .A2(n788), .ZN(n810) );
  OR2_X1 U812 ( .A1(n772), .A2(n592), .ZN(n788) );
  OR2_X1 U813 ( .A1(n811), .A2(n812), .ZN(n790) );
  AND2_X1 U814 ( .A1(n784), .A2(n786), .ZN(n812) );
  AND2_X1 U815 ( .A1(n813), .A2(n787), .ZN(n811) );
  OR2_X1 U816 ( .A1(n772), .A2(n621), .ZN(n787) );
  OR2_X1 U817 ( .A1(n786), .A2(n784), .ZN(n813) );
  OR2_X1 U818 ( .A1(n616), .A2(n771), .ZN(n784) );
  OR2_X1 U819 ( .A1(n814), .A2(n815), .ZN(n786) );
  AND2_X1 U820 ( .A1(n781), .A2(n783), .ZN(n815) );
  AND2_X1 U821 ( .A1(n782), .A2(n816), .ZN(n814) );
  OR2_X1 U822 ( .A1(n783), .A2(n781), .ZN(n816) );
  OR2_X1 U823 ( .A1(n613), .A2(n771), .ZN(n781) );
  OR2_X1 U824 ( .A1(n772), .A2(n616), .ZN(n783) );
  AND2_X1 U825 ( .A1(n777), .A2(n774), .ZN(n782) );
  OR3_X1 U826 ( .A1(n656), .A2(n771), .A3(n770), .ZN(n774) );
  OR2_X1 U827 ( .A1(n658), .A2(n772), .ZN(n770) );
  OR3_X1 U828 ( .A1(n658), .A2(n771), .A3(n779), .ZN(n777) );
  OR2_X1 U829 ( .A1(n772), .A2(n613), .ZN(n779) );
  OR2_X1 U830 ( .A1(n557), .A2(n771), .ZN(n800) );
  INV_X1 U831 ( .A(b_0_), .ZN(n771) );
  XOR2_X1 U832 ( .A(b_7_), .B(a_7_), .Z(Result_add_7_) );
  OR3_X1 U833 ( .A1(n817), .A2(n818), .A3(n612), .ZN(Result_add_6_) );
  AND2_X1 U834 ( .A1(n615), .A2(Result_mul_15_), .ZN(n612) );
  AND3_X1 U835 ( .A1(n819), .A2(n658), .A3(b_6_), .ZN(n818) );
  INV_X1 U836 ( .A(a_6_), .ZN(n658) );
  AND2_X1 U837 ( .A1(n820), .A2(n639), .ZN(n817) );
  INV_X1 U838 ( .A(b_6_), .ZN(n639) );
  XOR2_X1 U839 ( .A(a_6_), .B(Result_mul_15_), .Z(n820) );
  OR3_X1 U840 ( .A1(n821), .A2(n822), .A3(n823), .ZN(Result_add_5_) );
  AND2_X1 U841 ( .A1(n662), .A2(n824), .ZN(n823) );
  INV_X1 U842 ( .A(n688), .ZN(n662) );
  AND2_X1 U843 ( .A1(n825), .A2(n567), .ZN(n822) );
  XOR2_X1 U844 ( .A(n824), .B(a_5_), .Z(n825) );
  AND3_X1 U845 ( .A1(n826), .A2(n613), .A3(b_5_), .ZN(n821) );
  XNOR2_X1 U846 ( .A(n827), .B(n828), .ZN(Result_add_4_) );
  AND2_X1 U847 ( .A1(n699), .A2(n829), .ZN(n828) );
  OR3_X1 U848 ( .A1(n830), .A2(n831), .A3(n832), .ZN(Result_add_3_) );
  AND2_X1 U849 ( .A1(n833), .A2(n733), .ZN(n832) );
  INV_X1 U850 ( .A(n591), .ZN(n733) );
  AND2_X1 U851 ( .A1(n834), .A2(n521), .ZN(n831) );
  XOR2_X1 U852 ( .A(a_3_), .B(n833), .Z(n834) );
  INV_X1 U853 ( .A(n835), .ZN(n833) );
  AND3_X1 U854 ( .A1(n835), .A2(n621), .A3(b_3_), .ZN(n830) );
  XNOR2_X1 U855 ( .A(n836), .B(n837), .ZN(Result_add_2_) );
  AND2_X1 U856 ( .A1(n549), .A2(n838), .ZN(n837) );
  OR3_X1 U857 ( .A1(n839), .A2(n840), .A3(n841), .ZN(Result_add_1_) );
  INV_X1 U858 ( .A(n842), .ZN(n841) );
  OR2_X1 U859 ( .A1(n843), .A2(n795), .ZN(n842) );
  AND2_X1 U860 ( .A1(n844), .A2(n772), .ZN(n840) );
  XOR2_X1 U861 ( .A(n557), .B(n843), .Z(n844) );
  AND3_X1 U862 ( .A1(n843), .A2(n557), .A3(b_1_), .ZN(n839) );
  XOR2_X1 U863 ( .A(n845), .B(n846), .Z(Result_add_0_) );
  XOR2_X1 U864 ( .A(n522), .B(b_0_), .Z(n846) );
  INV_X1 U865 ( .A(a_0_), .ZN(n522) );
  OR2_X1 U866 ( .A1(n847), .A2(n848), .ZN(n845) );
  AND2_X1 U867 ( .A1(n557), .A2(n772), .ZN(n848) );
  AND2_X1 U868 ( .A1(n843), .A2(n795), .ZN(n847) );
  OR2_X1 U869 ( .A1(n772), .A2(n557), .ZN(n795) );
  INV_X1 U870 ( .A(a_1_), .ZN(n557) );
  INV_X1 U871 ( .A(b_1_), .ZN(n772) );
  OR2_X1 U872 ( .A1(n849), .A2(n850), .ZN(n843) );
  INV_X1 U873 ( .A(n838), .ZN(n850) );
  OR2_X1 U874 ( .A1(a_2_), .A2(b_2_), .ZN(n838) );
  AND2_X1 U875 ( .A1(n836), .A2(n549), .ZN(n849) );
  OR2_X1 U876 ( .A1(n720), .A2(n592), .ZN(n549) );
  INV_X1 U877 ( .A(a_2_), .ZN(n592) );
  INV_X1 U878 ( .A(b_2_), .ZN(n720) );
  OR2_X1 U879 ( .A1(n851), .A2(n852), .ZN(n836) );
  AND2_X1 U880 ( .A1(n621), .A2(n521), .ZN(n852) );
  AND2_X1 U881 ( .A1(n835), .A2(n591), .ZN(n851) );
  OR2_X1 U882 ( .A1(n521), .A2(n621), .ZN(n591) );
  INV_X1 U883 ( .A(a_3_), .ZN(n621) );
  INV_X1 U884 ( .A(b_3_), .ZN(n521) );
  OR2_X1 U885 ( .A1(n853), .A2(n854), .ZN(n835) );
  INV_X1 U886 ( .A(n829), .ZN(n854) );
  OR2_X1 U887 ( .A1(a_4_), .A2(b_4_), .ZN(n829) );
  AND2_X1 U888 ( .A1(n827), .A2(n699), .ZN(n853) );
  OR2_X1 U889 ( .A1(n616), .A2(n539), .ZN(n699) );
  INV_X1 U890 ( .A(b_4_), .ZN(n539) );
  INV_X1 U891 ( .A(a_4_), .ZN(n616) );
  OR2_X1 U892 ( .A1(n855), .A2(n856), .ZN(n827) );
  AND2_X1 U893 ( .A1(n613), .A2(n567), .ZN(n856) );
  AND2_X1 U894 ( .A1(n826), .A2(n688), .ZN(n855) );
  OR2_X1 U895 ( .A1(n613), .A2(n567), .ZN(n688) );
  INV_X1 U896 ( .A(b_5_), .ZN(n567) );
  INV_X1 U897 ( .A(a_5_), .ZN(n613) );
  INV_X1 U898 ( .A(n824), .ZN(n826) );
  OR2_X1 U899 ( .A1(n857), .A2(n615), .ZN(n824) );
  AND2_X1 U900 ( .A1(a_6_), .A2(b_6_), .ZN(n615) );
  AND2_X1 U901 ( .A1(Result_mul_15_), .A2(n858), .ZN(n857) );
  OR2_X1 U902 ( .A1(a_6_), .A2(b_6_), .ZN(n858) );
  INV_X1 U903 ( .A(n819), .ZN(Result_mul_15_) );
  OR2_X1 U904 ( .A1(n656), .A2(n596), .ZN(n819) );
  INV_X1 U905 ( .A(b_7_), .ZN(n596) );
  INV_X1 U906 ( .A(a_7_), .ZN(n656) );
endmodule

