module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, 
        test_se, test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, 
        test_si4, test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, 
        test_so7, test_si8, test_so8, test_si9, test_so9, test_si10, test_so10
 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961, test_so1, test_so2, test_so3, test_so4, test_so5,
         test_so6, test_so7, test_so8, test_so9, test_so10;
  wire   g100, g101, g102, g103, g104, g1170, g1173, g1176, g1179, g1182,
         g1185, g1188, g1191, g1194, g1197, g1203, g18, g1960, g1961, g27, g28,
         g29, g30, g31, g41, g42, g43, g44, g45, g46, g47, g48, g5816, g82,
         g83, g84, g85, g8561, g8562, g8563, g8564, g8565, g8566, g86, g87,
         g872, g873, g88, g886, g889, g89, g892, g895, g898, g90, g901, g904,
         g907, g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g9451,
         g95, g96, g99, test_so10, g10722, g10664, g1289, g8943, g1882, n1663,
         g255, g312, g11257, g452, g7032, g123, g6830, g207, g8920, g713,
         g4340, g1153, n1686, g4239, g1744, g6538, g1558, g8887, g695, g11372,
         g461, n1594, g8260, g940, g11391, g976, g8432, g709, n1719, g6088,
         g1092, g6478, g1574, g6795, g1864, g11320, g369, g6500, g1580, g5392,
         g1736, g10663, n1637, g10782, n3065, g6216, g1424, g1737, g10858,
         g1672, g5914, g1077, g7590, g1231, g6656, g4, g6728, g5126, g1104,
         n1658, g7290, g1304, g6841, g243, g8041, g1499, g8766, g1444, n3064,
         g8019, g6545, g1543, g256, g315, g6533, g1534, g8820, g622, n1713,
         g8941, g1927, g10859, g1660, g6922, g278, g8772, g1436, g8433, g718,
         g6526, g10793, g554, g11333, g496, n1689, g11392, g981, n1720, g794,
         g829, g6093, g1095, g8889, g704, g7302, g1265, g6525, g1786, g8429,
         g682, g7292, g1296, g6621, g7134, n3062, g260, g327, g6333, g1389,
         n1603, g6826, g1371, g1955, g1956, g10860, g1675, g11483, g354, g6392,
         g113, g7626, g639, n1692, g10866, g1684, g8193, g1639, g6983, g1791,
         n1702, g6839, g248, g4076, g1707, g4293, g1759, g11482, g351, g6507,
         g1604, g6096, g1098, g8250, g932, g8282, g1896, g8435, g736, g6924,
         g1019, g6819, n3061, g746, g745, g6244, g1419, n1602, g6627, g32,
         n1865, g6071, g1086, g8046, g1486, g10707, g1730, g6198, g1504, g8051,
         g1470, g8024, g822, g10862, g1678, g8050, g174, g7133, g1766, g7930,
         g1801, g6832, g186, g11308, g959, g6918, g8769, g1407, g6909, g1868,
         g4940, g5404, g1718, n1611, g11265, g396, g6930, g1015, g10726, n1650,
         g4891, n3059, n1874, g6224, g1415, g7586, g1227, g10770, g1721, n3058,
         n3057, g6934, g284, g11256, g426, g6824, g219, g1360, n3056, g6126,
         g806, g8767, g1428, g6546, g1564, g4238, g1741, g6823, g225, g6928,
         g281, g11602, g1308, g9721, g611, n1609, g4890, n3055, n1586, g1217,
         g6524, g1589, g8045, g1466, g6469, g1571, g6471, g1861, g6821, n3054,
         g11514, g1448, g4480, g1133, n1706, g11610, g1333, g7843, g153,
         g11310, g962, g5536, g11331, g486, n1621, g11380, g471, n1606, g6838,
         g1397, g8288, g1950, g755, g756, n3053, g10855, g1101, g549, g10898,
         g105, g10865, g1669, g6822, g6528, g1531, g6180, g1458, n1703, g10718,
         g572, g6912, g1011, g10719, n3051, g6234, g1411, g6099, g1074, g11259,
         g444, g8039, g1474, g6059, g1080, g5396, g1713, n1610, g262, g333,
         g6906, g269, g11266, g401, g11294, g1857, n1682, g5421, g9, g8649,
         g664, g11312, g965, g6840, g1400, g254, g309, g7202, g814, g6834,
         g231, g10795, g557, g875, g869, g6831, g1383, g8060, g158, g4893,
         g627, n1701, g7244, g1023, g6026, g259, n3050, g11608, g1327, g7660,
         g654, g6911, g293, g11640, g1346, g8777, g1633, g4274, g1753, g1508,
         n1707, g7297, g1240, g11326, g538, g11269, g416, g11325, g542, g10864,
         g1681, g11290, g374, g10798, g563, g8284, g1914, g11328, g530, g10800,
         g575, g8944, g1936, n1694, g7183, g4465, g1356, g1317, g11484, g357,
         g11263, g386, g6501, g1601, g6757, g166, g11334, g501, n1690, g6042,
         g8384, g1840, g6653, g257, g318, g5763, g5849, n3048, g6929, g302,
         g11488, g342, g7299, g1250, g4330, g1163, g1958, n3047, g7257, g1032,
         g8775, g1432, g5770, g1453, n1628, g11486, g363, g261, g330, g4338,
         g1157, g4500, n3046, g10721, n3045, g8147, g928, g6038, g11337, g516,
         n1620, g6045, g7191, g826, g861, g8774, g1627, g7293, g1292, g6907,
         g290, g4903, n3044, n1873, g6123, g6506, g1583, g11376, g466, n1646,
         g6542, g1561, g6551, g1546, g6901, g287, g10797, g560, g8505, g617,
         n1645, n1631, g11647, g336, g11340, g456, n1641, g253, g305, n1681,
         g11625, g345, g636, g8, g6502, N599, g6049, g8945, g1945, n1697,
         g4231, g1738, g8040, g1478, n3042, g6155, g1690, n1653, g8043, g1482,
         g5173, g1110, n1677, g6916, g296, g10861, g1663, g8431, g700, g4309,
         g1762, g11485, g360, g6334, g192, g10767, g1657, g8923, g722, n1693,
         g7189, g10799, g566, g6747, n3041, g6080, g1089, g3381, g5910, g1071,
         g11393, g986, n1722, g11349, g971, g6439, g143, g9266, g1814, n1608,
         g1212, g8940, g1918, g7705, g9269, g1822, n1643, g6820, g237, g8042,
         g1462, g6759, g178, g11487, g366, g802, g837, g9124, g599, n1644,
         g11293, g1854, g11298, g944, g8287, g1941, g8047, g170, g6205, g1520,
         n1710, g8885, g686, n1676, g11305, g953, g5556, n3040, g2478, g1765,
         g10711, g1733, g7303, g5194, g1610, g7541, g1796, n1626, g11607,
         g1324, g6541, g1540, g6827, n3038, g11332, g491, n1691, g4902, n3037,
         g6828, g213, g6516, g1781, n1659, g8938, g1900, n1675, g7298, g1245,
         n3036, g6672, n3035, g8048, g148, g798, g833, g8285, g1923, n1718,
         g8254, g936, g11604, g1314, g849, g11636, g1336, g6910, g272, g8173,
         g1806, g8245, n1716, g8281, g1887, g10724, n3034, g11314, g968, g4905,
         n3033, g4484, g1137, n1597, g8937, g1891, n1657, g7300, g1255, g6002,
         n1588, g874, g9110, g591, n1607, g8926, g731, n1696, g8631, g7632,
         g1218, g9150, g605, n1593, g6531, g6786, g182, g11303, g950, g4477,
         g1129, n1705, g857, g11258, g448, g9272, g1828, n1605, g10773, g1727,
         g6470, g1592, g5083, g1703, g8286, g1932, g8773, g1624, g6054, g11260,
         g440, g11338, g476, n1599, g5918, g119, n1613, g8922, g668, n1662,
         g8049, g139, g4342, g1149, n1685, g10720, n3031, g6755, n3030, g6897,
         g263, g7709, g818, g4255, g1747, g5543, n1622, g6915, g275, g6513,
         g1524, g6480, g1577, g6733, g810, g11264, g391, g8973, g658, n1615,
         g6833, g1386, g5996, n1587, g4473, g1125, n1708, g5755, g201, n1619,
         g7295, g1280, n1862, g6068, g1083, g7137, g650, n1709, g8779, g1636,
         g853, g11270, g421, g5529, g11306, g956, g11291, g378, g4283, g1756,
         g841, g6894, g1027, g6902, g1003, g8765, g1403, g4498, g1145, n1617,
         g5148, g1107, n1614, g7581, g1223, g11267, g406, g10936, g1811,
         g10784, n3029, g10765, g1654, g6332, g197, n1678, g6479, g1595, g6537,
         g1537, g8434, g727, g6908, g6243, n1717, g11324, g481, n1680, n1647,
         g11609, g1330, g845, g8244, g8194, g1512, n3027, g8052, g1490, g4325,
         g1166, g11481, g348, n3026, g7301, g1260, g6035, g8059, g131, n3025,
         g6015, g258, g11330, g521, n1698, g11605, g1318, g8921, g1872, n1616,
         g8883, g677, n1656, n3024, g6523, g1549, g11300, g947, g9555, g1834,
         n1655, g6481, g1598, g4471, g1121, n1618, g11606, g1321, g11335, g506,
         n1600, g10791, g546, g8939, g1909, g6529, g1552, g10776, g1687, g6514,
         g1586, g324, g4490, g1141, n1660, g11639, g1341, g4089, g1710, g10785,
         n3023, g6179, n3022, g8053, g135, g11329, g525, n1695, g6515, g1607,
         g321, g7204, g11443, g1275, g11603, g8770, g1615, g11292, g382, g6331,
         n3020, g6900, g266, g7294, g1284, n1864, g6829, n3019, g8428, g673,
         n3018, g8054, g162, g11268, g411, g11262, g431, n1876, g8283, g1905,
         g6193, g1515, n1627, g8776, g1630, g7143, g6898, g991, n1871, g7291,
         g1300, g11478, g339, g6000, g4264, g1750, g8768, g1440, g10863, g1666,
         g6522, g1528, g11641, g1351, n1721, g10780, n3017, g8044, g127, n1704,
         g11579, g1618, g7296, g1235, g6923, g299, g11261, g435, n1878, g6638,
         g6534, g1555, g6895, g995, g8771, g1621, g4506, n3016, g7441, g643,
         n1612, g8055, g1494, g6468, g1567, g8430, g691, g11327, g534, g6508,
         g1776, n1715, g10717, g569, g4334, g1160, n1585, g6679, g1, g11336,
         g511, n1679, g10771, g1724, g5445, g12, g8559, g1878, g7219, g5390,
         n1654, n1512, n1486, n1485, n1545, n1530, n1420, n1855, n1239, n1566,
         n1567, n1479, n1480, n1478, n1137, n1195, n1404, n1229, n1262, n1227,
         n1450, n916, n822, n958, n918, n1159, n812, n1056, n1258, n817, n837,
         n804, n1016, n1380, n926, n1385, n1391, n1564, n1231, n1226, n1232,
         n1260, n1107, n1154, n1093, n1214, n931, n962, n902, n1193, n1153,
         n1125, n1099, n917, n857, n806, n808, n1097, n1123, n1151, n1090,
         n1161, n967, n921, n898, n1055, n1150, n1096, n1098, n1213, n1152,
         n836, n838, Tg1_OUT1, Tg1_OUT2, Tg1_OUT3, Tg1_OUT4, Tg1_OUT5,
         Tg1_OUT6, Tg1_OUT7, Tg1_OUT8, Tg2_OUT1, Tg2_OUT2, Tg2_OUT3, Tg2_OUT4,
         Tg2_OUT5, Tg2_OUT6, Tg2_OUT7, Tg2_OUT8, test_se_NOT, Trigger_select,
         n1, n6, n19, n51, n59, n60, n72, n78, n102, n145, n147, n179, n180,
         n233, n238, n256, n363, n366, n386, n438, n493, n495, n628, n633,
         n650, n652, n655, n656, n660, n661, n665, n666, n3084, n3085, n3107,
         n3108, n3128, n3129, n3130, n3136, n3175, n3193, n3194, n3200, n3218,
         n3219, n3220, n3221, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3300, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3365, n3366, n3367, n3368, n3369,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, U1586_n1, U1754_n1, U1798_n1, U1839_n1,
         U1843_n1, U1877_n1, U1908_n1, U1909_n1, U1987_n1, U2031_n1, U2035_n1,
         U2418_n1, U2468_n1, U2478_n1, U2488_n1, U2533_n1, U2534_n1, U2639_n1,
         U2641_n1, U2654_n1, U2658_n1, U2683_n1, U2699_n1, U2846_n1, U2847_n1,
         U2848_n1, U2859_n1, U2860_n1, U2861_n1, U2867_n1, U2879_n1, U2881_n1,
         U2882_n1, U2883_n1, U2884_n1, U2885_n1, U2886_n1, U2887_n1, U2888_n1,
         U2889_n1, U2890_n1, U2891_n1, U2892_n1, U2893_n1, U2894_n1, U2895_n1,
         U2896_n1, U2897_n1, U2898_n1, U2899_n1, U2900_n1, U2901_n1, U2902_n1,
         U3090_n1, U3092_n1, U3094_n1, U3096_n1, U3098_n1, U3124_n1, U3171_n1;
  assign g11489 = 1'b0;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g4205 = g1170;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4206 = g1197;
  assign g4208 = g1203;
  assign g2355 = g18;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g7744 = g27;
  assign g6285 = g28;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g8271 = g5816;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6920 = g8561;
  assign g6926 = g8562;
  assign g6932 = g8563;
  assign g6942 = g8564;
  assign g6949 = g8565;
  assign g6955 = g8566;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g5101 = g872;
  assign g8061 = g872;
  assign g5105 = g873;
  assign g8062 = g873;
  assign g6270 = g88;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g6271 = g89;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g6272 = g90;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g6273 = g91;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g6274 = g92;
  assign g4204 = g922;
  assign g4196 = g925;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g9961 = g9451;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g8984 = test_so10;

  SDFFX1 DFF_0_Q_reg ( .D(n1), .SI(test_si1), .SE(n3475), .CLK(n3515), .Q(
        g1289), .QN(n3323) );
  SDFFX1 DFF_1_Q_reg ( .D(g8943), .SI(g1289), .SE(n3430), .CLK(n3537), .Q(
        g1882), .QN(n1663) );
  SDFFX1 DFF_2_Q_reg ( .D(g255), .SI(g1882), .SE(n3393), .CLK(n3555), .Q(g312), 
        .QN(n3276) );
  SDFFX1 DFF_3_Q_reg ( .D(g11257), .SI(g312), .SE(n3454), .CLK(n3525), .Q(g452) );
  SDFFX1 DFF_4_Q_reg ( .D(g7032), .SI(g452), .SE(n3464), .CLK(n3520), .Q(g123)
         );
  SDFFX1 DFF_5_Q_reg ( .D(g6830), .SI(g123), .SE(n3463), .CLK(n3520), .Q(g207), 
        .QN(n3358) );
  SDFFX1 DFF_6_Q_reg ( .D(g8920), .SI(g207), .SE(n3467), .CLK(n3519), .Q(g713), 
        .QN(n3348) );
  SDFFX1 DFF_7_Q_reg ( .D(g4340), .SI(g713), .SE(n3467), .CLK(n3519), .Q(g1153), .QN(n1686) );
  SDFFX1 DFF_9_Q_reg ( .D(g4239), .SI(g1153), .SE(n3397), .CLK(n3553), .Q(
        g1744) );
  SDFFX1 DFF_10_Q_reg ( .D(g6538), .SI(g1744), .SE(n3397), .CLK(n3554), .Q(
        g1558) );
  SDFFX1 DFF_11_Q_reg ( .D(g8887), .SI(g1558), .SE(n3459), .CLK(n3523), .Q(
        g695), .QN(n3329) );
  SDFFX1 DFF_12_Q_reg ( .D(g11372), .SI(g695), .SE(n3458), .CLK(n3523), .Q(
        g461), .QN(n1594) );
  SDFFX1 DFF_13_Q_reg ( .D(g8260), .SI(g461), .SE(n3442), .CLK(n3531), .Q(g940) );
  SDFFX1 DFF_14_Q_reg ( .D(g11391), .SI(g940), .SE(n3442), .CLK(n3531), .Q(
        g976), .QN(n3372) );
  SDFFX1 DFF_15_Q_reg ( .D(g8432), .SI(g976), .SE(n3468), .CLK(n3518), .Q(g709), .QN(n1719) );
  SDFFX1 DFF_16_Q_reg ( .D(g6088), .SI(g709), .SE(n3436), .CLK(n3534), .Q(
        g1092) );
  SDFFX1 DFF_17_Q_reg ( .D(g6478), .SI(g1092), .SE(n3418), .CLK(n3543), .Q(
        g1574) );
  SDFFX1 DFF_18_Q_reg ( .D(g6795), .SI(g1574), .SE(n3418), .CLK(n3543), .Q(
        g1864), .QN(n3316) );
  SDFFX1 DFF_19_Q_reg ( .D(g11320), .SI(g1864), .SE(n3396), .CLK(n3554), .Q(
        g369), .QN(n3374) );
  SDFFX1 DFF_20_Q_reg ( .D(g6500), .SI(g369), .SE(n3435), .CLK(n3534), .Q(
        g1580) );
  SDFFX1 DFF_21_Q_reg ( .D(g5392), .SI(g1580), .SE(n3435), .CLK(n3535), .Q(
        g1736) );
  SDFFX1 DFF_22_Q_reg ( .D(g10663), .SI(g1736), .SE(n3435), .CLK(n3535), .Q(
        n1637) );
  SDFFX1 DFF_23_Q_reg ( .D(g10782), .SI(n1637), .SE(n3435), .CLK(n3535), .Q(
        n3065) );
  SDFFX1 DFF_24_Q_reg ( .D(g6216), .SI(n3065), .SE(n3434), .CLK(n3535), .Q(
        g1424) );
  SDFFX1 DFF_25_Q_reg ( .D(g1736), .SI(g1424), .SE(n3434), .CLK(n3535), .Q(
        g1737), .QN(n3328) );
  SDFFX1 DFF_26_Q_reg ( .D(g10858), .SI(g1737), .SE(n3419), .CLK(n3542), .Q(
        g1672) );
  SDFFX1 DFF_27_Q_reg ( .D(g5914), .SI(g1672), .SE(n3446), .CLK(n3529), .Q(
        g1077) );
  SDFFX1 DFF_28_Q_reg ( .D(g7590), .SI(g1077), .SE(n3408), .CLK(n3548), .Q(
        g1231), .QN(n3361) );
  SDFFX1 DFF_29_Q_reg ( .D(g6656), .SI(g1231), .SE(n3466), .CLK(n3519), .Q(g4)
         );
  SDFFX1 DFF_30_Q_reg ( .D(g6728), .SI(g4), .SE(n3466), .CLK(n3519), .Q(g4177)
         );
  SDFFX1 DFF_31_Q_reg ( .D(g5126), .SI(g4177), .SE(n3466), .CLK(n3519), .Q(
        g1104), .QN(n1658) );
  SDFFX1 DFF_32_Q_reg ( .D(g7290), .SI(g1104), .SE(n3461), .CLK(n3522), .Q(
        g1304), .QN(n3235) );
  SDFFX1 DFF_33_Q_reg ( .D(g6841), .SI(g1304), .SE(n3430), .CLK(n3537), .Q(
        g243) );
  SDFFX1 DFF_34_Q_reg ( .D(g8041), .SI(g243), .SE(n3466), .CLK(n3519), .Q(
        g1499), .QN(n3271) );
  SDFFX1 DFF_36_Q_reg ( .D(g8766), .SI(g1499), .SE(n3438), .CLK(n3533), .Q(
        g1444), .QN(n3311) );
  SDFFX1 DFF_37_Q_reg ( .D(n19), .SI(g1444), .SE(n3438), .CLK(n3533), .Q(n3064) );
  SDFFX1 DFF_38_Q_reg ( .D(g8019), .SI(n3064), .SE(n3395), .CLK(n3555), .Q(
        g4180), .QN(n3363) );
  SDFFX1 DFF_39_Q_reg ( .D(g6545), .SI(g4180), .SE(n3395), .CLK(n3555), .Q(
        g1543) );
  SDFFX1 DFF_41_Q_reg ( .D(g256), .SI(g1543), .SE(n3463), .CLK(n3520), .Q(g315), .QN(n3295) );
  SDFFX1 DFF_42_Q_reg ( .D(g6533), .SI(g315), .SE(n3417), .CLK(n3543), .Q(
        g1534) );
  SDFFX1 DFF_43_Q_reg ( .D(g8820), .SI(g1534), .SE(n3417), .CLK(n3543), .Q(
        g622), .QN(n1713) );
  SDFFX1 DFF_44_Q_reg ( .D(g8941), .SI(g622), .SE(n3393), .CLK(n3555), .Q(
        g1927), .QN(n3347) );
  SDFFX1 DFF_45_Q_reg ( .D(g10859), .SI(g1927), .SE(n3457), .CLK(n3523), .Q(
        g1660) );
  SDFFX1 DFF_46_Q_reg ( .D(g6922), .SI(g1660), .SE(n3457), .CLK(n3523), .Q(
        g278) );
  SDFFX1 DFF_47_Q_reg ( .D(g8772), .SI(g278), .SE(n3438), .CLK(n3533), .Q(
        g1436), .QN(n3308) );
  SDFFX1 DFF_48_Q_reg ( .D(g8433), .SI(g1436), .SE(n3468), .CLK(n3518), .Q(
        g718), .QN(n3175) );
  SDFFX1 DFF_49_Q_reg ( .D(g6526), .SI(g718), .SE(n3427), .CLK(n3539), .Q(
        g8985) );
  SDFFX1 DFF_50_Q_reg ( .D(g10793), .SI(g8985), .SE(n3423), .CLK(n3541), .Q(
        g554) );
  SDFFX1 DFF_51_Q_reg ( .D(g11333), .SI(g554), .SE(n3422), .CLK(n3541), .Q(
        g496), .QN(n1689) );
  SDFFX1 DFF_52_Q_reg ( .D(g11392), .SI(g496), .SE(n3469), .CLK(n3517), .Q(
        g981), .QN(n1720) );
  SDFFX1 DFF_53_Q_reg ( .D(n3376), .SI(g981), .SE(n3470), .CLK(n3517), .Q(
        g3007) );
  SDFFX1 DFF_54_Q_reg ( .D(g1713), .SI(g3007), .SE(n3415), .CLK(n3545), .Q(
        test_so1), .QN(n3388) );
  SDFFX1 DFF_55_Q_reg ( .D(g794), .SI(test_si2), .SE(n3440), .CLK(n3532), .Q(
        g829) );
  SDFFX1 DFF_56_Q_reg ( .D(g6093), .SI(g829), .SE(n3390), .CLK(n3557), .Q(
        g1095) );
  SDFFX1 DFF_57_Q_reg ( .D(g8889), .SI(g1095), .SE(n3390), .CLK(n3557), .Q(
        g704), .QN(n3275) );
  SDFFX1 DFF_58_Q_reg ( .D(g7302), .SI(g704), .SE(n3461), .CLK(n3522), .Q(
        g1265), .QN(n3231) );
  SDFFX1 DFF_59_Q_reg ( .D(g6525), .SI(g1265), .SE(n3406), .CLK(n3549), .Q(
        g1786), .QN(n3332) );
  SDFFX1 DFF_60_Q_reg ( .D(g8429), .SI(g1786), .SE(n3467), .CLK(n3518), .Q(
        g682), .QN(n3344) );
  SDFFX1 DFF_61_Q_reg ( .D(g7292), .SI(g682), .SE(n3460), .CLK(n3522), .Q(
        g1296), .QN(n3233) );
  SDFFX1 DFF_62_Q_reg ( .D(g104), .SI(g1296), .SE(n3460), .CLK(n3522), .Q(
        g2602) );
  SDFFX1 DFF_63_Q_reg ( .D(g6621), .SI(g2602), .SE(n3427), .CLK(n3539), .Q(
        g8977) );
  SDFFX1 DFF_64_Q_reg ( .D(g7134), .SI(g8977), .SE(n3433), .CLK(n3536), .Q(
        n3062), .QN(n5996) );
  SDFFX1 DFF_65_Q_reg ( .D(g260), .SI(n3062), .SE(n3432), .CLK(n3536), .Q(g327), .QN(n3261) );
  SDFFX1 DFF_66_Q_reg ( .D(g6333), .SI(g327), .SE(n3432), .CLK(n3536), .Q(
        g1389), .QN(n1603) );
  SDFFX1 DFF_67_Q_reg ( .D(g6826), .SI(g1389), .SE(n3432), .CLK(n3536), .Q(
        g1371) );
  SDFFX1 DFF_68_Q_reg ( .D(g1955), .SI(g1371), .SE(n3432), .CLK(n3536), .Q(
        g1956) );
  SDFFX1 DFF_69_Q_reg ( .D(g10860), .SI(g1956), .SE(n3399), .CLK(n3552), .Q(
        g1675) );
  SDFFX1 DFF_70_Q_reg ( .D(g11483), .SI(g1675), .SE(n3443), .CLK(n3531), .Q(
        g354) );
  SDFFX1 DFF_71_Q_reg ( .D(g6392), .SI(g354), .SE(n3443), .CLK(n3531), .Q(g113) );
  SDFFX1 DFF_72_Q_reg ( .D(g7626), .SI(g113), .SE(n3459), .CLK(n3523), .Q(g639), .QN(n1692) );
  SDFFX1 DFF_73_Q_reg ( .D(g10866), .SI(g639), .SE(n3401), .CLK(n3551), .Q(
        g1684) );
  SDFFX1 DFF_74_Q_reg ( .D(g8193), .SI(g1684), .SE(n3451), .CLK(n3527), .Q(
        g1639) );
  SDFFX1 DFF_75_Q_reg ( .D(g6983), .SI(g1639), .SE(n3406), .CLK(n3549), .Q(
        g1791), .QN(n1702) );
  SDFFX1 DFF_76_Q_reg ( .D(g6839), .SI(g1791), .SE(n3431), .CLK(n3536), .Q(
        g248) );
  SDFFX1 DFF_77_Q_reg ( .D(g4076), .SI(g248), .SE(n3431), .CLK(n3537), .Q(
        g1707), .QN(n3327) );
  SDFFX1 DFF_78_Q_reg ( .D(g4293), .SI(g1707), .SE(n3396), .CLK(n3554), .Q(
        g1759) );
  SDFFX1 DFF_79_Q_reg ( .D(g11482), .SI(g1759), .SE(n3392), .CLK(n3556), .Q(
        g351) );
  SDFFX1 DFF_80_Q_reg ( .D(g1956), .SI(g351), .SE(n3392), .CLK(n3556), .Q(
        g1957) );
  SDFFX1 DFF_81_Q_reg ( .D(g6507), .SI(g1957), .SE(n3391), .CLK(n3556), .Q(
        g1604) );
  SDFFX1 DFF_82_Q_reg ( .D(g6096), .SI(g1604), .SE(n3445), .CLK(n3530), .Q(
        g1098) );
  SDFFX1 DFF_83_Q_reg ( .D(g8250), .SI(g1098), .SE(n3442), .CLK(n3531), .Q(
        g932) );
  SDFFX1 DFF_85_Q_reg ( .D(g8282), .SI(g932), .SE(n3451), .CLK(n3526), .Q(
        g1896), .QN(n3343) );
  SDFFX1 DFF_86_Q_reg ( .D(g8435), .SI(g1896), .SE(n3468), .CLK(n3518), .Q(
        g736), .QN(n3287) );
  SDFFX1 DFF_87_Q_reg ( .D(g6924), .SI(g736), .SE(n3445), .CLK(n3530), .Q(
        g1019), .QN(n3221) );
  SDFFX1 DFF_88_Q_reg ( .D(g6819), .SI(g1019), .SE(n3444), .CLK(n3530), .Q(
        n3061), .QN(n6000) );
  SDFFX1 DFF_89_Q_reg ( .D(g746), .SI(n3061), .SE(n3428), .CLK(n3538), .Q(g745), .QN(n3128) );
  SDFFX1 DFF_90_Q_reg ( .D(g6244), .SI(g745), .SE(n3428), .CLK(n3538), .Q(
        g1419), .QN(n1602) );
  SDFFX1 DFF_91_Q_reg ( .D(g6627), .SI(g1419), .SE(n3427), .CLK(n3539), .Q(
        g8979) );
  SDFFX1 DFF_92_Q_reg ( .D(n3375), .SI(g8979), .SE(n3465), .CLK(n3520), .Q(g32), .QN(n3389) );
  SDFFX1 DFF_93_Q_reg ( .D(g3007), .SI(g32), .SE(n3465), .CLK(n3520), .Q(n1865), .QN(n6002) );
  SDFFX1 DFF_94_Q_reg ( .D(g6071), .SI(n1865), .SE(n3464), .CLK(n3520), .Q(
        g1086) );
  SDFFX1 DFF_95_Q_reg ( .D(g8046), .SI(g1086), .SE(n3465), .CLK(n3519), .Q(
        g1486), .QN(n3244) );
  SDFFX1 DFF_96_Q_reg ( .D(g10707), .SI(g1486), .SE(n3419), .CLK(n3543), .Q(
        g1730) );
  SDFFX1 DFF_97_Q_reg ( .D(g6198), .SI(g1730), .SE(n3419), .CLK(n3543), .Q(
        g1504) );
  SDFFX1 DFF_98_Q_reg ( .D(g8051), .SI(g1504), .SE(n3450), .CLK(n3527), .Q(
        g1470), .QN(n3282) );
  SDFFX1 DFF_99_Q_reg ( .D(g8024), .SI(g1470), .SE(n3425), .CLK(n3539), .Q(
        g822), .QN(n3335) );
  SDFFX1 DFF_100_Q_reg ( .D(g29), .SI(g822), .SE(n3425), .CLK(n3540), .Q(g2609) );
  SDFFX1 DFF_101_Q_reg ( .D(g10862), .SI(g2609), .SE(n3393), .CLK(n3556), .Q(
        g1678) );
  SDFFX1 DFF_102_Q_reg ( .D(g8050), .SI(g1678), .SE(n3457), .CLK(n3524), .Q(
        g174), .QN(n3321) );
  SDFFX1 DFF_103_Q_reg ( .D(g7133), .SI(g174), .SE(n3414), .CLK(n3545), .Q(
        g1766), .QN(n3340) );
  SDFFX1 DFF_104_Q_reg ( .D(g7930), .SI(g1766), .SE(n3405), .CLK(n3549), .Q(
        g1801), .QN(n3319) );
  SDFFX1 DFF_105_Q_reg ( .D(g6832), .SI(g1801), .SE(n3405), .CLK(n3549), .Q(
        g186) );
  SDFFX1 DFF_106_Q_reg ( .D(g11308), .SI(g186), .SE(n3392), .CLK(n3556), .Q(
        g959) );
  SDFFX1 DFF_108_Q_reg ( .D(g6918), .SI(g959), .SE(n3390), .CLK(n3557), .Q(
        test_so2), .QN(n3385) );
  SDFFX1 DFF_109_Q_reg ( .D(g8769), .SI(test_si3), .SE(n3402), .CLK(n3551), 
        .Q(g1407) );
  SDFFX1 DFF_111_Q_reg ( .D(g6909), .SI(g1407), .SE(n3423), .CLK(n3540), .Q(
        g1868) );
  SDFFX1 DFF_112_Q_reg ( .D(g4940), .SI(g1868), .SE(n3423), .CLK(n3541), .Q(
        g4173), .QN(n3351) );
  SDFFX1 DFF_113_Q_reg ( .D(g5404), .SI(g4173), .SE(n3423), .CLK(n3541), .Q(
        g1718), .QN(n1611) );
  SDFFX1 DFF_114_Q_reg ( .D(g11265), .SI(g1718), .SE(n3455), .CLK(n3524), .Q(
        g396), .QN(n3258) );
  SDFFX1 DFF_115_Q_reg ( .D(g6930), .SI(g396), .SE(n3433), .CLK(n3535), .Q(
        g1015), .QN(n3220) );
  SDFFX1 DFF_116_Q_reg ( .D(g10726), .SI(g1015), .SE(n3433), .CLK(n3535), .Q(
        n1650) );
  SDFFX1 DFF_117_Q_reg ( .D(g4891), .SI(n1650), .SE(n3433), .CLK(n3535), .Q(
        n3059), .QN(n1874) );
  SDFFX1 DFF_118_Q_reg ( .D(g6224), .SI(n3059), .SE(n3428), .CLK(n3538), .Q(
        g1415), .QN(n3136) );
  SDFFX1 DFF_119_Q_reg ( .D(g7586), .SI(g1415), .SE(n3474), .CLK(n3515), .Q(
        g1227), .QN(n3129) );
  SDFFX1 DFF_120_Q_reg ( .D(g10770), .SI(g1227), .SE(n3474), .CLK(n3515), .Q(
        g1721) );
  SDFFX1 DFF_121_Q_reg ( .D(g2986), .SI(g1721), .SE(n3392), .CLK(n3556), .Q(
        n3058) );
  SDFFX1 DFF_122_Q_reg ( .D(n3381), .SI(n3058), .SE(n3392), .CLK(n3556), .Q(
        n3057) );
  SDFFX1 DFF_123_Q_reg ( .D(g6934), .SI(n3057), .SE(n3390), .CLK(n3557), .Q(
        g284) );
  SDFFX1 DFF_124_Q_reg ( .D(g11256), .SI(g284), .SE(n3470), .CLK(n3517), .Q(
        g426), .QN(n3294) );
  SDFFX1 DFF_125_Q_reg ( .D(g6824), .SI(g426), .SE(n3432), .CLK(n3536), .Q(
        g219), .QN(n3360) );
  SDFFX1 DFF_126_Q_reg ( .D(g1360), .SI(g219), .SE(n3413), .CLK(n3545), .Q(
        n3056) );
  SDFFX1 DFF_127_Q_reg ( .D(g6126), .SI(n3056), .SE(n3440), .CLK(n3532), .Q(
        g806), .QN(n3339) );
  SDFFX1 DFF_128_Q_reg ( .D(g8767), .SI(g806), .SE(n3402), .CLK(n3551), .Q(
        g1428), .QN(n3310) );
  SDFFX1 DFF_129_Q_reg ( .D(g102), .SI(g1428), .SE(n3402), .CLK(n3551), .Q(
        g2605) );
  SDFFX1 DFF_130_Q_reg ( .D(g6546), .SI(g2605), .SE(n3391), .CLK(n3556), .Q(
        g1564) );
  SDFFX1 DFF_131_Q_reg ( .D(g4238), .SI(g1564), .SE(n3391), .CLK(n3557), .Q(
        g1741) );
  SDFFX1 DFF_132_Q_reg ( .D(g6823), .SI(g1741), .SE(n3472), .CLK(n3516), .Q(
        g225), .QN(n3357) );
  SDFFX1 DFF_133_Q_reg ( .D(g6928), .SI(g225), .SE(n3391), .CLK(n3557), .Q(
        g281) );
  SDFFX1 DFF_134_Q_reg ( .D(g11602), .SI(g281), .SE(n3391), .CLK(n3557), .Q(
        g1308) );
  SDFFX1 DFF_135_Q_reg ( .D(g9721), .SI(g1308), .SE(n3471), .CLK(n3517), .Q(
        g611), .QN(n1609) );
  SDFFX1 DFF_136_Q_reg ( .D(g4890), .SI(g611), .SE(n3416), .CLK(n3544), .Q(
        n3055) );
  SDFFX1 DFF_137_Q_reg ( .D(n1586), .SI(n3055), .SE(n3416), .CLK(n3544), .Q(
        g1217) );
  SDFFX1 DFF_138_Q_reg ( .D(g6524), .SI(g1217), .SE(n3401), .CLK(n3551), .Q(
        g1589) );
  SDFFX1 DFF_139_Q_reg ( .D(g8045), .SI(g1589), .SE(n3450), .CLK(n3527), .Q(
        g1466), .QN(n3248) );
  SDFFX1 DFF_140_Q_reg ( .D(g6469), .SI(g1466), .SE(n3418), .CLK(n3543), .Q(
        g1571) );
  SDFFX1 DFF_141_Q_reg ( .D(g6471), .SI(g1571), .SE(n3424), .CLK(n3540), .Q(
        g1861), .QN(n3318) );
  SDFFX1 DFF_142_Q_reg ( .D(g6821), .SI(g1861), .SE(n3423), .CLK(n3540), .Q(
        n3054), .QN(n5999) );
  SDFFX1 DFF_143_Q_reg ( .D(g11514), .SI(n3054), .SE(n3439), .CLK(n3533), .Q(
        g1448), .QN(n3250) );
  SDFFX1 DFF_145_Q_reg ( .D(g4480), .SI(g1448), .SE(n3438), .CLK(n3533), .Q(
        g1133), .QN(n1706) );
  SDFFX1 DFF_146_Q_reg ( .D(g11610), .SI(g1133), .SE(n3464), .CLK(n3520), .Q(
        g1333) );
  SDFFX1 DFF_147_Q_reg ( .D(g7843), .SI(g1333), .SE(n3464), .CLK(n3520), .Q(
        g153), .QN(n3268) );
  SDFFX1 DFF_148_Q_reg ( .D(g11310), .SI(g153), .SE(n3444), .CLK(n3530), .Q(
        g962) );
  SDFFX1 DFF_149_Q_reg ( .D(g5536), .SI(g962), .SE(n3444), .CLK(n3530), .Q(
        g4175) );
  SDFFX1 DFF_150_Q_reg ( .D(g28), .SI(g4175), .SE(n3443), .CLK(n3530), .Q(
        g2603) );
  SDFFX1 DFF_151_Q_reg ( .D(g11331), .SI(g2603), .SE(n3443), .CLK(n3530), .Q(
        g486), .QN(n1621) );
  SDFFX1 DFF_152_Q_reg ( .D(g11380), .SI(g486), .SE(n3436), .CLK(n3534), .Q(
        g471), .QN(n1606) );
  SDFFX1 DFF_153_Q_reg ( .D(g6838), .SI(g471), .SE(n3431), .CLK(n3536), .Q(
        g1397) );
  SDFFX1 DFF_154_Q_reg ( .D(g103), .SI(g1397), .SE(n3431), .CLK(n3536), .Q(
        g2606) );
  SDFFX1 DFF_155_Q_reg ( .D(g8288), .SI(g2606), .SE(n3452), .CLK(n3526), .Q(
        g1950) );
  SDFFX1 DFF_156_Q_reg ( .D(g755), .SI(g1950), .SE(n3429), .CLK(n3538), .Q(
        g756) );
  SDFFX1 DFF_157_Q_reg ( .D(n256), .SI(g756), .SE(n3433), .CLK(n3536), .Q(
        n3053) );
  SDFFX1 DFF_159_Q_reg ( .D(g10855), .SI(g1101), .SE(n3413), .CLK(n3546), .Q(
        g549) );
  SDFFX1 DFF_161_Q_reg ( .D(g10898), .SI(g549), .SE(n3472), .CLK(n3516), .Q(
        g105), .QN(n3373) );
  SDFFX1 DFF_162_Q_reg ( .D(g10865), .SI(g105), .SE(n3472), .CLK(n3516), .Q(
        g1669) );
  SDFFX1 DFF_163_Q_reg ( .D(g6822), .SI(g1669), .SE(n3472), .CLK(n3516), .Q(
        test_so3) );
  SDFFX1 DFF_164_Q_reg ( .D(g6528), .SI(test_si4), .SE(n3418), .CLK(n3543), 
        .Q(g1531) );
  SDFFX1 DFF_165_Q_reg ( .D(g6180), .SI(g1531), .SE(n3450), .CLK(n3527), .Q(
        g1458), .QN(n1703) );
  SDFFX1 DFF_166_Q_reg ( .D(g10718), .SI(g1458), .SE(n3419), .CLK(n3542), .Q(
        g572) );
  SDFFX1 DFF_167_Q_reg ( .D(g6912), .SI(g572), .SE(n3436), .CLK(n3534), .Q(
        g1011), .QN(n3255) );
  SDFFX1 DFF_168_Q_reg ( .D(g10719), .SI(g1011), .SE(n3435), .CLK(n3534), .Q(
        n3051) );
  SDFFX1 DFF_169_Q_reg ( .D(g6234), .SI(n3051), .SE(n3435), .CLK(n3534), .Q(
        g1411) );
  SDFFX1 DFF_170_Q_reg ( .D(g6099), .SI(g1411), .SE(n3434), .CLK(n3535), .Q(
        g1074) );
  SDFFX1 DFF_171_Q_reg ( .D(g11259), .SI(g1074), .SE(n3454), .CLK(n3525), .Q(
        g444) );
  SDFFX1 DFF_172_Q_reg ( .D(g8039), .SI(g444), .SE(n3472), .CLK(n3516), .Q(
        g1474), .QN(n3281) );
  SDFFX1 DFF_173_Q_reg ( .D(g6059), .SI(g1474), .SE(n3419), .CLK(n3542), .Q(
        g1080) );
  SDFFX1 DFF_174_Q_reg ( .D(g5396), .SI(g1080), .SE(n3415), .CLK(n3545), .Q(
        g1713), .QN(n1610) );
  SDFFX1 DFF_175_Q_reg ( .D(g262), .SI(g1713), .SE(n3415), .CLK(n3545), .Q(
        g333), .QN(n3278) );
  SDFFX1 DFF_176_Q_reg ( .D(g6906), .SI(g333), .SE(n3400), .CLK(n3552), .Q(
        g269) );
  SDFFX1 DFF_177_Q_reg ( .D(g11266), .SI(g269), .SE(n3455), .CLK(n3524), .Q(
        g401), .QN(n3262) );
  SDFFX1 DFF_178_Q_reg ( .D(g11294), .SI(g401), .SE(n3474), .CLK(n3515), .Q(
        g1857), .QN(n1682) );
  SDFFX1 DFF_179_Q_reg ( .D(g5421), .SI(g1857), .SE(n3473), .CLK(n3515), .Q(g9) );
  SDFFX1 DFF_180_Q_reg ( .D(g8649), .SI(g9), .SE(n3468), .CLK(n3518), .Q(g664), 
        .QN(n3336) );
  SDFFX1 DFF_181_Q_reg ( .D(g11312), .SI(g664), .SE(n3421), .CLK(n3542), .Q(
        g965) );
  SDFFX1 DFF_182_Q_reg ( .D(g6840), .SI(g965), .SE(n3431), .CLK(n3537), .Q(
        g1400) );
  SDFFX1 DFF_183_Q_reg ( .D(g254), .SI(g1400), .SE(n3410), .CLK(n3547), .Q(
        g309), .QN(n3085) );
  SDFFX1 DFF_184_Q_reg ( .D(g7202), .SI(g309), .SE(n3439), .CLK(n3532), .Q(
        g814), .QN(n3338) );
  SDFFX1 DFF_185_Q_reg ( .D(g6834), .SI(g814), .SE(n3423), .CLK(n3540), .Q(
        g231), .QN(n3359) );
  SDFFX1 DFF_186_Q_reg ( .D(g10795), .SI(g231), .SE(n3437), .CLK(n3533), .Q(
        g557) );
  SDFFX1 DFF_187_Q_reg ( .D(g103), .SI(g557), .SE(n3437), .CLK(n3534), .Q(
        g2612) );
  SDFFX1 DFF_188_Q_reg ( .D(g875), .SI(g2612), .SE(n3404), .CLK(n3550), .Q(
        g869) );
  SDFFX1 DFF_189_Q_reg ( .D(g6831), .SI(g869), .SE(n3404), .CLK(n3550), .Q(
        g1383) );
  SDFFX1 DFF_190_Q_reg ( .D(g8060), .SI(g1383), .SE(n3456), .CLK(n3524), .Q(
        g158), .QN(n3247) );
  SDFFX1 DFF_191_Q_reg ( .D(g4893), .SI(g158), .SE(n3433), .CLK(n3536), .Q(
        g627), .QN(n1701) );
  SDFFX1 DFF_192_Q_reg ( .D(g7244), .SI(g627), .SE(n3441), .CLK(n3531), .Q(
        g1023), .QN(n3200) );
  SDFFX1 DFF_193_Q_reg ( .D(g6026), .SI(g1023), .SE(n3441), .CLK(n3531), .Q(
        g259) );
  SDFFX1 DFF_194_Q_reg ( .D(g3069), .SI(g259), .SE(n3441), .CLK(n3532), .Q(
        n3050) );
  SDFFX1 DFF_195_Q_reg ( .D(g11608), .SI(n3050), .SE(n3406), .CLK(n3549), .Q(
        g1327) );
  SDFFX1 DFF_196_Q_reg ( .D(g7660), .SI(g1327), .SE(n3459), .CLK(n3522), .Q(
        g654), .QN(n3315) );
  SDFFX1 DFF_197_Q_reg ( .D(g6911), .SI(g654), .SE(n3411), .CLK(n3546), .Q(
        g293) );
  SDFFX1 DFF_198_Q_reg ( .D(g11640), .SI(g293), .SE(n3408), .CLK(n3548), .Q(
        g1346) );
  SDFFX1 DFF_199_Q_reg ( .D(g8777), .SI(g1346), .SE(n3400), .CLK(n3552), .Q(
        g1633) );
  SDFFX1 DFF_200_Q_reg ( .D(g4274), .SI(g1633), .SE(n3396), .CLK(n3554), .Q(
        g1753) );
  SDFFX1 DFF_201_Q_reg ( .D(n3378), .SI(g1753), .SE(n3396), .CLK(n3554), .Q(
        g1508), .QN(n1707) );
  SDFFX1 DFF_202_Q_reg ( .D(g7297), .SI(g1508), .SE(n3462), .CLK(n3521), .Q(
        g1240), .QN(n3292) );
  SDFFX1 DFF_203_Q_reg ( .D(g11326), .SI(g1240), .SE(n3410), .CLK(n3547), .Q(
        g538), .QN(n3285) );
  SDFFX1 DFF_204_Q_reg ( .D(g11269), .SI(g538), .SE(n3455), .CLK(n3525), .Q(
        g416), .QN(n3236) );
  SDFFX1 DFF_205_Q_reg ( .D(g11325), .SI(g416), .SE(n3411), .CLK(n3547), .Q(
        g542), .QN(n3286) );
  SDFFX1 DFF_206_Q_reg ( .D(g10864), .SI(g542), .SE(n3411), .CLK(n3547), .Q(
        g1681) );
  SDFFX1 DFF_207_Q_reg ( .D(g11290), .SI(g1681), .SE(n3395), .CLK(n3554), .Q(
        g374), .QN(n3219) );
  SDFFX1 DFF_208_Q_reg ( .D(g10798), .SI(g374), .SE(n3395), .CLK(n3554), .Q(
        g563) );
  SDFFX1 DFF_209_Q_reg ( .D(g8284), .SI(g563), .SE(n3453), .CLK(n3525), .Q(
        g1914), .QN(n3224) );
  SDFFX1 DFF_210_Q_reg ( .D(g11328), .SI(g1914), .SE(n3410), .CLK(n3547), .Q(
        g530), .QN(n3283) );
  SDFFX1 DFF_211_Q_reg ( .D(g10800), .SI(g530), .SE(n3410), .CLK(n3547), .Q(
        g575) );
  SDFFX1 DFF_212_Q_reg ( .D(g8944), .SI(g575), .SE(n3451), .CLK(n3526), .Q(
        g1936), .QN(n1694) );
  SDFFX1 DFF_213_Q_reg ( .D(g7183), .SI(g1936), .SE(n3451), .CLK(n3527), .Q(
        g8978) );
  SDFFX1 DFF_214_Q_reg ( .D(g4465), .SI(g8978), .SE(n3451), .CLK(n3527), .Q(
        test_so4), .QN(n3387) );
  SDFFX1 DFF_215_Q_reg ( .D(g1356), .SI(test_si5), .SE(n3441), .CLK(n3532), 
        .Q(g1317), .QN(n3369) );
  SDFFX1 DFF_216_Q_reg ( .D(g11484), .SI(g1317), .SE(n3448), .CLK(n3528), .Q(
        g357) );
  SDFFX1 DFF_217_Q_reg ( .D(g11263), .SI(g357), .SE(n3448), .CLK(n3528), .Q(
        g386), .QN(n3260) );
  SDFFX1 DFF_218_Q_reg ( .D(g6501), .SI(g386), .SE(n3448), .CLK(n3528), .Q(
        g1601) );
  SDFFX1 DFF_220_Q_reg ( .D(g6757), .SI(g1601), .SE(n3448), .CLK(n3528), .Q(
        g166), .QN(n3245) );
  SDFFX1 DFF_221_Q_reg ( .D(g11334), .SI(g166), .SE(n3422), .CLK(n3541), .Q(
        g501), .QN(n1690) );
  SDFFX1 DFF_222_Q_reg ( .D(g6042), .SI(g501), .SE(n3430), .CLK(n3537), .Q(
        g262) );
  SDFFX1 DFF_223_Q_reg ( .D(g8384), .SI(g262), .SE(n3430), .CLK(n3537), .Q(
        g1840), .QN(n3288) );
  SDFFX1 DFF_224_Q_reg ( .D(g6653), .SI(g1840), .SE(n3426), .CLK(n3539), .Q(
        g8983) );
  SDFFX1 DFF_225_Q_reg ( .D(g257), .SI(g8983), .SE(n3426), .CLK(n3539), .Q(
        g318), .QN(n3259) );
  SDFFX1 DFF_226_Q_reg ( .D(g5763), .SI(g318), .SE(n3441), .CLK(n3532), .Q(
        g1356) );
  SDFFX1 DFF_227_Q_reg ( .D(g5849), .SI(g1356), .SE(n3440), .CLK(n3532), .Q(
        g794), .QN(n3346) );
  SDFFX1 DFF_228_Q_reg ( .D(g10722), .SI(g794), .SE(n3440), .CLK(n3532), .Q(
        n3048) );
  SDFFX1 DFF_229_Q_reg ( .D(g6929), .SI(n3048), .SE(n3411), .CLK(n3547), .Q(
        g302) );
  SDFFX1 DFF_230_Q_reg ( .D(g11488), .SI(g302), .SE(n3434), .CLK(n3535), .Q(
        g342) );
  SDFFX1 DFF_231_Q_reg ( .D(g7299), .SI(g342), .SE(n3462), .CLK(n3521), .Q(
        g1250), .QN(n3256) );
  SDFFX1 DFF_232_Q_reg ( .D(g4330), .SI(g1250), .SE(n3461), .CLK(n3521), .Q(
        g1163), .QN(n3265) );
  SDFFX1 DFF_233_Q_reg ( .D(g1958), .SI(g1163), .SE(n3398), .CLK(n3553), .Q(
        n3047), .QN(g5816) );
  SDFFX1 DFF_234_Q_reg ( .D(g7257), .SI(n3047), .SE(n3446), .CLK(n3529), .Q(
        g1032), .QN(n3368) );
  SDFFX1 DFF_235_Q_reg ( .D(g8775), .SI(g1032), .SE(n3445), .CLK(n3529), .Q(
        g1432), .QN(n3251) );
  SDFFX1 DFF_237_Q_reg ( .D(g5770), .SI(g1432), .SE(n3450), .CLK(n3527), .Q(
        g1453), .QN(n1628) );
  SDFFX1 DFF_238_Q_reg ( .D(g11486), .SI(g1453), .SE(n3458), .CLK(n3523), .Q(
        g363) );
  SDFFX1 DFF_239_Q_reg ( .D(g261), .SI(g363), .SE(n3458), .CLK(n3523), .Q(g330), .QN(n3084) );
  SDFFX1 DFF_240_Q_reg ( .D(g4338), .SI(g330), .SE(n3458), .CLK(n3523), .Q(
        g1157), .QN(n3263) );
  SDFFX1 DFF_241_Q_reg ( .D(g4500), .SI(g1157), .SE(n3458), .CLK(n3523), .Q(
        n3046), .QN(n6004) );
  SDFFX1 DFF_242_Q_reg ( .D(g10721), .SI(n3046), .SE(n3458), .CLK(n3523), .Q(
        n3045) );
  SDFFX1 DFF_243_Q_reg ( .D(g8147), .SI(n3045), .SE(n3442), .CLK(n3531), .Q(
        g928) );
  SDFFX1 DFF_244_Q_reg ( .D(g6038), .SI(g928), .SE(n3413), .CLK(n3546), .Q(
        g261) );
  SDFFX1 DFF_245_Q_reg ( .D(g11337), .SI(g261), .SE(n3412), .CLK(n3546), .Q(
        g516), .QN(n1620) );
  SDFFX1 DFF_246_Q_reg ( .D(g6045), .SI(g516), .SE(n3410), .CLK(n3547), .Q(
        g254) );
  SDFFX1 DFF_247_Q_reg ( .D(g7191), .SI(g254), .SE(n3394), .CLK(n3555), .Q(
        g4178), .QN(n3349) );
  SDFFX1 DFF_248_Q_reg ( .D(g826), .SI(g4178), .SE(n3425), .CLK(n3540), .Q(
        g861) );
  SDFFX1 DFF_249_Q_reg ( .D(g8774), .SI(g861), .SE(n3400), .CLK(n3552), .Q(
        g1627) );
  SDFFX1 DFF_250_Q_reg ( .D(g7293), .SI(g1627), .SE(n3460), .CLK(n3522), .Q(
        g1292), .QN(n3232) );
  SDFFX1 DFF_251_Q_reg ( .D(g6907), .SI(g1292), .SE(n3412), .CLK(n3546), .Q(
        g290) );
  SDFFX1 DFF_252_Q_reg ( .D(g4903), .SI(g290), .SE(n3412), .CLK(n3546), .Q(
        n3044), .QN(n1873) );
  SDFFX1 DFF_253_Q_reg ( .D(g6123), .SI(n3044), .SE(n3394), .CLK(n3555), .Q(
        g4176), .QN(n3350) );
  SDFFX1 DFF_254_Q_reg ( .D(g6506), .SI(g4176), .SE(n3434), .CLK(n3535), .Q(
        g1583) );
  SDFFX1 DFF_255_Q_reg ( .D(g11376), .SI(g1583), .SE(n3434), .CLK(n3535), .Q(
        g466), .QN(n1646) );
  SDFFX1 DFF_256_Q_reg ( .D(g6542), .SI(g466), .SE(n3402), .CLK(n3551), .Q(
        g1561) );
  SDFFX1 DFF_258_Q_reg ( .D(g6551), .SI(g1561), .SE(n3471), .CLK(n3516), .Q(
        g1546) );
  SDFFX1 DFF_259_Q_reg ( .D(g6901), .SI(g1546), .SE(n3447), .CLK(n3529), .Q(
        g287) );
  SDFFX1 DFF_260_Q_reg ( .D(g10797), .SI(g287), .SE(n3446), .CLK(n3529), .Q(
        g560) );
  SDFFX1 DFF_261_Q_reg ( .D(g8505), .SI(g560), .SE(n3417), .CLK(n3544), .Q(
        g617), .QN(n1645) );
  SDFFX1 DFF_262_Q_reg ( .D(n3379), .SI(g617), .SE(n3416), .CLK(n3544), .Q(
        n1631) );
  SDFFX1 DFF_263_Q_reg ( .D(g11647), .SI(n1631), .SE(n3463), .CLK(n3521), .Q(
        g336) );
  SDFFX1 DFF_264_Q_reg ( .D(g11340), .SI(g336), .SE(n3436), .CLK(n3534), .Q(
        g456), .QN(n1641) );
  SDFFX1 DFF_265_Q_reg ( .D(g253), .SI(g456), .SE(n3405), .CLK(n3550), .Q(g305), .QN(n1681) );
  SDFFX1 DFF_266_Q_reg ( .D(g11625), .SI(g305), .SE(n3446), .CLK(n3529), .Q(
        g345) );
  SDFFX1 DFF_267_Q_reg ( .D(g636), .SI(g345), .SE(n3470), .CLK(n3517), .Q(g8)
         );
  SDFFX1 DFF_268_Q_reg ( .D(g6502), .SI(g8), .SE(n3414), .CLK(n3545), .Q(
        test_so5), .QN(n3383) );
  SDFFX1 DFF_269_Q_reg ( .D(N599), .SI(test_si6), .SE(n3394), .CLK(n3555), .Q(
        g2648) );
  SDFFX1 DFF_270_Q_reg ( .D(g6049), .SI(g2648), .SE(n3393), .CLK(n3555), .Q(
        g255), .QN(n3334) );
  SDFFX1 DFF_271_Q_reg ( .D(g8945), .SI(g255), .SE(n3452), .CLK(n3526), .Q(
        g1945), .QN(n1697) );
  SDFFX1 DFF_272_Q_reg ( .D(g4231), .SI(g1945), .SE(n3397), .CLK(n3553), .Q(
        g1738) );
  SDFFX1 DFF_273_Q_reg ( .D(g8040), .SI(g1738), .SE(n3471), .CLK(n3516), .Q(
        g1478), .QN(n3314) );
  SDFFX1 DFF_275_Q_reg ( .D(n652), .SI(g1478), .SE(n3471), .CLK(n3516), .Q(
        n3042) );
  SDFFX1 DFF_276_Q_reg ( .D(g6155), .SI(n3042), .SE(n3431), .CLK(n3537), .Q(
        g1690), .QN(n1653) );
  SDFFX1 DFF_277_Q_reg ( .D(g8043), .SI(g1690), .SE(n3401), .CLK(n3552), .Q(
        g1482), .QN(n3249) );
  SDFFX1 DFF_278_Q_reg ( .D(g5173), .SI(g1482), .SE(n3401), .CLK(n3552), .Q(
        g1110), .QN(n1677) );
  SDFFX1 DFF_279_Q_reg ( .D(g6916), .SI(g1110), .SE(n3401), .CLK(n3552), .Q(
        g296) );
  SDFFX1 DFF_280_Q_reg ( .D(g10861), .SI(g296), .SE(n3469), .CLK(n3518), .Q(
        g1663) );
  SDFFX1 DFF_281_Q_reg ( .D(g8431), .SI(g1663), .SE(n3469), .CLK(n3518), .Q(
        g700), .QN(n3273) );
  SDFFX1 DFF_282_Q_reg ( .D(g4309), .SI(g700), .SE(n3396), .CLK(n3554), .Q(
        g1762) );
  SDFFX1 DFF_283_Q_reg ( .D(g11485), .SI(g1762), .SE(n3436), .CLK(n3534), .Q(
        g360) );
  SDFFX1 DFF_284_Q_reg ( .D(g6334), .SI(g360), .SE(n3432), .CLK(n3536), .Q(
        g192) );
  SDFFX1 DFF_285_Q_reg ( .D(g10767), .SI(g192), .SE(n3471), .CLK(n3517), .Q(
        g1657) );
  SDFFX1 DFF_286_Q_reg ( .D(g8923), .SI(g1657), .SE(n3471), .CLK(n3517), .Q(
        g722), .QN(n1693) );
  SDFFX1 DFF_287_Q_reg ( .D(g7189), .SI(g722), .SE(n3426), .CLK(n3539), .Q(
        g8980) );
  SDFFX1 DFF_288_Q_reg ( .D(g10799), .SI(g8980), .SE(n3457), .CLK(n3523), .Q(
        g566) );
  SDFFX1 DFF_289_Q_reg ( .D(g6747), .SI(g566), .SE(n3473), .CLK(n3516), .Q(
        n3041) );
  SDFFX1 DFF_290_Q_reg ( .D(g6080), .SI(n3041), .SE(n3473), .CLK(n3516), .Q(
        g1089) );
  SDFFX1 DFF_291_Q_reg ( .D(g3381), .SI(g1089), .SE(n3442), .CLK(n3531), .Q(
        g2986), .QN(n3107) );
  SDFFX1 DFF_292_Q_reg ( .D(g5910), .SI(g2986), .SE(n3441), .CLK(n3531), .Q(
        g1071) );
  SDFFX1 DFF_293_Q_reg ( .D(g11393), .SI(g1071), .SE(n3470), .CLK(n3517), .Q(
        g986), .QN(n1722) );
  SDFFX1 DFF_294_Q_reg ( .D(g11349), .SI(g986), .SE(n3470), .CLK(n3517), .Q(
        g971), .QN(n3371) );
  SDFFX1 DFF_295_Q_reg ( .D(g83), .SI(g971), .SE(n3469), .CLK(n3517), .Q(g1955) );
  SDFFX1 DFF_296_Q_reg ( .D(g6439), .SI(g1955), .SE(n3464), .CLK(n3520), .Q(
        g143), .QN(n3269) );
  SDFFX1 DFF_297_Q_reg ( .D(g9266), .SI(g143), .SE(n3429), .CLK(n3537), .Q(
        g1814), .QN(n1608) );
  SDFFX1 DFF_299_Q_reg ( .D(g1217), .SI(g1814), .SE(n3416), .CLK(n3544), .Q(
        g1212), .QN(n3362) );
  SDFFX1 DFF_300_Q_reg ( .D(g8940), .SI(g1212), .SE(n3430), .CLK(n3537), .Q(
        g1918), .QN(n3274) );
  SDFFX1 DFF_301_Q_reg ( .D(g7705), .SI(g1918), .SE(n3430), .CLK(n3537), .Q(
        g4179) );
  SDFFX1 DFF_302_Q_reg ( .D(g9269), .SI(g4179), .SE(n3429), .CLK(n3537), .Q(
        g1822), .QN(n1643) );
  SDFFX1 DFF_303_Q_reg ( .D(g6820), .SI(g1822), .SE(n3444), .CLK(n3530), .Q(
        g237) );
  SDFFX1 DFF_304_Q_reg ( .D(g756), .SI(g237), .SE(n3428), .CLK(n3538), .Q(g746), .QN(n3317) );
  SDFFX1 DFF_306_Q_reg ( .D(g8042), .SI(g746), .SE(n3450), .CLK(n3527), .Q(
        g1462), .QN(n3313) );
  SDFFX1 DFF_307_Q_reg ( .D(g6759), .SI(g1462), .SE(n3422), .CLK(n3541), .Q(
        g178) );
  SDFFX1 DFF_308_Q_reg ( .D(g11487), .SI(g178), .SE(n3445), .CLK(n3530), .Q(
        g366) );
  SDFFX1 DFF_309_Q_reg ( .D(g802), .SI(g366), .SE(n3440), .CLK(n3532), .Q(g837) );
  SDFFX1 DFF_310_Q_reg ( .D(g9124), .SI(g837), .SE(n3416), .CLK(n3544), .Q(
        g599), .QN(n1644) );
  SDFFX1 DFF_311_Q_reg ( .D(g11293), .SI(g599), .SE(n3474), .CLK(n3515), .Q(
        g1854) );
  SDFFX1 DFF_312_Q_reg ( .D(g11298), .SI(g1854), .SE(n3474), .CLK(n3515), .Q(
        g944) );
  SDFFX1 DFF_313_Q_reg ( .D(g8287), .SI(g944), .SE(n3453), .CLK(n3526), .Q(
        g1941), .QN(n3226) );
  SDFFX1 DFF_314_Q_reg ( .D(g8047), .SI(g1941), .SE(n3457), .CLK(n3524), .Q(
        g170), .QN(n3322) );
  SDFFX1 DFF_315_Q_reg ( .D(g6205), .SI(g170), .SE(n3428), .CLK(n3538), .Q(
        g1520), .QN(n1710) );
  SDFFX1 DFF_316_Q_reg ( .D(g8885), .SI(g1520), .SE(n3467), .CLK(n3518), .Q(
        g686), .QN(n1676) );
  SDFFX1 DFF_317_Q_reg ( .D(g11305), .SI(g686), .SE(n3398), .CLK(n3553), .Q(
        g953) );
  SDFFX1 DFF_318_Q_reg ( .D(g5556), .SI(g953), .SE(n3398), .CLK(n3553), .Q(
        g1958) );
  SDFFX1 DFF_319_Q_reg ( .D(g10664), .SI(g1958), .SE(n3398), .CLK(n3553), .Q(
        n3040) );
  SDFFX1 DFF_320_Q_reg ( .D(g2478), .SI(n3040), .SE(n3398), .CLK(n3553), .Q(
        g1765), .QN(n3366) );
  SDFFX1 DFF_321_Q_reg ( .D(g10711), .SI(g1765), .SE(n3397), .CLK(n3553), .Q(
        g1733) );
  SDFFX1 DFF_322_Q_reg ( .D(g7303), .SI(g1733), .SE(n3461), .CLK(n3522), .Q(
        test_so6), .QN(n3384) );
  SDFFX1 DFF_323_Q_reg ( .D(g5194), .SI(test_si7), .SE(n3420), .CLK(n3542), 
        .Q(g1610), .QN(n3365) );
  SDFFX1 DFF_324_Q_reg ( .D(g7541), .SI(g1610), .SE(n3406), .CLK(n3549), .Q(
        g1796), .QN(n1626) );
  SDFFX1 DFF_325_Q_reg ( .D(g11607), .SI(g1796), .SE(n3406), .CLK(n3549), .Q(
        g1324) );
  SDFFX1 DFF_326_Q_reg ( .D(g6541), .SI(g1324), .SE(n3407), .CLK(n3548), .Q(
        g1540) );
  SDFFX1 DFF_327_Q_reg ( .D(g6827), .SI(g1540), .SE(n3407), .CLK(n3548), .Q(
        n3038) );
  SDFFX1 DFF_328_Q_reg ( .D(n3380), .SI(n3038), .SE(n3392), .CLK(n3556), .Q(
        g3069), .QN(n3108) );
  SDFFX1 DFF_329_Q_reg ( .D(g11332), .SI(g3069), .SE(n3443), .CLK(n3530), .Q(
        g491), .QN(n1691) );
  SDFFX1 DFF_330_Q_reg ( .D(g4902), .SI(g491), .SE(n3424), .CLK(n3540), .Q(
        n3037) );
  SDFFX1 DFF_331_Q_reg ( .D(g6828), .SI(n3037), .SE(n3407), .CLK(n3548), .Q(
        g213) );
  SDFFX1 DFF_332_Q_reg ( .D(g6516), .SI(g213), .SE(n3407), .CLK(n3549), .Q(
        g1781), .QN(n1659) );
  SDFFX1 DFF_333_Q_reg ( .D(g8938), .SI(g1781), .SE(n3407), .CLK(n3549), .Q(
        g1900), .QN(n1675) );
  SDFFX1 DFF_334_Q_reg ( .D(g7298), .SI(g1900), .SE(n3462), .CLK(n3521), .Q(
        g1245), .QN(n3253) );
  SDFFX1 DFF_335_Q_reg ( .D(n6), .SI(g1245), .SE(n3462), .CLK(n3521), .Q(n3036), .QN(n6003) );
  SDFFX1 DFF_336_Q_reg ( .D(g6672), .SI(n3036), .SE(n3416), .CLK(n3544), .Q(
        n3035) );
  SDFFX1 DFF_337_Q_reg ( .D(g8048), .SI(n3035), .SE(n3422), .CLK(n3541), .Q(
        g148), .QN(n3270) );
  SDFFX1 DFF_338_Q_reg ( .D(g798), .SI(g148), .SE(n3400), .CLK(n3552), .Q(g833) );
  SDFFX1 DFF_339_Q_reg ( .D(g8285), .SI(g833), .SE(n3453), .CLK(n3526), .Q(
        g1923), .QN(n1718) );
  SDFFX1 DFF_340_Q_reg ( .D(g8254), .SI(g1923), .SE(n3442), .CLK(n3531), .Q(
        g936) );
  SDFFX1 DFF_342_Q_reg ( .D(g11604), .SI(g936), .SE(n3409), .CLK(n3548), .Q(
        g1314) );
  SDFFX1 DFF_343_Q_reg ( .D(g814), .SI(g1314), .SE(n3439), .CLK(n3532), .Q(
        g849) );
  SDFFX1 DFF_344_Q_reg ( .D(g11636), .SI(g849), .SE(n3439), .CLK(n3532), .Q(
        g1336), .QN(n3300) );
  SDFFX1 DFF_345_Q_reg ( .D(g6910), .SI(g1336), .SE(n3411), .CLK(n3546), .Q(
        g272) );
  SDFFX1 DFF_346_Q_reg ( .D(g8173), .SI(g272), .SE(n3403), .CLK(n3550), .Q(
        g1806), .QN(n3320) );
  SDFFX1 DFF_347_Q_reg ( .D(g8245), .SI(g1806), .SE(n3425), .CLK(n3540), .Q(
        g826), .QN(n1716) );
  SDFFX1 DFF_349_Q_reg ( .D(g8281), .SI(g826), .SE(n3452), .CLK(n3526), .Q(
        g1887), .QN(n3194) );
  SDFFX1 DFF_350_Q_reg ( .D(g10724), .SI(g1887), .SE(n3452), .CLK(n3526), .Q(
        n3034) );
  SDFFX1 DFF_351_Q_reg ( .D(g11314), .SI(n3034), .SE(n3424), .CLK(n3540), .Q(
        g968) );
  SDFFX1 DFF_352_Q_reg ( .D(g4905), .SI(g968), .SE(n3424), .CLK(n3540), .Q(
        n3033), .QN(n5998) );
  SDFFX1 DFF_353_Q_reg ( .D(g4484), .SI(n3033), .SE(n3424), .CLK(n3540), .Q(
        g1137), .QN(n1597) );
  SDFFX1 DFF_354_Q_reg ( .D(g8937), .SI(g1137), .SE(n3451), .CLK(n3526), .Q(
        g1891), .QN(n1657) );
  SDFFX1 DFF_355_Q_reg ( .D(g7300), .SI(g1891), .SE(n3461), .CLK(n3521), .Q(
        g1255), .QN(n3228) );
  SDFFX1 DFF_356_Q_reg ( .D(g6002), .SI(g1255), .SE(n3437), .CLK(n3534), .Q(
        g257) );
  SDFFX1 DFF_357_Q_reg ( .D(n1588), .SI(g257), .SE(n3437), .CLK(n3534), .Q(
        g874) );
  SDFFX1 DFF_358_Q_reg ( .D(g9110), .SI(g874), .SE(n3417), .CLK(n3544), .Q(
        g591), .QN(n1607) );
  SDFFX1 DFF_359_Q_reg ( .D(g8926), .SI(g591), .SE(n3390), .CLK(n3557), .Q(
        g731), .QN(n1696) );
  SDFFX1 DFF_360_Q_reg ( .D(g8631), .SI(g731), .SE(n3470), .CLK(n3517), .Q(
        g636) );
  SDFFX1 DFF_361_Q_reg ( .D(g7632), .SI(g636), .SE(n3475), .CLK(n3515), .Q(
        g1218), .QN(n3367) );
  SDFFX1 DFF_362_Q_reg ( .D(g9150), .SI(g1218), .SE(n3417), .CLK(n3543), .Q(
        g605), .QN(n1593) );
  SDFFX1 DFF_363_Q_reg ( .D(g6531), .SI(g605), .SE(n3417), .CLK(n3544), .Q(
        g8986) );
  SDFFX1 DFF_364_Q_reg ( .D(g6786), .SI(g8986), .SE(n3421), .CLK(n3541), .Q(
        g182), .QN(n3267) );
  SDFFX1 DFF_365_Q_reg ( .D(g11303), .SI(g182), .SE(n3421), .CLK(n3541), .Q(
        g950) );
  SDFFX1 DFF_366_Q_reg ( .D(g4477), .SI(g950), .SE(n3421), .CLK(n3541), .Q(
        g1129), .QN(n1705) );
  SDFFX1 DFF_367_Q_reg ( .D(g822), .SI(g1129), .SE(n3421), .CLK(n3542), .Q(
        g857) );
  SDFFX1 DFF_368_Q_reg ( .D(g11258), .SI(g857), .SE(n3454), .CLK(n3525), .Q(
        g448) );
  SDFFX1 DFF_369_Q_reg ( .D(g9272), .SI(g448), .SE(n3429), .CLK(n3537), .Q(
        g1828), .QN(n1605) );
  SDFFX1 DFF_370_Q_reg ( .D(g10773), .SI(g1828), .SE(n3402), .CLK(n3551), .Q(
        g1727) );
  SDFFX1 DFF_371_Q_reg ( .D(g6470), .SI(g1727), .SE(n3420), .CLK(n3542), .Q(
        g1592) );
  SDFFX1 DFF_372_Q_reg ( .D(g5083), .SI(g1592), .SE(n3420), .CLK(n3542), .Q(
        g1703), .QN(n3331) );
  SDFFX1 DFF_373_Q_reg ( .D(g8286), .SI(g1703), .SE(n3453), .CLK(n3526), .Q(
        g1932), .QN(n3227) );
  SDFFX1 DFF_374_Q_reg ( .D(g8773), .SI(g1932), .SE(n3401), .CLK(n3551), .Q(
        g1624) );
  SDFFX1 DFF_376_Q_reg ( .D(g6054), .SI(g1624), .SE(n3463), .CLK(n3521), .Q(
        test_so7) );
  SDFFX1 DFF_377_Q_reg ( .D(g101), .SI(test_si8), .SE(n3475), .CLK(n3515), .Q(
        g2601) );
  SDFFX1 DFF_378_Q_reg ( .D(g11260), .SI(g2601), .SE(n3454), .CLK(n3525), .Q(
        g440) );
  SDFFX1 DFF_379_Q_reg ( .D(g11338), .SI(g440), .SE(n3412), .CLK(n3546), .Q(
        g476), .QN(n1599) );
  SDFFX1 DFF_380_Q_reg ( .D(g5918), .SI(g476), .SE(n3412), .CLK(n3546), .Q(
        g119), .QN(n1613) );
  SDFFX1 DFF_381_Q_reg ( .D(g8922), .SI(g119), .SE(n3408), .CLK(n3548), .Q(
        g668), .QN(n1662) );
  SDFFX1 DFF_382_Q_reg ( .D(g8049), .SI(g668), .SE(n3448), .CLK(n3528), .Q(
        g139), .QN(n3242) );
  SDFFX1 DFF_383_Q_reg ( .D(g4342), .SI(g139), .SE(n3448), .CLK(n3528), .Q(
        g1149), .QN(n1685) );
  SDFFX1 DFF_384_Q_reg ( .D(g10720), .SI(g1149), .SE(n3447), .CLK(n3528), .Q(
        n3031) );
  SDFFX1 DFF_385_Q_reg ( .D(g6755), .SI(n3031), .SE(n3424), .CLK(n3540), .Q(
        n3030) );
  SDFFX1 DFF_386_Q_reg ( .D(g6897), .SI(n3030), .SE(n3400), .CLK(n3552), .Q(
        g263) );
  SDFFX1 DFF_387_Q_reg ( .D(g7709), .SI(g263), .SE(n3425), .CLK(n3539), .Q(
        g818), .QN(n3325) );
  SDFFX1 DFF_388_Q_reg ( .D(g4255), .SI(g818), .SE(n3394), .CLK(n3555), .Q(
        g1747) );
  SDFFX1 DFF_389_Q_reg ( .D(g5543), .SI(g1747), .SE(n3440), .CLK(n3532), .Q(
        g802), .QN(n1622) );
  SDFFX1 DFF_390_Q_reg ( .D(g6915), .SI(g802), .SE(n3456), .CLK(n3524), .Q(
        g275) );
  SDFFX1 DFF_391_Q_reg ( .D(g6513), .SI(g275), .SE(n3456), .CLK(n3524), .Q(
        g1524) );
  SDFFX1 DFF_392_Q_reg ( .D(g6480), .SI(g1524), .SE(n3456), .CLK(n3524), .Q(
        g1577) );
  SDFFX1 DFF_393_Q_reg ( .D(g6733), .SI(g1577), .SE(n3456), .CLK(n3524), .Q(
        g810), .QN(n3326) );
  SDFFX1 DFF_394_Q_reg ( .D(g11264), .SI(g810), .SE(n3455), .CLK(n3524), .Q(
        g391), .QN(n3296) );
  SDFFX1 DFF_395_Q_reg ( .D(g8973), .SI(g391), .SE(n3459), .CLK(n3523), .Q(
        g658), .QN(n1615) );
  SDFFX1 DFF_396_Q_reg ( .D(g6833), .SI(g658), .SE(n3405), .CLK(n3549), .Q(
        g1386), .QN(n3333) );
  SDFFX1 DFF_397_Q_reg ( .D(g5996), .SI(g1386), .SE(n3405), .CLK(n3550), .Q(
        g253) );
  SDFFX1 DFF_398_Q_reg ( .D(n1587), .SI(g253), .SE(n3405), .CLK(n3550), .Q(
        g875) );
  SDFFX1 DFF_399_Q_reg ( .D(g4473), .SI(g875), .SE(n3404), .CLK(n3550), .Q(
        g1125), .QN(n1708) );
  SDFFX1 DFF_400_Q_reg ( .D(g5755), .SI(g1125), .SE(n3404), .CLK(n3550), .Q(
        g201), .QN(n1619) );
  SDFFX1 DFF_401_Q_reg ( .D(g7295), .SI(g201), .SE(n3460), .CLK(n3522), .Q(
        g1280), .QN(n1862) );
  SDFFX1 DFF_402_Q_reg ( .D(g6068), .SI(g1280), .SE(n3459), .CLK(n3522), .Q(
        g1083) );
  SDFFX1 DFF_403_Q_reg ( .D(g7137), .SI(g1083), .SE(n3459), .CLK(n3522), .Q(
        g650), .QN(n1709) );
  SDFFX1 DFF_404_Q_reg ( .D(g8779), .SI(g650), .SE(n3444), .CLK(n3530), .Q(
        g1636) );
  SDFFX1 DFF_405_Q_reg ( .D(g818), .SI(g1636), .SE(n3444), .CLK(n3530), .Q(
        g853) );
  SDFFX1 DFF_406_Q_reg ( .D(g11270), .SI(g853), .SE(n3454), .CLK(n3525), .Q(
        g421), .QN(n3277) );
  SDFFX1 DFF_407_Q_reg ( .D(g5529), .SI(g421), .SE(n3399), .CLK(n3552), .Q(
        g4174), .QN(n3352) );
  SDFFX1 DFF_408_Q_reg ( .D(g11306), .SI(g4174), .SE(n3399), .CLK(n3552), .Q(
        g956) );
  SDFFX1 DFF_409_Q_reg ( .D(g11291), .SI(g956), .SE(n3399), .CLK(n3553), .Q(
        g378), .QN(n3218) );
  SDFFX1 DFF_410_Q_reg ( .D(g4283), .SI(g378), .SE(n3399), .CLK(n3553), .Q(
        g1756) );
  SDFFX1 DFF_411_Q_reg ( .D(g29), .SI(g1756), .SE(n3399), .CLK(n3553), .Q(
        g2604) );
  SDFFX1 DFF_412_Q_reg ( .D(g806), .SI(g2604), .SE(n3398), .CLK(n3553), .Q(
        g841) );
  SDFFX1 DFF_413_Q_reg ( .D(g6894), .SI(g841), .SE(n3463), .CLK(n3521), .Q(
        g1027), .QN(n3324) );
  SDFFX1 DFF_414_Q_reg ( .D(g6902), .SI(g1027), .SE(n3464), .CLK(n3520), .Q(
        g1003), .QN(n3293) );
  SDFFX1 DFF_415_Q_reg ( .D(g8765), .SI(g1003), .SE(n3421), .CLK(n3542), .Q(
        g1403), .QN(n3252) );
  SDFFX1 DFF_416_Q_reg ( .D(g4498), .SI(g1403), .SE(n3420), .CLK(n3542), .Q(
        g1145), .QN(n1617) );
  SDFFX1 DFF_417_Q_reg ( .D(g5148), .SI(g1145), .SE(n3413), .CLK(n3545), .Q(
        g1107), .QN(n1614) );
  SDFFX1 DFF_418_Q_reg ( .D(g7581), .SI(g1107), .SE(n3408), .CLK(n3548), .Q(
        g1223), .QN(n3130) );
  SDFFX1 DFF_419_Q_reg ( .D(g11267), .SI(g1223), .SE(n3455), .CLK(n3525), .Q(
        g406), .QN(n3230) );
  SDFFX1 DFF_420_Q_reg ( .D(g10936), .SI(g406), .SE(n3420), .CLK(n3542), .Q(
        g1811) );
  SDFFX1 DFF_421_Q_reg ( .D(g10784), .SI(g1811), .SE(n3420), .CLK(n3542), .Q(
        n3029) );
  SDFFX1 DFF_423_Q_reg ( .D(g10765), .SI(n3029), .SE(n3474), .CLK(n3515), .Q(
        g1654) );
  SDFFX1 DFF_424_Q_reg ( .D(g6332), .SI(g1654), .SE(n3473), .CLK(n3515), .Q(
        g197), .QN(n1678) );
  SDFFX1 DFF_425_Q_reg ( .D(g6479), .SI(g197), .SE(n3391), .CLK(n3556), .Q(
        g1595) );
  SDFFX1 DFF_426_Q_reg ( .D(g6537), .SI(g1595), .SE(n3465), .CLK(n3520), .Q(
        g1537) );
  SDFFX1 DFF_427_Q_reg ( .D(g8434), .SI(g1537), .SE(n3468), .CLK(n3518), .Q(
        g727), .QN(n3225) );
  SDFFX1 DFF_428_Q_reg ( .D(g6908), .SI(g727), .SE(n3473), .CLK(n3516), .Q(
        test_so8), .QN(n3386) );
  SDFFX1 DFF_429_Q_reg ( .D(g6243), .SI(test_si9), .SE(n3427), .CLK(n3538), 
        .Q(g798), .QN(n1717) );
  SDFFX1 DFF_430_Q_reg ( .D(g11324), .SI(g798), .SE(n3427), .CLK(n3538), .Q(
        g481), .QN(n1680) );
  SDFFX1 DFF_431_Q_reg ( .D(n438), .SI(g481), .SE(n3427), .CLK(n3538), .Q(
        g4172), .QN(n1647) );
  SDFFX1 DFF_432_Q_reg ( .D(g11609), .SI(g4172), .SE(n3404), .CLK(n3550), .Q(
        g1330) );
  SDFFX1 DFF_433_Q_reg ( .D(g810), .SI(g1330), .SE(n3404), .CLK(n3550), .Q(
        g845) );
  SDFFX1 DFF_434_Q_reg ( .D(g8244), .SI(g845), .SE(n3394), .CLK(n3555), .Q(
        g4181), .QN(n3345) );
  SDFFX1 DFF_435_Q_reg ( .D(g8194), .SI(g4181), .SE(n3394), .CLK(n3555), .Q(
        g1512) );
  SDFFX1 DFF_436_Q_reg ( .D(g113), .SI(g1512), .SE(n3443), .CLK(n3531), .Q(
        n3027) );
  SDFFX1 DFF_437_Q_reg ( .D(g8052), .SI(n3027), .SE(n3465), .CLK(n3519), .Q(
        g1490), .QN(n3312) );
  SDFFX1 DFF_438_Q_reg ( .D(g4325), .SI(g1490), .SE(n3465), .CLK(n3519), .Q(
        g1166), .QN(n3266) );
  SDFFX1 DFF_440_Q_reg ( .D(g11481), .SI(g1166), .SE(n3426), .CLK(n3539), .Q(
        g348) );
  SDFFX1 DFF_441_Q_reg ( .D(g874), .SI(g348), .SE(n3436), .CLK(n3534), .Q(
        n3026) );
  SDFFX1 DFF_442_Q_reg ( .D(g7301), .SI(n3026), .SE(n3461), .CLK(n3521), .Q(
        g1260), .QN(n3229) );
  SDFFX1 DFF_443_Q_reg ( .D(g6035), .SI(g1260), .SE(n3457), .CLK(n3524), .Q(
        g260) );
  SDFFX1 DFF_444_Q_reg ( .D(g8059), .SI(g260), .SE(n3447), .CLK(n3528), .Q(
        g131), .QN(n3241) );
  SDFFX1 DFF_445_Q_reg ( .D(g1854), .SI(g131), .SE(n3447), .CLK(n3529), .Q(
        n3025) );
  SDFFX1 DFF_446_Q_reg ( .D(g6015), .SI(n3025), .SE(n3446), .CLK(n3529), .Q(
        g258) );
  SDFFX1 DFF_447_Q_reg ( .D(g11330), .SI(g258), .SE(n3446), .CLK(n3529), .Q(
        g521), .QN(n1698) );
  SDFFX1 DFF_448_Q_reg ( .D(g11605), .SI(g521), .SE(n3403), .CLK(n3550), .Q(
        g1318) );
  SDFFX1 DFF_449_Q_reg ( .D(g8921), .SI(g1318), .SE(n3403), .CLK(n3550), .Q(
        g1872), .QN(n1616) );
  SDFFX1 DFF_450_Q_reg ( .D(g8883), .SI(g1872), .SE(n3403), .CLK(n3551), .Q(
        g677), .QN(n1656) );
  SDFFX1 DFF_451_Q_reg ( .D(g28), .SI(g677), .SE(n3403), .CLK(n3551), .Q(g2608) );
  SDFFX1 DFF_452_Q_reg ( .D(n60), .SI(g2608), .SE(n3403), .CLK(n3551), .Q(
        n3024) );
  SDFFX1 DFF_453_Q_reg ( .D(g6523), .SI(n3024), .SE(n3402), .CLK(n3551), .Q(
        g1549) );
  SDFFX1 DFF_454_Q_reg ( .D(g11300), .SI(g1549), .SE(n3400), .CLK(n3552), .Q(
        g947) );
  SDFFX1 DFF_455_Q_reg ( .D(g9555), .SI(g947), .SE(n3452), .CLK(n3526), .Q(
        g1834), .QN(n1655) );
  SDFFX1 DFF_456_Q_reg ( .D(g6481), .SI(g1834), .SE(n3438), .CLK(n3533), .Q(
        g1598) );
  SDFFX1 DFF_457_Q_reg ( .D(g4471), .SI(g1598), .SE(n3437), .CLK(n3533), .Q(
        g1121), .QN(n1618) );
  SDFFX1 DFF_458_Q_reg ( .D(g11606), .SI(g1121), .SE(n3406), .CLK(n3549), .Q(
        g1321) );
  SDFFX1 DFF_459_Q_reg ( .D(g11335), .SI(g1321), .SE(n3422), .CLK(n3541), .Q(
        g506), .QN(n1600) );
  SDFFX1 DFF_460_Q_reg ( .D(g10791), .SI(g506), .SE(n3422), .CLK(n3541), .Q(
        g546) );
  SDFFX1 DFF_461_Q_reg ( .D(g8939), .SI(g546), .SE(n3429), .CLK(n3538), .Q(
        g1909), .QN(n3330) );
  SDFFX1 DFF_462_Q_reg ( .D(g83), .SI(g1909), .SE(n3429), .CLK(n3538), .Q(g755) );
  SDFFX1 DFF_463_Q_reg ( .D(g6529), .SI(g755), .SE(n3449), .CLK(n3527), .Q(
        g1552) );
  SDFFX1 DFF_464_Q_reg ( .D(g101), .SI(g1552), .SE(n3449), .CLK(n3527), .Q(
        g2610) );
  SDFFX1 DFF_465_Q_reg ( .D(g10776), .SI(g2610), .SE(n3449), .CLK(n3527), .Q(
        g1687) );
  SDFFX1 DFF_466_Q_reg ( .D(g6514), .SI(g1687), .SE(n3449), .CLK(n3528), .Q(
        g1586) );
  SDFFX1 DFF_467_Q_reg ( .D(g259), .SI(g1586), .SE(n3449), .CLK(n3528), .Q(
        g324), .QN(n3257) );
  SDFFX1 DFF_468_Q_reg ( .D(g4490), .SI(g324), .SE(n3449), .CLK(n3528), .Q(
        g1141), .QN(n1660) );
  SDFFX1 DFF_470_Q_reg ( .D(g11639), .SI(g1141), .SE(n3415), .CLK(n3544), .Q(
        g1341), .QN(n3298) );
  SDFFX1 DFF_471_Q_reg ( .D(g4089), .SI(g1341), .SE(n3415), .CLK(n3544), .Q(
        g1710) );
  SDFFX1 DFF_472_Q_reg ( .D(g10785), .SI(g1710), .SE(n3415), .CLK(n3544), .Q(
        n3023) );
  SDFFX1 DFF_473_Q_reg ( .D(g6179), .SI(n3023), .SE(n3473), .CLK(n3515), .Q(
        n3022), .QN(n5997) );
  SDFFX1 DFF_474_Q_reg ( .D(g8053), .SI(n3022), .SE(n3447), .CLK(n3528), .Q(
        g135), .QN(n3243) );
  SDFFX1 DFF_475_Q_reg ( .D(g11329), .SI(g135), .SE(n3409), .CLK(n3547), .Q(
        g525), .QN(n1695) );
  SDFFX1 DFF_476_Q_reg ( .D(g104), .SI(g525), .SE(n3409), .CLK(n3547), .Q(
        g2607) );
  SDFFX1 DFF_477_Q_reg ( .D(g6515), .SI(g2607), .SE(n3409), .CLK(n3547), .Q(
        g1607) );
  SDFFX1 DFF_478_Q_reg ( .D(g258), .SI(g1607), .SE(n3409), .CLK(n3548), .Q(
        g321), .QN(n3297) );
  SDFFX1 DFF_479_Q_reg ( .D(g7204), .SI(g321), .SE(n3409), .CLK(n3548), .Q(
        g8982) );
  SDFFX1 DFF_480_Q_reg ( .D(g11443), .SI(g8982), .SE(n3462), .CLK(n3521), .Q(
        g1275), .QN(n3290) );
  SDFFX1 DFF_481_Q_reg ( .D(g11603), .SI(g1275), .SE(n3414), .CLK(n3545), .Q(
        test_so9) );
  SDFFX1 DFF_482_Q_reg ( .D(g8770), .SI(test_si10), .SE(n3437), .CLK(n3533), 
        .Q(g1615) );
  SDFFX1 DFF_483_Q_reg ( .D(g11292), .SI(g1615), .SE(n3396), .CLK(n3554), .Q(
        g382) );
  SDFFX1 DFF_484_Q_reg ( .D(g6331), .SI(g382), .SE(n3395), .CLK(n3554), .Q(
        n3020) );
  SDFFX1 DFF_485_Q_reg ( .D(g6900), .SI(n3020), .SE(n3395), .CLK(n3555), .Q(
        g266) );
  SDFFX1 DFF_486_Q_reg ( .D(g7294), .SI(g266), .SE(n3460), .CLK(n3522), .Q(
        g1284), .QN(n1864) );
  SDFFX1 DFF_487_Q_reg ( .D(g6829), .SI(g1284), .SE(n3407), .CLK(n3549), .Q(
        n3019) );
  SDFFX1 DFF_488_Q_reg ( .D(g8428), .SI(n3019), .SE(n3468), .CLK(n3518), .Q(
        g673), .QN(n3193) );
  SDFFX1 DFF_489_Q_reg ( .D(n386), .SI(g673), .SE(n3412), .CLK(n3546), .Q(
        n3018) );
  SDFFX1 DFF_490_Q_reg ( .D(g8054), .SI(n3018), .SE(n3456), .CLK(n3524), .Q(
        g162), .QN(n3246) );
  SDFFX1 DFF_491_Q_reg ( .D(g11268), .SI(g162), .SE(n3455), .CLK(n3525), .Q(
        g411), .QN(n3279) );
  SDFFX1 DFF_492_Q_reg ( .D(g11262), .SI(g411), .SE(n3453), .CLK(n3525), .Q(
        g431), .QN(n1876) );
  SDFFX1 DFF_493_Q_reg ( .D(g8283), .SI(g431), .SE(n3453), .CLK(n3525), .Q(
        g1905), .QN(n3342) );
  SDFFX1 DFF_494_Q_reg ( .D(g6193), .SI(g1905), .SE(n3428), .CLK(n3538), .Q(
        g1515), .QN(n1627) );
  SDFFX1 DFF_495_Q_reg ( .D(g8776), .SI(g1515), .SE(n3472), .CLK(n3516), .Q(
        g1630) );
  SDFFX1 DFF_496_Q_reg ( .D(g7143), .SI(g1630), .SE(n3426), .CLK(n3539), .Q(
        g8976) );
  SDFFX1 DFF_497_Q_reg ( .D(g6898), .SI(g8976), .SE(n3390), .CLK(n3557), .Q(
        g991), .QN(n1871) );
  SDFFX1 DFF_498_Q_reg ( .D(g7291), .SI(g991), .SE(n3460), .CLK(n3522), .Q(
        g1300), .QN(n3234) );
  SDFFX1 DFF_499_Q_reg ( .D(g11478), .SI(g1300), .SE(n3393), .CLK(n3556), .Q(
        g339) );
  SDFFX1 DFF_500_Q_reg ( .D(g6000), .SI(g339), .SE(n3463), .CLK(n3520), .Q(
        g256) );
  SDFFX1 DFF_501_Q_reg ( .D(g4264), .SI(g256), .SE(n3397), .CLK(n3554), .Q(
        g1750) );
  SDFFX1 DFF_502_Q_reg ( .D(g102), .SI(g1750), .SE(n3397), .CLK(n3554), .Q(
        g2611) );
  SDFFX1 DFF_503_Q_reg ( .D(g8768), .SI(g2611), .SE(n3438), .CLK(n3533), .Q(
        g1440), .QN(n3309) );
  SDFFX1 DFF_504_Q_reg ( .D(g10863), .SI(g1440), .SE(n3469), .CLK(n3517), .Q(
        g1666) );
  SDFFX1 DFF_505_Q_reg ( .D(g6522), .SI(g1666), .SE(n3469), .CLK(n3518), .Q(
        g1528) );
  SDFFX1 DFF_506_Q_reg ( .D(g11641), .SI(g1528), .SE(n3439), .CLK(n3533), .Q(
        g1351), .QN(n1721) );
  SDFFX1 DFF_507_Q_reg ( .D(g10780), .SI(g1351), .SE(n3439), .CLK(n3533), .Q(
        n3017) );
  SDFFX1 DFF_508_Q_reg ( .D(g8044), .SI(n3017), .SE(n3447), .CLK(n3529), .Q(
        g127), .QN(n1704) );
  SDFFX1 DFF_509_Q_reg ( .D(g11579), .SI(g127), .SE(n3467), .CLK(n3519), .Q(
        g1618) );
  SDFFX1 DFF_510_Q_reg ( .D(g7296), .SI(g1618), .SE(n3462), .CLK(n3521), .Q(
        g1235), .QN(n3254) );
  SDFFX1 DFF_511_Q_reg ( .D(g6923), .SI(g1235), .SE(n3411), .CLK(n3546), .Q(
        g299) );
  SDFFX1 DFF_512_Q_reg ( .D(g11261), .SI(g299), .SE(n3454), .CLK(n3525), .Q(
        g435), .QN(n1878) );
  SDFFX1 DFF_513_Q_reg ( .D(g6638), .SI(g435), .SE(n3426), .CLK(n3539), .Q(
        g8981) );
  SDFFX1 DFF_514_Q_reg ( .D(g6534), .SI(g8981), .SE(n3408), .CLK(n3548), .Q(
        g1555) );
  SDFFX1 DFF_515_Q_reg ( .D(g6895), .SI(g1555), .SE(n3408), .CLK(n3548), .Q(
        g995), .QN(n3291) );
  SDFFX1 DFF_516_Q_reg ( .D(g8771), .SI(g995), .SE(n3466), .CLK(n3519), .Q(
        g1621) );
  SDFFX1 DFF_517_Q_reg ( .D(g4506), .SI(g1621), .SE(n3466), .CLK(n3519), .Q(
        n3016), .QN(n6001) );
  SDFFX1 DFF_518_Q_reg ( .D(g7441), .SI(n3016), .SE(n3393), .CLK(n3556), .Q(
        g643), .QN(n1612) );
  SDFFX1 DFF_519_Q_reg ( .D(g8055), .SI(g643), .SE(n3450), .CLK(n3527), .Q(
        g1494), .QN(n3280) );
  SDFFX1 DFF_520_Q_reg ( .D(g6468), .SI(g1494), .SE(n3418), .CLK(n3543), .Q(
        g1567) );
  SDFFX1 DFF_521_Q_reg ( .D(g8430), .SI(g1567), .SE(n3467), .CLK(n3518), .Q(
        g691), .QN(n3341) );
  SDFFX1 DFF_522_Q_reg ( .D(g11327), .SI(g691), .SE(n3410), .CLK(n3547), .Q(
        g534), .QN(n3284) );
  SDFFX1 DFF_523_Q_reg ( .D(g6508), .SI(g534), .SE(n3414), .CLK(n3545), .Q(
        g1776), .QN(n1715) );
  SDFFX1 DFF_524_Q_reg ( .D(g10717), .SI(g1776), .SE(n3414), .CLK(n3545), .Q(
        g569) );
  SDFFX1 DFF_525_Q_reg ( .D(g4334), .SI(g569), .SE(n3414), .CLK(n3545), .Q(
        g1160), .QN(n3264) );
  SDFFX1 DFF_526_Q_reg ( .D(n1585), .SI(g1160), .SE(n3413), .CLK(n3545), .Q(
        g1360) );
  SDFFX1 DFF_528_Q_reg ( .D(g6679), .SI(g1360), .SE(n3445), .CLK(n3529), .Q(g1) );
  SDFFX1 DFF_529_Q_reg ( .D(g11336), .SI(g1), .SE(n3445), .CLK(n3529), .Q(g511), .QN(n1679) );
  SDFFX1 DFF_530_Q_reg ( .D(g10771), .SI(g511), .SE(n3419), .CLK(n3543), .Q(
        g1724) );
  SDFFX1 DFF_531_Q_reg ( .D(g5445), .SI(g1724), .SE(n3418), .CLK(n3543), .Q(
        g12) );
  SDFFX1 DFF_532_Q_reg ( .D(g8559), .SI(g12), .SE(n3452), .CLK(n3526), .Q(
        g1878), .QN(n3337) );
  SDFFX1 DFF_533_Q_reg ( .D(g7219), .SI(g1878), .SE(n3425), .CLK(n3539), .Q(
        test_so10) );
  SDFFX1 DFF_158_Q_reg ( .D(g5390), .SI(n3053), .SE(n3413), .CLK(n3546), .Q(
        g1101), .QN(n1654) );
  AND2X2 Tg1_Trojan1 ( .IN1(g6179), .IN2(n60), .Q(Tg1_OUT1) );
  AND2X2 Tg1_Trojan2 ( .IN1(n59), .IN2(n233), .Q(Tg1_OUT2) );
  AND2X2 Tg1_Trojan3 ( .IN1(n1226), .IN2(n72), .Q(Tg1_OUT3) );
  AND2X2 Tg1_Trojan4 ( .IN1(g5556), .IN2(n898), .Q(Tg1_OUT4) );
  AND4X1 Tg1_Trojan1234 ( .IN1(Tg1_OUT1), .IN2(Tg1_OUT2), .IN3(Tg1_OUT3), 
        .IN4(Tg1_OUT4) );
  NOR2X0 Tg1_Trojan5 ( .IN1(n1391), .IN2(n931), .QN(Tg1_OUT5) );
  NOR2X0 Tg1_Trojan6 ( .IN1(n857), .IN2(n902), .QN(Tg1_OUT6) );
  NOR2X0 Tg1_Trojan7 ( .IN1(n1239), .IN2(n1239), .QN(Tg1_OUT7) );
  NOR2X0 Tg1_Trojan8 ( .IN1(n1055), .IN2(n1016), .QN(Tg1_OUT8) );
  AND4X1 Tg1_Trojan5678 ( .IN1(Tg1_OUT5), .IN2(Tg1_OUT6), .IN3(Tg1_OUT7), 
        .IN4(Tg1_OUT8) );
  AND2X2 Tg2_Trojan1 ( .IN1(n78), .IN2(n51), .Q(Tg2_OUT1) );
  AND2X2 Tg2_Trojan2 ( .IN1(n51), .IN2(n51), .Q(Tg2_OUT2) );
  AND2X2 Tg2_Trojan3 ( .IN1(n51), .IN2(n51), .Q(Tg2_OUT3) );
  AND2X2 Tg2_Trojan4 ( .IN1(n51), .IN2(n51), .Q(Tg2_OUT4) );
  AND4X1 Tg2_Trojan1234 ( .IN1(Tg2_OUT1), .IN2(Tg2_OUT2), .IN3(Tg2_OUT3), 
        .IN4(Tg2_OUT4) );
  AND2X2 Tg2_Trojan5 ( .IN1(n1161), .IN2(n1154), .Q(Tg2_OUT5) );
  AND2X2 Tg2_Trojan6 ( .IN1(n179), .IN2(n145), .Q(Tg2_OUT6) );
  AND2X2 Tg2_Trojan7 ( .IN1(n147), .IN2(n1107), .Q(Tg2_OUT7) );
  AND2X2 Tg2_Trojan8 ( .IN1(n363), .IN2(n238), .Q(Tg2_OUT8) );
  AND4X1 Tg2_Trojan5678 ( .IN1(Tg2_OUT5), .IN2(Tg2_OUT6), .IN3(Tg2_OUT7), 
        .IN4(Tg2_OUT8) );
  INVX0 TrojanINVtest_se ( .INP(n3475), .ZN(test_se_NOT) );
  AND2X2 Trojan_Trigger ( .IN1(1'b1), .IN2(test_se_NOT), .Q(Trigger_select) );
  MUX21X2 Trojan_Paylaod ( .IN1(g1200), .IN2(n495), .S(Trigger_select), .Q(
        g4207) );
  NBUFFX2 U3406 ( .INP(n3566), .Z(n3516) );
  NBUFFX2 U3407 ( .INP(n3566), .Z(n3517) );
  NBUFFX2 U3408 ( .INP(n3566), .Z(n3515) );
  NBUFFX2 U3409 ( .INP(n3563), .Z(n3528) );
  NBUFFX2 U3410 ( .INP(n3565), .Z(n3521) );
  NBUFFX2 U3411 ( .INP(n3559), .Z(n3550) );
  NBUFFX2 U3412 ( .INP(n3560), .Z(n3547) );
  NBUFFX2 U3413 ( .INP(n3560), .Z(n3546) );
  NBUFFX2 U3414 ( .INP(n3560), .Z(n3544) );
  NBUFFX2 U3415 ( .INP(n3564), .Z(n3524) );
  NBUFFX2 U3416 ( .INP(n3561), .Z(n3540) );
  NBUFFX2 U3417 ( .INP(n3561), .Z(n3538) );
  NBUFFX2 U3418 ( .INP(n3564), .Z(n3526) );
  NBUFFX2 U3419 ( .INP(n3563), .Z(n3530) );
  NBUFFX2 U3420 ( .INP(n3558), .Z(n3556) );
  NBUFFX2 U3421 ( .INP(n3564), .Z(n3527) );
  NBUFFX2 U3422 ( .INP(n3559), .Z(n3551) );
  NBUFFX2 U3423 ( .INP(n3559), .Z(n3552) );
  NBUFFX2 U3424 ( .INP(n3562), .Z(n3536) );
  NBUFFX2 U3425 ( .INP(n3559), .Z(n3549) );
  NBUFFX2 U3426 ( .INP(n3563), .Z(n3532) );
  NBUFFX2 U3427 ( .INP(n3560), .Z(n3545) );
  NBUFFX2 U3428 ( .INP(n3561), .Z(n3541) );
  NBUFFX2 U3429 ( .INP(n3561), .Z(n3539) );
  NBUFFX2 U3430 ( .INP(n3562), .Z(n3533) );
  NBUFFX2 U3431 ( .INP(n3565), .Z(n3522) );
  NBUFFX2 U3432 ( .INP(n3559), .Z(n3548) );
  NBUFFX2 U3433 ( .INP(n3563), .Z(n3529) );
  NBUFFX2 U3434 ( .INP(n3561), .Z(n3542) );
  NBUFFX2 U3435 ( .INP(n3562), .Z(n3535) );
  NBUFFX2 U3436 ( .INP(n3560), .Z(n3543) );
  NBUFFX2 U3437 ( .INP(n3562), .Z(n3534) );
  NBUFFX2 U3438 ( .INP(n3565), .Z(n3518) );
  NBUFFX2 U3439 ( .INP(n3563), .Z(n3531) );
  NBUFFX2 U3440 ( .INP(n3564), .Z(n3523) );
  NBUFFX2 U3441 ( .INP(n3558), .Z(n3554) );
  NBUFFX2 U3442 ( .INP(n3558), .Z(n3553) );
  NBUFFX2 U3443 ( .INP(n3565), .Z(n3519) );
  NBUFFX2 U3444 ( .INP(n3565), .Z(n3520) );
  NBUFFX2 U3445 ( .INP(n3564), .Z(n3525) );
  NBUFFX2 U3446 ( .INP(n3558), .Z(n3555) );
  NBUFFX2 U3447 ( .INP(n3562), .Z(n3537) );
  NBUFFX2 U3448 ( .INP(n3558), .Z(n3557) );
  NBUFFX2 U3449 ( .INP(n3504), .Z(n3390) );
  NBUFFX2 U3450 ( .INP(n3504), .Z(n3391) );
  NBUFFX2 U3451 ( .INP(n3503), .Z(n3392) );
  NBUFFX2 U3452 ( .INP(n3503), .Z(n3393) );
  NBUFFX2 U3453 ( .INP(n3503), .Z(n3394) );
  NBUFFX2 U3454 ( .INP(n3502), .Z(n3395) );
  NBUFFX2 U3455 ( .INP(n3502), .Z(n3396) );
  NBUFFX2 U3456 ( .INP(n3502), .Z(n3397) );
  NBUFFX2 U3457 ( .INP(n3501), .Z(n3398) );
  NBUFFX2 U3458 ( .INP(n3501), .Z(n3399) );
  NBUFFX2 U3459 ( .INP(n3501), .Z(n3400) );
  NBUFFX2 U3460 ( .INP(n3500), .Z(n3401) );
  NBUFFX2 U3461 ( .INP(n3500), .Z(n3402) );
  NBUFFX2 U3462 ( .INP(n3500), .Z(n3403) );
  NBUFFX2 U3463 ( .INP(n3499), .Z(n3404) );
  NBUFFX2 U3464 ( .INP(n3499), .Z(n3405) );
  NBUFFX2 U3465 ( .INP(n3499), .Z(n3406) );
  NBUFFX2 U3466 ( .INP(n3498), .Z(n3407) );
  NBUFFX2 U3467 ( .INP(n3498), .Z(n3408) );
  NBUFFX2 U3468 ( .INP(n3498), .Z(n3409) );
  NBUFFX2 U3469 ( .INP(n3497), .Z(n3410) );
  NBUFFX2 U3470 ( .INP(n3497), .Z(n3411) );
  NBUFFX2 U3471 ( .INP(n3497), .Z(n3412) );
  NBUFFX2 U3472 ( .INP(n3496), .Z(n3413) );
  NBUFFX2 U3473 ( .INP(n3496), .Z(n3414) );
  NBUFFX2 U3474 ( .INP(n3496), .Z(n3415) );
  NBUFFX2 U3475 ( .INP(n3495), .Z(n3416) );
  NBUFFX2 U3476 ( .INP(n3495), .Z(n3417) );
  NBUFFX2 U3477 ( .INP(n3495), .Z(n3418) );
  NBUFFX2 U3478 ( .INP(n3494), .Z(n3419) );
  NBUFFX2 U3479 ( .INP(n3494), .Z(n3420) );
  NBUFFX2 U3480 ( .INP(n3494), .Z(n3421) );
  NBUFFX2 U3481 ( .INP(n3493), .Z(n3422) );
  NBUFFX2 U3482 ( .INP(n3493), .Z(n3423) );
  NBUFFX2 U3483 ( .INP(n3493), .Z(n3424) );
  NBUFFX2 U3484 ( .INP(n3492), .Z(n3425) );
  NBUFFX2 U3485 ( .INP(n3492), .Z(n3426) );
  NBUFFX2 U3486 ( .INP(n3492), .Z(n3427) );
  NBUFFX2 U3487 ( .INP(n3491), .Z(n3428) );
  NBUFFX2 U3488 ( .INP(n3491), .Z(n3429) );
  NBUFFX2 U3489 ( .INP(n3491), .Z(n3430) );
  NBUFFX2 U3490 ( .INP(n3490), .Z(n3431) );
  NBUFFX2 U3491 ( .INP(n3490), .Z(n3432) );
  NBUFFX2 U3492 ( .INP(n3490), .Z(n3433) );
  NBUFFX2 U3493 ( .INP(n3489), .Z(n3434) );
  NBUFFX2 U3494 ( .INP(n3489), .Z(n3435) );
  NBUFFX2 U3495 ( .INP(n3489), .Z(n3436) );
  NBUFFX2 U3496 ( .INP(n3488), .Z(n3437) );
  NBUFFX2 U3497 ( .INP(n3488), .Z(n3438) );
  NBUFFX2 U3498 ( .INP(n3488), .Z(n3439) );
  NBUFFX2 U3499 ( .INP(n3487), .Z(n3440) );
  NBUFFX2 U3500 ( .INP(n3487), .Z(n3441) );
  NBUFFX2 U3501 ( .INP(n3487), .Z(n3442) );
  NBUFFX2 U3502 ( .INP(n3486), .Z(n3443) );
  NBUFFX2 U3503 ( .INP(n3486), .Z(n3444) );
  NBUFFX2 U3504 ( .INP(n3486), .Z(n3445) );
  NBUFFX2 U3505 ( .INP(n3485), .Z(n3446) );
  NBUFFX2 U3506 ( .INP(n3485), .Z(n3447) );
  NBUFFX2 U3507 ( .INP(n3485), .Z(n3448) );
  NBUFFX2 U3508 ( .INP(n3484), .Z(n3449) );
  NBUFFX2 U3509 ( .INP(n3484), .Z(n3450) );
  NBUFFX2 U3510 ( .INP(n3484), .Z(n3451) );
  NBUFFX2 U3511 ( .INP(n3483), .Z(n3452) );
  NBUFFX2 U3512 ( .INP(n3483), .Z(n3453) );
  NBUFFX2 U3513 ( .INP(n3483), .Z(n3454) );
  NBUFFX2 U3514 ( .INP(n3482), .Z(n3455) );
  NBUFFX2 U3515 ( .INP(n3482), .Z(n3456) );
  NBUFFX2 U3516 ( .INP(n3482), .Z(n3457) );
  NBUFFX2 U3517 ( .INP(n3481), .Z(n3458) );
  NBUFFX2 U3518 ( .INP(n3481), .Z(n3459) );
  NBUFFX2 U3519 ( .INP(n3481), .Z(n3460) );
  NBUFFX2 U3520 ( .INP(n3480), .Z(n3461) );
  NBUFFX2 U3521 ( .INP(n3480), .Z(n3462) );
  NBUFFX2 U3522 ( .INP(n3480), .Z(n3463) );
  NBUFFX2 U3523 ( .INP(n3479), .Z(n3464) );
  NBUFFX2 U3524 ( .INP(n3479), .Z(n3465) );
  NBUFFX2 U3525 ( .INP(n3479), .Z(n3466) );
  NBUFFX2 U3526 ( .INP(n3478), .Z(n3467) );
  NBUFFX2 U3527 ( .INP(n3478), .Z(n3468) );
  NBUFFX2 U3528 ( .INP(n3478), .Z(n3469) );
  NBUFFX2 U3529 ( .INP(n3477), .Z(n3470) );
  NBUFFX2 U3530 ( .INP(n3477), .Z(n3471) );
  NBUFFX2 U3531 ( .INP(n3477), .Z(n3472) );
  NBUFFX2 U3532 ( .INP(n3476), .Z(n3473) );
  NBUFFX2 U3533 ( .INP(n3476), .Z(n3474) );
  NBUFFX2 U3534 ( .INP(n3476), .Z(n3475) );
  NBUFFX2 U3535 ( .INP(n3514), .Z(n3476) );
  NBUFFX2 U3536 ( .INP(n3514), .Z(n3477) );
  NBUFFX2 U3537 ( .INP(n3513), .Z(n3478) );
  NBUFFX2 U3538 ( .INP(n3513), .Z(n3479) );
  NBUFFX2 U3539 ( .INP(n3513), .Z(n3480) );
  NBUFFX2 U3540 ( .INP(n3512), .Z(n3481) );
  NBUFFX2 U3541 ( .INP(n3512), .Z(n3482) );
  NBUFFX2 U3542 ( .INP(n3512), .Z(n3483) );
  NBUFFX2 U3543 ( .INP(n3511), .Z(n3484) );
  NBUFFX2 U3544 ( .INP(n3511), .Z(n3485) );
  NBUFFX2 U3545 ( .INP(n3511), .Z(n3486) );
  NBUFFX2 U3546 ( .INP(n3510), .Z(n3487) );
  NBUFFX2 U3547 ( .INP(n3510), .Z(n3488) );
  NBUFFX2 U3548 ( .INP(n3510), .Z(n3489) );
  NBUFFX2 U3549 ( .INP(n3509), .Z(n3490) );
  NBUFFX2 U3550 ( .INP(n3509), .Z(n3491) );
  NBUFFX2 U3551 ( .INP(n3509), .Z(n3492) );
  NBUFFX2 U3552 ( .INP(n3508), .Z(n3493) );
  NBUFFX2 U3553 ( .INP(n3508), .Z(n3494) );
  NBUFFX2 U3554 ( .INP(n3508), .Z(n3495) );
  NBUFFX2 U3555 ( .INP(n3507), .Z(n3496) );
  NBUFFX2 U3556 ( .INP(n3507), .Z(n3497) );
  NBUFFX2 U3557 ( .INP(n3507), .Z(n3498) );
  NBUFFX2 U3558 ( .INP(n3506), .Z(n3499) );
  NBUFFX2 U3559 ( .INP(n3506), .Z(n3500) );
  NBUFFX2 U3560 ( .INP(n3506), .Z(n3501) );
  NBUFFX2 U3561 ( .INP(n3505), .Z(n3502) );
  NBUFFX2 U3562 ( .INP(n3505), .Z(n3503) );
  NBUFFX2 U3563 ( .INP(n3505), .Z(n3504) );
  NBUFFX2 U3564 ( .INP(test_se), .Z(n3505) );
  NBUFFX2 U3565 ( .INP(n3510), .Z(n3506) );
  NBUFFX2 U3566 ( .INP(n3487), .Z(n3507) );
  NBUFFX2 U3567 ( .INP(n3488), .Z(n3508) );
  NBUFFX2 U3568 ( .INP(n3489), .Z(n3509) );
  NBUFFX2 U3569 ( .INP(test_se), .Z(n3510) );
  NBUFFX2 U3570 ( .INP(test_se), .Z(n3511) );
  NBUFFX2 U3571 ( .INP(n3504), .Z(n3512) );
  NBUFFX2 U3572 ( .INP(test_se), .Z(n3513) );
  NBUFFX2 U3573 ( .INP(n3505), .Z(n3514) );
  NBUFFX2 U3574 ( .INP(n3569), .Z(n3558) );
  NBUFFX2 U3575 ( .INP(n3569), .Z(n3559) );
  NBUFFX2 U3576 ( .INP(n3569), .Z(n3560) );
  NBUFFX2 U3577 ( .INP(n3568), .Z(n3561) );
  NBUFFX2 U3578 ( .INP(n3568), .Z(n3562) );
  NBUFFX2 U3579 ( .INP(n3568), .Z(n3563) );
  NBUFFX2 U3580 ( .INP(n3567), .Z(n3564) );
  NBUFFX2 U3581 ( .INP(n3567), .Z(n3565) );
  NBUFFX2 U3582 ( .INP(n3567), .Z(n3566) );
  NBUFFX2 U3583 ( .INP(CK), .Z(n3567) );
  NBUFFX2 U3584 ( .INP(CK), .Z(n3568) );
  NBUFFX2 U3585 ( .INP(CK), .Z(n3569) );
  OR2X1 U3587 ( .IN1(n3570), .IN2(n3571), .Q(n962) );
  AND2X1 U3588 ( .IN1(n3572), .IN2(n1696), .Q(n3571) );
  AND2X1 U3589 ( .IN1(n3573), .IN2(g731), .Q(n3570) );
  OR2X1 U3590 ( .IN1(n3574), .IN2(n3575), .Q(n917) );
  AND2X1 U3591 ( .IN1(n3576), .IN2(n1697), .Q(n3575) );
  AND2X1 U3592 ( .IN1(n3577), .IN2(g1945), .Q(n3574) );
  AND2X1 U3593 ( .IN1(n804), .IN2(n3578), .Q(n838) );
  INVX0 U3594 ( .INP(n3579), .ZN(n665) );
  INVX0 U3595 ( .INP(n3580), .ZN(n655) );
  INVX0 U3596 ( .INP(n3581), .ZN(n628) );
  INVX0 U3597 ( .INP(n3582), .ZN(n438) );
  OR2X1 U3598 ( .IN1(n3583), .IN2(n3317), .Q(n3582) );
  AND2X1 U3599 ( .IN1(n3584), .IN2(n3585), .Q(n3583) );
  OR2X1 U3600 ( .IN1(g750), .IN2(n1647), .Q(n3584) );
  INVX0 U3601 ( .INP(n3586), .ZN(n386) );
  INVX0 U3602 ( .INP(n3587), .ZN(n3376) );
  INVX0 U3603 ( .INP(n3588), .ZN(n256) );
  INVX0 U3604 ( .INP(n3589), .ZN(n180) );
  OR2X1 U3605 ( .IN1(n3590), .IN2(n3591), .Q(n1588) );
  OR2X1 U3606 ( .IN1(g42), .IN2(n3592), .Q(n3591) );
  OR2X1 U3607 ( .IN1(n3592), .IN2(n3593), .Q(n1587) );
  OR2X1 U3608 ( .IN1(n3594), .IN2(n3593), .Q(n1586) );
  OR2X1 U3609 ( .IN1(n3590), .IN2(n3595), .Q(n1585) );
  OR2X1 U3610 ( .IN1(g42), .IN2(n3594), .Q(n3595) );
  OR2X1 U3611 ( .IN1(n3351), .IN2(n3352), .Q(n1214) );
  INVX0 U3612 ( .INP(n3596), .ZN(n1) );
  AND2X1 U3613 ( .IN1(n3323), .IN2(n3362), .Q(n3596) );
  AND2X1 U3614 ( .IN1(g18), .IN2(n3597), .Q(g9721) );
  OR2X1 U3615 ( .IN1(n3598), .IN2(n3599), .Q(n3597) );
  AND2X1 U3616 ( .IN1(n3600), .IN2(g611), .Q(n3599) );
  INVX0 U3617 ( .INP(n3601), .ZN(n3600) );
  AND2X1 U3618 ( .IN1(n1609), .IN2(n3601), .Q(n3598) );
  OR2X1 U3619 ( .IN1(n3602), .IN2(n3603), .Q(n3601) );
  AND2X1 U3620 ( .IN1(n3604), .IN2(n3605), .Q(n3602) );
  OR2X1 U3621 ( .IN1(n3606), .IN2(g617), .Q(n3605) );
  AND2X1 U3622 ( .IN1(n3607), .IN2(n3608), .Q(n3606) );
  AND2X1 U3623 ( .IN1(n3609), .IN2(g18), .Q(g9555) );
  AND2X1 U3624 ( .IN1(n3610), .IN2(n3611), .Q(n3609) );
  OR2X1 U3625 ( .IN1(n806), .IN2(g1834), .Q(n3611) );
  INVX0 U3626 ( .INP(n3612), .ZN(n3610) );
  AND2X1 U3627 ( .IN1(g1834), .IN2(n3613), .Q(n3612) );
  AND2X1 U3628 ( .IN1(n808), .IN2(n926), .Q(n3613) );
  OR2X1 U3629 ( .IN1(n3614), .IN2(g1840), .Q(n808) );
  AND2X1 U3630 ( .IN1(n366), .IN2(n3615), .Q(n3614) );
  INVX0 U3631 ( .INP(n3616), .ZN(n366) );
  OR2X1 U3632 ( .IN1(n3617), .IN2(n3618), .Q(g9451) );
  OR2X1 U3633 ( .IN1(g31), .IN2(g30), .Q(n3618) );
  AND2X1 U3634 ( .IN1(n3619), .IN2(g18), .Q(g9272) );
  AND2X1 U3635 ( .IN1(n3620), .IN2(n3621), .Q(n3619) );
  OR2X1 U3636 ( .IN1(n1605), .IN2(n3622), .Q(n3621) );
  INVX0 U3637 ( .INP(n3623), .ZN(n3620) );
  AND2X1 U3638 ( .IN1(n1605), .IN2(n3624), .Q(n3623) );
  AND2X1 U3639 ( .IN1(n3625), .IN2(n3622), .Q(n3624) );
  OR2X1 U3640 ( .IN1(n3626), .IN2(n3615), .Q(n3622) );
  AND2X1 U3641 ( .IN1(n3627), .IN2(n3628), .Q(n3626) );
  OR2X1 U3642 ( .IN1(n1643), .IN2(n817), .Q(n3628) );
  AND2X1 U3643 ( .IN1(n3629), .IN2(g18), .Q(g9269) );
  AND2X1 U3644 ( .IN1(n3630), .IN2(n3631), .Q(n3629) );
  OR2X1 U3645 ( .IN1(n3632), .IN2(g1822), .Q(n3631) );
  INVX0 U3646 ( .INP(n3633), .ZN(n3632) );
  OR2X1 U3647 ( .IN1(n1643), .IN2(n3633), .Q(n3630) );
  OR2X1 U3648 ( .IN1(n3634), .IN2(n3615), .Q(n3633) );
  AND2X1 U3649 ( .IN1(n3635), .IN2(n3636), .Q(n3634) );
  AND2X1 U3650 ( .IN1(n822), .IN2(n3637), .Q(n3635) );
  AND2X1 U3651 ( .IN1(n3638), .IN2(g18), .Q(g9266) );
  AND2X1 U3652 ( .IN1(n3639), .IN2(n3640), .Q(n3638) );
  OR2X1 U3653 ( .IN1(n3641), .IN2(g1814), .Q(n3640) );
  INVX0 U3654 ( .INP(n3642), .ZN(n3641) );
  OR2X1 U3655 ( .IN1(n1608), .IN2(n3642), .Q(n3639) );
  OR2X1 U3656 ( .IN1(n3643), .IN2(n3615), .Q(n3642) );
  AND2X1 U3657 ( .IN1(n3644), .IN2(n3636), .Q(n3643) );
  OR2X1 U3658 ( .IN1(n817), .IN2(g1822), .Q(n3636) );
  AND2X1 U3659 ( .IN1(n3645), .IN2(n3616), .Q(n3644) );
  AND2X1 U3660 ( .IN1(n3646), .IN2(g18), .Q(g9150) );
  AND2X1 U3661 ( .IN1(n3647), .IN2(n3648), .Q(n3646) );
  OR2X1 U3662 ( .IN1(n3649), .IN2(n3650), .Q(n3648) );
  OR2X1 U3663 ( .IN1(n3651), .IN2(g605), .Q(n3650) );
  INVX0 U3664 ( .INP(n3652), .ZN(n3649) );
  OR2X1 U3665 ( .IN1(n1593), .IN2(n3652), .Q(n3647) );
  OR2X1 U3666 ( .IN1(n3653), .IN2(n3608), .Q(n3652) );
  AND2X1 U3667 ( .IN1(n3654), .IN2(n3655), .Q(n3653) );
  AND2X1 U3668 ( .IN1(n3656), .IN2(n3657), .Q(n3655) );
  OR2X1 U3669 ( .IN1(n1644), .IN2(n3658), .Q(n3656) );
  AND2X1 U3670 ( .IN1(n3659), .IN2(n3660), .Q(n3654) );
  OR2X1 U3671 ( .IN1(n3661), .IN2(g622), .Q(n3660) );
  OR2X1 U3672 ( .IN1(g605), .IN2(n3662), .Q(n3659) );
  AND2X1 U3673 ( .IN1(g18), .IN2(n3663), .Q(g9124) );
  OR2X1 U3674 ( .IN1(n3664), .IN2(n3665), .Q(n3663) );
  AND2X1 U3675 ( .IN1(n1644), .IN2(n3666), .Q(n3665) );
  INVX0 U3676 ( .INP(n836), .ZN(n3666) );
  AND2X1 U3677 ( .IN1(n836), .IN2(g599), .Q(n3664) );
  AND2X1 U3678 ( .IN1(g18), .IN2(n3667), .Q(g9110) );
  OR2X1 U3679 ( .IN1(n3668), .IN2(n3669), .Q(n3667) );
  AND2X1 U3680 ( .IN1(n3670), .IN2(g591), .Q(n3669) );
  AND2X1 U3681 ( .IN1(n1607), .IN2(n3671), .Q(n3668) );
  INVX0 U3682 ( .INP(n3670), .ZN(n3671) );
  AND2X1 U3683 ( .IN1(n837), .IN2(n3672), .Q(n3670) );
  OR2X1 U3684 ( .IN1(n3608), .IN2(n3673), .Q(n3672) );
  AND2X1 U3685 ( .IN1(n3662), .IN2(n3661), .Q(n3673) );
  OR2X1 U3686 ( .IN1(n3658), .IN2(n3674), .Q(n837) );
  OR2X1 U3687 ( .IN1(g599), .IN2(n3608), .Q(n3674) );
  OR2X1 U3688 ( .IN1(n3675), .IN2(n3676), .Q(g8973) );
  AND2X1 U3689 ( .IN1(n3677), .IN2(n3678), .Q(n3675) );
  AND2X1 U3690 ( .IN1(n3679), .IN2(n3680), .Q(n3677) );
  OR2X1 U3691 ( .IN1(n3681), .IN2(g658), .Q(n3680) );
  INVX0 U3692 ( .INP(n3682), .ZN(n3681) );
  OR2X1 U3693 ( .IN1(n1615), .IN2(n3682), .Q(n3679) );
  OR2X1 U3694 ( .IN1(n3683), .IN2(n3684), .Q(n3682) );
  AND2X1 U3695 ( .IN1(n3336), .IN2(n3685), .Q(n3683) );
  OR2X1 U3696 ( .IN1(n3686), .IN2(n3687), .Q(g8945) );
  AND2X1 U3697 ( .IN1(n3688), .IN2(n3689), .Q(n3686) );
  AND2X1 U3698 ( .IN1(n3690), .IN2(n3691), .Q(n3688) );
  OR2X1 U3699 ( .IN1(n3692), .IN2(g1945), .Q(n3691) );
  OR2X1 U3700 ( .IN1(n1697), .IN2(n3693), .Q(n3690) );
  INVX0 U3701 ( .INP(n3692), .ZN(n3693) );
  OR2X1 U3702 ( .IN1(n3694), .IN2(n3695), .Q(n3692) );
  AND2X1 U3703 ( .IN1(n3696), .IN2(n3697), .Q(n3695) );
  AND2X1 U3704 ( .IN1(n3698), .IN2(n3699), .Q(n3696) );
  INVX0 U3705 ( .INP(n3700), .ZN(n3699) );
  OR2X1 U3706 ( .IN1(n3576), .IN2(n3577), .Q(n3698) );
  INVX0 U3707 ( .INP(n857), .ZN(n3577) );
  OR2X1 U3708 ( .IN1(n1694), .IN2(n3701), .Q(n857) );
  INVX0 U3709 ( .INP(n3702), .ZN(n3576) );
  OR2X1 U3710 ( .IN1(n3703), .IN2(n3704), .Q(n3702) );
  OR2X1 U3711 ( .IN1(g1927), .IN2(n3705), .Q(n3704) );
  OR2X1 U3712 ( .IN1(g1918), .IN2(g1909), .Q(n3705) );
  OR2X1 U3713 ( .IN1(n3706), .IN2(n3707), .Q(n3703) );
  OR2X1 U3714 ( .IN1(g1900), .IN2(g1936), .Q(n3707) );
  AND2X1 U3715 ( .IN1(n3708), .IN2(g1950), .Q(n3694) );
  OR2X1 U3716 ( .IN1(n3709), .IN2(n3687), .Q(g8944) );
  AND2X1 U3717 ( .IN1(n3710), .IN2(n3689), .Q(n3709) );
  AND2X1 U3718 ( .IN1(n3711), .IN2(n3712), .Q(n3710) );
  INVX0 U3719 ( .INP(n3713), .ZN(n3712) );
  AND2X1 U3720 ( .IN1(n3714), .IN2(n1694), .Q(n3713) );
  OR2X1 U3721 ( .IN1(n1694), .IN2(n3714), .Q(n3711) );
  OR2X1 U3722 ( .IN1(n3715), .IN2(n3700), .Q(n3714) );
  AND2X1 U3723 ( .IN1(n3716), .IN2(n3717), .Q(n3715) );
  OR2X1 U3724 ( .IN1(g1927), .IN2(n3718), .Q(n3717) );
  AND2X1 U3725 ( .IN1(n3719), .IN2(n3720), .Q(n3716) );
  OR2X1 U3726 ( .IN1(n3701), .IN2(n3708), .Q(n3720) );
  OR2X1 U3727 ( .IN1(n3721), .IN2(n3722), .Q(n3701) );
  OR2X1 U3728 ( .IN1(n3723), .IN2(n3724), .Q(n3722) );
  INVX0 U3729 ( .INP(n921), .ZN(n3724) );
  OR2X1 U3730 ( .IN1(n1675), .IN2(n3725), .Q(n3721) );
  OR2X1 U3731 ( .IN1(n3330), .IN2(n3274), .Q(n3725) );
  OR2X1 U3732 ( .IN1(n3226), .IN2(n3697), .Q(n3719) );
  OR2X1 U3733 ( .IN1(n3726), .IN2(n3687), .Q(g8943) );
  AND2X1 U3734 ( .IN1(n3727), .IN2(n3689), .Q(n3726) );
  AND2X1 U3735 ( .IN1(n3728), .IN2(n3729), .Q(n3727) );
  OR2X1 U3736 ( .IN1(n3730), .IN2(g1882), .Q(n3729) );
  INVX0 U3737 ( .INP(n3731), .ZN(n3730) );
  OR2X1 U3738 ( .IN1(n1663), .IN2(n3731), .Q(n3728) );
  OR2X1 U3739 ( .IN1(n3700), .IN2(n3732), .Q(n3731) );
  OR2X1 U3740 ( .IN1(n3733), .IN2(n3734), .Q(n3732) );
  AND2X1 U3741 ( .IN1(n3735), .IN2(n3697), .Q(n3734) );
  OR2X1 U3742 ( .IN1(n3736), .IN2(n3737), .Q(n3735) );
  AND2X1 U3743 ( .IN1(n3738), .IN2(g1872), .Q(n3737) );
  AND2X1 U3744 ( .IN1(n1616), .IN2(n3739), .Q(n3736) );
  AND2X1 U3745 ( .IN1(n3194), .IN2(n3708), .Q(n3733) );
  OR2X1 U3746 ( .IN1(n3740), .IN2(n3687), .Q(g8941) );
  AND2X1 U3747 ( .IN1(n3741), .IN2(n3689), .Q(n3740) );
  AND2X1 U3748 ( .IN1(n3742), .IN2(n3743), .Q(n3741) );
  OR2X1 U3749 ( .IN1(n3744), .IN2(g1927), .Q(n3743) );
  INVX0 U3750 ( .INP(n3745), .ZN(n3744) );
  OR2X1 U3751 ( .IN1(n3347), .IN2(n3745), .Q(n3742) );
  OR2X1 U3752 ( .IN1(n3746), .IN2(n3700), .Q(n3745) );
  AND2X1 U3753 ( .IN1(n3747), .IN2(n3748), .Q(n3746) );
  OR2X1 U3754 ( .IN1(n3274), .IN2(n3749), .Q(n3748) );
  AND2X1 U3755 ( .IN1(n3750), .IN2(n3718), .Q(n3747) );
  OR2X1 U3756 ( .IN1(g1918), .IN2(n3751), .Q(n3718) );
  OR2X1 U3757 ( .IN1(n3697), .IN2(n3227), .Q(n3750) );
  OR2X1 U3758 ( .IN1(n3752), .IN2(n3687), .Q(g8940) );
  AND2X1 U3759 ( .IN1(n3753), .IN2(n3689), .Q(n3752) );
  AND2X1 U3760 ( .IN1(n3754), .IN2(n3755), .Q(n3753) );
  OR2X1 U3761 ( .IN1(n3756), .IN2(g1918), .Q(n3755) );
  INVX0 U3762 ( .INP(n3757), .ZN(n3756) );
  OR2X1 U3763 ( .IN1(n3274), .IN2(n3757), .Q(n3754) );
  OR2X1 U3764 ( .IN1(n3758), .IN2(n3700), .Q(n3757) );
  AND2X1 U3765 ( .IN1(n3759), .IN2(n3760), .Q(n3758) );
  OR2X1 U3766 ( .IN1(n3697), .IN2(n1718), .Q(n3760) );
  AND2X1 U3767 ( .IN1(n3749), .IN2(n3751), .Q(n3759) );
  OR2X1 U3768 ( .IN1(n3761), .IN2(n3762), .Q(n3751) );
  OR2X1 U3769 ( .IN1(g1900), .IN2(g1909), .Q(n3762) );
  OR2X1 U3770 ( .IN1(n3763), .IN2(n3764), .Q(n3749) );
  OR2X1 U3771 ( .IN1(n3330), .IN2(n1675), .Q(n3764) );
  OR2X1 U3772 ( .IN1(n3765), .IN2(n3687), .Q(g8939) );
  AND2X1 U3773 ( .IN1(n3766), .IN2(n3689), .Q(n3765) );
  AND2X1 U3774 ( .IN1(n3767), .IN2(n3768), .Q(n3766) );
  OR2X1 U3775 ( .IN1(n3769), .IN2(g1909), .Q(n3768) );
  INVX0 U3776 ( .INP(n3770), .ZN(n3769) );
  OR2X1 U3777 ( .IN1(n3330), .IN2(n3770), .Q(n3767) );
  OR2X1 U3778 ( .IN1(n3771), .IN2(n3700), .Q(n3770) );
  AND2X1 U3779 ( .IN1(n3772), .IN2(n3773), .Q(n3771) );
  OR2X1 U3780 ( .IN1(n3697), .IN2(n3224), .Q(n3773) );
  AND2X1 U3781 ( .IN1(n3774), .IN2(n3775), .Q(n3772) );
  OR2X1 U3782 ( .IN1(n1675), .IN2(n3763), .Q(n3775) );
  OR2X1 U3783 ( .IN1(g1900), .IN2(n3761), .Q(n3774) );
  OR2X1 U3784 ( .IN1(n3776), .IN2(n3687), .Q(g8938) );
  AND2X1 U3785 ( .IN1(n3777), .IN2(n3689), .Q(n3776) );
  AND2X1 U3786 ( .IN1(n3778), .IN2(n3779), .Q(n3777) );
  INVX0 U3787 ( .INP(n3780), .ZN(n3779) );
  AND2X1 U3788 ( .IN1(n3781), .IN2(n1675), .Q(n3780) );
  OR2X1 U3789 ( .IN1(n1675), .IN2(n3781), .Q(n3778) );
  OR2X1 U3790 ( .IN1(n3782), .IN2(n3700), .Q(n3781) );
  AND2X1 U3791 ( .IN1(n3783), .IN2(n3784), .Q(n3782) );
  AND2X1 U3792 ( .IN1(n3761), .IN2(n3763), .Q(n3784) );
  OR2X1 U3793 ( .IN1(n3708), .IN2(n3785), .Q(n3763) );
  OR2X1 U3794 ( .IN1(n1657), .IN2(n3723), .Q(n3785) );
  OR2X1 U3795 ( .IN1(n3708), .IN2(n3706), .Q(n3761) );
  OR2X1 U3796 ( .IN1(n3786), .IN2(g1891), .Q(n3706) );
  OR2X1 U3797 ( .IN1(n3697), .IN2(n3342), .Q(n3783) );
  OR2X1 U3798 ( .IN1(n3787), .IN2(n3687), .Q(g8937) );
  AND2X1 U3799 ( .IN1(n3788), .IN2(n3689), .Q(n3787) );
  AND2X1 U3800 ( .IN1(n3789), .IN2(n3790), .Q(n3788) );
  OR2X1 U3801 ( .IN1(g1891), .IN2(n3791), .Q(n3790) );
  INVX0 U3802 ( .INP(n3792), .ZN(n3791) );
  OR2X1 U3803 ( .IN1(n1657), .IN2(n3792), .Q(n3789) );
  AND2X1 U3804 ( .IN1(n3793), .IN2(n3794), .Q(n3792) );
  OR2X1 U3805 ( .IN1(n3795), .IN2(n3708), .Q(n3794) );
  OR2X1 U3806 ( .IN1(n3796), .IN2(n3700), .Q(n3795) );
  AND2X1 U3807 ( .IN1(n3723), .IN2(n3786), .Q(n3796) );
  OR2X1 U3808 ( .IN1(g1882), .IN2(n3797), .Q(n3786) );
  OR2X1 U3809 ( .IN1(n3739), .IN2(g1872), .Q(n3797) );
  INVX0 U3810 ( .INP(n3738), .ZN(n3739) );
  OR2X1 U3811 ( .IN1(n3738), .IN2(n3798), .Q(n3723) );
  OR2X1 U3812 ( .IN1(n1663), .IN2(n1616), .Q(n3798) );
  AND2X1 U3813 ( .IN1(n3799), .IN2(n3627), .Q(n3738) );
  AND2X1 U3814 ( .IN1(n3800), .IN2(n3637), .Q(n3627) );
  OR2X1 U3815 ( .IN1(g1828), .IN2(n3645), .Q(n3800) );
  OR2X1 U3816 ( .IN1(g1822), .IN2(n1608), .Q(n3799) );
  OR2X1 U3817 ( .IN1(n3697), .IN2(n3343), .Q(n3793) );
  OR2X1 U3818 ( .IN1(n3801), .IN2(n3676), .Q(g8926) );
  AND2X1 U3819 ( .IN1(n3802), .IN2(n3678), .Q(n3801) );
  AND2X1 U3820 ( .IN1(n3803), .IN2(n3804), .Q(n3802) );
  OR2X1 U3821 ( .IN1(n898), .IN2(g731), .Q(n3804) );
  OR2X1 U3822 ( .IN1(n1696), .IN2(n3805), .Q(n3803) );
  INVX0 U3823 ( .INP(n898), .ZN(n3805) );
  OR2X1 U3824 ( .IN1(n3806), .IN2(n3807), .Q(n898) );
  AND2X1 U3825 ( .IN1(n3808), .IN2(n3809), .Q(n3807) );
  AND2X1 U3826 ( .IN1(n3810), .IN2(n3811), .Q(n3808) );
  INVX0 U3827 ( .INP(n3684), .ZN(n3811) );
  OR2X1 U3828 ( .IN1(n3572), .IN2(n3573), .Q(n3810) );
  INVX0 U3829 ( .INP(n902), .ZN(n3573) );
  OR2X1 U3830 ( .IN1(n1693), .IN2(n3812), .Q(n902) );
  INVX0 U3831 ( .INP(n3813), .ZN(n3572) );
  OR2X1 U3832 ( .IN1(n3814), .IN2(n3815), .Q(n3813) );
  OR2X1 U3833 ( .IN1(g713), .IN2(n3816), .Q(n3815) );
  OR2X1 U3834 ( .IN1(g704), .IN2(g695), .Q(n3816) );
  OR2X1 U3835 ( .IN1(n3817), .IN2(n3818), .Q(n3814) );
  OR2X1 U3836 ( .IN1(g686), .IN2(g722), .Q(n3818) );
  AND2X1 U3837 ( .IN1(n3685), .IN2(g736), .Q(n3806) );
  OR2X1 U3838 ( .IN1(n3819), .IN2(n3676), .Q(g8923) );
  AND2X1 U3839 ( .IN1(n3820), .IN2(n3678), .Q(n3819) );
  AND2X1 U3840 ( .IN1(n3821), .IN2(n3822), .Q(n3820) );
  INVX0 U3841 ( .INP(n3823), .ZN(n3822) );
  AND2X1 U3842 ( .IN1(n3824), .IN2(n1693), .Q(n3823) );
  OR2X1 U3843 ( .IN1(n1693), .IN2(n3824), .Q(n3821) );
  OR2X1 U3844 ( .IN1(n3825), .IN2(n3684), .Q(n3824) );
  AND2X1 U3845 ( .IN1(n3826), .IN2(n3827), .Q(n3825) );
  OR2X1 U3846 ( .IN1(g713), .IN2(n3828), .Q(n3827) );
  AND2X1 U3847 ( .IN1(n3829), .IN2(n3830), .Q(n3826) );
  OR2X1 U3848 ( .IN1(n3812), .IN2(n3685), .Q(n3830) );
  OR2X1 U3849 ( .IN1(n3831), .IN2(n3832), .Q(n3812) );
  OR2X1 U3850 ( .IN1(n3833), .IN2(n3834), .Q(n3832) );
  INVX0 U3851 ( .INP(n967), .ZN(n3834) );
  OR2X1 U3852 ( .IN1(n1676), .IN2(n3835), .Q(n3831) );
  OR2X1 U3853 ( .IN1(n3329), .IN2(n3275), .Q(n3835) );
  OR2X1 U3854 ( .IN1(n3225), .IN2(n3809), .Q(n3829) );
  OR2X1 U3855 ( .IN1(n3836), .IN2(n3676), .Q(g8922) );
  AND2X1 U3856 ( .IN1(n3837), .IN2(n3678), .Q(n3836) );
  AND2X1 U3857 ( .IN1(n3838), .IN2(n3839), .Q(n3837) );
  OR2X1 U3858 ( .IN1(n3840), .IN2(g668), .Q(n3839) );
  INVX0 U3859 ( .INP(n3841), .ZN(n3840) );
  OR2X1 U3860 ( .IN1(n1662), .IN2(n3841), .Q(n3838) );
  OR2X1 U3861 ( .IN1(n3684), .IN2(n3842), .Q(n3841) );
  OR2X1 U3862 ( .IN1(n3843), .IN2(n3844), .Q(n3842) );
  AND2X1 U3863 ( .IN1(n3845), .IN2(n3809), .Q(n3844) );
  OR2X1 U3864 ( .IN1(n3846), .IN2(n3847), .Q(n3845) );
  AND2X1 U3865 ( .IN1(n3848), .IN2(g658), .Q(n3847) );
  AND2X1 U3866 ( .IN1(n1615), .IN2(n3849), .Q(n3846) );
  AND2X1 U3867 ( .IN1(n3193), .IN2(n3685), .Q(n3843) );
  OR2X1 U3868 ( .IN1(n3850), .IN2(n3687), .Q(g8921) );
  AND2X1 U3869 ( .IN1(n3851), .IN2(n3852), .Q(n3687) );
  INVX0 U3870 ( .INP(n3853), .ZN(n3852) );
  OR2X1 U3871 ( .IN1(n3689), .IN2(n3854), .Q(n3853) );
  AND2X1 U3872 ( .IN1(n916), .IN2(n3625), .Q(n3851) );
  AND2X1 U3873 ( .IN1(n3855), .IN2(n3689), .Q(n3850) );
  AND2X1 U3874 ( .IN1(n3615), .IN2(n3625), .Q(n3689) );
  INVX0 U3875 ( .INP(n812), .ZN(n3615) );
  AND2X1 U3876 ( .IN1(n3856), .IN2(n3857), .Q(n3855) );
  OR2X1 U3877 ( .IN1(n3858), .IN2(g1872), .Q(n3857) );
  INVX0 U3878 ( .INP(n3859), .ZN(n3858) );
  OR2X1 U3879 ( .IN1(n1616), .IN2(n3859), .Q(n3856) );
  OR2X1 U3880 ( .IN1(n3860), .IN2(n3700), .Q(n3859) );
  AND2X1 U3881 ( .IN1(n918), .IN2(n3697), .Q(n3700) );
  INVX0 U3882 ( .INP(n3708), .ZN(n3697) );
  OR2X1 U3883 ( .IN1(n633), .IN2(n3861), .Q(n918) );
  AND2X1 U3884 ( .IN1(n3862), .IN2(n3616), .Q(n3861) );
  OR2X1 U3885 ( .IN1(g1840), .IN2(n3863), .Q(n3616) );
  OR2X1 U3886 ( .IN1(n1655), .IN2(n1608), .Q(n3863) );
  OR2X1 U3887 ( .IN1(n3864), .IN2(n1682), .Q(n3862) );
  AND2X1 U3888 ( .IN1(n1643), .IN2(n1605), .Q(n3864) );
  AND2X1 U3889 ( .IN1(n3337), .IN2(n3708), .Q(n3860) );
  OR2X1 U3890 ( .IN1(n3865), .IN2(n363), .Q(n3708) );
  AND2X1 U3891 ( .IN1(n926), .IN2(g1840), .Q(n3865) );
  OR2X1 U3892 ( .IN1(n3866), .IN2(n3676), .Q(g8920) );
  AND2X1 U3893 ( .IN1(n3867), .IN2(n3678), .Q(n3866) );
  AND2X1 U3894 ( .IN1(n3868), .IN2(n3869), .Q(n3867) );
  OR2X1 U3895 ( .IN1(n3870), .IN2(g713), .Q(n3869) );
  INVX0 U3896 ( .INP(n931), .ZN(n3870) );
  OR2X1 U3897 ( .IN1(n3348), .IN2(n931), .Q(n3868) );
  OR2X1 U3898 ( .IN1(n3871), .IN2(n3684), .Q(n931) );
  AND2X1 U3899 ( .IN1(n3872), .IN2(n3873), .Q(n3871) );
  OR2X1 U3900 ( .IN1(n3275), .IN2(n3874), .Q(n3873) );
  AND2X1 U3901 ( .IN1(n3875), .IN2(n3828), .Q(n3872) );
  OR2X1 U3902 ( .IN1(g704), .IN2(n3876), .Q(n3828) );
  OR2X1 U3903 ( .IN1(n3809), .IN2(n3175), .Q(n3875) );
  OR2X1 U3904 ( .IN1(n3877), .IN2(n3676), .Q(g8889) );
  AND2X1 U3905 ( .IN1(n3878), .IN2(n3678), .Q(n3877) );
  AND2X1 U3906 ( .IN1(n3879), .IN2(n3880), .Q(n3878) );
  OR2X1 U3907 ( .IN1(n78), .IN2(g704), .Q(n3880) );
  INVX0 U3908 ( .INP(n3881), .ZN(n78) );
  OR2X1 U3909 ( .IN1(n3275), .IN2(n3881), .Q(n3879) );
  OR2X1 U3910 ( .IN1(n3882), .IN2(n3684), .Q(n3881) );
  AND2X1 U3911 ( .IN1(n3883), .IN2(n3884), .Q(n3882) );
  OR2X1 U3912 ( .IN1(n3809), .IN2(n1719), .Q(n3884) );
  AND2X1 U3913 ( .IN1(n3874), .IN2(n3876), .Q(n3883) );
  OR2X1 U3914 ( .IN1(n3885), .IN2(n3886), .Q(n3876) );
  OR2X1 U3915 ( .IN1(g686), .IN2(g695), .Q(n3886) );
  OR2X1 U3916 ( .IN1(n3887), .IN2(n3888), .Q(n3874) );
  OR2X1 U3917 ( .IN1(n3329), .IN2(n1676), .Q(n3888) );
  OR2X1 U3918 ( .IN1(n3889), .IN2(n3676), .Q(g8887) );
  AND2X1 U3919 ( .IN1(n3890), .IN2(n3678), .Q(n3889) );
  AND2X1 U3920 ( .IN1(n3891), .IN2(n3892), .Q(n3890) );
  OR2X1 U3921 ( .IN1(n3893), .IN2(g695), .Q(n3892) );
  INVX0 U3922 ( .INP(n3894), .ZN(n3893) );
  OR2X1 U3923 ( .IN1(n3329), .IN2(n3894), .Q(n3891) );
  OR2X1 U3924 ( .IN1(n3895), .IN2(n3684), .Q(n3894) );
  AND2X1 U3925 ( .IN1(n3896), .IN2(n3897), .Q(n3895) );
  OR2X1 U3926 ( .IN1(n3809), .IN2(n3273), .Q(n3897) );
  AND2X1 U3927 ( .IN1(n3898), .IN2(n3899), .Q(n3896) );
  OR2X1 U3928 ( .IN1(n1676), .IN2(n3887), .Q(n3899) );
  OR2X1 U3929 ( .IN1(g686), .IN2(n3885), .Q(n3898) );
  OR2X1 U3930 ( .IN1(n3900), .IN2(n3676), .Q(g8885) );
  AND2X1 U3931 ( .IN1(n3901), .IN2(n3678), .Q(n3900) );
  AND2X1 U3932 ( .IN1(n3902), .IN2(n3903), .Q(n3901) );
  INVX0 U3933 ( .INP(n3904), .ZN(n3903) );
  AND2X1 U3934 ( .IN1(n3905), .IN2(n1676), .Q(n3904) );
  OR2X1 U3935 ( .IN1(n1676), .IN2(n3905), .Q(n3902) );
  OR2X1 U3936 ( .IN1(n3906), .IN2(n3684), .Q(n3905) );
  AND2X1 U3937 ( .IN1(n3907), .IN2(n3908), .Q(n3906) );
  AND2X1 U3938 ( .IN1(n3885), .IN2(n3887), .Q(n3908) );
  OR2X1 U3939 ( .IN1(n3685), .IN2(n3909), .Q(n3887) );
  OR2X1 U3940 ( .IN1(n1656), .IN2(n3833), .Q(n3909) );
  OR2X1 U3941 ( .IN1(n3685), .IN2(n3817), .Q(n3885) );
  OR2X1 U3942 ( .IN1(n3910), .IN2(g677), .Q(n3817) );
  OR2X1 U3943 ( .IN1(n3809), .IN2(n3341), .Q(n3907) );
  OR2X1 U3944 ( .IN1(n3911), .IN2(n3676), .Q(g8883) );
  INVX0 U3945 ( .INP(n3912), .ZN(n3676) );
  OR2X1 U3946 ( .IN1(n3913), .IN2(n3914), .Q(n3912) );
  OR2X1 U3947 ( .IN1(n3651), .IN2(n3578), .Q(n3914) );
  OR2X1 U3948 ( .IN1(n3678), .IN2(n3607), .Q(n3913) );
  AND2X1 U3949 ( .IN1(n3915), .IN2(n3678), .Q(n3911) );
  AND2X1 U3950 ( .IN1(n3916), .IN2(n3917), .Q(n3915) );
  OR2X1 U3951 ( .IN1(g677), .IN2(n3918), .Q(n3917) );
  INVX0 U3952 ( .INP(n3919), .ZN(n3918) );
  OR2X1 U3953 ( .IN1(n1656), .IN2(n3919), .Q(n3916) );
  AND2X1 U3954 ( .IN1(n3920), .IN2(n3921), .Q(n3919) );
  OR2X1 U3955 ( .IN1(n3922), .IN2(n3685), .Q(n3921) );
  INVX0 U3956 ( .INP(n3809), .ZN(n3685) );
  OR2X1 U3957 ( .IN1(n3923), .IN2(n3684), .Q(n3922) );
  AND2X1 U3958 ( .IN1(n958), .IN2(n3809), .Q(n3684) );
  OR2X1 U3959 ( .IN1(n3924), .IN2(n3925), .Q(n958) );
  AND2X1 U3960 ( .IN1(n3926), .IN2(n3661), .Q(n3924) );
  OR2X1 U3961 ( .IN1(n3927), .IN2(n1692), .Q(n3926) );
  AND2X1 U3962 ( .IN1(n1644), .IN2(n1593), .Q(n3927) );
  AND2X1 U3963 ( .IN1(n3833), .IN2(n3910), .Q(n3923) );
  OR2X1 U3964 ( .IN1(g668), .IN2(n3928), .Q(n3910) );
  OR2X1 U3965 ( .IN1(n3849), .IN2(g658), .Q(n3928) );
  OR2X1 U3966 ( .IN1(n3848), .IN2(n3929), .Q(n3833) );
  OR2X1 U3967 ( .IN1(n1662), .IN2(n1615), .Q(n3929) );
  INVX0 U3968 ( .INP(n3849), .ZN(n3848) );
  OR2X1 U3969 ( .IN1(n3930), .IN2(n3931), .Q(n3849) );
  AND2X1 U3970 ( .IN1(n3932), .IN2(n1593), .Q(n3931) );
  AND2X1 U3971 ( .IN1(n1644), .IN2(n3933), .Q(n3930) );
  OR2X1 U3972 ( .IN1(n3809), .IN2(n3344), .Q(n3920) );
  AND2X1 U3973 ( .IN1(n3934), .IN2(n3935), .Q(n3809) );
  OR2X1 U3974 ( .IN1(n3936), .IN2(n1607), .Q(n3934) );
  OR2X1 U3975 ( .IN1(n3937), .IN2(n3603), .Q(g8820) );
  AND2X1 U3976 ( .IN1(n1713), .IN2(n3938), .Q(n3603) );
  AND2X1 U3977 ( .IN1(n804), .IN2(n3607), .Q(n3938) );
  INVX0 U3978 ( .INP(n3661), .ZN(n3607) );
  AND2X1 U3979 ( .IN1(n3939), .IN2(g622), .Q(n3937) );
  OR2X1 U3980 ( .IN1(n3940), .IN2(n3678), .Q(n3939) );
  AND2X1 U3981 ( .IN1(n3608), .IN2(n3941), .Q(n3678) );
  INVX0 U3982 ( .INP(n804), .ZN(n3608) );
  AND2X1 U3983 ( .IN1(n3941), .IN2(n3661), .Q(n3940) );
  OR2X1 U3984 ( .IN1(n1609), .IN2(n3942), .Q(n3661) );
  OR2X1 U3985 ( .IN1(n3943), .IN2(n3944), .Q(g8779) );
  AND2X1 U3986 ( .IN1(n3945), .IN2(n3946), .Q(n3944) );
  AND2X1 U3987 ( .IN1(n495), .IN2(g1636), .Q(n3943) );
  OR2X1 U3988 ( .IN1(n3947), .IN2(n3948), .Q(g8777) );
  AND2X1 U3989 ( .IN1(n3949), .IN2(n3946), .Q(n3948) );
  AND2X1 U3990 ( .IN1(n495), .IN2(g1633), .Q(n3947) );
  OR2X1 U3991 ( .IN1(n3950), .IN2(n3951), .Q(g8776) );
  AND2X1 U3992 ( .IN1(n3952), .IN2(n3946), .Q(n3951) );
  AND2X1 U3993 ( .IN1(n495), .IN2(g1630), .Q(n3950) );
  AND2X1 U3994 ( .IN1(n3953), .IN2(g109), .Q(g8775) );
  OR2X1 U3995 ( .IN1(n3954), .IN2(n3955), .Q(n3953) );
  INVX0 U3996 ( .INP(n3956), .ZN(n3955) );
  OR2X1 U3997 ( .IN1(n3957), .IN2(n3308), .Q(n3956) );
  AND2X1 U3998 ( .IN1(n3308), .IN2(n3957), .Q(n3954) );
  OR2X1 U3999 ( .IN1(n3958), .IN2(n3959), .Q(g8774) );
  AND2X1 U4000 ( .IN1(n3957), .IN2(n3946), .Q(n3959) );
  OR2X1 U4001 ( .IN1(n3960), .IN2(n3961), .Q(n3957) );
  AND2X1 U4002 ( .IN1(n3962), .IN2(n3963), .Q(n3960) );
  AND2X1 U4003 ( .IN1(n3964), .IN2(n3965), .Q(n3962) );
  INVX0 U4004 ( .INP(n3966), .ZN(n3965) );
  AND2X1 U4005 ( .IN1(n3967), .IN2(n1706), .Q(n3966) );
  OR2X1 U4006 ( .IN1(n1706), .IN2(n3967), .Q(n3964) );
  OR2X1 U4007 ( .IN1(n3968), .IN2(n3969), .Q(n3967) );
  AND2X1 U4008 ( .IN1(n495), .IN2(g1627), .Q(n3958) );
  OR2X1 U4009 ( .IN1(n3970), .IN2(n3971), .Q(g8773) );
  AND2X1 U4010 ( .IN1(n3972), .IN2(n3946), .Q(n3971) );
  AND2X1 U4011 ( .IN1(n495), .IN2(g1624), .Q(n3970) );
  AND2X1 U4012 ( .IN1(n3973), .IN2(g109), .Q(g8772) );
  OR2X1 U4013 ( .IN1(n3974), .IN2(n3975), .Q(n3973) );
  INVX0 U4014 ( .INP(n3976), .ZN(n3975) );
  OR2X1 U4015 ( .IN1(n3952), .IN2(n3309), .Q(n3976) );
  AND2X1 U4016 ( .IN1(n3309), .IN2(n3952), .Q(n3974) );
  OR2X1 U4017 ( .IN1(n3977), .IN2(n3978), .Q(n3952) );
  AND2X1 U4018 ( .IN1(n3979), .IN2(n3963), .Q(n3977) );
  AND2X1 U4019 ( .IN1(n3980), .IN2(n3981), .Q(n3979) );
  OR2X1 U4020 ( .IN1(n3982), .IN2(g1137), .Q(n3981) );
  INVX0 U4021 ( .INP(n3983), .ZN(n3982) );
  OR2X1 U4022 ( .IN1(n1597), .IN2(n3983), .Q(n3980) );
  OR2X1 U4023 ( .IN1(n3984), .IN2(n3969), .Q(n3983) );
  OR2X1 U4024 ( .IN1(n1658), .IN2(n1614), .Q(n3969) );
  OR2X1 U4025 ( .IN1(n3985), .IN2(n3986), .Q(g8771) );
  AND2X1 U4026 ( .IN1(n3987), .IN2(n3946), .Q(n3986) );
  AND2X1 U4027 ( .IN1(n495), .IN2(g1621), .Q(n3985) );
  OR2X1 U4028 ( .IN1(n3988), .IN2(n3989), .Q(g8770) );
  AND2X1 U4029 ( .IN1(n3990), .IN2(n3946), .Q(n3989) );
  AND2X1 U4030 ( .IN1(n495), .IN2(g1615), .Q(n3988) );
  AND2X1 U4031 ( .IN1(n3991), .IN2(g109), .Q(g8769) );
  OR2X1 U4032 ( .IN1(n3992), .IN2(n3993), .Q(n3991) );
  INVX0 U4033 ( .INP(n3994), .ZN(n3993) );
  OR2X1 U4034 ( .IN1(n3990), .IN2(n3310), .Q(n3994) );
  AND2X1 U4035 ( .IN1(n3310), .IN2(n3990), .Q(n3992) );
  OR2X1 U4036 ( .IN1(n3995), .IN2(n3996), .Q(n3990) );
  AND2X1 U4037 ( .IN1(n3997), .IN2(n3963), .Q(n3995) );
  AND2X1 U4038 ( .IN1(n3998), .IN2(n3999), .Q(n3997) );
  INVX0 U4039 ( .INP(n4000), .ZN(n3999) );
  AND2X1 U4040 ( .IN1(n4001), .IN2(n1618), .Q(n4000) );
  OR2X1 U4041 ( .IN1(n1618), .IN2(n4001), .Q(n3998) );
  OR2X1 U4042 ( .IN1(n3984), .IN2(n4002), .Q(n4001) );
  AND2X1 U4043 ( .IN1(n4003), .IN2(g109), .Q(g8768) );
  OR2X1 U4044 ( .IN1(n4004), .IN2(n4005), .Q(n4003) );
  INVX0 U4045 ( .INP(n4006), .ZN(n4005) );
  OR2X1 U4046 ( .IN1(n3949), .IN2(n3311), .Q(n4006) );
  AND2X1 U4047 ( .IN1(n3311), .IN2(n3949), .Q(n4004) );
  OR2X1 U4048 ( .IN1(n4007), .IN2(n4008), .Q(n3949) );
  AND2X1 U4049 ( .IN1(n4009), .IN2(n3963), .Q(n4007) );
  AND2X1 U4050 ( .IN1(n4010), .IN2(n4011), .Q(n4009) );
  INVX0 U4051 ( .INP(n4012), .ZN(n4011) );
  AND2X1 U4052 ( .IN1(n4013), .IN2(n1660), .Q(n4012) );
  OR2X1 U4053 ( .IN1(n1660), .IN2(n4013), .Q(n4010) );
  OR2X1 U4054 ( .IN1(g1101), .IN2(n4014), .Q(n4013) );
  OR2X1 U4055 ( .IN1(n1677), .IN2(n4015), .Q(n4014) );
  AND2X1 U4056 ( .IN1(n4016), .IN2(g109), .Q(g8767) );
  OR2X1 U4057 ( .IN1(n4017), .IN2(n4018), .Q(n4016) );
  AND2X1 U4058 ( .IN1(n4019), .IN2(g1403), .Q(n4018) );
  INVX0 U4059 ( .INP(n3987), .ZN(n4019) );
  AND2X1 U4060 ( .IN1(n3252), .IN2(n3987), .Q(n4017) );
  OR2X1 U4061 ( .IN1(n4020), .IN2(n4021), .Q(n3987) );
  AND2X1 U4062 ( .IN1(n4022), .IN2(n3963), .Q(n4020) );
  AND2X1 U4063 ( .IN1(n4023), .IN2(n4024), .Q(n4022) );
  INVX0 U4064 ( .INP(n4025), .ZN(n4024) );
  AND2X1 U4065 ( .IN1(n4026), .IN2(n1708), .Q(n4025) );
  OR2X1 U4066 ( .IN1(n1708), .IN2(n4026), .Q(n4023) );
  OR2X1 U4067 ( .IN1(n3968), .IN2(n4027), .Q(n4026) );
  AND2X1 U4068 ( .IN1(n4028), .IN2(g109), .Q(g8766) );
  OR2X1 U4069 ( .IN1(n4029), .IN2(n4030), .Q(n4028) );
  AND2X1 U4070 ( .IN1(n4031), .IN2(g1448), .Q(n4030) );
  INVX0 U4071 ( .INP(n3945), .ZN(n4031) );
  AND2X1 U4072 ( .IN1(n3250), .IN2(n3945), .Q(n4029) );
  OR2X1 U4073 ( .IN1(n4032), .IN2(n4033), .Q(n3945) );
  AND2X1 U4074 ( .IN1(n4034), .IN2(n3963), .Q(n4032) );
  AND2X1 U4075 ( .IN1(n4035), .IN2(n4036), .Q(n4034) );
  INVX0 U4076 ( .INP(n4037), .ZN(n4036) );
  AND2X1 U4077 ( .IN1(n4038), .IN2(n1617), .Q(n4037) );
  OR2X1 U4078 ( .IN1(n1617), .IN2(n4038), .Q(n4035) );
  OR2X1 U4079 ( .IN1(n4015), .IN2(n4039), .Q(n4038) );
  OR2X1 U4080 ( .IN1(n1677), .IN2(n1654), .Q(n4039) );
  AND2X1 U4081 ( .IN1(n4040), .IN2(g109), .Q(g8765) );
  OR2X1 U4082 ( .IN1(n4041), .IN2(n4042), .Q(n4040) );
  INVX0 U4083 ( .INP(n4043), .ZN(n4042) );
  OR2X1 U4084 ( .IN1(n3972), .IN2(n3251), .Q(n4043) );
  AND2X1 U4085 ( .IN1(n3251), .IN2(n3972), .Q(n4041) );
  OR2X1 U4086 ( .IN1(n4044), .IN2(n4045), .Q(n3972) );
  AND2X1 U4087 ( .IN1(n4046), .IN2(n3963), .Q(n4044) );
  AND2X1 U4088 ( .IN1(n4047), .IN2(n4048), .Q(n4046) );
  INVX0 U4089 ( .INP(n4049), .ZN(n4048) );
  AND2X1 U4090 ( .IN1(n4050), .IN2(n1705), .Q(n4049) );
  OR2X1 U4091 ( .IN1(n1705), .IN2(n4050), .Q(n4047) );
  OR2X1 U4092 ( .IN1(n3984), .IN2(n4027), .Q(n4050) );
  OR2X1 U4093 ( .IN1(n1614), .IN2(g1104), .Q(n4027) );
  OR2X1 U4094 ( .IN1(n3651), .IN2(n4051), .Q(g8649) );
  OR2X1 U4095 ( .IN1(n4052), .IN2(n4053), .Q(n4051) );
  AND2X1 U4096 ( .IN1(n1016), .IN2(g664), .Q(n4053) );
  AND2X1 U4097 ( .IN1(n4054), .IN2(g736), .Q(n4052) );
  OR2X1 U4098 ( .IN1(n4055), .IN2(n4056), .Q(g8631) );
  AND2X1 U4099 ( .IN1(n4057), .IN2(n3941), .Q(n4056) );
  OR2X1 U4100 ( .IN1(n4058), .IN2(n4059), .Q(n4057) );
  AND2X1 U4101 ( .IN1(n4060), .IN2(g636), .Q(n4059) );
  OR2X1 U4102 ( .IN1(n3588), .IN2(n4061), .Q(n4060) );
  OR2X1 U4103 ( .IN1(n4062), .IN2(n4063), .Q(n4061) );
  AND2X1 U4104 ( .IN1(n4064), .IN2(n4065), .Q(n4063) );
  OR2X1 U4105 ( .IN1(n4066), .IN2(n4067), .Q(n4065) );
  OR2X1 U4106 ( .IN1(n4068), .IN2(n4069), .Q(n4067) );
  AND2X1 U4107 ( .IN1(n4070), .IN2(n1692), .Q(n4069) );
  AND2X1 U4108 ( .IN1(n1609), .IN2(n3658), .Q(n4070) );
  AND2X1 U4109 ( .IN1(n3662), .IN2(g639), .Q(n4068) );
  AND2X1 U4110 ( .IN1(g622), .IN2(g255), .Q(n4066) );
  OR2X1 U4111 ( .IN1(n4071), .IN2(n4072), .Q(n4064) );
  OR2X1 U4112 ( .IN1(n3334), .IN2(n1713), .Q(n4072) );
  OR2X1 U4113 ( .IN1(n4073), .IN2(n4074), .Q(n4071) );
  AND2X1 U4114 ( .IN1(n1692), .IN2(n4075), .Q(n4074) );
  OR2X1 U4115 ( .IN1(n4076), .IN2(g611), .Q(n4075) );
  AND2X1 U4116 ( .IN1(n3932), .IN2(g639), .Q(n4073) );
  AND2X1 U4117 ( .IN1(n4077), .IN2(n4078), .Q(n4062) );
  AND2X1 U4118 ( .IN1(n3658), .IN2(n3942), .Q(n4078) );
  AND2X1 U4119 ( .IN1(n1609), .IN2(n1644), .Q(n4077) );
  OR2X1 U4120 ( .IN1(n3379), .IN2(n1874), .Q(n3588) );
  AND2X1 U4121 ( .IN1(n4079), .IN2(n1713), .Q(n4058) );
  AND2X1 U4122 ( .IN1(n3651), .IN2(n4080), .Q(n4055) );
  OR2X1 U4123 ( .IN1(n4081), .IN2(n4082), .Q(n4080) );
  OR2X1 U4124 ( .IN1(n1716), .IN2(n4083), .Q(n4082) );
  AND2X1 U4125 ( .IN1(n4084), .IN2(n4085), .Q(n4083) );
  OR2X1 U4126 ( .IN1(n3326), .IN2(n3338), .Q(n4085) );
  OR2X1 U4127 ( .IN1(n3325), .IN2(n3335), .Q(n4084) );
  AND2X1 U4128 ( .IN1(n4086), .IN2(n4087), .Q(n4081) );
  OR2X1 U4129 ( .IN1(n1622), .IN2(n3339), .Q(n4086) );
  OR2X1 U4130 ( .IN1(n4088), .IN2(n4089), .Q(g8566) );
  AND2X1 U4131 ( .IN1(g1690), .IN2(g1687), .Q(n4089) );
  AND2X1 U4132 ( .IN1(n1653), .IN2(g1669), .Q(n4088) );
  OR2X1 U4133 ( .IN1(n4090), .IN2(n4091), .Q(g8565) );
  AND2X1 U4134 ( .IN1(g1690), .IN2(g1684), .Q(n4091) );
  AND2X1 U4135 ( .IN1(n1653), .IN2(g1666), .Q(n4090) );
  OR2X1 U4136 ( .IN1(n4092), .IN2(n4093), .Q(g8564) );
  AND2X1 U4137 ( .IN1(g1690), .IN2(g1681), .Q(n4093) );
  AND2X1 U4138 ( .IN1(n1653), .IN2(g1663), .Q(n4092) );
  OR2X1 U4139 ( .IN1(n4094), .IN2(n4095), .Q(g8563) );
  AND2X1 U4140 ( .IN1(g1690), .IN2(g1678), .Q(n4095) );
  AND2X1 U4141 ( .IN1(n1653), .IN2(g1660), .Q(n4094) );
  OR2X1 U4142 ( .IN1(n4096), .IN2(n4097), .Q(g8562) );
  AND2X1 U4143 ( .IN1(g1690), .IN2(g1675), .Q(n4097) );
  AND2X1 U4144 ( .IN1(n1653), .IN2(g1657), .Q(n4096) );
  OR2X1 U4145 ( .IN1(n4098), .IN2(n4099), .Q(g8561) );
  AND2X1 U4146 ( .IN1(g1690), .IN2(g1672), .Q(n4099) );
  AND2X1 U4147 ( .IN1(n1653), .IN2(g1654), .Q(n4098) );
  OR2X1 U4148 ( .IN1(n4100), .IN2(n4101), .Q(g8559) );
  OR2X1 U4149 ( .IN1(n4102), .IN2(n4103), .Q(n4101) );
  AND2X1 U4150 ( .IN1(n4104), .IN2(g1878), .Q(n4103) );
  AND2X1 U4151 ( .IN1(g18), .IN2(n4105), .Q(g8505) );
  OR2X1 U4152 ( .IN1(n4106), .IN2(n4107), .Q(n4105) );
  AND2X1 U4153 ( .IN1(n4108), .IN2(g617), .Q(n4107) );
  AND2X1 U4154 ( .IN1(n1645), .IN2(n4109), .Q(n4106) );
  INVX0 U4155 ( .INP(n4108), .ZN(n4109) );
  AND2X1 U4156 ( .IN1(n4110), .IN2(n4111), .Q(n4108) );
  OR2X1 U4157 ( .IN1(n1016), .IN2(n3287), .Q(n4111) );
  OR2X1 U4158 ( .IN1(n3936), .IN2(n3942), .Q(n4110) );
  OR2X1 U4159 ( .IN1(n1607), .IN2(g617), .Q(n3942) );
  OR2X1 U4160 ( .IN1(n4112), .IN2(n4113), .Q(n3936) );
  OR2X1 U4161 ( .IN1(n3925), .IN2(g611), .Q(n4113) );
  OR2X1 U4162 ( .IN1(g605), .IN2(g599), .Q(n4112) );
  OR2X1 U4163 ( .IN1(n4114), .IN2(n4115), .Q(g8435) );
  AND2X1 U4164 ( .IN1(n4054), .IN2(g727), .Q(n4115) );
  AND2X1 U4165 ( .IN1(n4116), .IN2(g736), .Q(n4114) );
  OR2X1 U4166 ( .IN1(n4117), .IN2(n4118), .Q(g8434) );
  AND2X1 U4167 ( .IN1(n4054), .IN2(g718), .Q(n4118) );
  AND2X1 U4168 ( .IN1(n4116), .IN2(g727), .Q(n4117) );
  OR2X1 U4169 ( .IN1(n4119), .IN2(n4120), .Q(g8433) );
  AND2X1 U4170 ( .IN1(n4054), .IN2(g709), .Q(n4120) );
  AND2X1 U4171 ( .IN1(n4116), .IN2(g718), .Q(n4119) );
  OR2X1 U4172 ( .IN1(n4121), .IN2(n4122), .Q(g8432) );
  AND2X1 U4173 ( .IN1(n4054), .IN2(g700), .Q(n4122) );
  AND2X1 U4174 ( .IN1(n4116), .IN2(g709), .Q(n4121) );
  OR2X1 U4175 ( .IN1(n4123), .IN2(n4124), .Q(g8431) );
  AND2X1 U4176 ( .IN1(n4054), .IN2(g691), .Q(n4124) );
  AND2X1 U4177 ( .IN1(n4116), .IN2(g700), .Q(n4123) );
  OR2X1 U4178 ( .IN1(n4125), .IN2(n4126), .Q(g8430) );
  AND2X1 U4179 ( .IN1(n4054), .IN2(g682), .Q(n4126) );
  AND2X1 U4180 ( .IN1(n4116), .IN2(g691), .Q(n4125) );
  OR2X1 U4181 ( .IN1(n4127), .IN2(n4128), .Q(g8429) );
  AND2X1 U4182 ( .IN1(n4054), .IN2(g673), .Q(n4128) );
  AND2X1 U4183 ( .IN1(n4116), .IN2(g682), .Q(n4127) );
  OR2X1 U4184 ( .IN1(n4129), .IN2(n4130), .Q(g8428) );
  AND2X1 U4185 ( .IN1(n4054), .IN2(g664), .Q(n4130) );
  INVX0 U4186 ( .INP(n1016), .ZN(n4054) );
  AND2X1 U4187 ( .IN1(n4116), .IN2(g673), .Q(n4129) );
  AND2X1 U4188 ( .IN1(n3941), .IN2(n1016), .Q(n4116) );
  OR2X1 U4189 ( .IN1(g611), .IN2(n3935), .Q(n1016) );
  OR2X1 U4190 ( .IN1(n1645), .IN2(n3925), .Q(n3935) );
  AND2X1 U4191 ( .IN1(g18), .IN2(n4131), .Q(g8384) );
  OR2X1 U4192 ( .IN1(n4132), .IN2(n4133), .Q(n4131) );
  AND2X1 U4193 ( .IN1(n4134), .IN2(g1840), .Q(n4133) );
  INVX0 U4194 ( .INP(n4135), .ZN(n4134) );
  AND2X1 U4195 ( .IN1(n3288), .IN2(n4135), .Q(n4132) );
  OR2X1 U4196 ( .IN1(n4102), .IN2(n363), .Q(n4135) );
  INVX0 U4197 ( .INP(n4136), .ZN(n363) );
  OR2X1 U4198 ( .IN1(n4137), .IN2(n4138), .Q(n4136) );
  OR2X1 U4199 ( .IN1(n633), .IN2(g1822), .Q(n4138) );
  AND2X1 U4200 ( .IN1(n4139), .IN2(g1950), .Q(n4102) );
  OR2X1 U4201 ( .IN1(g82), .IN2(g8986), .Q(g8352) );
  OR2X1 U4202 ( .IN1(g82), .IN2(g8985), .Q(g8349) );
  OR2X1 U4203 ( .IN1(g82), .IN2(g8976), .Q(g8347) );
  OR2X1 U4204 ( .IN1(g82), .IN2(test_so10), .Q(g8340) );
  OR2X1 U4205 ( .IN1(g82), .IN2(g8983), .Q(g8335) );
  OR2X1 U4206 ( .IN1(g82), .IN2(g8982), .Q(g8331) );
  OR2X1 U4207 ( .IN1(g82), .IN2(g8981), .Q(g8328) );
  OR2X1 U4208 ( .IN1(g82), .IN2(g8980), .Q(g8323) );
  OR2X1 U4209 ( .IN1(g82), .IN2(g8979), .Q(g8318) );
  OR2X1 U4210 ( .IN1(g82), .IN2(g8978), .Q(g8316) );
  OR2X1 U4211 ( .IN1(g82), .IN2(g8977), .Q(g8313) );
  OR2X1 U4212 ( .IN1(n4140), .IN2(n4141), .Q(g8288) );
  AND2X1 U4213 ( .IN1(n4139), .IN2(g1941), .Q(n4141) );
  AND2X1 U4214 ( .IN1(n4142), .IN2(g1950), .Q(n4140) );
  OR2X1 U4215 ( .IN1(n4143), .IN2(n4144), .Q(g8287) );
  AND2X1 U4216 ( .IN1(n4139), .IN2(g1932), .Q(n4144) );
  AND2X1 U4217 ( .IN1(n4142), .IN2(g1941), .Q(n4143) );
  OR2X1 U4218 ( .IN1(n4145), .IN2(n4146), .Q(g8286) );
  AND2X1 U4219 ( .IN1(n4139), .IN2(g1923), .Q(n4146) );
  AND2X1 U4220 ( .IN1(n4142), .IN2(g1932), .Q(n4145) );
  OR2X1 U4221 ( .IN1(n4147), .IN2(n4148), .Q(g8285) );
  AND2X1 U4222 ( .IN1(n4139), .IN2(g1914), .Q(n4148) );
  AND2X1 U4223 ( .IN1(n4142), .IN2(g1923), .Q(n4147) );
  OR2X1 U4224 ( .IN1(n4149), .IN2(n4150), .Q(g8284) );
  AND2X1 U4225 ( .IN1(n4139), .IN2(g1905), .Q(n4150) );
  AND2X1 U4226 ( .IN1(n4142), .IN2(g1914), .Q(n4149) );
  OR2X1 U4227 ( .IN1(n4151), .IN2(n4152), .Q(g8283) );
  AND2X1 U4228 ( .IN1(n4139), .IN2(g1896), .Q(n4152) );
  AND2X1 U4229 ( .IN1(n4142), .IN2(g1905), .Q(n4151) );
  OR2X1 U4230 ( .IN1(n4153), .IN2(n4154), .Q(g8282) );
  AND2X1 U4231 ( .IN1(n4139), .IN2(g1887), .Q(n4154) );
  AND2X1 U4232 ( .IN1(n4142), .IN2(g1896), .Q(n4153) );
  OR2X1 U4233 ( .IN1(n4155), .IN2(n4156), .Q(g8281) );
  AND2X1 U4234 ( .IN1(n4139), .IN2(g1878), .Q(n4156) );
  INVX0 U4235 ( .INP(n4104), .ZN(n4139) );
  AND2X1 U4236 ( .IN1(n4142), .IN2(g1887), .Q(n4155) );
  AND2X1 U4237 ( .IN1(n3625), .IN2(n4104), .Q(n4142) );
  OR2X1 U4238 ( .IN1(g1834), .IN2(n4157), .Q(n4104) );
  OR2X1 U4239 ( .IN1(n3288), .IN2(n633), .Q(n4157) );
  INVX0 U4240 ( .INP(n926), .ZN(n633) );
  AND2X1 U4241 ( .IN1(n4158), .IN2(g940), .Q(g8260) );
  AND2X1 U4242 ( .IN1(n4158), .IN2(g936), .Q(g8254) );
  AND2X1 U4243 ( .IN1(n4158), .IN2(g932), .Q(g8250) );
  AND2X1 U4244 ( .IN1(n4159), .IN2(n4160), .Q(g8245) );
  AND2X1 U4245 ( .IN1(n4161), .IN2(n4162), .Q(n4159) );
  INVX0 U4246 ( .INP(n4163), .ZN(n4162) );
  AND2X1 U4247 ( .IN1(n4164), .IN2(n1716), .Q(n4163) );
  OR2X1 U4248 ( .IN1(n1716), .IN2(n4164), .Q(n4161) );
  AND2X1 U4249 ( .IN1(n4165), .IN2(n4166), .Q(g8244) );
  AND2X1 U4250 ( .IN1(n4167), .IN2(n4168), .Q(n4165) );
  OR2X1 U4251 ( .IN1(n4169), .IN2(g4181), .Q(n4167) );
  AND2X1 U4252 ( .IN1(n1093), .IN2(g4180), .Q(n4169) );
  OR2X1 U4253 ( .IN1(n4170), .IN2(n4171), .Q(g8194) );
  AND2X1 U4254 ( .IN1(n4172), .IN2(n3946), .Q(n4171) );
  AND2X1 U4255 ( .IN1(n4173), .IN2(n4174), .Q(n4172) );
  INVX0 U4256 ( .INP(n4175), .ZN(n4174) );
  AND2X1 U4257 ( .IN1(n4176), .IN2(n6001), .Q(n4175) );
  OR2X1 U4258 ( .IN1(n6001), .IN2(n4176), .Q(n4173) );
  OR2X1 U4259 ( .IN1(n4002), .IN2(n4177), .Q(n4176) );
  OR2X1 U4260 ( .IN1(n1677), .IN2(g1101), .Q(n4177) );
  AND2X1 U4261 ( .IN1(n495), .IN2(g1512), .Q(n4170) );
  OR2X1 U4262 ( .IN1(n4178), .IN2(n4179), .Q(g8193) );
  AND2X1 U4263 ( .IN1(n4180), .IN2(n3946), .Q(n4179) );
  OR2X1 U4264 ( .IN1(n4181), .IN2(n4182), .Q(n4180) );
  AND2X1 U4265 ( .IN1(n4183), .IN2(n3387), .Q(n4182) );
  INVX0 U4266 ( .INP(n4184), .ZN(n4183) );
  AND2X1 U4267 ( .IN1(test_so4), .IN2(n4184), .Q(n4181) );
  OR2X1 U4268 ( .IN1(n3968), .IN2(n4002), .Q(n4184) );
  OR2X1 U4269 ( .IN1(n1658), .IN2(g1107), .Q(n4002) );
  OR2X1 U4270 ( .IN1(g1110), .IN2(g1101), .Q(n3968) );
  AND2X1 U4271 ( .IN1(n495), .IN2(g1639), .Q(n4178) );
  AND2X1 U4272 ( .IN1(n1610), .IN2(n4185), .Q(g8173) );
  OR2X1 U4273 ( .IN1(n4186), .IN2(n4187), .Q(n4185) );
  AND2X1 U4274 ( .IN1(n4188), .IN2(g1806), .Q(n4187) );
  OR2X1 U4275 ( .IN1(n493), .IN2(n1055), .Q(n4188) );
  AND2X1 U4276 ( .IN1(n4189), .IN2(n1056), .Q(n4186) );
  AND2X1 U4277 ( .IN1(n1055), .IN2(g1801), .Q(n4189) );
  OR2X1 U4278 ( .IN1(n3589), .IN2(n4190), .Q(n1055) );
  OR2X1 U4279 ( .IN1(n3320), .IN2(n3319), .Q(n4190) );
  OR2X1 U4280 ( .IN1(n1626), .IN2(n4191), .Q(n3589) );
  AND2X1 U4281 ( .IN1(n4158), .IN2(g928), .Q(g8147) );
  AND2X1 U4282 ( .IN1(g109), .IN2(n4192), .Q(n4158) );
  OR2X1 U4283 ( .IN1(n4193), .IN2(n4194), .Q(n4192) );
  OR2X1 U4284 ( .IN1(g881), .IN2(n3027), .Q(n4193) );
  AND2X1 U4285 ( .IN1(n4195), .IN2(g109), .Q(g8060) );
  OR2X1 U4286 ( .IN1(n4196), .IN2(n4197), .Q(n4195) );
  AND2X1 U4287 ( .IN1(n4198), .IN2(g162), .Q(n4197) );
  INVX0 U4288 ( .INP(g6002), .ZN(n4198) );
  AND2X1 U4289 ( .IN1(n3246), .IN2(g6002), .Q(n4196) );
  AND2X1 U4290 ( .IN1(n4199), .IN2(g109), .Q(g8059) );
  AND2X1 U4291 ( .IN1(n4200), .IN2(n4201), .Q(n4199) );
  OR2X1 U4292 ( .IN1(g135), .IN2(g6042), .Q(n4201) );
  OR2X1 U4293 ( .IN1(n3243), .IN2(n4202), .Q(n4200) );
  INVX0 U4294 ( .INP(g6042), .ZN(n4202) );
  AND2X1 U4295 ( .IN1(n4203), .IN2(g109), .Q(g8055) );
  OR2X1 U4296 ( .IN1(n4204), .IN2(n4205), .Q(n4203) );
  INVX0 U4297 ( .INP(n4206), .ZN(n4205) );
  OR2X1 U4298 ( .IN1(n4207), .IN2(n3312), .Q(n4206) );
  AND2X1 U4299 ( .IN1(n3312), .IN2(n4207), .Q(n4204) );
  AND2X1 U4300 ( .IN1(n4208), .IN2(g109), .Q(g8054) );
  OR2X1 U4301 ( .IN1(n4209), .IN2(n4210), .Q(n4208) );
  INVX0 U4302 ( .INP(n4211), .ZN(n4210) );
  OR2X1 U4303 ( .IN1(g6015), .IN2(n3321), .Q(n4211) );
  AND2X1 U4304 ( .IN1(n3321), .IN2(g6015), .Q(n4209) );
  AND2X1 U4305 ( .IN1(n4212), .IN2(g109), .Q(g8053) );
  AND2X1 U4306 ( .IN1(n4213), .IN2(n4214), .Q(n4212) );
  OR2X1 U4307 ( .IN1(g139), .IN2(g6045), .Q(n4214) );
  OR2X1 U4308 ( .IN1(n3242), .IN2(n4215), .Q(n4213) );
  INVX0 U4309 ( .INP(g6045), .ZN(n4215) );
  AND2X1 U4310 ( .IN1(n4216), .IN2(g109), .Q(g8052) );
  OR2X1 U4311 ( .IN1(n4217), .IN2(n4218), .Q(n4216) );
  AND2X1 U4312 ( .IN1(n4219), .IN2(g1486), .Q(n4218) );
  INVX0 U4313 ( .INP(n4220), .ZN(n4219) );
  AND2X1 U4314 ( .IN1(n3244), .IN2(n4220), .Q(n4217) );
  AND2X1 U4315 ( .IN1(n4221), .IN2(g109), .Q(g8051) );
  AND2X1 U4316 ( .IN1(n4222), .IN2(n4223), .Q(n4221) );
  OR2X1 U4317 ( .IN1(g1466), .IN2(n4224), .Q(n4223) );
  OR2X1 U4318 ( .IN1(n3248), .IN2(n4225), .Q(n4222) );
  INVX0 U4319 ( .INP(n4224), .ZN(n4225) );
  AND2X1 U4320 ( .IN1(n4226), .IN2(g109), .Q(g8050) );
  OR2X1 U4321 ( .IN1(n4227), .IN2(n4228), .Q(n4226) );
  INVX0 U4322 ( .INP(n4229), .ZN(n4228) );
  OR2X1 U4323 ( .IN1(g6026), .IN2(n3322), .Q(n4229) );
  AND2X1 U4324 ( .IN1(n3322), .IN2(g6026), .Q(n4227) );
  AND2X1 U4325 ( .IN1(n4230), .IN2(g109), .Q(g8049) );
  AND2X1 U4326 ( .IN1(n4231), .IN2(n4232), .Q(n4230) );
  OR2X1 U4327 ( .IN1(g166), .IN2(g6049), .Q(n4232) );
  OR2X1 U4328 ( .IN1(n3245), .IN2(n4233), .Q(n4231) );
  INVX0 U4329 ( .INP(g6049), .ZN(n4233) );
  AND2X1 U4330 ( .IN1(n4234), .IN2(g109), .Q(g8048) );
  OR2X1 U4331 ( .IN1(n4235), .IN2(n4236), .Q(n4234) );
  AND2X1 U4332 ( .IN1(n4237), .IN2(g153), .Q(n4236) );
  INVX0 U4333 ( .INP(g5996), .ZN(n4237) );
  AND2X1 U4334 ( .IN1(n3268), .IN2(g5996), .Q(n4235) );
  AND2X1 U4335 ( .IN1(n4238), .IN2(g109), .Q(g8047) );
  OR2X1 U4336 ( .IN1(n4239), .IN2(n4240), .Q(n4238) );
  AND2X1 U4337 ( .IN1(n4241), .IN2(g127), .Q(n4240) );
  INVX0 U4338 ( .INP(g6035), .ZN(n4241) );
  AND2X1 U4339 ( .IN1(n1704), .IN2(g6035), .Q(n4239) );
  AND2X1 U4340 ( .IN1(n4242), .IN2(g109), .Q(g8046) );
  OR2X1 U4341 ( .IN1(n4243), .IN2(n4244), .Q(n4242) );
  AND2X1 U4342 ( .IN1(n4245), .IN2(g1482), .Q(n4244) );
  INVX0 U4343 ( .INP(n4246), .ZN(n4245) );
  AND2X1 U4344 ( .IN1(n3249), .IN2(n4246), .Q(n4243) );
  AND2X1 U4345 ( .IN1(n4247), .IN2(g109), .Q(g8045) );
  AND2X1 U4346 ( .IN1(n4248), .IN2(n4249), .Q(n4247) );
  OR2X1 U4347 ( .IN1(g1462), .IN2(n4250), .Q(n4249) );
  OR2X1 U4348 ( .IN1(n3313), .IN2(n4251), .Q(n4248) );
  INVX0 U4349 ( .INP(n4250), .ZN(n4251) );
  AND2X1 U4350 ( .IN1(n4252), .IN2(g109), .Q(g8044) );
  OR2X1 U4351 ( .IN1(n4253), .IN2(n4254), .Q(n4252) );
  AND2X1 U4352 ( .IN1(n4255), .IN2(g131), .Q(n4254) );
  INVX0 U4353 ( .INP(g6038), .ZN(n4255) );
  AND2X1 U4354 ( .IN1(n3241), .IN2(g6038), .Q(n4253) );
  AND2X1 U4355 ( .IN1(n4256), .IN2(g109), .Q(g8043) );
  OR2X1 U4356 ( .IN1(n4257), .IN2(n4258), .Q(n4256) );
  INVX0 U4357 ( .INP(n4259), .ZN(n4258) );
  OR2X1 U4358 ( .IN1(n4260), .IN2(n3314), .Q(n4259) );
  AND2X1 U4359 ( .IN1(n3314), .IN2(n4260), .Q(n4257) );
  AND2X1 U4360 ( .IN1(n4261), .IN2(g109), .Q(g8042) );
  AND2X1 U4361 ( .IN1(n4262), .IN2(n4263), .Q(n4261) );
  OR2X1 U4362 ( .IN1(g1458), .IN2(n4264), .Q(n4263) );
  OR2X1 U4363 ( .IN1(n1703), .IN2(n4265), .Q(n4262) );
  INVX0 U4364 ( .INP(n4264), .ZN(n4265) );
  AND2X1 U4365 ( .IN1(n4266), .IN2(g109), .Q(g8041) );
  OR2X1 U4366 ( .IN1(n4267), .IN2(n4268), .Q(n4266) );
  AND2X1 U4367 ( .IN1(n4269), .IN2(g1494), .Q(n4268) );
  AND2X1 U4368 ( .IN1(n3280), .IN2(n4270), .Q(n4267) );
  AND2X1 U4369 ( .IN1(n4271), .IN2(g109), .Q(g8040) );
  OR2X1 U4370 ( .IN1(n4272), .IN2(n4273), .Q(n4271) );
  AND2X1 U4371 ( .IN1(n4274), .IN2(g1474), .Q(n4273) );
  AND2X1 U4372 ( .IN1(n3281), .IN2(n4275), .Q(n4272) );
  AND2X1 U4373 ( .IN1(n4276), .IN2(g109), .Q(g8039) );
  OR2X1 U4374 ( .IN1(n4277), .IN2(n4278), .Q(n4276) );
  INVX0 U4375 ( .INP(n4279), .ZN(n4278) );
  OR2X1 U4376 ( .IN1(n4280), .IN2(n3282), .Q(n4279) );
  AND2X1 U4377 ( .IN1(n3282), .IN2(n4280), .Q(n4277) );
  AND2X1 U4378 ( .IN1(n4281), .IN2(n4160), .Q(g8024) );
  AND2X1 U4379 ( .IN1(n4164), .IN2(n4282), .Q(n4281) );
  OR2X1 U4380 ( .IN1(n1090), .IN2(g822), .Q(n4282) );
  OR2X1 U4381 ( .IN1(n3335), .IN2(n4283), .Q(n4164) );
  INVX0 U4382 ( .INP(n1090), .ZN(n4283) );
  AND2X1 U4383 ( .IN1(n4284), .IN2(n4166), .Q(g8019) );
  AND2X1 U4384 ( .IN1(n4285), .IN2(n4286), .Q(n4284) );
  OR2X1 U4385 ( .IN1(n1093), .IN2(g4180), .Q(n4286) );
  OR2X1 U4386 ( .IN1(n3363), .IN2(n4287), .Q(n4285) );
  AND2X1 U4387 ( .IN1(n4288), .IN2(n1610), .Q(g7930) );
  AND2X1 U4388 ( .IN1(n4289), .IN2(n4290), .Q(n4288) );
  OR2X1 U4389 ( .IN1(n1056), .IN2(g1801), .Q(n4290) );
  OR2X1 U4390 ( .IN1(n3319), .IN2(n4291), .Q(n4289) );
  AND2X1 U4391 ( .IN1(n4292), .IN2(g109), .Q(g7843) );
  OR2X1 U4392 ( .IN1(n4293), .IN2(n4294), .Q(n4292) );
  AND2X1 U4393 ( .IN1(n4295), .IN2(g158), .Q(n4294) );
  INVX0 U4394 ( .INP(g6000), .ZN(n4295) );
  AND2X1 U4395 ( .IN1(n3247), .IN2(g6000), .Q(n4293) );
  INVX0 U4396 ( .INP(n4296), .ZN(g7709) );
  OR2X1 U4397 ( .IN1(n4297), .IN2(n4298), .Q(n4296) );
  OR2X1 U4398 ( .IN1(n1090), .IN2(n1096), .Q(n4297) );
  AND2X1 U4399 ( .IN1(n4299), .IN2(n4166), .Q(g7705) );
  AND2X1 U4400 ( .IN1(n4287), .IN2(n4300), .Q(n4299) );
  INVX0 U4401 ( .INP(n1098), .ZN(n4300) );
  OR2X1 U4402 ( .IN1(n4301), .IN2(n4302), .Q(g7660) );
  OR2X1 U4403 ( .IN1(n3604), .IN2(n3651), .Q(n4302) );
  INVX0 U4404 ( .INP(n4303), .ZN(n4301) );
  OR2X1 U4405 ( .IN1(n4304), .IN2(n3315), .Q(n4303) );
  AND2X1 U4406 ( .IN1(n4305), .IN2(n4306), .Q(g7632) );
  INVX0 U4407 ( .INP(n4307), .ZN(n4305) );
  OR2X1 U4408 ( .IN1(n4308), .IN2(n4309), .Q(n4307) );
  AND2X1 U4409 ( .IN1(n4310), .IN2(n3367), .Q(n4308) );
  OR2X1 U4410 ( .IN1(n3651), .IN2(n4311), .Q(g7626) );
  OR2X1 U4411 ( .IN1(n4312), .IN2(n4313), .Q(n4311) );
  AND2X1 U4412 ( .IN1(n4314), .IN2(n1692), .Q(n4313) );
  AND2X1 U4413 ( .IN1(n3604), .IN2(n4315), .Q(n4314) );
  OR2X1 U4414 ( .IN1(n3578), .IN2(n4316), .Q(n4315) );
  OR2X1 U4415 ( .IN1(n3932), .IN2(n4076), .Q(n4316) );
  INVX0 U4416 ( .INP(n3658), .ZN(n4076) );
  OR2X1 U4417 ( .IN1(n1593), .IN2(n1607), .Q(n3658) );
  INVX0 U4418 ( .INP(n3662), .ZN(n3932) );
  OR2X1 U4419 ( .IN1(n1644), .IN2(g591), .Q(n3662) );
  OR2X1 U4420 ( .IN1(n4317), .IN2(n4079), .Q(n3578) );
  INVX0 U4421 ( .INP(n3657), .ZN(n4079) );
  OR2X1 U4422 ( .IN1(g599), .IN2(n4318), .Q(n3657) );
  OR2X1 U4423 ( .IN1(n1593), .IN2(g591), .Q(n4318) );
  AND2X1 U4424 ( .IN1(n1593), .IN2(g599), .Q(n4317) );
  AND2X1 U4425 ( .IN1(n3925), .IN2(g639), .Q(n4312) );
  AND2X1 U4426 ( .IN1(n4306), .IN2(n4319), .Q(g7590) );
  INVX0 U4427 ( .INP(n4320), .ZN(n4319) );
  AND2X1 U4428 ( .IN1(n4321), .IN2(n3361), .Q(n4320) );
  AND2X1 U4429 ( .IN1(n4306), .IN2(n4322), .Q(g7586) );
  OR2X1 U4430 ( .IN1(n4323), .IN2(n1107), .Q(n4322) );
  AND2X1 U4431 ( .IN1(n4309), .IN2(n4324), .Q(n1107) );
  AND2X1 U4432 ( .IN1(g1223), .IN2(n4325), .Q(n4324) );
  AND2X1 U4433 ( .IN1(n4321), .IN2(g1227), .Q(n4323) );
  OR2X1 U4434 ( .IN1(n4310), .IN2(n4326), .Q(n4321) );
  OR2X1 U4435 ( .IN1(n4327), .IN2(n4325), .Q(n4326) );
  AND2X1 U4436 ( .IN1(n4328), .IN2(n4306), .Q(g7581) );
  AND2X1 U4437 ( .IN1(n4329), .IN2(n4330), .Q(n4328) );
  OR2X1 U4438 ( .IN1(n4309), .IN2(g1223), .Q(n4330) );
  INVX0 U4439 ( .INP(n4331), .ZN(n4309) );
  OR2X1 U4440 ( .IN1(n3130), .IN2(n4331), .Q(n4329) );
  OR2X1 U4441 ( .IN1(n4310), .IN2(n4332), .Q(n4331) );
  OR2X1 U4442 ( .IN1(n3367), .IN2(n4327), .Q(n4332) );
  AND2X1 U4443 ( .IN1(n4333), .IN2(n1610), .Q(g7541) );
  AND2X1 U4444 ( .IN1(n4334), .IN2(n4335), .Q(n4333) );
  OR2X1 U4445 ( .IN1(n1626), .IN2(n4291), .Q(n4335) );
  INVX0 U4446 ( .INP(n1056), .ZN(n4291) );
  OR2X1 U4447 ( .IN1(n179), .IN2(g1796), .Q(n4334) );
  INVX0 U4448 ( .INP(n4336), .ZN(n179) );
  OR2X1 U4449 ( .IN1(n4337), .IN2(n4338), .Q(g7441) );
  OR2X1 U4450 ( .IN1(n4339), .IN2(n3651), .Q(n4338) );
  AND2X1 U4451 ( .IN1(n1701), .IN2(g643), .Q(n4337) );
  OR2X1 U4452 ( .IN1(n4340), .IN2(n4341), .Q(g7303) );
  AND2X1 U4453 ( .IN1(n4342), .IN2(g1265), .Q(n4341) );
  AND2X1 U4454 ( .IN1(n4343), .IN2(test_so6), .Q(n4340) );
  OR2X1 U4455 ( .IN1(n4344), .IN2(n4345), .Q(g7302) );
  AND2X1 U4456 ( .IN1(n4342), .IN2(g1260), .Q(n4345) );
  AND2X1 U4457 ( .IN1(n4343), .IN2(g1265), .Q(n4344) );
  OR2X1 U4458 ( .IN1(n4346), .IN2(n4347), .Q(g7301) );
  AND2X1 U4459 ( .IN1(n4342), .IN2(g1255), .Q(n4347) );
  AND2X1 U4460 ( .IN1(n4343), .IN2(g1260), .Q(n4346) );
  OR2X1 U4461 ( .IN1(n4348), .IN2(n4349), .Q(g7300) );
  AND2X1 U4462 ( .IN1(n4342), .IN2(g1250), .Q(n4349) );
  AND2X1 U4463 ( .IN1(n4343), .IN2(g1255), .Q(n4348) );
  OR2X1 U4464 ( .IN1(n4350), .IN2(n4351), .Q(g7299) );
  AND2X1 U4465 ( .IN1(n4342), .IN2(g1245), .Q(n4351) );
  AND2X1 U4466 ( .IN1(n4343), .IN2(g1250), .Q(n4350) );
  OR2X1 U4467 ( .IN1(n4352), .IN2(n4353), .Q(g7298) );
  AND2X1 U4468 ( .IN1(n4342), .IN2(g1240), .Q(n4353) );
  AND2X1 U4469 ( .IN1(n4343), .IN2(g1245), .Q(n4352) );
  OR2X1 U4470 ( .IN1(n4354), .IN2(n4355), .Q(g7297) );
  AND2X1 U4471 ( .IN1(n4342), .IN2(g1235), .Q(n4355) );
  AND2X1 U4472 ( .IN1(n4343), .IN2(g1240), .Q(n4354) );
  OR2X1 U4473 ( .IN1(n4356), .IN2(n4357), .Q(g7296) );
  AND2X1 U4474 ( .IN1(n4342), .IN2(g1275), .Q(n4357) );
  AND2X1 U4475 ( .IN1(n4343), .IN2(g1235), .Q(n4356) );
  OR2X1 U4476 ( .IN1(n4358), .IN2(n4359), .Q(g7295) );
  AND2X1 U4477 ( .IN1(n4342), .IN2(g1284), .Q(n4359) );
  AND2X1 U4478 ( .IN1(n4343), .IN2(g1280), .Q(n4358) );
  OR2X1 U4479 ( .IN1(n4360), .IN2(n4361), .Q(g7294) );
  AND2X1 U4480 ( .IN1(n4342), .IN2(g1292), .Q(n4361) );
  AND2X1 U4481 ( .IN1(n4343), .IN2(g1284), .Q(n4360) );
  OR2X1 U4482 ( .IN1(n4362), .IN2(n4363), .Q(g7293) );
  AND2X1 U4483 ( .IN1(n4342), .IN2(g1296), .Q(n4363) );
  AND2X1 U4484 ( .IN1(n4343), .IN2(g1292), .Q(n4362) );
  OR2X1 U4485 ( .IN1(n4364), .IN2(n4365), .Q(g7292) );
  AND2X1 U4486 ( .IN1(n4342), .IN2(g1300), .Q(n4365) );
  AND2X1 U4487 ( .IN1(n4343), .IN2(g1296), .Q(n4364) );
  OR2X1 U4488 ( .IN1(n4366), .IN2(n4367), .Q(g7291) );
  AND2X1 U4489 ( .IN1(n4342), .IN2(g1304), .Q(n4367) );
  AND2X1 U4490 ( .IN1(n4343), .IN2(g1300), .Q(n4366) );
  OR2X1 U4491 ( .IN1(n4368), .IN2(n4369), .Q(g7290) );
  AND2X1 U4492 ( .IN1(n4342), .IN2(test_so6), .Q(n4369) );
  AND2X1 U4493 ( .IN1(n4343), .IN2(g1304), .Q(n4368) );
  OR2X1 U4494 ( .IN1(n4370), .IN2(n4371), .Q(g7257) );
  AND2X1 U4495 ( .IN1(n495), .IN2(g1032), .Q(n4371) );
  AND2X1 U4496 ( .IN1(n3946), .IN2(g1077), .Q(n4370) );
  OR2X1 U4497 ( .IN1(n4372), .IN2(n4373), .Q(g7244) );
  AND2X1 U4498 ( .IN1(n495), .IN2(g1023), .Q(n4373) );
  AND2X1 U4499 ( .IN1(n3946), .IN2(g1071), .Q(n4372) );
  OR2X1 U4500 ( .IN1(n4374), .IN2(test_so10), .Q(g7219) );
  OR2X1 U4501 ( .IN1(n4374), .IN2(g8982), .Q(g7204) );
  AND2X1 U4502 ( .IN1(n4375), .IN2(n4160), .Q(g7202) );
  AND2X1 U4503 ( .IN1(n1097), .IN2(n4376), .Q(n4375) );
  OR2X1 U4504 ( .IN1(n1123), .IN2(g814), .Q(n4376) );
  OR2X1 U4505 ( .IN1(n3338), .IN2(n4377), .Q(n1097) );
  INVX0 U4506 ( .INP(n1123), .ZN(n4377) );
  AND2X1 U4507 ( .IN1(n4378), .IN2(n4166), .Q(g7191) );
  AND2X1 U4508 ( .IN1(n1099), .IN2(n4379), .Q(n4378) );
  OR2X1 U4509 ( .IN1(n1125), .IN2(g4178), .Q(n4379) );
  OR2X1 U4510 ( .IN1(n3349), .IN2(n4380), .Q(n1099) );
  OR2X1 U4511 ( .IN1(n4374), .IN2(g8980), .Q(g7189) );
  OR2X1 U4512 ( .IN1(n4374), .IN2(g8978), .Q(g7183) );
  OR2X1 U4513 ( .IN1(n4374), .IN2(g8976), .Q(g7143) );
  AND2X1 U4514 ( .IN1(n4381), .IN2(n4382), .Q(g7137) );
  OR2X1 U4515 ( .IN1(n4383), .IN2(n4304), .Q(n4382) );
  INVX0 U4516 ( .INP(n4384), .ZN(n4383) );
  OR2X1 U4517 ( .IN1(n4385), .IN2(n1709), .Q(n4384) );
  AND2X1 U4518 ( .IN1(n4381), .IN2(n4386), .Q(g7134) );
  OR2X1 U4519 ( .IN1(n4387), .IN2(n4385), .Q(n4386) );
  INVX0 U4520 ( .INP(n4388), .ZN(n4387) );
  OR2X1 U4521 ( .IN1(n4339), .IN2(n5996), .Q(n4388) );
  AND2X1 U4522 ( .IN1(n3941), .IN2(n3925), .Q(n4381) );
  INVX0 U4523 ( .INP(n3604), .ZN(n3925) );
  AND2X1 U4524 ( .IN1(n4304), .IN2(n3315), .Q(n3604) );
  AND2X1 U4525 ( .IN1(n4385), .IN2(n1709), .Q(n4304) );
  AND2X1 U4526 ( .IN1(n4339), .IN2(n5996), .Q(n4385) );
  AND2X1 U4527 ( .IN1(g627), .IN2(n1612), .Q(n4339) );
  OR2X1 U4528 ( .IN1(n4389), .IN2(g1713), .Q(g7133) );
  AND2X1 U4529 ( .IN1(n4390), .IN2(n4391), .Q(n4389) );
  OR2X1 U4530 ( .IN1(n3382), .IN2(g1766), .Q(n4390) );
  OR2X1 U4531 ( .IN1(n4392), .IN2(n233), .Q(g7032) );
  INVX0 U4532 ( .INP(n4393), .ZN(n233) );
  OR2X1 U4533 ( .IN1(n4394), .IN2(n4395), .Q(n4393) );
  OR2X1 U4534 ( .IN1(n4396), .IN2(n4397), .Q(n4395) );
  OR2X1 U4535 ( .IN1(n4398), .IN2(n4399), .Q(n4397) );
  OR2X1 U4536 ( .IN1(g143), .IN2(g148), .Q(n4399) );
  OR2X1 U4537 ( .IN1(g158), .IN2(g153), .Q(n4398) );
  OR2X1 U4538 ( .IN1(n4400), .IN2(n4401), .Q(n4396) );
  OR2X1 U4539 ( .IN1(g135), .IN2(g162), .Q(n4401) );
  OR2X1 U4540 ( .IN1(g131), .IN2(g139), .Q(n4400) );
  OR2X1 U4541 ( .IN1(n4402), .IN2(n4403), .Q(n4394) );
  OR2X1 U4542 ( .IN1(n4404), .IN2(n4405), .Q(n4403) );
  OR2X1 U4543 ( .IN1(g119), .IN2(g127), .Q(n4405) );
  INVX0 U4544 ( .INP(n4406), .ZN(n4404) );
  AND2X1 U4545 ( .IN1(g6786), .IN2(n1137), .Q(n4406) );
  OR2X1 U4546 ( .IN1(n4407), .IN2(n4408), .Q(n4402) );
  OR2X1 U4547 ( .IN1(n3267), .IN2(n3245), .Q(n4408) );
  OR2X1 U4548 ( .IN1(n3322), .IN2(n3321), .Q(n4407) );
  AND2X1 U4549 ( .IN1(g109), .IN2(g123), .Q(n4392) );
  AND2X1 U4550 ( .IN1(n1610), .IN2(n4409), .Q(g6983) );
  OR2X1 U4551 ( .IN1(n4410), .IN2(n4411), .Q(n4409) );
  AND2X1 U4552 ( .IN1(n4336), .IN2(g1791), .Q(n4411) );
  OR2X1 U4553 ( .IN1(n493), .IN2(n4191), .Q(n4336) );
  AND2X1 U4554 ( .IN1(n4412), .IN2(n238), .Q(n4410) );
  AND2X1 U4555 ( .IN1(n4191), .IN2(g1786), .Q(n4412) );
  OR2X1 U4556 ( .IN1(n4413), .IN2(n4414), .Q(n4191) );
  OR2X1 U4557 ( .IN1(n1659), .IN2(n4415), .Q(n4414) );
  OR2X1 U4558 ( .IN1(n4416), .IN2(n4417), .Q(g6934) );
  INVX0 U4559 ( .INP(n4418), .ZN(n4417) );
  OR2X1 U4560 ( .IN1(n4419), .IN2(n3322), .Q(n4418) );
  AND2X1 U4561 ( .IN1(n4419), .IN2(g284), .Q(n4416) );
  OR2X1 U4562 ( .IN1(n4420), .IN2(n4421), .Q(g6930) );
  AND2X1 U4563 ( .IN1(n495), .IN2(g1015), .Q(n4421) );
  AND2X1 U4564 ( .IN1(n3946), .IN2(g1074), .Q(n4420) );
  OR2X1 U4565 ( .IN1(n4422), .IN2(n4423), .Q(g6929) );
  AND2X1 U4566 ( .IN1(n4424), .IN2(g143), .Q(n4423) );
  AND2X1 U4567 ( .IN1(n4419), .IN2(g302), .Q(n4422) );
  OR2X1 U4568 ( .IN1(n4425), .IN2(n4426), .Q(g6928) );
  INVX0 U4569 ( .INP(n4427), .ZN(n4426) );
  OR2X1 U4570 ( .IN1(n4419), .IN2(n3321), .Q(n4427) );
  AND2X1 U4571 ( .IN1(n4419), .IN2(g281), .Q(n4425) );
  OR2X1 U4572 ( .IN1(n4428), .IN2(n4429), .Q(g6924) );
  AND2X1 U4573 ( .IN1(n495), .IN2(g1019), .Q(n4429) );
  AND2X1 U4574 ( .IN1(n3946), .IN2(g1098), .Q(n4428) );
  OR2X1 U4575 ( .IN1(n4430), .IN2(n4431), .Q(g6923) );
  AND2X1 U4576 ( .IN1(n4424), .IN2(g166), .Q(n4431) );
  AND2X1 U4577 ( .IN1(n4419), .IN2(g299), .Q(n4430) );
  OR2X1 U4578 ( .IN1(n4432), .IN2(n4433), .Q(g6922) );
  AND2X1 U4579 ( .IN1(n4424), .IN2(g162), .Q(n4433) );
  AND2X1 U4580 ( .IN1(n4419), .IN2(g278), .Q(n4432) );
  OR2X1 U4581 ( .IN1(n4434), .IN2(n4435), .Q(g6918) );
  AND2X1 U4582 ( .IN1(test_so2), .IN2(n495), .Q(n4435) );
  AND2X1 U4583 ( .IN1(n3946), .IN2(g1095), .Q(n4434) );
  OR2X1 U4584 ( .IN1(n4436), .IN2(n4437), .Q(g6916) );
  AND2X1 U4585 ( .IN1(n4424), .IN2(g139), .Q(n4437) );
  AND2X1 U4586 ( .IN1(n4419), .IN2(g296), .Q(n4436) );
  OR2X1 U4587 ( .IN1(n4438), .IN2(n4439), .Q(g6915) );
  AND2X1 U4588 ( .IN1(n4424), .IN2(g158), .Q(n4439) );
  AND2X1 U4589 ( .IN1(n4419), .IN2(g275), .Q(n4438) );
  OR2X1 U4590 ( .IN1(n4440), .IN2(n4441), .Q(g6912) );
  AND2X1 U4591 ( .IN1(n495), .IN2(g1011), .Q(n4441) );
  AND2X1 U4592 ( .IN1(n3946), .IN2(g1092), .Q(n4440) );
  OR2X1 U4593 ( .IN1(n4442), .IN2(n4443), .Q(g6911) );
  AND2X1 U4594 ( .IN1(n4424), .IN2(g135), .Q(n4443) );
  AND2X1 U4595 ( .IN1(n4419), .IN2(g293), .Q(n4442) );
  OR2X1 U4596 ( .IN1(n4444), .IN2(n4445), .Q(g6910) );
  AND2X1 U4597 ( .IN1(n4424), .IN2(g153), .Q(n4445) );
  AND2X1 U4598 ( .IN1(n4419), .IN2(g272), .Q(n4444) );
  OR2X1 U4599 ( .IN1(n4446), .IN2(n4447), .Q(g6909) );
  AND2X1 U4600 ( .IN1(n4448), .IN2(g1868), .Q(n4446) );
  OR2X1 U4601 ( .IN1(n4449), .IN2(n4450), .Q(g6908) );
  AND2X1 U4602 ( .IN1(test_so8), .IN2(n495), .Q(n4450) );
  AND2X1 U4603 ( .IN1(n3946), .IN2(g1089), .Q(n4449) );
  OR2X1 U4604 ( .IN1(n4451), .IN2(n4452), .Q(g6907) );
  AND2X1 U4605 ( .IN1(n4424), .IN2(g131), .Q(n4452) );
  AND2X1 U4606 ( .IN1(n4419), .IN2(g290), .Q(n4451) );
  OR2X1 U4607 ( .IN1(n4453), .IN2(n4454), .Q(g6906) );
  AND2X1 U4608 ( .IN1(n4424), .IN2(g148), .Q(n4454) );
  AND2X1 U4609 ( .IN1(n4419), .IN2(g269), .Q(n4453) );
  OR2X1 U4610 ( .IN1(n4455), .IN2(n4456), .Q(g6902) );
  AND2X1 U4611 ( .IN1(n495), .IN2(g1003), .Q(n4456) );
  AND2X1 U4612 ( .IN1(n3946), .IN2(g1086), .Q(n4455) );
  OR2X1 U4613 ( .IN1(n4457), .IN2(n4458), .Q(g6901) );
  AND2X1 U4614 ( .IN1(n4424), .IN2(g127), .Q(n4458) );
  AND2X1 U4615 ( .IN1(n4419), .IN2(g287), .Q(n4457) );
  OR2X1 U4616 ( .IN1(n4459), .IN2(n4460), .Q(g6900) );
  AND2X1 U4617 ( .IN1(n4424), .IN2(g178), .Q(n4460) );
  AND2X1 U4618 ( .IN1(n4419), .IN2(g266), .Q(n4459) );
  OR2X1 U4619 ( .IN1(n4461), .IN2(n4462), .Q(g6898) );
  AND2X1 U4620 ( .IN1(n495), .IN2(g991), .Q(n4462) );
  AND2X1 U4621 ( .IN1(n3946), .IN2(g1083), .Q(n4461) );
  OR2X1 U4622 ( .IN1(n4463), .IN2(n4464), .Q(g6897) );
  AND2X1 U4623 ( .IN1(n4424), .IN2(g182), .Q(n4464) );
  AND2X1 U4624 ( .IN1(n4419), .IN2(g263), .Q(n4463) );
  INVX0 U4625 ( .INP(n4424), .ZN(n4419) );
  OR2X1 U4626 ( .IN1(n650), .IN2(n4465), .Q(n4424) );
  AND2X1 U4627 ( .IN1(n1613), .IN2(n1137), .Q(n4465) );
  AND2X1 U4628 ( .IN1(n3022), .IN2(g18), .Q(n1137) );
  OR2X1 U4629 ( .IN1(n4466), .IN2(n4467), .Q(g6895) );
  AND2X1 U4630 ( .IN1(n495), .IN2(g995), .Q(n4467) );
  AND2X1 U4631 ( .IN1(n3946), .IN2(g1080), .Q(n4466) );
  OR2X1 U4632 ( .IN1(n4468), .IN2(n4469), .Q(g6894) );
  AND2X1 U4633 ( .IN1(n495), .IN2(g1027), .Q(n4469) );
  AND2X1 U4634 ( .IN1(test_so7), .IN2(n3946), .Q(n4468) );
  AND2X1 U4635 ( .IN1(n4470), .IN2(n4471), .Q(g6842) );
  AND2X1 U4636 ( .IN1(g109), .IN2(g1400), .Q(g6841) );
  AND2X1 U4637 ( .IN1(g109), .IN2(g248), .Q(g6840) );
  AND2X1 U4638 ( .IN1(g109), .IN2(g1397), .Q(g6839) );
  AND2X1 U4639 ( .IN1(g109), .IN2(n3054), .Q(g6834) );
  AND2X1 U4640 ( .IN1(g109), .IN2(n3019), .Q(g6830) );
  AND2X1 U4641 ( .IN1(g109), .IN2(n3038), .Q(g6828) );
  AND2X1 U4642 ( .IN1(g109), .IN2(n3061), .Q(g6820) );
  INVX0 U4643 ( .INP(n4472), .ZN(g6795) );
  OR2X1 U4644 ( .IN1(n4447), .IN2(n4473), .Q(n4472) );
  AND2X1 U4645 ( .IN1(n4474), .IN2(n4448), .Q(n4473) );
  INVX0 U4646 ( .INP(n102), .ZN(n4448) );
  AND2X1 U4647 ( .IN1(n4475), .IN2(n3316), .Q(n102) );
  OR2X1 U4648 ( .IN1(n4475), .IN2(n3316), .Q(n4474) );
  OR2X1 U4649 ( .IN1(n3381), .IN2(n3033), .Q(g6755) );
  AND2X1 U4650 ( .IN1(n4476), .IN2(n5997), .Q(g6747) );
  AND2X1 U4651 ( .IN1(n4477), .IN2(g109), .Q(n4476) );
  OR2X1 U4652 ( .IN1(n3041), .IN2(n3024), .Q(n4477) );
  INVX0 U4653 ( .INP(n4478), .ZN(g6733) );
  OR2X1 U4654 ( .IN1(n4479), .IN2(n4298), .Q(n4478) );
  OR2X1 U4655 ( .IN1(n1123), .IN2(n1150), .Q(n4479) );
  AND2X1 U4656 ( .IN1(n4480), .IN2(n4166), .Q(g6728) );
  AND2X1 U4657 ( .IN1(n4380), .IN2(n4481), .Q(n4480) );
  INVX0 U4658 ( .INP(n1152), .ZN(n4481) );
  INVX0 U4659 ( .INP(n1125), .ZN(n4380) );
  OR2X1 U4660 ( .IN1(n4482), .IN2(n4483), .Q(g6679) );
  AND2X1 U4661 ( .IN1(g109), .IN2(g1), .Q(n4483) );
  AND2X1 U4662 ( .IN1(n1154), .IN2(n147), .Q(n4482) );
  INVX0 U4663 ( .INP(n4484), .ZN(n147) );
  OR2X1 U4664 ( .IN1(n4485), .IN2(n4486), .Q(n4484) );
  OR2X1 U4665 ( .IN1(n4487), .IN2(n4488), .Q(n4486) );
  OR2X1 U4666 ( .IN1(g1411), .IN2(g1403), .Q(n4488) );
  OR2X1 U4667 ( .IN1(g1415), .IN2(g1407), .Q(n4487) );
  OR2X1 U4668 ( .IN1(n4489), .IN2(n4490), .Q(n4485) );
  OR2X1 U4669 ( .IN1(n3309), .IN2(n3308), .Q(n4490) );
  OR2X1 U4670 ( .IN1(n3311), .IN2(n3310), .Q(n4489) );
  AND2X1 U4671 ( .IN1(n4491), .IN2(n4492), .Q(n1154) );
  AND2X1 U4672 ( .IN1(g6234), .IN2(n4493), .Q(n4492) );
  AND2X1 U4673 ( .IN1(g1419), .IN2(n1159), .Q(n4493) );
  INVX0 U4674 ( .INP(n4494), .ZN(n4491) );
  OR2X1 U4675 ( .IN1(n4495), .IN2(n4496), .Q(n4494) );
  OR2X1 U4676 ( .IN1(n1710), .IN2(n1627), .Q(n4496) );
  OR2X1 U4677 ( .IN1(n3251), .IN2(n3250), .Q(n4495) );
  OR2X1 U4678 ( .IN1(n3379), .IN2(g627), .Q(g6672) );
  OR2X1 U4679 ( .IN1(n4497), .IN2(n4498), .Q(g6656) );
  AND2X1 U4680 ( .IN1(g109), .IN2(g4), .Q(n4498) );
  AND2X1 U4681 ( .IN1(n1161), .IN2(n145), .Q(n4497) );
  INVX0 U4682 ( .INP(n4499), .ZN(n145) );
  OR2X1 U4683 ( .IN1(n4500), .IN2(n4501), .Q(n4499) );
  OR2X1 U4684 ( .IN1(n4502), .IN2(n4503), .Q(n4501) );
  OR2X1 U4685 ( .IN1(g1482), .IN2(g1499), .Q(n4503) );
  OR2X1 U4686 ( .IN1(g1486), .IN2(g1466), .Q(n4502) );
  OR2X1 U4687 ( .IN1(n4504), .IN2(n4505), .Q(n4500) );
  OR2X1 U4688 ( .IN1(n3312), .IN2(g1458), .Q(n4505) );
  OR2X1 U4689 ( .IN1(n3314), .IN2(n3313), .Q(n4504) );
  AND2X1 U4690 ( .IN1(n4506), .IN2(n4507), .Q(n1161) );
  AND2X1 U4691 ( .IN1(n1159), .IN2(n4508), .Q(n4507) );
  AND2X1 U4692 ( .IN1(g1453), .IN2(n3378), .Q(n4508) );
  AND2X1 U4693 ( .IN1(g1504), .IN2(g109), .Q(n3378) );
  INVX0 U4694 ( .INP(n4509), .ZN(n4506) );
  OR2X1 U4695 ( .IN1(n4510), .IN2(n4511), .Q(n4509) );
  OR2X1 U4696 ( .IN1(n3280), .IN2(n1707), .Q(n4511) );
  OR2X1 U4697 ( .IN1(n3282), .IN2(n3281), .Q(n4510) );
  AND2X1 U4698 ( .IN1(n3585), .IN2(g8983), .Q(g6653) );
  AND2X1 U4699 ( .IN1(n3585), .IN2(g8981), .Q(g6638) );
  AND2X1 U4700 ( .IN1(n3585), .IN2(g8979), .Q(g6627) );
  AND2X1 U4701 ( .IN1(n3585), .IN2(g8977), .Q(g6621) );
  OR2X1 U4702 ( .IN1(n4512), .IN2(n4513), .Q(g6551) );
  INVX0 U4703 ( .INP(n4514), .ZN(n4513) );
  OR2X1 U4704 ( .IN1(n4515), .IN2(n3314), .Q(n4514) );
  AND2X1 U4705 ( .IN1(n4515), .IN2(g1546), .Q(n4512) );
  OR2X1 U4706 ( .IN1(n4516), .IN2(n4517), .Q(g6546) );
  AND2X1 U4707 ( .IN1(n4518), .IN2(g1453), .Q(n4517) );
  AND2X1 U4708 ( .IN1(n4515), .IN2(g1564), .Q(n4516) );
  OR2X1 U4709 ( .IN1(n4519), .IN2(n4520), .Q(g6545) );
  AND2X1 U4710 ( .IN1(n4518), .IN2(g1482), .Q(n4520) );
  AND2X1 U4711 ( .IN1(n4515), .IN2(g1543), .Q(n4519) );
  OR2X1 U4712 ( .IN1(n4521), .IN2(n4522), .Q(g6542) );
  AND2X1 U4713 ( .IN1(n4518), .IN2(g1458), .Q(n4522) );
  AND2X1 U4714 ( .IN1(n4515), .IN2(g1561), .Q(n4521) );
  OR2X1 U4715 ( .IN1(n4523), .IN2(n4524), .Q(g6541) );
  AND2X1 U4716 ( .IN1(n4518), .IN2(g1486), .Q(n4524) );
  AND2X1 U4717 ( .IN1(n4515), .IN2(g1540), .Q(n4523) );
  OR2X1 U4718 ( .IN1(n4525), .IN2(n4526), .Q(g6538) );
  AND2X1 U4719 ( .IN1(n4518), .IN2(g1462), .Q(n4526) );
  AND2X1 U4720 ( .IN1(n4515), .IN2(g1558), .Q(n4525) );
  OR2X1 U4721 ( .IN1(n4527), .IN2(n4528), .Q(g6537) );
  AND2X1 U4722 ( .IN1(n4518), .IN2(g1490), .Q(n4528) );
  AND2X1 U4723 ( .IN1(n4515), .IN2(g1537), .Q(n4527) );
  OR2X1 U4724 ( .IN1(n4529), .IN2(n4530), .Q(g6534) );
  AND2X1 U4725 ( .IN1(n4518), .IN2(g1466), .Q(n4530) );
  AND2X1 U4726 ( .IN1(n4515), .IN2(g1555), .Q(n4529) );
  OR2X1 U4727 ( .IN1(n4531), .IN2(n4532), .Q(g6533) );
  AND2X1 U4728 ( .IN1(n4518), .IN2(g1494), .Q(n4532) );
  AND2X1 U4729 ( .IN1(n4515), .IN2(g1534), .Q(n4531) );
  AND2X1 U4730 ( .IN1(n3585), .IN2(g8986), .Q(g6531) );
  OR2X1 U4731 ( .IN1(n4533), .IN2(n4534), .Q(g6529) );
  INVX0 U4732 ( .INP(n4535), .ZN(n4534) );
  OR2X1 U4733 ( .IN1(n4515), .IN2(n3282), .Q(n4535) );
  AND2X1 U4734 ( .IN1(n4515), .IN2(g1552), .Q(n4533) );
  OR2X1 U4735 ( .IN1(n4536), .IN2(n4537), .Q(g6528) );
  AND2X1 U4736 ( .IN1(n4518), .IN2(g1499), .Q(n4537) );
  AND2X1 U4737 ( .IN1(n4515), .IN2(g1531), .Q(n4536) );
  AND2X1 U4738 ( .IN1(n3585), .IN2(g8985), .Q(g6526) );
  AND2X1 U4739 ( .IN1(n4538), .IN2(n1610), .Q(g6525) );
  AND2X1 U4740 ( .IN1(n4539), .IN2(n4540), .Q(n4538) );
  OR2X1 U4741 ( .IN1(n238), .IN2(g1786), .Q(n4540) );
  INVX0 U4742 ( .INP(n4541), .ZN(n238) );
  OR2X1 U4743 ( .IN1(n3332), .IN2(n4541), .Q(n4539) );
  OR2X1 U4744 ( .IN1(n4542), .IN2(n4543), .Q(g6524) );
  INVX0 U4745 ( .INP(n4544), .ZN(n4543) );
  OR2X1 U4746 ( .IN1(n4515), .IN2(n3310), .Q(n4544) );
  AND2X1 U4747 ( .IN1(n4515), .IN2(g1589), .Q(n4542) );
  OR2X1 U4748 ( .IN1(n4545), .IN2(n4546), .Q(g6523) );
  AND2X1 U4749 ( .IN1(n4518), .IN2(g1474), .Q(n4546) );
  AND2X1 U4750 ( .IN1(n4515), .IN2(g1549), .Q(n4545) );
  OR2X1 U4751 ( .IN1(n4547), .IN2(n4548), .Q(g6522) );
  AND2X1 U4752 ( .IN1(n4518), .IN2(g1504), .Q(n4548) );
  AND2X1 U4753 ( .IN1(n4515), .IN2(g1528), .Q(n4547) );
  AND2X1 U4754 ( .IN1(n4549), .IN2(n1610), .Q(g6516) );
  AND2X1 U4755 ( .IN1(n4550), .IN2(n4541), .Q(n4549) );
  OR2X1 U4756 ( .IN1(n1659), .IN2(n4551), .Q(n4541) );
  INVX0 U4757 ( .INP(n4552), .ZN(n4550) );
  AND2X1 U4758 ( .IN1(n4551), .IN2(n1659), .Q(n4552) );
  OR2X1 U4759 ( .IN1(n4553), .IN2(n4554), .Q(g6515) );
  AND2X1 U4760 ( .IN1(n4518), .IN2(g1448), .Q(n4554) );
  AND2X1 U4761 ( .IN1(n4515), .IN2(g1607), .Q(n4553) );
  OR2X1 U4762 ( .IN1(n4555), .IN2(n4556), .Q(g6514) );
  AND2X1 U4763 ( .IN1(n4518), .IN2(g1407), .Q(n4556) );
  AND2X1 U4764 ( .IN1(n4515), .IN2(g1586), .Q(n4555) );
  OR2X1 U4765 ( .IN1(n4557), .IN2(n4558), .Q(g6513) );
  AND2X1 U4766 ( .IN1(n4518), .IN2(g1508), .Q(n4558) );
  AND2X1 U4767 ( .IN1(n4515), .IN2(g1524), .Q(n4557) );
  AND2X1 U4768 ( .IN1(n1610), .IN2(n4559), .Q(g6508) );
  OR2X1 U4769 ( .IN1(n4560), .IN2(n4561), .Q(n4559) );
  AND2X1 U4770 ( .IN1(n4551), .IN2(g1776), .Q(n4561) );
  OR2X1 U4771 ( .IN1(n493), .IN2(n4415), .Q(n4551) );
  AND2X1 U4772 ( .IN1(n4562), .IN2(n4563), .Q(n4560) );
  AND2X1 U4773 ( .IN1(test_so5), .IN2(n4415), .Q(n4562) );
  OR2X1 U4774 ( .IN1(n4564), .IN2(n4565), .Q(g6507) );
  INVX0 U4775 ( .INP(n4566), .ZN(n4565) );
  OR2X1 U4776 ( .IN1(n4515), .IN2(n3311), .Q(n4566) );
  AND2X1 U4777 ( .IN1(n4515), .IN2(g1604), .Q(n4564) );
  OR2X1 U4778 ( .IN1(n4567), .IN2(n4568), .Q(g6506) );
  AND2X1 U4779 ( .IN1(n4518), .IN2(g1424), .Q(n4568) );
  AND2X1 U4780 ( .IN1(n4515), .IN2(g1583), .Q(n4567) );
  AND2X1 U4781 ( .IN1(n1610), .IN2(n4569), .Q(g6502) );
  OR2X1 U4782 ( .IN1(n4570), .IN2(n4571), .Q(n4569) );
  AND2X1 U4783 ( .IN1(n4563), .IN2(n3383), .Q(n4571) );
  INVX0 U4784 ( .INP(n4391), .ZN(n4563) );
  AND2X1 U4785 ( .IN1(test_so5), .IN2(n4391), .Q(n4570) );
  OR2X1 U4786 ( .IN1(n3340), .IN2(n493), .Q(n4391) );
  OR2X1 U4787 ( .IN1(n4572), .IN2(n4573), .Q(g6501) );
  INVX0 U4788 ( .INP(n4574), .ZN(n4573) );
  OR2X1 U4789 ( .IN1(n4515), .IN2(n3309), .Q(n4574) );
  AND2X1 U4790 ( .IN1(n4515), .IN2(g1601), .Q(n4572) );
  OR2X1 U4791 ( .IN1(n4575), .IN2(n4576), .Q(g6500) );
  AND2X1 U4792 ( .IN1(n4518), .IN2(g1411), .Q(n4576) );
  AND2X1 U4793 ( .IN1(n4515), .IN2(g1580), .Q(n4575) );
  OR2X1 U4794 ( .IN1(n4577), .IN2(n4578), .Q(g6481) );
  INVX0 U4795 ( .INP(n4579), .ZN(n4578) );
  OR2X1 U4796 ( .IN1(n4515), .IN2(n3308), .Q(n4579) );
  AND2X1 U4797 ( .IN1(n4515), .IN2(g1598), .Q(n4577) );
  OR2X1 U4798 ( .IN1(n4580), .IN2(n4581), .Q(g6480) );
  AND2X1 U4799 ( .IN1(n4518), .IN2(g1419), .Q(n4581) );
  AND2X1 U4800 ( .IN1(n4515), .IN2(g1577), .Q(n4580) );
  OR2X1 U4801 ( .IN1(n4582), .IN2(n4583), .Q(g6479) );
  INVX0 U4802 ( .INP(n4584), .ZN(n4583) );
  OR2X1 U4803 ( .IN1(n4515), .IN2(n3251), .Q(n4584) );
  AND2X1 U4804 ( .IN1(n4515), .IN2(g1595), .Q(n4582) );
  OR2X1 U4805 ( .IN1(n4585), .IN2(n4586), .Q(g6478) );
  AND2X1 U4806 ( .IN1(n4518), .IN2(g1515), .Q(n4586) );
  AND2X1 U4807 ( .IN1(n4515), .IN2(g1574), .Q(n4585) );
  AND2X1 U4808 ( .IN1(n4587), .IN2(n4588), .Q(g6471) );
  OR2X1 U4809 ( .IN1(n4589), .IN2(n4475), .Q(n4588) );
  AND2X1 U4810 ( .IN1(n3033), .IN2(n3318), .Q(n4475) );
  AND2X1 U4811 ( .IN1(n5998), .IN2(g1861), .Q(n4589) );
  OR2X1 U4812 ( .IN1(n4590), .IN2(n4591), .Q(g6470) );
  AND2X1 U4813 ( .IN1(n4518), .IN2(g1403), .Q(n4591) );
  AND2X1 U4814 ( .IN1(n4515), .IN2(g1592), .Q(n4590) );
  OR2X1 U4815 ( .IN1(n4592), .IN2(n4593), .Q(g6469) );
  AND2X1 U4816 ( .IN1(n4518), .IN2(g1520), .Q(n4593) );
  AND2X1 U4817 ( .IN1(n4515), .IN2(g1571), .Q(n4592) );
  OR2X1 U4818 ( .IN1(n4594), .IN2(n4595), .Q(g6468) );
  AND2X1 U4819 ( .IN1(n4518), .IN2(g1415), .Q(n4595) );
  AND2X1 U4820 ( .IN1(n4515), .IN2(g1567), .Q(n4594) );
  INVX0 U4821 ( .INP(n4518), .ZN(n4515) );
  OR2X1 U4822 ( .IN1(n1159), .IN2(n650), .Q(n4518) );
  AND2X1 U4823 ( .IN1(n4596), .IN2(g109), .Q(g6439) );
  OR2X1 U4824 ( .IN1(n4597), .IN2(n4598), .Q(n4596) );
  AND2X1 U4825 ( .IN1(n4599), .IN2(n4600), .Q(n4598) );
  INVX0 U4826 ( .INP(n4601), .ZN(n4597) );
  OR2X1 U4827 ( .IN1(n4600), .IN2(n4599), .Q(n4601) );
  OR2X1 U4828 ( .IN1(n4602), .IN2(n4603), .Q(n4599) );
  AND2X1 U4829 ( .IN1(n3267), .IN2(g153), .Q(n4603) );
  AND2X1 U4830 ( .IN1(n3268), .IN2(g182), .Q(n4602) );
  INVX0 U4831 ( .INP(n4604), .ZN(n4600) );
  OR2X1 U4832 ( .IN1(n4605), .IN2(n4606), .Q(n4604) );
  AND2X1 U4833 ( .IN1(n3269), .IN2(g148), .Q(n4606) );
  AND2X1 U4834 ( .IN1(n3270), .IN2(g143), .Q(n4605) );
  AND2X1 U4835 ( .IN1(n4607), .IN2(n4608), .Q(g6392) );
  INVX0 U4836 ( .INP(n4609), .ZN(n4607) );
  AND2X1 U4837 ( .IN1(g109), .IN2(g881), .Q(n4609) );
  AND2X1 U4838 ( .IN1(g109), .IN2(g1389), .Q(g6334) );
  AND2X1 U4839 ( .IN1(g109), .IN2(n3020), .Q(g6332) );
  OR2X1 U4840 ( .IN1(n4298), .IN2(n4610), .Q(g6243) );
  OR2X1 U4841 ( .IN1(n4611), .IN2(n4612), .Q(n4610) );
  INVX0 U4842 ( .INP(n4613), .ZN(n4612) );
  OR2X1 U4843 ( .IN1(g798), .IN2(n3346), .Q(n4613) );
  AND2X1 U4844 ( .IN1(n3346), .IN2(g798), .Q(n4611) );
  AND2X1 U4845 ( .IN1(g109), .IN2(g1520), .Q(g6224) );
  AND2X1 U4846 ( .IN1(g109), .IN2(g1515), .Q(g6205) );
  AND2X1 U4847 ( .IN1(g109), .IN2(g1453), .Q(g6180) );
  AND2X1 U4848 ( .IN1(n60), .IN2(n3041), .Q(g6179) );
  AND2X1 U4849 ( .IN1(n4614), .IN2(g6331), .Q(n60) );
  OR2X1 U4850 ( .IN1(n4615), .IN2(n4616), .Q(g6155) );
  AND2X1 U4851 ( .IN1(n4617), .IN2(n1653), .Q(n4616) );
  AND2X1 U4852 ( .IN1(g1700), .IN2(g1707), .Q(n4617) );
  AND2X1 U4853 ( .IN1(g4076), .IN2(g1690), .Q(n4615) );
  AND2X1 U4854 ( .IN1(n4618), .IN2(n4160), .Q(g6126) );
  INVX0 U4855 ( .INP(n4298), .ZN(n4160) );
  AND2X1 U4856 ( .IN1(n1151), .IN2(n4619), .Q(n4618) );
  INVX0 U4857 ( .INP(n4620), .ZN(n4619) );
  AND2X1 U4858 ( .IN1(n4621), .IN2(n3339), .Q(n4620) );
  OR2X1 U4859 ( .IN1(n3339), .IN2(n4621), .Q(n1151) );
  AND2X1 U4860 ( .IN1(n4622), .IN2(n4166), .Q(g6123) );
  AND2X1 U4861 ( .IN1(n1153), .IN2(n4623), .Q(n4622) );
  OR2X1 U4862 ( .IN1(n1193), .IN2(g4176), .Q(n4623) );
  OR2X1 U4863 ( .IN1(n3350), .IN2(n4624), .Q(n1153) );
  OR2X1 U4864 ( .IN1(n4625), .IN2(n4626), .Q(g6099) );
  AND2X1 U4865 ( .IN1(n4627), .IN2(g1074), .Q(n4626) );
  AND2X1 U4866 ( .IN1(n4628), .IN2(g342), .Q(n4625) );
  OR2X1 U4867 ( .IN1(n4629), .IN2(n4630), .Q(g6096) );
  AND2X1 U4868 ( .IN1(n4627), .IN2(g1098), .Q(n4630) );
  AND2X1 U4869 ( .IN1(n4628), .IN2(g366), .Q(n4629) );
  OR2X1 U4870 ( .IN1(n4631), .IN2(n4632), .Q(g6093) );
  AND2X1 U4871 ( .IN1(n4627), .IN2(g1095), .Q(n4632) );
  AND2X1 U4872 ( .IN1(n4628), .IN2(g363), .Q(n4631) );
  OR2X1 U4873 ( .IN1(n4633), .IN2(n4634), .Q(g6088) );
  AND2X1 U4874 ( .IN1(n4627), .IN2(g1092), .Q(n4634) );
  AND2X1 U4875 ( .IN1(n4628), .IN2(g360), .Q(n4633) );
  OR2X1 U4876 ( .IN1(n4635), .IN2(n4636), .Q(g6080) );
  AND2X1 U4877 ( .IN1(n4627), .IN2(g1089), .Q(n4636) );
  AND2X1 U4878 ( .IN1(n4628), .IN2(g357), .Q(n4635) );
  OR2X1 U4879 ( .IN1(n4637), .IN2(n4638), .Q(g6071) );
  AND2X1 U4880 ( .IN1(n4627), .IN2(g1086), .Q(n4638) );
  AND2X1 U4881 ( .IN1(n4628), .IN2(g354), .Q(n4637) );
  OR2X1 U4882 ( .IN1(n4639), .IN2(n4640), .Q(g6068) );
  AND2X1 U4883 ( .IN1(n4627), .IN2(g1083), .Q(n4640) );
  AND2X1 U4884 ( .IN1(n4628), .IN2(g351), .Q(n4639) );
  OR2X1 U4885 ( .IN1(n4641), .IN2(n4642), .Q(g6059) );
  AND2X1 U4886 ( .IN1(n4627), .IN2(g1080), .Q(n4642) );
  AND2X1 U4887 ( .IN1(n4628), .IN2(g348), .Q(n4641) );
  OR2X1 U4888 ( .IN1(n4643), .IN2(n4644), .Q(g6054) );
  AND2X1 U4889 ( .IN1(test_so7), .IN2(n4627), .Q(n4644) );
  AND2X1 U4890 ( .IN1(n4628), .IN2(g336), .Q(n4643) );
  OR2X1 U4891 ( .IN1(n4645), .IN2(n4646), .Q(g6049) );
  AND2X1 U4892 ( .IN1(n3963), .IN2(g549), .Q(n4646) );
  OR2X1 U4893 ( .IN1(n4647), .IN2(n4648), .Q(g6045) );
  AND2X1 U4894 ( .IN1(n3963), .IN2(g575), .Q(n4648) );
  OR2X1 U4895 ( .IN1(n4649), .IN2(n4650), .Q(g6042) );
  AND2X1 U4896 ( .IN1(n3963), .IN2(g572), .Q(n4650) );
  OR2X1 U4897 ( .IN1(n4651), .IN2(n4033), .Q(g6038) );
  AND2X1 U4898 ( .IN1(n3963), .IN2(g569), .Q(n4651) );
  OR2X1 U4899 ( .IN1(n4652), .IN2(n4008), .Q(g6035) );
  AND2X1 U4900 ( .IN1(n3963), .IN2(g566), .Q(n4652) );
  OR2X1 U4901 ( .IN1(n4653), .IN2(n3978), .Q(g6026) );
  AND2X1 U4902 ( .IN1(n3963), .IN2(g563), .Q(n4653) );
  OR2X1 U4903 ( .IN1(n4654), .IN2(n3961), .Q(g6015) );
  AND2X1 U4904 ( .IN1(n3963), .IN2(g560), .Q(n4654) );
  OR2X1 U4905 ( .IN1(n4655), .IN2(n4045), .Q(g6002) );
  AND2X1 U4906 ( .IN1(n3963), .IN2(g557), .Q(n4655) );
  OR2X1 U4907 ( .IN1(n4656), .IN2(n4021), .Q(g6000) );
  AND2X1 U4908 ( .IN1(n3963), .IN2(g554), .Q(n4656) );
  OR2X1 U4909 ( .IN1(n4657), .IN2(n3996), .Q(g5996) );
  AND2X1 U4910 ( .IN1(n3963), .IN2(g546), .Q(n4657) );
  OR2X1 U4911 ( .IN1(n4658), .IN2(n1195), .Q(g5918) );
  AND2X1 U4912 ( .IN1(g109), .IN2(g119), .Q(n4658) );
  OR2X1 U4913 ( .IN1(n4659), .IN2(n4660), .Q(g5914) );
  AND2X1 U4914 ( .IN1(n4627), .IN2(g1077), .Q(n4660) );
  AND2X1 U4915 ( .IN1(n4628), .IN2(g345), .Q(n4659) );
  OR2X1 U4916 ( .IN1(n4661), .IN2(n4662), .Q(g5910) );
  AND2X1 U4917 ( .IN1(n4627), .IN2(g1071), .Q(n4662) );
  AND2X1 U4918 ( .IN1(n4628), .IN2(g339), .Q(n4661) );
  AND2X1 U4919 ( .IN1(n4663), .IN2(g109), .Q(g5770) );
  OR2X1 U4920 ( .IN1(n4664), .IN2(n4665), .Q(n4663) );
  AND2X1 U4921 ( .IN1(n4666), .IN2(n4667), .Q(n4665) );
  INVX0 U4922 ( .INP(n4668), .ZN(n4664) );
  OR2X1 U4923 ( .IN1(n4667), .IN2(n4666), .Q(n4668) );
  OR2X1 U4924 ( .IN1(n4669), .IN2(n4670), .Q(n4666) );
  AND2X1 U4925 ( .IN1(n1628), .IN2(g1508), .Q(n4670) );
  AND2X1 U4926 ( .IN1(n1707), .IN2(g1453), .Q(n4669) );
  INVX0 U4927 ( .INP(n4671), .ZN(n4667) );
  OR2X1 U4928 ( .IN1(n4672), .IN2(n4673), .Q(n4671) );
  AND2X1 U4929 ( .IN1(n3271), .IN2(g1494), .Q(n4673) );
  AND2X1 U4930 ( .IN1(n3280), .IN2(g1499), .Q(n4672) );
  AND2X1 U4931 ( .IN1(n4674), .IN2(n4675), .Q(g5763) );
  OR2X1 U4932 ( .IN1(n6003), .IN2(n650), .Q(n4674) );
  OR2X1 U4933 ( .IN1(n4676), .IN2(n4677), .Q(g5755) );
  AND2X1 U4934 ( .IN1(n4678), .IN2(n1678), .Q(n4677) );
  AND2X1 U4935 ( .IN1(n4679), .IN2(n4680), .Q(n4678) );
  OR2X1 U4936 ( .IN1(n4681), .IN2(n4682), .Q(n4680) );
  AND2X1 U4937 ( .IN1(n1619), .IN2(g109), .Q(n4681) );
  OR2X1 U4938 ( .IN1(g6331), .IN2(n4683), .Q(n4679) );
  AND2X1 U4939 ( .IN1(g201), .IN2(g109), .Q(g6331) );
  AND2X1 U4940 ( .IN1(g6333), .IN2(n4684), .Q(n4676) );
  OR2X1 U4941 ( .IN1(n4685), .IN2(n4686), .Q(n4684) );
  AND2X1 U4942 ( .IN1(n4683), .IN2(g201), .Q(n4686) );
  AND2X1 U4943 ( .IN1(n4682), .IN2(n1619), .Q(n4685) );
  INVX0 U4944 ( .INP(n4683), .ZN(n4682) );
  OR2X1 U4945 ( .IN1(n4687), .IN2(n4688), .Q(n4683) );
  AND2X1 U4946 ( .IN1(n3333), .IN2(g1389), .Q(n4688) );
  AND2X1 U4947 ( .IN1(n1603), .IN2(n4689), .Q(n4687) );
  OR2X1 U4948 ( .IN1(n59), .IN2(g1386), .Q(n4689) );
  AND2X1 U4949 ( .IN1(n4614), .IN2(n1619), .Q(n59) );
  INVX0 U4950 ( .INP(n4690), .ZN(n4614) );
  OR2X1 U4951 ( .IN1(n4691), .IN2(n4692), .Q(n4690) );
  OR2X1 U4952 ( .IN1(n4693), .IN2(n4694), .Q(n4692) );
  OR2X1 U4953 ( .IN1(n4695), .IN2(n4696), .Q(n4694) );
  OR2X1 U4954 ( .IN1(g1383), .IN2(n3020), .Q(n4696) );
  OR2X1 U4955 ( .IN1(n3019), .IN2(n4697), .Q(n4695) );
  OR2X1 U4956 ( .IN1(g1371), .IN2(n3038), .Q(n4697) );
  INVX0 U4957 ( .INP(n4698), .ZN(n4693) );
  AND2X1 U4958 ( .IN1(n4699), .IN2(n4700), .Q(n4698) );
  AND2X1 U4959 ( .IN1(n5999), .IN2(n4701), .Q(n4700) );
  AND2X1 U4960 ( .IN1(n3360), .IN2(n6000), .Q(n4701) );
  AND2X1 U4961 ( .IN1(n3359), .IN2(n4702), .Q(n4699) );
  AND2X1 U4962 ( .IN1(n3357), .IN2(n3358), .Q(n4702) );
  OR2X1 U4963 ( .IN1(n4703), .IN2(n4704), .Q(n4691) );
  OR2X1 U4964 ( .IN1(n4705), .IN2(n4706), .Q(n4704) );
  OR2X1 U4965 ( .IN1(g186), .IN2(n4707), .Q(n4706) );
  OR2X1 U4966 ( .IN1(g213), .IN2(g237), .Q(n4707) );
  OR2X1 U4967 ( .IN1(g1386), .IN2(n4708), .Q(n4705) );
  OR2X1 U4968 ( .IN1(g192), .IN2(g243), .Q(n4708) );
  OR2X1 U4969 ( .IN1(n4709), .IN2(n4710), .Q(n4703) );
  OR2X1 U4970 ( .IN1(g1397), .IN2(n4711), .Q(n4710) );
  OR2X1 U4971 ( .IN1(g1400), .IN2(g197), .Q(n4711) );
  OR2X1 U4972 ( .IN1(g1389), .IN2(n4712), .Q(n4709) );
  OR2X1 U4973 ( .IN1(test_so3), .IN2(g248), .Q(n4712) );
  AND2X1 U4974 ( .IN1(g197), .IN2(g109), .Q(g6333) );
  AND2X1 U4975 ( .IN1(n4713), .IN2(g744), .Q(g5659) );
  AND2X1 U4976 ( .IN1(g743), .IN2(g109), .Q(n4713) );
  AND2X1 U4977 ( .IN1(n4714), .IN2(g742), .Q(g5658) );
  AND2X1 U4978 ( .IN1(g741), .IN2(g109), .Q(n4714) );
  AND2X1 U4979 ( .IN1(n4715), .IN2(n4716), .Q(g5556) );
  AND2X1 U4980 ( .IN1(n4717), .IN2(n4718), .Q(n4716) );
  AND2X1 U4981 ( .IN1(g1806), .IN2(g1707), .Q(n4718) );
  AND2X1 U4982 ( .IN1(g1690), .IN2(g1801), .Q(n4717) );
  INVX0 U4983 ( .INP(n4719), .ZN(n4715) );
  OR2X1 U4984 ( .IN1(n4720), .IN2(n4721), .Q(n4719) );
  OR2X1 U4985 ( .IN1(n4415), .IN2(n1626), .Q(n4721) );
  OR2X1 U4986 ( .IN1(n1715), .IN2(n4722), .Q(n4415) );
  OR2X1 U4987 ( .IN1(g1781), .IN2(n4413), .Q(n4720) );
  AND2X1 U4988 ( .IN1(n4723), .IN2(n4621), .Q(g5543) );
  OR2X1 U4989 ( .IN1(n1622), .IN2(n4087), .Q(n4621) );
  OR2X1 U4990 ( .IN1(n1717), .IN2(n3346), .Q(n4087) );
  INVX0 U4991 ( .INP(n4724), .ZN(n4723) );
  AND2X1 U4992 ( .IN1(n4725), .IN2(n4726), .Q(n4724) );
  OR2X1 U4993 ( .IN1(g5849), .IN2(n1717), .Q(n4726) );
  OR2X1 U4994 ( .IN1(n3346), .IN2(n4298), .Q(g5849) );
  OR2X1 U4995 ( .IN1(n4298), .IN2(n1622), .Q(n4725) );
  OR2X1 U4996 ( .IN1(n650), .IN2(n4727), .Q(n4298) );
  OR2X1 U4997 ( .IN1(n3317), .IN2(n3128), .Q(n4727) );
  AND2X1 U4998 ( .IN1(n4728), .IN2(n4166), .Q(g5536) );
  AND2X1 U4999 ( .IN1(n4624), .IN2(n4729), .Q(n4728) );
  INVX0 U5000 ( .INP(n1213), .ZN(n4729) );
  INVX0 U5001 ( .INP(n1193), .ZN(n4624) );
  OR2X1 U5002 ( .IN1(n4730), .IN2(n4731), .Q(g5529) );
  AND2X1 U5003 ( .IN1(n4732), .IN2(n3352), .Q(n4731) );
  AND2X1 U5004 ( .IN1(n4166), .IN2(g4173), .Q(n4732) );
  AND2X1 U5005 ( .IN1(g4940), .IN2(g4174), .Q(n4730) );
  OR2X1 U5006 ( .IN1(n4733), .IN2(n1195), .Q(g5445) );
  AND2X1 U5007 ( .IN1(g109), .IN2(g12), .Q(n4733) );
  OR2X1 U5008 ( .IN1(n4734), .IN2(n1195), .Q(g5421) );
  AND2X1 U5009 ( .IN1(g109), .IN2(g9), .Q(n4734) );
  OR2X1 U5010 ( .IN1(n4735), .IN2(n4736), .Q(g5404) );
  AND2X1 U5011 ( .IN1(n495), .IN2(g1718), .Q(n4736) );
  AND2X1 U5012 ( .IN1(n3946), .IN2(g1713), .Q(n4735) );
  OR2X1 U5013 ( .IN1(n4737), .IN2(n4738), .Q(g5396) );
  AND2X1 U5014 ( .IN1(n495), .IN2(g1713), .Q(n4738) );
  AND2X1 U5015 ( .IN1(n3946), .IN2(g1710), .Q(n4737) );
  AND2X1 U5016 ( .IN1(n4739), .IN2(g1101), .Q(g5390) );
  AND2X1 U5017 ( .IN1(n4739), .IN2(g1110), .Q(g5173) );
  AND2X1 U5018 ( .IN1(n4739), .IN2(g1107), .Q(g5148) );
  AND2X1 U5019 ( .IN1(n4739), .IN2(g1104), .Q(g5126) );
  INVX0 U5020 ( .INP(n4740), .ZN(n4739) );
  OR2X1 U5021 ( .IN1(n650), .IN2(n3056), .Q(n4740) );
  AND2X1 U5022 ( .IN1(n4741), .IN2(n4742), .Q(g5083) );
  AND2X1 U5023 ( .IN1(n495), .IN2(n4470), .Q(n4741) );
  INVX0 U5024 ( .INP(g4089), .ZN(n4470) );
  AND2X1 U5025 ( .IN1(n4166), .IN2(n3351), .Q(g4940) );
  AND2X1 U5026 ( .IN1(n3388), .IN2(g109), .Q(n4166) );
  AND2X1 U5027 ( .IN1(n4743), .IN2(n3018), .Q(g4905) );
  AND2X1 U5028 ( .IN1(n4743), .IN2(n3037), .Q(g4903) );
  AND2X1 U5029 ( .IN1(n4743), .IN2(n3030), .Q(g4902) );
  INVX0 U5030 ( .INP(n3381), .ZN(n4743) );
  AND2X1 U5031 ( .IN1(n4744), .IN2(n3053), .Q(g4893) );
  AND2X1 U5032 ( .IN1(n4744), .IN2(n3055), .Q(g4891) );
  AND2X1 U5033 ( .IN1(n4744), .IN2(n3035), .Q(g4890) );
  INVX0 U5034 ( .INP(n3379), .ZN(n4744) );
  OR2X1 U5035 ( .IN1(n4745), .IN2(n3651), .Q(n3379) );
  INVX0 U5036 ( .INP(n3941), .ZN(n3651) );
  OR2X1 U5037 ( .IN1(n3933), .IN2(n4746), .Q(n3941) );
  OR2X1 U5038 ( .IN1(g599), .IN2(g611), .Q(n4746) );
  OR2X1 U5039 ( .IN1(g605), .IN2(g591), .Q(n3933) );
  AND2X1 U5040 ( .IN1(n1607), .IN2(g611), .Q(n4745) );
  INVX0 U5041 ( .INP(n4747), .ZN(g4506) );
  OR2X1 U5042 ( .IN1(n650), .IN2(n6001), .Q(n4747) );
  INVX0 U5043 ( .INP(n4748), .ZN(g4500) );
  OR2X1 U5044 ( .IN1(n3946), .IN2(n6004), .Q(n4748) );
  INVX0 U5045 ( .INP(n4749), .ZN(g4498) );
  OR2X1 U5046 ( .IN1(n650), .IN2(n1617), .Q(n4749) );
  INVX0 U5047 ( .INP(n4750), .ZN(g4490) );
  OR2X1 U5048 ( .IN1(n650), .IN2(n1660), .Q(n4750) );
  AND2X1 U5049 ( .IN1(g109), .IN2(g1137), .Q(g4484) );
  INVX0 U5050 ( .INP(n4751), .ZN(g4480) );
  OR2X1 U5051 ( .IN1(n650), .IN2(n1706), .Q(n4751) );
  INVX0 U5052 ( .INP(n4752), .ZN(g4477) );
  OR2X1 U5053 ( .IN1(n650), .IN2(n1705), .Q(n4752) );
  INVX0 U5054 ( .INP(n4753), .ZN(g4473) );
  OR2X1 U5055 ( .IN1(n650), .IN2(n1708), .Q(n4753) );
  INVX0 U5056 ( .INP(n4754), .ZN(g4471) );
  OR2X1 U5057 ( .IN1(n650), .IN2(n1618), .Q(n4754) );
  AND2X1 U5058 ( .IN1(test_so4), .IN2(g109), .Q(g4465) );
  AND2X1 U5059 ( .IN1(g109), .IN2(g1149), .Q(g4342) );
  AND2X1 U5060 ( .IN1(g109), .IN2(g1153), .Q(g4340) );
  OR2X1 U5061 ( .IN1(n4755), .IN2(n4756), .Q(g4309) );
  AND2X1 U5062 ( .IN1(n4757), .IN2(g1762), .Q(n4756) );
  AND2X1 U5063 ( .IN1(n4758), .IN2(g1806), .Q(n4755) );
  OR2X1 U5064 ( .IN1(n4759), .IN2(n4760), .Q(g4293) );
  AND2X1 U5065 ( .IN1(n4757), .IN2(g1759), .Q(n4760) );
  AND2X1 U5066 ( .IN1(n4758), .IN2(g1801), .Q(n4759) );
  OR2X1 U5067 ( .IN1(n4761), .IN2(n4762), .Q(g4283) );
  AND2X1 U5068 ( .IN1(n4757), .IN2(g1756), .Q(n4762) );
  AND2X1 U5069 ( .IN1(n4758), .IN2(g1796), .Q(n4761) );
  OR2X1 U5070 ( .IN1(n4763), .IN2(n4764), .Q(g4274) );
  AND2X1 U5071 ( .IN1(n4757), .IN2(g1753), .Q(n4764) );
  AND2X1 U5072 ( .IN1(n4758), .IN2(g1791), .Q(n4763) );
  OR2X1 U5073 ( .IN1(n4765), .IN2(n4766), .Q(g4264) );
  AND2X1 U5074 ( .IN1(n4757), .IN2(g1750), .Q(n4766) );
  AND2X1 U5075 ( .IN1(n4758), .IN2(g1786), .Q(n4765) );
  OR2X1 U5076 ( .IN1(n4767), .IN2(n4768), .Q(g4255) );
  AND2X1 U5077 ( .IN1(n4757), .IN2(g1747), .Q(n4768) );
  AND2X1 U5078 ( .IN1(n4758), .IN2(g1781), .Q(n4767) );
  OR2X1 U5079 ( .IN1(n4769), .IN2(n4770), .Q(g4239) );
  AND2X1 U5080 ( .IN1(n4757), .IN2(g1744), .Q(n4770) );
  AND2X1 U5081 ( .IN1(n4758), .IN2(g1776), .Q(n4769) );
  OR2X1 U5082 ( .IN1(n4771), .IN2(n4772), .Q(g4238) );
  AND2X1 U5083 ( .IN1(n4757), .IN2(g1741), .Q(n4772) );
  AND2X1 U5084 ( .IN1(n4758), .IN2(test_so5), .Q(n4771) );
  OR2X1 U5085 ( .IN1(n4773), .IN2(n4774), .Q(g4231) );
  AND2X1 U5086 ( .IN1(n4757), .IN2(g1738), .Q(n4774) );
  AND2X1 U5087 ( .IN1(n4758), .IN2(g1766), .Q(n4773) );
  OR2X1 U5088 ( .IN1(n652), .IN2(n3042), .Q(g4089) );
  INVX0 U5089 ( .INP(g1700), .ZN(n652) );
  AND2X1 U5090 ( .IN1(g1700), .IN2(n3327), .Q(g4076) );
  AND2X1 U5091 ( .IN1(n4775), .IN2(n4776), .Q(g3381) );
  AND2X1 U5092 ( .IN1(g936), .IN2(g940), .Q(n4776) );
  AND2X1 U5093 ( .IN1(g932), .IN2(g928), .Q(n4775) );
  INVX0 U5094 ( .INP(g23), .ZN(g3327) );
  AND2X1 U5095 ( .IN1(n3365), .IN2(n3328), .Q(g2478) );
  OR2X1 U5096 ( .IN1(n4777), .IN2(n4778), .Q(g11647) );
  AND2X1 U5097 ( .IN1(n4374), .IN2(n4779), .Q(n4778) );
  OR2X1 U5098 ( .IN1(n4780), .IN2(n4781), .Q(n4779) );
  AND2X1 U5099 ( .IN1(n4782), .IN2(n4783), .Q(n4781) );
  AND2X1 U5100 ( .IN1(n4784), .IN2(n4785), .Q(n4780) );
  AND2X1 U5101 ( .IN1(n3585), .IN2(g336), .Q(n4777) );
  AND2X1 U5102 ( .IN1(n4786), .IN2(n4787), .Q(g11641) );
  INVX0 U5103 ( .INP(n4788), .ZN(n4786) );
  AND2X1 U5104 ( .IN1(n4789), .IN2(n4790), .Q(n4788) );
  OR2X1 U5105 ( .IN1(n1226), .IN2(n1721), .Q(n4790) );
  AND2X1 U5106 ( .IN1(n6), .IN2(n3380), .Q(n1226) );
  OR2X1 U5107 ( .IN1(n4791), .IN2(n3380), .Q(n4789) );
  AND2X1 U5108 ( .IN1(g1351), .IN2(n1229), .Q(n3380) );
  AND2X1 U5109 ( .IN1(n4792), .IN2(n4787), .Q(g11640) );
  OR2X1 U5110 ( .IN1(n4793), .IN2(n4794), .Q(n4792) );
  AND2X1 U5111 ( .IN1(n1232), .IN2(n1231), .Q(n4794) );
  AND2X1 U5112 ( .IN1(n4791), .IN2(g1346), .Q(n4793) );
  OR2X1 U5113 ( .IN1(n1227), .IN2(n4795), .Q(n4791) );
  INVX0 U5114 ( .INP(n1229), .ZN(n4795) );
  AND2X1 U5115 ( .IN1(g1341), .IN2(n4796), .Q(n1229) );
  AND2X1 U5116 ( .IN1(g1336), .IN2(g1346), .Q(n4796) );
  AND2X1 U5117 ( .IN1(n4797), .IN2(n4787), .Q(g11639) );
  AND2X1 U5118 ( .IN1(n4798), .IN2(n4799), .Q(n4797) );
  OR2X1 U5119 ( .IN1(n1231), .IN2(g1341), .Q(n4799) );
  OR2X1 U5120 ( .IN1(n3298), .IN2(n4800), .Q(n4798) );
  INVX0 U5121 ( .INP(n1231), .ZN(n4800) );
  AND2X1 U5122 ( .IN1(n4801), .IN2(n4787), .Q(g11636) );
  OR2X1 U5123 ( .IN1(n4802), .IN2(n4306), .Q(n4787) );
  AND2X1 U5124 ( .IN1(g109), .IN2(n3362), .Q(n4306) );
  AND2X1 U5125 ( .IN1(n4803), .IN2(g109), .Q(n4802) );
  OR2X1 U5126 ( .IN1(n4804), .IN2(n3036), .Q(n4803) );
  AND2X1 U5127 ( .IN1(n4805), .IN2(n4806), .Q(n4801) );
  OR2X1 U5128 ( .IN1(n6), .IN2(g1336), .Q(n4806) );
  INVX0 U5129 ( .INP(n1227), .ZN(n6) );
  OR2X1 U5130 ( .IN1(n3300), .IN2(n1227), .Q(n4805) );
  OR2X1 U5131 ( .IN1(n4807), .IN2(n4808), .Q(g11625) );
  AND2X1 U5132 ( .IN1(n4374), .IN2(n4809), .Q(n4808) );
  AND2X1 U5133 ( .IN1(n4810), .IN2(n4811), .Q(n4809) );
  OR2X1 U5134 ( .IN1(n4784), .IN2(n4783), .Q(n4811) );
  INVX0 U5135 ( .INP(n4812), .ZN(n4783) );
  INVX0 U5136 ( .INP(n4813), .ZN(n4784) );
  OR2X1 U5137 ( .IN1(n4812), .IN2(n4813), .Q(n4810) );
  AND2X1 U5138 ( .IN1(n4814), .IN2(n4815), .Q(n4813) );
  OR2X1 U5139 ( .IN1(n4816), .IN2(n4817), .Q(n4815) );
  INVX0 U5140 ( .INP(n4818), .ZN(n4814) );
  AND2X1 U5141 ( .IN1(n4817), .IN2(n4816), .Q(n4818) );
  AND2X1 U5142 ( .IN1(n4819), .IN2(n4820), .Q(n4816) );
  INVX0 U5143 ( .INP(n4821), .ZN(n4820) );
  AND2X1 U5144 ( .IN1(n4822), .IN2(n4823), .Q(n4821) );
  OR2X1 U5145 ( .IN1(n4823), .IN2(n4822), .Q(n4819) );
  OR2X1 U5146 ( .IN1(n4824), .IN2(n4825), .Q(n4822) );
  INVX0 U5147 ( .INP(n4826), .ZN(n4825) );
  OR2X1 U5148 ( .IN1(n4827), .IN2(n4828), .Q(n4826) );
  AND2X1 U5149 ( .IN1(n4828), .IN2(n4827), .Q(n4824) );
  AND2X1 U5150 ( .IN1(n4829), .IN2(n4830), .Q(n4827) );
  OR2X1 U5151 ( .IN1(n4831), .IN2(n4832), .Q(n4830) );
  INVX0 U5152 ( .INP(n4833), .ZN(n4829) );
  AND2X1 U5153 ( .IN1(n4832), .IN2(n4831), .Q(n4833) );
  INVX0 U5154 ( .INP(n4834), .ZN(n4831) );
  OR2X1 U5155 ( .IN1(n4835), .IN2(n4836), .Q(n4828) );
  INVX0 U5156 ( .INP(n4837), .ZN(n4836) );
  OR2X1 U5157 ( .IN1(n4838), .IN2(n4839), .Q(n4837) );
  AND2X1 U5158 ( .IN1(n4839), .IN2(n4838), .Q(n4835) );
  INVX0 U5159 ( .INP(n4840), .ZN(n4838) );
  AND2X1 U5160 ( .IN1(n4841), .IN2(n4842), .Q(n4823) );
  INVX0 U5161 ( .INP(n4843), .ZN(n4842) );
  AND2X1 U5162 ( .IN1(n4844), .IN2(n4845), .Q(n4843) );
  OR2X1 U5163 ( .IN1(n4845), .IN2(n4844), .Q(n4841) );
  OR2X1 U5164 ( .IN1(n4846), .IN2(n4847), .Q(n4844) );
  INVX0 U5165 ( .INP(n4848), .ZN(n4847) );
  OR2X1 U5166 ( .IN1(n4849), .IN2(n4850), .Q(n4848) );
  AND2X1 U5167 ( .IN1(n4850), .IN2(n4849), .Q(n4846) );
  INVX0 U5168 ( .INP(n4851), .ZN(n4849) );
  AND2X1 U5169 ( .IN1(n4852), .IN2(n4853), .Q(n4845) );
  OR2X1 U5170 ( .IN1(n4854), .IN2(n4855), .Q(n4853) );
  INVX0 U5171 ( .INP(n4856), .ZN(n4854) );
  OR2X1 U5172 ( .IN1(n4857), .IN2(n4856), .Q(n4852) );
  INVX0 U5173 ( .INP(n4855), .ZN(n4857) );
  OR2X1 U5174 ( .IN1(n4858), .IN2(n4859), .Q(n4812) );
  AND2X1 U5175 ( .IN1(n4860), .IN2(n1239), .Q(n4859) );
  OR2X1 U5176 ( .IN1(n4861), .IN2(n4862), .Q(n4860) );
  AND2X1 U5177 ( .IN1(n4863), .IN2(n4864), .Q(n4862) );
  INVX0 U5178 ( .INP(n4865), .ZN(n4861) );
  OR2X1 U5179 ( .IN1(n4864), .IN2(n4863), .Q(n4865) );
  OR2X1 U5180 ( .IN1(n4866), .IN2(g471), .Q(n4864) );
  AND2X1 U5181 ( .IN1(n51), .IN2(g305), .Q(n4858) );
  AND2X1 U5182 ( .IN1(n3585), .IN2(g345), .Q(n4807) );
  OR2X1 U5183 ( .IN1(n4867), .IN2(n4868), .Q(g11610) );
  AND2X1 U5184 ( .IN1(n4869), .IN2(g1333), .Q(n4868) );
  AND2X1 U5185 ( .IN1(n4870), .IN2(g1806), .Q(n4867) );
  OR2X1 U5186 ( .IN1(n4871), .IN2(n4872), .Q(g11609) );
  AND2X1 U5187 ( .IN1(n4869), .IN2(g1330), .Q(n4872) );
  AND2X1 U5188 ( .IN1(n4870), .IN2(g1801), .Q(n4871) );
  OR2X1 U5189 ( .IN1(n4873), .IN2(n4874), .Q(g11608) );
  AND2X1 U5190 ( .IN1(n4869), .IN2(g1327), .Q(n4874) );
  AND2X1 U5191 ( .IN1(n4870), .IN2(g1796), .Q(n4873) );
  OR2X1 U5192 ( .IN1(n4875), .IN2(n4876), .Q(g11607) );
  AND2X1 U5193 ( .IN1(n4869), .IN2(g1324), .Q(n4876) );
  AND2X1 U5194 ( .IN1(n4870), .IN2(g1791), .Q(n4875) );
  OR2X1 U5195 ( .IN1(n4877), .IN2(n4878), .Q(g11606) );
  AND2X1 U5196 ( .IN1(n4869), .IN2(g1321), .Q(n4878) );
  AND2X1 U5197 ( .IN1(n4870), .IN2(g1786), .Q(n4877) );
  OR2X1 U5198 ( .IN1(n4879), .IN2(n4880), .Q(g11605) );
  AND2X1 U5199 ( .IN1(n4869), .IN2(g1318), .Q(n4880) );
  AND2X1 U5200 ( .IN1(n4870), .IN2(g1781), .Q(n4879) );
  OR2X1 U5201 ( .IN1(n4881), .IN2(n4882), .Q(g11604) );
  AND2X1 U5202 ( .IN1(n4869), .IN2(g1314), .Q(n4882) );
  AND2X1 U5203 ( .IN1(n4870), .IN2(g1776), .Q(n4881) );
  OR2X1 U5204 ( .IN1(n4883), .IN2(n4884), .Q(g11603) );
  AND2X1 U5205 ( .IN1(n4870), .IN2(test_so5), .Q(n4884) );
  AND2X1 U5206 ( .IN1(test_so9), .IN2(n4869), .Q(n4883) );
  OR2X1 U5207 ( .IN1(n4885), .IN2(n4886), .Q(g11602) );
  AND2X1 U5208 ( .IN1(n4869), .IN2(g1308), .Q(n4886) );
  AND2X1 U5209 ( .IN1(n4870), .IN2(g1766), .Q(n4885) );
  INVX0 U5210 ( .INP(n4869), .ZN(n4870) );
  OR2X1 U5211 ( .IN1(n3369), .IN2(n1227), .Q(n4869) );
  OR2X1 U5212 ( .IN1(n4310), .IN2(n4887), .Q(n1227) );
  OR2X1 U5213 ( .IN1(n4888), .IN2(n4889), .Q(n4887) );
  AND2X1 U5214 ( .IN1(n4890), .IN2(n4891), .Q(n4888) );
  AND2X1 U5215 ( .IN1(n4892), .IN2(n4893), .Q(n4891) );
  AND2X1 U5216 ( .IN1(n4894), .IN2(n4895), .Q(n4893) );
  OR2X1 U5217 ( .IN1(n4896), .IN2(n4897), .Q(n4895) );
  AND2X1 U5218 ( .IN1(n3228), .IN2(n3385), .Q(n4897) );
  AND2X1 U5219 ( .IN1(test_so2), .IN2(g1255), .Q(n4896) );
  AND2X1 U5220 ( .IN1(n4898), .IN2(n4899), .Q(n4894) );
  OR2X1 U5221 ( .IN1(n4900), .IN2(n4901), .Q(n4899) );
  AND2X1 U5222 ( .IN1(n3200), .IN2(n3384), .Q(n4901) );
  AND2X1 U5223 ( .IN1(test_so6), .IN2(g1023), .Q(n4900) );
  OR2X1 U5224 ( .IN1(n4902), .IN2(n4903), .Q(n4898) );
  AND2X1 U5225 ( .IN1(n4904), .IN2(n4905), .Q(n4903) );
  AND2X1 U5226 ( .IN1(n4906), .IN2(n4907), .Q(n4902) );
  INVX0 U5227 ( .INP(n4904), .ZN(n4907) );
  AND2X1 U5228 ( .IN1(n4908), .IN2(n4909), .Q(n4892) );
  OR2X1 U5229 ( .IN1(n4910), .IN2(n4911), .Q(n4909) );
  AND2X1 U5230 ( .IN1(n3253), .IN2(n3386), .Q(n4911) );
  AND2X1 U5231 ( .IN1(test_so8), .IN2(g1245), .Q(n4910) );
  AND2X1 U5232 ( .IN1(n4912), .IN2(n4913), .Q(n4908) );
  OR2X1 U5233 ( .IN1(n3255), .IN2(g1250), .Q(n4913) );
  OR2X1 U5234 ( .IN1(n3256), .IN2(g1011), .Q(n4912) );
  AND2X1 U5235 ( .IN1(n4914), .IN2(n4915), .Q(n4890) );
  AND2X1 U5236 ( .IN1(n4916), .IN2(n4917), .Q(n4915) );
  AND2X1 U5237 ( .IN1(n4918), .IN2(n4919), .Q(n4917) );
  OR2X1 U5238 ( .IN1(n3221), .IN2(g1260), .Q(n4919) );
  OR2X1 U5239 ( .IN1(n3229), .IN2(g1019), .Q(n4918) );
  AND2X1 U5240 ( .IN1(n4920), .IN2(n4921), .Q(n4916) );
  AND2X1 U5241 ( .IN1(n4922), .IN2(n4923), .Q(n4921) );
  OR2X1 U5242 ( .IN1(n1871), .IN2(g1235), .Q(n4923) );
  OR2X1 U5243 ( .IN1(n3254), .IN2(g991), .Q(n4922) );
  AND2X1 U5244 ( .IN1(n4924), .IN2(n4925), .Q(n4920) );
  OR2X1 U5245 ( .IN1(n3290), .IN2(g995), .Q(n4925) );
  OR2X1 U5246 ( .IN1(n3291), .IN2(g1275), .Q(n4924) );
  AND2X1 U5247 ( .IN1(n4926), .IN2(n4927), .Q(n4914) );
  AND2X1 U5248 ( .IN1(n4928), .IN2(n4929), .Q(n4927) );
  OR2X1 U5249 ( .IN1(n3292), .IN2(g1003), .Q(n4929) );
  OR2X1 U5250 ( .IN1(n3293), .IN2(g1240), .Q(n4928) );
  AND2X1 U5251 ( .IN1(n4930), .IN2(n4931), .Q(n4926) );
  OR2X1 U5252 ( .IN1(n3220), .IN2(g1265), .Q(n4931) );
  OR2X1 U5253 ( .IN1(n3231), .IN2(g1015), .Q(n4930) );
  OR2X1 U5254 ( .IN1(n4932), .IN2(n4933), .Q(g11579) );
  AND2X1 U5255 ( .IN1(n4934), .IN2(n3946), .Q(n4933) );
  AND2X1 U5256 ( .IN1(n4935), .IN2(n4936), .Q(n4934) );
  OR2X1 U5257 ( .IN1(g1610), .IN2(n4937), .Q(n4936) );
  INVX0 U5258 ( .INP(n4938), .ZN(n4935) );
  AND2X1 U5259 ( .IN1(g1610), .IN2(n4937), .Q(n4938) );
  OR2X1 U5260 ( .IN1(n4939), .IN2(n4940), .Q(n4937) );
  AND2X1 U5261 ( .IN1(n1260), .IN2(n4941), .Q(n4940) );
  AND2X1 U5262 ( .IN1(n4942), .IN2(n4943), .Q(n4939) );
  OR2X1 U5263 ( .IN1(n1258), .IN2(n4944), .Q(n4943) );
  INVX0 U5264 ( .INP(n1262), .ZN(n4944) );
  OR2X1 U5265 ( .IN1(n4945), .IN2(n4946), .Q(n1262) );
  AND2X1 U5266 ( .IN1(n4946), .IN2(n4945), .Q(n1258) );
  INVX0 U5267 ( .INP(n4947), .ZN(n4945) );
  OR2X1 U5268 ( .IN1(n4948), .IN2(n4949), .Q(n4947) );
  AND2X1 U5269 ( .IN1(n1685), .IN2(n4950), .Q(n4949) );
  OR2X1 U5270 ( .IN1(n4951), .IN2(g1153), .Q(n4950) );
  AND2X1 U5271 ( .IN1(n4952), .IN2(n4953), .Q(n4951) );
  AND2X1 U5272 ( .IN1(n4954), .IN2(n4955), .Q(n4953) );
  AND2X1 U5273 ( .IN1(n4956), .IN2(n4957), .Q(n4955) );
  AND2X1 U5274 ( .IN1(n1597), .IN2(n3387), .Q(n4957) );
  AND2X1 U5275 ( .IN1(n1618), .IN2(n1617), .Q(n4956) );
  AND2X1 U5276 ( .IN1(n4958), .IN2(n1706), .Q(n4954) );
  AND2X1 U5277 ( .IN1(n1705), .IN2(n1660), .Q(n4958) );
  AND2X1 U5278 ( .IN1(n4959), .IN2(n4960), .Q(n4952) );
  AND2X1 U5279 ( .IN1(n4961), .IN2(n3264), .Q(n4960) );
  AND2X1 U5280 ( .IN1(n3263), .IN2(n1708), .Q(n4961) );
  AND2X1 U5281 ( .IN1(n4962), .IN2(n6001), .Q(n4959) );
  AND2X1 U5282 ( .IN1(n3266), .IN2(n3265), .Q(n4962) );
  AND2X1 U5283 ( .IN1(n1686), .IN2(g1149), .Q(n4948) );
  OR2X1 U5284 ( .IN1(n4015), .IN2(n3984), .Q(n4946) );
  OR2X1 U5285 ( .IN1(n1654), .IN2(g1110), .Q(n3984) );
  OR2X1 U5286 ( .IN1(g1107), .IN2(g1104), .Q(n4015) );
  AND2X1 U5287 ( .IN1(n495), .IN2(g1618), .Q(n4932) );
  AND2X1 U5288 ( .IN1(n4963), .IN2(n4964), .Q(g11514) );
  OR2X1 U5289 ( .IN1(n4965), .IN2(n4966), .Q(n4964) );
  AND2X1 U5290 ( .IN1(n4967), .IN2(n4968), .Q(n4966) );
  OR2X1 U5291 ( .IN1(g1419), .IN2(n4942), .Q(n4968) );
  OR2X1 U5292 ( .IN1(n1602), .IN2(n4941), .Q(n4967) );
  OR2X1 U5293 ( .IN1(n4969), .IN2(n4970), .Q(n4963) );
  AND2X1 U5294 ( .IN1(g6193), .IN2(n4942), .Q(n4970) );
  AND2X1 U5295 ( .IN1(g1419), .IN2(g109), .Q(g6193) );
  AND2X1 U5296 ( .IN1(n4971), .IN2(g109), .Q(n4969) );
  OR2X1 U5297 ( .IN1(n4972), .IN2(n4973), .Q(n4971) );
  INVX0 U5298 ( .INP(n4965), .ZN(n4973) );
  AND2X1 U5299 ( .IN1(n4974), .IN2(n4975), .Q(n4965) );
  OR2X1 U5300 ( .IN1(n1627), .IN2(n4976), .Q(n4975) );
  AND2X1 U5301 ( .IN1(n4977), .IN2(n4978), .Q(n4976) );
  OR2X1 U5302 ( .IN1(n3136), .IN2(g1448), .Q(n4978) );
  OR2X1 U5303 ( .IN1(n3250), .IN2(g1415), .Q(n4977) );
  OR2X1 U5304 ( .IN1(g1515), .IN2(n4979), .Q(n4974) );
  OR2X1 U5305 ( .IN1(n4980), .IN2(n4981), .Q(n4979) );
  AND2X1 U5306 ( .IN1(n3136), .IN2(g1448), .Q(n4981) );
  AND2X1 U5307 ( .IN1(n3250), .IN2(g1415), .Q(n4980) );
  AND2X1 U5308 ( .IN1(n1602), .IN2(n4941), .Q(n4972) );
  INVX0 U5309 ( .INP(n4942), .ZN(n4941) );
  OR2X1 U5310 ( .IN1(n4982), .IN2(n4983), .Q(n4942) );
  AND2X1 U5311 ( .IN1(n4984), .IN2(n3963), .Q(n4983) );
  OR2X1 U5312 ( .IN1(n4985), .IN2(n4986), .Q(n4984) );
  AND2X1 U5313 ( .IN1(n4987), .IN2(n4988), .Q(n4986) );
  OR2X1 U5314 ( .IN1(g10726), .IN2(n4989), .Q(n4987) );
  INVX0 U5315 ( .INP(n4990), .ZN(n4985) );
  OR2X1 U5316 ( .IN1(n4988), .IN2(g1811), .Q(n4990) );
  OR2X1 U5317 ( .IN1(n4991), .IN2(n4992), .Q(n4988) );
  OR2X1 U5318 ( .IN1(n3029), .IN2(n3023), .Q(n4992) );
  OR2X1 U5319 ( .IN1(n3017), .IN2(n3065), .Q(n4991) );
  AND2X1 U5320 ( .IN1(g18), .IN2(g201), .Q(n4982) );
  OR2X1 U5321 ( .IN1(n4993), .IN2(n4994), .Q(g11488) );
  AND2X1 U5322 ( .IN1(n4374), .IN2(n4851), .Q(n4994) );
  OR2X1 U5323 ( .IN1(n4995), .IN2(n4996), .Q(n4851) );
  AND2X1 U5324 ( .IN1(n4997), .IN2(n1239), .Q(n4996) );
  OR2X1 U5325 ( .IN1(n4998), .IN2(n4999), .Q(n4997) );
  INVX0 U5326 ( .INP(n5000), .ZN(n4999) );
  OR2X1 U5327 ( .IN1(n5001), .IN2(g516), .Q(n5000) );
  AND2X1 U5328 ( .IN1(n5001), .IN2(g516), .Q(n4998) );
  OR2X1 U5329 ( .IN1(n4866), .IN2(n1606), .Q(n5001) );
  OR2X1 U5330 ( .IN1(g466), .IN2(n5002), .Q(n4866) );
  OR2X1 U5331 ( .IN1(n1641), .IN2(g461), .Q(n5002) );
  AND2X1 U5332 ( .IN1(n51), .IN2(g309), .Q(n4995) );
  AND2X1 U5333 ( .IN1(n3585), .IN2(g342), .Q(n4993) );
  OR2X1 U5334 ( .IN1(n5003), .IN2(n5004), .Q(g11487) );
  AND2X1 U5335 ( .IN1(n4374), .IN2(n4850), .Q(n5004) );
  OR2X1 U5336 ( .IN1(n5005), .IN2(n5006), .Q(n4850) );
  AND2X1 U5337 ( .IN1(n5007), .IN2(n1239), .Q(n5006) );
  OR2X1 U5338 ( .IN1(n5008), .IN2(n5009), .Q(n5007) );
  AND2X1 U5339 ( .IN1(n5010), .IN2(n1679), .Q(n5009) );
  AND2X1 U5340 ( .IN1(n5011), .IN2(n1594), .Q(n5010) );
  AND2X1 U5341 ( .IN1(n5012), .IN2(g511), .Q(n5008) );
  OR2X1 U5342 ( .IN1(g461), .IN2(n5013), .Q(n5012) );
  AND2X1 U5343 ( .IN1(n51), .IN2(g333), .Q(n5005) );
  AND2X1 U5344 ( .IN1(n3585), .IN2(g366), .Q(n5003) );
  OR2X1 U5345 ( .IN1(n5014), .IN2(n5015), .Q(g11486) );
  AND2X1 U5346 ( .IN1(n4374), .IN2(n4856), .Q(n5015) );
  OR2X1 U5347 ( .IN1(n5016), .IN2(n5017), .Q(n4856) );
  AND2X1 U5348 ( .IN1(n5018), .IN2(n1239), .Q(n5017) );
  OR2X1 U5349 ( .IN1(n5019), .IN2(n5020), .Q(n5018) );
  AND2X1 U5350 ( .IN1(n5021), .IN2(n1600), .Q(n5020) );
  AND2X1 U5351 ( .IN1(n5022), .IN2(n1606), .Q(n5021) );
  AND2X1 U5352 ( .IN1(n5023), .IN2(g506), .Q(n5019) );
  OR2X1 U5353 ( .IN1(g471), .IN2(n5024), .Q(n5023) );
  AND2X1 U5354 ( .IN1(n51), .IN2(g330), .Q(n5016) );
  AND2X1 U5355 ( .IN1(n3585), .IN2(g363), .Q(n5014) );
  OR2X1 U5356 ( .IN1(n5025), .IN2(n5026), .Q(g11485) );
  AND2X1 U5357 ( .IN1(n4374), .IN2(n4840), .Q(n5026) );
  OR2X1 U5358 ( .IN1(n5027), .IN2(n5028), .Q(n4840) );
  AND2X1 U5359 ( .IN1(n5029), .IN2(n1239), .Q(n5028) );
  OR2X1 U5360 ( .IN1(n5030), .IN2(n5031), .Q(n5029) );
  AND2X1 U5361 ( .IN1(n5032), .IN2(n1690), .Q(n5031) );
  AND2X1 U5362 ( .IN1(n5033), .IN2(g461), .Q(n5032) );
  AND2X1 U5363 ( .IN1(n5034), .IN2(g501), .Q(n5030) );
  OR2X1 U5364 ( .IN1(n1594), .IN2(n5035), .Q(n5034) );
  AND2X1 U5365 ( .IN1(n51), .IN2(g327), .Q(n5027) );
  AND2X1 U5366 ( .IN1(n3585), .IN2(g360), .Q(n5025) );
  OR2X1 U5367 ( .IN1(n5036), .IN2(n5037), .Q(g11484) );
  AND2X1 U5368 ( .IN1(n4374), .IN2(n4839), .Q(n5037) );
  OR2X1 U5369 ( .IN1(n5038), .IN2(n5039), .Q(n4839) );
  AND2X1 U5370 ( .IN1(n5040), .IN2(n1239), .Q(n5039) );
  AND2X1 U5371 ( .IN1(n5041), .IN2(n5042), .Q(n5040) );
  OR2X1 U5372 ( .IN1(n5043), .IN2(g496), .Q(n5042) );
  INVX0 U5373 ( .INP(n5044), .ZN(n5043) );
  OR2X1 U5374 ( .IN1(n1689), .IN2(n5044), .Q(n5041) );
  OR2X1 U5375 ( .IN1(n5045), .IN2(n5046), .Q(n5044) );
  OR2X1 U5376 ( .IN1(g461), .IN2(g471), .Q(n5046) );
  AND2X1 U5377 ( .IN1(n51), .IN2(g324), .Q(n5038) );
  AND2X1 U5378 ( .IN1(n3585), .IN2(g357), .Q(n5036) );
  OR2X1 U5379 ( .IN1(n5047), .IN2(n5048), .Q(g11483) );
  AND2X1 U5380 ( .IN1(n4374), .IN2(n4834), .Q(n5048) );
  OR2X1 U5381 ( .IN1(n5049), .IN2(n5050), .Q(n4834) );
  AND2X1 U5382 ( .IN1(n5051), .IN2(n1239), .Q(n5050) );
  OR2X1 U5383 ( .IN1(n5052), .IN2(n5053), .Q(n5051) );
  AND2X1 U5384 ( .IN1(n5054), .IN2(n1691), .Q(n5053) );
  AND2X1 U5385 ( .IN1(n5033), .IN2(n1594), .Q(n5054) );
  INVX0 U5386 ( .INP(n5035), .ZN(n5033) );
  AND2X1 U5387 ( .IN1(n5055), .IN2(g491), .Q(n5052) );
  OR2X1 U5388 ( .IN1(g461), .IN2(n5035), .Q(n5055) );
  OR2X1 U5389 ( .IN1(g456), .IN2(n5056), .Q(n5035) );
  OR2X1 U5390 ( .IN1(n1646), .IN2(g471), .Q(n5056) );
  AND2X1 U5391 ( .IN1(n51), .IN2(g321), .Q(n5049) );
  AND2X1 U5392 ( .IN1(n3585), .IN2(g354), .Q(n5047) );
  OR2X1 U5393 ( .IN1(n5057), .IN2(n5058), .Q(g11482) );
  AND2X1 U5394 ( .IN1(n4374), .IN2(n4817), .Q(n5058) );
  OR2X1 U5395 ( .IN1(n5059), .IN2(n5060), .Q(n4817) );
  AND2X1 U5396 ( .IN1(n5061), .IN2(n1239), .Q(n5060) );
  OR2X1 U5397 ( .IN1(n5062), .IN2(n5063), .Q(n5061) );
  AND2X1 U5398 ( .IN1(n5064), .IN2(n1621), .Q(n5063) );
  AND2X1 U5399 ( .IN1(n5065), .IN2(g456), .Q(n5064) );
  AND2X1 U5400 ( .IN1(n5066), .IN2(g486), .Q(n5062) );
  OR2X1 U5401 ( .IN1(n1641), .IN2(n5067), .Q(n5066) );
  AND2X1 U5402 ( .IN1(n51), .IN2(g318), .Q(n5059) );
  AND2X1 U5403 ( .IN1(n3585), .IN2(g351), .Q(n5057) );
  OR2X1 U5404 ( .IN1(n5068), .IN2(n5069), .Q(g11481) );
  AND2X1 U5405 ( .IN1(n4374), .IN2(n4832), .Q(n5069) );
  OR2X1 U5406 ( .IN1(n5070), .IN2(n5071), .Q(n4832) );
  AND2X1 U5407 ( .IN1(n5072), .IN2(n1239), .Q(n5071) );
  OR2X1 U5408 ( .IN1(n5073), .IN2(n5074), .Q(n5072) );
  AND2X1 U5409 ( .IN1(n5075), .IN2(n1680), .Q(n5074) );
  AND2X1 U5410 ( .IN1(n1641), .IN2(n5065), .Q(n5075) );
  INVX0 U5411 ( .INP(n5067), .ZN(n5065) );
  AND2X1 U5412 ( .IN1(n5076), .IN2(g481), .Q(n5073) );
  OR2X1 U5413 ( .IN1(n5067), .IN2(g456), .Q(n5076) );
  OR2X1 U5414 ( .IN1(g471), .IN2(n5077), .Q(n5067) );
  OR2X1 U5415 ( .IN1(n1594), .IN2(g466), .Q(n5077) );
  AND2X1 U5416 ( .IN1(n51), .IN2(g315), .Q(n5070) );
  AND2X1 U5417 ( .IN1(n3585), .IN2(g348), .Q(n5068) );
  OR2X1 U5418 ( .IN1(n5078), .IN2(n5079), .Q(g11478) );
  AND2X1 U5419 ( .IN1(n4374), .IN2(n4855), .Q(n5079) );
  OR2X1 U5420 ( .IN1(n5080), .IN2(n5081), .Q(n4855) );
  AND2X1 U5421 ( .IN1(n5082), .IN2(n1239), .Q(n5081) );
  OR2X1 U5422 ( .IN1(n5083), .IN2(n5084), .Q(n5082) );
  AND2X1 U5423 ( .IN1(n5085), .IN2(n1599), .Q(n5084) );
  AND2X1 U5424 ( .IN1(n5011), .IN2(g461), .Q(n5085) );
  INVX0 U5425 ( .INP(n5013), .ZN(n5011) );
  AND2X1 U5426 ( .IN1(n5086), .IN2(g476), .Q(n5083) );
  OR2X1 U5427 ( .IN1(n1594), .IN2(n5013), .Q(n5086) );
  OR2X1 U5428 ( .IN1(g456), .IN2(n5087), .Q(n5013) );
  OR2X1 U5429 ( .IN1(n1606), .IN2(g466), .Q(n5087) );
  AND2X1 U5430 ( .IN1(n51), .IN2(g312), .Q(n5080) );
  AND2X1 U5431 ( .IN1(n3585), .IN2(g339), .Q(n5078) );
  INVX0 U5432 ( .INP(n4374), .ZN(n3585) );
  AND2X1 U5433 ( .IN1(g750), .IN2(n1647), .Q(n4374) );
  OR2X1 U5434 ( .IN1(n5088), .IN2(n5089), .Q(g11443) );
  AND2X1 U5435 ( .IN1(n4343), .IN2(g1275), .Q(n5089) );
  AND2X1 U5436 ( .IN1(g109), .IN2(n4310), .Q(n4343) );
  AND2X1 U5437 ( .IN1(n4342), .IN2(n4904), .Q(n5088) );
  OR2X1 U5438 ( .IN1(n5090), .IN2(n5091), .Q(n4904) );
  AND2X1 U5439 ( .IN1(n5092), .IN2(n4327), .Q(n5091) );
  INVX0 U5440 ( .INP(n4889), .ZN(n4327) );
  OR2X1 U5441 ( .IN1(n5093), .IN2(n5094), .Q(n5092) );
  AND2X1 U5442 ( .IN1(n1862), .IN2(n5095), .Q(n5094) );
  OR2X1 U5443 ( .IN1(n5096), .IN2(g1284), .Q(n5095) );
  AND2X1 U5444 ( .IN1(n5097), .IN2(n5098), .Q(n5096) );
  AND2X1 U5445 ( .IN1(n5099), .IN2(n5100), .Q(n5098) );
  AND2X1 U5446 ( .IN1(n5101), .IN2(n5102), .Q(n5100) );
  AND2X1 U5447 ( .IN1(n3228), .IN2(n3384), .Q(n5102) );
  AND2X1 U5448 ( .IN1(n3231), .IN2(n3229), .Q(n5101) );
  AND2X1 U5449 ( .IN1(n5103), .IN2(n3234), .Q(n5099) );
  AND2X1 U5450 ( .IN1(n3233), .IN2(n3232), .Q(n5103) );
  AND2X1 U5451 ( .IN1(n5104), .IN2(n5105), .Q(n5097) );
  AND2X1 U5452 ( .IN1(n5106), .IN2(n3254), .Q(n5105) );
  AND2X1 U5453 ( .IN1(n3253), .IN2(n3235), .Q(n5106) );
  AND2X1 U5454 ( .IN1(n5107), .IN2(n3292), .Q(n5104) );
  AND2X1 U5455 ( .IN1(n3290), .IN2(n3256), .Q(n5107) );
  AND2X1 U5456 ( .IN1(n1864), .IN2(g1280), .Q(n5093) );
  AND2X1 U5457 ( .IN1(n4905), .IN2(n4889), .Q(n5090) );
  OR2X1 U5458 ( .IN1(n3361), .IN2(n4325), .Q(n4889) );
  OR2X1 U5459 ( .IN1(n3129), .IN2(n5108), .Q(n4325) );
  OR2X1 U5460 ( .IN1(n3367), .IN2(n3130), .Q(n5108) );
  INVX0 U5461 ( .INP(n4906), .ZN(n4905) );
  OR2X1 U5462 ( .IN1(n5109), .IN2(n5110), .Q(n4906) );
  AND2X1 U5463 ( .IN1(n5111), .IN2(g1027), .Q(n5110) );
  AND2X1 U5464 ( .IN1(n4785), .IN2(g1032), .Q(n5111) );
  AND2X1 U5465 ( .IN1(n3324), .IN2(n5112), .Q(n5109) );
  OR2X1 U5466 ( .IN1(n3368), .IN2(n4782), .Q(n5112) );
  INVX0 U5467 ( .INP(n4310), .ZN(n4342) );
  OR2X1 U5468 ( .IN1(g1713), .IN2(n5113), .Q(n4310) );
  OR2X1 U5469 ( .IN1(n3323), .IN2(n495), .Q(n5113) );
  AND2X1 U5470 ( .IN1(n5114), .IN2(n5115), .Q(g11393) );
  OR2X1 U5471 ( .IN1(n5116), .IN2(n3587), .Q(n5115) );
  OR2X1 U5472 ( .IN1(n1722), .IN2(n5117), .Q(n3587) );
  AND2X1 U5473 ( .IN1(n5118), .IN2(n5119), .Q(n5114) );
  OR2X1 U5474 ( .IN1(n5120), .IN2(g986), .Q(n5118) );
  INVX0 U5475 ( .INP(n5121), .ZN(n5120) );
  AND2X1 U5476 ( .IN1(n5122), .IN2(n5119), .Q(g11392) );
  OR2X1 U5477 ( .IN1(n5123), .IN2(n5124), .Q(n5122) );
  AND2X1 U5478 ( .IN1(n5125), .IN2(n5117), .Q(n5124) );
  INVX0 U5479 ( .INP(n5126), .ZN(n5125) );
  AND2X1 U5480 ( .IN1(n5121), .IN2(g981), .Q(n5123) );
  OR2X1 U5481 ( .IN1(n5117), .IN2(n5116), .Q(n5121) );
  OR2X1 U5482 ( .IN1(n1720), .IN2(n5127), .Q(n5117) );
  AND2X1 U5483 ( .IN1(n5128), .IN2(n5129), .Q(g11391) );
  OR2X1 U5484 ( .IN1(n5130), .IN2(g976), .Q(n5129) );
  AND2X1 U5485 ( .IN1(n19), .IN2(g971), .Q(n5130) );
  AND2X1 U5486 ( .IN1(n5126), .IN2(n5119), .Q(n5128) );
  OR2X1 U5487 ( .IN1(n5116), .IN2(n5127), .Q(n5126) );
  OR2X1 U5488 ( .IN1(n3372), .IN2(n3371), .Q(n5127) );
  AND2X1 U5489 ( .IN1(n5131), .IN2(n5132), .Q(g11380) );
  OR2X1 U5490 ( .IN1(n5133), .IN2(g471), .Q(n5132) );
  AND2X1 U5491 ( .IN1(n5134), .IN2(n5022), .Q(n5133) );
  AND2X1 U5492 ( .IN1(n5131), .IN2(n5135), .Q(g11376) );
  OR2X1 U5493 ( .IN1(n5136), .IN2(n5137), .Q(n5135) );
  AND2X1 U5494 ( .IN1(n5138), .IN2(g466), .Q(n5137) );
  OR2X1 U5495 ( .IN1(n5024), .IN2(n5139), .Q(n5138) );
  AND2X1 U5496 ( .IN1(n5140), .IN2(n5141), .Q(n5136) );
  AND2X1 U5497 ( .IN1(g461), .IN2(g456), .Q(n5141) );
  AND2X1 U5498 ( .IN1(n5134), .IN2(n5024), .Q(n5140) );
  AND2X1 U5499 ( .IN1(n5142), .IN2(n5131), .Q(g11372) );
  AND2X1 U5500 ( .IN1(n5143), .IN2(n5144), .Q(n5142) );
  OR2X1 U5501 ( .IN1(n5145), .IN2(g461), .Q(n5144) );
  OR2X1 U5502 ( .IN1(n1594), .IN2(n5146), .Q(n5143) );
  INVX0 U5503 ( .INP(n5145), .ZN(n5146) );
  AND2X1 U5504 ( .IN1(g456), .IN2(n5134), .Q(n5145) );
  AND2X1 U5505 ( .IN1(n5147), .IN2(n5119), .Q(g11349) );
  OR2X1 U5506 ( .IN1(n5148), .IN2(n3377), .Q(n5119) );
  AND2X1 U5507 ( .IN1(g109), .IN2(n5149), .Q(n3377) );
  OR2X1 U5508 ( .IN1(n3064), .IN2(n5150), .Q(n5149) );
  AND2X1 U5509 ( .IN1(g3007), .IN2(n6002), .Q(n5150) );
  AND2X1 U5510 ( .IN1(n5151), .IN2(n5152), .Q(n5147) );
  OR2X1 U5511 ( .IN1(n19), .IN2(g971), .Q(n5152) );
  INVX0 U5512 ( .INP(n5116), .ZN(n19) );
  OR2X1 U5513 ( .IN1(n3371), .IN2(n5116), .Q(n5151) );
  OR2X1 U5514 ( .IN1(n5153), .IN2(n5154), .Q(n5116) );
  OR2X1 U5515 ( .IN1(n51), .IN2(n5155), .Q(n5154) );
  AND2X1 U5516 ( .IN1(n5156), .IN2(n5157), .Q(n5155) );
  AND2X1 U5517 ( .IN1(n5158), .IN2(n5159), .Q(n5157) );
  AND2X1 U5518 ( .IN1(n5160), .IN2(n5161), .Q(n5159) );
  AND2X1 U5519 ( .IN1(n5162), .IN2(n5163), .Q(n5161) );
  OR2X1 U5520 ( .IN1(n3276), .IN2(g421), .Q(n5163) );
  OR2X1 U5521 ( .IN1(n3277), .IN2(g312), .Q(n5162) );
  AND2X1 U5522 ( .IN1(n5164), .IN2(n5165), .Q(n5160) );
  AND2X1 U5523 ( .IN1(n5166), .IN2(n5167), .Q(n5165) );
  OR2X1 U5524 ( .IN1(n3278), .IN2(g411), .Q(n5167) );
  OR2X1 U5525 ( .IN1(n3279), .IN2(g333), .Q(n5166) );
  AND2X1 U5526 ( .IN1(n5168), .IN2(n5169), .Q(n5164) );
  OR2X1 U5527 ( .IN1(n3261), .IN2(g401), .Q(n5169) );
  OR2X1 U5528 ( .IN1(n3262), .IN2(g327), .Q(n5168) );
  AND2X1 U5529 ( .IN1(n5170), .IN2(n5171), .Q(n5158) );
  AND2X1 U5530 ( .IN1(n5172), .IN2(n5173), .Q(n5171) );
  OR2X1 U5531 ( .IN1(n3085), .IN2(g416), .Q(n5173) );
  OR2X1 U5532 ( .IN1(n3236), .IN2(g309), .Q(n5172) );
  AND2X1 U5533 ( .IN1(n5174), .IN2(n5175), .Q(n5170) );
  OR2X1 U5534 ( .IN1(g305), .IN2(n5176), .Q(n5175) );
  OR2X1 U5535 ( .IN1(n1681), .IN2(n5177), .Q(n5174) );
  AND2X1 U5536 ( .IN1(n5178), .IN2(n5179), .Q(n5156) );
  AND2X1 U5537 ( .IN1(n5180), .IN2(n5181), .Q(n5179) );
  AND2X1 U5538 ( .IN1(n5182), .IN2(n5183), .Q(n5181) );
  OR2X1 U5539 ( .IN1(n3257), .IN2(g396), .Q(n5183) );
  OR2X1 U5540 ( .IN1(n3258), .IN2(g324), .Q(n5182) );
  AND2X1 U5541 ( .IN1(n5184), .IN2(n5185), .Q(n5180) );
  AND2X1 U5542 ( .IN1(n5186), .IN2(n5187), .Q(n5185) );
  OR2X1 U5543 ( .IN1(n3294), .IN2(g315), .Q(n5187) );
  OR2X1 U5544 ( .IN1(n3295), .IN2(g426), .Q(n5186) );
  AND2X1 U5545 ( .IN1(n5188), .IN2(n5189), .Q(n5184) );
  OR2X1 U5546 ( .IN1(n3084), .IN2(g406), .Q(n5189) );
  OR2X1 U5547 ( .IN1(n3230), .IN2(g330), .Q(n5188) );
  AND2X1 U5548 ( .IN1(n5190), .IN2(n5191), .Q(n5178) );
  AND2X1 U5549 ( .IN1(n5192), .IN2(n5193), .Q(n5191) );
  OR2X1 U5550 ( .IN1(n3296), .IN2(g321), .Q(n5193) );
  OR2X1 U5551 ( .IN1(n3297), .IN2(g391), .Q(n5192) );
  AND2X1 U5552 ( .IN1(n5194), .IN2(n5195), .Q(n5190) );
  OR2X1 U5553 ( .IN1(n3259), .IN2(g386), .Q(n5195) );
  OR2X1 U5554 ( .IN1(n3260), .IN2(g318), .Q(n5194) );
  AND2X1 U5555 ( .IN1(n5196), .IN2(n5131), .Q(g11340) );
  INVX0 U5556 ( .INP(n5197), .ZN(n5131) );
  OR2X1 U5557 ( .IN1(n650), .IN2(n3026), .Q(n5197) );
  AND2X1 U5558 ( .IN1(n5198), .IN2(n5199), .Q(n5196) );
  OR2X1 U5559 ( .IN1(n5134), .IN2(g456), .Q(n5199) );
  INVX0 U5560 ( .INP(n5139), .ZN(n5134) );
  OR2X1 U5561 ( .IN1(n1641), .IN2(n5139), .Q(n5198) );
  OR2X1 U5562 ( .IN1(n51), .IN2(n5200), .Q(n5139) );
  AND2X1 U5563 ( .IN1(n5022), .IN2(g471), .Q(n5200) );
  INVX0 U5564 ( .INP(n5024), .ZN(n5022) );
  OR2X1 U5565 ( .IN1(n1594), .IN2(n5045), .Q(n5024) );
  OR2X1 U5566 ( .IN1(n1646), .IN2(n1641), .Q(n5045) );
  OR2X1 U5567 ( .IN1(n5201), .IN2(n5202), .Q(g11338) );
  AND2X1 U5568 ( .IN1(n1239), .IN2(g516), .Q(n5202) );
  AND2X1 U5569 ( .IN1(n51), .IN2(g476), .Q(n5201) );
  OR2X1 U5570 ( .IN1(n5203), .IN2(n5204), .Q(g11337) );
  AND2X1 U5571 ( .IN1(n1239), .IN2(g511), .Q(n5204) );
  AND2X1 U5572 ( .IN1(n51), .IN2(g516), .Q(n5203) );
  OR2X1 U5573 ( .IN1(n5205), .IN2(n5206), .Q(g11336) );
  AND2X1 U5574 ( .IN1(n1239), .IN2(g506), .Q(n5206) );
  AND2X1 U5575 ( .IN1(n51), .IN2(g511), .Q(n5205) );
  OR2X1 U5576 ( .IN1(n5207), .IN2(n5208), .Q(g11335) );
  AND2X1 U5577 ( .IN1(n1239), .IN2(g501), .Q(n5208) );
  AND2X1 U5578 ( .IN1(n51), .IN2(g506), .Q(n5207) );
  OR2X1 U5579 ( .IN1(n5209), .IN2(n5210), .Q(g11334) );
  AND2X1 U5580 ( .IN1(n1239), .IN2(g496), .Q(n5210) );
  AND2X1 U5581 ( .IN1(n51), .IN2(g501), .Q(n5209) );
  OR2X1 U5582 ( .IN1(n5211), .IN2(n5212), .Q(g11333) );
  AND2X1 U5583 ( .IN1(n1239), .IN2(g491), .Q(n5212) );
  AND2X1 U5584 ( .IN1(n51), .IN2(g496), .Q(n5211) );
  OR2X1 U5585 ( .IN1(n5213), .IN2(n5214), .Q(g11332) );
  AND2X1 U5586 ( .IN1(n1239), .IN2(g486), .Q(n5214) );
  AND2X1 U5587 ( .IN1(n51), .IN2(g491), .Q(n5213) );
  OR2X1 U5588 ( .IN1(n5215), .IN2(n5216), .Q(g11331) );
  AND2X1 U5589 ( .IN1(n1239), .IN2(g481), .Q(n5216) );
  AND2X1 U5590 ( .IN1(n51), .IN2(g486), .Q(n5215) );
  OR2X1 U5591 ( .IN1(n5217), .IN2(n5218), .Q(g11330) );
  AND2X1 U5592 ( .IN1(n1239), .IN2(g525), .Q(n5218) );
  AND2X1 U5593 ( .IN1(n51), .IN2(g521), .Q(n5217) );
  OR2X1 U5594 ( .IN1(n5219), .IN2(n5220), .Q(g11329) );
  AND2X1 U5595 ( .IN1(n1239), .IN2(g530), .Q(n5220) );
  AND2X1 U5596 ( .IN1(n51), .IN2(g525), .Q(n5219) );
  OR2X1 U5597 ( .IN1(n5221), .IN2(n5222), .Q(g11328) );
  AND2X1 U5598 ( .IN1(n1239), .IN2(g534), .Q(n5222) );
  AND2X1 U5599 ( .IN1(n51), .IN2(g530), .Q(n5221) );
  OR2X1 U5600 ( .IN1(n5223), .IN2(n5224), .Q(g11327) );
  AND2X1 U5601 ( .IN1(n1239), .IN2(g538), .Q(n5224) );
  AND2X1 U5602 ( .IN1(n51), .IN2(g534), .Q(n5223) );
  OR2X1 U5603 ( .IN1(n5225), .IN2(n5226), .Q(g11326) );
  AND2X1 U5604 ( .IN1(n1239), .IN2(g542), .Q(n5226) );
  AND2X1 U5605 ( .IN1(n51), .IN2(g538), .Q(n5225) );
  OR2X1 U5606 ( .IN1(n5227), .IN2(n5228), .Q(g11325) );
  AND2X1 U5607 ( .IN1(n1239), .IN2(g476), .Q(n5228) );
  AND2X1 U5608 ( .IN1(n51), .IN2(g542), .Q(n5227) );
  OR2X1 U5609 ( .IN1(n5229), .IN2(n5230), .Q(g11324) );
  AND2X1 U5610 ( .IN1(n4863), .IN2(n1239), .Q(n5230) );
  OR2X1 U5611 ( .IN1(n5231), .IN2(n5232), .Q(n4863) );
  AND2X1 U5612 ( .IN1(n1698), .IN2(n5233), .Q(n5232) );
  OR2X1 U5613 ( .IN1(n5234), .IN2(g525), .Q(n5233) );
  AND2X1 U5614 ( .IN1(n5235), .IN2(n5236), .Q(n5234) );
  AND2X1 U5615 ( .IN1(n5237), .IN2(n5238), .Q(n5236) );
  AND2X1 U5616 ( .IN1(n5239), .IN2(n5240), .Q(n5238) );
  AND2X1 U5617 ( .IN1(n1600), .IN2(n1599), .Q(n5240) );
  AND2X1 U5618 ( .IN1(n1621), .IN2(n1620), .Q(n5239) );
  AND2X1 U5619 ( .IN1(n5241), .IN2(n1689), .Q(n5237) );
  AND2X1 U5620 ( .IN1(n1680), .IN2(n1679), .Q(n5241) );
  AND2X1 U5621 ( .IN1(n5242), .IN2(n5243), .Q(n5235) );
  AND2X1 U5622 ( .IN1(n5244), .IN2(n3283), .Q(n5243) );
  AND2X1 U5623 ( .IN1(n1691), .IN2(n1690), .Q(n5244) );
  AND2X1 U5624 ( .IN1(n5245), .IN2(n3286), .Q(n5242) );
  AND2X1 U5625 ( .IN1(n3285), .IN2(n3284), .Q(n5245) );
  AND2X1 U5626 ( .IN1(n1695), .IN2(g521), .Q(n5231) );
  AND2X1 U5627 ( .IN1(n51), .IN2(g481), .Q(n5229) );
  AND2X1 U5628 ( .IN1(n5246), .IN2(n5148), .Q(g11320) );
  AND2X1 U5629 ( .IN1(n5247), .IN2(n5248), .Q(n5246) );
  OR2X1 U5630 ( .IN1(n5249), .IN2(g369), .Q(n5247) );
  AND2X1 U5631 ( .IN1(n1239), .IN2(n5153), .Q(n5249) );
  OR2X1 U5632 ( .IN1(n5250), .IN2(n5251), .Q(g11314) );
  AND2X1 U5633 ( .IN1(n5252), .IN2(g968), .Q(n5251) );
  AND2X1 U5634 ( .IN1(n1855), .IN2(g861), .Q(n5250) );
  OR2X1 U5635 ( .IN1(n5253), .IN2(n5254), .Q(g11312) );
  AND2X1 U5636 ( .IN1(g965), .IN2(n5252), .Q(n5254) );
  AND2X1 U5637 ( .IN1(n1855), .IN2(g857), .Q(n5253) );
  OR2X1 U5638 ( .IN1(n5255), .IN2(n5256), .Q(g11310) );
  AND2X1 U5639 ( .IN1(g962), .IN2(n5252), .Q(n5256) );
  AND2X1 U5640 ( .IN1(n1855), .IN2(g853), .Q(n5255) );
  OR2X1 U5641 ( .IN1(n5257), .IN2(n5258), .Q(g11308) );
  AND2X1 U5642 ( .IN1(n5252), .IN2(g959), .Q(n5258) );
  AND2X1 U5643 ( .IN1(n1855), .IN2(g849), .Q(n5257) );
  OR2X1 U5644 ( .IN1(n5259), .IN2(n5260), .Q(g11306) );
  AND2X1 U5645 ( .IN1(n5252), .IN2(g956), .Q(n5260) );
  AND2X1 U5646 ( .IN1(n1855), .IN2(g845), .Q(n5259) );
  OR2X1 U5647 ( .IN1(n5261), .IN2(n5262), .Q(g11305) );
  AND2X1 U5648 ( .IN1(n5252), .IN2(g953), .Q(n5262) );
  AND2X1 U5649 ( .IN1(n1855), .IN2(g841), .Q(n5261) );
  OR2X1 U5650 ( .IN1(n5263), .IN2(n5264), .Q(g11303) );
  AND2X1 U5651 ( .IN1(n5252), .IN2(g950), .Q(n5264) );
  AND2X1 U5652 ( .IN1(n1855), .IN2(g837), .Q(n5263) );
  OR2X1 U5653 ( .IN1(n5265), .IN2(n5266), .Q(g11300) );
  AND2X1 U5654 ( .IN1(n5252), .IN2(g947), .Q(n5266) );
  AND2X1 U5655 ( .IN1(n1855), .IN2(g833), .Q(n5265) );
  OR2X1 U5656 ( .IN1(n5267), .IN2(n5268), .Q(g11298) );
  AND2X1 U5657 ( .IN1(n1855), .IN2(g829), .Q(n5268) );
  AND2X1 U5658 ( .IN1(n5252), .IN2(g944), .Q(n5267) );
  INVX0 U5659 ( .INP(n1855), .ZN(n5252) );
  OR2X1 U5660 ( .IN1(n5269), .IN2(n5270), .Q(g11294) );
  OR2X1 U5661 ( .IN1(n5271), .IN2(n5272), .Q(n5270) );
  AND2X1 U5662 ( .IN1(n5273), .IN2(n1682), .Q(n5272) );
  AND2X1 U5663 ( .IN1(n926), .IN2(n5274), .Q(n5273) );
  OR2X1 U5664 ( .IN1(n5275), .IN2(n5276), .Q(n5274) );
  INVX0 U5665 ( .INP(n5277), .ZN(n5276) );
  AND2X1 U5666 ( .IN1(n822), .IN2(n817), .Q(n5277) );
  OR2X1 U5667 ( .IN1(n1605), .IN2(n1608), .Q(n817) );
  OR2X1 U5668 ( .IN1(n3854), .IN2(n5278), .Q(n5275) );
  AND2X1 U5669 ( .IN1(n4587), .IN2(g1857), .Q(n5271) );
  INVX0 U5670 ( .INP(n4447), .ZN(n4587) );
  OR2X1 U5671 ( .IN1(n926), .IN2(n4100), .Q(n4447) );
  AND2X1 U5672 ( .IN1(n5279), .IN2(n4100), .Q(n5269) );
  AND2X1 U5673 ( .IN1(n5280), .IN2(n5281), .Q(n5279) );
  OR2X1 U5674 ( .IN1(n1653), .IN2(n5282), .Q(n5281) );
  OR2X1 U5675 ( .IN1(n5283), .IN2(n5284), .Q(n5282) );
  AND2X1 U5676 ( .IN1(n5285), .IN2(n5286), .Q(n5284) );
  OR2X1 U5677 ( .IN1(n5287), .IN2(n5288), .Q(n5286) );
  OR2X1 U5678 ( .IN1(n5289), .IN2(n5290), .Q(n5285) );
  AND2X1 U5679 ( .IN1(n5291), .IN2(n5292), .Q(n5283) );
  INVX0 U5680 ( .INP(n5293), .ZN(n5292) );
  OR2X1 U5681 ( .IN1(n5294), .IN2(n5295), .Q(n5291) );
  OR2X1 U5682 ( .IN1(g1690), .IN2(n5296), .Q(n5280) );
  OR2X1 U5683 ( .IN1(n5297), .IN2(n5298), .Q(n5296) );
  AND2X1 U5684 ( .IN1(n5299), .IN2(n4413), .Q(n5298) );
  OR2X1 U5685 ( .IN1(n1702), .IN2(n3332), .Q(n4413) );
  OR2X1 U5686 ( .IN1(n1626), .IN2(n3319), .Q(n5299) );
  AND2X1 U5687 ( .IN1(n5300), .IN2(n4722), .Q(n5297) );
  OR2X1 U5688 ( .IN1(n3340), .IN2(n3383), .Q(n4722) );
  OR2X1 U5689 ( .IN1(n1659), .IN2(n1715), .Q(n5300) );
  OR2X1 U5690 ( .IN1(n5301), .IN2(n5302), .Q(g11293) );
  AND2X1 U5691 ( .IN1(n5303), .IN2(n4100), .Q(n5302) );
  OR2X1 U5692 ( .IN1(n5304), .IN2(n5305), .Q(n5303) );
  AND2X1 U5693 ( .IN1(n1653), .IN2(n3320), .Q(n5305) );
  AND2X1 U5694 ( .IN1(n5289), .IN2(g1690), .Q(n5304) );
  AND2X1 U5695 ( .IN1(n5306), .IN2(n3625), .Q(n5301) );
  OR2X1 U5696 ( .IN1(n5307), .IN2(n3854), .Q(n5306) );
  INVX0 U5697 ( .INP(n3637), .ZN(n3854) );
  OR2X1 U5698 ( .IN1(g1814), .IN2(n5308), .Q(n3637) );
  OR2X1 U5699 ( .IN1(n1605), .IN2(g1822), .Q(n5308) );
  AND2X1 U5700 ( .IN1(n5309), .IN2(g1854), .Q(n5307) );
  OR2X1 U5701 ( .IN1(n5310), .IN2(n5311), .Q(n5309) );
  OR2X1 U5702 ( .IN1(n5312), .IN2(n3586), .Q(n5311) );
  OR2X1 U5703 ( .IN1(n3381), .IN2(n1873), .Q(n3586) );
  OR2X1 U5704 ( .IN1(n5313), .IN2(n4100), .Q(n3381) );
  INVX0 U5705 ( .INP(n3625), .ZN(n4100) );
  OR2X1 U5706 ( .IN1(n5314), .IN2(n5315), .Q(n3625) );
  OR2X1 U5707 ( .IN1(g1814), .IN2(g1834), .Q(n5315) );
  OR2X1 U5708 ( .IN1(g1828), .IN2(g1822), .Q(n5314) );
  AND2X1 U5709 ( .IN1(n1608), .IN2(g1834), .Q(n5313) );
  AND2X1 U5710 ( .IN1(n5316), .IN2(n5317), .Q(n5312) );
  AND2X1 U5711 ( .IN1(n822), .IN2(n3645), .Q(n5317) );
  OR2X1 U5712 ( .IN1(n1643), .IN2(g1828), .Q(n822) );
  AND2X1 U5713 ( .IN1(n1380), .IN2(n4137), .Q(n5316) );
  OR2X1 U5714 ( .IN1(n5318), .IN2(n5319), .Q(n4137) );
  OR2X1 U5715 ( .IN1(g1828), .IN2(g1834), .Q(n5319) );
  OR2X1 U5716 ( .IN1(n1608), .IN2(g1840), .Q(n5318) );
  OR2X1 U5717 ( .IN1(n5320), .IN2(n5321), .Q(n5310) );
  AND2X1 U5718 ( .IN1(n1682), .IN2(n5322), .Q(n5321) );
  AND2X1 U5719 ( .IN1(n5323), .IN2(n5324), .Q(n5322) );
  INVX0 U5720 ( .INP(n5325), .ZN(n5324) );
  AND2X1 U5721 ( .IN1(n5326), .IN2(n1380), .Q(n5325) );
  OR2X1 U5722 ( .IN1(n1380), .IN2(n5326), .Q(n5323) );
  AND2X1 U5723 ( .IN1(n5327), .IN2(g1857), .Q(n5320) );
  OR2X1 U5724 ( .IN1(n5328), .IN2(n5329), .Q(n5327) );
  AND2X1 U5725 ( .IN1(n5330), .IN2(n3645), .Q(n5329) );
  AND2X1 U5726 ( .IN1(n5278), .IN2(n5326), .Q(n5328) );
  INVX0 U5727 ( .INP(n3645), .ZN(n5278) );
  OR2X1 U5728 ( .IN1(n1643), .IN2(g1814), .Q(n3645) );
  AND2X1 U5729 ( .IN1(n5148), .IN2(n5331), .Q(g11292) );
  OR2X1 U5730 ( .IN1(n5332), .IN2(g382), .Q(n5331) );
  AND2X1 U5731 ( .IN1(n5148), .IN2(n5333), .Q(g11291) );
  OR2X1 U5732 ( .IN1(n5334), .IN2(n5335), .Q(n5333) );
  INVX0 U5733 ( .INP(n5336), .ZN(n5335) );
  OR2X1 U5734 ( .IN1(n5332), .IN2(n3218), .Q(n5336) );
  AND2X1 U5735 ( .IN1(n1239), .IN2(n5337), .Q(n5332) );
  INVX0 U5736 ( .INP(n5338), .ZN(n5337) );
  OR2X1 U5737 ( .IN1(n1420), .IN2(n1385), .Q(n5338) );
  AND2X1 U5738 ( .IN1(n5339), .IN2(n5340), .Q(n5334) );
  AND2X1 U5739 ( .IN1(n1385), .IN2(g374), .Q(n5339) );
  OR2X1 U5740 ( .IN1(n3218), .IN2(n5341), .Q(n1385) );
  OR2X1 U5741 ( .IN1(n3374), .IN2(n3219), .Q(n5341) );
  AND2X1 U5742 ( .IN1(n5342), .IN2(n5148), .Q(g11290) );
  INVX0 U5743 ( .INP(n5343), .ZN(n5148) );
  OR2X1 U5744 ( .IN1(n650), .IN2(g869), .Q(n5343) );
  AND2X1 U5745 ( .IN1(n5344), .IN2(n5345), .Q(n5342) );
  OR2X1 U5746 ( .IN1(n5340), .IN2(g374), .Q(n5345) );
  INVX0 U5747 ( .INP(n5248), .ZN(n5340) );
  OR2X1 U5748 ( .IN1(n3219), .IN2(n5248), .Q(n5344) );
  OR2X1 U5749 ( .IN1(n51), .IN2(n5346), .Q(n5248) );
  OR2X1 U5750 ( .IN1(n3374), .IN2(n1420), .Q(n5346) );
  OR2X1 U5751 ( .IN1(n5347), .IN2(n5348), .Q(g11270) );
  AND2X1 U5752 ( .IN1(n1239), .IN2(g416), .Q(n5348) );
  AND2X1 U5753 ( .IN1(n51), .IN2(g421), .Q(n5347) );
  OR2X1 U5754 ( .IN1(n5349), .IN2(n5350), .Q(g11269) );
  AND2X1 U5755 ( .IN1(n1239), .IN2(g411), .Q(n5350) );
  AND2X1 U5756 ( .IN1(n51), .IN2(g416), .Q(n5349) );
  OR2X1 U5757 ( .IN1(n5351), .IN2(n5352), .Q(g11268) );
  AND2X1 U5758 ( .IN1(n1239), .IN2(g406), .Q(n5352) );
  AND2X1 U5759 ( .IN1(n51), .IN2(g411), .Q(n5351) );
  OR2X1 U5760 ( .IN1(n5353), .IN2(n5354), .Q(g11267) );
  AND2X1 U5761 ( .IN1(n1239), .IN2(g401), .Q(n5354) );
  AND2X1 U5762 ( .IN1(n51), .IN2(g406), .Q(n5353) );
  OR2X1 U5763 ( .IN1(n5355), .IN2(n5356), .Q(g11266) );
  AND2X1 U5764 ( .IN1(n1239), .IN2(g396), .Q(n5356) );
  AND2X1 U5765 ( .IN1(n51), .IN2(g401), .Q(n5355) );
  OR2X1 U5766 ( .IN1(n5357), .IN2(n5358), .Q(g11265) );
  AND2X1 U5767 ( .IN1(n1239), .IN2(g391), .Q(n5358) );
  AND2X1 U5768 ( .IN1(n51), .IN2(g396), .Q(n5357) );
  OR2X1 U5769 ( .IN1(n5359), .IN2(n5360), .Q(g11264) );
  AND2X1 U5770 ( .IN1(n1239), .IN2(g386), .Q(n5360) );
  AND2X1 U5771 ( .IN1(n51), .IN2(g391), .Q(n5359) );
  OR2X1 U5772 ( .IN1(n5361), .IN2(n5362), .Q(g11263) );
  AND2X1 U5773 ( .IN1(n1239), .IN2(g426), .Q(n5362) );
  AND2X1 U5774 ( .IN1(n51), .IN2(g386), .Q(n5361) );
  OR2X1 U5775 ( .IN1(n5363), .IN2(n5364), .Q(g11262) );
  AND2X1 U5776 ( .IN1(n1239), .IN2(g435), .Q(n5364) );
  AND2X1 U5777 ( .IN1(n51), .IN2(g431), .Q(n5363) );
  OR2X1 U5778 ( .IN1(n5365), .IN2(n5366), .Q(g11261) );
  AND2X1 U5779 ( .IN1(n1239), .IN2(g440), .Q(n5366) );
  AND2X1 U5780 ( .IN1(n51), .IN2(g435), .Q(n5365) );
  OR2X1 U5781 ( .IN1(n5367), .IN2(n5368), .Q(g11260) );
  AND2X1 U5782 ( .IN1(n1239), .IN2(g444), .Q(n5368) );
  AND2X1 U5783 ( .IN1(n51), .IN2(g440), .Q(n5367) );
  OR2X1 U5784 ( .IN1(n5369), .IN2(n5370), .Q(g11259) );
  AND2X1 U5785 ( .IN1(n1239), .IN2(g448), .Q(n5370) );
  AND2X1 U5786 ( .IN1(n51), .IN2(g444), .Q(n5369) );
  OR2X1 U5787 ( .IN1(n5371), .IN2(n5372), .Q(g11258) );
  AND2X1 U5788 ( .IN1(n1239), .IN2(g452), .Q(n5372) );
  AND2X1 U5789 ( .IN1(n51), .IN2(g448), .Q(n5371) );
  OR2X1 U5790 ( .IN1(n5373), .IN2(n5374), .Q(g11257) );
  AND2X1 U5791 ( .IN1(n1239), .IN2(g421), .Q(n5374) );
  AND2X1 U5792 ( .IN1(n51), .IN2(g452), .Q(n5373) );
  OR2X1 U5793 ( .IN1(n5375), .IN2(n5376), .Q(g11256) );
  AND2X1 U5794 ( .IN1(n5177), .IN2(n1239), .Q(n5376) );
  INVX0 U5795 ( .INP(n5176), .ZN(n5177) );
  OR2X1 U5796 ( .IN1(n5377), .IN2(n5378), .Q(n5176) );
  AND2X1 U5797 ( .IN1(n5379), .IN2(n1420), .Q(n5378) );
  OR2X1 U5798 ( .IN1(n5380), .IN2(n5381), .Q(n5379) );
  AND2X1 U5799 ( .IN1(n5382), .IN2(n1878), .Q(n5381) );
  AND2X1 U5800 ( .IN1(n1876), .IN2(n5383), .Q(n5382) );
  OR2X1 U5801 ( .IN1(n5384), .IN2(n5385), .Q(n5383) );
  OR2X1 U5802 ( .IN1(n5386), .IN2(n5387), .Q(n5385) );
  OR2X1 U5803 ( .IN1(g391), .IN2(n5388), .Q(n5387) );
  OR2X1 U5804 ( .IN1(g386), .IN2(g426), .Q(n5388) );
  OR2X1 U5805 ( .IN1(g396), .IN2(n5389), .Q(n5386) );
  OR2X1 U5806 ( .IN1(g448), .IN2(g452), .Q(n5389) );
  OR2X1 U5807 ( .IN1(n5390), .IN2(n5391), .Q(n5384) );
  OR2X1 U5808 ( .IN1(g444), .IN2(n5392), .Q(n5391) );
  OR2X1 U5809 ( .IN1(g406), .IN2(g440), .Q(n5392) );
  OR2X1 U5810 ( .IN1(n5393), .IN2(n5394), .Q(n5390) );
  OR2X1 U5811 ( .IN1(g421), .IN2(g416), .Q(n5394) );
  OR2X1 U5812 ( .IN1(g411), .IN2(g401), .Q(n5393) );
  AND2X1 U5813 ( .IN1(g431), .IN2(g435), .Q(n5380) );
  AND2X1 U5814 ( .IN1(n1681), .IN2(n5153), .Q(n5377) );
  INVX0 U5815 ( .INP(n1420), .ZN(n5153) );
  AND2X1 U5816 ( .IN1(n51), .IN2(g426), .Q(n5375) );
  INVX0 U5817 ( .INP(n1239), .ZN(n51) );
  OR2X1 U5818 ( .IN1(n5395), .IN2(n5396), .Q(n1239) );
  OR2X1 U5819 ( .IN1(n5397), .IN2(n5398), .Q(n5396) );
  OR2X1 U5820 ( .IN1(g849), .IN2(g845), .Q(n5398) );
  OR2X1 U5821 ( .IN1(g853), .IN2(n5399), .Q(n5397) );
  OR2X1 U5822 ( .IN1(g841), .IN2(g857), .Q(n5399) );
  OR2X1 U5823 ( .IN1(n5400), .IN2(n5401), .Q(n5395) );
  OR2X1 U5824 ( .IN1(g837), .IN2(g861), .Q(n5401) );
  OR2X1 U5825 ( .IN1(g833), .IN2(n5402), .Q(n5400) );
  OR2X1 U5826 ( .IN1(n5403), .IN2(g829), .Q(n5402) );
  AND2X1 U5827 ( .IN1(n5404), .IN2(n5405), .Q(n5403) );
  OR2X1 U5828 ( .IN1(n650), .IN2(n5406), .Q(n5405) );
  AND2X1 U5829 ( .IN1(n5407), .IN2(n5408), .Q(n5406) );
  INVX0 U5830 ( .INP(n5409), .ZN(n5404) );
  OR2X1 U5831 ( .IN1(n5410), .IN2(n5411), .Q(n5409) );
  AND2X1 U5832 ( .IN1(g10628), .IN2(n5412), .Q(g11206) );
  AND2X1 U5833 ( .IN1(n5413), .IN2(n5414), .Q(g11163) );
  INVX0 U5834 ( .INP(n5415), .ZN(n5414) );
  AND2X1 U5835 ( .IN1(n5412), .IN2(n3375), .Q(n5415) );
  OR2X1 U5836 ( .IN1(n5412), .IN2(n3375), .Q(n5413) );
  INVX0 U5837 ( .INP(n5416), .ZN(n5412) );
  OR2X1 U5838 ( .IN1(n5417), .IN2(n5418), .Q(n5416) );
  OR2X1 U5839 ( .IN1(n5419), .IN2(n5420), .Q(n5418) );
  AND2X1 U5840 ( .IN1(n4804), .IN2(g10724), .Q(n5420) );
  INVX0 U5841 ( .INP(n4675), .ZN(n4804) );
  OR2X1 U5842 ( .IN1(n3050), .IN2(n5421), .Q(n4675) );
  OR2X1 U5843 ( .IN1(n3108), .IN2(n650), .Q(n5421) );
  AND2X1 U5844 ( .IN1(n5422), .IN2(g109), .Q(n5419) );
  OR2X1 U5845 ( .IN1(n5423), .IN2(n5424), .Q(n5422) );
  OR2X1 U5846 ( .IN1(n5425), .IN2(n5426), .Q(n5424) );
  AND2X1 U5847 ( .IN1(g10664), .IN2(g2648), .Q(n5426) );
  AND2X1 U5848 ( .IN1(n5410), .IN2(n3036), .Q(n5425) );
  AND2X1 U5849 ( .IN1(n3373), .IN2(g10726), .Q(n5423) );
  AND2X1 U5850 ( .IN1(g5392), .IN2(g10663), .Q(n5417) );
  AND2X1 U5851 ( .IN1(g109), .IN2(n4758), .Q(g5392) );
  INVX0 U5852 ( .INP(n4757), .ZN(n4758) );
  OR2X1 U5853 ( .IN1(n3365), .IN2(n3366), .Q(n4757) );
  OR2X1 U5854 ( .IN1(n5427), .IN2(n5428), .Q(g10936) );
  AND2X1 U5855 ( .IN1(n1391), .IN2(n3382), .Q(n5428) );
  OR2X1 U5856 ( .IN1(n5429), .IN2(n5430), .Q(n1391) );
  INVX0 U5857 ( .INP(n5431), .ZN(n5430) );
  AND2X1 U5858 ( .IN1(n5408), .IN2(n5410), .Q(n5431) );
  OR2X1 U5859 ( .IN1(g10721), .IN2(n4989), .Q(n5429) );
  AND2X1 U5860 ( .IN1(n493), .IN2(g1811), .Q(n5427) );
  OR2X1 U5861 ( .IN1(n5432), .IN2(n5433), .Q(g10898) );
  AND2X1 U5862 ( .IN1(n5434), .IN2(n3946), .Q(n5433) );
  OR2X1 U5863 ( .IN1(n4782), .IN2(n5435), .Q(n5434) );
  OR2X1 U5864 ( .IN1(n5436), .IN2(n5437), .Q(n5435) );
  AND2X1 U5865 ( .IN1(n5438), .IN2(n5439), .Q(n5437) );
  INVX0 U5866 ( .INP(n5440), .ZN(n5436) );
  OR2X1 U5867 ( .IN1(n5439), .IN2(n5438), .Q(n5440) );
  OR2X1 U5868 ( .IN1(n5441), .IN2(n5442), .Q(n5438) );
  AND2X1 U5869 ( .IN1(n3221), .IN2(n3386), .Q(n5442) );
  AND2X1 U5870 ( .IN1(test_so8), .IN2(g1019), .Q(n5441) );
  INVX0 U5871 ( .INP(n5443), .ZN(n5439) );
  OR2X1 U5872 ( .IN1(n5444), .IN2(n5445), .Q(n5443) );
  AND2X1 U5873 ( .IN1(n5446), .IN2(n3291), .Q(n5445) );
  AND2X1 U5874 ( .IN1(n5447), .IN2(n5448), .Q(n5446) );
  OR2X1 U5875 ( .IN1(n5449), .IN2(n5450), .Q(n5448) );
  OR2X1 U5876 ( .IN1(n5451), .IN2(n5452), .Q(n5447) );
  AND2X1 U5877 ( .IN1(n5453), .IN2(g995), .Q(n5444) );
  OR2X1 U5878 ( .IN1(n5454), .IN2(n5455), .Q(n5453) );
  AND2X1 U5879 ( .IN1(n5449), .IN2(n5450), .Q(n5455) );
  INVX0 U5880 ( .INP(n5452), .ZN(n5449) );
  AND2X1 U5881 ( .IN1(n5451), .IN2(n5452), .Q(n5454) );
  AND2X1 U5882 ( .IN1(n5456), .IN2(n5457), .Q(n5452) );
  OR2X1 U5883 ( .IN1(n5458), .IN2(n5459), .Q(n5457) );
  INVX0 U5884 ( .INP(n5460), .ZN(n5458) );
  OR2X1 U5885 ( .IN1(n5461), .IN2(n5460), .Q(n5456) );
  OR2X1 U5886 ( .IN1(n5462), .IN2(n5463), .Q(n5460) );
  AND2X1 U5887 ( .IN1(n3200), .IN2(g1015), .Q(n5463) );
  AND2X1 U5888 ( .IN1(n3220), .IN2(g1023), .Q(n5462) );
  INVX0 U5889 ( .INP(n5459), .ZN(n5461) );
  OR2X1 U5890 ( .IN1(n5464), .IN2(n5465), .Q(n5459) );
  AND2X1 U5891 ( .IN1(n3255), .IN2(n3385), .Q(n5465) );
  AND2X1 U5892 ( .IN1(test_so2), .IN2(g1011), .Q(n5464) );
  INVX0 U5893 ( .INP(n5450), .ZN(n5451) );
  AND2X1 U5894 ( .IN1(n5466), .IN2(n5467), .Q(n5450) );
  OR2X1 U5895 ( .IN1(n5468), .IN2(n1871), .Q(n5467) );
  INVX0 U5896 ( .INP(n5469), .ZN(n5468) );
  OR2X1 U5897 ( .IN1(n5469), .IN2(g991), .Q(n5466) );
  OR2X1 U5898 ( .IN1(n5470), .IN2(n5471), .Q(n5469) );
  AND2X1 U5899 ( .IN1(n3293), .IN2(g1027), .Q(n5471) );
  AND2X1 U5900 ( .IN1(n3324), .IN2(g1003), .Q(n5470) );
  INVX0 U5901 ( .INP(n4785), .ZN(n4782) );
  OR2X1 U5902 ( .IN1(g10663), .IN2(n4989), .Q(n4785) );
  INVX0 U5903 ( .INP(n5472), .ZN(n4989) );
  OR2X1 U5904 ( .IN1(n3593), .IN2(n5473), .Q(n5472) );
  OR2X1 U5905 ( .IN1(g46), .IN2(n5474), .Q(n5473) );
  OR2X1 U5906 ( .IN1(n5475), .IN2(n3590), .Q(n3593) );
  OR2X1 U5907 ( .IN1(n5476), .IN2(n5477), .Q(n3590) );
  OR2X1 U5908 ( .IN1(g48), .IN2(g45), .Q(n5476) );
  AND2X1 U5909 ( .IN1(n495), .IN2(g105), .Q(n5432) );
  OR2X1 U5910 ( .IN1(n5478), .IN2(n5479), .Q(g10866) );
  AND2X1 U5911 ( .IN1(n495), .IN2(g1684), .Q(n5478) );
  OR2X1 U5912 ( .IN1(n5480), .IN2(n5481), .Q(g10865) );
  AND2X1 U5913 ( .IN1(n5482), .IN2(n4628), .Q(n5481) );
  AND2X1 U5914 ( .IN1(n1404), .IN2(n5483), .Q(n5482) );
  OR2X1 U5915 ( .IN1(n650), .IN2(g10722), .Q(n5483) );
  AND2X1 U5916 ( .IN1(n4627), .IN2(g1669), .Q(n5480) );
  OR2X1 U5917 ( .IN1(n5484), .IN2(n5485), .Q(g10864) );
  AND2X1 U5918 ( .IN1(n495), .IN2(g1681), .Q(n5484) );
  OR2X1 U5919 ( .IN1(n5486), .IN2(n5487), .Q(g10863) );
  AND2X1 U5920 ( .IN1(n5488), .IN2(n4628), .Q(n5487) );
  AND2X1 U5921 ( .IN1(n5489), .IN2(n5490), .Q(n5488) );
  OR2X1 U5922 ( .IN1(n5411), .IN2(g1718), .Q(n5489) );
  AND2X1 U5923 ( .IN1(n4627), .IN2(g1666), .Q(n5486) );
  OR2X1 U5924 ( .IN1(n5491), .IN2(n5492), .Q(g10862) );
  AND2X1 U5925 ( .IN1(n495), .IN2(g1678), .Q(n5491) );
  OR2X1 U5926 ( .IN1(n5493), .IN2(n5494), .Q(g10861) );
  AND2X1 U5927 ( .IN1(n5495), .IN2(n4628), .Q(n5494) );
  AND2X1 U5928 ( .IN1(n4627), .IN2(g1663), .Q(n5493) );
  OR2X1 U5929 ( .IN1(n5496), .IN2(n5497), .Q(g10860) );
  AND2X1 U5930 ( .IN1(n495), .IN2(g1675), .Q(n5496) );
  OR2X1 U5931 ( .IN1(n5498), .IN2(n5499), .Q(g10859) );
  AND2X1 U5932 ( .IN1(n5500), .IN2(n4628), .Q(n5499) );
  AND2X1 U5933 ( .IN1(n4627), .IN2(g1660), .Q(n5498) );
  OR2X1 U5934 ( .IN1(n5501), .IN2(n5502), .Q(g10858) );
  AND2X1 U5935 ( .IN1(n495), .IN2(g1672), .Q(n5501) );
  OR2X1 U5936 ( .IN1(n5503), .IN2(n5504), .Q(g10855) );
  AND2X1 U5937 ( .IN1(n5495), .IN2(n3946), .Q(n5504) );
  OR2X1 U5938 ( .IN1(n5505), .IN2(n5506), .Q(n5495) );
  AND2X1 U5939 ( .IN1(n4264), .IN2(n5507), .Q(n5506) );
  OR2X1 U5940 ( .IN1(n4645), .IN2(n5508), .Q(n4264) );
  AND2X1 U5941 ( .IN1(n3963), .IN2(g1512), .Q(n5508) );
  AND2X1 U5942 ( .IN1(g18), .IN2(g192), .Q(n4645) );
  AND2X1 U5943 ( .IN1(n5509), .IN2(n5490), .Q(n5505) );
  OR2X1 U5944 ( .IN1(n5510), .IN2(g1718), .Q(n5509) );
  AND2X1 U5945 ( .IN1(n495), .IN2(g549), .Q(n5503) );
  OR2X1 U5946 ( .IN1(n3375), .IN2(n3580), .Q(g10801) );
  AND2X1 U5947 ( .IN1(n5511), .IN2(n5512), .Q(n3375) );
  INVX0 U5948 ( .INP(n5513), .ZN(n5512) );
  AND2X1 U5949 ( .IN1(n5514), .IN2(n5515), .Q(n5513) );
  OR2X1 U5950 ( .IN1(n5515), .IN2(n5514), .Q(n5511) );
  OR2X1 U5951 ( .IN1(n5516), .IN2(n5517), .Q(n5514) );
  AND2X1 U5952 ( .IN1(n5518), .IN2(n5519), .Q(n5517) );
  AND2X1 U5953 ( .IN1(n5520), .IN2(n5521), .Q(n5519) );
  OR2X1 U5954 ( .IN1(n5522), .IN2(n5523), .Q(n5521) );
  OR2X1 U5955 ( .IN1(n5524), .IN2(n5525), .Q(n5520) );
  AND2X1 U5956 ( .IN1(n5526), .IN2(n72), .Q(n5516) );
  INVX0 U5957 ( .INP(n5518), .ZN(n72) );
  OR2X1 U5958 ( .IN1(n5527), .IN2(n5528), .Q(n5518) );
  AND2X1 U5959 ( .IN1(g10722), .IN2(n5287), .Q(n5528) );
  INVX0 U5960 ( .INP(g10721), .ZN(n5287) );
  AND2X1 U5961 ( .IN1(g10721), .IN2(n5288), .Q(n5527) );
  INVX0 U5962 ( .INP(g10722), .ZN(n5288) );
  OR2X1 U5963 ( .IN1(n5529), .IN2(n5530), .Q(n5526) );
  AND2X1 U5964 ( .IN1(n5522), .IN2(n5523), .Q(n5530) );
  AND2X1 U5965 ( .IN1(n5524), .IN2(n5525), .Q(n5529) );
  INVX0 U5966 ( .INP(n5522), .ZN(n5525) );
  AND2X1 U5967 ( .IN1(n5531), .IN2(n3389), .Q(n5522) );
  INVX0 U5968 ( .INP(n5523), .ZN(n5524) );
  OR2X1 U5969 ( .IN1(n5407), .IN2(n5532), .Q(n5523) );
  OR2X1 U5970 ( .IN1(n5533), .IN2(n5534), .Q(n5532) );
  AND2X1 U5971 ( .IN1(n5293), .IN2(n5295), .Q(n5534) );
  AND2X1 U5972 ( .IN1(g10663), .IN2(g10664), .Q(n5293) );
  AND2X1 U5973 ( .IN1(n5535), .IN2(g10726), .Q(n5533) );
  OR2X1 U5974 ( .IN1(n5536), .IN2(n5537), .Q(n5535) );
  AND2X1 U5975 ( .IN1(g10663), .IN2(n5538), .Q(n5537) );
  AND2X1 U5976 ( .IN1(g10664), .IN2(n5539), .Q(n5536) );
  AND2X1 U5977 ( .IN1(n5539), .IN2(n5540), .Q(n5407) );
  AND2X1 U5978 ( .IN1(n5295), .IN2(n5538), .Q(n5540) );
  INVX0 U5979 ( .INP(g10664), .ZN(n5538) );
  INVX0 U5980 ( .INP(g10663), .ZN(n5539) );
  OR2X1 U5981 ( .IN1(n5408), .IN2(n5541), .Q(n5515) );
  OR2X1 U5982 ( .IN1(n5542), .IN2(n5543), .Q(n5541) );
  AND2X1 U5983 ( .IN1(n5544), .IN2(n5294), .Q(n5543) );
  AND2X1 U5984 ( .IN1(g10719), .IN2(g10720), .Q(n5544) );
  AND2X1 U5985 ( .IN1(n5545), .IN2(g10724), .Q(n5542) );
  OR2X1 U5986 ( .IN1(n5546), .IN2(n5547), .Q(n5545) );
  AND2X1 U5987 ( .IN1(g10720), .IN2(n5289), .Q(n5547) );
  AND2X1 U5988 ( .IN1(g10719), .IN2(n5290), .Q(n5546) );
  AND2X1 U5989 ( .IN1(n5289), .IN2(n5548), .Q(n5408) );
  AND2X1 U5990 ( .IN1(n5294), .IN2(n5290), .Q(n5548) );
  INVX0 U5991 ( .INP(g10720), .ZN(n5290) );
  OR2X1 U5992 ( .IN1(n5549), .IN2(n5550), .Q(g10800) );
  AND2X1 U5993 ( .IN1(n5500), .IN2(n3946), .Q(n5550) );
  OR2X1 U5994 ( .IN1(n5551), .IN2(n5552), .Q(n5500) );
  AND2X1 U5995 ( .IN1(n4250), .IN2(n5507), .Q(n5552) );
  OR2X1 U5996 ( .IN1(n4647), .IN2(n5553), .Q(n4250) );
  AND2X1 U5997 ( .IN1(n3963), .IN2(g1636), .Q(n5553) );
  AND2X1 U5998 ( .IN1(g18), .IN2(g248), .Q(n4647) );
  AND2X1 U5999 ( .IN1(n5554), .IN2(n5490), .Q(n5551) );
  OR2X1 U6000 ( .IN1(g10719), .IN2(n5555), .Q(n5554) );
  AND2X1 U6001 ( .IN1(n495), .IN2(g575), .Q(n5549) );
  OR2X1 U6002 ( .IN1(n5556), .IN2(n5557), .Q(g10799) );
  AND2X1 U6003 ( .IN1(n495), .IN2(g566), .Q(n5556) );
  OR2X1 U6004 ( .IN1(n5558), .IN2(n5479), .Q(g10798) );
  AND2X1 U6005 ( .IN1(n5559), .IN2(n3946), .Q(n5479) );
  OR2X1 U6006 ( .IN1(n5560), .IN2(n5561), .Q(n5559) );
  AND2X1 U6007 ( .IN1(n1404), .IN2(n5326), .Q(n5561) );
  AND2X1 U6008 ( .IN1(n5507), .IN2(n4260), .Q(n5560) );
  OR2X1 U6009 ( .IN1(n5562), .IN2(n3978), .Q(n4260) );
  INVX0 U6010 ( .INP(n5563), .ZN(n3978) );
  OR2X1 U6011 ( .IN1(n3357), .IN2(n3963), .Q(n5563) );
  AND2X1 U6012 ( .IN1(n3963), .IN2(g1624), .Q(n5562) );
  AND2X1 U6013 ( .IN1(n495), .IN2(g563), .Q(n5558) );
  OR2X1 U6014 ( .IN1(n5564), .IN2(n5485), .Q(g10797) );
  AND2X1 U6015 ( .IN1(n5565), .IN2(n3946), .Q(n5485) );
  OR2X1 U6016 ( .IN1(n5566), .IN2(n5567), .Q(n5565) );
  AND2X1 U6017 ( .IN1(n1404), .IN2(n5410), .Q(n5567) );
  AND2X1 U6018 ( .IN1(n5507), .IN2(n4246), .Q(n5566) );
  OR2X1 U6019 ( .IN1(n5568), .IN2(n3961), .Q(n4246) );
  INVX0 U6020 ( .INP(n5569), .ZN(n3961) );
  OR2X1 U6021 ( .IN1(n3360), .IN2(n3963), .Q(n5569) );
  AND2X1 U6022 ( .IN1(n3963), .IN2(g1621), .Q(n5568) );
  AND2X1 U6023 ( .IN1(n495), .IN2(g560), .Q(n5564) );
  OR2X1 U6024 ( .IN1(n5570), .IN2(n5492), .Q(g10795) );
  AND2X1 U6025 ( .IN1(n5571), .IN2(n3946), .Q(n5492) );
  OR2X1 U6026 ( .IN1(n5572), .IN2(n5573), .Q(n5571) );
  AND2X1 U6027 ( .IN1(n1404), .IN2(n5411), .Q(n5573) );
  AND2X1 U6028 ( .IN1(n5507), .IN2(n4220), .Q(n5572) );
  OR2X1 U6029 ( .IN1(n5574), .IN2(n4045), .Q(n4220) );
  AND2X1 U6030 ( .IN1(g213), .IN2(g18), .Q(n4045) );
  AND2X1 U6031 ( .IN1(n3963), .IN2(g1615), .Q(n5574) );
  AND2X1 U6032 ( .IN1(n495), .IN2(g557), .Q(n5570) );
  OR2X1 U6033 ( .IN1(n5575), .IN2(n5497), .Q(g10793) );
  AND2X1 U6034 ( .IN1(n3946), .IN2(n5576), .Q(n5497) );
  AND2X1 U6035 ( .IN1(n5577), .IN2(n5578), .Q(n5576) );
  OR2X1 U6036 ( .IN1(n4207), .IN2(n5490), .Q(n5578) );
  OR2X1 U6037 ( .IN1(n5579), .IN2(n4021), .Q(n4207) );
  INVX0 U6038 ( .INP(n5580), .ZN(n4021) );
  OR2X1 U6039 ( .IN1(n3358), .IN2(n3963), .Q(n5580) );
  AND2X1 U6040 ( .IN1(n3963), .IN2(g1639), .Q(n5579) );
  OR2X1 U6041 ( .IN1(n5581), .IN2(n5507), .Q(n5577) );
  OR2X1 U6042 ( .IN1(n5555), .IN2(g10720), .Q(n5581) );
  OR2X1 U6043 ( .IN1(n650), .IN2(g1718), .Q(n5555) );
  AND2X1 U6044 ( .IN1(n495), .IN2(g554), .Q(n5575) );
  OR2X1 U6045 ( .IN1(n5582), .IN2(n5502), .Q(g10791) );
  INVX0 U6046 ( .INP(n5583), .ZN(n5502) );
  OR2X1 U6047 ( .IN1(n495), .IN2(n5584), .Q(n5583) );
  AND2X1 U6048 ( .IN1(n5585), .IN2(n5586), .Q(n5584) );
  OR2X1 U6049 ( .IN1(n5587), .IN2(n5588), .Q(n5586) );
  OR2X1 U6050 ( .IN1(n650), .IN2(n5289), .Q(n5588) );
  INVX0 U6051 ( .INP(g10719), .ZN(n5289) );
  OR2X1 U6052 ( .IN1(n4269), .IN2(n5490), .Q(n5585) );
  INVX0 U6053 ( .INP(n4270), .ZN(n4269) );
  OR2X1 U6054 ( .IN1(n5589), .IN2(n3996), .Q(n4270) );
  AND2X1 U6055 ( .IN1(g186), .IN2(g18), .Q(n3996) );
  AND2X1 U6056 ( .IN1(n3963), .IN2(g1618), .Q(n5589) );
  AND2X1 U6057 ( .IN1(n495), .IN2(g546), .Q(n5582) );
  AND2X1 U6058 ( .IN1(n493), .IN2(n3023), .Q(g10785) );
  AND2X1 U6059 ( .IN1(n493), .IN2(n3029), .Q(g10784) );
  AND2X1 U6060 ( .IN1(n493), .IN2(n3065), .Q(g10782) );
  AND2X1 U6061 ( .IN1(n493), .IN2(n3017), .Q(g10780) );
  INVX0 U6062 ( .INP(n3382), .ZN(n493) );
  AND2X1 U6063 ( .IN1(n3331), .IN2(g1696), .Q(n3382) );
  OR2X1 U6064 ( .IN1(n5590), .IN2(n5557), .Q(g10776) );
  INVX0 U6065 ( .INP(n5591), .ZN(n5557) );
  OR2X1 U6066 ( .IN1(n495), .IN2(n5592), .Q(n5591) );
  AND2X1 U6067 ( .IN1(n5593), .IN2(n5594), .Q(n5592) );
  OR2X1 U6068 ( .IN1(n5295), .IN2(n5587), .Q(n5594) );
  INVX0 U6069 ( .INP(g10726), .ZN(n5295) );
  AND2X1 U6070 ( .IN1(n5595), .IN2(n5596), .Q(n5593) );
  INVX0 U6071 ( .INP(n1450), .ZN(n5596) );
  OR2X1 U6072 ( .IN1(n4274), .IN2(n5490), .Q(n5595) );
  INVX0 U6073 ( .INP(n4275), .ZN(n4274) );
  OR2X1 U6074 ( .IN1(n5597), .IN2(n4008), .Q(n4275) );
  INVX0 U6075 ( .INP(n5598), .ZN(n4008) );
  OR2X1 U6076 ( .IN1(n3359), .IN2(n3963), .Q(n5598) );
  AND2X1 U6077 ( .IN1(n3963), .IN2(g1627), .Q(n5597) );
  AND2X1 U6078 ( .IN1(n495), .IN2(g1687), .Q(n5590) );
  OR2X1 U6079 ( .IN1(n5599), .IN2(n5600), .Q(g10773) );
  AND2X1 U6080 ( .IN1(n4742), .IN2(g1727), .Q(n5600) );
  AND2X1 U6081 ( .IN1(n5601), .IN2(n5411), .Q(n5599) );
  OR2X1 U6082 ( .IN1(n5602), .IN2(n5603), .Q(g10771) );
  AND2X1 U6083 ( .IN1(n5510), .IN2(n5601), .Q(n5603) );
  AND2X1 U6084 ( .IN1(g109), .IN2(g10720), .Q(n5510) );
  AND2X1 U6085 ( .IN1(n4742), .IN2(g1724), .Q(n5602) );
  OR2X1 U6086 ( .IN1(n5604), .IN2(n5605), .Q(g10770) );
  AND2X1 U6087 ( .IN1(n5606), .IN2(n5601), .Q(n5605) );
  AND2X1 U6088 ( .IN1(g109), .IN2(g10719), .Q(n5606) );
  AND2X1 U6089 ( .IN1(n4742), .IN2(g1721), .Q(n5604) );
  OR2X1 U6090 ( .IN1(n5607), .IN2(n5608), .Q(g10767) );
  AND2X1 U6091 ( .IN1(n5609), .IN2(n4628), .Q(n5608) );
  AND2X1 U6092 ( .IN1(n4627), .IN2(g1657), .Q(n5607) );
  OR2X1 U6093 ( .IN1(n5610), .IN2(n5611), .Q(g10765) );
  AND2X1 U6094 ( .IN1(n4628), .IN2(n5612), .Q(n5611) );
  INVX0 U6095 ( .INP(n4627), .ZN(n4628) );
  AND2X1 U6096 ( .IN1(n4627), .IN2(g1654), .Q(n5610) );
  OR2X1 U6097 ( .IN1(g1696), .IN2(n3331), .Q(n4627) );
  OR2X1 U6098 ( .IN1(n5613), .IN2(n5614), .Q(g10718) );
  AND2X1 U6099 ( .IN1(n5609), .IN2(n3946), .Q(n5614) );
  OR2X1 U6100 ( .IN1(n5615), .IN2(n5616), .Q(n5609) );
  AND2X1 U6101 ( .IN1(n4224), .IN2(n5507), .Q(n5616) );
  OR2X1 U6102 ( .IN1(n4649), .IN2(n5617), .Q(n4224) );
  AND2X1 U6103 ( .IN1(n3963), .IN2(g1633), .Q(n5617) );
  AND2X1 U6104 ( .IN1(g18), .IN2(g243), .Q(n4649) );
  AND2X1 U6105 ( .IN1(n5618), .IN2(n5490), .Q(n5615) );
  INVX0 U6106 ( .INP(n5507), .ZN(n5490) );
  OR2X1 U6107 ( .IN1(n5619), .IN2(g1718), .Q(n5618) );
  AND2X1 U6108 ( .IN1(g10664), .IN2(g109), .Q(n5619) );
  AND2X1 U6109 ( .IN1(n495), .IN2(g572), .Q(n5613) );
  OR2X1 U6110 ( .IN1(n5620), .IN2(n5621), .Q(g10717) );
  AND2X1 U6111 ( .IN1(n5612), .IN2(n3946), .Q(n5621) );
  OR2X1 U6112 ( .IN1(n5622), .IN2(n5623), .Q(n5612) );
  OR2X1 U6113 ( .IN1(n1450), .IN2(n5624), .Q(n5623) );
  AND2X1 U6114 ( .IN1(n5507), .IN2(n4280), .Q(n5624) );
  OR2X1 U6115 ( .IN1(n5625), .IN2(n4033), .Q(n4280) );
  AND2X1 U6116 ( .IN1(g237), .IN2(g18), .Q(n4033) );
  AND2X1 U6117 ( .IN1(n3963), .IN2(g1630), .Q(n5625) );
  INVX0 U6118 ( .INP(g18), .ZN(n3963) );
  AND2X1 U6119 ( .IN1(n1404), .IN2(g10663), .Q(n5622) );
  INVX0 U6120 ( .INP(n5587), .ZN(n1404) );
  OR2X1 U6121 ( .IN1(n5507), .IN2(g1718), .Q(n5587) );
  AND2X1 U6122 ( .IN1(n1611), .IN2(n6004), .Q(n5507) );
  AND2X1 U6123 ( .IN1(n495), .IN2(g569), .Q(n5620) );
  INVX0 U6124 ( .INP(n3946), .ZN(n495) );
  AND2X1 U6125 ( .IN1(n4471), .IN2(n3331), .Q(n3946) );
  OR2X1 U6126 ( .IN1(n5626), .IN2(n5627), .Q(g10711) );
  AND2X1 U6127 ( .IN1(n5601), .IN2(n5326), .Q(n5627) );
  INVX0 U6128 ( .INP(n5330), .ZN(n5326) );
  AND2X1 U6129 ( .IN1(g109), .IN2(n5294), .Q(n5330) );
  INVX0 U6130 ( .INP(g10724), .ZN(n5294) );
  AND2X1 U6131 ( .IN1(n4742), .IN2(g1733), .Q(n5626) );
  OR2X1 U6132 ( .IN1(n5628), .IN2(n5629), .Q(g10707) );
  AND2X1 U6133 ( .IN1(n4742), .IN2(g1730), .Q(n5629) );
  AND2X1 U6134 ( .IN1(n5601), .IN2(n5410), .Q(n5628) );
  INVX0 U6135 ( .INP(n4742), .ZN(n5601) );
  OR2X1 U6136 ( .IN1(n3331), .IN2(n4471), .Q(n4742) );
  INVX0 U6137 ( .INP(g1696), .ZN(n4471) );
  OR2X1 U6138 ( .IN1(n5630), .IN2(n5631), .Q(g10664) );
  OR2X1 U6139 ( .IN1(n5632), .IN2(n5633), .Q(n5631) );
  OR2X1 U6140 ( .IN1(n5634), .IN2(n5635), .Q(n5633) );
  OR2X1 U6141 ( .IN1(n5636), .IN2(n5637), .Q(n5635) );
  AND2X1 U6142 ( .IN1(g1191), .IN2(n5638), .Q(n5637) );
  AND2X1 U6143 ( .IN1(n5639), .IN2(n5640), .Q(n5636) );
  AND2X1 U6144 ( .IN1(n5641), .IN2(n5642), .Q(n5639) );
  INVX0 U6145 ( .INP(n5643), .ZN(n5642) );
  OR2X1 U6146 ( .IN1(n5644), .IN2(n5645), .Q(n5643) );
  OR2X1 U6147 ( .IN1(n1480), .IN2(n1479), .Q(n5644) );
  AND2X1 U6148 ( .IN1(n5646), .IN2(n1478), .Q(n5641) );
  AND2X1 U6149 ( .IN1(n5647), .IN2(n5648), .Q(n5646) );
  OR2X1 U6150 ( .IN1(n5649), .IN2(n5650), .Q(n5647) );
  AND2X1 U6151 ( .IN1(n5651), .IN2(n5652), .Q(n5649) );
  AND2X1 U6152 ( .IN1(test_so9), .IN2(n5653), .Q(n5634) );
  OR2X1 U6153 ( .IN1(n5654), .IN2(n5655), .Q(n5632) );
  AND2X1 U6154 ( .IN1(n5645), .IN2(g1741), .Q(n5655) );
  AND2X1 U6155 ( .IN1(n1486), .IN2(g1546), .Q(n5654) );
  OR2X1 U6156 ( .IN1(n5656), .IN2(n5657), .Q(n5630) );
  OR2X1 U6157 ( .IN1(n5658), .IN2(n5659), .Q(n5657) );
  AND2X1 U6158 ( .IN1(n1485), .IN2(g1589), .Q(n5659) );
  AND2X1 U6159 ( .IN1(n5531), .IN2(n3040), .Q(n5658) );
  OR2X1 U6160 ( .IN1(n5660), .IN2(n5661), .Q(n5656) );
  OR2X1 U6161 ( .IN1(n5662), .IN2(n5663), .Q(n5661) );
  AND2X1 U6162 ( .IN1(g919), .IN2(n5664), .Q(n5663) );
  AND2X1 U6163 ( .IN1(n5665), .IN2(g284), .Q(n5662) );
  AND2X1 U6164 ( .IN1(n5666), .IN2(g947), .Q(n5660) );
  INVX0 U6165 ( .INP(n5667), .ZN(g10628) );
  OR2X1 U6166 ( .IN1(n5668), .IN2(n5669), .Q(n5667) );
  AND2X1 U6167 ( .IN1(n5411), .IN2(n4194), .Q(n5669) );
  INVX0 U6168 ( .INP(n4608), .ZN(n4194) );
  OR2X1 U6169 ( .IN1(n3058), .IN2(n5670), .Q(n4608) );
  OR2X1 U6170 ( .IN1(n3107), .IN2(n650), .Q(n5670) );
  INVX0 U6171 ( .INP(g109), .ZN(n650) );
  AND2X1 U6172 ( .IN1(g109), .IN2(g10721), .Q(n5411) );
  AND2X1 U6173 ( .IN1(n5671), .IN2(g109), .Q(n5668) );
  OR2X1 U6174 ( .IN1(n5672), .IN2(n5673), .Q(n5671) );
  OR2X1 U6175 ( .IN1(n5674), .IN2(n5675), .Q(n5673) );
  AND2X1 U6176 ( .IN1(g881), .IN2(g10720), .Q(n5675) );
  AND2X1 U6177 ( .IN1(g877), .IN2(g10719), .Q(n5674) );
  OR2X1 U6178 ( .IN1(n5676), .IN2(n5677), .Q(n5672) );
  AND2X1 U6179 ( .IN1(n3064), .IN2(n5410), .Q(n5677) );
  AND2X1 U6180 ( .IN1(g109), .IN2(g10722), .Q(n5410) );
  OR2X1 U6181 ( .IN1(n5678), .IN2(n5679), .Q(g10722) );
  OR2X1 U6182 ( .IN1(n5680), .IN2(n5681), .Q(n5679) );
  OR2X1 U6183 ( .IN1(n5682), .IN2(n5683), .Q(n5681) );
  OR2X1 U6184 ( .IN1(n5684), .IN2(n5685), .Q(n5683) );
  AND2X1 U6185 ( .IN1(n1486), .IN2(g1534), .Q(n5685) );
  AND2X1 U6186 ( .IN1(n1485), .IN2(g1577), .Q(n5684) );
  OR2X1 U6187 ( .IN1(n5686), .IN2(n5687), .Q(n5682) );
  OR2X1 U6188 ( .IN1(n5688), .IN2(n5689), .Q(n5687) );
  AND2X1 U6189 ( .IN1(n1512), .IN2(g1203), .Q(n5689) );
  AND2X1 U6190 ( .IN1(n1480), .IN2(g1601), .Q(n5688) );
  AND2X1 U6191 ( .IN1(n1479), .IN2(g1558), .Q(n5686) );
  OR2X1 U6192 ( .IN1(n5690), .IN2(n5691), .Q(n5680) );
  OR2X1 U6193 ( .IN1(n5692), .IN2(n5693), .Q(n5691) );
  AND2X1 U6194 ( .IN1(n5531), .IN2(n3048), .Q(n5693) );
  AND2X1 U6195 ( .IN1(n5694), .IN2(g1753), .Q(n5692) );
  OR2X1 U6196 ( .IN1(n5695), .IN2(n5696), .Q(n5690) );
  OR2X1 U6197 ( .IN1(n5697), .IN2(n5698), .Q(n5696) );
  AND2X1 U6198 ( .IN1(g1179), .IN2(n5638), .Q(n5698) );
  AND2X1 U6199 ( .IN1(n5699), .IN2(g1324), .Q(n5697) );
  AND2X1 U6200 ( .IN1(n5645), .IN2(g1730), .Q(n5695) );
  OR2X1 U6201 ( .IN1(n5700), .IN2(n5701), .Q(n5678) );
  OR2X1 U6202 ( .IN1(n5702), .IN2(n5703), .Q(n5701) );
  OR2X1 U6203 ( .IN1(n5704), .IN2(n5705), .Q(n5703) );
  AND2X1 U6204 ( .IN1(n5653), .IN2(g1351), .Q(n5705) );
  AND2X1 U6205 ( .IN1(n5666), .IN2(g986), .Q(n5704) );
  OR2X1 U6206 ( .IN1(n5706), .IN2(n5707), .Q(n5702) );
  OR2X1 U6207 ( .IN1(n5708), .IN2(n5709), .Q(n5707) );
  AND2X1 U6208 ( .IN1(n5710), .IN2(g296), .Q(n5709) );
  AND2X1 U6209 ( .IN1(n5665), .IN2(g272), .Q(n5708) );
  AND2X1 U6210 ( .IN1(g907), .IN2(n5664), .Q(n5706) );
  OR2X1 U6211 ( .IN1(n5711), .IN2(n5712), .Q(n5700) );
  OR2X1 U6212 ( .IN1(n5713), .IN2(n5714), .Q(n5712) );
  OR2X1 U6213 ( .IN1(n5715), .IN2(n5716), .Q(n5714) );
  AND2X1 U6214 ( .IN1(n5717), .IN2(g8), .Q(n5716) );
  AND2X1 U6215 ( .IN1(g895), .IN2(n5718), .Q(n5715) );
  AND2X1 U6216 ( .IN1(n5719), .IN2(n1631), .Q(n5713) );
  OR2X1 U6217 ( .IN1(n5720), .IN2(n5721), .Q(n5711) );
  OR2X1 U6218 ( .IN1(n5722), .IN2(n5723), .Q(n5721) );
  AND2X1 U6219 ( .IN1(n5724), .IN2(g940), .Q(n5723) );
  AND2X1 U6220 ( .IN1(n3579), .IN2(g959), .Q(n5720) );
  AND2X1 U6221 ( .IN1(n5725), .IN2(n6002), .Q(n5676) );
  AND2X1 U6222 ( .IN1(g10724), .IN2(g3007), .Q(n5725) );
  OR2X1 U6223 ( .IN1(g10726), .IN2(n3580), .Q(g10465) );
  OR2X1 U6224 ( .IN1(n5726), .IN2(n5727), .Q(g10726) );
  OR2X1 U6225 ( .IN1(n5728), .IN2(n5729), .Q(n5727) );
  OR2X1 U6226 ( .IN1(n5730), .IN2(n5731), .Q(n5729) );
  OR2X1 U6227 ( .IN1(n5732), .IN2(n5733), .Q(n5731) );
  AND2X1 U6228 ( .IN1(n1485), .IN2(g1583), .Q(n5733) );
  AND2X1 U6229 ( .IN1(n1479), .IN2(g1564), .Q(n5732) );
  AND2X1 U6230 ( .IN1(n1486), .IN2(g1540), .Q(n5730) );
  OR2X1 U6231 ( .IN1(n5734), .IN2(n5735), .Q(n5728) );
  OR2X1 U6232 ( .IN1(n5736), .IN2(n5737), .Q(n5735) );
  AND2X1 U6233 ( .IN1(n5531), .IN2(n1650), .Q(n5737) );
  AND2X1 U6234 ( .IN1(n5694), .IN2(g1759), .Q(n5736) );
  AND2X1 U6235 ( .IN1(n1480), .IN2(g1607), .Q(n5734) );
  OR2X1 U6236 ( .IN1(n5738), .IN2(n5739), .Q(n5726) );
  OR2X1 U6237 ( .IN1(n5740), .IN2(n5741), .Q(n5739) );
  OR2X1 U6238 ( .IN1(n5742), .IN2(n5743), .Q(n5741) );
  AND2X1 U6239 ( .IN1(n5699), .IN2(g1330), .Q(n5743) );
  AND2X1 U6240 ( .IN1(g1185), .IN2(n5638), .Q(n5740) );
  OR2X1 U6241 ( .IN1(n5744), .IN2(n5745), .Q(n5738) );
  OR2X1 U6242 ( .IN1(n5746), .IN2(n5747), .Q(n5745) );
  AND2X1 U6243 ( .IN1(g913), .IN2(n5664), .Q(n5747) );
  AND2X1 U6244 ( .IN1(n5710), .IN2(g302), .Q(n5746) );
  OR2X1 U6245 ( .IN1(n5748), .IN2(n5749), .Q(n5744) );
  AND2X1 U6246 ( .IN1(n5665), .IN2(g278), .Q(n5749) );
  AND2X1 U6247 ( .IN1(n3579), .IN2(g965), .Q(n5748) );
  OR2X1 U6248 ( .IN1(g10724), .IN2(n3580), .Q(g10463) );
  OR2X1 U6249 ( .IN1(n5750), .IN2(n5751), .Q(g10724) );
  OR2X1 U6250 ( .IN1(n5752), .IN2(n5753), .Q(n5751) );
  OR2X1 U6251 ( .IN1(n5754), .IN2(n5755), .Q(n5753) );
  OR2X1 U6252 ( .IN1(n5756), .IN2(n5757), .Q(n5755) );
  AND2X1 U6253 ( .IN1(n1486), .IN2(g1537), .Q(n5757) );
  AND2X1 U6254 ( .IN1(n1485), .IN2(g1580), .Q(n5756) );
  OR2X1 U6255 ( .IN1(n5758), .IN2(n5759), .Q(n5754) );
  INVX0 U6256 ( .INP(n5760), .ZN(n5759) );
  AND2X1 U6257 ( .IN1(n5717), .IN2(n3025), .Q(n5758) );
  OR2X1 U6258 ( .IN1(n5761), .IN2(n5762), .Q(n5752) );
  OR2X1 U6259 ( .IN1(n5763), .IN2(n5764), .Q(n5762) );
  AND2X1 U6260 ( .IN1(n1479), .IN2(g1561), .Q(n5764) );
  AND2X1 U6261 ( .IN1(n1480), .IN2(g1604), .Q(n5763) );
  OR2X1 U6262 ( .IN1(n5765), .IN2(n5766), .Q(n5761) );
  AND2X1 U6263 ( .IN1(n5531), .IN2(n3034), .Q(n5766) );
  AND2X1 U6264 ( .IN1(n5694), .IN2(g1756), .Q(n5765) );
  OR2X1 U6265 ( .IN1(n5767), .IN2(n5768), .Q(n5750) );
  OR2X1 U6266 ( .IN1(n5769), .IN2(n5770), .Q(n5768) );
  OR2X1 U6267 ( .IN1(n5771), .IN2(n5772), .Q(n5770) );
  AND2X1 U6268 ( .IN1(n5645), .IN2(g1733), .Q(n5772) );
  AND2X1 U6269 ( .IN1(g1182), .IN2(n5638), .Q(n5771) );
  OR2X1 U6270 ( .IN1(n5773), .IN2(n5774), .Q(n5769) );
  AND2X1 U6271 ( .IN1(n5699), .IN2(g1327), .Q(n5774) );
  AND2X1 U6272 ( .IN1(g910), .IN2(n5664), .Q(n5773) );
  OR2X1 U6273 ( .IN1(n5775), .IN2(n5776), .Q(n5767) );
  OR2X1 U6274 ( .IN1(n5777), .IN2(n5778), .Q(n5776) );
  AND2X1 U6275 ( .IN1(n5710), .IN2(g299), .Q(n5778) );
  AND2X1 U6276 ( .IN1(n5665), .IN2(g275), .Q(n5777) );
  OR2X1 U6277 ( .IN1(n5779), .IN2(n5780), .Q(n5775) );
  AND2X1 U6278 ( .IN1(n5719), .IN2(n3057), .Q(n5780) );
  AND2X1 U6279 ( .IN1(n3579), .IN2(g962), .Q(n5779) );
  OR2X1 U6280 ( .IN1(g10721), .IN2(n3580), .Q(g10459) );
  OR2X1 U6281 ( .IN1(n5781), .IN2(n5782), .Q(g10721) );
  OR2X1 U6282 ( .IN1(n5783), .IN2(n5784), .Q(n5782) );
  OR2X1 U6283 ( .IN1(n5785), .IN2(n5786), .Q(n5784) );
  OR2X1 U6284 ( .IN1(n5787), .IN2(n5788), .Q(n5786) );
  AND2X1 U6285 ( .IN1(n1486), .IN2(g1531), .Q(n5788) );
  AND2X1 U6286 ( .IN1(n1485), .IN2(g1574), .Q(n5787) );
  OR2X1 U6287 ( .IN1(n5789), .IN2(n5790), .Q(n5785) );
  OR2X1 U6288 ( .IN1(n5791), .IN2(n5792), .Q(n5790) );
  AND2X1 U6289 ( .IN1(g1200), .IN2(n1512), .Q(n5792) );
  AND2X1 U6290 ( .IN1(n1480), .IN2(g1598), .Q(n5791) );
  AND2X1 U6291 ( .IN1(n1479), .IN2(g1555), .Q(n5789) );
  OR2X1 U6292 ( .IN1(n5793), .IN2(n5794), .Q(n5783) );
  OR2X1 U6293 ( .IN1(n5795), .IN2(n5796), .Q(n5794) );
  AND2X1 U6294 ( .IN1(n5531), .IN2(n3045), .Q(n5796) );
  AND2X1 U6295 ( .IN1(n5694), .IN2(g1750), .Q(n5795) );
  OR2X1 U6296 ( .IN1(n5797), .IN2(n5798), .Q(n5793) );
  OR2X1 U6297 ( .IN1(n5799), .IN2(n5800), .Q(n5798) );
  AND2X1 U6298 ( .IN1(g1176), .IN2(n5638), .Q(n5800) );
  AND2X1 U6299 ( .IN1(n5699), .IN2(g1321), .Q(n5799) );
  AND2X1 U6300 ( .IN1(n5645), .IN2(g1727), .Q(n5797) );
  OR2X1 U6301 ( .IN1(n5801), .IN2(n5802), .Q(n5781) );
  OR2X1 U6302 ( .IN1(n5803), .IN2(n5804), .Q(n5802) );
  OR2X1 U6303 ( .IN1(n5805), .IN2(n5806), .Q(n5804) );
  AND2X1 U6304 ( .IN1(n5653), .IN2(g1346), .Q(n5806) );
  AND2X1 U6305 ( .IN1(n5666), .IN2(g981), .Q(n5805) );
  OR2X1 U6306 ( .IN1(n5807), .IN2(n5808), .Q(n5803) );
  OR2X1 U6307 ( .IN1(n5809), .IN2(n5810), .Q(n5808) );
  AND2X1 U6308 ( .IN1(n5710), .IN2(g293), .Q(n5810) );
  AND2X1 U6309 ( .IN1(n5665), .IN2(g269), .Q(n5809) );
  AND2X1 U6310 ( .IN1(g904), .IN2(n5664), .Q(n5807) );
  OR2X1 U6311 ( .IN1(n5811), .IN2(n5812), .Q(n5801) );
  OR2X1 U6312 ( .IN1(n5813), .IN2(n5814), .Q(n5812) );
  OR2X1 U6313 ( .IN1(n5815), .IN2(n5816), .Q(n5814) );
  AND2X1 U6314 ( .IN1(n5717), .IN2(g1), .Q(n5816) );
  AND2X1 U6315 ( .IN1(g892), .IN2(n5718), .Q(n5815) );
  AND2X1 U6316 ( .IN1(n5719), .IN2(g9), .Q(n5813) );
  OR2X1 U6317 ( .IN1(n5817), .IN2(n5818), .Q(n5811) );
  OR2X1 U6318 ( .IN1(n5722), .IN2(n5819), .Q(n5818) );
  AND2X1 U6319 ( .IN1(n5724), .IN2(g936), .Q(n5819) );
  AND2X1 U6320 ( .IN1(n3579), .IN2(g956), .Q(n5817) );
  OR2X1 U6321 ( .IN1(g10720), .IN2(n3580), .Q(g10457) );
  OR2X1 U6322 ( .IN1(n5820), .IN2(n5821), .Q(g10720) );
  OR2X1 U6323 ( .IN1(n5822), .IN2(n5823), .Q(n5821) );
  OR2X1 U6324 ( .IN1(n5824), .IN2(n5825), .Q(n5823) );
  OR2X1 U6325 ( .IN1(n5826), .IN2(n5827), .Q(n5825) );
  AND2X1 U6326 ( .IN1(n1486), .IN2(g1528), .Q(n5827) );
  AND2X1 U6327 ( .IN1(n1485), .IN2(g1571), .Q(n5826) );
  OR2X1 U6328 ( .IN1(n5828), .IN2(n5829), .Q(n5824) );
  OR2X1 U6329 ( .IN1(n5830), .IN2(n5831), .Q(n5829) );
  AND2X1 U6330 ( .IN1(n1530), .IN2(g925), .Q(n5831) );
  AND2X1 U6331 ( .IN1(g1197), .IN2(n1512), .Q(n5830) );
  AND2X1 U6332 ( .IN1(n1479), .IN2(g1552), .Q(n5828) );
  OR2X1 U6333 ( .IN1(n5832), .IN2(n5833), .Q(n5822) );
  OR2X1 U6334 ( .IN1(n5834), .IN2(n5835), .Q(n5833) );
  OR2X1 U6335 ( .IN1(n5836), .IN2(n5837), .Q(n5835) );
  AND2X1 U6336 ( .IN1(n5531), .IN2(n3031), .Q(n5837) );
  AND2X1 U6337 ( .IN1(n5694), .IN2(g1747), .Q(n5836) );
  AND2X1 U6338 ( .IN1(n1480), .IN2(g1595), .Q(n5834) );
  OR2X1 U6339 ( .IN1(n5838), .IN2(n5839), .Q(n5832) );
  OR2X1 U6340 ( .IN1(n5840), .IN2(n5841), .Q(n5839) );
  AND2X1 U6341 ( .IN1(g1173), .IN2(n5638), .Q(n5841) );
  AND2X1 U6342 ( .IN1(n5699), .IN2(g1318), .Q(n5840) );
  AND2X1 U6343 ( .IN1(n5645), .IN2(g1724), .Q(n5838) );
  OR2X1 U6344 ( .IN1(n5842), .IN2(n5843), .Q(n5820) );
  OR2X1 U6345 ( .IN1(n5844), .IN2(n5845), .Q(n5843) );
  OR2X1 U6346 ( .IN1(n5846), .IN2(n5847), .Q(n5845) );
  AND2X1 U6347 ( .IN1(n5653), .IN2(g1341), .Q(n5847) );
  AND2X1 U6348 ( .IN1(n5666), .IN2(g976), .Q(n5846) );
  OR2X1 U6349 ( .IN1(n5848), .IN2(n5849), .Q(n5844) );
  OR2X1 U6350 ( .IN1(n5850), .IN2(n5851), .Q(n5849) );
  AND2X1 U6351 ( .IN1(n5710), .IN2(g290), .Q(n5851) );
  AND2X1 U6352 ( .IN1(n5665), .IN2(g266), .Q(n5850) );
  AND2X1 U6353 ( .IN1(g901), .IN2(n5664), .Q(n5848) );
  OR2X1 U6354 ( .IN1(n5852), .IN2(n5853), .Q(n5842) );
  OR2X1 U6355 ( .IN1(n5854), .IN2(n5855), .Q(n5853) );
  OR2X1 U6356 ( .IN1(n5856), .IN2(n5857), .Q(n5855) );
  AND2X1 U6357 ( .IN1(n5717), .IN2(g4), .Q(n5857) );
  AND2X1 U6358 ( .IN1(g889), .IN2(n5718), .Q(n5856) );
  AND2X1 U6359 ( .IN1(n5719), .IN2(g12), .Q(n5854) );
  OR2X1 U6360 ( .IN1(n5858), .IN2(n5859), .Q(n5852) );
  OR2X1 U6361 ( .IN1(n5722), .IN2(n5860), .Q(n5859) );
  AND2X1 U6362 ( .IN1(n5724), .IN2(g932), .Q(n5860) );
  AND2X1 U6363 ( .IN1(n3579), .IN2(g953), .Q(n5858) );
  OR2X1 U6364 ( .IN1(g10719), .IN2(n3580), .Q(g10455) );
  OR2X1 U6365 ( .IN1(n5861), .IN2(n5862), .Q(g10719) );
  OR2X1 U6366 ( .IN1(n5863), .IN2(n5864), .Q(n5862) );
  OR2X1 U6367 ( .IN1(n5865), .IN2(n5866), .Q(n5864) );
  OR2X1 U6368 ( .IN1(n5867), .IN2(n5868), .Q(n5866) );
  AND2X1 U6369 ( .IN1(n1486), .IN2(g1524), .Q(n5868) );
  AND2X1 U6370 ( .IN1(n1485), .IN2(g1567), .Q(n5867) );
  OR2X1 U6371 ( .IN1(n5869), .IN2(n5870), .Q(n5865) );
  OR2X1 U6372 ( .IN1(n5871), .IN2(n5872), .Q(n5870) );
  AND2X1 U6373 ( .IN1(g922), .IN2(n1530), .Q(n5872) );
  AND2X1 U6374 ( .IN1(g1194), .IN2(n1512), .Q(n5871) );
  AND2X1 U6375 ( .IN1(n1479), .IN2(g1549), .Q(n5869) );
  OR2X1 U6376 ( .IN1(n5873), .IN2(n5874), .Q(n5863) );
  OR2X1 U6377 ( .IN1(n5875), .IN2(n5876), .Q(n5874) );
  OR2X1 U6378 ( .IN1(n5877), .IN2(n5878), .Q(n5876) );
  AND2X1 U6379 ( .IN1(n5531), .IN2(n3051), .Q(n5878) );
  AND2X1 U6380 ( .IN1(n5694), .IN2(g1744), .Q(n5877) );
  AND2X1 U6381 ( .IN1(n1480), .IN2(g1592), .Q(n5875) );
  OR2X1 U6382 ( .IN1(n5879), .IN2(n5880), .Q(n5873) );
  OR2X1 U6383 ( .IN1(n5881), .IN2(n5882), .Q(n5880) );
  AND2X1 U6384 ( .IN1(g1170), .IN2(n5638), .Q(n5882) );
  AND2X1 U6385 ( .IN1(n5699), .IN2(g1314), .Q(n5881) );
  AND2X1 U6386 ( .IN1(n5645), .IN2(g1721), .Q(n5879) );
  OR2X1 U6387 ( .IN1(n5883), .IN2(n5884), .Q(n5861) );
  OR2X1 U6388 ( .IN1(n5885), .IN2(n5886), .Q(n5884) );
  OR2X1 U6389 ( .IN1(n5887), .IN2(n5888), .Q(n5886) );
  OR2X1 U6390 ( .IN1(n5889), .IN2(n5890), .Q(n5888) );
  AND2X1 U6391 ( .IN1(n5666), .IN2(g971), .Q(n5890) );
  AND2X1 U6392 ( .IN1(g898), .IN2(n5664), .Q(n5889) );
  AND2X1 U6393 ( .IN1(n5653), .IN2(g1336), .Q(n5887) );
  OR2X1 U6394 ( .IN1(n5891), .IN2(n5892), .Q(n5885) );
  OR2X1 U6395 ( .IN1(n5893), .IN2(n5894), .Q(n5892) );
  AND2X1 U6396 ( .IN1(n5665), .IN2(g263), .Q(n5894) );
  AND2X1 U6397 ( .IN1(n5719), .IN2(g119), .Q(n5893) );
  AND2X1 U6398 ( .IN1(n5710), .IN2(g287), .Q(n5891) );
  INVX0 U6399 ( .INP(n5895), .ZN(n5710) );
  OR2X1 U6400 ( .IN1(n5896), .IN2(n5897), .Q(n5883) );
  OR2X1 U6401 ( .IN1(n5898), .IN2(n5899), .Q(n5897) );
  OR2X1 U6402 ( .IN1(n5900), .IN2(n5901), .Q(n5899) );
  AND2X1 U6403 ( .IN1(g886), .IN2(n5718), .Q(n5901) );
  AND2X1 U6404 ( .IN1(n3579), .IN2(g950), .Q(n5900) );
  AND2X1 U6405 ( .IN1(n5717), .IN2(g123), .Q(n5898) );
  OR2X1 U6406 ( .IN1(n5902), .IN2(n5903), .Q(n5896) );
  OR2X1 U6407 ( .IN1(n656), .IN2(n5722), .Q(n5903) );
  INVX0 U6408 ( .INP(n5904), .ZN(n5722) );
  OR2X1 U6409 ( .IN1(n5905), .IN2(n5760), .Q(n5904) );
  OR2X1 U6410 ( .IN1(n5906), .IN2(n5717), .Q(n5760) );
  AND2X1 U6411 ( .IN1(g42), .IN2(n5907), .Q(n5717) );
  OR2X1 U6412 ( .IN1(n5908), .IN2(n5909), .Q(n5906) );
  OR2X1 U6413 ( .IN1(n3581), .IN2(n5910), .Q(n5909) );
  OR2X1 U6414 ( .IN1(n5911), .IN2(n5912), .Q(n3581) );
  OR2X1 U6415 ( .IN1(n5913), .IN2(n5914), .Q(n5912) );
  OR2X1 U6416 ( .IN1(n5724), .IN2(n5531), .Q(n5914) );
  OR2X1 U6417 ( .IN1(n5915), .IN2(n5718), .Q(n5913) );
  INVX0 U6418 ( .INP(n5916), .ZN(n5718) );
  OR2X1 U6419 ( .IN1(n5917), .IN2(n5918), .Q(n5916) );
  OR2X1 U6420 ( .IN1(g44), .IN2(n5919), .Q(n5918) );
  OR2X1 U6421 ( .IN1(n5920), .IN2(n5921), .Q(n5911) );
  OR2X1 U6422 ( .IN1(n5664), .IN2(n3579), .Q(n5921) );
  AND2X1 U6423 ( .IN1(n5922), .IN2(n666), .Q(n3579) );
  OR2X1 U6424 ( .IN1(n1530), .IN2(n5666), .Q(n5920) );
  OR2X1 U6425 ( .IN1(n5719), .IN2(n656), .Q(n5908) );
  AND2X1 U6426 ( .IN1(n5475), .IN2(n5907), .Q(n5719) );
  INVX0 U6427 ( .INP(n5923), .ZN(n5907) );
  OR2X1 U6428 ( .IN1(n5924), .IN2(n5925), .Q(n5923) );
  OR2X1 U6429 ( .IN1(n5650), .IN2(n5919), .Q(n5925) );
  OR2X1 U6430 ( .IN1(g45), .IN2(g44), .Q(n5924) );
  OR2X1 U6431 ( .IN1(n1512), .IN2(n5653), .Q(n5905) );
  AND2X1 U6432 ( .IN1(n5724), .IN2(g928), .Q(n5902) );
  INVX0 U6433 ( .INP(n5926), .ZN(n5724) );
  OR2X1 U6434 ( .IN1(n5917), .IN2(n5927), .Q(n5926) );
  OR2X1 U6435 ( .IN1(g43), .IN2(n5928), .Q(n5927) );
  OR2X1 U6436 ( .IN1(n5929), .IN2(n5930), .Q(n5917) );
  OR2X1 U6437 ( .IN1(g10663), .IN2(n3580), .Q(g10377) );
  OR2X1 U6438 ( .IN1(g30), .IN2(n5531), .Q(n3580) );
  OR2X1 U6439 ( .IN1(n5931), .IN2(n5932), .Q(g10663) );
  OR2X1 U6440 ( .IN1(n5933), .IN2(n5934), .Q(n5932) );
  OR2X1 U6441 ( .IN1(n5935), .IN2(n5936), .Q(n5934) );
  OR2X1 U6442 ( .IN1(n5937), .IN2(n5938), .Q(n5936) );
  AND2X1 U6443 ( .IN1(n1486), .IN2(g1543), .Q(n5938) );
  AND2X1 U6444 ( .IN1(n1485), .IN2(g1586), .Q(n5937) );
  OR2X1 U6445 ( .IN1(n5939), .IN2(n5940), .Q(n5935) );
  AND2X1 U6446 ( .IN1(n5742), .IN2(n5648), .Q(n5940) );
  AND2X1 U6447 ( .IN1(n1478), .IN2(n5941), .Q(n5742) );
  INVX0 U6448 ( .INP(n5910), .ZN(n5941) );
  OR2X1 U6449 ( .IN1(n5942), .IN2(n5943), .Q(n5910) );
  OR2X1 U6450 ( .IN1(n5699), .IN2(n5944), .Q(n5943) );
  OR2X1 U6451 ( .IN1(n5645), .IN2(n5638), .Q(n5944) );
  OR2X1 U6452 ( .IN1(n5694), .IN2(n5945), .Q(n5942) );
  OR2X1 U6453 ( .IN1(n1567), .IN2(n1566), .Q(n5945) );
  OR2X1 U6454 ( .IN1(n5946), .IN2(n1479), .Q(n1566) );
  AND2X1 U6455 ( .IN1(n5947), .IN2(n661), .Q(n5946) );
  OR2X1 U6456 ( .IN1(n5948), .IN2(n1480), .Q(n1567) );
  AND2X1 U6457 ( .IN1(n661), .IN2(n5922), .Q(n1480) );
  AND2X1 U6458 ( .IN1(n661), .IN2(n5949), .Q(n5948) );
  INVX0 U6459 ( .INP(n5650), .ZN(n661) );
  AND2X1 U6460 ( .IN1(n5653), .IN2(g1308), .Q(n5939) );
  INVX0 U6461 ( .INP(n5648), .ZN(n5653) );
  OR2X1 U6462 ( .IN1(n5950), .IN2(n5652), .Q(n5648) );
  OR2X1 U6463 ( .IN1(n5951), .IN2(n5952), .Q(n5933) );
  OR2X1 U6464 ( .IN1(n5953), .IN2(n5954), .Q(n5952) );
  AND2X1 U6465 ( .IN1(n5694), .IN2(g1762), .Q(n5954) );
  AND2X1 U6466 ( .IN1(n5475), .IN2(n5955), .Q(n5694) );
  AND2X1 U6467 ( .IN1(n5645), .IN2(g1738), .Q(n5953) );
  AND2X1 U6468 ( .IN1(g42), .IN2(n5955), .Q(n5645) );
  INVX0 U6469 ( .INP(n5956), .ZN(n5955) );
  OR2X1 U6470 ( .IN1(n5957), .IN2(n5958), .Q(n5956) );
  OR2X1 U6471 ( .IN1(n5919), .IN2(n5928), .Q(n5958) );
  OR2X1 U6472 ( .IN1(n5959), .IN2(n5950), .Q(n5957) );
  AND2X1 U6473 ( .IN1(n5531), .IN2(n1637), .Q(n5951) );
  OR2X1 U6474 ( .IN1(n5960), .IN2(n5961), .Q(n5931) );
  OR2X1 U6475 ( .IN1(n5962), .IN2(n5963), .Q(n5961) );
  OR2X1 U6476 ( .IN1(n5964), .IN2(n5965), .Q(n5963) );
  AND2X1 U6477 ( .IN1(n5699), .IN2(g1333), .Q(n5965) );
  AND2X1 U6478 ( .IN1(n660), .IN2(n5922), .Q(n5699) );
  INVX0 U6479 ( .INP(n5966), .ZN(n5922) );
  OR2X1 U6480 ( .IN1(n5477), .IN2(n5967), .Q(n5966) );
  OR2X1 U6481 ( .IN1(g42), .IN2(n5959), .Q(n5967) );
  INVX0 U6482 ( .INP(n5950), .ZN(n660) );
  AND2X1 U6483 ( .IN1(n5666), .IN2(g944), .Q(n5964) );
  AND2X1 U6484 ( .IN1(n5949), .IN2(n666), .Q(n5666) );
  INVX0 U6485 ( .INP(n5652), .ZN(n5949) );
  OR2X1 U6486 ( .IN1(n5477), .IN2(n5930), .Q(n5652) );
  OR2X1 U6487 ( .IN1(n5475), .IN2(n5959), .Q(n5930) );
  INVX0 U6488 ( .INP(g45), .ZN(n5959) );
  OR2X1 U6489 ( .IN1(g44), .IN2(g43), .Q(n5477) );
  AND2X1 U6490 ( .IN1(g1188), .IN2(n5638), .Q(n5962) );
  INVX0 U6491 ( .INP(n5640), .ZN(n5638) );
  OR2X1 U6492 ( .IN1(n5950), .IN2(n5651), .Q(n5640) );
  OR2X1 U6493 ( .IN1(n5968), .IN2(n3594), .Q(n5950) );
  OR2X1 U6494 ( .IN1(n5969), .IN2(n5970), .Q(n3594) );
  OR2X1 U6495 ( .IN1(g46), .IN2(n3617), .Q(n5970) );
  OR2X1 U6496 ( .IN1(n5971), .IN2(n5972), .Q(n5960) );
  OR2X1 U6497 ( .IN1(n5973), .IN2(n5974), .Q(n5972) );
  AND2X1 U6498 ( .IN1(g916), .IN2(n5664), .Q(n5974) );
  AND2X1 U6499 ( .IN1(n5947), .IN2(n666), .Q(n5664) );
  INVX0 U6500 ( .INP(n5929), .ZN(n666) );
  OR2X1 U6501 ( .IN1(n5968), .IN2(n3592), .Q(n5929) );
  OR2X1 U6502 ( .IN1(n5474), .IN2(n5975), .Q(n3592) );
  INVX0 U6503 ( .INP(n5651), .ZN(n5947) );
  OR2X1 U6504 ( .IN1(n5976), .IN2(n5977), .Q(n5651) );
  OR2X1 U6505 ( .IN1(n5475), .IN2(n5919), .Q(n5977) );
  INVX0 U6506 ( .INP(g42), .ZN(n5475) );
  AND2X1 U6507 ( .IN1(n5665), .IN2(g281), .Q(n5973) );
  AND2X1 U6508 ( .IN1(n5895), .IN2(n5915), .Q(n5665) );
  INVX0 U6509 ( .INP(n5978), .ZN(n5915) );
  OR2X1 U6510 ( .IN1(n5976), .IN2(n5979), .Q(n5978) );
  OR2X1 U6511 ( .IN1(g43), .IN2(n5650), .Q(n5979) );
  OR2X1 U6512 ( .IN1(n5980), .IN2(n5981), .Q(n5895) );
  OR2X1 U6513 ( .IN1(n5650), .IN2(n5976), .Q(n5981) );
  OR2X1 U6514 ( .IN1(n5474), .IN2(n5982), .Q(n5650) );
  OR2X1 U6515 ( .IN1(g46), .IN2(n5968), .Q(n5982) );
  OR2X1 U6516 ( .IN1(n3617), .IN2(g47), .Q(n5474) );
  OR2X1 U6517 ( .IN1(g43), .IN2(g42), .Q(n5980) );
  OR2X1 U6518 ( .IN1(n1564), .IN2(n656), .Q(n5971) );
  INVX0 U6519 ( .INP(n5983), .ZN(n656) );
  OR2X1 U6520 ( .IN1(n5984), .IN2(n5985), .Q(n5983) );
  OR2X1 U6521 ( .IN1(n5969), .IN2(n5975), .Q(n5985) );
  INVX0 U6522 ( .INP(g46), .ZN(n5975) );
  INVX0 U6523 ( .INP(g47), .ZN(n5969) );
  OR2X1 U6524 ( .IN1(n5968), .IN2(n5986), .Q(n5984) );
  OR2X1 U6525 ( .IN1(n1545), .IN2(n3617), .Q(n5986) );
  AND2X1 U6526 ( .IN1(n5987), .IN2(n5988), .Q(n3617) );
  OR2X1 U6527 ( .IN1(n5968), .IN2(n5531), .Q(n5988) );
  OR2X1 U6528 ( .IN1(g31), .IN2(n5989), .Q(n5531) );
  OR2X1 U6529 ( .IN1(n5990), .IN2(g30), .Q(n5987) );
  OR2X1 U6530 ( .IN1(g41), .IN2(g48), .Q(n5990) );
  OR2X1 U6531 ( .IN1(n5976), .IN2(n5991), .Q(n1545) );
  OR2X1 U6532 ( .IN1(g42), .IN2(n5919), .Q(n5991) );
  INVX0 U6533 ( .INP(g43), .ZN(n5919) );
  OR2X1 U6534 ( .IN1(g45), .IN2(n5928), .Q(n5976) );
  INVX0 U6535 ( .INP(g44), .ZN(n5928) );
  OR2X1 U6536 ( .IN1(g41), .IN2(n5989), .Q(n5968) );
  INVX0 U6537 ( .INP(g48), .ZN(n5989) );
  OR2X1 U6538 ( .IN1(n5992), .IN2(n5993), .Q(N599) );
  INVX0 U6539 ( .INP(n5994), .ZN(n5993) );
  OR2X1 U6540 ( .IN1(n4168), .IN2(test_so1), .Q(n5994) );
  AND2X1 U6541 ( .IN1(test_so1), .IN2(n4168), .Q(n5992) );
  OR2X1 U6542 ( .IN1(n4287), .IN2(n5995), .Q(n4168) );
  OR2X1 U6543 ( .IN1(n3363), .IN2(n3345), .Q(n5995) );
  INVX0 U6544 ( .INP(n1093), .ZN(n4287) );
  OR2X1 U1550_U1 ( .IN1(g10722), .IN2(n655), .Q(g10461) );
  OR2X1 U1551_U1 ( .IN1(g10664), .IN2(n655), .Q(g10379) );
  INVX0 U1586_U2 ( .INP(n3377), .ZN(U1586_n1) );
  AND2X1 U1586_U1 ( .IN1(n19), .IN2(U1586_n1), .Q(n1855) );
  INVX0 U1754_U2 ( .INP(n1545), .ZN(U1754_n1) );
  AND2X1 U1754_U1 ( .IN1(n661), .IN2(U1754_n1), .Q(n1479) );
  INVX0 U1798_U2 ( .INP(n1480), .ZN(U1798_n1) );
  AND2X1 U1798_U1 ( .IN1(n1567), .IN2(U1798_n1), .Q(n1485) );
  INVX0 U1839_U2 ( .INP(n1479), .ZN(U1839_n1) );
  AND2X1 U1839_U1 ( .IN1(n1566), .IN2(U1839_n1), .Q(n1486) );
  INVX0 U1843_U2 ( .INP(n656), .ZN(U1843_n1) );
  AND2X1 U1843_U1 ( .IN1(n628), .IN2(U1843_n1), .Q(n1478) );
  INVX0 U1877_U2 ( .INP(n650), .ZN(U1877_n1) );
  AND2X1 U1877_U1 ( .IN1(n1137), .IN2(U1877_n1), .Q(n1195) );
  INVX0 U1908_U2 ( .INP(n1545), .ZN(U1908_n1) );
  AND2X1 U1908_U1 ( .IN1(n660), .IN2(U1908_n1), .Q(n1512) );
  INVX0 U1909_U2 ( .INP(n1545), .ZN(U1909_n1) );
  AND2X1 U1909_U1 ( .IN1(n666), .IN2(U1909_n1), .Q(n1530) );
  INVX0 U1987_U2 ( .INP(n366), .ZN(U1987_n1) );
  AND2X1 U1987_U1 ( .IN1(n822), .IN2(U1987_n1), .Q(n916) );
  INVX0 U2031_U2 ( .INP(n493), .ZN(U2031_n1) );
  AND2X1 U2031_U1 ( .IN1(n180), .IN2(U2031_n1), .Q(n1056) );
  INVX0 U2035_U2 ( .INP(g109), .ZN(U2035_n1) );
  AND2X1 U2035_U1 ( .IN1(n1404), .IN2(U2035_n1), .Q(n1450) );
  INVX0 U2418_U2 ( .INP(n665), .ZN(U2418_n1) );
  AND2X1 U2418_U1 ( .IN1(g968), .IN2(U2418_n1), .Q(n1564) );
  INVX0 U2468_U2 ( .INP(n1227), .ZN(U2468_n1) );
  AND2X1 U2468_U1 ( .IN1(g1336), .IN2(U2468_n1), .Q(n1231) );
  INVX0 U2478_U2 ( .INP(n1229), .ZN(U2478_n1) );
  AND2X1 U2478_U1 ( .IN1(g1341), .IN2(U2478_n1), .Q(n1232) );
  INVX0 U2488_U2 ( .INP(n1258), .ZN(U2488_n1) );
  AND2X1 U2488_U1 ( .IN1(n1262), .IN2(U2488_n1), .Q(n1260) );
  INVX0 U2533_U2 ( .INP(n650), .ZN(U2533_n1) );
  AND2X1 U2533_U1 ( .IN1(g178), .IN2(U2533_n1), .Q(g6786) );
  INVX0 U2534_U2 ( .INP(n650), .ZN(U2534_n1) );
  AND2X1 U2534_U1 ( .IN1(g1424), .IN2(U2534_n1), .Q(g6234) );
  INVX0 U2639_U2 ( .INP(n958), .ZN(U2639_n1) );
  AND2X1 U2639_U1 ( .IN1(n962), .IN2(U2639_n1), .Q(n804) );
  INVX0 U2641_U2 ( .INP(g1868), .ZN(U2641_n1) );
  AND2X1 U2641_U1 ( .IN1(n102), .IN2(U2641_n1), .Q(n926) );
  INVX0 U2654_U2 ( .INP(g750), .ZN(U2654_n1) );
  AND2X1 U2654_U1 ( .IN1(g746), .IN2(U2654_n1), .Q(g4171) );
  INVX0 U2658_U2 ( .INP(n918), .ZN(U2658_n1) );
  AND2X1 U2658_U1 ( .IN1(n917), .IN2(U2658_n1), .Q(n812) );
  INVX0 U2683_U2 ( .INP(n1385), .ZN(U2683_n1) );
  AND2X1 U2683_U1 ( .IN1(g382), .IN2(U2683_n1), .Q(n1420) );
  INVX0 U2699_U2 ( .INP(n633), .ZN(U2699_n1) );
  AND2X1 U2699_U1 ( .IN1(n808), .IN2(U2699_n1), .Q(n806) );
  INVX0 U2846_U2 ( .INP(n1214), .ZN(U2846_n1) );
  AND2X1 U2846_U1 ( .IN1(g4175), .IN2(U2846_n1), .Q(n1193) );
  INVX0 U2847_U2 ( .INP(n1153), .ZN(U2847_n1) );
  AND2X1 U2847_U1 ( .IN1(g4177), .IN2(U2847_n1), .Q(n1125) );
  INVX0 U2848_U2 ( .INP(n1099), .ZN(U2848_n1) );
  AND2X1 U2848_U1 ( .IN1(g4179), .IN2(U2848_n1), .Q(n1093) );
  INVX0 U2859_U2 ( .INP(g12), .ZN(U2859_n1) );
  AND2X1 U2859_U1 ( .IN1(n1137), .IN2(U2859_n1), .Q(n1159) );
  INVX0 U2860_U2 ( .INP(n1151), .ZN(U2860_n1) );
  AND2X1 U2860_U1 ( .IN1(g810), .IN2(U2860_n1), .Q(n1123) );
  INVX0 U2861_U2 ( .INP(n1097), .ZN(U2861_n1) );
  AND2X1 U2861_U1 ( .IN1(g818), .IN2(U2861_n1), .Q(n1090) );
  INVX0 U2867_U2 ( .INP(g1834), .ZN(U2867_n1) );
  AND2X1 U2867_U1 ( .IN1(n817), .IN2(U2867_n1), .Q(n1380) );
  INVX0 U2879_U2 ( .INP(n1656), .ZN(U2879_n1) );
  AND2X1 U2879_U1 ( .IN1(g713), .IN2(U2879_n1), .Q(n967) );
  INVX0 U2881_U2 ( .INP(n1657), .ZN(U2881_n1) );
  AND2X1 U2881_U1 ( .IN1(g1927), .IN2(U2881_n1), .Q(n921) );
  INVX0 U2882_U2 ( .INP(n650), .ZN(U2882_n1) );
  AND2X1 U2882_U1 ( .IN1(g1160), .IN2(U2882_n1), .Q(g4334) );
  INVX0 U2883_U2 ( .INP(n650), .ZN(U2883_n1) );
  AND2X1 U2883_U1 ( .IN1(g1166), .IN2(U2883_n1), .Q(g4325) );
  INVX0 U2884_U2 ( .INP(n650), .ZN(U2884_n1) );
  AND2X1 U2884_U1 ( .IN1(g148), .IN2(U2884_n1), .Q(g6759) );
  INVX0 U2885_U2 ( .INP(n650), .ZN(U2885_n1) );
  AND2X1 U2885_U1 ( .IN1(g1157), .IN2(U2885_n1), .Q(g4338) );
  INVX0 U2886_U2 ( .INP(n650), .ZN(U2886_n1) );
  AND2X1 U2886_U1 ( .IN1(g1163), .IN2(U2886_n1), .Q(g4330) );
  INVX0 U2887_U2 ( .INP(n650), .ZN(U2887_n1) );
  AND2X1 U2887_U1 ( .IN1(g237), .IN2(U2887_n1), .Q(g6821) );
  INVX0 U2888_U2 ( .INP(n650), .ZN(U2888_n1) );
  AND2X1 U2888_U1 ( .IN1(g1499), .IN2(U2888_n1), .Q(g6198) );
  INVX0 U2889_U2 ( .INP(n650), .ZN(U2889_n1) );
  AND2X1 U2889_U1 ( .IN1(g1411), .IN2(U2889_n1), .Q(g6244) );
  INVX0 U2890_U2 ( .INP(n650), .ZN(U2890_n1) );
  AND2X1 U2890_U1 ( .IN1(g225), .IN2(U2890_n1), .Q(g6826) );
  INVX0 U2891_U2 ( .INP(n650), .ZN(U2891_n1) );
  AND2X1 U2891_U1 ( .IN1(g1407), .IN2(U2891_n1), .Q(g6216) );
  INVX0 U2892_U2 ( .INP(n650), .ZN(U2892_n1) );
  AND2X1 U2892_U1 ( .IN1(g213), .IN2(U2892_n1), .Q(g6829) );
  INVX0 U2893_U2 ( .INP(n650), .ZN(U2893_n1) );
  AND2X1 U2893_U1 ( .IN1(g186), .IN2(U2893_n1), .Q(g6833) );
  INVX0 U2894_U2 ( .INP(n650), .ZN(U2894_n1) );
  AND2X1 U2894_U1 ( .IN1(g219), .IN2(U2894_n1), .Q(g6827) );
  INVX0 U2895_U2 ( .INP(n650), .ZN(U2895_n1) );
  AND2X1 U2895_U1 ( .IN1(g143), .IN2(U2895_n1), .Q(g6757) );
  INVX0 U2896_U2 ( .INP(n650), .ZN(U2896_n1) );
  AND2X1 U2896_U1 ( .IN1(g207), .IN2(U2896_n1), .Q(g6831) );
  INVX0 U2897_U2 ( .INP(n650), .ZN(U2897_n1) );
  AND2X1 U2897_U1 ( .IN1(g231), .IN2(U2897_n1), .Q(g6822) );
  INVX0 U2898_U2 ( .INP(n650), .ZN(U2898_n1) );
  AND2X1 U2898_U1 ( .IN1(g192), .IN2(U2898_n1), .Q(g6838) );
  INVX0 U2899_U2 ( .INP(n650), .ZN(U2899_n1) );
  AND2X1 U2899_U1 ( .IN1(test_so3), .IN2(U2899_n1), .Q(g6823) );
  INVX0 U2900_U2 ( .INP(n650), .ZN(U2900_n1) );
  AND2X1 U2900_U1 ( .IN1(g1371), .IN2(U2900_n1), .Q(g6824) );
  INVX0 U2901_U2 ( .INP(n650), .ZN(U2901_n1) );
  AND2X1 U2901_U1 ( .IN1(g1383), .IN2(U2901_n1), .Q(g6832) );
  INVX0 U2902_U2 ( .INP(n650), .ZN(U2902_n1) );
  AND2X1 U2902_U1 ( .IN1(g243), .IN2(U2902_n1), .Q(g6819) );
  INVX0 U3090_U2 ( .INP(g810), .ZN(U3090_n1) );
  AND2X1 U3090_U1 ( .IN1(n1151), .IN2(U3090_n1), .Q(n1150) );
  INVX0 U3092_U2 ( .INP(g818), .ZN(U3092_n1) );
  AND2X1 U3092_U1 ( .IN1(n1097), .IN2(U3092_n1), .Q(n1096) );
  INVX0 U3094_U2 ( .INP(g4179), .ZN(U3094_n1) );
  AND2X1 U3094_U1 ( .IN1(n1099), .IN2(U3094_n1), .Q(n1098) );
  INVX0 U3096_U2 ( .INP(g4175), .ZN(U3096_n1) );
  AND2X1 U3096_U1 ( .IN1(n1214), .IN2(U3096_n1), .Q(n1213) );
  INVX0 U3098_U2 ( .INP(g4177), .ZN(U3098_n1) );
  AND2X1 U3098_U1 ( .IN1(n1153), .IN2(U3098_n1), .Q(n1152) );
  INVX0 U3124_U2 ( .INP(n838), .ZN(U3124_n1) );
  AND2X1 U3124_U1 ( .IN1(n837), .IN2(U3124_n1), .Q(n836) );
  INVX0 U3171_U2 ( .INP(n3382), .ZN(U3171_n1) );
  AND2X1 U3171_U1 ( .IN1(g1610), .IN2(U3171_n1), .Q(g5194) );
endmodule

