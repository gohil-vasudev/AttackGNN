module add_mul_sub_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, operation_0_, operation_1_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_
 );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783;

  INV_X1 U2374 ( .A(n2414), .ZN(n2342) );
  INV_X2 U2375 ( .A(n2342), .ZN(n2343) );
  INV_X1 U2376 ( .A(n2413), .ZN(n2344) );
  INV_X2 U2377 ( .A(n2344), .ZN(n2345) );
  INV_X1 U2378 ( .A(n2412), .ZN(n2346) );
  INV_X2 U2379 ( .A(n2346), .ZN(n2347) );
  INV_X1 U2380 ( .A(n2352), .ZN(n2348) );
  INV_X2 U2381 ( .A(n2348), .ZN(n2349) );
  NOR2_X2 U2382 ( .A1(n4579), .A2(n2428), .ZN(n2840) );
  NAND2_X1 U2383 ( .A1(n2350), .A2(n2351), .ZN(Result_9_) );
  NAND2_X1 U2384 ( .A1(n2349), .A2(n2353), .ZN(n2351) );
  XOR2_X1 U2385 ( .A(n2354), .B(n2355), .Z(n2353) );
  NAND2_X1 U2386 ( .A1(n2356), .A2(n2357), .ZN(n2355) );
  NAND2_X1 U2387 ( .A1(n2358), .A2(n2359), .ZN(n2354) );
  NAND2_X1 U2388 ( .A1(n2360), .A2(n2361), .ZN(n2359) );
  NAND2_X1 U2389 ( .A1(n2362), .A2(n2363), .ZN(n2360) );
  NAND2_X1 U2390 ( .A1(n2350), .A2(n2364), .ZN(Result_8_) );
  NAND2_X1 U2391 ( .A1(n2349), .A2(n2365), .ZN(n2364) );
  XOR2_X1 U2392 ( .A(n2366), .B(n2367), .Z(n2365) );
  NAND2_X1 U2393 ( .A1(n2350), .A2(n2368), .ZN(Result_7_) );
  NAND2_X1 U2394 ( .A1(n2349), .A2(n2369), .ZN(n2368) );
  XOR2_X1 U2395 ( .A(n2370), .B(n2371), .Z(n2369) );
  NAND2_X1 U2396 ( .A1(n2367), .A2(n2366), .ZN(n2371) );
  NAND2_X1 U2397 ( .A1(n2372), .A2(n2373), .ZN(n2370) );
  NAND2_X1 U2398 ( .A1(n2374), .A2(n2375), .ZN(n2373) );
  NAND2_X1 U2399 ( .A1(n2376), .A2(n2377), .ZN(n2374) );
  NAND2_X1 U2400 ( .A1(n2350), .A2(n2378), .ZN(Result_6_) );
  NAND2_X1 U2401 ( .A1(n2349), .A2(n2379), .ZN(n2378) );
  XOR2_X1 U2402 ( .A(n2380), .B(n2381), .Z(n2379) );
  NAND2_X1 U2403 ( .A1(n2350), .A2(n2382), .ZN(Result_5_) );
  NAND2_X1 U2404 ( .A1(n2349), .A2(n2383), .ZN(n2382) );
  XOR2_X1 U2405 ( .A(n2384), .B(n2385), .Z(n2383) );
  NAND2_X1 U2406 ( .A1(n2381), .A2(n2380), .ZN(n2385) );
  NAND2_X1 U2407 ( .A1(n2386), .A2(n2387), .ZN(n2384) );
  NAND2_X1 U2408 ( .A1(n2388), .A2(n2389), .ZN(n2387) );
  NAND2_X1 U2409 ( .A1(n2390), .A2(n2391), .ZN(n2388) );
  NAND2_X1 U2410 ( .A1(n2350), .A2(n2392), .ZN(Result_4_) );
  NAND2_X1 U2411 ( .A1(n2393), .A2(n2349), .ZN(n2392) );
  XOR2_X1 U2412 ( .A(n2394), .B(n2395), .Z(n2393) );
  NAND2_X1 U2413 ( .A1(n2350), .A2(n2396), .ZN(Result_3_) );
  NAND2_X1 U2414 ( .A1(n2349), .A2(n2397), .ZN(n2396) );
  XOR2_X1 U2415 ( .A(n2398), .B(n2399), .Z(n2397) );
  NAND2_X1 U2416 ( .A1(n2395), .A2(n2394), .ZN(n2399) );
  NAND2_X1 U2417 ( .A1(n2400), .A2(n2401), .ZN(n2398) );
  NAND2_X1 U2418 ( .A1(n2402), .A2(n2403), .ZN(n2401) );
  NAND2_X1 U2419 ( .A1(n2404), .A2(n2405), .ZN(n2402) );
  NAND2_X1 U2420 ( .A1(n2406), .A2(n2407), .ZN(Result_31_) );
  NAND2_X1 U2421 ( .A1(n2408), .A2(n2349), .ZN(n2407) );
  NAND2_X1 U2422 ( .A1(n2409), .A2(n2410), .ZN(n2406) );
  INV_X1 U2423 ( .A(n2411), .ZN(n2410) );
  NOR3_X1 U2424 ( .A1(n2347), .A2(n2345), .A3(n2343), .ZN(n2411) );
  NAND2_X1 U2425 ( .A1(n2415), .A2(n2416), .ZN(n2409) );
  NAND3_X1 U2426 ( .A1(n2417), .A2(n2418), .A3(n2419), .ZN(Result_30_) );
  NAND3_X1 U2427 ( .A1(a_14_), .A2(n2420), .A3(n2349), .ZN(n2419) );
  NAND2_X1 U2428 ( .A1(b_14_), .A2(n2421), .ZN(n2418) );
  NAND3_X1 U2429 ( .A1(n2422), .A2(n2423), .A3(n2424), .ZN(n2421) );
  NAND2_X1 U2430 ( .A1(n2349), .A2(n2425), .ZN(n2424) );
  NAND2_X1 U2431 ( .A1(n2416), .A2(n2426), .ZN(n2425) );
  NAND2_X1 U2432 ( .A1(n2427), .A2(n2428), .ZN(n2423) );
  NAND2_X1 U2433 ( .A1(a_14_), .A2(n2429), .ZN(n2422) );
  NAND2_X1 U2434 ( .A1(n2430), .A2(n2431), .ZN(n2417) );
  NAND2_X1 U2435 ( .A1(n2432), .A2(n2433), .ZN(n2430) );
  NAND2_X1 U2436 ( .A1(n2429), .A2(n2428), .ZN(n2433) );
  NAND3_X1 U2437 ( .A1(n2434), .A2(n2435), .A3(n2436), .ZN(n2429) );
  NAND2_X1 U2438 ( .A1(n2345), .A2(n2437), .ZN(n2436) );
  NAND2_X1 U2439 ( .A1(n2343), .A2(n2408), .ZN(n2435) );
  INV_X1 U2440 ( .A(n2438), .ZN(n2408) );
  NAND2_X1 U2441 ( .A1(n2347), .A2(n2420), .ZN(n2434) );
  NAND2_X1 U2442 ( .A1(a_14_), .A2(n2439), .ZN(n2432) );
  NAND2_X1 U2443 ( .A1(n2440), .A2(n2441), .ZN(n2439) );
  NAND2_X1 U2444 ( .A1(n2349), .A2(b_15_), .ZN(n2441) );
  INV_X1 U2445 ( .A(n2427), .ZN(n2440) );
  NAND3_X1 U2446 ( .A1(n2442), .A2(n2443), .A3(n2444), .ZN(n2427) );
  NAND2_X1 U2447 ( .A1(n2345), .A2(n2416), .ZN(n2444) );
  NAND2_X1 U2448 ( .A1(n2343), .A2(n2438), .ZN(n2443) );
  NAND2_X1 U2449 ( .A1(n2347), .A2(n2415), .ZN(n2442) );
  NAND2_X1 U2450 ( .A1(n2350), .A2(n2445), .ZN(Result_2_) );
  NAND2_X1 U2451 ( .A1(n2446), .A2(n2349), .ZN(n2445) );
  XOR2_X1 U2452 ( .A(n2447), .B(n2448), .Z(n2446) );
  NAND3_X1 U2453 ( .A1(n2449), .A2(n2450), .A3(n2451), .ZN(Result_29_) );
  NAND2_X1 U2454 ( .A1(n2452), .A2(n2349), .ZN(n2451) );
  XNOR2_X1 U2455 ( .A(n2453), .B(n2454), .ZN(n2452) );
  XOR2_X1 U2456 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND2_X1 U2457 ( .A1(n2457), .A2(n2458), .ZN(n2450) );
  NAND3_X1 U2458 ( .A1(n2459), .A2(n2460), .A3(n2461), .ZN(n2457) );
  NAND2_X1 U2459 ( .A1(n2345), .A2(n2462), .ZN(n2461) );
  NAND2_X1 U2460 ( .A1(n2343), .A2(n2463), .ZN(n2460) );
  NAND2_X1 U2461 ( .A1(n2347), .A2(n2464), .ZN(n2459) );
  NAND2_X1 U2462 ( .A1(n2465), .A2(n2466), .ZN(n2449) );
  NAND3_X1 U2463 ( .A1(n2467), .A2(n2468), .A3(n2469), .ZN(n2466) );
  NAND2_X1 U2464 ( .A1(n2345), .A2(n2470), .ZN(n2469) );
  NAND2_X1 U2465 ( .A1(n2471), .A2(n2343), .ZN(n2468) );
  INV_X1 U2466 ( .A(n2463), .ZN(n2471) );
  NAND2_X1 U2467 ( .A1(n2347), .A2(n2472), .ZN(n2467) );
  INV_X1 U2468 ( .A(n2458), .ZN(n2465) );
  NAND2_X1 U2469 ( .A1(n2473), .A2(n2474), .ZN(n2458) );
  NAND3_X1 U2470 ( .A1(n2475), .A2(n2476), .A3(n2477), .ZN(Result_28_) );
  NAND2_X1 U2471 ( .A1(n2478), .A2(n2349), .ZN(n2477) );
  XOR2_X1 U2472 ( .A(n2479), .B(n2480), .Z(n2478) );
  XOR2_X1 U2473 ( .A(n2481), .B(n2482), .Z(n2479) );
  NAND2_X1 U2474 ( .A1(n2483), .A2(n2484), .ZN(n2476) );
  NAND3_X1 U2475 ( .A1(n2485), .A2(n2486), .A3(n2487), .ZN(n2483) );
  NAND2_X1 U2476 ( .A1(n2345), .A2(n2488), .ZN(n2487) );
  NAND2_X1 U2477 ( .A1(n2343), .A2(n2489), .ZN(n2486) );
  NAND2_X1 U2478 ( .A1(n2347), .A2(n2490), .ZN(n2485) );
  NAND2_X1 U2479 ( .A1(n2491), .A2(n2492), .ZN(n2475) );
  NAND3_X1 U2480 ( .A1(n2493), .A2(n2494), .A3(n2495), .ZN(n2492) );
  NAND2_X1 U2481 ( .A1(n2345), .A2(n2496), .ZN(n2495) );
  NAND2_X1 U2482 ( .A1(n2497), .A2(n2343), .ZN(n2494) );
  INV_X1 U2483 ( .A(n2489), .ZN(n2497) );
  NAND2_X1 U2484 ( .A1(n2347), .A2(n2498), .ZN(n2493) );
  INV_X1 U2485 ( .A(n2484), .ZN(n2491) );
  NAND2_X1 U2486 ( .A1(n2499), .A2(n2500), .ZN(n2484) );
  NAND3_X1 U2487 ( .A1(n2501), .A2(n2502), .A3(n2503), .ZN(Result_27_) );
  NAND2_X1 U2488 ( .A1(n2504), .A2(n2349), .ZN(n2503) );
  XOR2_X1 U2489 ( .A(n2505), .B(n2506), .Z(n2504) );
  XOR2_X1 U2490 ( .A(n2507), .B(n2508), .Z(n2505) );
  NAND2_X1 U2491 ( .A1(n2509), .A2(n2510), .ZN(n2502) );
  NAND3_X1 U2492 ( .A1(n2511), .A2(n2512), .A3(n2513), .ZN(n2509) );
  NAND2_X1 U2493 ( .A1(n2345), .A2(n2514), .ZN(n2513) );
  NAND2_X1 U2494 ( .A1(n2343), .A2(n2515), .ZN(n2512) );
  NAND2_X1 U2495 ( .A1(n2347), .A2(n2516), .ZN(n2511) );
  NAND2_X1 U2496 ( .A1(n2517), .A2(n2518), .ZN(n2501) );
  NAND3_X1 U2497 ( .A1(n2519), .A2(n2520), .A3(n2521), .ZN(n2518) );
  NAND2_X1 U2498 ( .A1(n2345), .A2(n2522), .ZN(n2521) );
  NAND2_X1 U2499 ( .A1(n2523), .A2(n2343), .ZN(n2520) );
  INV_X1 U2500 ( .A(n2515), .ZN(n2523) );
  NAND2_X1 U2501 ( .A1(n2347), .A2(n2524), .ZN(n2519) );
  INV_X1 U2502 ( .A(n2510), .ZN(n2517) );
  NAND2_X1 U2503 ( .A1(n2525), .A2(n2526), .ZN(n2510) );
  NAND3_X1 U2504 ( .A1(n2527), .A2(n2528), .A3(n2529), .ZN(Result_26_) );
  NAND2_X1 U2505 ( .A1(n2349), .A2(n2530), .ZN(n2529) );
  XNOR2_X1 U2506 ( .A(n2531), .B(n2532), .ZN(n2530) );
  XOR2_X1 U2507 ( .A(n2533), .B(n2534), .Z(n2532) );
  NAND2_X1 U2508 ( .A1(n2535), .A2(n2536), .ZN(n2528) );
  NAND3_X1 U2509 ( .A1(n2537), .A2(n2538), .A3(n2539), .ZN(n2535) );
  NAND2_X1 U2510 ( .A1(n2345), .A2(n2540), .ZN(n2539) );
  NAND2_X1 U2511 ( .A1(n2343), .A2(n2541), .ZN(n2538) );
  NAND2_X1 U2512 ( .A1(n2347), .A2(n2542), .ZN(n2537) );
  NAND2_X1 U2513 ( .A1(n2543), .A2(n2544), .ZN(n2527) );
  NAND3_X1 U2514 ( .A1(n2545), .A2(n2546), .A3(n2547), .ZN(n2544) );
  NAND2_X1 U2515 ( .A1(n2345), .A2(n2548), .ZN(n2547) );
  NAND2_X1 U2516 ( .A1(n2549), .A2(n2343), .ZN(n2546) );
  INV_X1 U2517 ( .A(n2541), .ZN(n2549) );
  NAND2_X1 U2518 ( .A1(n2347), .A2(n2550), .ZN(n2545) );
  INV_X1 U2519 ( .A(n2536), .ZN(n2543) );
  NAND2_X1 U2520 ( .A1(n2551), .A2(n2552), .ZN(n2536) );
  NAND3_X1 U2521 ( .A1(n2553), .A2(n2554), .A3(n2555), .ZN(Result_25_) );
  NAND2_X1 U2522 ( .A1(n2349), .A2(n2556), .ZN(n2555) );
  XNOR2_X1 U2523 ( .A(n2557), .B(n2558), .ZN(n2556) );
  XNOR2_X1 U2524 ( .A(n2559), .B(n2560), .ZN(n2558) );
  NAND2_X1 U2525 ( .A1(n2561), .A2(n2562), .ZN(n2554) );
  NAND3_X1 U2526 ( .A1(n2563), .A2(n2564), .A3(n2565), .ZN(n2562) );
  NAND2_X1 U2527 ( .A1(n2345), .A2(n2566), .ZN(n2565) );
  NAND2_X1 U2528 ( .A1(n2567), .A2(n2343), .ZN(n2564) );
  NAND2_X1 U2529 ( .A1(n2347), .A2(n2568), .ZN(n2563) );
  NAND2_X1 U2530 ( .A1(n2569), .A2(n2570), .ZN(n2553) );
  NAND3_X1 U2531 ( .A1(n2571), .A2(n2572), .A3(n2573), .ZN(n2570) );
  NAND2_X1 U2532 ( .A1(n2345), .A2(n2574), .ZN(n2573) );
  NAND2_X1 U2533 ( .A1(n2343), .A2(n2575), .ZN(n2572) );
  NAND2_X1 U2534 ( .A1(n2347), .A2(n2576), .ZN(n2571) );
  INV_X1 U2535 ( .A(n2561), .ZN(n2569) );
  XNOR2_X1 U2536 ( .A(n2577), .B(b_9_), .ZN(n2561) );
  NAND3_X1 U2537 ( .A1(n2578), .A2(n2579), .A3(n2580), .ZN(Result_24_) );
  NAND2_X1 U2538 ( .A1(n2581), .A2(n2349), .ZN(n2580) );
  XOR2_X1 U2539 ( .A(n2582), .B(n2583), .Z(n2581) );
  XOR2_X1 U2540 ( .A(n2584), .B(n2585), .Z(n2582) );
  NAND2_X1 U2541 ( .A1(n2586), .A2(n2587), .ZN(n2579) );
  NAND3_X1 U2542 ( .A1(n2588), .A2(n2589), .A3(n2590), .ZN(n2586) );
  NAND2_X1 U2543 ( .A1(n2345), .A2(n2591), .ZN(n2590) );
  NAND2_X1 U2544 ( .A1(n2343), .A2(n2592), .ZN(n2589) );
  NAND2_X1 U2545 ( .A1(n2347), .A2(n2593), .ZN(n2588) );
  NAND2_X1 U2546 ( .A1(n2594), .A2(n2595), .ZN(n2578) );
  NAND3_X1 U2547 ( .A1(n2596), .A2(n2597), .A3(n2598), .ZN(n2595) );
  NAND2_X1 U2548 ( .A1(n2345), .A2(n2599), .ZN(n2598) );
  NAND2_X1 U2549 ( .A1(n2600), .A2(n2343), .ZN(n2597) );
  NAND2_X1 U2550 ( .A1(n2347), .A2(n2601), .ZN(n2596) );
  INV_X1 U2551 ( .A(n2587), .ZN(n2594) );
  NAND2_X1 U2552 ( .A1(n2602), .A2(n2603), .ZN(n2587) );
  NAND3_X1 U2553 ( .A1(n2604), .A2(n2605), .A3(n2606), .ZN(Result_23_) );
  NAND2_X1 U2554 ( .A1(n2607), .A2(n2349), .ZN(n2606) );
  XNOR2_X1 U2555 ( .A(n2608), .B(n2609), .ZN(n2607) );
  XOR2_X1 U2556 ( .A(n2610), .B(n2611), .Z(n2609) );
  NAND2_X1 U2557 ( .A1(n2612), .A2(n2613), .ZN(n2605) );
  NAND3_X1 U2558 ( .A1(n2614), .A2(n2615), .A3(n2616), .ZN(n2613) );
  NAND2_X1 U2559 ( .A1(n2345), .A2(n2617), .ZN(n2616) );
  NAND2_X1 U2560 ( .A1(n2618), .A2(n2343), .ZN(n2615) );
  INV_X1 U2561 ( .A(n2619), .ZN(n2618) );
  NAND2_X1 U2562 ( .A1(n2347), .A2(n2620), .ZN(n2614) );
  NAND2_X1 U2563 ( .A1(n2621), .A2(n2622), .ZN(n2604) );
  NAND3_X1 U2564 ( .A1(n2623), .A2(n2624), .A3(n2625), .ZN(n2622) );
  NAND2_X1 U2565 ( .A1(n2345), .A2(n2626), .ZN(n2625) );
  NAND2_X1 U2566 ( .A1(n2343), .A2(n2619), .ZN(n2624) );
  NAND2_X1 U2567 ( .A1(n2347), .A2(n2627), .ZN(n2623) );
  INV_X1 U2568 ( .A(n2612), .ZN(n2621) );
  XNOR2_X1 U2569 ( .A(n2628), .B(b_7_), .ZN(n2612) );
  NAND3_X1 U2570 ( .A1(n2629), .A2(n2630), .A3(n2631), .ZN(Result_22_) );
  NAND2_X1 U2571 ( .A1(n2349), .A2(n2632), .ZN(n2631) );
  XNOR2_X1 U2572 ( .A(n2633), .B(n2634), .ZN(n2632) );
  XNOR2_X1 U2573 ( .A(n2635), .B(n2636), .ZN(n2634) );
  NAND2_X1 U2574 ( .A1(n2637), .A2(n2638), .ZN(n2630) );
  NAND3_X1 U2575 ( .A1(n2639), .A2(n2640), .A3(n2641), .ZN(n2637) );
  NAND2_X1 U2576 ( .A1(n2345), .A2(n2642), .ZN(n2641) );
  NAND2_X1 U2577 ( .A1(n2343), .A2(n2643), .ZN(n2640) );
  NAND2_X1 U2578 ( .A1(n2347), .A2(n2644), .ZN(n2639) );
  NAND2_X1 U2579 ( .A1(n2645), .A2(n2646), .ZN(n2629) );
  NAND3_X1 U2580 ( .A1(n2647), .A2(n2648), .A3(n2649), .ZN(n2646) );
  NAND2_X1 U2581 ( .A1(n2345), .A2(n2650), .ZN(n2649) );
  NAND2_X1 U2582 ( .A1(n2651), .A2(n2343), .ZN(n2648) );
  INV_X1 U2583 ( .A(n2643), .ZN(n2651) );
  NAND2_X1 U2584 ( .A1(n2347), .A2(n2652), .ZN(n2647) );
  INV_X1 U2585 ( .A(n2638), .ZN(n2645) );
  NAND2_X1 U2586 ( .A1(n2653), .A2(n2654), .ZN(n2638) );
  NAND3_X1 U2587 ( .A1(n2655), .A2(n2656), .A3(n2657), .ZN(Result_21_) );
  NAND2_X1 U2588 ( .A1(n2349), .A2(n2658), .ZN(n2657) );
  XNOR2_X1 U2589 ( .A(n2659), .B(n2660), .ZN(n2658) );
  XNOR2_X1 U2590 ( .A(n2661), .B(n2662), .ZN(n2660) );
  NAND2_X1 U2591 ( .A1(n2663), .A2(n2664), .ZN(n2656) );
  NAND3_X1 U2592 ( .A1(n2665), .A2(n2666), .A3(n2667), .ZN(n2664) );
  NAND2_X1 U2593 ( .A1(n2345), .A2(n2668), .ZN(n2667) );
  NAND2_X1 U2594 ( .A1(n2669), .A2(n2343), .ZN(n2666) );
  INV_X1 U2595 ( .A(n2670), .ZN(n2669) );
  NAND2_X1 U2596 ( .A1(n2347), .A2(n2671), .ZN(n2665) );
  NAND2_X1 U2597 ( .A1(n2672), .A2(n2673), .ZN(n2655) );
  NAND3_X1 U2598 ( .A1(n2674), .A2(n2675), .A3(n2676), .ZN(n2673) );
  NAND2_X1 U2599 ( .A1(n2345), .A2(n2677), .ZN(n2676) );
  NAND2_X1 U2600 ( .A1(n2343), .A2(n2670), .ZN(n2675) );
  NAND2_X1 U2601 ( .A1(n2347), .A2(n2678), .ZN(n2674) );
  INV_X1 U2602 ( .A(n2663), .ZN(n2672) );
  XNOR2_X1 U2603 ( .A(n2679), .B(b_5_), .ZN(n2663) );
  NAND3_X1 U2604 ( .A1(n2680), .A2(n2681), .A3(n2682), .ZN(Result_20_) );
  NAND2_X1 U2605 ( .A1(n2349), .A2(n2683), .ZN(n2682) );
  XNOR2_X1 U2606 ( .A(n2684), .B(n2685), .ZN(n2683) );
  XNOR2_X1 U2607 ( .A(n2686), .B(n2687), .ZN(n2685) );
  NAND2_X1 U2608 ( .A1(n2688), .A2(n2689), .ZN(n2681) );
  NAND3_X1 U2609 ( .A1(n2690), .A2(n2691), .A3(n2692), .ZN(n2688) );
  NAND2_X1 U2610 ( .A1(n2345), .A2(n2693), .ZN(n2692) );
  NAND2_X1 U2611 ( .A1(n2343), .A2(n2694), .ZN(n2691) );
  NAND2_X1 U2612 ( .A1(n2347), .A2(n2695), .ZN(n2690) );
  NAND2_X1 U2613 ( .A1(n2696), .A2(n2697), .ZN(n2680) );
  NAND3_X1 U2614 ( .A1(n2698), .A2(n2699), .A3(n2700), .ZN(n2697) );
  NAND2_X1 U2615 ( .A1(n2345), .A2(n2701), .ZN(n2700) );
  NAND2_X1 U2616 ( .A1(n2702), .A2(n2343), .ZN(n2699) );
  INV_X1 U2617 ( .A(n2694), .ZN(n2702) );
  NAND2_X1 U2618 ( .A1(n2347), .A2(n2703), .ZN(n2698) );
  INV_X1 U2619 ( .A(n2689), .ZN(n2696) );
  NAND2_X1 U2620 ( .A1(n2704), .A2(n2705), .ZN(n2689) );
  NAND2_X1 U2621 ( .A1(n2350), .A2(n2706), .ZN(Result_1_) );
  NAND2_X1 U2622 ( .A1(n2349), .A2(n2707), .ZN(n2706) );
  XOR2_X1 U2623 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND2_X1 U2624 ( .A1(n2448), .A2(n2447), .ZN(n2709) );
  NAND2_X1 U2625 ( .A1(n2710), .A2(n2711), .ZN(n2708) );
  NAND3_X1 U2626 ( .A1(n2712), .A2(n2713), .A3(n2714), .ZN(n2711) );
  NAND3_X1 U2627 ( .A1(n2715), .A2(n2716), .A3(n2717), .ZN(Result_19_) );
  NAND2_X1 U2628 ( .A1(n2349), .A2(n2718), .ZN(n2717) );
  XNOR2_X1 U2629 ( .A(n2719), .B(n2720), .ZN(n2718) );
  NAND2_X1 U2630 ( .A1(n2721), .A2(n2722), .ZN(n2719) );
  NAND2_X1 U2631 ( .A1(n2723), .A2(n2724), .ZN(n2716) );
  NAND3_X1 U2632 ( .A1(n2725), .A2(n2726), .A3(n2727), .ZN(n2724) );
  NAND2_X1 U2633 ( .A1(n2345), .A2(n2728), .ZN(n2727) );
  NAND2_X1 U2634 ( .A1(n2729), .A2(n2343), .ZN(n2726) );
  INV_X1 U2635 ( .A(n2730), .ZN(n2729) );
  NAND2_X1 U2636 ( .A1(n2347), .A2(n2731), .ZN(n2725) );
  NAND2_X1 U2637 ( .A1(n2732), .A2(n2733), .ZN(n2715) );
  NAND3_X1 U2638 ( .A1(n2734), .A2(n2735), .A3(n2736), .ZN(n2733) );
  NAND2_X1 U2639 ( .A1(n2345), .A2(n2737), .ZN(n2736) );
  NAND2_X1 U2640 ( .A1(n2343), .A2(n2730), .ZN(n2735) );
  NAND2_X1 U2641 ( .A1(n2347), .A2(n2738), .ZN(n2734) );
  INV_X1 U2642 ( .A(n2723), .ZN(n2732) );
  XNOR2_X1 U2643 ( .A(n2739), .B(b_3_), .ZN(n2723) );
  NAND3_X1 U2644 ( .A1(n2740), .A2(n2741), .A3(n2742), .ZN(Result_18_) );
  NAND2_X1 U2645 ( .A1(n2743), .A2(n2349), .ZN(n2742) );
  XNOR2_X1 U2646 ( .A(n2744), .B(n2745), .ZN(n2743) );
  XOR2_X1 U2647 ( .A(n2746), .B(n2747), .Z(n2745) );
  NAND2_X1 U2648 ( .A1(a_2_), .A2(b_15_), .ZN(n2747) );
  NAND2_X1 U2649 ( .A1(n2748), .A2(n2749), .ZN(n2741) );
  NAND3_X1 U2650 ( .A1(n2750), .A2(n2751), .A3(n2752), .ZN(n2748) );
  NAND2_X1 U2651 ( .A1(n2345), .A2(n2753), .ZN(n2752) );
  NAND2_X1 U2652 ( .A1(n2343), .A2(n2754), .ZN(n2751) );
  NAND2_X1 U2653 ( .A1(n2347), .A2(n2755), .ZN(n2750) );
  NAND2_X1 U2654 ( .A1(n2756), .A2(n2757), .ZN(n2740) );
  NAND3_X1 U2655 ( .A1(n2758), .A2(n2759), .A3(n2760), .ZN(n2757) );
  NAND2_X1 U2656 ( .A1(n2345), .A2(n2761), .ZN(n2760) );
  NAND2_X1 U2657 ( .A1(n2762), .A2(n2343), .ZN(n2759) );
  INV_X1 U2658 ( .A(n2754), .ZN(n2762) );
  NAND2_X1 U2659 ( .A1(n2347), .A2(n2763), .ZN(n2758) );
  INV_X1 U2660 ( .A(n2749), .ZN(n2756) );
  NAND2_X1 U2661 ( .A1(n2764), .A2(n2765), .ZN(n2749) );
  NAND3_X1 U2662 ( .A1(n2766), .A2(n2767), .A3(n2768), .ZN(Result_17_) );
  NAND2_X1 U2663 ( .A1(n2769), .A2(n2349), .ZN(n2768) );
  XNOR2_X1 U2664 ( .A(n2770), .B(n2771), .ZN(n2769) );
  XOR2_X1 U2665 ( .A(n2772), .B(n2773), .Z(n2771) );
  NAND2_X1 U2666 ( .A1(a_1_), .A2(b_15_), .ZN(n2773) );
  NAND2_X1 U2667 ( .A1(n2774), .A2(n2775), .ZN(n2767) );
  NAND3_X1 U2668 ( .A1(n2776), .A2(n2777), .A3(n2778), .ZN(n2775) );
  NAND2_X1 U2669 ( .A1(n2345), .A2(n2779), .ZN(n2778) );
  NAND2_X1 U2670 ( .A1(n2780), .A2(n2343), .ZN(n2777) );
  NAND2_X1 U2671 ( .A1(n2347), .A2(n2781), .ZN(n2776) );
  NAND2_X1 U2672 ( .A1(n2782), .A2(n2783), .ZN(n2766) );
  NAND3_X1 U2673 ( .A1(n2784), .A2(n2785), .A3(n2786), .ZN(n2783) );
  NAND2_X1 U2674 ( .A1(n2345), .A2(n2787), .ZN(n2786) );
  NAND2_X1 U2675 ( .A1(n2343), .A2(n2788), .ZN(n2785) );
  NAND2_X1 U2676 ( .A1(n2347), .A2(n2789), .ZN(n2784) );
  INV_X1 U2677 ( .A(n2774), .ZN(n2782) );
  XNOR2_X1 U2678 ( .A(n2790), .B(b_1_), .ZN(n2774) );
  NAND3_X1 U2679 ( .A1(n2791), .A2(n2792), .A3(n2793), .ZN(Result_16_) );
  NAND2_X1 U2680 ( .A1(n2349), .A2(n2794), .ZN(n2793) );
  XNOR2_X1 U2681 ( .A(n2795), .B(n2796), .ZN(n2794) );
  XOR2_X1 U2682 ( .A(n2797), .B(n2798), .Z(n2796) );
  NAND2_X1 U2683 ( .A1(a_0_), .A2(b_15_), .ZN(n2798) );
  NAND2_X1 U2684 ( .A1(n2799), .A2(n2800), .ZN(n2792) );
  NAND3_X1 U2685 ( .A1(n2801), .A2(n2802), .A3(n2803), .ZN(n2799) );
  NAND2_X1 U2686 ( .A1(n2345), .A2(n2804), .ZN(n2803) );
  NAND2_X1 U2687 ( .A1(n2805), .A2(n2343), .ZN(n2802) );
  INV_X1 U2688 ( .A(n2806), .ZN(n2805) );
  NAND2_X1 U2689 ( .A1(n2347), .A2(n2807), .ZN(n2801) );
  NAND2_X1 U2690 ( .A1(n2808), .A2(n2809), .ZN(n2791) );
  NAND3_X1 U2691 ( .A1(n2810), .A2(n2811), .A3(n2812), .ZN(n2809) );
  NAND2_X1 U2692 ( .A1(n2345), .A2(n2813), .ZN(n2812) );
  NAND2_X1 U2693 ( .A1(n2343), .A2(n2806), .ZN(n2811) );
  NAND2_X1 U2694 ( .A1(n2814), .A2(n2815), .ZN(n2806) );
  NAND2_X1 U2695 ( .A1(n2780), .A2(n2816), .ZN(n2815) );
  INV_X1 U2696 ( .A(n2788), .ZN(n2780) );
  NAND2_X1 U2697 ( .A1(n2764), .A2(n2817), .ZN(n2788) );
  NAND2_X1 U2698 ( .A1(n2765), .A2(n2754), .ZN(n2817) );
  NAND2_X1 U2699 ( .A1(n2818), .A2(n2819), .ZN(n2754) );
  NAND2_X1 U2700 ( .A1(n2820), .A2(n2730), .ZN(n2819) );
  NAND2_X1 U2701 ( .A1(n2704), .A2(n2821), .ZN(n2730) );
  NAND2_X1 U2702 ( .A1(n2705), .A2(n2694), .ZN(n2821) );
  NAND2_X1 U2703 ( .A1(n2822), .A2(n2823), .ZN(n2694) );
  NAND2_X1 U2704 ( .A1(n2824), .A2(n2670), .ZN(n2823) );
  NAND2_X1 U2705 ( .A1(n2653), .A2(n2825), .ZN(n2670) );
  NAND2_X1 U2706 ( .A1(n2654), .A2(n2643), .ZN(n2825) );
  NAND2_X1 U2707 ( .A1(n2826), .A2(n2827), .ZN(n2643) );
  NAND2_X1 U2708 ( .A1(n2828), .A2(n2619), .ZN(n2827) );
  NAND2_X1 U2709 ( .A1(n2602), .A2(n2829), .ZN(n2619) );
  NAND2_X1 U2710 ( .A1(n2603), .A2(n2592), .ZN(n2829) );
  INV_X1 U2711 ( .A(n2600), .ZN(n2592) );
  NOR2_X1 U2712 ( .A1(n2830), .A2(n2831), .ZN(n2600) );
  NOR2_X1 U2713 ( .A1(n2832), .A2(n2567), .ZN(n2831) );
  INV_X1 U2714 ( .A(n2575), .ZN(n2567) );
  NAND2_X1 U2715 ( .A1(n2551), .A2(n2833), .ZN(n2575) );
  NAND2_X1 U2716 ( .A1(n2552), .A2(n2541), .ZN(n2833) );
  NAND2_X1 U2717 ( .A1(n2525), .A2(n2834), .ZN(n2541) );
  NAND2_X1 U2718 ( .A1(n2526), .A2(n2515), .ZN(n2834) );
  NAND2_X1 U2719 ( .A1(n2499), .A2(n2835), .ZN(n2515) );
  NAND2_X1 U2720 ( .A1(n2500), .A2(n2489), .ZN(n2835) );
  NAND2_X1 U2721 ( .A1(n2473), .A2(n2836), .ZN(n2489) );
  NAND2_X1 U2722 ( .A1(n2474), .A2(n2463), .ZN(n2836) );
  NAND2_X1 U2723 ( .A1(n2837), .A2(n2838), .ZN(n2463) );
  NAND2_X1 U2724 ( .A1(b_14_), .A2(n2839), .ZN(n2838) );
  NAND2_X1 U2725 ( .A1(n2428), .A2(n2438), .ZN(n2839) );
  NAND2_X1 U2726 ( .A1(a_15_), .A2(b_15_), .ZN(n2438) );
  NAND2_X1 U2727 ( .A1(n2840), .A2(b_15_), .ZN(n2837) );
  NAND2_X1 U2728 ( .A1(n2841), .A2(n2842), .ZN(n2474) );
  NAND2_X1 U2729 ( .A1(n2843), .A2(n2844), .ZN(n2500) );
  NAND2_X1 U2730 ( .A1(n2845), .A2(n2846), .ZN(n2526) );
  INV_X1 U2731 ( .A(n2847), .ZN(n2525) );
  NAND2_X1 U2732 ( .A1(n2848), .A2(n2849), .ZN(n2552) );
  NOR2_X1 U2733 ( .A1(b_9_), .A2(a_9_), .ZN(n2832) );
  NAND2_X1 U2734 ( .A1(n2850), .A2(n2851), .ZN(n2603) );
  NAND2_X1 U2735 ( .A1(n2852), .A2(n2628), .ZN(n2828) );
  NAND2_X1 U2736 ( .A1(n2853), .A2(n2854), .ZN(n2654) );
  NAND2_X1 U2737 ( .A1(n2855), .A2(n2679), .ZN(n2824) );
  NAND2_X1 U2738 ( .A1(n2856), .A2(n2857), .ZN(n2705) );
  NAND2_X1 U2739 ( .A1(n2858), .A2(n2739), .ZN(n2820) );
  NAND2_X1 U2740 ( .A1(n2859), .A2(n2860), .ZN(n2765) );
  NAND2_X1 U2741 ( .A1(n2861), .A2(n2790), .ZN(n2814) );
  NOR2_X1 U2742 ( .A1(operation_0_), .A2(operation_1_), .ZN(n2414) );
  NAND2_X1 U2743 ( .A1(n2347), .A2(n2862), .ZN(n2810) );
  INV_X1 U2744 ( .A(n2800), .ZN(n2808) );
  NAND2_X1 U2745 ( .A1(n2863), .A2(n2864), .ZN(n2800) );
  NAND2_X1 U2746 ( .A1(n2865), .A2(n2866), .ZN(n2864) );
  NAND2_X1 U2747 ( .A1(n2350), .A2(n2867), .ZN(Result_15_) );
  NAND2_X1 U2748 ( .A1(n2868), .A2(n2349), .ZN(n2867) );
  XOR2_X1 U2749 ( .A(n2869), .B(n2870), .Z(n2868) );
  NAND2_X1 U2750 ( .A1(n2350), .A2(n2871), .ZN(Result_14_) );
  NAND3_X1 U2751 ( .A1(n2872), .A2(n2873), .A3(n2349), .ZN(n2871) );
  NAND2_X1 U2752 ( .A1(n2874), .A2(n2875), .ZN(n2872) );
  NAND2_X1 U2753 ( .A1(n2870), .A2(n2869), .ZN(n2875) );
  XNOR2_X1 U2754 ( .A(n2876), .B(n2877), .ZN(n2874) );
  NAND2_X1 U2755 ( .A1(n2350), .A2(n2878), .ZN(Result_13_) );
  NAND2_X1 U2756 ( .A1(n2349), .A2(n2879), .ZN(n2878) );
  XOR2_X1 U2757 ( .A(n2873), .B(n2880), .Z(n2879) );
  NAND2_X1 U2758 ( .A1(n2881), .A2(n2882), .ZN(n2880) );
  NAND2_X1 U2759 ( .A1(n2883), .A2(n2884), .ZN(n2882) );
  INV_X1 U2760 ( .A(n2885), .ZN(n2883) );
  NOR2_X1 U2761 ( .A1(n2877), .A2(n2876), .ZN(n2885) );
  NAND2_X1 U2762 ( .A1(n2350), .A2(n2886), .ZN(Result_12_) );
  NAND2_X1 U2763 ( .A1(n2887), .A2(n2349), .ZN(n2886) );
  XOR2_X1 U2764 ( .A(n2888), .B(n2889), .Z(n2887) );
  NAND2_X1 U2765 ( .A1(n2350), .A2(n2890), .ZN(Result_11_) );
  NAND2_X1 U2766 ( .A1(n2349), .A2(n2891), .ZN(n2890) );
  XNOR2_X1 U2767 ( .A(n2892), .B(n2893), .ZN(n2891) );
  NAND2_X1 U2768 ( .A1(n2889), .A2(n2888), .ZN(n2893) );
  NOR2_X1 U2769 ( .A1(n2894), .A2(n2895), .ZN(n2892) );
  INV_X1 U2770 ( .A(n2896), .ZN(n2895) );
  NOR2_X1 U2771 ( .A1(n2897), .A2(n2898), .ZN(n2894) );
  INV_X1 U2772 ( .A(n2899), .ZN(n2897) );
  NAND2_X1 U2773 ( .A1(n2900), .A2(n2901), .ZN(n2899) );
  NAND2_X1 U2774 ( .A1(n2350), .A2(n2902), .ZN(Result_10_) );
  NAND2_X1 U2775 ( .A1(n2903), .A2(n2349), .ZN(n2902) );
  XOR2_X1 U2776 ( .A(n2357), .B(n2356), .Z(n2903) );
  NAND2_X1 U2777 ( .A1(n2350), .A2(n2904), .ZN(Result_0_) );
  NAND2_X1 U2778 ( .A1(n2349), .A2(n2905), .ZN(n2904) );
  NAND2_X1 U2779 ( .A1(n2906), .A2(n2907), .ZN(n2905) );
  NAND3_X1 U2780 ( .A1(n2710), .A2(n2447), .A3(n2448), .ZN(n2907) );
  XOR2_X1 U2781 ( .A(n2908), .B(n2909), .Z(n2448) );
  NAND3_X1 U2782 ( .A1(n2910), .A2(n2400), .A3(n2911), .ZN(n2447) );
  NAND3_X1 U2783 ( .A1(n2395), .A2(n2394), .A3(n2912), .ZN(n2911) );
  NAND3_X1 U2784 ( .A1(n2913), .A2(n2386), .A3(n2914), .ZN(n2394) );
  NAND3_X1 U2785 ( .A1(n2381), .A2(n2380), .A3(n2915), .ZN(n2914) );
  NAND3_X1 U2786 ( .A1(n2916), .A2(n2372), .A3(n2917), .ZN(n2380) );
  NAND3_X1 U2787 ( .A1(n2367), .A2(n2366), .A3(n2918), .ZN(n2917) );
  NAND3_X1 U2788 ( .A1(n2919), .A2(n2358), .A3(n2920), .ZN(n2366) );
  NAND3_X1 U2789 ( .A1(n2356), .A2(n2357), .A3(n2921), .ZN(n2920) );
  NAND3_X1 U2790 ( .A1(n2922), .A2(n2896), .A3(n2923), .ZN(n2357) );
  NAND2_X1 U2791 ( .A1(n2924), .A2(n2925), .ZN(n2923) );
  NAND3_X1 U2792 ( .A1(n2898), .A2(n2900), .A3(n2901), .ZN(n2896) );
  NAND3_X1 U2793 ( .A1(n2898), .A2(n2889), .A3(n2888), .ZN(n2922) );
  XOR2_X1 U2794 ( .A(n2900), .B(n2901), .Z(n2888) );
  XNOR2_X1 U2795 ( .A(n2926), .B(n2927), .ZN(n2901) );
  XNOR2_X1 U2796 ( .A(n2928), .B(n2929), .ZN(n2927) );
  NAND2_X1 U2797 ( .A1(n2930), .A2(n2931), .ZN(n2900) );
  NAND3_X1 U2798 ( .A1(a_0_), .A2(n2932), .A3(b_12_), .ZN(n2931) );
  INV_X1 U2799 ( .A(n2933), .ZN(n2932) );
  NOR2_X1 U2800 ( .A1(n2934), .A2(n2935), .ZN(n2933) );
  NAND2_X1 U2801 ( .A1(n2935), .A2(n2934), .ZN(n2930) );
  NAND3_X1 U2802 ( .A1(n2936), .A2(n2881), .A3(n2937), .ZN(n2889) );
  INV_X1 U2803 ( .A(n2938), .ZN(n2937) );
  NOR2_X1 U2804 ( .A1(n2873), .A2(n2884), .ZN(n2938) );
  NAND3_X1 U2805 ( .A1(n2939), .A2(n2869), .A3(n2870), .ZN(n2873) );
  XNOR2_X1 U2806 ( .A(n2940), .B(n2941), .ZN(n2870) );
  XOR2_X1 U2807 ( .A(n2942), .B(n2943), .Z(n2941) );
  NAND2_X1 U2808 ( .A1(b_14_), .A2(a_0_), .ZN(n2943) );
  NAND2_X1 U2809 ( .A1(n2944), .A2(n2945), .ZN(n2869) );
  NAND3_X1 U2810 ( .A1(b_15_), .A2(n2946), .A3(a_0_), .ZN(n2945) );
  INV_X1 U2811 ( .A(n2947), .ZN(n2946) );
  NOR2_X1 U2812 ( .A1(n2797), .A2(n2795), .ZN(n2947) );
  NAND2_X1 U2813 ( .A1(n2795), .A2(n2797), .ZN(n2944) );
  NAND2_X1 U2814 ( .A1(n2948), .A2(n2949), .ZN(n2797) );
  INV_X1 U2815 ( .A(n2950), .ZN(n2949) );
  NOR3_X1 U2816 ( .A1(n2951), .A2(n2952), .A3(n2790), .ZN(n2950) );
  NOR2_X1 U2817 ( .A1(n2772), .A2(n2770), .ZN(n2952) );
  NAND2_X1 U2818 ( .A1(n2770), .A2(n2772), .ZN(n2948) );
  NAND2_X1 U2819 ( .A1(n2953), .A2(n2954), .ZN(n2772) );
  INV_X1 U2820 ( .A(n2955), .ZN(n2954) );
  NOR3_X1 U2821 ( .A1(n2951), .A2(n2956), .A3(n2860), .ZN(n2955) );
  NOR2_X1 U2822 ( .A1(n2746), .A2(n2744), .ZN(n2956) );
  NAND2_X1 U2823 ( .A1(n2744), .A2(n2746), .ZN(n2953) );
  NAND2_X1 U2824 ( .A1(n2721), .A2(n2957), .ZN(n2746) );
  NAND2_X1 U2825 ( .A1(n2720), .A2(n2722), .ZN(n2957) );
  NAND2_X1 U2826 ( .A1(n2958), .A2(n2959), .ZN(n2722) );
  NAND2_X1 U2827 ( .A1(a_3_), .A2(b_15_), .ZN(n2959) );
  XNOR2_X1 U2828 ( .A(n2960), .B(n2961), .ZN(n2720) );
  XNOR2_X1 U2829 ( .A(n2962), .B(n2963), .ZN(n2960) );
  NOR2_X1 U2830 ( .A1(n2857), .A2(n2431), .ZN(n2963) );
  INV_X1 U2831 ( .A(n2964), .ZN(n2721) );
  NOR2_X1 U2832 ( .A1(n2739), .A2(n2958), .ZN(n2964) );
  NOR2_X1 U2833 ( .A1(n2965), .A2(n2966), .ZN(n2958) );
  INV_X1 U2834 ( .A(n2967), .ZN(n2966) );
  NAND2_X1 U2835 ( .A1(n2684), .A2(n2968), .ZN(n2967) );
  NAND2_X1 U2836 ( .A1(n2686), .A2(n2687), .ZN(n2968) );
  XNOR2_X1 U2837 ( .A(n2969), .B(n2970), .ZN(n2684) );
  XOR2_X1 U2838 ( .A(n2971), .B(n2972), .Z(n2970) );
  NAND2_X1 U2839 ( .A1(b_14_), .A2(a_5_), .ZN(n2972) );
  NOR2_X1 U2840 ( .A1(n2687), .A2(n2686), .ZN(n2965) );
  NOR2_X1 U2841 ( .A1(n2973), .A2(n2974), .ZN(n2686) );
  INV_X1 U2842 ( .A(n2975), .ZN(n2974) );
  NAND2_X1 U2843 ( .A1(n2659), .A2(n2976), .ZN(n2975) );
  NAND2_X1 U2844 ( .A1(n2661), .A2(n2662), .ZN(n2976) );
  XOR2_X1 U2845 ( .A(n2977), .B(n2978), .Z(n2659) );
  XOR2_X1 U2846 ( .A(n2979), .B(n2980), .Z(n2977) );
  NOR2_X1 U2847 ( .A1(n2854), .A2(n2431), .ZN(n2980) );
  NOR2_X1 U2848 ( .A1(n2662), .A2(n2661), .ZN(n2973) );
  NOR2_X1 U2849 ( .A1(n2981), .A2(n2982), .ZN(n2661) );
  INV_X1 U2850 ( .A(n2983), .ZN(n2982) );
  NAND2_X1 U2851 ( .A1(n2633), .A2(n2984), .ZN(n2983) );
  NAND2_X1 U2852 ( .A1(n2635), .A2(n2636), .ZN(n2984) );
  XOR2_X1 U2853 ( .A(n2985), .B(n2986), .Z(n2633) );
  XNOR2_X1 U2854 ( .A(n2987), .B(n2988), .ZN(n2986) );
  NAND2_X1 U2855 ( .A1(b_14_), .A2(a_7_), .ZN(n2988) );
  NOR2_X1 U2856 ( .A1(n2636), .A2(n2635), .ZN(n2981) );
  NOR2_X1 U2857 ( .A1(n2989), .A2(n2990), .ZN(n2635) );
  INV_X1 U2858 ( .A(n2991), .ZN(n2990) );
  NAND2_X1 U2859 ( .A1(n2608), .A2(n2992), .ZN(n2991) );
  NAND2_X1 U2860 ( .A1(n2993), .A2(n2611), .ZN(n2992) );
  XNOR2_X1 U2861 ( .A(n2994), .B(n2995), .ZN(n2608) );
  XNOR2_X1 U2862 ( .A(n2996), .B(n2997), .ZN(n2994) );
  NOR2_X1 U2863 ( .A1(n2851), .A2(n2431), .ZN(n2997) );
  NOR2_X1 U2864 ( .A1(n2611), .A2(n2993), .ZN(n2989) );
  INV_X1 U2865 ( .A(n2610), .ZN(n2993) );
  NAND2_X1 U2866 ( .A1(n2998), .A2(n2999), .ZN(n2610) );
  NAND2_X1 U2867 ( .A1(n2583), .A2(n3000), .ZN(n2999) );
  INV_X1 U2868 ( .A(n3001), .ZN(n3000) );
  NOR2_X1 U2869 ( .A1(n2584), .A2(n2585), .ZN(n3001) );
  XOR2_X1 U2870 ( .A(n3002), .B(n3003), .Z(n2583) );
  XOR2_X1 U2871 ( .A(n3004), .B(n3005), .Z(n3002) );
  NOR2_X1 U2872 ( .A1(n2577), .A2(n2431), .ZN(n3005) );
  NAND2_X1 U2873 ( .A1(n2585), .A2(n2584), .ZN(n2998) );
  NAND2_X1 U2874 ( .A1(n3006), .A2(n3007), .ZN(n2584) );
  NAND2_X1 U2875 ( .A1(n2557), .A2(n3008), .ZN(n3007) );
  NAND2_X1 U2876 ( .A1(n2559), .A2(n2560), .ZN(n3008) );
  XNOR2_X1 U2877 ( .A(n3009), .B(n3010), .ZN(n2557) );
  NAND2_X1 U2878 ( .A1(n3011), .A2(n3012), .ZN(n3009) );
  INV_X1 U2879 ( .A(n3013), .ZN(n3006) );
  NOR2_X1 U2880 ( .A1(n2560), .A2(n2559), .ZN(n3013) );
  NOR2_X1 U2881 ( .A1(n3014), .A2(n3015), .ZN(n2559) );
  INV_X1 U2882 ( .A(n3016), .ZN(n3015) );
  NAND2_X1 U2883 ( .A1(n2531), .A2(n3017), .ZN(n3016) );
  NAND2_X1 U2884 ( .A1(n3018), .A2(n2534), .ZN(n3017) );
  XNOR2_X1 U2885 ( .A(n3019), .B(n3020), .ZN(n2531) );
  NAND2_X1 U2886 ( .A1(n3021), .A2(n3022), .ZN(n3019) );
  NOR2_X1 U2887 ( .A1(n2534), .A2(n3018), .ZN(n3014) );
  INV_X1 U2888 ( .A(n2533), .ZN(n3018) );
  NAND2_X1 U2889 ( .A1(n3023), .A2(n3024), .ZN(n2533) );
  NAND2_X1 U2890 ( .A1(n2506), .A2(n3025), .ZN(n3024) );
  INV_X1 U2891 ( .A(n3026), .ZN(n3025) );
  NOR2_X1 U2892 ( .A1(n2507), .A2(n2508), .ZN(n3026) );
  XNOR2_X1 U2893 ( .A(n3027), .B(n3028), .ZN(n2506) );
  XNOR2_X1 U2894 ( .A(n3029), .B(n3030), .ZN(n3027) );
  NAND2_X1 U2895 ( .A1(n2508), .A2(n2507), .ZN(n3023) );
  NAND2_X1 U2896 ( .A1(n3031), .A2(n3032), .ZN(n2507) );
  NAND2_X1 U2897 ( .A1(n2482), .A2(n3033), .ZN(n3032) );
  NAND2_X1 U2898 ( .A1(n2480), .A2(n2481), .ZN(n3033) );
  NOR2_X1 U2899 ( .A1(n2844), .A2(n2951), .ZN(n2482) );
  INV_X1 U2900 ( .A(n3034), .ZN(n3031) );
  NOR2_X1 U2901 ( .A1(n2481), .A2(n2480), .ZN(n3034) );
  XOR2_X1 U2902 ( .A(n3035), .B(n3036), .Z(n2480) );
  XOR2_X1 U2903 ( .A(n3037), .B(n3038), .Z(n3036) );
  NAND2_X1 U2904 ( .A1(n3039), .A2(n3040), .ZN(n2481) );
  NAND2_X1 U2905 ( .A1(n3041), .A2(n2455), .ZN(n3040) );
  NAND2_X1 U2906 ( .A1(a_13_), .A2(b_15_), .ZN(n2455) );
  NAND2_X1 U2907 ( .A1(n2453), .A2(n2456), .ZN(n3041) );
  INV_X1 U2908 ( .A(n3042), .ZN(n3039) );
  NOR2_X1 U2909 ( .A1(n2456), .A2(n2453), .ZN(n3042) );
  NOR3_X1 U2910 ( .A1(n2431), .A2(n2951), .A3(n3043), .ZN(n2453) );
  NAND2_X1 U2911 ( .A1(n3044), .A2(n3045), .ZN(n2456) );
  NAND2_X1 U2912 ( .A1(b_13_), .A2(n3046), .ZN(n3045) );
  NAND2_X1 U2913 ( .A1(n2426), .A2(n3047), .ZN(n3046) );
  NAND2_X1 U2914 ( .A1(a_15_), .A2(n2431), .ZN(n3047) );
  NAND2_X1 U2915 ( .A1(b_14_), .A2(n3048), .ZN(n3044) );
  NAND2_X1 U2916 ( .A1(n3049), .A2(n3050), .ZN(n3048) );
  NAND2_X1 U2917 ( .A1(a_14_), .A2(n2841), .ZN(n3050) );
  NOR2_X1 U2918 ( .A1(n2846), .A2(n2951), .ZN(n2508) );
  NAND2_X1 U2919 ( .A1(a_10_), .A2(b_15_), .ZN(n2534) );
  NAND2_X1 U2920 ( .A1(a_9_), .A2(b_15_), .ZN(n2560) );
  NOR2_X1 U2921 ( .A1(n2851), .A2(n2951), .ZN(n2585) );
  NAND2_X1 U2922 ( .A1(a_7_), .A2(b_15_), .ZN(n2611) );
  NAND2_X1 U2923 ( .A1(a_6_), .A2(b_15_), .ZN(n2636) );
  NAND2_X1 U2924 ( .A1(a_5_), .A2(b_15_), .ZN(n2662) );
  NAND2_X1 U2925 ( .A1(a_4_), .A2(b_15_), .ZN(n2687) );
  XNOR2_X1 U2926 ( .A(n3051), .B(n3052), .ZN(n2744) );
  XNOR2_X1 U2927 ( .A(n3053), .B(n3054), .ZN(n3051) );
  NOR2_X1 U2928 ( .A1(n2739), .A2(n2431), .ZN(n3054) );
  XNOR2_X1 U2929 ( .A(n3055), .B(n3056), .ZN(n2770) );
  XNOR2_X1 U2930 ( .A(n3057), .B(n3058), .ZN(n3055) );
  NOR2_X1 U2931 ( .A1(n2860), .A2(n2431), .ZN(n3058) );
  XOR2_X1 U2932 ( .A(n3059), .B(n3060), .Z(n2795) );
  XNOR2_X1 U2933 ( .A(n3061), .B(n3062), .ZN(n3060) );
  NAND2_X1 U2934 ( .A1(b_14_), .A2(a_1_), .ZN(n3062) );
  XOR2_X1 U2935 ( .A(n2876), .B(n2877), .Z(n2939) );
  INV_X1 U2936 ( .A(n3063), .ZN(n2881) );
  NOR3_X1 U2937 ( .A1(n2877), .A2(n2876), .A3(n2884), .ZN(n3063) );
  NAND2_X1 U2938 ( .A1(n3064), .A2(n2936), .ZN(n2884) );
  NAND2_X1 U2939 ( .A1(n3065), .A2(n3066), .ZN(n3064) );
  INV_X1 U2940 ( .A(n3067), .ZN(n3066) );
  XOR2_X1 U2941 ( .A(n3068), .B(n2935), .Z(n3065) );
  NOR2_X1 U2942 ( .A1(n3069), .A2(n3070), .ZN(n2876) );
  NOR3_X1 U2943 ( .A1(n2865), .A2(n3071), .A3(n2431), .ZN(n3070) );
  NOR2_X1 U2944 ( .A1(n2942), .A2(n2940), .ZN(n3071) );
  INV_X1 U2945 ( .A(n3072), .ZN(n3069) );
  NAND2_X1 U2946 ( .A1(n2940), .A2(n2942), .ZN(n3072) );
  NAND2_X1 U2947 ( .A1(n3073), .A2(n3074), .ZN(n2942) );
  NAND3_X1 U2948 ( .A1(a_1_), .A2(n3075), .A3(b_14_), .ZN(n3074) );
  NAND2_X1 U2949 ( .A1(n3061), .A2(n3059), .ZN(n3075) );
  INV_X1 U2950 ( .A(n3076), .ZN(n3073) );
  NOR2_X1 U2951 ( .A1(n3059), .A2(n3061), .ZN(n3076) );
  NOR2_X1 U2952 ( .A1(n3077), .A2(n3078), .ZN(n3061) );
  NOR3_X1 U2953 ( .A1(n2860), .A2(n3079), .A3(n2431), .ZN(n3078) );
  INV_X1 U2954 ( .A(n3080), .ZN(n3079) );
  NAND2_X1 U2955 ( .A1(n3057), .A2(n3056), .ZN(n3080) );
  NOR2_X1 U2956 ( .A1(n3056), .A2(n3057), .ZN(n3077) );
  NOR2_X1 U2957 ( .A1(n3081), .A2(n3082), .ZN(n3057) );
  NOR3_X1 U2958 ( .A1(n2739), .A2(n3083), .A3(n2431), .ZN(n3082) );
  INV_X1 U2959 ( .A(n3084), .ZN(n3083) );
  NAND2_X1 U2960 ( .A1(n3053), .A2(n3052), .ZN(n3084) );
  NOR2_X1 U2961 ( .A1(n3052), .A2(n3053), .ZN(n3081) );
  NOR2_X1 U2962 ( .A1(n3085), .A2(n3086), .ZN(n3053) );
  INV_X1 U2963 ( .A(n3087), .ZN(n3086) );
  NAND3_X1 U2964 ( .A1(a_4_), .A2(n3088), .A3(b_14_), .ZN(n3087) );
  NAND2_X1 U2965 ( .A1(n2962), .A2(n2961), .ZN(n3088) );
  NOR2_X1 U2966 ( .A1(n2961), .A2(n2962), .ZN(n3085) );
  NOR2_X1 U2967 ( .A1(n3089), .A2(n3090), .ZN(n2962) );
  NOR3_X1 U2968 ( .A1(n2679), .A2(n3091), .A3(n2431), .ZN(n3090) );
  NOR2_X1 U2969 ( .A1(n2971), .A2(n2969), .ZN(n3091) );
  INV_X1 U2970 ( .A(n3092), .ZN(n3089) );
  NAND2_X1 U2971 ( .A1(n2969), .A2(n2971), .ZN(n3092) );
  NAND2_X1 U2972 ( .A1(n3093), .A2(n3094), .ZN(n2971) );
  NAND3_X1 U2973 ( .A1(a_6_), .A2(n3095), .A3(b_14_), .ZN(n3094) );
  INV_X1 U2974 ( .A(n3096), .ZN(n3095) );
  NOR2_X1 U2975 ( .A1(n2979), .A2(n2978), .ZN(n3096) );
  NAND2_X1 U2976 ( .A1(n2978), .A2(n2979), .ZN(n3093) );
  NAND2_X1 U2977 ( .A1(n3097), .A2(n3098), .ZN(n2979) );
  NAND3_X1 U2978 ( .A1(a_7_), .A2(n3099), .A3(b_14_), .ZN(n3098) );
  NAND2_X1 U2979 ( .A1(n2987), .A2(n2985), .ZN(n3099) );
  INV_X1 U2980 ( .A(n3100), .ZN(n3097) );
  NOR2_X1 U2981 ( .A1(n2985), .A2(n2987), .ZN(n3100) );
  NOR2_X1 U2982 ( .A1(n3101), .A2(n3102), .ZN(n2987) );
  NOR3_X1 U2983 ( .A1(n2851), .A2(n3103), .A3(n2431), .ZN(n3102) );
  INV_X1 U2984 ( .A(n3104), .ZN(n3103) );
  NAND2_X1 U2985 ( .A1(n2996), .A2(n2995), .ZN(n3104) );
  NOR2_X1 U2986 ( .A1(n2995), .A2(n2996), .ZN(n3101) );
  NOR2_X1 U2987 ( .A1(n3105), .A2(n3106), .ZN(n2996) );
  NOR3_X1 U2988 ( .A1(n2577), .A2(n3107), .A3(n2431), .ZN(n3106) );
  NOR2_X1 U2989 ( .A1(n3004), .A2(n3003), .ZN(n3107) );
  INV_X1 U2990 ( .A(n3108), .ZN(n3105) );
  NAND2_X1 U2991 ( .A1(n3003), .A2(n3004), .ZN(n3108) );
  NAND2_X1 U2992 ( .A1(n3011), .A2(n3109), .ZN(n3004) );
  NAND2_X1 U2993 ( .A1(n3010), .A2(n3012), .ZN(n3109) );
  NAND2_X1 U2994 ( .A1(n3110), .A2(n3111), .ZN(n3012) );
  NAND2_X1 U2995 ( .A1(b_14_), .A2(a_10_), .ZN(n3111) );
  INV_X1 U2996 ( .A(n3112), .ZN(n3110) );
  XOR2_X1 U2997 ( .A(n3113), .B(n3114), .Z(n3010) );
  XOR2_X1 U2998 ( .A(n3115), .B(n3116), .Z(n3113) );
  NAND2_X1 U2999 ( .A1(a_10_), .A2(n3112), .ZN(n3011) );
  NAND2_X1 U3000 ( .A1(n3021), .A2(n3117), .ZN(n3112) );
  NAND2_X1 U3001 ( .A1(n3020), .A2(n3022), .ZN(n3117) );
  NAND2_X1 U3002 ( .A1(n3118), .A2(n3119), .ZN(n3022) );
  NAND2_X1 U3003 ( .A1(b_14_), .A2(a_11_), .ZN(n3119) );
  XNOR2_X1 U3004 ( .A(n3120), .B(n3121), .ZN(n3020) );
  XNOR2_X1 U3005 ( .A(n3122), .B(n3123), .ZN(n3121) );
  INV_X1 U3006 ( .A(n3124), .ZN(n3021) );
  NOR2_X1 U3007 ( .A1(n2846), .A2(n3118), .ZN(n3124) );
  NOR2_X1 U3008 ( .A1(n3125), .A2(n3126), .ZN(n3118) );
  INV_X1 U3009 ( .A(n3127), .ZN(n3126) );
  NAND2_X1 U3010 ( .A1(n3029), .A2(n3128), .ZN(n3127) );
  NAND2_X1 U3011 ( .A1(n3030), .A2(n3028), .ZN(n3128) );
  NOR2_X1 U3012 ( .A1(n2431), .A2(n2844), .ZN(n3029) );
  NOR2_X1 U3013 ( .A1(n3028), .A2(n3030), .ZN(n3125) );
  NOR2_X1 U3014 ( .A1(n3129), .A2(n3130), .ZN(n3030) );
  INV_X1 U3015 ( .A(n3131), .ZN(n3130) );
  NAND2_X1 U3016 ( .A1(n3035), .A2(n3132), .ZN(n3131) );
  NAND2_X1 U3017 ( .A1(n3133), .A2(n3037), .ZN(n3132) );
  NOR2_X1 U3018 ( .A1(n2431), .A2(n2842), .ZN(n3035) );
  NOR2_X1 U3019 ( .A1(n3037), .A2(n3133), .ZN(n3129) );
  INV_X1 U3020 ( .A(n3038), .ZN(n3133) );
  NAND2_X1 U3021 ( .A1(n3134), .A2(n3135), .ZN(n3038) );
  NAND2_X1 U3022 ( .A1(b_12_), .A2(n3136), .ZN(n3135) );
  NAND2_X1 U3023 ( .A1(n2426), .A2(n3137), .ZN(n3136) );
  NAND2_X1 U3024 ( .A1(a_15_), .A2(n2841), .ZN(n3137) );
  NAND2_X1 U3025 ( .A1(b_13_), .A2(n3138), .ZN(n3134) );
  NAND2_X1 U3026 ( .A1(n3049), .A2(n3139), .ZN(n3138) );
  NAND2_X1 U3027 ( .A1(a_14_), .A2(n2843), .ZN(n3139) );
  NAND3_X1 U3028 ( .A1(b_13_), .A2(b_14_), .A3(n2840), .ZN(n3037) );
  XNOR2_X1 U3029 ( .A(n2473), .B(n3140), .ZN(n3028) );
  XOR2_X1 U3030 ( .A(n3141), .B(n3142), .Z(n3140) );
  XNOR2_X1 U3031 ( .A(n3143), .B(n3144), .ZN(n3003) );
  NAND2_X1 U3032 ( .A1(n3145), .A2(n3146), .ZN(n3143) );
  XNOR2_X1 U3033 ( .A(n3147), .B(n3148), .ZN(n2995) );
  XNOR2_X1 U3034 ( .A(n3149), .B(n3150), .ZN(n3148) );
  XOR2_X1 U3035 ( .A(n3151), .B(n3152), .Z(n2985) );
  XNOR2_X1 U3036 ( .A(n3153), .B(n3154), .ZN(n3152) );
  XOR2_X1 U3037 ( .A(n3155), .B(n3156), .Z(n2978) );
  XNOR2_X1 U3038 ( .A(n3157), .B(n3158), .ZN(n3156) );
  NAND2_X1 U3039 ( .A1(b_13_), .A2(a_7_), .ZN(n3158) );
  XOR2_X1 U3040 ( .A(n3159), .B(n3160), .Z(n2969) );
  XNOR2_X1 U3041 ( .A(n3161), .B(n3162), .ZN(n3160) );
  NAND2_X1 U3042 ( .A1(b_13_), .A2(a_6_), .ZN(n3162) );
  XOR2_X1 U3043 ( .A(n3163), .B(n3164), .Z(n2961) );
  XOR2_X1 U3044 ( .A(n3165), .B(n3166), .Z(n3164) );
  NAND2_X1 U3045 ( .A1(b_13_), .A2(a_5_), .ZN(n3166) );
  XOR2_X1 U3046 ( .A(n3167), .B(n3168), .Z(n3052) );
  XOR2_X1 U3047 ( .A(n3169), .B(n3170), .Z(n3168) );
  NAND2_X1 U3048 ( .A1(b_13_), .A2(a_4_), .ZN(n3170) );
  XNOR2_X1 U3049 ( .A(n3171), .B(n3172), .ZN(n3056) );
  XOR2_X1 U3050 ( .A(n3173), .B(n3174), .Z(n3171) );
  NOR2_X1 U3051 ( .A1(n2739), .A2(n2841), .ZN(n3174) );
  XOR2_X1 U3052 ( .A(n3175), .B(n3176), .Z(n3059) );
  XNOR2_X1 U3053 ( .A(n3177), .B(n3178), .ZN(n3176) );
  XOR2_X1 U3054 ( .A(n3179), .B(n3180), .Z(n2940) );
  XOR2_X1 U3055 ( .A(n3181), .B(n3182), .Z(n3179) );
  NOR2_X1 U3056 ( .A1(n2790), .A2(n2841), .ZN(n3182) );
  XOR2_X1 U3057 ( .A(n3183), .B(n3184), .Z(n2877) );
  NAND2_X1 U3058 ( .A1(n3185), .A2(n3186), .ZN(n3183) );
  NAND2_X1 U3059 ( .A1(n3187), .A2(n3067), .ZN(n2936) );
  NAND2_X1 U3060 ( .A1(n3185), .A2(n3188), .ZN(n3067) );
  NAND2_X1 U3061 ( .A1(n3184), .A2(n3186), .ZN(n3188) );
  NAND2_X1 U3062 ( .A1(n3189), .A2(n3190), .ZN(n3186) );
  NAND2_X1 U3063 ( .A1(b_13_), .A2(a_0_), .ZN(n3190) );
  XNOR2_X1 U3064 ( .A(n3191), .B(n3192), .ZN(n3184) );
  XNOR2_X1 U3065 ( .A(n3193), .B(n3194), .ZN(n3192) );
  NAND2_X1 U3066 ( .A1(a_0_), .A2(n3195), .ZN(n3185) );
  INV_X1 U3067 ( .A(n3189), .ZN(n3195) );
  NOR2_X1 U3068 ( .A1(n3196), .A2(n3197), .ZN(n3189) );
  NOR3_X1 U3069 ( .A1(n2790), .A2(n3198), .A3(n2841), .ZN(n3197) );
  NOR2_X1 U3070 ( .A1(n3181), .A2(n3180), .ZN(n3198) );
  INV_X1 U3071 ( .A(n3199), .ZN(n3196) );
  NAND2_X1 U3072 ( .A1(n3180), .A2(n3181), .ZN(n3199) );
  NAND2_X1 U3073 ( .A1(n3200), .A2(n3201), .ZN(n3181) );
  NAND2_X1 U3074 ( .A1(n3178), .A2(n3202), .ZN(n3201) );
  INV_X1 U3075 ( .A(n3203), .ZN(n3202) );
  NOR2_X1 U3076 ( .A1(n3177), .A2(n3175), .ZN(n3203) );
  NOR2_X1 U3077 ( .A1(n2841), .A2(n2860), .ZN(n3178) );
  NAND2_X1 U3078 ( .A1(n3175), .A2(n3177), .ZN(n3200) );
  NAND2_X1 U3079 ( .A1(n3204), .A2(n3205), .ZN(n3177) );
  INV_X1 U3080 ( .A(n3206), .ZN(n3205) );
  NOR3_X1 U3081 ( .A1(n2739), .A2(n3207), .A3(n2841), .ZN(n3206) );
  NOR2_X1 U3082 ( .A1(n3173), .A2(n3172), .ZN(n3207) );
  NAND2_X1 U3083 ( .A1(n3172), .A2(n3173), .ZN(n3204) );
  NAND2_X1 U3084 ( .A1(n3208), .A2(n3209), .ZN(n3173) );
  NAND3_X1 U3085 ( .A1(a_4_), .A2(n3210), .A3(b_13_), .ZN(n3209) );
  INV_X1 U3086 ( .A(n3211), .ZN(n3210) );
  NOR2_X1 U3087 ( .A1(n3169), .A2(n3167), .ZN(n3211) );
  NAND2_X1 U3088 ( .A1(n3167), .A2(n3169), .ZN(n3208) );
  NAND2_X1 U3089 ( .A1(n3212), .A2(n3213), .ZN(n3169) );
  INV_X1 U3090 ( .A(n3214), .ZN(n3213) );
  NOR3_X1 U3091 ( .A1(n2679), .A2(n3215), .A3(n2841), .ZN(n3214) );
  NOR2_X1 U3092 ( .A1(n3165), .A2(n3163), .ZN(n3215) );
  NAND2_X1 U3093 ( .A1(n3163), .A2(n3165), .ZN(n3212) );
  NAND2_X1 U3094 ( .A1(n3216), .A2(n3217), .ZN(n3165) );
  NAND3_X1 U3095 ( .A1(a_6_), .A2(n3218), .A3(b_13_), .ZN(n3217) );
  NAND2_X1 U3096 ( .A1(n3161), .A2(n3159), .ZN(n3218) );
  INV_X1 U3097 ( .A(n3219), .ZN(n3216) );
  NOR2_X1 U3098 ( .A1(n3159), .A2(n3161), .ZN(n3219) );
  NOR2_X1 U3099 ( .A1(n3220), .A2(n3221), .ZN(n3161) );
  NOR3_X1 U3100 ( .A1(n2628), .A2(n3222), .A3(n2841), .ZN(n3221) );
  INV_X1 U3101 ( .A(n3223), .ZN(n3222) );
  NAND2_X1 U3102 ( .A1(n3157), .A2(n3155), .ZN(n3223) );
  NOR2_X1 U3103 ( .A1(n3155), .A2(n3157), .ZN(n3220) );
  NOR2_X1 U3104 ( .A1(n3224), .A2(n3225), .ZN(n3157) );
  INV_X1 U3105 ( .A(n3226), .ZN(n3225) );
  NAND2_X1 U3106 ( .A1(n3154), .A2(n3227), .ZN(n3226) );
  NAND2_X1 U3107 ( .A1(n3151), .A2(n3153), .ZN(n3227) );
  NOR2_X1 U3108 ( .A1(n2841), .A2(n2851), .ZN(n3154) );
  NOR2_X1 U3109 ( .A1(n3153), .A2(n3151), .ZN(n3224) );
  XNOR2_X1 U3110 ( .A(n3228), .B(n3229), .ZN(n3151) );
  XOR2_X1 U3111 ( .A(n3230), .B(n3231), .Z(n3228) );
  NOR2_X1 U3112 ( .A1(n2577), .A2(n2843), .ZN(n3231) );
  NAND2_X1 U3113 ( .A1(n3232), .A2(n3233), .ZN(n3153) );
  NAND2_X1 U3114 ( .A1(n3147), .A2(n3234), .ZN(n3233) );
  NAND2_X1 U3115 ( .A1(n3150), .A2(n3149), .ZN(n3234) );
  XNOR2_X1 U3116 ( .A(n3235), .B(n3236), .ZN(n3147) );
  XNOR2_X1 U3117 ( .A(n3237), .B(n3238), .ZN(n3236) );
  INV_X1 U3118 ( .A(n3239), .ZN(n3232) );
  NOR2_X1 U3119 ( .A1(n3149), .A2(n3150), .ZN(n3239) );
  NOR2_X1 U3120 ( .A1(n2841), .A2(n2577), .ZN(n3150) );
  NAND2_X1 U3121 ( .A1(n3145), .A2(n3240), .ZN(n3149) );
  NAND2_X1 U3122 ( .A1(n3144), .A2(n3146), .ZN(n3240) );
  NAND2_X1 U3123 ( .A1(n3241), .A2(n3242), .ZN(n3146) );
  NAND2_X1 U3124 ( .A1(b_13_), .A2(a_10_), .ZN(n3242) );
  INV_X1 U3125 ( .A(n3243), .ZN(n3241) );
  XNOR2_X1 U3126 ( .A(n3244), .B(n3245), .ZN(n3144) );
  XNOR2_X1 U3127 ( .A(n3246), .B(n3247), .ZN(n3244) );
  NAND2_X1 U3128 ( .A1(a_10_), .A2(n3243), .ZN(n3145) );
  NAND2_X1 U3129 ( .A1(n3248), .A2(n3249), .ZN(n3243) );
  NAND2_X1 U3130 ( .A1(n3116), .A2(n3250), .ZN(n3249) );
  INV_X1 U3131 ( .A(n3251), .ZN(n3250) );
  NOR2_X1 U3132 ( .A1(n3115), .A2(n3114), .ZN(n3251) );
  NOR2_X1 U3133 ( .A1(n2841), .A2(n2846), .ZN(n3116) );
  NAND2_X1 U3134 ( .A1(n3114), .A2(n3115), .ZN(n3248) );
  NAND2_X1 U3135 ( .A1(n3252), .A2(n3253), .ZN(n3115) );
  NAND2_X1 U3136 ( .A1(n3123), .A2(n3254), .ZN(n3253) );
  NAND2_X1 U3137 ( .A1(n3120), .A2(n3122), .ZN(n3254) );
  NOR2_X1 U3138 ( .A1(n2841), .A2(n2844), .ZN(n3123) );
  INV_X1 U3139 ( .A(n3255), .ZN(n3252) );
  NOR2_X1 U3140 ( .A1(n3122), .A2(n3120), .ZN(n3255) );
  XOR2_X1 U3141 ( .A(n3256), .B(n3257), .Z(n3120) );
  XOR2_X1 U3142 ( .A(n3258), .B(n3259), .Z(n3257) );
  NAND2_X1 U3143 ( .A1(n3260), .A2(n3261), .ZN(n3122) );
  NAND2_X1 U3144 ( .A1(n3262), .A2(n3141), .ZN(n3261) );
  NAND3_X1 U3145 ( .A1(b_12_), .A2(b_13_), .A3(n2840), .ZN(n3141) );
  NAND2_X1 U3146 ( .A1(n3263), .A2(n3142), .ZN(n3262) );
  INV_X1 U3147 ( .A(n2473), .ZN(n3263) );
  NAND2_X1 U3148 ( .A1(n3264), .A2(n2473), .ZN(n3260) );
  NAND2_X1 U3149 ( .A1(b_13_), .A2(a_13_), .ZN(n2473) );
  INV_X1 U3150 ( .A(n3142), .ZN(n3264) );
  NAND2_X1 U3151 ( .A1(n3265), .A2(n3266), .ZN(n3142) );
  NAND2_X1 U3152 ( .A1(b_11_), .A2(n3267), .ZN(n3266) );
  NAND2_X1 U3153 ( .A1(n2426), .A2(n3268), .ZN(n3267) );
  NAND2_X1 U3154 ( .A1(a_15_), .A2(n2843), .ZN(n3268) );
  NAND2_X1 U3155 ( .A1(b_12_), .A2(n3269), .ZN(n3265) );
  NAND2_X1 U3156 ( .A1(n3049), .A2(n3270), .ZN(n3269) );
  NAND2_X1 U3157 ( .A1(a_14_), .A2(n2845), .ZN(n3270) );
  XNOR2_X1 U3158 ( .A(n3271), .B(n3272), .ZN(n3114) );
  XOR2_X1 U3159 ( .A(n2499), .B(n3273), .Z(n3271) );
  XOR2_X1 U3160 ( .A(n3274), .B(n3275), .Z(n3155) );
  XNOR2_X1 U3161 ( .A(n3276), .B(n3277), .ZN(n3274) );
  NOR2_X1 U3162 ( .A1(n2851), .A2(n2843), .ZN(n3277) );
  XOR2_X1 U3163 ( .A(n3278), .B(n3279), .Z(n3159) );
  XNOR2_X1 U3164 ( .A(n3280), .B(n3281), .ZN(n3278) );
  NOR2_X1 U3165 ( .A1(n2628), .A2(n2843), .ZN(n3281) );
  XNOR2_X1 U3166 ( .A(n3282), .B(n3283), .ZN(n3163) );
  XNOR2_X1 U3167 ( .A(n3284), .B(n3285), .ZN(n3282) );
  NOR2_X1 U3168 ( .A1(n2854), .A2(n2843), .ZN(n3285) );
  XOR2_X1 U3169 ( .A(n3286), .B(n3287), .Z(n3167) );
  XNOR2_X1 U3170 ( .A(n3288), .B(n3289), .ZN(n3287) );
  NAND2_X1 U3171 ( .A1(b_12_), .A2(a_5_), .ZN(n3289) );
  XNOR2_X1 U3172 ( .A(n3290), .B(n3291), .ZN(n3172) );
  XOR2_X1 U3173 ( .A(n3292), .B(n3293), .Z(n3291) );
  NAND2_X1 U3174 ( .A1(b_12_), .A2(a_4_), .ZN(n3293) );
  XOR2_X1 U3175 ( .A(n3294), .B(n3295), .Z(n3175) );
  XNOR2_X1 U3176 ( .A(n3296), .B(n3297), .ZN(n3295) );
  NAND2_X1 U3177 ( .A1(b_12_), .A2(a_3_), .ZN(n3297) );
  XOR2_X1 U3178 ( .A(n3298), .B(n3299), .Z(n3180) );
  XNOR2_X1 U3179 ( .A(n3300), .B(n3301), .ZN(n3299) );
  NAND2_X1 U3180 ( .A1(b_12_), .A2(a_2_), .ZN(n3301) );
  XOR2_X1 U3181 ( .A(n3302), .B(n3068), .Z(n3187) );
  XNOR2_X1 U3182 ( .A(n2934), .B(n3303), .ZN(n3068) );
  NOR2_X1 U3183 ( .A1(n2865), .A2(n2843), .ZN(n3303) );
  NAND2_X1 U3184 ( .A1(n3304), .A2(n3305), .ZN(n2934) );
  NAND2_X1 U3185 ( .A1(n3194), .A2(n3306), .ZN(n3305) );
  INV_X1 U3186 ( .A(n3307), .ZN(n3306) );
  NOR2_X1 U3187 ( .A1(n3193), .A2(n3191), .ZN(n3307) );
  NOR2_X1 U3188 ( .A1(n2843), .A2(n2790), .ZN(n3194) );
  NAND2_X1 U3189 ( .A1(n3191), .A2(n3193), .ZN(n3304) );
  NAND2_X1 U3190 ( .A1(n3308), .A2(n3309), .ZN(n3193) );
  NAND3_X1 U3191 ( .A1(a_2_), .A2(n3310), .A3(b_12_), .ZN(n3309) );
  NAND2_X1 U3192 ( .A1(n3300), .A2(n3298), .ZN(n3310) );
  INV_X1 U3193 ( .A(n3311), .ZN(n3308) );
  NOR2_X1 U3194 ( .A1(n3298), .A2(n3300), .ZN(n3311) );
  NOR2_X1 U3195 ( .A1(n3312), .A2(n3313), .ZN(n3300) );
  NOR3_X1 U3196 ( .A1(n2739), .A2(n3314), .A3(n2843), .ZN(n3313) );
  INV_X1 U3197 ( .A(n3315), .ZN(n3314) );
  NAND2_X1 U3198 ( .A1(n3296), .A2(n3294), .ZN(n3315) );
  NOR2_X1 U3199 ( .A1(n3294), .A2(n3296), .ZN(n3312) );
  NOR2_X1 U3200 ( .A1(n3316), .A2(n3317), .ZN(n3296) );
  NOR3_X1 U3201 ( .A1(n2857), .A2(n3318), .A3(n2843), .ZN(n3317) );
  NOR2_X1 U3202 ( .A1(n3292), .A2(n3290), .ZN(n3318) );
  INV_X1 U3203 ( .A(n3319), .ZN(n3316) );
  NAND2_X1 U3204 ( .A1(n3290), .A2(n3292), .ZN(n3319) );
  NAND2_X1 U3205 ( .A1(n3320), .A2(n3321), .ZN(n3292) );
  NAND3_X1 U3206 ( .A1(a_5_), .A2(n3322), .A3(b_12_), .ZN(n3321) );
  NAND2_X1 U3207 ( .A1(n3288), .A2(n3286), .ZN(n3322) );
  INV_X1 U3208 ( .A(n3323), .ZN(n3320) );
  NOR2_X1 U3209 ( .A1(n3286), .A2(n3288), .ZN(n3323) );
  NOR2_X1 U3210 ( .A1(n3324), .A2(n3325), .ZN(n3288) );
  INV_X1 U3211 ( .A(n3326), .ZN(n3325) );
  NAND3_X1 U3212 ( .A1(a_6_), .A2(n3327), .A3(b_12_), .ZN(n3326) );
  NAND2_X1 U3213 ( .A1(n3284), .A2(n3283), .ZN(n3327) );
  NOR2_X1 U3214 ( .A1(n3283), .A2(n3284), .ZN(n3324) );
  NOR2_X1 U3215 ( .A1(n3328), .A2(n3329), .ZN(n3284) );
  INV_X1 U3216 ( .A(n3330), .ZN(n3329) );
  NAND3_X1 U3217 ( .A1(a_7_), .A2(n3331), .A3(b_12_), .ZN(n3330) );
  NAND2_X1 U3218 ( .A1(n3280), .A2(n3279), .ZN(n3331) );
  NOR2_X1 U3219 ( .A1(n3279), .A2(n3280), .ZN(n3328) );
  NOR2_X1 U3220 ( .A1(n3332), .A2(n3333), .ZN(n3280) );
  NOR3_X1 U3221 ( .A1(n2851), .A2(n3334), .A3(n2843), .ZN(n3333) );
  INV_X1 U3222 ( .A(n3335), .ZN(n3334) );
  NAND2_X1 U3223 ( .A1(n3276), .A2(n3275), .ZN(n3335) );
  NOR2_X1 U3224 ( .A1(n3275), .A2(n3276), .ZN(n3332) );
  NOR2_X1 U3225 ( .A1(n3336), .A2(n3337), .ZN(n3276) );
  NOR3_X1 U3226 ( .A1(n2577), .A2(n3338), .A3(n2843), .ZN(n3337) );
  INV_X1 U3227 ( .A(n3339), .ZN(n3338) );
  NAND2_X1 U3228 ( .A1(n3229), .A2(n3230), .ZN(n3339) );
  NOR2_X1 U3229 ( .A1(n3230), .A2(n3229), .ZN(n3336) );
  XOR2_X1 U3230 ( .A(n3340), .B(n3341), .Z(n3229) );
  NAND2_X1 U3231 ( .A1(n3342), .A2(n3343), .ZN(n3340) );
  NAND2_X1 U3232 ( .A1(n3344), .A2(n3345), .ZN(n3230) );
  NAND2_X1 U3233 ( .A1(n3235), .A2(n3346), .ZN(n3345) );
  INV_X1 U3234 ( .A(n3347), .ZN(n3346) );
  NOR2_X1 U3235 ( .A1(n3238), .A2(n3237), .ZN(n3347) );
  XOR2_X1 U3236 ( .A(n3348), .B(n3349), .Z(n3235) );
  XOR2_X1 U3237 ( .A(n3350), .B(n2847), .Z(n3348) );
  NAND2_X1 U3238 ( .A1(n3237), .A2(n3238), .ZN(n3344) );
  NAND2_X1 U3239 ( .A1(b_12_), .A2(a_10_), .ZN(n3238) );
  NOR2_X1 U3240 ( .A1(n3351), .A2(n3352), .ZN(n3237) );
  INV_X1 U3241 ( .A(n3353), .ZN(n3352) );
  NAND2_X1 U3242 ( .A1(n3246), .A2(n3354), .ZN(n3353) );
  NAND2_X1 U3243 ( .A1(n3247), .A2(n3245), .ZN(n3354) );
  NOR2_X1 U3244 ( .A1(n2843), .A2(n2846), .ZN(n3246) );
  NOR2_X1 U3245 ( .A1(n3245), .A2(n3247), .ZN(n3351) );
  NOR2_X1 U3246 ( .A1(n3355), .A2(n3356), .ZN(n3247) );
  NOR2_X1 U3247 ( .A1(n2499), .A2(n3357), .ZN(n3356) );
  INV_X1 U3248 ( .A(n3358), .ZN(n3357) );
  NAND2_X1 U3249 ( .A1(n3273), .A2(n3272), .ZN(n3358) );
  NAND2_X1 U3250 ( .A1(b_12_), .A2(a_12_), .ZN(n2499) );
  NOR2_X1 U3251 ( .A1(n3272), .A2(n3273), .ZN(n3355) );
  NOR2_X1 U3252 ( .A1(n3359), .A2(n3360), .ZN(n3273) );
  INV_X1 U3253 ( .A(n3361), .ZN(n3360) );
  NAND2_X1 U3254 ( .A1(n3256), .A2(n3362), .ZN(n3361) );
  NAND2_X1 U3255 ( .A1(n3363), .A2(n3258), .ZN(n3362) );
  NOR2_X1 U3256 ( .A1(n2843), .A2(n2842), .ZN(n3256) );
  NOR2_X1 U3257 ( .A1(n3258), .A2(n3363), .ZN(n3359) );
  INV_X1 U3258 ( .A(n3259), .ZN(n3363) );
  NAND2_X1 U3259 ( .A1(n3364), .A2(n3365), .ZN(n3259) );
  NAND2_X1 U3260 ( .A1(b_10_), .A2(n3366), .ZN(n3365) );
  NAND2_X1 U3261 ( .A1(n2426), .A2(n3367), .ZN(n3366) );
  NAND2_X1 U3262 ( .A1(a_15_), .A2(n2845), .ZN(n3367) );
  NAND2_X1 U3263 ( .A1(b_11_), .A2(n3368), .ZN(n3364) );
  NAND2_X1 U3264 ( .A1(n3049), .A2(n3369), .ZN(n3368) );
  NAND2_X1 U3265 ( .A1(a_14_), .A2(n2848), .ZN(n3369) );
  NAND3_X1 U3266 ( .A1(b_11_), .A2(b_12_), .A3(n2840), .ZN(n3258) );
  XNOR2_X1 U3267 ( .A(n3370), .B(n3371), .ZN(n3272) );
  XOR2_X1 U3268 ( .A(n3372), .B(n3373), .Z(n3370) );
  XNOR2_X1 U3269 ( .A(n3374), .B(n3375), .ZN(n3245) );
  XOR2_X1 U3270 ( .A(n3376), .B(n3377), .Z(n3374) );
  XOR2_X1 U3271 ( .A(n3378), .B(n3379), .Z(n3275) );
  XOR2_X1 U3272 ( .A(n3380), .B(n3381), .Z(n3379) );
  NAND2_X1 U3273 ( .A1(b_11_), .A2(a_9_), .ZN(n3381) );
  XOR2_X1 U3274 ( .A(n3382), .B(n3383), .Z(n3279) );
  XOR2_X1 U3275 ( .A(n3384), .B(n3385), .Z(n3383) );
  NAND2_X1 U3276 ( .A1(b_11_), .A2(a_8_), .ZN(n3385) );
  XNOR2_X1 U3277 ( .A(n3386), .B(n3387), .ZN(n3283) );
  XOR2_X1 U3278 ( .A(n3388), .B(n3389), .Z(n3386) );
  NOR2_X1 U3279 ( .A1(n2628), .A2(n2845), .ZN(n3389) );
  XOR2_X1 U3280 ( .A(n3390), .B(n3391), .Z(n3286) );
  XOR2_X1 U3281 ( .A(n3392), .B(n3393), .Z(n3391) );
  NAND2_X1 U3282 ( .A1(b_11_), .A2(a_6_), .ZN(n3393) );
  XNOR2_X1 U3283 ( .A(n3394), .B(n3395), .ZN(n3290) );
  XOR2_X1 U3284 ( .A(n3396), .B(n3397), .Z(n3395) );
  NAND2_X1 U3285 ( .A1(b_11_), .A2(a_5_), .ZN(n3397) );
  XOR2_X1 U3286 ( .A(n3398), .B(n3399), .Z(n3294) );
  XNOR2_X1 U3287 ( .A(n3400), .B(n3401), .ZN(n3398) );
  XOR2_X1 U3288 ( .A(n3402), .B(n3403), .Z(n3298) );
  XOR2_X1 U3289 ( .A(n3404), .B(n3405), .Z(n3402) );
  XOR2_X1 U3290 ( .A(n3406), .B(n3407), .Z(n3191) );
  XOR2_X1 U3291 ( .A(n3408), .B(n3409), .Z(n3406) );
  NOR2_X1 U3292 ( .A1(n2860), .A2(n2845), .ZN(n3409) );
  INV_X1 U3293 ( .A(n2935), .ZN(n3302) );
  XOR2_X1 U3294 ( .A(n3410), .B(n3411), .Z(n2935) );
  XNOR2_X1 U3295 ( .A(n3412), .B(n3413), .ZN(n3411) );
  XOR2_X1 U3296 ( .A(n2925), .B(n2924), .Z(n2898) );
  XNOR2_X1 U3297 ( .A(n3414), .B(n3415), .ZN(n2924) );
  NAND2_X1 U3298 ( .A1(n3416), .A2(n3417), .ZN(n3414) );
  NAND2_X1 U3299 ( .A1(n3418), .A2(n3419), .ZN(n2925) );
  NAND2_X1 U3300 ( .A1(n2929), .A2(n3420), .ZN(n3419) );
  NAND2_X1 U3301 ( .A1(n2926), .A2(n2928), .ZN(n3420) );
  NOR2_X1 U3302 ( .A1(n2845), .A2(n2865), .ZN(n2929) );
  INV_X1 U3303 ( .A(n3421), .ZN(n3418) );
  NOR2_X1 U3304 ( .A1(n2928), .A2(n2926), .ZN(n3421) );
  XNOR2_X1 U3305 ( .A(n3422), .B(n3423), .ZN(n2926) );
  XNOR2_X1 U3306 ( .A(n3424), .B(n3425), .ZN(n3423) );
  NAND2_X1 U3307 ( .A1(b_10_), .A2(a_1_), .ZN(n3425) );
  NAND2_X1 U3308 ( .A1(n3426), .A2(n3427), .ZN(n2928) );
  NAND2_X1 U3309 ( .A1(n3410), .A2(n3428), .ZN(n3427) );
  INV_X1 U3310 ( .A(n3429), .ZN(n3428) );
  NOR2_X1 U3311 ( .A1(n3413), .A2(n3412), .ZN(n3429) );
  XOR2_X1 U3312 ( .A(n3430), .B(n3431), .Z(n3410) );
  XNOR2_X1 U3313 ( .A(n3432), .B(n3433), .ZN(n3430) );
  NAND2_X1 U3314 ( .A1(n3412), .A2(n3413), .ZN(n3426) );
  NAND2_X1 U3315 ( .A1(b_11_), .A2(a_1_), .ZN(n3413) );
  NOR2_X1 U3316 ( .A1(n3434), .A2(n3435), .ZN(n3412) );
  NOR3_X1 U3317 ( .A1(n2860), .A2(n3436), .A3(n2845), .ZN(n3435) );
  NOR2_X1 U3318 ( .A1(n3408), .A2(n3407), .ZN(n3436) );
  INV_X1 U3319 ( .A(n3437), .ZN(n3434) );
  NAND2_X1 U3320 ( .A1(n3407), .A2(n3408), .ZN(n3437) );
  NAND2_X1 U3321 ( .A1(n3438), .A2(n3439), .ZN(n3408) );
  NAND2_X1 U3322 ( .A1(n3405), .A2(n3440), .ZN(n3439) );
  NAND2_X1 U3323 ( .A1(n3403), .A2(n3441), .ZN(n3440) );
  INV_X1 U3324 ( .A(n3404), .ZN(n3441) );
  NOR2_X1 U3325 ( .A1(n2845), .A2(n2739), .ZN(n3405) );
  NAND2_X1 U3326 ( .A1(n3442), .A2(n3404), .ZN(n3438) );
  NAND2_X1 U3327 ( .A1(n3443), .A2(n3444), .ZN(n3404) );
  NAND2_X1 U3328 ( .A1(n3401), .A2(n3445), .ZN(n3444) );
  NAND2_X1 U3329 ( .A1(n3400), .A2(n3399), .ZN(n3445) );
  NOR2_X1 U3330 ( .A1(n2845), .A2(n2857), .ZN(n3401) );
  INV_X1 U3331 ( .A(n3446), .ZN(n3443) );
  NOR2_X1 U3332 ( .A1(n3399), .A2(n3400), .ZN(n3446) );
  NOR2_X1 U3333 ( .A1(n3447), .A2(n3448), .ZN(n3400) );
  NOR3_X1 U3334 ( .A1(n2679), .A2(n3449), .A3(n2845), .ZN(n3448) );
  NOR2_X1 U3335 ( .A1(n3394), .A2(n3396), .ZN(n3449) );
  INV_X1 U3336 ( .A(n3450), .ZN(n3447) );
  NAND2_X1 U3337 ( .A1(n3394), .A2(n3396), .ZN(n3450) );
  NAND2_X1 U3338 ( .A1(n3451), .A2(n3452), .ZN(n3396) );
  NAND3_X1 U3339 ( .A1(a_6_), .A2(n3453), .A3(b_11_), .ZN(n3452) );
  INV_X1 U3340 ( .A(n3454), .ZN(n3453) );
  NOR2_X1 U3341 ( .A1(n3390), .A2(n3392), .ZN(n3454) );
  NAND2_X1 U3342 ( .A1(n3390), .A2(n3392), .ZN(n3451) );
  NAND2_X1 U3343 ( .A1(n3455), .A2(n3456), .ZN(n3392) );
  INV_X1 U3344 ( .A(n3457), .ZN(n3456) );
  NOR3_X1 U3345 ( .A1(n2628), .A2(n3458), .A3(n2845), .ZN(n3457) );
  NOR2_X1 U3346 ( .A1(n3387), .A2(n3388), .ZN(n3458) );
  NAND2_X1 U3347 ( .A1(n3387), .A2(n3388), .ZN(n3455) );
  NAND2_X1 U3348 ( .A1(n3459), .A2(n3460), .ZN(n3388) );
  INV_X1 U3349 ( .A(n3461), .ZN(n3460) );
  NOR3_X1 U3350 ( .A1(n2851), .A2(n3462), .A3(n2845), .ZN(n3461) );
  NOR2_X1 U3351 ( .A1(n3384), .A2(n3382), .ZN(n3462) );
  NAND2_X1 U3352 ( .A1(n3382), .A2(n3384), .ZN(n3459) );
  NAND2_X1 U3353 ( .A1(n3463), .A2(n3464), .ZN(n3384) );
  INV_X1 U3354 ( .A(n3465), .ZN(n3464) );
  NOR3_X1 U3355 ( .A1(n2577), .A2(n3466), .A3(n2845), .ZN(n3465) );
  NOR2_X1 U3356 ( .A1(n3380), .A2(n3378), .ZN(n3466) );
  NAND2_X1 U3357 ( .A1(n3378), .A2(n3380), .ZN(n3463) );
  NAND2_X1 U3358 ( .A1(n3342), .A2(n3467), .ZN(n3380) );
  NAND2_X1 U3359 ( .A1(n3341), .A2(n3343), .ZN(n3467) );
  NAND2_X1 U3360 ( .A1(n3468), .A2(n3469), .ZN(n3343) );
  INV_X1 U3361 ( .A(n3470), .ZN(n3469) );
  NAND2_X1 U3362 ( .A1(b_11_), .A2(a_10_), .ZN(n3468) );
  XNOR2_X1 U3363 ( .A(n3471), .B(n3472), .ZN(n3341) );
  NAND2_X1 U3364 ( .A1(n3473), .A2(n3474), .ZN(n3471) );
  NAND2_X1 U3365 ( .A1(n3470), .A2(a_10_), .ZN(n3342) );
  NOR2_X1 U3366 ( .A1(n3475), .A2(n3476), .ZN(n3470) );
  INV_X1 U3367 ( .A(n3477), .ZN(n3476) );
  NAND2_X1 U3368 ( .A1(n3349), .A2(n3478), .ZN(n3477) );
  NAND2_X1 U3369 ( .A1(n2847), .A2(n3350), .ZN(n3478) );
  XOR2_X1 U3370 ( .A(n3479), .B(n3480), .Z(n3349) );
  XNOR2_X1 U3371 ( .A(n3481), .B(n3482), .ZN(n3479) );
  NOR2_X1 U3372 ( .A1(n3350), .A2(n2847), .ZN(n3475) );
  NOR2_X1 U3373 ( .A1(n2845), .A2(n2846), .ZN(n2847) );
  NAND2_X1 U3374 ( .A1(n3483), .A2(n3484), .ZN(n3350) );
  NAND2_X1 U3375 ( .A1(n3376), .A2(n3485), .ZN(n3484) );
  INV_X1 U3376 ( .A(n3486), .ZN(n3485) );
  NOR2_X1 U3377 ( .A1(n3377), .A2(n3375), .ZN(n3486) );
  NOR2_X1 U3378 ( .A1(n2845), .A2(n2844), .ZN(n3376) );
  NAND2_X1 U3379 ( .A1(n3375), .A2(n3377), .ZN(n3483) );
  NAND2_X1 U3380 ( .A1(n3487), .A2(n3488), .ZN(n3377) );
  NAND2_X1 U3381 ( .A1(n3371), .A2(n3489), .ZN(n3488) );
  INV_X1 U3382 ( .A(n3490), .ZN(n3489) );
  NOR2_X1 U3383 ( .A1(n3372), .A2(n3373), .ZN(n3490) );
  NOR2_X1 U3384 ( .A1(n2845), .A2(n2842), .ZN(n3371) );
  NAND2_X1 U3385 ( .A1(n3373), .A2(n3372), .ZN(n3487) );
  NAND2_X1 U3386 ( .A1(n3491), .A2(n3492), .ZN(n3372) );
  NAND2_X1 U3387 ( .A1(b_10_), .A2(n3493), .ZN(n3492) );
  NAND2_X1 U3388 ( .A1(n3049), .A2(n3494), .ZN(n3493) );
  NAND2_X1 U3389 ( .A1(a_14_), .A2(n3495), .ZN(n3494) );
  NAND2_X1 U3390 ( .A1(b_9_), .A2(n3496), .ZN(n3491) );
  NAND2_X1 U3391 ( .A1(n2426), .A2(n3497), .ZN(n3496) );
  NAND2_X1 U3392 ( .A1(a_15_), .A2(n2848), .ZN(n3497) );
  NOR3_X1 U3393 ( .A1(n2848), .A2(n2845), .A3(n3043), .ZN(n3373) );
  XNOR2_X1 U3394 ( .A(n3498), .B(n3499), .ZN(n3375) );
  XOR2_X1 U3395 ( .A(n3500), .B(n3501), .Z(n3499) );
  XOR2_X1 U3396 ( .A(n3502), .B(n3503), .Z(n3378) );
  XOR2_X1 U3397 ( .A(n3504), .B(n2551), .Z(n3502) );
  XNOR2_X1 U3398 ( .A(n3505), .B(n3506), .ZN(n3382) );
  XOR2_X1 U3399 ( .A(n3507), .B(n3508), .Z(n3506) );
  NAND2_X1 U3400 ( .A1(b_10_), .A2(a_9_), .ZN(n3508) );
  XNOR2_X1 U3401 ( .A(n3509), .B(n3510), .ZN(n3387) );
  XOR2_X1 U3402 ( .A(n3511), .B(n3512), .Z(n3510) );
  NAND2_X1 U3403 ( .A1(b_10_), .A2(a_8_), .ZN(n3512) );
  XNOR2_X1 U3404 ( .A(n3513), .B(n3514), .ZN(n3390) );
  XNOR2_X1 U3405 ( .A(n3515), .B(n3516), .ZN(n3513) );
  NOR2_X1 U3406 ( .A1(n2628), .A2(n2848), .ZN(n3516) );
  XNOR2_X1 U3407 ( .A(n3517), .B(n3518), .ZN(n3394) );
  XOR2_X1 U3408 ( .A(n3519), .B(n3520), .Z(n3518) );
  NAND2_X1 U3409 ( .A1(b_10_), .A2(a_6_), .ZN(n3520) );
  XOR2_X1 U3410 ( .A(n3521), .B(n3522), .Z(n3399) );
  XOR2_X1 U3411 ( .A(n3523), .B(n3524), .Z(n3522) );
  NAND2_X1 U3412 ( .A1(b_10_), .A2(a_5_), .ZN(n3524) );
  INV_X1 U3413 ( .A(n3403), .ZN(n3442) );
  XOR2_X1 U3414 ( .A(n3525), .B(n3526), .Z(n3403) );
  XOR2_X1 U3415 ( .A(n3527), .B(n3528), .Z(n3526) );
  NAND2_X1 U3416 ( .A1(b_10_), .A2(a_4_), .ZN(n3528) );
  XNOR2_X1 U3417 ( .A(n3529), .B(n3530), .ZN(n3407) );
  XOR2_X1 U3418 ( .A(n3531), .B(n3532), .Z(n3530) );
  XOR2_X1 U3419 ( .A(n2363), .B(n2362), .Z(n2356) );
  NAND3_X1 U3420 ( .A1(n2362), .A2(n2363), .A3(n2921), .ZN(n2358) );
  INV_X1 U3421 ( .A(n2361), .ZN(n2921) );
  NAND2_X1 U3422 ( .A1(n3533), .A2(n2919), .ZN(n2361) );
  NAND2_X1 U3423 ( .A1(n3534), .A2(n3535), .ZN(n3533) );
  XOR2_X1 U3424 ( .A(n3536), .B(n3537), .Z(n3535) );
  NAND2_X1 U3425 ( .A1(n3416), .A2(n3538), .ZN(n2363) );
  NAND2_X1 U3426 ( .A1(n3415), .A2(n3417), .ZN(n3538) );
  NAND2_X1 U3427 ( .A1(n3539), .A2(n3540), .ZN(n3417) );
  NAND2_X1 U3428 ( .A1(b_10_), .A2(a_0_), .ZN(n3540) );
  XOR2_X1 U3429 ( .A(n3541), .B(n3542), .Z(n3415) );
  XOR2_X1 U3430 ( .A(n3543), .B(n3544), .Z(n3541) );
  NOR2_X1 U3431 ( .A1(n2790), .A2(n3495), .ZN(n3544) );
  NAND2_X1 U3432 ( .A1(a_0_), .A2(n3545), .ZN(n3416) );
  INV_X1 U3433 ( .A(n3539), .ZN(n3545) );
  NOR2_X1 U3434 ( .A1(n3546), .A2(n3547), .ZN(n3539) );
  NOR3_X1 U3435 ( .A1(n2790), .A2(n3548), .A3(n2848), .ZN(n3547) );
  INV_X1 U3436 ( .A(n3549), .ZN(n3548) );
  NAND2_X1 U3437 ( .A1(n3424), .A2(n3422), .ZN(n3549) );
  NOR2_X1 U3438 ( .A1(n3422), .A2(n3424), .ZN(n3546) );
  NOR2_X1 U3439 ( .A1(n3550), .A2(n3551), .ZN(n3424) );
  INV_X1 U3440 ( .A(n3552), .ZN(n3551) );
  NAND2_X1 U3441 ( .A1(n3433), .A2(n3553), .ZN(n3552) );
  NAND2_X1 U3442 ( .A1(n3432), .A2(n3431), .ZN(n3553) );
  NOR2_X1 U3443 ( .A1(n2848), .A2(n2860), .ZN(n3433) );
  NOR2_X1 U3444 ( .A1(n3431), .A2(n3432), .ZN(n3550) );
  NOR2_X1 U3445 ( .A1(n3554), .A2(n3555), .ZN(n3432) );
  NOR2_X1 U3446 ( .A1(n3532), .A2(n3556), .ZN(n3555) );
  NOR2_X1 U3447 ( .A1(n3531), .A2(n3529), .ZN(n3556) );
  NAND2_X1 U3448 ( .A1(b_10_), .A2(a_3_), .ZN(n3532) );
  INV_X1 U3449 ( .A(n3557), .ZN(n3554) );
  NAND2_X1 U3450 ( .A1(n3529), .A2(n3531), .ZN(n3557) );
  NAND2_X1 U3451 ( .A1(n3558), .A2(n3559), .ZN(n3531) );
  NAND3_X1 U3452 ( .A1(a_4_), .A2(n3560), .A3(b_10_), .ZN(n3559) );
  INV_X1 U3453 ( .A(n3561), .ZN(n3560) );
  NOR2_X1 U3454 ( .A1(n3527), .A2(n3525), .ZN(n3561) );
  NAND2_X1 U3455 ( .A1(n3525), .A2(n3527), .ZN(n3558) );
  NAND2_X1 U3456 ( .A1(n3562), .A2(n3563), .ZN(n3527) );
  INV_X1 U3457 ( .A(n3564), .ZN(n3563) );
  NOR3_X1 U3458 ( .A1(n2679), .A2(n3565), .A3(n2848), .ZN(n3564) );
  NOR2_X1 U3459 ( .A1(n3523), .A2(n3521), .ZN(n3565) );
  NAND2_X1 U3460 ( .A1(n3521), .A2(n3523), .ZN(n3562) );
  NAND2_X1 U3461 ( .A1(n3566), .A2(n3567), .ZN(n3523) );
  INV_X1 U3462 ( .A(n3568), .ZN(n3567) );
  NOR3_X1 U3463 ( .A1(n2854), .A2(n3569), .A3(n2848), .ZN(n3568) );
  NOR2_X1 U3464 ( .A1(n3519), .A2(n3517), .ZN(n3569) );
  NAND2_X1 U3465 ( .A1(n3517), .A2(n3519), .ZN(n3566) );
  NAND2_X1 U3466 ( .A1(n3570), .A2(n3571), .ZN(n3519) );
  NAND3_X1 U3467 ( .A1(a_7_), .A2(n3572), .A3(b_10_), .ZN(n3571) );
  NAND2_X1 U3468 ( .A1(n3515), .A2(n3514), .ZN(n3572) );
  INV_X1 U3469 ( .A(n3573), .ZN(n3570) );
  NOR2_X1 U3470 ( .A1(n3514), .A2(n3515), .ZN(n3573) );
  NOR2_X1 U3471 ( .A1(n3574), .A2(n3575), .ZN(n3515) );
  NOR3_X1 U3472 ( .A1(n2851), .A2(n3576), .A3(n2848), .ZN(n3575) );
  NOR2_X1 U3473 ( .A1(n3511), .A2(n3509), .ZN(n3576) );
  INV_X1 U3474 ( .A(n3577), .ZN(n3574) );
  NAND2_X1 U3475 ( .A1(n3509), .A2(n3511), .ZN(n3577) );
  NAND2_X1 U3476 ( .A1(n3578), .A2(n3579), .ZN(n3511) );
  NAND3_X1 U3477 ( .A1(a_9_), .A2(n3580), .A3(b_10_), .ZN(n3579) );
  INV_X1 U3478 ( .A(n3581), .ZN(n3580) );
  NOR2_X1 U3479 ( .A1(n3507), .A2(n3505), .ZN(n3581) );
  NAND2_X1 U3480 ( .A1(n3505), .A2(n3507), .ZN(n3578) );
  NAND2_X1 U3481 ( .A1(n3582), .A2(n3583), .ZN(n3507) );
  NAND2_X1 U3482 ( .A1(n3503), .A2(n3584), .ZN(n3583) );
  NAND2_X1 U3483 ( .A1(n3504), .A2(n2551), .ZN(n3584) );
  INV_X1 U3484 ( .A(n3585), .ZN(n2551) );
  INV_X1 U3485 ( .A(n3586), .ZN(n3504) );
  XNOR2_X1 U3486 ( .A(n3587), .B(n3588), .ZN(n3503) );
  NAND2_X1 U3487 ( .A1(n3589), .A2(n3590), .ZN(n3587) );
  NAND2_X1 U3488 ( .A1(n3585), .A2(n3586), .ZN(n3582) );
  NAND2_X1 U3489 ( .A1(n3473), .A2(n3591), .ZN(n3586) );
  NAND2_X1 U3490 ( .A1(n3472), .A2(n3474), .ZN(n3591) );
  NAND2_X1 U3491 ( .A1(n3592), .A2(n3593), .ZN(n3474) );
  NAND2_X1 U3492 ( .A1(b_10_), .A2(a_11_), .ZN(n3593) );
  XNOR2_X1 U3493 ( .A(n3594), .B(n3595), .ZN(n3472) );
  XNOR2_X1 U3494 ( .A(n3596), .B(n3597), .ZN(n3594) );
  INV_X1 U3495 ( .A(n3598), .ZN(n3473) );
  NOR2_X1 U3496 ( .A1(n2846), .A2(n3592), .ZN(n3598) );
  NOR2_X1 U3497 ( .A1(n3599), .A2(n3600), .ZN(n3592) );
  INV_X1 U3498 ( .A(n3601), .ZN(n3600) );
  NAND2_X1 U3499 ( .A1(n3481), .A2(n3602), .ZN(n3601) );
  NAND2_X1 U3500 ( .A1(n3482), .A2(n3480), .ZN(n3602) );
  NOR2_X1 U3501 ( .A1(n2848), .A2(n2844), .ZN(n3481) );
  NOR2_X1 U3502 ( .A1(n3480), .A2(n3482), .ZN(n3599) );
  NOR2_X1 U3503 ( .A1(n3603), .A2(n3604), .ZN(n3482) );
  INV_X1 U3504 ( .A(n3605), .ZN(n3604) );
  NAND2_X1 U3505 ( .A1(n3498), .A2(n3606), .ZN(n3605) );
  NAND2_X1 U3506 ( .A1(n3607), .A2(n3500), .ZN(n3606) );
  NOR2_X1 U3507 ( .A1(n2848), .A2(n2842), .ZN(n3498) );
  NOR2_X1 U3508 ( .A1(n3500), .A2(n3607), .ZN(n3603) );
  INV_X1 U3509 ( .A(n3501), .ZN(n3607) );
  NAND2_X1 U3510 ( .A1(n3608), .A2(n3609), .ZN(n3501) );
  NAND2_X1 U3511 ( .A1(b_8_), .A2(n3610), .ZN(n3609) );
  NAND2_X1 U3512 ( .A1(n2426), .A2(n3611), .ZN(n3610) );
  NAND2_X1 U3513 ( .A1(a_15_), .A2(n3495), .ZN(n3611) );
  NAND2_X1 U3514 ( .A1(b_9_), .A2(n3612), .ZN(n3608) );
  NAND2_X1 U3515 ( .A1(n3049), .A2(n3613), .ZN(n3612) );
  NAND2_X1 U3516 ( .A1(a_14_), .A2(n2850), .ZN(n3613) );
  NAND3_X1 U3517 ( .A1(b_9_), .A2(b_10_), .A3(n2840), .ZN(n3500) );
  XOR2_X1 U3518 ( .A(n3614), .B(n3615), .Z(n3480) );
  XOR2_X1 U3519 ( .A(n3616), .B(n3617), .Z(n3615) );
  NOR2_X1 U3520 ( .A1(n2848), .A2(n2849), .ZN(n3585) );
  XNOR2_X1 U3521 ( .A(n3618), .B(n3619), .ZN(n3505) );
  NAND2_X1 U3522 ( .A1(n3620), .A2(n3621), .ZN(n3618) );
  XOR2_X1 U3523 ( .A(n3622), .B(n3623), .Z(n3509) );
  XNOR2_X1 U3524 ( .A(n3624), .B(n2830), .ZN(n3623) );
  XNOR2_X1 U3525 ( .A(n3625), .B(n3626), .ZN(n3514) );
  XOR2_X1 U3526 ( .A(n3627), .B(n3628), .Z(n3626) );
  XOR2_X1 U3527 ( .A(n3629), .B(n3630), .Z(n3517) );
  XOR2_X1 U3528 ( .A(n3631), .B(n3632), .Z(n3629) );
  NOR2_X1 U3529 ( .A1(n2628), .A2(n3495), .ZN(n3632) );
  XNOR2_X1 U3530 ( .A(n3633), .B(n3634), .ZN(n3521) );
  XNOR2_X1 U3531 ( .A(n3635), .B(n3636), .ZN(n3634) );
  XOR2_X1 U3532 ( .A(n3637), .B(n3638), .Z(n3525) );
  XNOR2_X1 U3533 ( .A(n3639), .B(n3640), .ZN(n3637) );
  XNOR2_X1 U3534 ( .A(n3641), .B(n3642), .ZN(n3529) );
  NAND2_X1 U3535 ( .A1(n3643), .A2(n3644), .ZN(n3641) );
  XOR2_X1 U3536 ( .A(n3645), .B(n3646), .Z(n3431) );
  XOR2_X1 U3537 ( .A(n3647), .B(n3648), .Z(n3646) );
  NAND2_X1 U3538 ( .A1(b_9_), .A2(a_3_), .ZN(n3648) );
  XOR2_X1 U3539 ( .A(n3649), .B(n3650), .Z(n3422) );
  XOR2_X1 U3540 ( .A(n3651), .B(n3652), .Z(n3650) );
  NAND2_X1 U3541 ( .A1(b_9_), .A2(a_2_), .ZN(n3652) );
  XOR2_X1 U3542 ( .A(n3653), .B(n3654), .Z(n2362) );
  XNOR2_X1 U3543 ( .A(n3655), .B(n3656), .ZN(n3654) );
  NAND2_X1 U3544 ( .A1(b_9_), .A2(a_0_), .ZN(n3656) );
  NAND2_X1 U3545 ( .A1(n3657), .A2(n3658), .ZN(n2919) );
  INV_X1 U3546 ( .A(n3534), .ZN(n3658) );
  NOR2_X1 U3547 ( .A1(n3659), .A2(n3660), .ZN(n3534) );
  INV_X1 U3548 ( .A(n3661), .ZN(n3660) );
  NAND3_X1 U3549 ( .A1(a_0_), .A2(n3662), .A3(b_9_), .ZN(n3661) );
  NAND2_X1 U3550 ( .A1(n3655), .A2(n3653), .ZN(n3662) );
  NOR2_X1 U3551 ( .A1(n3653), .A2(n3655), .ZN(n3659) );
  NOR2_X1 U3552 ( .A1(n3663), .A2(n3664), .ZN(n3655) );
  NOR3_X1 U3553 ( .A1(n2790), .A2(n3665), .A3(n3495), .ZN(n3664) );
  NOR2_X1 U3554 ( .A1(n3543), .A2(n3542), .ZN(n3665) );
  INV_X1 U3555 ( .A(n3666), .ZN(n3663) );
  NAND2_X1 U3556 ( .A1(n3542), .A2(n3543), .ZN(n3666) );
  NAND2_X1 U3557 ( .A1(n3667), .A2(n3668), .ZN(n3543) );
  NAND3_X1 U3558 ( .A1(a_2_), .A2(n3669), .A3(b_9_), .ZN(n3668) );
  INV_X1 U3559 ( .A(n3670), .ZN(n3669) );
  NOR2_X1 U3560 ( .A1(n3651), .A2(n3649), .ZN(n3670) );
  NAND2_X1 U3561 ( .A1(n3649), .A2(n3651), .ZN(n3667) );
  NAND2_X1 U3562 ( .A1(n3671), .A2(n3672), .ZN(n3651) );
  INV_X1 U3563 ( .A(n3673), .ZN(n3672) );
  NOR3_X1 U3564 ( .A1(n2739), .A2(n3674), .A3(n3495), .ZN(n3673) );
  NOR2_X1 U3565 ( .A1(n3647), .A2(n3645), .ZN(n3674) );
  NAND2_X1 U3566 ( .A1(n3645), .A2(n3647), .ZN(n3671) );
  NAND2_X1 U3567 ( .A1(n3643), .A2(n3675), .ZN(n3647) );
  NAND2_X1 U3568 ( .A1(n3642), .A2(n3644), .ZN(n3675) );
  NAND2_X1 U3569 ( .A1(n3676), .A2(n3677), .ZN(n3644) );
  NAND2_X1 U3570 ( .A1(b_9_), .A2(a_4_), .ZN(n3677) );
  XNOR2_X1 U3571 ( .A(n3678), .B(n3679), .ZN(n3642) );
  XOR2_X1 U3572 ( .A(n3680), .B(n3681), .Z(n3679) );
  INV_X1 U3573 ( .A(n3682), .ZN(n3643) );
  NOR2_X1 U3574 ( .A1(n2857), .A2(n3676), .ZN(n3682) );
  NOR2_X1 U3575 ( .A1(n3683), .A2(n3684), .ZN(n3676) );
  NOR2_X1 U3576 ( .A1(n3639), .A2(n3685), .ZN(n3684) );
  NOR2_X1 U3577 ( .A1(n3640), .A2(n3638), .ZN(n3685) );
  NAND2_X1 U3578 ( .A1(b_9_), .A2(a_5_), .ZN(n3639) );
  INV_X1 U3579 ( .A(n3686), .ZN(n3683) );
  NAND2_X1 U3580 ( .A1(n3638), .A2(n3640), .ZN(n3686) );
  NAND2_X1 U3581 ( .A1(n3687), .A2(n3688), .ZN(n3640) );
  NAND2_X1 U3582 ( .A1(n3636), .A2(n3689), .ZN(n3688) );
  INV_X1 U3583 ( .A(n3690), .ZN(n3689) );
  NOR2_X1 U3584 ( .A1(n3635), .A2(n3633), .ZN(n3690) );
  NOR2_X1 U3585 ( .A1(n3495), .A2(n2854), .ZN(n3636) );
  NAND2_X1 U3586 ( .A1(n3633), .A2(n3635), .ZN(n3687) );
  NAND2_X1 U3587 ( .A1(n3691), .A2(n3692), .ZN(n3635) );
  INV_X1 U3588 ( .A(n3693), .ZN(n3692) );
  NOR3_X1 U3589 ( .A1(n2628), .A2(n3694), .A3(n3495), .ZN(n3693) );
  NOR2_X1 U3590 ( .A1(n3631), .A2(n3630), .ZN(n3694) );
  NAND2_X1 U3591 ( .A1(n3630), .A2(n3631), .ZN(n3691) );
  NAND2_X1 U3592 ( .A1(n3695), .A2(n3696), .ZN(n3631) );
  NAND2_X1 U3593 ( .A1(n3628), .A2(n3697), .ZN(n3696) );
  INV_X1 U3594 ( .A(n3698), .ZN(n3697) );
  NOR2_X1 U3595 ( .A1(n3625), .A2(n3627), .ZN(n3698) );
  NOR2_X1 U3596 ( .A1(n3495), .A2(n2851), .ZN(n3628) );
  NAND2_X1 U3597 ( .A1(n3627), .A2(n3625), .ZN(n3695) );
  XNOR2_X1 U3598 ( .A(n3699), .B(n3700), .ZN(n3625) );
  XOR2_X1 U3599 ( .A(n3701), .B(n3702), .Z(n3700) );
  NAND2_X1 U3600 ( .A1(b_8_), .A2(a_9_), .ZN(n3702) );
  NOR2_X1 U3601 ( .A1(n3703), .A2(n3704), .ZN(n3627) );
  INV_X1 U3602 ( .A(n3705), .ZN(n3704) );
  NAND2_X1 U3603 ( .A1(n3622), .A2(n3706), .ZN(n3705) );
  NAND2_X1 U3604 ( .A1(n2830), .A2(n3624), .ZN(n3706) );
  XOR2_X1 U3605 ( .A(n3707), .B(n3708), .Z(n3622) );
  NAND2_X1 U3606 ( .A1(n3709), .A2(n3710), .ZN(n3707) );
  NOR2_X1 U3607 ( .A1(n3624), .A2(n2830), .ZN(n3703) );
  NOR2_X1 U3608 ( .A1(n3495), .A2(n2577), .ZN(n2830) );
  NAND2_X1 U3609 ( .A1(n3620), .A2(n3711), .ZN(n3624) );
  NAND2_X1 U3610 ( .A1(n3619), .A2(n3621), .ZN(n3711) );
  NAND2_X1 U3611 ( .A1(n3712), .A2(n3713), .ZN(n3621) );
  NAND2_X1 U3612 ( .A1(b_9_), .A2(a_10_), .ZN(n3713) );
  INV_X1 U3613 ( .A(n3714), .ZN(n3712) );
  XNOR2_X1 U3614 ( .A(n3715), .B(n3716), .ZN(n3619) );
  NAND2_X1 U3615 ( .A1(n3717), .A2(n3718), .ZN(n3715) );
  NAND2_X1 U3616 ( .A1(a_10_), .A2(n3714), .ZN(n3620) );
  NAND2_X1 U3617 ( .A1(n3589), .A2(n3719), .ZN(n3714) );
  NAND2_X1 U3618 ( .A1(n3588), .A2(n3590), .ZN(n3719) );
  NAND2_X1 U3619 ( .A1(n3720), .A2(n3721), .ZN(n3590) );
  NAND2_X1 U3620 ( .A1(b_9_), .A2(a_11_), .ZN(n3721) );
  XNOR2_X1 U3621 ( .A(n3722), .B(n3723), .ZN(n3588) );
  XNOR2_X1 U3622 ( .A(n3724), .B(n3725), .ZN(n3722) );
  INV_X1 U3623 ( .A(n3726), .ZN(n3589) );
  NOR2_X1 U3624 ( .A1(n2846), .A2(n3720), .ZN(n3726) );
  NOR2_X1 U3625 ( .A1(n3727), .A2(n3728), .ZN(n3720) );
  INV_X1 U3626 ( .A(n3729), .ZN(n3728) );
  NAND2_X1 U3627 ( .A1(n3596), .A2(n3730), .ZN(n3729) );
  NAND2_X1 U3628 ( .A1(n3597), .A2(n3595), .ZN(n3730) );
  NOR2_X1 U3629 ( .A1(n3495), .A2(n2844), .ZN(n3596) );
  NOR2_X1 U3630 ( .A1(n3595), .A2(n3597), .ZN(n3727) );
  NOR2_X1 U3631 ( .A1(n3731), .A2(n3732), .ZN(n3597) );
  INV_X1 U3632 ( .A(n3733), .ZN(n3732) );
  NAND2_X1 U3633 ( .A1(n3614), .A2(n3734), .ZN(n3733) );
  NAND2_X1 U3634 ( .A1(n3735), .A2(n3616), .ZN(n3734) );
  NOR2_X1 U3635 ( .A1(n3495), .A2(n2842), .ZN(n3614) );
  NOR2_X1 U3636 ( .A1(n3616), .A2(n3735), .ZN(n3731) );
  INV_X1 U3637 ( .A(n3617), .ZN(n3735) );
  NAND2_X1 U3638 ( .A1(n3736), .A2(n3737), .ZN(n3617) );
  NAND2_X1 U3639 ( .A1(b_7_), .A2(n3738), .ZN(n3737) );
  NAND2_X1 U3640 ( .A1(n2426), .A2(n3739), .ZN(n3738) );
  NAND2_X1 U3641 ( .A1(a_15_), .A2(n2850), .ZN(n3739) );
  NAND2_X1 U3642 ( .A1(b_8_), .A2(n3740), .ZN(n3736) );
  NAND2_X1 U3643 ( .A1(n3049), .A2(n3741), .ZN(n3740) );
  NAND2_X1 U3644 ( .A1(a_14_), .A2(n2852), .ZN(n3741) );
  NAND3_X1 U3645 ( .A1(b_8_), .A2(b_9_), .A3(n2840), .ZN(n3616) );
  XOR2_X1 U3646 ( .A(n3742), .B(n3743), .Z(n3595) );
  XOR2_X1 U3647 ( .A(n3744), .B(n3745), .Z(n3743) );
  XNOR2_X1 U3648 ( .A(n3746), .B(n3747), .ZN(n3630) );
  XOR2_X1 U3649 ( .A(n3748), .B(n3749), .Z(n3746) );
  XNOR2_X1 U3650 ( .A(n3750), .B(n3751), .ZN(n3633) );
  XOR2_X1 U3651 ( .A(n3752), .B(n3753), .Z(n3751) );
  NAND2_X1 U3652 ( .A1(b_8_), .A2(a_7_), .ZN(n3753) );
  XOR2_X1 U3653 ( .A(n3754), .B(n3755), .Z(n3638) );
  XNOR2_X1 U3654 ( .A(n3756), .B(n3757), .ZN(n3755) );
  NAND2_X1 U3655 ( .A1(b_8_), .A2(a_6_), .ZN(n3757) );
  XNOR2_X1 U3656 ( .A(n3758), .B(n3759), .ZN(n3645) );
  XNOR2_X1 U3657 ( .A(n3760), .B(n3761), .ZN(n3758) );
  XNOR2_X1 U3658 ( .A(n3762), .B(n3763), .ZN(n3649) );
  XNOR2_X1 U3659 ( .A(n3764), .B(n3765), .ZN(n3762) );
  XOR2_X1 U3660 ( .A(n3766), .B(n3767), .Z(n3542) );
  XOR2_X1 U3661 ( .A(n3768), .B(n3769), .Z(n3766) );
  XOR2_X1 U3662 ( .A(n3770), .B(n3771), .Z(n3653) );
  XNOR2_X1 U3663 ( .A(n3772), .B(n3773), .ZN(n3771) );
  XNOR2_X1 U3664 ( .A(n3536), .B(n3537), .ZN(n3657) );
  NAND2_X1 U3665 ( .A1(n3774), .A2(n3775), .ZN(n3536) );
  XOR2_X1 U3666 ( .A(n2376), .B(n2377), .Z(n2367) );
  NAND3_X1 U3667 ( .A1(n2376), .A2(n2377), .A3(n2918), .ZN(n2372) );
  INV_X1 U3668 ( .A(n2375), .ZN(n2918) );
  NAND2_X1 U3669 ( .A1(n3776), .A2(n2916), .ZN(n2375) );
  NAND2_X1 U3670 ( .A1(n3777), .A2(n3778), .ZN(n3776) );
  XOR2_X1 U3671 ( .A(n3779), .B(n3780), .Z(n3777) );
  NAND2_X1 U3672 ( .A1(n3774), .A2(n3781), .ZN(n2377) );
  NAND2_X1 U3673 ( .A1(n3537), .A2(n3775), .ZN(n3781) );
  NAND2_X1 U3674 ( .A1(n3782), .A2(n3783), .ZN(n3775) );
  NAND2_X1 U3675 ( .A1(b_8_), .A2(a_0_), .ZN(n3783) );
  INV_X1 U3676 ( .A(n3784), .ZN(n3782) );
  XNOR2_X1 U3677 ( .A(n3785), .B(n3786), .ZN(n3537) );
  XNOR2_X1 U3678 ( .A(n3787), .B(n3788), .ZN(n3785) );
  NOR2_X1 U3679 ( .A1(n2790), .A2(n2852), .ZN(n3788) );
  NAND2_X1 U3680 ( .A1(a_0_), .A2(n3784), .ZN(n3774) );
  NAND2_X1 U3681 ( .A1(n3789), .A2(n3790), .ZN(n3784) );
  NAND2_X1 U3682 ( .A1(n3773), .A2(n3791), .ZN(n3790) );
  INV_X1 U3683 ( .A(n3792), .ZN(n3791) );
  NOR2_X1 U3684 ( .A1(n3772), .A2(n3770), .ZN(n3792) );
  NOR2_X1 U3685 ( .A1(n2850), .A2(n2790), .ZN(n3773) );
  NAND2_X1 U3686 ( .A1(n3770), .A2(n3772), .ZN(n3789) );
  NAND2_X1 U3687 ( .A1(n3793), .A2(n3794), .ZN(n3772) );
  NAND2_X1 U3688 ( .A1(n3769), .A2(n3795), .ZN(n3794) );
  INV_X1 U3689 ( .A(n3796), .ZN(n3795) );
  NOR2_X1 U3690 ( .A1(n3768), .A2(n3767), .ZN(n3796) );
  NOR2_X1 U3691 ( .A1(n2850), .A2(n2860), .ZN(n3769) );
  NAND2_X1 U3692 ( .A1(n3767), .A2(n3768), .ZN(n3793) );
  NAND2_X1 U3693 ( .A1(n3797), .A2(n3798), .ZN(n3768) );
  NAND2_X1 U3694 ( .A1(n3765), .A2(n3799), .ZN(n3798) );
  NAND2_X1 U3695 ( .A1(n3763), .A2(n3764), .ZN(n3799) );
  NOR2_X1 U3696 ( .A1(n2850), .A2(n2739), .ZN(n3765) );
  INV_X1 U3697 ( .A(n3800), .ZN(n3797) );
  NOR2_X1 U3698 ( .A1(n3763), .A2(n3764), .ZN(n3800) );
  NOR2_X1 U3699 ( .A1(n3801), .A2(n3802), .ZN(n3764) );
  INV_X1 U3700 ( .A(n3803), .ZN(n3802) );
  NAND2_X1 U3701 ( .A1(n3761), .A2(n3804), .ZN(n3803) );
  NAND2_X1 U3702 ( .A1(n3760), .A2(n3759), .ZN(n3804) );
  NOR2_X1 U3703 ( .A1(n2850), .A2(n2857), .ZN(n3761) );
  NOR2_X1 U3704 ( .A1(n3759), .A2(n3760), .ZN(n3801) );
  NOR2_X1 U3705 ( .A1(n3805), .A2(n3806), .ZN(n3760) );
  NOR2_X1 U3706 ( .A1(n3681), .A2(n3807), .ZN(n3806) );
  NOR2_X1 U3707 ( .A1(n3680), .A2(n3678), .ZN(n3807) );
  NAND2_X1 U3708 ( .A1(b_8_), .A2(a_5_), .ZN(n3681) );
  INV_X1 U3709 ( .A(n3808), .ZN(n3805) );
  NAND2_X1 U3710 ( .A1(n3678), .A2(n3680), .ZN(n3808) );
  NAND2_X1 U3711 ( .A1(n3809), .A2(n3810), .ZN(n3680) );
  NAND3_X1 U3712 ( .A1(a_6_), .A2(n3811), .A3(b_8_), .ZN(n3810) );
  NAND2_X1 U3713 ( .A1(n3756), .A2(n3754), .ZN(n3811) );
  INV_X1 U3714 ( .A(n3812), .ZN(n3809) );
  NOR2_X1 U3715 ( .A1(n3754), .A2(n3756), .ZN(n3812) );
  NOR2_X1 U3716 ( .A1(n3813), .A2(n3814), .ZN(n3756) );
  INV_X1 U3717 ( .A(n3815), .ZN(n3814) );
  NAND3_X1 U3718 ( .A1(a_7_), .A2(n3816), .A3(b_8_), .ZN(n3815) );
  NAND2_X1 U3719 ( .A1(n3750), .A2(n3752), .ZN(n3816) );
  NOR2_X1 U3720 ( .A1(n3750), .A2(n3752), .ZN(n3813) );
  NAND2_X1 U3721 ( .A1(n3817), .A2(n3818), .ZN(n3752) );
  NAND2_X1 U3722 ( .A1(n3747), .A2(n3819), .ZN(n3818) );
  NAND2_X1 U3723 ( .A1(n3749), .A2(n3748), .ZN(n3819) );
  INV_X1 U3724 ( .A(n3820), .ZN(n3748) );
  INV_X1 U3725 ( .A(n2602), .ZN(n3749) );
  XOR2_X1 U3726 ( .A(n3821), .B(n3822), .Z(n3747) );
  XOR2_X1 U3727 ( .A(n3823), .B(n3824), .Z(n3822) );
  NAND2_X1 U3728 ( .A1(b_7_), .A2(a_9_), .ZN(n3824) );
  NAND2_X1 U3729 ( .A1(n3820), .A2(n2602), .ZN(n3817) );
  NAND2_X1 U3730 ( .A1(b_8_), .A2(a_8_), .ZN(n2602) );
  NOR2_X1 U3731 ( .A1(n3825), .A2(n3826), .ZN(n3820) );
  NOR3_X1 U3732 ( .A1(n2577), .A2(n3827), .A3(n2850), .ZN(n3826) );
  NOR2_X1 U3733 ( .A1(n3699), .A2(n3701), .ZN(n3827) );
  INV_X1 U3734 ( .A(n3828), .ZN(n3825) );
  NAND2_X1 U3735 ( .A1(n3699), .A2(n3701), .ZN(n3828) );
  NAND2_X1 U3736 ( .A1(n3709), .A2(n3829), .ZN(n3701) );
  NAND2_X1 U3737 ( .A1(n3708), .A2(n3710), .ZN(n3829) );
  NAND2_X1 U3738 ( .A1(n3830), .A2(n3831), .ZN(n3710) );
  NAND2_X1 U3739 ( .A1(b_8_), .A2(a_10_), .ZN(n3831) );
  INV_X1 U3740 ( .A(n3832), .ZN(n3830) );
  XNOR2_X1 U3741 ( .A(n3833), .B(n3834), .ZN(n3708) );
  NAND2_X1 U3742 ( .A1(n3835), .A2(n3836), .ZN(n3833) );
  NAND2_X1 U3743 ( .A1(a_10_), .A2(n3832), .ZN(n3709) );
  NAND2_X1 U3744 ( .A1(n3717), .A2(n3837), .ZN(n3832) );
  NAND2_X1 U3745 ( .A1(n3716), .A2(n3718), .ZN(n3837) );
  NAND2_X1 U3746 ( .A1(n3838), .A2(n3839), .ZN(n3718) );
  NAND2_X1 U3747 ( .A1(b_8_), .A2(a_11_), .ZN(n3839) );
  XNOR2_X1 U3748 ( .A(n3840), .B(n3841), .ZN(n3716) );
  XNOR2_X1 U3749 ( .A(n3842), .B(n3843), .ZN(n3840) );
  INV_X1 U3750 ( .A(n3844), .ZN(n3717) );
  NOR2_X1 U3751 ( .A1(n2846), .A2(n3838), .ZN(n3844) );
  NOR2_X1 U3752 ( .A1(n3845), .A2(n3846), .ZN(n3838) );
  INV_X1 U3753 ( .A(n3847), .ZN(n3846) );
  NAND2_X1 U3754 ( .A1(n3724), .A2(n3848), .ZN(n3847) );
  NAND2_X1 U3755 ( .A1(n3725), .A2(n3723), .ZN(n3848) );
  NOR2_X1 U3756 ( .A1(n2850), .A2(n2844), .ZN(n3724) );
  NOR2_X1 U3757 ( .A1(n3723), .A2(n3725), .ZN(n3845) );
  NOR2_X1 U3758 ( .A1(n3849), .A2(n3850), .ZN(n3725) );
  INV_X1 U3759 ( .A(n3851), .ZN(n3850) );
  NAND2_X1 U3760 ( .A1(n3742), .A2(n3852), .ZN(n3851) );
  NAND2_X1 U3761 ( .A1(n3853), .A2(n3744), .ZN(n3852) );
  NOR2_X1 U3762 ( .A1(n2850), .A2(n2842), .ZN(n3742) );
  NOR2_X1 U3763 ( .A1(n3744), .A2(n3853), .ZN(n3849) );
  INV_X1 U3764 ( .A(n3745), .ZN(n3853) );
  NAND2_X1 U3765 ( .A1(n3854), .A2(n3855), .ZN(n3745) );
  NAND2_X1 U3766 ( .A1(b_6_), .A2(n3856), .ZN(n3855) );
  NAND2_X1 U3767 ( .A1(n2426), .A2(n3857), .ZN(n3856) );
  NAND2_X1 U3768 ( .A1(a_15_), .A2(n2852), .ZN(n3857) );
  NAND2_X1 U3769 ( .A1(b_7_), .A2(n3858), .ZN(n3854) );
  NAND2_X1 U3770 ( .A1(n3049), .A2(n3859), .ZN(n3858) );
  NAND2_X1 U3771 ( .A1(a_14_), .A2(n2853), .ZN(n3859) );
  NAND3_X1 U3772 ( .A1(b_7_), .A2(b_8_), .A3(n2840), .ZN(n3744) );
  XOR2_X1 U3773 ( .A(n3860), .B(n3861), .Z(n3723) );
  XOR2_X1 U3774 ( .A(n3862), .B(n3863), .Z(n3861) );
  XNOR2_X1 U3775 ( .A(n3864), .B(n3865), .ZN(n3699) );
  NAND2_X1 U3776 ( .A1(n3866), .A2(n3867), .ZN(n3864) );
  XNOR2_X1 U3777 ( .A(n3868), .B(n3869), .ZN(n3750) );
  XOR2_X1 U3778 ( .A(n3870), .B(n3871), .Z(n3868) );
  XOR2_X1 U3779 ( .A(n3872), .B(n3873), .Z(n3754) );
  XOR2_X1 U3780 ( .A(n3874), .B(n3875), .Z(n3872) );
  XOR2_X1 U3781 ( .A(n3876), .B(n3877), .Z(n3678) );
  NOR2_X1 U3782 ( .A1(n3878), .A2(n3879), .ZN(n3877) );
  NOR2_X1 U3783 ( .A1(n3880), .A2(n3881), .ZN(n3878) );
  NOR2_X1 U3784 ( .A1(n2854), .A2(n2852), .ZN(n3881) );
  INV_X1 U3785 ( .A(n3882), .ZN(n3880) );
  XOR2_X1 U3786 ( .A(n3883), .B(n3884), .Z(n3759) );
  XOR2_X1 U3787 ( .A(n3885), .B(n3886), .Z(n3884) );
  NAND2_X1 U3788 ( .A1(b_7_), .A2(a_5_), .ZN(n3886) );
  XNOR2_X1 U3789 ( .A(n3887), .B(n3888), .ZN(n3763) );
  XNOR2_X1 U3790 ( .A(n3889), .B(n3890), .ZN(n3888) );
  NAND2_X1 U3791 ( .A1(b_7_), .A2(a_4_), .ZN(n3890) );
  XNOR2_X1 U3792 ( .A(n3891), .B(n3892), .ZN(n3767) );
  XNOR2_X1 U3793 ( .A(n3893), .B(n3894), .ZN(n3891) );
  NOR2_X1 U3794 ( .A1(n2739), .A2(n2852), .ZN(n3894) );
  XOR2_X1 U3795 ( .A(n3895), .B(n3896), .Z(n3770) );
  XNOR2_X1 U3796 ( .A(n3897), .B(n3898), .ZN(n3896) );
  NAND2_X1 U3797 ( .A1(b_7_), .A2(a_2_), .ZN(n3898) );
  XNOR2_X1 U3798 ( .A(n3899), .B(n3900), .ZN(n2376) );
  XNOR2_X1 U3799 ( .A(n3901), .B(n3902), .ZN(n3899) );
  NOR2_X1 U3800 ( .A1(n2865), .A2(n2852), .ZN(n3902) );
  NAND2_X1 U3801 ( .A1(n3903), .A2(n3904), .ZN(n2916) );
  INV_X1 U3802 ( .A(n3778), .ZN(n3904) );
  NOR2_X1 U3803 ( .A1(n3905), .A2(n3906), .ZN(n3778) );
  INV_X1 U3804 ( .A(n3907), .ZN(n3906) );
  NAND3_X1 U3805 ( .A1(a_0_), .A2(n3908), .A3(b_7_), .ZN(n3907) );
  NAND2_X1 U3806 ( .A1(n3901), .A2(n3900), .ZN(n3908) );
  NOR2_X1 U3807 ( .A1(n3900), .A2(n3901), .ZN(n3905) );
  NOR2_X1 U3808 ( .A1(n3909), .A2(n3910), .ZN(n3901) );
  NOR3_X1 U3809 ( .A1(n2790), .A2(n3911), .A3(n2852), .ZN(n3910) );
  INV_X1 U3810 ( .A(n3912), .ZN(n3911) );
  NAND2_X1 U3811 ( .A1(n3786), .A2(n3787), .ZN(n3912) );
  NOR2_X1 U3812 ( .A1(n3786), .A2(n3787), .ZN(n3909) );
  NOR2_X1 U3813 ( .A1(n3913), .A2(n3914), .ZN(n3787) );
  NOR3_X1 U3814 ( .A1(n2860), .A2(n3915), .A3(n2852), .ZN(n3914) );
  INV_X1 U3815 ( .A(n3916), .ZN(n3915) );
  NAND2_X1 U3816 ( .A1(n3895), .A2(n3897), .ZN(n3916) );
  NOR2_X1 U3817 ( .A1(n3895), .A2(n3897), .ZN(n3913) );
  NOR2_X1 U3818 ( .A1(n3917), .A2(n3918), .ZN(n3897) );
  INV_X1 U3819 ( .A(n3919), .ZN(n3918) );
  NAND3_X1 U3820 ( .A1(a_3_), .A2(n3920), .A3(b_7_), .ZN(n3919) );
  NAND2_X1 U3821 ( .A1(n3892), .A2(n3893), .ZN(n3920) );
  NOR2_X1 U3822 ( .A1(n3892), .A2(n3893), .ZN(n3917) );
  NOR2_X1 U3823 ( .A1(n3921), .A2(n3922), .ZN(n3893) );
  NOR3_X1 U3824 ( .A1(n2857), .A2(n3923), .A3(n2852), .ZN(n3922) );
  INV_X1 U3825 ( .A(n3924), .ZN(n3923) );
  NAND2_X1 U3826 ( .A1(n3889), .A2(n3887), .ZN(n3924) );
  NOR2_X1 U3827 ( .A1(n3887), .A2(n3889), .ZN(n3921) );
  NOR2_X1 U3828 ( .A1(n3925), .A2(n3926), .ZN(n3889) );
  NOR3_X1 U3829 ( .A1(n2679), .A2(n3927), .A3(n2852), .ZN(n3926) );
  NOR2_X1 U3830 ( .A1(n3883), .A2(n3885), .ZN(n3927) );
  INV_X1 U3831 ( .A(n3928), .ZN(n3925) );
  NAND2_X1 U3832 ( .A1(n3883), .A2(n3885), .ZN(n3928) );
  NAND2_X1 U3833 ( .A1(n3929), .A2(n3930), .ZN(n3885) );
  NAND2_X1 U3834 ( .A1(n3876), .A2(n3931), .ZN(n3930) );
  NAND2_X1 U3835 ( .A1(n3882), .A2(n3932), .ZN(n3931) );
  NAND2_X1 U3836 ( .A1(b_7_), .A2(a_6_), .ZN(n3932) );
  XNOR2_X1 U3837 ( .A(n3933), .B(n3934), .ZN(n3876) );
  XOR2_X1 U3838 ( .A(n3935), .B(n3936), .Z(n3934) );
  INV_X1 U3839 ( .A(n3879), .ZN(n3929) );
  NOR2_X1 U3840 ( .A1(n3882), .A2(n2854), .ZN(n3879) );
  NAND2_X1 U3841 ( .A1(n3937), .A2(n3938), .ZN(n3882) );
  NAND2_X1 U3842 ( .A1(n3873), .A2(n3939), .ZN(n3938) );
  NAND2_X1 U3843 ( .A1(n3875), .A2(n3874), .ZN(n3939) );
  XNOR2_X1 U3844 ( .A(n3940), .B(n3941), .ZN(n3873) );
  XNOR2_X1 U3845 ( .A(n3942), .B(n3943), .ZN(n3941) );
  NAND2_X1 U3846 ( .A1(b_6_), .A2(a_8_), .ZN(n3943) );
  INV_X1 U3847 ( .A(n3944), .ZN(n3937) );
  NOR2_X1 U3848 ( .A1(n3874), .A2(n3875), .ZN(n3944) );
  INV_X1 U3849 ( .A(n2826), .ZN(n3875) );
  NAND2_X1 U3850 ( .A1(b_7_), .A2(a_7_), .ZN(n2826) );
  NAND2_X1 U3851 ( .A1(n3945), .A2(n3946), .ZN(n3874) );
  NAND2_X1 U3852 ( .A1(n3871), .A2(n3947), .ZN(n3946) );
  INV_X1 U3853 ( .A(n3948), .ZN(n3947) );
  NOR2_X1 U3854 ( .A1(n3869), .A2(n3870), .ZN(n3948) );
  NOR2_X1 U3855 ( .A1(n2852), .A2(n2851), .ZN(n3871) );
  NAND2_X1 U3856 ( .A1(n3869), .A2(n3870), .ZN(n3945) );
  NAND2_X1 U3857 ( .A1(n3949), .A2(n3950), .ZN(n3870) );
  INV_X1 U3858 ( .A(n3951), .ZN(n3950) );
  NOR3_X1 U3859 ( .A1(n2577), .A2(n3952), .A3(n2852), .ZN(n3951) );
  NOR2_X1 U3860 ( .A1(n3821), .A2(n3823), .ZN(n3952) );
  NAND2_X1 U3861 ( .A1(n3821), .A2(n3823), .ZN(n3949) );
  NAND2_X1 U3862 ( .A1(n3866), .A2(n3953), .ZN(n3823) );
  NAND2_X1 U3863 ( .A1(n3865), .A2(n3867), .ZN(n3953) );
  NAND2_X1 U3864 ( .A1(n3954), .A2(n3955), .ZN(n3867) );
  NAND2_X1 U3865 ( .A1(b_7_), .A2(a_10_), .ZN(n3955) );
  INV_X1 U3866 ( .A(n3956), .ZN(n3954) );
  XNOR2_X1 U3867 ( .A(n3957), .B(n3958), .ZN(n3865) );
  NAND2_X1 U3868 ( .A1(n3959), .A2(n3960), .ZN(n3957) );
  NAND2_X1 U3869 ( .A1(a_10_), .A2(n3956), .ZN(n3866) );
  NAND2_X1 U3870 ( .A1(n3835), .A2(n3961), .ZN(n3956) );
  NAND2_X1 U3871 ( .A1(n3834), .A2(n3836), .ZN(n3961) );
  NAND2_X1 U3872 ( .A1(n3962), .A2(n3963), .ZN(n3836) );
  NAND2_X1 U3873 ( .A1(b_7_), .A2(a_11_), .ZN(n3963) );
  XNOR2_X1 U3874 ( .A(n3964), .B(n3965), .ZN(n3834) );
  XNOR2_X1 U3875 ( .A(n3966), .B(n3967), .ZN(n3964) );
  INV_X1 U3876 ( .A(n3968), .ZN(n3835) );
  NOR2_X1 U3877 ( .A1(n2846), .A2(n3962), .ZN(n3968) );
  NOR2_X1 U3878 ( .A1(n3969), .A2(n3970), .ZN(n3962) );
  INV_X1 U3879 ( .A(n3971), .ZN(n3970) );
  NAND2_X1 U3880 ( .A1(n3842), .A2(n3972), .ZN(n3971) );
  NAND2_X1 U3881 ( .A1(n3843), .A2(n3841), .ZN(n3972) );
  NOR2_X1 U3882 ( .A1(n2852), .A2(n2844), .ZN(n3842) );
  NOR2_X1 U3883 ( .A1(n3841), .A2(n3843), .ZN(n3969) );
  NOR2_X1 U3884 ( .A1(n3973), .A2(n3974), .ZN(n3843) );
  INV_X1 U3885 ( .A(n3975), .ZN(n3974) );
  NAND2_X1 U3886 ( .A1(n3860), .A2(n3976), .ZN(n3975) );
  NAND2_X1 U3887 ( .A1(n3977), .A2(n3862), .ZN(n3976) );
  NOR2_X1 U3888 ( .A1(n2852), .A2(n2842), .ZN(n3860) );
  NOR2_X1 U3889 ( .A1(n3862), .A2(n3977), .ZN(n3973) );
  INV_X1 U3890 ( .A(n3863), .ZN(n3977) );
  NAND2_X1 U3891 ( .A1(n3978), .A2(n3979), .ZN(n3863) );
  NAND2_X1 U3892 ( .A1(b_5_), .A2(n3980), .ZN(n3979) );
  NAND2_X1 U3893 ( .A1(n2426), .A2(n3981), .ZN(n3980) );
  NAND2_X1 U3894 ( .A1(a_15_), .A2(n2853), .ZN(n3981) );
  NAND2_X1 U3895 ( .A1(b_6_), .A2(n3982), .ZN(n3978) );
  NAND2_X1 U3896 ( .A1(n3049), .A2(n3983), .ZN(n3982) );
  NAND2_X1 U3897 ( .A1(a_14_), .A2(n2855), .ZN(n3983) );
  NAND3_X1 U3898 ( .A1(b_6_), .A2(b_7_), .A3(n2840), .ZN(n3862) );
  XOR2_X1 U3899 ( .A(n3984), .B(n3985), .Z(n3841) );
  XOR2_X1 U3900 ( .A(n3986), .B(n3987), .Z(n3985) );
  XNOR2_X1 U3901 ( .A(n3988), .B(n3989), .ZN(n3821) );
  NAND2_X1 U3902 ( .A1(n3990), .A2(n3991), .ZN(n3988) );
  XNOR2_X1 U3903 ( .A(n3992), .B(n3993), .ZN(n3869) );
  XOR2_X1 U3904 ( .A(n3994), .B(n3995), .Z(n3993) );
  NAND2_X1 U3905 ( .A1(b_6_), .A2(a_9_), .ZN(n3995) );
  XNOR2_X1 U3906 ( .A(n3996), .B(n3997), .ZN(n3883) );
  XOR2_X1 U3907 ( .A(n3998), .B(n3999), .Z(n3996) );
  XOR2_X1 U3908 ( .A(n4000), .B(n4001), .Z(n3887) );
  XNOR2_X1 U3909 ( .A(n4002), .B(n4003), .ZN(n4001) );
  XOR2_X1 U3910 ( .A(n4004), .B(n4005), .Z(n3892) );
  XNOR2_X1 U3911 ( .A(n4006), .B(n4007), .ZN(n4004) );
  XOR2_X1 U3912 ( .A(n4008), .B(n4009), .Z(n3895) );
  XNOR2_X1 U3913 ( .A(n4010), .B(n4011), .ZN(n4008) );
  XOR2_X1 U3914 ( .A(n4012), .B(n4013), .Z(n3786) );
  XNOR2_X1 U3915 ( .A(n4014), .B(n4015), .ZN(n4012) );
  XOR2_X1 U3916 ( .A(n4016), .B(n4017), .Z(n3900) );
  XNOR2_X1 U3917 ( .A(n4018), .B(n4019), .ZN(n4016) );
  NOR2_X1 U3918 ( .A1(n2790), .A2(n2853), .ZN(n4019) );
  XOR2_X1 U3919 ( .A(n4020), .B(n3780), .Z(n3903) );
  XOR2_X1 U3920 ( .A(n4021), .B(n4022), .Z(n3780) );
  NOR2_X1 U3921 ( .A1(n2865), .A2(n2853), .ZN(n4022) );
  XOR2_X1 U3922 ( .A(n2391), .B(n2390), .Z(n2381) );
  NAND3_X1 U3923 ( .A1(n2390), .A2(n2391), .A3(n2915), .ZN(n2386) );
  INV_X1 U3924 ( .A(n2389), .ZN(n2915) );
  NAND2_X1 U3925 ( .A1(n4023), .A2(n2913), .ZN(n2389) );
  NAND2_X1 U3926 ( .A1(n4024), .A2(n4025), .ZN(n4023) );
  XOR2_X1 U3927 ( .A(n4026), .B(n4027), .Z(n4024) );
  NAND2_X1 U3928 ( .A1(n4028), .A2(n4029), .ZN(n2391) );
  NAND3_X1 U3929 ( .A1(a_0_), .A2(n4030), .A3(b_6_), .ZN(n4029) );
  NAND2_X1 U3930 ( .A1(n4021), .A2(n4020), .ZN(n4030) );
  INV_X1 U3931 ( .A(n4031), .ZN(n4021) );
  NAND2_X1 U3932 ( .A1(n3779), .A2(n4031), .ZN(n4028) );
  NAND2_X1 U3933 ( .A1(n4032), .A2(n4033), .ZN(n4031) );
  NAND3_X1 U3934 ( .A1(a_1_), .A2(n4034), .A3(b_6_), .ZN(n4033) );
  NAND2_X1 U3935 ( .A1(n4017), .A2(n4018), .ZN(n4034) );
  INV_X1 U3936 ( .A(n4035), .ZN(n4032) );
  NOR2_X1 U3937 ( .A1(n4017), .A2(n4018), .ZN(n4035) );
  NOR2_X1 U3938 ( .A1(n4036), .A2(n4037), .ZN(n4018) );
  INV_X1 U3939 ( .A(n4038), .ZN(n4037) );
  NAND2_X1 U3940 ( .A1(n4015), .A2(n4039), .ZN(n4038) );
  NAND2_X1 U3941 ( .A1(n4014), .A2(n4013), .ZN(n4039) );
  NOR2_X1 U3942 ( .A1(n2853), .A2(n2860), .ZN(n4015) );
  NOR2_X1 U3943 ( .A1(n4013), .A2(n4014), .ZN(n4036) );
  NOR2_X1 U3944 ( .A1(n4040), .A2(n4041), .ZN(n4014) );
  INV_X1 U3945 ( .A(n4042), .ZN(n4041) );
  NAND2_X1 U3946 ( .A1(n4011), .A2(n4043), .ZN(n4042) );
  NAND2_X1 U3947 ( .A1(n4010), .A2(n4009), .ZN(n4043) );
  NOR2_X1 U3948 ( .A1(n2853), .A2(n2739), .ZN(n4011) );
  NOR2_X1 U3949 ( .A1(n4009), .A2(n4010), .ZN(n4040) );
  NOR2_X1 U3950 ( .A1(n4044), .A2(n4045), .ZN(n4010) );
  INV_X1 U3951 ( .A(n4046), .ZN(n4045) );
  NAND2_X1 U3952 ( .A1(n4007), .A2(n4047), .ZN(n4046) );
  NAND2_X1 U3953 ( .A1(n4006), .A2(n4005), .ZN(n4047) );
  NOR2_X1 U3954 ( .A1(n2853), .A2(n2857), .ZN(n4007) );
  NOR2_X1 U3955 ( .A1(n4005), .A2(n4006), .ZN(n4044) );
  NOR2_X1 U3956 ( .A1(n4048), .A2(n4049), .ZN(n4006) );
  INV_X1 U3957 ( .A(n4050), .ZN(n4049) );
  NAND2_X1 U3958 ( .A1(n4003), .A2(n4051), .ZN(n4050) );
  NAND2_X1 U3959 ( .A1(n4000), .A2(n4002), .ZN(n4051) );
  NOR2_X1 U3960 ( .A1(n2853), .A2(n2679), .ZN(n4003) );
  NOR2_X1 U3961 ( .A1(n4000), .A2(n4002), .ZN(n4048) );
  NAND2_X1 U3962 ( .A1(n4052), .A2(n4053), .ZN(n4002) );
  NAND2_X1 U3963 ( .A1(n3997), .A2(n4054), .ZN(n4053) );
  NAND2_X1 U3964 ( .A1(n3999), .A2(n3998), .ZN(n4054) );
  INV_X1 U3965 ( .A(n2653), .ZN(n3999) );
  XOR2_X1 U3966 ( .A(n4055), .B(n4056), .Z(n3997) );
  XOR2_X1 U3967 ( .A(n4057), .B(n4058), .Z(n4056) );
  NAND2_X1 U3968 ( .A1(b_5_), .A2(a_7_), .ZN(n4058) );
  NAND2_X1 U3969 ( .A1(n4059), .A2(n2653), .ZN(n4052) );
  NAND2_X1 U3970 ( .A1(b_6_), .A2(a_6_), .ZN(n2653) );
  INV_X1 U3971 ( .A(n3998), .ZN(n4059) );
  NAND2_X1 U3972 ( .A1(n4060), .A2(n4061), .ZN(n3998) );
  INV_X1 U3973 ( .A(n4062), .ZN(n4061) );
  NOR2_X1 U3974 ( .A1(n3936), .A2(n4063), .ZN(n4062) );
  NOR2_X1 U3975 ( .A1(n3933), .A2(n3935), .ZN(n4063) );
  NAND2_X1 U3976 ( .A1(b_6_), .A2(a_7_), .ZN(n3936) );
  NAND2_X1 U3977 ( .A1(n3933), .A2(n3935), .ZN(n4060) );
  NAND2_X1 U3978 ( .A1(n4064), .A2(n4065), .ZN(n3935) );
  NAND3_X1 U3979 ( .A1(a_8_), .A2(n4066), .A3(b_6_), .ZN(n4065) );
  NAND2_X1 U3980 ( .A1(n3942), .A2(n3940), .ZN(n4066) );
  INV_X1 U3981 ( .A(n4067), .ZN(n4064) );
  NOR2_X1 U3982 ( .A1(n3940), .A2(n3942), .ZN(n4067) );
  NOR2_X1 U3983 ( .A1(n4068), .A2(n4069), .ZN(n3942) );
  NOR3_X1 U3984 ( .A1(n2577), .A2(n4070), .A3(n2853), .ZN(n4069) );
  NOR2_X1 U3985 ( .A1(n3994), .A2(n3992), .ZN(n4070) );
  INV_X1 U3986 ( .A(n4071), .ZN(n4068) );
  NAND2_X1 U3987 ( .A1(n3992), .A2(n3994), .ZN(n4071) );
  NAND2_X1 U3988 ( .A1(n3990), .A2(n4072), .ZN(n3994) );
  NAND2_X1 U3989 ( .A1(n3989), .A2(n3991), .ZN(n4072) );
  NAND2_X1 U3990 ( .A1(n4073), .A2(n4074), .ZN(n3991) );
  NAND2_X1 U3991 ( .A1(b_6_), .A2(a_10_), .ZN(n4074) );
  INV_X1 U3992 ( .A(n4075), .ZN(n4073) );
  XNOR2_X1 U3993 ( .A(n4076), .B(n4077), .ZN(n3989) );
  NAND2_X1 U3994 ( .A1(n4078), .A2(n4079), .ZN(n4076) );
  NAND2_X1 U3995 ( .A1(a_10_), .A2(n4075), .ZN(n3990) );
  NAND2_X1 U3996 ( .A1(n3959), .A2(n4080), .ZN(n4075) );
  NAND2_X1 U3997 ( .A1(n3958), .A2(n3960), .ZN(n4080) );
  NAND2_X1 U3998 ( .A1(n4081), .A2(n4082), .ZN(n3960) );
  NAND2_X1 U3999 ( .A1(b_6_), .A2(a_11_), .ZN(n4082) );
  XNOR2_X1 U4000 ( .A(n4083), .B(n4084), .ZN(n3958) );
  XNOR2_X1 U4001 ( .A(n4085), .B(n4086), .ZN(n4083) );
  INV_X1 U4002 ( .A(n4087), .ZN(n3959) );
  NOR2_X1 U4003 ( .A1(n2846), .A2(n4081), .ZN(n4087) );
  NOR2_X1 U4004 ( .A1(n4088), .A2(n4089), .ZN(n4081) );
  INV_X1 U4005 ( .A(n4090), .ZN(n4089) );
  NAND2_X1 U4006 ( .A1(n3966), .A2(n4091), .ZN(n4090) );
  NAND2_X1 U4007 ( .A1(n3967), .A2(n3965), .ZN(n4091) );
  NOR2_X1 U4008 ( .A1(n2853), .A2(n2844), .ZN(n3966) );
  NOR2_X1 U4009 ( .A1(n3965), .A2(n3967), .ZN(n4088) );
  NOR2_X1 U4010 ( .A1(n4092), .A2(n4093), .ZN(n3967) );
  INV_X1 U4011 ( .A(n4094), .ZN(n4093) );
  NAND2_X1 U4012 ( .A1(n3984), .A2(n4095), .ZN(n4094) );
  NAND2_X1 U4013 ( .A1(n4096), .A2(n3986), .ZN(n4095) );
  NOR2_X1 U4014 ( .A1(n2853), .A2(n2842), .ZN(n3984) );
  NOR2_X1 U4015 ( .A1(n3986), .A2(n4096), .ZN(n4092) );
  INV_X1 U4016 ( .A(n3987), .ZN(n4096) );
  NAND2_X1 U4017 ( .A1(n4097), .A2(n4098), .ZN(n3987) );
  NAND2_X1 U4018 ( .A1(b_4_), .A2(n4099), .ZN(n4098) );
  NAND2_X1 U4019 ( .A1(n2426), .A2(n4100), .ZN(n4099) );
  NAND2_X1 U4020 ( .A1(a_15_), .A2(n2855), .ZN(n4100) );
  NAND2_X1 U4021 ( .A1(b_5_), .A2(n4101), .ZN(n4097) );
  NAND2_X1 U4022 ( .A1(n3049), .A2(n4102), .ZN(n4101) );
  NAND2_X1 U4023 ( .A1(a_14_), .A2(n2856), .ZN(n4102) );
  NAND3_X1 U4024 ( .A1(b_5_), .A2(b_6_), .A3(n2840), .ZN(n3986) );
  XOR2_X1 U4025 ( .A(n4103), .B(n4104), .Z(n3965) );
  XOR2_X1 U4026 ( .A(n4105), .B(n4106), .Z(n4104) );
  XNOR2_X1 U4027 ( .A(n4107), .B(n4108), .ZN(n3992) );
  NAND2_X1 U4028 ( .A1(n4109), .A2(n4110), .ZN(n4107) );
  XNOR2_X1 U4029 ( .A(n4111), .B(n4112), .ZN(n3940) );
  XOR2_X1 U4030 ( .A(n4113), .B(n4114), .Z(n4111) );
  NOR2_X1 U4031 ( .A1(n2577), .A2(n2855), .ZN(n4114) );
  XNOR2_X1 U4032 ( .A(n4115), .B(n4116), .ZN(n3933) );
  XOR2_X1 U4033 ( .A(n4117), .B(n4118), .Z(n4116) );
  NAND2_X1 U4034 ( .A1(b_5_), .A2(a_8_), .ZN(n4118) );
  XOR2_X1 U4035 ( .A(n4119), .B(n4120), .Z(n4000) );
  XOR2_X1 U4036 ( .A(n4121), .B(n4122), .Z(n4120) );
  NAND2_X1 U4037 ( .A1(b_5_), .A2(a_6_), .ZN(n4122) );
  XNOR2_X1 U4038 ( .A(n4123), .B(n4124), .ZN(n4005) );
  XOR2_X1 U4039 ( .A(n4125), .B(n2822), .Z(n4123) );
  XNOR2_X1 U4040 ( .A(n4126), .B(n4127), .ZN(n4009) );
  XOR2_X1 U4041 ( .A(n4128), .B(n4129), .Z(n4126) );
  NOR2_X1 U4042 ( .A1(n2857), .A2(n2855), .ZN(n4129) );
  XNOR2_X1 U4043 ( .A(n4130), .B(n4131), .ZN(n4013) );
  XOR2_X1 U4044 ( .A(n4132), .B(n4133), .Z(n4130) );
  NOR2_X1 U4045 ( .A1(n2739), .A2(n2855), .ZN(n4133) );
  XNOR2_X1 U4046 ( .A(n4134), .B(n4135), .ZN(n4017) );
  XOR2_X1 U4047 ( .A(n4136), .B(n4137), .Z(n4134) );
  NOR2_X1 U4048 ( .A1(n2860), .A2(n2855), .ZN(n4137) );
  INV_X1 U4049 ( .A(n4020), .ZN(n3779) );
  XNOR2_X1 U4050 ( .A(n4138), .B(n4139), .ZN(n4020) );
  XNOR2_X1 U4051 ( .A(n4140), .B(n4141), .ZN(n4139) );
  NAND2_X1 U4052 ( .A1(b_5_), .A2(a_1_), .ZN(n4141) );
  XNOR2_X1 U4053 ( .A(n4142), .B(n4143), .ZN(n2390) );
  XNOR2_X1 U4054 ( .A(n4144), .B(n4145), .ZN(n4142) );
  NOR2_X1 U4055 ( .A1(n2865), .A2(n2855), .ZN(n4145) );
  NAND2_X1 U4056 ( .A1(n4146), .A2(n4147), .ZN(n2913) );
  INV_X1 U4057 ( .A(n4025), .ZN(n4147) );
  NOR2_X1 U4058 ( .A1(n4148), .A2(n4149), .ZN(n4025) );
  INV_X1 U4059 ( .A(n4150), .ZN(n4149) );
  NAND3_X1 U4060 ( .A1(a_0_), .A2(n4151), .A3(b_5_), .ZN(n4150) );
  NAND2_X1 U4061 ( .A1(n4144), .A2(n4143), .ZN(n4151) );
  NOR2_X1 U4062 ( .A1(n4143), .A2(n4144), .ZN(n4148) );
  NOR2_X1 U4063 ( .A1(n4152), .A2(n4153), .ZN(n4144) );
  NOR3_X1 U4064 ( .A1(n2790), .A2(n4154), .A3(n2855), .ZN(n4153) );
  INV_X1 U4065 ( .A(n4155), .ZN(n4154) );
  NAND2_X1 U4066 ( .A1(n4138), .A2(n4140), .ZN(n4155) );
  NOR2_X1 U4067 ( .A1(n4138), .A2(n4140), .ZN(n4152) );
  NOR2_X1 U4068 ( .A1(n4156), .A2(n4157), .ZN(n4140) );
  NOR3_X1 U4069 ( .A1(n2860), .A2(n4158), .A3(n2855), .ZN(n4157) );
  NOR2_X1 U4070 ( .A1(n4136), .A2(n4135), .ZN(n4158) );
  INV_X1 U4071 ( .A(n4159), .ZN(n4156) );
  NAND2_X1 U4072 ( .A1(n4135), .A2(n4136), .ZN(n4159) );
  NAND2_X1 U4073 ( .A1(n4160), .A2(n4161), .ZN(n4136) );
  INV_X1 U4074 ( .A(n4162), .ZN(n4161) );
  NOR3_X1 U4075 ( .A1(n2739), .A2(n4163), .A3(n2855), .ZN(n4162) );
  NOR2_X1 U4076 ( .A1(n4131), .A2(n4132), .ZN(n4163) );
  NAND2_X1 U4077 ( .A1(n4131), .A2(n4132), .ZN(n4160) );
  NAND2_X1 U4078 ( .A1(n4164), .A2(n4165), .ZN(n4132) );
  NAND3_X1 U4079 ( .A1(a_4_), .A2(n4166), .A3(b_5_), .ZN(n4165) );
  INV_X1 U4080 ( .A(n4167), .ZN(n4166) );
  NOR2_X1 U4081 ( .A1(n4127), .A2(n4128), .ZN(n4167) );
  NAND2_X1 U4082 ( .A1(n4127), .A2(n4128), .ZN(n4164) );
  NAND2_X1 U4083 ( .A1(n4168), .A2(n4169), .ZN(n4128) );
  NAND2_X1 U4084 ( .A1(n4124), .A2(n4170), .ZN(n4169) );
  NAND2_X1 U4085 ( .A1(n4125), .A2(n2822), .ZN(n4170) );
  XOR2_X1 U4086 ( .A(n4171), .B(n4172), .Z(n4124) );
  XOR2_X1 U4087 ( .A(n4173), .B(n4174), .Z(n4172) );
  INV_X1 U4088 ( .A(n4175), .ZN(n4168) );
  NOR2_X1 U4089 ( .A1(n2822), .A2(n4125), .ZN(n4175) );
  NOR2_X1 U4090 ( .A1(n4176), .A2(n4177), .ZN(n4125) );
  NOR3_X1 U4091 ( .A1(n2854), .A2(n4178), .A3(n2855), .ZN(n4177) );
  NOR2_X1 U4092 ( .A1(n4119), .A2(n4121), .ZN(n4178) );
  INV_X1 U4093 ( .A(n4179), .ZN(n4176) );
  NAND2_X1 U4094 ( .A1(n4119), .A2(n4121), .ZN(n4179) );
  NAND2_X1 U4095 ( .A1(n4180), .A2(n4181), .ZN(n4121) );
  INV_X1 U4096 ( .A(n4182), .ZN(n4181) );
  NOR3_X1 U4097 ( .A1(n2628), .A2(n4183), .A3(n2855), .ZN(n4182) );
  NOR2_X1 U4098 ( .A1(n4055), .A2(n4057), .ZN(n4183) );
  NAND2_X1 U4099 ( .A1(n4055), .A2(n4057), .ZN(n4180) );
  NAND2_X1 U4100 ( .A1(n4184), .A2(n4185), .ZN(n4057) );
  NAND3_X1 U4101 ( .A1(a_8_), .A2(n4186), .A3(b_5_), .ZN(n4185) );
  INV_X1 U4102 ( .A(n4187), .ZN(n4186) );
  NOR2_X1 U4103 ( .A1(n4117), .A2(n4115), .ZN(n4187) );
  NAND2_X1 U4104 ( .A1(n4115), .A2(n4117), .ZN(n4184) );
  NAND2_X1 U4105 ( .A1(n4188), .A2(n4189), .ZN(n4117) );
  INV_X1 U4106 ( .A(n4190), .ZN(n4189) );
  NOR3_X1 U4107 ( .A1(n2577), .A2(n4191), .A3(n2855), .ZN(n4190) );
  NOR2_X1 U4108 ( .A1(n4112), .A2(n4113), .ZN(n4191) );
  NAND2_X1 U4109 ( .A1(n4112), .A2(n4113), .ZN(n4188) );
  NAND2_X1 U4110 ( .A1(n4109), .A2(n4192), .ZN(n4113) );
  NAND2_X1 U4111 ( .A1(n4108), .A2(n4110), .ZN(n4192) );
  NAND2_X1 U4112 ( .A1(n4193), .A2(n4194), .ZN(n4110) );
  NAND2_X1 U4113 ( .A1(b_5_), .A2(a_10_), .ZN(n4194) );
  INV_X1 U4114 ( .A(n4195), .ZN(n4193) );
  XOR2_X1 U4115 ( .A(n4196), .B(n4197), .Z(n4108) );
  XOR2_X1 U4116 ( .A(n4198), .B(n4199), .Z(n4196) );
  NAND2_X1 U4117 ( .A1(a_10_), .A2(n4195), .ZN(n4109) );
  NAND2_X1 U4118 ( .A1(n4078), .A2(n4200), .ZN(n4195) );
  NAND2_X1 U4119 ( .A1(n4077), .A2(n4079), .ZN(n4200) );
  NAND2_X1 U4120 ( .A1(n4201), .A2(n4202), .ZN(n4079) );
  NAND2_X1 U4121 ( .A1(b_5_), .A2(a_11_), .ZN(n4202) );
  XNOR2_X1 U4122 ( .A(n4203), .B(n4204), .ZN(n4077) );
  XNOR2_X1 U4123 ( .A(n4205), .B(n4206), .ZN(n4203) );
  INV_X1 U4124 ( .A(n4207), .ZN(n4078) );
  NOR2_X1 U4125 ( .A1(n2846), .A2(n4201), .ZN(n4207) );
  NOR2_X1 U4126 ( .A1(n4208), .A2(n4209), .ZN(n4201) );
  INV_X1 U4127 ( .A(n4210), .ZN(n4209) );
  NAND2_X1 U4128 ( .A1(n4085), .A2(n4211), .ZN(n4210) );
  NAND2_X1 U4129 ( .A1(n4086), .A2(n4084), .ZN(n4211) );
  NOR2_X1 U4130 ( .A1(n2855), .A2(n2844), .ZN(n4085) );
  NOR2_X1 U4131 ( .A1(n4084), .A2(n4086), .ZN(n4208) );
  NOR2_X1 U4132 ( .A1(n4212), .A2(n4213), .ZN(n4086) );
  INV_X1 U4133 ( .A(n4214), .ZN(n4213) );
  NAND2_X1 U4134 ( .A1(n4103), .A2(n4215), .ZN(n4214) );
  NAND2_X1 U4135 ( .A1(n4216), .A2(n4105), .ZN(n4215) );
  NOR2_X1 U4136 ( .A1(n2855), .A2(n2842), .ZN(n4103) );
  NOR2_X1 U4137 ( .A1(n4105), .A2(n4216), .ZN(n4212) );
  INV_X1 U4138 ( .A(n4106), .ZN(n4216) );
  NAND2_X1 U4139 ( .A1(n4217), .A2(n4218), .ZN(n4106) );
  NAND2_X1 U4140 ( .A1(b_3_), .A2(n4219), .ZN(n4218) );
  NAND2_X1 U4141 ( .A1(n2426), .A2(n4220), .ZN(n4219) );
  NAND2_X1 U4142 ( .A1(a_15_), .A2(n2856), .ZN(n4220) );
  NAND2_X1 U4143 ( .A1(b_4_), .A2(n4221), .ZN(n4217) );
  NAND2_X1 U4144 ( .A1(n3049), .A2(n4222), .ZN(n4221) );
  NAND2_X1 U4145 ( .A1(a_14_), .A2(n2858), .ZN(n4222) );
  NAND3_X1 U4146 ( .A1(b_4_), .A2(b_5_), .A3(n2840), .ZN(n4105) );
  XOR2_X1 U4147 ( .A(n4223), .B(n4224), .Z(n4084) );
  XOR2_X1 U4148 ( .A(n4225), .B(n4226), .Z(n4224) );
  XNOR2_X1 U4149 ( .A(n4227), .B(n4228), .ZN(n4112) );
  XOR2_X1 U4150 ( .A(n4229), .B(n4230), .Z(n4227) );
  XNOR2_X1 U4151 ( .A(n4231), .B(n4232), .ZN(n4115) );
  XNOR2_X1 U4152 ( .A(n4233), .B(n4234), .ZN(n4231) );
  XNOR2_X1 U4153 ( .A(n4235), .B(n4236), .ZN(n4055) );
  XNOR2_X1 U4154 ( .A(n4237), .B(n4238), .ZN(n4235) );
  XNOR2_X1 U4155 ( .A(n4239), .B(n4240), .ZN(n4119) );
  XNOR2_X1 U4156 ( .A(n4241), .B(n4242), .ZN(n4239) );
  NAND2_X1 U4157 ( .A1(b_5_), .A2(a_5_), .ZN(n2822) );
  XOR2_X1 U4158 ( .A(n4243), .B(n4244), .Z(n4127) );
  XOR2_X1 U4159 ( .A(n4245), .B(n4246), .Z(n4243) );
  XOR2_X1 U4160 ( .A(n4247), .B(n4248), .Z(n4131) );
  XOR2_X1 U4161 ( .A(n4249), .B(n4250), .Z(n4248) );
  XNOR2_X1 U4162 ( .A(n4251), .B(n4252), .ZN(n4135) );
  XNOR2_X1 U4163 ( .A(n4253), .B(n4254), .ZN(n4252) );
  XNOR2_X1 U4164 ( .A(n4255), .B(n4256), .ZN(n4138) );
  XOR2_X1 U4165 ( .A(n4257), .B(n4258), .Z(n4256) );
  XOR2_X1 U4166 ( .A(n4259), .B(n4260), .Z(n4143) );
  XNOR2_X1 U4167 ( .A(n4261), .B(n4262), .ZN(n4259) );
  NOR2_X1 U4168 ( .A1(n2790), .A2(n2856), .ZN(n4262) );
  XOR2_X1 U4169 ( .A(n4263), .B(n4026), .Z(n4146) );
  XNOR2_X1 U4170 ( .A(n4264), .B(n4265), .ZN(n4026) );
  NOR2_X1 U4171 ( .A1(n2865), .A2(n2856), .ZN(n4265) );
  XOR2_X1 U4172 ( .A(n2405), .B(n2404), .Z(n2395) );
  NAND3_X1 U4173 ( .A1(n2404), .A2(n2405), .A3(n2912), .ZN(n2400) );
  INV_X1 U4174 ( .A(n2403), .ZN(n2912) );
  NAND2_X1 U4175 ( .A1(n4266), .A2(n2910), .ZN(n2403) );
  NAND2_X1 U4176 ( .A1(n4267), .A2(n4268), .ZN(n4266) );
  XOR2_X1 U4177 ( .A(n4269), .B(n4270), .Z(n4268) );
  INV_X1 U4178 ( .A(n4271), .ZN(n4267) );
  NAND2_X1 U4179 ( .A1(n4272), .A2(n4273), .ZN(n2405) );
  NAND3_X1 U4180 ( .A1(a_0_), .A2(n4274), .A3(b_4_), .ZN(n4273) );
  NAND2_X1 U4181 ( .A1(n4275), .A2(n4263), .ZN(n4274) );
  INV_X1 U4182 ( .A(n4264), .ZN(n4275) );
  NAND2_X1 U4183 ( .A1(n4027), .A2(n4264), .ZN(n4272) );
  NAND2_X1 U4184 ( .A1(n4276), .A2(n4277), .ZN(n4264) );
  NAND3_X1 U4185 ( .A1(a_1_), .A2(n4278), .A3(b_4_), .ZN(n4277) );
  NAND2_X1 U4186 ( .A1(n4260), .A2(n4261), .ZN(n4278) );
  INV_X1 U4187 ( .A(n4279), .ZN(n4276) );
  NOR2_X1 U4188 ( .A1(n4260), .A2(n4261), .ZN(n4279) );
  NOR2_X1 U4189 ( .A1(n4280), .A2(n4281), .ZN(n4261) );
  INV_X1 U4190 ( .A(n4282), .ZN(n4281) );
  NAND2_X1 U4191 ( .A1(n4258), .A2(n4283), .ZN(n4282) );
  NAND2_X1 U4192 ( .A1(n4257), .A2(n4255), .ZN(n4283) );
  NOR2_X1 U4193 ( .A1(n2856), .A2(n2860), .ZN(n4258) );
  NOR2_X1 U4194 ( .A1(n4255), .A2(n4257), .ZN(n4280) );
  NOR2_X1 U4195 ( .A1(n4284), .A2(n4285), .ZN(n4257) );
  INV_X1 U4196 ( .A(n4286), .ZN(n4285) );
  NAND2_X1 U4197 ( .A1(n4254), .A2(n4287), .ZN(n4286) );
  NAND2_X1 U4198 ( .A1(n4251), .A2(n4253), .ZN(n4287) );
  NOR2_X1 U4199 ( .A1(n2856), .A2(n2739), .ZN(n4254) );
  NOR2_X1 U4200 ( .A1(n4251), .A2(n4253), .ZN(n4284) );
  NAND2_X1 U4201 ( .A1(n4288), .A2(n4289), .ZN(n4253) );
  NAND2_X1 U4202 ( .A1(n4247), .A2(n4290), .ZN(n4289) );
  NAND2_X1 U4203 ( .A1(n4250), .A2(n4291), .ZN(n4290) );
  XNOR2_X1 U4204 ( .A(n4292), .B(n4293), .ZN(n4247) );
  XNOR2_X1 U4205 ( .A(n4294), .B(n4295), .ZN(n4293) );
  NAND2_X1 U4206 ( .A1(b_3_), .A2(a_5_), .ZN(n4295) );
  NAND2_X1 U4207 ( .A1(n4249), .A2(n2704), .ZN(n4288) );
  INV_X1 U4208 ( .A(n4250), .ZN(n2704) );
  NOR2_X1 U4209 ( .A1(n2856), .A2(n2857), .ZN(n4250) );
  INV_X1 U4210 ( .A(n4291), .ZN(n4249) );
  NAND2_X1 U4211 ( .A1(n4296), .A2(n4297), .ZN(n4291) );
  NAND2_X1 U4212 ( .A1(n4246), .A2(n4298), .ZN(n4297) );
  INV_X1 U4213 ( .A(n4299), .ZN(n4298) );
  NOR2_X1 U4214 ( .A1(n4245), .A2(n4244), .ZN(n4299) );
  NOR2_X1 U4215 ( .A1(n2856), .A2(n2679), .ZN(n4246) );
  NAND2_X1 U4216 ( .A1(n4244), .A2(n4245), .ZN(n4296) );
  NAND2_X1 U4217 ( .A1(n4300), .A2(n4301), .ZN(n4245) );
  NAND2_X1 U4218 ( .A1(n4174), .A2(n4302), .ZN(n4301) );
  NAND2_X1 U4219 ( .A1(n4173), .A2(n4171), .ZN(n4302) );
  INV_X1 U4220 ( .A(n4303), .ZN(n4171) );
  INV_X1 U4221 ( .A(n4304), .ZN(n4173) );
  NOR2_X1 U4222 ( .A1(n2856), .A2(n2854), .ZN(n4174) );
  NAND2_X1 U4223 ( .A1(n4303), .A2(n4304), .ZN(n4300) );
  NAND2_X1 U4224 ( .A1(n4305), .A2(n4306), .ZN(n4304) );
  NAND2_X1 U4225 ( .A1(n4242), .A2(n4307), .ZN(n4306) );
  NAND2_X1 U4226 ( .A1(n4241), .A2(n4240), .ZN(n4307) );
  NOR2_X1 U4227 ( .A1(n2856), .A2(n2628), .ZN(n4242) );
  INV_X1 U4228 ( .A(n4308), .ZN(n4305) );
  NOR2_X1 U4229 ( .A1(n4240), .A2(n4241), .ZN(n4308) );
  NOR2_X1 U4230 ( .A1(n4309), .A2(n4310), .ZN(n4241) );
  INV_X1 U4231 ( .A(n4311), .ZN(n4310) );
  NAND2_X1 U4232 ( .A1(n4238), .A2(n4312), .ZN(n4311) );
  NAND2_X1 U4233 ( .A1(n4237), .A2(n4236), .ZN(n4312) );
  NOR2_X1 U4234 ( .A1(n2856), .A2(n2851), .ZN(n4238) );
  NOR2_X1 U4235 ( .A1(n4236), .A2(n4237), .ZN(n4309) );
  NOR2_X1 U4236 ( .A1(n4313), .A2(n4314), .ZN(n4237) );
  INV_X1 U4237 ( .A(n4315), .ZN(n4314) );
  NAND2_X1 U4238 ( .A1(n4233), .A2(n4316), .ZN(n4315) );
  NAND2_X1 U4239 ( .A1(n4232), .A2(n4234), .ZN(n4316) );
  NOR2_X1 U4240 ( .A1(n2856), .A2(n2577), .ZN(n4233) );
  NOR2_X1 U4241 ( .A1(n4232), .A2(n4234), .ZN(n4313) );
  NOR2_X1 U4242 ( .A1(n4317), .A2(n4318), .ZN(n4234) );
  INV_X1 U4243 ( .A(n4319), .ZN(n4318) );
  NAND2_X1 U4244 ( .A1(n4230), .A2(n4320), .ZN(n4319) );
  NAND2_X1 U4245 ( .A1(n4321), .A2(n4228), .ZN(n4320) );
  NOR2_X1 U4246 ( .A1(n2856), .A2(n2849), .ZN(n4230) );
  NOR2_X1 U4247 ( .A1(n4228), .A2(n4321), .ZN(n4317) );
  INV_X1 U4248 ( .A(n4229), .ZN(n4321) );
  NAND2_X1 U4249 ( .A1(n4322), .A2(n4323), .ZN(n4229) );
  NAND2_X1 U4250 ( .A1(n4199), .A2(n4324), .ZN(n4323) );
  NAND2_X1 U4251 ( .A1(n4325), .A2(n4326), .ZN(n4324) );
  INV_X1 U4252 ( .A(n4198), .ZN(n4326) );
  INV_X1 U4253 ( .A(n4197), .ZN(n4325) );
  NOR2_X1 U4254 ( .A1(n2856), .A2(n2846), .ZN(n4199) );
  NAND2_X1 U4255 ( .A1(n4197), .A2(n4198), .ZN(n4322) );
  NAND2_X1 U4256 ( .A1(n4327), .A2(n4328), .ZN(n4198) );
  NAND2_X1 U4257 ( .A1(n4205), .A2(n4329), .ZN(n4328) );
  NAND2_X1 U4258 ( .A1(n4206), .A2(n4204), .ZN(n4329) );
  NOR2_X1 U4259 ( .A1(n2856), .A2(n2844), .ZN(n4205) );
  INV_X1 U4260 ( .A(n4330), .ZN(n4327) );
  NOR2_X1 U4261 ( .A1(n4204), .A2(n4206), .ZN(n4330) );
  NOR2_X1 U4262 ( .A1(n4331), .A2(n4332), .ZN(n4206) );
  INV_X1 U4263 ( .A(n4333), .ZN(n4332) );
  NAND2_X1 U4264 ( .A1(n4223), .A2(n4334), .ZN(n4333) );
  NAND2_X1 U4265 ( .A1(n4335), .A2(n4225), .ZN(n4334) );
  NOR2_X1 U4266 ( .A1(n2856), .A2(n2842), .ZN(n4223) );
  NOR2_X1 U4267 ( .A1(n4225), .A2(n4335), .ZN(n4331) );
  INV_X1 U4268 ( .A(n4226), .ZN(n4335) );
  NAND2_X1 U4269 ( .A1(n4336), .A2(n4337), .ZN(n4226) );
  NAND2_X1 U4270 ( .A1(b_2_), .A2(n4338), .ZN(n4337) );
  NAND2_X1 U4271 ( .A1(n2426), .A2(n4339), .ZN(n4338) );
  NAND2_X1 U4272 ( .A1(a_15_), .A2(n2858), .ZN(n4339) );
  NAND2_X1 U4273 ( .A1(b_3_), .A2(n4340), .ZN(n4336) );
  NAND2_X1 U4274 ( .A1(n3049), .A2(n4341), .ZN(n4340) );
  NAND2_X1 U4275 ( .A1(a_14_), .A2(n2859), .ZN(n4341) );
  NAND3_X1 U4276 ( .A1(b_3_), .A2(b_4_), .A3(n2840), .ZN(n4225) );
  XOR2_X1 U4277 ( .A(n4342), .B(n4343), .Z(n4204) );
  XOR2_X1 U4278 ( .A(n4344), .B(n4345), .Z(n4343) );
  XNOR2_X1 U4279 ( .A(n4346), .B(n4347), .ZN(n4197) );
  XNOR2_X1 U4280 ( .A(n4348), .B(n4349), .ZN(n4346) );
  XOR2_X1 U4281 ( .A(n4350), .B(n4351), .Z(n4228) );
  NAND2_X1 U4282 ( .A1(n4352), .A2(n4353), .ZN(n4350) );
  XOR2_X1 U4283 ( .A(n4354), .B(n4355), .Z(n4232) );
  NAND2_X1 U4284 ( .A1(n4356), .A2(n4357), .ZN(n4354) );
  XNOR2_X1 U4285 ( .A(n4358), .B(n4359), .ZN(n4236) );
  XOR2_X1 U4286 ( .A(n4360), .B(n4361), .Z(n4358) );
  NOR2_X1 U4287 ( .A1(n2577), .A2(n2858), .ZN(n4361) );
  XNOR2_X1 U4288 ( .A(n4362), .B(n4363), .ZN(n4240) );
  XOR2_X1 U4289 ( .A(n4364), .B(n4365), .Z(n4362) );
  NOR2_X1 U4290 ( .A1(n2851), .A2(n2858), .ZN(n4365) );
  XNOR2_X1 U4291 ( .A(n4366), .B(n4367), .ZN(n4303) );
  XOR2_X1 U4292 ( .A(n4368), .B(n4369), .Z(n4367) );
  NAND2_X1 U4293 ( .A1(b_3_), .A2(a_7_), .ZN(n4369) );
  XNOR2_X1 U4294 ( .A(n4370), .B(n4371), .ZN(n4244) );
  XNOR2_X1 U4295 ( .A(n4372), .B(n4373), .ZN(n4370) );
  NOR2_X1 U4296 ( .A1(n2854), .A2(n2858), .ZN(n4373) );
  XOR2_X1 U4297 ( .A(n4374), .B(n4375), .Z(n4251) );
  XNOR2_X1 U4298 ( .A(n4376), .B(n4377), .ZN(n4374) );
  NOR2_X1 U4299 ( .A1(n2857), .A2(n2858), .ZN(n4377) );
  XNOR2_X1 U4300 ( .A(n4378), .B(n4379), .ZN(n4255) );
  XNOR2_X1 U4301 ( .A(n4380), .B(n2818), .ZN(n4379) );
  XNOR2_X1 U4302 ( .A(n4381), .B(n4382), .ZN(n4260) );
  XOR2_X1 U4303 ( .A(n4383), .B(n4384), .Z(n4381) );
  NOR2_X1 U4304 ( .A1(n2860), .A2(n2858), .ZN(n4384) );
  INV_X1 U4305 ( .A(n4263), .ZN(n4027) );
  XNOR2_X1 U4306 ( .A(n4385), .B(n4386), .ZN(n4263) );
  XNOR2_X1 U4307 ( .A(n4387), .B(n4388), .ZN(n4386) );
  NAND2_X1 U4308 ( .A1(b_3_), .A2(a_1_), .ZN(n4388) );
  XNOR2_X1 U4309 ( .A(n4389), .B(n4390), .ZN(n2404) );
  XOR2_X1 U4310 ( .A(n4391), .B(n4392), .Z(n4389) );
  NAND2_X1 U4311 ( .A1(b_3_), .A2(a_0_), .ZN(n4391) );
  NAND2_X1 U4312 ( .A1(n4393), .A2(n4271), .ZN(n2910) );
  NAND2_X1 U4313 ( .A1(n4394), .A2(n4395), .ZN(n4271) );
  NAND3_X1 U4314 ( .A1(a_0_), .A2(n4396), .A3(b_3_), .ZN(n4395) );
  NAND2_X1 U4315 ( .A1(n4390), .A2(n4392), .ZN(n4396) );
  INV_X1 U4316 ( .A(n4397), .ZN(n4394) );
  NOR2_X1 U4317 ( .A1(n4390), .A2(n4392), .ZN(n4397) );
  NOR2_X1 U4318 ( .A1(n4398), .A2(n4399), .ZN(n4392) );
  NOR3_X1 U4319 ( .A1(n2790), .A2(n4400), .A3(n2858), .ZN(n4399) );
  INV_X1 U4320 ( .A(n4401), .ZN(n4400) );
  NAND2_X1 U4321 ( .A1(n4385), .A2(n4387), .ZN(n4401) );
  NOR2_X1 U4322 ( .A1(n4385), .A2(n4387), .ZN(n4398) );
  NOR2_X1 U4323 ( .A1(n4402), .A2(n4403), .ZN(n4387) );
  INV_X1 U4324 ( .A(n4404), .ZN(n4403) );
  NAND3_X1 U4325 ( .A1(a_2_), .A2(n4405), .A3(b_3_), .ZN(n4404) );
  NAND2_X1 U4326 ( .A1(n4382), .A2(n4383), .ZN(n4405) );
  NOR2_X1 U4327 ( .A1(n4383), .A2(n4382), .ZN(n4402) );
  XNOR2_X1 U4328 ( .A(n4406), .B(n4407), .ZN(n4382) );
  XOR2_X1 U4329 ( .A(n4408), .B(n4409), .Z(n4406) );
  NAND2_X1 U4330 ( .A1(n4410), .A2(n4411), .ZN(n4383) );
  NAND2_X1 U4331 ( .A1(n4378), .A2(n4412), .ZN(n4411) );
  INV_X1 U4332 ( .A(n4413), .ZN(n4412) );
  NOR2_X1 U4333 ( .A1(n2818), .A2(n4380), .ZN(n4413) );
  XNOR2_X1 U4334 ( .A(n4414), .B(n4415), .ZN(n4378) );
  XOR2_X1 U4335 ( .A(n4416), .B(n4417), .Z(n4414) );
  NAND2_X1 U4336 ( .A1(n4380), .A2(n2818), .ZN(n4410) );
  NAND2_X1 U4337 ( .A1(b_3_), .A2(a_3_), .ZN(n2818) );
  NOR2_X1 U4338 ( .A1(n4418), .A2(n4419), .ZN(n4380) );
  NOR3_X1 U4339 ( .A1(n2857), .A2(n4420), .A3(n2858), .ZN(n4419) );
  INV_X1 U4340 ( .A(n4421), .ZN(n4420) );
  NAND2_X1 U4341 ( .A1(n4375), .A2(n4376), .ZN(n4421) );
  NOR2_X1 U4342 ( .A1(n4375), .A2(n4376), .ZN(n4418) );
  NOR2_X1 U4343 ( .A1(n4422), .A2(n4423), .ZN(n4376) );
  NOR3_X1 U4344 ( .A1(n2679), .A2(n4424), .A3(n2858), .ZN(n4423) );
  INV_X1 U4345 ( .A(n4425), .ZN(n4424) );
  NAND2_X1 U4346 ( .A1(n4292), .A2(n4294), .ZN(n4425) );
  NOR2_X1 U4347 ( .A1(n4292), .A2(n4294), .ZN(n4422) );
  NOR2_X1 U4348 ( .A1(n4426), .A2(n4427), .ZN(n4294) );
  NOR3_X1 U4349 ( .A1(n2854), .A2(n4428), .A3(n2858), .ZN(n4427) );
  INV_X1 U4350 ( .A(n4429), .ZN(n4428) );
  NAND2_X1 U4351 ( .A1(n4371), .A2(n4372), .ZN(n4429) );
  NOR2_X1 U4352 ( .A1(n4371), .A2(n4372), .ZN(n4426) );
  NOR2_X1 U4353 ( .A1(n4430), .A2(n4431), .ZN(n4372) );
  NOR3_X1 U4354 ( .A1(n2628), .A2(n4432), .A3(n2858), .ZN(n4431) );
  NOR2_X1 U4355 ( .A1(n4366), .A2(n4368), .ZN(n4432) );
  INV_X1 U4356 ( .A(n4433), .ZN(n4430) );
  NAND2_X1 U4357 ( .A1(n4366), .A2(n4368), .ZN(n4433) );
  NAND2_X1 U4358 ( .A1(n4434), .A2(n4435), .ZN(n4368) );
  NAND3_X1 U4359 ( .A1(a_8_), .A2(n4436), .A3(b_3_), .ZN(n4435) );
  INV_X1 U4360 ( .A(n4437), .ZN(n4436) );
  NOR2_X1 U4361 ( .A1(n4363), .A2(n4364), .ZN(n4437) );
  NAND2_X1 U4362 ( .A1(n4363), .A2(n4364), .ZN(n4434) );
  NAND2_X1 U4363 ( .A1(n4438), .A2(n4439), .ZN(n4364) );
  NAND3_X1 U4364 ( .A1(a_9_), .A2(n4440), .A3(b_3_), .ZN(n4439) );
  INV_X1 U4365 ( .A(n4441), .ZN(n4440) );
  NOR2_X1 U4366 ( .A1(n4359), .A2(n4360), .ZN(n4441) );
  NAND2_X1 U4367 ( .A1(n4359), .A2(n4360), .ZN(n4438) );
  NAND2_X1 U4368 ( .A1(n4356), .A2(n4442), .ZN(n4360) );
  NAND2_X1 U4369 ( .A1(n4355), .A2(n4357), .ZN(n4442) );
  NAND2_X1 U4370 ( .A1(n4443), .A2(n4444), .ZN(n4357) );
  NAND2_X1 U4371 ( .A1(b_3_), .A2(a_10_), .ZN(n4444) );
  INV_X1 U4372 ( .A(n4445), .ZN(n4443) );
  XNOR2_X1 U4373 ( .A(n4446), .B(n4447), .ZN(n4355) );
  XNOR2_X1 U4374 ( .A(n4448), .B(n4449), .ZN(n4447) );
  NAND2_X1 U4375 ( .A1(a_10_), .A2(n4445), .ZN(n4356) );
  NAND2_X1 U4376 ( .A1(n4352), .A2(n4450), .ZN(n4445) );
  NAND2_X1 U4377 ( .A1(n4351), .A2(n4353), .ZN(n4450) );
  NAND2_X1 U4378 ( .A1(n4451), .A2(n4452), .ZN(n4353) );
  NAND2_X1 U4379 ( .A1(b_3_), .A2(a_11_), .ZN(n4452) );
  XOR2_X1 U4380 ( .A(n4453), .B(n4454), .Z(n4351) );
  XOR2_X1 U4381 ( .A(n4455), .B(n4456), .Z(n4453) );
  INV_X1 U4382 ( .A(n4457), .ZN(n4352) );
  NOR2_X1 U4383 ( .A1(n2846), .A2(n4451), .ZN(n4457) );
  NOR2_X1 U4384 ( .A1(n4458), .A2(n4459), .ZN(n4451) );
  INV_X1 U4385 ( .A(n4460), .ZN(n4459) );
  NAND2_X1 U4386 ( .A1(n4348), .A2(n4461), .ZN(n4460) );
  NAND2_X1 U4387 ( .A1(n4349), .A2(n4347), .ZN(n4461) );
  NOR2_X1 U4388 ( .A1(n2858), .A2(n2844), .ZN(n4348) );
  NOR2_X1 U4389 ( .A1(n4347), .A2(n4349), .ZN(n4458) );
  NOR2_X1 U4390 ( .A1(n4462), .A2(n4463), .ZN(n4349) );
  INV_X1 U4391 ( .A(n4464), .ZN(n4463) );
  NAND2_X1 U4392 ( .A1(n4342), .A2(n4465), .ZN(n4464) );
  NAND2_X1 U4393 ( .A1(n4466), .A2(n4344), .ZN(n4465) );
  NOR2_X1 U4394 ( .A1(n2858), .A2(n2842), .ZN(n4342) );
  NOR2_X1 U4395 ( .A1(n4344), .A2(n4466), .ZN(n4462) );
  INV_X1 U4396 ( .A(n4345), .ZN(n4466) );
  NAND2_X1 U4397 ( .A1(n4467), .A2(n4468), .ZN(n4345) );
  NAND2_X1 U4398 ( .A1(b_1_), .A2(n4469), .ZN(n4468) );
  NAND2_X1 U4399 ( .A1(n2426), .A2(n4470), .ZN(n4469) );
  NAND2_X1 U4400 ( .A1(a_15_), .A2(n2859), .ZN(n4470) );
  NAND2_X1 U4401 ( .A1(b_2_), .A2(n4471), .ZN(n4467) );
  NAND2_X1 U4402 ( .A1(n3049), .A2(n4472), .ZN(n4471) );
  NAND2_X1 U4403 ( .A1(a_14_), .A2(n2861), .ZN(n4472) );
  NAND3_X1 U4404 ( .A1(b_2_), .A2(b_3_), .A3(n2840), .ZN(n4344) );
  XOR2_X1 U4405 ( .A(n4473), .B(n4474), .Z(n4347) );
  XNOR2_X1 U4406 ( .A(n4475), .B(n4476), .ZN(n4474) );
  XOR2_X1 U4407 ( .A(n4477), .B(n4478), .Z(n4359) );
  XOR2_X1 U4408 ( .A(n4479), .B(n4480), .Z(n4477) );
  XOR2_X1 U4409 ( .A(n4481), .B(n4482), .Z(n4363) );
  XOR2_X1 U4410 ( .A(n4483), .B(n4484), .Z(n4481) );
  XOR2_X1 U4411 ( .A(n4485), .B(n4486), .Z(n4366) );
  XOR2_X1 U4412 ( .A(n4487), .B(n4488), .Z(n4485) );
  XNOR2_X1 U4413 ( .A(n4489), .B(n4490), .ZN(n4371) );
  XOR2_X1 U4414 ( .A(n4491), .B(n4492), .Z(n4489) );
  XNOR2_X1 U4415 ( .A(n4493), .B(n4494), .ZN(n4292) );
  XOR2_X1 U4416 ( .A(n4495), .B(n4496), .Z(n4493) );
  XNOR2_X1 U4417 ( .A(n4497), .B(n4498), .ZN(n4375) );
  XOR2_X1 U4418 ( .A(n4499), .B(n4500), .Z(n4497) );
  XNOR2_X1 U4419 ( .A(n4501), .B(n4502), .ZN(n4385) );
  XNOR2_X1 U4420 ( .A(n2764), .B(n4503), .ZN(n4501) );
  XNOR2_X1 U4421 ( .A(n4504), .B(n4505), .ZN(n4390) );
  XOR2_X1 U4422 ( .A(n4506), .B(n4507), .Z(n4504) );
  NOR2_X1 U4423 ( .A1(n2790), .A2(n2859), .ZN(n4507) );
  XNOR2_X1 U4424 ( .A(n4269), .B(n4270), .ZN(n4393) );
  NAND2_X1 U4425 ( .A1(n4508), .A2(n4509), .ZN(n4269) );
  NAND2_X1 U4426 ( .A1(n4510), .A2(n4511), .ZN(n2710) );
  XOR2_X1 U4427 ( .A(n2714), .B(n2713), .Z(n4510) );
  INV_X1 U4428 ( .A(n2863), .ZN(n2714) );
  NAND2_X1 U4429 ( .A1(b_0_), .A2(a_0_), .ZN(n2863) );
  NAND2_X1 U4430 ( .A1(a_0_), .A2(n4512), .ZN(n2906) );
  NAND2_X1 U4431 ( .A1(n2713), .A2(n4513), .ZN(n4512) );
  NAND2_X1 U4432 ( .A1(n2712), .A2(b_0_), .ZN(n4513) );
  INV_X1 U4433 ( .A(n4511), .ZN(n2712) );
  NAND2_X1 U4434 ( .A1(n2909), .A2(n2908), .ZN(n4511) );
  NAND2_X1 U4435 ( .A1(n4508), .A2(n4514), .ZN(n2908) );
  NAND2_X1 U4436 ( .A1(n4270), .A2(n4509), .ZN(n4514) );
  NAND2_X1 U4437 ( .A1(n4515), .A2(n4516), .ZN(n4509) );
  NAND2_X1 U4438 ( .A1(b_2_), .A2(a_0_), .ZN(n4516) );
  XOR2_X1 U4439 ( .A(n4517), .B(n4518), .Z(n4270) );
  NOR2_X1 U4440 ( .A1(n2860), .A2(n2866), .ZN(n4518) );
  XOR2_X1 U4441 ( .A(n2816), .B(n4519), .Z(n4517) );
  INV_X1 U4442 ( .A(n4520), .ZN(n4508) );
  NOR2_X1 U4443 ( .A1(n2865), .A2(n4515), .ZN(n4520) );
  NOR2_X1 U4444 ( .A1(n4521), .A2(n4522), .ZN(n4515) );
  NOR3_X1 U4445 ( .A1(n2790), .A2(n4523), .A3(n2859), .ZN(n4522) );
  NOR2_X1 U4446 ( .A1(n4506), .A2(n4505), .ZN(n4523) );
  INV_X1 U4447 ( .A(n4524), .ZN(n4521) );
  NAND2_X1 U4448 ( .A1(n4505), .A2(n4506), .ZN(n4524) );
  NAND2_X1 U4449 ( .A1(n4525), .A2(n4526), .ZN(n4506) );
  INV_X1 U4450 ( .A(n4527), .ZN(n4526) );
  NOR2_X1 U4451 ( .A1(n2764), .A2(n4528), .ZN(n4527) );
  NOR2_X1 U4452 ( .A1(n4503), .A2(n4502), .ZN(n4528) );
  NAND2_X1 U4453 ( .A1(b_2_), .A2(a_2_), .ZN(n2764) );
  NAND2_X1 U4454 ( .A1(n4502), .A2(n4503), .ZN(n4525) );
  NAND2_X1 U4455 ( .A1(n4529), .A2(n4530), .ZN(n4503) );
  NAND2_X1 U4456 ( .A1(n4409), .A2(n4531), .ZN(n4530) );
  INV_X1 U4457 ( .A(n4532), .ZN(n4531) );
  NOR2_X1 U4458 ( .A1(n4408), .A2(n4407), .ZN(n4532) );
  NOR2_X1 U4459 ( .A1(n2859), .A2(n2739), .ZN(n4409) );
  NAND2_X1 U4460 ( .A1(n4407), .A2(n4408), .ZN(n4529) );
  NAND2_X1 U4461 ( .A1(n4533), .A2(n4534), .ZN(n4408) );
  NAND2_X1 U4462 ( .A1(n4416), .A2(n4535), .ZN(n4534) );
  INV_X1 U4463 ( .A(n4536), .ZN(n4535) );
  NOR2_X1 U4464 ( .A1(n4417), .A2(n4415), .ZN(n4536) );
  NOR2_X1 U4465 ( .A1(n2859), .A2(n2857), .ZN(n4416) );
  NAND2_X1 U4466 ( .A1(n4415), .A2(n4417), .ZN(n4533) );
  NAND2_X1 U4467 ( .A1(n4537), .A2(n4538), .ZN(n4417) );
  NAND2_X1 U4468 ( .A1(n4500), .A2(n4539), .ZN(n4538) );
  INV_X1 U4469 ( .A(n4540), .ZN(n4539) );
  NOR2_X1 U4470 ( .A1(n4499), .A2(n4498), .ZN(n4540) );
  NOR2_X1 U4471 ( .A1(n2859), .A2(n2679), .ZN(n4500) );
  NAND2_X1 U4472 ( .A1(n4498), .A2(n4499), .ZN(n4537) );
  NAND2_X1 U4473 ( .A1(n4541), .A2(n4542), .ZN(n4499) );
  NAND2_X1 U4474 ( .A1(n4495), .A2(n4543), .ZN(n4542) );
  INV_X1 U4475 ( .A(n4544), .ZN(n4543) );
  NOR2_X1 U4476 ( .A1(n4496), .A2(n4494), .ZN(n4544) );
  NOR2_X1 U4477 ( .A1(n2859), .A2(n2854), .ZN(n4495) );
  NAND2_X1 U4478 ( .A1(n4494), .A2(n4496), .ZN(n4541) );
  NAND2_X1 U4479 ( .A1(n4545), .A2(n4546), .ZN(n4496) );
  NAND2_X1 U4480 ( .A1(n4492), .A2(n4547), .ZN(n4546) );
  INV_X1 U4481 ( .A(n4548), .ZN(n4547) );
  NOR2_X1 U4482 ( .A1(n4491), .A2(n4490), .ZN(n4548) );
  NOR2_X1 U4483 ( .A1(n2859), .A2(n2628), .ZN(n4492) );
  NAND2_X1 U4484 ( .A1(n4490), .A2(n4491), .ZN(n4545) );
  NAND2_X1 U4485 ( .A1(n4549), .A2(n4550), .ZN(n4491) );
  NAND2_X1 U4486 ( .A1(n4487), .A2(n4551), .ZN(n4550) );
  INV_X1 U4487 ( .A(n4552), .ZN(n4551) );
  NOR2_X1 U4488 ( .A1(n4488), .A2(n4486), .ZN(n4552) );
  NOR2_X1 U4489 ( .A1(n2859), .A2(n2851), .ZN(n4487) );
  NAND2_X1 U4490 ( .A1(n4486), .A2(n4488), .ZN(n4549) );
  NAND2_X1 U4491 ( .A1(n4553), .A2(n4554), .ZN(n4488) );
  NAND2_X1 U4492 ( .A1(n4484), .A2(n4555), .ZN(n4554) );
  INV_X1 U4493 ( .A(n4556), .ZN(n4555) );
  NOR2_X1 U4494 ( .A1(n4483), .A2(n4482), .ZN(n4556) );
  NOR2_X1 U4495 ( .A1(n2859), .A2(n2577), .ZN(n4484) );
  NAND2_X1 U4496 ( .A1(n4482), .A2(n4483), .ZN(n4553) );
  NAND2_X1 U4497 ( .A1(n4557), .A2(n4558), .ZN(n4483) );
  NAND2_X1 U4498 ( .A1(n4479), .A2(n4559), .ZN(n4558) );
  INV_X1 U4499 ( .A(n4560), .ZN(n4559) );
  NOR2_X1 U4500 ( .A1(n4480), .A2(n4478), .ZN(n4560) );
  NOR2_X1 U4501 ( .A1(n2859), .A2(n2849), .ZN(n4479) );
  NAND2_X1 U4502 ( .A1(n4478), .A2(n4480), .ZN(n4557) );
  NAND2_X1 U4503 ( .A1(n4561), .A2(n4562), .ZN(n4480) );
  NAND2_X1 U4504 ( .A1(n4449), .A2(n4563), .ZN(n4562) );
  INV_X1 U4505 ( .A(n4564), .ZN(n4563) );
  NOR2_X1 U4506 ( .A1(n4448), .A2(n4446), .ZN(n4564) );
  NOR2_X1 U4507 ( .A1(n2859), .A2(n2846), .ZN(n4449) );
  NAND2_X1 U4508 ( .A1(n4446), .A2(n4448), .ZN(n4561) );
  NAND2_X1 U4509 ( .A1(n4565), .A2(n4566), .ZN(n4448) );
  NAND2_X1 U4510 ( .A1(n4455), .A2(n4567), .ZN(n4566) );
  INV_X1 U4511 ( .A(n4568), .ZN(n4567) );
  NOR2_X1 U4512 ( .A1(n4454), .A2(n4456), .ZN(n4568) );
  NOR2_X1 U4513 ( .A1(n2859), .A2(n2844), .ZN(n4455) );
  NAND2_X1 U4514 ( .A1(n4454), .A2(n4456), .ZN(n4565) );
  NAND2_X1 U4515 ( .A1(n4569), .A2(n4570), .ZN(n4456) );
  NAND2_X1 U4516 ( .A1(n4473), .A2(n4571), .ZN(n4570) );
  INV_X1 U4517 ( .A(n4572), .ZN(n4571) );
  NOR2_X1 U4518 ( .A1(n4476), .A2(n4475), .ZN(n4572) );
  NOR2_X1 U4519 ( .A1(n2859), .A2(n2842), .ZN(n4473) );
  NAND2_X1 U4520 ( .A1(n4475), .A2(n4476), .ZN(n4569) );
  NAND2_X1 U4521 ( .A1(n4573), .A2(n4574), .ZN(n4476) );
  NAND2_X1 U4522 ( .A1(b_0_), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U4523 ( .A1(n2426), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U4524 ( .A1(a_15_), .A2(n2861), .ZN(n4576) );
  NAND2_X1 U4525 ( .A1(a_15_), .A2(n2428), .ZN(n2426) );
  NAND2_X1 U4526 ( .A1(b_1_), .A2(n4577), .ZN(n4573) );
  NAND2_X1 U4527 ( .A1(n3049), .A2(n4578), .ZN(n4577) );
  NAND2_X1 U4528 ( .A1(a_14_), .A2(n2866), .ZN(n4578) );
  NAND2_X1 U4529 ( .A1(a_14_), .A2(n4579), .ZN(n3049) );
  NOR3_X1 U4530 ( .A1(n2861), .A2(n2859), .A3(n3043), .ZN(n4475) );
  INV_X1 U4531 ( .A(n2840), .ZN(n3043) );
  XNOR2_X1 U4532 ( .A(n4580), .B(n4581), .ZN(n4454) );
  XNOR2_X1 U4533 ( .A(n4582), .B(n4583), .ZN(n4581) );
  NAND2_X1 U4534 ( .A1(b_0_), .A2(a_14_), .ZN(n4580) );
  XNOR2_X1 U4535 ( .A(n4584), .B(n4585), .ZN(n4446) );
  NAND2_X1 U4536 ( .A1(n4586), .A2(n4587), .ZN(n4584) );
  NAND2_X1 U4537 ( .A1(n4588), .A2(n4589), .ZN(n4587) );
  NAND2_X1 U4538 ( .A1(b_1_), .A2(a_12_), .ZN(n4588) );
  XOR2_X1 U4539 ( .A(n4590), .B(n4591), .Z(n4478) );
  XOR2_X1 U4540 ( .A(n4592), .B(n4593), .Z(n4591) );
  NAND2_X1 U4541 ( .A1(b_1_), .A2(a_11_), .ZN(n4590) );
  XOR2_X1 U4542 ( .A(n4594), .B(n4595), .Z(n4482) );
  XNOR2_X1 U4543 ( .A(n4596), .B(n4597), .ZN(n4595) );
  NAND2_X1 U4544 ( .A1(b_1_), .A2(a_10_), .ZN(n4594) );
  XOR2_X1 U4545 ( .A(n4598), .B(n4599), .Z(n4486) );
  NOR2_X1 U4546 ( .A1(n2577), .A2(n2861), .ZN(n4599) );
  XOR2_X1 U4547 ( .A(n4600), .B(n4601), .Z(n4598) );
  XOR2_X1 U4548 ( .A(n4602), .B(n4603), .Z(n4490) );
  XNOR2_X1 U4549 ( .A(n4604), .B(n4605), .ZN(n4603) );
  NAND2_X1 U4550 ( .A1(b_1_), .A2(a_8_), .ZN(n4602) );
  XOR2_X1 U4551 ( .A(n4606), .B(n4607), .Z(n4494) );
  NOR2_X1 U4552 ( .A1(n2628), .A2(n2861), .ZN(n4607) );
  XOR2_X1 U4553 ( .A(n4608), .B(n4609), .Z(n4606) );
  XOR2_X1 U4554 ( .A(n4610), .B(n4611), .Z(n4498) );
  XNOR2_X1 U4555 ( .A(n4612), .B(n4613), .ZN(n4611) );
  NAND2_X1 U4556 ( .A1(b_1_), .A2(a_6_), .ZN(n4610) );
  XOR2_X1 U4557 ( .A(n4614), .B(n4615), .Z(n4415) );
  NOR2_X1 U4558 ( .A1(n2679), .A2(n2861), .ZN(n4615) );
  XOR2_X1 U4559 ( .A(n4616), .B(n4617), .Z(n4614) );
  XOR2_X1 U4560 ( .A(n4618), .B(n4619), .Z(n4407) );
  XNOR2_X1 U4561 ( .A(n4620), .B(n4621), .ZN(n4619) );
  NAND2_X1 U4562 ( .A1(b_1_), .A2(a_4_), .ZN(n4618) );
  XOR2_X1 U4563 ( .A(n4622), .B(n4623), .Z(n4502) );
  NOR2_X1 U4564 ( .A1(n2739), .A2(n2861), .ZN(n4623) );
  XOR2_X1 U4565 ( .A(n4624), .B(n4625), .Z(n4622) );
  XOR2_X1 U4566 ( .A(n4626), .B(n4627), .Z(n4505) );
  XNOR2_X1 U4567 ( .A(n4628), .B(n4629), .ZN(n4627) );
  NAND2_X1 U4568 ( .A1(b_1_), .A2(a_2_), .ZN(n4626) );
  XOR2_X1 U4569 ( .A(n4630), .B(n4631), .Z(n2909) );
  XNOR2_X1 U4570 ( .A(n4632), .B(n4633), .ZN(n4631) );
  NAND2_X1 U4571 ( .A1(b_0_), .A2(a_1_), .ZN(n4630) );
  NOR2_X1 U4572 ( .A1(n4634), .A2(n4635), .ZN(n2713) );
  INV_X1 U4573 ( .A(n4636), .ZN(n4635) );
  NAND3_X1 U4574 ( .A1(a_1_), .A2(n4637), .A3(b_0_), .ZN(n4636) );
  NAND2_X1 U4575 ( .A1(n4633), .A2(n4632), .ZN(n4637) );
  NOR2_X1 U4576 ( .A1(n4632), .A2(n4633), .ZN(n4634) );
  NOR2_X1 U4577 ( .A1(n4638), .A2(n4639), .ZN(n4633) );
  NOR3_X1 U4578 ( .A1(n2860), .A2(n4640), .A3(n2866), .ZN(n4639) );
  INV_X1 U4579 ( .A(n4641), .ZN(n4640) );
  NAND2_X1 U4580 ( .A1(n4519), .A2(n2816), .ZN(n4641) );
  NOR2_X1 U4581 ( .A1(n2816), .A2(n4519), .ZN(n4638) );
  NOR2_X1 U4582 ( .A1(n4642), .A2(n4643), .ZN(n4519) );
  INV_X1 U4583 ( .A(n4644), .ZN(n4643) );
  NAND3_X1 U4584 ( .A1(a_2_), .A2(n4645), .A3(b_1_), .ZN(n4644) );
  NAND2_X1 U4585 ( .A1(n4629), .A2(n4628), .ZN(n4645) );
  NOR2_X1 U4586 ( .A1(n4628), .A2(n4629), .ZN(n4642) );
  NOR2_X1 U4587 ( .A1(n4646), .A2(n4647), .ZN(n4629) );
  NOR3_X1 U4588 ( .A1(n2739), .A2(n4648), .A3(n2861), .ZN(n4647) );
  INV_X1 U4589 ( .A(n4649), .ZN(n4648) );
  NAND2_X1 U4590 ( .A1(n4625), .A2(n4624), .ZN(n4649) );
  NOR2_X1 U4591 ( .A1(n4624), .A2(n4625), .ZN(n4646) );
  NOR2_X1 U4592 ( .A1(n4650), .A2(n4651), .ZN(n4625) );
  INV_X1 U4593 ( .A(n4652), .ZN(n4651) );
  NAND3_X1 U4594 ( .A1(a_4_), .A2(n4653), .A3(b_1_), .ZN(n4652) );
  NAND2_X1 U4595 ( .A1(n4621), .A2(n4620), .ZN(n4653) );
  NOR2_X1 U4596 ( .A1(n4620), .A2(n4621), .ZN(n4650) );
  NOR2_X1 U4597 ( .A1(n4654), .A2(n4655), .ZN(n4621) );
  NOR3_X1 U4598 ( .A1(n2679), .A2(n4656), .A3(n2861), .ZN(n4655) );
  INV_X1 U4599 ( .A(n4657), .ZN(n4656) );
  NAND2_X1 U4600 ( .A1(n4617), .A2(n4616), .ZN(n4657) );
  NOR2_X1 U4601 ( .A1(n4616), .A2(n4617), .ZN(n4654) );
  NOR2_X1 U4602 ( .A1(n4658), .A2(n4659), .ZN(n4617) );
  INV_X1 U4603 ( .A(n4660), .ZN(n4659) );
  NAND3_X1 U4604 ( .A1(a_6_), .A2(n4661), .A3(b_1_), .ZN(n4660) );
  NAND2_X1 U4605 ( .A1(n4613), .A2(n4612), .ZN(n4661) );
  NOR2_X1 U4606 ( .A1(n4612), .A2(n4613), .ZN(n4658) );
  NOR2_X1 U4607 ( .A1(n4662), .A2(n4663), .ZN(n4613) );
  NOR3_X1 U4608 ( .A1(n2628), .A2(n4664), .A3(n2861), .ZN(n4663) );
  INV_X1 U4609 ( .A(n4665), .ZN(n4664) );
  NAND2_X1 U4610 ( .A1(n4609), .A2(n4608), .ZN(n4665) );
  NOR2_X1 U4611 ( .A1(n4608), .A2(n4609), .ZN(n4662) );
  NOR2_X1 U4612 ( .A1(n4666), .A2(n4667), .ZN(n4609) );
  INV_X1 U4613 ( .A(n4668), .ZN(n4667) );
  NAND3_X1 U4614 ( .A1(a_8_), .A2(n4669), .A3(b_1_), .ZN(n4668) );
  NAND2_X1 U4615 ( .A1(n4605), .A2(n4604), .ZN(n4669) );
  NOR2_X1 U4616 ( .A1(n4604), .A2(n4605), .ZN(n4666) );
  NOR2_X1 U4617 ( .A1(n4670), .A2(n4671), .ZN(n4605) );
  NOR3_X1 U4618 ( .A1(n2577), .A2(n4672), .A3(n2861), .ZN(n4671) );
  INV_X1 U4619 ( .A(n4673), .ZN(n4672) );
  NAND2_X1 U4620 ( .A1(n4601), .A2(n4600), .ZN(n4673) );
  NOR2_X1 U4621 ( .A1(n4600), .A2(n4601), .ZN(n4670) );
  NOR2_X1 U4622 ( .A1(n4674), .A2(n4675), .ZN(n4601) );
  NOR3_X1 U4623 ( .A1(n2849), .A2(n4676), .A3(n2861), .ZN(n4675) );
  NOR2_X1 U4624 ( .A1(n4597), .A2(n4596), .ZN(n4676) );
  INV_X1 U4625 ( .A(n4677), .ZN(n4674) );
  NAND2_X1 U4626 ( .A1(n4596), .A2(n4597), .ZN(n4677) );
  NAND2_X1 U4627 ( .A1(n4678), .A2(n4679), .ZN(n4597) );
  NAND3_X1 U4628 ( .A1(a_11_), .A2(n4680), .A3(b_1_), .ZN(n4679) );
  NAND2_X1 U4629 ( .A1(n4593), .A2(n4681), .ZN(n4680) );
  INV_X1 U4630 ( .A(n4682), .ZN(n4593) );
  NAND2_X1 U4631 ( .A1(n4592), .A2(n4682), .ZN(n4678) );
  NAND2_X1 U4632 ( .A1(n4586), .A2(n4683), .ZN(n4682) );
  NAND2_X1 U4633 ( .A1(n4684), .A2(n4585), .ZN(n4683) );
  NAND2_X1 U4634 ( .A1(n4583), .A2(n4685), .ZN(n4585) );
  NAND3_X1 U4635 ( .A1(b_0_), .A2(a_14_), .A3(n4582), .ZN(n4685) );
  NOR2_X1 U4636 ( .A1(n2861), .A2(n2842), .ZN(n4582) );
  NAND3_X1 U4637 ( .A1(b_1_), .A2(b_0_), .A3(n2840), .ZN(n4583) );
  INV_X1 U4638 ( .A(a_15_), .ZN(n4579) );
  NAND2_X1 U4639 ( .A1(n4589), .A2(n2844), .ZN(n4684) );
  INV_X1 U4640 ( .A(n4686), .ZN(n4589) );
  NAND3_X1 U4641 ( .A1(b_1_), .A2(a_12_), .A3(n4686), .ZN(n4586) );
  NOR2_X1 U4642 ( .A1(n2866), .A2(n2842), .ZN(n4686) );
  INV_X1 U4643 ( .A(n4681), .ZN(n4592) );
  NAND2_X1 U4644 ( .A1(b_0_), .A2(a_12_), .ZN(n4681) );
  NOR2_X1 U4645 ( .A1(n2866), .A2(n2846), .ZN(n4596) );
  NAND2_X1 U4646 ( .A1(b_0_), .A2(a_10_), .ZN(n4600) );
  NAND2_X1 U4647 ( .A1(b_0_), .A2(a_9_), .ZN(n4604) );
  NAND2_X1 U4648 ( .A1(b_0_), .A2(a_8_), .ZN(n4608) );
  NAND2_X1 U4649 ( .A1(b_0_), .A2(a_7_), .ZN(n4612) );
  NAND2_X1 U4650 ( .A1(b_0_), .A2(a_6_), .ZN(n4616) );
  NAND2_X1 U4651 ( .A1(b_0_), .A2(a_5_), .ZN(n4620) );
  NAND2_X1 U4652 ( .A1(b_0_), .A2(a_4_), .ZN(n4624) );
  NAND2_X1 U4653 ( .A1(b_0_), .A2(a_3_), .ZN(n4628) );
  NAND2_X1 U4654 ( .A1(b_1_), .A2(a_1_), .ZN(n2816) );
  NAND2_X1 U4655 ( .A1(b_1_), .A2(a_0_), .ZN(n4632) );
  NOR2_X1 U4656 ( .A1(n4687), .A2(n4688), .ZN(n2352) );
  INV_X1 U4657 ( .A(n4689), .ZN(n2350) );
  NAND2_X1 U4658 ( .A1(n4690), .A2(n4691), .ZN(n4689) );
  NAND2_X1 U4659 ( .A1(n2347), .A2(n4692), .ZN(n4691) );
  NAND2_X1 U4660 ( .A1(n4693), .A2(n4694), .ZN(n4692) );
  NAND2_X1 U4661 ( .A1(b_0_), .A2(n4695), .ZN(n4694) );
  NAND2_X1 U4662 ( .A1(a_0_), .A2(n2862), .ZN(n4695) );
  NAND2_X1 U4663 ( .A1(n2807), .A2(n2865), .ZN(n4693) );
  INV_X1 U4664 ( .A(n2862), .ZN(n2807) );
  NAND2_X1 U4665 ( .A1(n4696), .A2(n4697), .ZN(n2862) );
  NAND2_X1 U4666 ( .A1(n4698), .A2(n2861), .ZN(n4697) );
  INV_X1 U4667 ( .A(b_1_), .ZN(n2861) );
  NAND2_X1 U4668 ( .A1(n2789), .A2(n2790), .ZN(n4698) );
  INV_X1 U4669 ( .A(n2781), .ZN(n2789) );
  NAND2_X1 U4670 ( .A1(a_1_), .A2(n2781), .ZN(n4696) );
  NAND2_X1 U4671 ( .A1(n4699), .A2(n4700), .ZN(n2781) );
  NAND2_X1 U4672 ( .A1(n4701), .A2(n2859), .ZN(n4700) );
  INV_X1 U4673 ( .A(b_2_), .ZN(n2859) );
  NAND2_X1 U4674 ( .A1(n2755), .A2(n2860), .ZN(n4701) );
  INV_X1 U4675 ( .A(n2763), .ZN(n2755) );
  NAND2_X1 U4676 ( .A1(a_2_), .A2(n2763), .ZN(n4699) );
  NAND2_X1 U4677 ( .A1(n4702), .A2(n4703), .ZN(n2763) );
  NAND2_X1 U4678 ( .A1(n4704), .A2(n2858), .ZN(n4703) );
  INV_X1 U4679 ( .A(b_3_), .ZN(n2858) );
  NAND2_X1 U4680 ( .A1(n2738), .A2(n2739), .ZN(n4704) );
  INV_X1 U4681 ( .A(n2731), .ZN(n2738) );
  NAND2_X1 U4682 ( .A1(a_3_), .A2(n2731), .ZN(n4702) );
  NAND2_X1 U4683 ( .A1(n4705), .A2(n4706), .ZN(n2731) );
  NAND2_X1 U4684 ( .A1(n4707), .A2(n2856), .ZN(n4706) );
  INV_X1 U4685 ( .A(b_4_), .ZN(n2856) );
  NAND2_X1 U4686 ( .A1(n2695), .A2(n2857), .ZN(n4707) );
  INV_X1 U4687 ( .A(n2703), .ZN(n2695) );
  NAND2_X1 U4688 ( .A1(a_4_), .A2(n2703), .ZN(n4705) );
  NAND2_X1 U4689 ( .A1(n4708), .A2(n4709), .ZN(n2703) );
  NAND2_X1 U4690 ( .A1(n4710), .A2(n2855), .ZN(n4709) );
  INV_X1 U4691 ( .A(b_5_), .ZN(n2855) );
  NAND2_X1 U4692 ( .A1(n2678), .A2(n2679), .ZN(n4710) );
  INV_X1 U4693 ( .A(n2671), .ZN(n2678) );
  NAND2_X1 U4694 ( .A1(a_5_), .A2(n2671), .ZN(n4708) );
  NAND2_X1 U4695 ( .A1(n4711), .A2(n4712), .ZN(n2671) );
  NAND2_X1 U4696 ( .A1(n4713), .A2(n2853), .ZN(n4712) );
  INV_X1 U4697 ( .A(b_6_), .ZN(n2853) );
  NAND2_X1 U4698 ( .A1(n2644), .A2(n2854), .ZN(n4713) );
  INV_X1 U4699 ( .A(n2652), .ZN(n2644) );
  NAND2_X1 U4700 ( .A1(a_6_), .A2(n2652), .ZN(n4711) );
  NAND2_X1 U4701 ( .A1(n4714), .A2(n4715), .ZN(n2652) );
  NAND2_X1 U4702 ( .A1(n4716), .A2(n2852), .ZN(n4715) );
  INV_X1 U4703 ( .A(b_7_), .ZN(n2852) );
  NAND2_X1 U4704 ( .A1(n2627), .A2(n2628), .ZN(n4716) );
  INV_X1 U4705 ( .A(n2620), .ZN(n2627) );
  NAND2_X1 U4706 ( .A1(a_7_), .A2(n2620), .ZN(n4714) );
  NAND2_X1 U4707 ( .A1(n4717), .A2(n4718), .ZN(n2620) );
  NAND2_X1 U4708 ( .A1(n4719), .A2(n2850), .ZN(n4718) );
  INV_X1 U4709 ( .A(b_8_), .ZN(n2850) );
  NAND2_X1 U4710 ( .A1(n2593), .A2(n2851), .ZN(n4719) );
  INV_X1 U4711 ( .A(n2601), .ZN(n2593) );
  NAND2_X1 U4712 ( .A1(a_8_), .A2(n2601), .ZN(n4717) );
  NAND2_X1 U4713 ( .A1(n4720), .A2(n4721), .ZN(n2601) );
  NAND2_X1 U4714 ( .A1(n4722), .A2(n3495), .ZN(n4721) );
  INV_X1 U4715 ( .A(b_9_), .ZN(n3495) );
  NAND2_X1 U4716 ( .A1(n2576), .A2(n2577), .ZN(n4722) );
  INV_X1 U4717 ( .A(n2568), .ZN(n2576) );
  NAND2_X1 U4718 ( .A1(a_9_), .A2(n2568), .ZN(n4720) );
  NAND2_X1 U4719 ( .A1(n4723), .A2(n4724), .ZN(n2568) );
  NAND2_X1 U4720 ( .A1(n4725), .A2(n2848), .ZN(n4724) );
  INV_X1 U4721 ( .A(b_10_), .ZN(n2848) );
  NAND2_X1 U4722 ( .A1(n2542), .A2(n2849), .ZN(n4725) );
  INV_X1 U4723 ( .A(n2550), .ZN(n2542) );
  NAND2_X1 U4724 ( .A1(a_10_), .A2(n2550), .ZN(n4723) );
  NAND2_X1 U4725 ( .A1(n4726), .A2(n4727), .ZN(n2550) );
  NAND2_X1 U4726 ( .A1(n4728), .A2(n2845), .ZN(n4727) );
  INV_X1 U4727 ( .A(b_11_), .ZN(n2845) );
  NAND2_X1 U4728 ( .A1(n2516), .A2(n2846), .ZN(n4728) );
  INV_X1 U4729 ( .A(n2524), .ZN(n2516) );
  NAND2_X1 U4730 ( .A1(a_11_), .A2(n2524), .ZN(n4726) );
  NAND2_X1 U4731 ( .A1(n4729), .A2(n4730), .ZN(n2524) );
  NAND2_X1 U4732 ( .A1(n4731), .A2(n2843), .ZN(n4730) );
  INV_X1 U4733 ( .A(b_12_), .ZN(n2843) );
  NAND2_X1 U4734 ( .A1(n2490), .A2(n2844), .ZN(n4731) );
  INV_X1 U4735 ( .A(n2498), .ZN(n2490) );
  NAND2_X1 U4736 ( .A1(a_12_), .A2(n2498), .ZN(n4729) );
  NAND2_X1 U4737 ( .A1(n4732), .A2(n4733), .ZN(n2498) );
  NAND2_X1 U4738 ( .A1(n4734), .A2(n2841), .ZN(n4733) );
  INV_X1 U4739 ( .A(b_13_), .ZN(n2841) );
  NAND2_X1 U4740 ( .A1(n2464), .A2(n2842), .ZN(n4734) );
  INV_X1 U4741 ( .A(n2472), .ZN(n2464) );
  NAND2_X1 U4742 ( .A1(a_13_), .A2(n2472), .ZN(n4732) );
  NAND2_X1 U4743 ( .A1(n4735), .A2(n4736), .ZN(n2472) );
  NAND2_X1 U4744 ( .A1(n4737), .A2(n2431), .ZN(n4736) );
  INV_X1 U4745 ( .A(b_14_), .ZN(n2431) );
  NAND2_X1 U4746 ( .A1(n2420), .A2(n2428), .ZN(n4737) );
  NAND2_X1 U4747 ( .A1(a_14_), .A2(n2415), .ZN(n4735) );
  INV_X1 U4748 ( .A(n2420), .ZN(n2415) );
  NOR2_X1 U4749 ( .A1(n2951), .A2(a_15_), .ZN(n2420) );
  NOR2_X1 U4750 ( .A1(n4688), .A2(operation_0_), .ZN(n2412) );
  INV_X1 U4751 ( .A(operation_1_), .ZN(n4688) );
  NAND2_X1 U4752 ( .A1(n2345), .A2(n4738), .ZN(n4690) );
  NAND2_X1 U4753 ( .A1(n4739), .A2(n4740), .ZN(n4738) );
  NAND2_X1 U4754 ( .A1(n4741), .A2(n2866), .ZN(n4740) );
  INV_X1 U4755 ( .A(b_0_), .ZN(n2866) );
  NAND2_X1 U4756 ( .A1(n2865), .A2(n2813), .ZN(n4741) );
  INV_X1 U4757 ( .A(a_0_), .ZN(n2865) );
  NAND2_X1 U4758 ( .A1(n2804), .A2(a_0_), .ZN(n4739) );
  INV_X1 U4759 ( .A(n2813), .ZN(n2804) );
  NAND2_X1 U4760 ( .A1(n4742), .A2(n4743), .ZN(n2813) );
  NAND2_X1 U4761 ( .A1(b_1_), .A2(n4744), .ZN(n4743) );
  NAND2_X1 U4762 ( .A1(n2787), .A2(a_1_), .ZN(n4744) );
  INV_X1 U4763 ( .A(n2779), .ZN(n2787) );
  NAND2_X1 U4764 ( .A1(n2779), .A2(n2790), .ZN(n4742) );
  INV_X1 U4765 ( .A(a_1_), .ZN(n2790) );
  NAND2_X1 U4766 ( .A1(n4745), .A2(n4746), .ZN(n2779) );
  NAND2_X1 U4767 ( .A1(b_2_), .A2(n4747), .ZN(n4746) );
  NAND2_X1 U4768 ( .A1(n2753), .A2(a_2_), .ZN(n4747) );
  INV_X1 U4769 ( .A(n2761), .ZN(n2753) );
  NAND2_X1 U4770 ( .A1(n2761), .A2(n2860), .ZN(n4745) );
  INV_X1 U4771 ( .A(a_2_), .ZN(n2860) );
  NAND2_X1 U4772 ( .A1(n4748), .A2(n4749), .ZN(n2761) );
  NAND2_X1 U4773 ( .A1(b_3_), .A2(n4750), .ZN(n4749) );
  NAND2_X1 U4774 ( .A1(n2737), .A2(a_3_), .ZN(n4750) );
  INV_X1 U4775 ( .A(n2728), .ZN(n2737) );
  NAND2_X1 U4776 ( .A1(n2728), .A2(n2739), .ZN(n4748) );
  INV_X1 U4777 ( .A(a_3_), .ZN(n2739) );
  NAND2_X1 U4778 ( .A1(n4751), .A2(n4752), .ZN(n2728) );
  NAND2_X1 U4779 ( .A1(b_4_), .A2(n4753), .ZN(n4752) );
  NAND2_X1 U4780 ( .A1(n2693), .A2(a_4_), .ZN(n4753) );
  INV_X1 U4781 ( .A(n2701), .ZN(n2693) );
  NAND2_X1 U4782 ( .A1(n2701), .A2(n2857), .ZN(n4751) );
  INV_X1 U4783 ( .A(a_4_), .ZN(n2857) );
  NAND2_X1 U4784 ( .A1(n4754), .A2(n4755), .ZN(n2701) );
  NAND2_X1 U4785 ( .A1(b_5_), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U4786 ( .A1(n2677), .A2(a_5_), .ZN(n4756) );
  INV_X1 U4787 ( .A(n2668), .ZN(n2677) );
  NAND2_X1 U4788 ( .A1(n2668), .A2(n2679), .ZN(n4754) );
  INV_X1 U4789 ( .A(a_5_), .ZN(n2679) );
  NAND2_X1 U4790 ( .A1(n4757), .A2(n4758), .ZN(n2668) );
  NAND2_X1 U4791 ( .A1(b_6_), .A2(n4759), .ZN(n4758) );
  NAND2_X1 U4792 ( .A1(n2642), .A2(a_6_), .ZN(n4759) );
  INV_X1 U4793 ( .A(n2650), .ZN(n2642) );
  NAND2_X1 U4794 ( .A1(n2650), .A2(n2854), .ZN(n4757) );
  INV_X1 U4795 ( .A(a_6_), .ZN(n2854) );
  NAND2_X1 U4796 ( .A1(n4760), .A2(n4761), .ZN(n2650) );
  NAND2_X1 U4797 ( .A1(b_7_), .A2(n4762), .ZN(n4761) );
  NAND2_X1 U4798 ( .A1(n2626), .A2(a_7_), .ZN(n4762) );
  INV_X1 U4799 ( .A(n2617), .ZN(n2626) );
  NAND2_X1 U4800 ( .A1(n2617), .A2(n2628), .ZN(n4760) );
  INV_X1 U4801 ( .A(a_7_), .ZN(n2628) );
  NAND2_X1 U4802 ( .A1(n4763), .A2(n4764), .ZN(n2617) );
  NAND2_X1 U4803 ( .A1(b_8_), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U4804 ( .A1(n2591), .A2(a_8_), .ZN(n4765) );
  INV_X1 U4805 ( .A(n2599), .ZN(n2591) );
  NAND2_X1 U4806 ( .A1(n2599), .A2(n2851), .ZN(n4763) );
  INV_X1 U4807 ( .A(a_8_), .ZN(n2851) );
  NAND2_X1 U4808 ( .A1(n4766), .A2(n4767), .ZN(n2599) );
  NAND2_X1 U4809 ( .A1(b_9_), .A2(n4768), .ZN(n4767) );
  NAND2_X1 U4810 ( .A1(n2574), .A2(a_9_), .ZN(n4768) );
  INV_X1 U4811 ( .A(n2566), .ZN(n2574) );
  NAND2_X1 U4812 ( .A1(n2566), .A2(n2577), .ZN(n4766) );
  INV_X1 U4813 ( .A(a_9_), .ZN(n2577) );
  NAND2_X1 U4814 ( .A1(n4769), .A2(n4770), .ZN(n2566) );
  NAND2_X1 U4815 ( .A1(b_10_), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U4816 ( .A1(n2540), .A2(a_10_), .ZN(n4771) );
  INV_X1 U4817 ( .A(n2548), .ZN(n2540) );
  NAND2_X1 U4818 ( .A1(n2548), .A2(n2849), .ZN(n4769) );
  INV_X1 U4819 ( .A(a_10_), .ZN(n2849) );
  NAND2_X1 U4820 ( .A1(n4772), .A2(n4773), .ZN(n2548) );
  NAND2_X1 U4821 ( .A1(b_11_), .A2(n4774), .ZN(n4773) );
  NAND2_X1 U4822 ( .A1(n2514), .A2(a_11_), .ZN(n4774) );
  INV_X1 U4823 ( .A(n2522), .ZN(n2514) );
  NAND2_X1 U4824 ( .A1(n2522), .A2(n2846), .ZN(n4772) );
  INV_X1 U4825 ( .A(a_11_), .ZN(n2846) );
  NAND2_X1 U4826 ( .A1(n4775), .A2(n4776), .ZN(n2522) );
  NAND2_X1 U4827 ( .A1(b_12_), .A2(n4777), .ZN(n4776) );
  NAND2_X1 U4828 ( .A1(n2488), .A2(a_12_), .ZN(n4777) );
  INV_X1 U4829 ( .A(n2496), .ZN(n2488) );
  NAND2_X1 U4830 ( .A1(n2496), .A2(n2844), .ZN(n4775) );
  INV_X1 U4831 ( .A(a_12_), .ZN(n2844) );
  NAND2_X1 U4832 ( .A1(n4778), .A2(n4779), .ZN(n2496) );
  NAND2_X1 U4833 ( .A1(b_13_), .A2(n4780), .ZN(n4779) );
  NAND2_X1 U4834 ( .A1(n2462), .A2(a_13_), .ZN(n4780) );
  INV_X1 U4835 ( .A(n2470), .ZN(n2462) );
  NAND2_X1 U4836 ( .A1(n2470), .A2(n2842), .ZN(n4778) );
  INV_X1 U4837 ( .A(a_13_), .ZN(n2842) );
  NAND2_X1 U4838 ( .A1(n4781), .A2(n4782), .ZN(n2470) );
  NAND2_X1 U4839 ( .A1(b_14_), .A2(n4783), .ZN(n4782) );
  NAND2_X1 U4840 ( .A1(n2437), .A2(a_14_), .ZN(n4783) );
  INV_X1 U4841 ( .A(n2416), .ZN(n2437) );
  NAND2_X1 U4842 ( .A1(n2416), .A2(n2428), .ZN(n4781) );
  INV_X1 U4843 ( .A(a_14_), .ZN(n2428) );
  NAND2_X1 U4844 ( .A1(a_15_), .A2(n2951), .ZN(n2416) );
  INV_X1 U4845 ( .A(b_15_), .ZN(n2951) );
  NOR2_X1 U4846 ( .A1(n4687), .A2(operation_1_), .ZN(n2413) );
  INV_X1 U4847 ( .A(operation_0_), .ZN(n4687) );
endmodule

