module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n307_, new_n309_, new_n310_, new_n312_, new_n313_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n325_, new_n327_, new_n328_, new_n330_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n341_, new_n343_, new_n345_, new_n346_, new_n348_, new_n349_, new_n351_, new_n353_, new_n355_, new_n356_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n392_, new_n393_, new_n395_, new_n396_, new_n398_, new_n399_, new_n401_, new_n402_, new_n404_, new_n405_, new_n406_, new_n408_, new_n410_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n427_, new_n428_, new_n429_, new_n430_, new_n432_, new_n434_, new_n435_, new_n437_, new_n438_, new_n439_, new_n440_, new_n442_, new_n443_, new_n444_, new_n446_, new_n448_, new_n449_;
  INV_X1 g000 ( .A(G1GAT), .ZN(new_n138_) );
  XOR2_X1 g001 ( .A(G155GAT), .B(KEYINPUT3), .Z(new_n139_) );
  XNOR2_X1 g002 ( .A(G141GAT), .B(KEYINPUT2), .ZN(new_n140_) );
  XNOR2_X1 g003 ( .A(new_n139_), .B(new_n140_), .ZN(new_n141_) );
  XNOR2_X1 g004 ( .A(G57GAT), .B(KEYINPUT1), .ZN(new_n142_) );
  AND2_X1 g005 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n143_) );
  XNOR2_X1 g006 ( .A(new_n142_), .B(new_n143_), .ZN(new_n144_) );
  XNOR2_X1 g007 ( .A(new_n141_), .B(new_n144_), .ZN(new_n145_) );
  XNOR2_X1 g008 ( .A(G120GAT), .B(G127GAT), .ZN(new_n146_) );
  XNOR2_X1 g009 ( .A(G113GAT), .B(KEYINPUT0), .ZN(new_n147_) );
  XNOR2_X1 g010 ( .A(new_n146_), .B(new_n147_), .ZN(new_n148_) );
  XNOR2_X1 g011 ( .A(new_n148_), .B(new_n138_), .ZN(new_n149_) );
  XNOR2_X1 g012 ( .A(new_n145_), .B(new_n149_), .ZN(new_n150_) );
  XNOR2_X1 g013 ( .A(G29GAT), .B(G134GAT), .ZN(new_n151_) );
  XOR2_X1 g014 ( .A(new_n150_), .B(new_n151_), .Z(new_n152_) );
  XOR2_X1 g015 ( .A(G85GAT), .B(G162GAT), .Z(new_n153_) );
  XNOR2_X1 g016 ( .A(new_n152_), .B(new_n153_), .ZN(new_n154_) );
  XNOR2_X1 g017 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(new_n155_) );
  XNOR2_X1 g018 ( .A(G148GAT), .B(KEYINPUT6), .ZN(new_n156_) );
  XNOR2_X1 g019 ( .A(new_n155_), .B(new_n156_), .ZN(new_n157_) );
  XOR2_X1 g020 ( .A(new_n154_), .B(new_n157_), .Z(new_n158_) );
  INV_X1 g021 ( .A(new_n158_), .ZN(new_n159_) );
  INV_X1 g022 ( .A(G197GAT), .ZN(new_n160_) );
  XNOR2_X1 g023 ( .A(G211GAT), .B(G218GAT), .ZN(new_n161_) );
  XNOR2_X1 g024 ( .A(G204GAT), .B(KEYINPUT21), .ZN(new_n162_) );
  XNOR2_X1 g025 ( .A(new_n161_), .B(new_n162_), .ZN(new_n163_) );
  XNOR2_X1 g026 ( .A(new_n163_), .B(new_n160_), .ZN(new_n164_) );
  XOR2_X1 g027 ( .A(new_n164_), .B(new_n141_), .Z(new_n165_) );
  XOR2_X1 g028 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(new_n166_) );
  XNOR2_X1 g029 ( .A(G22GAT), .B(KEYINPUT22), .ZN(new_n167_) );
  XNOR2_X1 g030 ( .A(new_n166_), .B(new_n167_), .ZN(new_n168_) );
  INV_X1 g031 ( .A(G78GAT), .ZN(new_n169_) );
  INV_X1 g032 ( .A(G106GAT), .ZN(new_n170_) );
  AND2_X1 g033 ( .A1(new_n169_), .A2(new_n170_), .ZN(new_n171_) );
  AND2_X1 g034 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n172_) );
  OR2_X1 g035 ( .A1(new_n172_), .A2(G148GAT), .ZN(new_n173_) );
  OR2_X1 g036 ( .A1(new_n173_), .A2(new_n171_), .ZN(new_n174_) );
  INV_X1 g037 ( .A(G148GAT), .ZN(new_n175_) );
  XOR2_X1 g038 ( .A(G78GAT), .B(G106GAT), .Z(new_n176_) );
  OR2_X1 g039 ( .A1(new_n176_), .A2(new_n175_), .ZN(new_n177_) );
  AND2_X1 g040 ( .A1(new_n174_), .A2(new_n177_), .ZN(new_n178_) );
  XOR2_X1 g041 ( .A(new_n178_), .B(new_n168_), .Z(new_n179_) );
  XNOR2_X1 g042 ( .A(new_n165_), .B(new_n179_), .ZN(new_n180_) );
  XNOR2_X1 g043 ( .A(G50GAT), .B(G162GAT), .ZN(new_n181_) );
  XNOR2_X1 g044 ( .A(new_n180_), .B(new_n181_), .ZN(new_n182_) );
  AND2_X1 g045 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n183_) );
  XOR2_X1 g046 ( .A(new_n182_), .B(new_n183_), .Z(new_n184_) );
  XOR2_X1 g047 ( .A(new_n148_), .B(G15GAT), .Z(new_n185_) );
  AND2_X1 g048 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n186_) );
  XOR2_X1 g049 ( .A(new_n185_), .B(new_n186_), .Z(new_n187_) );
  XOR2_X1 g050 ( .A(G176GAT), .B(G183GAT), .Z(new_n188_) );
  XNOR2_X1 g051 ( .A(G71GAT), .B(KEYINPUT20), .ZN(new_n189_) );
  XOR2_X1 g052 ( .A(new_n188_), .B(new_n189_), .Z(new_n190_) );
  XNOR2_X1 g053 ( .A(new_n187_), .B(new_n190_), .ZN(new_n191_) );
  XNOR2_X1 g054 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(new_n192_) );
  XNOR2_X1 g055 ( .A(G169GAT), .B(KEYINPUT19), .ZN(new_n193_) );
  XNOR2_X1 g056 ( .A(new_n192_), .B(new_n193_), .ZN(new_n194_) );
  XNOR2_X1 g057 ( .A(G134GAT), .B(G190GAT), .ZN(new_n195_) );
  XNOR2_X1 g058 ( .A(G43GAT), .B(G99GAT), .ZN(new_n196_) );
  XNOR2_X1 g059 ( .A(new_n195_), .B(new_n196_), .ZN(new_n197_) );
  XNOR2_X1 g060 ( .A(new_n194_), .B(new_n197_), .ZN(new_n198_) );
  XOR2_X1 g061 ( .A(new_n191_), .B(new_n198_), .Z(new_n199_) );
  AND2_X1 g062 ( .A1(new_n184_), .A2(new_n199_), .ZN(new_n200_) );
  XNOR2_X1 g063 ( .A(new_n200_), .B(KEYINPUT26), .ZN(new_n201_) );
  XOR2_X1 g064 ( .A(G36GAT), .B(G190GAT), .Z(new_n202_) );
  XNOR2_X1 g065 ( .A(new_n164_), .B(new_n202_), .ZN(new_n203_) );
  INV_X1 g066 ( .A(G92GAT), .ZN(new_n204_) );
  XNOR2_X1 g067 ( .A(G64GAT), .B(G176GAT), .ZN(new_n205_) );
  XNOR2_X1 g068 ( .A(new_n205_), .B(new_n204_), .ZN(new_n206_) );
  AND2_X1 g069 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n207_) );
  XNOR2_X1 g070 ( .A(new_n206_), .B(new_n207_), .ZN(new_n208_) );
  XOR2_X1 g071 ( .A(G8GAT), .B(G183GAT), .Z(new_n209_) );
  XOR2_X1 g072 ( .A(new_n208_), .B(new_n209_), .Z(new_n210_) );
  XNOR2_X1 g073 ( .A(new_n210_), .B(new_n203_), .ZN(new_n211_) );
  XOR2_X1 g074 ( .A(new_n211_), .B(new_n194_), .Z(new_n212_) );
  XOR2_X1 g075 ( .A(new_n212_), .B(KEYINPUT27), .Z(new_n213_) );
  AND2_X1 g076 ( .A1(new_n201_), .A2(new_n213_), .ZN(new_n214_) );
  INV_X1 g077 ( .A(new_n199_), .ZN(new_n215_) );
  INV_X1 g078 ( .A(new_n212_), .ZN(new_n216_) );
  AND2_X1 g079 ( .A1(new_n215_), .A2(new_n216_), .ZN(new_n217_) );
  OR2_X1 g080 ( .A1(new_n217_), .A2(new_n184_), .ZN(new_n218_) );
  XNOR2_X1 g081 ( .A(new_n218_), .B(KEYINPUT25), .ZN(new_n219_) );
  OR2_X1 g082 ( .A1(new_n214_), .A2(new_n219_), .ZN(new_n220_) );
  AND2_X1 g083 ( .A1(new_n220_), .A2(new_n159_), .ZN(new_n221_) );
  XOR2_X1 g084 ( .A(new_n184_), .B(KEYINPUT28), .Z(new_n222_) );
  AND2_X1 g085 ( .A1(new_n213_), .A2(new_n158_), .ZN(new_n223_) );
  AND2_X1 g086 ( .A1(new_n223_), .A2(new_n199_), .ZN(new_n224_) );
  AND2_X1 g087 ( .A1(new_n224_), .A2(new_n222_), .ZN(new_n225_) );
  OR2_X1 g088 ( .A1(new_n221_), .A2(new_n225_), .ZN(new_n226_) );
  XNOR2_X1 g089 ( .A(G106GAT), .B(G218GAT), .ZN(new_n227_) );
  XNOR2_X1 g090 ( .A(new_n151_), .B(new_n227_), .ZN(new_n228_) );
  INV_X1 g091 ( .A(G43GAT), .ZN(new_n229_) );
  INV_X1 g092 ( .A(KEYINPUT8), .ZN(new_n230_) );
  AND2_X1 g093 ( .A1(new_n229_), .A2(new_n230_), .ZN(new_n231_) );
  AND2_X1 g094 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n232_) );
  OR2_X1 g095 ( .A1(new_n232_), .A2(KEYINPUT7), .ZN(new_n233_) );
  OR2_X1 g096 ( .A1(new_n233_), .A2(new_n231_), .ZN(new_n234_) );
  INV_X1 g097 ( .A(KEYINPUT7), .ZN(new_n235_) );
  XOR2_X1 g098 ( .A(G43GAT), .B(KEYINPUT8), .Z(new_n236_) );
  OR2_X1 g099 ( .A1(new_n236_), .A2(new_n235_), .ZN(new_n237_) );
  AND2_X1 g100 ( .A1(new_n234_), .A2(new_n237_), .ZN(new_n238_) );
  INV_X1 g101 ( .A(G85GAT), .ZN(new_n239_) );
  INV_X1 g102 ( .A(G99GAT), .ZN(new_n240_) );
  AND2_X1 g103 ( .A1(new_n239_), .A2(new_n240_), .ZN(new_n241_) );
  AND2_X1 g104 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n242_) );
  OR2_X1 g105 ( .A1(new_n242_), .A2(G92GAT), .ZN(new_n243_) );
  OR2_X1 g106 ( .A1(new_n243_), .A2(new_n241_), .ZN(new_n244_) );
  XOR2_X1 g107 ( .A(G85GAT), .B(G99GAT), .Z(new_n245_) );
  OR2_X1 g108 ( .A1(new_n245_), .A2(new_n204_), .ZN(new_n246_) );
  AND2_X1 g109 ( .A1(new_n244_), .A2(new_n246_), .ZN(new_n247_) );
  XNOR2_X1 g110 ( .A(new_n238_), .B(new_n247_), .ZN(new_n248_) );
  XNOR2_X1 g111 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(new_n249_) );
  AND2_X1 g112 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n250_) );
  XNOR2_X1 g113 ( .A(new_n249_), .B(new_n250_), .ZN(new_n251_) );
  XNOR2_X1 g114 ( .A(new_n251_), .B(KEYINPUT9), .ZN(new_n252_) );
  XNOR2_X1 g115 ( .A(new_n248_), .B(new_n252_), .ZN(new_n253_) );
  XNOR2_X1 g116 ( .A(new_n253_), .B(new_n228_), .ZN(new_n254_) );
  XNOR2_X1 g117 ( .A(new_n254_), .B(new_n181_), .ZN(new_n255_) );
  XNOR2_X1 g118 ( .A(new_n255_), .B(new_n202_), .ZN(new_n256_) );
  INV_X1 g119 ( .A(new_n256_), .ZN(new_n257_) );
  XNOR2_X1 g120 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(new_n258_) );
  XNOR2_X1 g121 ( .A(G64GAT), .B(KEYINPUT15), .ZN(new_n259_) );
  XNOR2_X1 g122 ( .A(new_n258_), .B(new_n259_), .ZN(new_n260_) );
  XNOR2_X1 g123 ( .A(G78GAT), .B(G155GAT), .ZN(new_n261_) );
  XNOR2_X1 g124 ( .A(G127GAT), .B(G211GAT), .ZN(new_n262_) );
  XNOR2_X1 g125 ( .A(new_n261_), .B(new_n262_), .ZN(new_n263_) );
  XNOR2_X1 g126 ( .A(new_n260_), .B(new_n263_), .ZN(new_n264_) );
  XNOR2_X1 g127 ( .A(G15GAT), .B(G22GAT), .ZN(new_n265_) );
  XNOR2_X1 g128 ( .A(new_n265_), .B(new_n138_), .ZN(new_n266_) );
  XNOR2_X1 g129 ( .A(G57GAT), .B(G71GAT), .ZN(new_n267_) );
  XOR2_X1 g130 ( .A(new_n267_), .B(KEYINPUT13), .Z(new_n268_) );
  XNOR2_X1 g131 ( .A(new_n268_), .B(new_n266_), .ZN(new_n269_) );
  XOR2_X1 g132 ( .A(new_n269_), .B(new_n264_), .Z(new_n270_) );
  XNOR2_X1 g133 ( .A(new_n270_), .B(new_n209_), .ZN(new_n271_) );
  AND2_X1 g134 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n272_) );
  XOR2_X1 g135 ( .A(new_n271_), .B(new_n272_), .Z(new_n273_) );
  INV_X1 g136 ( .A(new_n273_), .ZN(new_n274_) );
  AND2_X1 g137 ( .A1(new_n257_), .A2(new_n274_), .ZN(new_n275_) );
  XNOR2_X1 g138 ( .A(new_n275_), .B(KEYINPUT16), .ZN(new_n276_) );
  AND2_X1 g139 ( .A1(new_n226_), .A2(new_n276_), .ZN(new_n277_) );
  INV_X1 g140 ( .A(new_n268_), .ZN(new_n278_) );
  XOR2_X1 g141 ( .A(G120GAT), .B(G204GAT), .Z(new_n279_) );
  XNOR2_X1 g142 ( .A(new_n178_), .B(new_n247_), .ZN(new_n280_) );
  XOR2_X1 g143 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(new_n281_) );
  AND2_X1 g144 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n282_) );
  XNOR2_X1 g145 ( .A(new_n281_), .B(new_n282_), .ZN(new_n283_) );
  XNOR2_X1 g146 ( .A(new_n283_), .B(KEYINPUT32), .ZN(new_n284_) );
  XNOR2_X1 g147 ( .A(new_n280_), .B(new_n284_), .ZN(new_n285_) );
  XNOR2_X1 g148 ( .A(new_n285_), .B(new_n205_), .ZN(new_n286_) );
  XNOR2_X1 g149 ( .A(new_n286_), .B(new_n279_), .ZN(new_n287_) );
  XNOR2_X1 g150 ( .A(new_n287_), .B(new_n278_), .ZN(new_n288_) );
  XNOR2_X1 g151 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(new_n289_) );
  XNOR2_X1 g152 ( .A(G8GAT), .B(G169GAT), .ZN(new_n290_) );
  XNOR2_X1 g153 ( .A(new_n289_), .B(new_n290_), .ZN(new_n291_) );
  XNOR2_X1 g154 ( .A(G113GAT), .B(G197GAT), .ZN(new_n292_) );
  XNOR2_X1 g155 ( .A(G29GAT), .B(G141GAT), .ZN(new_n293_) );
  XOR2_X1 g156 ( .A(new_n292_), .B(new_n293_), .Z(new_n294_) );
  XNOR2_X1 g157 ( .A(new_n294_), .B(new_n291_), .ZN(new_n295_) );
  XNOR2_X1 g158 ( .A(new_n238_), .B(new_n266_), .ZN(new_n296_) );
  XOR2_X1 g159 ( .A(new_n296_), .B(new_n295_), .Z(new_n297_) );
  XOR2_X1 g160 ( .A(G36GAT), .B(G50GAT), .Z(new_n298_) );
  AND2_X1 g161 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n299_) );
  XNOR2_X1 g162 ( .A(new_n298_), .B(new_n299_), .ZN(new_n300_) );
  XOR2_X1 g163 ( .A(new_n297_), .B(new_n300_), .Z(new_n301_) );
  AND2_X1 g164 ( .A1(new_n288_), .A2(new_n301_), .ZN(new_n302_) );
  AND2_X1 g165 ( .A1(new_n277_), .A2(new_n302_), .ZN(new_n303_) );
  AND2_X1 g166 ( .A1(new_n303_), .A2(new_n158_), .ZN(new_n304_) );
  XNOR2_X1 g167 ( .A(new_n304_), .B(KEYINPUT34), .ZN(new_n305_) );
  XNOR2_X1 g168 ( .A(new_n305_), .B(new_n138_), .ZN(G1324GAT) );
  AND2_X1 g169 ( .A1(new_n303_), .A2(new_n216_), .ZN(new_n307_) );
  XOR2_X1 g170 ( .A(new_n307_), .B(G8GAT), .Z(G1325GAT) );
  AND2_X1 g171 ( .A1(new_n303_), .A2(new_n215_), .ZN(new_n309_) );
  XNOR2_X1 g172 ( .A(G15GAT), .B(KEYINPUT35), .ZN(new_n310_) );
  XNOR2_X1 g173 ( .A(new_n309_), .B(new_n310_), .ZN(G1326GAT) );
  INV_X1 g174 ( .A(new_n222_), .ZN(new_n312_) );
  AND2_X1 g175 ( .A1(new_n303_), .A2(new_n312_), .ZN(new_n313_) );
  XOR2_X1 g176 ( .A(new_n313_), .B(G22GAT), .Z(G1327GAT) );
  XOR2_X1 g177 ( .A(new_n256_), .B(KEYINPUT36), .Z(new_n315_) );
  INV_X1 g178 ( .A(new_n315_), .ZN(new_n316_) );
  AND2_X1 g179 ( .A1(new_n316_), .A2(new_n273_), .ZN(new_n317_) );
  AND2_X1 g180 ( .A1(new_n226_), .A2(new_n317_), .ZN(new_n318_) );
  XOR2_X1 g181 ( .A(new_n318_), .B(KEYINPUT37), .Z(new_n319_) );
  AND2_X1 g182 ( .A1(new_n319_), .A2(new_n302_), .ZN(new_n320_) );
  XNOR2_X1 g183 ( .A(new_n320_), .B(KEYINPUT38), .ZN(new_n321_) );
  AND2_X1 g184 ( .A1(new_n321_), .A2(new_n158_), .ZN(new_n322_) );
  XNOR2_X1 g185 ( .A(G29GAT), .B(KEYINPUT39), .ZN(new_n323_) );
  XNOR2_X1 g186 ( .A(new_n322_), .B(new_n323_), .ZN(G1328GAT) );
  AND2_X1 g187 ( .A1(new_n321_), .A2(new_n216_), .ZN(new_n325_) );
  XOR2_X1 g188 ( .A(new_n325_), .B(G36GAT), .Z(G1329GAT) );
  AND2_X1 g189 ( .A1(new_n321_), .A2(new_n215_), .ZN(new_n327_) );
  XNOR2_X1 g190 ( .A(new_n327_), .B(KEYINPUT40), .ZN(new_n328_) );
  XNOR2_X1 g191 ( .A(new_n328_), .B(new_n229_), .ZN(G1330GAT) );
  AND2_X1 g192 ( .A1(new_n321_), .A2(new_n312_), .ZN(new_n330_) );
  XOR2_X1 g193 ( .A(new_n330_), .B(G50GAT), .Z(G1331GAT) );
  INV_X1 g194 ( .A(new_n301_), .ZN(new_n332_) );
  INV_X1 g195 ( .A(KEYINPUT41), .ZN(new_n333_) );
  XNOR2_X1 g196 ( .A(new_n288_), .B(new_n333_), .ZN(new_n334_) );
  INV_X1 g197 ( .A(new_n334_), .ZN(new_n335_) );
  AND2_X1 g198 ( .A1(new_n335_), .A2(new_n332_), .ZN(new_n336_) );
  AND2_X1 g199 ( .A1(new_n277_), .A2(new_n336_), .ZN(new_n337_) );
  AND2_X1 g200 ( .A1(new_n337_), .A2(new_n158_), .ZN(new_n338_) );
  XOR2_X1 g201 ( .A(G57GAT), .B(KEYINPUT42), .Z(new_n339_) );
  XNOR2_X1 g202 ( .A(new_n338_), .B(new_n339_), .ZN(G1332GAT) );
  AND2_X1 g203 ( .A1(new_n337_), .A2(new_n216_), .ZN(new_n341_) );
  XOR2_X1 g204 ( .A(new_n341_), .B(G64GAT), .Z(G1333GAT) );
  AND2_X1 g205 ( .A1(new_n337_), .A2(new_n215_), .ZN(new_n343_) );
  XOR2_X1 g206 ( .A(new_n343_), .B(G71GAT), .Z(G1334GAT) );
  AND2_X1 g207 ( .A1(new_n337_), .A2(new_n312_), .ZN(new_n345_) );
  XNOR2_X1 g208 ( .A(G78GAT), .B(KEYINPUT43), .ZN(new_n346_) );
  XNOR2_X1 g209 ( .A(new_n345_), .B(new_n346_), .ZN(G1335GAT) );
  AND2_X1 g210 ( .A1(new_n319_), .A2(new_n336_), .ZN(new_n348_) );
  AND2_X1 g211 ( .A1(new_n348_), .A2(new_n158_), .ZN(new_n349_) );
  XNOR2_X1 g212 ( .A(new_n349_), .B(new_n239_), .ZN(G1336GAT) );
  AND2_X1 g213 ( .A1(new_n348_), .A2(new_n216_), .ZN(new_n351_) );
  XNOR2_X1 g214 ( .A(new_n351_), .B(new_n204_), .ZN(G1337GAT) );
  AND2_X1 g215 ( .A1(new_n348_), .A2(new_n215_), .ZN(new_n353_) );
  XNOR2_X1 g216 ( .A(new_n353_), .B(new_n240_), .ZN(G1338GAT) );
  AND2_X1 g217 ( .A1(new_n348_), .A2(new_n312_), .ZN(new_n355_) );
  XNOR2_X1 g218 ( .A(new_n355_), .B(KEYINPUT44), .ZN(new_n356_) );
  XNOR2_X1 g219 ( .A(new_n356_), .B(new_n170_), .ZN(G1339GAT) );
  INV_X1 g220 ( .A(KEYINPUT46), .ZN(new_n358_) );
  OR2_X1 g221 ( .A1(new_n334_), .A2(new_n332_), .ZN(new_n359_) );
  AND2_X1 g222 ( .A1(new_n359_), .A2(new_n358_), .ZN(new_n360_) );
  INV_X1 g223 ( .A(new_n360_), .ZN(new_n361_) );
  OR2_X1 g224 ( .A1(new_n359_), .A2(new_n358_), .ZN(new_n362_) );
  AND2_X1 g225 ( .A1(new_n257_), .A2(new_n273_), .ZN(new_n363_) );
  AND2_X1 g226 ( .A1(new_n362_), .A2(new_n363_), .ZN(new_n364_) );
  AND2_X1 g227 ( .A1(new_n364_), .A2(new_n361_), .ZN(new_n365_) );
  INV_X1 g228 ( .A(new_n365_), .ZN(new_n366_) );
  AND2_X1 g229 ( .A1(new_n366_), .A2(KEYINPUT47), .ZN(new_n367_) );
  INV_X1 g230 ( .A(KEYINPUT47), .ZN(new_n368_) );
  AND2_X1 g231 ( .A1(new_n365_), .A2(new_n368_), .ZN(new_n369_) );
  INV_X1 g232 ( .A(KEYINPUT45), .ZN(new_n370_) );
  OR2_X1 g233 ( .A1(new_n315_), .A2(new_n273_), .ZN(new_n371_) );
  INV_X1 g234 ( .A(new_n371_), .ZN(new_n372_) );
  OR2_X1 g235 ( .A1(new_n372_), .A2(new_n370_), .ZN(new_n373_) );
  OR2_X1 g236 ( .A1(new_n371_), .A2(KEYINPUT45), .ZN(new_n374_) );
  AND2_X1 g237 ( .A1(new_n288_), .A2(new_n332_), .ZN(new_n375_) );
  AND2_X1 g238 ( .A1(new_n374_), .A2(new_n375_), .ZN(new_n376_) );
  AND2_X1 g239 ( .A1(new_n376_), .A2(new_n373_), .ZN(new_n377_) );
  OR2_X1 g240 ( .A1(new_n369_), .A2(new_n377_), .ZN(new_n378_) );
  OR2_X1 g241 ( .A1(new_n378_), .A2(new_n367_), .ZN(new_n379_) );
  INV_X1 g242 ( .A(new_n379_), .ZN(new_n380_) );
  AND2_X1 g243 ( .A1(new_n380_), .A2(KEYINPUT48), .ZN(new_n381_) );
  INV_X1 g244 ( .A(new_n381_), .ZN(new_n382_) );
  INV_X1 g245 ( .A(KEYINPUT48), .ZN(new_n383_) );
  AND2_X1 g246 ( .A1(new_n379_), .A2(new_n383_), .ZN(new_n384_) );
  INV_X1 g247 ( .A(new_n384_), .ZN(new_n385_) );
  AND2_X1 g248 ( .A1(new_n385_), .A2(new_n223_), .ZN(new_n386_) );
  AND2_X1 g249 ( .A1(new_n386_), .A2(new_n382_), .ZN(new_n387_) );
  AND2_X1 g250 ( .A1(new_n222_), .A2(new_n215_), .ZN(new_n388_) );
  AND2_X1 g251 ( .A1(new_n387_), .A2(new_n388_), .ZN(new_n389_) );
  AND2_X1 g252 ( .A1(new_n389_), .A2(new_n301_), .ZN(new_n390_) );
  XOR2_X1 g253 ( .A(new_n390_), .B(G113GAT), .Z(G1340GAT) );
  AND2_X1 g254 ( .A1(new_n389_), .A2(new_n335_), .ZN(new_n392_) );
  XNOR2_X1 g255 ( .A(G120GAT), .B(KEYINPUT49), .ZN(new_n393_) );
  XNOR2_X1 g256 ( .A(new_n392_), .B(new_n393_), .ZN(G1341GAT) );
  AND2_X1 g257 ( .A1(new_n389_), .A2(new_n274_), .ZN(new_n395_) );
  XNOR2_X1 g258 ( .A(new_n395_), .B(KEYINPUT50), .ZN(new_n396_) );
  XOR2_X1 g259 ( .A(new_n396_), .B(G127GAT), .Z(G1342GAT) );
  AND2_X1 g260 ( .A1(new_n389_), .A2(new_n256_), .ZN(new_n398_) );
  XNOR2_X1 g261 ( .A(G134GAT), .B(KEYINPUT51), .ZN(new_n399_) );
  XNOR2_X1 g262 ( .A(new_n398_), .B(new_n399_), .ZN(G1343GAT) );
  AND2_X1 g263 ( .A1(new_n387_), .A2(new_n201_), .ZN(new_n401_) );
  AND2_X1 g264 ( .A1(new_n401_), .A2(new_n301_), .ZN(new_n402_) );
  XOR2_X1 g265 ( .A(new_n402_), .B(G141GAT), .Z(G1344GAT) );
  AND2_X1 g266 ( .A1(new_n401_), .A2(new_n335_), .ZN(new_n404_) );
  XOR2_X1 g267 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(new_n405_) );
  XNOR2_X1 g268 ( .A(new_n404_), .B(new_n405_), .ZN(new_n406_) );
  XNOR2_X1 g269 ( .A(new_n406_), .B(new_n175_), .ZN(G1345GAT) );
  AND2_X1 g270 ( .A1(new_n401_), .A2(new_n274_), .ZN(new_n408_) );
  XOR2_X1 g271 ( .A(new_n408_), .B(G155GAT), .Z(G1346GAT) );
  AND2_X1 g272 ( .A1(new_n401_), .A2(new_n256_), .ZN(new_n410_) );
  XOR2_X1 g273 ( .A(new_n410_), .B(G162GAT), .Z(G1347GAT) );
  INV_X1 g274 ( .A(KEYINPUT55), .ZN(new_n412_) );
  INV_X1 g275 ( .A(new_n184_), .ZN(new_n413_) );
  INV_X1 g276 ( .A(KEYINPUT54), .ZN(new_n414_) );
  OR2_X1 g277 ( .A1(new_n384_), .A2(new_n212_), .ZN(new_n415_) );
  OR2_X1 g278 ( .A1(new_n415_), .A2(new_n381_), .ZN(new_n416_) );
  INV_X1 g279 ( .A(new_n416_), .ZN(new_n417_) );
  OR2_X1 g280 ( .A1(new_n417_), .A2(new_n414_), .ZN(new_n418_) );
  OR2_X1 g281 ( .A1(new_n416_), .A2(KEYINPUT54), .ZN(new_n419_) );
  AND2_X1 g282 ( .A1(new_n419_), .A2(new_n159_), .ZN(new_n420_) );
  AND2_X1 g283 ( .A1(new_n420_), .A2(new_n418_), .ZN(new_n421_) );
  AND2_X1 g284 ( .A1(new_n421_), .A2(new_n413_), .ZN(new_n422_) );
  XNOR2_X1 g285 ( .A(new_n422_), .B(new_n412_), .ZN(new_n423_) );
  AND2_X1 g286 ( .A1(new_n423_), .A2(new_n215_), .ZN(new_n424_) );
  AND2_X1 g287 ( .A1(new_n424_), .A2(new_n301_), .ZN(new_n425_) );
  XOR2_X1 g288 ( .A(new_n425_), .B(G169GAT), .Z(G1348GAT) );
  INV_X1 g289 ( .A(G176GAT), .ZN(new_n427_) );
  AND2_X1 g290 ( .A1(new_n424_), .A2(new_n335_), .ZN(new_n428_) );
  XOR2_X1 g291 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(new_n429_) );
  XNOR2_X1 g292 ( .A(new_n428_), .B(new_n429_), .ZN(new_n430_) );
  XNOR2_X1 g293 ( .A(new_n430_), .B(new_n427_), .ZN(G1349GAT) );
  AND2_X1 g294 ( .A1(new_n424_), .A2(new_n274_), .ZN(new_n432_) );
  XOR2_X1 g295 ( .A(new_n432_), .B(G183GAT), .Z(G1350GAT) );
  AND2_X1 g296 ( .A1(new_n424_), .A2(new_n256_), .ZN(new_n434_) );
  XOR2_X1 g297 ( .A(G190GAT), .B(KEYINPUT58), .Z(new_n435_) );
  XNOR2_X1 g298 ( .A(new_n434_), .B(new_n435_), .ZN(G1351GAT) );
  AND2_X1 g299 ( .A1(new_n421_), .A2(new_n201_), .ZN(new_n437_) );
  AND2_X1 g300 ( .A1(new_n437_), .A2(new_n301_), .ZN(new_n438_) );
  XOR2_X1 g301 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(new_n439_) );
  XNOR2_X1 g302 ( .A(new_n438_), .B(new_n439_), .ZN(new_n440_) );
  XNOR2_X1 g303 ( .A(new_n440_), .B(new_n160_), .ZN(G1352GAT) );
  INV_X1 g304 ( .A(new_n288_), .ZN(new_n442_) );
  AND2_X1 g305 ( .A1(new_n437_), .A2(new_n442_), .ZN(new_n443_) );
  XNOR2_X1 g306 ( .A(G204GAT), .B(KEYINPUT61), .ZN(new_n444_) );
  XNOR2_X1 g307 ( .A(new_n443_), .B(new_n444_), .ZN(G1353GAT) );
  AND2_X1 g308 ( .A1(new_n437_), .A2(new_n274_), .ZN(new_n446_) );
  XOR2_X1 g309 ( .A(new_n446_), .B(G211GAT), .Z(G1354GAT) );
  AND2_X1 g310 ( .A1(new_n437_), .A2(new_n316_), .ZN(new_n448_) );
  XNOR2_X1 g311 ( .A(new_n448_), .B(KEYINPUT62), .ZN(new_n449_) );
  XOR2_X1 g312 ( .A(new_n449_), .B(G218GAT), .Z(G1355GAT) );
endmodule


