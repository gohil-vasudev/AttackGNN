module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n173_, new_n220_, new_n419_, new_n214_, new_n451_, new_n424_, new_n114_, new_n188_, new_n240_, new_n413_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n462_, new_n317_, new_n344_, new_n287_, new_n427_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n110_, new_n315_, new_n124_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n350_, new_n117_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n150_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n351_, new_n325_, new_n180_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n423_, new_n205_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n256_, new_n452_, new_n381_, new_n388_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n436_, new_n397_, new_n399_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n161_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n113_, new_n371_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n460_, new_n130_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n126_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n125_, new_n145_, new_n253_, new_n403_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n182_, new_n407_, new_n480_, new_n151_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n428_, new_n199_, new_n146_, new_n360_, new_n302_, new_n191_, new_n225_, new_n387_, new_n476_, new_n112_, new_n121_, new_n415_, new_n221_, new_n243_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n459_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n340_, new_n147_, new_n285_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n332_, new_n453_, new_n163_, new_n148_, new_n440_, new_n122_, new_n111_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n115_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n134_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n278_, new_n304_, new_n217_, new_n269_, new_n129_, new_n412_, new_n327_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n128_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n455_, new_n120_, new_n406_, new_n356_, new_n229_, new_n464_, new_n204_, new_n181_, new_n135_, new_n405_;

not g000 ( new_n108_, N69 );
not g001 ( new_n109_, keyIn_0_9 );
or g002 ( new_n110_, new_n109_, N63 );
or g003 ( new_n111_, new_n110_, new_n108_ );
not g004 ( new_n112_, N63 );
and g005 ( new_n113_, new_n112_, N69 );
or g006 ( new_n114_, new_n113_, keyIn_0_9 );
and g007 ( new_n115_, new_n111_, new_n114_ );
not g008 ( new_n116_, keyIn_0_5 );
not g009 ( new_n117_, N89 );
and g010 ( new_n118_, new_n116_, new_n117_ );
not g011 ( new_n119_, N95 );
and g012 ( new_n120_, keyIn_0_5, N89 );
or g013 ( new_n121_, new_n120_, new_n119_ );
or g014 ( new_n122_, new_n121_, new_n118_ );
not g015 ( new_n123_, N30 );
or g016 ( new_n124_, new_n123_, N24 );
and g017 ( new_n125_, new_n124_, keyIn_0_8 );
not g018 ( new_n126_, keyIn_0_8 );
not g019 ( new_n127_, N24 );
and g020 ( new_n128_, new_n126_, new_n127_ );
and g021 ( new_n129_, new_n128_, N30 );
or g022 ( new_n130_, new_n125_, new_n129_ );
and g023 ( new_n131_, new_n130_, new_n122_ );
and g024 ( new_n132_, new_n131_, new_n115_ );
not g025 ( new_n133_, keyIn_0_7 );
not g026 ( new_n134_, N17 );
or g027 ( new_n135_, new_n134_, N11 );
and g028 ( new_n136_, new_n135_, new_n133_ );
not g029 ( new_n137_, N11 );
and g030 ( new_n138_, new_n137_, keyIn_0_7 );
and g031 ( new_n139_, new_n138_, N17 );
or g032 ( new_n140_, new_n136_, new_n139_ );
not g033 ( new_n141_, N56 );
or g034 ( new_n142_, new_n141_, N50 );
not g035 ( new_n143_, N82 );
or g036 ( new_n144_, new_n143_, N76 );
not g037 ( new_n145_, N4 );
or g038 ( new_n146_, new_n145_, N1 );
and g039 ( new_n147_, new_n144_, new_n146_ );
and g040 ( new_n148_, new_n147_, new_n142_ );
and g041 ( new_n149_, new_n140_, new_n148_ );
not g042 ( new_n150_, N43 );
xor g043 ( new_n151_, keyIn_0_2, N37 );
or g044 ( new_n152_, new_n151_, new_n150_ );
not g045 ( new_n153_, N108 );
not g046 ( new_n154_, keyIn_0_10 );
or g047 ( new_n155_, new_n154_, N102 );
or g048 ( new_n156_, new_n155_, new_n153_ );
not g049 ( new_n157_, N102 );
and g050 ( new_n158_, new_n157_, N108 );
or g051 ( new_n159_, new_n158_, keyIn_0_10 );
and g052 ( new_n160_, new_n156_, new_n159_ );
and g053 ( new_n161_, new_n160_, new_n152_ );
and g054 ( new_n162_, new_n149_, new_n161_ );
and g055 ( new_n163_, new_n132_, new_n162_ );
xor g056 ( N223, new_n163_, keyIn_0_20 );
xnor g057 ( new_n165_, new_n163_, keyIn_0_18 );
xnor g058 ( new_n166_, new_n165_, new_n140_ );
xor g059 ( new_n167_, new_n166_, keyIn_0_21 );
not g060 ( new_n168_, N21 );
and g061 ( new_n169_, new_n168_, N17 );
and g062 ( new_n170_, new_n167_, new_n169_ );
xor g063 ( new_n171_, new_n170_, keyIn_0_29 );
xnor g064 ( new_n172_, new_n165_, new_n144_ );
not g065 ( new_n173_, N86 );
and g066 ( new_n174_, new_n173_, N82 );
not g067 ( new_n175_, new_n174_ );
or g068 ( new_n176_, new_n172_, new_n175_ );
not g069 ( new_n177_, new_n115_ );
or g070 ( new_n178_, new_n165_, new_n177_ );
not g071 ( new_n179_, keyIn_0_18 );
and g072 ( new_n180_, new_n177_, new_n179_ );
not g073 ( new_n181_, new_n180_ );
and g074 ( new_n182_, new_n178_, new_n181_ );
not g075 ( new_n183_, N73 );
xnor g076 ( new_n184_, keyIn_0_4, N69 );
and g077 ( new_n185_, new_n184_, new_n183_ );
not g078 ( new_n186_, new_n185_ );
or g079 ( new_n187_, new_n182_, new_n186_ );
and g080 ( new_n188_, new_n187_, new_n176_ );
xnor g081 ( new_n189_, new_n165_, new_n142_ );
or g082 ( new_n190_, new_n141_, N60 );
xor g083 ( new_n191_, new_n190_, keyIn_0_13 );
or g084 ( new_n192_, new_n189_, new_n191_ );
not g085 ( new_n193_, new_n130_ );
or g086 ( new_n194_, new_n165_, new_n193_ );
and g087 ( new_n195_, new_n193_, new_n179_ );
not g088 ( new_n196_, new_n195_ );
and g089 ( new_n197_, new_n194_, new_n196_ );
not g090 ( new_n198_, N34 );
xor g091 ( new_n199_, keyIn_0_1, N30 );
not g092 ( new_n200_, new_n199_ );
and g093 ( new_n201_, new_n200_, new_n198_ );
not g094 ( new_n202_, new_n201_ );
or g095 ( new_n203_, new_n197_, new_n202_ );
and g096 ( new_n204_, new_n203_, new_n192_ );
xnor g097 ( new_n205_, new_n165_, new_n122_ );
or g098 ( new_n206_, new_n119_, N99 );
or g099 ( new_n207_, new_n205_, new_n206_ );
xnor g100 ( new_n208_, new_n165_, new_n160_ );
or g101 ( new_n209_, new_n153_, N112 );
xor g102 ( new_n210_, new_n209_, keyIn_0_17 );
not g103 ( new_n211_, new_n210_ );
or g104 ( new_n212_, new_n208_, new_n211_ );
and g105 ( new_n213_, new_n207_, new_n212_ );
and g106 ( new_n214_, new_n204_, new_n213_ );
and g107 ( new_n215_, new_n214_, new_n188_ );
xor g108 ( new_n216_, new_n165_, new_n146_ );
not g109 ( new_n217_, N8 );
xor g110 ( new_n218_, keyIn_0_0, N4 );
and g111 ( new_n219_, new_n218_, new_n217_ );
xnor g112 ( new_n220_, new_n219_, keyIn_0_6 );
and g113 ( new_n221_, new_n216_, new_n220_ );
xnor g114 ( new_n222_, new_n221_, keyIn_0_27 );
xor g115 ( new_n223_, new_n165_, new_n152_ );
not g116 ( new_n224_, N47 );
xor g117 ( new_n225_, keyIn_0_3, N43 );
and g118 ( new_n226_, new_n225_, new_n224_ );
xnor g119 ( new_n227_, new_n226_, keyIn_0_12 );
and g120 ( new_n228_, new_n223_, new_n227_ );
xnor g121 ( new_n229_, new_n228_, keyIn_0_30 );
and g122 ( new_n230_, new_n222_, new_n229_ );
and g123 ( new_n231_, new_n215_, new_n230_ );
and g124 ( new_n232_, new_n231_, new_n171_ );
xnor g125 ( new_n233_, new_n232_, keyIn_0_32 );
xnor g126 ( N329, new_n233_, keyIn_0_38 );
not g127 ( new_n235_, keyIn_0_42 );
not g128 ( new_n236_, keyIn_0_37 );
xnor g129 ( new_n237_, new_n233_, new_n236_ );
xor g130 ( new_n238_, new_n237_, new_n187_ );
xnor g131 ( new_n239_, new_n238_, new_n235_ );
not g132 ( new_n240_, new_n182_ );
not g133 ( new_n241_, N79 );
and g134 ( new_n242_, new_n184_, new_n241_ );
xor g135 ( new_n243_, new_n242_, keyIn_0_14 );
and g136 ( new_n244_, new_n240_, new_n243_ );
xnor g137 ( new_n245_, new_n244_, keyIn_0_35 );
not g138 ( new_n246_, new_n245_ );
and g139 ( new_n247_, new_n239_, new_n246_ );
not g140 ( new_n248_, new_n247_ );
or g141 ( new_n249_, new_n248_, keyIn_0_46 );
not g142 ( new_n250_, keyIn_0_46 );
or g143 ( new_n251_, new_n247_, new_n250_ );
not g144 ( new_n252_, new_n171_ );
xnor g145 ( new_n253_, new_n237_, new_n252_ );
not g146 ( new_n254_, new_n253_ );
and g147 ( new_n255_, new_n254_, keyIn_0_40 );
not g148 ( new_n256_, keyIn_0_40 );
and g149 ( new_n257_, new_n253_, new_n256_ );
not g150 ( new_n258_, N27 );
and g151 ( new_n259_, new_n258_, N17 );
and g152 ( new_n260_, new_n167_, new_n259_ );
xnor g153 ( new_n261_, new_n260_, keyIn_0_33 );
or g154 ( new_n262_, new_n257_, new_n261_ );
or g155 ( new_n263_, new_n262_, new_n255_ );
xor g156 ( new_n264_, new_n237_, new_n192_ );
or g157 ( new_n265_, new_n141_, N66 );
or g158 ( new_n266_, new_n189_, new_n265_ );
or g159 ( new_n267_, new_n264_, new_n266_ );
not g160 ( new_n268_, new_n176_ );
xnor g161 ( new_n269_, new_n237_, new_n268_ );
not g162 ( new_n270_, N92 );
and g163 ( new_n271_, new_n270_, N82 );
xnor g164 ( new_n272_, new_n271_, keyIn_0_15 );
or g165 ( new_n273_, new_n172_, new_n272_ );
xnor g166 ( new_n274_, new_n273_, keyIn_0_36 );
or g167 ( new_n275_, new_n269_, new_n274_ );
not g168 ( new_n276_, new_n203_ );
xnor g169 ( new_n277_, new_n237_, new_n276_ );
or g170 ( new_n278_, new_n199_, N40 );
xor g171 ( new_n279_, new_n278_, keyIn_0_11 );
or g172 ( new_n280_, new_n197_, new_n279_ );
xnor g173 ( new_n281_, new_n280_, keyIn_0_34 );
or g174 ( new_n282_, new_n277_, new_n281_ );
and g175 ( new_n283_, new_n275_, new_n282_ );
and g176 ( new_n284_, new_n283_, new_n267_ );
and g177 ( new_n285_, new_n263_, new_n284_ );
and g178 ( new_n286_, new_n285_, new_n251_ );
and g179 ( new_n287_, new_n286_, new_n249_ );
xnor g180 ( new_n288_, new_n237_, new_n229_ );
xnor g181 ( new_n289_, new_n288_, keyIn_0_41 );
not g182 ( new_n290_, N53 );
and g183 ( new_n291_, new_n225_, new_n290_ );
and g184 ( new_n292_, new_n223_, new_n291_ );
and g185 ( new_n293_, new_n289_, new_n292_ );
xnor g186 ( new_n294_, new_n293_, keyIn_0_45 );
xor g187 ( new_n295_, new_n237_, new_n207_ );
or g188 ( new_n296_, new_n119_, N105 );
xor g189 ( new_n297_, new_n296_, keyIn_0_16 );
or g190 ( new_n298_, new_n205_, new_n297_ );
or g191 ( new_n299_, new_n295_, new_n298_ );
xor g192 ( new_n300_, new_n299_, keyIn_0_47 );
xnor g193 ( new_n301_, new_n237_, new_n212_ );
not g194 ( new_n302_, new_n301_ );
and g195 ( new_n303_, new_n302_, keyIn_0_43 );
not g196 ( new_n304_, keyIn_0_43 );
and g197 ( new_n305_, new_n301_, new_n304_ );
or g198 ( new_n306_, new_n153_, N115 );
or g199 ( new_n307_, new_n208_, new_n306_ );
xnor g200 ( new_n308_, new_n307_, keyIn_0_31 );
or g201 ( new_n309_, new_n305_, new_n308_ );
or g202 ( new_n310_, new_n309_, new_n303_ );
xnor g203 ( new_n311_, new_n237_, new_n222_ );
not g204 ( new_n312_, new_n311_ );
and g205 ( new_n313_, new_n312_, keyIn_0_39 );
not g206 ( new_n314_, keyIn_0_39 );
and g207 ( new_n315_, new_n311_, new_n314_ );
not g208 ( new_n316_, N14 );
and g209 ( new_n317_, new_n218_, new_n316_ );
and g210 ( new_n318_, new_n216_, new_n317_ );
xor g211 ( new_n319_, new_n318_, keyIn_0_28 );
or g212 ( new_n320_, new_n315_, new_n319_ );
or g213 ( new_n321_, new_n320_, new_n313_ );
and g214 ( new_n322_, new_n310_, new_n321_ );
and g215 ( new_n323_, new_n322_, new_n300_ );
and g216 ( new_n324_, new_n323_, new_n294_ );
and g217 ( new_n325_, new_n324_, new_n287_ );
xnor g218 ( N370, new_n325_, keyIn_0_48 );
not g219 ( new_n327_, keyIn_0_49 );
not g220 ( new_n328_, keyIn_0_48 );
xnor g221 ( new_n329_, new_n325_, new_n328_ );
and g222 ( new_n330_, new_n329_, new_n327_ );
not g223 ( new_n331_, new_n330_ );
or g224 ( new_n332_, new_n329_, new_n327_ );
and g225 ( new_n333_, new_n332_, N105 );
and g226 ( new_n334_, new_n333_, new_n331_ );
xnor g227 ( new_n335_, new_n334_, keyIn_0_52 );
not g228 ( new_n336_, N99 );
or g229 ( new_n337_, new_n233_, new_n336_ );
xor g230 ( new_n338_, new_n163_, keyIn_0_19 );
or g231 ( new_n339_, new_n338_, new_n117_ );
and g232 ( new_n340_, new_n339_, N95 );
and g233 ( new_n341_, new_n337_, new_n340_ );
and g234 ( new_n342_, new_n335_, new_n341_ );
xnor g235 ( new_n343_, new_n342_, keyIn_0_55 );
and g236 ( new_n344_, new_n332_, N66 );
and g237 ( new_n345_, new_n344_, new_n331_ );
not g238 ( new_n346_, new_n345_ );
and g239 ( new_n347_, new_n346_, keyIn_0_50 );
not g240 ( new_n348_, keyIn_0_50 );
and g241 ( new_n349_, new_n345_, new_n348_ );
not g242 ( new_n350_, new_n233_ );
and g243 ( new_n351_, new_n350_, N60 );
not g244 ( new_n352_, new_n351_ );
not g245 ( new_n353_, keyIn_0_24 );
not g246 ( new_n354_, new_n338_ );
and g247 ( new_n355_, new_n354_, N50 );
and g248 ( new_n356_, new_n355_, new_n353_ );
not g249 ( new_n357_, new_n356_ );
or g250 ( new_n358_, new_n355_, new_n353_ );
and g251 ( new_n359_, new_n358_, N56 );
and g252 ( new_n360_, new_n359_, new_n357_ );
and g253 ( new_n361_, new_n352_, new_n360_ );
not g254 ( new_n362_, new_n361_ );
or g255 ( new_n363_, new_n349_, new_n362_ );
or g256 ( new_n364_, new_n363_, new_n347_ );
and g257 ( new_n365_, new_n332_, N53 );
and g258 ( new_n366_, new_n365_, new_n331_ );
and g259 ( new_n367_, new_n350_, N47 );
and g260 ( new_n368_, new_n354_, N37 );
xnor g261 ( new_n369_, new_n368_, keyIn_0_23 );
or g262 ( new_n370_, new_n369_, new_n150_ );
or g263 ( new_n371_, new_n367_, new_n370_ );
or g264 ( new_n372_, new_n366_, new_n371_ );
and g265 ( new_n373_, new_n364_, new_n372_ );
and g266 ( new_n374_, new_n332_, N79 );
and g267 ( new_n375_, new_n374_, new_n331_ );
xnor g268 ( new_n376_, new_n375_, keyIn_0_51 );
and g269 ( new_n377_, new_n350_, N73 );
not g270 ( new_n378_, new_n377_ );
not g271 ( new_n379_, keyIn_0_25 );
and g272 ( new_n380_, new_n354_, N63 );
and g273 ( new_n381_, new_n380_, new_n379_ );
not g274 ( new_n382_, new_n381_ );
or g275 ( new_n383_, new_n380_, new_n379_ );
and g276 ( new_n384_, new_n383_, N69 );
and g277 ( new_n385_, new_n384_, new_n382_ );
and g278 ( new_n386_, new_n378_, new_n385_ );
not g279 ( new_n387_, new_n386_ );
or g280 ( new_n388_, new_n376_, new_n387_ );
and g281 ( new_n389_, new_n332_, N40 );
and g282 ( new_n390_, new_n389_, new_n331_ );
and g283 ( new_n391_, new_n350_, N34 );
and g284 ( new_n392_, new_n354_, N24 );
or g285 ( new_n393_, new_n392_, new_n123_ );
or g286 ( new_n394_, new_n391_, new_n393_ );
or g287 ( new_n395_, new_n390_, new_n394_ );
and g288 ( new_n396_, new_n332_, N27 );
and g289 ( new_n397_, new_n396_, new_n331_ );
and g290 ( new_n398_, new_n350_, N21 );
not g291 ( new_n399_, new_n398_ );
not g292 ( new_n400_, keyIn_0_22 );
and g293 ( new_n401_, new_n354_, N11 );
and g294 ( new_n402_, new_n401_, new_n400_ );
not g295 ( new_n403_, new_n402_ );
or g296 ( new_n404_, new_n401_, new_n400_ );
and g297 ( new_n405_, new_n404_, N17 );
and g298 ( new_n406_, new_n405_, new_n403_ );
and g299 ( new_n407_, new_n399_, new_n406_ );
not g300 ( new_n408_, new_n407_ );
or g301 ( new_n409_, new_n397_, new_n408_ );
and g302 ( new_n410_, new_n395_, new_n409_ );
and g303 ( new_n411_, new_n388_, new_n410_ );
and g304 ( new_n412_, N370, keyIn_0_49 );
or g305 ( new_n413_, new_n412_, new_n270_ );
or g306 ( new_n414_, new_n413_, new_n330_ );
or g307 ( new_n415_, new_n233_, new_n173_ );
and g308 ( new_n416_, new_n354_, N76 );
not g309 ( new_n417_, new_n416_ );
or g310 ( new_n418_, new_n417_, keyIn_0_26 );
not g311 ( new_n419_, keyIn_0_26 );
or g312 ( new_n420_, new_n416_, new_n419_ );
and g313 ( new_n421_, new_n420_, N82 );
and g314 ( new_n422_, new_n421_, new_n418_ );
and g315 ( new_n423_, new_n415_, new_n422_ );
and g316 ( new_n424_, new_n414_, new_n423_ );
xnor g317 ( new_n425_, new_n424_, keyIn_0_54 );
not g318 ( new_n426_, new_n425_ );
and g319 ( new_n427_, new_n332_, N115 );
and g320 ( new_n428_, new_n427_, new_n331_ );
and g321 ( new_n429_, new_n350_, N112 );
xor g322 ( new_n430_, new_n429_, keyIn_0_44 );
and g323 ( new_n431_, new_n354_, N102 );
or g324 ( new_n432_, new_n431_, new_n153_ );
or g325 ( new_n433_, new_n430_, new_n432_ );
or g326 ( new_n434_, new_n428_, new_n433_ );
xnor g327 ( new_n435_, new_n434_, keyIn_0_56 );
and g328 ( new_n436_, new_n426_, new_n435_ );
and g329 ( new_n437_, new_n436_, new_n411_ );
and g330 ( new_n438_, new_n437_, new_n373_ );
and g331 ( new_n439_, new_n438_, new_n343_ );
xnor g332 ( new_n440_, new_n439_, keyIn_0_58 );
and g333 ( new_n441_, new_n332_, N14 );
and g334 ( new_n442_, new_n441_, new_n331_ );
and g335 ( new_n443_, new_n350_, N8 );
and g336 ( new_n444_, new_n354_, N1 );
or g337 ( new_n445_, new_n444_, new_n145_ );
or g338 ( new_n446_, new_n443_, new_n445_ );
or g339 ( new_n447_, new_n442_, new_n446_ );
xnor g340 ( new_n448_, new_n447_, keyIn_0_53 );
xnor g341 ( new_n449_, new_n448_, keyIn_0_57 );
and g342 ( N421, new_n440_, new_n449_ );
not g343 ( new_n451_, new_n372_ );
and g344 ( new_n452_, new_n451_, new_n395_ );
xnor g345 ( new_n453_, new_n452_, keyIn_0_60 );
not g346 ( new_n454_, new_n453_ );
and g347 ( new_n455_, new_n364_, new_n410_ );
and g348 ( new_n456_, new_n454_, new_n455_ );
xor g349 ( N430, new_n456_, keyIn_0_62 );
not g350 ( new_n458_, keyIn_0_61 );
not g351 ( new_n459_, keyIn_0_59 );
and g352 ( new_n460_, new_n425_, new_n459_ );
not g353 ( new_n461_, new_n460_ );
or g354 ( new_n462_, new_n425_, new_n459_ );
and g355 ( new_n463_, new_n373_, new_n462_ );
and g356 ( new_n464_, new_n463_, new_n461_ );
not g357 ( new_n465_, new_n464_ );
or g358 ( new_n466_, new_n465_, new_n458_ );
or g359 ( new_n467_, new_n464_, keyIn_0_61 );
not g360 ( new_n468_, new_n373_ );
not g361 ( new_n469_, new_n395_ );
or g362 ( new_n470_, new_n388_, new_n469_ );
or g363 ( new_n471_, new_n468_, new_n470_ );
and g364 ( new_n472_, new_n471_, new_n410_ );
and g365 ( new_n473_, new_n467_, new_n472_ );
and g366 ( new_n474_, new_n473_, new_n466_ );
xnor g367 ( N431, new_n474_, keyIn_0_63 );
not g368 ( new_n476_, new_n343_ );
and g369 ( new_n477_, new_n372_, new_n395_ );
and g370 ( new_n478_, new_n426_, new_n477_ );
and g371 ( new_n479_, new_n476_, new_n478_ );
not g372 ( new_n480_, new_n471_ );
not g373 ( new_n481_, new_n409_ );
or g374 ( new_n482_, new_n453_, new_n481_ );
or g375 ( new_n483_, new_n480_, new_n482_ );
or g376 ( N432, new_n483_, new_n479_ );
endmodule