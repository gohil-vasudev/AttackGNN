module add_mul_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, 
        a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, 
        a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, 
        b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, 
        b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, 
        b_28_, b_29_, b_30_, b_31_, operation, Result_0_, Result_1_, Result_2_, 
        Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, 
        Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, 
        Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, 
        Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, 
        Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, Result_32_, 
        Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, Result_38_, 
        Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, Result_44_, 
        Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, Result_50_, 
        Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, Result_56_, 
        Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, Result_62_, 
        Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963;

  AND2_X1 U7512 ( .A1(operation), .A2(n7448), .ZN(Result_9_) );
  XOR2_X1 U7513 ( .A(n7449), .B(n7450), .Z(n7448) );
  AND2_X1 U7514 ( .A1(n7451), .A2(n7452), .ZN(n7450) );
  OR2_X1 U7515 ( .A1(n7453), .A2(n7454), .ZN(n7452) );
  AND2_X1 U7516 ( .A1(n7455), .A2(n7456), .ZN(n7454) );
  INV_X1 U7517 ( .A(n7457), .ZN(n7451) );
  AND2_X1 U7518 ( .A1(n7458), .A2(operation), .ZN(Result_8_) );
  XOR2_X1 U7519 ( .A(n7459), .B(n7460), .Z(n7458) );
  AND2_X1 U7520 ( .A1(operation), .A2(n7461), .ZN(Result_7_) );
  XOR2_X1 U7521 ( .A(n7462), .B(n7463), .Z(n7461) );
  AND2_X1 U7522 ( .A1(n7464), .A2(n7465), .ZN(n7463) );
  OR2_X1 U7523 ( .A1(n7466), .A2(n7467), .ZN(n7465) );
  AND2_X1 U7524 ( .A1(n7468), .A2(n7469), .ZN(n7467) );
  INV_X1 U7525 ( .A(n7470), .ZN(n7464) );
  AND2_X1 U7526 ( .A1(n7471), .A2(operation), .ZN(Result_6_) );
  XOR2_X1 U7527 ( .A(n7472), .B(n7473), .Z(n7471) );
  OR2_X1 U7528 ( .A1(n7474), .A2(n7475), .ZN(Result_63_) );
  AND2_X1 U7529 ( .A1(n7476), .A2(operation), .ZN(n7475) );
  AND2_X1 U7530 ( .A1(n7477), .A2(n7478), .ZN(n7474) );
  XNOR2_X1 U7531 ( .A(n7479), .B(a_31_), .ZN(n7477) );
  OR2_X1 U7532 ( .A1(n7480), .A2(n7481), .ZN(Result_62_) );
  AND2_X1 U7533 ( .A1(n7482), .A2(n7478), .ZN(n7481) );
  XOR2_X1 U7534 ( .A(n7476), .B(n7483), .Z(n7482) );
  XNOR2_X1 U7535 ( .A(n7484), .B(a_30_), .ZN(n7483) );
  AND2_X1 U7536 ( .A1(operation), .A2(n7485), .ZN(n7480) );
  OR2_X1 U7537 ( .A1(n7486), .A2(n7487), .ZN(n7485) );
  AND2_X1 U7538 ( .A1(b_31_), .A2(n7488), .ZN(n7487) );
  OR2_X1 U7539 ( .A1(n7489), .A2(n7490), .ZN(n7488) );
  AND2_X1 U7540 ( .A1(a_30_), .A2(n7484), .ZN(n7489) );
  AND2_X1 U7541 ( .A1(b_30_), .A2(n7491), .ZN(n7486) );
  OR2_X1 U7542 ( .A1(n7492), .A2(n7493), .ZN(n7491) );
  AND2_X1 U7543 ( .A1(a_31_), .A2(n7479), .ZN(n7492) );
  OR2_X1 U7544 ( .A1(n7494), .A2(n7495), .ZN(Result_61_) );
  AND2_X1 U7545 ( .A1(n7496), .A2(n7478), .ZN(n7495) );
  OR2_X1 U7546 ( .A1(n7497), .A2(n7498), .ZN(n7496) );
  AND2_X1 U7547 ( .A1(n7499), .A2(n7500), .ZN(n7498) );
  XNOR2_X1 U7548 ( .A(n7501), .B(a_29_), .ZN(n7499) );
  AND2_X1 U7549 ( .A1(n7502), .A2(n7503), .ZN(n7497) );
  OR2_X1 U7550 ( .A1(n7504), .A2(n7505), .ZN(n7502) );
  AND2_X1 U7551 ( .A1(n7506), .A2(operation), .ZN(n7494) );
  XOR2_X1 U7552 ( .A(n7507), .B(n7508), .Z(n7506) );
  XNOR2_X1 U7553 ( .A(n7509), .B(n7510), .ZN(n7508) );
  OR2_X1 U7554 ( .A1(n7511), .A2(n7512), .ZN(Result_60_) );
  AND2_X1 U7555 ( .A1(n7513), .A2(operation), .ZN(n7512) );
  XNOR2_X1 U7556 ( .A(n7514), .B(n7515), .ZN(n7513) );
  XOR2_X1 U7557 ( .A(n7516), .B(n7517), .Z(n7515) );
  AND2_X1 U7558 ( .A1(n7518), .A2(n7478), .ZN(n7511) );
  XNOR2_X1 U7559 ( .A(n7519), .B(n7520), .ZN(n7518) );
  AND2_X1 U7560 ( .A1(n7521), .A2(n7522), .ZN(n7520) );
  OR2_X1 U7561 ( .A1(b_28_), .A2(a_28_), .ZN(n7522) );
  AND2_X1 U7562 ( .A1(operation), .A2(n7523), .ZN(Result_5_) );
  XOR2_X1 U7563 ( .A(n7524), .B(n7525), .Z(n7523) );
  AND2_X1 U7564 ( .A1(n7526), .A2(n7527), .ZN(n7525) );
  OR2_X1 U7565 ( .A1(n7528), .A2(n7529), .ZN(n7527) );
  AND2_X1 U7566 ( .A1(n7530), .A2(n7531), .ZN(n7529) );
  INV_X1 U7567 ( .A(n7532), .ZN(n7526) );
  OR2_X1 U7568 ( .A1(n7533), .A2(n7534), .ZN(Result_59_) );
  AND2_X1 U7569 ( .A1(n7535), .A2(n7478), .ZN(n7534) );
  OR2_X1 U7570 ( .A1(n7536), .A2(n7537), .ZN(n7535) );
  AND2_X1 U7571 ( .A1(n7538), .A2(n7539), .ZN(n7537) );
  XNOR2_X1 U7572 ( .A(n7540), .B(a_27_), .ZN(n7538) );
  AND2_X1 U7573 ( .A1(n7541), .A2(n7542), .ZN(n7536) );
  OR2_X1 U7574 ( .A1(n7543), .A2(n7544), .ZN(n7542) );
  INV_X1 U7575 ( .A(n7539), .ZN(n7541) );
  AND2_X1 U7576 ( .A1(n7545), .A2(operation), .ZN(n7533) );
  XNOR2_X1 U7577 ( .A(n7546), .B(n7547), .ZN(n7545) );
  XOR2_X1 U7578 ( .A(n7548), .B(n7549), .Z(n7547) );
  OR2_X1 U7579 ( .A1(n7550), .A2(n7551), .ZN(Result_58_) );
  AND2_X1 U7580 ( .A1(n7552), .A2(operation), .ZN(n7551) );
  XNOR2_X1 U7581 ( .A(n7553), .B(n7554), .ZN(n7552) );
  XOR2_X1 U7582 ( .A(n7555), .B(n7556), .Z(n7554) );
  AND2_X1 U7583 ( .A1(n7557), .A2(n7478), .ZN(n7550) );
  XNOR2_X1 U7584 ( .A(n7558), .B(n7559), .ZN(n7557) );
  AND2_X1 U7585 ( .A1(n7560), .A2(n7561), .ZN(n7559) );
  OR2_X1 U7586 ( .A1(b_26_), .A2(a_26_), .ZN(n7561) );
  OR2_X1 U7587 ( .A1(n7562), .A2(n7563), .ZN(Result_57_) );
  AND2_X1 U7588 ( .A1(n7564), .A2(n7478), .ZN(n7563) );
  OR2_X1 U7589 ( .A1(n7565), .A2(n7566), .ZN(n7564) );
  AND2_X1 U7590 ( .A1(n7567), .A2(n7568), .ZN(n7566) );
  XNOR2_X1 U7591 ( .A(n7569), .B(a_25_), .ZN(n7567) );
  AND2_X1 U7592 ( .A1(n7570), .A2(n7571), .ZN(n7565) );
  OR2_X1 U7593 ( .A1(n7572), .A2(n7573), .ZN(n7571) );
  INV_X1 U7594 ( .A(n7568), .ZN(n7570) );
  AND2_X1 U7595 ( .A1(n7574), .A2(operation), .ZN(n7562) );
  XNOR2_X1 U7596 ( .A(n7575), .B(n7576), .ZN(n7574) );
  XOR2_X1 U7597 ( .A(n7577), .B(n7578), .Z(n7576) );
  OR2_X1 U7598 ( .A1(n7579), .A2(n7580), .ZN(Result_56_) );
  AND2_X1 U7599 ( .A1(n7581), .A2(operation), .ZN(n7580) );
  XNOR2_X1 U7600 ( .A(n7582), .B(n7583), .ZN(n7581) );
  XOR2_X1 U7601 ( .A(n7584), .B(n7585), .Z(n7583) );
  AND2_X1 U7602 ( .A1(n7586), .A2(n7478), .ZN(n7579) );
  XNOR2_X1 U7603 ( .A(n7587), .B(n7588), .ZN(n7586) );
  AND2_X1 U7604 ( .A1(n7589), .A2(n7590), .ZN(n7588) );
  OR2_X1 U7605 ( .A1(b_24_), .A2(a_24_), .ZN(n7590) );
  OR2_X1 U7606 ( .A1(n7591), .A2(n7592), .ZN(Result_55_) );
  AND2_X1 U7607 ( .A1(n7593), .A2(n7478), .ZN(n7592) );
  OR2_X1 U7608 ( .A1(n7594), .A2(n7595), .ZN(n7593) );
  AND2_X1 U7609 ( .A1(n7596), .A2(n7597), .ZN(n7595) );
  XNOR2_X1 U7610 ( .A(n7598), .B(a_23_), .ZN(n7596) );
  AND2_X1 U7611 ( .A1(n7599), .A2(n7600), .ZN(n7594) );
  OR2_X1 U7612 ( .A1(n7601), .A2(n7602), .ZN(n7600) );
  INV_X1 U7613 ( .A(n7597), .ZN(n7599) );
  AND2_X1 U7614 ( .A1(n7603), .A2(operation), .ZN(n7591) );
  XNOR2_X1 U7615 ( .A(n7604), .B(n7605), .ZN(n7603) );
  XOR2_X1 U7616 ( .A(n7606), .B(n7607), .Z(n7605) );
  OR2_X1 U7617 ( .A1(n7608), .A2(n7609), .ZN(Result_54_) );
  AND2_X1 U7618 ( .A1(n7610), .A2(operation), .ZN(n7609) );
  XNOR2_X1 U7619 ( .A(n7611), .B(n7612), .ZN(n7610) );
  XOR2_X1 U7620 ( .A(n7613), .B(n7614), .Z(n7612) );
  AND2_X1 U7621 ( .A1(n7615), .A2(n7478), .ZN(n7608) );
  XOR2_X1 U7622 ( .A(n7616), .B(n7617), .Z(n7615) );
  OR2_X1 U7623 ( .A1(n7618), .A2(n7619), .ZN(n7617) );
  OR2_X1 U7624 ( .A1(n7620), .A2(n7621), .ZN(Result_53_) );
  AND2_X1 U7625 ( .A1(n7622), .A2(n7478), .ZN(n7621) );
  OR2_X1 U7626 ( .A1(n7623), .A2(n7624), .ZN(n7622) );
  AND2_X1 U7627 ( .A1(n7625), .A2(n7626), .ZN(n7624) );
  XNOR2_X1 U7628 ( .A(n7627), .B(a_21_), .ZN(n7625) );
  AND2_X1 U7629 ( .A1(n7628), .A2(n7629), .ZN(n7623) );
  OR2_X1 U7630 ( .A1(n7630), .A2(n7631), .ZN(n7629) );
  INV_X1 U7631 ( .A(n7626), .ZN(n7628) );
  AND2_X1 U7632 ( .A1(n7632), .A2(operation), .ZN(n7620) );
  XNOR2_X1 U7633 ( .A(n7633), .B(n7634), .ZN(n7632) );
  XOR2_X1 U7634 ( .A(n7635), .B(n7636), .Z(n7634) );
  OR2_X1 U7635 ( .A1(n7637), .A2(n7638), .ZN(Result_52_) );
  AND2_X1 U7636 ( .A1(n7639), .A2(operation), .ZN(n7638) );
  XNOR2_X1 U7637 ( .A(n7640), .B(n7641), .ZN(n7639) );
  XOR2_X1 U7638 ( .A(n7642), .B(n7643), .Z(n7641) );
  AND2_X1 U7639 ( .A1(n7644), .A2(n7478), .ZN(n7637) );
  XOR2_X1 U7640 ( .A(n7645), .B(n7646), .Z(n7644) );
  OR2_X1 U7641 ( .A1(n7647), .A2(n7648), .ZN(n7646) );
  OR2_X1 U7642 ( .A1(n7649), .A2(n7650), .ZN(Result_51_) );
  AND2_X1 U7643 ( .A1(n7651), .A2(n7478), .ZN(n7650) );
  OR2_X1 U7644 ( .A1(n7652), .A2(n7653), .ZN(n7651) );
  AND2_X1 U7645 ( .A1(n7654), .A2(n7655), .ZN(n7653) );
  XNOR2_X1 U7646 ( .A(n7656), .B(a_19_), .ZN(n7654) );
  AND2_X1 U7647 ( .A1(n7657), .A2(n7658), .ZN(n7652) );
  OR2_X1 U7648 ( .A1(n7659), .A2(n7660), .ZN(n7658) );
  INV_X1 U7649 ( .A(n7655), .ZN(n7657) );
  AND2_X1 U7650 ( .A1(n7661), .A2(operation), .ZN(n7649) );
  XNOR2_X1 U7651 ( .A(n7662), .B(n7663), .ZN(n7661) );
  XOR2_X1 U7652 ( .A(n7664), .B(n7665), .Z(n7663) );
  OR2_X1 U7653 ( .A1(n7666), .A2(n7667), .ZN(Result_50_) );
  AND2_X1 U7654 ( .A1(n7668), .A2(operation), .ZN(n7667) );
  XNOR2_X1 U7655 ( .A(n7669), .B(n7670), .ZN(n7668) );
  XOR2_X1 U7656 ( .A(n7671), .B(n7672), .Z(n7670) );
  AND2_X1 U7657 ( .A1(n7673), .A2(n7478), .ZN(n7666) );
  XOR2_X1 U7658 ( .A(n7674), .B(n7675), .Z(n7673) );
  OR2_X1 U7659 ( .A1(n7676), .A2(n7677), .ZN(n7675) );
  AND2_X1 U7660 ( .A1(n7678), .A2(operation), .ZN(Result_4_) );
  XOR2_X1 U7661 ( .A(n7679), .B(n7680), .Z(n7678) );
  OR2_X1 U7662 ( .A1(n7681), .A2(n7682), .ZN(Result_49_) );
  AND2_X1 U7663 ( .A1(n7683), .A2(n7478), .ZN(n7682) );
  OR2_X1 U7664 ( .A1(n7684), .A2(n7685), .ZN(n7683) );
  AND2_X1 U7665 ( .A1(n7686), .A2(n7687), .ZN(n7685) );
  XNOR2_X1 U7666 ( .A(n7688), .B(a_17_), .ZN(n7686) );
  AND2_X1 U7667 ( .A1(n7689), .A2(n7690), .ZN(n7684) );
  OR2_X1 U7668 ( .A1(n7691), .A2(n7692), .ZN(n7690) );
  INV_X1 U7669 ( .A(n7687), .ZN(n7689) );
  AND2_X1 U7670 ( .A1(n7693), .A2(operation), .ZN(n7681) );
  XNOR2_X1 U7671 ( .A(n7694), .B(n7695), .ZN(n7693) );
  XOR2_X1 U7672 ( .A(n7696), .B(n7697), .Z(n7695) );
  OR2_X1 U7673 ( .A1(n7698), .A2(n7699), .ZN(Result_48_) );
  AND2_X1 U7674 ( .A1(n7700), .A2(operation), .ZN(n7699) );
  XNOR2_X1 U7675 ( .A(n7701), .B(n7702), .ZN(n7700) );
  XOR2_X1 U7676 ( .A(n7703), .B(n7704), .Z(n7702) );
  AND2_X1 U7677 ( .A1(n7705), .A2(n7478), .ZN(n7698) );
  XOR2_X1 U7678 ( .A(n7706), .B(n7707), .Z(n7705) );
  OR2_X1 U7679 ( .A1(n7708), .A2(n7709), .ZN(n7707) );
  OR2_X1 U7680 ( .A1(n7710), .A2(n7711), .ZN(Result_47_) );
  AND2_X1 U7681 ( .A1(n7712), .A2(n7478), .ZN(n7711) );
  OR2_X1 U7682 ( .A1(n7713), .A2(n7714), .ZN(n7712) );
  AND2_X1 U7683 ( .A1(n7715), .A2(n7716), .ZN(n7714) );
  XNOR2_X1 U7684 ( .A(n7717), .B(a_15_), .ZN(n7715) );
  AND2_X1 U7685 ( .A1(n7718), .A2(n7719), .ZN(n7713) );
  OR2_X1 U7686 ( .A1(n7720), .A2(n7721), .ZN(n7719) );
  INV_X1 U7687 ( .A(n7716), .ZN(n7718) );
  AND2_X1 U7688 ( .A1(n7722), .A2(operation), .ZN(n7710) );
  XNOR2_X1 U7689 ( .A(n7723), .B(n7724), .ZN(n7722) );
  XOR2_X1 U7690 ( .A(n7725), .B(n7726), .Z(n7724) );
  OR2_X1 U7691 ( .A1(n7727), .A2(n7728), .ZN(Result_46_) );
  AND2_X1 U7692 ( .A1(n7729), .A2(operation), .ZN(n7728) );
  XNOR2_X1 U7693 ( .A(n7730), .B(n7731), .ZN(n7729) );
  XOR2_X1 U7694 ( .A(n7732), .B(n7733), .Z(n7731) );
  AND2_X1 U7695 ( .A1(n7734), .A2(n7478), .ZN(n7727) );
  XOR2_X1 U7696 ( .A(n7735), .B(n7736), .Z(n7734) );
  OR2_X1 U7697 ( .A1(n7737), .A2(n7738), .ZN(n7736) );
  OR2_X1 U7698 ( .A1(n7739), .A2(n7740), .ZN(Result_45_) );
  AND2_X1 U7699 ( .A1(n7741), .A2(n7478), .ZN(n7740) );
  OR2_X1 U7700 ( .A1(n7742), .A2(n7743), .ZN(n7741) );
  AND2_X1 U7701 ( .A1(n7744), .A2(n7745), .ZN(n7743) );
  XNOR2_X1 U7702 ( .A(n7746), .B(a_13_), .ZN(n7744) );
  AND2_X1 U7703 ( .A1(n7747), .A2(n7748), .ZN(n7742) );
  OR2_X1 U7704 ( .A1(n7749), .A2(n7750), .ZN(n7748) );
  INV_X1 U7705 ( .A(n7745), .ZN(n7747) );
  AND2_X1 U7706 ( .A1(n7751), .A2(operation), .ZN(n7739) );
  XNOR2_X1 U7707 ( .A(n7752), .B(n7753), .ZN(n7751) );
  XOR2_X1 U7708 ( .A(n7754), .B(n7755), .Z(n7753) );
  OR2_X1 U7709 ( .A1(n7756), .A2(n7757), .ZN(Result_44_) );
  AND2_X1 U7710 ( .A1(n7758), .A2(operation), .ZN(n7757) );
  XNOR2_X1 U7711 ( .A(n7759), .B(n7760), .ZN(n7758) );
  XOR2_X1 U7712 ( .A(n7761), .B(n7762), .Z(n7760) );
  AND2_X1 U7713 ( .A1(n7763), .A2(n7478), .ZN(n7756) );
  XOR2_X1 U7714 ( .A(n7764), .B(n7765), .Z(n7763) );
  OR2_X1 U7715 ( .A1(n7766), .A2(n7767), .ZN(n7765) );
  OR2_X1 U7716 ( .A1(n7768), .A2(n7769), .ZN(Result_43_) );
  AND2_X1 U7717 ( .A1(n7770), .A2(n7478), .ZN(n7769) );
  OR2_X1 U7718 ( .A1(n7771), .A2(n7772), .ZN(n7770) );
  AND2_X1 U7719 ( .A1(n7773), .A2(n7774), .ZN(n7772) );
  XNOR2_X1 U7720 ( .A(n7775), .B(a_11_), .ZN(n7773) );
  AND2_X1 U7721 ( .A1(n7776), .A2(n7777), .ZN(n7771) );
  OR2_X1 U7722 ( .A1(n7778), .A2(n7779), .ZN(n7777) );
  INV_X1 U7723 ( .A(n7774), .ZN(n7776) );
  AND2_X1 U7724 ( .A1(n7780), .A2(operation), .ZN(n7768) );
  XNOR2_X1 U7725 ( .A(n7781), .B(n7782), .ZN(n7780) );
  XOR2_X1 U7726 ( .A(n7783), .B(n7784), .Z(n7782) );
  OR2_X1 U7727 ( .A1(n7785), .A2(n7786), .ZN(Result_42_) );
  AND2_X1 U7728 ( .A1(n7787), .A2(operation), .ZN(n7786) );
  XNOR2_X1 U7729 ( .A(n7788), .B(n7789), .ZN(n7787) );
  XOR2_X1 U7730 ( .A(n7790), .B(n7791), .Z(n7789) );
  AND2_X1 U7731 ( .A1(n7792), .A2(n7478), .ZN(n7785) );
  XOR2_X1 U7732 ( .A(n7793), .B(n7794), .Z(n7792) );
  OR2_X1 U7733 ( .A1(n7795), .A2(n7796), .ZN(n7794) );
  OR2_X1 U7734 ( .A1(n7797), .A2(n7798), .ZN(Result_41_) );
  AND2_X1 U7735 ( .A1(n7799), .A2(n7478), .ZN(n7798) );
  OR2_X1 U7736 ( .A1(n7800), .A2(n7801), .ZN(n7799) );
  AND2_X1 U7737 ( .A1(n7802), .A2(n7803), .ZN(n7801) );
  XNOR2_X1 U7738 ( .A(n7804), .B(a_9_), .ZN(n7802) );
  AND2_X1 U7739 ( .A1(n7805), .A2(n7806), .ZN(n7800) );
  OR2_X1 U7740 ( .A1(n7807), .A2(n7808), .ZN(n7806) );
  INV_X1 U7741 ( .A(n7803), .ZN(n7805) );
  AND2_X1 U7742 ( .A1(n7809), .A2(operation), .ZN(n7797) );
  XNOR2_X1 U7743 ( .A(n7810), .B(n7811), .ZN(n7809) );
  XOR2_X1 U7744 ( .A(n7812), .B(n7813), .Z(n7811) );
  OR2_X1 U7745 ( .A1(n7814), .A2(n7815), .ZN(Result_40_) );
  AND2_X1 U7746 ( .A1(n7816), .A2(operation), .ZN(n7815) );
  XNOR2_X1 U7747 ( .A(n7817), .B(n7818), .ZN(n7816) );
  XOR2_X1 U7748 ( .A(n7819), .B(n7820), .Z(n7818) );
  AND2_X1 U7749 ( .A1(n7821), .A2(n7478), .ZN(n7814) );
  XOR2_X1 U7750 ( .A(n7822), .B(n7823), .Z(n7821) );
  OR2_X1 U7751 ( .A1(n7824), .A2(n7825), .ZN(n7823) );
  AND2_X1 U7752 ( .A1(operation), .A2(n7826), .ZN(Result_3_) );
  XOR2_X1 U7753 ( .A(n7827), .B(n7828), .Z(n7826) );
  AND2_X1 U7754 ( .A1(n7829), .A2(n7830), .ZN(n7828) );
  OR2_X1 U7755 ( .A1(n7831), .A2(n7832), .ZN(n7830) );
  AND2_X1 U7756 ( .A1(n7833), .A2(n7834), .ZN(n7832) );
  INV_X1 U7757 ( .A(n7835), .ZN(n7829) );
  OR2_X1 U7758 ( .A1(n7836), .A2(n7837), .ZN(Result_39_) );
  AND2_X1 U7759 ( .A1(n7838), .A2(n7478), .ZN(n7837) );
  OR2_X1 U7760 ( .A1(n7839), .A2(n7840), .ZN(n7838) );
  AND2_X1 U7761 ( .A1(n7841), .A2(n7842), .ZN(n7840) );
  XNOR2_X1 U7762 ( .A(n7843), .B(a_7_), .ZN(n7841) );
  AND2_X1 U7763 ( .A1(n7844), .A2(n7845), .ZN(n7839) );
  OR2_X1 U7764 ( .A1(n7846), .A2(n7847), .ZN(n7845) );
  INV_X1 U7765 ( .A(n7842), .ZN(n7844) );
  AND2_X1 U7766 ( .A1(n7848), .A2(operation), .ZN(n7836) );
  XNOR2_X1 U7767 ( .A(n7849), .B(n7850), .ZN(n7848) );
  XOR2_X1 U7768 ( .A(n7851), .B(n7852), .Z(n7850) );
  OR2_X1 U7769 ( .A1(n7853), .A2(n7854), .ZN(Result_38_) );
  AND2_X1 U7770 ( .A1(n7855), .A2(operation), .ZN(n7854) );
  XNOR2_X1 U7771 ( .A(n7856), .B(n7857), .ZN(n7855) );
  XOR2_X1 U7772 ( .A(n7858), .B(n7859), .Z(n7857) );
  AND2_X1 U7773 ( .A1(n7860), .A2(n7478), .ZN(n7853) );
  XOR2_X1 U7774 ( .A(n7861), .B(n7862), .Z(n7860) );
  OR2_X1 U7775 ( .A1(n7863), .A2(n7864), .ZN(n7862) );
  OR2_X1 U7776 ( .A1(n7865), .A2(n7866), .ZN(Result_37_) );
  AND2_X1 U7777 ( .A1(n7867), .A2(n7478), .ZN(n7866) );
  OR2_X1 U7778 ( .A1(n7868), .A2(n7869), .ZN(n7867) );
  AND2_X1 U7779 ( .A1(n7870), .A2(n7871), .ZN(n7869) );
  XNOR2_X1 U7780 ( .A(n7872), .B(a_5_), .ZN(n7870) );
  AND2_X1 U7781 ( .A1(n7873), .A2(n7874), .ZN(n7868) );
  OR2_X1 U7782 ( .A1(n7875), .A2(n7876), .ZN(n7874) );
  INV_X1 U7783 ( .A(n7871), .ZN(n7873) );
  AND2_X1 U7784 ( .A1(n7877), .A2(operation), .ZN(n7865) );
  XNOR2_X1 U7785 ( .A(n7878), .B(n7879), .ZN(n7877) );
  XOR2_X1 U7786 ( .A(n7880), .B(n7881), .Z(n7879) );
  OR2_X1 U7787 ( .A1(n7882), .A2(n7883), .ZN(Result_36_) );
  AND2_X1 U7788 ( .A1(n7884), .A2(operation), .ZN(n7883) );
  XNOR2_X1 U7789 ( .A(n7885), .B(n7886), .ZN(n7884) );
  XOR2_X1 U7790 ( .A(n7887), .B(n7888), .Z(n7886) );
  AND2_X1 U7791 ( .A1(n7889), .A2(n7478), .ZN(n7882) );
  XOR2_X1 U7792 ( .A(n7890), .B(n7891), .Z(n7889) );
  OR2_X1 U7793 ( .A1(n7892), .A2(n7893), .ZN(n7891) );
  OR2_X1 U7794 ( .A1(n7894), .A2(n7895), .ZN(Result_35_) );
  AND2_X1 U7795 ( .A1(n7896), .A2(n7478), .ZN(n7895) );
  OR2_X1 U7796 ( .A1(n7897), .A2(n7898), .ZN(n7896) );
  AND2_X1 U7797 ( .A1(n7899), .A2(n7900), .ZN(n7898) );
  XNOR2_X1 U7798 ( .A(n7901), .B(a_3_), .ZN(n7899) );
  AND2_X1 U7799 ( .A1(n7902), .A2(n7903), .ZN(n7897) );
  OR2_X1 U7800 ( .A1(n7904), .A2(n7905), .ZN(n7903) );
  INV_X1 U7801 ( .A(n7900), .ZN(n7902) );
  AND2_X1 U7802 ( .A1(n7906), .A2(operation), .ZN(n7894) );
  XNOR2_X1 U7803 ( .A(n7907), .B(n7908), .ZN(n7906) );
  XOR2_X1 U7804 ( .A(n7909), .B(n7910), .Z(n7908) );
  OR2_X1 U7805 ( .A1(n7911), .A2(n7912), .ZN(Result_34_) );
  AND2_X1 U7806 ( .A1(n7913), .A2(operation), .ZN(n7912) );
  XNOR2_X1 U7807 ( .A(n7914), .B(n7915), .ZN(n7913) );
  XOR2_X1 U7808 ( .A(n7916), .B(n7917), .Z(n7915) );
  AND2_X1 U7809 ( .A1(n7918), .A2(n7478), .ZN(n7911) );
  XOR2_X1 U7810 ( .A(n7919), .B(n7920), .Z(n7918) );
  OR2_X1 U7811 ( .A1(n7921), .A2(n7922), .ZN(n7920) );
  OR2_X1 U7812 ( .A1(n7923), .A2(n7924), .ZN(Result_33_) );
  AND2_X1 U7813 ( .A1(n7925), .A2(n7478), .ZN(n7924) );
  OR2_X1 U7814 ( .A1(n7926), .A2(n7927), .ZN(n7925) );
  AND2_X1 U7815 ( .A1(n7928), .A2(n7929), .ZN(n7927) );
  XNOR2_X1 U7816 ( .A(n7930), .B(a_1_), .ZN(n7928) );
  AND2_X1 U7817 ( .A1(n7931), .A2(n7932), .ZN(n7926) );
  OR2_X1 U7818 ( .A1(n7933), .A2(n7934), .ZN(n7932) );
  INV_X1 U7819 ( .A(n7929), .ZN(n7931) );
  AND2_X1 U7820 ( .A1(n7935), .A2(operation), .ZN(n7923) );
  XNOR2_X1 U7821 ( .A(n7936), .B(n7937), .ZN(n7935) );
  XOR2_X1 U7822 ( .A(n7938), .B(n7939), .Z(n7937) );
  OR2_X1 U7823 ( .A1(n7940), .A2(n7941), .ZN(Result_32_) );
  AND2_X1 U7824 ( .A1(n7942), .A2(operation), .ZN(n7941) );
  XNOR2_X1 U7825 ( .A(n7943), .B(n7944), .ZN(n7942) );
  XOR2_X1 U7826 ( .A(n7945), .B(n7946), .Z(n7944) );
  AND2_X1 U7827 ( .A1(n7947), .A2(n7478), .ZN(n7940) );
  INV_X1 U7828 ( .A(operation), .ZN(n7478) );
  XOR2_X1 U7829 ( .A(n7948), .B(n7949), .Z(n7947) );
  XNOR2_X1 U7830 ( .A(n7950), .B(n7951), .ZN(n7949) );
  OR2_X1 U7831 ( .A1(n7952), .A2(n7933), .ZN(n7948) );
  AND2_X1 U7832 ( .A1(n7953), .A2(n7930), .ZN(n7933) );
  AND2_X1 U7833 ( .A1(n7929), .A2(n7954), .ZN(n7952) );
  OR2_X1 U7834 ( .A1(n7955), .A2(n7921), .ZN(n7929) );
  AND2_X1 U7835 ( .A1(n7956), .A2(n7957), .ZN(n7921) );
  AND2_X1 U7836 ( .A1(n7919), .A2(n7958), .ZN(n7955) );
  OR2_X1 U7837 ( .A1(n7959), .A2(n7904), .ZN(n7919) );
  AND2_X1 U7838 ( .A1(n7960), .A2(n7901), .ZN(n7904) );
  AND2_X1 U7839 ( .A1(n7900), .A2(n7961), .ZN(n7959) );
  OR2_X1 U7840 ( .A1(n7962), .A2(n7892), .ZN(n7900) );
  AND2_X1 U7841 ( .A1(n7963), .A2(n7964), .ZN(n7892) );
  AND2_X1 U7842 ( .A1(n7890), .A2(n7965), .ZN(n7962) );
  OR2_X1 U7843 ( .A1(n7966), .A2(n7875), .ZN(n7890) );
  AND2_X1 U7844 ( .A1(n7967), .A2(n7872), .ZN(n7875) );
  AND2_X1 U7845 ( .A1(n7871), .A2(n7968), .ZN(n7966) );
  OR2_X1 U7846 ( .A1(n7969), .A2(n7863), .ZN(n7871) );
  AND2_X1 U7847 ( .A1(n7970), .A2(n7971), .ZN(n7863) );
  AND2_X1 U7848 ( .A1(n7861), .A2(n7972), .ZN(n7969) );
  OR2_X1 U7849 ( .A1(n7973), .A2(n7846), .ZN(n7861) );
  AND2_X1 U7850 ( .A1(n7974), .A2(n7843), .ZN(n7846) );
  AND2_X1 U7851 ( .A1(n7842), .A2(n7975), .ZN(n7973) );
  OR2_X1 U7852 ( .A1(n7976), .A2(n7824), .ZN(n7842) );
  AND2_X1 U7853 ( .A1(n7977), .A2(n7978), .ZN(n7824) );
  AND2_X1 U7854 ( .A1(n7822), .A2(n7979), .ZN(n7976) );
  OR2_X1 U7855 ( .A1(n7980), .A2(n7807), .ZN(n7822) );
  AND2_X1 U7856 ( .A1(n7981), .A2(n7804), .ZN(n7807) );
  AND2_X1 U7857 ( .A1(n7803), .A2(n7982), .ZN(n7980) );
  OR2_X1 U7858 ( .A1(n7983), .A2(n7795), .ZN(n7803) );
  AND2_X1 U7859 ( .A1(n7984), .A2(n7985), .ZN(n7795) );
  AND2_X1 U7860 ( .A1(n7793), .A2(n7986), .ZN(n7983) );
  OR2_X1 U7861 ( .A1(n7987), .A2(n7778), .ZN(n7793) );
  AND2_X1 U7862 ( .A1(n7988), .A2(n7775), .ZN(n7778) );
  AND2_X1 U7863 ( .A1(n7774), .A2(n7989), .ZN(n7987) );
  OR2_X1 U7864 ( .A1(n7990), .A2(n7766), .ZN(n7774) );
  AND2_X1 U7865 ( .A1(n7991), .A2(n7992), .ZN(n7766) );
  AND2_X1 U7866 ( .A1(n7764), .A2(n7993), .ZN(n7990) );
  OR2_X1 U7867 ( .A1(n7994), .A2(n7749), .ZN(n7764) );
  AND2_X1 U7868 ( .A1(n7995), .A2(n7746), .ZN(n7749) );
  AND2_X1 U7869 ( .A1(n7745), .A2(n7996), .ZN(n7994) );
  OR2_X1 U7870 ( .A1(n7997), .A2(n7737), .ZN(n7745) );
  AND2_X1 U7871 ( .A1(n7998), .A2(n7999), .ZN(n7737) );
  AND2_X1 U7872 ( .A1(n7735), .A2(n8000), .ZN(n7997) );
  OR2_X1 U7873 ( .A1(n8001), .A2(n7720), .ZN(n7735) );
  AND2_X1 U7874 ( .A1(n8002), .A2(n7717), .ZN(n7720) );
  AND2_X1 U7875 ( .A1(n7716), .A2(n8003), .ZN(n8001) );
  OR2_X1 U7876 ( .A1(n8004), .A2(n7708), .ZN(n7716) );
  AND2_X1 U7877 ( .A1(n8005), .A2(n8006), .ZN(n7708) );
  AND2_X1 U7878 ( .A1(n7706), .A2(n8007), .ZN(n8004) );
  OR2_X1 U7879 ( .A1(n8008), .A2(n7691), .ZN(n7706) );
  AND2_X1 U7880 ( .A1(n8009), .A2(n7688), .ZN(n7691) );
  AND2_X1 U7881 ( .A1(n7687), .A2(n8010), .ZN(n8008) );
  OR2_X1 U7882 ( .A1(n8011), .A2(n7676), .ZN(n7687) );
  AND2_X1 U7883 ( .A1(n8012), .A2(n8013), .ZN(n7676) );
  AND2_X1 U7884 ( .A1(n7674), .A2(n8014), .ZN(n8011) );
  OR2_X1 U7885 ( .A1(n8015), .A2(n7659), .ZN(n7674) );
  AND2_X1 U7886 ( .A1(n8016), .A2(n7656), .ZN(n7659) );
  AND2_X1 U7887 ( .A1(n7655), .A2(n8017), .ZN(n8015) );
  OR2_X1 U7888 ( .A1(n8018), .A2(n7647), .ZN(n7655) );
  AND2_X1 U7889 ( .A1(n8019), .A2(n8020), .ZN(n7647) );
  AND2_X1 U7890 ( .A1(n7645), .A2(n8021), .ZN(n8018) );
  OR2_X1 U7891 ( .A1(n8022), .A2(n7630), .ZN(n7645) );
  AND2_X1 U7892 ( .A1(n8023), .A2(n7627), .ZN(n7630) );
  AND2_X1 U7893 ( .A1(n7626), .A2(n8024), .ZN(n8022) );
  OR2_X1 U7894 ( .A1(n8025), .A2(n7618), .ZN(n7626) );
  AND2_X1 U7895 ( .A1(n8026), .A2(n8027), .ZN(n7618) );
  AND2_X1 U7896 ( .A1(n7616), .A2(n8028), .ZN(n8025) );
  OR2_X1 U7897 ( .A1(n8029), .A2(n7601), .ZN(n7616) );
  AND2_X1 U7898 ( .A1(n8030), .A2(n7598), .ZN(n7601) );
  AND2_X1 U7899 ( .A1(n7597), .A2(n8031), .ZN(n8029) );
  OR2_X1 U7900 ( .A1(n8032), .A2(n8033), .ZN(n7597) );
  AND2_X1 U7901 ( .A1(n8034), .A2(n8035), .ZN(n8033) );
  AND2_X1 U7902 ( .A1(n7587), .A2(n7589), .ZN(n8032) );
  OR2_X1 U7903 ( .A1(n8036), .A2(n7572), .ZN(n7587) );
  AND2_X1 U7904 ( .A1(n8037), .A2(n7569), .ZN(n7572) );
  AND2_X1 U7905 ( .A1(n7568), .A2(n8038), .ZN(n8036) );
  OR2_X1 U7906 ( .A1(n8039), .A2(n8040), .ZN(n7568) );
  AND2_X1 U7907 ( .A1(n8041), .A2(n8042), .ZN(n8040) );
  AND2_X1 U7908 ( .A1(n7558), .A2(n7560), .ZN(n8039) );
  OR2_X1 U7909 ( .A1(n8043), .A2(n7543), .ZN(n7558) );
  AND2_X1 U7910 ( .A1(n8044), .A2(n7540), .ZN(n7543) );
  AND2_X1 U7911 ( .A1(n7539), .A2(n8045), .ZN(n8043) );
  OR2_X1 U7912 ( .A1(n8046), .A2(n8047), .ZN(n7539) );
  AND2_X1 U7913 ( .A1(n8048), .A2(n8049), .ZN(n8047) );
  AND2_X1 U7914 ( .A1(n7519), .A2(n7521), .ZN(n8046) );
  OR2_X1 U7915 ( .A1(n8050), .A2(n7504), .ZN(n7519) );
  AND2_X1 U7916 ( .A1(n8051), .A2(n7501), .ZN(n7504) );
  AND2_X1 U7917 ( .A1(n7500), .A2(n8052), .ZN(n8050) );
  INV_X1 U7918 ( .A(n7503), .ZN(n7500) );
  OR2_X1 U7919 ( .A1(n8053), .A2(n8054), .ZN(n7503) );
  AND2_X1 U7920 ( .A1(b_30_), .A2(n8055), .ZN(n8054) );
  OR2_X1 U7921 ( .A1(a_30_), .A2(n7476), .ZN(n8055) );
  AND2_X1 U7922 ( .A1(a_31_), .A2(b_31_), .ZN(n7476) );
  AND2_X1 U7923 ( .A1(operation), .A2(n8056), .ZN(Result_31_) );
  XNOR2_X1 U7924 ( .A(n8057), .B(n8058), .ZN(n8056) );
  AND3_X1 U7925 ( .A1(n8059), .A2(n8060), .A3(operation), .ZN(Result_30_) );
  OR2_X1 U7926 ( .A1(n8061), .A2(n8062), .ZN(n8059) );
  AND2_X1 U7927 ( .A1(n8063), .A2(n8058), .ZN(n8061) );
  AND2_X1 U7928 ( .A1(n8064), .A2(operation), .ZN(Result_2_) );
  XOR2_X1 U7929 ( .A(n8065), .B(n8066), .Z(n8064) );
  AND2_X1 U7930 ( .A1(operation), .A2(n8067), .ZN(Result_29_) );
  XNOR2_X1 U7931 ( .A(n8060), .B(n8068), .ZN(n8067) );
  AND2_X1 U7932 ( .A1(n8069), .A2(n8070), .ZN(n8068) );
  INV_X1 U7933 ( .A(n8071), .ZN(n8060) );
  AND2_X1 U7934 ( .A1(n8072), .A2(operation), .ZN(Result_28_) );
  XOR2_X1 U7935 ( .A(n8073), .B(n8074), .Z(n8072) );
  AND2_X1 U7936 ( .A1(n8075), .A2(n8076), .ZN(n8074) );
  INV_X1 U7937 ( .A(n8077), .ZN(n8076) );
  AND2_X1 U7938 ( .A1(n8078), .A2(operation), .ZN(Result_27_) );
  XOR2_X1 U7939 ( .A(n8079), .B(n8080), .Z(n8078) );
  AND2_X1 U7940 ( .A1(n8081), .A2(n8082), .ZN(n8080) );
  INV_X1 U7941 ( .A(n8083), .ZN(n8082) );
  AND2_X1 U7942 ( .A1(n8084), .A2(operation), .ZN(Result_26_) );
  XOR2_X1 U7943 ( .A(n8085), .B(n8086), .Z(n8084) );
  AND2_X1 U7944 ( .A1(n8087), .A2(n8088), .ZN(n8086) );
  INV_X1 U7945 ( .A(n8089), .ZN(n8088) );
  AND2_X1 U7946 ( .A1(n8090), .A2(operation), .ZN(Result_25_) );
  XOR2_X1 U7947 ( .A(n8091), .B(n8092), .Z(n8090) );
  AND2_X1 U7948 ( .A1(n8093), .A2(n8094), .ZN(n8092) );
  INV_X1 U7949 ( .A(n8095), .ZN(n8093) );
  AND2_X1 U7950 ( .A1(n8096), .A2(operation), .ZN(Result_24_) );
  XOR2_X1 U7951 ( .A(n8097), .B(n8098), .Z(n8096) );
  AND2_X1 U7952 ( .A1(n8099), .A2(n8100), .ZN(n8098) );
  AND2_X1 U7953 ( .A1(n8101), .A2(operation), .ZN(Result_23_) );
  XOR2_X1 U7954 ( .A(n8102), .B(n8103), .Z(n8101) );
  AND2_X1 U7955 ( .A1(n8104), .A2(n8105), .ZN(n8103) );
  AND2_X1 U7956 ( .A1(n8106), .A2(operation), .ZN(Result_22_) );
  XOR2_X1 U7957 ( .A(n8107), .B(n8108), .Z(n8106) );
  AND2_X1 U7958 ( .A1(n8109), .A2(n8110), .ZN(n8108) );
  AND2_X1 U7959 ( .A1(n8111), .A2(operation), .ZN(Result_21_) );
  XOR2_X1 U7960 ( .A(n8112), .B(n8113), .Z(n8111) );
  AND2_X1 U7961 ( .A1(n8114), .A2(n8115), .ZN(n8113) );
  INV_X1 U7962 ( .A(n8116), .ZN(n8114) );
  AND2_X1 U7963 ( .A1(n8117), .A2(operation), .ZN(Result_20_) );
  XOR2_X1 U7964 ( .A(n8118), .B(n8119), .Z(n8117) );
  AND2_X1 U7965 ( .A1(n8120), .A2(n8121), .ZN(n8119) );
  AND2_X1 U7966 ( .A1(operation), .A2(n8122), .ZN(Result_1_) );
  XOR2_X1 U7967 ( .A(n8123), .B(n8124), .Z(n8122) );
  AND2_X1 U7968 ( .A1(n8125), .A2(n8126), .ZN(n8124) );
  OR2_X1 U7969 ( .A1(n8127), .A2(n8128), .ZN(n8126) );
  AND2_X1 U7970 ( .A1(n8129), .A2(n8130), .ZN(n8127) );
  INV_X1 U7971 ( .A(n8131), .ZN(n8125) );
  AND2_X1 U7972 ( .A1(n8132), .A2(operation), .ZN(Result_19_) );
  XOR2_X1 U7973 ( .A(n8133), .B(n8134), .Z(n8132) );
  AND2_X1 U7974 ( .A1(n8135), .A2(n8136), .ZN(n8134) );
  AND2_X1 U7975 ( .A1(n8137), .A2(operation), .ZN(Result_18_) );
  XOR2_X1 U7976 ( .A(n8138), .B(n8139), .Z(n8137) );
  AND2_X1 U7977 ( .A1(n8140), .A2(n8141), .ZN(n8139) );
  AND2_X1 U7978 ( .A1(n8142), .A2(operation), .ZN(Result_17_) );
  XOR2_X1 U7979 ( .A(n8143), .B(n8144), .Z(n8142) );
  AND2_X1 U7980 ( .A1(n8145), .A2(n8146), .ZN(n8144) );
  AND2_X1 U7981 ( .A1(n8147), .A2(operation), .ZN(Result_16_) );
  XOR2_X1 U7982 ( .A(n8148), .B(n8149), .Z(n8147) );
  AND2_X1 U7983 ( .A1(n8150), .A2(n8151), .ZN(n8149) );
  AND2_X1 U7984 ( .A1(n8152), .A2(operation), .ZN(Result_15_) );
  XOR2_X1 U7985 ( .A(n8153), .B(n8154), .Z(n8152) );
  AND2_X1 U7986 ( .A1(n8155), .A2(n8156), .ZN(n8154) );
  AND2_X1 U7987 ( .A1(n8157), .A2(operation), .ZN(Result_14_) );
  XOR2_X1 U7988 ( .A(n8158), .B(n8159), .Z(n8157) );
  AND2_X1 U7989 ( .A1(n8160), .A2(n8161), .ZN(n8159) );
  INV_X1 U7990 ( .A(n8162), .ZN(n8161) );
  OR2_X1 U7991 ( .A1(n8163), .A2(n8164), .ZN(n8160) );
  AND2_X1 U7992 ( .A1(n8165), .A2(n8166), .ZN(n8163) );
  AND2_X1 U7993 ( .A1(n8167), .A2(operation), .ZN(Result_13_) );
  XOR2_X1 U7994 ( .A(n8168), .B(n8169), .Z(n8167) );
  AND2_X1 U7995 ( .A1(n8170), .A2(n8171), .ZN(n8169) );
  INV_X1 U7996 ( .A(n8172), .ZN(n8171) );
  OR2_X1 U7997 ( .A1(n8173), .A2(n8174), .ZN(n8170) );
  AND2_X1 U7998 ( .A1(n8175), .A2(n8176), .ZN(n8173) );
  AND2_X1 U7999 ( .A1(n8177), .A2(operation), .ZN(Result_12_) );
  XOR2_X1 U8000 ( .A(n8178), .B(n8179), .Z(n8177) );
  AND2_X1 U8001 ( .A1(operation), .A2(n8180), .ZN(Result_11_) );
  XOR2_X1 U8002 ( .A(n8181), .B(n8182), .Z(n8180) );
  AND2_X1 U8003 ( .A1(n8183), .A2(n8184), .ZN(n8182) );
  INV_X1 U8004 ( .A(n8185), .ZN(n8184) );
  OR2_X1 U8005 ( .A1(n8186), .A2(n8187), .ZN(n8183) );
  AND2_X1 U8006 ( .A1(n8188), .A2(n8189), .ZN(n8186) );
  AND2_X1 U8007 ( .A1(n8190), .A2(operation), .ZN(Result_10_) );
  XOR2_X1 U8008 ( .A(n8191), .B(n8192), .Z(n8190) );
  AND2_X1 U8009 ( .A1(operation), .A2(n8193), .ZN(Result_0_) );
  OR3_X1 U8010 ( .A1(n8131), .A2(n8194), .A3(n8195), .ZN(n8193) );
  AND2_X1 U8011 ( .A1(n8196), .A2(a_0_), .ZN(n8195) );
  AND2_X1 U8012 ( .A1(n8123), .A2(n8128), .ZN(n8194) );
  AND2_X1 U8013 ( .A1(n8065), .A2(n8066), .ZN(n8123) );
  XNOR2_X1 U8014 ( .A(n8130), .B(n8197), .ZN(n8066) );
  OR2_X1 U8015 ( .A1(n8198), .A2(n8199), .ZN(n8065) );
  OR2_X1 U8016 ( .A1(n8200), .A2(n7835), .ZN(n8198) );
  AND3_X1 U8017 ( .A1(n7834), .A2(n7833), .A3(n7831), .ZN(n7835) );
  INV_X1 U8018 ( .A(n8201), .ZN(n7833) );
  AND2_X1 U8019 ( .A1(n7827), .A2(n7831), .ZN(n8200) );
  INV_X1 U8020 ( .A(n8202), .ZN(n7831) );
  OR2_X1 U8021 ( .A1(n8203), .A2(n8199), .ZN(n8202) );
  INV_X1 U8022 ( .A(n8204), .ZN(n8199) );
  OR2_X1 U8023 ( .A1(n8205), .A2(n8206), .ZN(n8204) );
  AND2_X1 U8024 ( .A1(n8205), .A2(n8206), .ZN(n8203) );
  OR2_X1 U8025 ( .A1(n8207), .A2(n8208), .ZN(n8206) );
  AND2_X1 U8026 ( .A1(n8209), .A2(n8210), .ZN(n8208) );
  AND2_X1 U8027 ( .A1(n8211), .A2(n8212), .ZN(n8207) );
  OR2_X1 U8028 ( .A1(n8210), .A2(n8209), .ZN(n8212) );
  XOR2_X1 U8029 ( .A(n8213), .B(n8214), .Z(n8205) );
  XOR2_X1 U8030 ( .A(n8215), .B(n8216), .Z(n8214) );
  AND2_X1 U8031 ( .A1(n7679), .A2(n7680), .ZN(n7827) );
  XNOR2_X1 U8032 ( .A(n7834), .B(n8201), .ZN(n7680) );
  OR2_X1 U8033 ( .A1(n8217), .A2(n8218), .ZN(n8201) );
  AND2_X1 U8034 ( .A1(n8219), .A2(n8220), .ZN(n8218) );
  AND2_X1 U8035 ( .A1(n8221), .A2(n8222), .ZN(n8217) );
  OR2_X1 U8036 ( .A1(n8220), .A2(n8219), .ZN(n8222) );
  XNOR2_X1 U8037 ( .A(n8211), .B(n8223), .ZN(n7834) );
  XOR2_X1 U8038 ( .A(n8210), .B(n8209), .Z(n8223) );
  OR2_X1 U8039 ( .A1(n7901), .A2(n7950), .ZN(n8209) );
  OR2_X1 U8040 ( .A1(n8224), .A2(n8225), .ZN(n8210) );
  AND2_X1 U8041 ( .A1(n8226), .A2(n8227), .ZN(n8225) );
  AND2_X1 U8042 ( .A1(n8228), .A2(n8229), .ZN(n8224) );
  OR2_X1 U8043 ( .A1(n8227), .A2(n8226), .ZN(n8229) );
  XOR2_X1 U8044 ( .A(n8230), .B(n8231), .Z(n8211) );
  XOR2_X1 U8045 ( .A(n8232), .B(n8233), .Z(n8231) );
  OR2_X1 U8046 ( .A1(n8234), .A2(n8235), .ZN(n7679) );
  OR2_X1 U8047 ( .A1(n8236), .A2(n7532), .ZN(n8234) );
  AND3_X1 U8048 ( .A1(n7531), .A2(n7530), .A3(n7528), .ZN(n7532) );
  INV_X1 U8049 ( .A(n8237), .ZN(n7530) );
  AND2_X1 U8050 ( .A1(n7524), .A2(n7528), .ZN(n8236) );
  INV_X1 U8051 ( .A(n8238), .ZN(n7528) );
  OR2_X1 U8052 ( .A1(n8239), .A2(n8235), .ZN(n8238) );
  INV_X1 U8053 ( .A(n8240), .ZN(n8235) );
  OR2_X1 U8054 ( .A1(n8241), .A2(n8242), .ZN(n8240) );
  AND2_X1 U8055 ( .A1(n8241), .A2(n8242), .ZN(n8239) );
  OR2_X1 U8056 ( .A1(n8243), .A2(n8244), .ZN(n8242) );
  AND2_X1 U8057 ( .A1(n8245), .A2(n8246), .ZN(n8244) );
  AND2_X1 U8058 ( .A1(n8247), .A2(n8248), .ZN(n8243) );
  OR2_X1 U8059 ( .A1(n8246), .A2(n8245), .ZN(n8248) );
  XOR2_X1 U8060 ( .A(n8221), .B(n8249), .Z(n8241) );
  XOR2_X1 U8061 ( .A(n8220), .B(n8219), .Z(n8249) );
  OR2_X1 U8062 ( .A1(n7964), .A2(n7950), .ZN(n8219) );
  OR2_X1 U8063 ( .A1(n8250), .A2(n8251), .ZN(n8220) );
  AND2_X1 U8064 ( .A1(n8252), .A2(n8253), .ZN(n8251) );
  AND2_X1 U8065 ( .A1(n8254), .A2(n8255), .ZN(n8250) );
  OR2_X1 U8066 ( .A1(n8253), .A2(n8252), .ZN(n8255) );
  XOR2_X1 U8067 ( .A(n8228), .B(n8256), .Z(n8221) );
  XOR2_X1 U8068 ( .A(n8227), .B(n8226), .Z(n8256) );
  OR2_X1 U8069 ( .A1(n7901), .A2(n7953), .ZN(n8226) );
  OR2_X1 U8070 ( .A1(n8257), .A2(n8258), .ZN(n8227) );
  AND2_X1 U8071 ( .A1(n8259), .A2(n8260), .ZN(n8258) );
  AND2_X1 U8072 ( .A1(n8261), .A2(n8262), .ZN(n8257) );
  OR2_X1 U8073 ( .A1(n8260), .A2(n8259), .ZN(n8262) );
  XNOR2_X1 U8074 ( .A(n8263), .B(n8264), .ZN(n8228) );
  XNOR2_X1 U8075 ( .A(n7958), .B(n8265), .ZN(n8263) );
  AND2_X1 U8076 ( .A1(n7472), .A2(n7473), .ZN(n7524) );
  XNOR2_X1 U8077 ( .A(n7531), .B(n8237), .ZN(n7473) );
  OR2_X1 U8078 ( .A1(n8266), .A2(n8267), .ZN(n8237) );
  AND2_X1 U8079 ( .A1(n8268), .A2(n8269), .ZN(n8267) );
  AND2_X1 U8080 ( .A1(n8270), .A2(n8271), .ZN(n8266) );
  OR2_X1 U8081 ( .A1(n8269), .A2(n8268), .ZN(n8271) );
  XNOR2_X1 U8082 ( .A(n8247), .B(n8272), .ZN(n7531) );
  XOR2_X1 U8083 ( .A(n8246), .B(n8245), .Z(n8272) );
  OR2_X1 U8084 ( .A1(n7872), .A2(n7950), .ZN(n8245) );
  OR2_X1 U8085 ( .A1(n8273), .A2(n8274), .ZN(n8246) );
  AND2_X1 U8086 ( .A1(n8275), .A2(n8276), .ZN(n8274) );
  AND2_X1 U8087 ( .A1(n8277), .A2(n8278), .ZN(n8273) );
  OR2_X1 U8088 ( .A1(n8276), .A2(n8275), .ZN(n8278) );
  XOR2_X1 U8089 ( .A(n8254), .B(n8279), .Z(n8247) );
  XOR2_X1 U8090 ( .A(n8253), .B(n8252), .Z(n8279) );
  OR2_X1 U8091 ( .A1(n7964), .A2(n7953), .ZN(n8252) );
  OR2_X1 U8092 ( .A1(n8280), .A2(n8281), .ZN(n8253) );
  AND2_X1 U8093 ( .A1(n8282), .A2(n8283), .ZN(n8281) );
  AND2_X1 U8094 ( .A1(n8284), .A2(n8285), .ZN(n8280) );
  OR2_X1 U8095 ( .A1(n8283), .A2(n8282), .ZN(n8285) );
  XOR2_X1 U8096 ( .A(n8261), .B(n8286), .Z(n8254) );
  XOR2_X1 U8097 ( .A(n8260), .B(n8259), .Z(n8286) );
  OR2_X1 U8098 ( .A1(n7901), .A2(n7956), .ZN(n8259) );
  OR2_X1 U8099 ( .A1(n8287), .A2(n8288), .ZN(n8260) );
  AND2_X1 U8100 ( .A1(n7961), .A2(n8289), .ZN(n8288) );
  AND2_X1 U8101 ( .A1(n8290), .A2(n8291), .ZN(n8287) );
  OR2_X1 U8102 ( .A1(n8289), .A2(n7961), .ZN(n8291) );
  INV_X1 U8103 ( .A(n7905), .ZN(n7961) );
  XOR2_X1 U8104 ( .A(n8292), .B(n8293), .Z(n8261) );
  XOR2_X1 U8105 ( .A(n8294), .B(n8295), .Z(n8293) );
  OR2_X1 U8106 ( .A1(n8296), .A2(n8297), .ZN(n7472) );
  OR2_X1 U8107 ( .A1(n8298), .A2(n7470), .ZN(n8296) );
  AND3_X1 U8108 ( .A1(n7469), .A2(n7468), .A3(n7466), .ZN(n7470) );
  INV_X1 U8109 ( .A(n8299), .ZN(n7468) );
  AND2_X1 U8110 ( .A1(n7462), .A2(n7466), .ZN(n8298) );
  INV_X1 U8111 ( .A(n8300), .ZN(n7466) );
  OR2_X1 U8112 ( .A1(n8301), .A2(n8297), .ZN(n8300) );
  INV_X1 U8113 ( .A(n8302), .ZN(n8297) );
  OR2_X1 U8114 ( .A1(n8303), .A2(n8304), .ZN(n8302) );
  AND2_X1 U8115 ( .A1(n8303), .A2(n8304), .ZN(n8301) );
  OR2_X1 U8116 ( .A1(n8305), .A2(n8306), .ZN(n8304) );
  AND2_X1 U8117 ( .A1(n8307), .A2(n8308), .ZN(n8306) );
  AND2_X1 U8118 ( .A1(n8309), .A2(n8310), .ZN(n8305) );
  OR2_X1 U8119 ( .A1(n8308), .A2(n8307), .ZN(n8310) );
  XOR2_X1 U8120 ( .A(n8270), .B(n8311), .Z(n8303) );
  XOR2_X1 U8121 ( .A(n8269), .B(n8268), .Z(n8311) );
  OR2_X1 U8122 ( .A1(n7971), .A2(n7950), .ZN(n8268) );
  OR2_X1 U8123 ( .A1(n8312), .A2(n8313), .ZN(n8269) );
  AND2_X1 U8124 ( .A1(n8314), .A2(n8315), .ZN(n8313) );
  AND2_X1 U8125 ( .A1(n8316), .A2(n8317), .ZN(n8312) );
  OR2_X1 U8126 ( .A1(n8315), .A2(n8314), .ZN(n8317) );
  XOR2_X1 U8127 ( .A(n8277), .B(n8318), .Z(n8270) );
  XOR2_X1 U8128 ( .A(n8276), .B(n8275), .Z(n8318) );
  OR2_X1 U8129 ( .A1(n7872), .A2(n7953), .ZN(n8275) );
  OR2_X1 U8130 ( .A1(n8319), .A2(n8320), .ZN(n8276) );
  AND2_X1 U8131 ( .A1(n8321), .A2(n8322), .ZN(n8320) );
  AND2_X1 U8132 ( .A1(n8323), .A2(n8324), .ZN(n8319) );
  OR2_X1 U8133 ( .A1(n8322), .A2(n8321), .ZN(n8324) );
  XOR2_X1 U8134 ( .A(n8284), .B(n8325), .Z(n8277) );
  XOR2_X1 U8135 ( .A(n8283), .B(n8282), .Z(n8325) );
  OR2_X1 U8136 ( .A1(n7964), .A2(n7956), .ZN(n8282) );
  OR2_X1 U8137 ( .A1(n8326), .A2(n8327), .ZN(n8283) );
  AND2_X1 U8138 ( .A1(n8328), .A2(n8329), .ZN(n8327) );
  AND2_X1 U8139 ( .A1(n8330), .A2(n8331), .ZN(n8326) );
  OR2_X1 U8140 ( .A1(n8329), .A2(n8328), .ZN(n8331) );
  XOR2_X1 U8141 ( .A(n8290), .B(n8332), .Z(n8284) );
  XNOR2_X1 U8142 ( .A(n8289), .B(n7905), .ZN(n8332) );
  AND2_X1 U8143 ( .A1(b_3_), .A2(a_3_), .ZN(n7905) );
  OR2_X1 U8144 ( .A1(n8333), .A2(n8334), .ZN(n8289) );
  AND2_X1 U8145 ( .A1(n8335), .A2(n8336), .ZN(n8334) );
  AND2_X1 U8146 ( .A1(n8337), .A2(n8338), .ZN(n8333) );
  OR2_X1 U8147 ( .A1(n8336), .A2(n8335), .ZN(n8338) );
  XOR2_X1 U8148 ( .A(n8339), .B(n8340), .Z(n8290) );
  XOR2_X1 U8149 ( .A(n8341), .B(n8342), .Z(n8340) );
  AND2_X1 U8150 ( .A1(n7459), .A2(n7460), .ZN(n7462) );
  XNOR2_X1 U8151 ( .A(n7469), .B(n8299), .ZN(n7460) );
  OR2_X1 U8152 ( .A1(n8343), .A2(n8344), .ZN(n8299) );
  AND2_X1 U8153 ( .A1(n8345), .A2(n8346), .ZN(n8344) );
  AND2_X1 U8154 ( .A1(n8347), .A2(n8348), .ZN(n8343) );
  OR2_X1 U8155 ( .A1(n8346), .A2(n8345), .ZN(n8348) );
  XNOR2_X1 U8156 ( .A(n8309), .B(n8349), .ZN(n7469) );
  XOR2_X1 U8157 ( .A(n8308), .B(n8307), .Z(n8349) );
  OR2_X1 U8158 ( .A1(n7843), .A2(n7950), .ZN(n8307) );
  OR2_X1 U8159 ( .A1(n8350), .A2(n8351), .ZN(n8308) );
  AND2_X1 U8160 ( .A1(n8352), .A2(n8353), .ZN(n8351) );
  AND2_X1 U8161 ( .A1(n8354), .A2(n8355), .ZN(n8350) );
  OR2_X1 U8162 ( .A1(n8353), .A2(n8352), .ZN(n8355) );
  XOR2_X1 U8163 ( .A(n8316), .B(n8356), .Z(n8309) );
  XOR2_X1 U8164 ( .A(n8315), .B(n8314), .Z(n8356) );
  OR2_X1 U8165 ( .A1(n7971), .A2(n7953), .ZN(n8314) );
  OR2_X1 U8166 ( .A1(n8357), .A2(n8358), .ZN(n8315) );
  AND2_X1 U8167 ( .A1(n8359), .A2(n8360), .ZN(n8358) );
  AND2_X1 U8168 ( .A1(n8361), .A2(n8362), .ZN(n8357) );
  OR2_X1 U8169 ( .A1(n8360), .A2(n8359), .ZN(n8362) );
  XOR2_X1 U8170 ( .A(n8323), .B(n8363), .Z(n8316) );
  XOR2_X1 U8171 ( .A(n8322), .B(n8321), .Z(n8363) );
  OR2_X1 U8172 ( .A1(n7872), .A2(n7956), .ZN(n8321) );
  OR2_X1 U8173 ( .A1(n8364), .A2(n8365), .ZN(n8322) );
  AND2_X1 U8174 ( .A1(n8366), .A2(n8367), .ZN(n8365) );
  AND2_X1 U8175 ( .A1(n8368), .A2(n8369), .ZN(n8364) );
  OR2_X1 U8176 ( .A1(n8367), .A2(n8366), .ZN(n8369) );
  XOR2_X1 U8177 ( .A(n8330), .B(n8370), .Z(n8323) );
  XOR2_X1 U8178 ( .A(n8329), .B(n8328), .Z(n8370) );
  OR2_X1 U8179 ( .A1(n7964), .A2(n7960), .ZN(n8328) );
  OR2_X1 U8180 ( .A1(n8371), .A2(n8372), .ZN(n8329) );
  AND2_X1 U8181 ( .A1(n8373), .A2(n7965), .ZN(n8372) );
  AND2_X1 U8182 ( .A1(n8374), .A2(n8375), .ZN(n8371) );
  OR2_X1 U8183 ( .A1(n7965), .A2(n8373), .ZN(n8375) );
  XOR2_X1 U8184 ( .A(n8337), .B(n8376), .Z(n8330) );
  XOR2_X1 U8185 ( .A(n8336), .B(n8335), .Z(n8376) );
  OR2_X1 U8186 ( .A1(n7901), .A2(n7963), .ZN(n8335) );
  OR2_X1 U8187 ( .A1(n8377), .A2(n8378), .ZN(n8336) );
  AND2_X1 U8188 ( .A1(n8379), .A2(n8380), .ZN(n8378) );
  AND2_X1 U8189 ( .A1(n8381), .A2(n8382), .ZN(n8377) );
  OR2_X1 U8190 ( .A1(n8380), .A2(n8379), .ZN(n8382) );
  XOR2_X1 U8191 ( .A(n8383), .B(n8384), .Z(n8337) );
  XOR2_X1 U8192 ( .A(n8385), .B(n8386), .Z(n8384) );
  OR2_X1 U8193 ( .A1(n8387), .A2(n8388), .ZN(n7459) );
  OR2_X1 U8194 ( .A1(n8389), .A2(n7457), .ZN(n8387) );
  AND3_X1 U8195 ( .A1(n7456), .A2(n7455), .A3(n7453), .ZN(n7457) );
  INV_X1 U8196 ( .A(n8390), .ZN(n7455) );
  AND2_X1 U8197 ( .A1(n7449), .A2(n7453), .ZN(n8389) );
  INV_X1 U8198 ( .A(n8391), .ZN(n7453) );
  OR2_X1 U8199 ( .A1(n8392), .A2(n8388), .ZN(n8391) );
  INV_X1 U8200 ( .A(n8393), .ZN(n8388) );
  OR2_X1 U8201 ( .A1(n8394), .A2(n8395), .ZN(n8393) );
  AND2_X1 U8202 ( .A1(n8394), .A2(n8395), .ZN(n8392) );
  OR2_X1 U8203 ( .A1(n8396), .A2(n8397), .ZN(n8395) );
  AND2_X1 U8204 ( .A1(n8398), .A2(n8399), .ZN(n8397) );
  AND2_X1 U8205 ( .A1(n8400), .A2(n8401), .ZN(n8396) );
  OR2_X1 U8206 ( .A1(n8399), .A2(n8398), .ZN(n8401) );
  XOR2_X1 U8207 ( .A(n8347), .B(n8402), .Z(n8394) );
  XOR2_X1 U8208 ( .A(n8346), .B(n8345), .Z(n8402) );
  OR2_X1 U8209 ( .A1(n7978), .A2(n7950), .ZN(n8345) );
  OR2_X1 U8210 ( .A1(n8403), .A2(n8404), .ZN(n8346) );
  AND2_X1 U8211 ( .A1(n8405), .A2(n8406), .ZN(n8404) );
  AND2_X1 U8212 ( .A1(n8407), .A2(n8408), .ZN(n8403) );
  OR2_X1 U8213 ( .A1(n8406), .A2(n8405), .ZN(n8408) );
  XOR2_X1 U8214 ( .A(n8354), .B(n8409), .Z(n8347) );
  XOR2_X1 U8215 ( .A(n8353), .B(n8352), .Z(n8409) );
  OR2_X1 U8216 ( .A1(n7843), .A2(n7953), .ZN(n8352) );
  OR2_X1 U8217 ( .A1(n8410), .A2(n8411), .ZN(n8353) );
  AND2_X1 U8218 ( .A1(n8412), .A2(n8413), .ZN(n8411) );
  AND2_X1 U8219 ( .A1(n8414), .A2(n8415), .ZN(n8410) );
  OR2_X1 U8220 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  XOR2_X1 U8221 ( .A(n8361), .B(n8416), .Z(n8354) );
  XOR2_X1 U8222 ( .A(n8360), .B(n8359), .Z(n8416) );
  OR2_X1 U8223 ( .A1(n7971), .A2(n7956), .ZN(n8359) );
  OR2_X1 U8224 ( .A1(n8417), .A2(n8418), .ZN(n8360) );
  AND2_X1 U8225 ( .A1(n8419), .A2(n8420), .ZN(n8418) );
  AND2_X1 U8226 ( .A1(n8421), .A2(n8422), .ZN(n8417) );
  OR2_X1 U8227 ( .A1(n8420), .A2(n8419), .ZN(n8422) );
  XOR2_X1 U8228 ( .A(n8368), .B(n8423), .Z(n8361) );
  XOR2_X1 U8229 ( .A(n8367), .B(n8366), .Z(n8423) );
  OR2_X1 U8230 ( .A1(n7872), .A2(n7960), .ZN(n8366) );
  OR2_X1 U8231 ( .A1(n8424), .A2(n8425), .ZN(n8367) );
  AND2_X1 U8232 ( .A1(n8426), .A2(n8427), .ZN(n8425) );
  AND2_X1 U8233 ( .A1(n8428), .A2(n8429), .ZN(n8424) );
  OR2_X1 U8234 ( .A1(n8427), .A2(n8426), .ZN(n8429) );
  XNOR2_X1 U8235 ( .A(n8430), .B(n8374), .ZN(n8368) );
  XOR2_X1 U8236 ( .A(n8381), .B(n8431), .Z(n8374) );
  XOR2_X1 U8237 ( .A(n8380), .B(n8379), .Z(n8431) );
  OR2_X1 U8238 ( .A1(n7901), .A2(n7967), .ZN(n8379) );
  OR2_X1 U8239 ( .A1(n8432), .A2(n8433), .ZN(n8380) );
  AND2_X1 U8240 ( .A1(n8434), .A2(n8435), .ZN(n8433) );
  AND2_X1 U8241 ( .A1(n8436), .A2(n8437), .ZN(n8432) );
  OR2_X1 U8242 ( .A1(n8435), .A2(n8434), .ZN(n8437) );
  XOR2_X1 U8243 ( .A(n8438), .B(n8439), .Z(n8381) );
  XOR2_X1 U8244 ( .A(n8440), .B(n8441), .Z(n8439) );
  XNOR2_X1 U8245 ( .A(n7965), .B(n8373), .ZN(n8430) );
  OR2_X1 U8246 ( .A1(n8442), .A2(n8443), .ZN(n8373) );
  AND2_X1 U8247 ( .A1(n8444), .A2(n8445), .ZN(n8443) );
  AND2_X1 U8248 ( .A1(n8446), .A2(n8447), .ZN(n8442) );
  OR2_X1 U8249 ( .A1(n8445), .A2(n8444), .ZN(n8447) );
  INV_X1 U8250 ( .A(n7893), .ZN(n7965) );
  AND2_X1 U8251 ( .A1(b_4_), .A2(a_4_), .ZN(n7893) );
  AND2_X1 U8252 ( .A1(n8191), .A2(n8192), .ZN(n7449) );
  XNOR2_X1 U8253 ( .A(n7456), .B(n8390), .ZN(n8192) );
  OR2_X1 U8254 ( .A1(n8448), .A2(n8449), .ZN(n8390) );
  AND2_X1 U8255 ( .A1(n8450), .A2(n8451), .ZN(n8449) );
  AND2_X1 U8256 ( .A1(n8452), .A2(n8453), .ZN(n8448) );
  OR2_X1 U8257 ( .A1(n8451), .A2(n8450), .ZN(n8453) );
  XNOR2_X1 U8258 ( .A(n8400), .B(n8454), .ZN(n7456) );
  XOR2_X1 U8259 ( .A(n8399), .B(n8398), .Z(n8454) );
  OR2_X1 U8260 ( .A1(n7804), .A2(n7950), .ZN(n8398) );
  OR2_X1 U8261 ( .A1(n8455), .A2(n8456), .ZN(n8399) );
  AND2_X1 U8262 ( .A1(n8457), .A2(n8458), .ZN(n8456) );
  AND2_X1 U8263 ( .A1(n8459), .A2(n8460), .ZN(n8455) );
  OR2_X1 U8264 ( .A1(n8458), .A2(n8457), .ZN(n8460) );
  XOR2_X1 U8265 ( .A(n8407), .B(n8461), .Z(n8400) );
  XOR2_X1 U8266 ( .A(n8406), .B(n8405), .Z(n8461) );
  OR2_X1 U8267 ( .A1(n7978), .A2(n7953), .ZN(n8405) );
  OR2_X1 U8268 ( .A1(n8462), .A2(n8463), .ZN(n8406) );
  AND2_X1 U8269 ( .A1(n8464), .A2(n8465), .ZN(n8463) );
  AND2_X1 U8270 ( .A1(n8466), .A2(n8467), .ZN(n8462) );
  OR2_X1 U8271 ( .A1(n8465), .A2(n8464), .ZN(n8467) );
  XOR2_X1 U8272 ( .A(n8414), .B(n8468), .Z(n8407) );
  XOR2_X1 U8273 ( .A(n8413), .B(n8412), .Z(n8468) );
  OR2_X1 U8274 ( .A1(n7843), .A2(n7956), .ZN(n8412) );
  OR2_X1 U8275 ( .A1(n8469), .A2(n8470), .ZN(n8413) );
  AND2_X1 U8276 ( .A1(n8471), .A2(n8472), .ZN(n8470) );
  AND2_X1 U8277 ( .A1(n8473), .A2(n8474), .ZN(n8469) );
  OR2_X1 U8278 ( .A1(n8472), .A2(n8471), .ZN(n8474) );
  XOR2_X1 U8279 ( .A(n8421), .B(n8475), .Z(n8414) );
  XOR2_X1 U8280 ( .A(n8420), .B(n8419), .Z(n8475) );
  OR2_X1 U8281 ( .A1(n7971), .A2(n7960), .ZN(n8419) );
  OR2_X1 U8282 ( .A1(n8476), .A2(n8477), .ZN(n8420) );
  AND2_X1 U8283 ( .A1(n8478), .A2(n8479), .ZN(n8477) );
  AND2_X1 U8284 ( .A1(n8480), .A2(n8481), .ZN(n8476) );
  OR2_X1 U8285 ( .A1(n8479), .A2(n8478), .ZN(n8481) );
  XOR2_X1 U8286 ( .A(n8428), .B(n8482), .Z(n8421) );
  XOR2_X1 U8287 ( .A(n8427), .B(n8426), .Z(n8482) );
  OR2_X1 U8288 ( .A1(n7872), .A2(n7963), .ZN(n8426) );
  OR2_X1 U8289 ( .A1(n8483), .A2(n8484), .ZN(n8427) );
  AND2_X1 U8290 ( .A1(n7968), .A2(n8485), .ZN(n8484) );
  AND2_X1 U8291 ( .A1(n8486), .A2(n8487), .ZN(n8483) );
  OR2_X1 U8292 ( .A1(n8485), .A2(n7968), .ZN(n8487) );
  INV_X1 U8293 ( .A(n7876), .ZN(n7968) );
  XOR2_X1 U8294 ( .A(n8446), .B(n8488), .Z(n8428) );
  XOR2_X1 U8295 ( .A(n8445), .B(n8444), .Z(n8488) );
  OR2_X1 U8296 ( .A1(n7964), .A2(n7967), .ZN(n8444) );
  OR2_X1 U8297 ( .A1(n8489), .A2(n8490), .ZN(n8445) );
  AND2_X1 U8298 ( .A1(n8491), .A2(n8492), .ZN(n8490) );
  AND2_X1 U8299 ( .A1(n8493), .A2(n8494), .ZN(n8489) );
  OR2_X1 U8300 ( .A1(n8492), .A2(n8491), .ZN(n8494) );
  XOR2_X1 U8301 ( .A(n8436), .B(n8495), .Z(n8446) );
  XOR2_X1 U8302 ( .A(n8435), .B(n8434), .Z(n8495) );
  OR2_X1 U8303 ( .A1(n7901), .A2(n7970), .ZN(n8434) );
  OR2_X1 U8304 ( .A1(n8496), .A2(n8497), .ZN(n8435) );
  AND2_X1 U8305 ( .A1(n8498), .A2(n8499), .ZN(n8497) );
  AND2_X1 U8306 ( .A1(n8500), .A2(n8501), .ZN(n8496) );
  OR2_X1 U8307 ( .A1(n8499), .A2(n8498), .ZN(n8501) );
  XOR2_X1 U8308 ( .A(n8502), .B(n8503), .Z(n8436) );
  XOR2_X1 U8309 ( .A(n8504), .B(n8505), .Z(n8503) );
  OR2_X1 U8310 ( .A1(n8506), .A2(n8507), .ZN(n8191) );
  OR2_X1 U8311 ( .A1(n8508), .A2(n8185), .ZN(n8507) );
  AND3_X1 U8312 ( .A1(n8189), .A2(n8188), .A3(n8187), .ZN(n8185) );
  INV_X1 U8313 ( .A(n8509), .ZN(n8188) );
  AND2_X1 U8314 ( .A1(n8181), .A2(n8187), .ZN(n8508) );
  INV_X1 U8315 ( .A(n8510), .ZN(n8187) );
  OR2_X1 U8316 ( .A1(n8511), .A2(n8506), .ZN(n8510) );
  AND2_X1 U8317 ( .A1(n8512), .A2(n8513), .ZN(n8511) );
  AND2_X1 U8318 ( .A1(n8178), .A2(n8179), .ZN(n8181) );
  XNOR2_X1 U8319 ( .A(n8189), .B(n8509), .ZN(n8179) );
  OR2_X1 U8320 ( .A1(n8514), .A2(n8515), .ZN(n8509) );
  AND2_X1 U8321 ( .A1(n8516), .A2(n8517), .ZN(n8515) );
  AND2_X1 U8322 ( .A1(n8518), .A2(n8519), .ZN(n8514) );
  OR2_X1 U8323 ( .A1(n8517), .A2(n8516), .ZN(n8519) );
  XNOR2_X1 U8324 ( .A(n8520), .B(n8521), .ZN(n8189) );
  XOR2_X1 U8325 ( .A(n8522), .B(n8523), .Z(n8521) );
  OR2_X1 U8326 ( .A1(n8524), .A2(n8525), .ZN(n8178) );
  OR2_X1 U8327 ( .A1(n8526), .A2(n8172), .ZN(n8525) );
  AND3_X1 U8328 ( .A1(n8176), .A2(n8175), .A3(n8174), .ZN(n8172) );
  INV_X1 U8329 ( .A(n8527), .ZN(n8175) );
  AND2_X1 U8330 ( .A1(n8174), .A2(n8168), .ZN(n8526) );
  OR2_X1 U8331 ( .A1(n8528), .A2(n8162), .ZN(n8168) );
  AND3_X1 U8332 ( .A1(n8166), .A2(n8164), .A3(n8165), .ZN(n8162) );
  AND2_X1 U8333 ( .A1(n8164), .A2(n8158), .ZN(n8528) );
  OR2_X1 U8334 ( .A1(n8529), .A2(n8530), .ZN(n8158) );
  INV_X1 U8335 ( .A(n8156), .ZN(n8530) );
  OR3_X1 U8336 ( .A1(n8531), .A2(n8532), .A3(n8533), .ZN(n8156) );
  AND2_X1 U8337 ( .A1(n8153), .A2(n8155), .ZN(n8529) );
  INV_X1 U8338 ( .A(n8534), .ZN(n8155) );
  AND2_X1 U8339 ( .A1(n8535), .A2(n8532), .ZN(n8534) );
  XNOR2_X1 U8340 ( .A(n8166), .B(n8165), .ZN(n8532) );
  INV_X1 U8341 ( .A(n8536), .ZN(n8165) );
  OR2_X1 U8342 ( .A1(n8537), .A2(n8538), .ZN(n8536) );
  AND2_X1 U8343 ( .A1(n8539), .A2(n8540), .ZN(n8538) );
  AND2_X1 U8344 ( .A1(n8541), .A2(n8542), .ZN(n8537) );
  OR2_X1 U8345 ( .A1(n8540), .A2(n8539), .ZN(n8542) );
  XNOR2_X1 U8346 ( .A(n8543), .B(n8544), .ZN(n8166) );
  XOR2_X1 U8347 ( .A(n8545), .B(n8546), .Z(n8544) );
  OR2_X1 U8348 ( .A1(n8533), .A2(n8531), .ZN(n8535) );
  OR2_X1 U8349 ( .A1(n8547), .A2(n8548), .ZN(n8153) );
  INV_X1 U8350 ( .A(n8150), .ZN(n8548) );
  OR3_X1 U8351 ( .A1(n8549), .A2(n8550), .A3(n8551), .ZN(n8150) );
  AND2_X1 U8352 ( .A1(n8148), .A2(n8151), .ZN(n8547) );
  INV_X1 U8353 ( .A(n8552), .ZN(n8151) );
  AND2_X1 U8354 ( .A1(n8553), .A2(n8550), .ZN(n8552) );
  XNOR2_X1 U8355 ( .A(n8531), .B(n8533), .ZN(n8550) );
  OR2_X1 U8356 ( .A1(n8554), .A2(n8555), .ZN(n8533) );
  AND2_X1 U8357 ( .A1(n8556), .A2(n8557), .ZN(n8555) );
  AND2_X1 U8358 ( .A1(n8558), .A2(n8559), .ZN(n8554) );
  OR2_X1 U8359 ( .A1(n8556), .A2(n8557), .ZN(n8559) );
  XOR2_X1 U8360 ( .A(n8541), .B(n8560), .Z(n8531) );
  XOR2_X1 U8361 ( .A(n8540), .B(n8539), .Z(n8560) );
  OR2_X1 U8362 ( .A1(n7950), .A2(n7717), .ZN(n8539) );
  OR2_X1 U8363 ( .A1(n8561), .A2(n8562), .ZN(n8540) );
  AND2_X1 U8364 ( .A1(n8563), .A2(n8564), .ZN(n8562) );
  AND2_X1 U8365 ( .A1(n8565), .A2(n8566), .ZN(n8561) );
  OR2_X1 U8366 ( .A1(n8564), .A2(n8563), .ZN(n8566) );
  XOR2_X1 U8367 ( .A(n8567), .B(n8568), .Z(n8541) );
  XOR2_X1 U8368 ( .A(n8569), .B(n8570), .Z(n8568) );
  OR2_X1 U8369 ( .A1(n8551), .A2(n8549), .ZN(n8553) );
  OR2_X1 U8370 ( .A1(n8571), .A2(n8572), .ZN(n8148) );
  INV_X1 U8371 ( .A(n8145), .ZN(n8572) );
  OR3_X1 U8372 ( .A1(n8573), .A2(n8574), .A3(n8575), .ZN(n8145) );
  AND2_X1 U8373 ( .A1(n8143), .A2(n8146), .ZN(n8571) );
  INV_X1 U8374 ( .A(n8576), .ZN(n8146) );
  AND2_X1 U8375 ( .A1(n8577), .A2(n8574), .ZN(n8576) );
  XNOR2_X1 U8376 ( .A(n8549), .B(n8551), .ZN(n8574) );
  OR2_X1 U8377 ( .A1(n8578), .A2(n8579), .ZN(n8551) );
  AND2_X1 U8378 ( .A1(n8580), .A2(n8581), .ZN(n8579) );
  AND2_X1 U8379 ( .A1(n8582), .A2(n8583), .ZN(n8578) );
  OR2_X1 U8380 ( .A1(n8580), .A2(n8581), .ZN(n8583) );
  XOR2_X1 U8381 ( .A(n8558), .B(n8584), .Z(n8549) );
  XOR2_X1 U8382 ( .A(n8557), .B(n8556), .Z(n8584) );
  OR2_X1 U8383 ( .A1(n7950), .A2(n8006), .ZN(n8556) );
  OR2_X1 U8384 ( .A1(n8585), .A2(n8586), .ZN(n8557) );
  AND2_X1 U8385 ( .A1(n8587), .A2(n8588), .ZN(n8586) );
  AND2_X1 U8386 ( .A1(n8589), .A2(n8590), .ZN(n8585) );
  OR2_X1 U8387 ( .A1(n8587), .A2(n8588), .ZN(n8590) );
  XOR2_X1 U8388 ( .A(n8565), .B(n8591), .Z(n8558) );
  XOR2_X1 U8389 ( .A(n8564), .B(n8563), .Z(n8591) );
  OR2_X1 U8390 ( .A1(n7953), .A2(n7717), .ZN(n8563) );
  OR2_X1 U8391 ( .A1(n8592), .A2(n8593), .ZN(n8564) );
  AND2_X1 U8392 ( .A1(n8594), .A2(n8595), .ZN(n8593) );
  AND2_X1 U8393 ( .A1(n8596), .A2(n8597), .ZN(n8592) );
  OR2_X1 U8394 ( .A1(n8595), .A2(n8594), .ZN(n8597) );
  XOR2_X1 U8395 ( .A(n8598), .B(n8599), .Z(n8565) );
  XOR2_X1 U8396 ( .A(n8600), .B(n8601), .Z(n8599) );
  OR2_X1 U8397 ( .A1(n8575), .A2(n8573), .ZN(n8577) );
  OR2_X1 U8398 ( .A1(n8602), .A2(n8603), .ZN(n8143) );
  INV_X1 U8399 ( .A(n8141), .ZN(n8603) );
  OR3_X1 U8400 ( .A1(n8604), .A2(n8605), .A3(n8606), .ZN(n8141) );
  AND2_X1 U8401 ( .A1(n8138), .A2(n8140), .ZN(n8602) );
  INV_X1 U8402 ( .A(n8607), .ZN(n8140) );
  AND2_X1 U8403 ( .A1(n8608), .A2(n8605), .ZN(n8607) );
  XNOR2_X1 U8404 ( .A(n8573), .B(n8575), .ZN(n8605) );
  OR2_X1 U8405 ( .A1(n8609), .A2(n8610), .ZN(n8575) );
  AND2_X1 U8406 ( .A1(n8611), .A2(n8612), .ZN(n8610) );
  AND2_X1 U8407 ( .A1(n8613), .A2(n8614), .ZN(n8609) );
  OR2_X1 U8408 ( .A1(n8611), .A2(n8612), .ZN(n8614) );
  XOR2_X1 U8409 ( .A(n8582), .B(n8615), .Z(n8573) );
  XOR2_X1 U8410 ( .A(n8581), .B(n8580), .Z(n8615) );
  OR2_X1 U8411 ( .A1(n7950), .A2(n7688), .ZN(n8580) );
  OR2_X1 U8412 ( .A1(n8616), .A2(n8617), .ZN(n8581) );
  AND2_X1 U8413 ( .A1(n8618), .A2(n8619), .ZN(n8617) );
  AND2_X1 U8414 ( .A1(n8620), .A2(n8621), .ZN(n8616) );
  OR2_X1 U8415 ( .A1(n8618), .A2(n8619), .ZN(n8621) );
  XOR2_X1 U8416 ( .A(n8589), .B(n8622), .Z(n8582) );
  XOR2_X1 U8417 ( .A(n8588), .B(n8587), .Z(n8622) );
  OR2_X1 U8418 ( .A1(n7953), .A2(n8006), .ZN(n8587) );
  OR2_X1 U8419 ( .A1(n8623), .A2(n8624), .ZN(n8588) );
  AND2_X1 U8420 ( .A1(n8625), .A2(n8626), .ZN(n8624) );
  AND2_X1 U8421 ( .A1(n8627), .A2(n8628), .ZN(n8623) );
  OR2_X1 U8422 ( .A1(n8625), .A2(n8626), .ZN(n8628) );
  XOR2_X1 U8423 ( .A(n8596), .B(n8629), .Z(n8589) );
  XOR2_X1 U8424 ( .A(n8595), .B(n8594), .Z(n8629) );
  OR2_X1 U8425 ( .A1(n7956), .A2(n7717), .ZN(n8594) );
  OR2_X1 U8426 ( .A1(n8630), .A2(n8631), .ZN(n8595) );
  AND2_X1 U8427 ( .A1(n8632), .A2(n8633), .ZN(n8631) );
  AND2_X1 U8428 ( .A1(n8634), .A2(n8635), .ZN(n8630) );
  OR2_X1 U8429 ( .A1(n8633), .A2(n8632), .ZN(n8635) );
  XOR2_X1 U8430 ( .A(n8636), .B(n8637), .Z(n8596) );
  XOR2_X1 U8431 ( .A(n8638), .B(n8639), .Z(n8637) );
  OR2_X1 U8432 ( .A1(n8606), .A2(n8604), .ZN(n8608) );
  OR2_X1 U8433 ( .A1(n8640), .A2(n8641), .ZN(n8138) );
  INV_X1 U8434 ( .A(n8135), .ZN(n8641) );
  OR3_X1 U8435 ( .A1(n8642), .A2(n8643), .A3(n8644), .ZN(n8135) );
  AND2_X1 U8436 ( .A1(n8133), .A2(n8136), .ZN(n8640) );
  INV_X1 U8437 ( .A(n8645), .ZN(n8136) );
  AND2_X1 U8438 ( .A1(n8646), .A2(n8643), .ZN(n8645) );
  XNOR2_X1 U8439 ( .A(n8604), .B(n8606), .ZN(n8643) );
  OR2_X1 U8440 ( .A1(n8647), .A2(n8648), .ZN(n8606) );
  AND2_X1 U8441 ( .A1(n8649), .A2(n8650), .ZN(n8648) );
  AND2_X1 U8442 ( .A1(n8651), .A2(n8652), .ZN(n8647) );
  OR2_X1 U8443 ( .A1(n8649), .A2(n8650), .ZN(n8652) );
  XOR2_X1 U8444 ( .A(n8613), .B(n8653), .Z(n8604) );
  XOR2_X1 U8445 ( .A(n8612), .B(n8611), .Z(n8653) );
  OR2_X1 U8446 ( .A1(n7950), .A2(n8013), .ZN(n8611) );
  OR2_X1 U8447 ( .A1(n8654), .A2(n8655), .ZN(n8612) );
  AND2_X1 U8448 ( .A1(n8656), .A2(n8657), .ZN(n8655) );
  AND2_X1 U8449 ( .A1(n8658), .A2(n8659), .ZN(n8654) );
  OR2_X1 U8450 ( .A1(n8656), .A2(n8657), .ZN(n8659) );
  XOR2_X1 U8451 ( .A(n8620), .B(n8660), .Z(n8613) );
  XOR2_X1 U8452 ( .A(n8619), .B(n8618), .Z(n8660) );
  OR2_X1 U8453 ( .A1(n7953), .A2(n7688), .ZN(n8618) );
  OR2_X1 U8454 ( .A1(n8661), .A2(n8662), .ZN(n8619) );
  AND2_X1 U8455 ( .A1(n8663), .A2(n8664), .ZN(n8662) );
  AND2_X1 U8456 ( .A1(n8665), .A2(n8666), .ZN(n8661) );
  OR2_X1 U8457 ( .A1(n8663), .A2(n8664), .ZN(n8666) );
  XOR2_X1 U8458 ( .A(n8627), .B(n8667), .Z(n8620) );
  XOR2_X1 U8459 ( .A(n8626), .B(n8625), .Z(n8667) );
  OR2_X1 U8460 ( .A1(n7956), .A2(n8006), .ZN(n8625) );
  OR2_X1 U8461 ( .A1(n8668), .A2(n8669), .ZN(n8626) );
  AND2_X1 U8462 ( .A1(n8670), .A2(n8671), .ZN(n8669) );
  AND2_X1 U8463 ( .A1(n8672), .A2(n8673), .ZN(n8668) );
  OR2_X1 U8464 ( .A1(n8670), .A2(n8671), .ZN(n8673) );
  XOR2_X1 U8465 ( .A(n8634), .B(n8674), .Z(n8627) );
  XOR2_X1 U8466 ( .A(n8633), .B(n8632), .Z(n8674) );
  OR2_X1 U8467 ( .A1(n7960), .A2(n7717), .ZN(n8632) );
  OR2_X1 U8468 ( .A1(n8675), .A2(n8676), .ZN(n8633) );
  AND2_X1 U8469 ( .A1(n8677), .A2(n8678), .ZN(n8676) );
  AND2_X1 U8470 ( .A1(n8679), .A2(n8680), .ZN(n8675) );
  OR2_X1 U8471 ( .A1(n8678), .A2(n8677), .ZN(n8680) );
  XOR2_X1 U8472 ( .A(n8681), .B(n8682), .Z(n8634) );
  XOR2_X1 U8473 ( .A(n8683), .B(n8684), .Z(n8682) );
  OR2_X1 U8474 ( .A1(n8644), .A2(n8642), .ZN(n8646) );
  OR2_X1 U8475 ( .A1(n8685), .A2(n8686), .ZN(n8133) );
  INV_X1 U8476 ( .A(n8120), .ZN(n8686) );
  OR3_X1 U8477 ( .A1(n8687), .A2(n8688), .A3(n8689), .ZN(n8120) );
  AND2_X1 U8478 ( .A1(n8118), .A2(n8121), .ZN(n8685) );
  INV_X1 U8479 ( .A(n8690), .ZN(n8121) );
  AND2_X1 U8480 ( .A1(n8691), .A2(n8688), .ZN(n8690) );
  XNOR2_X1 U8481 ( .A(n8642), .B(n8644), .ZN(n8688) );
  OR2_X1 U8482 ( .A1(n8692), .A2(n8693), .ZN(n8644) );
  AND2_X1 U8483 ( .A1(n8694), .A2(n8695), .ZN(n8693) );
  AND2_X1 U8484 ( .A1(n8696), .A2(n8697), .ZN(n8692) );
  OR2_X1 U8485 ( .A1(n8694), .A2(n8695), .ZN(n8697) );
  XOR2_X1 U8486 ( .A(n8651), .B(n8698), .Z(n8642) );
  XOR2_X1 U8487 ( .A(n8650), .B(n8649), .Z(n8698) );
  OR2_X1 U8488 ( .A1(n7950), .A2(n7656), .ZN(n8649) );
  OR2_X1 U8489 ( .A1(n8699), .A2(n8700), .ZN(n8650) );
  AND2_X1 U8490 ( .A1(n8701), .A2(n8702), .ZN(n8700) );
  AND2_X1 U8491 ( .A1(n8703), .A2(n8704), .ZN(n8699) );
  OR2_X1 U8492 ( .A1(n8701), .A2(n8702), .ZN(n8704) );
  XOR2_X1 U8493 ( .A(n8658), .B(n8705), .Z(n8651) );
  XOR2_X1 U8494 ( .A(n8657), .B(n8656), .Z(n8705) );
  OR2_X1 U8495 ( .A1(n7953), .A2(n8013), .ZN(n8656) );
  OR2_X1 U8496 ( .A1(n8706), .A2(n8707), .ZN(n8657) );
  AND2_X1 U8497 ( .A1(n8708), .A2(n8709), .ZN(n8707) );
  AND2_X1 U8498 ( .A1(n8710), .A2(n8711), .ZN(n8706) );
  OR2_X1 U8499 ( .A1(n8708), .A2(n8709), .ZN(n8711) );
  XOR2_X1 U8500 ( .A(n8665), .B(n8712), .Z(n8658) );
  XOR2_X1 U8501 ( .A(n8664), .B(n8663), .Z(n8712) );
  OR2_X1 U8502 ( .A1(n7956), .A2(n7688), .ZN(n8663) );
  OR2_X1 U8503 ( .A1(n8713), .A2(n8714), .ZN(n8664) );
  AND2_X1 U8504 ( .A1(n8715), .A2(n8716), .ZN(n8714) );
  AND2_X1 U8505 ( .A1(n8717), .A2(n8718), .ZN(n8713) );
  OR2_X1 U8506 ( .A1(n8715), .A2(n8716), .ZN(n8718) );
  XOR2_X1 U8507 ( .A(n8672), .B(n8719), .Z(n8665) );
  XOR2_X1 U8508 ( .A(n8671), .B(n8670), .Z(n8719) );
  OR2_X1 U8509 ( .A1(n7960), .A2(n8006), .ZN(n8670) );
  OR2_X1 U8510 ( .A1(n8720), .A2(n8721), .ZN(n8671) );
  AND2_X1 U8511 ( .A1(n8722), .A2(n8723), .ZN(n8721) );
  AND2_X1 U8512 ( .A1(n8724), .A2(n8725), .ZN(n8720) );
  OR2_X1 U8513 ( .A1(n8722), .A2(n8723), .ZN(n8725) );
  XOR2_X1 U8514 ( .A(n8679), .B(n8726), .Z(n8672) );
  XOR2_X1 U8515 ( .A(n8678), .B(n8677), .Z(n8726) );
  OR2_X1 U8516 ( .A1(n7963), .A2(n7717), .ZN(n8677) );
  OR2_X1 U8517 ( .A1(n8727), .A2(n8728), .ZN(n8678) );
  AND2_X1 U8518 ( .A1(n8729), .A2(n8730), .ZN(n8728) );
  AND2_X1 U8519 ( .A1(n8731), .A2(n8732), .ZN(n8727) );
  OR2_X1 U8520 ( .A1(n8730), .A2(n8729), .ZN(n8732) );
  XOR2_X1 U8521 ( .A(n8733), .B(n8734), .Z(n8679) );
  XOR2_X1 U8522 ( .A(n8735), .B(n8736), .Z(n8734) );
  OR2_X1 U8523 ( .A1(n8689), .A2(n8687), .ZN(n8691) );
  OR2_X1 U8524 ( .A1(n8737), .A2(n8116), .ZN(n8118) );
  AND3_X1 U8525 ( .A1(n8738), .A2(n8739), .A3(n8740), .ZN(n8116) );
  AND2_X1 U8526 ( .A1(n8115), .A2(n8112), .ZN(n8737) );
  OR2_X1 U8527 ( .A1(n8741), .A2(n8742), .ZN(n8112) );
  INV_X1 U8528 ( .A(n8110), .ZN(n8742) );
  OR3_X1 U8529 ( .A1(n8743), .A2(n8744), .A3(n8745), .ZN(n8110) );
  AND2_X1 U8530 ( .A1(n8107), .A2(n8109), .ZN(n8741) );
  INV_X1 U8531 ( .A(n8746), .ZN(n8109) );
  AND2_X1 U8532 ( .A1(n8747), .A2(n8744), .ZN(n8746) );
  XNOR2_X1 U8533 ( .A(n8738), .B(n8740), .ZN(n8744) );
  OR2_X1 U8534 ( .A1(n8745), .A2(n8743), .ZN(n8747) );
  OR2_X1 U8535 ( .A1(n8748), .A2(n8749), .ZN(n8107) );
  INV_X1 U8536 ( .A(n8104), .ZN(n8749) );
  OR3_X1 U8537 ( .A1(n8750), .A2(n8751), .A3(n8752), .ZN(n8104) );
  AND2_X1 U8538 ( .A1(n8102), .A2(n8105), .ZN(n8748) );
  INV_X1 U8539 ( .A(n8753), .ZN(n8105) );
  AND2_X1 U8540 ( .A1(n8754), .A2(n8751), .ZN(n8753) );
  XNOR2_X1 U8541 ( .A(n8743), .B(n8745), .ZN(n8751) );
  OR2_X1 U8542 ( .A1(n8755), .A2(n8756), .ZN(n8745) );
  AND2_X1 U8543 ( .A1(n8757), .A2(n8758), .ZN(n8756) );
  AND2_X1 U8544 ( .A1(n8759), .A2(n8760), .ZN(n8755) );
  OR2_X1 U8545 ( .A1(n8757), .A2(n8758), .ZN(n8760) );
  XOR2_X1 U8546 ( .A(n8761), .B(n8762), .Z(n8743) );
  XOR2_X1 U8547 ( .A(n8763), .B(n8764), .Z(n8762) );
  OR2_X1 U8548 ( .A1(n8752), .A2(n8750), .ZN(n8754) );
  OR2_X1 U8549 ( .A1(n8765), .A2(n8766), .ZN(n8102) );
  INV_X1 U8550 ( .A(n8099), .ZN(n8766) );
  OR3_X1 U8551 ( .A1(n8767), .A2(n8768), .A3(n8769), .ZN(n8099) );
  AND2_X1 U8552 ( .A1(n8097), .A2(n8100), .ZN(n8765) );
  INV_X1 U8553 ( .A(n8770), .ZN(n8100) );
  AND2_X1 U8554 ( .A1(n8771), .A2(n8768), .ZN(n8770) );
  XNOR2_X1 U8555 ( .A(n8750), .B(n8752), .ZN(n8768) );
  OR2_X1 U8556 ( .A1(n8772), .A2(n8773), .ZN(n8752) );
  AND2_X1 U8557 ( .A1(n8774), .A2(n8775), .ZN(n8773) );
  AND2_X1 U8558 ( .A1(n8776), .A2(n8777), .ZN(n8772) );
  OR2_X1 U8559 ( .A1(n8774), .A2(n8775), .ZN(n8777) );
  XOR2_X1 U8560 ( .A(n8759), .B(n8778), .Z(n8750) );
  XOR2_X1 U8561 ( .A(n8758), .B(n8757), .Z(n8778) );
  OR2_X1 U8562 ( .A1(n7950), .A2(n7598), .ZN(n8757) );
  OR2_X1 U8563 ( .A1(n8779), .A2(n8780), .ZN(n8758) );
  AND2_X1 U8564 ( .A1(n8781), .A2(n8782), .ZN(n8780) );
  AND2_X1 U8565 ( .A1(n8783), .A2(n8784), .ZN(n8779) );
  OR2_X1 U8566 ( .A1(n8781), .A2(n8782), .ZN(n8784) );
  XOR2_X1 U8567 ( .A(n8785), .B(n8786), .Z(n8759) );
  XOR2_X1 U8568 ( .A(n8787), .B(n8788), .Z(n8786) );
  OR2_X1 U8569 ( .A1(n8769), .A2(n8767), .ZN(n8771) );
  OR2_X1 U8570 ( .A1(n8789), .A2(n8095), .ZN(n8097) );
  AND3_X1 U8571 ( .A1(n8790), .A2(n8791), .A3(n8792), .ZN(n8095) );
  AND2_X1 U8572 ( .A1(n8094), .A2(n8091), .ZN(n8789) );
  OR2_X1 U8573 ( .A1(n8793), .A2(n8089), .ZN(n8091) );
  AND2_X1 U8574 ( .A1(n8794), .A2(n8795), .ZN(n8089) );
  AND2_X1 U8575 ( .A1(n8087), .A2(n8085), .ZN(n8793) );
  OR2_X1 U8576 ( .A1(n8796), .A2(n8083), .ZN(n8085) );
  AND3_X1 U8577 ( .A1(n8797), .A2(n8798), .A3(n8799), .ZN(n8083) );
  AND2_X1 U8578 ( .A1(n8081), .A2(n8079), .ZN(n8796) );
  OR2_X1 U8579 ( .A1(n8800), .A2(n8077), .ZN(n8079) );
  AND3_X1 U8580 ( .A1(n8801), .A2(n8802), .A3(n8803), .ZN(n8077) );
  AND2_X1 U8581 ( .A1(n8075), .A2(n8073), .ZN(n8800) );
  OR2_X1 U8582 ( .A1(n8804), .A2(n8805), .ZN(n8073) );
  INV_X1 U8583 ( .A(n8070), .ZN(n8805) );
  OR3_X1 U8584 ( .A1(n8806), .A2(n8807), .A3(n8808), .ZN(n8070) );
  XNOR2_X1 U8585 ( .A(n8801), .B(n8803), .ZN(n8806) );
  AND2_X1 U8586 ( .A1(n8071), .A2(n8069), .ZN(n8804) );
  OR2_X1 U8587 ( .A1(n8809), .A2(n8810), .ZN(n8069) );
  XNOR2_X1 U8588 ( .A(n8811), .B(n8801), .ZN(n8810) );
  INV_X1 U8589 ( .A(n8812), .ZN(n8809) );
  OR2_X1 U8590 ( .A1(n8808), .A2(n8807), .ZN(n8812) );
  AND3_X1 U8591 ( .A1(n8058), .A2(n8062), .A3(n8063), .ZN(n8071) );
  INV_X1 U8592 ( .A(n8057), .ZN(n8063) );
  OR2_X1 U8593 ( .A1(n8813), .A2(n8814), .ZN(n8057) );
  AND2_X1 U8594 ( .A1(n7946), .A2(n7945), .ZN(n8814) );
  AND2_X1 U8595 ( .A1(n7943), .A2(n8815), .ZN(n8813) );
  OR2_X1 U8596 ( .A1(n7946), .A2(n7945), .ZN(n8815) );
  OR2_X1 U8597 ( .A1(n8816), .A2(n8817), .ZN(n7945) );
  AND2_X1 U8598 ( .A1(n7939), .A2(n7938), .ZN(n8817) );
  AND2_X1 U8599 ( .A1(n7936), .A2(n8818), .ZN(n8816) );
  OR2_X1 U8600 ( .A1(n7939), .A2(n7938), .ZN(n8818) );
  OR2_X1 U8601 ( .A1(n8819), .A2(n8820), .ZN(n7938) );
  AND2_X1 U8602 ( .A1(n7917), .A2(n7916), .ZN(n8820) );
  AND2_X1 U8603 ( .A1(n7914), .A2(n8821), .ZN(n8819) );
  OR2_X1 U8604 ( .A1(n7917), .A2(n7916), .ZN(n8821) );
  OR2_X1 U8605 ( .A1(n8822), .A2(n8823), .ZN(n7916) );
  AND2_X1 U8606 ( .A1(n7910), .A2(n7909), .ZN(n8823) );
  AND2_X1 U8607 ( .A1(n7907), .A2(n8824), .ZN(n8822) );
  OR2_X1 U8608 ( .A1(n7910), .A2(n7909), .ZN(n8824) );
  OR2_X1 U8609 ( .A1(n8825), .A2(n8826), .ZN(n7909) );
  AND2_X1 U8610 ( .A1(n7888), .A2(n7887), .ZN(n8826) );
  AND2_X1 U8611 ( .A1(n7885), .A2(n8827), .ZN(n8825) );
  OR2_X1 U8612 ( .A1(n7888), .A2(n7887), .ZN(n8827) );
  OR2_X1 U8613 ( .A1(n8828), .A2(n8829), .ZN(n7887) );
  AND2_X1 U8614 ( .A1(n7881), .A2(n7880), .ZN(n8829) );
  AND2_X1 U8615 ( .A1(n7878), .A2(n8830), .ZN(n8828) );
  OR2_X1 U8616 ( .A1(n7881), .A2(n7880), .ZN(n8830) );
  OR2_X1 U8617 ( .A1(n8831), .A2(n8832), .ZN(n7880) );
  AND2_X1 U8618 ( .A1(n7859), .A2(n7858), .ZN(n8832) );
  AND2_X1 U8619 ( .A1(n7856), .A2(n8833), .ZN(n8831) );
  OR2_X1 U8620 ( .A1(n7859), .A2(n7858), .ZN(n8833) );
  OR2_X1 U8621 ( .A1(n8834), .A2(n8835), .ZN(n7858) );
  AND2_X1 U8622 ( .A1(n7852), .A2(n7851), .ZN(n8835) );
  AND2_X1 U8623 ( .A1(n7849), .A2(n8836), .ZN(n8834) );
  OR2_X1 U8624 ( .A1(n7852), .A2(n7851), .ZN(n8836) );
  OR2_X1 U8625 ( .A1(n8837), .A2(n8838), .ZN(n7851) );
  AND2_X1 U8626 ( .A1(n7820), .A2(n7819), .ZN(n8838) );
  AND2_X1 U8627 ( .A1(n7817), .A2(n8839), .ZN(n8837) );
  OR2_X1 U8628 ( .A1(n7820), .A2(n7819), .ZN(n8839) );
  OR2_X1 U8629 ( .A1(n8840), .A2(n8841), .ZN(n7819) );
  AND2_X1 U8630 ( .A1(n7813), .A2(n7812), .ZN(n8841) );
  AND2_X1 U8631 ( .A1(n7810), .A2(n8842), .ZN(n8840) );
  OR2_X1 U8632 ( .A1(n7813), .A2(n7812), .ZN(n8842) );
  OR2_X1 U8633 ( .A1(n8843), .A2(n8844), .ZN(n7812) );
  AND2_X1 U8634 ( .A1(n7791), .A2(n7790), .ZN(n8844) );
  AND2_X1 U8635 ( .A1(n7788), .A2(n8845), .ZN(n8843) );
  OR2_X1 U8636 ( .A1(n7791), .A2(n7790), .ZN(n8845) );
  OR2_X1 U8637 ( .A1(n8846), .A2(n8847), .ZN(n7790) );
  AND2_X1 U8638 ( .A1(n7784), .A2(n7783), .ZN(n8847) );
  AND2_X1 U8639 ( .A1(n7781), .A2(n8848), .ZN(n8846) );
  OR2_X1 U8640 ( .A1(n7784), .A2(n7783), .ZN(n8848) );
  OR2_X1 U8641 ( .A1(n8849), .A2(n8850), .ZN(n7783) );
  AND2_X1 U8642 ( .A1(n7762), .A2(n7761), .ZN(n8850) );
  AND2_X1 U8643 ( .A1(n7759), .A2(n8851), .ZN(n8849) );
  OR2_X1 U8644 ( .A1(n7762), .A2(n7761), .ZN(n8851) );
  OR2_X1 U8645 ( .A1(n8852), .A2(n8853), .ZN(n7761) );
  AND2_X1 U8646 ( .A1(n7755), .A2(n7754), .ZN(n8853) );
  AND2_X1 U8647 ( .A1(n7752), .A2(n8854), .ZN(n8852) );
  OR2_X1 U8648 ( .A1(n7755), .A2(n7754), .ZN(n8854) );
  OR2_X1 U8649 ( .A1(n8855), .A2(n8856), .ZN(n7754) );
  AND2_X1 U8650 ( .A1(n7733), .A2(n7732), .ZN(n8856) );
  AND2_X1 U8651 ( .A1(n7730), .A2(n8857), .ZN(n8855) );
  OR2_X1 U8652 ( .A1(n7733), .A2(n7732), .ZN(n8857) );
  OR2_X1 U8653 ( .A1(n8858), .A2(n8859), .ZN(n7732) );
  AND2_X1 U8654 ( .A1(n7726), .A2(n7725), .ZN(n8859) );
  AND2_X1 U8655 ( .A1(n7723), .A2(n8860), .ZN(n8858) );
  OR2_X1 U8656 ( .A1(n7726), .A2(n7725), .ZN(n8860) );
  OR2_X1 U8657 ( .A1(n8861), .A2(n8862), .ZN(n7725) );
  AND2_X1 U8658 ( .A1(n7704), .A2(n7703), .ZN(n8862) );
  AND2_X1 U8659 ( .A1(n7701), .A2(n8863), .ZN(n8861) );
  OR2_X1 U8660 ( .A1(n7704), .A2(n7703), .ZN(n8863) );
  OR2_X1 U8661 ( .A1(n8864), .A2(n8865), .ZN(n7703) );
  AND2_X1 U8662 ( .A1(n7697), .A2(n7696), .ZN(n8865) );
  AND2_X1 U8663 ( .A1(n7694), .A2(n8866), .ZN(n8864) );
  OR2_X1 U8664 ( .A1(n7697), .A2(n7696), .ZN(n8866) );
  OR2_X1 U8665 ( .A1(n8867), .A2(n8868), .ZN(n7696) );
  AND2_X1 U8666 ( .A1(n7672), .A2(n7671), .ZN(n8868) );
  AND2_X1 U8667 ( .A1(n7669), .A2(n8869), .ZN(n8867) );
  OR2_X1 U8668 ( .A1(n7672), .A2(n7671), .ZN(n8869) );
  OR2_X1 U8669 ( .A1(n8870), .A2(n8871), .ZN(n7671) );
  AND2_X1 U8670 ( .A1(n7665), .A2(n7664), .ZN(n8871) );
  AND2_X1 U8671 ( .A1(n7662), .A2(n8872), .ZN(n8870) );
  OR2_X1 U8672 ( .A1(n7665), .A2(n7664), .ZN(n8872) );
  OR2_X1 U8673 ( .A1(n8873), .A2(n8874), .ZN(n7664) );
  AND2_X1 U8674 ( .A1(n7643), .A2(n7642), .ZN(n8874) );
  AND2_X1 U8675 ( .A1(n7640), .A2(n8875), .ZN(n8873) );
  OR2_X1 U8676 ( .A1(n7643), .A2(n7642), .ZN(n8875) );
  OR2_X1 U8677 ( .A1(n8876), .A2(n8877), .ZN(n7642) );
  AND2_X1 U8678 ( .A1(n7636), .A2(n7635), .ZN(n8877) );
  AND2_X1 U8679 ( .A1(n7633), .A2(n8878), .ZN(n8876) );
  OR2_X1 U8680 ( .A1(n7636), .A2(n7635), .ZN(n8878) );
  OR2_X1 U8681 ( .A1(n8879), .A2(n8880), .ZN(n7635) );
  AND2_X1 U8682 ( .A1(n7614), .A2(n7613), .ZN(n8880) );
  AND2_X1 U8683 ( .A1(n7611), .A2(n8881), .ZN(n8879) );
  OR2_X1 U8684 ( .A1(n7614), .A2(n7613), .ZN(n8881) );
  OR2_X1 U8685 ( .A1(n8882), .A2(n8883), .ZN(n7613) );
  AND2_X1 U8686 ( .A1(n7607), .A2(n7606), .ZN(n8883) );
  AND2_X1 U8687 ( .A1(n7604), .A2(n8884), .ZN(n8882) );
  OR2_X1 U8688 ( .A1(n7607), .A2(n7606), .ZN(n8884) );
  OR2_X1 U8689 ( .A1(n8885), .A2(n8886), .ZN(n7606) );
  AND2_X1 U8690 ( .A1(n7585), .A2(n7584), .ZN(n8886) );
  AND2_X1 U8691 ( .A1(n7582), .A2(n8887), .ZN(n8885) );
  OR2_X1 U8692 ( .A1(n7585), .A2(n7584), .ZN(n8887) );
  OR2_X1 U8693 ( .A1(n8888), .A2(n8889), .ZN(n7584) );
  AND2_X1 U8694 ( .A1(n7578), .A2(n7577), .ZN(n8889) );
  AND2_X1 U8695 ( .A1(n7575), .A2(n8890), .ZN(n8888) );
  OR2_X1 U8696 ( .A1(n7578), .A2(n7577), .ZN(n8890) );
  OR2_X1 U8697 ( .A1(n8891), .A2(n8892), .ZN(n7577) );
  AND2_X1 U8698 ( .A1(n7556), .A2(n7555), .ZN(n8892) );
  AND2_X1 U8699 ( .A1(n7553), .A2(n8893), .ZN(n8891) );
  OR2_X1 U8700 ( .A1(n7556), .A2(n7555), .ZN(n8893) );
  OR2_X1 U8701 ( .A1(n8894), .A2(n8895), .ZN(n7555) );
  AND2_X1 U8702 ( .A1(n7549), .A2(n7548), .ZN(n8895) );
  AND2_X1 U8703 ( .A1(n7546), .A2(n8896), .ZN(n8894) );
  OR2_X1 U8704 ( .A1(n7549), .A2(n7548), .ZN(n8896) );
  OR2_X1 U8705 ( .A1(n8897), .A2(n8898), .ZN(n7548) );
  AND2_X1 U8706 ( .A1(n7517), .A2(n7516), .ZN(n8898) );
  AND2_X1 U8707 ( .A1(n7514), .A2(n8899), .ZN(n8897) );
  OR2_X1 U8708 ( .A1(n7517), .A2(n7516), .ZN(n8899) );
  OR2_X1 U8709 ( .A1(n8900), .A2(n8901), .ZN(n7516) );
  AND2_X1 U8710 ( .A1(n7507), .A2(n7510), .ZN(n8901) );
  AND2_X1 U8711 ( .A1(n7509), .A2(n8902), .ZN(n8900) );
  OR2_X1 U8712 ( .A1(n7507), .A2(n7510), .ZN(n8902) );
  OR2_X1 U8713 ( .A1(n8051), .A2(n7479), .ZN(n7510) );
  INV_X1 U8714 ( .A(n8903), .ZN(n7507) );
  AND2_X1 U8715 ( .A1(b_30_), .A2(n8053), .ZN(n8903) );
  AND2_X1 U8716 ( .A1(n8904), .A2(b_31_), .ZN(n8053) );
  INV_X1 U8717 ( .A(n8905), .ZN(n7509) );
  OR2_X1 U8718 ( .A1(n8906), .A2(n8907), .ZN(n8905) );
  AND2_X1 U8719 ( .A1(b_30_), .A2(n8908), .ZN(n8907) );
  OR2_X1 U8720 ( .A1(n8909), .A2(n7490), .ZN(n8908) );
  AND2_X1 U8721 ( .A1(a_30_), .A2(n7501), .ZN(n8909) );
  AND2_X1 U8722 ( .A1(b_29_), .A2(n8910), .ZN(n8906) );
  OR2_X1 U8723 ( .A1(n8911), .A2(n7493), .ZN(n8910) );
  AND2_X1 U8724 ( .A1(a_31_), .A2(n7484), .ZN(n8911) );
  OR2_X1 U8725 ( .A1(n8048), .A2(n7479), .ZN(n7517) );
  XNOR2_X1 U8726 ( .A(n8912), .B(n8913), .ZN(n7514) );
  XNOR2_X1 U8727 ( .A(n8914), .B(n8915), .ZN(n8913) );
  OR2_X1 U8728 ( .A1(n8044), .A2(n7479), .ZN(n7549) );
  XOR2_X1 U8729 ( .A(n8916), .B(n8917), .Z(n7546) );
  XOR2_X1 U8730 ( .A(n8918), .B(n8919), .Z(n8917) );
  OR2_X1 U8731 ( .A1(n8041), .A2(n7479), .ZN(n7556) );
  XOR2_X1 U8732 ( .A(n8920), .B(n8921), .Z(n7553) );
  XOR2_X1 U8733 ( .A(n8922), .B(n8923), .Z(n8921) );
  OR2_X1 U8734 ( .A1(n8037), .A2(n7479), .ZN(n7578) );
  XOR2_X1 U8735 ( .A(n8924), .B(n8925), .Z(n7575) );
  XOR2_X1 U8736 ( .A(n8926), .B(n8927), .Z(n8925) );
  OR2_X1 U8737 ( .A1(n8034), .A2(n7479), .ZN(n7585) );
  XOR2_X1 U8738 ( .A(n8928), .B(n8929), .Z(n7582) );
  XOR2_X1 U8739 ( .A(n8930), .B(n8931), .Z(n8929) );
  OR2_X1 U8740 ( .A1(n8030), .A2(n7479), .ZN(n7607) );
  XOR2_X1 U8741 ( .A(n8932), .B(n8933), .Z(n7604) );
  XOR2_X1 U8742 ( .A(n8934), .B(n8935), .Z(n8933) );
  OR2_X1 U8743 ( .A1(n8026), .A2(n7479), .ZN(n7614) );
  XOR2_X1 U8744 ( .A(n8936), .B(n8937), .Z(n7611) );
  XOR2_X1 U8745 ( .A(n8938), .B(n8939), .Z(n8937) );
  OR2_X1 U8746 ( .A1(n8023), .A2(n7479), .ZN(n7636) );
  XOR2_X1 U8747 ( .A(n8940), .B(n8941), .Z(n7633) );
  XOR2_X1 U8748 ( .A(n8942), .B(n8943), .Z(n8941) );
  OR2_X1 U8749 ( .A1(n8019), .A2(n7479), .ZN(n7643) );
  XOR2_X1 U8750 ( .A(n8944), .B(n8945), .Z(n7640) );
  XOR2_X1 U8751 ( .A(n8946), .B(n8947), .Z(n8945) );
  OR2_X1 U8752 ( .A1(n8016), .A2(n7479), .ZN(n7665) );
  XOR2_X1 U8753 ( .A(n8948), .B(n8949), .Z(n7662) );
  XOR2_X1 U8754 ( .A(n8950), .B(n8951), .Z(n8949) );
  OR2_X1 U8755 ( .A1(n8012), .A2(n7479), .ZN(n7672) );
  XOR2_X1 U8756 ( .A(n8952), .B(n8953), .Z(n7669) );
  XOR2_X1 U8757 ( .A(n8954), .B(n8955), .Z(n8953) );
  OR2_X1 U8758 ( .A1(n8009), .A2(n7479), .ZN(n7697) );
  XOR2_X1 U8759 ( .A(n8956), .B(n8957), .Z(n7694) );
  XOR2_X1 U8760 ( .A(n8958), .B(n8959), .Z(n8957) );
  OR2_X1 U8761 ( .A1(n8005), .A2(n7479), .ZN(n7704) );
  XOR2_X1 U8762 ( .A(n8960), .B(n8961), .Z(n7701) );
  XOR2_X1 U8763 ( .A(n8962), .B(n8963), .Z(n8961) );
  OR2_X1 U8764 ( .A1(n8002), .A2(n7479), .ZN(n7726) );
  XOR2_X1 U8765 ( .A(n8964), .B(n8965), .Z(n7723) );
  XOR2_X1 U8766 ( .A(n8966), .B(n8967), .Z(n8965) );
  OR2_X1 U8767 ( .A1(n7998), .A2(n7479), .ZN(n7733) );
  XOR2_X1 U8768 ( .A(n8968), .B(n8969), .Z(n7730) );
  XOR2_X1 U8769 ( .A(n8970), .B(n8971), .Z(n8969) );
  OR2_X1 U8770 ( .A1(n7995), .A2(n7479), .ZN(n7755) );
  XOR2_X1 U8771 ( .A(n8972), .B(n8973), .Z(n7752) );
  XOR2_X1 U8772 ( .A(n8974), .B(n8975), .Z(n8973) );
  OR2_X1 U8773 ( .A1(n7991), .A2(n7479), .ZN(n7762) );
  XOR2_X1 U8774 ( .A(n8976), .B(n8977), .Z(n7759) );
  XOR2_X1 U8775 ( .A(n8978), .B(n8979), .Z(n8977) );
  OR2_X1 U8776 ( .A1(n7988), .A2(n7479), .ZN(n7784) );
  XOR2_X1 U8777 ( .A(n8980), .B(n8981), .Z(n7781) );
  XOR2_X1 U8778 ( .A(n8982), .B(n8983), .Z(n8981) );
  OR2_X1 U8779 ( .A1(n7984), .A2(n7479), .ZN(n7791) );
  XOR2_X1 U8780 ( .A(n8984), .B(n8985), .Z(n7788) );
  XOR2_X1 U8781 ( .A(n8986), .B(n8987), .Z(n8985) );
  OR2_X1 U8782 ( .A1(n7981), .A2(n7479), .ZN(n7813) );
  XOR2_X1 U8783 ( .A(n8988), .B(n8989), .Z(n7810) );
  XOR2_X1 U8784 ( .A(n8990), .B(n8991), .Z(n8989) );
  OR2_X1 U8785 ( .A1(n7977), .A2(n7479), .ZN(n7820) );
  XOR2_X1 U8786 ( .A(n8992), .B(n8993), .Z(n7817) );
  XOR2_X1 U8787 ( .A(n8994), .B(n8995), .Z(n8993) );
  OR2_X1 U8788 ( .A1(n7974), .A2(n7479), .ZN(n7852) );
  XOR2_X1 U8789 ( .A(n8996), .B(n8997), .Z(n7849) );
  XOR2_X1 U8790 ( .A(n8998), .B(n8999), .Z(n8997) );
  OR2_X1 U8791 ( .A1(n7970), .A2(n7479), .ZN(n7859) );
  XOR2_X1 U8792 ( .A(n9000), .B(n9001), .Z(n7856) );
  XOR2_X1 U8793 ( .A(n9002), .B(n9003), .Z(n9001) );
  OR2_X1 U8794 ( .A1(n7967), .A2(n7479), .ZN(n7881) );
  XOR2_X1 U8795 ( .A(n9004), .B(n9005), .Z(n7878) );
  XOR2_X1 U8796 ( .A(n9006), .B(n9007), .Z(n9005) );
  OR2_X1 U8797 ( .A1(n7963), .A2(n7479), .ZN(n7888) );
  XOR2_X1 U8798 ( .A(n9008), .B(n9009), .Z(n7885) );
  XOR2_X1 U8799 ( .A(n9010), .B(n9011), .Z(n9009) );
  OR2_X1 U8800 ( .A1(n7960), .A2(n7479), .ZN(n7910) );
  XOR2_X1 U8801 ( .A(n9012), .B(n9013), .Z(n7907) );
  XOR2_X1 U8802 ( .A(n9014), .B(n9015), .Z(n9013) );
  OR2_X1 U8803 ( .A1(n7956), .A2(n7479), .ZN(n7917) );
  XOR2_X1 U8804 ( .A(n9016), .B(n9017), .Z(n7914) );
  XOR2_X1 U8805 ( .A(n9018), .B(n9019), .Z(n9017) );
  OR2_X1 U8806 ( .A1(n7953), .A2(n7479), .ZN(n7939) );
  XOR2_X1 U8807 ( .A(n9020), .B(n9021), .Z(n7936) );
  XOR2_X1 U8808 ( .A(n9022), .B(n9023), .Z(n9021) );
  OR2_X1 U8809 ( .A1(n7950), .A2(n7479), .ZN(n7946) );
  INV_X1 U8810 ( .A(b_31_), .ZN(n7479) );
  XOR2_X1 U8811 ( .A(n9024), .B(n9025), .Z(n7943) );
  XOR2_X1 U8812 ( .A(n9026), .B(n9027), .Z(n9025) );
  XOR2_X1 U8813 ( .A(n8807), .B(n8808), .Z(n8062) );
  OR2_X1 U8814 ( .A1(n9028), .A2(n9029), .ZN(n8808) );
  AND2_X1 U8815 ( .A1(n9030), .A2(n9031), .ZN(n9029) );
  AND2_X1 U8816 ( .A1(n9032), .A2(n9033), .ZN(n9028) );
  OR2_X1 U8817 ( .A1(n9030), .A2(n9031), .ZN(n9033) );
  XOR2_X1 U8818 ( .A(n9034), .B(n9035), .Z(n8807) );
  XOR2_X1 U8819 ( .A(n9036), .B(n9037), .Z(n9035) );
  XNOR2_X1 U8820 ( .A(n9032), .B(n9038), .ZN(n8058) );
  XOR2_X1 U8821 ( .A(n9031), .B(n9030), .Z(n9038) );
  OR2_X1 U8822 ( .A1(n7950), .A2(n7484), .ZN(n9030) );
  OR2_X1 U8823 ( .A1(n9039), .A2(n9040), .ZN(n9031) );
  AND2_X1 U8824 ( .A1(n9024), .A2(n9027), .ZN(n9040) );
  AND2_X1 U8825 ( .A1(n9041), .A2(n9026), .ZN(n9039) );
  OR2_X1 U8826 ( .A1(n9042), .A2(n9043), .ZN(n9026) );
  AND2_X1 U8827 ( .A1(n9020), .A2(n9023), .ZN(n9043) );
  AND2_X1 U8828 ( .A1(n9044), .A2(n9022), .ZN(n9042) );
  OR2_X1 U8829 ( .A1(n9045), .A2(n9046), .ZN(n9022) );
  AND2_X1 U8830 ( .A1(n9016), .A2(n9019), .ZN(n9046) );
  AND2_X1 U8831 ( .A1(n9047), .A2(n9018), .ZN(n9045) );
  OR2_X1 U8832 ( .A1(n9048), .A2(n9049), .ZN(n9018) );
  AND2_X1 U8833 ( .A1(n9012), .A2(n9015), .ZN(n9049) );
  AND2_X1 U8834 ( .A1(n9050), .A2(n9014), .ZN(n9048) );
  OR2_X1 U8835 ( .A1(n9051), .A2(n9052), .ZN(n9014) );
  AND2_X1 U8836 ( .A1(n9008), .A2(n9011), .ZN(n9052) );
  AND2_X1 U8837 ( .A1(n9053), .A2(n9010), .ZN(n9051) );
  OR2_X1 U8838 ( .A1(n9054), .A2(n9055), .ZN(n9010) );
  AND2_X1 U8839 ( .A1(n9004), .A2(n9007), .ZN(n9055) );
  AND2_X1 U8840 ( .A1(n9056), .A2(n9006), .ZN(n9054) );
  OR2_X1 U8841 ( .A1(n9057), .A2(n9058), .ZN(n9006) );
  AND2_X1 U8842 ( .A1(n9000), .A2(n9003), .ZN(n9058) );
  AND2_X1 U8843 ( .A1(n9059), .A2(n9002), .ZN(n9057) );
  OR2_X1 U8844 ( .A1(n9060), .A2(n9061), .ZN(n9002) );
  AND2_X1 U8845 ( .A1(n8996), .A2(n8999), .ZN(n9061) );
  AND2_X1 U8846 ( .A1(n9062), .A2(n8998), .ZN(n9060) );
  OR2_X1 U8847 ( .A1(n9063), .A2(n9064), .ZN(n8998) );
  AND2_X1 U8848 ( .A1(n8992), .A2(n8995), .ZN(n9064) );
  AND2_X1 U8849 ( .A1(n9065), .A2(n8994), .ZN(n9063) );
  OR2_X1 U8850 ( .A1(n9066), .A2(n9067), .ZN(n8994) );
  AND2_X1 U8851 ( .A1(n8988), .A2(n8991), .ZN(n9067) );
  AND2_X1 U8852 ( .A1(n9068), .A2(n8990), .ZN(n9066) );
  OR2_X1 U8853 ( .A1(n9069), .A2(n9070), .ZN(n8990) );
  AND2_X1 U8854 ( .A1(n8984), .A2(n8987), .ZN(n9070) );
  AND2_X1 U8855 ( .A1(n9071), .A2(n8986), .ZN(n9069) );
  OR2_X1 U8856 ( .A1(n9072), .A2(n9073), .ZN(n8986) );
  AND2_X1 U8857 ( .A1(n8980), .A2(n8983), .ZN(n9073) );
  AND2_X1 U8858 ( .A1(n9074), .A2(n8982), .ZN(n9072) );
  OR2_X1 U8859 ( .A1(n9075), .A2(n9076), .ZN(n8982) );
  AND2_X1 U8860 ( .A1(n8976), .A2(n8979), .ZN(n9076) );
  AND2_X1 U8861 ( .A1(n9077), .A2(n8978), .ZN(n9075) );
  OR2_X1 U8862 ( .A1(n9078), .A2(n9079), .ZN(n8978) );
  AND2_X1 U8863 ( .A1(n8972), .A2(n8975), .ZN(n9079) );
  AND2_X1 U8864 ( .A1(n9080), .A2(n8974), .ZN(n9078) );
  OR2_X1 U8865 ( .A1(n9081), .A2(n9082), .ZN(n8974) );
  AND2_X1 U8866 ( .A1(n8968), .A2(n8971), .ZN(n9082) );
  AND2_X1 U8867 ( .A1(n9083), .A2(n8970), .ZN(n9081) );
  OR2_X1 U8868 ( .A1(n9084), .A2(n9085), .ZN(n8970) );
  AND2_X1 U8869 ( .A1(n8964), .A2(n8967), .ZN(n9085) );
  AND2_X1 U8870 ( .A1(n9086), .A2(n8966), .ZN(n9084) );
  OR2_X1 U8871 ( .A1(n9087), .A2(n9088), .ZN(n8966) );
  AND2_X1 U8872 ( .A1(n8960), .A2(n8963), .ZN(n9088) );
  AND2_X1 U8873 ( .A1(n9089), .A2(n8962), .ZN(n9087) );
  OR2_X1 U8874 ( .A1(n9090), .A2(n9091), .ZN(n8962) );
  AND2_X1 U8875 ( .A1(n8956), .A2(n8959), .ZN(n9091) );
  AND2_X1 U8876 ( .A1(n9092), .A2(n8958), .ZN(n9090) );
  OR2_X1 U8877 ( .A1(n9093), .A2(n9094), .ZN(n8958) );
  AND2_X1 U8878 ( .A1(n8952), .A2(n8955), .ZN(n9094) );
  AND2_X1 U8879 ( .A1(n9095), .A2(n8954), .ZN(n9093) );
  OR2_X1 U8880 ( .A1(n9096), .A2(n9097), .ZN(n8954) );
  AND2_X1 U8881 ( .A1(n8948), .A2(n8951), .ZN(n9097) );
  AND2_X1 U8882 ( .A1(n9098), .A2(n8950), .ZN(n9096) );
  OR2_X1 U8883 ( .A1(n9099), .A2(n9100), .ZN(n8950) );
  AND2_X1 U8884 ( .A1(n8944), .A2(n8947), .ZN(n9100) );
  AND2_X1 U8885 ( .A1(n9101), .A2(n8946), .ZN(n9099) );
  OR2_X1 U8886 ( .A1(n9102), .A2(n9103), .ZN(n8946) );
  AND2_X1 U8887 ( .A1(n8940), .A2(n8943), .ZN(n9103) );
  AND2_X1 U8888 ( .A1(n9104), .A2(n8942), .ZN(n9102) );
  OR2_X1 U8889 ( .A1(n9105), .A2(n9106), .ZN(n8942) );
  AND2_X1 U8890 ( .A1(n8936), .A2(n8939), .ZN(n9106) );
  AND2_X1 U8891 ( .A1(n9107), .A2(n8938), .ZN(n9105) );
  OR2_X1 U8892 ( .A1(n9108), .A2(n9109), .ZN(n8938) );
  AND2_X1 U8893 ( .A1(n8932), .A2(n8935), .ZN(n9109) );
  AND2_X1 U8894 ( .A1(n9110), .A2(n8934), .ZN(n9108) );
  OR2_X1 U8895 ( .A1(n9111), .A2(n9112), .ZN(n8934) );
  AND2_X1 U8896 ( .A1(n8928), .A2(n8931), .ZN(n9112) );
  AND2_X1 U8897 ( .A1(n9113), .A2(n8930), .ZN(n9111) );
  OR2_X1 U8898 ( .A1(n9114), .A2(n9115), .ZN(n8930) );
  AND2_X1 U8899 ( .A1(n8924), .A2(n8927), .ZN(n9115) );
  AND2_X1 U8900 ( .A1(n9116), .A2(n8926), .ZN(n9114) );
  OR2_X1 U8901 ( .A1(n9117), .A2(n9118), .ZN(n8926) );
  AND2_X1 U8902 ( .A1(n8920), .A2(n8923), .ZN(n9118) );
  AND2_X1 U8903 ( .A1(n9119), .A2(n8922), .ZN(n9117) );
  OR2_X1 U8904 ( .A1(n9120), .A2(n9121), .ZN(n8922) );
  AND2_X1 U8905 ( .A1(n8916), .A2(n8919), .ZN(n9121) );
  AND2_X1 U8906 ( .A1(n9122), .A2(n8918), .ZN(n9120) );
  OR2_X1 U8907 ( .A1(n9123), .A2(n9124), .ZN(n8918) );
  AND2_X1 U8908 ( .A1(n8912), .A2(n9125), .ZN(n9124) );
  AND2_X1 U8909 ( .A1(n9126), .A2(n9127), .ZN(n9123) );
  OR2_X1 U8910 ( .A1(n9125), .A2(n8912), .ZN(n9127) );
  OR2_X1 U8911 ( .A1(n8051), .A2(n7484), .ZN(n8912) );
  INV_X1 U8912 ( .A(n8915), .ZN(n9125) );
  AND3_X1 U8913 ( .A1(n8904), .A2(b_29_), .A3(b_30_), .ZN(n8915) );
  INV_X1 U8914 ( .A(n8914), .ZN(n9126) );
  OR2_X1 U8915 ( .A1(n9128), .A2(n9129), .ZN(n8914) );
  AND2_X1 U8916 ( .A1(b_29_), .A2(n9130), .ZN(n9129) );
  OR2_X1 U8917 ( .A1(n9131), .A2(n7490), .ZN(n9130) );
  AND2_X1 U8918 ( .A1(a_30_), .A2(n8049), .ZN(n9131) );
  AND2_X1 U8919 ( .A1(b_28_), .A2(n9132), .ZN(n9128) );
  OR2_X1 U8920 ( .A1(n9133), .A2(n7493), .ZN(n9132) );
  AND2_X1 U8921 ( .A1(a_31_), .A2(n7501), .ZN(n9133) );
  OR2_X1 U8922 ( .A1(n8919), .A2(n8916), .ZN(n9122) );
  XOR2_X1 U8923 ( .A(n7505), .B(n9134), .Z(n8916) );
  XNOR2_X1 U8924 ( .A(n9135), .B(n9136), .ZN(n9134) );
  OR2_X1 U8925 ( .A1(n8048), .A2(n7484), .ZN(n8919) );
  OR2_X1 U8926 ( .A1(n8923), .A2(n8920), .ZN(n9119) );
  XOR2_X1 U8927 ( .A(n9137), .B(n9138), .Z(n8920) );
  XOR2_X1 U8928 ( .A(n9139), .B(n9140), .Z(n9138) );
  OR2_X1 U8929 ( .A1(n8044), .A2(n7484), .ZN(n8923) );
  OR2_X1 U8930 ( .A1(n8927), .A2(n8924), .ZN(n9116) );
  XOR2_X1 U8931 ( .A(n9141), .B(n9142), .Z(n8924) );
  XOR2_X1 U8932 ( .A(n9143), .B(n9144), .Z(n9142) );
  OR2_X1 U8933 ( .A1(n8041), .A2(n7484), .ZN(n8927) );
  OR2_X1 U8934 ( .A1(n8931), .A2(n8928), .ZN(n9113) );
  XOR2_X1 U8935 ( .A(n9145), .B(n9146), .Z(n8928) );
  XOR2_X1 U8936 ( .A(n9147), .B(n9148), .Z(n9146) );
  OR2_X1 U8937 ( .A1(n8037), .A2(n7484), .ZN(n8931) );
  OR2_X1 U8938 ( .A1(n8935), .A2(n8932), .ZN(n9110) );
  XOR2_X1 U8939 ( .A(n9149), .B(n9150), .Z(n8932) );
  XOR2_X1 U8940 ( .A(n9151), .B(n9152), .Z(n9150) );
  OR2_X1 U8941 ( .A1(n8034), .A2(n7484), .ZN(n8935) );
  OR2_X1 U8942 ( .A1(n8939), .A2(n8936), .ZN(n9107) );
  XOR2_X1 U8943 ( .A(n9153), .B(n9154), .Z(n8936) );
  XOR2_X1 U8944 ( .A(n9155), .B(n9156), .Z(n9154) );
  OR2_X1 U8945 ( .A1(n8030), .A2(n7484), .ZN(n8939) );
  OR2_X1 U8946 ( .A1(n8943), .A2(n8940), .ZN(n9104) );
  XOR2_X1 U8947 ( .A(n9157), .B(n9158), .Z(n8940) );
  XOR2_X1 U8948 ( .A(n9159), .B(n9160), .Z(n9158) );
  OR2_X1 U8949 ( .A1(n8026), .A2(n7484), .ZN(n8943) );
  OR2_X1 U8950 ( .A1(n8947), .A2(n8944), .ZN(n9101) );
  XOR2_X1 U8951 ( .A(n9161), .B(n9162), .Z(n8944) );
  XOR2_X1 U8952 ( .A(n9163), .B(n9164), .Z(n9162) );
  OR2_X1 U8953 ( .A1(n8023), .A2(n7484), .ZN(n8947) );
  OR2_X1 U8954 ( .A1(n8951), .A2(n8948), .ZN(n9098) );
  XOR2_X1 U8955 ( .A(n9165), .B(n9166), .Z(n8948) );
  XOR2_X1 U8956 ( .A(n9167), .B(n9168), .Z(n9166) );
  OR2_X1 U8957 ( .A1(n8019), .A2(n7484), .ZN(n8951) );
  OR2_X1 U8958 ( .A1(n8955), .A2(n8952), .ZN(n9095) );
  XOR2_X1 U8959 ( .A(n9169), .B(n9170), .Z(n8952) );
  XOR2_X1 U8960 ( .A(n9171), .B(n9172), .Z(n9170) );
  OR2_X1 U8961 ( .A1(n8016), .A2(n7484), .ZN(n8955) );
  OR2_X1 U8962 ( .A1(n8959), .A2(n8956), .ZN(n9092) );
  XOR2_X1 U8963 ( .A(n9173), .B(n9174), .Z(n8956) );
  XOR2_X1 U8964 ( .A(n9175), .B(n9176), .Z(n9174) );
  OR2_X1 U8965 ( .A1(n8012), .A2(n7484), .ZN(n8959) );
  OR2_X1 U8966 ( .A1(n8963), .A2(n8960), .ZN(n9089) );
  XOR2_X1 U8967 ( .A(n9177), .B(n9178), .Z(n8960) );
  XOR2_X1 U8968 ( .A(n9179), .B(n9180), .Z(n9178) );
  OR2_X1 U8969 ( .A1(n8009), .A2(n7484), .ZN(n8963) );
  OR2_X1 U8970 ( .A1(n8967), .A2(n8964), .ZN(n9086) );
  XOR2_X1 U8971 ( .A(n9181), .B(n9182), .Z(n8964) );
  XOR2_X1 U8972 ( .A(n9183), .B(n9184), .Z(n9182) );
  OR2_X1 U8973 ( .A1(n8005), .A2(n7484), .ZN(n8967) );
  OR2_X1 U8974 ( .A1(n8971), .A2(n8968), .ZN(n9083) );
  XOR2_X1 U8975 ( .A(n9185), .B(n9186), .Z(n8968) );
  XOR2_X1 U8976 ( .A(n9187), .B(n9188), .Z(n9186) );
  OR2_X1 U8977 ( .A1(n8002), .A2(n7484), .ZN(n8971) );
  OR2_X1 U8978 ( .A1(n8975), .A2(n8972), .ZN(n9080) );
  XOR2_X1 U8979 ( .A(n9189), .B(n9190), .Z(n8972) );
  XOR2_X1 U8980 ( .A(n9191), .B(n9192), .Z(n9190) );
  OR2_X1 U8981 ( .A1(n7998), .A2(n7484), .ZN(n8975) );
  OR2_X1 U8982 ( .A1(n8979), .A2(n8976), .ZN(n9077) );
  XOR2_X1 U8983 ( .A(n9193), .B(n9194), .Z(n8976) );
  XOR2_X1 U8984 ( .A(n9195), .B(n9196), .Z(n9194) );
  OR2_X1 U8985 ( .A1(n7995), .A2(n7484), .ZN(n8979) );
  OR2_X1 U8986 ( .A1(n8983), .A2(n8980), .ZN(n9074) );
  XOR2_X1 U8987 ( .A(n9197), .B(n9198), .Z(n8980) );
  XOR2_X1 U8988 ( .A(n9199), .B(n9200), .Z(n9198) );
  OR2_X1 U8989 ( .A1(n7991), .A2(n7484), .ZN(n8983) );
  OR2_X1 U8990 ( .A1(n8987), .A2(n8984), .ZN(n9071) );
  XOR2_X1 U8991 ( .A(n9201), .B(n9202), .Z(n8984) );
  XOR2_X1 U8992 ( .A(n9203), .B(n9204), .Z(n9202) );
  OR2_X1 U8993 ( .A1(n7988), .A2(n7484), .ZN(n8987) );
  OR2_X1 U8994 ( .A1(n8991), .A2(n8988), .ZN(n9068) );
  XOR2_X1 U8995 ( .A(n9205), .B(n9206), .Z(n8988) );
  XOR2_X1 U8996 ( .A(n9207), .B(n9208), .Z(n9206) );
  OR2_X1 U8997 ( .A1(n7984), .A2(n7484), .ZN(n8991) );
  OR2_X1 U8998 ( .A1(n8995), .A2(n8992), .ZN(n9065) );
  XOR2_X1 U8999 ( .A(n9209), .B(n9210), .Z(n8992) );
  XOR2_X1 U9000 ( .A(n9211), .B(n9212), .Z(n9210) );
  OR2_X1 U9001 ( .A1(n7981), .A2(n7484), .ZN(n8995) );
  OR2_X1 U9002 ( .A1(n8999), .A2(n8996), .ZN(n9062) );
  XOR2_X1 U9003 ( .A(n9213), .B(n9214), .Z(n8996) );
  XOR2_X1 U9004 ( .A(n9215), .B(n9216), .Z(n9214) );
  OR2_X1 U9005 ( .A1(n7977), .A2(n7484), .ZN(n8999) );
  OR2_X1 U9006 ( .A1(n9003), .A2(n9000), .ZN(n9059) );
  XOR2_X1 U9007 ( .A(n9217), .B(n9218), .Z(n9000) );
  XOR2_X1 U9008 ( .A(n9219), .B(n9220), .Z(n9218) );
  OR2_X1 U9009 ( .A1(n7974), .A2(n7484), .ZN(n9003) );
  OR2_X1 U9010 ( .A1(n9007), .A2(n9004), .ZN(n9056) );
  XOR2_X1 U9011 ( .A(n9221), .B(n9222), .Z(n9004) );
  XOR2_X1 U9012 ( .A(n9223), .B(n9224), .Z(n9222) );
  OR2_X1 U9013 ( .A1(n7970), .A2(n7484), .ZN(n9007) );
  OR2_X1 U9014 ( .A1(n9011), .A2(n9008), .ZN(n9053) );
  XOR2_X1 U9015 ( .A(n9225), .B(n9226), .Z(n9008) );
  XOR2_X1 U9016 ( .A(n9227), .B(n9228), .Z(n9226) );
  OR2_X1 U9017 ( .A1(n7967), .A2(n7484), .ZN(n9011) );
  OR2_X1 U9018 ( .A1(n9015), .A2(n9012), .ZN(n9050) );
  XOR2_X1 U9019 ( .A(n9229), .B(n9230), .Z(n9012) );
  XOR2_X1 U9020 ( .A(n9231), .B(n9232), .Z(n9230) );
  OR2_X1 U9021 ( .A1(n7963), .A2(n7484), .ZN(n9015) );
  OR2_X1 U9022 ( .A1(n9019), .A2(n9016), .ZN(n9047) );
  XOR2_X1 U9023 ( .A(n9233), .B(n9234), .Z(n9016) );
  XOR2_X1 U9024 ( .A(n9235), .B(n9236), .Z(n9234) );
  OR2_X1 U9025 ( .A1(n7960), .A2(n7484), .ZN(n9019) );
  OR2_X1 U9026 ( .A1(n9023), .A2(n9020), .ZN(n9044) );
  XOR2_X1 U9027 ( .A(n9237), .B(n9238), .Z(n9020) );
  XOR2_X1 U9028 ( .A(n9239), .B(n9240), .Z(n9238) );
  OR2_X1 U9029 ( .A1(n7956), .A2(n7484), .ZN(n9023) );
  OR2_X1 U9030 ( .A1(n9027), .A2(n9024), .ZN(n9041) );
  XNOR2_X1 U9031 ( .A(n9241), .B(n9242), .ZN(n9024) );
  XNOR2_X1 U9032 ( .A(n9243), .B(n9244), .ZN(n9241) );
  OR2_X1 U9033 ( .A1(n7953), .A2(n7484), .ZN(n9027) );
  INV_X1 U9034 ( .A(b_30_), .ZN(n7484) );
  XOR2_X1 U9035 ( .A(n9245), .B(n9246), .Z(n9032) );
  XOR2_X1 U9036 ( .A(n9247), .B(n9248), .Z(n9246) );
  OR2_X1 U9037 ( .A1(n9249), .A2(n8802), .ZN(n8075) );
  XNOR2_X1 U9038 ( .A(n8797), .B(n9250), .ZN(n8802) );
  AND2_X1 U9039 ( .A1(n8803), .A2(n8801), .ZN(n9249) );
  XNOR2_X1 U9040 ( .A(n9251), .B(n9252), .ZN(n8801) );
  XOR2_X1 U9041 ( .A(n9253), .B(n9254), .Z(n9252) );
  INV_X1 U9042 ( .A(n8811), .ZN(n8803) );
  OR2_X1 U9043 ( .A1(n9255), .A2(n9256), .ZN(n8811) );
  AND2_X1 U9044 ( .A1(n9037), .A2(n9036), .ZN(n9256) );
  AND2_X1 U9045 ( .A1(n9034), .A2(n9257), .ZN(n9255) );
  OR2_X1 U9046 ( .A1(n9036), .A2(n9037), .ZN(n9257) );
  OR2_X1 U9047 ( .A1(n7950), .A2(n7501), .ZN(n9037) );
  OR2_X1 U9048 ( .A1(n9258), .A2(n9259), .ZN(n9036) );
  AND2_X1 U9049 ( .A1(n9248), .A2(n9247), .ZN(n9259) );
  AND2_X1 U9050 ( .A1(n9245), .A2(n9260), .ZN(n9258) );
  OR2_X1 U9051 ( .A1(n9247), .A2(n9248), .ZN(n9260) );
  OR2_X1 U9052 ( .A1(n7953), .A2(n7501), .ZN(n9248) );
  OR2_X1 U9053 ( .A1(n9261), .A2(n9262), .ZN(n9247) );
  AND2_X1 U9054 ( .A1(n9244), .A2(n9243), .ZN(n9262) );
  AND2_X1 U9055 ( .A1(n9242), .A2(n9263), .ZN(n9261) );
  OR2_X1 U9056 ( .A1(n9243), .A2(n9244), .ZN(n9263) );
  OR2_X1 U9057 ( .A1(n9264), .A2(n9265), .ZN(n9244) );
  AND2_X1 U9058 ( .A1(n9240), .A2(n9239), .ZN(n9265) );
  AND2_X1 U9059 ( .A1(n9237), .A2(n9266), .ZN(n9264) );
  OR2_X1 U9060 ( .A1(n9239), .A2(n9240), .ZN(n9266) );
  OR2_X1 U9061 ( .A1(n7960), .A2(n7501), .ZN(n9240) );
  OR2_X1 U9062 ( .A1(n9267), .A2(n9268), .ZN(n9239) );
  AND2_X1 U9063 ( .A1(n9236), .A2(n9235), .ZN(n9268) );
  AND2_X1 U9064 ( .A1(n9233), .A2(n9269), .ZN(n9267) );
  OR2_X1 U9065 ( .A1(n9235), .A2(n9236), .ZN(n9269) );
  OR2_X1 U9066 ( .A1(n7963), .A2(n7501), .ZN(n9236) );
  OR2_X1 U9067 ( .A1(n9270), .A2(n9271), .ZN(n9235) );
  AND2_X1 U9068 ( .A1(n9232), .A2(n9231), .ZN(n9271) );
  AND2_X1 U9069 ( .A1(n9229), .A2(n9272), .ZN(n9270) );
  OR2_X1 U9070 ( .A1(n9231), .A2(n9232), .ZN(n9272) );
  OR2_X1 U9071 ( .A1(n7967), .A2(n7501), .ZN(n9232) );
  OR2_X1 U9072 ( .A1(n9273), .A2(n9274), .ZN(n9231) );
  AND2_X1 U9073 ( .A1(n9228), .A2(n9227), .ZN(n9274) );
  AND2_X1 U9074 ( .A1(n9225), .A2(n9275), .ZN(n9273) );
  OR2_X1 U9075 ( .A1(n9227), .A2(n9228), .ZN(n9275) );
  OR2_X1 U9076 ( .A1(n7970), .A2(n7501), .ZN(n9228) );
  OR2_X1 U9077 ( .A1(n9276), .A2(n9277), .ZN(n9227) );
  AND2_X1 U9078 ( .A1(n9224), .A2(n9223), .ZN(n9277) );
  AND2_X1 U9079 ( .A1(n9221), .A2(n9278), .ZN(n9276) );
  OR2_X1 U9080 ( .A1(n9223), .A2(n9224), .ZN(n9278) );
  OR2_X1 U9081 ( .A1(n7974), .A2(n7501), .ZN(n9224) );
  OR2_X1 U9082 ( .A1(n9279), .A2(n9280), .ZN(n9223) );
  AND2_X1 U9083 ( .A1(n9220), .A2(n9219), .ZN(n9280) );
  AND2_X1 U9084 ( .A1(n9217), .A2(n9281), .ZN(n9279) );
  OR2_X1 U9085 ( .A1(n9219), .A2(n9220), .ZN(n9281) );
  OR2_X1 U9086 ( .A1(n7977), .A2(n7501), .ZN(n9220) );
  OR2_X1 U9087 ( .A1(n9282), .A2(n9283), .ZN(n9219) );
  AND2_X1 U9088 ( .A1(n9216), .A2(n9215), .ZN(n9283) );
  AND2_X1 U9089 ( .A1(n9213), .A2(n9284), .ZN(n9282) );
  OR2_X1 U9090 ( .A1(n9215), .A2(n9216), .ZN(n9284) );
  OR2_X1 U9091 ( .A1(n7981), .A2(n7501), .ZN(n9216) );
  OR2_X1 U9092 ( .A1(n9285), .A2(n9286), .ZN(n9215) );
  AND2_X1 U9093 ( .A1(n9212), .A2(n9211), .ZN(n9286) );
  AND2_X1 U9094 ( .A1(n9209), .A2(n9287), .ZN(n9285) );
  OR2_X1 U9095 ( .A1(n9211), .A2(n9212), .ZN(n9287) );
  OR2_X1 U9096 ( .A1(n7984), .A2(n7501), .ZN(n9212) );
  OR2_X1 U9097 ( .A1(n9288), .A2(n9289), .ZN(n9211) );
  AND2_X1 U9098 ( .A1(n9208), .A2(n9207), .ZN(n9289) );
  AND2_X1 U9099 ( .A1(n9205), .A2(n9290), .ZN(n9288) );
  OR2_X1 U9100 ( .A1(n9207), .A2(n9208), .ZN(n9290) );
  OR2_X1 U9101 ( .A1(n7988), .A2(n7501), .ZN(n9208) );
  OR2_X1 U9102 ( .A1(n9291), .A2(n9292), .ZN(n9207) );
  AND2_X1 U9103 ( .A1(n9204), .A2(n9203), .ZN(n9292) );
  AND2_X1 U9104 ( .A1(n9201), .A2(n9293), .ZN(n9291) );
  OR2_X1 U9105 ( .A1(n9203), .A2(n9204), .ZN(n9293) );
  OR2_X1 U9106 ( .A1(n7991), .A2(n7501), .ZN(n9204) );
  OR2_X1 U9107 ( .A1(n9294), .A2(n9295), .ZN(n9203) );
  AND2_X1 U9108 ( .A1(n9200), .A2(n9199), .ZN(n9295) );
  AND2_X1 U9109 ( .A1(n9197), .A2(n9296), .ZN(n9294) );
  OR2_X1 U9110 ( .A1(n9199), .A2(n9200), .ZN(n9296) );
  OR2_X1 U9111 ( .A1(n7995), .A2(n7501), .ZN(n9200) );
  OR2_X1 U9112 ( .A1(n9297), .A2(n9298), .ZN(n9199) );
  AND2_X1 U9113 ( .A1(n9196), .A2(n9195), .ZN(n9298) );
  AND2_X1 U9114 ( .A1(n9193), .A2(n9299), .ZN(n9297) );
  OR2_X1 U9115 ( .A1(n9195), .A2(n9196), .ZN(n9299) );
  OR2_X1 U9116 ( .A1(n7998), .A2(n7501), .ZN(n9196) );
  OR2_X1 U9117 ( .A1(n9300), .A2(n9301), .ZN(n9195) );
  AND2_X1 U9118 ( .A1(n9192), .A2(n9191), .ZN(n9301) );
  AND2_X1 U9119 ( .A1(n9189), .A2(n9302), .ZN(n9300) );
  OR2_X1 U9120 ( .A1(n9191), .A2(n9192), .ZN(n9302) );
  OR2_X1 U9121 ( .A1(n8002), .A2(n7501), .ZN(n9192) );
  OR2_X1 U9122 ( .A1(n9303), .A2(n9304), .ZN(n9191) );
  AND2_X1 U9123 ( .A1(n9188), .A2(n9187), .ZN(n9304) );
  AND2_X1 U9124 ( .A1(n9185), .A2(n9305), .ZN(n9303) );
  OR2_X1 U9125 ( .A1(n9187), .A2(n9188), .ZN(n9305) );
  OR2_X1 U9126 ( .A1(n8005), .A2(n7501), .ZN(n9188) );
  OR2_X1 U9127 ( .A1(n9306), .A2(n9307), .ZN(n9187) );
  AND2_X1 U9128 ( .A1(n9184), .A2(n9183), .ZN(n9307) );
  AND2_X1 U9129 ( .A1(n9181), .A2(n9308), .ZN(n9306) );
  OR2_X1 U9130 ( .A1(n9183), .A2(n9184), .ZN(n9308) );
  OR2_X1 U9131 ( .A1(n8009), .A2(n7501), .ZN(n9184) );
  OR2_X1 U9132 ( .A1(n9309), .A2(n9310), .ZN(n9183) );
  AND2_X1 U9133 ( .A1(n9180), .A2(n9179), .ZN(n9310) );
  AND2_X1 U9134 ( .A1(n9177), .A2(n9311), .ZN(n9309) );
  OR2_X1 U9135 ( .A1(n9179), .A2(n9180), .ZN(n9311) );
  OR2_X1 U9136 ( .A1(n8012), .A2(n7501), .ZN(n9180) );
  OR2_X1 U9137 ( .A1(n9312), .A2(n9313), .ZN(n9179) );
  AND2_X1 U9138 ( .A1(n9176), .A2(n9175), .ZN(n9313) );
  AND2_X1 U9139 ( .A1(n9173), .A2(n9314), .ZN(n9312) );
  OR2_X1 U9140 ( .A1(n9175), .A2(n9176), .ZN(n9314) );
  OR2_X1 U9141 ( .A1(n8016), .A2(n7501), .ZN(n9176) );
  OR2_X1 U9142 ( .A1(n9315), .A2(n9316), .ZN(n9175) );
  AND2_X1 U9143 ( .A1(n9172), .A2(n9171), .ZN(n9316) );
  AND2_X1 U9144 ( .A1(n9169), .A2(n9317), .ZN(n9315) );
  OR2_X1 U9145 ( .A1(n9171), .A2(n9172), .ZN(n9317) );
  OR2_X1 U9146 ( .A1(n8019), .A2(n7501), .ZN(n9172) );
  OR2_X1 U9147 ( .A1(n9318), .A2(n9319), .ZN(n9171) );
  AND2_X1 U9148 ( .A1(n9168), .A2(n9167), .ZN(n9319) );
  AND2_X1 U9149 ( .A1(n9165), .A2(n9320), .ZN(n9318) );
  OR2_X1 U9150 ( .A1(n9167), .A2(n9168), .ZN(n9320) );
  OR2_X1 U9151 ( .A1(n8023), .A2(n7501), .ZN(n9168) );
  OR2_X1 U9152 ( .A1(n9321), .A2(n9322), .ZN(n9167) );
  AND2_X1 U9153 ( .A1(n9164), .A2(n9163), .ZN(n9322) );
  AND2_X1 U9154 ( .A1(n9161), .A2(n9323), .ZN(n9321) );
  OR2_X1 U9155 ( .A1(n9163), .A2(n9164), .ZN(n9323) );
  OR2_X1 U9156 ( .A1(n8026), .A2(n7501), .ZN(n9164) );
  OR2_X1 U9157 ( .A1(n9324), .A2(n9325), .ZN(n9163) );
  AND2_X1 U9158 ( .A1(n9160), .A2(n9159), .ZN(n9325) );
  AND2_X1 U9159 ( .A1(n9157), .A2(n9326), .ZN(n9324) );
  OR2_X1 U9160 ( .A1(n9159), .A2(n9160), .ZN(n9326) );
  OR2_X1 U9161 ( .A1(n8030), .A2(n7501), .ZN(n9160) );
  OR2_X1 U9162 ( .A1(n9327), .A2(n9328), .ZN(n9159) );
  AND2_X1 U9163 ( .A1(n9156), .A2(n9155), .ZN(n9328) );
  AND2_X1 U9164 ( .A1(n9153), .A2(n9329), .ZN(n9327) );
  OR2_X1 U9165 ( .A1(n9155), .A2(n9156), .ZN(n9329) );
  OR2_X1 U9166 ( .A1(n8034), .A2(n7501), .ZN(n9156) );
  OR2_X1 U9167 ( .A1(n9330), .A2(n9331), .ZN(n9155) );
  AND2_X1 U9168 ( .A1(n9152), .A2(n9151), .ZN(n9331) );
  AND2_X1 U9169 ( .A1(n9149), .A2(n9332), .ZN(n9330) );
  OR2_X1 U9170 ( .A1(n9151), .A2(n9152), .ZN(n9332) );
  OR2_X1 U9171 ( .A1(n8037), .A2(n7501), .ZN(n9152) );
  OR2_X1 U9172 ( .A1(n9333), .A2(n9334), .ZN(n9151) );
  AND2_X1 U9173 ( .A1(n9148), .A2(n9147), .ZN(n9334) );
  AND2_X1 U9174 ( .A1(n9145), .A2(n9335), .ZN(n9333) );
  OR2_X1 U9175 ( .A1(n9147), .A2(n9148), .ZN(n9335) );
  OR2_X1 U9176 ( .A1(n8041), .A2(n7501), .ZN(n9148) );
  OR2_X1 U9177 ( .A1(n9336), .A2(n9337), .ZN(n9147) );
  AND2_X1 U9178 ( .A1(n9144), .A2(n9143), .ZN(n9337) );
  AND2_X1 U9179 ( .A1(n9141), .A2(n9338), .ZN(n9336) );
  OR2_X1 U9180 ( .A1(n9143), .A2(n9144), .ZN(n9338) );
  OR2_X1 U9181 ( .A1(n8044), .A2(n7501), .ZN(n9144) );
  OR2_X1 U9182 ( .A1(n9339), .A2(n9340), .ZN(n9143) );
  AND2_X1 U9183 ( .A1(n9140), .A2(n9139), .ZN(n9340) );
  AND2_X1 U9184 ( .A1(n9137), .A2(n9341), .ZN(n9339) );
  OR2_X1 U9185 ( .A1(n9139), .A2(n9140), .ZN(n9341) );
  OR2_X1 U9186 ( .A1(n8048), .A2(n7501), .ZN(n9140) );
  OR2_X1 U9187 ( .A1(n9342), .A2(n9343), .ZN(n9139) );
  AND2_X1 U9188 ( .A1(n8052), .A2(n9344), .ZN(n9343) );
  AND2_X1 U9189 ( .A1(n9345), .A2(n9346), .ZN(n9342) );
  OR2_X1 U9190 ( .A1(n9344), .A2(n8052), .ZN(n9346) );
  INV_X1 U9191 ( .A(n7505), .ZN(n8052) );
  AND2_X1 U9192 ( .A1(a_29_), .A2(b_29_), .ZN(n7505) );
  INV_X1 U9193 ( .A(n9136), .ZN(n9344) );
  AND3_X1 U9194 ( .A1(n8904), .A2(b_29_), .A3(b_28_), .ZN(n9136) );
  INV_X1 U9195 ( .A(n9135), .ZN(n9345) );
  OR2_X1 U9196 ( .A1(n9347), .A2(n9348), .ZN(n9135) );
  AND2_X1 U9197 ( .A1(b_28_), .A2(n9349), .ZN(n9348) );
  OR2_X1 U9198 ( .A1(n9350), .A2(n7490), .ZN(n9349) );
  AND2_X1 U9199 ( .A1(a_30_), .A2(n7540), .ZN(n9350) );
  AND2_X1 U9200 ( .A1(b_27_), .A2(n9351), .ZN(n9347) );
  OR2_X1 U9201 ( .A1(n9352), .A2(n7493), .ZN(n9351) );
  AND2_X1 U9202 ( .A1(a_31_), .A2(n8049), .ZN(n9352) );
  XNOR2_X1 U9203 ( .A(n9353), .B(n9354), .ZN(n9137) );
  XNOR2_X1 U9204 ( .A(n9355), .B(n9356), .ZN(n9354) );
  XOR2_X1 U9205 ( .A(n9357), .B(n9358), .Z(n9141) );
  XOR2_X1 U9206 ( .A(n9359), .B(n7521), .Z(n9358) );
  XOR2_X1 U9207 ( .A(n9360), .B(n9361), .Z(n9145) );
  XOR2_X1 U9208 ( .A(n9362), .B(n9363), .Z(n9361) );
  XOR2_X1 U9209 ( .A(n9364), .B(n9365), .Z(n9149) );
  XOR2_X1 U9210 ( .A(n9366), .B(n9367), .Z(n9365) );
  XOR2_X1 U9211 ( .A(n9368), .B(n9369), .Z(n9153) );
  XOR2_X1 U9212 ( .A(n9370), .B(n9371), .Z(n9369) );
  XOR2_X1 U9213 ( .A(n9372), .B(n9373), .Z(n9157) );
  XOR2_X1 U9214 ( .A(n9374), .B(n9375), .Z(n9373) );
  XOR2_X1 U9215 ( .A(n9376), .B(n9377), .Z(n9161) );
  XOR2_X1 U9216 ( .A(n9378), .B(n9379), .Z(n9377) );
  XOR2_X1 U9217 ( .A(n9380), .B(n9381), .Z(n9165) );
  XOR2_X1 U9218 ( .A(n9382), .B(n9383), .Z(n9381) );
  XOR2_X1 U9219 ( .A(n9384), .B(n9385), .Z(n9169) );
  XOR2_X1 U9220 ( .A(n9386), .B(n9387), .Z(n9385) );
  XOR2_X1 U9221 ( .A(n9388), .B(n9389), .Z(n9173) );
  XOR2_X1 U9222 ( .A(n9390), .B(n9391), .Z(n9389) );
  XOR2_X1 U9223 ( .A(n9392), .B(n9393), .Z(n9177) );
  XOR2_X1 U9224 ( .A(n9394), .B(n9395), .Z(n9393) );
  XOR2_X1 U9225 ( .A(n9396), .B(n9397), .Z(n9181) );
  XOR2_X1 U9226 ( .A(n9398), .B(n9399), .Z(n9397) );
  XOR2_X1 U9227 ( .A(n9400), .B(n9401), .Z(n9185) );
  XOR2_X1 U9228 ( .A(n9402), .B(n9403), .Z(n9401) );
  XOR2_X1 U9229 ( .A(n9404), .B(n9405), .Z(n9189) );
  XOR2_X1 U9230 ( .A(n9406), .B(n9407), .Z(n9405) );
  XOR2_X1 U9231 ( .A(n9408), .B(n9409), .Z(n9193) );
  XOR2_X1 U9232 ( .A(n9410), .B(n9411), .Z(n9409) );
  XOR2_X1 U9233 ( .A(n9412), .B(n9413), .Z(n9197) );
  XOR2_X1 U9234 ( .A(n9414), .B(n9415), .Z(n9413) );
  XOR2_X1 U9235 ( .A(n9416), .B(n9417), .Z(n9201) );
  XOR2_X1 U9236 ( .A(n9418), .B(n9419), .Z(n9417) );
  XOR2_X1 U9237 ( .A(n9420), .B(n9421), .Z(n9205) );
  XOR2_X1 U9238 ( .A(n9422), .B(n9423), .Z(n9421) );
  XOR2_X1 U9239 ( .A(n9424), .B(n9425), .Z(n9209) );
  XOR2_X1 U9240 ( .A(n9426), .B(n9427), .Z(n9425) );
  XOR2_X1 U9241 ( .A(n9428), .B(n9429), .Z(n9213) );
  XOR2_X1 U9242 ( .A(n9430), .B(n9431), .Z(n9429) );
  XOR2_X1 U9243 ( .A(n9432), .B(n9433), .Z(n9217) );
  XOR2_X1 U9244 ( .A(n9434), .B(n9435), .Z(n9433) );
  XOR2_X1 U9245 ( .A(n9436), .B(n9437), .Z(n9221) );
  XOR2_X1 U9246 ( .A(n9438), .B(n9439), .Z(n9437) );
  XOR2_X1 U9247 ( .A(n9440), .B(n9441), .Z(n9225) );
  XOR2_X1 U9248 ( .A(n9442), .B(n9443), .Z(n9441) );
  XOR2_X1 U9249 ( .A(n9444), .B(n9445), .Z(n9229) );
  XOR2_X1 U9250 ( .A(n9446), .B(n9447), .Z(n9445) );
  XOR2_X1 U9251 ( .A(n9448), .B(n9449), .Z(n9233) );
  XOR2_X1 U9252 ( .A(n9450), .B(n9451), .Z(n9449) );
  XOR2_X1 U9253 ( .A(n9452), .B(n9453), .Z(n9237) );
  XOR2_X1 U9254 ( .A(n9454), .B(n9455), .Z(n9453) );
  OR2_X1 U9255 ( .A1(n7956), .A2(n7501), .ZN(n9243) );
  INV_X1 U9256 ( .A(b_29_), .ZN(n7501) );
  XOR2_X1 U9257 ( .A(n9456), .B(n9457), .Z(n9242) );
  XOR2_X1 U9258 ( .A(n9458), .B(n9459), .Z(n9457) );
  XNOR2_X1 U9259 ( .A(n9460), .B(n9461), .ZN(n9245) );
  XNOR2_X1 U9260 ( .A(n9462), .B(n9463), .ZN(n9460) );
  XOR2_X1 U9261 ( .A(n9464), .B(n9465), .Z(n9034) );
  XOR2_X1 U9262 ( .A(n9466), .B(n9467), .Z(n9465) );
  OR2_X1 U9263 ( .A1(n9468), .A2(n8799), .ZN(n8081) );
  INV_X1 U9264 ( .A(n9469), .ZN(n8799) );
  OR2_X1 U9265 ( .A1(n9470), .A2(n8795), .ZN(n9469) );
  AND2_X1 U9266 ( .A1(n9471), .A2(n9472), .ZN(n9470) );
  AND2_X1 U9267 ( .A1(n8798), .A2(n8797), .ZN(n9468) );
  XNOR2_X1 U9268 ( .A(n9473), .B(n9474), .ZN(n8797) );
  XOR2_X1 U9269 ( .A(n9475), .B(n9476), .Z(n9474) );
  INV_X1 U9270 ( .A(n9250), .ZN(n8798) );
  OR2_X1 U9271 ( .A1(n9477), .A2(n9478), .ZN(n9250) );
  AND2_X1 U9272 ( .A1(n9254), .A2(n9253), .ZN(n9478) );
  AND2_X1 U9273 ( .A1(n9251), .A2(n9479), .ZN(n9477) );
  OR2_X1 U9274 ( .A1(n9253), .A2(n9254), .ZN(n9479) );
  OR2_X1 U9275 ( .A1(n7950), .A2(n8049), .ZN(n9254) );
  OR2_X1 U9276 ( .A1(n9480), .A2(n9481), .ZN(n9253) );
  AND2_X1 U9277 ( .A1(n9467), .A2(n9466), .ZN(n9481) );
  AND2_X1 U9278 ( .A1(n9464), .A2(n9482), .ZN(n9480) );
  OR2_X1 U9279 ( .A1(n9466), .A2(n9467), .ZN(n9482) );
  OR2_X1 U9280 ( .A1(n7953), .A2(n8049), .ZN(n9467) );
  OR2_X1 U9281 ( .A1(n9483), .A2(n9484), .ZN(n9466) );
  AND2_X1 U9282 ( .A1(n9463), .A2(n9462), .ZN(n9484) );
  AND2_X1 U9283 ( .A1(n9461), .A2(n9485), .ZN(n9483) );
  OR2_X1 U9284 ( .A1(n9462), .A2(n9463), .ZN(n9485) );
  OR2_X1 U9285 ( .A1(n9486), .A2(n9487), .ZN(n9463) );
  AND2_X1 U9286 ( .A1(n9459), .A2(n9458), .ZN(n9487) );
  AND2_X1 U9287 ( .A1(n9456), .A2(n9488), .ZN(n9486) );
  OR2_X1 U9288 ( .A1(n9458), .A2(n9459), .ZN(n9488) );
  OR2_X1 U9289 ( .A1(n7960), .A2(n8049), .ZN(n9459) );
  OR2_X1 U9290 ( .A1(n9489), .A2(n9490), .ZN(n9458) );
  AND2_X1 U9291 ( .A1(n9455), .A2(n9454), .ZN(n9490) );
  AND2_X1 U9292 ( .A1(n9452), .A2(n9491), .ZN(n9489) );
  OR2_X1 U9293 ( .A1(n9454), .A2(n9455), .ZN(n9491) );
  OR2_X1 U9294 ( .A1(n7963), .A2(n8049), .ZN(n9455) );
  OR2_X1 U9295 ( .A1(n9492), .A2(n9493), .ZN(n9454) );
  AND2_X1 U9296 ( .A1(n9451), .A2(n9450), .ZN(n9493) );
  AND2_X1 U9297 ( .A1(n9448), .A2(n9494), .ZN(n9492) );
  OR2_X1 U9298 ( .A1(n9450), .A2(n9451), .ZN(n9494) );
  OR2_X1 U9299 ( .A1(n7967), .A2(n8049), .ZN(n9451) );
  OR2_X1 U9300 ( .A1(n9495), .A2(n9496), .ZN(n9450) );
  AND2_X1 U9301 ( .A1(n9447), .A2(n9446), .ZN(n9496) );
  AND2_X1 U9302 ( .A1(n9444), .A2(n9497), .ZN(n9495) );
  OR2_X1 U9303 ( .A1(n9446), .A2(n9447), .ZN(n9497) );
  OR2_X1 U9304 ( .A1(n7970), .A2(n8049), .ZN(n9447) );
  OR2_X1 U9305 ( .A1(n9498), .A2(n9499), .ZN(n9446) );
  AND2_X1 U9306 ( .A1(n9443), .A2(n9442), .ZN(n9499) );
  AND2_X1 U9307 ( .A1(n9440), .A2(n9500), .ZN(n9498) );
  OR2_X1 U9308 ( .A1(n9442), .A2(n9443), .ZN(n9500) );
  OR2_X1 U9309 ( .A1(n7974), .A2(n8049), .ZN(n9443) );
  OR2_X1 U9310 ( .A1(n9501), .A2(n9502), .ZN(n9442) );
  AND2_X1 U9311 ( .A1(n9439), .A2(n9438), .ZN(n9502) );
  AND2_X1 U9312 ( .A1(n9436), .A2(n9503), .ZN(n9501) );
  OR2_X1 U9313 ( .A1(n9438), .A2(n9439), .ZN(n9503) );
  OR2_X1 U9314 ( .A1(n7977), .A2(n8049), .ZN(n9439) );
  OR2_X1 U9315 ( .A1(n9504), .A2(n9505), .ZN(n9438) );
  AND2_X1 U9316 ( .A1(n9435), .A2(n9434), .ZN(n9505) );
  AND2_X1 U9317 ( .A1(n9432), .A2(n9506), .ZN(n9504) );
  OR2_X1 U9318 ( .A1(n9434), .A2(n9435), .ZN(n9506) );
  OR2_X1 U9319 ( .A1(n7981), .A2(n8049), .ZN(n9435) );
  OR2_X1 U9320 ( .A1(n9507), .A2(n9508), .ZN(n9434) );
  AND2_X1 U9321 ( .A1(n9431), .A2(n9430), .ZN(n9508) );
  AND2_X1 U9322 ( .A1(n9428), .A2(n9509), .ZN(n9507) );
  OR2_X1 U9323 ( .A1(n9430), .A2(n9431), .ZN(n9509) );
  OR2_X1 U9324 ( .A1(n7984), .A2(n8049), .ZN(n9431) );
  OR2_X1 U9325 ( .A1(n9510), .A2(n9511), .ZN(n9430) );
  AND2_X1 U9326 ( .A1(n9427), .A2(n9426), .ZN(n9511) );
  AND2_X1 U9327 ( .A1(n9424), .A2(n9512), .ZN(n9510) );
  OR2_X1 U9328 ( .A1(n9426), .A2(n9427), .ZN(n9512) );
  OR2_X1 U9329 ( .A1(n7988), .A2(n8049), .ZN(n9427) );
  OR2_X1 U9330 ( .A1(n9513), .A2(n9514), .ZN(n9426) );
  AND2_X1 U9331 ( .A1(n9423), .A2(n9422), .ZN(n9514) );
  AND2_X1 U9332 ( .A1(n9420), .A2(n9515), .ZN(n9513) );
  OR2_X1 U9333 ( .A1(n9422), .A2(n9423), .ZN(n9515) );
  OR2_X1 U9334 ( .A1(n7991), .A2(n8049), .ZN(n9423) );
  OR2_X1 U9335 ( .A1(n9516), .A2(n9517), .ZN(n9422) );
  AND2_X1 U9336 ( .A1(n9419), .A2(n9418), .ZN(n9517) );
  AND2_X1 U9337 ( .A1(n9416), .A2(n9518), .ZN(n9516) );
  OR2_X1 U9338 ( .A1(n9418), .A2(n9419), .ZN(n9518) );
  OR2_X1 U9339 ( .A1(n7995), .A2(n8049), .ZN(n9419) );
  OR2_X1 U9340 ( .A1(n9519), .A2(n9520), .ZN(n9418) );
  AND2_X1 U9341 ( .A1(n9415), .A2(n9414), .ZN(n9520) );
  AND2_X1 U9342 ( .A1(n9412), .A2(n9521), .ZN(n9519) );
  OR2_X1 U9343 ( .A1(n9414), .A2(n9415), .ZN(n9521) );
  OR2_X1 U9344 ( .A1(n7998), .A2(n8049), .ZN(n9415) );
  OR2_X1 U9345 ( .A1(n9522), .A2(n9523), .ZN(n9414) );
  AND2_X1 U9346 ( .A1(n9411), .A2(n9410), .ZN(n9523) );
  AND2_X1 U9347 ( .A1(n9408), .A2(n9524), .ZN(n9522) );
  OR2_X1 U9348 ( .A1(n9410), .A2(n9411), .ZN(n9524) );
  OR2_X1 U9349 ( .A1(n8002), .A2(n8049), .ZN(n9411) );
  OR2_X1 U9350 ( .A1(n9525), .A2(n9526), .ZN(n9410) );
  AND2_X1 U9351 ( .A1(n9407), .A2(n9406), .ZN(n9526) );
  AND2_X1 U9352 ( .A1(n9404), .A2(n9527), .ZN(n9525) );
  OR2_X1 U9353 ( .A1(n9406), .A2(n9407), .ZN(n9527) );
  OR2_X1 U9354 ( .A1(n8005), .A2(n8049), .ZN(n9407) );
  OR2_X1 U9355 ( .A1(n9528), .A2(n9529), .ZN(n9406) );
  AND2_X1 U9356 ( .A1(n9403), .A2(n9402), .ZN(n9529) );
  AND2_X1 U9357 ( .A1(n9400), .A2(n9530), .ZN(n9528) );
  OR2_X1 U9358 ( .A1(n9402), .A2(n9403), .ZN(n9530) );
  OR2_X1 U9359 ( .A1(n8009), .A2(n8049), .ZN(n9403) );
  OR2_X1 U9360 ( .A1(n9531), .A2(n9532), .ZN(n9402) );
  AND2_X1 U9361 ( .A1(n9399), .A2(n9398), .ZN(n9532) );
  AND2_X1 U9362 ( .A1(n9396), .A2(n9533), .ZN(n9531) );
  OR2_X1 U9363 ( .A1(n9398), .A2(n9399), .ZN(n9533) );
  OR2_X1 U9364 ( .A1(n8012), .A2(n8049), .ZN(n9399) );
  OR2_X1 U9365 ( .A1(n9534), .A2(n9535), .ZN(n9398) );
  AND2_X1 U9366 ( .A1(n9395), .A2(n9394), .ZN(n9535) );
  AND2_X1 U9367 ( .A1(n9392), .A2(n9536), .ZN(n9534) );
  OR2_X1 U9368 ( .A1(n9394), .A2(n9395), .ZN(n9536) );
  OR2_X1 U9369 ( .A1(n8016), .A2(n8049), .ZN(n9395) );
  OR2_X1 U9370 ( .A1(n9537), .A2(n9538), .ZN(n9394) );
  AND2_X1 U9371 ( .A1(n9391), .A2(n9390), .ZN(n9538) );
  AND2_X1 U9372 ( .A1(n9388), .A2(n9539), .ZN(n9537) );
  OR2_X1 U9373 ( .A1(n9390), .A2(n9391), .ZN(n9539) );
  OR2_X1 U9374 ( .A1(n8019), .A2(n8049), .ZN(n9391) );
  OR2_X1 U9375 ( .A1(n9540), .A2(n9541), .ZN(n9390) );
  AND2_X1 U9376 ( .A1(n9387), .A2(n9386), .ZN(n9541) );
  AND2_X1 U9377 ( .A1(n9384), .A2(n9542), .ZN(n9540) );
  OR2_X1 U9378 ( .A1(n9386), .A2(n9387), .ZN(n9542) );
  OR2_X1 U9379 ( .A1(n8023), .A2(n8049), .ZN(n9387) );
  OR2_X1 U9380 ( .A1(n9543), .A2(n9544), .ZN(n9386) );
  AND2_X1 U9381 ( .A1(n9383), .A2(n9382), .ZN(n9544) );
  AND2_X1 U9382 ( .A1(n9380), .A2(n9545), .ZN(n9543) );
  OR2_X1 U9383 ( .A1(n9382), .A2(n9383), .ZN(n9545) );
  OR2_X1 U9384 ( .A1(n8026), .A2(n8049), .ZN(n9383) );
  OR2_X1 U9385 ( .A1(n9546), .A2(n9547), .ZN(n9382) );
  AND2_X1 U9386 ( .A1(n9379), .A2(n9378), .ZN(n9547) );
  AND2_X1 U9387 ( .A1(n9376), .A2(n9548), .ZN(n9546) );
  OR2_X1 U9388 ( .A1(n9378), .A2(n9379), .ZN(n9548) );
  OR2_X1 U9389 ( .A1(n8030), .A2(n8049), .ZN(n9379) );
  OR2_X1 U9390 ( .A1(n9549), .A2(n9550), .ZN(n9378) );
  AND2_X1 U9391 ( .A1(n9375), .A2(n9374), .ZN(n9550) );
  AND2_X1 U9392 ( .A1(n9372), .A2(n9551), .ZN(n9549) );
  OR2_X1 U9393 ( .A1(n9374), .A2(n9375), .ZN(n9551) );
  OR2_X1 U9394 ( .A1(n8034), .A2(n8049), .ZN(n9375) );
  OR2_X1 U9395 ( .A1(n9552), .A2(n9553), .ZN(n9374) );
  AND2_X1 U9396 ( .A1(n9371), .A2(n9370), .ZN(n9553) );
  AND2_X1 U9397 ( .A1(n9368), .A2(n9554), .ZN(n9552) );
  OR2_X1 U9398 ( .A1(n9370), .A2(n9371), .ZN(n9554) );
  OR2_X1 U9399 ( .A1(n8037), .A2(n8049), .ZN(n9371) );
  OR2_X1 U9400 ( .A1(n9555), .A2(n9556), .ZN(n9370) );
  AND2_X1 U9401 ( .A1(n9367), .A2(n9366), .ZN(n9556) );
  AND2_X1 U9402 ( .A1(n9364), .A2(n9557), .ZN(n9555) );
  OR2_X1 U9403 ( .A1(n9366), .A2(n9367), .ZN(n9557) );
  OR2_X1 U9404 ( .A1(n8041), .A2(n8049), .ZN(n9367) );
  OR2_X1 U9405 ( .A1(n9558), .A2(n9559), .ZN(n9366) );
  AND2_X1 U9406 ( .A1(n9363), .A2(n9362), .ZN(n9559) );
  AND2_X1 U9407 ( .A1(n9360), .A2(n9560), .ZN(n9558) );
  OR2_X1 U9408 ( .A1(n9362), .A2(n9363), .ZN(n9560) );
  OR2_X1 U9409 ( .A1(n8044), .A2(n8049), .ZN(n9363) );
  OR2_X1 U9410 ( .A1(n9561), .A2(n9562), .ZN(n9362) );
  AND2_X1 U9411 ( .A1(n7521), .A2(n9359), .ZN(n9562) );
  AND2_X1 U9412 ( .A1(n9357), .A2(n9563), .ZN(n9561) );
  OR2_X1 U9413 ( .A1(n9359), .A2(n7521), .ZN(n9563) );
  OR2_X1 U9414 ( .A1(n8048), .A2(n8049), .ZN(n7521) );
  OR2_X1 U9415 ( .A1(n9564), .A2(n9565), .ZN(n9359) );
  AND2_X1 U9416 ( .A1(n9353), .A2(n9566), .ZN(n9565) );
  AND2_X1 U9417 ( .A1(n9567), .A2(n9568), .ZN(n9564) );
  OR2_X1 U9418 ( .A1(n9566), .A2(n9353), .ZN(n9568) );
  OR2_X1 U9419 ( .A1(n8051), .A2(n8049), .ZN(n9353) );
  INV_X1 U9420 ( .A(n9356), .ZN(n9566) );
  AND3_X1 U9421 ( .A1(n8904), .A2(b_28_), .A3(b_27_), .ZN(n9356) );
  INV_X1 U9422 ( .A(n9355), .ZN(n9567) );
  OR2_X1 U9423 ( .A1(n9569), .A2(n9570), .ZN(n9355) );
  AND2_X1 U9424 ( .A1(b_27_), .A2(n9571), .ZN(n9570) );
  OR2_X1 U9425 ( .A1(n9572), .A2(n7490), .ZN(n9571) );
  AND2_X1 U9426 ( .A1(a_30_), .A2(n8042), .ZN(n9572) );
  AND2_X1 U9427 ( .A1(b_26_), .A2(n9573), .ZN(n9569) );
  OR2_X1 U9428 ( .A1(n9574), .A2(n7493), .ZN(n9573) );
  AND2_X1 U9429 ( .A1(a_31_), .A2(n7540), .ZN(n9574) );
  XNOR2_X1 U9430 ( .A(n9575), .B(n9576), .ZN(n9357) );
  XNOR2_X1 U9431 ( .A(n9577), .B(n9578), .ZN(n9576) );
  XOR2_X1 U9432 ( .A(n9579), .B(n9580), .Z(n9360) );
  XOR2_X1 U9433 ( .A(n9581), .B(n9582), .Z(n9580) );
  XOR2_X1 U9434 ( .A(n9583), .B(n9584), .Z(n9364) );
  XNOR2_X1 U9435 ( .A(n9585), .B(n7544), .ZN(n9584) );
  XOR2_X1 U9436 ( .A(n9586), .B(n9587), .Z(n9368) );
  XOR2_X1 U9437 ( .A(n9588), .B(n9589), .Z(n9587) );
  XOR2_X1 U9438 ( .A(n9590), .B(n9591), .Z(n9372) );
  XOR2_X1 U9439 ( .A(n9592), .B(n9593), .Z(n9591) );
  XOR2_X1 U9440 ( .A(n9594), .B(n9595), .Z(n9376) );
  XOR2_X1 U9441 ( .A(n9596), .B(n9597), .Z(n9595) );
  XOR2_X1 U9442 ( .A(n9598), .B(n9599), .Z(n9380) );
  XOR2_X1 U9443 ( .A(n9600), .B(n9601), .Z(n9599) );
  XOR2_X1 U9444 ( .A(n9602), .B(n9603), .Z(n9384) );
  XOR2_X1 U9445 ( .A(n9604), .B(n9605), .Z(n9603) );
  XOR2_X1 U9446 ( .A(n9606), .B(n9607), .Z(n9388) );
  XOR2_X1 U9447 ( .A(n9608), .B(n9609), .Z(n9607) );
  XOR2_X1 U9448 ( .A(n9610), .B(n9611), .Z(n9392) );
  XOR2_X1 U9449 ( .A(n9612), .B(n9613), .Z(n9611) );
  XOR2_X1 U9450 ( .A(n9614), .B(n9615), .Z(n9396) );
  XOR2_X1 U9451 ( .A(n9616), .B(n9617), .Z(n9615) );
  XOR2_X1 U9452 ( .A(n9618), .B(n9619), .Z(n9400) );
  XOR2_X1 U9453 ( .A(n9620), .B(n9621), .Z(n9619) );
  XOR2_X1 U9454 ( .A(n9622), .B(n9623), .Z(n9404) );
  XOR2_X1 U9455 ( .A(n9624), .B(n9625), .Z(n9623) );
  XOR2_X1 U9456 ( .A(n9626), .B(n9627), .Z(n9408) );
  XOR2_X1 U9457 ( .A(n9628), .B(n9629), .Z(n9627) );
  XOR2_X1 U9458 ( .A(n9630), .B(n9631), .Z(n9412) );
  XOR2_X1 U9459 ( .A(n9632), .B(n9633), .Z(n9631) );
  XOR2_X1 U9460 ( .A(n9634), .B(n9635), .Z(n9416) );
  XOR2_X1 U9461 ( .A(n9636), .B(n9637), .Z(n9635) );
  XOR2_X1 U9462 ( .A(n9638), .B(n9639), .Z(n9420) );
  XOR2_X1 U9463 ( .A(n9640), .B(n9641), .Z(n9639) );
  XOR2_X1 U9464 ( .A(n9642), .B(n9643), .Z(n9424) );
  XOR2_X1 U9465 ( .A(n9644), .B(n9645), .Z(n9643) );
  XOR2_X1 U9466 ( .A(n9646), .B(n9647), .Z(n9428) );
  XOR2_X1 U9467 ( .A(n9648), .B(n9649), .Z(n9647) );
  XOR2_X1 U9468 ( .A(n9650), .B(n9651), .Z(n9432) );
  XOR2_X1 U9469 ( .A(n9652), .B(n9653), .Z(n9651) );
  XOR2_X1 U9470 ( .A(n9654), .B(n9655), .Z(n9436) );
  XOR2_X1 U9471 ( .A(n9656), .B(n9657), .Z(n9655) );
  XOR2_X1 U9472 ( .A(n9658), .B(n9659), .Z(n9440) );
  XOR2_X1 U9473 ( .A(n9660), .B(n9661), .Z(n9659) );
  XOR2_X1 U9474 ( .A(n9662), .B(n9663), .Z(n9444) );
  XOR2_X1 U9475 ( .A(n9664), .B(n9665), .Z(n9663) );
  XNOR2_X1 U9476 ( .A(n9666), .B(n9667), .ZN(n9448) );
  XNOR2_X1 U9477 ( .A(n9668), .B(n9669), .ZN(n9666) );
  XOR2_X1 U9478 ( .A(n9670), .B(n9671), .Z(n9452) );
  XOR2_X1 U9479 ( .A(n9672), .B(n9673), .Z(n9671) );
  XOR2_X1 U9480 ( .A(n9674), .B(n9675), .Z(n9456) );
  XOR2_X1 U9481 ( .A(n9676), .B(n9677), .Z(n9675) );
  OR2_X1 U9482 ( .A1(n7956), .A2(n8049), .ZN(n9462) );
  INV_X1 U9483 ( .A(b_28_), .ZN(n8049) );
  XOR2_X1 U9484 ( .A(n9678), .B(n9679), .Z(n9461) );
  XOR2_X1 U9485 ( .A(n9680), .B(n9681), .Z(n9679) );
  XNOR2_X1 U9486 ( .A(n9682), .B(n9683), .ZN(n9464) );
  XNOR2_X1 U9487 ( .A(n9684), .B(n9685), .ZN(n9682) );
  XOR2_X1 U9488 ( .A(n9686), .B(n9687), .Z(n9251) );
  XOR2_X1 U9489 ( .A(n9688), .B(n9689), .Z(n9687) );
  OR2_X1 U9490 ( .A1(n8795), .A2(n8794), .ZN(n8087) );
  XNOR2_X1 U9491 ( .A(n8790), .B(n9690), .ZN(n8794) );
  INV_X1 U9492 ( .A(n9691), .ZN(n8795) );
  OR2_X1 U9493 ( .A1(n9471), .A2(n9472), .ZN(n9691) );
  OR2_X1 U9494 ( .A1(n9692), .A2(n9693), .ZN(n9472) );
  AND2_X1 U9495 ( .A1(n9473), .A2(n9476), .ZN(n9693) );
  AND2_X1 U9496 ( .A1(n9694), .A2(n9475), .ZN(n9692) );
  OR2_X1 U9497 ( .A1(n9695), .A2(n9696), .ZN(n9475) );
  AND2_X1 U9498 ( .A1(n9686), .A2(n9689), .ZN(n9696) );
  AND2_X1 U9499 ( .A1(n9697), .A2(n9688), .ZN(n9695) );
  OR2_X1 U9500 ( .A1(n9698), .A2(n9699), .ZN(n9688) );
  AND2_X1 U9501 ( .A1(n9685), .A2(n9684), .ZN(n9699) );
  AND2_X1 U9502 ( .A1(n9683), .A2(n9700), .ZN(n9698) );
  OR2_X1 U9503 ( .A1(n9684), .A2(n9685), .ZN(n9700) );
  OR2_X1 U9504 ( .A1(n9701), .A2(n9702), .ZN(n9685) );
  AND2_X1 U9505 ( .A1(n9681), .A2(n9680), .ZN(n9702) );
  AND2_X1 U9506 ( .A1(n9678), .A2(n9703), .ZN(n9701) );
  OR2_X1 U9507 ( .A1(n9680), .A2(n9681), .ZN(n9703) );
  OR2_X1 U9508 ( .A1(n7960), .A2(n7540), .ZN(n9681) );
  OR2_X1 U9509 ( .A1(n9704), .A2(n9705), .ZN(n9680) );
  AND2_X1 U9510 ( .A1(n9677), .A2(n9676), .ZN(n9705) );
  AND2_X1 U9511 ( .A1(n9674), .A2(n9706), .ZN(n9704) );
  OR2_X1 U9512 ( .A1(n9676), .A2(n9677), .ZN(n9706) );
  OR2_X1 U9513 ( .A1(n7963), .A2(n7540), .ZN(n9677) );
  OR2_X1 U9514 ( .A1(n9707), .A2(n9708), .ZN(n9676) );
  AND2_X1 U9515 ( .A1(n9673), .A2(n9672), .ZN(n9708) );
  AND2_X1 U9516 ( .A1(n9670), .A2(n9709), .ZN(n9707) );
  OR2_X1 U9517 ( .A1(n9672), .A2(n9673), .ZN(n9709) );
  OR2_X1 U9518 ( .A1(n7967), .A2(n7540), .ZN(n9673) );
  OR2_X1 U9519 ( .A1(n9710), .A2(n9711), .ZN(n9672) );
  AND2_X1 U9520 ( .A1(n9669), .A2(n9668), .ZN(n9711) );
  AND2_X1 U9521 ( .A1(n9667), .A2(n9712), .ZN(n9710) );
  OR2_X1 U9522 ( .A1(n9668), .A2(n9669), .ZN(n9712) );
  OR2_X1 U9523 ( .A1(n9713), .A2(n9714), .ZN(n9669) );
  AND2_X1 U9524 ( .A1(n9665), .A2(n9664), .ZN(n9714) );
  AND2_X1 U9525 ( .A1(n9662), .A2(n9715), .ZN(n9713) );
  OR2_X1 U9526 ( .A1(n9664), .A2(n9665), .ZN(n9715) );
  OR2_X1 U9527 ( .A1(n7974), .A2(n7540), .ZN(n9665) );
  OR2_X1 U9528 ( .A1(n9716), .A2(n9717), .ZN(n9664) );
  AND2_X1 U9529 ( .A1(n9661), .A2(n9660), .ZN(n9717) );
  AND2_X1 U9530 ( .A1(n9658), .A2(n9718), .ZN(n9716) );
  OR2_X1 U9531 ( .A1(n9660), .A2(n9661), .ZN(n9718) );
  OR2_X1 U9532 ( .A1(n7977), .A2(n7540), .ZN(n9661) );
  OR2_X1 U9533 ( .A1(n9719), .A2(n9720), .ZN(n9660) );
  AND2_X1 U9534 ( .A1(n9657), .A2(n9656), .ZN(n9720) );
  AND2_X1 U9535 ( .A1(n9654), .A2(n9721), .ZN(n9719) );
  OR2_X1 U9536 ( .A1(n9656), .A2(n9657), .ZN(n9721) );
  OR2_X1 U9537 ( .A1(n7981), .A2(n7540), .ZN(n9657) );
  OR2_X1 U9538 ( .A1(n9722), .A2(n9723), .ZN(n9656) );
  AND2_X1 U9539 ( .A1(n9653), .A2(n9652), .ZN(n9723) );
  AND2_X1 U9540 ( .A1(n9650), .A2(n9724), .ZN(n9722) );
  OR2_X1 U9541 ( .A1(n9652), .A2(n9653), .ZN(n9724) );
  OR2_X1 U9542 ( .A1(n7984), .A2(n7540), .ZN(n9653) );
  OR2_X1 U9543 ( .A1(n9725), .A2(n9726), .ZN(n9652) );
  AND2_X1 U9544 ( .A1(n9649), .A2(n9648), .ZN(n9726) );
  AND2_X1 U9545 ( .A1(n9646), .A2(n9727), .ZN(n9725) );
  OR2_X1 U9546 ( .A1(n9648), .A2(n9649), .ZN(n9727) );
  OR2_X1 U9547 ( .A1(n7988), .A2(n7540), .ZN(n9649) );
  OR2_X1 U9548 ( .A1(n9728), .A2(n9729), .ZN(n9648) );
  AND2_X1 U9549 ( .A1(n9645), .A2(n9644), .ZN(n9729) );
  AND2_X1 U9550 ( .A1(n9642), .A2(n9730), .ZN(n9728) );
  OR2_X1 U9551 ( .A1(n9644), .A2(n9645), .ZN(n9730) );
  OR2_X1 U9552 ( .A1(n7991), .A2(n7540), .ZN(n9645) );
  OR2_X1 U9553 ( .A1(n9731), .A2(n9732), .ZN(n9644) );
  AND2_X1 U9554 ( .A1(n9641), .A2(n9640), .ZN(n9732) );
  AND2_X1 U9555 ( .A1(n9638), .A2(n9733), .ZN(n9731) );
  OR2_X1 U9556 ( .A1(n9640), .A2(n9641), .ZN(n9733) );
  OR2_X1 U9557 ( .A1(n7995), .A2(n7540), .ZN(n9641) );
  OR2_X1 U9558 ( .A1(n9734), .A2(n9735), .ZN(n9640) );
  AND2_X1 U9559 ( .A1(n9637), .A2(n9636), .ZN(n9735) );
  AND2_X1 U9560 ( .A1(n9634), .A2(n9736), .ZN(n9734) );
  OR2_X1 U9561 ( .A1(n9636), .A2(n9637), .ZN(n9736) );
  OR2_X1 U9562 ( .A1(n7998), .A2(n7540), .ZN(n9637) );
  OR2_X1 U9563 ( .A1(n9737), .A2(n9738), .ZN(n9636) );
  AND2_X1 U9564 ( .A1(n9633), .A2(n9632), .ZN(n9738) );
  AND2_X1 U9565 ( .A1(n9630), .A2(n9739), .ZN(n9737) );
  OR2_X1 U9566 ( .A1(n9632), .A2(n9633), .ZN(n9739) );
  OR2_X1 U9567 ( .A1(n8002), .A2(n7540), .ZN(n9633) );
  OR2_X1 U9568 ( .A1(n9740), .A2(n9741), .ZN(n9632) );
  AND2_X1 U9569 ( .A1(n9629), .A2(n9628), .ZN(n9741) );
  AND2_X1 U9570 ( .A1(n9626), .A2(n9742), .ZN(n9740) );
  OR2_X1 U9571 ( .A1(n9628), .A2(n9629), .ZN(n9742) );
  OR2_X1 U9572 ( .A1(n8005), .A2(n7540), .ZN(n9629) );
  OR2_X1 U9573 ( .A1(n9743), .A2(n9744), .ZN(n9628) );
  AND2_X1 U9574 ( .A1(n9625), .A2(n9624), .ZN(n9744) );
  AND2_X1 U9575 ( .A1(n9622), .A2(n9745), .ZN(n9743) );
  OR2_X1 U9576 ( .A1(n9624), .A2(n9625), .ZN(n9745) );
  OR2_X1 U9577 ( .A1(n8009), .A2(n7540), .ZN(n9625) );
  OR2_X1 U9578 ( .A1(n9746), .A2(n9747), .ZN(n9624) );
  AND2_X1 U9579 ( .A1(n9621), .A2(n9620), .ZN(n9747) );
  AND2_X1 U9580 ( .A1(n9618), .A2(n9748), .ZN(n9746) );
  OR2_X1 U9581 ( .A1(n9620), .A2(n9621), .ZN(n9748) );
  OR2_X1 U9582 ( .A1(n8012), .A2(n7540), .ZN(n9621) );
  OR2_X1 U9583 ( .A1(n9749), .A2(n9750), .ZN(n9620) );
  AND2_X1 U9584 ( .A1(n9617), .A2(n9616), .ZN(n9750) );
  AND2_X1 U9585 ( .A1(n9614), .A2(n9751), .ZN(n9749) );
  OR2_X1 U9586 ( .A1(n9616), .A2(n9617), .ZN(n9751) );
  OR2_X1 U9587 ( .A1(n8016), .A2(n7540), .ZN(n9617) );
  OR2_X1 U9588 ( .A1(n9752), .A2(n9753), .ZN(n9616) );
  AND2_X1 U9589 ( .A1(n9613), .A2(n9612), .ZN(n9753) );
  AND2_X1 U9590 ( .A1(n9610), .A2(n9754), .ZN(n9752) );
  OR2_X1 U9591 ( .A1(n9612), .A2(n9613), .ZN(n9754) );
  OR2_X1 U9592 ( .A1(n8019), .A2(n7540), .ZN(n9613) );
  OR2_X1 U9593 ( .A1(n9755), .A2(n9756), .ZN(n9612) );
  AND2_X1 U9594 ( .A1(n9609), .A2(n9608), .ZN(n9756) );
  AND2_X1 U9595 ( .A1(n9606), .A2(n9757), .ZN(n9755) );
  OR2_X1 U9596 ( .A1(n9608), .A2(n9609), .ZN(n9757) );
  OR2_X1 U9597 ( .A1(n8023), .A2(n7540), .ZN(n9609) );
  OR2_X1 U9598 ( .A1(n9758), .A2(n9759), .ZN(n9608) );
  AND2_X1 U9599 ( .A1(n9605), .A2(n9604), .ZN(n9759) );
  AND2_X1 U9600 ( .A1(n9602), .A2(n9760), .ZN(n9758) );
  OR2_X1 U9601 ( .A1(n9604), .A2(n9605), .ZN(n9760) );
  OR2_X1 U9602 ( .A1(n8026), .A2(n7540), .ZN(n9605) );
  OR2_X1 U9603 ( .A1(n9761), .A2(n9762), .ZN(n9604) );
  AND2_X1 U9604 ( .A1(n9601), .A2(n9600), .ZN(n9762) );
  AND2_X1 U9605 ( .A1(n9598), .A2(n9763), .ZN(n9761) );
  OR2_X1 U9606 ( .A1(n9600), .A2(n9601), .ZN(n9763) );
  OR2_X1 U9607 ( .A1(n8030), .A2(n7540), .ZN(n9601) );
  OR2_X1 U9608 ( .A1(n9764), .A2(n9765), .ZN(n9600) );
  AND2_X1 U9609 ( .A1(n9597), .A2(n9596), .ZN(n9765) );
  AND2_X1 U9610 ( .A1(n9594), .A2(n9766), .ZN(n9764) );
  OR2_X1 U9611 ( .A1(n9596), .A2(n9597), .ZN(n9766) );
  OR2_X1 U9612 ( .A1(n8034), .A2(n7540), .ZN(n9597) );
  OR2_X1 U9613 ( .A1(n9767), .A2(n9768), .ZN(n9596) );
  AND2_X1 U9614 ( .A1(n9593), .A2(n9592), .ZN(n9768) );
  AND2_X1 U9615 ( .A1(n9590), .A2(n9769), .ZN(n9767) );
  OR2_X1 U9616 ( .A1(n9592), .A2(n9593), .ZN(n9769) );
  OR2_X1 U9617 ( .A1(n8037), .A2(n7540), .ZN(n9593) );
  OR2_X1 U9618 ( .A1(n9770), .A2(n9771), .ZN(n9592) );
  AND2_X1 U9619 ( .A1(n9589), .A2(n9588), .ZN(n9771) );
  AND2_X1 U9620 ( .A1(n9586), .A2(n9772), .ZN(n9770) );
  OR2_X1 U9621 ( .A1(n9588), .A2(n9589), .ZN(n9772) );
  OR2_X1 U9622 ( .A1(n8041), .A2(n7540), .ZN(n9589) );
  OR2_X1 U9623 ( .A1(n9773), .A2(n9774), .ZN(n9588) );
  AND2_X1 U9624 ( .A1(n8045), .A2(n9585), .ZN(n9774) );
  AND2_X1 U9625 ( .A1(n9583), .A2(n9775), .ZN(n9773) );
  OR2_X1 U9626 ( .A1(n9585), .A2(n8045), .ZN(n9775) );
  INV_X1 U9627 ( .A(n7544), .ZN(n8045) );
  AND2_X1 U9628 ( .A1(a_27_), .A2(b_27_), .ZN(n7544) );
  OR2_X1 U9629 ( .A1(n9776), .A2(n9777), .ZN(n9585) );
  AND2_X1 U9630 ( .A1(n9582), .A2(n9581), .ZN(n9777) );
  AND2_X1 U9631 ( .A1(n9579), .A2(n9778), .ZN(n9776) );
  OR2_X1 U9632 ( .A1(n9581), .A2(n9582), .ZN(n9778) );
  OR2_X1 U9633 ( .A1(n8048), .A2(n7540), .ZN(n9582) );
  OR2_X1 U9634 ( .A1(n9779), .A2(n9780), .ZN(n9581) );
  AND2_X1 U9635 ( .A1(n9575), .A2(n9781), .ZN(n9780) );
  AND2_X1 U9636 ( .A1(n9782), .A2(n9783), .ZN(n9779) );
  OR2_X1 U9637 ( .A1(n9781), .A2(n9575), .ZN(n9783) );
  OR2_X1 U9638 ( .A1(n8051), .A2(n7540), .ZN(n9575) );
  INV_X1 U9639 ( .A(n9578), .ZN(n9781) );
  AND3_X1 U9640 ( .A1(n8904), .A2(b_27_), .A3(b_26_), .ZN(n9578) );
  INV_X1 U9641 ( .A(n9577), .ZN(n9782) );
  OR2_X1 U9642 ( .A1(n9784), .A2(n9785), .ZN(n9577) );
  AND2_X1 U9643 ( .A1(b_26_), .A2(n9786), .ZN(n9785) );
  OR2_X1 U9644 ( .A1(n9787), .A2(n7490), .ZN(n9786) );
  AND2_X1 U9645 ( .A1(a_30_), .A2(n7569), .ZN(n9787) );
  AND2_X1 U9646 ( .A1(b_25_), .A2(n9788), .ZN(n9784) );
  OR2_X1 U9647 ( .A1(n9789), .A2(n7493), .ZN(n9788) );
  AND2_X1 U9648 ( .A1(a_31_), .A2(n8042), .ZN(n9789) );
  XNOR2_X1 U9649 ( .A(n9790), .B(n9791), .ZN(n9579) );
  XNOR2_X1 U9650 ( .A(n9792), .B(n9793), .ZN(n9791) );
  XOR2_X1 U9651 ( .A(n9794), .B(n9795), .Z(n9583) );
  XOR2_X1 U9652 ( .A(n9796), .B(n9797), .Z(n9795) );
  XOR2_X1 U9653 ( .A(n9798), .B(n9799), .Z(n9586) );
  XOR2_X1 U9654 ( .A(n9800), .B(n9801), .Z(n9799) );
  XOR2_X1 U9655 ( .A(n9802), .B(n9803), .Z(n9590) );
  XOR2_X1 U9656 ( .A(n9804), .B(n7560), .Z(n9803) );
  XOR2_X1 U9657 ( .A(n9805), .B(n9806), .Z(n9594) );
  XOR2_X1 U9658 ( .A(n9807), .B(n9808), .Z(n9806) );
  XOR2_X1 U9659 ( .A(n9809), .B(n9810), .Z(n9598) );
  XOR2_X1 U9660 ( .A(n9811), .B(n9812), .Z(n9810) );
  XOR2_X1 U9661 ( .A(n9813), .B(n9814), .Z(n9602) );
  XOR2_X1 U9662 ( .A(n9815), .B(n9816), .Z(n9814) );
  XOR2_X1 U9663 ( .A(n9817), .B(n9818), .Z(n9606) );
  XOR2_X1 U9664 ( .A(n9819), .B(n9820), .Z(n9818) );
  XOR2_X1 U9665 ( .A(n9821), .B(n9822), .Z(n9610) );
  XOR2_X1 U9666 ( .A(n9823), .B(n9824), .Z(n9822) );
  XOR2_X1 U9667 ( .A(n9825), .B(n9826), .Z(n9614) );
  XOR2_X1 U9668 ( .A(n9827), .B(n9828), .Z(n9826) );
  XOR2_X1 U9669 ( .A(n9829), .B(n9830), .Z(n9618) );
  XOR2_X1 U9670 ( .A(n9831), .B(n9832), .Z(n9830) );
  XOR2_X1 U9671 ( .A(n9833), .B(n9834), .Z(n9622) );
  XOR2_X1 U9672 ( .A(n9835), .B(n9836), .Z(n9834) );
  XOR2_X1 U9673 ( .A(n9837), .B(n9838), .Z(n9626) );
  XOR2_X1 U9674 ( .A(n9839), .B(n9840), .Z(n9838) );
  XOR2_X1 U9675 ( .A(n9841), .B(n9842), .Z(n9630) );
  XOR2_X1 U9676 ( .A(n9843), .B(n9844), .Z(n9842) );
  XOR2_X1 U9677 ( .A(n9845), .B(n9846), .Z(n9634) );
  XOR2_X1 U9678 ( .A(n9847), .B(n9848), .Z(n9846) );
  XOR2_X1 U9679 ( .A(n9849), .B(n9850), .Z(n9638) );
  XOR2_X1 U9680 ( .A(n9851), .B(n9852), .Z(n9850) );
  XOR2_X1 U9681 ( .A(n9853), .B(n9854), .Z(n9642) );
  XOR2_X1 U9682 ( .A(n9855), .B(n9856), .Z(n9854) );
  XOR2_X1 U9683 ( .A(n9857), .B(n9858), .Z(n9646) );
  XOR2_X1 U9684 ( .A(n9859), .B(n9860), .Z(n9858) );
  XOR2_X1 U9685 ( .A(n9861), .B(n9862), .Z(n9650) );
  XOR2_X1 U9686 ( .A(n9863), .B(n9864), .Z(n9862) );
  XOR2_X1 U9687 ( .A(n9865), .B(n9866), .Z(n9654) );
  XOR2_X1 U9688 ( .A(n9867), .B(n9868), .Z(n9866) );
  XOR2_X1 U9689 ( .A(n9869), .B(n9870), .Z(n9658) );
  XOR2_X1 U9690 ( .A(n9871), .B(n9872), .Z(n9870) );
  XOR2_X1 U9691 ( .A(n9873), .B(n9874), .Z(n9662) );
  XOR2_X1 U9692 ( .A(n9875), .B(n9876), .Z(n9874) );
  OR2_X1 U9693 ( .A1(n7970), .A2(n7540), .ZN(n9668) );
  XOR2_X1 U9694 ( .A(n9877), .B(n9878), .Z(n9667) );
  XOR2_X1 U9695 ( .A(n9879), .B(n9880), .Z(n9878) );
  XNOR2_X1 U9696 ( .A(n9881), .B(n9882), .ZN(n9670) );
  XNOR2_X1 U9697 ( .A(n9883), .B(n9884), .ZN(n9881) );
  XOR2_X1 U9698 ( .A(n9885), .B(n9886), .Z(n9674) );
  XOR2_X1 U9699 ( .A(n9887), .B(n9888), .Z(n9886) );
  XOR2_X1 U9700 ( .A(n9889), .B(n9890), .Z(n9678) );
  XOR2_X1 U9701 ( .A(n9891), .B(n9892), .Z(n9890) );
  OR2_X1 U9702 ( .A1(n7956), .A2(n7540), .ZN(n9684) );
  XOR2_X1 U9703 ( .A(n9893), .B(n9894), .Z(n9683) );
  XOR2_X1 U9704 ( .A(n9895), .B(n9896), .Z(n9894) );
  OR2_X1 U9705 ( .A1(n9686), .A2(n9689), .ZN(n9697) );
  OR2_X1 U9706 ( .A1(n7953), .A2(n7540), .ZN(n9689) );
  XOR2_X1 U9707 ( .A(n9897), .B(n9898), .Z(n9686) );
  XOR2_X1 U9708 ( .A(n9899), .B(n9900), .Z(n9898) );
  OR2_X1 U9709 ( .A1(n9473), .A2(n9476), .ZN(n9694) );
  OR2_X1 U9710 ( .A1(n7950), .A2(n7540), .ZN(n9476) );
  INV_X1 U9711 ( .A(b_27_), .ZN(n7540) );
  XOR2_X1 U9712 ( .A(n9901), .B(n9902), .Z(n9473) );
  XOR2_X1 U9713 ( .A(n9903), .B(n9904), .Z(n9902) );
  XOR2_X1 U9714 ( .A(n9905), .B(n9906), .Z(n9471) );
  XOR2_X1 U9715 ( .A(n9907), .B(n9908), .Z(n9906) );
  OR2_X1 U9716 ( .A1(n9909), .A2(n8791), .ZN(n8094) );
  XOR2_X1 U9717 ( .A(n8767), .B(n8769), .Z(n8791) );
  OR2_X1 U9718 ( .A1(n9910), .A2(n9911), .ZN(n8769) );
  AND2_X1 U9719 ( .A1(n9912), .A2(n9913), .ZN(n9911) );
  AND2_X1 U9720 ( .A1(n9914), .A2(n9915), .ZN(n9910) );
  OR2_X1 U9721 ( .A1(n9912), .A2(n9913), .ZN(n9915) );
  XOR2_X1 U9722 ( .A(n8776), .B(n9916), .Z(n8767) );
  XOR2_X1 U9723 ( .A(n8775), .B(n8774), .Z(n9916) );
  OR2_X1 U9724 ( .A1(n7950), .A2(n8035), .ZN(n8774) );
  OR2_X1 U9725 ( .A1(n9917), .A2(n9918), .ZN(n8775) );
  AND2_X1 U9726 ( .A1(n9919), .A2(n9920), .ZN(n9918) );
  AND2_X1 U9727 ( .A1(n9921), .A2(n9922), .ZN(n9917) );
  OR2_X1 U9728 ( .A1(n9919), .A2(n9920), .ZN(n9922) );
  XOR2_X1 U9729 ( .A(n8783), .B(n9923), .Z(n8776) );
  XOR2_X1 U9730 ( .A(n8782), .B(n8781), .Z(n9923) );
  OR2_X1 U9731 ( .A1(n7953), .A2(n7598), .ZN(n8781) );
  OR2_X1 U9732 ( .A1(n9924), .A2(n9925), .ZN(n8782) );
  AND2_X1 U9733 ( .A1(n9926), .A2(n9927), .ZN(n9925) );
  AND2_X1 U9734 ( .A1(n9928), .A2(n9929), .ZN(n9924) );
  OR2_X1 U9735 ( .A1(n9926), .A2(n9927), .ZN(n9929) );
  XOR2_X1 U9736 ( .A(n9930), .B(n9931), .Z(n8783) );
  XOR2_X1 U9737 ( .A(n9932), .B(n9933), .Z(n9931) );
  AND2_X1 U9738 ( .A1(n8792), .A2(n8790), .ZN(n9909) );
  XNOR2_X1 U9739 ( .A(n9914), .B(n9934), .ZN(n8790) );
  XOR2_X1 U9740 ( .A(n9913), .B(n9912), .Z(n9934) );
  OR2_X1 U9741 ( .A1(n7950), .A2(n7569), .ZN(n9912) );
  OR2_X1 U9742 ( .A1(n9935), .A2(n9936), .ZN(n9913) );
  AND2_X1 U9743 ( .A1(n9937), .A2(n9938), .ZN(n9936) );
  AND2_X1 U9744 ( .A1(n9939), .A2(n9940), .ZN(n9935) );
  OR2_X1 U9745 ( .A1(n9937), .A2(n9938), .ZN(n9940) );
  XNOR2_X1 U9746 ( .A(n9941), .B(n9921), .ZN(n9914) );
  XOR2_X1 U9747 ( .A(n9928), .B(n9942), .Z(n9921) );
  XOR2_X1 U9748 ( .A(n9927), .B(n9926), .Z(n9942) );
  OR2_X1 U9749 ( .A1(n7956), .A2(n7598), .ZN(n9926) );
  OR2_X1 U9750 ( .A1(n9943), .A2(n9944), .ZN(n9927) );
  AND2_X1 U9751 ( .A1(n9945), .A2(n9946), .ZN(n9944) );
  AND2_X1 U9752 ( .A1(n9947), .A2(n9948), .ZN(n9943) );
  OR2_X1 U9753 ( .A1(n9945), .A2(n9946), .ZN(n9948) );
  XOR2_X1 U9754 ( .A(n9949), .B(n9950), .Z(n9928) );
  XOR2_X1 U9755 ( .A(n9951), .B(n9952), .Z(n9950) );
  XNOR2_X1 U9756 ( .A(n9920), .B(n9919), .ZN(n9941) );
  OR2_X1 U9757 ( .A1(n9953), .A2(n9954), .ZN(n9919) );
  AND2_X1 U9758 ( .A1(n9955), .A2(n9956), .ZN(n9954) );
  AND2_X1 U9759 ( .A1(n9957), .A2(n9958), .ZN(n9953) );
  OR2_X1 U9760 ( .A1(n9955), .A2(n9956), .ZN(n9958) );
  OR2_X1 U9761 ( .A1(n7953), .A2(n8035), .ZN(n9920) );
  INV_X1 U9762 ( .A(n9690), .ZN(n8792) );
  OR2_X1 U9763 ( .A1(n9959), .A2(n9960), .ZN(n9690) );
  AND2_X1 U9764 ( .A1(n9908), .A2(n9907), .ZN(n9960) );
  AND2_X1 U9765 ( .A1(n9905), .A2(n9961), .ZN(n9959) );
  OR2_X1 U9766 ( .A1(n9907), .A2(n9908), .ZN(n9961) );
  OR2_X1 U9767 ( .A1(n7950), .A2(n8042), .ZN(n9908) );
  OR2_X1 U9768 ( .A1(n9962), .A2(n9963), .ZN(n9907) );
  AND2_X1 U9769 ( .A1(n9904), .A2(n9903), .ZN(n9963) );
  AND2_X1 U9770 ( .A1(n9901), .A2(n9964), .ZN(n9962) );
  OR2_X1 U9771 ( .A1(n9903), .A2(n9904), .ZN(n9964) );
  OR2_X1 U9772 ( .A1(n7953), .A2(n8042), .ZN(n9904) );
  OR2_X1 U9773 ( .A1(n9965), .A2(n9966), .ZN(n9903) );
  AND2_X1 U9774 ( .A1(n9900), .A2(n9899), .ZN(n9966) );
  AND2_X1 U9775 ( .A1(n9897), .A2(n9967), .ZN(n9965) );
  OR2_X1 U9776 ( .A1(n9899), .A2(n9900), .ZN(n9967) );
  OR2_X1 U9777 ( .A1(n7956), .A2(n8042), .ZN(n9900) );
  OR2_X1 U9778 ( .A1(n9968), .A2(n9969), .ZN(n9899) );
  AND2_X1 U9779 ( .A1(n9896), .A2(n9895), .ZN(n9969) );
  AND2_X1 U9780 ( .A1(n9893), .A2(n9970), .ZN(n9968) );
  OR2_X1 U9781 ( .A1(n9895), .A2(n9896), .ZN(n9970) );
  OR2_X1 U9782 ( .A1(n7960), .A2(n8042), .ZN(n9896) );
  OR2_X1 U9783 ( .A1(n9971), .A2(n9972), .ZN(n9895) );
  AND2_X1 U9784 ( .A1(n9892), .A2(n9891), .ZN(n9972) );
  AND2_X1 U9785 ( .A1(n9889), .A2(n9973), .ZN(n9971) );
  OR2_X1 U9786 ( .A1(n9891), .A2(n9892), .ZN(n9973) );
  OR2_X1 U9787 ( .A1(n7963), .A2(n8042), .ZN(n9892) );
  OR2_X1 U9788 ( .A1(n9974), .A2(n9975), .ZN(n9891) );
  AND2_X1 U9789 ( .A1(n9888), .A2(n9887), .ZN(n9975) );
  AND2_X1 U9790 ( .A1(n9885), .A2(n9976), .ZN(n9974) );
  OR2_X1 U9791 ( .A1(n9887), .A2(n9888), .ZN(n9976) );
  OR2_X1 U9792 ( .A1(n7967), .A2(n8042), .ZN(n9888) );
  OR2_X1 U9793 ( .A1(n9977), .A2(n9978), .ZN(n9887) );
  AND2_X1 U9794 ( .A1(n9884), .A2(n9883), .ZN(n9978) );
  AND2_X1 U9795 ( .A1(n9882), .A2(n9979), .ZN(n9977) );
  OR2_X1 U9796 ( .A1(n9883), .A2(n9884), .ZN(n9979) );
  OR2_X1 U9797 ( .A1(n9980), .A2(n9981), .ZN(n9884) );
  AND2_X1 U9798 ( .A1(n9880), .A2(n9879), .ZN(n9981) );
  AND2_X1 U9799 ( .A1(n9877), .A2(n9982), .ZN(n9980) );
  OR2_X1 U9800 ( .A1(n9879), .A2(n9880), .ZN(n9982) );
  OR2_X1 U9801 ( .A1(n7974), .A2(n8042), .ZN(n9880) );
  OR2_X1 U9802 ( .A1(n9983), .A2(n9984), .ZN(n9879) );
  AND2_X1 U9803 ( .A1(n9876), .A2(n9875), .ZN(n9984) );
  AND2_X1 U9804 ( .A1(n9873), .A2(n9985), .ZN(n9983) );
  OR2_X1 U9805 ( .A1(n9875), .A2(n9876), .ZN(n9985) );
  OR2_X1 U9806 ( .A1(n7977), .A2(n8042), .ZN(n9876) );
  OR2_X1 U9807 ( .A1(n9986), .A2(n9987), .ZN(n9875) );
  AND2_X1 U9808 ( .A1(n9872), .A2(n9871), .ZN(n9987) );
  AND2_X1 U9809 ( .A1(n9869), .A2(n9988), .ZN(n9986) );
  OR2_X1 U9810 ( .A1(n9871), .A2(n9872), .ZN(n9988) );
  OR2_X1 U9811 ( .A1(n7981), .A2(n8042), .ZN(n9872) );
  OR2_X1 U9812 ( .A1(n9989), .A2(n9990), .ZN(n9871) );
  AND2_X1 U9813 ( .A1(n9868), .A2(n9867), .ZN(n9990) );
  AND2_X1 U9814 ( .A1(n9865), .A2(n9991), .ZN(n9989) );
  OR2_X1 U9815 ( .A1(n9867), .A2(n9868), .ZN(n9991) );
  OR2_X1 U9816 ( .A1(n7984), .A2(n8042), .ZN(n9868) );
  OR2_X1 U9817 ( .A1(n9992), .A2(n9993), .ZN(n9867) );
  AND2_X1 U9818 ( .A1(n9864), .A2(n9863), .ZN(n9993) );
  AND2_X1 U9819 ( .A1(n9861), .A2(n9994), .ZN(n9992) );
  OR2_X1 U9820 ( .A1(n9863), .A2(n9864), .ZN(n9994) );
  OR2_X1 U9821 ( .A1(n7988), .A2(n8042), .ZN(n9864) );
  OR2_X1 U9822 ( .A1(n9995), .A2(n9996), .ZN(n9863) );
  AND2_X1 U9823 ( .A1(n9860), .A2(n9859), .ZN(n9996) );
  AND2_X1 U9824 ( .A1(n9857), .A2(n9997), .ZN(n9995) );
  OR2_X1 U9825 ( .A1(n9859), .A2(n9860), .ZN(n9997) );
  OR2_X1 U9826 ( .A1(n7991), .A2(n8042), .ZN(n9860) );
  OR2_X1 U9827 ( .A1(n9998), .A2(n9999), .ZN(n9859) );
  AND2_X1 U9828 ( .A1(n9856), .A2(n9855), .ZN(n9999) );
  AND2_X1 U9829 ( .A1(n9853), .A2(n10000), .ZN(n9998) );
  OR2_X1 U9830 ( .A1(n9855), .A2(n9856), .ZN(n10000) );
  OR2_X1 U9831 ( .A1(n7995), .A2(n8042), .ZN(n9856) );
  OR2_X1 U9832 ( .A1(n10001), .A2(n10002), .ZN(n9855) );
  AND2_X1 U9833 ( .A1(n9852), .A2(n9851), .ZN(n10002) );
  AND2_X1 U9834 ( .A1(n9849), .A2(n10003), .ZN(n10001) );
  OR2_X1 U9835 ( .A1(n9851), .A2(n9852), .ZN(n10003) );
  OR2_X1 U9836 ( .A1(n7998), .A2(n8042), .ZN(n9852) );
  OR2_X1 U9837 ( .A1(n10004), .A2(n10005), .ZN(n9851) );
  AND2_X1 U9838 ( .A1(n9848), .A2(n9847), .ZN(n10005) );
  AND2_X1 U9839 ( .A1(n9845), .A2(n10006), .ZN(n10004) );
  OR2_X1 U9840 ( .A1(n9847), .A2(n9848), .ZN(n10006) );
  OR2_X1 U9841 ( .A1(n8002), .A2(n8042), .ZN(n9848) );
  OR2_X1 U9842 ( .A1(n10007), .A2(n10008), .ZN(n9847) );
  AND2_X1 U9843 ( .A1(n9844), .A2(n9843), .ZN(n10008) );
  AND2_X1 U9844 ( .A1(n9841), .A2(n10009), .ZN(n10007) );
  OR2_X1 U9845 ( .A1(n9843), .A2(n9844), .ZN(n10009) );
  OR2_X1 U9846 ( .A1(n8005), .A2(n8042), .ZN(n9844) );
  OR2_X1 U9847 ( .A1(n10010), .A2(n10011), .ZN(n9843) );
  AND2_X1 U9848 ( .A1(n9840), .A2(n9839), .ZN(n10011) );
  AND2_X1 U9849 ( .A1(n9837), .A2(n10012), .ZN(n10010) );
  OR2_X1 U9850 ( .A1(n9839), .A2(n9840), .ZN(n10012) );
  OR2_X1 U9851 ( .A1(n8009), .A2(n8042), .ZN(n9840) );
  OR2_X1 U9852 ( .A1(n10013), .A2(n10014), .ZN(n9839) );
  AND2_X1 U9853 ( .A1(n9836), .A2(n9835), .ZN(n10014) );
  AND2_X1 U9854 ( .A1(n9833), .A2(n10015), .ZN(n10013) );
  OR2_X1 U9855 ( .A1(n9835), .A2(n9836), .ZN(n10015) );
  OR2_X1 U9856 ( .A1(n8012), .A2(n8042), .ZN(n9836) );
  OR2_X1 U9857 ( .A1(n10016), .A2(n10017), .ZN(n9835) );
  AND2_X1 U9858 ( .A1(n9832), .A2(n9831), .ZN(n10017) );
  AND2_X1 U9859 ( .A1(n9829), .A2(n10018), .ZN(n10016) );
  OR2_X1 U9860 ( .A1(n9831), .A2(n9832), .ZN(n10018) );
  OR2_X1 U9861 ( .A1(n8016), .A2(n8042), .ZN(n9832) );
  OR2_X1 U9862 ( .A1(n10019), .A2(n10020), .ZN(n9831) );
  AND2_X1 U9863 ( .A1(n9828), .A2(n9827), .ZN(n10020) );
  AND2_X1 U9864 ( .A1(n9825), .A2(n10021), .ZN(n10019) );
  OR2_X1 U9865 ( .A1(n9827), .A2(n9828), .ZN(n10021) );
  OR2_X1 U9866 ( .A1(n8019), .A2(n8042), .ZN(n9828) );
  OR2_X1 U9867 ( .A1(n10022), .A2(n10023), .ZN(n9827) );
  AND2_X1 U9868 ( .A1(n9824), .A2(n9823), .ZN(n10023) );
  AND2_X1 U9869 ( .A1(n9821), .A2(n10024), .ZN(n10022) );
  OR2_X1 U9870 ( .A1(n9823), .A2(n9824), .ZN(n10024) );
  OR2_X1 U9871 ( .A1(n8023), .A2(n8042), .ZN(n9824) );
  OR2_X1 U9872 ( .A1(n10025), .A2(n10026), .ZN(n9823) );
  AND2_X1 U9873 ( .A1(n9820), .A2(n9819), .ZN(n10026) );
  AND2_X1 U9874 ( .A1(n9817), .A2(n10027), .ZN(n10025) );
  OR2_X1 U9875 ( .A1(n9819), .A2(n9820), .ZN(n10027) );
  OR2_X1 U9876 ( .A1(n8026), .A2(n8042), .ZN(n9820) );
  OR2_X1 U9877 ( .A1(n10028), .A2(n10029), .ZN(n9819) );
  AND2_X1 U9878 ( .A1(n9816), .A2(n9815), .ZN(n10029) );
  AND2_X1 U9879 ( .A1(n9813), .A2(n10030), .ZN(n10028) );
  OR2_X1 U9880 ( .A1(n9815), .A2(n9816), .ZN(n10030) );
  OR2_X1 U9881 ( .A1(n8030), .A2(n8042), .ZN(n9816) );
  OR2_X1 U9882 ( .A1(n10031), .A2(n10032), .ZN(n9815) );
  AND2_X1 U9883 ( .A1(n9812), .A2(n9811), .ZN(n10032) );
  AND2_X1 U9884 ( .A1(n9809), .A2(n10033), .ZN(n10031) );
  OR2_X1 U9885 ( .A1(n9811), .A2(n9812), .ZN(n10033) );
  OR2_X1 U9886 ( .A1(n8034), .A2(n8042), .ZN(n9812) );
  OR2_X1 U9887 ( .A1(n10034), .A2(n10035), .ZN(n9811) );
  AND2_X1 U9888 ( .A1(n9808), .A2(n9807), .ZN(n10035) );
  AND2_X1 U9889 ( .A1(n9805), .A2(n10036), .ZN(n10034) );
  OR2_X1 U9890 ( .A1(n9807), .A2(n9808), .ZN(n10036) );
  OR2_X1 U9891 ( .A1(n8037), .A2(n8042), .ZN(n9808) );
  OR2_X1 U9892 ( .A1(n10037), .A2(n10038), .ZN(n9807) );
  AND2_X1 U9893 ( .A1(n7560), .A2(n9804), .ZN(n10038) );
  AND2_X1 U9894 ( .A1(n9802), .A2(n10039), .ZN(n10037) );
  OR2_X1 U9895 ( .A1(n9804), .A2(n7560), .ZN(n10039) );
  OR2_X1 U9896 ( .A1(n8041), .A2(n8042), .ZN(n7560) );
  OR2_X1 U9897 ( .A1(n10040), .A2(n10041), .ZN(n9804) );
  AND2_X1 U9898 ( .A1(n9801), .A2(n9800), .ZN(n10041) );
  AND2_X1 U9899 ( .A1(n9798), .A2(n10042), .ZN(n10040) );
  OR2_X1 U9900 ( .A1(n9800), .A2(n9801), .ZN(n10042) );
  OR2_X1 U9901 ( .A1(n8044), .A2(n8042), .ZN(n9801) );
  OR2_X1 U9902 ( .A1(n10043), .A2(n10044), .ZN(n9800) );
  AND2_X1 U9903 ( .A1(n9797), .A2(n9796), .ZN(n10044) );
  AND2_X1 U9904 ( .A1(n9794), .A2(n10045), .ZN(n10043) );
  OR2_X1 U9905 ( .A1(n9796), .A2(n9797), .ZN(n10045) );
  OR2_X1 U9906 ( .A1(n8048), .A2(n8042), .ZN(n9797) );
  OR2_X1 U9907 ( .A1(n10046), .A2(n10047), .ZN(n9796) );
  AND2_X1 U9908 ( .A1(n9790), .A2(n10048), .ZN(n10047) );
  AND2_X1 U9909 ( .A1(n10049), .A2(n10050), .ZN(n10046) );
  OR2_X1 U9910 ( .A1(n10048), .A2(n9790), .ZN(n10050) );
  OR2_X1 U9911 ( .A1(n8051), .A2(n8042), .ZN(n9790) );
  INV_X1 U9912 ( .A(n9793), .ZN(n10048) );
  AND3_X1 U9913 ( .A1(n8904), .A2(b_25_), .A3(b_26_), .ZN(n9793) );
  INV_X1 U9914 ( .A(n9792), .ZN(n10049) );
  OR2_X1 U9915 ( .A1(n10051), .A2(n10052), .ZN(n9792) );
  AND2_X1 U9916 ( .A1(b_25_), .A2(n10053), .ZN(n10052) );
  OR2_X1 U9917 ( .A1(n10054), .A2(n7490), .ZN(n10053) );
  AND2_X1 U9918 ( .A1(a_30_), .A2(n8035), .ZN(n10054) );
  AND2_X1 U9919 ( .A1(b_24_), .A2(n10055), .ZN(n10051) );
  OR2_X1 U9920 ( .A1(n10056), .A2(n7493), .ZN(n10055) );
  AND2_X1 U9921 ( .A1(a_31_), .A2(n7569), .ZN(n10056) );
  XNOR2_X1 U9922 ( .A(n10057), .B(n10058), .ZN(n9794) );
  XNOR2_X1 U9923 ( .A(n10059), .B(n10060), .ZN(n10058) );
  XOR2_X1 U9924 ( .A(n10061), .B(n10062), .Z(n9798) );
  XOR2_X1 U9925 ( .A(n10063), .B(n10064), .Z(n10062) );
  XOR2_X1 U9926 ( .A(n10065), .B(n10066), .Z(n9802) );
  XOR2_X1 U9927 ( .A(n10067), .B(n10068), .Z(n10066) );
  XOR2_X1 U9928 ( .A(n10069), .B(n10070), .Z(n9805) );
  XOR2_X1 U9929 ( .A(n10071), .B(n10072), .Z(n10070) );
  XOR2_X1 U9930 ( .A(n10073), .B(n10074), .Z(n9809) );
  XNOR2_X1 U9931 ( .A(n10075), .B(n7573), .ZN(n10074) );
  XOR2_X1 U9932 ( .A(n10076), .B(n10077), .Z(n9813) );
  XOR2_X1 U9933 ( .A(n10078), .B(n10079), .Z(n10077) );
  XOR2_X1 U9934 ( .A(n10080), .B(n10081), .Z(n9817) );
  XOR2_X1 U9935 ( .A(n10082), .B(n10083), .Z(n10081) );
  XOR2_X1 U9936 ( .A(n10084), .B(n10085), .Z(n9821) );
  XOR2_X1 U9937 ( .A(n10086), .B(n10087), .Z(n10085) );
  XOR2_X1 U9938 ( .A(n10088), .B(n10089), .Z(n9825) );
  XOR2_X1 U9939 ( .A(n10090), .B(n10091), .Z(n10089) );
  XOR2_X1 U9940 ( .A(n10092), .B(n10093), .Z(n9829) );
  XOR2_X1 U9941 ( .A(n10094), .B(n10095), .Z(n10093) );
  XOR2_X1 U9942 ( .A(n10096), .B(n10097), .Z(n9833) );
  XOR2_X1 U9943 ( .A(n10098), .B(n10099), .Z(n10097) );
  XOR2_X1 U9944 ( .A(n10100), .B(n10101), .Z(n9837) );
  XOR2_X1 U9945 ( .A(n10102), .B(n10103), .Z(n10101) );
  XOR2_X1 U9946 ( .A(n10104), .B(n10105), .Z(n9841) );
  XOR2_X1 U9947 ( .A(n10106), .B(n10107), .Z(n10105) );
  XOR2_X1 U9948 ( .A(n10108), .B(n10109), .Z(n9845) );
  XOR2_X1 U9949 ( .A(n10110), .B(n10111), .Z(n10109) );
  XOR2_X1 U9950 ( .A(n10112), .B(n10113), .Z(n9849) );
  XOR2_X1 U9951 ( .A(n10114), .B(n10115), .Z(n10113) );
  XOR2_X1 U9952 ( .A(n10116), .B(n10117), .Z(n9853) );
  XOR2_X1 U9953 ( .A(n10118), .B(n10119), .Z(n10117) );
  XOR2_X1 U9954 ( .A(n10120), .B(n10121), .Z(n9857) );
  XOR2_X1 U9955 ( .A(n10122), .B(n10123), .Z(n10121) );
  XOR2_X1 U9956 ( .A(n10124), .B(n10125), .Z(n9861) );
  XOR2_X1 U9957 ( .A(n10126), .B(n10127), .Z(n10125) );
  XOR2_X1 U9958 ( .A(n10128), .B(n10129), .Z(n9865) );
  XOR2_X1 U9959 ( .A(n10130), .B(n10131), .Z(n10129) );
  XNOR2_X1 U9960 ( .A(n10132), .B(n10133), .ZN(n9869) );
  XNOR2_X1 U9961 ( .A(n10134), .B(n10135), .ZN(n10132) );
  XOR2_X1 U9962 ( .A(n10136), .B(n10137), .Z(n9873) );
  XOR2_X1 U9963 ( .A(n10138), .B(n10139), .Z(n10137) );
  XOR2_X1 U9964 ( .A(n10140), .B(n10141), .Z(n9877) );
  XOR2_X1 U9965 ( .A(n10142), .B(n10143), .Z(n10141) );
  OR2_X1 U9966 ( .A1(n7970), .A2(n8042), .ZN(n9883) );
  INV_X1 U9967 ( .A(b_26_), .ZN(n8042) );
  XOR2_X1 U9968 ( .A(n10144), .B(n10145), .Z(n9882) );
  XOR2_X1 U9969 ( .A(n10146), .B(n10147), .Z(n10145) );
  XNOR2_X1 U9970 ( .A(n10148), .B(n10149), .ZN(n9885) );
  XNOR2_X1 U9971 ( .A(n10150), .B(n10151), .ZN(n10148) );
  XOR2_X1 U9972 ( .A(n10152), .B(n10153), .Z(n9889) );
  XOR2_X1 U9973 ( .A(n10154), .B(n10155), .Z(n10153) );
  XOR2_X1 U9974 ( .A(n10156), .B(n10157), .Z(n9893) );
  XOR2_X1 U9975 ( .A(n10158), .B(n10159), .Z(n10157) );
  XOR2_X1 U9976 ( .A(n10160), .B(n10161), .Z(n9897) );
  XOR2_X1 U9977 ( .A(n10162), .B(n10163), .Z(n10161) );
  XOR2_X1 U9978 ( .A(n10164), .B(n10165), .Z(n9901) );
  XOR2_X1 U9979 ( .A(n10166), .B(n10167), .Z(n10165) );
  XOR2_X1 U9980 ( .A(n9939), .B(n10168), .Z(n9905) );
  XOR2_X1 U9981 ( .A(n9938), .B(n9937), .Z(n10168) );
  OR2_X1 U9982 ( .A1(n7953), .A2(n7569), .ZN(n9937) );
  OR2_X1 U9983 ( .A1(n10169), .A2(n10170), .ZN(n9938) );
  AND2_X1 U9984 ( .A1(n10167), .A2(n10166), .ZN(n10170) );
  AND2_X1 U9985 ( .A1(n10164), .A2(n10171), .ZN(n10169) );
  OR2_X1 U9986 ( .A1(n10167), .A2(n10166), .ZN(n10171) );
  OR2_X1 U9987 ( .A1(n10172), .A2(n10173), .ZN(n10166) );
  AND2_X1 U9988 ( .A1(n10163), .A2(n10162), .ZN(n10173) );
  AND2_X1 U9989 ( .A1(n10160), .A2(n10174), .ZN(n10172) );
  OR2_X1 U9990 ( .A1(n10163), .A2(n10162), .ZN(n10174) );
  OR2_X1 U9991 ( .A1(n10175), .A2(n10176), .ZN(n10162) );
  AND2_X1 U9992 ( .A1(n10159), .A2(n10158), .ZN(n10176) );
  AND2_X1 U9993 ( .A1(n10156), .A2(n10177), .ZN(n10175) );
  OR2_X1 U9994 ( .A1(n10159), .A2(n10158), .ZN(n10177) );
  OR2_X1 U9995 ( .A1(n10178), .A2(n10179), .ZN(n10158) );
  AND2_X1 U9996 ( .A1(n10155), .A2(n10154), .ZN(n10179) );
  AND2_X1 U9997 ( .A1(n10152), .A2(n10180), .ZN(n10178) );
  OR2_X1 U9998 ( .A1(n10155), .A2(n10154), .ZN(n10180) );
  OR2_X1 U9999 ( .A1(n10181), .A2(n10182), .ZN(n10154) );
  AND2_X1 U10000 ( .A1(n10151), .A2(n10150), .ZN(n10182) );
  AND2_X1 U10001 ( .A1(n10149), .A2(n10183), .ZN(n10181) );
  OR2_X1 U10002 ( .A1(n10151), .A2(n10150), .ZN(n10183) );
  OR2_X1 U10003 ( .A1(n7970), .A2(n7569), .ZN(n10150) );
  OR2_X1 U10004 ( .A1(n10184), .A2(n10185), .ZN(n10151) );
  AND2_X1 U10005 ( .A1(n10147), .A2(n10146), .ZN(n10185) );
  AND2_X1 U10006 ( .A1(n10144), .A2(n10186), .ZN(n10184) );
  OR2_X1 U10007 ( .A1(n10147), .A2(n10146), .ZN(n10186) );
  OR2_X1 U10008 ( .A1(n10187), .A2(n10188), .ZN(n10146) );
  AND2_X1 U10009 ( .A1(n10143), .A2(n10142), .ZN(n10188) );
  AND2_X1 U10010 ( .A1(n10140), .A2(n10189), .ZN(n10187) );
  OR2_X1 U10011 ( .A1(n10143), .A2(n10142), .ZN(n10189) );
  OR2_X1 U10012 ( .A1(n10190), .A2(n10191), .ZN(n10142) );
  AND2_X1 U10013 ( .A1(n10139), .A2(n10138), .ZN(n10191) );
  AND2_X1 U10014 ( .A1(n10136), .A2(n10192), .ZN(n10190) );
  OR2_X1 U10015 ( .A1(n10139), .A2(n10138), .ZN(n10192) );
  OR2_X1 U10016 ( .A1(n10193), .A2(n10194), .ZN(n10138) );
  AND2_X1 U10017 ( .A1(n10135), .A2(n10134), .ZN(n10194) );
  AND2_X1 U10018 ( .A1(n10133), .A2(n10195), .ZN(n10193) );
  OR2_X1 U10019 ( .A1(n10135), .A2(n10134), .ZN(n10195) );
  OR2_X1 U10020 ( .A1(n7984), .A2(n7569), .ZN(n10134) );
  OR2_X1 U10021 ( .A1(n10196), .A2(n10197), .ZN(n10135) );
  AND2_X1 U10022 ( .A1(n10131), .A2(n10130), .ZN(n10197) );
  AND2_X1 U10023 ( .A1(n10128), .A2(n10198), .ZN(n10196) );
  OR2_X1 U10024 ( .A1(n10131), .A2(n10130), .ZN(n10198) );
  OR2_X1 U10025 ( .A1(n10199), .A2(n10200), .ZN(n10130) );
  AND2_X1 U10026 ( .A1(n10127), .A2(n10126), .ZN(n10200) );
  AND2_X1 U10027 ( .A1(n10124), .A2(n10201), .ZN(n10199) );
  OR2_X1 U10028 ( .A1(n10127), .A2(n10126), .ZN(n10201) );
  OR2_X1 U10029 ( .A1(n10202), .A2(n10203), .ZN(n10126) );
  AND2_X1 U10030 ( .A1(n10123), .A2(n10122), .ZN(n10203) );
  AND2_X1 U10031 ( .A1(n10120), .A2(n10204), .ZN(n10202) );
  OR2_X1 U10032 ( .A1(n10123), .A2(n10122), .ZN(n10204) );
  OR2_X1 U10033 ( .A1(n10205), .A2(n10206), .ZN(n10122) );
  AND2_X1 U10034 ( .A1(n10119), .A2(n10118), .ZN(n10206) );
  AND2_X1 U10035 ( .A1(n10116), .A2(n10207), .ZN(n10205) );
  OR2_X1 U10036 ( .A1(n10119), .A2(n10118), .ZN(n10207) );
  OR2_X1 U10037 ( .A1(n10208), .A2(n10209), .ZN(n10118) );
  AND2_X1 U10038 ( .A1(n10115), .A2(n10114), .ZN(n10209) );
  AND2_X1 U10039 ( .A1(n10112), .A2(n10210), .ZN(n10208) );
  OR2_X1 U10040 ( .A1(n10115), .A2(n10114), .ZN(n10210) );
  OR2_X1 U10041 ( .A1(n10211), .A2(n10212), .ZN(n10114) );
  AND2_X1 U10042 ( .A1(n10111), .A2(n10110), .ZN(n10212) );
  AND2_X1 U10043 ( .A1(n10108), .A2(n10213), .ZN(n10211) );
  OR2_X1 U10044 ( .A1(n10111), .A2(n10110), .ZN(n10213) );
  OR2_X1 U10045 ( .A1(n10214), .A2(n10215), .ZN(n10110) );
  AND2_X1 U10046 ( .A1(n10107), .A2(n10106), .ZN(n10215) );
  AND2_X1 U10047 ( .A1(n10104), .A2(n10216), .ZN(n10214) );
  OR2_X1 U10048 ( .A1(n10107), .A2(n10106), .ZN(n10216) );
  OR2_X1 U10049 ( .A1(n10217), .A2(n10218), .ZN(n10106) );
  AND2_X1 U10050 ( .A1(n10103), .A2(n10102), .ZN(n10218) );
  AND2_X1 U10051 ( .A1(n10100), .A2(n10219), .ZN(n10217) );
  OR2_X1 U10052 ( .A1(n10103), .A2(n10102), .ZN(n10219) );
  OR2_X1 U10053 ( .A1(n10220), .A2(n10221), .ZN(n10102) );
  AND2_X1 U10054 ( .A1(n10099), .A2(n10098), .ZN(n10221) );
  AND2_X1 U10055 ( .A1(n10096), .A2(n10222), .ZN(n10220) );
  OR2_X1 U10056 ( .A1(n10099), .A2(n10098), .ZN(n10222) );
  OR2_X1 U10057 ( .A1(n10223), .A2(n10224), .ZN(n10098) );
  AND2_X1 U10058 ( .A1(n10095), .A2(n10094), .ZN(n10224) );
  AND2_X1 U10059 ( .A1(n10092), .A2(n10225), .ZN(n10223) );
  OR2_X1 U10060 ( .A1(n10095), .A2(n10094), .ZN(n10225) );
  OR2_X1 U10061 ( .A1(n10226), .A2(n10227), .ZN(n10094) );
  AND2_X1 U10062 ( .A1(n10091), .A2(n10090), .ZN(n10227) );
  AND2_X1 U10063 ( .A1(n10088), .A2(n10228), .ZN(n10226) );
  OR2_X1 U10064 ( .A1(n10091), .A2(n10090), .ZN(n10228) );
  OR2_X1 U10065 ( .A1(n10229), .A2(n10230), .ZN(n10090) );
  AND2_X1 U10066 ( .A1(n10087), .A2(n10086), .ZN(n10230) );
  AND2_X1 U10067 ( .A1(n10084), .A2(n10231), .ZN(n10229) );
  OR2_X1 U10068 ( .A1(n10087), .A2(n10086), .ZN(n10231) );
  OR2_X1 U10069 ( .A1(n10232), .A2(n10233), .ZN(n10086) );
  AND2_X1 U10070 ( .A1(n10083), .A2(n10082), .ZN(n10233) );
  AND2_X1 U10071 ( .A1(n10080), .A2(n10234), .ZN(n10232) );
  OR2_X1 U10072 ( .A1(n10083), .A2(n10082), .ZN(n10234) );
  OR2_X1 U10073 ( .A1(n10235), .A2(n10236), .ZN(n10082) );
  AND2_X1 U10074 ( .A1(n10079), .A2(n10078), .ZN(n10236) );
  AND2_X1 U10075 ( .A1(n10076), .A2(n10237), .ZN(n10235) );
  OR2_X1 U10076 ( .A1(n10079), .A2(n10078), .ZN(n10237) );
  OR2_X1 U10077 ( .A1(n10238), .A2(n10239), .ZN(n10078) );
  AND2_X1 U10078 ( .A1(n8038), .A2(n10075), .ZN(n10239) );
  AND2_X1 U10079 ( .A1(n10073), .A2(n10240), .ZN(n10238) );
  OR2_X1 U10080 ( .A1(n8038), .A2(n10075), .ZN(n10240) );
  OR2_X1 U10081 ( .A1(n10241), .A2(n10242), .ZN(n10075) );
  AND2_X1 U10082 ( .A1(n10072), .A2(n10071), .ZN(n10242) );
  AND2_X1 U10083 ( .A1(n10069), .A2(n10243), .ZN(n10241) );
  OR2_X1 U10084 ( .A1(n10072), .A2(n10071), .ZN(n10243) );
  OR2_X1 U10085 ( .A1(n10244), .A2(n10245), .ZN(n10071) );
  AND2_X1 U10086 ( .A1(n10068), .A2(n10067), .ZN(n10245) );
  AND2_X1 U10087 ( .A1(n10065), .A2(n10246), .ZN(n10244) );
  OR2_X1 U10088 ( .A1(n10068), .A2(n10067), .ZN(n10246) );
  OR2_X1 U10089 ( .A1(n10247), .A2(n10248), .ZN(n10067) );
  AND2_X1 U10090 ( .A1(n10064), .A2(n10063), .ZN(n10248) );
  AND2_X1 U10091 ( .A1(n10061), .A2(n10249), .ZN(n10247) );
  OR2_X1 U10092 ( .A1(n10064), .A2(n10063), .ZN(n10249) );
  OR2_X1 U10093 ( .A1(n10250), .A2(n10251), .ZN(n10063) );
  AND2_X1 U10094 ( .A1(n10057), .A2(n10252), .ZN(n10251) );
  AND2_X1 U10095 ( .A1(n10253), .A2(n10254), .ZN(n10250) );
  OR2_X1 U10096 ( .A1(n10057), .A2(n10252), .ZN(n10254) );
  INV_X1 U10097 ( .A(n10060), .ZN(n10252) );
  AND3_X1 U10098 ( .A1(n8904), .A2(b_24_), .A3(b_25_), .ZN(n10060) );
  OR2_X1 U10099 ( .A1(n8051), .A2(n7569), .ZN(n10057) );
  INV_X1 U10100 ( .A(n10059), .ZN(n10253) );
  OR2_X1 U10101 ( .A1(n10255), .A2(n10256), .ZN(n10059) );
  AND2_X1 U10102 ( .A1(b_24_), .A2(n10257), .ZN(n10256) );
  OR2_X1 U10103 ( .A1(n10258), .A2(n7490), .ZN(n10257) );
  AND2_X1 U10104 ( .A1(a_30_), .A2(n7598), .ZN(n10258) );
  AND2_X1 U10105 ( .A1(b_23_), .A2(n10259), .ZN(n10255) );
  OR2_X1 U10106 ( .A1(n10260), .A2(n7493), .ZN(n10259) );
  AND2_X1 U10107 ( .A1(a_31_), .A2(n8035), .ZN(n10260) );
  OR2_X1 U10108 ( .A1(n8048), .A2(n7569), .ZN(n10064) );
  XNOR2_X1 U10109 ( .A(n10261), .B(n10262), .ZN(n10061) );
  XNOR2_X1 U10110 ( .A(n10263), .B(n10264), .ZN(n10262) );
  OR2_X1 U10111 ( .A1(n8044), .A2(n7569), .ZN(n10068) );
  XOR2_X1 U10112 ( .A(n10265), .B(n10266), .Z(n10065) );
  XOR2_X1 U10113 ( .A(n10267), .B(n10268), .Z(n10266) );
  OR2_X1 U10114 ( .A1(n8041), .A2(n7569), .ZN(n10072) );
  XOR2_X1 U10115 ( .A(n10269), .B(n10270), .Z(n10069) );
  XOR2_X1 U10116 ( .A(n10271), .B(n10272), .Z(n10270) );
  INV_X1 U10117 ( .A(n7573), .ZN(n8038) );
  AND2_X1 U10118 ( .A1(a_25_), .A2(b_25_), .ZN(n7573) );
  XOR2_X1 U10119 ( .A(n10273), .B(n10274), .Z(n10073) );
  XOR2_X1 U10120 ( .A(n10275), .B(n10276), .Z(n10274) );
  OR2_X1 U10121 ( .A1(n8034), .A2(n7569), .ZN(n10079) );
  XOR2_X1 U10122 ( .A(n10277), .B(n10278), .Z(n10076) );
  XOR2_X1 U10123 ( .A(n10279), .B(n10280), .Z(n10278) );
  OR2_X1 U10124 ( .A1(n8030), .A2(n7569), .ZN(n10083) );
  XOR2_X1 U10125 ( .A(n10281), .B(n10282), .Z(n10080) );
  XOR2_X1 U10126 ( .A(n10283), .B(n7589), .Z(n10282) );
  OR2_X1 U10127 ( .A1(n8026), .A2(n7569), .ZN(n10087) );
  XOR2_X1 U10128 ( .A(n10284), .B(n10285), .Z(n10084) );
  XOR2_X1 U10129 ( .A(n10286), .B(n10287), .Z(n10285) );
  OR2_X1 U10130 ( .A1(n8023), .A2(n7569), .ZN(n10091) );
  XOR2_X1 U10131 ( .A(n10288), .B(n10289), .Z(n10088) );
  XOR2_X1 U10132 ( .A(n10290), .B(n10291), .Z(n10289) );
  OR2_X1 U10133 ( .A1(n8019), .A2(n7569), .ZN(n10095) );
  XOR2_X1 U10134 ( .A(n10292), .B(n10293), .Z(n10092) );
  XOR2_X1 U10135 ( .A(n10294), .B(n10295), .Z(n10293) );
  OR2_X1 U10136 ( .A1(n8016), .A2(n7569), .ZN(n10099) );
  XOR2_X1 U10137 ( .A(n10296), .B(n10297), .Z(n10096) );
  XOR2_X1 U10138 ( .A(n10298), .B(n10299), .Z(n10297) );
  OR2_X1 U10139 ( .A1(n8012), .A2(n7569), .ZN(n10103) );
  XOR2_X1 U10140 ( .A(n10300), .B(n10301), .Z(n10100) );
  XOR2_X1 U10141 ( .A(n10302), .B(n10303), .Z(n10301) );
  OR2_X1 U10142 ( .A1(n8009), .A2(n7569), .ZN(n10107) );
  XOR2_X1 U10143 ( .A(n10304), .B(n10305), .Z(n10104) );
  XOR2_X1 U10144 ( .A(n10306), .B(n10307), .Z(n10305) );
  OR2_X1 U10145 ( .A1(n8005), .A2(n7569), .ZN(n10111) );
  XOR2_X1 U10146 ( .A(n10308), .B(n10309), .Z(n10108) );
  XOR2_X1 U10147 ( .A(n10310), .B(n10311), .Z(n10309) );
  OR2_X1 U10148 ( .A1(n8002), .A2(n7569), .ZN(n10115) );
  XOR2_X1 U10149 ( .A(n10312), .B(n10313), .Z(n10112) );
  XOR2_X1 U10150 ( .A(n10314), .B(n10315), .Z(n10313) );
  OR2_X1 U10151 ( .A1(n7998), .A2(n7569), .ZN(n10119) );
  XOR2_X1 U10152 ( .A(n10316), .B(n10317), .Z(n10116) );
  XOR2_X1 U10153 ( .A(n10318), .B(n10319), .Z(n10317) );
  OR2_X1 U10154 ( .A1(n7995), .A2(n7569), .ZN(n10123) );
  XOR2_X1 U10155 ( .A(n10320), .B(n10321), .Z(n10120) );
  XOR2_X1 U10156 ( .A(n10322), .B(n10323), .Z(n10321) );
  OR2_X1 U10157 ( .A1(n7991), .A2(n7569), .ZN(n10127) );
  XOR2_X1 U10158 ( .A(n10324), .B(n10325), .Z(n10124) );
  XOR2_X1 U10159 ( .A(n10326), .B(n10327), .Z(n10325) );
  OR2_X1 U10160 ( .A1(n7988), .A2(n7569), .ZN(n10131) );
  XOR2_X1 U10161 ( .A(n10328), .B(n10329), .Z(n10128) );
  XOR2_X1 U10162 ( .A(n10330), .B(n10331), .Z(n10329) );
  XOR2_X1 U10163 ( .A(n10332), .B(n10333), .Z(n10133) );
  XOR2_X1 U10164 ( .A(n10334), .B(n10335), .Z(n10333) );
  OR2_X1 U10165 ( .A1(n7981), .A2(n7569), .ZN(n10139) );
  XNOR2_X1 U10166 ( .A(n10336), .B(n10337), .ZN(n10136) );
  XNOR2_X1 U10167 ( .A(n10338), .B(n10339), .ZN(n10336) );
  OR2_X1 U10168 ( .A1(n7977), .A2(n7569), .ZN(n10143) );
  XOR2_X1 U10169 ( .A(n10340), .B(n10341), .Z(n10140) );
  XOR2_X1 U10170 ( .A(n10342), .B(n10343), .Z(n10341) );
  OR2_X1 U10171 ( .A1(n7974), .A2(n7569), .ZN(n10147) );
  XOR2_X1 U10172 ( .A(n10344), .B(n10345), .Z(n10144) );
  XOR2_X1 U10173 ( .A(n10346), .B(n10347), .Z(n10345) );
  XOR2_X1 U10174 ( .A(n10348), .B(n10349), .Z(n10149) );
  XOR2_X1 U10175 ( .A(n10350), .B(n10351), .Z(n10349) );
  OR2_X1 U10176 ( .A1(n7967), .A2(n7569), .ZN(n10155) );
  XNOR2_X1 U10177 ( .A(n10352), .B(n10353), .ZN(n10152) );
  XNOR2_X1 U10178 ( .A(n10354), .B(n10355), .ZN(n10352) );
  OR2_X1 U10179 ( .A1(n7963), .A2(n7569), .ZN(n10159) );
  XOR2_X1 U10180 ( .A(n10356), .B(n10357), .Z(n10156) );
  XOR2_X1 U10181 ( .A(n10358), .B(n10359), .Z(n10357) );
  OR2_X1 U10182 ( .A1(n7960), .A2(n7569), .ZN(n10163) );
  XOR2_X1 U10183 ( .A(n10360), .B(n10361), .Z(n10160) );
  XOR2_X1 U10184 ( .A(n10362), .B(n10363), .Z(n10361) );
  OR2_X1 U10185 ( .A1(n7956), .A2(n7569), .ZN(n10167) );
  INV_X1 U10186 ( .A(b_25_), .ZN(n7569) );
  XNOR2_X1 U10187 ( .A(n10364), .B(n10365), .ZN(n10164) );
  XNOR2_X1 U10188 ( .A(n10366), .B(n10367), .ZN(n10364) );
  XOR2_X1 U10189 ( .A(n9957), .B(n10368), .Z(n9939) );
  XOR2_X1 U10190 ( .A(n9956), .B(n9955), .Z(n10368) );
  OR2_X1 U10191 ( .A1(n7956), .A2(n8035), .ZN(n9955) );
  OR2_X1 U10192 ( .A1(n10369), .A2(n10370), .ZN(n9956) );
  AND2_X1 U10193 ( .A1(n10367), .A2(n10366), .ZN(n10370) );
  AND2_X1 U10194 ( .A1(n10365), .A2(n10371), .ZN(n10369) );
  OR2_X1 U10195 ( .A1(n10367), .A2(n10366), .ZN(n10371) );
  OR2_X1 U10196 ( .A1(n7960), .A2(n8035), .ZN(n10366) );
  OR2_X1 U10197 ( .A1(n10372), .A2(n10373), .ZN(n10367) );
  AND2_X1 U10198 ( .A1(n10363), .A2(n10362), .ZN(n10373) );
  AND2_X1 U10199 ( .A1(n10360), .A2(n10374), .ZN(n10372) );
  OR2_X1 U10200 ( .A1(n10363), .A2(n10362), .ZN(n10374) );
  OR2_X1 U10201 ( .A1(n10375), .A2(n10376), .ZN(n10362) );
  AND2_X1 U10202 ( .A1(n10359), .A2(n10358), .ZN(n10376) );
  AND2_X1 U10203 ( .A1(n10356), .A2(n10377), .ZN(n10375) );
  OR2_X1 U10204 ( .A1(n10359), .A2(n10358), .ZN(n10377) );
  OR2_X1 U10205 ( .A1(n10378), .A2(n10379), .ZN(n10358) );
  AND2_X1 U10206 ( .A1(n10355), .A2(n10354), .ZN(n10379) );
  AND2_X1 U10207 ( .A1(n10353), .A2(n10380), .ZN(n10378) );
  OR2_X1 U10208 ( .A1(n10355), .A2(n10354), .ZN(n10380) );
  OR2_X1 U10209 ( .A1(n7970), .A2(n8035), .ZN(n10354) );
  OR2_X1 U10210 ( .A1(n10381), .A2(n10382), .ZN(n10355) );
  AND2_X1 U10211 ( .A1(n10351), .A2(n10350), .ZN(n10382) );
  AND2_X1 U10212 ( .A1(n10348), .A2(n10383), .ZN(n10381) );
  OR2_X1 U10213 ( .A1(n10351), .A2(n10350), .ZN(n10383) );
  OR2_X1 U10214 ( .A1(n10384), .A2(n10385), .ZN(n10350) );
  AND2_X1 U10215 ( .A1(n10347), .A2(n10346), .ZN(n10385) );
  AND2_X1 U10216 ( .A1(n10344), .A2(n10386), .ZN(n10384) );
  OR2_X1 U10217 ( .A1(n10347), .A2(n10346), .ZN(n10386) );
  OR2_X1 U10218 ( .A1(n10387), .A2(n10388), .ZN(n10346) );
  AND2_X1 U10219 ( .A1(n10343), .A2(n10342), .ZN(n10388) );
  AND2_X1 U10220 ( .A1(n10340), .A2(n10389), .ZN(n10387) );
  OR2_X1 U10221 ( .A1(n10343), .A2(n10342), .ZN(n10389) );
  OR2_X1 U10222 ( .A1(n10390), .A2(n10391), .ZN(n10342) );
  AND2_X1 U10223 ( .A1(n10339), .A2(n10338), .ZN(n10391) );
  AND2_X1 U10224 ( .A1(n10337), .A2(n10392), .ZN(n10390) );
  OR2_X1 U10225 ( .A1(n10339), .A2(n10338), .ZN(n10392) );
  OR2_X1 U10226 ( .A1(n7984), .A2(n8035), .ZN(n10338) );
  OR2_X1 U10227 ( .A1(n10393), .A2(n10394), .ZN(n10339) );
  AND2_X1 U10228 ( .A1(n10335), .A2(n10334), .ZN(n10394) );
  AND2_X1 U10229 ( .A1(n10332), .A2(n10395), .ZN(n10393) );
  OR2_X1 U10230 ( .A1(n10335), .A2(n10334), .ZN(n10395) );
  OR2_X1 U10231 ( .A1(n10396), .A2(n10397), .ZN(n10334) );
  AND2_X1 U10232 ( .A1(n10331), .A2(n10330), .ZN(n10397) );
  AND2_X1 U10233 ( .A1(n10328), .A2(n10398), .ZN(n10396) );
  OR2_X1 U10234 ( .A1(n10331), .A2(n10330), .ZN(n10398) );
  OR2_X1 U10235 ( .A1(n10399), .A2(n10400), .ZN(n10330) );
  AND2_X1 U10236 ( .A1(n10327), .A2(n10326), .ZN(n10400) );
  AND2_X1 U10237 ( .A1(n10324), .A2(n10401), .ZN(n10399) );
  OR2_X1 U10238 ( .A1(n10327), .A2(n10326), .ZN(n10401) );
  OR2_X1 U10239 ( .A1(n10402), .A2(n10403), .ZN(n10326) );
  AND2_X1 U10240 ( .A1(n10323), .A2(n10322), .ZN(n10403) );
  AND2_X1 U10241 ( .A1(n10320), .A2(n10404), .ZN(n10402) );
  OR2_X1 U10242 ( .A1(n10323), .A2(n10322), .ZN(n10404) );
  OR2_X1 U10243 ( .A1(n10405), .A2(n10406), .ZN(n10322) );
  AND2_X1 U10244 ( .A1(n10319), .A2(n10318), .ZN(n10406) );
  AND2_X1 U10245 ( .A1(n10316), .A2(n10407), .ZN(n10405) );
  OR2_X1 U10246 ( .A1(n10319), .A2(n10318), .ZN(n10407) );
  OR2_X1 U10247 ( .A1(n10408), .A2(n10409), .ZN(n10318) );
  AND2_X1 U10248 ( .A1(n10315), .A2(n10314), .ZN(n10409) );
  AND2_X1 U10249 ( .A1(n10312), .A2(n10410), .ZN(n10408) );
  OR2_X1 U10250 ( .A1(n10315), .A2(n10314), .ZN(n10410) );
  OR2_X1 U10251 ( .A1(n10411), .A2(n10412), .ZN(n10314) );
  AND2_X1 U10252 ( .A1(n10311), .A2(n10310), .ZN(n10412) );
  AND2_X1 U10253 ( .A1(n10308), .A2(n10413), .ZN(n10411) );
  OR2_X1 U10254 ( .A1(n10311), .A2(n10310), .ZN(n10413) );
  OR2_X1 U10255 ( .A1(n10414), .A2(n10415), .ZN(n10310) );
  AND2_X1 U10256 ( .A1(n10307), .A2(n10306), .ZN(n10415) );
  AND2_X1 U10257 ( .A1(n10304), .A2(n10416), .ZN(n10414) );
  OR2_X1 U10258 ( .A1(n10307), .A2(n10306), .ZN(n10416) );
  OR2_X1 U10259 ( .A1(n10417), .A2(n10418), .ZN(n10306) );
  AND2_X1 U10260 ( .A1(n10303), .A2(n10302), .ZN(n10418) );
  AND2_X1 U10261 ( .A1(n10300), .A2(n10419), .ZN(n10417) );
  OR2_X1 U10262 ( .A1(n10303), .A2(n10302), .ZN(n10419) );
  OR2_X1 U10263 ( .A1(n10420), .A2(n10421), .ZN(n10302) );
  AND2_X1 U10264 ( .A1(n10299), .A2(n10298), .ZN(n10421) );
  AND2_X1 U10265 ( .A1(n10296), .A2(n10422), .ZN(n10420) );
  OR2_X1 U10266 ( .A1(n10299), .A2(n10298), .ZN(n10422) );
  OR2_X1 U10267 ( .A1(n10423), .A2(n10424), .ZN(n10298) );
  AND2_X1 U10268 ( .A1(n10295), .A2(n10294), .ZN(n10424) );
  AND2_X1 U10269 ( .A1(n10292), .A2(n10425), .ZN(n10423) );
  OR2_X1 U10270 ( .A1(n10295), .A2(n10294), .ZN(n10425) );
  OR2_X1 U10271 ( .A1(n10426), .A2(n10427), .ZN(n10294) );
  AND2_X1 U10272 ( .A1(n10291), .A2(n10290), .ZN(n10427) );
  AND2_X1 U10273 ( .A1(n10288), .A2(n10428), .ZN(n10426) );
  OR2_X1 U10274 ( .A1(n10291), .A2(n10290), .ZN(n10428) );
  OR2_X1 U10275 ( .A1(n10429), .A2(n10430), .ZN(n10290) );
  AND2_X1 U10276 ( .A1(n10287), .A2(n10286), .ZN(n10430) );
  AND2_X1 U10277 ( .A1(n10284), .A2(n10431), .ZN(n10429) );
  OR2_X1 U10278 ( .A1(n10287), .A2(n10286), .ZN(n10431) );
  OR2_X1 U10279 ( .A1(n10432), .A2(n10433), .ZN(n10286) );
  AND2_X1 U10280 ( .A1(n7589), .A2(n10283), .ZN(n10433) );
  AND2_X1 U10281 ( .A1(n10281), .A2(n10434), .ZN(n10432) );
  OR2_X1 U10282 ( .A1(n7589), .A2(n10283), .ZN(n10434) );
  OR2_X1 U10283 ( .A1(n10435), .A2(n10436), .ZN(n10283) );
  AND2_X1 U10284 ( .A1(n10280), .A2(n10279), .ZN(n10436) );
  AND2_X1 U10285 ( .A1(n10277), .A2(n10437), .ZN(n10435) );
  OR2_X1 U10286 ( .A1(n10280), .A2(n10279), .ZN(n10437) );
  OR2_X1 U10287 ( .A1(n10438), .A2(n10439), .ZN(n10279) );
  AND2_X1 U10288 ( .A1(n10276), .A2(n10275), .ZN(n10439) );
  AND2_X1 U10289 ( .A1(n10273), .A2(n10440), .ZN(n10438) );
  OR2_X1 U10290 ( .A1(n10276), .A2(n10275), .ZN(n10440) );
  OR2_X1 U10291 ( .A1(n10441), .A2(n10442), .ZN(n10275) );
  AND2_X1 U10292 ( .A1(n10272), .A2(n10271), .ZN(n10442) );
  AND2_X1 U10293 ( .A1(n10269), .A2(n10443), .ZN(n10441) );
  OR2_X1 U10294 ( .A1(n10272), .A2(n10271), .ZN(n10443) );
  OR2_X1 U10295 ( .A1(n10444), .A2(n10445), .ZN(n10271) );
  AND2_X1 U10296 ( .A1(n10268), .A2(n10267), .ZN(n10445) );
  AND2_X1 U10297 ( .A1(n10265), .A2(n10446), .ZN(n10444) );
  OR2_X1 U10298 ( .A1(n10268), .A2(n10267), .ZN(n10446) );
  OR2_X1 U10299 ( .A1(n10447), .A2(n10448), .ZN(n10267) );
  AND2_X1 U10300 ( .A1(n10261), .A2(n10449), .ZN(n10448) );
  AND2_X1 U10301 ( .A1(n10450), .A2(n10451), .ZN(n10447) );
  OR2_X1 U10302 ( .A1(n10261), .A2(n10449), .ZN(n10451) );
  INV_X1 U10303 ( .A(n10264), .ZN(n10449) );
  AND3_X1 U10304 ( .A1(n8904), .A2(b_23_), .A3(b_24_), .ZN(n10264) );
  OR2_X1 U10305 ( .A1(n8051), .A2(n8035), .ZN(n10261) );
  INV_X1 U10306 ( .A(n10263), .ZN(n10450) );
  OR2_X1 U10307 ( .A1(n10452), .A2(n10453), .ZN(n10263) );
  AND2_X1 U10308 ( .A1(b_23_), .A2(n10454), .ZN(n10453) );
  OR2_X1 U10309 ( .A1(n10455), .A2(n7490), .ZN(n10454) );
  AND2_X1 U10310 ( .A1(a_30_), .A2(n8027), .ZN(n10455) );
  AND2_X1 U10311 ( .A1(b_22_), .A2(n10456), .ZN(n10452) );
  OR2_X1 U10312 ( .A1(n10457), .A2(n7493), .ZN(n10456) );
  AND2_X1 U10313 ( .A1(a_31_), .A2(n7598), .ZN(n10457) );
  OR2_X1 U10314 ( .A1(n8048), .A2(n8035), .ZN(n10268) );
  XNOR2_X1 U10315 ( .A(n10458), .B(n10459), .ZN(n10265) );
  XNOR2_X1 U10316 ( .A(n10460), .B(n10461), .ZN(n10459) );
  OR2_X1 U10317 ( .A1(n8044), .A2(n8035), .ZN(n10272) );
  XOR2_X1 U10318 ( .A(n10462), .B(n10463), .Z(n10269) );
  XOR2_X1 U10319 ( .A(n10464), .B(n10465), .Z(n10463) );
  OR2_X1 U10320 ( .A1(n8041), .A2(n8035), .ZN(n10276) );
  XOR2_X1 U10321 ( .A(n10466), .B(n10467), .Z(n10273) );
  XOR2_X1 U10322 ( .A(n10468), .B(n10469), .Z(n10467) );
  OR2_X1 U10323 ( .A1(n8037), .A2(n8035), .ZN(n10280) );
  XOR2_X1 U10324 ( .A(n10470), .B(n10471), .Z(n10277) );
  XOR2_X1 U10325 ( .A(n10472), .B(n10473), .Z(n10471) );
  OR2_X1 U10326 ( .A1(n8034), .A2(n8035), .ZN(n7589) );
  XOR2_X1 U10327 ( .A(n10474), .B(n10475), .Z(n10281) );
  XOR2_X1 U10328 ( .A(n10476), .B(n10477), .Z(n10475) );
  OR2_X1 U10329 ( .A1(n8030), .A2(n8035), .ZN(n10287) );
  XOR2_X1 U10330 ( .A(n10478), .B(n10479), .Z(n10284) );
  XOR2_X1 U10331 ( .A(n10480), .B(n10481), .Z(n10479) );
  OR2_X1 U10332 ( .A1(n8026), .A2(n8035), .ZN(n10291) );
  XOR2_X1 U10333 ( .A(n10482), .B(n10483), .Z(n10288) );
  XNOR2_X1 U10334 ( .A(n10484), .B(n7602), .ZN(n10483) );
  OR2_X1 U10335 ( .A1(n8023), .A2(n8035), .ZN(n10295) );
  XOR2_X1 U10336 ( .A(n10485), .B(n10486), .Z(n10292) );
  XOR2_X1 U10337 ( .A(n10487), .B(n10488), .Z(n10486) );
  OR2_X1 U10338 ( .A1(n8019), .A2(n8035), .ZN(n10299) );
  XOR2_X1 U10339 ( .A(n10489), .B(n10490), .Z(n10296) );
  XOR2_X1 U10340 ( .A(n10491), .B(n10492), .Z(n10490) );
  OR2_X1 U10341 ( .A1(n8016), .A2(n8035), .ZN(n10303) );
  XOR2_X1 U10342 ( .A(n10493), .B(n10494), .Z(n10300) );
  XOR2_X1 U10343 ( .A(n10495), .B(n10496), .Z(n10494) );
  OR2_X1 U10344 ( .A1(n8012), .A2(n8035), .ZN(n10307) );
  XOR2_X1 U10345 ( .A(n10497), .B(n10498), .Z(n10304) );
  XOR2_X1 U10346 ( .A(n10499), .B(n10500), .Z(n10498) );
  OR2_X1 U10347 ( .A1(n8009), .A2(n8035), .ZN(n10311) );
  XOR2_X1 U10348 ( .A(n10501), .B(n10502), .Z(n10308) );
  XOR2_X1 U10349 ( .A(n10503), .B(n10504), .Z(n10502) );
  OR2_X1 U10350 ( .A1(n8005), .A2(n8035), .ZN(n10315) );
  XOR2_X1 U10351 ( .A(n10505), .B(n10506), .Z(n10312) );
  XOR2_X1 U10352 ( .A(n10507), .B(n10508), .Z(n10506) );
  OR2_X1 U10353 ( .A1(n8002), .A2(n8035), .ZN(n10319) );
  XOR2_X1 U10354 ( .A(n10509), .B(n10510), .Z(n10316) );
  XOR2_X1 U10355 ( .A(n10511), .B(n10512), .Z(n10510) );
  OR2_X1 U10356 ( .A1(n7998), .A2(n8035), .ZN(n10323) );
  XOR2_X1 U10357 ( .A(n10513), .B(n10514), .Z(n10320) );
  XOR2_X1 U10358 ( .A(n10515), .B(n10516), .Z(n10514) );
  OR2_X1 U10359 ( .A1(n7995), .A2(n8035), .ZN(n10327) );
  XNOR2_X1 U10360 ( .A(n10517), .B(n10518), .ZN(n10324) );
  XNOR2_X1 U10361 ( .A(n10519), .B(n10520), .ZN(n10517) );
  OR2_X1 U10362 ( .A1(n7991), .A2(n8035), .ZN(n10331) );
  XOR2_X1 U10363 ( .A(n10521), .B(n10522), .Z(n10328) );
  XOR2_X1 U10364 ( .A(n10523), .B(n10524), .Z(n10522) );
  OR2_X1 U10365 ( .A1(n7988), .A2(n8035), .ZN(n10335) );
  XOR2_X1 U10366 ( .A(n10525), .B(n10526), .Z(n10332) );
  XOR2_X1 U10367 ( .A(n10527), .B(n10528), .Z(n10526) );
  XOR2_X1 U10368 ( .A(n10529), .B(n10530), .Z(n10337) );
  XOR2_X1 U10369 ( .A(n10531), .B(n10532), .Z(n10530) );
  OR2_X1 U10370 ( .A1(n7981), .A2(n8035), .ZN(n10343) );
  XNOR2_X1 U10371 ( .A(n10533), .B(n10534), .ZN(n10340) );
  XNOR2_X1 U10372 ( .A(n10535), .B(n10536), .ZN(n10533) );
  OR2_X1 U10373 ( .A1(n7977), .A2(n8035), .ZN(n10347) );
  XOR2_X1 U10374 ( .A(n10537), .B(n10538), .Z(n10344) );
  XOR2_X1 U10375 ( .A(n10539), .B(n10540), .Z(n10538) );
  OR2_X1 U10376 ( .A1(n7974), .A2(n8035), .ZN(n10351) );
  XOR2_X1 U10377 ( .A(n10541), .B(n10542), .Z(n10348) );
  XOR2_X1 U10378 ( .A(n10543), .B(n10544), .Z(n10542) );
  XOR2_X1 U10379 ( .A(n10545), .B(n10546), .Z(n10353) );
  XOR2_X1 U10380 ( .A(n10547), .B(n10548), .Z(n10546) );
  OR2_X1 U10381 ( .A1(n7967), .A2(n8035), .ZN(n10359) );
  XNOR2_X1 U10382 ( .A(n10549), .B(n10550), .ZN(n10356) );
  XNOR2_X1 U10383 ( .A(n10551), .B(n10552), .ZN(n10549) );
  OR2_X1 U10384 ( .A1(n7963), .A2(n8035), .ZN(n10363) );
  INV_X1 U10385 ( .A(b_24_), .ZN(n8035) );
  XOR2_X1 U10386 ( .A(n10553), .B(n10554), .Z(n10360) );
  XOR2_X1 U10387 ( .A(n10555), .B(n10556), .Z(n10554) );
  XOR2_X1 U10388 ( .A(n10557), .B(n10558), .Z(n10365) );
  XOR2_X1 U10389 ( .A(n10559), .B(n10560), .Z(n10558) );
  XOR2_X1 U10390 ( .A(n9947), .B(n10561), .Z(n9957) );
  XOR2_X1 U10391 ( .A(n9946), .B(n9945), .Z(n10561) );
  OR2_X1 U10392 ( .A1(n7960), .A2(n7598), .ZN(n9945) );
  OR2_X1 U10393 ( .A1(n10562), .A2(n10563), .ZN(n9946) );
  AND2_X1 U10394 ( .A1(n10560), .A2(n10559), .ZN(n10563) );
  AND2_X1 U10395 ( .A1(n10557), .A2(n10564), .ZN(n10562) );
  OR2_X1 U10396 ( .A1(n10560), .A2(n10559), .ZN(n10564) );
  OR2_X1 U10397 ( .A1(n10565), .A2(n10566), .ZN(n10559) );
  AND2_X1 U10398 ( .A1(n10556), .A2(n10555), .ZN(n10566) );
  AND2_X1 U10399 ( .A1(n10553), .A2(n10567), .ZN(n10565) );
  OR2_X1 U10400 ( .A1(n10556), .A2(n10555), .ZN(n10567) );
  OR2_X1 U10401 ( .A1(n10568), .A2(n10569), .ZN(n10555) );
  AND2_X1 U10402 ( .A1(n10552), .A2(n10551), .ZN(n10569) );
  AND2_X1 U10403 ( .A1(n10550), .A2(n10570), .ZN(n10568) );
  OR2_X1 U10404 ( .A1(n10552), .A2(n10551), .ZN(n10570) );
  OR2_X1 U10405 ( .A1(n7970), .A2(n7598), .ZN(n10551) );
  OR2_X1 U10406 ( .A1(n10571), .A2(n10572), .ZN(n10552) );
  AND2_X1 U10407 ( .A1(n10548), .A2(n10547), .ZN(n10572) );
  AND2_X1 U10408 ( .A1(n10545), .A2(n10573), .ZN(n10571) );
  OR2_X1 U10409 ( .A1(n10548), .A2(n10547), .ZN(n10573) );
  OR2_X1 U10410 ( .A1(n10574), .A2(n10575), .ZN(n10547) );
  AND2_X1 U10411 ( .A1(n10544), .A2(n10543), .ZN(n10575) );
  AND2_X1 U10412 ( .A1(n10541), .A2(n10576), .ZN(n10574) );
  OR2_X1 U10413 ( .A1(n10544), .A2(n10543), .ZN(n10576) );
  OR2_X1 U10414 ( .A1(n10577), .A2(n10578), .ZN(n10543) );
  AND2_X1 U10415 ( .A1(n10540), .A2(n10539), .ZN(n10578) );
  AND2_X1 U10416 ( .A1(n10537), .A2(n10579), .ZN(n10577) );
  OR2_X1 U10417 ( .A1(n10540), .A2(n10539), .ZN(n10579) );
  OR2_X1 U10418 ( .A1(n10580), .A2(n10581), .ZN(n10539) );
  AND2_X1 U10419 ( .A1(n10536), .A2(n10535), .ZN(n10581) );
  AND2_X1 U10420 ( .A1(n10534), .A2(n10582), .ZN(n10580) );
  OR2_X1 U10421 ( .A1(n10536), .A2(n10535), .ZN(n10582) );
  OR2_X1 U10422 ( .A1(n7984), .A2(n7598), .ZN(n10535) );
  OR2_X1 U10423 ( .A1(n10583), .A2(n10584), .ZN(n10536) );
  AND2_X1 U10424 ( .A1(n10532), .A2(n10531), .ZN(n10584) );
  AND2_X1 U10425 ( .A1(n10529), .A2(n10585), .ZN(n10583) );
  OR2_X1 U10426 ( .A1(n10532), .A2(n10531), .ZN(n10585) );
  OR2_X1 U10427 ( .A1(n10586), .A2(n10587), .ZN(n10531) );
  AND2_X1 U10428 ( .A1(n10528), .A2(n10527), .ZN(n10587) );
  AND2_X1 U10429 ( .A1(n10525), .A2(n10588), .ZN(n10586) );
  OR2_X1 U10430 ( .A1(n10528), .A2(n10527), .ZN(n10588) );
  OR2_X1 U10431 ( .A1(n10589), .A2(n10590), .ZN(n10527) );
  AND2_X1 U10432 ( .A1(n10524), .A2(n10523), .ZN(n10590) );
  AND2_X1 U10433 ( .A1(n10521), .A2(n10591), .ZN(n10589) );
  OR2_X1 U10434 ( .A1(n10524), .A2(n10523), .ZN(n10591) );
  OR2_X1 U10435 ( .A1(n10592), .A2(n10593), .ZN(n10523) );
  AND2_X1 U10436 ( .A1(n10520), .A2(n10519), .ZN(n10593) );
  AND2_X1 U10437 ( .A1(n10518), .A2(n10594), .ZN(n10592) );
  OR2_X1 U10438 ( .A1(n10520), .A2(n10519), .ZN(n10594) );
  OR2_X1 U10439 ( .A1(n7998), .A2(n7598), .ZN(n10519) );
  OR2_X1 U10440 ( .A1(n10595), .A2(n10596), .ZN(n10520) );
  AND2_X1 U10441 ( .A1(n10516), .A2(n10515), .ZN(n10596) );
  AND2_X1 U10442 ( .A1(n10513), .A2(n10597), .ZN(n10595) );
  OR2_X1 U10443 ( .A1(n10516), .A2(n10515), .ZN(n10597) );
  OR2_X1 U10444 ( .A1(n10598), .A2(n10599), .ZN(n10515) );
  AND2_X1 U10445 ( .A1(n10512), .A2(n10511), .ZN(n10599) );
  AND2_X1 U10446 ( .A1(n10509), .A2(n10600), .ZN(n10598) );
  OR2_X1 U10447 ( .A1(n10512), .A2(n10511), .ZN(n10600) );
  OR2_X1 U10448 ( .A1(n10601), .A2(n10602), .ZN(n10511) );
  AND2_X1 U10449 ( .A1(n10508), .A2(n10507), .ZN(n10602) );
  AND2_X1 U10450 ( .A1(n10505), .A2(n10603), .ZN(n10601) );
  OR2_X1 U10451 ( .A1(n10508), .A2(n10507), .ZN(n10603) );
  OR2_X1 U10452 ( .A1(n10604), .A2(n10605), .ZN(n10507) );
  AND2_X1 U10453 ( .A1(n10504), .A2(n10503), .ZN(n10605) );
  AND2_X1 U10454 ( .A1(n10501), .A2(n10606), .ZN(n10604) );
  OR2_X1 U10455 ( .A1(n10504), .A2(n10503), .ZN(n10606) );
  OR2_X1 U10456 ( .A1(n10607), .A2(n10608), .ZN(n10503) );
  AND2_X1 U10457 ( .A1(n10500), .A2(n10499), .ZN(n10608) );
  AND2_X1 U10458 ( .A1(n10497), .A2(n10609), .ZN(n10607) );
  OR2_X1 U10459 ( .A1(n10500), .A2(n10499), .ZN(n10609) );
  OR2_X1 U10460 ( .A1(n10610), .A2(n10611), .ZN(n10499) );
  AND2_X1 U10461 ( .A1(n10496), .A2(n10495), .ZN(n10611) );
  AND2_X1 U10462 ( .A1(n10493), .A2(n10612), .ZN(n10610) );
  OR2_X1 U10463 ( .A1(n10496), .A2(n10495), .ZN(n10612) );
  OR2_X1 U10464 ( .A1(n10613), .A2(n10614), .ZN(n10495) );
  AND2_X1 U10465 ( .A1(n10492), .A2(n10491), .ZN(n10614) );
  AND2_X1 U10466 ( .A1(n10489), .A2(n10615), .ZN(n10613) );
  OR2_X1 U10467 ( .A1(n10492), .A2(n10491), .ZN(n10615) );
  OR2_X1 U10468 ( .A1(n10616), .A2(n10617), .ZN(n10491) );
  AND2_X1 U10469 ( .A1(n10488), .A2(n10487), .ZN(n10617) );
  AND2_X1 U10470 ( .A1(n10485), .A2(n10618), .ZN(n10616) );
  OR2_X1 U10471 ( .A1(n10488), .A2(n10487), .ZN(n10618) );
  OR2_X1 U10472 ( .A1(n10619), .A2(n10620), .ZN(n10487) );
  AND2_X1 U10473 ( .A1(n8031), .A2(n10484), .ZN(n10620) );
  AND2_X1 U10474 ( .A1(n10482), .A2(n10621), .ZN(n10619) );
  OR2_X1 U10475 ( .A1(n8031), .A2(n10484), .ZN(n10621) );
  OR2_X1 U10476 ( .A1(n10622), .A2(n10623), .ZN(n10484) );
  AND2_X1 U10477 ( .A1(n10481), .A2(n10480), .ZN(n10623) );
  AND2_X1 U10478 ( .A1(n10478), .A2(n10624), .ZN(n10622) );
  OR2_X1 U10479 ( .A1(n10481), .A2(n10480), .ZN(n10624) );
  OR2_X1 U10480 ( .A1(n10625), .A2(n10626), .ZN(n10480) );
  AND2_X1 U10481 ( .A1(n10477), .A2(n10476), .ZN(n10626) );
  AND2_X1 U10482 ( .A1(n10474), .A2(n10627), .ZN(n10625) );
  OR2_X1 U10483 ( .A1(n10477), .A2(n10476), .ZN(n10627) );
  OR2_X1 U10484 ( .A1(n10628), .A2(n10629), .ZN(n10476) );
  AND2_X1 U10485 ( .A1(n10473), .A2(n10472), .ZN(n10629) );
  AND2_X1 U10486 ( .A1(n10470), .A2(n10630), .ZN(n10628) );
  OR2_X1 U10487 ( .A1(n10473), .A2(n10472), .ZN(n10630) );
  OR2_X1 U10488 ( .A1(n10631), .A2(n10632), .ZN(n10472) );
  AND2_X1 U10489 ( .A1(n10469), .A2(n10468), .ZN(n10632) );
  AND2_X1 U10490 ( .A1(n10466), .A2(n10633), .ZN(n10631) );
  OR2_X1 U10491 ( .A1(n10469), .A2(n10468), .ZN(n10633) );
  OR2_X1 U10492 ( .A1(n10634), .A2(n10635), .ZN(n10468) );
  AND2_X1 U10493 ( .A1(n10465), .A2(n10464), .ZN(n10635) );
  AND2_X1 U10494 ( .A1(n10462), .A2(n10636), .ZN(n10634) );
  OR2_X1 U10495 ( .A1(n10465), .A2(n10464), .ZN(n10636) );
  OR2_X1 U10496 ( .A1(n10637), .A2(n10638), .ZN(n10464) );
  AND2_X1 U10497 ( .A1(n10458), .A2(n10639), .ZN(n10638) );
  AND2_X1 U10498 ( .A1(n10640), .A2(n10641), .ZN(n10637) );
  OR2_X1 U10499 ( .A1(n10458), .A2(n10639), .ZN(n10641) );
  INV_X1 U10500 ( .A(n10461), .ZN(n10639) );
  AND3_X1 U10501 ( .A1(n8904), .A2(b_23_), .A3(b_22_), .ZN(n10461) );
  OR2_X1 U10502 ( .A1(n8051), .A2(n7598), .ZN(n10458) );
  INV_X1 U10503 ( .A(n10460), .ZN(n10640) );
  OR2_X1 U10504 ( .A1(n10642), .A2(n10643), .ZN(n10460) );
  AND2_X1 U10505 ( .A1(b_22_), .A2(n10644), .ZN(n10643) );
  OR2_X1 U10506 ( .A1(n10645), .A2(n7490), .ZN(n10644) );
  AND2_X1 U10507 ( .A1(a_30_), .A2(n7627), .ZN(n10645) );
  AND2_X1 U10508 ( .A1(b_21_), .A2(n10646), .ZN(n10642) );
  OR2_X1 U10509 ( .A1(n10647), .A2(n7493), .ZN(n10646) );
  AND2_X1 U10510 ( .A1(a_31_), .A2(n8027), .ZN(n10647) );
  OR2_X1 U10511 ( .A1(n8048), .A2(n7598), .ZN(n10465) );
  XNOR2_X1 U10512 ( .A(n10648), .B(n10649), .ZN(n10462) );
  XNOR2_X1 U10513 ( .A(n10650), .B(n10651), .ZN(n10649) );
  OR2_X1 U10514 ( .A1(n8044), .A2(n7598), .ZN(n10469) );
  XOR2_X1 U10515 ( .A(n10652), .B(n10653), .Z(n10466) );
  XOR2_X1 U10516 ( .A(n10654), .B(n10655), .Z(n10653) );
  OR2_X1 U10517 ( .A1(n8041), .A2(n7598), .ZN(n10473) );
  XOR2_X1 U10518 ( .A(n10656), .B(n10657), .Z(n10470) );
  XOR2_X1 U10519 ( .A(n10658), .B(n10659), .Z(n10657) );
  OR2_X1 U10520 ( .A1(n8037), .A2(n7598), .ZN(n10477) );
  XOR2_X1 U10521 ( .A(n10660), .B(n10661), .Z(n10474) );
  XOR2_X1 U10522 ( .A(n10662), .B(n10663), .Z(n10661) );
  OR2_X1 U10523 ( .A1(n8034), .A2(n7598), .ZN(n10481) );
  XOR2_X1 U10524 ( .A(n10664), .B(n10665), .Z(n10478) );
  XOR2_X1 U10525 ( .A(n10666), .B(n10667), .Z(n10665) );
  INV_X1 U10526 ( .A(n7602), .ZN(n8031) );
  AND2_X1 U10527 ( .A1(a_23_), .A2(b_23_), .ZN(n7602) );
  XOR2_X1 U10528 ( .A(n10668), .B(n10669), .Z(n10482) );
  XOR2_X1 U10529 ( .A(n10670), .B(n10671), .Z(n10669) );
  OR2_X1 U10530 ( .A1(n8026), .A2(n7598), .ZN(n10488) );
  XOR2_X1 U10531 ( .A(n10672), .B(n10673), .Z(n10485) );
  XOR2_X1 U10532 ( .A(n10674), .B(n10675), .Z(n10673) );
  OR2_X1 U10533 ( .A1(n8023), .A2(n7598), .ZN(n10492) );
  XOR2_X1 U10534 ( .A(n10676), .B(n10677), .Z(n10489) );
  XNOR2_X1 U10535 ( .A(n10678), .B(n7619), .ZN(n10677) );
  OR2_X1 U10536 ( .A1(n8019), .A2(n7598), .ZN(n10496) );
  XOR2_X1 U10537 ( .A(n10679), .B(n10680), .Z(n10493) );
  XOR2_X1 U10538 ( .A(n10681), .B(n10682), .Z(n10680) );
  OR2_X1 U10539 ( .A1(n8016), .A2(n7598), .ZN(n10500) );
  XOR2_X1 U10540 ( .A(n10683), .B(n10684), .Z(n10497) );
  XOR2_X1 U10541 ( .A(n10685), .B(n10686), .Z(n10684) );
  OR2_X1 U10542 ( .A1(n8012), .A2(n7598), .ZN(n10504) );
  XOR2_X1 U10543 ( .A(n10687), .B(n10688), .Z(n10501) );
  XOR2_X1 U10544 ( .A(n10689), .B(n10690), .Z(n10688) );
  OR2_X1 U10545 ( .A1(n8009), .A2(n7598), .ZN(n10508) );
  XOR2_X1 U10546 ( .A(n10691), .B(n10692), .Z(n10505) );
  XOR2_X1 U10547 ( .A(n10693), .B(n10694), .Z(n10692) );
  OR2_X1 U10548 ( .A1(n8005), .A2(n7598), .ZN(n10512) );
  XOR2_X1 U10549 ( .A(n10695), .B(n10696), .Z(n10509) );
  XOR2_X1 U10550 ( .A(n10697), .B(n10698), .Z(n10696) );
  OR2_X1 U10551 ( .A1(n8002), .A2(n7598), .ZN(n10516) );
  XOR2_X1 U10552 ( .A(n10699), .B(n10700), .Z(n10513) );
  XOR2_X1 U10553 ( .A(n10701), .B(n10702), .Z(n10700) );
  XOR2_X1 U10554 ( .A(n10703), .B(n10704), .Z(n10518) );
  XOR2_X1 U10555 ( .A(n10705), .B(n10706), .Z(n10704) );
  OR2_X1 U10556 ( .A1(n7995), .A2(n7598), .ZN(n10524) );
  XOR2_X1 U10557 ( .A(n10707), .B(n10708), .Z(n10521) );
  XOR2_X1 U10558 ( .A(n10709), .B(n10710), .Z(n10708) );
  OR2_X1 U10559 ( .A1(n7991), .A2(n7598), .ZN(n10528) );
  XOR2_X1 U10560 ( .A(n10711), .B(n10712), .Z(n10525) );
  XOR2_X1 U10561 ( .A(n10713), .B(n10714), .Z(n10712) );
  OR2_X1 U10562 ( .A1(n7988), .A2(n7598), .ZN(n10532) );
  XOR2_X1 U10563 ( .A(n10715), .B(n10716), .Z(n10529) );
  XOR2_X1 U10564 ( .A(n10717), .B(n10718), .Z(n10716) );
  XOR2_X1 U10565 ( .A(n10719), .B(n10720), .Z(n10534) );
  XOR2_X1 U10566 ( .A(n10721), .B(n10722), .Z(n10720) );
  OR2_X1 U10567 ( .A1(n7981), .A2(n7598), .ZN(n10540) );
  XOR2_X1 U10568 ( .A(n10723), .B(n10724), .Z(n10537) );
  XOR2_X1 U10569 ( .A(n10725), .B(n10726), .Z(n10724) );
  OR2_X1 U10570 ( .A1(n7977), .A2(n7598), .ZN(n10544) );
  XOR2_X1 U10571 ( .A(n10727), .B(n10728), .Z(n10541) );
  XOR2_X1 U10572 ( .A(n10729), .B(n10730), .Z(n10728) );
  OR2_X1 U10573 ( .A1(n7974), .A2(n7598), .ZN(n10548) );
  XOR2_X1 U10574 ( .A(n10731), .B(n10732), .Z(n10545) );
  XOR2_X1 U10575 ( .A(n10733), .B(n10734), .Z(n10732) );
  XOR2_X1 U10576 ( .A(n10735), .B(n10736), .Z(n10550) );
  XOR2_X1 U10577 ( .A(n10737), .B(n10738), .Z(n10736) );
  OR2_X1 U10578 ( .A1(n7967), .A2(n7598), .ZN(n10556) );
  XOR2_X1 U10579 ( .A(n10739), .B(n10740), .Z(n10553) );
  XOR2_X1 U10580 ( .A(n10741), .B(n10742), .Z(n10740) );
  OR2_X1 U10581 ( .A1(n7963), .A2(n7598), .ZN(n10560) );
  INV_X1 U10582 ( .A(b_23_), .ZN(n7598) );
  XOR2_X1 U10583 ( .A(n10743), .B(n10744), .Z(n10557) );
  XOR2_X1 U10584 ( .A(n10745), .B(n10746), .Z(n10744) );
  XOR2_X1 U10585 ( .A(n10747), .B(n10748), .Z(n9947) );
  XOR2_X1 U10586 ( .A(n10749), .B(n10750), .Z(n10748) );
  OR2_X1 U10587 ( .A1(n10751), .A2(n8739), .ZN(n8115) );
  XOR2_X1 U10588 ( .A(n8687), .B(n8689), .Z(n8739) );
  OR2_X1 U10589 ( .A1(n10752), .A2(n10753), .ZN(n8689) );
  AND2_X1 U10590 ( .A1(n10754), .A2(n10755), .ZN(n10753) );
  AND2_X1 U10591 ( .A1(n10756), .A2(n10757), .ZN(n10752) );
  OR2_X1 U10592 ( .A1(n10754), .A2(n10755), .ZN(n10757) );
  XOR2_X1 U10593 ( .A(n8696), .B(n10758), .Z(n8687) );
  XOR2_X1 U10594 ( .A(n8695), .B(n8694), .Z(n10758) );
  OR2_X1 U10595 ( .A1(n7950), .A2(n8020), .ZN(n8694) );
  OR2_X1 U10596 ( .A1(n10759), .A2(n10760), .ZN(n8695) );
  AND2_X1 U10597 ( .A1(n10761), .A2(n10762), .ZN(n10760) );
  AND2_X1 U10598 ( .A1(n10763), .A2(n10764), .ZN(n10759) );
  OR2_X1 U10599 ( .A1(n10761), .A2(n10762), .ZN(n10764) );
  XOR2_X1 U10600 ( .A(n8703), .B(n10765), .Z(n8696) );
  XOR2_X1 U10601 ( .A(n8702), .B(n8701), .Z(n10765) );
  OR2_X1 U10602 ( .A1(n7953), .A2(n7656), .ZN(n8701) );
  OR2_X1 U10603 ( .A1(n10766), .A2(n10767), .ZN(n8702) );
  AND2_X1 U10604 ( .A1(n10768), .A2(n10769), .ZN(n10767) );
  AND2_X1 U10605 ( .A1(n10770), .A2(n10771), .ZN(n10766) );
  OR2_X1 U10606 ( .A1(n10768), .A2(n10769), .ZN(n10771) );
  XOR2_X1 U10607 ( .A(n8710), .B(n10772), .Z(n8703) );
  XOR2_X1 U10608 ( .A(n8709), .B(n8708), .Z(n10772) );
  OR2_X1 U10609 ( .A1(n7956), .A2(n8013), .ZN(n8708) );
  OR2_X1 U10610 ( .A1(n10773), .A2(n10774), .ZN(n8709) );
  AND2_X1 U10611 ( .A1(n10775), .A2(n10776), .ZN(n10774) );
  AND2_X1 U10612 ( .A1(n10777), .A2(n10778), .ZN(n10773) );
  OR2_X1 U10613 ( .A1(n10775), .A2(n10776), .ZN(n10778) );
  XOR2_X1 U10614 ( .A(n8717), .B(n10779), .Z(n8710) );
  XOR2_X1 U10615 ( .A(n8716), .B(n8715), .Z(n10779) );
  OR2_X1 U10616 ( .A1(n7960), .A2(n7688), .ZN(n8715) );
  OR2_X1 U10617 ( .A1(n10780), .A2(n10781), .ZN(n8716) );
  AND2_X1 U10618 ( .A1(n10782), .A2(n10783), .ZN(n10781) );
  AND2_X1 U10619 ( .A1(n10784), .A2(n10785), .ZN(n10780) );
  OR2_X1 U10620 ( .A1(n10782), .A2(n10783), .ZN(n10785) );
  XOR2_X1 U10621 ( .A(n8724), .B(n10786), .Z(n8717) );
  XOR2_X1 U10622 ( .A(n8723), .B(n8722), .Z(n10786) );
  OR2_X1 U10623 ( .A1(n7963), .A2(n8006), .ZN(n8722) );
  OR2_X1 U10624 ( .A1(n10787), .A2(n10788), .ZN(n8723) );
  AND2_X1 U10625 ( .A1(n10789), .A2(n10790), .ZN(n10788) );
  AND2_X1 U10626 ( .A1(n10791), .A2(n10792), .ZN(n10787) );
  OR2_X1 U10627 ( .A1(n10789), .A2(n10790), .ZN(n10792) );
  XOR2_X1 U10628 ( .A(n8731), .B(n10793), .Z(n8724) );
  XOR2_X1 U10629 ( .A(n8730), .B(n8729), .Z(n10793) );
  OR2_X1 U10630 ( .A1(n7967), .A2(n7717), .ZN(n8729) );
  OR2_X1 U10631 ( .A1(n10794), .A2(n10795), .ZN(n8730) );
  AND2_X1 U10632 ( .A1(n10796), .A2(n10797), .ZN(n10795) );
  AND2_X1 U10633 ( .A1(n10798), .A2(n10799), .ZN(n10794) );
  OR2_X1 U10634 ( .A1(n10797), .A2(n10796), .ZN(n10799) );
  XOR2_X1 U10635 ( .A(n10800), .B(n10801), .Z(n8731) );
  XOR2_X1 U10636 ( .A(n10802), .B(n10803), .Z(n10801) );
  AND2_X1 U10637 ( .A1(n8740), .A2(n8738), .ZN(n10751) );
  XNOR2_X1 U10638 ( .A(n10756), .B(n10804), .ZN(n8738) );
  XOR2_X1 U10639 ( .A(n10755), .B(n10754), .Z(n10804) );
  OR2_X1 U10640 ( .A1(n7950), .A2(n7627), .ZN(n10754) );
  OR2_X1 U10641 ( .A1(n10805), .A2(n10806), .ZN(n10755) );
  AND2_X1 U10642 ( .A1(n10807), .A2(n10808), .ZN(n10806) );
  AND2_X1 U10643 ( .A1(n10809), .A2(n10810), .ZN(n10805) );
  OR2_X1 U10644 ( .A1(n10807), .A2(n10808), .ZN(n10810) );
  XOR2_X1 U10645 ( .A(n10763), .B(n10811), .Z(n10756) );
  XOR2_X1 U10646 ( .A(n10762), .B(n10761), .Z(n10811) );
  OR2_X1 U10647 ( .A1(n7953), .A2(n8020), .ZN(n10761) );
  OR2_X1 U10648 ( .A1(n10812), .A2(n10813), .ZN(n10762) );
  AND2_X1 U10649 ( .A1(n10814), .A2(n10815), .ZN(n10813) );
  AND2_X1 U10650 ( .A1(n10816), .A2(n10817), .ZN(n10812) );
  OR2_X1 U10651 ( .A1(n10814), .A2(n10815), .ZN(n10817) );
  XOR2_X1 U10652 ( .A(n10770), .B(n10818), .Z(n10763) );
  XOR2_X1 U10653 ( .A(n10769), .B(n10768), .Z(n10818) );
  OR2_X1 U10654 ( .A1(n7956), .A2(n7656), .ZN(n10768) );
  OR2_X1 U10655 ( .A1(n10819), .A2(n10820), .ZN(n10769) );
  AND2_X1 U10656 ( .A1(n10821), .A2(n10822), .ZN(n10820) );
  AND2_X1 U10657 ( .A1(n10823), .A2(n10824), .ZN(n10819) );
  OR2_X1 U10658 ( .A1(n10821), .A2(n10822), .ZN(n10824) );
  XOR2_X1 U10659 ( .A(n10777), .B(n10825), .Z(n10770) );
  XOR2_X1 U10660 ( .A(n10776), .B(n10775), .Z(n10825) );
  OR2_X1 U10661 ( .A1(n7960), .A2(n8013), .ZN(n10775) );
  OR2_X1 U10662 ( .A1(n10826), .A2(n10827), .ZN(n10776) );
  AND2_X1 U10663 ( .A1(n10828), .A2(n10829), .ZN(n10827) );
  AND2_X1 U10664 ( .A1(n10830), .A2(n10831), .ZN(n10826) );
  OR2_X1 U10665 ( .A1(n10828), .A2(n10829), .ZN(n10831) );
  XOR2_X1 U10666 ( .A(n10784), .B(n10832), .Z(n10777) );
  XOR2_X1 U10667 ( .A(n10783), .B(n10782), .Z(n10832) );
  OR2_X1 U10668 ( .A1(n7963), .A2(n7688), .ZN(n10782) );
  OR2_X1 U10669 ( .A1(n10833), .A2(n10834), .ZN(n10783) );
  AND2_X1 U10670 ( .A1(n10835), .A2(n10836), .ZN(n10834) );
  AND2_X1 U10671 ( .A1(n10837), .A2(n10838), .ZN(n10833) );
  OR2_X1 U10672 ( .A1(n10835), .A2(n10836), .ZN(n10838) );
  XOR2_X1 U10673 ( .A(n10791), .B(n10839), .Z(n10784) );
  XOR2_X1 U10674 ( .A(n10790), .B(n10789), .Z(n10839) );
  OR2_X1 U10675 ( .A1(n7967), .A2(n8006), .ZN(n10789) );
  OR2_X1 U10676 ( .A1(n10840), .A2(n10841), .ZN(n10790) );
  AND2_X1 U10677 ( .A1(n10842), .A2(n10843), .ZN(n10841) );
  AND2_X1 U10678 ( .A1(n10844), .A2(n10845), .ZN(n10840) );
  OR2_X1 U10679 ( .A1(n10842), .A2(n10843), .ZN(n10845) );
  XOR2_X1 U10680 ( .A(n10798), .B(n10846), .Z(n10791) );
  XOR2_X1 U10681 ( .A(n10797), .B(n10796), .Z(n10846) );
  OR2_X1 U10682 ( .A1(n7970), .A2(n7717), .ZN(n10796) );
  OR2_X1 U10683 ( .A1(n10847), .A2(n10848), .ZN(n10797) );
  AND2_X1 U10684 ( .A1(n10849), .A2(n10850), .ZN(n10848) );
  AND2_X1 U10685 ( .A1(n10851), .A2(n10852), .ZN(n10847) );
  OR2_X1 U10686 ( .A1(n10850), .A2(n10849), .ZN(n10852) );
  XOR2_X1 U10687 ( .A(n10853), .B(n10854), .Z(n10798) );
  XOR2_X1 U10688 ( .A(n10855), .B(n10856), .Z(n10854) );
  INV_X1 U10689 ( .A(n10857), .ZN(n8740) );
  OR2_X1 U10690 ( .A1(n10858), .A2(n10859), .ZN(n10857) );
  AND2_X1 U10691 ( .A1(n8764), .A2(n8763), .ZN(n10859) );
  AND2_X1 U10692 ( .A1(n8761), .A2(n10860), .ZN(n10858) );
  OR2_X1 U10693 ( .A1(n8763), .A2(n8764), .ZN(n10860) );
  OR2_X1 U10694 ( .A1(n7950), .A2(n8027), .ZN(n8764) );
  OR2_X1 U10695 ( .A1(n10861), .A2(n10862), .ZN(n8763) );
  AND2_X1 U10696 ( .A1(n8788), .A2(n8787), .ZN(n10862) );
  AND2_X1 U10697 ( .A1(n8785), .A2(n10863), .ZN(n10861) );
  OR2_X1 U10698 ( .A1(n8787), .A2(n8788), .ZN(n10863) );
  OR2_X1 U10699 ( .A1(n7953), .A2(n8027), .ZN(n8788) );
  OR2_X1 U10700 ( .A1(n10864), .A2(n10865), .ZN(n8787) );
  AND2_X1 U10701 ( .A1(n9933), .A2(n9932), .ZN(n10865) );
  AND2_X1 U10702 ( .A1(n9930), .A2(n10866), .ZN(n10864) );
  OR2_X1 U10703 ( .A1(n9932), .A2(n9933), .ZN(n10866) );
  OR2_X1 U10704 ( .A1(n7956), .A2(n8027), .ZN(n9933) );
  OR2_X1 U10705 ( .A1(n10867), .A2(n10868), .ZN(n9932) );
  AND2_X1 U10706 ( .A1(n9952), .A2(n9951), .ZN(n10868) );
  AND2_X1 U10707 ( .A1(n9949), .A2(n10869), .ZN(n10867) );
  OR2_X1 U10708 ( .A1(n9951), .A2(n9952), .ZN(n10869) );
  OR2_X1 U10709 ( .A1(n7960), .A2(n8027), .ZN(n9952) );
  OR2_X1 U10710 ( .A1(n10870), .A2(n10871), .ZN(n9951) );
  AND2_X1 U10711 ( .A1(n10750), .A2(n10749), .ZN(n10871) );
  AND2_X1 U10712 ( .A1(n10747), .A2(n10872), .ZN(n10870) );
  OR2_X1 U10713 ( .A1(n10749), .A2(n10750), .ZN(n10872) );
  OR2_X1 U10714 ( .A1(n7963), .A2(n8027), .ZN(n10750) );
  OR2_X1 U10715 ( .A1(n10873), .A2(n10874), .ZN(n10749) );
  AND2_X1 U10716 ( .A1(n10746), .A2(n10745), .ZN(n10874) );
  AND2_X1 U10717 ( .A1(n10743), .A2(n10875), .ZN(n10873) );
  OR2_X1 U10718 ( .A1(n10745), .A2(n10746), .ZN(n10875) );
  OR2_X1 U10719 ( .A1(n7967), .A2(n8027), .ZN(n10746) );
  OR2_X1 U10720 ( .A1(n10876), .A2(n10877), .ZN(n10745) );
  AND2_X1 U10721 ( .A1(n10742), .A2(n10741), .ZN(n10877) );
  AND2_X1 U10722 ( .A1(n10739), .A2(n10878), .ZN(n10876) );
  OR2_X1 U10723 ( .A1(n10741), .A2(n10742), .ZN(n10878) );
  OR2_X1 U10724 ( .A1(n7970), .A2(n8027), .ZN(n10742) );
  OR2_X1 U10725 ( .A1(n10879), .A2(n10880), .ZN(n10741) );
  AND2_X1 U10726 ( .A1(n10738), .A2(n10737), .ZN(n10880) );
  AND2_X1 U10727 ( .A1(n10735), .A2(n10881), .ZN(n10879) );
  OR2_X1 U10728 ( .A1(n10737), .A2(n10738), .ZN(n10881) );
  OR2_X1 U10729 ( .A1(n7974), .A2(n8027), .ZN(n10738) );
  OR2_X1 U10730 ( .A1(n10882), .A2(n10883), .ZN(n10737) );
  AND2_X1 U10731 ( .A1(n10734), .A2(n10733), .ZN(n10883) );
  AND2_X1 U10732 ( .A1(n10731), .A2(n10884), .ZN(n10882) );
  OR2_X1 U10733 ( .A1(n10733), .A2(n10734), .ZN(n10884) );
  OR2_X1 U10734 ( .A1(n7977), .A2(n8027), .ZN(n10734) );
  OR2_X1 U10735 ( .A1(n10885), .A2(n10886), .ZN(n10733) );
  AND2_X1 U10736 ( .A1(n10730), .A2(n10729), .ZN(n10886) );
  AND2_X1 U10737 ( .A1(n10727), .A2(n10887), .ZN(n10885) );
  OR2_X1 U10738 ( .A1(n10729), .A2(n10730), .ZN(n10887) );
  OR2_X1 U10739 ( .A1(n7981), .A2(n8027), .ZN(n10730) );
  OR2_X1 U10740 ( .A1(n10888), .A2(n10889), .ZN(n10729) );
  AND2_X1 U10741 ( .A1(n10726), .A2(n10725), .ZN(n10889) );
  AND2_X1 U10742 ( .A1(n10723), .A2(n10890), .ZN(n10888) );
  OR2_X1 U10743 ( .A1(n10725), .A2(n10726), .ZN(n10890) );
  OR2_X1 U10744 ( .A1(n7984), .A2(n8027), .ZN(n10726) );
  OR2_X1 U10745 ( .A1(n10891), .A2(n10892), .ZN(n10725) );
  AND2_X1 U10746 ( .A1(n10722), .A2(n10721), .ZN(n10892) );
  AND2_X1 U10747 ( .A1(n10719), .A2(n10893), .ZN(n10891) );
  OR2_X1 U10748 ( .A1(n10721), .A2(n10722), .ZN(n10893) );
  OR2_X1 U10749 ( .A1(n7988), .A2(n8027), .ZN(n10722) );
  OR2_X1 U10750 ( .A1(n10894), .A2(n10895), .ZN(n10721) );
  AND2_X1 U10751 ( .A1(n10718), .A2(n10717), .ZN(n10895) );
  AND2_X1 U10752 ( .A1(n10715), .A2(n10896), .ZN(n10894) );
  OR2_X1 U10753 ( .A1(n10717), .A2(n10718), .ZN(n10896) );
  OR2_X1 U10754 ( .A1(n7991), .A2(n8027), .ZN(n10718) );
  OR2_X1 U10755 ( .A1(n10897), .A2(n10898), .ZN(n10717) );
  AND2_X1 U10756 ( .A1(n10714), .A2(n10713), .ZN(n10898) );
  AND2_X1 U10757 ( .A1(n10711), .A2(n10899), .ZN(n10897) );
  OR2_X1 U10758 ( .A1(n10713), .A2(n10714), .ZN(n10899) );
  OR2_X1 U10759 ( .A1(n7995), .A2(n8027), .ZN(n10714) );
  OR2_X1 U10760 ( .A1(n10900), .A2(n10901), .ZN(n10713) );
  AND2_X1 U10761 ( .A1(n10710), .A2(n10709), .ZN(n10901) );
  AND2_X1 U10762 ( .A1(n10707), .A2(n10902), .ZN(n10900) );
  OR2_X1 U10763 ( .A1(n10709), .A2(n10710), .ZN(n10902) );
  OR2_X1 U10764 ( .A1(n7998), .A2(n8027), .ZN(n10710) );
  OR2_X1 U10765 ( .A1(n10903), .A2(n10904), .ZN(n10709) );
  AND2_X1 U10766 ( .A1(n10706), .A2(n10705), .ZN(n10904) );
  AND2_X1 U10767 ( .A1(n10703), .A2(n10905), .ZN(n10903) );
  OR2_X1 U10768 ( .A1(n10705), .A2(n10706), .ZN(n10905) );
  OR2_X1 U10769 ( .A1(n8002), .A2(n8027), .ZN(n10706) );
  OR2_X1 U10770 ( .A1(n10906), .A2(n10907), .ZN(n10705) );
  AND2_X1 U10771 ( .A1(n10702), .A2(n10701), .ZN(n10907) );
  AND2_X1 U10772 ( .A1(n10699), .A2(n10908), .ZN(n10906) );
  OR2_X1 U10773 ( .A1(n10701), .A2(n10702), .ZN(n10908) );
  OR2_X1 U10774 ( .A1(n8005), .A2(n8027), .ZN(n10702) );
  OR2_X1 U10775 ( .A1(n10909), .A2(n10910), .ZN(n10701) );
  AND2_X1 U10776 ( .A1(n10698), .A2(n10697), .ZN(n10910) );
  AND2_X1 U10777 ( .A1(n10695), .A2(n10911), .ZN(n10909) );
  OR2_X1 U10778 ( .A1(n10697), .A2(n10698), .ZN(n10911) );
  OR2_X1 U10779 ( .A1(n8009), .A2(n8027), .ZN(n10698) );
  OR2_X1 U10780 ( .A1(n10912), .A2(n10913), .ZN(n10697) );
  AND2_X1 U10781 ( .A1(n10694), .A2(n10693), .ZN(n10913) );
  AND2_X1 U10782 ( .A1(n10691), .A2(n10914), .ZN(n10912) );
  OR2_X1 U10783 ( .A1(n10693), .A2(n10694), .ZN(n10914) );
  OR2_X1 U10784 ( .A1(n8012), .A2(n8027), .ZN(n10694) );
  OR2_X1 U10785 ( .A1(n10915), .A2(n10916), .ZN(n10693) );
  AND2_X1 U10786 ( .A1(n10690), .A2(n10689), .ZN(n10916) );
  AND2_X1 U10787 ( .A1(n10687), .A2(n10917), .ZN(n10915) );
  OR2_X1 U10788 ( .A1(n10689), .A2(n10690), .ZN(n10917) );
  OR2_X1 U10789 ( .A1(n8016), .A2(n8027), .ZN(n10690) );
  OR2_X1 U10790 ( .A1(n10918), .A2(n10919), .ZN(n10689) );
  AND2_X1 U10791 ( .A1(n10686), .A2(n10685), .ZN(n10919) );
  AND2_X1 U10792 ( .A1(n10683), .A2(n10920), .ZN(n10918) );
  OR2_X1 U10793 ( .A1(n10685), .A2(n10686), .ZN(n10920) );
  OR2_X1 U10794 ( .A1(n8019), .A2(n8027), .ZN(n10686) );
  OR2_X1 U10795 ( .A1(n10921), .A2(n10922), .ZN(n10685) );
  AND2_X1 U10796 ( .A1(n10682), .A2(n10681), .ZN(n10922) );
  AND2_X1 U10797 ( .A1(n10679), .A2(n10923), .ZN(n10921) );
  OR2_X1 U10798 ( .A1(n10681), .A2(n10682), .ZN(n10923) );
  OR2_X1 U10799 ( .A1(n8023), .A2(n8027), .ZN(n10682) );
  OR2_X1 U10800 ( .A1(n10924), .A2(n10925), .ZN(n10681) );
  AND2_X1 U10801 ( .A1(n8028), .A2(n10678), .ZN(n10925) );
  AND2_X1 U10802 ( .A1(n10676), .A2(n10926), .ZN(n10924) );
  OR2_X1 U10803 ( .A1(n10678), .A2(n8028), .ZN(n10926) );
  INV_X1 U10804 ( .A(n7619), .ZN(n8028) );
  AND2_X1 U10805 ( .A1(a_22_), .A2(b_22_), .ZN(n7619) );
  OR2_X1 U10806 ( .A1(n10927), .A2(n10928), .ZN(n10678) );
  AND2_X1 U10807 ( .A1(n10675), .A2(n10674), .ZN(n10928) );
  AND2_X1 U10808 ( .A1(n10672), .A2(n10929), .ZN(n10927) );
  OR2_X1 U10809 ( .A1(n10674), .A2(n10675), .ZN(n10929) );
  OR2_X1 U10810 ( .A1(n8030), .A2(n8027), .ZN(n10675) );
  OR2_X1 U10811 ( .A1(n10930), .A2(n10931), .ZN(n10674) );
  AND2_X1 U10812 ( .A1(n10671), .A2(n10670), .ZN(n10931) );
  AND2_X1 U10813 ( .A1(n10668), .A2(n10932), .ZN(n10930) );
  OR2_X1 U10814 ( .A1(n10670), .A2(n10671), .ZN(n10932) );
  OR2_X1 U10815 ( .A1(n8034), .A2(n8027), .ZN(n10671) );
  OR2_X1 U10816 ( .A1(n10933), .A2(n10934), .ZN(n10670) );
  AND2_X1 U10817 ( .A1(n10667), .A2(n10666), .ZN(n10934) );
  AND2_X1 U10818 ( .A1(n10664), .A2(n10935), .ZN(n10933) );
  OR2_X1 U10819 ( .A1(n10666), .A2(n10667), .ZN(n10935) );
  OR2_X1 U10820 ( .A1(n8037), .A2(n8027), .ZN(n10667) );
  OR2_X1 U10821 ( .A1(n10936), .A2(n10937), .ZN(n10666) );
  AND2_X1 U10822 ( .A1(n10663), .A2(n10662), .ZN(n10937) );
  AND2_X1 U10823 ( .A1(n10660), .A2(n10938), .ZN(n10936) );
  OR2_X1 U10824 ( .A1(n10662), .A2(n10663), .ZN(n10938) );
  OR2_X1 U10825 ( .A1(n8041), .A2(n8027), .ZN(n10663) );
  OR2_X1 U10826 ( .A1(n10939), .A2(n10940), .ZN(n10662) );
  AND2_X1 U10827 ( .A1(n10659), .A2(n10658), .ZN(n10940) );
  AND2_X1 U10828 ( .A1(n10656), .A2(n10941), .ZN(n10939) );
  OR2_X1 U10829 ( .A1(n10658), .A2(n10659), .ZN(n10941) );
  OR2_X1 U10830 ( .A1(n8044), .A2(n8027), .ZN(n10659) );
  OR2_X1 U10831 ( .A1(n10942), .A2(n10943), .ZN(n10658) );
  AND2_X1 U10832 ( .A1(n10655), .A2(n10654), .ZN(n10943) );
  AND2_X1 U10833 ( .A1(n10652), .A2(n10944), .ZN(n10942) );
  OR2_X1 U10834 ( .A1(n10654), .A2(n10655), .ZN(n10944) );
  OR2_X1 U10835 ( .A1(n8048), .A2(n8027), .ZN(n10655) );
  OR2_X1 U10836 ( .A1(n10945), .A2(n10946), .ZN(n10654) );
  AND2_X1 U10837 ( .A1(n10648), .A2(n10947), .ZN(n10946) );
  AND2_X1 U10838 ( .A1(n10948), .A2(n10949), .ZN(n10945) );
  OR2_X1 U10839 ( .A1(n10947), .A2(n10648), .ZN(n10949) );
  OR2_X1 U10840 ( .A1(n8051), .A2(n8027), .ZN(n10648) );
  INV_X1 U10841 ( .A(b_22_), .ZN(n8027) );
  INV_X1 U10842 ( .A(n10651), .ZN(n10947) );
  AND3_X1 U10843 ( .A1(n8904), .A2(b_21_), .A3(b_22_), .ZN(n10651) );
  INV_X1 U10844 ( .A(n10650), .ZN(n10948) );
  OR2_X1 U10845 ( .A1(n10950), .A2(n10951), .ZN(n10650) );
  AND2_X1 U10846 ( .A1(b_21_), .A2(n10952), .ZN(n10951) );
  OR2_X1 U10847 ( .A1(n10953), .A2(n7490), .ZN(n10952) );
  AND2_X1 U10848 ( .A1(a_30_), .A2(n8020), .ZN(n10953) );
  AND2_X1 U10849 ( .A1(b_20_), .A2(n10954), .ZN(n10950) );
  OR2_X1 U10850 ( .A1(n10955), .A2(n7493), .ZN(n10954) );
  AND2_X1 U10851 ( .A1(a_31_), .A2(n7627), .ZN(n10955) );
  XNOR2_X1 U10852 ( .A(n10956), .B(n10957), .ZN(n10652) );
  XNOR2_X1 U10853 ( .A(n10958), .B(n10959), .ZN(n10957) );
  XOR2_X1 U10854 ( .A(n10960), .B(n10961), .Z(n10656) );
  XOR2_X1 U10855 ( .A(n10962), .B(n10963), .Z(n10961) );
  XOR2_X1 U10856 ( .A(n10964), .B(n10965), .Z(n10660) );
  XOR2_X1 U10857 ( .A(n10966), .B(n10967), .Z(n10965) );
  XOR2_X1 U10858 ( .A(n10968), .B(n10969), .Z(n10664) );
  XOR2_X1 U10859 ( .A(n10970), .B(n10971), .Z(n10969) );
  XOR2_X1 U10860 ( .A(n10972), .B(n10973), .Z(n10668) );
  XOR2_X1 U10861 ( .A(n10974), .B(n10975), .Z(n10973) );
  XOR2_X1 U10862 ( .A(n10976), .B(n10977), .Z(n10672) );
  XOR2_X1 U10863 ( .A(n10978), .B(n10979), .Z(n10977) );
  XOR2_X1 U10864 ( .A(n10980), .B(n10981), .Z(n10676) );
  XOR2_X1 U10865 ( .A(n10982), .B(n10983), .Z(n10981) );
  XOR2_X1 U10866 ( .A(n10984), .B(n10985), .Z(n10679) );
  XOR2_X1 U10867 ( .A(n10986), .B(n10987), .Z(n10985) );
  XOR2_X1 U10868 ( .A(n10988), .B(n10989), .Z(n10683) );
  XNOR2_X1 U10869 ( .A(n10990), .B(n7631), .ZN(n10989) );
  XOR2_X1 U10870 ( .A(n10991), .B(n10992), .Z(n10687) );
  XOR2_X1 U10871 ( .A(n10993), .B(n10994), .Z(n10992) );
  XOR2_X1 U10872 ( .A(n10995), .B(n10996), .Z(n10691) );
  XOR2_X1 U10873 ( .A(n10997), .B(n10998), .Z(n10996) );
  XOR2_X1 U10874 ( .A(n10999), .B(n11000), .Z(n10695) );
  XOR2_X1 U10875 ( .A(n11001), .B(n11002), .Z(n11000) );
  XOR2_X1 U10876 ( .A(n11003), .B(n11004), .Z(n10699) );
  XOR2_X1 U10877 ( .A(n11005), .B(n11006), .Z(n11004) );
  XOR2_X1 U10878 ( .A(n11007), .B(n11008), .Z(n10703) );
  XOR2_X1 U10879 ( .A(n11009), .B(n11010), .Z(n11008) );
  XOR2_X1 U10880 ( .A(n11011), .B(n11012), .Z(n10707) );
  XOR2_X1 U10881 ( .A(n11013), .B(n11014), .Z(n11012) );
  XOR2_X1 U10882 ( .A(n11015), .B(n11016), .Z(n10711) );
  XOR2_X1 U10883 ( .A(n11017), .B(n11018), .Z(n11016) );
  XOR2_X1 U10884 ( .A(n11019), .B(n11020), .Z(n10715) );
  XOR2_X1 U10885 ( .A(n11021), .B(n11022), .Z(n11020) );
  XOR2_X1 U10886 ( .A(n11023), .B(n11024), .Z(n10719) );
  XOR2_X1 U10887 ( .A(n11025), .B(n11026), .Z(n11024) );
  XOR2_X1 U10888 ( .A(n11027), .B(n11028), .Z(n10723) );
  XOR2_X1 U10889 ( .A(n11029), .B(n11030), .Z(n11028) );
  XOR2_X1 U10890 ( .A(n11031), .B(n11032), .Z(n10727) );
  XOR2_X1 U10891 ( .A(n11033), .B(n11034), .Z(n11032) );
  XOR2_X1 U10892 ( .A(n11035), .B(n11036), .Z(n10731) );
  XOR2_X1 U10893 ( .A(n11037), .B(n11038), .Z(n11036) );
  XOR2_X1 U10894 ( .A(n11039), .B(n11040), .Z(n10735) );
  XOR2_X1 U10895 ( .A(n11041), .B(n11042), .Z(n11040) );
  XOR2_X1 U10896 ( .A(n11043), .B(n11044), .Z(n10739) );
  XOR2_X1 U10897 ( .A(n11045), .B(n11046), .Z(n11044) );
  XOR2_X1 U10898 ( .A(n11047), .B(n11048), .Z(n10743) );
  XOR2_X1 U10899 ( .A(n11049), .B(n11050), .Z(n11048) );
  XOR2_X1 U10900 ( .A(n11051), .B(n11052), .Z(n10747) );
  XOR2_X1 U10901 ( .A(n11053), .B(n11054), .Z(n11052) );
  XOR2_X1 U10902 ( .A(n11055), .B(n11056), .Z(n9949) );
  XOR2_X1 U10903 ( .A(n11057), .B(n11058), .Z(n11056) );
  XOR2_X1 U10904 ( .A(n11059), .B(n11060), .Z(n9930) );
  XOR2_X1 U10905 ( .A(n11061), .B(n11062), .Z(n11060) );
  XOR2_X1 U10906 ( .A(n11063), .B(n11064), .Z(n8785) );
  XOR2_X1 U10907 ( .A(n11065), .B(n11066), .Z(n11064) );
  XOR2_X1 U10908 ( .A(n10809), .B(n11067), .Z(n8761) );
  XOR2_X1 U10909 ( .A(n10808), .B(n10807), .Z(n11067) );
  OR2_X1 U10910 ( .A1(n7953), .A2(n7627), .ZN(n10807) );
  OR2_X1 U10911 ( .A1(n11068), .A2(n11069), .ZN(n10808) );
  AND2_X1 U10912 ( .A1(n11066), .A2(n11065), .ZN(n11069) );
  AND2_X1 U10913 ( .A1(n11063), .A2(n11070), .ZN(n11068) );
  OR2_X1 U10914 ( .A1(n11066), .A2(n11065), .ZN(n11070) );
  OR2_X1 U10915 ( .A1(n11071), .A2(n11072), .ZN(n11065) );
  AND2_X1 U10916 ( .A1(n11062), .A2(n11061), .ZN(n11072) );
  AND2_X1 U10917 ( .A1(n11059), .A2(n11073), .ZN(n11071) );
  OR2_X1 U10918 ( .A1(n11062), .A2(n11061), .ZN(n11073) );
  OR2_X1 U10919 ( .A1(n11074), .A2(n11075), .ZN(n11061) );
  AND2_X1 U10920 ( .A1(n11058), .A2(n11057), .ZN(n11075) );
  AND2_X1 U10921 ( .A1(n11055), .A2(n11076), .ZN(n11074) );
  OR2_X1 U10922 ( .A1(n11058), .A2(n11057), .ZN(n11076) );
  OR2_X1 U10923 ( .A1(n11077), .A2(n11078), .ZN(n11057) );
  AND2_X1 U10924 ( .A1(n11054), .A2(n11053), .ZN(n11078) );
  AND2_X1 U10925 ( .A1(n11051), .A2(n11079), .ZN(n11077) );
  OR2_X1 U10926 ( .A1(n11054), .A2(n11053), .ZN(n11079) );
  OR2_X1 U10927 ( .A1(n11080), .A2(n11081), .ZN(n11053) );
  AND2_X1 U10928 ( .A1(n11050), .A2(n11049), .ZN(n11081) );
  AND2_X1 U10929 ( .A1(n11047), .A2(n11082), .ZN(n11080) );
  OR2_X1 U10930 ( .A1(n11050), .A2(n11049), .ZN(n11082) );
  OR2_X1 U10931 ( .A1(n11083), .A2(n11084), .ZN(n11049) );
  AND2_X1 U10932 ( .A1(n11046), .A2(n11045), .ZN(n11084) );
  AND2_X1 U10933 ( .A1(n11043), .A2(n11085), .ZN(n11083) );
  OR2_X1 U10934 ( .A1(n11046), .A2(n11045), .ZN(n11085) );
  OR2_X1 U10935 ( .A1(n11086), .A2(n11087), .ZN(n11045) );
  AND2_X1 U10936 ( .A1(n11042), .A2(n11041), .ZN(n11087) );
  AND2_X1 U10937 ( .A1(n11039), .A2(n11088), .ZN(n11086) );
  OR2_X1 U10938 ( .A1(n11042), .A2(n11041), .ZN(n11088) );
  OR2_X1 U10939 ( .A1(n11089), .A2(n11090), .ZN(n11041) );
  AND2_X1 U10940 ( .A1(n11038), .A2(n11037), .ZN(n11090) );
  AND2_X1 U10941 ( .A1(n11035), .A2(n11091), .ZN(n11089) );
  OR2_X1 U10942 ( .A1(n11038), .A2(n11037), .ZN(n11091) );
  OR2_X1 U10943 ( .A1(n11092), .A2(n11093), .ZN(n11037) );
  AND2_X1 U10944 ( .A1(n11034), .A2(n11033), .ZN(n11093) );
  AND2_X1 U10945 ( .A1(n11031), .A2(n11094), .ZN(n11092) );
  OR2_X1 U10946 ( .A1(n11034), .A2(n11033), .ZN(n11094) );
  OR2_X1 U10947 ( .A1(n11095), .A2(n11096), .ZN(n11033) );
  AND2_X1 U10948 ( .A1(n11030), .A2(n11029), .ZN(n11096) );
  AND2_X1 U10949 ( .A1(n11027), .A2(n11097), .ZN(n11095) );
  OR2_X1 U10950 ( .A1(n11030), .A2(n11029), .ZN(n11097) );
  OR2_X1 U10951 ( .A1(n11098), .A2(n11099), .ZN(n11029) );
  AND2_X1 U10952 ( .A1(n11026), .A2(n11025), .ZN(n11099) );
  AND2_X1 U10953 ( .A1(n11023), .A2(n11100), .ZN(n11098) );
  OR2_X1 U10954 ( .A1(n11026), .A2(n11025), .ZN(n11100) );
  OR2_X1 U10955 ( .A1(n11101), .A2(n11102), .ZN(n11025) );
  AND2_X1 U10956 ( .A1(n11022), .A2(n11021), .ZN(n11102) );
  AND2_X1 U10957 ( .A1(n11019), .A2(n11103), .ZN(n11101) );
  OR2_X1 U10958 ( .A1(n11022), .A2(n11021), .ZN(n11103) );
  OR2_X1 U10959 ( .A1(n11104), .A2(n11105), .ZN(n11021) );
  AND2_X1 U10960 ( .A1(n11018), .A2(n11017), .ZN(n11105) );
  AND2_X1 U10961 ( .A1(n11015), .A2(n11106), .ZN(n11104) );
  OR2_X1 U10962 ( .A1(n11018), .A2(n11017), .ZN(n11106) );
  OR2_X1 U10963 ( .A1(n11107), .A2(n11108), .ZN(n11017) );
  AND2_X1 U10964 ( .A1(n11014), .A2(n11013), .ZN(n11108) );
  AND2_X1 U10965 ( .A1(n11011), .A2(n11109), .ZN(n11107) );
  OR2_X1 U10966 ( .A1(n11014), .A2(n11013), .ZN(n11109) );
  OR2_X1 U10967 ( .A1(n11110), .A2(n11111), .ZN(n11013) );
  AND2_X1 U10968 ( .A1(n11010), .A2(n11009), .ZN(n11111) );
  AND2_X1 U10969 ( .A1(n11007), .A2(n11112), .ZN(n11110) );
  OR2_X1 U10970 ( .A1(n11010), .A2(n11009), .ZN(n11112) );
  OR2_X1 U10971 ( .A1(n11113), .A2(n11114), .ZN(n11009) );
  AND2_X1 U10972 ( .A1(n11006), .A2(n11005), .ZN(n11114) );
  AND2_X1 U10973 ( .A1(n11003), .A2(n11115), .ZN(n11113) );
  OR2_X1 U10974 ( .A1(n11006), .A2(n11005), .ZN(n11115) );
  OR2_X1 U10975 ( .A1(n11116), .A2(n11117), .ZN(n11005) );
  AND2_X1 U10976 ( .A1(n11002), .A2(n11001), .ZN(n11117) );
  AND2_X1 U10977 ( .A1(n10999), .A2(n11118), .ZN(n11116) );
  OR2_X1 U10978 ( .A1(n11002), .A2(n11001), .ZN(n11118) );
  OR2_X1 U10979 ( .A1(n11119), .A2(n11120), .ZN(n11001) );
  AND2_X1 U10980 ( .A1(n10998), .A2(n10997), .ZN(n11120) );
  AND2_X1 U10981 ( .A1(n10995), .A2(n11121), .ZN(n11119) );
  OR2_X1 U10982 ( .A1(n10998), .A2(n10997), .ZN(n11121) );
  OR2_X1 U10983 ( .A1(n11122), .A2(n11123), .ZN(n10997) );
  AND2_X1 U10984 ( .A1(n10994), .A2(n10993), .ZN(n11123) );
  AND2_X1 U10985 ( .A1(n10991), .A2(n11124), .ZN(n11122) );
  OR2_X1 U10986 ( .A1(n10994), .A2(n10993), .ZN(n11124) );
  OR2_X1 U10987 ( .A1(n11125), .A2(n11126), .ZN(n10993) );
  AND2_X1 U10988 ( .A1(n8024), .A2(n10990), .ZN(n11126) );
  AND2_X1 U10989 ( .A1(n10988), .A2(n11127), .ZN(n11125) );
  OR2_X1 U10990 ( .A1(n8024), .A2(n10990), .ZN(n11127) );
  OR2_X1 U10991 ( .A1(n11128), .A2(n11129), .ZN(n10990) );
  AND2_X1 U10992 ( .A1(n10987), .A2(n10986), .ZN(n11129) );
  AND2_X1 U10993 ( .A1(n10984), .A2(n11130), .ZN(n11128) );
  OR2_X1 U10994 ( .A1(n10987), .A2(n10986), .ZN(n11130) );
  OR2_X1 U10995 ( .A1(n11131), .A2(n11132), .ZN(n10986) );
  AND2_X1 U10996 ( .A1(n10983), .A2(n10982), .ZN(n11132) );
  AND2_X1 U10997 ( .A1(n10980), .A2(n11133), .ZN(n11131) );
  OR2_X1 U10998 ( .A1(n10983), .A2(n10982), .ZN(n11133) );
  OR2_X1 U10999 ( .A1(n11134), .A2(n11135), .ZN(n10982) );
  AND2_X1 U11000 ( .A1(n10979), .A2(n10978), .ZN(n11135) );
  AND2_X1 U11001 ( .A1(n10976), .A2(n11136), .ZN(n11134) );
  OR2_X1 U11002 ( .A1(n10979), .A2(n10978), .ZN(n11136) );
  OR2_X1 U11003 ( .A1(n11137), .A2(n11138), .ZN(n10978) );
  AND2_X1 U11004 ( .A1(n10975), .A2(n10974), .ZN(n11138) );
  AND2_X1 U11005 ( .A1(n10972), .A2(n11139), .ZN(n11137) );
  OR2_X1 U11006 ( .A1(n10975), .A2(n10974), .ZN(n11139) );
  OR2_X1 U11007 ( .A1(n11140), .A2(n11141), .ZN(n10974) );
  AND2_X1 U11008 ( .A1(n10971), .A2(n10970), .ZN(n11141) );
  AND2_X1 U11009 ( .A1(n10968), .A2(n11142), .ZN(n11140) );
  OR2_X1 U11010 ( .A1(n10971), .A2(n10970), .ZN(n11142) );
  OR2_X1 U11011 ( .A1(n11143), .A2(n11144), .ZN(n10970) );
  AND2_X1 U11012 ( .A1(n10967), .A2(n10966), .ZN(n11144) );
  AND2_X1 U11013 ( .A1(n10964), .A2(n11145), .ZN(n11143) );
  OR2_X1 U11014 ( .A1(n10967), .A2(n10966), .ZN(n11145) );
  OR2_X1 U11015 ( .A1(n11146), .A2(n11147), .ZN(n10966) );
  AND2_X1 U11016 ( .A1(n10963), .A2(n10962), .ZN(n11147) );
  AND2_X1 U11017 ( .A1(n10960), .A2(n11148), .ZN(n11146) );
  OR2_X1 U11018 ( .A1(n10963), .A2(n10962), .ZN(n11148) );
  OR2_X1 U11019 ( .A1(n11149), .A2(n11150), .ZN(n10962) );
  AND2_X1 U11020 ( .A1(n10956), .A2(n11151), .ZN(n11150) );
  AND2_X1 U11021 ( .A1(n11152), .A2(n11153), .ZN(n11149) );
  OR2_X1 U11022 ( .A1(n10956), .A2(n11151), .ZN(n11153) );
  INV_X1 U11023 ( .A(n10959), .ZN(n11151) );
  AND3_X1 U11024 ( .A1(n8904), .A2(b_20_), .A3(b_21_), .ZN(n10959) );
  OR2_X1 U11025 ( .A1(n8051), .A2(n7627), .ZN(n10956) );
  INV_X1 U11026 ( .A(n10958), .ZN(n11152) );
  OR2_X1 U11027 ( .A1(n11154), .A2(n11155), .ZN(n10958) );
  AND2_X1 U11028 ( .A1(b_20_), .A2(n11156), .ZN(n11155) );
  OR2_X1 U11029 ( .A1(n11157), .A2(n7490), .ZN(n11156) );
  AND2_X1 U11030 ( .A1(a_30_), .A2(n7656), .ZN(n11157) );
  AND2_X1 U11031 ( .A1(b_19_), .A2(n11158), .ZN(n11154) );
  OR2_X1 U11032 ( .A1(n11159), .A2(n7493), .ZN(n11158) );
  AND2_X1 U11033 ( .A1(a_31_), .A2(n8020), .ZN(n11159) );
  OR2_X1 U11034 ( .A1(n8048), .A2(n7627), .ZN(n10963) );
  XNOR2_X1 U11035 ( .A(n11160), .B(n11161), .ZN(n10960) );
  XNOR2_X1 U11036 ( .A(n11162), .B(n11163), .ZN(n11161) );
  OR2_X1 U11037 ( .A1(n8044), .A2(n7627), .ZN(n10967) );
  XOR2_X1 U11038 ( .A(n11164), .B(n11165), .Z(n10964) );
  XOR2_X1 U11039 ( .A(n11166), .B(n11167), .Z(n11165) );
  OR2_X1 U11040 ( .A1(n8041), .A2(n7627), .ZN(n10971) );
  XOR2_X1 U11041 ( .A(n11168), .B(n11169), .Z(n10968) );
  XOR2_X1 U11042 ( .A(n11170), .B(n11171), .Z(n11169) );
  OR2_X1 U11043 ( .A1(n8037), .A2(n7627), .ZN(n10975) );
  XOR2_X1 U11044 ( .A(n11172), .B(n11173), .Z(n10972) );
  XOR2_X1 U11045 ( .A(n11174), .B(n11175), .Z(n11173) );
  OR2_X1 U11046 ( .A1(n8034), .A2(n7627), .ZN(n10979) );
  XOR2_X1 U11047 ( .A(n11176), .B(n11177), .Z(n10976) );
  XOR2_X1 U11048 ( .A(n11178), .B(n11179), .Z(n11177) );
  OR2_X1 U11049 ( .A1(n8030), .A2(n7627), .ZN(n10983) );
  XOR2_X1 U11050 ( .A(n11180), .B(n11181), .Z(n10980) );
  XOR2_X1 U11051 ( .A(n11182), .B(n11183), .Z(n11181) );
  OR2_X1 U11052 ( .A1(n8026), .A2(n7627), .ZN(n10987) );
  XOR2_X1 U11053 ( .A(n11184), .B(n11185), .Z(n10984) );
  XOR2_X1 U11054 ( .A(n11186), .B(n11187), .Z(n11185) );
  INV_X1 U11055 ( .A(n7631), .ZN(n8024) );
  AND2_X1 U11056 ( .A1(a_21_), .A2(b_21_), .ZN(n7631) );
  XOR2_X1 U11057 ( .A(n11188), .B(n11189), .Z(n10988) );
  XOR2_X1 U11058 ( .A(n11190), .B(n11191), .Z(n11189) );
  OR2_X1 U11059 ( .A1(n8019), .A2(n7627), .ZN(n10994) );
  XOR2_X1 U11060 ( .A(n11192), .B(n11193), .Z(n10991) );
  XOR2_X1 U11061 ( .A(n11194), .B(n11195), .Z(n11193) );
  OR2_X1 U11062 ( .A1(n8016), .A2(n7627), .ZN(n10998) );
  XNOR2_X1 U11063 ( .A(n11196), .B(n11197), .ZN(n10995) );
  XNOR2_X1 U11064 ( .A(n8021), .B(n11198), .ZN(n11196) );
  OR2_X1 U11065 ( .A1(n8012), .A2(n7627), .ZN(n11002) );
  XOR2_X1 U11066 ( .A(n11199), .B(n11200), .Z(n10999) );
  XOR2_X1 U11067 ( .A(n11201), .B(n11202), .Z(n11200) );
  OR2_X1 U11068 ( .A1(n8009), .A2(n7627), .ZN(n11006) );
  XOR2_X1 U11069 ( .A(n11203), .B(n11204), .Z(n11003) );
  XOR2_X1 U11070 ( .A(n11205), .B(n11206), .Z(n11204) );
  OR2_X1 U11071 ( .A1(n8005), .A2(n7627), .ZN(n11010) );
  XOR2_X1 U11072 ( .A(n11207), .B(n11208), .Z(n11007) );
  XOR2_X1 U11073 ( .A(n11209), .B(n11210), .Z(n11208) );
  OR2_X1 U11074 ( .A1(n8002), .A2(n7627), .ZN(n11014) );
  XOR2_X1 U11075 ( .A(n11211), .B(n11212), .Z(n11011) );
  XOR2_X1 U11076 ( .A(n11213), .B(n11214), .Z(n11212) );
  OR2_X1 U11077 ( .A1(n7998), .A2(n7627), .ZN(n11018) );
  XOR2_X1 U11078 ( .A(n11215), .B(n11216), .Z(n11015) );
  XOR2_X1 U11079 ( .A(n11217), .B(n11218), .Z(n11216) );
  OR2_X1 U11080 ( .A1(n7995), .A2(n7627), .ZN(n11022) );
  XOR2_X1 U11081 ( .A(n11219), .B(n11220), .Z(n11019) );
  XOR2_X1 U11082 ( .A(n11221), .B(n11222), .Z(n11220) );
  OR2_X1 U11083 ( .A1(n7991), .A2(n7627), .ZN(n11026) );
  XOR2_X1 U11084 ( .A(n11223), .B(n11224), .Z(n11023) );
  XOR2_X1 U11085 ( .A(n11225), .B(n11226), .Z(n11224) );
  OR2_X1 U11086 ( .A1(n7988), .A2(n7627), .ZN(n11030) );
  XOR2_X1 U11087 ( .A(n11227), .B(n11228), .Z(n11027) );
  XOR2_X1 U11088 ( .A(n11229), .B(n11230), .Z(n11228) );
  OR2_X1 U11089 ( .A1(n7984), .A2(n7627), .ZN(n11034) );
  XOR2_X1 U11090 ( .A(n11231), .B(n11232), .Z(n11031) );
  XOR2_X1 U11091 ( .A(n11233), .B(n11234), .Z(n11232) );
  OR2_X1 U11092 ( .A1(n7981), .A2(n7627), .ZN(n11038) );
  XOR2_X1 U11093 ( .A(n11235), .B(n11236), .Z(n11035) );
  XOR2_X1 U11094 ( .A(n11237), .B(n11238), .Z(n11236) );
  OR2_X1 U11095 ( .A1(n7977), .A2(n7627), .ZN(n11042) );
  XOR2_X1 U11096 ( .A(n11239), .B(n11240), .Z(n11039) );
  XOR2_X1 U11097 ( .A(n11241), .B(n11242), .Z(n11240) );
  OR2_X1 U11098 ( .A1(n7974), .A2(n7627), .ZN(n11046) );
  XOR2_X1 U11099 ( .A(n11243), .B(n11244), .Z(n11043) );
  XOR2_X1 U11100 ( .A(n11245), .B(n11246), .Z(n11244) );
  OR2_X1 U11101 ( .A1(n7970), .A2(n7627), .ZN(n11050) );
  XOR2_X1 U11102 ( .A(n11247), .B(n11248), .Z(n11047) );
  XOR2_X1 U11103 ( .A(n11249), .B(n11250), .Z(n11248) );
  OR2_X1 U11104 ( .A1(n7967), .A2(n7627), .ZN(n11054) );
  XOR2_X1 U11105 ( .A(n11251), .B(n11252), .Z(n11051) );
  XOR2_X1 U11106 ( .A(n11253), .B(n11254), .Z(n11252) );
  OR2_X1 U11107 ( .A1(n7963), .A2(n7627), .ZN(n11058) );
  XOR2_X1 U11108 ( .A(n11255), .B(n11256), .Z(n11055) );
  XOR2_X1 U11109 ( .A(n11257), .B(n11258), .Z(n11256) );
  OR2_X1 U11110 ( .A1(n7960), .A2(n7627), .ZN(n11062) );
  XOR2_X1 U11111 ( .A(n11259), .B(n11260), .Z(n11059) );
  XOR2_X1 U11112 ( .A(n11261), .B(n11262), .Z(n11260) );
  OR2_X1 U11113 ( .A1(n7956), .A2(n7627), .ZN(n11066) );
  INV_X1 U11114 ( .A(b_21_), .ZN(n7627) );
  XOR2_X1 U11115 ( .A(n11263), .B(n11264), .Z(n11063) );
  XOR2_X1 U11116 ( .A(n11265), .B(n11266), .Z(n11264) );
  XOR2_X1 U11117 ( .A(n10816), .B(n11267), .Z(n10809) );
  XOR2_X1 U11118 ( .A(n10815), .B(n10814), .Z(n11267) );
  OR2_X1 U11119 ( .A1(n7956), .A2(n8020), .ZN(n10814) );
  OR2_X1 U11120 ( .A1(n11268), .A2(n11269), .ZN(n10815) );
  AND2_X1 U11121 ( .A1(n11266), .A2(n11265), .ZN(n11269) );
  AND2_X1 U11122 ( .A1(n11263), .A2(n11270), .ZN(n11268) );
  OR2_X1 U11123 ( .A1(n11266), .A2(n11265), .ZN(n11270) );
  OR2_X1 U11124 ( .A1(n11271), .A2(n11272), .ZN(n11265) );
  AND2_X1 U11125 ( .A1(n11262), .A2(n11261), .ZN(n11272) );
  AND2_X1 U11126 ( .A1(n11259), .A2(n11273), .ZN(n11271) );
  OR2_X1 U11127 ( .A1(n11262), .A2(n11261), .ZN(n11273) );
  OR2_X1 U11128 ( .A1(n11274), .A2(n11275), .ZN(n11261) );
  AND2_X1 U11129 ( .A1(n11258), .A2(n11257), .ZN(n11275) );
  AND2_X1 U11130 ( .A1(n11255), .A2(n11276), .ZN(n11274) );
  OR2_X1 U11131 ( .A1(n11258), .A2(n11257), .ZN(n11276) );
  OR2_X1 U11132 ( .A1(n11277), .A2(n11278), .ZN(n11257) );
  AND2_X1 U11133 ( .A1(n11254), .A2(n11253), .ZN(n11278) );
  AND2_X1 U11134 ( .A1(n11251), .A2(n11279), .ZN(n11277) );
  OR2_X1 U11135 ( .A1(n11254), .A2(n11253), .ZN(n11279) );
  OR2_X1 U11136 ( .A1(n11280), .A2(n11281), .ZN(n11253) );
  AND2_X1 U11137 ( .A1(n11250), .A2(n11249), .ZN(n11281) );
  AND2_X1 U11138 ( .A1(n11247), .A2(n11282), .ZN(n11280) );
  OR2_X1 U11139 ( .A1(n11250), .A2(n11249), .ZN(n11282) );
  OR2_X1 U11140 ( .A1(n11283), .A2(n11284), .ZN(n11249) );
  AND2_X1 U11141 ( .A1(n11246), .A2(n11245), .ZN(n11284) );
  AND2_X1 U11142 ( .A1(n11243), .A2(n11285), .ZN(n11283) );
  OR2_X1 U11143 ( .A1(n11246), .A2(n11245), .ZN(n11285) );
  OR2_X1 U11144 ( .A1(n11286), .A2(n11287), .ZN(n11245) );
  AND2_X1 U11145 ( .A1(n11242), .A2(n11241), .ZN(n11287) );
  AND2_X1 U11146 ( .A1(n11239), .A2(n11288), .ZN(n11286) );
  OR2_X1 U11147 ( .A1(n11242), .A2(n11241), .ZN(n11288) );
  OR2_X1 U11148 ( .A1(n11289), .A2(n11290), .ZN(n11241) );
  AND2_X1 U11149 ( .A1(n11238), .A2(n11237), .ZN(n11290) );
  AND2_X1 U11150 ( .A1(n11235), .A2(n11291), .ZN(n11289) );
  OR2_X1 U11151 ( .A1(n11238), .A2(n11237), .ZN(n11291) );
  OR2_X1 U11152 ( .A1(n11292), .A2(n11293), .ZN(n11237) );
  AND2_X1 U11153 ( .A1(n11234), .A2(n11233), .ZN(n11293) );
  AND2_X1 U11154 ( .A1(n11231), .A2(n11294), .ZN(n11292) );
  OR2_X1 U11155 ( .A1(n11234), .A2(n11233), .ZN(n11294) );
  OR2_X1 U11156 ( .A1(n11295), .A2(n11296), .ZN(n11233) );
  AND2_X1 U11157 ( .A1(n11230), .A2(n11229), .ZN(n11296) );
  AND2_X1 U11158 ( .A1(n11227), .A2(n11297), .ZN(n11295) );
  OR2_X1 U11159 ( .A1(n11230), .A2(n11229), .ZN(n11297) );
  OR2_X1 U11160 ( .A1(n11298), .A2(n11299), .ZN(n11229) );
  AND2_X1 U11161 ( .A1(n11226), .A2(n11225), .ZN(n11299) );
  AND2_X1 U11162 ( .A1(n11223), .A2(n11300), .ZN(n11298) );
  OR2_X1 U11163 ( .A1(n11226), .A2(n11225), .ZN(n11300) );
  OR2_X1 U11164 ( .A1(n11301), .A2(n11302), .ZN(n11225) );
  AND2_X1 U11165 ( .A1(n11222), .A2(n11221), .ZN(n11302) );
  AND2_X1 U11166 ( .A1(n11219), .A2(n11303), .ZN(n11301) );
  OR2_X1 U11167 ( .A1(n11222), .A2(n11221), .ZN(n11303) );
  OR2_X1 U11168 ( .A1(n11304), .A2(n11305), .ZN(n11221) );
  AND2_X1 U11169 ( .A1(n11218), .A2(n11217), .ZN(n11305) );
  AND2_X1 U11170 ( .A1(n11215), .A2(n11306), .ZN(n11304) );
  OR2_X1 U11171 ( .A1(n11218), .A2(n11217), .ZN(n11306) );
  OR2_X1 U11172 ( .A1(n11307), .A2(n11308), .ZN(n11217) );
  AND2_X1 U11173 ( .A1(n11214), .A2(n11213), .ZN(n11308) );
  AND2_X1 U11174 ( .A1(n11211), .A2(n11309), .ZN(n11307) );
  OR2_X1 U11175 ( .A1(n11214), .A2(n11213), .ZN(n11309) );
  OR2_X1 U11176 ( .A1(n11310), .A2(n11311), .ZN(n11213) );
  AND2_X1 U11177 ( .A1(n11210), .A2(n11209), .ZN(n11311) );
  AND2_X1 U11178 ( .A1(n11207), .A2(n11312), .ZN(n11310) );
  OR2_X1 U11179 ( .A1(n11210), .A2(n11209), .ZN(n11312) );
  OR2_X1 U11180 ( .A1(n11313), .A2(n11314), .ZN(n11209) );
  AND2_X1 U11181 ( .A1(n11206), .A2(n11205), .ZN(n11314) );
  AND2_X1 U11182 ( .A1(n11203), .A2(n11315), .ZN(n11313) );
  OR2_X1 U11183 ( .A1(n11206), .A2(n11205), .ZN(n11315) );
  OR2_X1 U11184 ( .A1(n11316), .A2(n11317), .ZN(n11205) );
  AND2_X1 U11185 ( .A1(n11202), .A2(n11201), .ZN(n11317) );
  AND2_X1 U11186 ( .A1(n11199), .A2(n11318), .ZN(n11316) );
  OR2_X1 U11187 ( .A1(n11202), .A2(n11201), .ZN(n11318) );
  OR2_X1 U11188 ( .A1(n11319), .A2(n11320), .ZN(n11201) );
  AND2_X1 U11189 ( .A1(n11198), .A2(n8021), .ZN(n11320) );
  AND2_X1 U11190 ( .A1(n11197), .A2(n11321), .ZN(n11319) );
  OR2_X1 U11191 ( .A1(n11198), .A2(n8021), .ZN(n11321) );
  INV_X1 U11192 ( .A(n7648), .ZN(n8021) );
  AND2_X1 U11193 ( .A1(a_20_), .A2(b_20_), .ZN(n7648) );
  OR2_X1 U11194 ( .A1(n11322), .A2(n11323), .ZN(n11198) );
  AND2_X1 U11195 ( .A1(n11195), .A2(n11194), .ZN(n11323) );
  AND2_X1 U11196 ( .A1(n11192), .A2(n11324), .ZN(n11322) );
  OR2_X1 U11197 ( .A1(n11195), .A2(n11194), .ZN(n11324) );
  OR2_X1 U11198 ( .A1(n11325), .A2(n11326), .ZN(n11194) );
  AND2_X1 U11199 ( .A1(n11191), .A2(n11190), .ZN(n11326) );
  AND2_X1 U11200 ( .A1(n11188), .A2(n11327), .ZN(n11325) );
  OR2_X1 U11201 ( .A1(n11191), .A2(n11190), .ZN(n11327) );
  OR2_X1 U11202 ( .A1(n11328), .A2(n11329), .ZN(n11190) );
  AND2_X1 U11203 ( .A1(n11187), .A2(n11186), .ZN(n11329) );
  AND2_X1 U11204 ( .A1(n11184), .A2(n11330), .ZN(n11328) );
  OR2_X1 U11205 ( .A1(n11187), .A2(n11186), .ZN(n11330) );
  OR2_X1 U11206 ( .A1(n11331), .A2(n11332), .ZN(n11186) );
  AND2_X1 U11207 ( .A1(n11183), .A2(n11182), .ZN(n11332) );
  AND2_X1 U11208 ( .A1(n11180), .A2(n11333), .ZN(n11331) );
  OR2_X1 U11209 ( .A1(n11183), .A2(n11182), .ZN(n11333) );
  OR2_X1 U11210 ( .A1(n11334), .A2(n11335), .ZN(n11182) );
  AND2_X1 U11211 ( .A1(n11179), .A2(n11178), .ZN(n11335) );
  AND2_X1 U11212 ( .A1(n11176), .A2(n11336), .ZN(n11334) );
  OR2_X1 U11213 ( .A1(n11179), .A2(n11178), .ZN(n11336) );
  OR2_X1 U11214 ( .A1(n11337), .A2(n11338), .ZN(n11178) );
  AND2_X1 U11215 ( .A1(n11175), .A2(n11174), .ZN(n11338) );
  AND2_X1 U11216 ( .A1(n11172), .A2(n11339), .ZN(n11337) );
  OR2_X1 U11217 ( .A1(n11175), .A2(n11174), .ZN(n11339) );
  OR2_X1 U11218 ( .A1(n11340), .A2(n11341), .ZN(n11174) );
  AND2_X1 U11219 ( .A1(n11171), .A2(n11170), .ZN(n11341) );
  AND2_X1 U11220 ( .A1(n11168), .A2(n11342), .ZN(n11340) );
  OR2_X1 U11221 ( .A1(n11171), .A2(n11170), .ZN(n11342) );
  OR2_X1 U11222 ( .A1(n11343), .A2(n11344), .ZN(n11170) );
  AND2_X1 U11223 ( .A1(n11167), .A2(n11166), .ZN(n11344) );
  AND2_X1 U11224 ( .A1(n11164), .A2(n11345), .ZN(n11343) );
  OR2_X1 U11225 ( .A1(n11167), .A2(n11166), .ZN(n11345) );
  OR2_X1 U11226 ( .A1(n11346), .A2(n11347), .ZN(n11166) );
  AND2_X1 U11227 ( .A1(n11160), .A2(n11348), .ZN(n11347) );
  AND2_X1 U11228 ( .A1(n11349), .A2(n11350), .ZN(n11346) );
  OR2_X1 U11229 ( .A1(n11160), .A2(n11348), .ZN(n11350) );
  INV_X1 U11230 ( .A(n11163), .ZN(n11348) );
  AND3_X1 U11231 ( .A1(n8904), .A2(b_19_), .A3(b_20_), .ZN(n11163) );
  OR2_X1 U11232 ( .A1(n8051), .A2(n8020), .ZN(n11160) );
  INV_X1 U11233 ( .A(n11162), .ZN(n11349) );
  OR2_X1 U11234 ( .A1(n11351), .A2(n11352), .ZN(n11162) );
  AND2_X1 U11235 ( .A1(b_19_), .A2(n11353), .ZN(n11352) );
  OR2_X1 U11236 ( .A1(n11354), .A2(n7490), .ZN(n11353) );
  AND2_X1 U11237 ( .A1(a_30_), .A2(n8013), .ZN(n11354) );
  AND2_X1 U11238 ( .A1(b_18_), .A2(n11355), .ZN(n11351) );
  OR2_X1 U11239 ( .A1(n11356), .A2(n7493), .ZN(n11355) );
  AND2_X1 U11240 ( .A1(a_31_), .A2(n7656), .ZN(n11356) );
  OR2_X1 U11241 ( .A1(n8048), .A2(n8020), .ZN(n11167) );
  XNOR2_X1 U11242 ( .A(n11357), .B(n11358), .ZN(n11164) );
  XNOR2_X1 U11243 ( .A(n11359), .B(n11360), .ZN(n11358) );
  OR2_X1 U11244 ( .A1(n8044), .A2(n8020), .ZN(n11171) );
  XOR2_X1 U11245 ( .A(n11361), .B(n11362), .Z(n11168) );
  XOR2_X1 U11246 ( .A(n11363), .B(n11364), .Z(n11362) );
  OR2_X1 U11247 ( .A1(n8041), .A2(n8020), .ZN(n11175) );
  XOR2_X1 U11248 ( .A(n11365), .B(n11366), .Z(n11172) );
  XOR2_X1 U11249 ( .A(n11367), .B(n11368), .Z(n11366) );
  OR2_X1 U11250 ( .A1(n8037), .A2(n8020), .ZN(n11179) );
  XOR2_X1 U11251 ( .A(n11369), .B(n11370), .Z(n11176) );
  XOR2_X1 U11252 ( .A(n11371), .B(n11372), .Z(n11370) );
  OR2_X1 U11253 ( .A1(n8034), .A2(n8020), .ZN(n11183) );
  XOR2_X1 U11254 ( .A(n11373), .B(n11374), .Z(n11180) );
  XOR2_X1 U11255 ( .A(n11375), .B(n11376), .Z(n11374) );
  OR2_X1 U11256 ( .A1(n8030), .A2(n8020), .ZN(n11187) );
  XOR2_X1 U11257 ( .A(n11377), .B(n11378), .Z(n11184) );
  XOR2_X1 U11258 ( .A(n11379), .B(n11380), .Z(n11378) );
  OR2_X1 U11259 ( .A1(n8026), .A2(n8020), .ZN(n11191) );
  XOR2_X1 U11260 ( .A(n11381), .B(n11382), .Z(n11188) );
  XOR2_X1 U11261 ( .A(n11383), .B(n11384), .Z(n11382) );
  OR2_X1 U11262 ( .A1(n8023), .A2(n8020), .ZN(n11195) );
  XOR2_X1 U11263 ( .A(n11385), .B(n11386), .Z(n11192) );
  XOR2_X1 U11264 ( .A(n11387), .B(n11388), .Z(n11386) );
  XOR2_X1 U11265 ( .A(n11389), .B(n11390), .Z(n11197) );
  XOR2_X1 U11266 ( .A(n11391), .B(n11392), .Z(n11390) );
  OR2_X1 U11267 ( .A1(n8016), .A2(n8020), .ZN(n11202) );
  XOR2_X1 U11268 ( .A(n11393), .B(n11394), .Z(n11199) );
  XOR2_X1 U11269 ( .A(n11395), .B(n11396), .Z(n11394) );
  OR2_X1 U11270 ( .A1(n8012), .A2(n8020), .ZN(n11206) );
  XOR2_X1 U11271 ( .A(n11397), .B(n11398), .Z(n11203) );
  XNOR2_X1 U11272 ( .A(n11399), .B(n7660), .ZN(n11398) );
  OR2_X1 U11273 ( .A1(n8009), .A2(n8020), .ZN(n11210) );
  XOR2_X1 U11274 ( .A(n11400), .B(n11401), .Z(n11207) );
  XOR2_X1 U11275 ( .A(n11402), .B(n11403), .Z(n11401) );
  OR2_X1 U11276 ( .A1(n8005), .A2(n8020), .ZN(n11214) );
  XOR2_X1 U11277 ( .A(n11404), .B(n11405), .Z(n11211) );
  XOR2_X1 U11278 ( .A(n11406), .B(n11407), .Z(n11405) );
  OR2_X1 U11279 ( .A1(n8002), .A2(n8020), .ZN(n11218) );
  XOR2_X1 U11280 ( .A(n11408), .B(n11409), .Z(n11215) );
  XOR2_X1 U11281 ( .A(n11410), .B(n11411), .Z(n11409) );
  OR2_X1 U11282 ( .A1(n7998), .A2(n8020), .ZN(n11222) );
  XOR2_X1 U11283 ( .A(n11412), .B(n11413), .Z(n11219) );
  XOR2_X1 U11284 ( .A(n11414), .B(n11415), .Z(n11413) );
  OR2_X1 U11285 ( .A1(n7995), .A2(n8020), .ZN(n11226) );
  XOR2_X1 U11286 ( .A(n11416), .B(n11417), .Z(n11223) );
  XOR2_X1 U11287 ( .A(n11418), .B(n11419), .Z(n11417) );
  OR2_X1 U11288 ( .A1(n7991), .A2(n8020), .ZN(n11230) );
  XOR2_X1 U11289 ( .A(n11420), .B(n11421), .Z(n11227) );
  XOR2_X1 U11290 ( .A(n11422), .B(n11423), .Z(n11421) );
  OR2_X1 U11291 ( .A1(n7988), .A2(n8020), .ZN(n11234) );
  XOR2_X1 U11292 ( .A(n11424), .B(n11425), .Z(n11231) );
  XOR2_X1 U11293 ( .A(n11426), .B(n11427), .Z(n11425) );
  OR2_X1 U11294 ( .A1(n7984), .A2(n8020), .ZN(n11238) );
  XOR2_X1 U11295 ( .A(n11428), .B(n11429), .Z(n11235) );
  XOR2_X1 U11296 ( .A(n11430), .B(n11431), .Z(n11429) );
  OR2_X1 U11297 ( .A1(n7981), .A2(n8020), .ZN(n11242) );
  XOR2_X1 U11298 ( .A(n11432), .B(n11433), .Z(n11239) );
  XOR2_X1 U11299 ( .A(n11434), .B(n11435), .Z(n11433) );
  OR2_X1 U11300 ( .A1(n7977), .A2(n8020), .ZN(n11246) );
  XOR2_X1 U11301 ( .A(n11436), .B(n11437), .Z(n11243) );
  XOR2_X1 U11302 ( .A(n11438), .B(n11439), .Z(n11437) );
  OR2_X1 U11303 ( .A1(n7974), .A2(n8020), .ZN(n11250) );
  XOR2_X1 U11304 ( .A(n11440), .B(n11441), .Z(n11247) );
  XOR2_X1 U11305 ( .A(n11442), .B(n11443), .Z(n11441) );
  OR2_X1 U11306 ( .A1(n7970), .A2(n8020), .ZN(n11254) );
  XOR2_X1 U11307 ( .A(n11444), .B(n11445), .Z(n11251) );
  XOR2_X1 U11308 ( .A(n11446), .B(n11447), .Z(n11445) );
  OR2_X1 U11309 ( .A1(n7967), .A2(n8020), .ZN(n11258) );
  XOR2_X1 U11310 ( .A(n11448), .B(n11449), .Z(n11255) );
  XOR2_X1 U11311 ( .A(n11450), .B(n11451), .Z(n11449) );
  OR2_X1 U11312 ( .A1(n7963), .A2(n8020), .ZN(n11262) );
  XOR2_X1 U11313 ( .A(n11452), .B(n11453), .Z(n11259) );
  XOR2_X1 U11314 ( .A(n11454), .B(n11455), .Z(n11453) );
  OR2_X1 U11315 ( .A1(n7960), .A2(n8020), .ZN(n11266) );
  INV_X1 U11316 ( .A(b_20_), .ZN(n8020) );
  XOR2_X1 U11317 ( .A(n11456), .B(n11457), .Z(n11263) );
  XOR2_X1 U11318 ( .A(n11458), .B(n11459), .Z(n11457) );
  XOR2_X1 U11319 ( .A(n10823), .B(n11460), .Z(n10816) );
  XOR2_X1 U11320 ( .A(n10822), .B(n10821), .Z(n11460) );
  OR2_X1 U11321 ( .A1(n7960), .A2(n7656), .ZN(n10821) );
  OR2_X1 U11322 ( .A1(n11461), .A2(n11462), .ZN(n10822) );
  AND2_X1 U11323 ( .A1(n11459), .A2(n11458), .ZN(n11462) );
  AND2_X1 U11324 ( .A1(n11456), .A2(n11463), .ZN(n11461) );
  OR2_X1 U11325 ( .A1(n11459), .A2(n11458), .ZN(n11463) );
  OR2_X1 U11326 ( .A1(n11464), .A2(n11465), .ZN(n11458) );
  AND2_X1 U11327 ( .A1(n11455), .A2(n11454), .ZN(n11465) );
  AND2_X1 U11328 ( .A1(n11452), .A2(n11466), .ZN(n11464) );
  OR2_X1 U11329 ( .A1(n11455), .A2(n11454), .ZN(n11466) );
  OR2_X1 U11330 ( .A1(n11467), .A2(n11468), .ZN(n11454) );
  AND2_X1 U11331 ( .A1(n11451), .A2(n11450), .ZN(n11468) );
  AND2_X1 U11332 ( .A1(n11448), .A2(n11469), .ZN(n11467) );
  OR2_X1 U11333 ( .A1(n11451), .A2(n11450), .ZN(n11469) );
  OR2_X1 U11334 ( .A1(n11470), .A2(n11471), .ZN(n11450) );
  AND2_X1 U11335 ( .A1(n11447), .A2(n11446), .ZN(n11471) );
  AND2_X1 U11336 ( .A1(n11444), .A2(n11472), .ZN(n11470) );
  OR2_X1 U11337 ( .A1(n11447), .A2(n11446), .ZN(n11472) );
  OR2_X1 U11338 ( .A1(n11473), .A2(n11474), .ZN(n11446) );
  AND2_X1 U11339 ( .A1(n11443), .A2(n11442), .ZN(n11474) );
  AND2_X1 U11340 ( .A1(n11440), .A2(n11475), .ZN(n11473) );
  OR2_X1 U11341 ( .A1(n11443), .A2(n11442), .ZN(n11475) );
  OR2_X1 U11342 ( .A1(n11476), .A2(n11477), .ZN(n11442) );
  AND2_X1 U11343 ( .A1(n11439), .A2(n11438), .ZN(n11477) );
  AND2_X1 U11344 ( .A1(n11436), .A2(n11478), .ZN(n11476) );
  OR2_X1 U11345 ( .A1(n11439), .A2(n11438), .ZN(n11478) );
  OR2_X1 U11346 ( .A1(n11479), .A2(n11480), .ZN(n11438) );
  AND2_X1 U11347 ( .A1(n11435), .A2(n11434), .ZN(n11480) );
  AND2_X1 U11348 ( .A1(n11432), .A2(n11481), .ZN(n11479) );
  OR2_X1 U11349 ( .A1(n11435), .A2(n11434), .ZN(n11481) );
  OR2_X1 U11350 ( .A1(n11482), .A2(n11483), .ZN(n11434) );
  AND2_X1 U11351 ( .A1(n11431), .A2(n11430), .ZN(n11483) );
  AND2_X1 U11352 ( .A1(n11428), .A2(n11484), .ZN(n11482) );
  OR2_X1 U11353 ( .A1(n11431), .A2(n11430), .ZN(n11484) );
  OR2_X1 U11354 ( .A1(n11485), .A2(n11486), .ZN(n11430) );
  AND2_X1 U11355 ( .A1(n11427), .A2(n11426), .ZN(n11486) );
  AND2_X1 U11356 ( .A1(n11424), .A2(n11487), .ZN(n11485) );
  OR2_X1 U11357 ( .A1(n11427), .A2(n11426), .ZN(n11487) );
  OR2_X1 U11358 ( .A1(n11488), .A2(n11489), .ZN(n11426) );
  AND2_X1 U11359 ( .A1(n11423), .A2(n11422), .ZN(n11489) );
  AND2_X1 U11360 ( .A1(n11420), .A2(n11490), .ZN(n11488) );
  OR2_X1 U11361 ( .A1(n11423), .A2(n11422), .ZN(n11490) );
  OR2_X1 U11362 ( .A1(n11491), .A2(n11492), .ZN(n11422) );
  AND2_X1 U11363 ( .A1(n11419), .A2(n11418), .ZN(n11492) );
  AND2_X1 U11364 ( .A1(n11416), .A2(n11493), .ZN(n11491) );
  OR2_X1 U11365 ( .A1(n11419), .A2(n11418), .ZN(n11493) );
  OR2_X1 U11366 ( .A1(n11494), .A2(n11495), .ZN(n11418) );
  AND2_X1 U11367 ( .A1(n11415), .A2(n11414), .ZN(n11495) );
  AND2_X1 U11368 ( .A1(n11412), .A2(n11496), .ZN(n11494) );
  OR2_X1 U11369 ( .A1(n11415), .A2(n11414), .ZN(n11496) );
  OR2_X1 U11370 ( .A1(n11497), .A2(n11498), .ZN(n11414) );
  AND2_X1 U11371 ( .A1(n11411), .A2(n11410), .ZN(n11498) );
  AND2_X1 U11372 ( .A1(n11408), .A2(n11499), .ZN(n11497) );
  OR2_X1 U11373 ( .A1(n11411), .A2(n11410), .ZN(n11499) );
  OR2_X1 U11374 ( .A1(n11500), .A2(n11501), .ZN(n11410) );
  AND2_X1 U11375 ( .A1(n11407), .A2(n11406), .ZN(n11501) );
  AND2_X1 U11376 ( .A1(n11404), .A2(n11502), .ZN(n11500) );
  OR2_X1 U11377 ( .A1(n11407), .A2(n11406), .ZN(n11502) );
  OR2_X1 U11378 ( .A1(n11503), .A2(n11504), .ZN(n11406) );
  AND2_X1 U11379 ( .A1(n11403), .A2(n11402), .ZN(n11504) );
  AND2_X1 U11380 ( .A1(n11400), .A2(n11505), .ZN(n11503) );
  OR2_X1 U11381 ( .A1(n11403), .A2(n11402), .ZN(n11505) );
  OR2_X1 U11382 ( .A1(n11506), .A2(n11507), .ZN(n11402) );
  AND2_X1 U11383 ( .A1(n8017), .A2(n11399), .ZN(n11507) );
  AND2_X1 U11384 ( .A1(n11397), .A2(n11508), .ZN(n11506) );
  OR2_X1 U11385 ( .A1(n8017), .A2(n11399), .ZN(n11508) );
  OR2_X1 U11386 ( .A1(n11509), .A2(n11510), .ZN(n11399) );
  AND2_X1 U11387 ( .A1(n11396), .A2(n11395), .ZN(n11510) );
  AND2_X1 U11388 ( .A1(n11393), .A2(n11511), .ZN(n11509) );
  OR2_X1 U11389 ( .A1(n11396), .A2(n11395), .ZN(n11511) );
  OR2_X1 U11390 ( .A1(n11512), .A2(n11513), .ZN(n11395) );
  AND2_X1 U11391 ( .A1(n11392), .A2(n11391), .ZN(n11513) );
  AND2_X1 U11392 ( .A1(n11389), .A2(n11514), .ZN(n11512) );
  OR2_X1 U11393 ( .A1(n11392), .A2(n11391), .ZN(n11514) );
  OR2_X1 U11394 ( .A1(n11515), .A2(n11516), .ZN(n11391) );
  AND2_X1 U11395 ( .A1(n11388), .A2(n11387), .ZN(n11516) );
  AND2_X1 U11396 ( .A1(n11385), .A2(n11517), .ZN(n11515) );
  OR2_X1 U11397 ( .A1(n11388), .A2(n11387), .ZN(n11517) );
  OR2_X1 U11398 ( .A1(n11518), .A2(n11519), .ZN(n11387) );
  AND2_X1 U11399 ( .A1(n11384), .A2(n11383), .ZN(n11519) );
  AND2_X1 U11400 ( .A1(n11381), .A2(n11520), .ZN(n11518) );
  OR2_X1 U11401 ( .A1(n11384), .A2(n11383), .ZN(n11520) );
  OR2_X1 U11402 ( .A1(n11521), .A2(n11522), .ZN(n11383) );
  AND2_X1 U11403 ( .A1(n11380), .A2(n11379), .ZN(n11522) );
  AND2_X1 U11404 ( .A1(n11377), .A2(n11523), .ZN(n11521) );
  OR2_X1 U11405 ( .A1(n11380), .A2(n11379), .ZN(n11523) );
  OR2_X1 U11406 ( .A1(n11524), .A2(n11525), .ZN(n11379) );
  AND2_X1 U11407 ( .A1(n11376), .A2(n11375), .ZN(n11525) );
  AND2_X1 U11408 ( .A1(n11373), .A2(n11526), .ZN(n11524) );
  OR2_X1 U11409 ( .A1(n11376), .A2(n11375), .ZN(n11526) );
  OR2_X1 U11410 ( .A1(n11527), .A2(n11528), .ZN(n11375) );
  AND2_X1 U11411 ( .A1(n11372), .A2(n11371), .ZN(n11528) );
  AND2_X1 U11412 ( .A1(n11369), .A2(n11529), .ZN(n11527) );
  OR2_X1 U11413 ( .A1(n11372), .A2(n11371), .ZN(n11529) );
  OR2_X1 U11414 ( .A1(n11530), .A2(n11531), .ZN(n11371) );
  AND2_X1 U11415 ( .A1(n11368), .A2(n11367), .ZN(n11531) );
  AND2_X1 U11416 ( .A1(n11365), .A2(n11532), .ZN(n11530) );
  OR2_X1 U11417 ( .A1(n11368), .A2(n11367), .ZN(n11532) );
  OR2_X1 U11418 ( .A1(n11533), .A2(n11534), .ZN(n11367) );
  AND2_X1 U11419 ( .A1(n11364), .A2(n11363), .ZN(n11534) );
  AND2_X1 U11420 ( .A1(n11361), .A2(n11535), .ZN(n11533) );
  OR2_X1 U11421 ( .A1(n11364), .A2(n11363), .ZN(n11535) );
  OR2_X1 U11422 ( .A1(n11536), .A2(n11537), .ZN(n11363) );
  AND2_X1 U11423 ( .A1(n11357), .A2(n11538), .ZN(n11537) );
  AND2_X1 U11424 ( .A1(n11539), .A2(n11540), .ZN(n11536) );
  OR2_X1 U11425 ( .A1(n11357), .A2(n11538), .ZN(n11540) );
  INV_X1 U11426 ( .A(n11360), .ZN(n11538) );
  AND3_X1 U11427 ( .A1(n8904), .A2(b_18_), .A3(b_19_), .ZN(n11360) );
  OR2_X1 U11428 ( .A1(n8051), .A2(n7656), .ZN(n11357) );
  INV_X1 U11429 ( .A(n11359), .ZN(n11539) );
  OR2_X1 U11430 ( .A1(n11541), .A2(n11542), .ZN(n11359) );
  AND2_X1 U11431 ( .A1(b_18_), .A2(n11543), .ZN(n11542) );
  OR2_X1 U11432 ( .A1(n11544), .A2(n7490), .ZN(n11543) );
  AND2_X1 U11433 ( .A1(a_30_), .A2(n7688), .ZN(n11544) );
  AND2_X1 U11434 ( .A1(b_17_), .A2(n11545), .ZN(n11541) );
  OR2_X1 U11435 ( .A1(n11546), .A2(n7493), .ZN(n11545) );
  AND2_X1 U11436 ( .A1(a_31_), .A2(n8013), .ZN(n11546) );
  OR2_X1 U11437 ( .A1(n8048), .A2(n7656), .ZN(n11364) );
  XNOR2_X1 U11438 ( .A(n11547), .B(n11548), .ZN(n11361) );
  XNOR2_X1 U11439 ( .A(n11549), .B(n11550), .ZN(n11548) );
  OR2_X1 U11440 ( .A1(n8044), .A2(n7656), .ZN(n11368) );
  XOR2_X1 U11441 ( .A(n11551), .B(n11552), .Z(n11365) );
  XOR2_X1 U11442 ( .A(n11553), .B(n11554), .Z(n11552) );
  OR2_X1 U11443 ( .A1(n8041), .A2(n7656), .ZN(n11372) );
  XOR2_X1 U11444 ( .A(n11555), .B(n11556), .Z(n11369) );
  XOR2_X1 U11445 ( .A(n11557), .B(n11558), .Z(n11556) );
  OR2_X1 U11446 ( .A1(n8037), .A2(n7656), .ZN(n11376) );
  XOR2_X1 U11447 ( .A(n11559), .B(n11560), .Z(n11373) );
  XOR2_X1 U11448 ( .A(n11561), .B(n11562), .Z(n11560) );
  OR2_X1 U11449 ( .A1(n8034), .A2(n7656), .ZN(n11380) );
  XOR2_X1 U11450 ( .A(n11563), .B(n11564), .Z(n11377) );
  XOR2_X1 U11451 ( .A(n11565), .B(n11566), .Z(n11564) );
  OR2_X1 U11452 ( .A1(n8030), .A2(n7656), .ZN(n11384) );
  XOR2_X1 U11453 ( .A(n11567), .B(n11568), .Z(n11381) );
  XOR2_X1 U11454 ( .A(n11569), .B(n11570), .Z(n11568) );
  OR2_X1 U11455 ( .A1(n8026), .A2(n7656), .ZN(n11388) );
  XOR2_X1 U11456 ( .A(n11571), .B(n11572), .Z(n11385) );
  XOR2_X1 U11457 ( .A(n11573), .B(n11574), .Z(n11572) );
  OR2_X1 U11458 ( .A1(n8023), .A2(n7656), .ZN(n11392) );
  XOR2_X1 U11459 ( .A(n11575), .B(n11576), .Z(n11389) );
  XOR2_X1 U11460 ( .A(n11577), .B(n11578), .Z(n11576) );
  OR2_X1 U11461 ( .A1(n8019), .A2(n7656), .ZN(n11396) );
  XOR2_X1 U11462 ( .A(n11579), .B(n11580), .Z(n11393) );
  XOR2_X1 U11463 ( .A(n11581), .B(n11582), .Z(n11580) );
  INV_X1 U11464 ( .A(n7660), .ZN(n8017) );
  AND2_X1 U11465 ( .A1(a_19_), .A2(b_19_), .ZN(n7660) );
  XOR2_X1 U11466 ( .A(n11583), .B(n11584), .Z(n11397) );
  XOR2_X1 U11467 ( .A(n11585), .B(n11586), .Z(n11584) );
  OR2_X1 U11468 ( .A1(n8012), .A2(n7656), .ZN(n11403) );
  XOR2_X1 U11469 ( .A(n11587), .B(n11588), .Z(n11400) );
  XOR2_X1 U11470 ( .A(n11589), .B(n11590), .Z(n11588) );
  OR2_X1 U11471 ( .A1(n8009), .A2(n7656), .ZN(n11407) );
  XNOR2_X1 U11472 ( .A(n11591), .B(n11592), .ZN(n11404) );
  XNOR2_X1 U11473 ( .A(n8014), .B(n11593), .ZN(n11591) );
  OR2_X1 U11474 ( .A1(n8005), .A2(n7656), .ZN(n11411) );
  XOR2_X1 U11475 ( .A(n11594), .B(n11595), .Z(n11408) );
  XOR2_X1 U11476 ( .A(n11596), .B(n11597), .Z(n11595) );
  OR2_X1 U11477 ( .A1(n8002), .A2(n7656), .ZN(n11415) );
  XOR2_X1 U11478 ( .A(n11598), .B(n11599), .Z(n11412) );
  XOR2_X1 U11479 ( .A(n11600), .B(n11601), .Z(n11599) );
  OR2_X1 U11480 ( .A1(n7998), .A2(n7656), .ZN(n11419) );
  XOR2_X1 U11481 ( .A(n11602), .B(n11603), .Z(n11416) );
  XOR2_X1 U11482 ( .A(n11604), .B(n11605), .Z(n11603) );
  OR2_X1 U11483 ( .A1(n7995), .A2(n7656), .ZN(n11423) );
  XOR2_X1 U11484 ( .A(n11606), .B(n11607), .Z(n11420) );
  XOR2_X1 U11485 ( .A(n11608), .B(n11609), .Z(n11607) );
  OR2_X1 U11486 ( .A1(n7991), .A2(n7656), .ZN(n11427) );
  XOR2_X1 U11487 ( .A(n11610), .B(n11611), .Z(n11424) );
  XOR2_X1 U11488 ( .A(n11612), .B(n11613), .Z(n11611) );
  OR2_X1 U11489 ( .A1(n7988), .A2(n7656), .ZN(n11431) );
  XOR2_X1 U11490 ( .A(n11614), .B(n11615), .Z(n11428) );
  XOR2_X1 U11491 ( .A(n11616), .B(n11617), .Z(n11615) );
  OR2_X1 U11492 ( .A1(n7984), .A2(n7656), .ZN(n11435) );
  XOR2_X1 U11493 ( .A(n11618), .B(n11619), .Z(n11432) );
  XOR2_X1 U11494 ( .A(n11620), .B(n11621), .Z(n11619) );
  OR2_X1 U11495 ( .A1(n7981), .A2(n7656), .ZN(n11439) );
  XOR2_X1 U11496 ( .A(n11622), .B(n11623), .Z(n11436) );
  XOR2_X1 U11497 ( .A(n11624), .B(n11625), .Z(n11623) );
  OR2_X1 U11498 ( .A1(n7977), .A2(n7656), .ZN(n11443) );
  XOR2_X1 U11499 ( .A(n11626), .B(n11627), .Z(n11440) );
  XOR2_X1 U11500 ( .A(n11628), .B(n11629), .Z(n11627) );
  OR2_X1 U11501 ( .A1(n7974), .A2(n7656), .ZN(n11447) );
  XOR2_X1 U11502 ( .A(n11630), .B(n11631), .Z(n11444) );
  XOR2_X1 U11503 ( .A(n11632), .B(n11633), .Z(n11631) );
  OR2_X1 U11504 ( .A1(n7970), .A2(n7656), .ZN(n11451) );
  XOR2_X1 U11505 ( .A(n11634), .B(n11635), .Z(n11448) );
  XOR2_X1 U11506 ( .A(n11636), .B(n11637), .Z(n11635) );
  OR2_X1 U11507 ( .A1(n7967), .A2(n7656), .ZN(n11455) );
  XOR2_X1 U11508 ( .A(n11638), .B(n11639), .Z(n11452) );
  XOR2_X1 U11509 ( .A(n11640), .B(n11641), .Z(n11639) );
  OR2_X1 U11510 ( .A1(n7963), .A2(n7656), .ZN(n11459) );
  INV_X1 U11511 ( .A(b_19_), .ZN(n7656) );
  XOR2_X1 U11512 ( .A(n11642), .B(n11643), .Z(n11456) );
  XOR2_X1 U11513 ( .A(n11644), .B(n11645), .Z(n11643) );
  XOR2_X1 U11514 ( .A(n10830), .B(n11646), .Z(n10823) );
  XOR2_X1 U11515 ( .A(n10829), .B(n10828), .Z(n11646) );
  OR2_X1 U11516 ( .A1(n7963), .A2(n8013), .ZN(n10828) );
  OR2_X1 U11517 ( .A1(n11647), .A2(n11648), .ZN(n10829) );
  AND2_X1 U11518 ( .A1(n11645), .A2(n11644), .ZN(n11648) );
  AND2_X1 U11519 ( .A1(n11642), .A2(n11649), .ZN(n11647) );
  OR2_X1 U11520 ( .A1(n11645), .A2(n11644), .ZN(n11649) );
  OR2_X1 U11521 ( .A1(n11650), .A2(n11651), .ZN(n11644) );
  AND2_X1 U11522 ( .A1(n11641), .A2(n11640), .ZN(n11651) );
  AND2_X1 U11523 ( .A1(n11638), .A2(n11652), .ZN(n11650) );
  OR2_X1 U11524 ( .A1(n11641), .A2(n11640), .ZN(n11652) );
  OR2_X1 U11525 ( .A1(n11653), .A2(n11654), .ZN(n11640) );
  AND2_X1 U11526 ( .A1(n11637), .A2(n11636), .ZN(n11654) );
  AND2_X1 U11527 ( .A1(n11634), .A2(n11655), .ZN(n11653) );
  OR2_X1 U11528 ( .A1(n11637), .A2(n11636), .ZN(n11655) );
  OR2_X1 U11529 ( .A1(n11656), .A2(n11657), .ZN(n11636) );
  AND2_X1 U11530 ( .A1(n11633), .A2(n11632), .ZN(n11657) );
  AND2_X1 U11531 ( .A1(n11630), .A2(n11658), .ZN(n11656) );
  OR2_X1 U11532 ( .A1(n11633), .A2(n11632), .ZN(n11658) );
  OR2_X1 U11533 ( .A1(n11659), .A2(n11660), .ZN(n11632) );
  AND2_X1 U11534 ( .A1(n11629), .A2(n11628), .ZN(n11660) );
  AND2_X1 U11535 ( .A1(n11626), .A2(n11661), .ZN(n11659) );
  OR2_X1 U11536 ( .A1(n11629), .A2(n11628), .ZN(n11661) );
  OR2_X1 U11537 ( .A1(n11662), .A2(n11663), .ZN(n11628) );
  AND2_X1 U11538 ( .A1(n11625), .A2(n11624), .ZN(n11663) );
  AND2_X1 U11539 ( .A1(n11622), .A2(n11664), .ZN(n11662) );
  OR2_X1 U11540 ( .A1(n11625), .A2(n11624), .ZN(n11664) );
  OR2_X1 U11541 ( .A1(n11665), .A2(n11666), .ZN(n11624) );
  AND2_X1 U11542 ( .A1(n11621), .A2(n11620), .ZN(n11666) );
  AND2_X1 U11543 ( .A1(n11618), .A2(n11667), .ZN(n11665) );
  OR2_X1 U11544 ( .A1(n11621), .A2(n11620), .ZN(n11667) );
  OR2_X1 U11545 ( .A1(n11668), .A2(n11669), .ZN(n11620) );
  AND2_X1 U11546 ( .A1(n11617), .A2(n11616), .ZN(n11669) );
  AND2_X1 U11547 ( .A1(n11614), .A2(n11670), .ZN(n11668) );
  OR2_X1 U11548 ( .A1(n11617), .A2(n11616), .ZN(n11670) );
  OR2_X1 U11549 ( .A1(n11671), .A2(n11672), .ZN(n11616) );
  AND2_X1 U11550 ( .A1(n11613), .A2(n11612), .ZN(n11672) );
  AND2_X1 U11551 ( .A1(n11610), .A2(n11673), .ZN(n11671) );
  OR2_X1 U11552 ( .A1(n11613), .A2(n11612), .ZN(n11673) );
  OR2_X1 U11553 ( .A1(n11674), .A2(n11675), .ZN(n11612) );
  AND2_X1 U11554 ( .A1(n11609), .A2(n11608), .ZN(n11675) );
  AND2_X1 U11555 ( .A1(n11606), .A2(n11676), .ZN(n11674) );
  OR2_X1 U11556 ( .A1(n11609), .A2(n11608), .ZN(n11676) );
  OR2_X1 U11557 ( .A1(n11677), .A2(n11678), .ZN(n11608) );
  AND2_X1 U11558 ( .A1(n11605), .A2(n11604), .ZN(n11678) );
  AND2_X1 U11559 ( .A1(n11602), .A2(n11679), .ZN(n11677) );
  OR2_X1 U11560 ( .A1(n11605), .A2(n11604), .ZN(n11679) );
  OR2_X1 U11561 ( .A1(n11680), .A2(n11681), .ZN(n11604) );
  AND2_X1 U11562 ( .A1(n11601), .A2(n11600), .ZN(n11681) );
  AND2_X1 U11563 ( .A1(n11598), .A2(n11682), .ZN(n11680) );
  OR2_X1 U11564 ( .A1(n11601), .A2(n11600), .ZN(n11682) );
  OR2_X1 U11565 ( .A1(n11683), .A2(n11684), .ZN(n11600) );
  AND2_X1 U11566 ( .A1(n11597), .A2(n11596), .ZN(n11684) );
  AND2_X1 U11567 ( .A1(n11594), .A2(n11685), .ZN(n11683) );
  OR2_X1 U11568 ( .A1(n11597), .A2(n11596), .ZN(n11685) );
  OR2_X1 U11569 ( .A1(n11686), .A2(n11687), .ZN(n11596) );
  AND2_X1 U11570 ( .A1(n11593), .A2(n8014), .ZN(n11687) );
  AND2_X1 U11571 ( .A1(n11592), .A2(n11688), .ZN(n11686) );
  OR2_X1 U11572 ( .A1(n11593), .A2(n8014), .ZN(n11688) );
  INV_X1 U11573 ( .A(n7677), .ZN(n8014) );
  AND2_X1 U11574 ( .A1(a_18_), .A2(b_18_), .ZN(n7677) );
  OR2_X1 U11575 ( .A1(n11689), .A2(n11690), .ZN(n11593) );
  AND2_X1 U11576 ( .A1(n11590), .A2(n11589), .ZN(n11690) );
  AND2_X1 U11577 ( .A1(n11587), .A2(n11691), .ZN(n11689) );
  OR2_X1 U11578 ( .A1(n11590), .A2(n11589), .ZN(n11691) );
  OR2_X1 U11579 ( .A1(n11692), .A2(n11693), .ZN(n11589) );
  AND2_X1 U11580 ( .A1(n11586), .A2(n11585), .ZN(n11693) );
  AND2_X1 U11581 ( .A1(n11583), .A2(n11694), .ZN(n11692) );
  OR2_X1 U11582 ( .A1(n11586), .A2(n11585), .ZN(n11694) );
  OR2_X1 U11583 ( .A1(n11695), .A2(n11696), .ZN(n11585) );
  AND2_X1 U11584 ( .A1(n11582), .A2(n11581), .ZN(n11696) );
  AND2_X1 U11585 ( .A1(n11579), .A2(n11697), .ZN(n11695) );
  OR2_X1 U11586 ( .A1(n11582), .A2(n11581), .ZN(n11697) );
  OR2_X1 U11587 ( .A1(n11698), .A2(n11699), .ZN(n11581) );
  AND2_X1 U11588 ( .A1(n11578), .A2(n11577), .ZN(n11699) );
  AND2_X1 U11589 ( .A1(n11575), .A2(n11700), .ZN(n11698) );
  OR2_X1 U11590 ( .A1(n11578), .A2(n11577), .ZN(n11700) );
  OR2_X1 U11591 ( .A1(n11701), .A2(n11702), .ZN(n11577) );
  AND2_X1 U11592 ( .A1(n11574), .A2(n11573), .ZN(n11702) );
  AND2_X1 U11593 ( .A1(n11571), .A2(n11703), .ZN(n11701) );
  OR2_X1 U11594 ( .A1(n11574), .A2(n11573), .ZN(n11703) );
  OR2_X1 U11595 ( .A1(n11704), .A2(n11705), .ZN(n11573) );
  AND2_X1 U11596 ( .A1(n11570), .A2(n11569), .ZN(n11705) );
  AND2_X1 U11597 ( .A1(n11567), .A2(n11706), .ZN(n11704) );
  OR2_X1 U11598 ( .A1(n11570), .A2(n11569), .ZN(n11706) );
  OR2_X1 U11599 ( .A1(n11707), .A2(n11708), .ZN(n11569) );
  AND2_X1 U11600 ( .A1(n11566), .A2(n11565), .ZN(n11708) );
  AND2_X1 U11601 ( .A1(n11563), .A2(n11709), .ZN(n11707) );
  OR2_X1 U11602 ( .A1(n11566), .A2(n11565), .ZN(n11709) );
  OR2_X1 U11603 ( .A1(n11710), .A2(n11711), .ZN(n11565) );
  AND2_X1 U11604 ( .A1(n11562), .A2(n11561), .ZN(n11711) );
  AND2_X1 U11605 ( .A1(n11559), .A2(n11712), .ZN(n11710) );
  OR2_X1 U11606 ( .A1(n11562), .A2(n11561), .ZN(n11712) );
  OR2_X1 U11607 ( .A1(n11713), .A2(n11714), .ZN(n11561) );
  AND2_X1 U11608 ( .A1(n11558), .A2(n11557), .ZN(n11714) );
  AND2_X1 U11609 ( .A1(n11555), .A2(n11715), .ZN(n11713) );
  OR2_X1 U11610 ( .A1(n11558), .A2(n11557), .ZN(n11715) );
  OR2_X1 U11611 ( .A1(n11716), .A2(n11717), .ZN(n11557) );
  AND2_X1 U11612 ( .A1(n11554), .A2(n11553), .ZN(n11717) );
  AND2_X1 U11613 ( .A1(n11551), .A2(n11718), .ZN(n11716) );
  OR2_X1 U11614 ( .A1(n11554), .A2(n11553), .ZN(n11718) );
  OR2_X1 U11615 ( .A1(n11719), .A2(n11720), .ZN(n11553) );
  AND2_X1 U11616 ( .A1(n11547), .A2(n11721), .ZN(n11720) );
  AND2_X1 U11617 ( .A1(n11722), .A2(n11723), .ZN(n11719) );
  OR2_X1 U11618 ( .A1(n11547), .A2(n11721), .ZN(n11723) );
  INV_X1 U11619 ( .A(n11550), .ZN(n11721) );
  AND3_X1 U11620 ( .A1(n8904), .A2(b_17_), .A3(b_18_), .ZN(n11550) );
  OR2_X1 U11621 ( .A1(n8051), .A2(n8013), .ZN(n11547) );
  INV_X1 U11622 ( .A(n11549), .ZN(n11722) );
  OR2_X1 U11623 ( .A1(n11724), .A2(n11725), .ZN(n11549) );
  AND2_X1 U11624 ( .A1(b_17_), .A2(n11726), .ZN(n11725) );
  OR2_X1 U11625 ( .A1(n11727), .A2(n7490), .ZN(n11726) );
  AND2_X1 U11626 ( .A1(a_30_), .A2(n8006), .ZN(n11727) );
  AND2_X1 U11627 ( .A1(b_16_), .A2(n11728), .ZN(n11724) );
  OR2_X1 U11628 ( .A1(n11729), .A2(n7493), .ZN(n11728) );
  AND2_X1 U11629 ( .A1(a_31_), .A2(n7688), .ZN(n11729) );
  OR2_X1 U11630 ( .A1(n8048), .A2(n8013), .ZN(n11554) );
  XNOR2_X1 U11631 ( .A(n11730), .B(n11731), .ZN(n11551) );
  XNOR2_X1 U11632 ( .A(n11732), .B(n11733), .ZN(n11731) );
  OR2_X1 U11633 ( .A1(n8044), .A2(n8013), .ZN(n11558) );
  XOR2_X1 U11634 ( .A(n11734), .B(n11735), .Z(n11555) );
  XOR2_X1 U11635 ( .A(n11736), .B(n11737), .Z(n11735) );
  OR2_X1 U11636 ( .A1(n8041), .A2(n8013), .ZN(n11562) );
  XOR2_X1 U11637 ( .A(n11738), .B(n11739), .Z(n11559) );
  XOR2_X1 U11638 ( .A(n11740), .B(n11741), .Z(n11739) );
  OR2_X1 U11639 ( .A1(n8037), .A2(n8013), .ZN(n11566) );
  XOR2_X1 U11640 ( .A(n11742), .B(n11743), .Z(n11563) );
  XOR2_X1 U11641 ( .A(n11744), .B(n11745), .Z(n11743) );
  OR2_X1 U11642 ( .A1(n8034), .A2(n8013), .ZN(n11570) );
  XOR2_X1 U11643 ( .A(n11746), .B(n11747), .Z(n11567) );
  XOR2_X1 U11644 ( .A(n11748), .B(n11749), .Z(n11747) );
  OR2_X1 U11645 ( .A1(n8030), .A2(n8013), .ZN(n11574) );
  XOR2_X1 U11646 ( .A(n11750), .B(n11751), .Z(n11571) );
  XOR2_X1 U11647 ( .A(n11752), .B(n11753), .Z(n11751) );
  OR2_X1 U11648 ( .A1(n8026), .A2(n8013), .ZN(n11578) );
  XOR2_X1 U11649 ( .A(n11754), .B(n11755), .Z(n11575) );
  XOR2_X1 U11650 ( .A(n11756), .B(n11757), .Z(n11755) );
  OR2_X1 U11651 ( .A1(n8023), .A2(n8013), .ZN(n11582) );
  XOR2_X1 U11652 ( .A(n11758), .B(n11759), .Z(n11579) );
  XOR2_X1 U11653 ( .A(n11760), .B(n11761), .Z(n11759) );
  OR2_X1 U11654 ( .A1(n8019), .A2(n8013), .ZN(n11586) );
  XOR2_X1 U11655 ( .A(n11762), .B(n11763), .Z(n11583) );
  XOR2_X1 U11656 ( .A(n11764), .B(n11765), .Z(n11763) );
  OR2_X1 U11657 ( .A1(n8016), .A2(n8013), .ZN(n11590) );
  XOR2_X1 U11658 ( .A(n11766), .B(n11767), .Z(n11587) );
  XOR2_X1 U11659 ( .A(n11768), .B(n11769), .Z(n11767) );
  XOR2_X1 U11660 ( .A(n11770), .B(n11771), .Z(n11592) );
  XOR2_X1 U11661 ( .A(n11772), .B(n11773), .Z(n11771) );
  OR2_X1 U11662 ( .A1(n8009), .A2(n8013), .ZN(n11597) );
  XOR2_X1 U11663 ( .A(n11774), .B(n11775), .Z(n11594) );
  XOR2_X1 U11664 ( .A(n11776), .B(n11777), .Z(n11775) );
  OR2_X1 U11665 ( .A1(n8005), .A2(n8013), .ZN(n11601) );
  XOR2_X1 U11666 ( .A(n11778), .B(n11779), .Z(n11598) );
  XNOR2_X1 U11667 ( .A(n11780), .B(n7692), .ZN(n11779) );
  OR2_X1 U11668 ( .A1(n8002), .A2(n8013), .ZN(n11605) );
  XOR2_X1 U11669 ( .A(n11781), .B(n11782), .Z(n11602) );
  XOR2_X1 U11670 ( .A(n11783), .B(n11784), .Z(n11782) );
  OR2_X1 U11671 ( .A1(n7998), .A2(n8013), .ZN(n11609) );
  XOR2_X1 U11672 ( .A(n11785), .B(n11786), .Z(n11606) );
  XOR2_X1 U11673 ( .A(n11787), .B(n11788), .Z(n11786) );
  OR2_X1 U11674 ( .A1(n7995), .A2(n8013), .ZN(n11613) );
  XOR2_X1 U11675 ( .A(n11789), .B(n11790), .Z(n11610) );
  XOR2_X1 U11676 ( .A(n11791), .B(n11792), .Z(n11790) );
  OR2_X1 U11677 ( .A1(n7991), .A2(n8013), .ZN(n11617) );
  XOR2_X1 U11678 ( .A(n11793), .B(n11794), .Z(n11614) );
  XOR2_X1 U11679 ( .A(n11795), .B(n11796), .Z(n11794) );
  OR2_X1 U11680 ( .A1(n7988), .A2(n8013), .ZN(n11621) );
  XOR2_X1 U11681 ( .A(n11797), .B(n11798), .Z(n11618) );
  XOR2_X1 U11682 ( .A(n11799), .B(n11800), .Z(n11798) );
  OR2_X1 U11683 ( .A1(n7984), .A2(n8013), .ZN(n11625) );
  XOR2_X1 U11684 ( .A(n11801), .B(n11802), .Z(n11622) );
  XOR2_X1 U11685 ( .A(n11803), .B(n11804), .Z(n11802) );
  OR2_X1 U11686 ( .A1(n7981), .A2(n8013), .ZN(n11629) );
  XOR2_X1 U11687 ( .A(n11805), .B(n11806), .Z(n11626) );
  XOR2_X1 U11688 ( .A(n11807), .B(n11808), .Z(n11806) );
  OR2_X1 U11689 ( .A1(n7977), .A2(n8013), .ZN(n11633) );
  XOR2_X1 U11690 ( .A(n11809), .B(n11810), .Z(n11630) );
  XOR2_X1 U11691 ( .A(n11811), .B(n11812), .Z(n11810) );
  OR2_X1 U11692 ( .A1(n7974), .A2(n8013), .ZN(n11637) );
  XOR2_X1 U11693 ( .A(n11813), .B(n11814), .Z(n11634) );
  XOR2_X1 U11694 ( .A(n11815), .B(n11816), .Z(n11814) );
  OR2_X1 U11695 ( .A1(n7970), .A2(n8013), .ZN(n11641) );
  XOR2_X1 U11696 ( .A(n11817), .B(n11818), .Z(n11638) );
  XOR2_X1 U11697 ( .A(n11819), .B(n11820), .Z(n11818) );
  OR2_X1 U11698 ( .A1(n7967), .A2(n8013), .ZN(n11645) );
  INV_X1 U11699 ( .A(b_18_), .ZN(n8013) );
  XOR2_X1 U11700 ( .A(n11821), .B(n11822), .Z(n11642) );
  XOR2_X1 U11701 ( .A(n11823), .B(n11824), .Z(n11822) );
  XOR2_X1 U11702 ( .A(n10837), .B(n11825), .Z(n10830) );
  XOR2_X1 U11703 ( .A(n10836), .B(n10835), .Z(n11825) );
  OR2_X1 U11704 ( .A1(n7967), .A2(n7688), .ZN(n10835) );
  OR2_X1 U11705 ( .A1(n11826), .A2(n11827), .ZN(n10836) );
  AND2_X1 U11706 ( .A1(n11824), .A2(n11823), .ZN(n11827) );
  AND2_X1 U11707 ( .A1(n11821), .A2(n11828), .ZN(n11826) );
  OR2_X1 U11708 ( .A1(n11824), .A2(n11823), .ZN(n11828) );
  OR2_X1 U11709 ( .A1(n11829), .A2(n11830), .ZN(n11823) );
  AND2_X1 U11710 ( .A1(n11820), .A2(n11819), .ZN(n11830) );
  AND2_X1 U11711 ( .A1(n11817), .A2(n11831), .ZN(n11829) );
  OR2_X1 U11712 ( .A1(n11820), .A2(n11819), .ZN(n11831) );
  OR2_X1 U11713 ( .A1(n11832), .A2(n11833), .ZN(n11819) );
  AND2_X1 U11714 ( .A1(n11816), .A2(n11815), .ZN(n11833) );
  AND2_X1 U11715 ( .A1(n11813), .A2(n11834), .ZN(n11832) );
  OR2_X1 U11716 ( .A1(n11816), .A2(n11815), .ZN(n11834) );
  OR2_X1 U11717 ( .A1(n11835), .A2(n11836), .ZN(n11815) );
  AND2_X1 U11718 ( .A1(n11812), .A2(n11811), .ZN(n11836) );
  AND2_X1 U11719 ( .A1(n11809), .A2(n11837), .ZN(n11835) );
  OR2_X1 U11720 ( .A1(n11812), .A2(n11811), .ZN(n11837) );
  OR2_X1 U11721 ( .A1(n11838), .A2(n11839), .ZN(n11811) );
  AND2_X1 U11722 ( .A1(n11808), .A2(n11807), .ZN(n11839) );
  AND2_X1 U11723 ( .A1(n11805), .A2(n11840), .ZN(n11838) );
  OR2_X1 U11724 ( .A1(n11808), .A2(n11807), .ZN(n11840) );
  OR2_X1 U11725 ( .A1(n11841), .A2(n11842), .ZN(n11807) );
  AND2_X1 U11726 ( .A1(n11804), .A2(n11803), .ZN(n11842) );
  AND2_X1 U11727 ( .A1(n11801), .A2(n11843), .ZN(n11841) );
  OR2_X1 U11728 ( .A1(n11804), .A2(n11803), .ZN(n11843) );
  OR2_X1 U11729 ( .A1(n11844), .A2(n11845), .ZN(n11803) );
  AND2_X1 U11730 ( .A1(n11800), .A2(n11799), .ZN(n11845) );
  AND2_X1 U11731 ( .A1(n11797), .A2(n11846), .ZN(n11844) );
  OR2_X1 U11732 ( .A1(n11800), .A2(n11799), .ZN(n11846) );
  OR2_X1 U11733 ( .A1(n11847), .A2(n11848), .ZN(n11799) );
  AND2_X1 U11734 ( .A1(n11796), .A2(n11795), .ZN(n11848) );
  AND2_X1 U11735 ( .A1(n11793), .A2(n11849), .ZN(n11847) );
  OR2_X1 U11736 ( .A1(n11796), .A2(n11795), .ZN(n11849) );
  OR2_X1 U11737 ( .A1(n11850), .A2(n11851), .ZN(n11795) );
  AND2_X1 U11738 ( .A1(n11792), .A2(n11791), .ZN(n11851) );
  AND2_X1 U11739 ( .A1(n11789), .A2(n11852), .ZN(n11850) );
  OR2_X1 U11740 ( .A1(n11792), .A2(n11791), .ZN(n11852) );
  OR2_X1 U11741 ( .A1(n11853), .A2(n11854), .ZN(n11791) );
  AND2_X1 U11742 ( .A1(n11788), .A2(n11787), .ZN(n11854) );
  AND2_X1 U11743 ( .A1(n11785), .A2(n11855), .ZN(n11853) );
  OR2_X1 U11744 ( .A1(n11788), .A2(n11787), .ZN(n11855) );
  OR2_X1 U11745 ( .A1(n11856), .A2(n11857), .ZN(n11787) );
  AND2_X1 U11746 ( .A1(n11784), .A2(n11783), .ZN(n11857) );
  AND2_X1 U11747 ( .A1(n11781), .A2(n11858), .ZN(n11856) );
  OR2_X1 U11748 ( .A1(n11784), .A2(n11783), .ZN(n11858) );
  OR2_X1 U11749 ( .A1(n11859), .A2(n11860), .ZN(n11783) );
  AND2_X1 U11750 ( .A1(n8010), .A2(n11780), .ZN(n11860) );
  AND2_X1 U11751 ( .A1(n11778), .A2(n11861), .ZN(n11859) );
  OR2_X1 U11752 ( .A1(n8010), .A2(n11780), .ZN(n11861) );
  OR2_X1 U11753 ( .A1(n11862), .A2(n11863), .ZN(n11780) );
  AND2_X1 U11754 ( .A1(n11777), .A2(n11776), .ZN(n11863) );
  AND2_X1 U11755 ( .A1(n11774), .A2(n11864), .ZN(n11862) );
  OR2_X1 U11756 ( .A1(n11777), .A2(n11776), .ZN(n11864) );
  OR2_X1 U11757 ( .A1(n11865), .A2(n11866), .ZN(n11776) );
  AND2_X1 U11758 ( .A1(n11773), .A2(n11772), .ZN(n11866) );
  AND2_X1 U11759 ( .A1(n11770), .A2(n11867), .ZN(n11865) );
  OR2_X1 U11760 ( .A1(n11773), .A2(n11772), .ZN(n11867) );
  OR2_X1 U11761 ( .A1(n11868), .A2(n11869), .ZN(n11772) );
  AND2_X1 U11762 ( .A1(n11769), .A2(n11768), .ZN(n11869) );
  AND2_X1 U11763 ( .A1(n11766), .A2(n11870), .ZN(n11868) );
  OR2_X1 U11764 ( .A1(n11769), .A2(n11768), .ZN(n11870) );
  OR2_X1 U11765 ( .A1(n11871), .A2(n11872), .ZN(n11768) );
  AND2_X1 U11766 ( .A1(n11765), .A2(n11764), .ZN(n11872) );
  AND2_X1 U11767 ( .A1(n11762), .A2(n11873), .ZN(n11871) );
  OR2_X1 U11768 ( .A1(n11765), .A2(n11764), .ZN(n11873) );
  OR2_X1 U11769 ( .A1(n11874), .A2(n11875), .ZN(n11764) );
  AND2_X1 U11770 ( .A1(n11761), .A2(n11760), .ZN(n11875) );
  AND2_X1 U11771 ( .A1(n11758), .A2(n11876), .ZN(n11874) );
  OR2_X1 U11772 ( .A1(n11761), .A2(n11760), .ZN(n11876) );
  OR2_X1 U11773 ( .A1(n11877), .A2(n11878), .ZN(n11760) );
  AND2_X1 U11774 ( .A1(n11757), .A2(n11756), .ZN(n11878) );
  AND2_X1 U11775 ( .A1(n11754), .A2(n11879), .ZN(n11877) );
  OR2_X1 U11776 ( .A1(n11757), .A2(n11756), .ZN(n11879) );
  OR2_X1 U11777 ( .A1(n11880), .A2(n11881), .ZN(n11756) );
  AND2_X1 U11778 ( .A1(n11753), .A2(n11752), .ZN(n11881) );
  AND2_X1 U11779 ( .A1(n11750), .A2(n11882), .ZN(n11880) );
  OR2_X1 U11780 ( .A1(n11753), .A2(n11752), .ZN(n11882) );
  OR2_X1 U11781 ( .A1(n11883), .A2(n11884), .ZN(n11752) );
  AND2_X1 U11782 ( .A1(n11749), .A2(n11748), .ZN(n11884) );
  AND2_X1 U11783 ( .A1(n11746), .A2(n11885), .ZN(n11883) );
  OR2_X1 U11784 ( .A1(n11749), .A2(n11748), .ZN(n11885) );
  OR2_X1 U11785 ( .A1(n11886), .A2(n11887), .ZN(n11748) );
  AND2_X1 U11786 ( .A1(n11745), .A2(n11744), .ZN(n11887) );
  AND2_X1 U11787 ( .A1(n11742), .A2(n11888), .ZN(n11886) );
  OR2_X1 U11788 ( .A1(n11745), .A2(n11744), .ZN(n11888) );
  OR2_X1 U11789 ( .A1(n11889), .A2(n11890), .ZN(n11744) );
  AND2_X1 U11790 ( .A1(n11741), .A2(n11740), .ZN(n11890) );
  AND2_X1 U11791 ( .A1(n11738), .A2(n11891), .ZN(n11889) );
  OR2_X1 U11792 ( .A1(n11741), .A2(n11740), .ZN(n11891) );
  OR2_X1 U11793 ( .A1(n11892), .A2(n11893), .ZN(n11740) );
  AND2_X1 U11794 ( .A1(n11737), .A2(n11736), .ZN(n11893) );
  AND2_X1 U11795 ( .A1(n11734), .A2(n11894), .ZN(n11892) );
  OR2_X1 U11796 ( .A1(n11737), .A2(n11736), .ZN(n11894) );
  OR2_X1 U11797 ( .A1(n11895), .A2(n11896), .ZN(n11736) );
  AND2_X1 U11798 ( .A1(n11730), .A2(n11897), .ZN(n11896) );
  AND2_X1 U11799 ( .A1(n11898), .A2(n11899), .ZN(n11895) );
  OR2_X1 U11800 ( .A1(n11730), .A2(n11897), .ZN(n11899) );
  INV_X1 U11801 ( .A(n11733), .ZN(n11897) );
  AND3_X1 U11802 ( .A1(n8904), .A2(b_16_), .A3(b_17_), .ZN(n11733) );
  OR2_X1 U11803 ( .A1(n8051), .A2(n7688), .ZN(n11730) );
  INV_X1 U11804 ( .A(n11732), .ZN(n11898) );
  OR2_X1 U11805 ( .A1(n11900), .A2(n11901), .ZN(n11732) );
  AND2_X1 U11806 ( .A1(b_16_), .A2(n11902), .ZN(n11901) );
  OR2_X1 U11807 ( .A1(n11903), .A2(n7490), .ZN(n11902) );
  AND2_X1 U11808 ( .A1(a_30_), .A2(n7717), .ZN(n11903) );
  AND2_X1 U11809 ( .A1(b_15_), .A2(n11904), .ZN(n11900) );
  OR2_X1 U11810 ( .A1(n11905), .A2(n7493), .ZN(n11904) );
  AND2_X1 U11811 ( .A1(a_31_), .A2(n8006), .ZN(n11905) );
  OR2_X1 U11812 ( .A1(n8048), .A2(n7688), .ZN(n11737) );
  XNOR2_X1 U11813 ( .A(n11906), .B(n11907), .ZN(n11734) );
  XNOR2_X1 U11814 ( .A(n11908), .B(n11909), .ZN(n11907) );
  OR2_X1 U11815 ( .A1(n8044), .A2(n7688), .ZN(n11741) );
  XOR2_X1 U11816 ( .A(n11910), .B(n11911), .Z(n11738) );
  XOR2_X1 U11817 ( .A(n11912), .B(n11913), .Z(n11911) );
  OR2_X1 U11818 ( .A1(n8041), .A2(n7688), .ZN(n11745) );
  XOR2_X1 U11819 ( .A(n11914), .B(n11915), .Z(n11742) );
  XOR2_X1 U11820 ( .A(n11916), .B(n11917), .Z(n11915) );
  OR2_X1 U11821 ( .A1(n8037), .A2(n7688), .ZN(n11749) );
  XOR2_X1 U11822 ( .A(n11918), .B(n11919), .Z(n11746) );
  XOR2_X1 U11823 ( .A(n11920), .B(n11921), .Z(n11919) );
  OR2_X1 U11824 ( .A1(n8034), .A2(n7688), .ZN(n11753) );
  XOR2_X1 U11825 ( .A(n11922), .B(n11923), .Z(n11750) );
  XOR2_X1 U11826 ( .A(n11924), .B(n11925), .Z(n11923) );
  OR2_X1 U11827 ( .A1(n8030), .A2(n7688), .ZN(n11757) );
  XOR2_X1 U11828 ( .A(n11926), .B(n11927), .Z(n11754) );
  XOR2_X1 U11829 ( .A(n11928), .B(n11929), .Z(n11927) );
  OR2_X1 U11830 ( .A1(n8026), .A2(n7688), .ZN(n11761) );
  XOR2_X1 U11831 ( .A(n11930), .B(n11931), .Z(n11758) );
  XOR2_X1 U11832 ( .A(n11932), .B(n11933), .Z(n11931) );
  OR2_X1 U11833 ( .A1(n8023), .A2(n7688), .ZN(n11765) );
  XOR2_X1 U11834 ( .A(n11934), .B(n11935), .Z(n11762) );
  XOR2_X1 U11835 ( .A(n11936), .B(n11937), .Z(n11935) );
  OR2_X1 U11836 ( .A1(n8019), .A2(n7688), .ZN(n11769) );
  XOR2_X1 U11837 ( .A(n11938), .B(n11939), .Z(n11766) );
  XOR2_X1 U11838 ( .A(n11940), .B(n11941), .Z(n11939) );
  OR2_X1 U11839 ( .A1(n8016), .A2(n7688), .ZN(n11773) );
  XOR2_X1 U11840 ( .A(n11942), .B(n11943), .Z(n11770) );
  XOR2_X1 U11841 ( .A(n11944), .B(n11945), .Z(n11943) );
  OR2_X1 U11842 ( .A1(n8012), .A2(n7688), .ZN(n11777) );
  XOR2_X1 U11843 ( .A(n11946), .B(n11947), .Z(n11774) );
  XOR2_X1 U11844 ( .A(n11948), .B(n11949), .Z(n11947) );
  INV_X1 U11845 ( .A(n7692), .ZN(n8010) );
  AND2_X1 U11846 ( .A1(a_17_), .A2(b_17_), .ZN(n7692) );
  XOR2_X1 U11847 ( .A(n11950), .B(n11951), .Z(n11778) );
  XOR2_X1 U11848 ( .A(n11952), .B(n11953), .Z(n11951) );
  OR2_X1 U11849 ( .A1(n8005), .A2(n7688), .ZN(n11784) );
  XOR2_X1 U11850 ( .A(n11954), .B(n11955), .Z(n11781) );
  XOR2_X1 U11851 ( .A(n11956), .B(n11957), .Z(n11955) );
  OR2_X1 U11852 ( .A1(n8002), .A2(n7688), .ZN(n11788) );
  XNOR2_X1 U11853 ( .A(n11958), .B(n11959), .ZN(n11785) );
  XNOR2_X1 U11854 ( .A(n8007), .B(n11960), .ZN(n11958) );
  OR2_X1 U11855 ( .A1(n7998), .A2(n7688), .ZN(n11792) );
  XOR2_X1 U11856 ( .A(n11961), .B(n11962), .Z(n11789) );
  XOR2_X1 U11857 ( .A(n11963), .B(n11964), .Z(n11962) );
  OR2_X1 U11858 ( .A1(n7995), .A2(n7688), .ZN(n11796) );
  XOR2_X1 U11859 ( .A(n11965), .B(n11966), .Z(n11793) );
  XOR2_X1 U11860 ( .A(n11967), .B(n11968), .Z(n11966) );
  OR2_X1 U11861 ( .A1(n7991), .A2(n7688), .ZN(n11800) );
  XOR2_X1 U11862 ( .A(n11969), .B(n11970), .Z(n11797) );
  XOR2_X1 U11863 ( .A(n11971), .B(n11972), .Z(n11970) );
  OR2_X1 U11864 ( .A1(n7988), .A2(n7688), .ZN(n11804) );
  XOR2_X1 U11865 ( .A(n11973), .B(n11974), .Z(n11801) );
  XOR2_X1 U11866 ( .A(n11975), .B(n11976), .Z(n11974) );
  OR2_X1 U11867 ( .A1(n7984), .A2(n7688), .ZN(n11808) );
  XOR2_X1 U11868 ( .A(n11977), .B(n11978), .Z(n11805) );
  XOR2_X1 U11869 ( .A(n11979), .B(n11980), .Z(n11978) );
  OR2_X1 U11870 ( .A1(n7981), .A2(n7688), .ZN(n11812) );
  XOR2_X1 U11871 ( .A(n11981), .B(n11982), .Z(n11809) );
  XOR2_X1 U11872 ( .A(n11983), .B(n11984), .Z(n11982) );
  OR2_X1 U11873 ( .A1(n7977), .A2(n7688), .ZN(n11816) );
  XOR2_X1 U11874 ( .A(n11985), .B(n11986), .Z(n11813) );
  XOR2_X1 U11875 ( .A(n11987), .B(n11988), .Z(n11986) );
  OR2_X1 U11876 ( .A1(n7974), .A2(n7688), .ZN(n11820) );
  XOR2_X1 U11877 ( .A(n11989), .B(n11990), .Z(n11817) );
  XOR2_X1 U11878 ( .A(n11991), .B(n11992), .Z(n11990) );
  OR2_X1 U11879 ( .A1(n7970), .A2(n7688), .ZN(n11824) );
  INV_X1 U11880 ( .A(b_17_), .ZN(n7688) );
  XOR2_X1 U11881 ( .A(n11993), .B(n11994), .Z(n11821) );
  XOR2_X1 U11882 ( .A(n11995), .B(n11996), .Z(n11994) );
  XOR2_X1 U11883 ( .A(n10844), .B(n11997), .Z(n10837) );
  XOR2_X1 U11884 ( .A(n10843), .B(n10842), .Z(n11997) );
  OR2_X1 U11885 ( .A1(n7970), .A2(n8006), .ZN(n10842) );
  OR2_X1 U11886 ( .A1(n11998), .A2(n11999), .ZN(n10843) );
  AND2_X1 U11887 ( .A1(n11996), .A2(n11995), .ZN(n11999) );
  AND2_X1 U11888 ( .A1(n11993), .A2(n12000), .ZN(n11998) );
  OR2_X1 U11889 ( .A1(n11996), .A2(n11995), .ZN(n12000) );
  OR2_X1 U11890 ( .A1(n12001), .A2(n12002), .ZN(n11995) );
  AND2_X1 U11891 ( .A1(n11992), .A2(n11991), .ZN(n12002) );
  AND2_X1 U11892 ( .A1(n11989), .A2(n12003), .ZN(n12001) );
  OR2_X1 U11893 ( .A1(n11992), .A2(n11991), .ZN(n12003) );
  OR2_X1 U11894 ( .A1(n12004), .A2(n12005), .ZN(n11991) );
  AND2_X1 U11895 ( .A1(n11988), .A2(n11987), .ZN(n12005) );
  AND2_X1 U11896 ( .A1(n11985), .A2(n12006), .ZN(n12004) );
  OR2_X1 U11897 ( .A1(n11988), .A2(n11987), .ZN(n12006) );
  OR2_X1 U11898 ( .A1(n12007), .A2(n12008), .ZN(n11987) );
  AND2_X1 U11899 ( .A1(n11984), .A2(n11983), .ZN(n12008) );
  AND2_X1 U11900 ( .A1(n11981), .A2(n12009), .ZN(n12007) );
  OR2_X1 U11901 ( .A1(n11984), .A2(n11983), .ZN(n12009) );
  OR2_X1 U11902 ( .A1(n12010), .A2(n12011), .ZN(n11983) );
  AND2_X1 U11903 ( .A1(n11980), .A2(n11979), .ZN(n12011) );
  AND2_X1 U11904 ( .A1(n11977), .A2(n12012), .ZN(n12010) );
  OR2_X1 U11905 ( .A1(n11980), .A2(n11979), .ZN(n12012) );
  OR2_X1 U11906 ( .A1(n12013), .A2(n12014), .ZN(n11979) );
  AND2_X1 U11907 ( .A1(n11976), .A2(n11975), .ZN(n12014) );
  AND2_X1 U11908 ( .A1(n11973), .A2(n12015), .ZN(n12013) );
  OR2_X1 U11909 ( .A1(n11976), .A2(n11975), .ZN(n12015) );
  OR2_X1 U11910 ( .A1(n12016), .A2(n12017), .ZN(n11975) );
  AND2_X1 U11911 ( .A1(n11969), .A2(n11972), .ZN(n12017) );
  AND2_X1 U11912 ( .A1(n12018), .A2(n11971), .ZN(n12016) );
  OR2_X1 U11913 ( .A1(n12019), .A2(n12020), .ZN(n11971) );
  AND2_X1 U11914 ( .A1(n11968), .A2(n11967), .ZN(n12020) );
  AND2_X1 U11915 ( .A1(n11965), .A2(n12021), .ZN(n12019) );
  OR2_X1 U11916 ( .A1(n11968), .A2(n11967), .ZN(n12021) );
  OR2_X1 U11917 ( .A1(n12022), .A2(n12023), .ZN(n11967) );
  AND2_X1 U11918 ( .A1(n11961), .A2(n11964), .ZN(n12023) );
  AND2_X1 U11919 ( .A1(n12024), .A2(n11963), .ZN(n12022) );
  OR2_X1 U11920 ( .A1(n12025), .A2(n12026), .ZN(n11963) );
  AND2_X1 U11921 ( .A1(n11959), .A2(n8007), .ZN(n12026) );
  AND2_X1 U11922 ( .A1(n12027), .A2(n11960), .ZN(n12025) );
  OR2_X1 U11923 ( .A1(n12028), .A2(n12029), .ZN(n11960) );
  AND2_X1 U11924 ( .A1(n11954), .A2(n11957), .ZN(n12029) );
  AND2_X1 U11925 ( .A1(n12030), .A2(n11956), .ZN(n12028) );
  OR2_X1 U11926 ( .A1(n12031), .A2(n12032), .ZN(n11956) );
  AND2_X1 U11927 ( .A1(n11950), .A2(n11953), .ZN(n12032) );
  AND2_X1 U11928 ( .A1(n12033), .A2(n11952), .ZN(n12031) );
  OR2_X1 U11929 ( .A1(n12034), .A2(n12035), .ZN(n11952) );
  AND2_X1 U11930 ( .A1(n11946), .A2(n11949), .ZN(n12035) );
  AND2_X1 U11931 ( .A1(n12036), .A2(n11948), .ZN(n12034) );
  OR2_X1 U11932 ( .A1(n12037), .A2(n12038), .ZN(n11948) );
  AND2_X1 U11933 ( .A1(n11942), .A2(n11945), .ZN(n12038) );
  AND2_X1 U11934 ( .A1(n12039), .A2(n11944), .ZN(n12037) );
  OR2_X1 U11935 ( .A1(n12040), .A2(n12041), .ZN(n11944) );
  AND2_X1 U11936 ( .A1(n11938), .A2(n11941), .ZN(n12041) );
  AND2_X1 U11937 ( .A1(n12042), .A2(n11940), .ZN(n12040) );
  OR2_X1 U11938 ( .A1(n12043), .A2(n12044), .ZN(n11940) );
  AND2_X1 U11939 ( .A1(n11934), .A2(n11937), .ZN(n12044) );
  AND2_X1 U11940 ( .A1(n12045), .A2(n11936), .ZN(n12043) );
  OR2_X1 U11941 ( .A1(n12046), .A2(n12047), .ZN(n11936) );
  AND2_X1 U11942 ( .A1(n11930), .A2(n11933), .ZN(n12047) );
  AND2_X1 U11943 ( .A1(n12048), .A2(n11932), .ZN(n12046) );
  OR2_X1 U11944 ( .A1(n12049), .A2(n12050), .ZN(n11932) );
  AND2_X1 U11945 ( .A1(n11926), .A2(n11929), .ZN(n12050) );
  AND2_X1 U11946 ( .A1(n12051), .A2(n11928), .ZN(n12049) );
  OR2_X1 U11947 ( .A1(n12052), .A2(n12053), .ZN(n11928) );
  AND2_X1 U11948 ( .A1(n11922), .A2(n11925), .ZN(n12053) );
  AND2_X1 U11949 ( .A1(n12054), .A2(n11924), .ZN(n12052) );
  OR2_X1 U11950 ( .A1(n12055), .A2(n12056), .ZN(n11924) );
  AND2_X1 U11951 ( .A1(n11918), .A2(n11921), .ZN(n12056) );
  AND2_X1 U11952 ( .A1(n12057), .A2(n11920), .ZN(n12055) );
  OR2_X1 U11953 ( .A1(n12058), .A2(n12059), .ZN(n11920) );
  AND2_X1 U11954 ( .A1(n11914), .A2(n11917), .ZN(n12059) );
  AND2_X1 U11955 ( .A1(n12060), .A2(n11916), .ZN(n12058) );
  OR2_X1 U11956 ( .A1(n12061), .A2(n12062), .ZN(n11916) );
  AND2_X1 U11957 ( .A1(n11910), .A2(n11913), .ZN(n12062) );
  AND2_X1 U11958 ( .A1(n12063), .A2(n11912), .ZN(n12061) );
  OR2_X1 U11959 ( .A1(n12064), .A2(n12065), .ZN(n11912) );
  AND2_X1 U11960 ( .A1(n11906), .A2(n12066), .ZN(n12065) );
  AND2_X1 U11961 ( .A1(n12067), .A2(n12068), .ZN(n12064) );
  OR2_X1 U11962 ( .A1(n11906), .A2(n12066), .ZN(n12068) );
  INV_X1 U11963 ( .A(n11909), .ZN(n12066) );
  AND3_X1 U11964 ( .A1(n8904), .A2(b_15_), .A3(b_16_), .ZN(n11909) );
  OR2_X1 U11965 ( .A1(n8051), .A2(n8006), .ZN(n11906) );
  INV_X1 U11966 ( .A(n11908), .ZN(n12067) );
  OR2_X1 U11967 ( .A1(n12069), .A2(n12070), .ZN(n11908) );
  AND2_X1 U11968 ( .A1(b_15_), .A2(n12071), .ZN(n12070) );
  OR2_X1 U11969 ( .A1(n12072), .A2(n7490), .ZN(n12071) );
  AND2_X1 U11970 ( .A1(a_30_), .A2(n7999), .ZN(n12072) );
  AND2_X1 U11971 ( .A1(b_14_), .A2(n12073), .ZN(n12069) );
  OR2_X1 U11972 ( .A1(n12074), .A2(n7493), .ZN(n12073) );
  AND2_X1 U11973 ( .A1(a_31_), .A2(n7717), .ZN(n12074) );
  OR2_X1 U11974 ( .A1(n11910), .A2(n11913), .ZN(n12063) );
  OR2_X1 U11975 ( .A1(n8048), .A2(n8006), .ZN(n11913) );
  XNOR2_X1 U11976 ( .A(n12075), .B(n12076), .ZN(n11910) );
  XNOR2_X1 U11977 ( .A(n12077), .B(n12078), .ZN(n12076) );
  OR2_X1 U11978 ( .A1(n11914), .A2(n11917), .ZN(n12060) );
  OR2_X1 U11979 ( .A1(n8044), .A2(n8006), .ZN(n11917) );
  XOR2_X1 U11980 ( .A(n12079), .B(n12080), .Z(n11914) );
  XOR2_X1 U11981 ( .A(n12081), .B(n12082), .Z(n12080) );
  OR2_X1 U11982 ( .A1(n11918), .A2(n11921), .ZN(n12057) );
  OR2_X1 U11983 ( .A1(n8041), .A2(n8006), .ZN(n11921) );
  XOR2_X1 U11984 ( .A(n12083), .B(n12084), .Z(n11918) );
  XOR2_X1 U11985 ( .A(n12085), .B(n12086), .Z(n12084) );
  OR2_X1 U11986 ( .A1(n11922), .A2(n11925), .ZN(n12054) );
  OR2_X1 U11987 ( .A1(n8037), .A2(n8006), .ZN(n11925) );
  XOR2_X1 U11988 ( .A(n12087), .B(n12088), .Z(n11922) );
  XOR2_X1 U11989 ( .A(n12089), .B(n12090), .Z(n12088) );
  OR2_X1 U11990 ( .A1(n11926), .A2(n11929), .ZN(n12051) );
  OR2_X1 U11991 ( .A1(n8034), .A2(n8006), .ZN(n11929) );
  XOR2_X1 U11992 ( .A(n12091), .B(n12092), .Z(n11926) );
  XOR2_X1 U11993 ( .A(n12093), .B(n12094), .Z(n12092) );
  OR2_X1 U11994 ( .A1(n11930), .A2(n11933), .ZN(n12048) );
  OR2_X1 U11995 ( .A1(n8030), .A2(n8006), .ZN(n11933) );
  XOR2_X1 U11996 ( .A(n12095), .B(n12096), .Z(n11930) );
  XOR2_X1 U11997 ( .A(n12097), .B(n12098), .Z(n12096) );
  OR2_X1 U11998 ( .A1(n11934), .A2(n11937), .ZN(n12045) );
  OR2_X1 U11999 ( .A1(n8026), .A2(n8006), .ZN(n11937) );
  XOR2_X1 U12000 ( .A(n12099), .B(n12100), .Z(n11934) );
  XOR2_X1 U12001 ( .A(n12101), .B(n12102), .Z(n12100) );
  OR2_X1 U12002 ( .A1(n11938), .A2(n11941), .ZN(n12042) );
  OR2_X1 U12003 ( .A1(n8023), .A2(n8006), .ZN(n11941) );
  XOR2_X1 U12004 ( .A(n12103), .B(n12104), .Z(n11938) );
  XOR2_X1 U12005 ( .A(n12105), .B(n12106), .Z(n12104) );
  OR2_X1 U12006 ( .A1(n11942), .A2(n11945), .ZN(n12039) );
  OR2_X1 U12007 ( .A1(n8019), .A2(n8006), .ZN(n11945) );
  XOR2_X1 U12008 ( .A(n12107), .B(n12108), .Z(n11942) );
  XOR2_X1 U12009 ( .A(n12109), .B(n12110), .Z(n12108) );
  OR2_X1 U12010 ( .A1(n11946), .A2(n11949), .ZN(n12036) );
  OR2_X1 U12011 ( .A1(n8016), .A2(n8006), .ZN(n11949) );
  XOR2_X1 U12012 ( .A(n12111), .B(n12112), .Z(n11946) );
  XOR2_X1 U12013 ( .A(n12113), .B(n12114), .Z(n12112) );
  OR2_X1 U12014 ( .A1(n11950), .A2(n11953), .ZN(n12033) );
  OR2_X1 U12015 ( .A1(n8012), .A2(n8006), .ZN(n11953) );
  XOR2_X1 U12016 ( .A(n12115), .B(n12116), .Z(n11950) );
  XOR2_X1 U12017 ( .A(n12117), .B(n12118), .Z(n12116) );
  OR2_X1 U12018 ( .A1(n11954), .A2(n11957), .ZN(n12030) );
  OR2_X1 U12019 ( .A1(n8009), .A2(n8006), .ZN(n11957) );
  XOR2_X1 U12020 ( .A(n12119), .B(n12120), .Z(n11954) );
  XOR2_X1 U12021 ( .A(n12121), .B(n12122), .Z(n12120) );
  OR2_X1 U12022 ( .A1(n11959), .A2(n8007), .ZN(n12027) );
  INV_X1 U12023 ( .A(n7709), .ZN(n8007) );
  AND2_X1 U12024 ( .A1(a_16_), .A2(b_16_), .ZN(n7709) );
  XOR2_X1 U12025 ( .A(n12123), .B(n12124), .Z(n11959) );
  XOR2_X1 U12026 ( .A(n12125), .B(n12126), .Z(n12124) );
  OR2_X1 U12027 ( .A1(n11961), .A2(n11964), .ZN(n12024) );
  OR2_X1 U12028 ( .A1(n8002), .A2(n8006), .ZN(n11964) );
  XOR2_X1 U12029 ( .A(n12127), .B(n12128), .Z(n11961) );
  XOR2_X1 U12030 ( .A(n12129), .B(n12130), .Z(n12128) );
  OR2_X1 U12031 ( .A1(n7998), .A2(n8006), .ZN(n11968) );
  XOR2_X1 U12032 ( .A(n12131), .B(n12132), .Z(n11965) );
  XNOR2_X1 U12033 ( .A(n12133), .B(n7721), .ZN(n12132) );
  OR2_X1 U12034 ( .A1(n11969), .A2(n11972), .ZN(n12018) );
  OR2_X1 U12035 ( .A1(n7995), .A2(n8006), .ZN(n11972) );
  XOR2_X1 U12036 ( .A(n12134), .B(n12135), .Z(n11969) );
  XOR2_X1 U12037 ( .A(n12136), .B(n12137), .Z(n12135) );
  OR2_X1 U12038 ( .A1(n7991), .A2(n8006), .ZN(n11976) );
  XOR2_X1 U12039 ( .A(n12138), .B(n12139), .Z(n11973) );
  XOR2_X1 U12040 ( .A(n12140), .B(n12141), .Z(n12139) );
  OR2_X1 U12041 ( .A1(n7988), .A2(n8006), .ZN(n11980) );
  XOR2_X1 U12042 ( .A(n12142), .B(n12143), .Z(n11977) );
  XOR2_X1 U12043 ( .A(n12144), .B(n12145), .Z(n12143) );
  OR2_X1 U12044 ( .A1(n7984), .A2(n8006), .ZN(n11984) );
  XOR2_X1 U12045 ( .A(n12146), .B(n12147), .Z(n11981) );
  XOR2_X1 U12046 ( .A(n12148), .B(n12149), .Z(n12147) );
  OR2_X1 U12047 ( .A1(n7981), .A2(n8006), .ZN(n11988) );
  XOR2_X1 U12048 ( .A(n12150), .B(n12151), .Z(n11985) );
  XOR2_X1 U12049 ( .A(n12152), .B(n12153), .Z(n12151) );
  OR2_X1 U12050 ( .A1(n7977), .A2(n8006), .ZN(n11992) );
  XOR2_X1 U12051 ( .A(n12154), .B(n12155), .Z(n11989) );
  XOR2_X1 U12052 ( .A(n12156), .B(n12157), .Z(n12155) );
  OR2_X1 U12053 ( .A1(n7974), .A2(n8006), .ZN(n11996) );
  INV_X1 U12054 ( .A(b_16_), .ZN(n8006) );
  XOR2_X1 U12055 ( .A(n12158), .B(n12159), .Z(n11993) );
  XOR2_X1 U12056 ( .A(n12160), .B(n12161), .Z(n12159) );
  XOR2_X1 U12057 ( .A(n10851), .B(n12162), .Z(n10844) );
  XOR2_X1 U12058 ( .A(n10850), .B(n10849), .Z(n12162) );
  OR2_X1 U12059 ( .A1(n7974), .A2(n7717), .ZN(n10849) );
  OR2_X1 U12060 ( .A1(n12163), .A2(n12164), .ZN(n10850) );
  AND2_X1 U12061 ( .A1(n12161), .A2(n12160), .ZN(n12164) );
  AND2_X1 U12062 ( .A1(n12158), .A2(n12165), .ZN(n12163) );
  OR2_X1 U12063 ( .A1(n12160), .A2(n12161), .ZN(n12165) );
  OR2_X1 U12064 ( .A1(n7977), .A2(n7717), .ZN(n12161) );
  OR2_X1 U12065 ( .A1(n12166), .A2(n12167), .ZN(n12160) );
  AND2_X1 U12066 ( .A1(n12157), .A2(n12156), .ZN(n12167) );
  AND2_X1 U12067 ( .A1(n12154), .A2(n12168), .ZN(n12166) );
  OR2_X1 U12068 ( .A1(n12156), .A2(n12157), .ZN(n12168) );
  OR2_X1 U12069 ( .A1(n7981), .A2(n7717), .ZN(n12157) );
  OR2_X1 U12070 ( .A1(n12169), .A2(n12170), .ZN(n12156) );
  AND2_X1 U12071 ( .A1(n12153), .A2(n12152), .ZN(n12170) );
  AND2_X1 U12072 ( .A1(n12150), .A2(n12171), .ZN(n12169) );
  OR2_X1 U12073 ( .A1(n12152), .A2(n12153), .ZN(n12171) );
  OR2_X1 U12074 ( .A1(n7984), .A2(n7717), .ZN(n12153) );
  OR2_X1 U12075 ( .A1(n12172), .A2(n12173), .ZN(n12152) );
  AND2_X1 U12076 ( .A1(n12149), .A2(n12148), .ZN(n12173) );
  AND2_X1 U12077 ( .A1(n12146), .A2(n12174), .ZN(n12172) );
  OR2_X1 U12078 ( .A1(n12148), .A2(n12149), .ZN(n12174) );
  OR2_X1 U12079 ( .A1(n7988), .A2(n7717), .ZN(n12149) );
  OR2_X1 U12080 ( .A1(n12175), .A2(n12176), .ZN(n12148) );
  AND2_X1 U12081 ( .A1(n12145), .A2(n12144), .ZN(n12176) );
  AND2_X1 U12082 ( .A1(n12142), .A2(n12177), .ZN(n12175) );
  OR2_X1 U12083 ( .A1(n12144), .A2(n12145), .ZN(n12177) );
  OR2_X1 U12084 ( .A1(n7991), .A2(n7717), .ZN(n12145) );
  OR2_X1 U12085 ( .A1(n12178), .A2(n12179), .ZN(n12144) );
  AND2_X1 U12086 ( .A1(n12141), .A2(n12140), .ZN(n12179) );
  AND2_X1 U12087 ( .A1(n12138), .A2(n12180), .ZN(n12178) );
  OR2_X1 U12088 ( .A1(n12140), .A2(n12141), .ZN(n12180) );
  OR2_X1 U12089 ( .A1(n7995), .A2(n7717), .ZN(n12141) );
  OR2_X1 U12090 ( .A1(n12181), .A2(n12182), .ZN(n12140) );
  AND2_X1 U12091 ( .A1(n12137), .A2(n12136), .ZN(n12182) );
  AND2_X1 U12092 ( .A1(n12134), .A2(n12183), .ZN(n12181) );
  OR2_X1 U12093 ( .A1(n12136), .A2(n12137), .ZN(n12183) );
  OR2_X1 U12094 ( .A1(n7998), .A2(n7717), .ZN(n12137) );
  OR2_X1 U12095 ( .A1(n12184), .A2(n12185), .ZN(n12136) );
  AND2_X1 U12096 ( .A1(n8003), .A2(n12133), .ZN(n12185) );
  AND2_X1 U12097 ( .A1(n12131), .A2(n12186), .ZN(n12184) );
  OR2_X1 U12098 ( .A1(n12133), .A2(n8003), .ZN(n12186) );
  INV_X1 U12099 ( .A(n7721), .ZN(n8003) );
  AND2_X1 U12100 ( .A1(a_15_), .A2(b_15_), .ZN(n7721) );
  OR2_X1 U12101 ( .A1(n12187), .A2(n12188), .ZN(n12133) );
  AND2_X1 U12102 ( .A1(n12130), .A2(n12129), .ZN(n12188) );
  AND2_X1 U12103 ( .A1(n12127), .A2(n12189), .ZN(n12187) );
  OR2_X1 U12104 ( .A1(n12129), .A2(n12130), .ZN(n12189) );
  OR2_X1 U12105 ( .A1(n8005), .A2(n7717), .ZN(n12130) );
  OR2_X1 U12106 ( .A1(n12190), .A2(n12191), .ZN(n12129) );
  AND2_X1 U12107 ( .A1(n12126), .A2(n12125), .ZN(n12191) );
  AND2_X1 U12108 ( .A1(n12123), .A2(n12192), .ZN(n12190) );
  OR2_X1 U12109 ( .A1(n12125), .A2(n12126), .ZN(n12192) );
  OR2_X1 U12110 ( .A1(n8009), .A2(n7717), .ZN(n12126) );
  OR2_X1 U12111 ( .A1(n12193), .A2(n12194), .ZN(n12125) );
  AND2_X1 U12112 ( .A1(n12122), .A2(n12121), .ZN(n12194) );
  AND2_X1 U12113 ( .A1(n12119), .A2(n12195), .ZN(n12193) );
  OR2_X1 U12114 ( .A1(n12121), .A2(n12122), .ZN(n12195) );
  OR2_X1 U12115 ( .A1(n8012), .A2(n7717), .ZN(n12122) );
  OR2_X1 U12116 ( .A1(n12196), .A2(n12197), .ZN(n12121) );
  AND2_X1 U12117 ( .A1(n12118), .A2(n12117), .ZN(n12197) );
  AND2_X1 U12118 ( .A1(n12115), .A2(n12198), .ZN(n12196) );
  OR2_X1 U12119 ( .A1(n12117), .A2(n12118), .ZN(n12198) );
  OR2_X1 U12120 ( .A1(n8016), .A2(n7717), .ZN(n12118) );
  OR2_X1 U12121 ( .A1(n12199), .A2(n12200), .ZN(n12117) );
  AND2_X1 U12122 ( .A1(n12114), .A2(n12113), .ZN(n12200) );
  AND2_X1 U12123 ( .A1(n12111), .A2(n12201), .ZN(n12199) );
  OR2_X1 U12124 ( .A1(n12113), .A2(n12114), .ZN(n12201) );
  OR2_X1 U12125 ( .A1(n8019), .A2(n7717), .ZN(n12114) );
  OR2_X1 U12126 ( .A1(n12202), .A2(n12203), .ZN(n12113) );
  AND2_X1 U12127 ( .A1(n12110), .A2(n12109), .ZN(n12203) );
  AND2_X1 U12128 ( .A1(n12107), .A2(n12204), .ZN(n12202) );
  OR2_X1 U12129 ( .A1(n12109), .A2(n12110), .ZN(n12204) );
  OR2_X1 U12130 ( .A1(n8023), .A2(n7717), .ZN(n12110) );
  OR2_X1 U12131 ( .A1(n12205), .A2(n12206), .ZN(n12109) );
  AND2_X1 U12132 ( .A1(n12106), .A2(n12105), .ZN(n12206) );
  AND2_X1 U12133 ( .A1(n12103), .A2(n12207), .ZN(n12205) );
  OR2_X1 U12134 ( .A1(n12105), .A2(n12106), .ZN(n12207) );
  OR2_X1 U12135 ( .A1(n8026), .A2(n7717), .ZN(n12106) );
  OR2_X1 U12136 ( .A1(n12208), .A2(n12209), .ZN(n12105) );
  AND2_X1 U12137 ( .A1(n12102), .A2(n12101), .ZN(n12209) );
  AND2_X1 U12138 ( .A1(n12099), .A2(n12210), .ZN(n12208) );
  OR2_X1 U12139 ( .A1(n12101), .A2(n12102), .ZN(n12210) );
  OR2_X1 U12140 ( .A1(n8030), .A2(n7717), .ZN(n12102) );
  OR2_X1 U12141 ( .A1(n12211), .A2(n12212), .ZN(n12101) );
  AND2_X1 U12142 ( .A1(n12098), .A2(n12097), .ZN(n12212) );
  AND2_X1 U12143 ( .A1(n12095), .A2(n12213), .ZN(n12211) );
  OR2_X1 U12144 ( .A1(n12097), .A2(n12098), .ZN(n12213) );
  OR2_X1 U12145 ( .A1(n8034), .A2(n7717), .ZN(n12098) );
  OR2_X1 U12146 ( .A1(n12214), .A2(n12215), .ZN(n12097) );
  AND2_X1 U12147 ( .A1(n12094), .A2(n12093), .ZN(n12215) );
  AND2_X1 U12148 ( .A1(n12091), .A2(n12216), .ZN(n12214) );
  OR2_X1 U12149 ( .A1(n12093), .A2(n12094), .ZN(n12216) );
  OR2_X1 U12150 ( .A1(n8037), .A2(n7717), .ZN(n12094) );
  OR2_X1 U12151 ( .A1(n12217), .A2(n12218), .ZN(n12093) );
  AND2_X1 U12152 ( .A1(n12090), .A2(n12089), .ZN(n12218) );
  AND2_X1 U12153 ( .A1(n12087), .A2(n12219), .ZN(n12217) );
  OR2_X1 U12154 ( .A1(n12089), .A2(n12090), .ZN(n12219) );
  OR2_X1 U12155 ( .A1(n8041), .A2(n7717), .ZN(n12090) );
  OR2_X1 U12156 ( .A1(n12220), .A2(n12221), .ZN(n12089) );
  AND2_X1 U12157 ( .A1(n12086), .A2(n12085), .ZN(n12221) );
  AND2_X1 U12158 ( .A1(n12083), .A2(n12222), .ZN(n12220) );
  OR2_X1 U12159 ( .A1(n12085), .A2(n12086), .ZN(n12222) );
  OR2_X1 U12160 ( .A1(n8044), .A2(n7717), .ZN(n12086) );
  OR2_X1 U12161 ( .A1(n12223), .A2(n12224), .ZN(n12085) );
  AND2_X1 U12162 ( .A1(n12082), .A2(n12081), .ZN(n12224) );
  AND2_X1 U12163 ( .A1(n12079), .A2(n12225), .ZN(n12223) );
  OR2_X1 U12164 ( .A1(n12081), .A2(n12082), .ZN(n12225) );
  OR2_X1 U12165 ( .A1(n8048), .A2(n7717), .ZN(n12082) );
  OR2_X1 U12166 ( .A1(n12226), .A2(n12227), .ZN(n12081) );
  AND2_X1 U12167 ( .A1(n12075), .A2(n12228), .ZN(n12227) );
  AND2_X1 U12168 ( .A1(n12229), .A2(n12230), .ZN(n12226) );
  OR2_X1 U12169 ( .A1(n12228), .A2(n12075), .ZN(n12230) );
  OR2_X1 U12170 ( .A1(n8051), .A2(n7717), .ZN(n12075) );
  INV_X1 U12171 ( .A(b_15_), .ZN(n7717) );
  INV_X1 U12172 ( .A(n12078), .ZN(n12228) );
  AND3_X1 U12173 ( .A1(n8904), .A2(b_14_), .A3(b_15_), .ZN(n12078) );
  INV_X1 U12174 ( .A(n12077), .ZN(n12229) );
  OR2_X1 U12175 ( .A1(n12231), .A2(n12232), .ZN(n12077) );
  AND2_X1 U12176 ( .A1(b_14_), .A2(n12233), .ZN(n12232) );
  OR2_X1 U12177 ( .A1(n12234), .A2(n7490), .ZN(n12233) );
  AND2_X1 U12178 ( .A1(a_30_), .A2(n7746), .ZN(n12234) );
  AND2_X1 U12179 ( .A1(b_13_), .A2(n12235), .ZN(n12231) );
  OR2_X1 U12180 ( .A1(n12236), .A2(n7493), .ZN(n12235) );
  AND2_X1 U12181 ( .A1(a_31_), .A2(n7999), .ZN(n12236) );
  XNOR2_X1 U12182 ( .A(n12237), .B(n12238), .ZN(n12079) );
  XNOR2_X1 U12183 ( .A(n12239), .B(n12240), .ZN(n12238) );
  XOR2_X1 U12184 ( .A(n12241), .B(n12242), .Z(n12083) );
  XOR2_X1 U12185 ( .A(n12243), .B(n12244), .Z(n12242) );
  XOR2_X1 U12186 ( .A(n12245), .B(n12246), .Z(n12087) );
  XOR2_X1 U12187 ( .A(n12247), .B(n12248), .Z(n12246) );
  XOR2_X1 U12188 ( .A(n12249), .B(n12250), .Z(n12091) );
  XOR2_X1 U12189 ( .A(n12251), .B(n12252), .Z(n12250) );
  XOR2_X1 U12190 ( .A(n12253), .B(n12254), .Z(n12095) );
  XOR2_X1 U12191 ( .A(n12255), .B(n12256), .Z(n12254) );
  XOR2_X1 U12192 ( .A(n12257), .B(n12258), .Z(n12099) );
  XOR2_X1 U12193 ( .A(n12259), .B(n12260), .Z(n12258) );
  XOR2_X1 U12194 ( .A(n12261), .B(n12262), .Z(n12103) );
  XOR2_X1 U12195 ( .A(n12263), .B(n12264), .Z(n12262) );
  XOR2_X1 U12196 ( .A(n12265), .B(n12266), .Z(n12107) );
  XOR2_X1 U12197 ( .A(n12267), .B(n12268), .Z(n12266) );
  XOR2_X1 U12198 ( .A(n12269), .B(n12270), .Z(n12111) );
  XOR2_X1 U12199 ( .A(n12271), .B(n12272), .Z(n12270) );
  XOR2_X1 U12200 ( .A(n12273), .B(n12274), .Z(n12115) );
  XOR2_X1 U12201 ( .A(n12275), .B(n12276), .Z(n12274) );
  XOR2_X1 U12202 ( .A(n12277), .B(n12278), .Z(n12119) );
  XOR2_X1 U12203 ( .A(n12279), .B(n12280), .Z(n12278) );
  XOR2_X1 U12204 ( .A(n12281), .B(n12282), .Z(n12123) );
  XOR2_X1 U12205 ( .A(n12283), .B(n12284), .Z(n12282) );
  XOR2_X1 U12206 ( .A(n12285), .B(n12286), .Z(n12127) );
  XOR2_X1 U12207 ( .A(n12287), .B(n12288), .Z(n12286) );
  XOR2_X1 U12208 ( .A(n12289), .B(n12290), .Z(n12131) );
  XOR2_X1 U12209 ( .A(n12291), .B(n12292), .Z(n12290) );
  XOR2_X1 U12210 ( .A(n12293), .B(n12294), .Z(n12134) );
  XOR2_X1 U12211 ( .A(n12295), .B(n12296), .Z(n12294) );
  XNOR2_X1 U12212 ( .A(n12297), .B(n12298), .ZN(n12138) );
  XNOR2_X1 U12213 ( .A(n8000), .B(n12299), .ZN(n12297) );
  XOR2_X1 U12214 ( .A(n12300), .B(n12301), .Z(n12142) );
  XOR2_X1 U12215 ( .A(n12302), .B(n12303), .Z(n12301) );
  XOR2_X1 U12216 ( .A(n12304), .B(n12305), .Z(n12146) );
  XOR2_X1 U12217 ( .A(n12306), .B(n12307), .Z(n12305) );
  XOR2_X1 U12218 ( .A(n12308), .B(n12309), .Z(n12150) );
  XOR2_X1 U12219 ( .A(n12310), .B(n12311), .Z(n12309) );
  XOR2_X1 U12220 ( .A(n12312), .B(n12313), .Z(n12154) );
  XOR2_X1 U12221 ( .A(n12314), .B(n12315), .Z(n12313) );
  XOR2_X1 U12222 ( .A(n12316), .B(n12317), .Z(n12158) );
  XOR2_X1 U12223 ( .A(n12318), .B(n12319), .Z(n12317) );
  XOR2_X1 U12224 ( .A(n12320), .B(n12321), .Z(n10851) );
  XOR2_X1 U12225 ( .A(n12322), .B(n12323), .Z(n12321) );
  XNOR2_X1 U12226 ( .A(n8176), .B(n8527), .ZN(n8164) );
  OR2_X1 U12227 ( .A1(n12324), .A2(n12325), .ZN(n8527) );
  AND2_X1 U12228 ( .A1(n8546), .A2(n8545), .ZN(n12325) );
  AND2_X1 U12229 ( .A1(n8543), .A2(n12326), .ZN(n12324) );
  OR2_X1 U12230 ( .A1(n8545), .A2(n8546), .ZN(n12326) );
  OR2_X1 U12231 ( .A1(n7950), .A2(n7999), .ZN(n8546) );
  OR2_X1 U12232 ( .A1(n12327), .A2(n12328), .ZN(n8545) );
  AND2_X1 U12233 ( .A1(n8570), .A2(n8569), .ZN(n12328) );
  AND2_X1 U12234 ( .A1(n8567), .A2(n12329), .ZN(n12327) );
  OR2_X1 U12235 ( .A1(n8569), .A2(n8570), .ZN(n12329) );
  OR2_X1 U12236 ( .A1(n7953), .A2(n7999), .ZN(n8570) );
  OR2_X1 U12237 ( .A1(n12330), .A2(n12331), .ZN(n8569) );
  AND2_X1 U12238 ( .A1(n8601), .A2(n8600), .ZN(n12331) );
  AND2_X1 U12239 ( .A1(n8598), .A2(n12332), .ZN(n12330) );
  OR2_X1 U12240 ( .A1(n8600), .A2(n8601), .ZN(n12332) );
  OR2_X1 U12241 ( .A1(n7956), .A2(n7999), .ZN(n8601) );
  OR2_X1 U12242 ( .A1(n12333), .A2(n12334), .ZN(n8600) );
  AND2_X1 U12243 ( .A1(n8639), .A2(n8638), .ZN(n12334) );
  AND2_X1 U12244 ( .A1(n8636), .A2(n12335), .ZN(n12333) );
  OR2_X1 U12245 ( .A1(n8638), .A2(n8639), .ZN(n12335) );
  OR2_X1 U12246 ( .A1(n7960), .A2(n7999), .ZN(n8639) );
  OR2_X1 U12247 ( .A1(n12336), .A2(n12337), .ZN(n8638) );
  AND2_X1 U12248 ( .A1(n8684), .A2(n8683), .ZN(n12337) );
  AND2_X1 U12249 ( .A1(n8681), .A2(n12338), .ZN(n12336) );
  OR2_X1 U12250 ( .A1(n8683), .A2(n8684), .ZN(n12338) );
  OR2_X1 U12251 ( .A1(n7963), .A2(n7999), .ZN(n8684) );
  OR2_X1 U12252 ( .A1(n12339), .A2(n12340), .ZN(n8683) );
  AND2_X1 U12253 ( .A1(n8736), .A2(n8735), .ZN(n12340) );
  AND2_X1 U12254 ( .A1(n8733), .A2(n12341), .ZN(n12339) );
  OR2_X1 U12255 ( .A1(n8735), .A2(n8736), .ZN(n12341) );
  OR2_X1 U12256 ( .A1(n7967), .A2(n7999), .ZN(n8736) );
  OR2_X1 U12257 ( .A1(n12342), .A2(n12343), .ZN(n8735) );
  AND2_X1 U12258 ( .A1(n10803), .A2(n10802), .ZN(n12343) );
  AND2_X1 U12259 ( .A1(n10800), .A2(n12344), .ZN(n12342) );
  OR2_X1 U12260 ( .A1(n10802), .A2(n10803), .ZN(n12344) );
  OR2_X1 U12261 ( .A1(n7970), .A2(n7999), .ZN(n10803) );
  OR2_X1 U12262 ( .A1(n12345), .A2(n12346), .ZN(n10802) );
  AND2_X1 U12263 ( .A1(n10856), .A2(n10855), .ZN(n12346) );
  AND2_X1 U12264 ( .A1(n10853), .A2(n12347), .ZN(n12345) );
  OR2_X1 U12265 ( .A1(n10855), .A2(n10856), .ZN(n12347) );
  OR2_X1 U12266 ( .A1(n7974), .A2(n7999), .ZN(n10856) );
  OR2_X1 U12267 ( .A1(n12348), .A2(n12349), .ZN(n10855) );
  AND2_X1 U12268 ( .A1(n12323), .A2(n12322), .ZN(n12349) );
  AND2_X1 U12269 ( .A1(n12320), .A2(n12350), .ZN(n12348) );
  OR2_X1 U12270 ( .A1(n12322), .A2(n12323), .ZN(n12350) );
  OR2_X1 U12271 ( .A1(n7977), .A2(n7999), .ZN(n12323) );
  OR2_X1 U12272 ( .A1(n12351), .A2(n12352), .ZN(n12322) );
  AND2_X1 U12273 ( .A1(n12319), .A2(n12318), .ZN(n12352) );
  AND2_X1 U12274 ( .A1(n12316), .A2(n12353), .ZN(n12351) );
  OR2_X1 U12275 ( .A1(n12318), .A2(n12319), .ZN(n12353) );
  OR2_X1 U12276 ( .A1(n7981), .A2(n7999), .ZN(n12319) );
  OR2_X1 U12277 ( .A1(n12354), .A2(n12355), .ZN(n12318) );
  AND2_X1 U12278 ( .A1(n12315), .A2(n12314), .ZN(n12355) );
  AND2_X1 U12279 ( .A1(n12312), .A2(n12356), .ZN(n12354) );
  OR2_X1 U12280 ( .A1(n12314), .A2(n12315), .ZN(n12356) );
  OR2_X1 U12281 ( .A1(n7984), .A2(n7999), .ZN(n12315) );
  OR2_X1 U12282 ( .A1(n12357), .A2(n12358), .ZN(n12314) );
  AND2_X1 U12283 ( .A1(n12311), .A2(n12310), .ZN(n12358) );
  AND2_X1 U12284 ( .A1(n12308), .A2(n12359), .ZN(n12357) );
  OR2_X1 U12285 ( .A1(n12310), .A2(n12311), .ZN(n12359) );
  OR2_X1 U12286 ( .A1(n7988), .A2(n7999), .ZN(n12311) );
  OR2_X1 U12287 ( .A1(n12360), .A2(n12361), .ZN(n12310) );
  AND2_X1 U12288 ( .A1(n12307), .A2(n12306), .ZN(n12361) );
  AND2_X1 U12289 ( .A1(n12304), .A2(n12362), .ZN(n12360) );
  OR2_X1 U12290 ( .A1(n12306), .A2(n12307), .ZN(n12362) );
  OR2_X1 U12291 ( .A1(n7991), .A2(n7999), .ZN(n12307) );
  OR2_X1 U12292 ( .A1(n12363), .A2(n12364), .ZN(n12306) );
  AND2_X1 U12293 ( .A1(n12303), .A2(n12302), .ZN(n12364) );
  AND2_X1 U12294 ( .A1(n12300), .A2(n12365), .ZN(n12363) );
  OR2_X1 U12295 ( .A1(n12302), .A2(n12303), .ZN(n12365) );
  OR2_X1 U12296 ( .A1(n7995), .A2(n7999), .ZN(n12303) );
  OR2_X1 U12297 ( .A1(n12366), .A2(n12367), .ZN(n12302) );
  AND2_X1 U12298 ( .A1(n12299), .A2(n8000), .ZN(n12367) );
  AND2_X1 U12299 ( .A1(n12298), .A2(n12368), .ZN(n12366) );
  OR2_X1 U12300 ( .A1(n8000), .A2(n12299), .ZN(n12368) );
  OR2_X1 U12301 ( .A1(n12369), .A2(n12370), .ZN(n12299) );
  AND2_X1 U12302 ( .A1(n12296), .A2(n12295), .ZN(n12370) );
  AND2_X1 U12303 ( .A1(n12293), .A2(n12371), .ZN(n12369) );
  OR2_X1 U12304 ( .A1(n12295), .A2(n12296), .ZN(n12371) );
  OR2_X1 U12305 ( .A1(n8002), .A2(n7999), .ZN(n12296) );
  OR2_X1 U12306 ( .A1(n12372), .A2(n12373), .ZN(n12295) );
  AND2_X1 U12307 ( .A1(n12292), .A2(n12291), .ZN(n12373) );
  AND2_X1 U12308 ( .A1(n12289), .A2(n12374), .ZN(n12372) );
  OR2_X1 U12309 ( .A1(n12291), .A2(n12292), .ZN(n12374) );
  OR2_X1 U12310 ( .A1(n8005), .A2(n7999), .ZN(n12292) );
  OR2_X1 U12311 ( .A1(n12375), .A2(n12376), .ZN(n12291) );
  AND2_X1 U12312 ( .A1(n12288), .A2(n12287), .ZN(n12376) );
  AND2_X1 U12313 ( .A1(n12285), .A2(n12377), .ZN(n12375) );
  OR2_X1 U12314 ( .A1(n12287), .A2(n12288), .ZN(n12377) );
  OR2_X1 U12315 ( .A1(n8009), .A2(n7999), .ZN(n12288) );
  OR2_X1 U12316 ( .A1(n12378), .A2(n12379), .ZN(n12287) );
  AND2_X1 U12317 ( .A1(n12284), .A2(n12283), .ZN(n12379) );
  AND2_X1 U12318 ( .A1(n12281), .A2(n12380), .ZN(n12378) );
  OR2_X1 U12319 ( .A1(n12283), .A2(n12284), .ZN(n12380) );
  OR2_X1 U12320 ( .A1(n8012), .A2(n7999), .ZN(n12284) );
  OR2_X1 U12321 ( .A1(n12381), .A2(n12382), .ZN(n12283) );
  AND2_X1 U12322 ( .A1(n12280), .A2(n12279), .ZN(n12382) );
  AND2_X1 U12323 ( .A1(n12277), .A2(n12383), .ZN(n12381) );
  OR2_X1 U12324 ( .A1(n12279), .A2(n12280), .ZN(n12383) );
  OR2_X1 U12325 ( .A1(n8016), .A2(n7999), .ZN(n12280) );
  OR2_X1 U12326 ( .A1(n12384), .A2(n12385), .ZN(n12279) );
  AND2_X1 U12327 ( .A1(n12276), .A2(n12275), .ZN(n12385) );
  AND2_X1 U12328 ( .A1(n12273), .A2(n12386), .ZN(n12384) );
  OR2_X1 U12329 ( .A1(n12275), .A2(n12276), .ZN(n12386) );
  OR2_X1 U12330 ( .A1(n8019), .A2(n7999), .ZN(n12276) );
  OR2_X1 U12331 ( .A1(n12387), .A2(n12388), .ZN(n12275) );
  AND2_X1 U12332 ( .A1(n12272), .A2(n12271), .ZN(n12388) );
  AND2_X1 U12333 ( .A1(n12269), .A2(n12389), .ZN(n12387) );
  OR2_X1 U12334 ( .A1(n12271), .A2(n12272), .ZN(n12389) );
  OR2_X1 U12335 ( .A1(n8023), .A2(n7999), .ZN(n12272) );
  OR2_X1 U12336 ( .A1(n12390), .A2(n12391), .ZN(n12271) );
  AND2_X1 U12337 ( .A1(n12268), .A2(n12267), .ZN(n12391) );
  AND2_X1 U12338 ( .A1(n12265), .A2(n12392), .ZN(n12390) );
  OR2_X1 U12339 ( .A1(n12267), .A2(n12268), .ZN(n12392) );
  OR2_X1 U12340 ( .A1(n8026), .A2(n7999), .ZN(n12268) );
  OR2_X1 U12341 ( .A1(n12393), .A2(n12394), .ZN(n12267) );
  AND2_X1 U12342 ( .A1(n12264), .A2(n12263), .ZN(n12394) );
  AND2_X1 U12343 ( .A1(n12261), .A2(n12395), .ZN(n12393) );
  OR2_X1 U12344 ( .A1(n12263), .A2(n12264), .ZN(n12395) );
  OR2_X1 U12345 ( .A1(n8030), .A2(n7999), .ZN(n12264) );
  OR2_X1 U12346 ( .A1(n12396), .A2(n12397), .ZN(n12263) );
  AND2_X1 U12347 ( .A1(n12260), .A2(n12259), .ZN(n12397) );
  AND2_X1 U12348 ( .A1(n12257), .A2(n12398), .ZN(n12396) );
  OR2_X1 U12349 ( .A1(n12259), .A2(n12260), .ZN(n12398) );
  OR2_X1 U12350 ( .A1(n8034), .A2(n7999), .ZN(n12260) );
  OR2_X1 U12351 ( .A1(n12399), .A2(n12400), .ZN(n12259) );
  AND2_X1 U12352 ( .A1(n12256), .A2(n12255), .ZN(n12400) );
  AND2_X1 U12353 ( .A1(n12253), .A2(n12401), .ZN(n12399) );
  OR2_X1 U12354 ( .A1(n12255), .A2(n12256), .ZN(n12401) );
  OR2_X1 U12355 ( .A1(n8037), .A2(n7999), .ZN(n12256) );
  OR2_X1 U12356 ( .A1(n12402), .A2(n12403), .ZN(n12255) );
  AND2_X1 U12357 ( .A1(n12252), .A2(n12251), .ZN(n12403) );
  AND2_X1 U12358 ( .A1(n12249), .A2(n12404), .ZN(n12402) );
  OR2_X1 U12359 ( .A1(n12251), .A2(n12252), .ZN(n12404) );
  OR2_X1 U12360 ( .A1(n8041), .A2(n7999), .ZN(n12252) );
  OR2_X1 U12361 ( .A1(n12405), .A2(n12406), .ZN(n12251) );
  AND2_X1 U12362 ( .A1(n12248), .A2(n12247), .ZN(n12406) );
  AND2_X1 U12363 ( .A1(n12245), .A2(n12407), .ZN(n12405) );
  OR2_X1 U12364 ( .A1(n12247), .A2(n12248), .ZN(n12407) );
  OR2_X1 U12365 ( .A1(n8044), .A2(n7999), .ZN(n12248) );
  OR2_X1 U12366 ( .A1(n12408), .A2(n12409), .ZN(n12247) );
  AND2_X1 U12367 ( .A1(n12244), .A2(n12243), .ZN(n12409) );
  AND2_X1 U12368 ( .A1(n12241), .A2(n12410), .ZN(n12408) );
  OR2_X1 U12369 ( .A1(n12243), .A2(n12244), .ZN(n12410) );
  OR2_X1 U12370 ( .A1(n8048), .A2(n7999), .ZN(n12244) );
  OR2_X1 U12371 ( .A1(n12411), .A2(n12412), .ZN(n12243) );
  AND2_X1 U12372 ( .A1(n12237), .A2(n12413), .ZN(n12412) );
  AND2_X1 U12373 ( .A1(n12414), .A2(n12415), .ZN(n12411) );
  OR2_X1 U12374 ( .A1(n12413), .A2(n12237), .ZN(n12415) );
  OR2_X1 U12375 ( .A1(n8051), .A2(n7999), .ZN(n12237) );
  INV_X1 U12376 ( .A(b_14_), .ZN(n7999) );
  INV_X1 U12377 ( .A(n12240), .ZN(n12413) );
  AND3_X1 U12378 ( .A1(n8904), .A2(b_13_), .A3(b_14_), .ZN(n12240) );
  INV_X1 U12379 ( .A(n12239), .ZN(n12414) );
  OR2_X1 U12380 ( .A1(n12416), .A2(n12417), .ZN(n12239) );
  AND2_X1 U12381 ( .A1(b_13_), .A2(n12418), .ZN(n12417) );
  OR2_X1 U12382 ( .A1(n12419), .A2(n7490), .ZN(n12418) );
  AND2_X1 U12383 ( .A1(a_30_), .A2(n7992), .ZN(n12419) );
  AND2_X1 U12384 ( .A1(b_12_), .A2(n12420), .ZN(n12416) );
  OR2_X1 U12385 ( .A1(n12421), .A2(n7493), .ZN(n12420) );
  AND2_X1 U12386 ( .A1(a_31_), .A2(n7746), .ZN(n12421) );
  XNOR2_X1 U12387 ( .A(n12422), .B(n12423), .ZN(n12241) );
  XNOR2_X1 U12388 ( .A(n12424), .B(n12425), .ZN(n12423) );
  XOR2_X1 U12389 ( .A(n12426), .B(n12427), .Z(n12245) );
  XOR2_X1 U12390 ( .A(n12428), .B(n12429), .Z(n12427) );
  XOR2_X1 U12391 ( .A(n12430), .B(n12431), .Z(n12249) );
  XOR2_X1 U12392 ( .A(n12432), .B(n12433), .Z(n12431) );
  XOR2_X1 U12393 ( .A(n12434), .B(n12435), .Z(n12253) );
  XOR2_X1 U12394 ( .A(n12436), .B(n12437), .Z(n12435) );
  XOR2_X1 U12395 ( .A(n12438), .B(n12439), .Z(n12257) );
  XOR2_X1 U12396 ( .A(n12440), .B(n12441), .Z(n12439) );
  XOR2_X1 U12397 ( .A(n12442), .B(n12443), .Z(n12261) );
  XOR2_X1 U12398 ( .A(n12444), .B(n12445), .Z(n12443) );
  XOR2_X1 U12399 ( .A(n12446), .B(n12447), .Z(n12265) );
  XOR2_X1 U12400 ( .A(n12448), .B(n12449), .Z(n12447) );
  XOR2_X1 U12401 ( .A(n12450), .B(n12451), .Z(n12269) );
  XOR2_X1 U12402 ( .A(n12452), .B(n12453), .Z(n12451) );
  XOR2_X1 U12403 ( .A(n12454), .B(n12455), .Z(n12273) );
  XOR2_X1 U12404 ( .A(n12456), .B(n12457), .Z(n12455) );
  XOR2_X1 U12405 ( .A(n12458), .B(n12459), .Z(n12277) );
  XOR2_X1 U12406 ( .A(n12460), .B(n12461), .Z(n12459) );
  XOR2_X1 U12407 ( .A(n12462), .B(n12463), .Z(n12281) );
  XOR2_X1 U12408 ( .A(n12464), .B(n12465), .Z(n12463) );
  XOR2_X1 U12409 ( .A(n12466), .B(n12467), .Z(n12285) );
  XOR2_X1 U12410 ( .A(n12468), .B(n12469), .Z(n12467) );
  XOR2_X1 U12411 ( .A(n12470), .B(n12471), .Z(n12289) );
  XOR2_X1 U12412 ( .A(n12472), .B(n12473), .Z(n12471) );
  XOR2_X1 U12413 ( .A(n12474), .B(n12475), .Z(n12293) );
  XOR2_X1 U12414 ( .A(n12476), .B(n12477), .Z(n12475) );
  INV_X1 U12415 ( .A(n7738), .ZN(n8000) );
  AND2_X1 U12416 ( .A1(a_14_), .A2(b_14_), .ZN(n7738) );
  XOR2_X1 U12417 ( .A(n12478), .B(n12479), .Z(n12298) );
  XOR2_X1 U12418 ( .A(n12480), .B(n12481), .Z(n12479) );
  XOR2_X1 U12419 ( .A(n12482), .B(n12483), .Z(n12300) );
  XOR2_X1 U12420 ( .A(n12484), .B(n12485), .Z(n12483) );
  XOR2_X1 U12421 ( .A(n12486), .B(n12487), .Z(n12304) );
  XNOR2_X1 U12422 ( .A(n12488), .B(n7750), .ZN(n12487) );
  XOR2_X1 U12423 ( .A(n12489), .B(n12490), .Z(n12308) );
  XOR2_X1 U12424 ( .A(n12491), .B(n12492), .Z(n12490) );
  XOR2_X1 U12425 ( .A(n12493), .B(n12494), .Z(n12312) );
  XOR2_X1 U12426 ( .A(n12495), .B(n12496), .Z(n12494) );
  XOR2_X1 U12427 ( .A(n12497), .B(n12498), .Z(n12316) );
  XOR2_X1 U12428 ( .A(n12499), .B(n12500), .Z(n12498) );
  XOR2_X1 U12429 ( .A(n12501), .B(n12502), .Z(n12320) );
  XOR2_X1 U12430 ( .A(n12503), .B(n12504), .Z(n12502) );
  XOR2_X1 U12431 ( .A(n12505), .B(n12506), .Z(n10853) );
  XOR2_X1 U12432 ( .A(n12507), .B(n12508), .Z(n12506) );
  XOR2_X1 U12433 ( .A(n12509), .B(n12510), .Z(n10800) );
  XOR2_X1 U12434 ( .A(n12511), .B(n12512), .Z(n12510) );
  XOR2_X1 U12435 ( .A(n12513), .B(n12514), .Z(n8733) );
  XOR2_X1 U12436 ( .A(n12515), .B(n12516), .Z(n12514) );
  XOR2_X1 U12437 ( .A(n12517), .B(n12518), .Z(n8681) );
  XOR2_X1 U12438 ( .A(n12519), .B(n12520), .Z(n12518) );
  XOR2_X1 U12439 ( .A(n12521), .B(n12522), .Z(n8636) );
  XOR2_X1 U12440 ( .A(n12523), .B(n12524), .Z(n12522) );
  XOR2_X1 U12441 ( .A(n12525), .B(n12526), .Z(n8598) );
  XOR2_X1 U12442 ( .A(n12527), .B(n12528), .Z(n12526) );
  XOR2_X1 U12443 ( .A(n12529), .B(n12530), .Z(n8567) );
  XOR2_X1 U12444 ( .A(n12531), .B(n12532), .Z(n12530) );
  XOR2_X1 U12445 ( .A(n12533), .B(n12534), .Z(n8543) );
  XOR2_X1 U12446 ( .A(n12535), .B(n12536), .Z(n12534) );
  XNOR2_X1 U12447 ( .A(n12537), .B(n12538), .ZN(n8176) );
  XOR2_X1 U12448 ( .A(n12539), .B(n12540), .Z(n12538) );
  INV_X1 U12449 ( .A(n12541), .ZN(n8174) );
  OR2_X1 U12450 ( .A1(n12542), .A2(n8524), .ZN(n12541) );
  AND2_X1 U12451 ( .A1(n12543), .A2(n12544), .ZN(n12542) );
  INV_X1 U12452 ( .A(n12545), .ZN(n8524) );
  OR2_X1 U12453 ( .A1(n12543), .A2(n12544), .ZN(n12545) );
  OR2_X1 U12454 ( .A1(n12546), .A2(n12547), .ZN(n12544) );
  AND2_X1 U12455 ( .A1(n12540), .A2(n12539), .ZN(n12547) );
  AND2_X1 U12456 ( .A1(n12537), .A2(n12548), .ZN(n12546) );
  OR2_X1 U12457 ( .A1(n12540), .A2(n12539), .ZN(n12548) );
  OR2_X1 U12458 ( .A1(n12549), .A2(n12550), .ZN(n12539) );
  AND2_X1 U12459 ( .A1(n12536), .A2(n12535), .ZN(n12550) );
  AND2_X1 U12460 ( .A1(n12533), .A2(n12551), .ZN(n12549) );
  OR2_X1 U12461 ( .A1(n12536), .A2(n12535), .ZN(n12551) );
  OR2_X1 U12462 ( .A1(n12552), .A2(n12553), .ZN(n12535) );
  AND2_X1 U12463 ( .A1(n12532), .A2(n12531), .ZN(n12553) );
  AND2_X1 U12464 ( .A1(n12529), .A2(n12554), .ZN(n12552) );
  OR2_X1 U12465 ( .A1(n12532), .A2(n12531), .ZN(n12554) );
  OR2_X1 U12466 ( .A1(n12555), .A2(n12556), .ZN(n12531) );
  AND2_X1 U12467 ( .A1(n12528), .A2(n12527), .ZN(n12556) );
  AND2_X1 U12468 ( .A1(n12525), .A2(n12557), .ZN(n12555) );
  OR2_X1 U12469 ( .A1(n12528), .A2(n12527), .ZN(n12557) );
  OR2_X1 U12470 ( .A1(n12558), .A2(n12559), .ZN(n12527) );
  AND2_X1 U12471 ( .A1(n12524), .A2(n12523), .ZN(n12559) );
  AND2_X1 U12472 ( .A1(n12521), .A2(n12560), .ZN(n12558) );
  OR2_X1 U12473 ( .A1(n12524), .A2(n12523), .ZN(n12560) );
  OR2_X1 U12474 ( .A1(n12561), .A2(n12562), .ZN(n12523) );
  AND2_X1 U12475 ( .A1(n12520), .A2(n12519), .ZN(n12562) );
  AND2_X1 U12476 ( .A1(n12517), .A2(n12563), .ZN(n12561) );
  OR2_X1 U12477 ( .A1(n12520), .A2(n12519), .ZN(n12563) );
  OR2_X1 U12478 ( .A1(n12564), .A2(n12565), .ZN(n12519) );
  AND2_X1 U12479 ( .A1(n12516), .A2(n12515), .ZN(n12565) );
  AND2_X1 U12480 ( .A1(n12513), .A2(n12566), .ZN(n12564) );
  OR2_X1 U12481 ( .A1(n12516), .A2(n12515), .ZN(n12566) );
  OR2_X1 U12482 ( .A1(n12567), .A2(n12568), .ZN(n12515) );
  AND2_X1 U12483 ( .A1(n12512), .A2(n12511), .ZN(n12568) );
  AND2_X1 U12484 ( .A1(n12509), .A2(n12569), .ZN(n12567) );
  OR2_X1 U12485 ( .A1(n12512), .A2(n12511), .ZN(n12569) );
  OR2_X1 U12486 ( .A1(n12570), .A2(n12571), .ZN(n12511) );
  AND2_X1 U12487 ( .A1(n12508), .A2(n12507), .ZN(n12571) );
  AND2_X1 U12488 ( .A1(n12505), .A2(n12572), .ZN(n12570) );
  OR2_X1 U12489 ( .A1(n12508), .A2(n12507), .ZN(n12572) );
  OR2_X1 U12490 ( .A1(n12573), .A2(n12574), .ZN(n12507) );
  AND2_X1 U12491 ( .A1(n12504), .A2(n12503), .ZN(n12574) );
  AND2_X1 U12492 ( .A1(n12501), .A2(n12575), .ZN(n12573) );
  OR2_X1 U12493 ( .A1(n12504), .A2(n12503), .ZN(n12575) );
  OR2_X1 U12494 ( .A1(n12576), .A2(n12577), .ZN(n12503) );
  AND2_X1 U12495 ( .A1(n12500), .A2(n12499), .ZN(n12577) );
  AND2_X1 U12496 ( .A1(n12497), .A2(n12578), .ZN(n12576) );
  OR2_X1 U12497 ( .A1(n12500), .A2(n12499), .ZN(n12578) );
  OR2_X1 U12498 ( .A1(n12579), .A2(n12580), .ZN(n12499) );
  AND2_X1 U12499 ( .A1(n12496), .A2(n12495), .ZN(n12580) );
  AND2_X1 U12500 ( .A1(n12493), .A2(n12581), .ZN(n12579) );
  OR2_X1 U12501 ( .A1(n12496), .A2(n12495), .ZN(n12581) );
  OR2_X1 U12502 ( .A1(n12582), .A2(n12583), .ZN(n12495) );
  AND2_X1 U12503 ( .A1(n12492), .A2(n12491), .ZN(n12583) );
  AND2_X1 U12504 ( .A1(n12489), .A2(n12584), .ZN(n12582) );
  OR2_X1 U12505 ( .A1(n12492), .A2(n12491), .ZN(n12584) );
  OR2_X1 U12506 ( .A1(n12585), .A2(n12586), .ZN(n12491) );
  AND2_X1 U12507 ( .A1(n7996), .A2(n12488), .ZN(n12586) );
  AND2_X1 U12508 ( .A1(n12486), .A2(n12587), .ZN(n12585) );
  OR2_X1 U12509 ( .A1(n7996), .A2(n12488), .ZN(n12587) );
  OR2_X1 U12510 ( .A1(n12588), .A2(n12589), .ZN(n12488) );
  AND2_X1 U12511 ( .A1(n12485), .A2(n12484), .ZN(n12589) );
  AND2_X1 U12512 ( .A1(n12482), .A2(n12590), .ZN(n12588) );
  OR2_X1 U12513 ( .A1(n12485), .A2(n12484), .ZN(n12590) );
  OR2_X1 U12514 ( .A1(n12591), .A2(n12592), .ZN(n12484) );
  AND2_X1 U12515 ( .A1(n12481), .A2(n12480), .ZN(n12592) );
  AND2_X1 U12516 ( .A1(n12478), .A2(n12593), .ZN(n12591) );
  OR2_X1 U12517 ( .A1(n12481), .A2(n12480), .ZN(n12593) );
  OR2_X1 U12518 ( .A1(n12594), .A2(n12595), .ZN(n12480) );
  AND2_X1 U12519 ( .A1(n12477), .A2(n12476), .ZN(n12595) );
  AND2_X1 U12520 ( .A1(n12474), .A2(n12596), .ZN(n12594) );
  OR2_X1 U12521 ( .A1(n12477), .A2(n12476), .ZN(n12596) );
  OR2_X1 U12522 ( .A1(n12597), .A2(n12598), .ZN(n12476) );
  AND2_X1 U12523 ( .A1(n12473), .A2(n12472), .ZN(n12598) );
  AND2_X1 U12524 ( .A1(n12470), .A2(n12599), .ZN(n12597) );
  OR2_X1 U12525 ( .A1(n12473), .A2(n12472), .ZN(n12599) );
  OR2_X1 U12526 ( .A1(n12600), .A2(n12601), .ZN(n12472) );
  AND2_X1 U12527 ( .A1(n12469), .A2(n12468), .ZN(n12601) );
  AND2_X1 U12528 ( .A1(n12466), .A2(n12602), .ZN(n12600) );
  OR2_X1 U12529 ( .A1(n12469), .A2(n12468), .ZN(n12602) );
  OR2_X1 U12530 ( .A1(n12603), .A2(n12604), .ZN(n12468) );
  AND2_X1 U12531 ( .A1(n12465), .A2(n12464), .ZN(n12604) );
  AND2_X1 U12532 ( .A1(n12462), .A2(n12605), .ZN(n12603) );
  OR2_X1 U12533 ( .A1(n12465), .A2(n12464), .ZN(n12605) );
  OR2_X1 U12534 ( .A1(n12606), .A2(n12607), .ZN(n12464) );
  AND2_X1 U12535 ( .A1(n12461), .A2(n12460), .ZN(n12607) );
  AND2_X1 U12536 ( .A1(n12458), .A2(n12608), .ZN(n12606) );
  OR2_X1 U12537 ( .A1(n12461), .A2(n12460), .ZN(n12608) );
  OR2_X1 U12538 ( .A1(n12609), .A2(n12610), .ZN(n12460) );
  AND2_X1 U12539 ( .A1(n12457), .A2(n12456), .ZN(n12610) );
  AND2_X1 U12540 ( .A1(n12454), .A2(n12611), .ZN(n12609) );
  OR2_X1 U12541 ( .A1(n12457), .A2(n12456), .ZN(n12611) );
  OR2_X1 U12542 ( .A1(n12612), .A2(n12613), .ZN(n12456) );
  AND2_X1 U12543 ( .A1(n12453), .A2(n12452), .ZN(n12613) );
  AND2_X1 U12544 ( .A1(n12450), .A2(n12614), .ZN(n12612) );
  OR2_X1 U12545 ( .A1(n12453), .A2(n12452), .ZN(n12614) );
  OR2_X1 U12546 ( .A1(n12615), .A2(n12616), .ZN(n12452) );
  AND2_X1 U12547 ( .A1(n12449), .A2(n12448), .ZN(n12616) );
  AND2_X1 U12548 ( .A1(n12446), .A2(n12617), .ZN(n12615) );
  OR2_X1 U12549 ( .A1(n12449), .A2(n12448), .ZN(n12617) );
  OR2_X1 U12550 ( .A1(n12618), .A2(n12619), .ZN(n12448) );
  AND2_X1 U12551 ( .A1(n12445), .A2(n12444), .ZN(n12619) );
  AND2_X1 U12552 ( .A1(n12442), .A2(n12620), .ZN(n12618) );
  OR2_X1 U12553 ( .A1(n12445), .A2(n12444), .ZN(n12620) );
  OR2_X1 U12554 ( .A1(n12621), .A2(n12622), .ZN(n12444) );
  AND2_X1 U12555 ( .A1(n12441), .A2(n12440), .ZN(n12622) );
  AND2_X1 U12556 ( .A1(n12438), .A2(n12623), .ZN(n12621) );
  OR2_X1 U12557 ( .A1(n12441), .A2(n12440), .ZN(n12623) );
  OR2_X1 U12558 ( .A1(n12624), .A2(n12625), .ZN(n12440) );
  AND2_X1 U12559 ( .A1(n12437), .A2(n12436), .ZN(n12625) );
  AND2_X1 U12560 ( .A1(n12434), .A2(n12626), .ZN(n12624) );
  OR2_X1 U12561 ( .A1(n12437), .A2(n12436), .ZN(n12626) );
  OR2_X1 U12562 ( .A1(n12627), .A2(n12628), .ZN(n12436) );
  AND2_X1 U12563 ( .A1(n12433), .A2(n12432), .ZN(n12628) );
  AND2_X1 U12564 ( .A1(n12430), .A2(n12629), .ZN(n12627) );
  OR2_X1 U12565 ( .A1(n12433), .A2(n12432), .ZN(n12629) );
  OR2_X1 U12566 ( .A1(n12630), .A2(n12631), .ZN(n12432) );
  AND2_X1 U12567 ( .A1(n12429), .A2(n12428), .ZN(n12631) );
  AND2_X1 U12568 ( .A1(n12426), .A2(n12632), .ZN(n12630) );
  OR2_X1 U12569 ( .A1(n12429), .A2(n12428), .ZN(n12632) );
  OR2_X1 U12570 ( .A1(n12633), .A2(n12634), .ZN(n12428) );
  AND2_X1 U12571 ( .A1(n12422), .A2(n12635), .ZN(n12634) );
  AND2_X1 U12572 ( .A1(n12636), .A2(n12637), .ZN(n12633) );
  OR2_X1 U12573 ( .A1(n12422), .A2(n12635), .ZN(n12637) );
  INV_X1 U12574 ( .A(n12425), .ZN(n12635) );
  AND3_X1 U12575 ( .A1(n8904), .A2(b_12_), .A3(b_13_), .ZN(n12425) );
  OR2_X1 U12576 ( .A1(n8051), .A2(n7746), .ZN(n12422) );
  INV_X1 U12577 ( .A(n12424), .ZN(n12636) );
  OR2_X1 U12578 ( .A1(n12638), .A2(n12639), .ZN(n12424) );
  AND2_X1 U12579 ( .A1(b_12_), .A2(n12640), .ZN(n12639) );
  OR2_X1 U12580 ( .A1(n12641), .A2(n7490), .ZN(n12640) );
  AND2_X1 U12581 ( .A1(a_30_), .A2(n7775), .ZN(n12641) );
  AND2_X1 U12582 ( .A1(b_11_), .A2(n12642), .ZN(n12638) );
  OR2_X1 U12583 ( .A1(n12643), .A2(n7493), .ZN(n12642) );
  AND2_X1 U12584 ( .A1(a_31_), .A2(n7992), .ZN(n12643) );
  OR2_X1 U12585 ( .A1(n8048), .A2(n7746), .ZN(n12429) );
  XNOR2_X1 U12586 ( .A(n12644), .B(n12645), .ZN(n12426) );
  XNOR2_X1 U12587 ( .A(n12646), .B(n12647), .ZN(n12645) );
  OR2_X1 U12588 ( .A1(n8044), .A2(n7746), .ZN(n12433) );
  XOR2_X1 U12589 ( .A(n12648), .B(n12649), .Z(n12430) );
  XOR2_X1 U12590 ( .A(n12650), .B(n12651), .Z(n12649) );
  OR2_X1 U12591 ( .A1(n8041), .A2(n7746), .ZN(n12437) );
  XOR2_X1 U12592 ( .A(n12652), .B(n12653), .Z(n12434) );
  XOR2_X1 U12593 ( .A(n12654), .B(n12655), .Z(n12653) );
  OR2_X1 U12594 ( .A1(n8037), .A2(n7746), .ZN(n12441) );
  XOR2_X1 U12595 ( .A(n12656), .B(n12657), .Z(n12438) );
  XOR2_X1 U12596 ( .A(n12658), .B(n12659), .Z(n12657) );
  OR2_X1 U12597 ( .A1(n8034), .A2(n7746), .ZN(n12445) );
  XOR2_X1 U12598 ( .A(n12660), .B(n12661), .Z(n12442) );
  XOR2_X1 U12599 ( .A(n12662), .B(n12663), .Z(n12661) );
  OR2_X1 U12600 ( .A1(n8030), .A2(n7746), .ZN(n12449) );
  XOR2_X1 U12601 ( .A(n12664), .B(n12665), .Z(n12446) );
  XOR2_X1 U12602 ( .A(n12666), .B(n12667), .Z(n12665) );
  OR2_X1 U12603 ( .A1(n8026), .A2(n7746), .ZN(n12453) );
  XOR2_X1 U12604 ( .A(n12668), .B(n12669), .Z(n12450) );
  XOR2_X1 U12605 ( .A(n12670), .B(n12671), .Z(n12669) );
  OR2_X1 U12606 ( .A1(n8023), .A2(n7746), .ZN(n12457) );
  XOR2_X1 U12607 ( .A(n12672), .B(n12673), .Z(n12454) );
  XOR2_X1 U12608 ( .A(n12674), .B(n12675), .Z(n12673) );
  OR2_X1 U12609 ( .A1(n8019), .A2(n7746), .ZN(n12461) );
  XOR2_X1 U12610 ( .A(n12676), .B(n12677), .Z(n12458) );
  XOR2_X1 U12611 ( .A(n12678), .B(n12679), .Z(n12677) );
  OR2_X1 U12612 ( .A1(n8016), .A2(n7746), .ZN(n12465) );
  XOR2_X1 U12613 ( .A(n12680), .B(n12681), .Z(n12462) );
  XOR2_X1 U12614 ( .A(n12682), .B(n12683), .Z(n12681) );
  OR2_X1 U12615 ( .A1(n8012), .A2(n7746), .ZN(n12469) );
  XOR2_X1 U12616 ( .A(n12684), .B(n12685), .Z(n12466) );
  XOR2_X1 U12617 ( .A(n12686), .B(n12687), .Z(n12685) );
  OR2_X1 U12618 ( .A1(n8009), .A2(n7746), .ZN(n12473) );
  XOR2_X1 U12619 ( .A(n12688), .B(n12689), .Z(n12470) );
  XOR2_X1 U12620 ( .A(n12690), .B(n12691), .Z(n12689) );
  OR2_X1 U12621 ( .A1(n8005), .A2(n7746), .ZN(n12477) );
  XOR2_X1 U12622 ( .A(n12692), .B(n12693), .Z(n12474) );
  XOR2_X1 U12623 ( .A(n12694), .B(n12695), .Z(n12693) );
  OR2_X1 U12624 ( .A1(n8002), .A2(n7746), .ZN(n12481) );
  XOR2_X1 U12625 ( .A(n12696), .B(n12697), .Z(n12478) );
  XOR2_X1 U12626 ( .A(n12698), .B(n12699), .Z(n12697) );
  OR2_X1 U12627 ( .A1(n7998), .A2(n7746), .ZN(n12485) );
  XOR2_X1 U12628 ( .A(n12700), .B(n12701), .Z(n12482) );
  XOR2_X1 U12629 ( .A(n12702), .B(n12703), .Z(n12701) );
  INV_X1 U12630 ( .A(n7750), .ZN(n7996) );
  AND2_X1 U12631 ( .A1(a_13_), .A2(b_13_), .ZN(n7750) );
  XOR2_X1 U12632 ( .A(n12704), .B(n12705), .Z(n12486) );
  XOR2_X1 U12633 ( .A(n12706), .B(n12707), .Z(n12705) );
  OR2_X1 U12634 ( .A1(n7991), .A2(n7746), .ZN(n12492) );
  XOR2_X1 U12635 ( .A(n12708), .B(n12709), .Z(n12489) );
  XOR2_X1 U12636 ( .A(n12710), .B(n12711), .Z(n12709) );
  OR2_X1 U12637 ( .A1(n7988), .A2(n7746), .ZN(n12496) );
  XNOR2_X1 U12638 ( .A(n12712), .B(n12713), .ZN(n12493) );
  XNOR2_X1 U12639 ( .A(n7993), .B(n12714), .ZN(n12712) );
  OR2_X1 U12640 ( .A1(n7984), .A2(n7746), .ZN(n12500) );
  XOR2_X1 U12641 ( .A(n12715), .B(n12716), .Z(n12497) );
  XOR2_X1 U12642 ( .A(n12717), .B(n12718), .Z(n12716) );
  OR2_X1 U12643 ( .A1(n7981), .A2(n7746), .ZN(n12504) );
  XOR2_X1 U12644 ( .A(n12719), .B(n12720), .Z(n12501) );
  XOR2_X1 U12645 ( .A(n12721), .B(n12722), .Z(n12720) );
  OR2_X1 U12646 ( .A1(n7977), .A2(n7746), .ZN(n12508) );
  XOR2_X1 U12647 ( .A(n12723), .B(n12724), .Z(n12505) );
  XOR2_X1 U12648 ( .A(n12725), .B(n12726), .Z(n12724) );
  OR2_X1 U12649 ( .A1(n7974), .A2(n7746), .ZN(n12512) );
  XOR2_X1 U12650 ( .A(n12727), .B(n12728), .Z(n12509) );
  XOR2_X1 U12651 ( .A(n12729), .B(n12730), .Z(n12728) );
  OR2_X1 U12652 ( .A1(n7970), .A2(n7746), .ZN(n12516) );
  XOR2_X1 U12653 ( .A(n12731), .B(n12732), .Z(n12513) );
  XOR2_X1 U12654 ( .A(n12733), .B(n12734), .Z(n12732) );
  OR2_X1 U12655 ( .A1(n7967), .A2(n7746), .ZN(n12520) );
  XOR2_X1 U12656 ( .A(n12735), .B(n12736), .Z(n12517) );
  XOR2_X1 U12657 ( .A(n12737), .B(n12738), .Z(n12736) );
  OR2_X1 U12658 ( .A1(n7963), .A2(n7746), .ZN(n12524) );
  XOR2_X1 U12659 ( .A(n12739), .B(n12740), .Z(n12521) );
  XOR2_X1 U12660 ( .A(n12741), .B(n12742), .Z(n12740) );
  OR2_X1 U12661 ( .A1(n7960), .A2(n7746), .ZN(n12528) );
  XOR2_X1 U12662 ( .A(n12743), .B(n12744), .Z(n12525) );
  XOR2_X1 U12663 ( .A(n12745), .B(n12746), .Z(n12744) );
  OR2_X1 U12664 ( .A1(n7956), .A2(n7746), .ZN(n12532) );
  XOR2_X1 U12665 ( .A(n12747), .B(n12748), .Z(n12529) );
  XOR2_X1 U12666 ( .A(n12749), .B(n12750), .Z(n12748) );
  OR2_X1 U12667 ( .A1(n7953), .A2(n7746), .ZN(n12536) );
  XOR2_X1 U12668 ( .A(n12751), .B(n12752), .Z(n12533) );
  XOR2_X1 U12669 ( .A(n12753), .B(n12754), .Z(n12752) );
  OR2_X1 U12670 ( .A1(n7950), .A2(n7746), .ZN(n12540) );
  INV_X1 U12671 ( .A(b_13_), .ZN(n7746) );
  XOR2_X1 U12672 ( .A(n12755), .B(n12756), .Z(n12537) );
  XOR2_X1 U12673 ( .A(n12757), .B(n12758), .Z(n12756) );
  XOR2_X1 U12674 ( .A(n8518), .B(n12759), .Z(n12543) );
  XOR2_X1 U12675 ( .A(n8517), .B(n8516), .Z(n12759) );
  OR2_X1 U12676 ( .A1(n7950), .A2(n7992), .ZN(n8516) );
  OR2_X1 U12677 ( .A1(n12760), .A2(n12761), .ZN(n8517) );
  AND2_X1 U12678 ( .A1(n12758), .A2(n12757), .ZN(n12761) );
  AND2_X1 U12679 ( .A1(n12755), .A2(n12762), .ZN(n12760) );
  OR2_X1 U12680 ( .A1(n12757), .A2(n12758), .ZN(n12762) );
  OR2_X1 U12681 ( .A1(n7953), .A2(n7992), .ZN(n12758) );
  OR2_X1 U12682 ( .A1(n12763), .A2(n12764), .ZN(n12757) );
  AND2_X1 U12683 ( .A1(n12754), .A2(n12753), .ZN(n12764) );
  AND2_X1 U12684 ( .A1(n12751), .A2(n12765), .ZN(n12763) );
  OR2_X1 U12685 ( .A1(n12753), .A2(n12754), .ZN(n12765) );
  OR2_X1 U12686 ( .A1(n7956), .A2(n7992), .ZN(n12754) );
  OR2_X1 U12687 ( .A1(n12766), .A2(n12767), .ZN(n12753) );
  AND2_X1 U12688 ( .A1(n12750), .A2(n12749), .ZN(n12767) );
  AND2_X1 U12689 ( .A1(n12747), .A2(n12768), .ZN(n12766) );
  OR2_X1 U12690 ( .A1(n12749), .A2(n12750), .ZN(n12768) );
  OR2_X1 U12691 ( .A1(n7960), .A2(n7992), .ZN(n12750) );
  OR2_X1 U12692 ( .A1(n12769), .A2(n12770), .ZN(n12749) );
  AND2_X1 U12693 ( .A1(n12746), .A2(n12745), .ZN(n12770) );
  AND2_X1 U12694 ( .A1(n12743), .A2(n12771), .ZN(n12769) );
  OR2_X1 U12695 ( .A1(n12745), .A2(n12746), .ZN(n12771) );
  OR2_X1 U12696 ( .A1(n7963), .A2(n7992), .ZN(n12746) );
  OR2_X1 U12697 ( .A1(n12772), .A2(n12773), .ZN(n12745) );
  AND2_X1 U12698 ( .A1(n12742), .A2(n12741), .ZN(n12773) );
  AND2_X1 U12699 ( .A1(n12739), .A2(n12774), .ZN(n12772) );
  OR2_X1 U12700 ( .A1(n12741), .A2(n12742), .ZN(n12774) );
  OR2_X1 U12701 ( .A1(n7967), .A2(n7992), .ZN(n12742) );
  OR2_X1 U12702 ( .A1(n12775), .A2(n12776), .ZN(n12741) );
  AND2_X1 U12703 ( .A1(n12738), .A2(n12737), .ZN(n12776) );
  AND2_X1 U12704 ( .A1(n12735), .A2(n12777), .ZN(n12775) );
  OR2_X1 U12705 ( .A1(n12737), .A2(n12738), .ZN(n12777) );
  OR2_X1 U12706 ( .A1(n7970), .A2(n7992), .ZN(n12738) );
  OR2_X1 U12707 ( .A1(n12778), .A2(n12779), .ZN(n12737) );
  AND2_X1 U12708 ( .A1(n12734), .A2(n12733), .ZN(n12779) );
  AND2_X1 U12709 ( .A1(n12731), .A2(n12780), .ZN(n12778) );
  OR2_X1 U12710 ( .A1(n12733), .A2(n12734), .ZN(n12780) );
  OR2_X1 U12711 ( .A1(n7974), .A2(n7992), .ZN(n12734) );
  OR2_X1 U12712 ( .A1(n12781), .A2(n12782), .ZN(n12733) );
  AND2_X1 U12713 ( .A1(n12730), .A2(n12729), .ZN(n12782) );
  AND2_X1 U12714 ( .A1(n12727), .A2(n12783), .ZN(n12781) );
  OR2_X1 U12715 ( .A1(n12729), .A2(n12730), .ZN(n12783) );
  OR2_X1 U12716 ( .A1(n7977), .A2(n7992), .ZN(n12730) );
  OR2_X1 U12717 ( .A1(n12784), .A2(n12785), .ZN(n12729) );
  AND2_X1 U12718 ( .A1(n12726), .A2(n12725), .ZN(n12785) );
  AND2_X1 U12719 ( .A1(n12723), .A2(n12786), .ZN(n12784) );
  OR2_X1 U12720 ( .A1(n12725), .A2(n12726), .ZN(n12786) );
  OR2_X1 U12721 ( .A1(n7981), .A2(n7992), .ZN(n12726) );
  OR2_X1 U12722 ( .A1(n12787), .A2(n12788), .ZN(n12725) );
  AND2_X1 U12723 ( .A1(n12722), .A2(n12721), .ZN(n12788) );
  AND2_X1 U12724 ( .A1(n12719), .A2(n12789), .ZN(n12787) );
  OR2_X1 U12725 ( .A1(n12721), .A2(n12722), .ZN(n12789) );
  OR2_X1 U12726 ( .A1(n7984), .A2(n7992), .ZN(n12722) );
  OR2_X1 U12727 ( .A1(n12790), .A2(n12791), .ZN(n12721) );
  AND2_X1 U12728 ( .A1(n12718), .A2(n12717), .ZN(n12791) );
  AND2_X1 U12729 ( .A1(n12715), .A2(n12792), .ZN(n12790) );
  OR2_X1 U12730 ( .A1(n12717), .A2(n12718), .ZN(n12792) );
  OR2_X1 U12731 ( .A1(n7988), .A2(n7992), .ZN(n12718) );
  OR2_X1 U12732 ( .A1(n12793), .A2(n12794), .ZN(n12717) );
  AND2_X1 U12733 ( .A1(n12714), .A2(n7993), .ZN(n12794) );
  AND2_X1 U12734 ( .A1(n12713), .A2(n12795), .ZN(n12793) );
  OR2_X1 U12735 ( .A1(n7993), .A2(n12714), .ZN(n12795) );
  OR2_X1 U12736 ( .A1(n12796), .A2(n12797), .ZN(n12714) );
  AND2_X1 U12737 ( .A1(n12711), .A2(n12710), .ZN(n12797) );
  AND2_X1 U12738 ( .A1(n12708), .A2(n12798), .ZN(n12796) );
  OR2_X1 U12739 ( .A1(n12710), .A2(n12711), .ZN(n12798) );
  OR2_X1 U12740 ( .A1(n7995), .A2(n7992), .ZN(n12711) );
  OR2_X1 U12741 ( .A1(n12799), .A2(n12800), .ZN(n12710) );
  AND2_X1 U12742 ( .A1(n12707), .A2(n12706), .ZN(n12800) );
  AND2_X1 U12743 ( .A1(n12704), .A2(n12801), .ZN(n12799) );
  OR2_X1 U12744 ( .A1(n12706), .A2(n12707), .ZN(n12801) );
  OR2_X1 U12745 ( .A1(n7998), .A2(n7992), .ZN(n12707) );
  OR2_X1 U12746 ( .A1(n12802), .A2(n12803), .ZN(n12706) );
  AND2_X1 U12747 ( .A1(n12703), .A2(n12702), .ZN(n12803) );
  AND2_X1 U12748 ( .A1(n12700), .A2(n12804), .ZN(n12802) );
  OR2_X1 U12749 ( .A1(n12702), .A2(n12703), .ZN(n12804) );
  OR2_X1 U12750 ( .A1(n8002), .A2(n7992), .ZN(n12703) );
  OR2_X1 U12751 ( .A1(n12805), .A2(n12806), .ZN(n12702) );
  AND2_X1 U12752 ( .A1(n12699), .A2(n12698), .ZN(n12806) );
  AND2_X1 U12753 ( .A1(n12696), .A2(n12807), .ZN(n12805) );
  OR2_X1 U12754 ( .A1(n12698), .A2(n12699), .ZN(n12807) );
  OR2_X1 U12755 ( .A1(n8005), .A2(n7992), .ZN(n12699) );
  OR2_X1 U12756 ( .A1(n12808), .A2(n12809), .ZN(n12698) );
  AND2_X1 U12757 ( .A1(n12695), .A2(n12694), .ZN(n12809) );
  AND2_X1 U12758 ( .A1(n12692), .A2(n12810), .ZN(n12808) );
  OR2_X1 U12759 ( .A1(n12694), .A2(n12695), .ZN(n12810) );
  OR2_X1 U12760 ( .A1(n8009), .A2(n7992), .ZN(n12695) );
  OR2_X1 U12761 ( .A1(n12811), .A2(n12812), .ZN(n12694) );
  AND2_X1 U12762 ( .A1(n12691), .A2(n12690), .ZN(n12812) );
  AND2_X1 U12763 ( .A1(n12688), .A2(n12813), .ZN(n12811) );
  OR2_X1 U12764 ( .A1(n12690), .A2(n12691), .ZN(n12813) );
  OR2_X1 U12765 ( .A1(n8012), .A2(n7992), .ZN(n12691) );
  OR2_X1 U12766 ( .A1(n12814), .A2(n12815), .ZN(n12690) );
  AND2_X1 U12767 ( .A1(n12687), .A2(n12686), .ZN(n12815) );
  AND2_X1 U12768 ( .A1(n12684), .A2(n12816), .ZN(n12814) );
  OR2_X1 U12769 ( .A1(n12686), .A2(n12687), .ZN(n12816) );
  OR2_X1 U12770 ( .A1(n8016), .A2(n7992), .ZN(n12687) );
  OR2_X1 U12771 ( .A1(n12817), .A2(n12818), .ZN(n12686) );
  AND2_X1 U12772 ( .A1(n12683), .A2(n12682), .ZN(n12818) );
  AND2_X1 U12773 ( .A1(n12680), .A2(n12819), .ZN(n12817) );
  OR2_X1 U12774 ( .A1(n12682), .A2(n12683), .ZN(n12819) );
  OR2_X1 U12775 ( .A1(n8019), .A2(n7992), .ZN(n12683) );
  OR2_X1 U12776 ( .A1(n12820), .A2(n12821), .ZN(n12682) );
  AND2_X1 U12777 ( .A1(n12679), .A2(n12678), .ZN(n12821) );
  AND2_X1 U12778 ( .A1(n12676), .A2(n12822), .ZN(n12820) );
  OR2_X1 U12779 ( .A1(n12678), .A2(n12679), .ZN(n12822) );
  OR2_X1 U12780 ( .A1(n8023), .A2(n7992), .ZN(n12679) );
  OR2_X1 U12781 ( .A1(n12823), .A2(n12824), .ZN(n12678) );
  AND2_X1 U12782 ( .A1(n12675), .A2(n12674), .ZN(n12824) );
  AND2_X1 U12783 ( .A1(n12672), .A2(n12825), .ZN(n12823) );
  OR2_X1 U12784 ( .A1(n12674), .A2(n12675), .ZN(n12825) );
  OR2_X1 U12785 ( .A1(n8026), .A2(n7992), .ZN(n12675) );
  OR2_X1 U12786 ( .A1(n12826), .A2(n12827), .ZN(n12674) );
  AND2_X1 U12787 ( .A1(n12671), .A2(n12670), .ZN(n12827) );
  AND2_X1 U12788 ( .A1(n12668), .A2(n12828), .ZN(n12826) );
  OR2_X1 U12789 ( .A1(n12670), .A2(n12671), .ZN(n12828) );
  OR2_X1 U12790 ( .A1(n8030), .A2(n7992), .ZN(n12671) );
  OR2_X1 U12791 ( .A1(n12829), .A2(n12830), .ZN(n12670) );
  AND2_X1 U12792 ( .A1(n12667), .A2(n12666), .ZN(n12830) );
  AND2_X1 U12793 ( .A1(n12664), .A2(n12831), .ZN(n12829) );
  OR2_X1 U12794 ( .A1(n12666), .A2(n12667), .ZN(n12831) );
  OR2_X1 U12795 ( .A1(n8034), .A2(n7992), .ZN(n12667) );
  OR2_X1 U12796 ( .A1(n12832), .A2(n12833), .ZN(n12666) );
  AND2_X1 U12797 ( .A1(n12663), .A2(n12662), .ZN(n12833) );
  AND2_X1 U12798 ( .A1(n12660), .A2(n12834), .ZN(n12832) );
  OR2_X1 U12799 ( .A1(n12662), .A2(n12663), .ZN(n12834) );
  OR2_X1 U12800 ( .A1(n8037), .A2(n7992), .ZN(n12663) );
  OR2_X1 U12801 ( .A1(n12835), .A2(n12836), .ZN(n12662) );
  AND2_X1 U12802 ( .A1(n12659), .A2(n12658), .ZN(n12836) );
  AND2_X1 U12803 ( .A1(n12656), .A2(n12837), .ZN(n12835) );
  OR2_X1 U12804 ( .A1(n12658), .A2(n12659), .ZN(n12837) );
  OR2_X1 U12805 ( .A1(n8041), .A2(n7992), .ZN(n12659) );
  OR2_X1 U12806 ( .A1(n12838), .A2(n12839), .ZN(n12658) );
  AND2_X1 U12807 ( .A1(n12655), .A2(n12654), .ZN(n12839) );
  AND2_X1 U12808 ( .A1(n12652), .A2(n12840), .ZN(n12838) );
  OR2_X1 U12809 ( .A1(n12654), .A2(n12655), .ZN(n12840) );
  OR2_X1 U12810 ( .A1(n8044), .A2(n7992), .ZN(n12655) );
  OR2_X1 U12811 ( .A1(n12841), .A2(n12842), .ZN(n12654) );
  AND2_X1 U12812 ( .A1(n12651), .A2(n12650), .ZN(n12842) );
  AND2_X1 U12813 ( .A1(n12648), .A2(n12843), .ZN(n12841) );
  OR2_X1 U12814 ( .A1(n12650), .A2(n12651), .ZN(n12843) );
  OR2_X1 U12815 ( .A1(n8048), .A2(n7992), .ZN(n12651) );
  OR2_X1 U12816 ( .A1(n12844), .A2(n12845), .ZN(n12650) );
  AND2_X1 U12817 ( .A1(n12644), .A2(n12846), .ZN(n12845) );
  AND2_X1 U12818 ( .A1(n12847), .A2(n12848), .ZN(n12844) );
  OR2_X1 U12819 ( .A1(n12846), .A2(n12644), .ZN(n12848) );
  OR2_X1 U12820 ( .A1(n8051), .A2(n7992), .ZN(n12644) );
  INV_X1 U12821 ( .A(b_12_), .ZN(n7992) );
  INV_X1 U12822 ( .A(n12647), .ZN(n12846) );
  AND3_X1 U12823 ( .A1(n8904), .A2(b_11_), .A3(b_12_), .ZN(n12647) );
  INV_X1 U12824 ( .A(n12646), .ZN(n12847) );
  OR2_X1 U12825 ( .A1(n12849), .A2(n12850), .ZN(n12646) );
  AND2_X1 U12826 ( .A1(b_11_), .A2(n12851), .ZN(n12850) );
  OR2_X1 U12827 ( .A1(n12852), .A2(n7490), .ZN(n12851) );
  AND2_X1 U12828 ( .A1(a_30_), .A2(n7985), .ZN(n12852) );
  AND2_X1 U12829 ( .A1(b_10_), .A2(n12853), .ZN(n12849) );
  OR2_X1 U12830 ( .A1(n12854), .A2(n7493), .ZN(n12853) );
  AND2_X1 U12831 ( .A1(a_31_), .A2(n7775), .ZN(n12854) );
  XNOR2_X1 U12832 ( .A(n12855), .B(n12856), .ZN(n12648) );
  XNOR2_X1 U12833 ( .A(n12857), .B(n12858), .ZN(n12856) );
  XOR2_X1 U12834 ( .A(n12859), .B(n12860), .Z(n12652) );
  XOR2_X1 U12835 ( .A(n12861), .B(n12862), .Z(n12860) );
  XOR2_X1 U12836 ( .A(n12863), .B(n12864), .Z(n12656) );
  XOR2_X1 U12837 ( .A(n12865), .B(n12866), .Z(n12864) );
  XOR2_X1 U12838 ( .A(n12867), .B(n12868), .Z(n12660) );
  XOR2_X1 U12839 ( .A(n12869), .B(n12870), .Z(n12868) );
  XOR2_X1 U12840 ( .A(n12871), .B(n12872), .Z(n12664) );
  XOR2_X1 U12841 ( .A(n12873), .B(n12874), .Z(n12872) );
  XOR2_X1 U12842 ( .A(n12875), .B(n12876), .Z(n12668) );
  XOR2_X1 U12843 ( .A(n12877), .B(n12878), .Z(n12876) );
  XOR2_X1 U12844 ( .A(n12879), .B(n12880), .Z(n12672) );
  XOR2_X1 U12845 ( .A(n12881), .B(n12882), .Z(n12880) );
  XOR2_X1 U12846 ( .A(n12883), .B(n12884), .Z(n12676) );
  XOR2_X1 U12847 ( .A(n12885), .B(n12886), .Z(n12884) );
  XOR2_X1 U12848 ( .A(n12887), .B(n12888), .Z(n12680) );
  XOR2_X1 U12849 ( .A(n12889), .B(n12890), .Z(n12888) );
  XOR2_X1 U12850 ( .A(n12891), .B(n12892), .Z(n12684) );
  XOR2_X1 U12851 ( .A(n12893), .B(n12894), .Z(n12892) );
  XOR2_X1 U12852 ( .A(n12895), .B(n12896), .Z(n12688) );
  XOR2_X1 U12853 ( .A(n12897), .B(n12898), .Z(n12896) );
  XOR2_X1 U12854 ( .A(n12899), .B(n12900), .Z(n12692) );
  XOR2_X1 U12855 ( .A(n12901), .B(n12902), .Z(n12900) );
  XOR2_X1 U12856 ( .A(n12903), .B(n12904), .Z(n12696) );
  XOR2_X1 U12857 ( .A(n12905), .B(n12906), .Z(n12904) );
  XOR2_X1 U12858 ( .A(n12907), .B(n12908), .Z(n12700) );
  XOR2_X1 U12859 ( .A(n12909), .B(n12910), .Z(n12908) );
  XOR2_X1 U12860 ( .A(n12911), .B(n12912), .Z(n12704) );
  XOR2_X1 U12861 ( .A(n12913), .B(n12914), .Z(n12912) );
  XOR2_X1 U12862 ( .A(n12915), .B(n12916), .Z(n12708) );
  XOR2_X1 U12863 ( .A(n12917), .B(n12918), .Z(n12916) );
  INV_X1 U12864 ( .A(n7767), .ZN(n7993) );
  AND2_X1 U12865 ( .A1(a_12_), .A2(b_12_), .ZN(n7767) );
  XOR2_X1 U12866 ( .A(n12919), .B(n12920), .Z(n12713) );
  XOR2_X1 U12867 ( .A(n12921), .B(n12922), .Z(n12920) );
  XOR2_X1 U12868 ( .A(n12923), .B(n12924), .Z(n12715) );
  XOR2_X1 U12869 ( .A(n12925), .B(n12926), .Z(n12924) );
  XOR2_X1 U12870 ( .A(n12927), .B(n12928), .Z(n12719) );
  XNOR2_X1 U12871 ( .A(n12929), .B(n7779), .ZN(n12928) );
  XOR2_X1 U12872 ( .A(n12930), .B(n12931), .Z(n12723) );
  XOR2_X1 U12873 ( .A(n12932), .B(n12933), .Z(n12931) );
  XOR2_X1 U12874 ( .A(n12934), .B(n12935), .Z(n12727) );
  XOR2_X1 U12875 ( .A(n12936), .B(n12937), .Z(n12935) );
  XOR2_X1 U12876 ( .A(n12938), .B(n12939), .Z(n12731) );
  XOR2_X1 U12877 ( .A(n12940), .B(n12941), .Z(n12939) );
  XOR2_X1 U12878 ( .A(n12942), .B(n12943), .Z(n12735) );
  XOR2_X1 U12879 ( .A(n12944), .B(n12945), .Z(n12943) );
  XOR2_X1 U12880 ( .A(n12946), .B(n12947), .Z(n12739) );
  XOR2_X1 U12881 ( .A(n12948), .B(n12949), .Z(n12947) );
  XOR2_X1 U12882 ( .A(n12950), .B(n12951), .Z(n12743) );
  XOR2_X1 U12883 ( .A(n12952), .B(n12953), .Z(n12951) );
  XOR2_X1 U12884 ( .A(n12954), .B(n12955), .Z(n12747) );
  XOR2_X1 U12885 ( .A(n12956), .B(n12957), .Z(n12955) );
  XOR2_X1 U12886 ( .A(n12958), .B(n12959), .Z(n12751) );
  XOR2_X1 U12887 ( .A(n12960), .B(n12961), .Z(n12959) );
  XOR2_X1 U12888 ( .A(n12962), .B(n12963), .Z(n12755) );
  XOR2_X1 U12889 ( .A(n12964), .B(n12965), .Z(n12963) );
  XOR2_X1 U12890 ( .A(n12966), .B(n12967), .Z(n8518) );
  XOR2_X1 U12891 ( .A(n12968), .B(n12969), .Z(n12967) );
  INV_X1 U12892 ( .A(n12970), .ZN(n8506) );
  OR2_X1 U12893 ( .A1(n8512), .A2(n8513), .ZN(n12970) );
  OR2_X1 U12894 ( .A1(n12971), .A2(n12972), .ZN(n8513) );
  AND2_X1 U12895 ( .A1(n8523), .A2(n8522), .ZN(n12972) );
  AND2_X1 U12896 ( .A1(n8520), .A2(n12973), .ZN(n12971) );
  OR2_X1 U12897 ( .A1(n8523), .A2(n8522), .ZN(n12973) );
  OR2_X1 U12898 ( .A1(n12974), .A2(n12975), .ZN(n8522) );
  AND2_X1 U12899 ( .A1(n12969), .A2(n12968), .ZN(n12975) );
  AND2_X1 U12900 ( .A1(n12966), .A2(n12976), .ZN(n12974) );
  OR2_X1 U12901 ( .A1(n12969), .A2(n12968), .ZN(n12976) );
  OR2_X1 U12902 ( .A1(n12977), .A2(n12978), .ZN(n12968) );
  AND2_X1 U12903 ( .A1(n12965), .A2(n12964), .ZN(n12978) );
  AND2_X1 U12904 ( .A1(n12962), .A2(n12979), .ZN(n12977) );
  OR2_X1 U12905 ( .A1(n12965), .A2(n12964), .ZN(n12979) );
  OR2_X1 U12906 ( .A1(n12980), .A2(n12981), .ZN(n12964) );
  AND2_X1 U12907 ( .A1(n12961), .A2(n12960), .ZN(n12981) );
  AND2_X1 U12908 ( .A1(n12958), .A2(n12982), .ZN(n12980) );
  OR2_X1 U12909 ( .A1(n12961), .A2(n12960), .ZN(n12982) );
  OR2_X1 U12910 ( .A1(n12983), .A2(n12984), .ZN(n12960) );
  AND2_X1 U12911 ( .A1(n12957), .A2(n12956), .ZN(n12984) );
  AND2_X1 U12912 ( .A1(n12954), .A2(n12985), .ZN(n12983) );
  OR2_X1 U12913 ( .A1(n12957), .A2(n12956), .ZN(n12985) );
  OR2_X1 U12914 ( .A1(n12986), .A2(n12987), .ZN(n12956) );
  AND2_X1 U12915 ( .A1(n12953), .A2(n12952), .ZN(n12987) );
  AND2_X1 U12916 ( .A1(n12950), .A2(n12988), .ZN(n12986) );
  OR2_X1 U12917 ( .A1(n12953), .A2(n12952), .ZN(n12988) );
  OR2_X1 U12918 ( .A1(n12989), .A2(n12990), .ZN(n12952) );
  AND2_X1 U12919 ( .A1(n12949), .A2(n12948), .ZN(n12990) );
  AND2_X1 U12920 ( .A1(n12946), .A2(n12991), .ZN(n12989) );
  OR2_X1 U12921 ( .A1(n12949), .A2(n12948), .ZN(n12991) );
  OR2_X1 U12922 ( .A1(n12992), .A2(n12993), .ZN(n12948) );
  AND2_X1 U12923 ( .A1(n12945), .A2(n12944), .ZN(n12993) );
  AND2_X1 U12924 ( .A1(n12942), .A2(n12994), .ZN(n12992) );
  OR2_X1 U12925 ( .A1(n12945), .A2(n12944), .ZN(n12994) );
  OR2_X1 U12926 ( .A1(n12995), .A2(n12996), .ZN(n12944) );
  AND2_X1 U12927 ( .A1(n12941), .A2(n12940), .ZN(n12996) );
  AND2_X1 U12928 ( .A1(n12938), .A2(n12997), .ZN(n12995) );
  OR2_X1 U12929 ( .A1(n12941), .A2(n12940), .ZN(n12997) );
  OR2_X1 U12930 ( .A1(n12998), .A2(n12999), .ZN(n12940) );
  AND2_X1 U12931 ( .A1(n12937), .A2(n12936), .ZN(n12999) );
  AND2_X1 U12932 ( .A1(n12934), .A2(n13000), .ZN(n12998) );
  OR2_X1 U12933 ( .A1(n12937), .A2(n12936), .ZN(n13000) );
  OR2_X1 U12934 ( .A1(n13001), .A2(n13002), .ZN(n12936) );
  AND2_X1 U12935 ( .A1(n12933), .A2(n12932), .ZN(n13002) );
  AND2_X1 U12936 ( .A1(n12930), .A2(n13003), .ZN(n13001) );
  OR2_X1 U12937 ( .A1(n12933), .A2(n12932), .ZN(n13003) );
  OR2_X1 U12938 ( .A1(n13004), .A2(n13005), .ZN(n12932) );
  AND2_X1 U12939 ( .A1(n7989), .A2(n12929), .ZN(n13005) );
  AND2_X1 U12940 ( .A1(n12927), .A2(n13006), .ZN(n13004) );
  OR2_X1 U12941 ( .A1(n7989), .A2(n12929), .ZN(n13006) );
  OR2_X1 U12942 ( .A1(n13007), .A2(n13008), .ZN(n12929) );
  AND2_X1 U12943 ( .A1(n12926), .A2(n12925), .ZN(n13008) );
  AND2_X1 U12944 ( .A1(n12923), .A2(n13009), .ZN(n13007) );
  OR2_X1 U12945 ( .A1(n12926), .A2(n12925), .ZN(n13009) );
  OR2_X1 U12946 ( .A1(n13010), .A2(n13011), .ZN(n12925) );
  AND2_X1 U12947 ( .A1(n12922), .A2(n12921), .ZN(n13011) );
  AND2_X1 U12948 ( .A1(n12919), .A2(n13012), .ZN(n13010) );
  OR2_X1 U12949 ( .A1(n12922), .A2(n12921), .ZN(n13012) );
  OR2_X1 U12950 ( .A1(n13013), .A2(n13014), .ZN(n12921) );
  AND2_X1 U12951 ( .A1(n12918), .A2(n12917), .ZN(n13014) );
  AND2_X1 U12952 ( .A1(n12915), .A2(n13015), .ZN(n13013) );
  OR2_X1 U12953 ( .A1(n12918), .A2(n12917), .ZN(n13015) );
  OR2_X1 U12954 ( .A1(n13016), .A2(n13017), .ZN(n12917) );
  AND2_X1 U12955 ( .A1(n12914), .A2(n12913), .ZN(n13017) );
  AND2_X1 U12956 ( .A1(n12911), .A2(n13018), .ZN(n13016) );
  OR2_X1 U12957 ( .A1(n12914), .A2(n12913), .ZN(n13018) );
  OR2_X1 U12958 ( .A1(n13019), .A2(n13020), .ZN(n12913) );
  AND2_X1 U12959 ( .A1(n12910), .A2(n12909), .ZN(n13020) );
  AND2_X1 U12960 ( .A1(n12907), .A2(n13021), .ZN(n13019) );
  OR2_X1 U12961 ( .A1(n12910), .A2(n12909), .ZN(n13021) );
  OR2_X1 U12962 ( .A1(n13022), .A2(n13023), .ZN(n12909) );
  AND2_X1 U12963 ( .A1(n12906), .A2(n12905), .ZN(n13023) );
  AND2_X1 U12964 ( .A1(n12903), .A2(n13024), .ZN(n13022) );
  OR2_X1 U12965 ( .A1(n12906), .A2(n12905), .ZN(n13024) );
  OR2_X1 U12966 ( .A1(n13025), .A2(n13026), .ZN(n12905) );
  AND2_X1 U12967 ( .A1(n12902), .A2(n12901), .ZN(n13026) );
  AND2_X1 U12968 ( .A1(n12899), .A2(n13027), .ZN(n13025) );
  OR2_X1 U12969 ( .A1(n12902), .A2(n12901), .ZN(n13027) );
  OR2_X1 U12970 ( .A1(n13028), .A2(n13029), .ZN(n12901) );
  AND2_X1 U12971 ( .A1(n12898), .A2(n12897), .ZN(n13029) );
  AND2_X1 U12972 ( .A1(n12895), .A2(n13030), .ZN(n13028) );
  OR2_X1 U12973 ( .A1(n12898), .A2(n12897), .ZN(n13030) );
  OR2_X1 U12974 ( .A1(n13031), .A2(n13032), .ZN(n12897) );
  AND2_X1 U12975 ( .A1(n12894), .A2(n12893), .ZN(n13032) );
  AND2_X1 U12976 ( .A1(n12891), .A2(n13033), .ZN(n13031) );
  OR2_X1 U12977 ( .A1(n12894), .A2(n12893), .ZN(n13033) );
  OR2_X1 U12978 ( .A1(n13034), .A2(n13035), .ZN(n12893) );
  AND2_X1 U12979 ( .A1(n12890), .A2(n12889), .ZN(n13035) );
  AND2_X1 U12980 ( .A1(n12887), .A2(n13036), .ZN(n13034) );
  OR2_X1 U12981 ( .A1(n12890), .A2(n12889), .ZN(n13036) );
  OR2_X1 U12982 ( .A1(n13037), .A2(n13038), .ZN(n12889) );
  AND2_X1 U12983 ( .A1(n12886), .A2(n12885), .ZN(n13038) );
  AND2_X1 U12984 ( .A1(n12883), .A2(n13039), .ZN(n13037) );
  OR2_X1 U12985 ( .A1(n12886), .A2(n12885), .ZN(n13039) );
  OR2_X1 U12986 ( .A1(n13040), .A2(n13041), .ZN(n12885) );
  AND2_X1 U12987 ( .A1(n12882), .A2(n12881), .ZN(n13041) );
  AND2_X1 U12988 ( .A1(n12879), .A2(n13042), .ZN(n13040) );
  OR2_X1 U12989 ( .A1(n12882), .A2(n12881), .ZN(n13042) );
  OR2_X1 U12990 ( .A1(n13043), .A2(n13044), .ZN(n12881) );
  AND2_X1 U12991 ( .A1(n12878), .A2(n12877), .ZN(n13044) );
  AND2_X1 U12992 ( .A1(n12875), .A2(n13045), .ZN(n13043) );
  OR2_X1 U12993 ( .A1(n12878), .A2(n12877), .ZN(n13045) );
  OR2_X1 U12994 ( .A1(n13046), .A2(n13047), .ZN(n12877) );
  AND2_X1 U12995 ( .A1(n12874), .A2(n12873), .ZN(n13047) );
  AND2_X1 U12996 ( .A1(n12871), .A2(n13048), .ZN(n13046) );
  OR2_X1 U12997 ( .A1(n12874), .A2(n12873), .ZN(n13048) );
  OR2_X1 U12998 ( .A1(n13049), .A2(n13050), .ZN(n12873) );
  AND2_X1 U12999 ( .A1(n12870), .A2(n12869), .ZN(n13050) );
  AND2_X1 U13000 ( .A1(n12867), .A2(n13051), .ZN(n13049) );
  OR2_X1 U13001 ( .A1(n12870), .A2(n12869), .ZN(n13051) );
  OR2_X1 U13002 ( .A1(n13052), .A2(n13053), .ZN(n12869) );
  AND2_X1 U13003 ( .A1(n12866), .A2(n12865), .ZN(n13053) );
  AND2_X1 U13004 ( .A1(n12863), .A2(n13054), .ZN(n13052) );
  OR2_X1 U13005 ( .A1(n12866), .A2(n12865), .ZN(n13054) );
  OR2_X1 U13006 ( .A1(n13055), .A2(n13056), .ZN(n12865) );
  AND2_X1 U13007 ( .A1(n12862), .A2(n12861), .ZN(n13056) );
  AND2_X1 U13008 ( .A1(n12859), .A2(n13057), .ZN(n13055) );
  OR2_X1 U13009 ( .A1(n12862), .A2(n12861), .ZN(n13057) );
  OR2_X1 U13010 ( .A1(n13058), .A2(n13059), .ZN(n12861) );
  AND2_X1 U13011 ( .A1(n12855), .A2(n13060), .ZN(n13059) );
  AND2_X1 U13012 ( .A1(n13061), .A2(n13062), .ZN(n13058) );
  OR2_X1 U13013 ( .A1(n12855), .A2(n13060), .ZN(n13062) );
  INV_X1 U13014 ( .A(n12858), .ZN(n13060) );
  AND3_X1 U13015 ( .A1(b_10_), .A2(n8904), .A3(b_11_), .ZN(n12858) );
  OR2_X1 U13016 ( .A1(n7775), .A2(n8051), .ZN(n12855) );
  INV_X1 U13017 ( .A(n12857), .ZN(n13061) );
  OR2_X1 U13018 ( .A1(n13063), .A2(n13064), .ZN(n12857) );
  AND2_X1 U13019 ( .A1(b_9_), .A2(n13065), .ZN(n13064) );
  OR2_X1 U13020 ( .A1(n13066), .A2(n7493), .ZN(n13065) );
  AND2_X1 U13021 ( .A1(a_31_), .A2(n7985), .ZN(n13066) );
  AND2_X1 U13022 ( .A1(b_10_), .A2(n13067), .ZN(n13063) );
  OR2_X1 U13023 ( .A1(n13068), .A2(n7490), .ZN(n13067) );
  AND2_X1 U13024 ( .A1(a_30_), .A2(n7804), .ZN(n13068) );
  OR2_X1 U13025 ( .A1(n7775), .A2(n8048), .ZN(n12862) );
  XNOR2_X1 U13026 ( .A(n13069), .B(n13070), .ZN(n12859) );
  XNOR2_X1 U13027 ( .A(n13071), .B(n13072), .ZN(n13070) );
  OR2_X1 U13028 ( .A1(n7775), .A2(n8044), .ZN(n12866) );
  XOR2_X1 U13029 ( .A(n13073), .B(n13074), .Z(n12863) );
  XOR2_X1 U13030 ( .A(n13075), .B(n13076), .Z(n13074) );
  OR2_X1 U13031 ( .A1(n7775), .A2(n8041), .ZN(n12870) );
  XOR2_X1 U13032 ( .A(n13077), .B(n13078), .Z(n12867) );
  XOR2_X1 U13033 ( .A(n13079), .B(n13080), .Z(n13078) );
  OR2_X1 U13034 ( .A1(n7775), .A2(n8037), .ZN(n12874) );
  XOR2_X1 U13035 ( .A(n13081), .B(n13082), .Z(n12871) );
  XOR2_X1 U13036 ( .A(n13083), .B(n13084), .Z(n13082) );
  OR2_X1 U13037 ( .A1(n7775), .A2(n8034), .ZN(n12878) );
  XOR2_X1 U13038 ( .A(n13085), .B(n13086), .Z(n12875) );
  XOR2_X1 U13039 ( .A(n13087), .B(n13088), .Z(n13086) );
  OR2_X1 U13040 ( .A1(n7775), .A2(n8030), .ZN(n12882) );
  XOR2_X1 U13041 ( .A(n13089), .B(n13090), .Z(n12879) );
  XOR2_X1 U13042 ( .A(n13091), .B(n13092), .Z(n13090) );
  OR2_X1 U13043 ( .A1(n7775), .A2(n8026), .ZN(n12886) );
  XOR2_X1 U13044 ( .A(n13093), .B(n13094), .Z(n12883) );
  XOR2_X1 U13045 ( .A(n13095), .B(n13096), .Z(n13094) );
  OR2_X1 U13046 ( .A1(n7775), .A2(n8023), .ZN(n12890) );
  XOR2_X1 U13047 ( .A(n13097), .B(n13098), .Z(n12887) );
  XOR2_X1 U13048 ( .A(n13099), .B(n13100), .Z(n13098) );
  OR2_X1 U13049 ( .A1(n7775), .A2(n8019), .ZN(n12894) );
  XOR2_X1 U13050 ( .A(n13101), .B(n13102), .Z(n12891) );
  XOR2_X1 U13051 ( .A(n13103), .B(n13104), .Z(n13102) );
  OR2_X1 U13052 ( .A1(n7775), .A2(n8016), .ZN(n12898) );
  XOR2_X1 U13053 ( .A(n13105), .B(n13106), .Z(n12895) );
  XOR2_X1 U13054 ( .A(n13107), .B(n13108), .Z(n13106) );
  OR2_X1 U13055 ( .A1(n7775), .A2(n8012), .ZN(n12902) );
  XOR2_X1 U13056 ( .A(n13109), .B(n13110), .Z(n12899) );
  XOR2_X1 U13057 ( .A(n13111), .B(n13112), .Z(n13110) );
  OR2_X1 U13058 ( .A1(n7775), .A2(n8009), .ZN(n12906) );
  XOR2_X1 U13059 ( .A(n13113), .B(n13114), .Z(n12903) );
  XOR2_X1 U13060 ( .A(n13115), .B(n13116), .Z(n13114) );
  OR2_X1 U13061 ( .A1(n7775), .A2(n8005), .ZN(n12910) );
  XOR2_X1 U13062 ( .A(n13117), .B(n13118), .Z(n12907) );
  XOR2_X1 U13063 ( .A(n13119), .B(n13120), .Z(n13118) );
  OR2_X1 U13064 ( .A1(n7775), .A2(n8002), .ZN(n12914) );
  XOR2_X1 U13065 ( .A(n13121), .B(n13122), .Z(n12911) );
  XOR2_X1 U13066 ( .A(n13123), .B(n13124), .Z(n13122) );
  OR2_X1 U13067 ( .A1(n7775), .A2(n7998), .ZN(n12918) );
  XOR2_X1 U13068 ( .A(n13125), .B(n13126), .Z(n12915) );
  XOR2_X1 U13069 ( .A(n13127), .B(n13128), .Z(n13126) );
  OR2_X1 U13070 ( .A1(n7775), .A2(n7995), .ZN(n12922) );
  XOR2_X1 U13071 ( .A(n13129), .B(n13130), .Z(n12919) );
  XOR2_X1 U13072 ( .A(n13131), .B(n13132), .Z(n13130) );
  OR2_X1 U13073 ( .A1(n7775), .A2(n7991), .ZN(n12926) );
  XOR2_X1 U13074 ( .A(n13133), .B(n13134), .Z(n12923) );
  XOR2_X1 U13075 ( .A(n13135), .B(n13136), .Z(n13134) );
  INV_X1 U13076 ( .A(n7779), .ZN(n7989) );
  AND2_X1 U13077 ( .A1(b_11_), .A2(a_11_), .ZN(n7779) );
  XOR2_X1 U13078 ( .A(n13137), .B(n13138), .Z(n12927) );
  XOR2_X1 U13079 ( .A(n13139), .B(n13140), .Z(n13138) );
  OR2_X1 U13080 ( .A1(n7775), .A2(n7984), .ZN(n12933) );
  XOR2_X1 U13081 ( .A(n13141), .B(n13142), .Z(n12930) );
  XOR2_X1 U13082 ( .A(n13143), .B(n13144), .Z(n13142) );
  OR2_X1 U13083 ( .A1(n7775), .A2(n7981), .ZN(n12937) );
  XNOR2_X1 U13084 ( .A(n13145), .B(n13146), .ZN(n12934) );
  XNOR2_X1 U13085 ( .A(n7986), .B(n13147), .ZN(n13145) );
  OR2_X1 U13086 ( .A1(n7775), .A2(n7977), .ZN(n12941) );
  XOR2_X1 U13087 ( .A(n13148), .B(n13149), .Z(n12938) );
  XOR2_X1 U13088 ( .A(n13150), .B(n13151), .Z(n13149) );
  OR2_X1 U13089 ( .A1(n7775), .A2(n7974), .ZN(n12945) );
  XOR2_X1 U13090 ( .A(n13152), .B(n13153), .Z(n12942) );
  XOR2_X1 U13091 ( .A(n13154), .B(n13155), .Z(n13153) );
  OR2_X1 U13092 ( .A1(n7775), .A2(n7970), .ZN(n12949) );
  XOR2_X1 U13093 ( .A(n13156), .B(n13157), .Z(n12946) );
  XOR2_X1 U13094 ( .A(n13158), .B(n13159), .Z(n13157) );
  OR2_X1 U13095 ( .A1(n7775), .A2(n7967), .ZN(n12953) );
  XOR2_X1 U13096 ( .A(n13160), .B(n13161), .Z(n12950) );
  XOR2_X1 U13097 ( .A(n13162), .B(n13163), .Z(n13161) );
  OR2_X1 U13098 ( .A1(n7775), .A2(n7963), .ZN(n12957) );
  XOR2_X1 U13099 ( .A(n13164), .B(n13165), .Z(n12954) );
  XOR2_X1 U13100 ( .A(n13166), .B(n13167), .Z(n13165) );
  OR2_X1 U13101 ( .A1(n7775), .A2(n7960), .ZN(n12961) );
  XOR2_X1 U13102 ( .A(n13168), .B(n13169), .Z(n12958) );
  XOR2_X1 U13103 ( .A(n13170), .B(n13171), .Z(n13169) );
  OR2_X1 U13104 ( .A1(n7775), .A2(n7956), .ZN(n12965) );
  XOR2_X1 U13105 ( .A(n13172), .B(n13173), .Z(n12962) );
  XOR2_X1 U13106 ( .A(n13174), .B(n13175), .Z(n13173) );
  OR2_X1 U13107 ( .A1(n7775), .A2(n7953), .ZN(n12969) );
  XOR2_X1 U13108 ( .A(n13176), .B(n13177), .Z(n12966) );
  XOR2_X1 U13109 ( .A(n13178), .B(n13179), .Z(n13177) );
  OR2_X1 U13110 ( .A1(n7775), .A2(n7950), .ZN(n8523) );
  INV_X1 U13111 ( .A(b_11_), .ZN(n7775) );
  XOR2_X1 U13112 ( .A(n13180), .B(n13181), .Z(n8520) );
  XOR2_X1 U13113 ( .A(n13182), .B(n13183), .Z(n13181) );
  XOR2_X1 U13114 ( .A(n8452), .B(n13184), .Z(n8512) );
  XOR2_X1 U13115 ( .A(n8451), .B(n8450), .Z(n13184) );
  OR2_X1 U13116 ( .A1(n7985), .A2(n7950), .ZN(n8450) );
  OR2_X1 U13117 ( .A1(n13185), .A2(n13186), .ZN(n8451) );
  AND2_X1 U13118 ( .A1(n13183), .A2(n13182), .ZN(n13186) );
  AND2_X1 U13119 ( .A1(n13180), .A2(n13187), .ZN(n13185) );
  OR2_X1 U13120 ( .A1(n13182), .A2(n13183), .ZN(n13187) );
  OR2_X1 U13121 ( .A1(n7985), .A2(n7953), .ZN(n13183) );
  OR2_X1 U13122 ( .A1(n13188), .A2(n13189), .ZN(n13182) );
  AND2_X1 U13123 ( .A1(n13179), .A2(n13178), .ZN(n13189) );
  AND2_X1 U13124 ( .A1(n13176), .A2(n13190), .ZN(n13188) );
  OR2_X1 U13125 ( .A1(n13178), .A2(n13179), .ZN(n13190) );
  OR2_X1 U13126 ( .A1(n7985), .A2(n7956), .ZN(n13179) );
  OR2_X1 U13127 ( .A1(n13191), .A2(n13192), .ZN(n13178) );
  AND2_X1 U13128 ( .A1(n13175), .A2(n13174), .ZN(n13192) );
  AND2_X1 U13129 ( .A1(n13172), .A2(n13193), .ZN(n13191) );
  OR2_X1 U13130 ( .A1(n13174), .A2(n13175), .ZN(n13193) );
  OR2_X1 U13131 ( .A1(n7985), .A2(n7960), .ZN(n13175) );
  OR2_X1 U13132 ( .A1(n13194), .A2(n13195), .ZN(n13174) );
  AND2_X1 U13133 ( .A1(n13171), .A2(n13170), .ZN(n13195) );
  AND2_X1 U13134 ( .A1(n13168), .A2(n13196), .ZN(n13194) );
  OR2_X1 U13135 ( .A1(n13170), .A2(n13171), .ZN(n13196) );
  OR2_X1 U13136 ( .A1(n7985), .A2(n7963), .ZN(n13171) );
  OR2_X1 U13137 ( .A1(n13197), .A2(n13198), .ZN(n13170) );
  AND2_X1 U13138 ( .A1(n13167), .A2(n13166), .ZN(n13198) );
  AND2_X1 U13139 ( .A1(n13164), .A2(n13199), .ZN(n13197) );
  OR2_X1 U13140 ( .A1(n13166), .A2(n13167), .ZN(n13199) );
  OR2_X1 U13141 ( .A1(n7985), .A2(n7967), .ZN(n13167) );
  OR2_X1 U13142 ( .A1(n13200), .A2(n13201), .ZN(n13166) );
  AND2_X1 U13143 ( .A1(n13163), .A2(n13162), .ZN(n13201) );
  AND2_X1 U13144 ( .A1(n13160), .A2(n13202), .ZN(n13200) );
  OR2_X1 U13145 ( .A1(n13162), .A2(n13163), .ZN(n13202) );
  OR2_X1 U13146 ( .A1(n7985), .A2(n7970), .ZN(n13163) );
  OR2_X1 U13147 ( .A1(n13203), .A2(n13204), .ZN(n13162) );
  AND2_X1 U13148 ( .A1(n13159), .A2(n13158), .ZN(n13204) );
  AND2_X1 U13149 ( .A1(n13156), .A2(n13205), .ZN(n13203) );
  OR2_X1 U13150 ( .A1(n13158), .A2(n13159), .ZN(n13205) );
  OR2_X1 U13151 ( .A1(n7985), .A2(n7974), .ZN(n13159) );
  OR2_X1 U13152 ( .A1(n13206), .A2(n13207), .ZN(n13158) );
  AND2_X1 U13153 ( .A1(n13155), .A2(n13154), .ZN(n13207) );
  AND2_X1 U13154 ( .A1(n13152), .A2(n13208), .ZN(n13206) );
  OR2_X1 U13155 ( .A1(n13154), .A2(n13155), .ZN(n13208) );
  OR2_X1 U13156 ( .A1(n7985), .A2(n7977), .ZN(n13155) );
  OR2_X1 U13157 ( .A1(n13209), .A2(n13210), .ZN(n13154) );
  AND2_X1 U13158 ( .A1(n13151), .A2(n13150), .ZN(n13210) );
  AND2_X1 U13159 ( .A1(n13148), .A2(n13211), .ZN(n13209) );
  OR2_X1 U13160 ( .A1(n13150), .A2(n13151), .ZN(n13211) );
  OR2_X1 U13161 ( .A1(n7985), .A2(n7981), .ZN(n13151) );
  OR2_X1 U13162 ( .A1(n13212), .A2(n13213), .ZN(n13150) );
  AND2_X1 U13163 ( .A1(n13147), .A2(n7986), .ZN(n13213) );
  AND2_X1 U13164 ( .A1(n13146), .A2(n13214), .ZN(n13212) );
  OR2_X1 U13165 ( .A1(n7986), .A2(n13147), .ZN(n13214) );
  OR2_X1 U13166 ( .A1(n13215), .A2(n13216), .ZN(n13147) );
  AND2_X1 U13167 ( .A1(n13144), .A2(n13143), .ZN(n13216) );
  AND2_X1 U13168 ( .A1(n13141), .A2(n13217), .ZN(n13215) );
  OR2_X1 U13169 ( .A1(n13143), .A2(n13144), .ZN(n13217) );
  OR2_X1 U13170 ( .A1(n7985), .A2(n7988), .ZN(n13144) );
  OR2_X1 U13171 ( .A1(n13218), .A2(n13219), .ZN(n13143) );
  AND2_X1 U13172 ( .A1(n13140), .A2(n13139), .ZN(n13219) );
  AND2_X1 U13173 ( .A1(n13137), .A2(n13220), .ZN(n13218) );
  OR2_X1 U13174 ( .A1(n13139), .A2(n13140), .ZN(n13220) );
  OR2_X1 U13175 ( .A1(n7985), .A2(n7991), .ZN(n13140) );
  OR2_X1 U13176 ( .A1(n13221), .A2(n13222), .ZN(n13139) );
  AND2_X1 U13177 ( .A1(n13136), .A2(n13135), .ZN(n13222) );
  AND2_X1 U13178 ( .A1(n13133), .A2(n13223), .ZN(n13221) );
  OR2_X1 U13179 ( .A1(n13135), .A2(n13136), .ZN(n13223) );
  OR2_X1 U13180 ( .A1(n7985), .A2(n7995), .ZN(n13136) );
  OR2_X1 U13181 ( .A1(n13224), .A2(n13225), .ZN(n13135) );
  AND2_X1 U13182 ( .A1(n13132), .A2(n13131), .ZN(n13225) );
  AND2_X1 U13183 ( .A1(n13129), .A2(n13226), .ZN(n13224) );
  OR2_X1 U13184 ( .A1(n13131), .A2(n13132), .ZN(n13226) );
  OR2_X1 U13185 ( .A1(n7985), .A2(n7998), .ZN(n13132) );
  OR2_X1 U13186 ( .A1(n13227), .A2(n13228), .ZN(n13131) );
  AND2_X1 U13187 ( .A1(n13128), .A2(n13127), .ZN(n13228) );
  AND2_X1 U13188 ( .A1(n13125), .A2(n13229), .ZN(n13227) );
  OR2_X1 U13189 ( .A1(n13127), .A2(n13128), .ZN(n13229) );
  OR2_X1 U13190 ( .A1(n7985), .A2(n8002), .ZN(n13128) );
  OR2_X1 U13191 ( .A1(n13230), .A2(n13231), .ZN(n13127) );
  AND2_X1 U13192 ( .A1(n13124), .A2(n13123), .ZN(n13231) );
  AND2_X1 U13193 ( .A1(n13121), .A2(n13232), .ZN(n13230) );
  OR2_X1 U13194 ( .A1(n13123), .A2(n13124), .ZN(n13232) );
  OR2_X1 U13195 ( .A1(n7985), .A2(n8005), .ZN(n13124) );
  OR2_X1 U13196 ( .A1(n13233), .A2(n13234), .ZN(n13123) );
  AND2_X1 U13197 ( .A1(n13120), .A2(n13119), .ZN(n13234) );
  AND2_X1 U13198 ( .A1(n13117), .A2(n13235), .ZN(n13233) );
  OR2_X1 U13199 ( .A1(n13119), .A2(n13120), .ZN(n13235) );
  OR2_X1 U13200 ( .A1(n7985), .A2(n8009), .ZN(n13120) );
  OR2_X1 U13201 ( .A1(n13236), .A2(n13237), .ZN(n13119) );
  AND2_X1 U13202 ( .A1(n13116), .A2(n13115), .ZN(n13237) );
  AND2_X1 U13203 ( .A1(n13113), .A2(n13238), .ZN(n13236) );
  OR2_X1 U13204 ( .A1(n13115), .A2(n13116), .ZN(n13238) );
  OR2_X1 U13205 ( .A1(n7985), .A2(n8012), .ZN(n13116) );
  OR2_X1 U13206 ( .A1(n13239), .A2(n13240), .ZN(n13115) );
  AND2_X1 U13207 ( .A1(n13109), .A2(n13112), .ZN(n13240) );
  AND2_X1 U13208 ( .A1(n13241), .A2(n13111), .ZN(n13239) );
  OR2_X1 U13209 ( .A1(n13242), .A2(n13243), .ZN(n13111) );
  AND2_X1 U13210 ( .A1(n13108), .A2(n13107), .ZN(n13243) );
  AND2_X1 U13211 ( .A1(n13105), .A2(n13244), .ZN(n13242) );
  OR2_X1 U13212 ( .A1(n13107), .A2(n13108), .ZN(n13244) );
  OR2_X1 U13213 ( .A1(n7985), .A2(n8019), .ZN(n13108) );
  OR2_X1 U13214 ( .A1(n13245), .A2(n13246), .ZN(n13107) );
  AND2_X1 U13215 ( .A1(n13101), .A2(n13104), .ZN(n13246) );
  AND2_X1 U13216 ( .A1(n13247), .A2(n13103), .ZN(n13245) );
  OR2_X1 U13217 ( .A1(n13248), .A2(n13249), .ZN(n13103) );
  AND2_X1 U13218 ( .A1(n13097), .A2(n13100), .ZN(n13249) );
  AND2_X1 U13219 ( .A1(n13250), .A2(n13099), .ZN(n13248) );
  OR2_X1 U13220 ( .A1(n13251), .A2(n13252), .ZN(n13099) );
  AND2_X1 U13221 ( .A1(n13093), .A2(n13096), .ZN(n13252) );
  AND2_X1 U13222 ( .A1(n13253), .A2(n13095), .ZN(n13251) );
  OR2_X1 U13223 ( .A1(n13254), .A2(n13255), .ZN(n13095) );
  AND2_X1 U13224 ( .A1(n13089), .A2(n13092), .ZN(n13255) );
  AND2_X1 U13225 ( .A1(n13256), .A2(n13091), .ZN(n13254) );
  OR2_X1 U13226 ( .A1(n13257), .A2(n13258), .ZN(n13091) );
  AND2_X1 U13227 ( .A1(n13085), .A2(n13088), .ZN(n13258) );
  AND2_X1 U13228 ( .A1(n13259), .A2(n13087), .ZN(n13257) );
  OR2_X1 U13229 ( .A1(n13260), .A2(n13261), .ZN(n13087) );
  AND2_X1 U13230 ( .A1(n13081), .A2(n13084), .ZN(n13261) );
  AND2_X1 U13231 ( .A1(n13262), .A2(n13083), .ZN(n13260) );
  OR2_X1 U13232 ( .A1(n13263), .A2(n13264), .ZN(n13083) );
  AND2_X1 U13233 ( .A1(n13077), .A2(n13080), .ZN(n13264) );
  AND2_X1 U13234 ( .A1(n13265), .A2(n13079), .ZN(n13263) );
  OR2_X1 U13235 ( .A1(n13266), .A2(n13267), .ZN(n13079) );
  AND2_X1 U13236 ( .A1(n13073), .A2(n13076), .ZN(n13267) );
  AND2_X1 U13237 ( .A1(n13268), .A2(n13075), .ZN(n13266) );
  OR2_X1 U13238 ( .A1(n13269), .A2(n13270), .ZN(n13075) );
  AND2_X1 U13239 ( .A1(n13069), .A2(n13271), .ZN(n13270) );
  AND2_X1 U13240 ( .A1(n13272), .A2(n13273), .ZN(n13269) );
  OR2_X1 U13241 ( .A1(n13271), .A2(n13069), .ZN(n13273) );
  OR2_X1 U13242 ( .A1(n7985), .A2(n8051), .ZN(n13069) );
  INV_X1 U13243 ( .A(n13072), .ZN(n13271) );
  AND3_X1 U13244 ( .A1(b_10_), .A2(b_9_), .A3(n8904), .ZN(n13072) );
  INV_X1 U13245 ( .A(n13071), .ZN(n13272) );
  OR2_X1 U13246 ( .A1(n13274), .A2(n13275), .ZN(n13071) );
  AND2_X1 U13247 ( .A1(b_9_), .A2(n13276), .ZN(n13275) );
  OR2_X1 U13248 ( .A1(n13277), .A2(n7490), .ZN(n13276) );
  AND2_X1 U13249 ( .A1(a_30_), .A2(n7978), .ZN(n13277) );
  AND2_X1 U13250 ( .A1(b_8_), .A2(n13278), .ZN(n13274) );
  OR2_X1 U13251 ( .A1(n13279), .A2(n7493), .ZN(n13278) );
  AND2_X1 U13252 ( .A1(a_31_), .A2(n7804), .ZN(n13279) );
  OR2_X1 U13253 ( .A1(n13076), .A2(n13073), .ZN(n13268) );
  XNOR2_X1 U13254 ( .A(n13280), .B(n13281), .ZN(n13073) );
  XNOR2_X1 U13255 ( .A(n13282), .B(n13283), .ZN(n13281) );
  OR2_X1 U13256 ( .A1(n7985), .A2(n8048), .ZN(n13076) );
  OR2_X1 U13257 ( .A1(n13080), .A2(n13077), .ZN(n13265) );
  XOR2_X1 U13258 ( .A(n13284), .B(n13285), .Z(n13077) );
  XOR2_X1 U13259 ( .A(n13286), .B(n13287), .Z(n13285) );
  OR2_X1 U13260 ( .A1(n7985), .A2(n8044), .ZN(n13080) );
  OR2_X1 U13261 ( .A1(n13084), .A2(n13081), .ZN(n13262) );
  XOR2_X1 U13262 ( .A(n13288), .B(n13289), .Z(n13081) );
  XOR2_X1 U13263 ( .A(n13290), .B(n13291), .Z(n13289) );
  OR2_X1 U13264 ( .A1(n7985), .A2(n8041), .ZN(n13084) );
  OR2_X1 U13265 ( .A1(n13088), .A2(n13085), .ZN(n13259) );
  XOR2_X1 U13266 ( .A(n13292), .B(n13293), .Z(n13085) );
  XOR2_X1 U13267 ( .A(n13294), .B(n13295), .Z(n13293) );
  OR2_X1 U13268 ( .A1(n7985), .A2(n8037), .ZN(n13088) );
  OR2_X1 U13269 ( .A1(n13092), .A2(n13089), .ZN(n13256) );
  XOR2_X1 U13270 ( .A(n13296), .B(n13297), .Z(n13089) );
  XOR2_X1 U13271 ( .A(n13298), .B(n13299), .Z(n13297) );
  OR2_X1 U13272 ( .A1(n7985), .A2(n8034), .ZN(n13092) );
  OR2_X1 U13273 ( .A1(n13096), .A2(n13093), .ZN(n13253) );
  XOR2_X1 U13274 ( .A(n13300), .B(n13301), .Z(n13093) );
  XOR2_X1 U13275 ( .A(n13302), .B(n13303), .Z(n13301) );
  OR2_X1 U13276 ( .A1(n7985), .A2(n8030), .ZN(n13096) );
  OR2_X1 U13277 ( .A1(n13100), .A2(n13097), .ZN(n13250) );
  XOR2_X1 U13278 ( .A(n13304), .B(n13305), .Z(n13097) );
  XOR2_X1 U13279 ( .A(n13306), .B(n13307), .Z(n13305) );
  OR2_X1 U13280 ( .A1(n7985), .A2(n8026), .ZN(n13100) );
  OR2_X1 U13281 ( .A1(n13104), .A2(n13101), .ZN(n13247) );
  XOR2_X1 U13282 ( .A(n13308), .B(n13309), .Z(n13101) );
  XOR2_X1 U13283 ( .A(n13310), .B(n13311), .Z(n13309) );
  OR2_X1 U13284 ( .A1(n7985), .A2(n8023), .ZN(n13104) );
  XOR2_X1 U13285 ( .A(n13312), .B(n13313), .Z(n13105) );
  XOR2_X1 U13286 ( .A(n13314), .B(n13315), .Z(n13313) );
  OR2_X1 U13287 ( .A1(n13112), .A2(n13109), .ZN(n13241) );
  XOR2_X1 U13288 ( .A(n13316), .B(n13317), .Z(n13109) );
  XOR2_X1 U13289 ( .A(n13318), .B(n13319), .Z(n13317) );
  OR2_X1 U13290 ( .A1(n7985), .A2(n8016), .ZN(n13112) );
  INV_X1 U13291 ( .A(b_10_), .ZN(n7985) );
  XOR2_X1 U13292 ( .A(n13320), .B(n13321), .Z(n13113) );
  XOR2_X1 U13293 ( .A(n13322), .B(n13323), .Z(n13321) );
  XOR2_X1 U13294 ( .A(n13324), .B(n13325), .Z(n13117) );
  XOR2_X1 U13295 ( .A(n13326), .B(n13327), .Z(n13325) );
  XOR2_X1 U13296 ( .A(n13328), .B(n13329), .Z(n13121) );
  XOR2_X1 U13297 ( .A(n13330), .B(n13331), .Z(n13329) );
  XOR2_X1 U13298 ( .A(n13332), .B(n13333), .Z(n13125) );
  XOR2_X1 U13299 ( .A(n13334), .B(n13335), .Z(n13333) );
  XOR2_X1 U13300 ( .A(n13336), .B(n13337), .Z(n13129) );
  XOR2_X1 U13301 ( .A(n13338), .B(n13339), .Z(n13337) );
  XOR2_X1 U13302 ( .A(n13340), .B(n13341), .Z(n13133) );
  XOR2_X1 U13303 ( .A(n13342), .B(n13343), .Z(n13341) );
  XOR2_X1 U13304 ( .A(n13344), .B(n13345), .Z(n13137) );
  XOR2_X1 U13305 ( .A(n13346), .B(n13347), .Z(n13345) );
  XOR2_X1 U13306 ( .A(n13348), .B(n13349), .Z(n13141) );
  XOR2_X1 U13307 ( .A(n13350), .B(n13351), .Z(n13349) );
  INV_X1 U13308 ( .A(n7796), .ZN(n7986) );
  AND2_X1 U13309 ( .A1(b_10_), .A2(a_10_), .ZN(n7796) );
  XOR2_X1 U13310 ( .A(n13352), .B(n13353), .Z(n13146) );
  XOR2_X1 U13311 ( .A(n13354), .B(n13355), .Z(n13353) );
  XOR2_X1 U13312 ( .A(n13356), .B(n13357), .Z(n13148) );
  XOR2_X1 U13313 ( .A(n13358), .B(n13359), .Z(n13357) );
  XOR2_X1 U13314 ( .A(n13360), .B(n13361), .Z(n13152) );
  XNOR2_X1 U13315 ( .A(n13362), .B(n7808), .ZN(n13361) );
  XOR2_X1 U13316 ( .A(n13363), .B(n13364), .Z(n13156) );
  XOR2_X1 U13317 ( .A(n13365), .B(n13366), .Z(n13364) );
  XOR2_X1 U13318 ( .A(n13367), .B(n13368), .Z(n13160) );
  XOR2_X1 U13319 ( .A(n13369), .B(n13370), .Z(n13368) );
  XOR2_X1 U13320 ( .A(n13371), .B(n13372), .Z(n13164) );
  XOR2_X1 U13321 ( .A(n13373), .B(n13374), .Z(n13372) );
  XOR2_X1 U13322 ( .A(n13375), .B(n13376), .Z(n13168) );
  XOR2_X1 U13323 ( .A(n13377), .B(n13378), .Z(n13376) );
  XOR2_X1 U13324 ( .A(n13379), .B(n13380), .Z(n13172) );
  XOR2_X1 U13325 ( .A(n13381), .B(n13382), .Z(n13380) );
  XOR2_X1 U13326 ( .A(n13383), .B(n13384), .Z(n13176) );
  XOR2_X1 U13327 ( .A(n13385), .B(n13386), .Z(n13384) );
  XOR2_X1 U13328 ( .A(n13387), .B(n13388), .Z(n13180) );
  XOR2_X1 U13329 ( .A(n13389), .B(n13390), .Z(n13388) );
  XOR2_X1 U13330 ( .A(n8459), .B(n13391), .Z(n8452) );
  XOR2_X1 U13331 ( .A(n8458), .B(n8457), .Z(n13391) );
  OR2_X1 U13332 ( .A1(n7804), .A2(n7953), .ZN(n8457) );
  OR2_X1 U13333 ( .A1(n13392), .A2(n13393), .ZN(n8458) );
  AND2_X1 U13334 ( .A1(n13390), .A2(n13389), .ZN(n13393) );
  AND2_X1 U13335 ( .A1(n13387), .A2(n13394), .ZN(n13392) );
  OR2_X1 U13336 ( .A1(n13389), .A2(n13390), .ZN(n13394) );
  OR2_X1 U13337 ( .A1(n7804), .A2(n7956), .ZN(n13390) );
  OR2_X1 U13338 ( .A1(n13395), .A2(n13396), .ZN(n13389) );
  AND2_X1 U13339 ( .A1(n13386), .A2(n13385), .ZN(n13396) );
  AND2_X1 U13340 ( .A1(n13383), .A2(n13397), .ZN(n13395) );
  OR2_X1 U13341 ( .A1(n13385), .A2(n13386), .ZN(n13397) );
  OR2_X1 U13342 ( .A1(n7804), .A2(n7960), .ZN(n13386) );
  OR2_X1 U13343 ( .A1(n13398), .A2(n13399), .ZN(n13385) );
  AND2_X1 U13344 ( .A1(n13382), .A2(n13381), .ZN(n13399) );
  AND2_X1 U13345 ( .A1(n13379), .A2(n13400), .ZN(n13398) );
  OR2_X1 U13346 ( .A1(n13381), .A2(n13382), .ZN(n13400) );
  OR2_X1 U13347 ( .A1(n7804), .A2(n7963), .ZN(n13382) );
  OR2_X1 U13348 ( .A1(n13401), .A2(n13402), .ZN(n13381) );
  AND2_X1 U13349 ( .A1(n13378), .A2(n13377), .ZN(n13402) );
  AND2_X1 U13350 ( .A1(n13375), .A2(n13403), .ZN(n13401) );
  OR2_X1 U13351 ( .A1(n13377), .A2(n13378), .ZN(n13403) );
  OR2_X1 U13352 ( .A1(n7804), .A2(n7967), .ZN(n13378) );
  OR2_X1 U13353 ( .A1(n13404), .A2(n13405), .ZN(n13377) );
  AND2_X1 U13354 ( .A1(n13374), .A2(n13373), .ZN(n13405) );
  AND2_X1 U13355 ( .A1(n13371), .A2(n13406), .ZN(n13404) );
  OR2_X1 U13356 ( .A1(n13373), .A2(n13374), .ZN(n13406) );
  OR2_X1 U13357 ( .A1(n7804), .A2(n7970), .ZN(n13374) );
  OR2_X1 U13358 ( .A1(n13407), .A2(n13408), .ZN(n13373) );
  AND2_X1 U13359 ( .A1(n13370), .A2(n13369), .ZN(n13408) );
  AND2_X1 U13360 ( .A1(n13367), .A2(n13409), .ZN(n13407) );
  OR2_X1 U13361 ( .A1(n13369), .A2(n13370), .ZN(n13409) );
  OR2_X1 U13362 ( .A1(n7804), .A2(n7974), .ZN(n13370) );
  OR2_X1 U13363 ( .A1(n13410), .A2(n13411), .ZN(n13369) );
  AND2_X1 U13364 ( .A1(n13366), .A2(n13365), .ZN(n13411) );
  AND2_X1 U13365 ( .A1(n13363), .A2(n13412), .ZN(n13410) );
  OR2_X1 U13366 ( .A1(n13365), .A2(n13366), .ZN(n13412) );
  OR2_X1 U13367 ( .A1(n7804), .A2(n7977), .ZN(n13366) );
  OR2_X1 U13368 ( .A1(n13413), .A2(n13414), .ZN(n13365) );
  AND2_X1 U13369 ( .A1(n7982), .A2(n13362), .ZN(n13414) );
  AND2_X1 U13370 ( .A1(n13360), .A2(n13415), .ZN(n13413) );
  OR2_X1 U13371 ( .A1(n13362), .A2(n7982), .ZN(n13415) );
  INV_X1 U13372 ( .A(n7808), .ZN(n7982) );
  AND2_X1 U13373 ( .A1(b_9_), .A2(a_9_), .ZN(n7808) );
  OR2_X1 U13374 ( .A1(n13416), .A2(n13417), .ZN(n13362) );
  AND2_X1 U13375 ( .A1(n13359), .A2(n13358), .ZN(n13417) );
  AND2_X1 U13376 ( .A1(n13356), .A2(n13418), .ZN(n13416) );
  OR2_X1 U13377 ( .A1(n13358), .A2(n13359), .ZN(n13418) );
  OR2_X1 U13378 ( .A1(n7804), .A2(n7984), .ZN(n13359) );
  OR2_X1 U13379 ( .A1(n13419), .A2(n13420), .ZN(n13358) );
  AND2_X1 U13380 ( .A1(n13355), .A2(n13354), .ZN(n13420) );
  AND2_X1 U13381 ( .A1(n13352), .A2(n13421), .ZN(n13419) );
  OR2_X1 U13382 ( .A1(n13354), .A2(n13355), .ZN(n13421) );
  OR2_X1 U13383 ( .A1(n7804), .A2(n7988), .ZN(n13355) );
  OR2_X1 U13384 ( .A1(n13422), .A2(n13423), .ZN(n13354) );
  AND2_X1 U13385 ( .A1(n13351), .A2(n13350), .ZN(n13423) );
  AND2_X1 U13386 ( .A1(n13348), .A2(n13424), .ZN(n13422) );
  OR2_X1 U13387 ( .A1(n13350), .A2(n13351), .ZN(n13424) );
  OR2_X1 U13388 ( .A1(n7804), .A2(n7991), .ZN(n13351) );
  OR2_X1 U13389 ( .A1(n13425), .A2(n13426), .ZN(n13350) );
  AND2_X1 U13390 ( .A1(n13347), .A2(n13346), .ZN(n13426) );
  AND2_X1 U13391 ( .A1(n13344), .A2(n13427), .ZN(n13425) );
  OR2_X1 U13392 ( .A1(n13346), .A2(n13347), .ZN(n13427) );
  OR2_X1 U13393 ( .A1(n7804), .A2(n7995), .ZN(n13347) );
  OR2_X1 U13394 ( .A1(n13428), .A2(n13429), .ZN(n13346) );
  AND2_X1 U13395 ( .A1(n13343), .A2(n13342), .ZN(n13429) );
  AND2_X1 U13396 ( .A1(n13340), .A2(n13430), .ZN(n13428) );
  OR2_X1 U13397 ( .A1(n13342), .A2(n13343), .ZN(n13430) );
  OR2_X1 U13398 ( .A1(n7804), .A2(n7998), .ZN(n13343) );
  OR2_X1 U13399 ( .A1(n13431), .A2(n13432), .ZN(n13342) );
  AND2_X1 U13400 ( .A1(n13339), .A2(n13338), .ZN(n13432) );
  AND2_X1 U13401 ( .A1(n13336), .A2(n13433), .ZN(n13431) );
  OR2_X1 U13402 ( .A1(n13338), .A2(n13339), .ZN(n13433) );
  OR2_X1 U13403 ( .A1(n7804), .A2(n8002), .ZN(n13339) );
  OR2_X1 U13404 ( .A1(n13434), .A2(n13435), .ZN(n13338) );
  AND2_X1 U13405 ( .A1(n13335), .A2(n13334), .ZN(n13435) );
  AND2_X1 U13406 ( .A1(n13332), .A2(n13436), .ZN(n13434) );
  OR2_X1 U13407 ( .A1(n13334), .A2(n13335), .ZN(n13436) );
  OR2_X1 U13408 ( .A1(n7804), .A2(n8005), .ZN(n13335) );
  OR2_X1 U13409 ( .A1(n13437), .A2(n13438), .ZN(n13334) );
  AND2_X1 U13410 ( .A1(n13331), .A2(n13330), .ZN(n13438) );
  AND2_X1 U13411 ( .A1(n13328), .A2(n13439), .ZN(n13437) );
  OR2_X1 U13412 ( .A1(n13330), .A2(n13331), .ZN(n13439) );
  OR2_X1 U13413 ( .A1(n7804), .A2(n8009), .ZN(n13331) );
  OR2_X1 U13414 ( .A1(n13440), .A2(n13441), .ZN(n13330) );
  AND2_X1 U13415 ( .A1(n13327), .A2(n13326), .ZN(n13441) );
  AND2_X1 U13416 ( .A1(n13324), .A2(n13442), .ZN(n13440) );
  OR2_X1 U13417 ( .A1(n13326), .A2(n13327), .ZN(n13442) );
  OR2_X1 U13418 ( .A1(n7804), .A2(n8012), .ZN(n13327) );
  OR2_X1 U13419 ( .A1(n13443), .A2(n13444), .ZN(n13326) );
  AND2_X1 U13420 ( .A1(n13323), .A2(n13322), .ZN(n13444) );
  AND2_X1 U13421 ( .A1(n13320), .A2(n13445), .ZN(n13443) );
  OR2_X1 U13422 ( .A1(n13322), .A2(n13323), .ZN(n13445) );
  OR2_X1 U13423 ( .A1(n7804), .A2(n8016), .ZN(n13323) );
  OR2_X1 U13424 ( .A1(n13446), .A2(n13447), .ZN(n13322) );
  AND2_X1 U13425 ( .A1(n13316), .A2(n13319), .ZN(n13447) );
  AND2_X1 U13426 ( .A1(n13448), .A2(n13318), .ZN(n13446) );
  OR2_X1 U13427 ( .A1(n13449), .A2(n13450), .ZN(n13318) );
  AND2_X1 U13428 ( .A1(n13315), .A2(n13314), .ZN(n13450) );
  AND2_X1 U13429 ( .A1(n13312), .A2(n13451), .ZN(n13449) );
  OR2_X1 U13430 ( .A1(n13314), .A2(n13315), .ZN(n13451) );
  OR2_X1 U13431 ( .A1(n7804), .A2(n8023), .ZN(n13315) );
  OR2_X1 U13432 ( .A1(n13452), .A2(n13453), .ZN(n13314) );
  AND2_X1 U13433 ( .A1(n13308), .A2(n13311), .ZN(n13453) );
  AND2_X1 U13434 ( .A1(n13454), .A2(n13310), .ZN(n13452) );
  OR2_X1 U13435 ( .A1(n13455), .A2(n13456), .ZN(n13310) );
  AND2_X1 U13436 ( .A1(n13304), .A2(n13307), .ZN(n13456) );
  AND2_X1 U13437 ( .A1(n13457), .A2(n13306), .ZN(n13455) );
  OR2_X1 U13438 ( .A1(n13458), .A2(n13459), .ZN(n13306) );
  AND2_X1 U13439 ( .A1(n13300), .A2(n13303), .ZN(n13459) );
  AND2_X1 U13440 ( .A1(n13460), .A2(n13302), .ZN(n13458) );
  OR2_X1 U13441 ( .A1(n13461), .A2(n13462), .ZN(n13302) );
  AND2_X1 U13442 ( .A1(n13296), .A2(n13299), .ZN(n13462) );
  AND2_X1 U13443 ( .A1(n13463), .A2(n13298), .ZN(n13461) );
  OR2_X1 U13444 ( .A1(n13464), .A2(n13465), .ZN(n13298) );
  AND2_X1 U13445 ( .A1(n13292), .A2(n13295), .ZN(n13465) );
  AND2_X1 U13446 ( .A1(n13466), .A2(n13294), .ZN(n13464) );
  OR2_X1 U13447 ( .A1(n13467), .A2(n13468), .ZN(n13294) );
  AND2_X1 U13448 ( .A1(n13288), .A2(n13291), .ZN(n13468) );
  AND2_X1 U13449 ( .A1(n13469), .A2(n13290), .ZN(n13467) );
  OR2_X1 U13450 ( .A1(n13470), .A2(n13471), .ZN(n13290) );
  AND2_X1 U13451 ( .A1(n13284), .A2(n13287), .ZN(n13471) );
  AND2_X1 U13452 ( .A1(n13472), .A2(n13286), .ZN(n13470) );
  OR2_X1 U13453 ( .A1(n13473), .A2(n13474), .ZN(n13286) );
  AND2_X1 U13454 ( .A1(n13280), .A2(n13475), .ZN(n13474) );
  AND2_X1 U13455 ( .A1(n13476), .A2(n13477), .ZN(n13473) );
  OR2_X1 U13456 ( .A1(n13475), .A2(n13280), .ZN(n13477) );
  OR2_X1 U13457 ( .A1(n7804), .A2(n8051), .ZN(n13280) );
  INV_X1 U13458 ( .A(n13283), .ZN(n13475) );
  AND3_X1 U13459 ( .A1(b_9_), .A2(n8904), .A3(b_8_), .ZN(n13283) );
  INV_X1 U13460 ( .A(n13282), .ZN(n13476) );
  OR2_X1 U13461 ( .A1(n13478), .A2(n13479), .ZN(n13282) );
  AND2_X1 U13462 ( .A1(b_8_), .A2(n13480), .ZN(n13479) );
  OR2_X1 U13463 ( .A1(n13481), .A2(n7490), .ZN(n13480) );
  AND2_X1 U13464 ( .A1(a_30_), .A2(n7843), .ZN(n13481) );
  AND2_X1 U13465 ( .A1(b_7_), .A2(n13482), .ZN(n13478) );
  OR2_X1 U13466 ( .A1(n13483), .A2(n7493), .ZN(n13482) );
  AND2_X1 U13467 ( .A1(a_31_), .A2(n7978), .ZN(n13483) );
  OR2_X1 U13468 ( .A1(n13287), .A2(n13284), .ZN(n13472) );
  XNOR2_X1 U13469 ( .A(n13484), .B(n13485), .ZN(n13284) );
  XNOR2_X1 U13470 ( .A(n13486), .B(n13487), .ZN(n13485) );
  OR2_X1 U13471 ( .A1(n7804), .A2(n8048), .ZN(n13287) );
  OR2_X1 U13472 ( .A1(n13291), .A2(n13288), .ZN(n13469) );
  XOR2_X1 U13473 ( .A(n13488), .B(n13489), .Z(n13288) );
  XOR2_X1 U13474 ( .A(n13490), .B(n13491), .Z(n13489) );
  OR2_X1 U13475 ( .A1(n7804), .A2(n8044), .ZN(n13291) );
  OR2_X1 U13476 ( .A1(n13295), .A2(n13292), .ZN(n13466) );
  XOR2_X1 U13477 ( .A(n13492), .B(n13493), .Z(n13292) );
  XOR2_X1 U13478 ( .A(n13494), .B(n13495), .Z(n13493) );
  OR2_X1 U13479 ( .A1(n7804), .A2(n8041), .ZN(n13295) );
  OR2_X1 U13480 ( .A1(n13299), .A2(n13296), .ZN(n13463) );
  XOR2_X1 U13481 ( .A(n13496), .B(n13497), .Z(n13296) );
  XOR2_X1 U13482 ( .A(n13498), .B(n13499), .Z(n13497) );
  OR2_X1 U13483 ( .A1(n7804), .A2(n8037), .ZN(n13299) );
  OR2_X1 U13484 ( .A1(n13303), .A2(n13300), .ZN(n13460) );
  XOR2_X1 U13485 ( .A(n13500), .B(n13501), .Z(n13300) );
  XOR2_X1 U13486 ( .A(n13502), .B(n13503), .Z(n13501) );
  OR2_X1 U13487 ( .A1(n7804), .A2(n8034), .ZN(n13303) );
  OR2_X1 U13488 ( .A1(n13307), .A2(n13304), .ZN(n13457) );
  XOR2_X1 U13489 ( .A(n13504), .B(n13505), .Z(n13304) );
  XOR2_X1 U13490 ( .A(n13506), .B(n13507), .Z(n13505) );
  OR2_X1 U13491 ( .A1(n7804), .A2(n8030), .ZN(n13307) );
  OR2_X1 U13492 ( .A1(n13311), .A2(n13308), .ZN(n13454) );
  XOR2_X1 U13493 ( .A(n13508), .B(n13509), .Z(n13308) );
  XOR2_X1 U13494 ( .A(n13510), .B(n13511), .Z(n13509) );
  OR2_X1 U13495 ( .A1(n7804), .A2(n8026), .ZN(n13311) );
  XOR2_X1 U13496 ( .A(n13512), .B(n13513), .Z(n13312) );
  XOR2_X1 U13497 ( .A(n13514), .B(n13515), .Z(n13513) );
  OR2_X1 U13498 ( .A1(n13319), .A2(n13316), .ZN(n13448) );
  XOR2_X1 U13499 ( .A(n13516), .B(n13517), .Z(n13316) );
  XOR2_X1 U13500 ( .A(n13518), .B(n13519), .Z(n13517) );
  OR2_X1 U13501 ( .A1(n7804), .A2(n8019), .ZN(n13319) );
  INV_X1 U13502 ( .A(b_9_), .ZN(n7804) );
  XOR2_X1 U13503 ( .A(n13520), .B(n13521), .Z(n13320) );
  XOR2_X1 U13504 ( .A(n13522), .B(n13523), .Z(n13521) );
  XOR2_X1 U13505 ( .A(n13524), .B(n13525), .Z(n13324) );
  XOR2_X1 U13506 ( .A(n13526), .B(n13527), .Z(n13525) );
  XOR2_X1 U13507 ( .A(n13528), .B(n13529), .Z(n13328) );
  XOR2_X1 U13508 ( .A(n13530), .B(n13531), .Z(n13529) );
  XOR2_X1 U13509 ( .A(n13532), .B(n13533), .Z(n13332) );
  XOR2_X1 U13510 ( .A(n13534), .B(n13535), .Z(n13533) );
  XOR2_X1 U13511 ( .A(n13536), .B(n13537), .Z(n13336) );
  XOR2_X1 U13512 ( .A(n13538), .B(n13539), .Z(n13537) );
  XOR2_X1 U13513 ( .A(n13540), .B(n13541), .Z(n13340) );
  XOR2_X1 U13514 ( .A(n13542), .B(n13543), .Z(n13541) );
  XOR2_X1 U13515 ( .A(n13544), .B(n13545), .Z(n13344) );
  XOR2_X1 U13516 ( .A(n13546), .B(n13547), .Z(n13545) );
  XOR2_X1 U13517 ( .A(n13548), .B(n13549), .Z(n13348) );
  XOR2_X1 U13518 ( .A(n13550), .B(n13551), .Z(n13549) );
  XOR2_X1 U13519 ( .A(n13552), .B(n13553), .Z(n13352) );
  XOR2_X1 U13520 ( .A(n13554), .B(n13555), .Z(n13553) );
  XOR2_X1 U13521 ( .A(n13556), .B(n13557), .Z(n13356) );
  XOR2_X1 U13522 ( .A(n13558), .B(n13559), .Z(n13557) );
  XOR2_X1 U13523 ( .A(n13560), .B(n13561), .Z(n13360) );
  XOR2_X1 U13524 ( .A(n13562), .B(n13563), .Z(n13561) );
  XOR2_X1 U13525 ( .A(n13564), .B(n13565), .Z(n13363) );
  XOR2_X1 U13526 ( .A(n13566), .B(n13567), .Z(n13565) );
  XNOR2_X1 U13527 ( .A(n13568), .B(n13569), .ZN(n13367) );
  XNOR2_X1 U13528 ( .A(n7979), .B(n13570), .ZN(n13568) );
  XOR2_X1 U13529 ( .A(n13571), .B(n13572), .Z(n13371) );
  XOR2_X1 U13530 ( .A(n13573), .B(n13574), .Z(n13572) );
  XOR2_X1 U13531 ( .A(n13575), .B(n13576), .Z(n13375) );
  XOR2_X1 U13532 ( .A(n13577), .B(n13578), .Z(n13576) );
  XOR2_X1 U13533 ( .A(n13579), .B(n13580), .Z(n13379) );
  XOR2_X1 U13534 ( .A(n13581), .B(n13582), .Z(n13580) );
  XOR2_X1 U13535 ( .A(n13583), .B(n13584), .Z(n13383) );
  XOR2_X1 U13536 ( .A(n13585), .B(n13586), .Z(n13584) );
  XOR2_X1 U13537 ( .A(n13587), .B(n13588), .Z(n13387) );
  XOR2_X1 U13538 ( .A(n13589), .B(n13590), .Z(n13588) );
  XOR2_X1 U13539 ( .A(n8466), .B(n13591), .Z(n8459) );
  XOR2_X1 U13540 ( .A(n8465), .B(n8464), .Z(n13591) );
  OR2_X1 U13541 ( .A1(n7978), .A2(n7956), .ZN(n8464) );
  OR2_X1 U13542 ( .A1(n13592), .A2(n13593), .ZN(n8465) );
  AND2_X1 U13543 ( .A1(n13590), .A2(n13589), .ZN(n13593) );
  AND2_X1 U13544 ( .A1(n13587), .A2(n13594), .ZN(n13592) );
  OR2_X1 U13545 ( .A1(n13589), .A2(n13590), .ZN(n13594) );
  OR2_X1 U13546 ( .A1(n7978), .A2(n7960), .ZN(n13590) );
  OR2_X1 U13547 ( .A1(n13595), .A2(n13596), .ZN(n13589) );
  AND2_X1 U13548 ( .A1(n13586), .A2(n13585), .ZN(n13596) );
  AND2_X1 U13549 ( .A1(n13583), .A2(n13597), .ZN(n13595) );
  OR2_X1 U13550 ( .A1(n13585), .A2(n13586), .ZN(n13597) );
  OR2_X1 U13551 ( .A1(n7978), .A2(n7963), .ZN(n13586) );
  OR2_X1 U13552 ( .A1(n13598), .A2(n13599), .ZN(n13585) );
  AND2_X1 U13553 ( .A1(n13582), .A2(n13581), .ZN(n13599) );
  AND2_X1 U13554 ( .A1(n13579), .A2(n13600), .ZN(n13598) );
  OR2_X1 U13555 ( .A1(n13581), .A2(n13582), .ZN(n13600) );
  OR2_X1 U13556 ( .A1(n7978), .A2(n7967), .ZN(n13582) );
  OR2_X1 U13557 ( .A1(n13601), .A2(n13602), .ZN(n13581) );
  AND2_X1 U13558 ( .A1(n13578), .A2(n13577), .ZN(n13602) );
  AND2_X1 U13559 ( .A1(n13575), .A2(n13603), .ZN(n13601) );
  OR2_X1 U13560 ( .A1(n13577), .A2(n13578), .ZN(n13603) );
  OR2_X1 U13561 ( .A1(n7978), .A2(n7970), .ZN(n13578) );
  OR2_X1 U13562 ( .A1(n13604), .A2(n13605), .ZN(n13577) );
  AND2_X1 U13563 ( .A1(n13574), .A2(n13573), .ZN(n13605) );
  AND2_X1 U13564 ( .A1(n13571), .A2(n13606), .ZN(n13604) );
  OR2_X1 U13565 ( .A1(n13573), .A2(n13574), .ZN(n13606) );
  OR2_X1 U13566 ( .A1(n7978), .A2(n7974), .ZN(n13574) );
  OR2_X1 U13567 ( .A1(n13607), .A2(n13608), .ZN(n13573) );
  AND2_X1 U13568 ( .A1(n13570), .A2(n7979), .ZN(n13608) );
  AND2_X1 U13569 ( .A1(n13569), .A2(n13609), .ZN(n13607) );
  OR2_X1 U13570 ( .A1(n7979), .A2(n13570), .ZN(n13609) );
  OR2_X1 U13571 ( .A1(n13610), .A2(n13611), .ZN(n13570) );
  AND2_X1 U13572 ( .A1(n13567), .A2(n13566), .ZN(n13611) );
  AND2_X1 U13573 ( .A1(n13564), .A2(n13612), .ZN(n13610) );
  OR2_X1 U13574 ( .A1(n13566), .A2(n13567), .ZN(n13612) );
  OR2_X1 U13575 ( .A1(n7978), .A2(n7981), .ZN(n13567) );
  OR2_X1 U13576 ( .A1(n13613), .A2(n13614), .ZN(n13566) );
  AND2_X1 U13577 ( .A1(n13563), .A2(n13562), .ZN(n13614) );
  AND2_X1 U13578 ( .A1(n13560), .A2(n13615), .ZN(n13613) );
  OR2_X1 U13579 ( .A1(n13562), .A2(n13563), .ZN(n13615) );
  OR2_X1 U13580 ( .A1(n7978), .A2(n7984), .ZN(n13563) );
  OR2_X1 U13581 ( .A1(n13616), .A2(n13617), .ZN(n13562) );
  AND2_X1 U13582 ( .A1(n13559), .A2(n13558), .ZN(n13617) );
  AND2_X1 U13583 ( .A1(n13556), .A2(n13618), .ZN(n13616) );
  OR2_X1 U13584 ( .A1(n13558), .A2(n13559), .ZN(n13618) );
  OR2_X1 U13585 ( .A1(n7978), .A2(n7988), .ZN(n13559) );
  OR2_X1 U13586 ( .A1(n13619), .A2(n13620), .ZN(n13558) );
  AND2_X1 U13587 ( .A1(n13555), .A2(n13554), .ZN(n13620) );
  AND2_X1 U13588 ( .A1(n13552), .A2(n13621), .ZN(n13619) );
  OR2_X1 U13589 ( .A1(n13554), .A2(n13555), .ZN(n13621) );
  OR2_X1 U13590 ( .A1(n7978), .A2(n7991), .ZN(n13555) );
  OR2_X1 U13591 ( .A1(n13622), .A2(n13623), .ZN(n13554) );
  AND2_X1 U13592 ( .A1(n13551), .A2(n13550), .ZN(n13623) );
  AND2_X1 U13593 ( .A1(n13548), .A2(n13624), .ZN(n13622) );
  OR2_X1 U13594 ( .A1(n13550), .A2(n13551), .ZN(n13624) );
  OR2_X1 U13595 ( .A1(n7978), .A2(n7995), .ZN(n13551) );
  OR2_X1 U13596 ( .A1(n13625), .A2(n13626), .ZN(n13550) );
  AND2_X1 U13597 ( .A1(n13547), .A2(n13546), .ZN(n13626) );
  AND2_X1 U13598 ( .A1(n13544), .A2(n13627), .ZN(n13625) );
  OR2_X1 U13599 ( .A1(n13546), .A2(n13547), .ZN(n13627) );
  OR2_X1 U13600 ( .A1(n7978), .A2(n7998), .ZN(n13547) );
  OR2_X1 U13601 ( .A1(n13628), .A2(n13629), .ZN(n13546) );
  AND2_X1 U13602 ( .A1(n13543), .A2(n13542), .ZN(n13629) );
  AND2_X1 U13603 ( .A1(n13540), .A2(n13630), .ZN(n13628) );
  OR2_X1 U13604 ( .A1(n13542), .A2(n13543), .ZN(n13630) );
  OR2_X1 U13605 ( .A1(n7978), .A2(n8002), .ZN(n13543) );
  OR2_X1 U13606 ( .A1(n13631), .A2(n13632), .ZN(n13542) );
  AND2_X1 U13607 ( .A1(n13539), .A2(n13538), .ZN(n13632) );
  AND2_X1 U13608 ( .A1(n13536), .A2(n13633), .ZN(n13631) );
  OR2_X1 U13609 ( .A1(n13538), .A2(n13539), .ZN(n13633) );
  OR2_X1 U13610 ( .A1(n7978), .A2(n8005), .ZN(n13539) );
  OR2_X1 U13611 ( .A1(n13634), .A2(n13635), .ZN(n13538) );
  AND2_X1 U13612 ( .A1(n13535), .A2(n13534), .ZN(n13635) );
  AND2_X1 U13613 ( .A1(n13532), .A2(n13636), .ZN(n13634) );
  OR2_X1 U13614 ( .A1(n13534), .A2(n13535), .ZN(n13636) );
  OR2_X1 U13615 ( .A1(n7978), .A2(n8009), .ZN(n13535) );
  OR2_X1 U13616 ( .A1(n13637), .A2(n13638), .ZN(n13534) );
  AND2_X1 U13617 ( .A1(n13531), .A2(n13530), .ZN(n13638) );
  AND2_X1 U13618 ( .A1(n13528), .A2(n13639), .ZN(n13637) );
  OR2_X1 U13619 ( .A1(n13530), .A2(n13531), .ZN(n13639) );
  OR2_X1 U13620 ( .A1(n7978), .A2(n8012), .ZN(n13531) );
  OR2_X1 U13621 ( .A1(n13640), .A2(n13641), .ZN(n13530) );
  AND2_X1 U13622 ( .A1(n13527), .A2(n13526), .ZN(n13641) );
  AND2_X1 U13623 ( .A1(n13524), .A2(n13642), .ZN(n13640) );
  OR2_X1 U13624 ( .A1(n13526), .A2(n13527), .ZN(n13642) );
  OR2_X1 U13625 ( .A1(n7978), .A2(n8016), .ZN(n13527) );
  OR2_X1 U13626 ( .A1(n13643), .A2(n13644), .ZN(n13526) );
  AND2_X1 U13627 ( .A1(n13523), .A2(n13522), .ZN(n13644) );
  AND2_X1 U13628 ( .A1(n13520), .A2(n13645), .ZN(n13643) );
  OR2_X1 U13629 ( .A1(n13522), .A2(n13523), .ZN(n13645) );
  OR2_X1 U13630 ( .A1(n7978), .A2(n8019), .ZN(n13523) );
  OR2_X1 U13631 ( .A1(n13646), .A2(n13647), .ZN(n13522) );
  AND2_X1 U13632 ( .A1(n13516), .A2(n13519), .ZN(n13647) );
  AND2_X1 U13633 ( .A1(n13648), .A2(n13518), .ZN(n13646) );
  OR2_X1 U13634 ( .A1(n13649), .A2(n13650), .ZN(n13518) );
  AND2_X1 U13635 ( .A1(n13515), .A2(n13514), .ZN(n13650) );
  AND2_X1 U13636 ( .A1(n13512), .A2(n13651), .ZN(n13649) );
  OR2_X1 U13637 ( .A1(n13514), .A2(n13515), .ZN(n13651) );
  OR2_X1 U13638 ( .A1(n7978), .A2(n8026), .ZN(n13515) );
  OR2_X1 U13639 ( .A1(n13652), .A2(n13653), .ZN(n13514) );
  AND2_X1 U13640 ( .A1(n13508), .A2(n13511), .ZN(n13653) );
  AND2_X1 U13641 ( .A1(n13654), .A2(n13510), .ZN(n13652) );
  OR2_X1 U13642 ( .A1(n13655), .A2(n13656), .ZN(n13510) );
  AND2_X1 U13643 ( .A1(n13504), .A2(n13507), .ZN(n13656) );
  AND2_X1 U13644 ( .A1(n13657), .A2(n13506), .ZN(n13655) );
  OR2_X1 U13645 ( .A1(n13658), .A2(n13659), .ZN(n13506) );
  AND2_X1 U13646 ( .A1(n13500), .A2(n13503), .ZN(n13659) );
  AND2_X1 U13647 ( .A1(n13660), .A2(n13502), .ZN(n13658) );
  OR2_X1 U13648 ( .A1(n13661), .A2(n13662), .ZN(n13502) );
  AND2_X1 U13649 ( .A1(n13496), .A2(n13499), .ZN(n13662) );
  AND2_X1 U13650 ( .A1(n13663), .A2(n13498), .ZN(n13661) );
  OR2_X1 U13651 ( .A1(n13664), .A2(n13665), .ZN(n13498) );
  AND2_X1 U13652 ( .A1(n13492), .A2(n13495), .ZN(n13665) );
  AND2_X1 U13653 ( .A1(n13666), .A2(n13494), .ZN(n13664) );
  OR2_X1 U13654 ( .A1(n13667), .A2(n13668), .ZN(n13494) );
  AND2_X1 U13655 ( .A1(n13488), .A2(n13491), .ZN(n13668) );
  AND2_X1 U13656 ( .A1(n13669), .A2(n13490), .ZN(n13667) );
  OR2_X1 U13657 ( .A1(n13670), .A2(n13671), .ZN(n13490) );
  AND2_X1 U13658 ( .A1(n13484), .A2(n13672), .ZN(n13671) );
  AND2_X1 U13659 ( .A1(n13673), .A2(n13674), .ZN(n13670) );
  OR2_X1 U13660 ( .A1(n13672), .A2(n13484), .ZN(n13674) );
  OR2_X1 U13661 ( .A1(n8051), .A2(n7978), .ZN(n13484) );
  INV_X1 U13662 ( .A(n13487), .ZN(n13672) );
  AND3_X1 U13663 ( .A1(n8904), .A2(b_8_), .A3(b_7_), .ZN(n13487) );
  INV_X1 U13664 ( .A(n13486), .ZN(n13673) );
  OR2_X1 U13665 ( .A1(n13675), .A2(n13676), .ZN(n13486) );
  AND2_X1 U13666 ( .A1(b_7_), .A2(n13677), .ZN(n13676) );
  OR2_X1 U13667 ( .A1(n13678), .A2(n7490), .ZN(n13677) );
  AND2_X1 U13668 ( .A1(a_30_), .A2(n7971), .ZN(n13678) );
  AND2_X1 U13669 ( .A1(b_6_), .A2(n13679), .ZN(n13675) );
  OR2_X1 U13670 ( .A1(n13680), .A2(n7493), .ZN(n13679) );
  AND2_X1 U13671 ( .A1(a_31_), .A2(n7843), .ZN(n13680) );
  OR2_X1 U13672 ( .A1(n13491), .A2(n13488), .ZN(n13669) );
  XNOR2_X1 U13673 ( .A(n13681), .B(n13682), .ZN(n13488) );
  XNOR2_X1 U13674 ( .A(n13683), .B(n13684), .ZN(n13682) );
  OR2_X1 U13675 ( .A1(n8048), .A2(n7978), .ZN(n13491) );
  OR2_X1 U13676 ( .A1(n13495), .A2(n13492), .ZN(n13666) );
  XOR2_X1 U13677 ( .A(n13685), .B(n13686), .Z(n13492) );
  XOR2_X1 U13678 ( .A(n13687), .B(n13688), .Z(n13686) );
  OR2_X1 U13679 ( .A1(n7978), .A2(n8044), .ZN(n13495) );
  OR2_X1 U13680 ( .A1(n13499), .A2(n13496), .ZN(n13663) );
  XOR2_X1 U13681 ( .A(n13689), .B(n13690), .Z(n13496) );
  XOR2_X1 U13682 ( .A(n13691), .B(n13692), .Z(n13690) );
  OR2_X1 U13683 ( .A1(n7978), .A2(n8041), .ZN(n13499) );
  OR2_X1 U13684 ( .A1(n13503), .A2(n13500), .ZN(n13660) );
  XOR2_X1 U13685 ( .A(n13693), .B(n13694), .Z(n13500) );
  XOR2_X1 U13686 ( .A(n13695), .B(n13696), .Z(n13694) );
  OR2_X1 U13687 ( .A1(n7978), .A2(n8037), .ZN(n13503) );
  OR2_X1 U13688 ( .A1(n13507), .A2(n13504), .ZN(n13657) );
  XOR2_X1 U13689 ( .A(n13697), .B(n13698), .Z(n13504) );
  XOR2_X1 U13690 ( .A(n13699), .B(n13700), .Z(n13698) );
  OR2_X1 U13691 ( .A1(n7978), .A2(n8034), .ZN(n13507) );
  OR2_X1 U13692 ( .A1(n13511), .A2(n13508), .ZN(n13654) );
  XOR2_X1 U13693 ( .A(n13701), .B(n13702), .Z(n13508) );
  XOR2_X1 U13694 ( .A(n13703), .B(n13704), .Z(n13702) );
  OR2_X1 U13695 ( .A1(n7978), .A2(n8030), .ZN(n13511) );
  XOR2_X1 U13696 ( .A(n13705), .B(n13706), .Z(n13512) );
  XOR2_X1 U13697 ( .A(n13707), .B(n13708), .Z(n13706) );
  OR2_X1 U13698 ( .A1(n13519), .A2(n13516), .ZN(n13648) );
  XOR2_X1 U13699 ( .A(n13709), .B(n13710), .Z(n13516) );
  XOR2_X1 U13700 ( .A(n13711), .B(n13712), .Z(n13710) );
  OR2_X1 U13701 ( .A1(n7978), .A2(n8023), .ZN(n13519) );
  INV_X1 U13702 ( .A(b_8_), .ZN(n7978) );
  XOR2_X1 U13703 ( .A(n13713), .B(n13714), .Z(n13520) );
  XOR2_X1 U13704 ( .A(n13715), .B(n13716), .Z(n13714) );
  XOR2_X1 U13705 ( .A(n13717), .B(n13718), .Z(n13524) );
  XOR2_X1 U13706 ( .A(n13719), .B(n13720), .Z(n13718) );
  XOR2_X1 U13707 ( .A(n13721), .B(n13722), .Z(n13528) );
  XOR2_X1 U13708 ( .A(n13723), .B(n13724), .Z(n13722) );
  XOR2_X1 U13709 ( .A(n13725), .B(n13726), .Z(n13532) );
  XOR2_X1 U13710 ( .A(n13727), .B(n13728), .Z(n13726) );
  XOR2_X1 U13711 ( .A(n13729), .B(n13730), .Z(n13536) );
  XOR2_X1 U13712 ( .A(n13731), .B(n13732), .Z(n13730) );
  XOR2_X1 U13713 ( .A(n13733), .B(n13734), .Z(n13540) );
  XOR2_X1 U13714 ( .A(n13735), .B(n13736), .Z(n13734) );
  XOR2_X1 U13715 ( .A(n13737), .B(n13738), .Z(n13544) );
  XOR2_X1 U13716 ( .A(n13739), .B(n13740), .Z(n13738) );
  XOR2_X1 U13717 ( .A(n13741), .B(n13742), .Z(n13548) );
  XOR2_X1 U13718 ( .A(n13743), .B(n13744), .Z(n13742) );
  XOR2_X1 U13719 ( .A(n13745), .B(n13746), .Z(n13552) );
  XOR2_X1 U13720 ( .A(n13747), .B(n13748), .Z(n13746) );
  XOR2_X1 U13721 ( .A(n13749), .B(n13750), .Z(n13556) );
  XOR2_X1 U13722 ( .A(n13751), .B(n13752), .Z(n13750) );
  XOR2_X1 U13723 ( .A(n13753), .B(n13754), .Z(n13560) );
  XOR2_X1 U13724 ( .A(n13755), .B(n13756), .Z(n13754) );
  XOR2_X1 U13725 ( .A(n13757), .B(n13758), .Z(n13564) );
  XOR2_X1 U13726 ( .A(n13759), .B(n13760), .Z(n13758) );
  INV_X1 U13727 ( .A(n7825), .ZN(n7979) );
  AND2_X1 U13728 ( .A1(b_8_), .A2(a_8_), .ZN(n7825) );
  XOR2_X1 U13729 ( .A(n13761), .B(n13762), .Z(n13569) );
  XOR2_X1 U13730 ( .A(n13763), .B(n13764), .Z(n13762) );
  XOR2_X1 U13731 ( .A(n13765), .B(n13766), .Z(n13571) );
  XOR2_X1 U13732 ( .A(n13767), .B(n13768), .Z(n13766) );
  XOR2_X1 U13733 ( .A(n13769), .B(n13770), .Z(n13575) );
  XNOR2_X1 U13734 ( .A(n13771), .B(n7847), .ZN(n13770) );
  XOR2_X1 U13735 ( .A(n13772), .B(n13773), .Z(n13579) );
  XOR2_X1 U13736 ( .A(n13774), .B(n13775), .Z(n13773) );
  XOR2_X1 U13737 ( .A(n13776), .B(n13777), .Z(n13583) );
  XOR2_X1 U13738 ( .A(n13778), .B(n13779), .Z(n13777) );
  XOR2_X1 U13739 ( .A(n13780), .B(n13781), .Z(n13587) );
  XOR2_X1 U13740 ( .A(n13782), .B(n13783), .Z(n13781) );
  XOR2_X1 U13741 ( .A(n8473), .B(n13784), .Z(n8466) );
  XOR2_X1 U13742 ( .A(n8472), .B(n8471), .Z(n13784) );
  OR2_X1 U13743 ( .A1(n7843), .A2(n7960), .ZN(n8471) );
  OR2_X1 U13744 ( .A1(n13785), .A2(n13786), .ZN(n8472) );
  AND2_X1 U13745 ( .A1(n13783), .A2(n13782), .ZN(n13786) );
  AND2_X1 U13746 ( .A1(n13780), .A2(n13787), .ZN(n13785) );
  OR2_X1 U13747 ( .A1(n13782), .A2(n13783), .ZN(n13787) );
  OR2_X1 U13748 ( .A1(n7843), .A2(n7963), .ZN(n13783) );
  OR2_X1 U13749 ( .A1(n13788), .A2(n13789), .ZN(n13782) );
  AND2_X1 U13750 ( .A1(n13779), .A2(n13778), .ZN(n13789) );
  AND2_X1 U13751 ( .A1(n13776), .A2(n13790), .ZN(n13788) );
  OR2_X1 U13752 ( .A1(n13778), .A2(n13779), .ZN(n13790) );
  OR2_X1 U13753 ( .A1(n7843), .A2(n7967), .ZN(n13779) );
  OR2_X1 U13754 ( .A1(n13791), .A2(n13792), .ZN(n13778) );
  AND2_X1 U13755 ( .A1(n13775), .A2(n13774), .ZN(n13792) );
  AND2_X1 U13756 ( .A1(n13772), .A2(n13793), .ZN(n13791) );
  OR2_X1 U13757 ( .A1(n13774), .A2(n13775), .ZN(n13793) );
  OR2_X1 U13758 ( .A1(n7843), .A2(n7970), .ZN(n13775) );
  OR2_X1 U13759 ( .A1(n13794), .A2(n13795), .ZN(n13774) );
  AND2_X1 U13760 ( .A1(n7975), .A2(n13771), .ZN(n13795) );
  AND2_X1 U13761 ( .A1(n13769), .A2(n13796), .ZN(n13794) );
  OR2_X1 U13762 ( .A1(n13771), .A2(n7975), .ZN(n13796) );
  INV_X1 U13763 ( .A(n7847), .ZN(n7975) );
  AND2_X1 U13764 ( .A1(b_7_), .A2(a_7_), .ZN(n7847) );
  OR2_X1 U13765 ( .A1(n13797), .A2(n13798), .ZN(n13771) );
  AND2_X1 U13766 ( .A1(n13768), .A2(n13767), .ZN(n13798) );
  AND2_X1 U13767 ( .A1(n13765), .A2(n13799), .ZN(n13797) );
  OR2_X1 U13768 ( .A1(n13767), .A2(n13768), .ZN(n13799) );
  OR2_X1 U13769 ( .A1(n7843), .A2(n7977), .ZN(n13768) );
  OR2_X1 U13770 ( .A1(n13800), .A2(n13801), .ZN(n13767) );
  AND2_X1 U13771 ( .A1(n13764), .A2(n13763), .ZN(n13801) );
  AND2_X1 U13772 ( .A1(n13761), .A2(n13802), .ZN(n13800) );
  OR2_X1 U13773 ( .A1(n13763), .A2(n13764), .ZN(n13802) );
  OR2_X1 U13774 ( .A1(n7843), .A2(n7981), .ZN(n13764) );
  OR2_X1 U13775 ( .A1(n13803), .A2(n13804), .ZN(n13763) );
  AND2_X1 U13776 ( .A1(n13760), .A2(n13759), .ZN(n13804) );
  AND2_X1 U13777 ( .A1(n13757), .A2(n13805), .ZN(n13803) );
  OR2_X1 U13778 ( .A1(n13759), .A2(n13760), .ZN(n13805) );
  OR2_X1 U13779 ( .A1(n7843), .A2(n7984), .ZN(n13760) );
  OR2_X1 U13780 ( .A1(n13806), .A2(n13807), .ZN(n13759) );
  AND2_X1 U13781 ( .A1(n13756), .A2(n13755), .ZN(n13807) );
  AND2_X1 U13782 ( .A1(n13753), .A2(n13808), .ZN(n13806) );
  OR2_X1 U13783 ( .A1(n13755), .A2(n13756), .ZN(n13808) );
  OR2_X1 U13784 ( .A1(n7843), .A2(n7988), .ZN(n13756) );
  OR2_X1 U13785 ( .A1(n13809), .A2(n13810), .ZN(n13755) );
  AND2_X1 U13786 ( .A1(n13752), .A2(n13751), .ZN(n13810) );
  AND2_X1 U13787 ( .A1(n13749), .A2(n13811), .ZN(n13809) );
  OR2_X1 U13788 ( .A1(n13751), .A2(n13752), .ZN(n13811) );
  OR2_X1 U13789 ( .A1(n7843), .A2(n7991), .ZN(n13752) );
  OR2_X1 U13790 ( .A1(n13812), .A2(n13813), .ZN(n13751) );
  AND2_X1 U13791 ( .A1(n13748), .A2(n13747), .ZN(n13813) );
  AND2_X1 U13792 ( .A1(n13745), .A2(n13814), .ZN(n13812) );
  OR2_X1 U13793 ( .A1(n13747), .A2(n13748), .ZN(n13814) );
  OR2_X1 U13794 ( .A1(n7843), .A2(n7995), .ZN(n13748) );
  OR2_X1 U13795 ( .A1(n13815), .A2(n13816), .ZN(n13747) );
  AND2_X1 U13796 ( .A1(n13744), .A2(n13743), .ZN(n13816) );
  AND2_X1 U13797 ( .A1(n13741), .A2(n13817), .ZN(n13815) );
  OR2_X1 U13798 ( .A1(n13743), .A2(n13744), .ZN(n13817) );
  OR2_X1 U13799 ( .A1(n7843), .A2(n7998), .ZN(n13744) );
  OR2_X1 U13800 ( .A1(n13818), .A2(n13819), .ZN(n13743) );
  AND2_X1 U13801 ( .A1(n13740), .A2(n13739), .ZN(n13819) );
  AND2_X1 U13802 ( .A1(n13737), .A2(n13820), .ZN(n13818) );
  OR2_X1 U13803 ( .A1(n13739), .A2(n13740), .ZN(n13820) );
  OR2_X1 U13804 ( .A1(n7843), .A2(n8002), .ZN(n13740) );
  OR2_X1 U13805 ( .A1(n13821), .A2(n13822), .ZN(n13739) );
  AND2_X1 U13806 ( .A1(n13736), .A2(n13735), .ZN(n13822) );
  AND2_X1 U13807 ( .A1(n13733), .A2(n13823), .ZN(n13821) );
  OR2_X1 U13808 ( .A1(n13735), .A2(n13736), .ZN(n13823) );
  OR2_X1 U13809 ( .A1(n7843), .A2(n8005), .ZN(n13736) );
  OR2_X1 U13810 ( .A1(n13824), .A2(n13825), .ZN(n13735) );
  AND2_X1 U13811 ( .A1(n13732), .A2(n13731), .ZN(n13825) );
  AND2_X1 U13812 ( .A1(n13729), .A2(n13826), .ZN(n13824) );
  OR2_X1 U13813 ( .A1(n13731), .A2(n13732), .ZN(n13826) );
  OR2_X1 U13814 ( .A1(n7843), .A2(n8009), .ZN(n13732) );
  OR2_X1 U13815 ( .A1(n13827), .A2(n13828), .ZN(n13731) );
  AND2_X1 U13816 ( .A1(n13728), .A2(n13727), .ZN(n13828) );
  AND2_X1 U13817 ( .A1(n13725), .A2(n13829), .ZN(n13827) );
  OR2_X1 U13818 ( .A1(n13727), .A2(n13728), .ZN(n13829) );
  OR2_X1 U13819 ( .A1(n7843), .A2(n8012), .ZN(n13728) );
  OR2_X1 U13820 ( .A1(n13830), .A2(n13831), .ZN(n13727) );
  AND2_X1 U13821 ( .A1(n13724), .A2(n13723), .ZN(n13831) );
  AND2_X1 U13822 ( .A1(n13721), .A2(n13832), .ZN(n13830) );
  OR2_X1 U13823 ( .A1(n13723), .A2(n13724), .ZN(n13832) );
  OR2_X1 U13824 ( .A1(n7843), .A2(n8016), .ZN(n13724) );
  OR2_X1 U13825 ( .A1(n13833), .A2(n13834), .ZN(n13723) );
  AND2_X1 U13826 ( .A1(n13720), .A2(n13719), .ZN(n13834) );
  AND2_X1 U13827 ( .A1(n13717), .A2(n13835), .ZN(n13833) );
  OR2_X1 U13828 ( .A1(n13719), .A2(n13720), .ZN(n13835) );
  OR2_X1 U13829 ( .A1(n7843), .A2(n8019), .ZN(n13720) );
  OR2_X1 U13830 ( .A1(n13836), .A2(n13837), .ZN(n13719) );
  AND2_X1 U13831 ( .A1(n13716), .A2(n13715), .ZN(n13837) );
  AND2_X1 U13832 ( .A1(n13713), .A2(n13838), .ZN(n13836) );
  OR2_X1 U13833 ( .A1(n13715), .A2(n13716), .ZN(n13838) );
  OR2_X1 U13834 ( .A1(n7843), .A2(n8023), .ZN(n13716) );
  OR2_X1 U13835 ( .A1(n13839), .A2(n13840), .ZN(n13715) );
  AND2_X1 U13836 ( .A1(n13709), .A2(n13712), .ZN(n13840) );
  AND2_X1 U13837 ( .A1(n13841), .A2(n13711), .ZN(n13839) );
  OR2_X1 U13838 ( .A1(n13842), .A2(n13843), .ZN(n13711) );
  AND2_X1 U13839 ( .A1(n13708), .A2(n13707), .ZN(n13843) );
  AND2_X1 U13840 ( .A1(n13705), .A2(n13844), .ZN(n13842) );
  OR2_X1 U13841 ( .A1(n13707), .A2(n13708), .ZN(n13844) );
  OR2_X1 U13842 ( .A1(n7843), .A2(n8030), .ZN(n13708) );
  OR2_X1 U13843 ( .A1(n13845), .A2(n13846), .ZN(n13707) );
  AND2_X1 U13844 ( .A1(n13701), .A2(n13704), .ZN(n13846) );
  AND2_X1 U13845 ( .A1(n13847), .A2(n13703), .ZN(n13845) );
  OR2_X1 U13846 ( .A1(n13848), .A2(n13849), .ZN(n13703) );
  AND2_X1 U13847 ( .A1(n13697), .A2(n13700), .ZN(n13849) );
  AND2_X1 U13848 ( .A1(n13850), .A2(n13699), .ZN(n13848) );
  OR2_X1 U13849 ( .A1(n13851), .A2(n13852), .ZN(n13699) );
  AND2_X1 U13850 ( .A1(n13693), .A2(n13696), .ZN(n13852) );
  AND2_X1 U13851 ( .A1(n13853), .A2(n13695), .ZN(n13851) );
  OR2_X1 U13852 ( .A1(n13854), .A2(n13855), .ZN(n13695) );
  AND2_X1 U13853 ( .A1(n13689), .A2(n13692), .ZN(n13855) );
  AND2_X1 U13854 ( .A1(n13856), .A2(n13691), .ZN(n13854) );
  OR2_X1 U13855 ( .A1(n13857), .A2(n13858), .ZN(n13691) );
  AND2_X1 U13856 ( .A1(n13685), .A2(n13688), .ZN(n13858) );
  AND2_X1 U13857 ( .A1(n13859), .A2(n13687), .ZN(n13857) );
  OR2_X1 U13858 ( .A1(n13860), .A2(n13861), .ZN(n13687) );
  AND2_X1 U13859 ( .A1(n13681), .A2(n13862), .ZN(n13861) );
  AND2_X1 U13860 ( .A1(n13863), .A2(n13864), .ZN(n13860) );
  OR2_X1 U13861 ( .A1(n13862), .A2(n13681), .ZN(n13864) );
  OR2_X1 U13862 ( .A1(n8051), .A2(n7843), .ZN(n13681) );
  INV_X1 U13863 ( .A(n13684), .ZN(n13862) );
  AND3_X1 U13864 ( .A1(n8904), .A2(b_7_), .A3(b_6_), .ZN(n13684) );
  INV_X1 U13865 ( .A(n13683), .ZN(n13863) );
  OR2_X1 U13866 ( .A1(n13865), .A2(n13866), .ZN(n13683) );
  AND2_X1 U13867 ( .A1(b_6_), .A2(n13867), .ZN(n13866) );
  OR2_X1 U13868 ( .A1(n13868), .A2(n7490), .ZN(n13867) );
  AND2_X1 U13869 ( .A1(a_30_), .A2(n7872), .ZN(n13868) );
  AND2_X1 U13870 ( .A1(b_5_), .A2(n13869), .ZN(n13865) );
  OR2_X1 U13871 ( .A1(n13870), .A2(n7493), .ZN(n13869) );
  AND2_X1 U13872 ( .A1(a_31_), .A2(n7971), .ZN(n13870) );
  OR2_X1 U13873 ( .A1(n13688), .A2(n13685), .ZN(n13859) );
  XNOR2_X1 U13874 ( .A(n13871), .B(n13872), .ZN(n13685) );
  XNOR2_X1 U13875 ( .A(n13873), .B(n13874), .ZN(n13872) );
  OR2_X1 U13876 ( .A1(n8048), .A2(n7843), .ZN(n13688) );
  OR2_X1 U13877 ( .A1(n13692), .A2(n13689), .ZN(n13856) );
  XOR2_X1 U13878 ( .A(n13875), .B(n13876), .Z(n13689) );
  XOR2_X1 U13879 ( .A(n13877), .B(n13878), .Z(n13876) );
  OR2_X1 U13880 ( .A1(n8044), .A2(n7843), .ZN(n13692) );
  OR2_X1 U13881 ( .A1(n13696), .A2(n13693), .ZN(n13853) );
  XOR2_X1 U13882 ( .A(n13879), .B(n13880), .Z(n13693) );
  XOR2_X1 U13883 ( .A(n13881), .B(n13882), .Z(n13880) );
  OR2_X1 U13884 ( .A1(n7843), .A2(n8041), .ZN(n13696) );
  OR2_X1 U13885 ( .A1(n13700), .A2(n13697), .ZN(n13850) );
  XOR2_X1 U13886 ( .A(n13883), .B(n13884), .Z(n13697) );
  XOR2_X1 U13887 ( .A(n13885), .B(n13886), .Z(n13884) );
  OR2_X1 U13888 ( .A1(n7843), .A2(n8037), .ZN(n13700) );
  OR2_X1 U13889 ( .A1(n13704), .A2(n13701), .ZN(n13847) );
  XOR2_X1 U13890 ( .A(n13887), .B(n13888), .Z(n13701) );
  XOR2_X1 U13891 ( .A(n13889), .B(n13890), .Z(n13888) );
  OR2_X1 U13892 ( .A1(n7843), .A2(n8034), .ZN(n13704) );
  XOR2_X1 U13893 ( .A(n13891), .B(n13892), .Z(n13705) );
  XOR2_X1 U13894 ( .A(n13893), .B(n13894), .Z(n13892) );
  OR2_X1 U13895 ( .A1(n13712), .A2(n13709), .ZN(n13841) );
  XOR2_X1 U13896 ( .A(n13895), .B(n13896), .Z(n13709) );
  XOR2_X1 U13897 ( .A(n13897), .B(n13898), .Z(n13896) );
  OR2_X1 U13898 ( .A1(n7843), .A2(n8026), .ZN(n13712) );
  INV_X1 U13899 ( .A(b_7_), .ZN(n7843) );
  XOR2_X1 U13900 ( .A(n13899), .B(n13900), .Z(n13713) );
  XOR2_X1 U13901 ( .A(n13901), .B(n13902), .Z(n13900) );
  XOR2_X1 U13902 ( .A(n13903), .B(n13904), .Z(n13717) );
  XOR2_X1 U13903 ( .A(n13905), .B(n13906), .Z(n13904) );
  XOR2_X1 U13904 ( .A(n13907), .B(n13908), .Z(n13721) );
  XOR2_X1 U13905 ( .A(n13909), .B(n13910), .Z(n13908) );
  XOR2_X1 U13906 ( .A(n13911), .B(n13912), .Z(n13725) );
  XOR2_X1 U13907 ( .A(n13913), .B(n13914), .Z(n13912) );
  XOR2_X1 U13908 ( .A(n13915), .B(n13916), .Z(n13729) );
  XOR2_X1 U13909 ( .A(n13917), .B(n13918), .Z(n13916) );
  XOR2_X1 U13910 ( .A(n13919), .B(n13920), .Z(n13733) );
  XOR2_X1 U13911 ( .A(n13921), .B(n13922), .Z(n13920) );
  XOR2_X1 U13912 ( .A(n13923), .B(n13924), .Z(n13737) );
  XOR2_X1 U13913 ( .A(n13925), .B(n13926), .Z(n13924) );
  XOR2_X1 U13914 ( .A(n13927), .B(n13928), .Z(n13741) );
  XOR2_X1 U13915 ( .A(n13929), .B(n13930), .Z(n13928) );
  XOR2_X1 U13916 ( .A(n13931), .B(n13932), .Z(n13745) );
  XOR2_X1 U13917 ( .A(n13933), .B(n13934), .Z(n13932) );
  XOR2_X1 U13918 ( .A(n13935), .B(n13936), .Z(n13749) );
  XOR2_X1 U13919 ( .A(n13937), .B(n13938), .Z(n13936) );
  XOR2_X1 U13920 ( .A(n13939), .B(n13940), .Z(n13753) );
  XOR2_X1 U13921 ( .A(n13941), .B(n13942), .Z(n13940) );
  XOR2_X1 U13922 ( .A(n13943), .B(n13944), .Z(n13757) );
  XOR2_X1 U13923 ( .A(n13945), .B(n13946), .Z(n13944) );
  XOR2_X1 U13924 ( .A(n13947), .B(n13948), .Z(n13761) );
  XOR2_X1 U13925 ( .A(n13949), .B(n13950), .Z(n13948) );
  XOR2_X1 U13926 ( .A(n13951), .B(n13952), .Z(n13765) );
  XOR2_X1 U13927 ( .A(n13953), .B(n13954), .Z(n13952) );
  XOR2_X1 U13928 ( .A(n13955), .B(n13956), .Z(n13769) );
  XOR2_X1 U13929 ( .A(n13957), .B(n13958), .Z(n13956) );
  XOR2_X1 U13930 ( .A(n13959), .B(n13960), .Z(n13772) );
  XOR2_X1 U13931 ( .A(n13961), .B(n13962), .Z(n13960) );
  XNOR2_X1 U13932 ( .A(n13963), .B(n13964), .ZN(n13776) );
  XNOR2_X1 U13933 ( .A(n7972), .B(n13965), .ZN(n13963) );
  XOR2_X1 U13934 ( .A(n13966), .B(n13967), .Z(n13780) );
  XOR2_X1 U13935 ( .A(n13968), .B(n13969), .Z(n13967) );
  XOR2_X1 U13936 ( .A(n8480), .B(n13970), .Z(n8473) );
  XOR2_X1 U13937 ( .A(n8479), .B(n8478), .Z(n13970) );
  OR2_X1 U13938 ( .A1(n7971), .A2(n7963), .ZN(n8478) );
  OR2_X1 U13939 ( .A1(n13971), .A2(n13972), .ZN(n8479) );
  AND2_X1 U13940 ( .A1(n13969), .A2(n13968), .ZN(n13972) );
  AND2_X1 U13941 ( .A1(n13966), .A2(n13973), .ZN(n13971) );
  OR2_X1 U13942 ( .A1(n13968), .A2(n13969), .ZN(n13973) );
  OR2_X1 U13943 ( .A1(n7971), .A2(n7967), .ZN(n13969) );
  OR2_X1 U13944 ( .A1(n13974), .A2(n13975), .ZN(n13968) );
  AND2_X1 U13945 ( .A1(n13965), .A2(n7972), .ZN(n13975) );
  AND2_X1 U13946 ( .A1(n13964), .A2(n13976), .ZN(n13974) );
  OR2_X1 U13947 ( .A1(n7972), .A2(n13965), .ZN(n13976) );
  OR2_X1 U13948 ( .A1(n13977), .A2(n13978), .ZN(n13965) );
  AND2_X1 U13949 ( .A1(n13962), .A2(n13961), .ZN(n13978) );
  AND2_X1 U13950 ( .A1(n13959), .A2(n13979), .ZN(n13977) );
  OR2_X1 U13951 ( .A1(n13961), .A2(n13962), .ZN(n13979) );
  OR2_X1 U13952 ( .A1(n7971), .A2(n7974), .ZN(n13962) );
  OR2_X1 U13953 ( .A1(n13980), .A2(n13981), .ZN(n13961) );
  AND2_X1 U13954 ( .A1(n13958), .A2(n13957), .ZN(n13981) );
  AND2_X1 U13955 ( .A1(n13955), .A2(n13982), .ZN(n13980) );
  OR2_X1 U13956 ( .A1(n13957), .A2(n13958), .ZN(n13982) );
  OR2_X1 U13957 ( .A1(n7971), .A2(n7977), .ZN(n13958) );
  OR2_X1 U13958 ( .A1(n13983), .A2(n13984), .ZN(n13957) );
  AND2_X1 U13959 ( .A1(n13954), .A2(n13953), .ZN(n13984) );
  AND2_X1 U13960 ( .A1(n13951), .A2(n13985), .ZN(n13983) );
  OR2_X1 U13961 ( .A1(n13953), .A2(n13954), .ZN(n13985) );
  OR2_X1 U13962 ( .A1(n7971), .A2(n7981), .ZN(n13954) );
  OR2_X1 U13963 ( .A1(n13986), .A2(n13987), .ZN(n13953) );
  AND2_X1 U13964 ( .A1(n13950), .A2(n13949), .ZN(n13987) );
  AND2_X1 U13965 ( .A1(n13947), .A2(n13988), .ZN(n13986) );
  OR2_X1 U13966 ( .A1(n13949), .A2(n13950), .ZN(n13988) );
  OR2_X1 U13967 ( .A1(n7971), .A2(n7984), .ZN(n13950) );
  OR2_X1 U13968 ( .A1(n13989), .A2(n13990), .ZN(n13949) );
  AND2_X1 U13969 ( .A1(n13946), .A2(n13945), .ZN(n13990) );
  AND2_X1 U13970 ( .A1(n13943), .A2(n13991), .ZN(n13989) );
  OR2_X1 U13971 ( .A1(n13945), .A2(n13946), .ZN(n13991) );
  OR2_X1 U13972 ( .A1(n7971), .A2(n7988), .ZN(n13946) );
  OR2_X1 U13973 ( .A1(n13992), .A2(n13993), .ZN(n13945) );
  AND2_X1 U13974 ( .A1(n13942), .A2(n13941), .ZN(n13993) );
  AND2_X1 U13975 ( .A1(n13939), .A2(n13994), .ZN(n13992) );
  OR2_X1 U13976 ( .A1(n13941), .A2(n13942), .ZN(n13994) );
  OR2_X1 U13977 ( .A1(n7971), .A2(n7991), .ZN(n13942) );
  OR2_X1 U13978 ( .A1(n13995), .A2(n13996), .ZN(n13941) );
  AND2_X1 U13979 ( .A1(n13938), .A2(n13937), .ZN(n13996) );
  AND2_X1 U13980 ( .A1(n13935), .A2(n13997), .ZN(n13995) );
  OR2_X1 U13981 ( .A1(n13937), .A2(n13938), .ZN(n13997) );
  OR2_X1 U13982 ( .A1(n7971), .A2(n7995), .ZN(n13938) );
  OR2_X1 U13983 ( .A1(n13998), .A2(n13999), .ZN(n13937) );
  AND2_X1 U13984 ( .A1(n13934), .A2(n13933), .ZN(n13999) );
  AND2_X1 U13985 ( .A1(n13931), .A2(n14000), .ZN(n13998) );
  OR2_X1 U13986 ( .A1(n13933), .A2(n13934), .ZN(n14000) );
  OR2_X1 U13987 ( .A1(n7971), .A2(n7998), .ZN(n13934) );
  OR2_X1 U13988 ( .A1(n14001), .A2(n14002), .ZN(n13933) );
  AND2_X1 U13989 ( .A1(n13930), .A2(n13929), .ZN(n14002) );
  AND2_X1 U13990 ( .A1(n13927), .A2(n14003), .ZN(n14001) );
  OR2_X1 U13991 ( .A1(n13929), .A2(n13930), .ZN(n14003) );
  OR2_X1 U13992 ( .A1(n7971), .A2(n8002), .ZN(n13930) );
  OR2_X1 U13993 ( .A1(n14004), .A2(n14005), .ZN(n13929) );
  AND2_X1 U13994 ( .A1(n13926), .A2(n13925), .ZN(n14005) );
  AND2_X1 U13995 ( .A1(n13923), .A2(n14006), .ZN(n14004) );
  OR2_X1 U13996 ( .A1(n13925), .A2(n13926), .ZN(n14006) );
  OR2_X1 U13997 ( .A1(n7971), .A2(n8005), .ZN(n13926) );
  OR2_X1 U13998 ( .A1(n14007), .A2(n14008), .ZN(n13925) );
  AND2_X1 U13999 ( .A1(n13922), .A2(n13921), .ZN(n14008) );
  AND2_X1 U14000 ( .A1(n13919), .A2(n14009), .ZN(n14007) );
  OR2_X1 U14001 ( .A1(n13921), .A2(n13922), .ZN(n14009) );
  OR2_X1 U14002 ( .A1(n7971), .A2(n8009), .ZN(n13922) );
  OR2_X1 U14003 ( .A1(n14010), .A2(n14011), .ZN(n13921) );
  AND2_X1 U14004 ( .A1(n13918), .A2(n13917), .ZN(n14011) );
  AND2_X1 U14005 ( .A1(n13915), .A2(n14012), .ZN(n14010) );
  OR2_X1 U14006 ( .A1(n13917), .A2(n13918), .ZN(n14012) );
  OR2_X1 U14007 ( .A1(n7971), .A2(n8012), .ZN(n13918) );
  OR2_X1 U14008 ( .A1(n14013), .A2(n14014), .ZN(n13917) );
  AND2_X1 U14009 ( .A1(n13914), .A2(n13913), .ZN(n14014) );
  AND2_X1 U14010 ( .A1(n13911), .A2(n14015), .ZN(n14013) );
  OR2_X1 U14011 ( .A1(n13913), .A2(n13914), .ZN(n14015) );
  OR2_X1 U14012 ( .A1(n7971), .A2(n8016), .ZN(n13914) );
  OR2_X1 U14013 ( .A1(n14016), .A2(n14017), .ZN(n13913) );
  AND2_X1 U14014 ( .A1(n13910), .A2(n13909), .ZN(n14017) );
  AND2_X1 U14015 ( .A1(n13907), .A2(n14018), .ZN(n14016) );
  OR2_X1 U14016 ( .A1(n13909), .A2(n13910), .ZN(n14018) );
  OR2_X1 U14017 ( .A1(n7971), .A2(n8019), .ZN(n13910) );
  OR2_X1 U14018 ( .A1(n14019), .A2(n14020), .ZN(n13909) );
  AND2_X1 U14019 ( .A1(n13906), .A2(n13905), .ZN(n14020) );
  AND2_X1 U14020 ( .A1(n13903), .A2(n14021), .ZN(n14019) );
  OR2_X1 U14021 ( .A1(n13905), .A2(n13906), .ZN(n14021) );
  OR2_X1 U14022 ( .A1(n7971), .A2(n8023), .ZN(n13906) );
  OR2_X1 U14023 ( .A1(n14022), .A2(n14023), .ZN(n13905) );
  AND2_X1 U14024 ( .A1(n13902), .A2(n13901), .ZN(n14023) );
  AND2_X1 U14025 ( .A1(n13899), .A2(n14024), .ZN(n14022) );
  OR2_X1 U14026 ( .A1(n13901), .A2(n13902), .ZN(n14024) );
  OR2_X1 U14027 ( .A1(n7971), .A2(n8026), .ZN(n13902) );
  OR2_X1 U14028 ( .A1(n14025), .A2(n14026), .ZN(n13901) );
  AND2_X1 U14029 ( .A1(n13895), .A2(n13898), .ZN(n14026) );
  AND2_X1 U14030 ( .A1(n14027), .A2(n13897), .ZN(n14025) );
  OR2_X1 U14031 ( .A1(n14028), .A2(n14029), .ZN(n13897) );
  AND2_X1 U14032 ( .A1(n13894), .A2(n13893), .ZN(n14029) );
  AND2_X1 U14033 ( .A1(n13891), .A2(n14030), .ZN(n14028) );
  OR2_X1 U14034 ( .A1(n13893), .A2(n13894), .ZN(n14030) );
  OR2_X1 U14035 ( .A1(n7971), .A2(n8034), .ZN(n13894) );
  OR2_X1 U14036 ( .A1(n14031), .A2(n14032), .ZN(n13893) );
  AND2_X1 U14037 ( .A1(n13887), .A2(n13890), .ZN(n14032) );
  AND2_X1 U14038 ( .A1(n14033), .A2(n13889), .ZN(n14031) );
  OR2_X1 U14039 ( .A1(n14034), .A2(n14035), .ZN(n13889) );
  AND2_X1 U14040 ( .A1(n13883), .A2(n13886), .ZN(n14035) );
  AND2_X1 U14041 ( .A1(n14036), .A2(n13885), .ZN(n14034) );
  OR2_X1 U14042 ( .A1(n14037), .A2(n14038), .ZN(n13885) );
  AND2_X1 U14043 ( .A1(n13879), .A2(n13882), .ZN(n14038) );
  AND2_X1 U14044 ( .A1(n14039), .A2(n13881), .ZN(n14037) );
  OR2_X1 U14045 ( .A1(n14040), .A2(n14041), .ZN(n13881) );
  AND2_X1 U14046 ( .A1(n13875), .A2(n13878), .ZN(n14041) );
  AND2_X1 U14047 ( .A1(n14042), .A2(n13877), .ZN(n14040) );
  OR2_X1 U14048 ( .A1(n14043), .A2(n14044), .ZN(n13877) );
  AND2_X1 U14049 ( .A1(n13871), .A2(n14045), .ZN(n14044) );
  AND2_X1 U14050 ( .A1(n14046), .A2(n14047), .ZN(n14043) );
  OR2_X1 U14051 ( .A1(n14045), .A2(n13871), .ZN(n14047) );
  OR2_X1 U14052 ( .A1(n8051), .A2(n7971), .ZN(n13871) );
  INV_X1 U14053 ( .A(n13874), .ZN(n14045) );
  AND3_X1 U14054 ( .A1(n8904), .A2(b_6_), .A3(b_5_), .ZN(n13874) );
  INV_X1 U14055 ( .A(n13873), .ZN(n14046) );
  OR2_X1 U14056 ( .A1(n14048), .A2(n14049), .ZN(n13873) );
  AND2_X1 U14057 ( .A1(b_5_), .A2(n14050), .ZN(n14049) );
  OR2_X1 U14058 ( .A1(n14051), .A2(n7490), .ZN(n14050) );
  AND2_X1 U14059 ( .A1(a_30_), .A2(n7964), .ZN(n14051) );
  AND2_X1 U14060 ( .A1(b_4_), .A2(n14052), .ZN(n14048) );
  OR2_X1 U14061 ( .A1(n14053), .A2(n7493), .ZN(n14052) );
  AND2_X1 U14062 ( .A1(a_31_), .A2(n7872), .ZN(n14053) );
  OR2_X1 U14063 ( .A1(n13878), .A2(n13875), .ZN(n14042) );
  XNOR2_X1 U14064 ( .A(n14054), .B(n14055), .ZN(n13875) );
  XNOR2_X1 U14065 ( .A(n14056), .B(n14057), .ZN(n14055) );
  OR2_X1 U14066 ( .A1(n8048), .A2(n7971), .ZN(n13878) );
  OR2_X1 U14067 ( .A1(n13882), .A2(n13879), .ZN(n14039) );
  XOR2_X1 U14068 ( .A(n14058), .B(n14059), .Z(n13879) );
  XOR2_X1 U14069 ( .A(n14060), .B(n14061), .Z(n14059) );
  OR2_X1 U14070 ( .A1(n8044), .A2(n7971), .ZN(n13882) );
  OR2_X1 U14071 ( .A1(n13886), .A2(n13883), .ZN(n14036) );
  XOR2_X1 U14072 ( .A(n14062), .B(n14063), .Z(n13883) );
  XOR2_X1 U14073 ( .A(n14064), .B(n14065), .Z(n14063) );
  OR2_X1 U14074 ( .A1(n8041), .A2(n7971), .ZN(n13886) );
  OR2_X1 U14075 ( .A1(n13890), .A2(n13887), .ZN(n14033) );
  XOR2_X1 U14076 ( .A(n14066), .B(n14067), .Z(n13887) );
  XOR2_X1 U14077 ( .A(n14068), .B(n14069), .Z(n14067) );
  OR2_X1 U14078 ( .A1(n7971), .A2(n8037), .ZN(n13890) );
  XOR2_X1 U14079 ( .A(n14070), .B(n14071), .Z(n13891) );
  XOR2_X1 U14080 ( .A(n14072), .B(n14073), .Z(n14071) );
  OR2_X1 U14081 ( .A1(n13898), .A2(n13895), .ZN(n14027) );
  XOR2_X1 U14082 ( .A(n14074), .B(n14075), .Z(n13895) );
  XOR2_X1 U14083 ( .A(n14076), .B(n14077), .Z(n14075) );
  OR2_X1 U14084 ( .A1(n7971), .A2(n8030), .ZN(n13898) );
  INV_X1 U14085 ( .A(b_6_), .ZN(n7971) );
  XOR2_X1 U14086 ( .A(n14078), .B(n14079), .Z(n13899) );
  XOR2_X1 U14087 ( .A(n14080), .B(n14081), .Z(n14079) );
  XOR2_X1 U14088 ( .A(n14082), .B(n14083), .Z(n13903) );
  XOR2_X1 U14089 ( .A(n14084), .B(n14085), .Z(n14083) );
  XOR2_X1 U14090 ( .A(n14086), .B(n14087), .Z(n13907) );
  XOR2_X1 U14091 ( .A(n14088), .B(n14089), .Z(n14087) );
  XOR2_X1 U14092 ( .A(n14090), .B(n14091), .Z(n13911) );
  XOR2_X1 U14093 ( .A(n14092), .B(n14093), .Z(n14091) );
  XOR2_X1 U14094 ( .A(n14094), .B(n14095), .Z(n13915) );
  XOR2_X1 U14095 ( .A(n14096), .B(n14097), .Z(n14095) );
  XOR2_X1 U14096 ( .A(n14098), .B(n14099), .Z(n13919) );
  XOR2_X1 U14097 ( .A(n14100), .B(n14101), .Z(n14099) );
  XOR2_X1 U14098 ( .A(n14102), .B(n14103), .Z(n13923) );
  XOR2_X1 U14099 ( .A(n14104), .B(n14105), .Z(n14103) );
  XOR2_X1 U14100 ( .A(n14106), .B(n14107), .Z(n13927) );
  XOR2_X1 U14101 ( .A(n14108), .B(n14109), .Z(n14107) );
  XOR2_X1 U14102 ( .A(n14110), .B(n14111), .Z(n13931) );
  XOR2_X1 U14103 ( .A(n14112), .B(n14113), .Z(n14111) );
  XOR2_X1 U14104 ( .A(n14114), .B(n14115), .Z(n13935) );
  XOR2_X1 U14105 ( .A(n14116), .B(n14117), .Z(n14115) );
  XOR2_X1 U14106 ( .A(n14118), .B(n14119), .Z(n13939) );
  XOR2_X1 U14107 ( .A(n14120), .B(n14121), .Z(n14119) );
  XOR2_X1 U14108 ( .A(n14122), .B(n14123), .Z(n13943) );
  XOR2_X1 U14109 ( .A(n14124), .B(n14125), .Z(n14123) );
  XOR2_X1 U14110 ( .A(n14126), .B(n14127), .Z(n13947) );
  XOR2_X1 U14111 ( .A(n14128), .B(n14129), .Z(n14127) );
  XOR2_X1 U14112 ( .A(n14130), .B(n14131), .Z(n13951) );
  XOR2_X1 U14113 ( .A(n14132), .B(n14133), .Z(n14131) );
  XOR2_X1 U14114 ( .A(n14134), .B(n14135), .Z(n13955) );
  XOR2_X1 U14115 ( .A(n14136), .B(n14137), .Z(n14135) );
  XOR2_X1 U14116 ( .A(n14138), .B(n14139), .Z(n13959) );
  XOR2_X1 U14117 ( .A(n14140), .B(n14141), .Z(n14139) );
  INV_X1 U14118 ( .A(n7864), .ZN(n7972) );
  AND2_X1 U14119 ( .A1(b_6_), .A2(a_6_), .ZN(n7864) );
  XOR2_X1 U14120 ( .A(n14142), .B(n14143), .Z(n13964) );
  XOR2_X1 U14121 ( .A(n14144), .B(n14145), .Z(n14143) );
  XOR2_X1 U14122 ( .A(n14146), .B(n14147), .Z(n13966) );
  XOR2_X1 U14123 ( .A(n14148), .B(n14149), .Z(n14147) );
  XOR2_X1 U14124 ( .A(n8486), .B(n14150), .Z(n8480) );
  XNOR2_X1 U14125 ( .A(n8485), .B(n7876), .ZN(n14150) );
  AND2_X1 U14126 ( .A1(b_5_), .A2(a_5_), .ZN(n7876) );
  OR2_X1 U14127 ( .A1(n14151), .A2(n14152), .ZN(n8485) );
  AND2_X1 U14128 ( .A1(n14149), .A2(n14148), .ZN(n14152) );
  AND2_X1 U14129 ( .A1(n14146), .A2(n14153), .ZN(n14151) );
  OR2_X1 U14130 ( .A1(n14148), .A2(n14149), .ZN(n14153) );
  OR2_X1 U14131 ( .A1(n7872), .A2(n7970), .ZN(n14149) );
  OR2_X1 U14132 ( .A1(n14154), .A2(n14155), .ZN(n14148) );
  AND2_X1 U14133 ( .A1(n14145), .A2(n14144), .ZN(n14155) );
  AND2_X1 U14134 ( .A1(n14142), .A2(n14156), .ZN(n14154) );
  OR2_X1 U14135 ( .A1(n14144), .A2(n14145), .ZN(n14156) );
  OR2_X1 U14136 ( .A1(n7872), .A2(n7974), .ZN(n14145) );
  OR2_X1 U14137 ( .A1(n14157), .A2(n14158), .ZN(n14144) );
  AND2_X1 U14138 ( .A1(n14141), .A2(n14140), .ZN(n14158) );
  AND2_X1 U14139 ( .A1(n14138), .A2(n14159), .ZN(n14157) );
  OR2_X1 U14140 ( .A1(n14140), .A2(n14141), .ZN(n14159) );
  OR2_X1 U14141 ( .A1(n7872), .A2(n7977), .ZN(n14141) );
  OR2_X1 U14142 ( .A1(n14160), .A2(n14161), .ZN(n14140) );
  AND2_X1 U14143 ( .A1(n14137), .A2(n14136), .ZN(n14161) );
  AND2_X1 U14144 ( .A1(n14134), .A2(n14162), .ZN(n14160) );
  OR2_X1 U14145 ( .A1(n14136), .A2(n14137), .ZN(n14162) );
  OR2_X1 U14146 ( .A1(n7872), .A2(n7981), .ZN(n14137) );
  OR2_X1 U14147 ( .A1(n14163), .A2(n14164), .ZN(n14136) );
  AND2_X1 U14148 ( .A1(n14133), .A2(n14132), .ZN(n14164) );
  AND2_X1 U14149 ( .A1(n14130), .A2(n14165), .ZN(n14163) );
  OR2_X1 U14150 ( .A1(n14132), .A2(n14133), .ZN(n14165) );
  OR2_X1 U14151 ( .A1(n7872), .A2(n7984), .ZN(n14133) );
  OR2_X1 U14152 ( .A1(n14166), .A2(n14167), .ZN(n14132) );
  AND2_X1 U14153 ( .A1(n14129), .A2(n14128), .ZN(n14167) );
  AND2_X1 U14154 ( .A1(n14126), .A2(n14168), .ZN(n14166) );
  OR2_X1 U14155 ( .A1(n14128), .A2(n14129), .ZN(n14168) );
  OR2_X1 U14156 ( .A1(n7872), .A2(n7988), .ZN(n14129) );
  OR2_X1 U14157 ( .A1(n14169), .A2(n14170), .ZN(n14128) );
  AND2_X1 U14158 ( .A1(n14125), .A2(n14124), .ZN(n14170) );
  AND2_X1 U14159 ( .A1(n14122), .A2(n14171), .ZN(n14169) );
  OR2_X1 U14160 ( .A1(n14124), .A2(n14125), .ZN(n14171) );
  OR2_X1 U14161 ( .A1(n7872), .A2(n7991), .ZN(n14125) );
  OR2_X1 U14162 ( .A1(n14172), .A2(n14173), .ZN(n14124) );
  AND2_X1 U14163 ( .A1(n14121), .A2(n14120), .ZN(n14173) );
  AND2_X1 U14164 ( .A1(n14118), .A2(n14174), .ZN(n14172) );
  OR2_X1 U14165 ( .A1(n14120), .A2(n14121), .ZN(n14174) );
  OR2_X1 U14166 ( .A1(n7872), .A2(n7995), .ZN(n14121) );
  OR2_X1 U14167 ( .A1(n14175), .A2(n14176), .ZN(n14120) );
  AND2_X1 U14168 ( .A1(n14117), .A2(n14116), .ZN(n14176) );
  AND2_X1 U14169 ( .A1(n14114), .A2(n14177), .ZN(n14175) );
  OR2_X1 U14170 ( .A1(n14116), .A2(n14117), .ZN(n14177) );
  OR2_X1 U14171 ( .A1(n7872), .A2(n7998), .ZN(n14117) );
  OR2_X1 U14172 ( .A1(n14178), .A2(n14179), .ZN(n14116) );
  AND2_X1 U14173 ( .A1(n14113), .A2(n14112), .ZN(n14179) );
  AND2_X1 U14174 ( .A1(n14110), .A2(n14180), .ZN(n14178) );
  OR2_X1 U14175 ( .A1(n14112), .A2(n14113), .ZN(n14180) );
  OR2_X1 U14176 ( .A1(n7872), .A2(n8002), .ZN(n14113) );
  OR2_X1 U14177 ( .A1(n14181), .A2(n14182), .ZN(n14112) );
  AND2_X1 U14178 ( .A1(n14109), .A2(n14108), .ZN(n14182) );
  AND2_X1 U14179 ( .A1(n14106), .A2(n14183), .ZN(n14181) );
  OR2_X1 U14180 ( .A1(n14108), .A2(n14109), .ZN(n14183) );
  OR2_X1 U14181 ( .A1(n7872), .A2(n8005), .ZN(n14109) );
  OR2_X1 U14182 ( .A1(n14184), .A2(n14185), .ZN(n14108) );
  AND2_X1 U14183 ( .A1(n14105), .A2(n14104), .ZN(n14185) );
  AND2_X1 U14184 ( .A1(n14102), .A2(n14186), .ZN(n14184) );
  OR2_X1 U14185 ( .A1(n14104), .A2(n14105), .ZN(n14186) );
  OR2_X1 U14186 ( .A1(n7872), .A2(n8009), .ZN(n14105) );
  OR2_X1 U14187 ( .A1(n14187), .A2(n14188), .ZN(n14104) );
  AND2_X1 U14188 ( .A1(n14101), .A2(n14100), .ZN(n14188) );
  AND2_X1 U14189 ( .A1(n14098), .A2(n14189), .ZN(n14187) );
  OR2_X1 U14190 ( .A1(n14100), .A2(n14101), .ZN(n14189) );
  OR2_X1 U14191 ( .A1(n7872), .A2(n8012), .ZN(n14101) );
  OR2_X1 U14192 ( .A1(n14190), .A2(n14191), .ZN(n14100) );
  AND2_X1 U14193 ( .A1(n14097), .A2(n14096), .ZN(n14191) );
  AND2_X1 U14194 ( .A1(n14094), .A2(n14192), .ZN(n14190) );
  OR2_X1 U14195 ( .A1(n14096), .A2(n14097), .ZN(n14192) );
  OR2_X1 U14196 ( .A1(n7872), .A2(n8016), .ZN(n14097) );
  OR2_X1 U14197 ( .A1(n14193), .A2(n14194), .ZN(n14096) );
  AND2_X1 U14198 ( .A1(n14093), .A2(n14092), .ZN(n14194) );
  AND2_X1 U14199 ( .A1(n14090), .A2(n14195), .ZN(n14193) );
  OR2_X1 U14200 ( .A1(n14092), .A2(n14093), .ZN(n14195) );
  OR2_X1 U14201 ( .A1(n7872), .A2(n8019), .ZN(n14093) );
  OR2_X1 U14202 ( .A1(n14196), .A2(n14197), .ZN(n14092) );
  AND2_X1 U14203 ( .A1(n14089), .A2(n14088), .ZN(n14197) );
  AND2_X1 U14204 ( .A1(n14086), .A2(n14198), .ZN(n14196) );
  OR2_X1 U14205 ( .A1(n14088), .A2(n14089), .ZN(n14198) );
  OR2_X1 U14206 ( .A1(n7872), .A2(n8023), .ZN(n14089) );
  OR2_X1 U14207 ( .A1(n14199), .A2(n14200), .ZN(n14088) );
  AND2_X1 U14208 ( .A1(n14085), .A2(n14084), .ZN(n14200) );
  AND2_X1 U14209 ( .A1(n14082), .A2(n14201), .ZN(n14199) );
  OR2_X1 U14210 ( .A1(n14084), .A2(n14085), .ZN(n14201) );
  OR2_X1 U14211 ( .A1(n7872), .A2(n8026), .ZN(n14085) );
  OR2_X1 U14212 ( .A1(n14202), .A2(n14203), .ZN(n14084) );
  AND2_X1 U14213 ( .A1(n14081), .A2(n14080), .ZN(n14203) );
  AND2_X1 U14214 ( .A1(n14078), .A2(n14204), .ZN(n14202) );
  OR2_X1 U14215 ( .A1(n14080), .A2(n14081), .ZN(n14204) );
  OR2_X1 U14216 ( .A1(n7872), .A2(n8030), .ZN(n14081) );
  OR2_X1 U14217 ( .A1(n14205), .A2(n14206), .ZN(n14080) );
  AND2_X1 U14218 ( .A1(n14074), .A2(n14077), .ZN(n14206) );
  AND2_X1 U14219 ( .A1(n14207), .A2(n14076), .ZN(n14205) );
  OR2_X1 U14220 ( .A1(n14208), .A2(n14209), .ZN(n14076) );
  AND2_X1 U14221 ( .A1(n14073), .A2(n14072), .ZN(n14209) );
  AND2_X1 U14222 ( .A1(n14070), .A2(n14210), .ZN(n14208) );
  OR2_X1 U14223 ( .A1(n14072), .A2(n14073), .ZN(n14210) );
  OR2_X1 U14224 ( .A1(n8037), .A2(n7872), .ZN(n14073) );
  OR2_X1 U14225 ( .A1(n14211), .A2(n14212), .ZN(n14072) );
  AND2_X1 U14226 ( .A1(n14066), .A2(n14069), .ZN(n14212) );
  AND2_X1 U14227 ( .A1(n14213), .A2(n14068), .ZN(n14211) );
  OR2_X1 U14228 ( .A1(n14214), .A2(n14215), .ZN(n14068) );
  AND2_X1 U14229 ( .A1(n14062), .A2(n14065), .ZN(n14215) );
  AND2_X1 U14230 ( .A1(n14216), .A2(n14064), .ZN(n14214) );
  OR2_X1 U14231 ( .A1(n14217), .A2(n14218), .ZN(n14064) );
  AND2_X1 U14232 ( .A1(n14058), .A2(n14061), .ZN(n14218) );
  AND2_X1 U14233 ( .A1(n14219), .A2(n14060), .ZN(n14217) );
  OR2_X1 U14234 ( .A1(n14220), .A2(n14221), .ZN(n14060) );
  AND2_X1 U14235 ( .A1(n14054), .A2(n14222), .ZN(n14221) );
  AND2_X1 U14236 ( .A1(n14223), .A2(n14224), .ZN(n14220) );
  OR2_X1 U14237 ( .A1(n14222), .A2(n14054), .ZN(n14224) );
  OR2_X1 U14238 ( .A1(n8051), .A2(n7872), .ZN(n14054) );
  INV_X1 U14239 ( .A(n14057), .ZN(n14222) );
  AND3_X1 U14240 ( .A1(n8904), .A2(b_5_), .A3(b_4_), .ZN(n14057) );
  INV_X1 U14241 ( .A(n14056), .ZN(n14223) );
  OR2_X1 U14242 ( .A1(n14225), .A2(n14226), .ZN(n14056) );
  AND2_X1 U14243 ( .A1(b_4_), .A2(n14227), .ZN(n14226) );
  OR2_X1 U14244 ( .A1(n14228), .A2(n7490), .ZN(n14227) );
  AND2_X1 U14245 ( .A1(a_30_), .A2(n7901), .ZN(n14228) );
  AND2_X1 U14246 ( .A1(b_3_), .A2(n14229), .ZN(n14225) );
  OR2_X1 U14247 ( .A1(n14230), .A2(n7493), .ZN(n14229) );
  AND2_X1 U14248 ( .A1(a_31_), .A2(n7964), .ZN(n14230) );
  OR2_X1 U14249 ( .A1(n14061), .A2(n14058), .ZN(n14219) );
  XNOR2_X1 U14250 ( .A(n14231), .B(n14232), .ZN(n14058) );
  XNOR2_X1 U14251 ( .A(n14233), .B(n14234), .ZN(n14232) );
  OR2_X1 U14252 ( .A1(n8048), .A2(n7872), .ZN(n14061) );
  OR2_X1 U14253 ( .A1(n14065), .A2(n14062), .ZN(n14216) );
  XOR2_X1 U14254 ( .A(n14235), .B(n14236), .Z(n14062) );
  XOR2_X1 U14255 ( .A(n14237), .B(n14238), .Z(n14236) );
  OR2_X1 U14256 ( .A1(n8044), .A2(n7872), .ZN(n14065) );
  OR2_X1 U14257 ( .A1(n14069), .A2(n14066), .ZN(n14213) );
  XOR2_X1 U14258 ( .A(n14239), .B(n14240), .Z(n14066) );
  XOR2_X1 U14259 ( .A(n14241), .B(n14242), .Z(n14240) );
  OR2_X1 U14260 ( .A1(n8041), .A2(n7872), .ZN(n14069) );
  XOR2_X1 U14261 ( .A(n14243), .B(n14244), .Z(n14070) );
  XOR2_X1 U14262 ( .A(n14245), .B(n14246), .Z(n14244) );
  OR2_X1 U14263 ( .A1(n14077), .A2(n14074), .ZN(n14207) );
  XOR2_X1 U14264 ( .A(n14247), .B(n14248), .Z(n14074) );
  XOR2_X1 U14265 ( .A(n14249), .B(n14250), .Z(n14248) );
  OR2_X1 U14266 ( .A1(n7872), .A2(n8034), .ZN(n14077) );
  INV_X1 U14267 ( .A(b_5_), .ZN(n7872) );
  XOR2_X1 U14268 ( .A(n14251), .B(n14252), .Z(n14078) );
  XOR2_X1 U14269 ( .A(n14253), .B(n14254), .Z(n14252) );
  XOR2_X1 U14270 ( .A(n14255), .B(n14256), .Z(n14082) );
  XOR2_X1 U14271 ( .A(n14257), .B(n14258), .Z(n14256) );
  XOR2_X1 U14272 ( .A(n14259), .B(n14260), .Z(n14086) );
  XOR2_X1 U14273 ( .A(n14261), .B(n14262), .Z(n14260) );
  XOR2_X1 U14274 ( .A(n14263), .B(n14264), .Z(n14090) );
  XOR2_X1 U14275 ( .A(n14265), .B(n14266), .Z(n14264) );
  XOR2_X1 U14276 ( .A(n14267), .B(n14268), .Z(n14094) );
  XOR2_X1 U14277 ( .A(n14269), .B(n14270), .Z(n14268) );
  XOR2_X1 U14278 ( .A(n14271), .B(n14272), .Z(n14098) );
  XOR2_X1 U14279 ( .A(n14273), .B(n14274), .Z(n14272) );
  XOR2_X1 U14280 ( .A(n14275), .B(n14276), .Z(n14102) );
  XOR2_X1 U14281 ( .A(n14277), .B(n14278), .Z(n14276) );
  XOR2_X1 U14282 ( .A(n14279), .B(n14280), .Z(n14106) );
  XOR2_X1 U14283 ( .A(n14281), .B(n14282), .Z(n14280) );
  XOR2_X1 U14284 ( .A(n14283), .B(n14284), .Z(n14110) );
  XOR2_X1 U14285 ( .A(n14285), .B(n14286), .Z(n14284) );
  XOR2_X1 U14286 ( .A(n14287), .B(n14288), .Z(n14114) );
  XOR2_X1 U14287 ( .A(n14289), .B(n14290), .Z(n14288) );
  XOR2_X1 U14288 ( .A(n14291), .B(n14292), .Z(n14118) );
  XOR2_X1 U14289 ( .A(n14293), .B(n14294), .Z(n14292) );
  XOR2_X1 U14290 ( .A(n14295), .B(n14296), .Z(n14122) );
  XOR2_X1 U14291 ( .A(n14297), .B(n14298), .Z(n14296) );
  XOR2_X1 U14292 ( .A(n14299), .B(n14300), .Z(n14126) );
  XOR2_X1 U14293 ( .A(n14301), .B(n14302), .Z(n14300) );
  XOR2_X1 U14294 ( .A(n14303), .B(n14304), .Z(n14130) );
  XOR2_X1 U14295 ( .A(n14305), .B(n14306), .Z(n14304) );
  XOR2_X1 U14296 ( .A(n14307), .B(n14308), .Z(n14134) );
  XOR2_X1 U14297 ( .A(n14309), .B(n14310), .Z(n14308) );
  XOR2_X1 U14298 ( .A(n14311), .B(n14312), .Z(n14138) );
  XOR2_X1 U14299 ( .A(n14313), .B(n14314), .Z(n14312) );
  XOR2_X1 U14300 ( .A(n14315), .B(n14316), .Z(n14142) );
  XOR2_X1 U14301 ( .A(n14317), .B(n14318), .Z(n14316) );
  XOR2_X1 U14302 ( .A(n14319), .B(n14320), .Z(n14146) );
  XOR2_X1 U14303 ( .A(n14321), .B(n14322), .Z(n14320) );
  XOR2_X1 U14304 ( .A(n8493), .B(n14323), .Z(n8486) );
  XOR2_X1 U14305 ( .A(n8492), .B(n8491), .Z(n14323) );
  OR2_X1 U14306 ( .A1(n7964), .A2(n7970), .ZN(n8491) );
  OR2_X1 U14307 ( .A1(n14324), .A2(n14325), .ZN(n8492) );
  AND2_X1 U14308 ( .A1(n14322), .A2(n14321), .ZN(n14325) );
  AND2_X1 U14309 ( .A1(n14319), .A2(n14326), .ZN(n14324) );
  OR2_X1 U14310 ( .A1(n14321), .A2(n14322), .ZN(n14326) );
  OR2_X1 U14311 ( .A1(n7964), .A2(n7974), .ZN(n14322) );
  OR2_X1 U14312 ( .A1(n14327), .A2(n14328), .ZN(n14321) );
  AND2_X1 U14313 ( .A1(n14318), .A2(n14317), .ZN(n14328) );
  AND2_X1 U14314 ( .A1(n14315), .A2(n14329), .ZN(n14327) );
  OR2_X1 U14315 ( .A1(n14317), .A2(n14318), .ZN(n14329) );
  OR2_X1 U14316 ( .A1(n7964), .A2(n7977), .ZN(n14318) );
  OR2_X1 U14317 ( .A1(n14330), .A2(n14331), .ZN(n14317) );
  AND2_X1 U14318 ( .A1(n14314), .A2(n14313), .ZN(n14331) );
  AND2_X1 U14319 ( .A1(n14311), .A2(n14332), .ZN(n14330) );
  OR2_X1 U14320 ( .A1(n14313), .A2(n14314), .ZN(n14332) );
  OR2_X1 U14321 ( .A1(n7964), .A2(n7981), .ZN(n14314) );
  OR2_X1 U14322 ( .A1(n14333), .A2(n14334), .ZN(n14313) );
  AND2_X1 U14323 ( .A1(n14310), .A2(n14309), .ZN(n14334) );
  AND2_X1 U14324 ( .A1(n14307), .A2(n14335), .ZN(n14333) );
  OR2_X1 U14325 ( .A1(n14309), .A2(n14310), .ZN(n14335) );
  OR2_X1 U14326 ( .A1(n7964), .A2(n7984), .ZN(n14310) );
  OR2_X1 U14327 ( .A1(n14336), .A2(n14337), .ZN(n14309) );
  AND2_X1 U14328 ( .A1(n14306), .A2(n14305), .ZN(n14337) );
  AND2_X1 U14329 ( .A1(n14303), .A2(n14338), .ZN(n14336) );
  OR2_X1 U14330 ( .A1(n14305), .A2(n14306), .ZN(n14338) );
  OR2_X1 U14331 ( .A1(n7964), .A2(n7988), .ZN(n14306) );
  OR2_X1 U14332 ( .A1(n14339), .A2(n14340), .ZN(n14305) );
  AND2_X1 U14333 ( .A1(n14302), .A2(n14301), .ZN(n14340) );
  AND2_X1 U14334 ( .A1(n14299), .A2(n14341), .ZN(n14339) );
  OR2_X1 U14335 ( .A1(n14301), .A2(n14302), .ZN(n14341) );
  OR2_X1 U14336 ( .A1(n7964), .A2(n7991), .ZN(n14302) );
  OR2_X1 U14337 ( .A1(n14342), .A2(n14343), .ZN(n14301) );
  AND2_X1 U14338 ( .A1(n14298), .A2(n14297), .ZN(n14343) );
  AND2_X1 U14339 ( .A1(n14295), .A2(n14344), .ZN(n14342) );
  OR2_X1 U14340 ( .A1(n14297), .A2(n14298), .ZN(n14344) );
  OR2_X1 U14341 ( .A1(n7964), .A2(n7995), .ZN(n14298) );
  OR2_X1 U14342 ( .A1(n14345), .A2(n14346), .ZN(n14297) );
  AND2_X1 U14343 ( .A1(n14294), .A2(n14293), .ZN(n14346) );
  AND2_X1 U14344 ( .A1(n14291), .A2(n14347), .ZN(n14345) );
  OR2_X1 U14345 ( .A1(n14293), .A2(n14294), .ZN(n14347) );
  OR2_X1 U14346 ( .A1(n7964), .A2(n7998), .ZN(n14294) );
  OR2_X1 U14347 ( .A1(n14348), .A2(n14349), .ZN(n14293) );
  AND2_X1 U14348 ( .A1(n14290), .A2(n14289), .ZN(n14349) );
  AND2_X1 U14349 ( .A1(n14287), .A2(n14350), .ZN(n14348) );
  OR2_X1 U14350 ( .A1(n14289), .A2(n14290), .ZN(n14350) );
  OR2_X1 U14351 ( .A1(n7964), .A2(n8002), .ZN(n14290) );
  OR2_X1 U14352 ( .A1(n14351), .A2(n14352), .ZN(n14289) );
  AND2_X1 U14353 ( .A1(n14286), .A2(n14285), .ZN(n14352) );
  AND2_X1 U14354 ( .A1(n14283), .A2(n14353), .ZN(n14351) );
  OR2_X1 U14355 ( .A1(n14285), .A2(n14286), .ZN(n14353) );
  OR2_X1 U14356 ( .A1(n7964), .A2(n8005), .ZN(n14286) );
  OR2_X1 U14357 ( .A1(n14354), .A2(n14355), .ZN(n14285) );
  AND2_X1 U14358 ( .A1(n14282), .A2(n14281), .ZN(n14355) );
  AND2_X1 U14359 ( .A1(n14279), .A2(n14356), .ZN(n14354) );
  OR2_X1 U14360 ( .A1(n14281), .A2(n14282), .ZN(n14356) );
  OR2_X1 U14361 ( .A1(n7964), .A2(n8009), .ZN(n14282) );
  OR2_X1 U14362 ( .A1(n14357), .A2(n14358), .ZN(n14281) );
  AND2_X1 U14363 ( .A1(n14278), .A2(n14277), .ZN(n14358) );
  AND2_X1 U14364 ( .A1(n14275), .A2(n14359), .ZN(n14357) );
  OR2_X1 U14365 ( .A1(n14277), .A2(n14278), .ZN(n14359) );
  OR2_X1 U14366 ( .A1(n7964), .A2(n8012), .ZN(n14278) );
  OR2_X1 U14367 ( .A1(n14360), .A2(n14361), .ZN(n14277) );
  AND2_X1 U14368 ( .A1(n14274), .A2(n14273), .ZN(n14361) );
  AND2_X1 U14369 ( .A1(n14271), .A2(n14362), .ZN(n14360) );
  OR2_X1 U14370 ( .A1(n14273), .A2(n14274), .ZN(n14362) );
  OR2_X1 U14371 ( .A1(n7964), .A2(n8016), .ZN(n14274) );
  OR2_X1 U14372 ( .A1(n14363), .A2(n14364), .ZN(n14273) );
  AND2_X1 U14373 ( .A1(n14270), .A2(n14269), .ZN(n14364) );
  AND2_X1 U14374 ( .A1(n14267), .A2(n14365), .ZN(n14363) );
  OR2_X1 U14375 ( .A1(n14269), .A2(n14270), .ZN(n14365) );
  OR2_X1 U14376 ( .A1(n7964), .A2(n8019), .ZN(n14270) );
  OR2_X1 U14377 ( .A1(n14366), .A2(n14367), .ZN(n14269) );
  AND2_X1 U14378 ( .A1(n14266), .A2(n14265), .ZN(n14367) );
  AND2_X1 U14379 ( .A1(n14263), .A2(n14368), .ZN(n14366) );
  OR2_X1 U14380 ( .A1(n14265), .A2(n14266), .ZN(n14368) );
  OR2_X1 U14381 ( .A1(n7964), .A2(n8023), .ZN(n14266) );
  OR2_X1 U14382 ( .A1(n14369), .A2(n14370), .ZN(n14265) );
  AND2_X1 U14383 ( .A1(n14262), .A2(n14261), .ZN(n14370) );
  AND2_X1 U14384 ( .A1(n14259), .A2(n14371), .ZN(n14369) );
  OR2_X1 U14385 ( .A1(n14261), .A2(n14262), .ZN(n14371) );
  OR2_X1 U14386 ( .A1(n7964), .A2(n8026), .ZN(n14262) );
  OR2_X1 U14387 ( .A1(n14372), .A2(n14373), .ZN(n14261) );
  AND2_X1 U14388 ( .A1(n14258), .A2(n14257), .ZN(n14373) );
  AND2_X1 U14389 ( .A1(n14255), .A2(n14374), .ZN(n14372) );
  OR2_X1 U14390 ( .A1(n14257), .A2(n14258), .ZN(n14374) );
  OR2_X1 U14391 ( .A1(n7964), .A2(n8030), .ZN(n14258) );
  OR2_X1 U14392 ( .A1(n14375), .A2(n14376), .ZN(n14257) );
  AND2_X1 U14393 ( .A1(n14254), .A2(n14253), .ZN(n14376) );
  AND2_X1 U14394 ( .A1(n14251), .A2(n14377), .ZN(n14375) );
  OR2_X1 U14395 ( .A1(n14253), .A2(n14254), .ZN(n14377) );
  OR2_X1 U14396 ( .A1(n8034), .A2(n7964), .ZN(n14254) );
  OR2_X1 U14397 ( .A1(n14378), .A2(n14379), .ZN(n14253) );
  AND2_X1 U14398 ( .A1(n14247), .A2(n14250), .ZN(n14379) );
  AND2_X1 U14399 ( .A1(n14380), .A2(n14249), .ZN(n14378) );
  OR2_X1 U14400 ( .A1(n14381), .A2(n14382), .ZN(n14249) );
  AND2_X1 U14401 ( .A1(n14246), .A2(n14245), .ZN(n14382) );
  AND2_X1 U14402 ( .A1(n14243), .A2(n14383), .ZN(n14381) );
  OR2_X1 U14403 ( .A1(n14245), .A2(n14246), .ZN(n14383) );
  OR2_X1 U14404 ( .A1(n8041), .A2(n7964), .ZN(n14246) );
  OR2_X1 U14405 ( .A1(n14384), .A2(n14385), .ZN(n14245) );
  AND2_X1 U14406 ( .A1(n14239), .A2(n14242), .ZN(n14385) );
  AND2_X1 U14407 ( .A1(n14386), .A2(n14241), .ZN(n14384) );
  OR2_X1 U14408 ( .A1(n14387), .A2(n14388), .ZN(n14241) );
  AND2_X1 U14409 ( .A1(n14235), .A2(n14238), .ZN(n14388) );
  AND2_X1 U14410 ( .A1(n14389), .A2(n14237), .ZN(n14387) );
  OR2_X1 U14411 ( .A1(n14390), .A2(n14391), .ZN(n14237) );
  AND2_X1 U14412 ( .A1(n14231), .A2(n14392), .ZN(n14391) );
  AND2_X1 U14413 ( .A1(n14393), .A2(n14394), .ZN(n14390) );
  OR2_X1 U14414 ( .A1(n14392), .A2(n14231), .ZN(n14394) );
  OR2_X1 U14415 ( .A1(n8051), .A2(n7964), .ZN(n14231) );
  INV_X1 U14416 ( .A(n14234), .ZN(n14392) );
  AND3_X1 U14417 ( .A1(n8904), .A2(b_4_), .A3(b_3_), .ZN(n14234) );
  INV_X1 U14418 ( .A(n14233), .ZN(n14393) );
  OR2_X1 U14419 ( .A1(n14395), .A2(n14396), .ZN(n14233) );
  AND2_X1 U14420 ( .A1(b_3_), .A2(n14397), .ZN(n14396) );
  OR2_X1 U14421 ( .A1(n14398), .A2(n7490), .ZN(n14397) );
  AND2_X1 U14422 ( .A1(a_30_), .A2(n7957), .ZN(n14398) );
  AND2_X1 U14423 ( .A1(b_2_), .A2(n14399), .ZN(n14395) );
  OR2_X1 U14424 ( .A1(n14400), .A2(n7493), .ZN(n14399) );
  AND2_X1 U14425 ( .A1(a_31_), .A2(n7901), .ZN(n14400) );
  OR2_X1 U14426 ( .A1(n14238), .A2(n14235), .ZN(n14389) );
  XNOR2_X1 U14427 ( .A(n14401), .B(n14402), .ZN(n14235) );
  XNOR2_X1 U14428 ( .A(n14403), .B(n14404), .ZN(n14402) );
  OR2_X1 U14429 ( .A1(n8048), .A2(n7964), .ZN(n14238) );
  OR2_X1 U14430 ( .A1(n14242), .A2(n14239), .ZN(n14386) );
  XOR2_X1 U14431 ( .A(n14405), .B(n14406), .Z(n14239) );
  XOR2_X1 U14432 ( .A(n14407), .B(n14408), .Z(n14406) );
  OR2_X1 U14433 ( .A1(n8044), .A2(n7964), .ZN(n14242) );
  XOR2_X1 U14434 ( .A(n14409), .B(n14410), .Z(n14243) );
  XOR2_X1 U14435 ( .A(n14411), .B(n14412), .Z(n14410) );
  OR2_X1 U14436 ( .A1(n14250), .A2(n14247), .ZN(n14380) );
  XOR2_X1 U14437 ( .A(n14413), .B(n14414), .Z(n14247) );
  XOR2_X1 U14438 ( .A(n14415), .B(n14416), .Z(n14414) );
  OR2_X1 U14439 ( .A1(n8037), .A2(n7964), .ZN(n14250) );
  INV_X1 U14440 ( .A(b_4_), .ZN(n7964) );
  XOR2_X1 U14441 ( .A(n14417), .B(n14418), .Z(n14251) );
  XOR2_X1 U14442 ( .A(n14419), .B(n14420), .Z(n14418) );
  XOR2_X1 U14443 ( .A(n14421), .B(n14422), .Z(n14255) );
  XOR2_X1 U14444 ( .A(n14423), .B(n14424), .Z(n14422) );
  XOR2_X1 U14445 ( .A(n14425), .B(n14426), .Z(n14259) );
  XOR2_X1 U14446 ( .A(n14427), .B(n14428), .Z(n14426) );
  XOR2_X1 U14447 ( .A(n14429), .B(n14430), .Z(n14263) );
  XOR2_X1 U14448 ( .A(n14431), .B(n14432), .Z(n14430) );
  XOR2_X1 U14449 ( .A(n14433), .B(n14434), .Z(n14267) );
  XOR2_X1 U14450 ( .A(n14435), .B(n14436), .Z(n14434) );
  XOR2_X1 U14451 ( .A(n14437), .B(n14438), .Z(n14271) );
  XOR2_X1 U14452 ( .A(n14439), .B(n14440), .Z(n14438) );
  XOR2_X1 U14453 ( .A(n14441), .B(n14442), .Z(n14275) );
  XOR2_X1 U14454 ( .A(n14443), .B(n14444), .Z(n14442) );
  XOR2_X1 U14455 ( .A(n14445), .B(n14446), .Z(n14279) );
  XOR2_X1 U14456 ( .A(n14447), .B(n14448), .Z(n14446) );
  XOR2_X1 U14457 ( .A(n14449), .B(n14450), .Z(n14283) );
  XOR2_X1 U14458 ( .A(n14451), .B(n14452), .Z(n14450) );
  XOR2_X1 U14459 ( .A(n14453), .B(n14454), .Z(n14287) );
  XOR2_X1 U14460 ( .A(n14455), .B(n14456), .Z(n14454) );
  XOR2_X1 U14461 ( .A(n14457), .B(n14458), .Z(n14291) );
  XOR2_X1 U14462 ( .A(n14459), .B(n14460), .Z(n14458) );
  XOR2_X1 U14463 ( .A(n14461), .B(n14462), .Z(n14295) );
  XOR2_X1 U14464 ( .A(n14463), .B(n14464), .Z(n14462) );
  XOR2_X1 U14465 ( .A(n14465), .B(n14466), .Z(n14299) );
  XOR2_X1 U14466 ( .A(n14467), .B(n14468), .Z(n14466) );
  XOR2_X1 U14467 ( .A(n14469), .B(n14470), .Z(n14303) );
  XOR2_X1 U14468 ( .A(n14471), .B(n14472), .Z(n14470) );
  XOR2_X1 U14469 ( .A(n14473), .B(n14474), .Z(n14307) );
  XOR2_X1 U14470 ( .A(n14475), .B(n14476), .Z(n14474) );
  XOR2_X1 U14471 ( .A(n14477), .B(n14478), .Z(n14311) );
  XOR2_X1 U14472 ( .A(n14479), .B(n14480), .Z(n14478) );
  XOR2_X1 U14473 ( .A(n14481), .B(n14482), .Z(n14315) );
  XOR2_X1 U14474 ( .A(n14483), .B(n14484), .Z(n14482) );
  XOR2_X1 U14475 ( .A(n14485), .B(n14486), .Z(n14319) );
  XOR2_X1 U14476 ( .A(n14487), .B(n14488), .Z(n14486) );
  XOR2_X1 U14477 ( .A(n8500), .B(n14489), .Z(n8493) );
  XOR2_X1 U14478 ( .A(n8499), .B(n8498), .Z(n14489) );
  OR2_X1 U14479 ( .A1(n7901), .A2(n7974), .ZN(n8498) );
  OR2_X1 U14480 ( .A1(n14490), .A2(n14491), .ZN(n8499) );
  AND2_X1 U14481 ( .A1(n14488), .A2(n14487), .ZN(n14491) );
  AND2_X1 U14482 ( .A1(n14485), .A2(n14492), .ZN(n14490) );
  OR2_X1 U14483 ( .A1(n14487), .A2(n14488), .ZN(n14492) );
  OR2_X1 U14484 ( .A1(n7901), .A2(n7977), .ZN(n14488) );
  OR2_X1 U14485 ( .A1(n14493), .A2(n14494), .ZN(n14487) );
  AND2_X1 U14486 ( .A1(n14484), .A2(n14483), .ZN(n14494) );
  AND2_X1 U14487 ( .A1(n14481), .A2(n14495), .ZN(n14493) );
  OR2_X1 U14488 ( .A1(n14483), .A2(n14484), .ZN(n14495) );
  OR2_X1 U14489 ( .A1(n7901), .A2(n7981), .ZN(n14484) );
  OR2_X1 U14490 ( .A1(n14496), .A2(n14497), .ZN(n14483) );
  AND2_X1 U14491 ( .A1(n14480), .A2(n14479), .ZN(n14497) );
  AND2_X1 U14492 ( .A1(n14477), .A2(n14498), .ZN(n14496) );
  OR2_X1 U14493 ( .A1(n14479), .A2(n14480), .ZN(n14498) );
  OR2_X1 U14494 ( .A1(n7901), .A2(n7984), .ZN(n14480) );
  OR2_X1 U14495 ( .A1(n14499), .A2(n14500), .ZN(n14479) );
  AND2_X1 U14496 ( .A1(n14476), .A2(n14475), .ZN(n14500) );
  AND2_X1 U14497 ( .A1(n14473), .A2(n14501), .ZN(n14499) );
  OR2_X1 U14498 ( .A1(n14475), .A2(n14476), .ZN(n14501) );
  OR2_X1 U14499 ( .A1(n7901), .A2(n7988), .ZN(n14476) );
  OR2_X1 U14500 ( .A1(n14502), .A2(n14503), .ZN(n14475) );
  AND2_X1 U14501 ( .A1(n14472), .A2(n14471), .ZN(n14503) );
  AND2_X1 U14502 ( .A1(n14469), .A2(n14504), .ZN(n14502) );
  OR2_X1 U14503 ( .A1(n14471), .A2(n14472), .ZN(n14504) );
  OR2_X1 U14504 ( .A1(n7901), .A2(n7991), .ZN(n14472) );
  OR2_X1 U14505 ( .A1(n14505), .A2(n14506), .ZN(n14471) );
  AND2_X1 U14506 ( .A1(n14468), .A2(n14467), .ZN(n14506) );
  AND2_X1 U14507 ( .A1(n14465), .A2(n14507), .ZN(n14505) );
  OR2_X1 U14508 ( .A1(n14467), .A2(n14468), .ZN(n14507) );
  OR2_X1 U14509 ( .A1(n7901), .A2(n7995), .ZN(n14468) );
  OR2_X1 U14510 ( .A1(n14508), .A2(n14509), .ZN(n14467) );
  AND2_X1 U14511 ( .A1(n14464), .A2(n14463), .ZN(n14509) );
  AND2_X1 U14512 ( .A1(n14461), .A2(n14510), .ZN(n14508) );
  OR2_X1 U14513 ( .A1(n14463), .A2(n14464), .ZN(n14510) );
  OR2_X1 U14514 ( .A1(n7901), .A2(n7998), .ZN(n14464) );
  OR2_X1 U14515 ( .A1(n14511), .A2(n14512), .ZN(n14463) );
  AND2_X1 U14516 ( .A1(n14460), .A2(n14459), .ZN(n14512) );
  AND2_X1 U14517 ( .A1(n14457), .A2(n14513), .ZN(n14511) );
  OR2_X1 U14518 ( .A1(n14459), .A2(n14460), .ZN(n14513) );
  OR2_X1 U14519 ( .A1(n7901), .A2(n8002), .ZN(n14460) );
  OR2_X1 U14520 ( .A1(n14514), .A2(n14515), .ZN(n14459) );
  AND2_X1 U14521 ( .A1(n14456), .A2(n14455), .ZN(n14515) );
  AND2_X1 U14522 ( .A1(n14453), .A2(n14516), .ZN(n14514) );
  OR2_X1 U14523 ( .A1(n14455), .A2(n14456), .ZN(n14516) );
  OR2_X1 U14524 ( .A1(n7901), .A2(n8005), .ZN(n14456) );
  OR2_X1 U14525 ( .A1(n14517), .A2(n14518), .ZN(n14455) );
  AND2_X1 U14526 ( .A1(n14452), .A2(n14451), .ZN(n14518) );
  AND2_X1 U14527 ( .A1(n14449), .A2(n14519), .ZN(n14517) );
  OR2_X1 U14528 ( .A1(n14451), .A2(n14452), .ZN(n14519) );
  OR2_X1 U14529 ( .A1(n7901), .A2(n8009), .ZN(n14452) );
  OR2_X1 U14530 ( .A1(n14520), .A2(n14521), .ZN(n14451) );
  AND2_X1 U14531 ( .A1(n14448), .A2(n14447), .ZN(n14521) );
  AND2_X1 U14532 ( .A1(n14445), .A2(n14522), .ZN(n14520) );
  OR2_X1 U14533 ( .A1(n14447), .A2(n14448), .ZN(n14522) );
  OR2_X1 U14534 ( .A1(n7901), .A2(n8012), .ZN(n14448) );
  OR2_X1 U14535 ( .A1(n14523), .A2(n14524), .ZN(n14447) );
  AND2_X1 U14536 ( .A1(n14444), .A2(n14443), .ZN(n14524) );
  AND2_X1 U14537 ( .A1(n14441), .A2(n14525), .ZN(n14523) );
  OR2_X1 U14538 ( .A1(n14443), .A2(n14444), .ZN(n14525) );
  OR2_X1 U14539 ( .A1(n7901), .A2(n8016), .ZN(n14444) );
  OR2_X1 U14540 ( .A1(n14526), .A2(n14527), .ZN(n14443) );
  AND2_X1 U14541 ( .A1(n14440), .A2(n14439), .ZN(n14527) );
  AND2_X1 U14542 ( .A1(n14437), .A2(n14528), .ZN(n14526) );
  OR2_X1 U14543 ( .A1(n14439), .A2(n14440), .ZN(n14528) );
  OR2_X1 U14544 ( .A1(n7901), .A2(n8019), .ZN(n14440) );
  OR2_X1 U14545 ( .A1(n14529), .A2(n14530), .ZN(n14439) );
  AND2_X1 U14546 ( .A1(n14436), .A2(n14435), .ZN(n14530) );
  AND2_X1 U14547 ( .A1(n14433), .A2(n14531), .ZN(n14529) );
  OR2_X1 U14548 ( .A1(n14435), .A2(n14436), .ZN(n14531) );
  OR2_X1 U14549 ( .A1(n7901), .A2(n8023), .ZN(n14436) );
  OR2_X1 U14550 ( .A1(n14532), .A2(n14533), .ZN(n14435) );
  AND2_X1 U14551 ( .A1(n14432), .A2(n14431), .ZN(n14533) );
  AND2_X1 U14552 ( .A1(n14429), .A2(n14534), .ZN(n14532) );
  OR2_X1 U14553 ( .A1(n14431), .A2(n14432), .ZN(n14534) );
  OR2_X1 U14554 ( .A1(n7901), .A2(n8026), .ZN(n14432) );
  OR2_X1 U14555 ( .A1(n14535), .A2(n14536), .ZN(n14431) );
  AND2_X1 U14556 ( .A1(n14428), .A2(n14427), .ZN(n14536) );
  AND2_X1 U14557 ( .A1(n14425), .A2(n14537), .ZN(n14535) );
  OR2_X1 U14558 ( .A1(n14427), .A2(n14428), .ZN(n14537) );
  OR2_X1 U14559 ( .A1(n8030), .A2(n7901), .ZN(n14428) );
  OR2_X1 U14560 ( .A1(n14538), .A2(n14539), .ZN(n14427) );
  AND2_X1 U14561 ( .A1(n14424), .A2(n14423), .ZN(n14539) );
  AND2_X1 U14562 ( .A1(n14421), .A2(n14540), .ZN(n14538) );
  OR2_X1 U14563 ( .A1(n14423), .A2(n14424), .ZN(n14540) );
  OR2_X1 U14564 ( .A1(n8034), .A2(n7901), .ZN(n14424) );
  OR2_X1 U14565 ( .A1(n14541), .A2(n14542), .ZN(n14423) );
  AND2_X1 U14566 ( .A1(n14420), .A2(n14419), .ZN(n14542) );
  AND2_X1 U14567 ( .A1(n14417), .A2(n14543), .ZN(n14541) );
  OR2_X1 U14568 ( .A1(n14419), .A2(n14420), .ZN(n14543) );
  OR2_X1 U14569 ( .A1(n8037), .A2(n7901), .ZN(n14420) );
  OR2_X1 U14570 ( .A1(n14544), .A2(n14545), .ZN(n14419) );
  AND2_X1 U14571 ( .A1(n14413), .A2(n14416), .ZN(n14545) );
  AND2_X1 U14572 ( .A1(n14546), .A2(n14415), .ZN(n14544) );
  OR2_X1 U14573 ( .A1(n14547), .A2(n14548), .ZN(n14415) );
  AND2_X1 U14574 ( .A1(n14412), .A2(n14411), .ZN(n14548) );
  AND2_X1 U14575 ( .A1(n14409), .A2(n14549), .ZN(n14547) );
  OR2_X1 U14576 ( .A1(n14411), .A2(n14412), .ZN(n14549) );
  OR2_X1 U14577 ( .A1(n8044), .A2(n7901), .ZN(n14412) );
  OR2_X1 U14578 ( .A1(n14550), .A2(n14551), .ZN(n14411) );
  AND2_X1 U14579 ( .A1(n14405), .A2(n14408), .ZN(n14551) );
  AND2_X1 U14580 ( .A1(n14552), .A2(n14407), .ZN(n14550) );
  OR2_X1 U14581 ( .A1(n14553), .A2(n14554), .ZN(n14407) );
  AND2_X1 U14582 ( .A1(n14401), .A2(n14555), .ZN(n14554) );
  AND2_X1 U14583 ( .A1(n14556), .A2(n14557), .ZN(n14553) );
  OR2_X1 U14584 ( .A1(n14555), .A2(n14401), .ZN(n14557) );
  OR2_X1 U14585 ( .A1(n8051), .A2(n7901), .ZN(n14401) );
  INV_X1 U14586 ( .A(n14404), .ZN(n14555) );
  AND3_X1 U14587 ( .A1(n8904), .A2(b_3_), .A3(b_2_), .ZN(n14404) );
  INV_X1 U14588 ( .A(n14403), .ZN(n14556) );
  OR2_X1 U14589 ( .A1(n14558), .A2(n14559), .ZN(n14403) );
  AND2_X1 U14590 ( .A1(b_2_), .A2(n14560), .ZN(n14559) );
  OR2_X1 U14591 ( .A1(n14561), .A2(n7490), .ZN(n14560) );
  AND2_X1 U14592 ( .A1(a_30_), .A2(n7930), .ZN(n14561) );
  AND2_X1 U14593 ( .A1(b_1_), .A2(n14562), .ZN(n14558) );
  OR2_X1 U14594 ( .A1(n14563), .A2(n7493), .ZN(n14562) );
  AND2_X1 U14595 ( .A1(a_31_), .A2(n7957), .ZN(n14563) );
  OR2_X1 U14596 ( .A1(n14408), .A2(n14405), .ZN(n14552) );
  XNOR2_X1 U14597 ( .A(n14564), .B(n14565), .ZN(n14405) );
  XNOR2_X1 U14598 ( .A(n14566), .B(n14567), .ZN(n14565) );
  OR2_X1 U14599 ( .A1(n8048), .A2(n7901), .ZN(n14408) );
  XOR2_X1 U14600 ( .A(n14568), .B(n14569), .Z(n14409) );
  XOR2_X1 U14601 ( .A(n14570), .B(n14571), .Z(n14569) );
  OR2_X1 U14602 ( .A1(n14416), .A2(n14413), .ZN(n14546) );
  XOR2_X1 U14603 ( .A(n14572), .B(n14573), .Z(n14413) );
  XOR2_X1 U14604 ( .A(n14574), .B(n14575), .Z(n14573) );
  OR2_X1 U14605 ( .A1(n8041), .A2(n7901), .ZN(n14416) );
  INV_X1 U14606 ( .A(b_3_), .ZN(n7901) );
  XOR2_X1 U14607 ( .A(n14576), .B(n14577), .Z(n14417) );
  XOR2_X1 U14608 ( .A(n14578), .B(n14579), .Z(n14577) );
  XOR2_X1 U14609 ( .A(n14580), .B(n14581), .Z(n14421) );
  XOR2_X1 U14610 ( .A(n14582), .B(n14583), .Z(n14581) );
  XOR2_X1 U14611 ( .A(n14584), .B(n14585), .Z(n14425) );
  XOR2_X1 U14612 ( .A(n14586), .B(n14587), .Z(n14585) );
  XOR2_X1 U14613 ( .A(n14588), .B(n14589), .Z(n14429) );
  XOR2_X1 U14614 ( .A(n14590), .B(n14591), .Z(n14589) );
  XOR2_X1 U14615 ( .A(n14592), .B(n14593), .Z(n14433) );
  XOR2_X1 U14616 ( .A(n14594), .B(n14595), .Z(n14593) );
  XOR2_X1 U14617 ( .A(n14596), .B(n14597), .Z(n14437) );
  XOR2_X1 U14618 ( .A(n14598), .B(n14599), .Z(n14597) );
  XOR2_X1 U14619 ( .A(n14600), .B(n14601), .Z(n14441) );
  XOR2_X1 U14620 ( .A(n14602), .B(n14603), .Z(n14601) );
  XOR2_X1 U14621 ( .A(n14604), .B(n14605), .Z(n14445) );
  XOR2_X1 U14622 ( .A(n14606), .B(n14607), .Z(n14605) );
  XOR2_X1 U14623 ( .A(n14608), .B(n14609), .Z(n14449) );
  XOR2_X1 U14624 ( .A(n14610), .B(n14611), .Z(n14609) );
  XOR2_X1 U14625 ( .A(n14612), .B(n14613), .Z(n14453) );
  XOR2_X1 U14626 ( .A(n14614), .B(n14615), .Z(n14613) );
  XOR2_X1 U14627 ( .A(n14616), .B(n14617), .Z(n14457) );
  XOR2_X1 U14628 ( .A(n14618), .B(n14619), .Z(n14617) );
  XOR2_X1 U14629 ( .A(n14620), .B(n14621), .Z(n14461) );
  XOR2_X1 U14630 ( .A(n14622), .B(n14623), .Z(n14621) );
  XOR2_X1 U14631 ( .A(n14624), .B(n14625), .Z(n14465) );
  XOR2_X1 U14632 ( .A(n14626), .B(n14627), .Z(n14625) );
  XOR2_X1 U14633 ( .A(n14628), .B(n14629), .Z(n14469) );
  XOR2_X1 U14634 ( .A(n14630), .B(n14631), .Z(n14629) );
  XOR2_X1 U14635 ( .A(n14632), .B(n14633), .Z(n14473) );
  XOR2_X1 U14636 ( .A(n14634), .B(n14635), .Z(n14633) );
  XOR2_X1 U14637 ( .A(n14636), .B(n14637), .Z(n14477) );
  XOR2_X1 U14638 ( .A(n14638), .B(n14639), .Z(n14637) );
  XOR2_X1 U14639 ( .A(n14640), .B(n14641), .Z(n14481) );
  XOR2_X1 U14640 ( .A(n14642), .B(n14643), .Z(n14641) );
  XOR2_X1 U14641 ( .A(n14644), .B(n14645), .Z(n14485) );
  XOR2_X1 U14642 ( .A(n14646), .B(n14647), .Z(n14645) );
  XOR2_X1 U14643 ( .A(n14648), .B(n14649), .Z(n8500) );
  XOR2_X1 U14644 ( .A(n14650), .B(n14651), .Z(n14649) );
  AND3_X1 U14645 ( .A1(n8130), .A2(n8128), .A3(n8129), .ZN(n8131) );
  INV_X1 U14646 ( .A(n8197), .ZN(n8129) );
  OR2_X1 U14647 ( .A1(n14652), .A2(n14653), .ZN(n8197) );
  AND2_X1 U14648 ( .A1(n8216), .A2(n8215), .ZN(n14653) );
  AND2_X1 U14649 ( .A1(n8213), .A2(n14654), .ZN(n14652) );
  OR2_X1 U14650 ( .A1(n8215), .A2(n8216), .ZN(n14654) );
  OR2_X1 U14651 ( .A1(n7957), .A2(n7950), .ZN(n8216) );
  OR2_X1 U14652 ( .A1(n14655), .A2(n14656), .ZN(n8215) );
  AND2_X1 U14653 ( .A1(n8233), .A2(n8232), .ZN(n14656) );
  AND2_X1 U14654 ( .A1(n8230), .A2(n14657), .ZN(n14655) );
  OR2_X1 U14655 ( .A1(n8232), .A2(n8233), .ZN(n14657) );
  OR2_X1 U14656 ( .A1(n7957), .A2(n7953), .ZN(n8233) );
  OR2_X1 U14657 ( .A1(n14658), .A2(n14659), .ZN(n8232) );
  AND2_X1 U14658 ( .A1(n8265), .A2(n7958), .ZN(n14659) );
  AND2_X1 U14659 ( .A1(n8264), .A2(n14660), .ZN(n14658) );
  OR2_X1 U14660 ( .A1(n7958), .A2(n8265), .ZN(n14660) );
  OR2_X1 U14661 ( .A1(n14661), .A2(n14662), .ZN(n8265) );
  AND2_X1 U14662 ( .A1(n8295), .A2(n8294), .ZN(n14662) );
  AND2_X1 U14663 ( .A1(n8292), .A2(n14663), .ZN(n14661) );
  OR2_X1 U14664 ( .A1(n8294), .A2(n8295), .ZN(n14663) );
  OR2_X1 U14665 ( .A1(n7957), .A2(n7960), .ZN(n8295) );
  OR2_X1 U14666 ( .A1(n14664), .A2(n14665), .ZN(n8294) );
  AND2_X1 U14667 ( .A1(n8342), .A2(n8341), .ZN(n14665) );
  AND2_X1 U14668 ( .A1(n8339), .A2(n14666), .ZN(n14664) );
  OR2_X1 U14669 ( .A1(n8341), .A2(n8342), .ZN(n14666) );
  OR2_X1 U14670 ( .A1(n7957), .A2(n7963), .ZN(n8342) );
  OR2_X1 U14671 ( .A1(n14667), .A2(n14668), .ZN(n8341) );
  AND2_X1 U14672 ( .A1(n8386), .A2(n8385), .ZN(n14668) );
  AND2_X1 U14673 ( .A1(n8383), .A2(n14669), .ZN(n14667) );
  OR2_X1 U14674 ( .A1(n8385), .A2(n8386), .ZN(n14669) );
  OR2_X1 U14675 ( .A1(n7957), .A2(n7967), .ZN(n8386) );
  OR2_X1 U14676 ( .A1(n14670), .A2(n14671), .ZN(n8385) );
  AND2_X1 U14677 ( .A1(n8441), .A2(n8440), .ZN(n14671) );
  AND2_X1 U14678 ( .A1(n8438), .A2(n14672), .ZN(n14670) );
  OR2_X1 U14679 ( .A1(n8440), .A2(n8441), .ZN(n14672) );
  OR2_X1 U14680 ( .A1(n7957), .A2(n7970), .ZN(n8441) );
  OR2_X1 U14681 ( .A1(n14673), .A2(n14674), .ZN(n8440) );
  AND2_X1 U14682 ( .A1(n8505), .A2(n8504), .ZN(n14674) );
  AND2_X1 U14683 ( .A1(n8502), .A2(n14675), .ZN(n14673) );
  OR2_X1 U14684 ( .A1(n8504), .A2(n8505), .ZN(n14675) );
  OR2_X1 U14685 ( .A1(n7957), .A2(n7974), .ZN(n8505) );
  OR2_X1 U14686 ( .A1(n14676), .A2(n14677), .ZN(n8504) );
  AND2_X1 U14687 ( .A1(n14651), .A2(n14650), .ZN(n14677) );
  AND2_X1 U14688 ( .A1(n14648), .A2(n14678), .ZN(n14676) );
  OR2_X1 U14689 ( .A1(n14650), .A2(n14651), .ZN(n14678) );
  OR2_X1 U14690 ( .A1(n7957), .A2(n7977), .ZN(n14651) );
  OR2_X1 U14691 ( .A1(n14679), .A2(n14680), .ZN(n14650) );
  AND2_X1 U14692 ( .A1(n14647), .A2(n14646), .ZN(n14680) );
  AND2_X1 U14693 ( .A1(n14644), .A2(n14681), .ZN(n14679) );
  OR2_X1 U14694 ( .A1(n14646), .A2(n14647), .ZN(n14681) );
  OR2_X1 U14695 ( .A1(n7957), .A2(n7981), .ZN(n14647) );
  OR2_X1 U14696 ( .A1(n14682), .A2(n14683), .ZN(n14646) );
  AND2_X1 U14697 ( .A1(n14643), .A2(n14642), .ZN(n14683) );
  AND2_X1 U14698 ( .A1(n14640), .A2(n14684), .ZN(n14682) );
  OR2_X1 U14699 ( .A1(n14642), .A2(n14643), .ZN(n14684) );
  OR2_X1 U14700 ( .A1(n7957), .A2(n7984), .ZN(n14643) );
  OR2_X1 U14701 ( .A1(n14685), .A2(n14686), .ZN(n14642) );
  AND2_X1 U14702 ( .A1(n14639), .A2(n14638), .ZN(n14686) );
  AND2_X1 U14703 ( .A1(n14636), .A2(n14687), .ZN(n14685) );
  OR2_X1 U14704 ( .A1(n14638), .A2(n14639), .ZN(n14687) );
  OR2_X1 U14705 ( .A1(n7957), .A2(n7988), .ZN(n14639) );
  OR2_X1 U14706 ( .A1(n14688), .A2(n14689), .ZN(n14638) );
  AND2_X1 U14707 ( .A1(n14635), .A2(n14634), .ZN(n14689) );
  AND2_X1 U14708 ( .A1(n14632), .A2(n14690), .ZN(n14688) );
  OR2_X1 U14709 ( .A1(n14634), .A2(n14635), .ZN(n14690) );
  OR2_X1 U14710 ( .A1(n7957), .A2(n7991), .ZN(n14635) );
  OR2_X1 U14711 ( .A1(n14691), .A2(n14692), .ZN(n14634) );
  AND2_X1 U14712 ( .A1(n14631), .A2(n14630), .ZN(n14692) );
  AND2_X1 U14713 ( .A1(n14628), .A2(n14693), .ZN(n14691) );
  OR2_X1 U14714 ( .A1(n14630), .A2(n14631), .ZN(n14693) );
  OR2_X1 U14715 ( .A1(n7957), .A2(n7995), .ZN(n14631) );
  OR2_X1 U14716 ( .A1(n14694), .A2(n14695), .ZN(n14630) );
  AND2_X1 U14717 ( .A1(n14627), .A2(n14626), .ZN(n14695) );
  AND2_X1 U14718 ( .A1(n14624), .A2(n14696), .ZN(n14694) );
  OR2_X1 U14719 ( .A1(n14626), .A2(n14627), .ZN(n14696) );
  OR2_X1 U14720 ( .A1(n7957), .A2(n7998), .ZN(n14627) );
  OR2_X1 U14721 ( .A1(n14697), .A2(n14698), .ZN(n14626) );
  AND2_X1 U14722 ( .A1(n14623), .A2(n14622), .ZN(n14698) );
  AND2_X1 U14723 ( .A1(n14620), .A2(n14699), .ZN(n14697) );
  OR2_X1 U14724 ( .A1(n14622), .A2(n14623), .ZN(n14699) );
  OR2_X1 U14725 ( .A1(n7957), .A2(n8002), .ZN(n14623) );
  OR2_X1 U14726 ( .A1(n14700), .A2(n14701), .ZN(n14622) );
  AND2_X1 U14727 ( .A1(n14619), .A2(n14618), .ZN(n14701) );
  AND2_X1 U14728 ( .A1(n14616), .A2(n14702), .ZN(n14700) );
  OR2_X1 U14729 ( .A1(n14618), .A2(n14619), .ZN(n14702) );
  OR2_X1 U14730 ( .A1(n7957), .A2(n8005), .ZN(n14619) );
  OR2_X1 U14731 ( .A1(n14703), .A2(n14704), .ZN(n14618) );
  AND2_X1 U14732 ( .A1(n14615), .A2(n14614), .ZN(n14704) );
  AND2_X1 U14733 ( .A1(n14612), .A2(n14705), .ZN(n14703) );
  OR2_X1 U14734 ( .A1(n14614), .A2(n14615), .ZN(n14705) );
  OR2_X1 U14735 ( .A1(n7957), .A2(n8009), .ZN(n14615) );
  OR2_X1 U14736 ( .A1(n14706), .A2(n14707), .ZN(n14614) );
  AND2_X1 U14737 ( .A1(n14611), .A2(n14610), .ZN(n14707) );
  AND2_X1 U14738 ( .A1(n14608), .A2(n14708), .ZN(n14706) );
  OR2_X1 U14739 ( .A1(n14610), .A2(n14611), .ZN(n14708) );
  OR2_X1 U14740 ( .A1(n7957), .A2(n8012), .ZN(n14611) );
  OR2_X1 U14741 ( .A1(n14709), .A2(n14710), .ZN(n14610) );
  AND2_X1 U14742 ( .A1(n14607), .A2(n14606), .ZN(n14710) );
  AND2_X1 U14743 ( .A1(n14604), .A2(n14711), .ZN(n14709) );
  OR2_X1 U14744 ( .A1(n14606), .A2(n14607), .ZN(n14711) );
  OR2_X1 U14745 ( .A1(n7957), .A2(n8016), .ZN(n14607) );
  OR2_X1 U14746 ( .A1(n14712), .A2(n14713), .ZN(n14606) );
  AND2_X1 U14747 ( .A1(n14603), .A2(n14602), .ZN(n14713) );
  AND2_X1 U14748 ( .A1(n14600), .A2(n14714), .ZN(n14712) );
  OR2_X1 U14749 ( .A1(n14602), .A2(n14603), .ZN(n14714) );
  OR2_X1 U14750 ( .A1(n7957), .A2(n8019), .ZN(n14603) );
  OR2_X1 U14751 ( .A1(n14715), .A2(n14716), .ZN(n14602) );
  AND2_X1 U14752 ( .A1(n14599), .A2(n14598), .ZN(n14716) );
  AND2_X1 U14753 ( .A1(n14596), .A2(n14717), .ZN(n14715) );
  OR2_X1 U14754 ( .A1(n14598), .A2(n14599), .ZN(n14717) );
  OR2_X1 U14755 ( .A1(n7957), .A2(n8023), .ZN(n14599) );
  OR2_X1 U14756 ( .A1(n14718), .A2(n14719), .ZN(n14598) );
  AND2_X1 U14757 ( .A1(n14595), .A2(n14594), .ZN(n14719) );
  AND2_X1 U14758 ( .A1(n14592), .A2(n14720), .ZN(n14718) );
  OR2_X1 U14759 ( .A1(n14594), .A2(n14595), .ZN(n14720) );
  OR2_X1 U14760 ( .A1(n8026), .A2(n7957), .ZN(n14595) );
  OR2_X1 U14761 ( .A1(n14721), .A2(n14722), .ZN(n14594) );
  AND2_X1 U14762 ( .A1(n14591), .A2(n14590), .ZN(n14722) );
  AND2_X1 U14763 ( .A1(n14588), .A2(n14723), .ZN(n14721) );
  OR2_X1 U14764 ( .A1(n14590), .A2(n14591), .ZN(n14723) );
  OR2_X1 U14765 ( .A1(n8030), .A2(n7957), .ZN(n14591) );
  OR2_X1 U14766 ( .A1(n14724), .A2(n14725), .ZN(n14590) );
  AND2_X1 U14767 ( .A1(n14587), .A2(n14586), .ZN(n14725) );
  AND2_X1 U14768 ( .A1(n14584), .A2(n14726), .ZN(n14724) );
  OR2_X1 U14769 ( .A1(n14586), .A2(n14587), .ZN(n14726) );
  OR2_X1 U14770 ( .A1(n8034), .A2(n7957), .ZN(n14587) );
  OR2_X1 U14771 ( .A1(n14727), .A2(n14728), .ZN(n14586) );
  AND2_X1 U14772 ( .A1(n14583), .A2(n14582), .ZN(n14728) );
  AND2_X1 U14773 ( .A1(n14580), .A2(n14729), .ZN(n14727) );
  OR2_X1 U14774 ( .A1(n14582), .A2(n14583), .ZN(n14729) );
  OR2_X1 U14775 ( .A1(n8037), .A2(n7957), .ZN(n14583) );
  OR2_X1 U14776 ( .A1(n14730), .A2(n14731), .ZN(n14582) );
  AND2_X1 U14777 ( .A1(n14579), .A2(n14578), .ZN(n14731) );
  AND2_X1 U14778 ( .A1(n14576), .A2(n14732), .ZN(n14730) );
  OR2_X1 U14779 ( .A1(n14578), .A2(n14579), .ZN(n14732) );
  OR2_X1 U14780 ( .A1(n8041), .A2(n7957), .ZN(n14579) );
  OR2_X1 U14781 ( .A1(n14733), .A2(n14734), .ZN(n14578) );
  AND2_X1 U14782 ( .A1(n14572), .A2(n14575), .ZN(n14734) );
  AND2_X1 U14783 ( .A1(n14735), .A2(n14574), .ZN(n14733) );
  OR2_X1 U14784 ( .A1(n14736), .A2(n14737), .ZN(n14574) );
  AND2_X1 U14785 ( .A1(n14571), .A2(n14570), .ZN(n14737) );
  AND2_X1 U14786 ( .A1(n14568), .A2(n14738), .ZN(n14736) );
  OR2_X1 U14787 ( .A1(n14570), .A2(n14571), .ZN(n14738) );
  OR2_X1 U14788 ( .A1(n8048), .A2(n7957), .ZN(n14571) );
  OR2_X1 U14789 ( .A1(n14739), .A2(n14740), .ZN(n14570) );
  AND2_X1 U14790 ( .A1(n14564), .A2(n14741), .ZN(n14740) );
  AND2_X1 U14791 ( .A1(n14742), .A2(n14743), .ZN(n14739) );
  OR2_X1 U14792 ( .A1(n14741), .A2(n14564), .ZN(n14743) );
  OR2_X1 U14793 ( .A1(n8051), .A2(n7957), .ZN(n14564) );
  INV_X1 U14794 ( .A(n14567), .ZN(n14741) );
  AND3_X1 U14795 ( .A1(n8904), .A2(b_2_), .A3(b_1_), .ZN(n14567) );
  INV_X1 U14796 ( .A(n14566), .ZN(n14742) );
  OR2_X1 U14797 ( .A1(n14744), .A2(n14745), .ZN(n14566) );
  AND2_X1 U14798 ( .A1(b_1_), .A2(n14746), .ZN(n14745) );
  OR2_X1 U14799 ( .A1(n14747), .A2(n7490), .ZN(n14746) );
  AND2_X1 U14800 ( .A1(n14748), .A2(a_30_), .ZN(n7490) );
  INV_X1 U14801 ( .A(a_31_), .ZN(n14748) );
  AND2_X1 U14802 ( .A1(a_30_), .A2(n7951), .ZN(n14747) );
  AND2_X1 U14803 ( .A1(b_0_), .A2(n14749), .ZN(n14744) );
  OR2_X1 U14804 ( .A1(n14750), .A2(n7493), .ZN(n14749) );
  AND2_X1 U14805 ( .A1(n14751), .A2(a_31_), .ZN(n7493) );
  AND2_X1 U14806 ( .A1(a_31_), .A2(n7930), .ZN(n14750) );
  XOR2_X1 U14807 ( .A(n14752), .B(n14753), .Z(n14568) );
  OR2_X1 U14808 ( .A1(n14754), .A2(n14755), .ZN(n14752) );
  AND2_X1 U14809 ( .A1(n14756), .A2(n14757), .ZN(n14754) );
  INV_X1 U14810 ( .A(n14758), .ZN(n14757) );
  OR2_X1 U14811 ( .A1(n14751), .A2(n7951), .ZN(n14756) );
  INV_X1 U14812 ( .A(a_30_), .ZN(n14751) );
  OR2_X1 U14813 ( .A1(n14575), .A2(n14572), .ZN(n14735) );
  XNOR2_X1 U14814 ( .A(n14759), .B(n14760), .ZN(n14572) );
  XNOR2_X1 U14815 ( .A(n14761), .B(n14762), .ZN(n14760) );
  OR2_X1 U14816 ( .A1(n8044), .A2(n7957), .ZN(n14575) );
  INV_X1 U14817 ( .A(b_2_), .ZN(n7957) );
  XNOR2_X1 U14818 ( .A(n14763), .B(n14764), .ZN(n14576) );
  XNOR2_X1 U14819 ( .A(n14765), .B(n14766), .ZN(n14763) );
  XNOR2_X1 U14820 ( .A(n14767), .B(n14768), .ZN(n14580) );
  XNOR2_X1 U14821 ( .A(n14769), .B(n14770), .ZN(n14767) );
  XNOR2_X1 U14822 ( .A(n14771), .B(n14772), .ZN(n14584) );
  XNOR2_X1 U14823 ( .A(n14773), .B(n14774), .ZN(n14771) );
  XNOR2_X1 U14824 ( .A(n14775), .B(n14776), .ZN(n14588) );
  XNOR2_X1 U14825 ( .A(n14777), .B(n14778), .ZN(n14775) );
  XNOR2_X1 U14826 ( .A(n14779), .B(n14780), .ZN(n14592) );
  XNOR2_X1 U14827 ( .A(n14781), .B(n14782), .ZN(n14779) );
  XNOR2_X1 U14828 ( .A(n14783), .B(n14784), .ZN(n14596) );
  XNOR2_X1 U14829 ( .A(n14785), .B(n14786), .ZN(n14783) );
  XNOR2_X1 U14830 ( .A(n14787), .B(n14788), .ZN(n14600) );
  XNOR2_X1 U14831 ( .A(n14789), .B(n14790), .ZN(n14787) );
  XNOR2_X1 U14832 ( .A(n14791), .B(n14792), .ZN(n14604) );
  XNOR2_X1 U14833 ( .A(n14793), .B(n14794), .ZN(n14791) );
  XNOR2_X1 U14834 ( .A(n14795), .B(n14796), .ZN(n14608) );
  XNOR2_X1 U14835 ( .A(n14797), .B(n14798), .ZN(n14795) );
  XNOR2_X1 U14836 ( .A(n14799), .B(n14800), .ZN(n14612) );
  XNOR2_X1 U14837 ( .A(n14801), .B(n14802), .ZN(n14799) );
  XNOR2_X1 U14838 ( .A(n14803), .B(n14804), .ZN(n14616) );
  XNOR2_X1 U14839 ( .A(n14805), .B(n14806), .ZN(n14803) );
  XNOR2_X1 U14840 ( .A(n14807), .B(n14808), .ZN(n14620) );
  XNOR2_X1 U14841 ( .A(n14809), .B(n14810), .ZN(n14807) );
  XNOR2_X1 U14842 ( .A(n14811), .B(n14812), .ZN(n14624) );
  XNOR2_X1 U14843 ( .A(n14813), .B(n14814), .ZN(n14811) );
  XNOR2_X1 U14844 ( .A(n14815), .B(n14816), .ZN(n14628) );
  XNOR2_X1 U14845 ( .A(n14817), .B(n14818), .ZN(n14815) );
  XNOR2_X1 U14846 ( .A(n14819), .B(n14820), .ZN(n14632) );
  XNOR2_X1 U14847 ( .A(n14821), .B(n14822), .ZN(n14819) );
  XNOR2_X1 U14848 ( .A(n14823), .B(n14824), .ZN(n14636) );
  XNOR2_X1 U14849 ( .A(n14825), .B(n14826), .ZN(n14823) );
  XNOR2_X1 U14850 ( .A(n14827), .B(n14828), .ZN(n14640) );
  XNOR2_X1 U14851 ( .A(n14829), .B(n14830), .ZN(n14827) );
  XNOR2_X1 U14852 ( .A(n14831), .B(n14832), .ZN(n14644) );
  XNOR2_X1 U14853 ( .A(n14833), .B(n14834), .ZN(n14831) );
  XNOR2_X1 U14854 ( .A(n14835), .B(n14836), .ZN(n14648) );
  XNOR2_X1 U14855 ( .A(n14837), .B(n14838), .ZN(n14835) );
  XOR2_X1 U14856 ( .A(n14839), .B(n14840), .Z(n8502) );
  XOR2_X1 U14857 ( .A(n14841), .B(n14842), .Z(n14840) );
  XOR2_X1 U14858 ( .A(n14843), .B(n14844), .Z(n8438) );
  XOR2_X1 U14859 ( .A(n14845), .B(n14846), .Z(n14844) );
  XOR2_X1 U14860 ( .A(n14847), .B(n14848), .Z(n8383) );
  XOR2_X1 U14861 ( .A(n14849), .B(n14850), .Z(n14848) );
  XOR2_X1 U14862 ( .A(n14851), .B(n14852), .Z(n8339) );
  XOR2_X1 U14863 ( .A(n14853), .B(n14854), .Z(n14852) );
  XOR2_X1 U14864 ( .A(n14855), .B(n14856), .Z(n8292) );
  XOR2_X1 U14865 ( .A(n14857), .B(n14858), .Z(n14856) );
  INV_X1 U14866 ( .A(n7922), .ZN(n7958) );
  AND2_X1 U14867 ( .A1(b_2_), .A2(a_2_), .ZN(n7922) );
  XOR2_X1 U14868 ( .A(n14859), .B(n14860), .Z(n8264) );
  XOR2_X1 U14869 ( .A(n14861), .B(n14862), .Z(n14860) );
  XOR2_X1 U14870 ( .A(n14863), .B(n14864), .Z(n8230) );
  XOR2_X1 U14871 ( .A(n14865), .B(n14866), .Z(n14864) );
  XOR2_X1 U14872 ( .A(n14867), .B(n14868), .Z(n8213) );
  XNOR2_X1 U14873 ( .A(n14869), .B(n7934), .ZN(n14868) );
  XOR2_X1 U14874 ( .A(n14870), .B(n8196), .Z(n8128) );
  INV_X1 U14875 ( .A(n14871), .ZN(n8196) );
  OR2_X1 U14876 ( .A1(n14872), .A2(n14873), .ZN(n14871) );
  AND2_X1 U14877 ( .A1(n14874), .A2(n14875), .ZN(n14873) );
  AND2_X1 U14878 ( .A1(n14876), .A2(n14877), .ZN(n14872) );
  OR2_X1 U14879 ( .A1(n14875), .A2(n14874), .ZN(n14876) );
  AND2_X1 U14880 ( .A1(b_0_), .A2(a_0_), .ZN(n14870) );
  XOR2_X1 U14881 ( .A(n14878), .B(n14874), .Z(n8130) );
  OR2_X1 U14882 ( .A1(n14879), .A2(n14880), .ZN(n14874) );
  AND2_X1 U14883 ( .A1(n14867), .A2(n14869), .ZN(n14880) );
  AND2_X1 U14884 ( .A1(n14881), .A2(n7954), .ZN(n14879) );
  INV_X1 U14885 ( .A(n7934), .ZN(n7954) );
  AND2_X1 U14886 ( .A1(b_1_), .A2(a_1_), .ZN(n7934) );
  OR2_X1 U14887 ( .A1(n14869), .A2(n14867), .ZN(n14881) );
  OR2_X1 U14888 ( .A1(n7951), .A2(n7956), .ZN(n14867) );
  OR2_X1 U14889 ( .A1(n14882), .A2(n14883), .ZN(n14869) );
  AND2_X1 U14890 ( .A1(n14863), .A2(n14865), .ZN(n14883) );
  AND2_X1 U14891 ( .A1(n14884), .A2(n14866), .ZN(n14882) );
  OR2_X1 U14892 ( .A1(n7951), .A2(n7960), .ZN(n14866) );
  OR2_X1 U14893 ( .A1(n14865), .A2(n14863), .ZN(n14884) );
  OR2_X1 U14894 ( .A1(n7930), .A2(n7956), .ZN(n14863) );
  INV_X1 U14895 ( .A(a_2_), .ZN(n7956) );
  OR2_X1 U14896 ( .A1(n14885), .A2(n14886), .ZN(n14865) );
  AND2_X1 U14897 ( .A1(n14859), .A2(n14861), .ZN(n14886) );
  AND2_X1 U14898 ( .A1(n14887), .A2(n14862), .ZN(n14885) );
  OR2_X1 U14899 ( .A1(n7951), .A2(n7963), .ZN(n14862) );
  OR2_X1 U14900 ( .A1(n14861), .A2(n14859), .ZN(n14887) );
  OR2_X1 U14901 ( .A1(n7930), .A2(n7960), .ZN(n14859) );
  INV_X1 U14902 ( .A(a_3_), .ZN(n7960) );
  OR2_X1 U14903 ( .A1(n14888), .A2(n14889), .ZN(n14861) );
  AND2_X1 U14904 ( .A1(n14855), .A2(n14857), .ZN(n14889) );
  AND2_X1 U14905 ( .A1(n14890), .A2(n14858), .ZN(n14888) );
  OR2_X1 U14906 ( .A1(n7951), .A2(n7967), .ZN(n14858) );
  OR2_X1 U14907 ( .A1(n14857), .A2(n14855), .ZN(n14890) );
  OR2_X1 U14908 ( .A1(n7930), .A2(n7963), .ZN(n14855) );
  INV_X1 U14909 ( .A(a_4_), .ZN(n7963) );
  OR2_X1 U14910 ( .A1(n14891), .A2(n14892), .ZN(n14857) );
  AND2_X1 U14911 ( .A1(n14851), .A2(n14853), .ZN(n14892) );
  AND2_X1 U14912 ( .A1(n14893), .A2(n14854), .ZN(n14891) );
  OR2_X1 U14913 ( .A1(n7951), .A2(n7970), .ZN(n14854) );
  OR2_X1 U14914 ( .A1(n14853), .A2(n14851), .ZN(n14893) );
  OR2_X1 U14915 ( .A1(n7930), .A2(n7967), .ZN(n14851) );
  INV_X1 U14916 ( .A(a_5_), .ZN(n7967) );
  OR2_X1 U14917 ( .A1(n14894), .A2(n14895), .ZN(n14853) );
  AND2_X1 U14918 ( .A1(n14847), .A2(n14849), .ZN(n14895) );
  AND2_X1 U14919 ( .A1(n14896), .A2(n14850), .ZN(n14894) );
  OR2_X1 U14920 ( .A1(n7951), .A2(n7974), .ZN(n14850) );
  OR2_X1 U14921 ( .A1(n14849), .A2(n14847), .ZN(n14896) );
  OR2_X1 U14922 ( .A1(n7930), .A2(n7970), .ZN(n14847) );
  INV_X1 U14923 ( .A(a_6_), .ZN(n7970) );
  OR2_X1 U14924 ( .A1(n14897), .A2(n14898), .ZN(n14849) );
  AND2_X1 U14925 ( .A1(n14843), .A2(n14845), .ZN(n14898) );
  AND2_X1 U14926 ( .A1(n14899), .A2(n14846), .ZN(n14897) );
  OR2_X1 U14927 ( .A1(n7951), .A2(n7977), .ZN(n14846) );
  OR2_X1 U14928 ( .A1(n14845), .A2(n14843), .ZN(n14899) );
  OR2_X1 U14929 ( .A1(n7930), .A2(n7974), .ZN(n14843) );
  INV_X1 U14930 ( .A(a_7_), .ZN(n7974) );
  OR2_X1 U14931 ( .A1(n14900), .A2(n14901), .ZN(n14845) );
  AND2_X1 U14932 ( .A1(n14839), .A2(n14841), .ZN(n14901) );
  AND2_X1 U14933 ( .A1(n14902), .A2(n14842), .ZN(n14900) );
  OR2_X1 U14934 ( .A1(n7951), .A2(n7981), .ZN(n14842) );
  OR2_X1 U14935 ( .A1(n14841), .A2(n14839), .ZN(n14902) );
  OR2_X1 U14936 ( .A1(n7930), .A2(n7977), .ZN(n14839) );
  INV_X1 U14937 ( .A(a_8_), .ZN(n7977) );
  OR2_X1 U14938 ( .A1(n14903), .A2(n14904), .ZN(n14841) );
  AND2_X1 U14939 ( .A1(n14836), .A2(n14838), .ZN(n14904) );
  AND2_X1 U14940 ( .A1(n14905), .A2(n14837), .ZN(n14903) );
  OR2_X1 U14941 ( .A1(n7951), .A2(n7984), .ZN(n14837) );
  OR2_X1 U14942 ( .A1(n14838), .A2(n14836), .ZN(n14905) );
  OR2_X1 U14943 ( .A1(n7930), .A2(n7981), .ZN(n14836) );
  INV_X1 U14944 ( .A(a_9_), .ZN(n7981) );
  OR2_X1 U14945 ( .A1(n14906), .A2(n14907), .ZN(n14838) );
  AND2_X1 U14946 ( .A1(n14832), .A2(n14834), .ZN(n14907) );
  AND2_X1 U14947 ( .A1(n14908), .A2(n14833), .ZN(n14906) );
  OR2_X1 U14948 ( .A1(n7951), .A2(n7988), .ZN(n14833) );
  OR2_X1 U14949 ( .A1(n14834), .A2(n14832), .ZN(n14908) );
  OR2_X1 U14950 ( .A1(n7930), .A2(n7984), .ZN(n14832) );
  INV_X1 U14951 ( .A(a_10_), .ZN(n7984) );
  OR2_X1 U14952 ( .A1(n14909), .A2(n14910), .ZN(n14834) );
  AND2_X1 U14953 ( .A1(n14828), .A2(n14830), .ZN(n14910) );
  AND2_X1 U14954 ( .A1(n14911), .A2(n14829), .ZN(n14909) );
  OR2_X1 U14955 ( .A1(n7951), .A2(n7991), .ZN(n14829) );
  OR2_X1 U14956 ( .A1(n14830), .A2(n14828), .ZN(n14911) );
  OR2_X1 U14957 ( .A1(n7930), .A2(n7988), .ZN(n14828) );
  INV_X1 U14958 ( .A(a_11_), .ZN(n7988) );
  OR2_X1 U14959 ( .A1(n14912), .A2(n14913), .ZN(n14830) );
  AND2_X1 U14960 ( .A1(n14824), .A2(n14826), .ZN(n14913) );
  AND2_X1 U14961 ( .A1(n14914), .A2(n14825), .ZN(n14912) );
  OR2_X1 U14962 ( .A1(n7951), .A2(n7995), .ZN(n14825) );
  OR2_X1 U14963 ( .A1(n14826), .A2(n14824), .ZN(n14914) );
  OR2_X1 U14964 ( .A1(n7930), .A2(n7991), .ZN(n14824) );
  INV_X1 U14965 ( .A(a_12_), .ZN(n7991) );
  OR2_X1 U14966 ( .A1(n14915), .A2(n14916), .ZN(n14826) );
  AND2_X1 U14967 ( .A1(n14820), .A2(n14822), .ZN(n14916) );
  AND2_X1 U14968 ( .A1(n14917), .A2(n14821), .ZN(n14915) );
  OR2_X1 U14969 ( .A1(n7951), .A2(n7998), .ZN(n14821) );
  OR2_X1 U14970 ( .A1(n14822), .A2(n14820), .ZN(n14917) );
  OR2_X1 U14971 ( .A1(n7930), .A2(n7995), .ZN(n14820) );
  INV_X1 U14972 ( .A(a_13_), .ZN(n7995) );
  OR2_X1 U14973 ( .A1(n14918), .A2(n14919), .ZN(n14822) );
  AND2_X1 U14974 ( .A1(n14816), .A2(n14818), .ZN(n14919) );
  AND2_X1 U14975 ( .A1(n14920), .A2(n14817), .ZN(n14918) );
  OR2_X1 U14976 ( .A1(n7951), .A2(n8002), .ZN(n14817) );
  OR2_X1 U14977 ( .A1(n14818), .A2(n14816), .ZN(n14920) );
  OR2_X1 U14978 ( .A1(n7930), .A2(n7998), .ZN(n14816) );
  INV_X1 U14979 ( .A(a_14_), .ZN(n7998) );
  OR2_X1 U14980 ( .A1(n14921), .A2(n14922), .ZN(n14818) );
  AND2_X1 U14981 ( .A1(n14812), .A2(n14814), .ZN(n14922) );
  AND2_X1 U14982 ( .A1(n14923), .A2(n14813), .ZN(n14921) );
  OR2_X1 U14983 ( .A1(n7951), .A2(n8005), .ZN(n14813) );
  OR2_X1 U14984 ( .A1(n14814), .A2(n14812), .ZN(n14923) );
  OR2_X1 U14985 ( .A1(n7930), .A2(n8002), .ZN(n14812) );
  INV_X1 U14986 ( .A(a_15_), .ZN(n8002) );
  OR2_X1 U14987 ( .A1(n14924), .A2(n14925), .ZN(n14814) );
  AND2_X1 U14988 ( .A1(n14808), .A2(n14810), .ZN(n14925) );
  AND2_X1 U14989 ( .A1(n14926), .A2(n14809), .ZN(n14924) );
  OR2_X1 U14990 ( .A1(n7951), .A2(n8009), .ZN(n14809) );
  OR2_X1 U14991 ( .A1(n14810), .A2(n14808), .ZN(n14926) );
  OR2_X1 U14992 ( .A1(n7930), .A2(n8005), .ZN(n14808) );
  INV_X1 U14993 ( .A(a_16_), .ZN(n8005) );
  OR2_X1 U14994 ( .A1(n14927), .A2(n14928), .ZN(n14810) );
  AND2_X1 U14995 ( .A1(n14804), .A2(n14806), .ZN(n14928) );
  AND2_X1 U14996 ( .A1(n14929), .A2(n14805), .ZN(n14927) );
  OR2_X1 U14997 ( .A1(n7951), .A2(n8012), .ZN(n14805) );
  OR2_X1 U14998 ( .A1(n14806), .A2(n14804), .ZN(n14929) );
  OR2_X1 U14999 ( .A1(n7930), .A2(n8009), .ZN(n14804) );
  INV_X1 U15000 ( .A(a_17_), .ZN(n8009) );
  OR2_X1 U15001 ( .A1(n14930), .A2(n14931), .ZN(n14806) );
  AND2_X1 U15002 ( .A1(n14800), .A2(n14802), .ZN(n14931) );
  AND2_X1 U15003 ( .A1(n14932), .A2(n14801), .ZN(n14930) );
  OR2_X1 U15004 ( .A1(n7951), .A2(n8016), .ZN(n14801) );
  OR2_X1 U15005 ( .A1(n14802), .A2(n14800), .ZN(n14932) );
  OR2_X1 U15006 ( .A1(n7930), .A2(n8012), .ZN(n14800) );
  INV_X1 U15007 ( .A(a_18_), .ZN(n8012) );
  OR2_X1 U15008 ( .A1(n14933), .A2(n14934), .ZN(n14802) );
  AND2_X1 U15009 ( .A1(n14796), .A2(n14798), .ZN(n14934) );
  AND2_X1 U15010 ( .A1(n14935), .A2(n14797), .ZN(n14933) );
  OR2_X1 U15011 ( .A1(n8019), .A2(n7951), .ZN(n14797) );
  OR2_X1 U15012 ( .A1(n14798), .A2(n14796), .ZN(n14935) );
  OR2_X1 U15013 ( .A1(n7930), .A2(n8016), .ZN(n14796) );
  INV_X1 U15014 ( .A(a_19_), .ZN(n8016) );
  OR2_X1 U15015 ( .A1(n14936), .A2(n14937), .ZN(n14798) );
  AND2_X1 U15016 ( .A1(n14792), .A2(n14794), .ZN(n14937) );
  AND2_X1 U15017 ( .A1(n14938), .A2(n14793), .ZN(n14936) );
  OR2_X1 U15018 ( .A1(n8023), .A2(n7951), .ZN(n14793) );
  OR2_X1 U15019 ( .A1(n14794), .A2(n14792), .ZN(n14938) );
  OR2_X1 U15020 ( .A1(n7930), .A2(n8019), .ZN(n14792) );
  INV_X1 U15021 ( .A(a_20_), .ZN(n8019) );
  OR2_X1 U15022 ( .A1(n14939), .A2(n14940), .ZN(n14794) );
  AND2_X1 U15023 ( .A1(n14788), .A2(n14790), .ZN(n14940) );
  AND2_X1 U15024 ( .A1(n14941), .A2(n14789), .ZN(n14939) );
  OR2_X1 U15025 ( .A1(n8026), .A2(n7951), .ZN(n14789) );
  OR2_X1 U15026 ( .A1(n14790), .A2(n14788), .ZN(n14941) );
  OR2_X1 U15027 ( .A1(n8023), .A2(n7930), .ZN(n14788) );
  INV_X1 U15028 ( .A(a_21_), .ZN(n8023) );
  OR2_X1 U15029 ( .A1(n14942), .A2(n14943), .ZN(n14790) );
  AND2_X1 U15030 ( .A1(n14784), .A2(n14786), .ZN(n14943) );
  AND2_X1 U15031 ( .A1(n14944), .A2(n14785), .ZN(n14942) );
  OR2_X1 U15032 ( .A1(n8030), .A2(n7951), .ZN(n14785) );
  OR2_X1 U15033 ( .A1(n14786), .A2(n14784), .ZN(n14944) );
  OR2_X1 U15034 ( .A1(n8026), .A2(n7930), .ZN(n14784) );
  INV_X1 U15035 ( .A(a_22_), .ZN(n8026) );
  OR2_X1 U15036 ( .A1(n14945), .A2(n14946), .ZN(n14786) );
  AND2_X1 U15037 ( .A1(n14780), .A2(n14782), .ZN(n14946) );
  AND2_X1 U15038 ( .A1(n14947), .A2(n14781), .ZN(n14945) );
  OR2_X1 U15039 ( .A1(n8034), .A2(n7951), .ZN(n14781) );
  OR2_X1 U15040 ( .A1(n14782), .A2(n14780), .ZN(n14947) );
  OR2_X1 U15041 ( .A1(n8030), .A2(n7930), .ZN(n14780) );
  INV_X1 U15042 ( .A(a_23_), .ZN(n8030) );
  OR2_X1 U15043 ( .A1(n14948), .A2(n14949), .ZN(n14782) );
  AND2_X1 U15044 ( .A1(n14776), .A2(n14778), .ZN(n14949) );
  AND2_X1 U15045 ( .A1(n14950), .A2(n14777), .ZN(n14948) );
  OR2_X1 U15046 ( .A1(n8037), .A2(n7951), .ZN(n14777) );
  OR2_X1 U15047 ( .A1(n14778), .A2(n14776), .ZN(n14950) );
  OR2_X1 U15048 ( .A1(n8034), .A2(n7930), .ZN(n14776) );
  INV_X1 U15049 ( .A(a_24_), .ZN(n8034) );
  OR2_X1 U15050 ( .A1(n14951), .A2(n14952), .ZN(n14778) );
  AND2_X1 U15051 ( .A1(n14772), .A2(n14774), .ZN(n14952) );
  AND2_X1 U15052 ( .A1(n14953), .A2(n14773), .ZN(n14951) );
  OR2_X1 U15053 ( .A1(n8041), .A2(n7951), .ZN(n14773) );
  OR2_X1 U15054 ( .A1(n14774), .A2(n14772), .ZN(n14953) );
  OR2_X1 U15055 ( .A1(n8037), .A2(n7930), .ZN(n14772) );
  INV_X1 U15056 ( .A(a_25_), .ZN(n8037) );
  OR2_X1 U15057 ( .A1(n14954), .A2(n14955), .ZN(n14774) );
  AND2_X1 U15058 ( .A1(n14768), .A2(n14770), .ZN(n14955) );
  AND2_X1 U15059 ( .A1(n14956), .A2(n14769), .ZN(n14954) );
  OR2_X1 U15060 ( .A1(n8044), .A2(n7951), .ZN(n14769) );
  OR2_X1 U15061 ( .A1(n14770), .A2(n14768), .ZN(n14956) );
  OR2_X1 U15062 ( .A1(n8041), .A2(n7930), .ZN(n14768) );
  INV_X1 U15063 ( .A(a_26_), .ZN(n8041) );
  OR2_X1 U15064 ( .A1(n14957), .A2(n14958), .ZN(n14770) );
  AND2_X1 U15065 ( .A1(n14764), .A2(n14766), .ZN(n14958) );
  AND2_X1 U15066 ( .A1(n14959), .A2(n14765), .ZN(n14957) );
  OR2_X1 U15067 ( .A1(n8048), .A2(n7951), .ZN(n14765) );
  OR2_X1 U15068 ( .A1(n14766), .A2(n14764), .ZN(n14959) );
  OR2_X1 U15069 ( .A1(n8044), .A2(n7930), .ZN(n14764) );
  INV_X1 U15070 ( .A(a_27_), .ZN(n8044) );
  OR2_X1 U15071 ( .A1(n14960), .A2(n14961), .ZN(n14766) );
  AND2_X1 U15072 ( .A1(n14759), .A2(n14762), .ZN(n14961) );
  AND2_X1 U15073 ( .A1(n14761), .A2(n14962), .ZN(n14960) );
  OR2_X1 U15074 ( .A1(n14762), .A2(n14759), .ZN(n14962) );
  OR2_X1 U15075 ( .A1(n8048), .A2(n7930), .ZN(n14759) );
  INV_X1 U15076 ( .A(a_28_), .ZN(n8048) );
  OR2_X1 U15077 ( .A1(n8051), .A2(n7951), .ZN(n14762) );
  INV_X1 U15078 ( .A(a_29_), .ZN(n8051) );
  INV_X1 U15079 ( .A(n14963), .ZN(n14761) );
  OR2_X1 U15080 ( .A1(n14755), .A2(n14753), .ZN(n14963) );
  AND3_X1 U15081 ( .A1(n8904), .A2(b_1_), .A3(b_0_), .ZN(n14753) );
  AND2_X1 U15082 ( .A1(a_30_), .A2(a_31_), .ZN(n8904) );
  AND3_X1 U15083 ( .A1(a_30_), .A2(b_0_), .A3(n14758), .ZN(n14755) );
  AND2_X1 U15084 ( .A1(a_29_), .A2(b_1_), .ZN(n14758) );
  XNOR2_X1 U15085 ( .A(n14875), .B(n14877), .ZN(n14878) );
  OR2_X1 U15086 ( .A1(n7930), .A2(n7950), .ZN(n14877) );
  INV_X1 U15087 ( .A(a_0_), .ZN(n7950) );
  INV_X1 U15088 ( .A(b_1_), .ZN(n7930) );
  OR2_X1 U15089 ( .A1(n7951), .A2(n7953), .ZN(n14875) );
  INV_X1 U15090 ( .A(a_1_), .ZN(n7953) );
  INV_X1 U15091 ( .A(b_0_), .ZN(n7951) );
endmodule

