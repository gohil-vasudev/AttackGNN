module add_mul_combine_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_mul_0_, 
        Result_mul_1_, Result_mul_2_, Result_mul_3_, Result_mul_4_, 
        Result_mul_5_, Result_mul_6_, Result_mul_7_, Result_mul_8_, 
        Result_mul_9_, Result_mul_10_, Result_mul_11_, Result_mul_12_, 
        Result_mul_13_, Result_mul_14_, Result_mul_15_, Result_add_0_, 
        Result_add_1_, Result_add_2_, Result_add_3_, Result_add_4_, 
        Result_add_5_, Result_add_6_, Result_add_7_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_;
  wire   n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884;

  XOR2_X1 U439 ( .A(n415), .B(n416), .Z(Result_mul_9_) );
  XOR2_X1 U440 ( .A(n417), .B(n418), .Z(n416) );
  NOR2_X1 U441 ( .A1(n419), .A2(n420), .ZN(n418) );
  XOR2_X1 U442 ( .A(n421), .B(n422), .Z(Result_mul_8_) );
  XOR2_X1 U443 ( .A(n423), .B(n424), .Z(n421) );
  XOR2_X1 U444 ( .A(n425), .B(n426), .Z(Result_mul_7_) );
  NOR2_X1 U445 ( .A1(n427), .A2(n428), .ZN(Result_mul_6_) );
  NOR2_X1 U446 ( .A1(n429), .A2(n430), .ZN(n428) );
  XOR2_X1 U447 ( .A(n427), .B(n431), .Z(Result_mul_5_) );
  NOR2_X1 U448 ( .A1(n432), .A2(n433), .ZN(n431) );
  NOR2_X1 U449 ( .A1(n434), .A2(n435), .ZN(n432) );
  XOR2_X1 U450 ( .A(n436), .B(n437), .Z(Result_mul_4_) );
  XNOR2_X1 U451 ( .A(n438), .B(n439), .ZN(Result_mul_3_) );
  NAND2_X1 U452 ( .A1(n440), .A2(n441), .ZN(n439) );
  XNOR2_X1 U453 ( .A(n442), .B(n443), .ZN(Result_mul_2_) );
  NAND2_X1 U454 ( .A1(n444), .A2(n445), .ZN(n442) );
  XOR2_X1 U455 ( .A(n446), .B(n447), .Z(Result_mul_1_) );
  NAND2_X1 U456 ( .A1(n448), .A2(n449), .ZN(n446) );
  XOR2_X1 U457 ( .A(n450), .B(n451), .Z(Result_mul_14_) );
  NAND2_X1 U458 ( .A1(b_7_), .A2(a_6_), .ZN(n451) );
  XNOR2_X1 U459 ( .A(n452), .B(n453), .ZN(Result_mul_13_) );
  XNOR2_X1 U460 ( .A(n454), .B(n455), .ZN(n453) );
  NAND2_X1 U461 ( .A1(b_7_), .A2(a_5_), .ZN(n454) );
  XNOR2_X1 U462 ( .A(n456), .B(n457), .ZN(Result_mul_12_) );
  NAND2_X1 U463 ( .A1(n458), .A2(n459), .ZN(n456) );
  XOR2_X1 U464 ( .A(n460), .B(n461), .Z(Result_mul_11_) );
  XNOR2_X1 U465 ( .A(n462), .B(n463), .ZN(n461) );
  NAND2_X1 U466 ( .A1(b_7_), .A2(a_3_), .ZN(n462) );
  XOR2_X1 U467 ( .A(n464), .B(n465), .Z(Result_mul_10_) );
  XOR2_X1 U468 ( .A(n466), .B(n467), .Z(n465) );
  NAND2_X1 U469 ( .A1(n468), .A2(n469), .ZN(Result_mul_0_) );
  NAND2_X1 U470 ( .A1(a_0_), .A2(n470), .ZN(n469) );
  NOR2_X1 U471 ( .A1(n471), .A2(n472), .ZN(n468) );
  NOR2_X1 U472 ( .A1(n447), .A2(n473), .ZN(n472) );
  INV_X1 U473 ( .A(n449), .ZN(n473) );
  NAND2_X1 U474 ( .A1(n474), .A2(n475), .ZN(n449) );
  OR2_X1 U475 ( .A1(n476), .A2(n477), .ZN(n475) );
  XNOR2_X1 U476 ( .A(n478), .B(n470), .ZN(n474) );
  AND2_X1 U477 ( .A1(n444), .A2(n479), .ZN(n447) );
  NAND2_X1 U478 ( .A1(n445), .A2(n443), .ZN(n479) );
  NAND2_X1 U479 ( .A1(n440), .A2(n480), .ZN(n443) );
  NAND2_X1 U480 ( .A1(n438), .A2(n441), .ZN(n480) );
  NAND2_X1 U481 ( .A1(n481), .A2(n482), .ZN(n441) );
  NAND2_X1 U482 ( .A1(n483), .A2(n484), .ZN(n482) );
  AND2_X1 U483 ( .A1(n437), .A2(n436), .ZN(n438) );
  NAND2_X1 U484 ( .A1(n485), .A2(n486), .ZN(n436) );
  NAND2_X1 U485 ( .A1(n427), .A2(n434), .ZN(n486) );
  AND2_X1 U486 ( .A1(n429), .A2(n430), .ZN(n427) );
  XOR2_X1 U487 ( .A(n487), .B(n488), .Z(n430) );
  NOR2_X1 U488 ( .A1(n426), .A2(n425), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n489), .B(n490), .ZN(n425) );
  NOR2_X1 U490 ( .A1(n491), .A2(n492), .ZN(n490) );
  NOR2_X1 U491 ( .A1(n493), .A2(n494), .ZN(n491) );
  NOR2_X1 U492 ( .A1(n495), .A2(n496), .ZN(n493) );
  AND2_X1 U493 ( .A1(n497), .A2(n498), .ZN(n426) );
  NAND2_X1 U494 ( .A1(n424), .A2(n499), .ZN(n498) );
  OR2_X1 U495 ( .A1(n422), .A2(n423), .ZN(n499) );
  NOR2_X1 U496 ( .A1(n496), .A2(n419), .ZN(n424) );
  NAND2_X1 U497 ( .A1(n422), .A2(n423), .ZN(n497) );
  NAND2_X1 U498 ( .A1(n500), .A2(n501), .ZN(n423) );
  NAND2_X1 U499 ( .A1(n502), .A2(a_1_), .ZN(n501) );
  NOR2_X1 U500 ( .A1(n503), .A2(n419), .ZN(n502) );
  NOR2_X1 U501 ( .A1(n415), .A2(n417), .ZN(n503) );
  NAND2_X1 U502 ( .A1(n415), .A2(n417), .ZN(n500) );
  NAND2_X1 U503 ( .A1(n504), .A2(n505), .ZN(n417) );
  NAND2_X1 U504 ( .A1(n467), .A2(n506), .ZN(n505) );
  NAND2_X1 U505 ( .A1(n466), .A2(n464), .ZN(n506) );
  NOR2_X1 U506 ( .A1(n419), .A2(n507), .ZN(n467) );
  OR2_X1 U507 ( .A1(n464), .A2(n466), .ZN(n504) );
  AND2_X1 U508 ( .A1(n508), .A2(n509), .ZN(n466) );
  NAND2_X1 U509 ( .A1(n510), .A2(b_7_), .ZN(n509) );
  NOR2_X1 U510 ( .A1(n511), .A2(n512), .ZN(n510) );
  NOR2_X1 U511 ( .A1(n460), .A2(n463), .ZN(n511) );
  NAND2_X1 U512 ( .A1(n460), .A2(n463), .ZN(n508) );
  NAND2_X1 U513 ( .A1(n458), .A2(n513), .ZN(n463) );
  NAND2_X1 U514 ( .A1(n457), .A2(n459), .ZN(n513) );
  NAND2_X1 U515 ( .A1(n514), .A2(n515), .ZN(n459) );
  NAND2_X1 U516 ( .A1(b_7_), .A2(a_4_), .ZN(n515) );
  INV_X1 U517 ( .A(n516), .ZN(n514) );
  XNOR2_X1 U518 ( .A(n517), .B(n518), .ZN(n457) );
  NAND2_X1 U519 ( .A1(n519), .A2(n520), .ZN(n517) );
  NAND2_X1 U520 ( .A1(a_4_), .A2(n516), .ZN(n458) );
  NAND2_X1 U521 ( .A1(n521), .A2(n522), .ZN(n516) );
  NAND2_X1 U522 ( .A1(n523), .A2(b_7_), .ZN(n522) );
  NOR2_X1 U523 ( .A1(n524), .A2(n525), .ZN(n523) );
  NOR2_X1 U524 ( .A1(n526), .A2(n452), .ZN(n524) );
  NAND2_X1 U525 ( .A1(n526), .A2(n452), .ZN(n521) );
  XOR2_X1 U526 ( .A(n527), .B(n528), .Z(n452) );
  NOR2_X1 U527 ( .A1(n529), .A2(n530), .ZN(n528) );
  XNOR2_X1 U528 ( .A(n531), .B(n532), .ZN(n460) );
  XNOR2_X1 U529 ( .A(n533), .B(n534), .ZN(n532) );
  XNOR2_X1 U530 ( .A(n535), .B(n536), .ZN(n464) );
  XOR2_X1 U531 ( .A(n537), .B(n538), .Z(n535) );
  NOR2_X1 U532 ( .A1(n512), .A2(n495), .ZN(n538) );
  XOR2_X1 U533 ( .A(n539), .B(n540), .Z(n415) );
  XOR2_X1 U534 ( .A(n541), .B(n542), .Z(n539) );
  XOR2_X1 U535 ( .A(n543), .B(n544), .Z(n422) );
  XOR2_X1 U536 ( .A(n545), .B(n546), .Z(n543) );
  NOR2_X1 U537 ( .A1(n433), .A2(n547), .ZN(n485) );
  AND2_X1 U538 ( .A1(n435), .A2(n434), .ZN(n433) );
  NOR2_X1 U539 ( .A1(n547), .A2(n548), .ZN(n434) );
  AND2_X1 U540 ( .A1(n549), .A2(n550), .ZN(n548) );
  NOR2_X1 U541 ( .A1(n550), .A2(n549), .ZN(n547) );
  AND2_X1 U542 ( .A1(n551), .A2(n552), .ZN(n549) );
  NAND2_X1 U543 ( .A1(n553), .A2(n554), .ZN(n552) );
  XNOR2_X1 U544 ( .A(n555), .B(n556), .ZN(n550) );
  XNOR2_X1 U545 ( .A(n557), .B(n558), .ZN(n556) );
  NOR2_X1 U546 ( .A1(n487), .A2(n488), .ZN(n435) );
  XOR2_X1 U547 ( .A(n559), .B(n553), .Z(n488) );
  XNOR2_X1 U548 ( .A(n560), .B(n561), .ZN(n553) );
  NAND2_X1 U549 ( .A1(n562), .A2(n563), .ZN(n560) );
  NAND2_X1 U550 ( .A1(n551), .A2(n554), .ZN(n559) );
  NAND2_X1 U551 ( .A1(n564), .A2(n565), .ZN(n554) );
  NAND2_X1 U552 ( .A1(a_0_), .A2(b_5_), .ZN(n565) );
  INV_X1 U553 ( .A(n566), .ZN(n564) );
  NAND2_X1 U554 ( .A1(a_0_), .A2(n566), .ZN(n551) );
  NAND2_X1 U555 ( .A1(n567), .A2(n568), .ZN(n566) );
  NAND2_X1 U556 ( .A1(n569), .A2(n570), .ZN(n568) );
  OR2_X1 U557 ( .A1(n571), .A2(n572), .ZN(n570) );
  NAND2_X1 U558 ( .A1(n572), .A2(n571), .ZN(n567) );
  NOR2_X1 U559 ( .A1(n492), .A2(n573), .ZN(n487) );
  AND2_X1 U560 ( .A1(n489), .A2(n574), .ZN(n573) );
  NAND2_X1 U561 ( .A1(n575), .A2(n576), .ZN(n574) );
  NAND2_X1 U562 ( .A1(a_0_), .A2(b_6_), .ZN(n576) );
  XOR2_X1 U563 ( .A(n577), .B(n572), .Z(n489) );
  XOR2_X1 U564 ( .A(n578), .B(n579), .Z(n572) );
  NOR2_X1 U565 ( .A1(n580), .A2(n581), .ZN(n579) );
  NOR2_X1 U566 ( .A1(n582), .A2(n583), .ZN(n580) );
  NOR2_X1 U567 ( .A1(n584), .A2(n507), .ZN(n583) );
  INV_X1 U568 ( .A(n585), .ZN(n582) );
  XOR2_X1 U569 ( .A(n569), .B(n571), .Z(n577) );
  NAND2_X1 U570 ( .A1(n586), .A2(n587), .ZN(n571) );
  NAND2_X1 U571 ( .A1(n588), .A2(a_2_), .ZN(n587) );
  NOR2_X1 U572 ( .A1(n589), .A2(n530), .ZN(n588) );
  NOR2_X1 U573 ( .A1(n590), .A2(n591), .ZN(n589) );
  NAND2_X1 U574 ( .A1(n591), .A2(n590), .ZN(n586) );
  NOR2_X1 U575 ( .A1(n420), .A2(n530), .ZN(n569) );
  NOR2_X1 U576 ( .A1(n496), .A2(n575), .ZN(n492) );
  INV_X1 U577 ( .A(n494), .ZN(n575) );
  NAND2_X1 U578 ( .A1(n592), .A2(n593), .ZN(n494) );
  NAND2_X1 U579 ( .A1(n546), .A2(n594), .ZN(n593) );
  OR2_X1 U580 ( .A1(n545), .A2(n544), .ZN(n594) );
  NOR2_X1 U581 ( .A1(n420), .A2(n495), .ZN(n546) );
  NAND2_X1 U582 ( .A1(n544), .A2(n545), .ZN(n592) );
  NAND2_X1 U583 ( .A1(n595), .A2(n596), .ZN(n545) );
  NAND2_X1 U584 ( .A1(n542), .A2(n597), .ZN(n596) );
  OR2_X1 U585 ( .A1(n540), .A2(n541), .ZN(n597) );
  NOR2_X1 U586 ( .A1(n507), .A2(n495), .ZN(n542) );
  NAND2_X1 U587 ( .A1(n540), .A2(n541), .ZN(n595) );
  NAND2_X1 U588 ( .A1(n598), .A2(n599), .ZN(n541) );
  NAND2_X1 U589 ( .A1(n600), .A2(b_6_), .ZN(n599) );
  NOR2_X1 U590 ( .A1(n601), .A2(n512), .ZN(n600) );
  NOR2_X1 U591 ( .A1(n536), .A2(n537), .ZN(n601) );
  NAND2_X1 U592 ( .A1(n536), .A2(n537), .ZN(n598) );
  NAND2_X1 U593 ( .A1(n602), .A2(n603), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n534), .A2(n604), .ZN(n603) );
  OR2_X1 U595 ( .A1(n533), .A2(n531), .ZN(n604) );
  NOR2_X1 U596 ( .A1(n495), .A2(n605), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n531), .A2(n533), .ZN(n602) );
  NAND2_X1 U598 ( .A1(n519), .A2(n606), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n518), .A2(n520), .ZN(n606) );
  NAND2_X1 U600 ( .A1(n607), .A2(n608), .ZN(n520) );
  INV_X1 U601 ( .A(n609), .ZN(n608) );
  NAND2_X1 U602 ( .A1(b_6_), .A2(a_5_), .ZN(n607) );
  XNOR2_X1 U603 ( .A(n610), .B(n611), .ZN(n518) );
  NOR2_X1 U604 ( .A1(n529), .A2(n584), .ZN(n611) );
  NAND2_X1 U605 ( .A1(n609), .A2(a_5_), .ZN(n519) );
  NOR2_X1 U606 ( .A1(n450), .A2(n610), .ZN(n609) );
  NAND2_X1 U607 ( .A1(b_6_), .A2(a_7_), .ZN(n450) );
  XNOR2_X1 U608 ( .A(n612), .B(n613), .ZN(n531) );
  XNOR2_X1 U609 ( .A(n614), .B(n615), .ZN(n612) );
  XNOR2_X1 U610 ( .A(n616), .B(n617), .ZN(n536) );
  NAND2_X1 U611 ( .A1(n618), .A2(n619), .ZN(n616) );
  XOR2_X1 U612 ( .A(n620), .B(n621), .Z(n540) );
  XOR2_X1 U613 ( .A(n622), .B(n623), .Z(n620) );
  NOR2_X1 U614 ( .A1(n530), .A2(n512), .ZN(n623) );
  XNOR2_X1 U615 ( .A(n591), .B(n624), .ZN(n544) );
  XOR2_X1 U616 ( .A(n590), .B(n625), .Z(n624) );
  NAND2_X1 U617 ( .A1(a_2_), .A2(b_5_), .ZN(n625) );
  NAND2_X1 U618 ( .A1(n626), .A2(n627), .ZN(n590) );
  NAND2_X1 U619 ( .A1(n628), .A2(a_3_), .ZN(n627) );
  NOR2_X1 U620 ( .A1(n629), .A2(n530), .ZN(n628) );
  NOR2_X1 U621 ( .A1(n621), .A2(n622), .ZN(n629) );
  NAND2_X1 U622 ( .A1(n621), .A2(n622), .ZN(n626) );
  NAND2_X1 U623 ( .A1(n618), .A2(n630), .ZN(n622) );
  NAND2_X1 U624 ( .A1(n617), .A2(n619), .ZN(n630) );
  NAND2_X1 U625 ( .A1(n631), .A2(n632), .ZN(n619) );
  NAND2_X1 U626 ( .A1(b_5_), .A2(a_4_), .ZN(n632) );
  INV_X1 U627 ( .A(n633), .ZN(n631) );
  XOR2_X1 U628 ( .A(n634), .B(n635), .Z(n617) );
  NOR2_X1 U629 ( .A1(n636), .A2(n637), .ZN(n635) );
  NOR2_X1 U630 ( .A1(n638), .A2(n639), .ZN(n636) );
  NOR2_X1 U631 ( .A1(n525), .A2(n584), .ZN(n639) );
  INV_X1 U632 ( .A(n640), .ZN(n638) );
  NAND2_X1 U633 ( .A1(a_4_), .A2(n633), .ZN(n618) );
  NAND2_X1 U634 ( .A1(n641), .A2(n642), .ZN(n633) );
  NAND2_X1 U635 ( .A1(n615), .A2(n643), .ZN(n642) );
  OR2_X1 U636 ( .A1(n613), .A2(n614), .ZN(n643) );
  NOR2_X1 U637 ( .A1(n644), .A2(n610), .ZN(n615) );
  NAND2_X1 U638 ( .A1(b_5_), .A2(a_6_), .ZN(n610) );
  NAND2_X1 U639 ( .A1(a_7_), .A2(b_4_), .ZN(n644) );
  NAND2_X1 U640 ( .A1(n614), .A2(n613), .ZN(n641) );
  XOR2_X1 U641 ( .A(n645), .B(n646), .Z(n613) );
  XNOR2_X1 U642 ( .A(n647), .B(n648), .ZN(n621) );
  XOR2_X1 U643 ( .A(n649), .B(n650), .Z(n647) );
  XOR2_X1 U644 ( .A(n651), .B(n652), .Z(n591) );
  XNOR2_X1 U645 ( .A(n653), .B(n654), .ZN(n651) );
  XNOR2_X1 U646 ( .A(n483), .B(n655), .ZN(n437) );
  NAND2_X1 U647 ( .A1(n656), .A2(n483), .ZN(n440) );
  AND2_X1 U648 ( .A1(n657), .A2(n658), .ZN(n483) );
  NAND2_X1 U649 ( .A1(n557), .A2(n659), .ZN(n658) );
  OR2_X1 U650 ( .A1(n555), .A2(n558), .ZN(n659) );
  AND2_X1 U651 ( .A1(n562), .A2(n660), .ZN(n557) );
  NAND2_X1 U652 ( .A1(n561), .A2(n563), .ZN(n660) );
  NAND2_X1 U653 ( .A1(n661), .A2(n662), .ZN(n563) );
  NAND2_X1 U654 ( .A1(a_1_), .A2(b_4_), .ZN(n662) );
  XNOR2_X1 U655 ( .A(n663), .B(n664), .ZN(n561) );
  XNOR2_X1 U656 ( .A(n665), .B(n666), .ZN(n663) );
  NOR2_X1 U657 ( .A1(n667), .A2(n507), .ZN(n666) );
  OR2_X1 U658 ( .A1(n420), .A2(n661), .ZN(n562) );
  NOR2_X1 U659 ( .A1(n581), .A2(n668), .ZN(n661) );
  AND2_X1 U660 ( .A1(n578), .A2(n669), .ZN(n668) );
  NAND2_X1 U661 ( .A1(n585), .A2(n670), .ZN(n669) );
  NAND2_X1 U662 ( .A1(a_2_), .A2(b_4_), .ZN(n670) );
  XNOR2_X1 U663 ( .A(n671), .B(n672), .ZN(n578) );
  XNOR2_X1 U664 ( .A(n673), .B(n674), .ZN(n672) );
  NOR2_X1 U665 ( .A1(n585), .A2(n507), .ZN(n581) );
  NAND2_X1 U666 ( .A1(n675), .A2(n676), .ZN(n585) );
  NAND2_X1 U667 ( .A1(n652), .A2(n677), .ZN(n676) );
  NAND2_X1 U668 ( .A1(n654), .A2(n653), .ZN(n677) );
  XOR2_X1 U669 ( .A(n678), .B(n679), .Z(n652) );
  NAND2_X1 U670 ( .A1(n680), .A2(n681), .ZN(n678) );
  OR2_X1 U671 ( .A1(n654), .A2(n653), .ZN(n675) );
  AND2_X1 U672 ( .A1(n682), .A2(n683), .ZN(n653) );
  NAND2_X1 U673 ( .A1(n684), .A2(n649), .ZN(n683) );
  OR2_X1 U674 ( .A1(n648), .A2(n650), .ZN(n684) );
  NAND2_X1 U675 ( .A1(n648), .A2(n650), .ZN(n682) );
  NOR2_X1 U676 ( .A1(n637), .A2(n685), .ZN(n650) );
  AND2_X1 U677 ( .A1(n634), .A2(n686), .ZN(n685) );
  NAND2_X1 U678 ( .A1(n640), .A2(n687), .ZN(n686) );
  NAND2_X1 U679 ( .A1(b_4_), .A2(a_5_), .ZN(n687) );
  AND2_X1 U680 ( .A1(n688), .A2(n689), .ZN(n634) );
  NAND2_X1 U681 ( .A1(n690), .A2(n691), .ZN(n689) );
  NAND2_X1 U682 ( .A1(b_3_), .A2(a_6_), .ZN(n690) );
  NOR2_X1 U683 ( .A1(n640), .A2(n525), .ZN(n637) );
  NAND2_X1 U684 ( .A1(n645), .A2(n646), .ZN(n640) );
  NOR2_X1 U685 ( .A1(n584), .A2(n692), .ZN(n646) );
  NOR2_X1 U686 ( .A1(n667), .A2(n529), .ZN(n645) );
  XNOR2_X1 U687 ( .A(n693), .B(n694), .ZN(n648) );
  NOR2_X1 U688 ( .A1(n695), .A2(n696), .ZN(n694) );
  NOR2_X1 U689 ( .A1(n697), .A2(n698), .ZN(n695) );
  NOR2_X1 U690 ( .A1(n667), .A2(n525), .ZN(n698) );
  INV_X1 U691 ( .A(n688), .ZN(n697) );
  NOR2_X1 U692 ( .A1(n512), .A2(n584), .ZN(n654) );
  NAND2_X1 U693 ( .A1(n555), .A2(n558), .ZN(n657) );
  NAND2_X1 U694 ( .A1(a_0_), .A2(b_4_), .ZN(n558) );
  XOR2_X1 U695 ( .A(n699), .B(n700), .Z(n555) );
  XOR2_X1 U696 ( .A(n701), .B(n702), .Z(n700) );
  NOR2_X1 U697 ( .A1(n655), .A2(n481), .ZN(n656) );
  XNOR2_X1 U698 ( .A(n703), .B(n704), .ZN(n481) );
  INV_X1 U699 ( .A(n484), .ZN(n655) );
  XOR2_X1 U700 ( .A(n705), .B(n706), .Z(n484) );
  XNOR2_X1 U701 ( .A(n707), .B(n708), .ZN(n706) );
  NAND2_X1 U702 ( .A1(a_0_), .A2(b_3_), .ZN(n708) );
  NAND2_X1 U703 ( .A1(n709), .A2(n710), .ZN(n445) );
  NAND2_X1 U704 ( .A1(n703), .A2(n704), .ZN(n710) );
  NAND2_X1 U705 ( .A1(n711), .A2(n703), .ZN(n444) );
  XNOR2_X1 U706 ( .A(n712), .B(n713), .ZN(n703) );
  NAND2_X1 U707 ( .A1(n714), .A2(n715), .ZN(n712) );
  NOR2_X1 U708 ( .A1(n716), .A2(n709), .ZN(n711) );
  XNOR2_X1 U709 ( .A(n477), .B(n476), .ZN(n709) );
  INV_X1 U710 ( .A(n704), .ZN(n716) );
  NAND2_X1 U711 ( .A1(n717), .A2(n718), .ZN(n704) );
  NAND2_X1 U712 ( .A1(n719), .A2(a_0_), .ZN(n718) );
  NOR2_X1 U713 ( .A1(n720), .A2(n667), .ZN(n719) );
  NOR2_X1 U714 ( .A1(n707), .A2(n705), .ZN(n720) );
  NAND2_X1 U715 ( .A1(n707), .A2(n705), .ZN(n717) );
  XOR2_X1 U716 ( .A(n721), .B(n722), .Z(n705) );
  XOR2_X1 U717 ( .A(n723), .B(n724), .Z(n721) );
  AND2_X1 U718 ( .A1(n725), .A2(n726), .ZN(n707) );
  NAND2_X1 U719 ( .A1(n701), .A2(n727), .ZN(n726) );
  NAND2_X1 U720 ( .A1(n702), .A2(n699), .ZN(n727) );
  AND2_X1 U721 ( .A1(n728), .A2(n729), .ZN(n701) );
  NAND2_X1 U722 ( .A1(n730), .A2(a_2_), .ZN(n729) );
  NOR2_X1 U723 ( .A1(n731), .A2(n667), .ZN(n730) );
  NOR2_X1 U724 ( .A1(n665), .A2(n664), .ZN(n731) );
  NAND2_X1 U725 ( .A1(n665), .A2(n664), .ZN(n728) );
  XOR2_X1 U726 ( .A(n732), .B(n733), .Z(n664) );
  XNOR2_X1 U727 ( .A(n734), .B(n735), .ZN(n732) );
  NAND2_X1 U728 ( .A1(a_3_), .A2(b_2_), .ZN(n734) );
  AND2_X1 U729 ( .A1(n736), .A2(n737), .ZN(n665) );
  NAND2_X1 U730 ( .A1(n738), .A2(n739), .ZN(n737) );
  NAND2_X1 U731 ( .A1(n671), .A2(n674), .ZN(n738) );
  OR2_X1 U732 ( .A1(n671), .A2(n674), .ZN(n736) );
  NAND2_X1 U733 ( .A1(n680), .A2(n740), .ZN(n674) );
  NAND2_X1 U734 ( .A1(n679), .A2(n681), .ZN(n740) );
  NAND2_X1 U735 ( .A1(n741), .A2(n742), .ZN(n681) );
  NAND2_X1 U736 ( .A1(a_4_), .A2(b_3_), .ZN(n742) );
  XNOR2_X1 U737 ( .A(n743), .B(n744), .ZN(n679) );
  NAND2_X1 U738 ( .A1(n745), .A2(n746), .ZN(n743) );
  OR2_X1 U739 ( .A1(n605), .A2(n741), .ZN(n680) );
  NOR2_X1 U740 ( .A1(n696), .A2(n747), .ZN(n741) );
  AND2_X1 U741 ( .A1(n693), .A2(n748), .ZN(n747) );
  NAND2_X1 U742 ( .A1(n688), .A2(n749), .ZN(n748) );
  NAND2_X1 U743 ( .A1(a_5_), .A2(b_3_), .ZN(n749) );
  XOR2_X1 U744 ( .A(n750), .B(n751), .Z(n693) );
  NOR2_X1 U745 ( .A1(n688), .A2(n525), .ZN(n696) );
  NAND2_X1 U746 ( .A1(n752), .A2(b_3_), .ZN(n688) );
  NOR2_X1 U747 ( .A1(n691), .A2(n692), .ZN(n752) );
  NAND2_X1 U748 ( .A1(b_2_), .A2(a_7_), .ZN(n691) );
  XNOR2_X1 U749 ( .A(n753), .B(n754), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n755), .A2(n756), .ZN(n753) );
  OR2_X1 U751 ( .A1(n699), .A2(n702), .ZN(n725) );
  NOR2_X1 U752 ( .A1(n420), .A2(n667), .ZN(n702) );
  XOR2_X1 U753 ( .A(n757), .B(n758), .Z(n699) );
  XOR2_X1 U754 ( .A(n759), .B(n760), .Z(n757) );
  INV_X1 U755 ( .A(n448), .ZN(n471) );
  NAND2_X1 U756 ( .A1(n761), .A2(n762), .ZN(n448) );
  NOR2_X1 U757 ( .A1(n477), .A2(n476), .ZN(n762) );
  XNOR2_X1 U758 ( .A(n763), .B(n764), .ZN(n476) );
  NOR2_X1 U759 ( .A1(n765), .A2(n766), .ZN(n764) );
  INV_X1 U760 ( .A(n767), .ZN(n766) );
  NOR2_X1 U761 ( .A1(n768), .A2(n769), .ZN(n765) );
  AND2_X1 U762 ( .A1(n714), .A2(n770), .ZN(n477) );
  NAND2_X1 U763 ( .A1(n713), .A2(n715), .ZN(n770) );
  NAND2_X1 U764 ( .A1(n771), .A2(n772), .ZN(n715) );
  NAND2_X1 U765 ( .A1(a_0_), .A2(b_2_), .ZN(n772) );
  INV_X1 U766 ( .A(n773), .ZN(n771) );
  XOR2_X1 U767 ( .A(n774), .B(n775), .Z(n713) );
  XNOR2_X1 U768 ( .A(n776), .B(n777), .ZN(n775) );
  NAND2_X1 U769 ( .A1(b_0_), .A2(a_2_), .ZN(n774) );
  NAND2_X1 U770 ( .A1(a_0_), .A2(n773), .ZN(n714) );
  NAND2_X1 U771 ( .A1(n778), .A2(n779), .ZN(n773) );
  NAND2_X1 U772 ( .A1(n724), .A2(n780), .ZN(n779) );
  OR2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n780) );
  NOR2_X1 U774 ( .A1(n420), .A2(n781), .ZN(n724) );
  NAND2_X1 U775 ( .A1(n722), .A2(n723), .ZN(n778) );
  NAND2_X1 U776 ( .A1(n782), .A2(n783), .ZN(n723) );
  NAND2_X1 U777 ( .A1(n760), .A2(n784), .ZN(n783) );
  OR2_X1 U778 ( .A1(n759), .A2(n758), .ZN(n784) );
  NAND2_X1 U779 ( .A1(n758), .A2(n759), .ZN(n782) );
  NAND2_X1 U780 ( .A1(n785), .A2(n786), .ZN(n759) );
  NAND2_X1 U781 ( .A1(n787), .A2(a_3_), .ZN(n786) );
  NOR2_X1 U782 ( .A1(n788), .A2(n781), .ZN(n787) );
  NOR2_X1 U783 ( .A1(n733), .A2(n735), .ZN(n788) );
  NAND2_X1 U784 ( .A1(n733), .A2(n735), .ZN(n785) );
  NAND2_X1 U785 ( .A1(n755), .A2(n789), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n754), .A2(n756), .ZN(n789) );
  NAND2_X1 U787 ( .A1(n790), .A2(n791), .ZN(n756) );
  NAND2_X1 U788 ( .A1(a_4_), .A2(b_2_), .ZN(n791) );
  INV_X1 U789 ( .A(n792), .ZN(n790) );
  XOR2_X1 U790 ( .A(n793), .B(n794), .Z(n754) );
  AND2_X1 U791 ( .A1(n795), .A2(n796), .ZN(n794) );
  NAND2_X1 U792 ( .A1(a_4_), .A2(n792), .ZN(n755) );
  NAND2_X1 U793 ( .A1(n745), .A2(n797), .ZN(n792) );
  NAND2_X1 U794 ( .A1(n744), .A2(n746), .ZN(n797) );
  NAND2_X1 U795 ( .A1(n798), .A2(n799), .ZN(n746) );
  NAND2_X1 U796 ( .A1(a_5_), .A2(b_2_), .ZN(n799) );
  AND2_X1 U797 ( .A1(n795), .A2(n800), .ZN(n744) );
  NAND2_X1 U798 ( .A1(n801), .A2(n802), .ZN(n800) );
  NAND2_X1 U799 ( .A1(b_0_), .A2(a_7_), .ZN(n802) );
  NAND2_X1 U800 ( .A1(b_1_), .A2(a_6_), .ZN(n801) );
  OR2_X1 U801 ( .A1(n798), .A2(n525), .ZN(n745) );
  NAND2_X1 U802 ( .A1(n750), .A2(n751), .ZN(n798) );
  NOR2_X1 U803 ( .A1(n692), .A2(n781), .ZN(n750) );
  XOR2_X1 U804 ( .A(n803), .B(n804), .Z(n733) );
  XOR2_X1 U805 ( .A(n805), .B(n806), .Z(n803) );
  XOR2_X1 U806 ( .A(n807), .B(n808), .Z(n758) );
  XNOR2_X1 U807 ( .A(n809), .B(n810), .ZN(n808) );
  NAND2_X1 U808 ( .A1(b_0_), .A2(a_4_), .ZN(n807) );
  XOR2_X1 U809 ( .A(n811), .B(n812), .Z(n722) );
  NOR2_X1 U810 ( .A1(n813), .A2(n814), .ZN(n812) );
  INV_X1 U811 ( .A(n815), .ZN(n814) );
  NOR2_X1 U812 ( .A1(n816), .A2(n817), .ZN(n813) );
  NOR2_X1 U813 ( .A1(n818), .A2(n470), .ZN(n761) );
  NAND2_X1 U814 ( .A1(n767), .A2(n819), .ZN(n470) );
  NAND2_X1 U815 ( .A1(n820), .A2(n763), .ZN(n819) );
  NAND2_X1 U816 ( .A1(n821), .A2(n822), .ZN(n763) );
  NAND2_X1 U817 ( .A1(n823), .A2(b_0_), .ZN(n822) );
  NOR2_X1 U818 ( .A1(n824), .A2(n507), .ZN(n823) );
  NOR2_X1 U819 ( .A1(n776), .A2(n777), .ZN(n824) );
  NAND2_X1 U820 ( .A1(n776), .A2(n777), .ZN(n821) );
  NAND2_X1 U821 ( .A1(n815), .A2(n825), .ZN(n777) );
  NAND2_X1 U822 ( .A1(n826), .A2(n811), .ZN(n825) );
  NAND2_X1 U823 ( .A1(n827), .A2(n828), .ZN(n811) );
  NAND2_X1 U824 ( .A1(n829), .A2(b_0_), .ZN(n828) );
  NOR2_X1 U825 ( .A1(n830), .A2(n605), .ZN(n829) );
  NOR2_X1 U826 ( .A1(n810), .A2(n809), .ZN(n830) );
  NAND2_X1 U827 ( .A1(n810), .A2(n809), .ZN(n827) );
  NAND2_X1 U828 ( .A1(n831), .A2(n832), .ZN(n809) );
  NAND2_X1 U829 ( .A1(n804), .A2(n833), .ZN(n832) );
  OR2_X1 U830 ( .A1(n806), .A2(n805), .ZN(n833) );
  AND2_X1 U831 ( .A1(b_0_), .A2(a_5_), .ZN(n804) );
  NAND2_X1 U832 ( .A1(n805), .A2(n806), .ZN(n831) );
  NAND2_X1 U833 ( .A1(n834), .A2(n795), .ZN(n806) );
  NAND2_X1 U834 ( .A1(n796), .A2(n751), .ZN(n795) );
  NOR2_X1 U835 ( .A1(n835), .A2(n529), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n793), .A2(n796), .ZN(n834) );
  AND2_X1 U837 ( .A1(b_0_), .A2(a_6_), .ZN(n796) );
  NOR2_X1 U838 ( .A1(n835), .A2(n525), .ZN(n793) );
  NOR2_X1 U839 ( .A1(n605), .A2(n835), .ZN(n805) );
  NOR2_X1 U840 ( .A1(n512), .A2(n835), .ZN(n810) );
  NAND2_X1 U841 ( .A1(n836), .A2(n507), .ZN(n826) );
  NAND2_X1 U842 ( .A1(n817), .A2(n816), .ZN(n815) );
  INV_X1 U843 ( .A(n836), .ZN(n816) );
  NAND2_X1 U844 ( .A1(b_0_), .A2(a_3_), .ZN(n836) );
  NOR2_X1 U845 ( .A1(n835), .A2(n507), .ZN(n817) );
  NAND2_X1 U846 ( .A1(n837), .A2(n496), .ZN(n820) );
  NAND2_X1 U847 ( .A1(n769), .A2(n768), .ZN(n767) );
  INV_X1 U848 ( .A(n837), .ZN(n768) );
  NAND2_X1 U849 ( .A1(b_0_), .A2(a_1_), .ZN(n837) );
  NOR2_X1 U850 ( .A1(n835), .A2(n496), .ZN(n769) );
  INV_X1 U851 ( .A(a_0_), .ZN(n496) );
  XNOR2_X1 U852 ( .A(n419), .B(a_7_), .ZN(Result_add_7_) );
  NAND2_X1 U853 ( .A1(n838), .A2(n455), .ZN(Result_add_6_) );
  INV_X1 U854 ( .A(n526), .ZN(n455) );
  NOR2_X1 U855 ( .A1(n839), .A2(n840), .ZN(n526) );
  NOR2_X1 U856 ( .A1(n841), .A2(n842), .ZN(n838) );
  NOR2_X1 U857 ( .A1(n495), .A2(n843), .ZN(n842) );
  NAND2_X1 U858 ( .A1(n839), .A2(n692), .ZN(n843) );
  INV_X1 U859 ( .A(Result_mul_15_), .ZN(n839) );
  NOR2_X1 U860 ( .A1(b_6_), .A2(n844), .ZN(n841) );
  XNOR2_X1 U861 ( .A(Result_mul_15_), .B(a_6_), .ZN(n844) );
  NAND2_X1 U862 ( .A1(n845), .A2(n846), .ZN(Result_add_5_) );
  NAND2_X1 U863 ( .A1(n614), .A2(n847), .ZN(n846) );
  NOR2_X1 U864 ( .A1(n848), .A2(n849), .ZN(n845) );
  NOR2_X1 U865 ( .A1(b_5_), .A2(n850), .ZN(n849) );
  XNOR2_X1 U866 ( .A(n525), .B(n851), .ZN(n850) );
  NOR2_X1 U867 ( .A1(n530), .A2(n852), .ZN(n848) );
  NAND2_X1 U868 ( .A1(n851), .A2(n525), .ZN(n852) );
  INV_X1 U869 ( .A(n847), .ZN(n851) );
  XNOR2_X1 U870 ( .A(n853), .B(n854), .ZN(Result_add_4_) );
  NAND2_X1 U871 ( .A1(n649), .A2(n855), .ZN(n853) );
  NAND2_X1 U872 ( .A1(n856), .A2(n857), .ZN(Result_add_3_) );
  NAND2_X1 U873 ( .A1(n673), .A2(n858), .ZN(n857) );
  NOR2_X1 U874 ( .A1(n859), .A2(n860), .ZN(n856) );
  NOR2_X1 U875 ( .A1(b_3_), .A2(n861), .ZN(n860) );
  XNOR2_X1 U876 ( .A(a_3_), .B(n858), .ZN(n861) );
  NOR2_X1 U877 ( .A1(n667), .A2(n862), .ZN(n859) );
  OR2_X1 U878 ( .A1(n858), .A2(a_3_), .ZN(n862) );
  XNOR2_X1 U879 ( .A(n863), .B(n864), .ZN(Result_add_2_) );
  NOR2_X1 U880 ( .A1(n865), .A2(n760), .ZN(n864) );
  NAND2_X1 U881 ( .A1(n866), .A2(n867), .ZN(Result_add_1_) );
  NAND2_X1 U882 ( .A1(n868), .A2(n869), .ZN(n867) );
  OR2_X1 U883 ( .A1(n776), .A2(n870), .ZN(n868) );
  NAND2_X1 U884 ( .A1(n871), .A2(n872), .ZN(n866) );
  XNOR2_X1 U885 ( .A(n835), .B(a_1_), .ZN(n871) );
  XOR2_X1 U886 ( .A(n873), .B(n874), .Z(Result_add_0_) );
  NOR2_X1 U887 ( .A1(n875), .A2(n478), .ZN(n874) );
  INV_X1 U888 ( .A(n818), .ZN(n478) );
  NAND2_X1 U889 ( .A1(a_0_), .A2(b_0_), .ZN(n818) );
  NOR2_X1 U890 ( .A1(b_0_), .A2(a_0_), .ZN(n875) );
  NOR2_X1 U891 ( .A1(n870), .A2(n876), .ZN(n873) );
  NOR2_X1 U892 ( .A1(n776), .A2(n869), .ZN(n876) );
  INV_X1 U893 ( .A(n872), .ZN(n869) );
  NOR2_X1 U894 ( .A1(n760), .A2(n877), .ZN(n872) );
  NOR2_X1 U895 ( .A1(n865), .A2(n863), .ZN(n877) );
  AND2_X1 U896 ( .A1(n739), .A2(n878), .ZN(n863) );
  NAND2_X1 U897 ( .A1(n879), .A2(n858), .ZN(n878) );
  NAND2_X1 U898 ( .A1(n649), .A2(n880), .ZN(n858) );
  NAND2_X1 U899 ( .A1(n855), .A2(n854), .ZN(n880) );
  OR2_X1 U900 ( .A1(n614), .A2(n881), .ZN(n854) );
  AND2_X1 U901 ( .A1(n882), .A2(n847), .ZN(n881) );
  NAND2_X1 U902 ( .A1(n840), .A2(n883), .ZN(n847) );
  NAND2_X1 U903 ( .A1(Result_mul_15_), .A2(n884), .ZN(n883) );
  NAND2_X1 U904 ( .A1(n495), .A2(n692), .ZN(n884) );
  NOR2_X1 U905 ( .A1(n419), .A2(n529), .ZN(Result_mul_15_) );
  INV_X1 U906 ( .A(a_7_), .ZN(n529) );
  INV_X1 U907 ( .A(b_7_), .ZN(n419) );
  INV_X1 U908 ( .A(n527), .ZN(n840) );
  NOR2_X1 U909 ( .A1(n495), .A2(n692), .ZN(n527) );
  INV_X1 U910 ( .A(a_6_), .ZN(n692) );
  INV_X1 U911 ( .A(b_6_), .ZN(n495) );
  NAND2_X1 U912 ( .A1(n530), .A2(n525), .ZN(n882) );
  NOR2_X1 U913 ( .A1(n530), .A2(n525), .ZN(n614) );
  INV_X1 U914 ( .A(a_5_), .ZN(n525) );
  INV_X1 U915 ( .A(b_5_), .ZN(n530) );
  NAND2_X1 U916 ( .A1(n584), .A2(n605), .ZN(n855) );
  INV_X1 U917 ( .A(a_4_), .ZN(n605) );
  INV_X1 U918 ( .A(b_4_), .ZN(n584) );
  NAND2_X1 U919 ( .A1(b_4_), .A2(a_4_), .ZN(n649) );
  NAND2_X1 U920 ( .A1(n667), .A2(n512), .ZN(n879) );
  INV_X1 U921 ( .A(n673), .ZN(n739) );
  NOR2_X1 U922 ( .A1(n512), .A2(n667), .ZN(n673) );
  INV_X1 U923 ( .A(b_3_), .ZN(n667) );
  INV_X1 U924 ( .A(a_3_), .ZN(n512) );
  NOR2_X1 U925 ( .A1(b_2_), .A2(a_2_), .ZN(n865) );
  NOR2_X1 U926 ( .A1(n507), .A2(n781), .ZN(n760) );
  INV_X1 U927 ( .A(b_2_), .ZN(n781) );
  INV_X1 U928 ( .A(a_2_), .ZN(n507) );
  NOR2_X1 U929 ( .A1(n420), .A2(n835), .ZN(n776) );
  INV_X1 U930 ( .A(b_1_), .ZN(n835) );
  INV_X1 U931 ( .A(a_1_), .ZN(n420) );
  NOR2_X1 U932 ( .A1(b_1_), .A2(a_1_), .ZN(n870) );
endmodule

