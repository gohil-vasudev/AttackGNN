module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n318_, new_n155_, new_n384_, new_n163_, new_n236_, new_n238_, new_n148_, new_n321_, new_n122_, new_n324_, new_n250_, new_n113_, new_n111_, new_n288_, new_n158_, new_n371_, new_n252_, new_n202_, new_n262_, new_n296_, new_n160_, new_n308_, new_n271_, new_n274_, new_n372_, new_n242_, new_n368_, new_n232_, new_n218_, new_n115_, new_n258_, new_n307_, new_n190_, new_n176_, new_n305_, new_n156_, new_n223_, new_n283_, new_n306_, new_n291_, new_n366_, new_n261_, new_n241_, new_n309_, new_n186_, new_n339_, new_n213_, new_n134_, new_n197_, new_n205_, new_n323_, new_n141_, new_n365_, new_n259_, new_n362_, new_n386_, new_n206_, new_n109_, new_n254_, new_n227_, new_n355_, new_n353_, new_n222_, new_n265_, new_n246_, new_n170_, new_n256_, new_n328_, new_n266_, new_n367_, new_n278_, new_n304_, new_n381_, new_n130_, new_n173_, new_n220_, new_n268_, new_n217_, new_n269_, new_n374_, new_n376_, new_n194_, new_n380_, new_n214_, new_n116_, new_n129_, new_n138_, new_n142_, new_n299_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n139_, new_n240_, new_n314_, new_n352_, new_n118_, new_n363_, new_n165_, new_n123_, new_n127_, new_n211_, new_n126_, new_n342_, new_n327_, new_n216_, new_n177_, new_n196_, new_n280_, new_n264_, new_n319_, new_n235_, new_n273_, new_n224_, new_n301_, new_n169_, new_n270_, new_n338_, new_n383_, new_n317_, new_n210_, new_n343_, new_n143_, new_n344_, new_n207_, new_n125_, new_n145_, new_n267_, new_n287_, new_n253_, new_n140_, new_n336_, new_n247_, new_n377_, new_n237_, new_n330_, new_n375_, new_n234_, new_n149_, new_n294_, new_n187_, new_n260_, new_n311_, new_n251_, new_n189_, new_n300_, new_n292_, new_n195_, new_n263_, new_n215_, new_n331_, new_n334_, new_n152_, new_n341_, new_n378_, new_n157_, new_n182_, new_n153_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n133_, new_n277_, new_n245_, new_n212_, new_n151_, new_n286_, new_n335_, new_n347_, new_n364_, new_n193_, new_n219_, new_n231_, new_n313_, new_n239_, new_n382_, new_n272_, new_n282_, new_n346_, new_n198_, new_n201_, new_n128_, new_n192_, new_n199_, new_n146_, new_n358_, new_n208_, new_n348_, new_n360_, new_n159_, new_n110_, new_n228_, new_n315_, new_n322_, new_n302_, new_n191_, new_n124_, new_n289_, new_n326_, new_n179_, new_n225_, new_n164_, new_n230_, new_n175_, new_n226_, new_n281_, new_n185_, new_n373_, new_n112_, new_n171_, new_n248_, new_n350_, new_n117_, new_n121_, new_n167_, new_n221_, new_n243_, new_n385_, new_n200_, new_n345_, new_n298_, new_n184_, new_n131_, new_n255_, new_n329_, new_n249_, new_n136_, new_n233_, new_n284_, new_n119_, new_n293_, new_n178_, new_n168_, new_n174_, new_n297_, new_n279_, new_n361_, new_n150_, new_n295_, new_n359_, new_n120_, new_n132_, new_n354_, new_n166_, new_n108_, new_n137_, new_n162_, new_n183_, new_n303_, new_n161_, new_n340_, new_n147_, new_n285_, new_n356_, new_n333_, new_n229_, new_n209_, new_n337_, new_n351_, new_n290_, new_n203_, new_n316_, new_n204_, new_n325_, new_n181_, new_n135_, new_n180_, new_n276_, new_n332_;

not g000 ( new_n108_, keyIn_0_36 );
not g001 ( new_n109_, keyIn_0_21 );
xnor g002 ( new_n110_, keyIn_0_4, N24 );
and g003 ( new_n111_, new_n110_, N30 );
xnor g004 ( new_n112_, new_n111_, new_n109_ );
not g005 ( new_n113_, keyIn_0_26 );
xnor g006 ( new_n114_, keyIn_0_14, N89 );
and g007 ( new_n115_, new_n114_, N95 );
xnor g008 ( new_n116_, new_n115_, new_n113_ );
not g009 ( new_n117_, N4 );
xnor g010 ( new_n118_, keyIn_0_0, N1 );
or g011 ( new_n119_, new_n118_, new_n117_ );
xnor g012 ( new_n120_, new_n119_, keyIn_0_18 );
and g013 ( new_n121_, new_n120_, new_n112_, new_n116_ );
not g014 ( new_n122_, keyIn_0_25 );
xnor g015 ( new_n123_, keyIn_0_12, N76 );
and g016 ( new_n124_, new_n123_, N82 );
xnor g017 ( new_n125_, new_n124_, new_n122_ );
not g018 ( new_n126_, keyIn_0_27 );
and g019 ( new_n127_, keyIn_0_16, N102 );
not g020 ( new_n128_, new_n127_ );
or g021 ( new_n129_, keyIn_0_16, N102 );
and g022 ( new_n130_, new_n128_, N108, new_n129_ );
xnor g023 ( new_n131_, new_n130_, new_n126_ );
and g024 ( new_n132_, new_n125_, new_n131_ );
xnor g025 ( new_n133_, keyIn_0_10, N63 );
and g026 ( new_n134_, new_n133_, N69 );
xnor g027 ( new_n135_, new_n134_, keyIn_0_24 );
not g028 ( new_n136_, keyIn_0_20 );
or g029 ( new_n137_, keyIn_0_2, N11 );
and g030 ( new_n138_, keyIn_0_2, N11 );
not g031 ( new_n139_, new_n138_ );
and g032 ( new_n140_, new_n139_, N17, new_n137_ );
xnor g033 ( new_n141_, new_n140_, new_n136_ );
and g034 ( new_n142_, new_n135_, new_n141_ );
not g035 ( new_n143_, keyIn_0_22 );
xnor g036 ( new_n144_, keyIn_0_6, N37 );
and g037 ( new_n145_, new_n144_, N43 );
xnor g038 ( new_n146_, new_n145_, new_n143_ );
not g039 ( new_n147_, keyIn_0_23 );
not g040 ( new_n148_, N56 );
xnor g041 ( new_n149_, keyIn_0_8, N50 );
or g042 ( new_n150_, new_n149_, new_n148_ );
xnor g043 ( new_n151_, new_n150_, new_n147_ );
and g044 ( new_n152_, new_n151_, new_n146_ );
and g045 ( new_n153_, new_n121_, new_n152_, new_n132_, new_n142_ );
xnor g046 ( N223, new_n153_, new_n108_ );
not g047 ( new_n155_, keyIn_0_50 );
not g048 ( new_n156_, keyIn_0_41 );
not g049 ( new_n157_, keyIn_0_37 );
xnor g050 ( new_n158_, N223, new_n157_ );
xnor g051 ( new_n159_, new_n158_, new_n146_ );
xnor g052 ( new_n160_, new_n159_, new_n156_ );
xnor g053 ( new_n161_, keyIn_0_7, N43 );
not g054 ( new_n162_, new_n161_ );
or g055 ( new_n163_, new_n162_, N47 );
xnor g056 ( new_n164_, new_n163_, keyIn_0_30 );
and g057 ( new_n165_, new_n160_, new_n164_ );
xnor g058 ( new_n166_, new_n165_, new_n155_ );
not g059 ( new_n167_, keyIn_0_48 );
not g060 ( new_n168_, keyIn_0_39 );
xnor g061 ( new_n169_, new_n158_, new_n141_ );
xnor g062 ( new_n170_, new_n169_, new_n168_ );
xnor g063 ( new_n171_, keyIn_0_3, N17 );
or g064 ( new_n172_, new_n171_, N21 );
xor g065 ( new_n173_, new_n172_, keyIn_0_28 );
and g066 ( new_n174_, new_n170_, new_n173_ );
xnor g067 ( new_n175_, new_n174_, new_n167_ );
not g068 ( new_n176_, keyIn_0_47 );
xor g069 ( new_n177_, keyIn_0_1, N4 );
or g070 ( new_n178_, new_n177_, N8 );
xnor g071 ( new_n179_, new_n178_, keyIn_0_19 );
not g072 ( new_n180_, new_n179_ );
not g073 ( new_n181_, keyIn_0_38 );
xnor g074 ( new_n182_, new_n158_, new_n120_ );
or g075 ( new_n183_, new_n182_, new_n181_ );
xnor g076 ( new_n184_, N223, keyIn_0_37 );
and g077 ( new_n185_, new_n184_, new_n120_ );
not g078 ( new_n186_, new_n120_ );
and g079 ( new_n187_, new_n158_, new_n186_ );
or g080 ( new_n188_, new_n185_, new_n187_, keyIn_0_38 );
and g081 ( new_n189_, new_n183_, new_n180_, new_n188_ );
xnor g082 ( new_n190_, new_n189_, new_n176_ );
and g083 ( new_n191_, new_n166_, new_n175_, new_n190_ );
not g084 ( new_n192_, keyIn_0_42 );
xnor g085 ( new_n193_, new_n158_, new_n151_ );
xnor g086 ( new_n194_, new_n193_, new_n192_ );
xor g087 ( new_n195_, keyIn_0_9, N56 );
not g088 ( new_n196_, new_n195_ );
or g089 ( new_n197_, new_n196_, N60 );
xnor g090 ( new_n198_, new_n197_, keyIn_0_31 );
and g091 ( new_n199_, new_n194_, new_n198_ );
xnor g092 ( new_n200_, new_n199_, keyIn_0_51 );
not g093 ( new_n201_, keyIn_0_52 );
xnor g094 ( new_n202_, new_n184_, new_n135_ );
xnor g095 ( new_n203_, new_n202_, keyIn_0_43 );
xnor g096 ( new_n204_, keyIn_0_11, N69 );
or g097 ( new_n205_, new_n204_, N73 );
xor g098 ( new_n206_, new_n205_, keyIn_0_32 );
and g099 ( new_n207_, new_n203_, new_n206_ );
xnor g100 ( new_n208_, new_n207_, new_n201_ );
and g101 ( new_n209_, new_n200_, new_n208_ );
xnor g102 ( new_n210_, new_n158_, new_n131_ );
xnor g103 ( new_n211_, new_n210_, keyIn_0_46 );
not g104 ( new_n212_, N112 );
xnor g105 ( new_n213_, keyIn_0_17, N108 );
and g106 ( new_n214_, new_n213_, new_n212_ );
xor g107 ( new_n215_, new_n214_, keyIn_0_35 );
and g108 ( new_n216_, new_n211_, new_n215_ );
xnor g109 ( new_n217_, new_n216_, keyIn_0_55 );
not g110 ( new_n218_, keyIn_0_54 );
xnor g111 ( new_n219_, new_n158_, new_n116_ );
xnor g112 ( new_n220_, new_n219_, keyIn_0_45 );
not g113 ( new_n221_, N99 );
xnor g114 ( new_n222_, keyIn_0_15, N95 );
and g115 ( new_n223_, new_n222_, new_n221_ );
xnor g116 ( new_n224_, new_n223_, keyIn_0_34 );
and g117 ( new_n225_, new_n220_, new_n224_ );
xnor g118 ( new_n226_, new_n225_, new_n218_ );
and g119 ( new_n227_, new_n217_, new_n226_ );
not g120 ( new_n228_, keyIn_0_53 );
xnor g121 ( new_n229_, new_n158_, new_n125_ );
xnor g122 ( new_n230_, new_n229_, keyIn_0_44 );
not g123 ( new_n231_, N86 );
or g124 ( new_n232_, keyIn_0_13, N82 );
and g125 ( new_n233_, keyIn_0_13, N82 );
not g126 ( new_n234_, new_n233_ );
and g127 ( new_n235_, new_n234_, new_n231_, new_n232_ );
xor g128 ( new_n236_, new_n235_, keyIn_0_33 );
not g129 ( new_n237_, new_n236_ );
and g130 ( new_n238_, new_n230_, new_n237_ );
or g131 ( new_n239_, new_n238_, new_n228_ );
not g132 ( new_n240_, new_n230_ );
or g133 ( new_n241_, new_n240_, keyIn_0_53, new_n236_ );
not g134 ( new_n242_, N34 );
xor g135 ( new_n243_, keyIn_0_5, N30 );
and g136 ( new_n244_, new_n243_, new_n242_ );
xnor g137 ( new_n245_, new_n244_, keyIn_0_29 );
not g138 ( new_n246_, keyIn_0_40 );
xnor g139 ( new_n247_, new_n158_, new_n112_ );
xnor g140 ( new_n248_, new_n247_, new_n246_ );
not g141 ( new_n249_, new_n248_ );
or g142 ( new_n250_, new_n249_, keyIn_0_49, new_n245_ );
not g143 ( new_n251_, keyIn_0_49 );
not g144 ( new_n252_, new_n245_ );
and g145 ( new_n253_, new_n248_, new_n252_ );
or g146 ( new_n254_, new_n253_, new_n251_ );
and g147 ( new_n255_, new_n239_, new_n254_, new_n241_, new_n250_ );
and g148 ( new_n256_, new_n191_, new_n209_, new_n227_, new_n255_ );
xnor g149 ( N329, new_n256_, keyIn_0_60 );
not g150 ( new_n258_, keyIn_0_62 );
xnor g151 ( new_n259_, N329, keyIn_0_61 );
xnor g152 ( new_n260_, new_n259_, new_n217_ );
not g153 ( new_n261_, N115 );
and g154 ( new_n262_, new_n211_, new_n261_, new_n213_ );
xor g155 ( new_n263_, new_n262_, keyIn_0_59 );
or g156 ( new_n264_, new_n260_, new_n263_ );
xnor g157 ( new_n265_, new_n259_, new_n200_ );
not g158 ( new_n266_, new_n194_ );
or g159 ( new_n267_, new_n266_, N66, new_n196_ );
or g160 ( new_n268_, new_n265_, new_n267_ );
xnor g161 ( new_n269_, new_n259_, new_n226_ );
not g162 ( new_n270_, N105 );
and g163 ( new_n271_, new_n220_, new_n270_, new_n222_ );
xnor g164 ( new_n272_, new_n271_, keyIn_0_58 );
or g165 ( new_n273_, new_n269_, new_n272_ );
and g166 ( new_n274_, new_n264_, new_n268_, new_n273_ );
and g167 ( new_n275_, new_n254_, new_n250_ );
xnor g168 ( new_n276_, new_n259_, new_n275_ );
not g169 ( new_n277_, new_n243_ );
or g170 ( new_n278_, new_n249_, N40, new_n277_ );
or g171 ( new_n279_, new_n276_, new_n278_ );
xnor g172 ( new_n280_, new_n259_, new_n166_ );
not g173 ( new_n281_, new_n160_ );
or g174 ( new_n282_, new_n281_, N53, new_n162_ );
or g175 ( new_n283_, new_n280_, new_n282_ );
and g176 ( new_n284_, new_n279_, new_n283_ );
and g177 ( new_n285_, new_n239_, new_n241_ );
xnor g178 ( new_n286_, new_n259_, new_n285_ );
not g179 ( new_n287_, N92 );
and g180 ( new_n288_, new_n230_, new_n287_, new_n232_, new_n234_ );
xor g181 ( new_n289_, new_n288_, keyIn_0_57 );
or g182 ( new_n290_, new_n286_, new_n289_ );
xnor g183 ( new_n291_, new_n259_, new_n208_ );
not g184 ( new_n292_, N79 );
not g185 ( new_n293_, new_n204_ );
and g186 ( new_n294_, new_n203_, new_n292_, new_n293_ );
xor g187 ( new_n295_, new_n294_, keyIn_0_56 );
or g188 ( new_n296_, new_n291_, new_n295_ );
and g189 ( new_n297_, new_n290_, new_n296_ );
xnor g190 ( new_n298_, new_n259_, new_n190_ );
xnor g191 ( new_n299_, new_n182_, new_n181_ );
or g192 ( new_n300_, new_n299_, N14, new_n177_ );
or g193 ( new_n301_, new_n298_, new_n300_ );
xnor g194 ( new_n302_, new_n259_, new_n175_ );
not g195 ( new_n303_, new_n170_ );
or g196 ( new_n304_, new_n303_, N27, new_n171_ );
or g197 ( new_n305_, new_n302_, new_n304_ );
and g198 ( new_n306_, new_n301_, new_n305_ );
and g199 ( new_n307_, new_n274_, new_n284_, new_n297_, new_n306_ );
or g200 ( new_n308_, new_n307_, new_n258_ );
and g201 ( new_n309_, new_n290_, new_n296_, new_n301_, new_n305_ );
and g202 ( new_n310_, new_n309_, new_n258_, new_n274_, new_n284_ );
not g203 ( new_n311_, new_n310_ );
and g204 ( N370, new_n308_, new_n311_ );
not g205 ( new_n313_, keyIn_0_63 );
and g206 ( new_n314_, new_n308_, N27, new_n311_ );
not g207 ( new_n315_, N17 );
and g208 ( new_n316_, N329, N21 );
and g209 ( new_n317_, N223, N11 );
or g210 ( new_n318_, new_n316_, new_n315_, new_n317_ );
or g211 ( new_n319_, new_n314_, new_n318_ );
and g212 ( new_n320_, new_n308_, N40, new_n311_ );
not g213 ( new_n321_, N30 );
and g214 ( new_n322_, N329, N34 );
and g215 ( new_n323_, N223, N24 );
or g216 ( new_n324_, new_n322_, new_n321_, new_n323_ );
or g217 ( new_n325_, new_n320_, new_n324_ );
and g218 ( new_n326_, new_n308_, N53, new_n311_ );
not g219 ( new_n327_, N43 );
and g220 ( new_n328_, N329, N47 );
and g221 ( new_n329_, N223, N37 );
or g222 ( new_n330_, new_n328_, new_n327_, new_n329_ );
or g223 ( new_n331_, new_n326_, new_n330_ );
and g224 ( new_n332_, new_n308_, N66, new_n311_ );
and g225 ( new_n333_, N329, N60 );
and g226 ( new_n334_, N223, N50 );
or g227 ( new_n335_, new_n333_, new_n148_, new_n334_ );
or g228 ( new_n336_, new_n332_, new_n335_ );
and g229 ( new_n337_, new_n319_, new_n325_, new_n331_, new_n336_ );
and g230 ( new_n338_, new_n308_, N105, new_n311_ );
not g231 ( new_n339_, N95 );
and g232 ( new_n340_, N329, N99 );
and g233 ( new_n341_, N223, N89 );
or g234 ( new_n342_, new_n340_, new_n339_, new_n341_ );
or g235 ( new_n343_, new_n338_, new_n342_ );
and g236 ( new_n344_, new_n308_, N115, new_n311_ );
not g237 ( new_n345_, N108 );
and g238 ( new_n346_, N329, N112 );
and g239 ( new_n347_, N223, N102 );
or g240 ( new_n348_, new_n346_, new_n345_, new_n347_ );
or g241 ( new_n349_, new_n344_, new_n348_ );
and g242 ( new_n350_, new_n308_, N79, new_n311_ );
not g243 ( new_n351_, N69 );
and g244 ( new_n352_, N329, N73 );
and g245 ( new_n353_, N223, N63 );
or g246 ( new_n354_, new_n352_, new_n351_, new_n353_ );
or g247 ( new_n355_, new_n350_, new_n354_ );
and g248 ( new_n356_, new_n308_, N92, new_n311_ );
not g249 ( new_n357_, N82 );
and g250 ( new_n358_, N329, N86 );
and g251 ( new_n359_, N223, N76 );
or g252 ( new_n360_, new_n358_, new_n357_, new_n359_ );
or g253 ( new_n361_, new_n356_, new_n360_ );
and g254 ( new_n362_, new_n343_, new_n349_, new_n355_, new_n361_ );
and g255 ( new_n363_, new_n337_, new_n362_ );
xnor g256 ( new_n364_, new_n363_, new_n313_ );
and g257 ( new_n365_, N370, N14 );
and g258 ( new_n366_, N329, N8 );
and g259 ( new_n367_, N223, N1 );
or g260 ( new_n368_, new_n365_, new_n117_, new_n366_, new_n367_ );
and g261 ( N421, new_n364_, new_n368_ );
not g262 ( N430, new_n337_ );
and g263 ( new_n371_, new_n319_, new_n325_ );
not g264 ( new_n372_, new_n371_ );
not g265 ( new_n373_, new_n361_ );
and g266 ( new_n374_, new_n373_, new_n331_, new_n336_ );
not g267 ( new_n375_, new_n350_ );
not g268 ( new_n376_, new_n354_ );
and g269 ( new_n377_, new_n336_, new_n375_, new_n376_ );
and g270 ( new_n378_, new_n377_, new_n325_, new_n331_ );
or g271 ( N431, new_n378_, new_n372_, new_n374_ );
not g272 ( new_n380_, new_n319_ );
not g273 ( new_n381_, new_n331_ );
not g274 ( new_n382_, new_n338_ );
not g275 ( new_n383_, new_n342_ );
and g276 ( new_n384_, new_n361_, new_n382_, new_n383_ );
or g277 ( new_n385_, new_n377_, new_n384_, new_n381_ );
and g278 ( new_n386_, new_n385_, new_n325_ );
or g279 ( N432, new_n386_, new_n380_ );
endmodule