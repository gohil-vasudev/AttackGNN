module add_mul_comp_sub_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, 
        a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, 
        b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, 
        b_13_, b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   Result_9_, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543;
  assign Result_8_ = Result_9_;
  assign Result_6_ = Result_9_;
  assign Result_4_ = Result_9_;
  assign Result_2_ = Result_9_;
  assign Result_15_ = Result_9_;
  assign Result_13_ = Result_9_;
  assign Result_11_ = Result_9_;
  assign Result_0_ = Result_9_;
  assign Result_10_ = Result_9_;
  assign Result_12_ = Result_9_;
  assign Result_14_ = Result_9_;
  assign Result_1_ = Result_9_;
  assign Result_3_ = Result_9_;
  assign Result_5_ = Result_9_;
  assign Result_7_ = Result_9_;

  INV_X1 U289 ( .A(n272), .ZN(Result_31_) );
  AND2_X1 U290 ( .A1(n273), .A2(n274), .ZN(n272) );
  OR2_X1 U291 ( .A1(n275), .A2(n276), .ZN(Result_30_) );
  AND2_X1 U292 ( .A1(n277), .A2(n278), .ZN(n276) );
  OR2_X1 U293 ( .A1(n279), .A2(n280), .ZN(n278) );
  AND2_X1 U294 ( .A1(Result_9_), .A2(n274), .ZN(n280) );
  INV_X1 U295 ( .A(n281), .ZN(n274) );
  AND2_X1 U296 ( .A1(n282), .A2(n283), .ZN(n279) );
  INV_X1 U297 ( .A(n284), .ZN(n283) );
  AND2_X1 U298 ( .A1(a_15_), .A2(b_15_), .ZN(n284) );
  AND2_X1 U299 ( .A1(n285), .A2(n286), .ZN(n275) );
  OR2_X1 U300 ( .A1(n287), .A2(n288), .ZN(n286) );
  AND2_X1 U301 ( .A1(n281), .A2(Result_9_), .ZN(n288) );
  AND3_X1 U302 ( .A1(b_15_), .A2(a_15_), .A3(n282), .ZN(n287) );
  INV_X1 U303 ( .A(n277), .ZN(n285) );
  OR2_X1 U304 ( .A1(n289), .A2(n290), .ZN(n277) );
  INV_X1 U305 ( .A(n291), .ZN(n290) );
  OR2_X1 U306 ( .A1(n292), .A2(n293), .ZN(Result_29_) );
  AND2_X1 U307 ( .A1(n294), .A2(Result_9_), .ZN(n293) );
  XOR2_X1 U308 ( .A(n295), .B(n296), .Z(n294) );
  AND2_X1 U309 ( .A1(n282), .A2(n297), .ZN(n292) );
  XOR2_X1 U310 ( .A(n296), .B(n298), .Z(n297) );
  OR2_X1 U311 ( .A1(n299), .A2(n300), .ZN(n296) );
  INV_X1 U312 ( .A(n301), .ZN(n300) );
  OR2_X1 U313 ( .A1(n302), .A2(n303), .ZN(Result_28_) );
  AND2_X1 U314 ( .A1(n304), .A2(Result_9_), .ZN(n303) );
  XOR2_X1 U315 ( .A(n305), .B(n306), .Z(n304) );
  AND2_X1 U316 ( .A1(n307), .A2(n282), .ZN(n302) );
  XNOR2_X1 U317 ( .A(n306), .B(n308), .ZN(n307) );
  OR2_X1 U318 ( .A1(n309), .A2(n310), .ZN(n306) );
  INV_X1 U319 ( .A(n311), .ZN(n310) );
  OR2_X1 U320 ( .A1(n312), .A2(n313), .ZN(Result_27_) );
  AND2_X1 U321 ( .A1(n314), .A2(Result_9_), .ZN(n313) );
  XOR2_X1 U322 ( .A(n315), .B(n316), .Z(n314) );
  AND2_X1 U323 ( .A1(n317), .A2(n282), .ZN(n312) );
  XNOR2_X1 U324 ( .A(n316), .B(n318), .ZN(n317) );
  OR2_X1 U325 ( .A1(n319), .A2(n320), .ZN(n316) );
  INV_X1 U326 ( .A(n321), .ZN(n320) );
  OR2_X1 U327 ( .A1(n322), .A2(n323), .ZN(Result_26_) );
  AND2_X1 U328 ( .A1(n324), .A2(Result_9_), .ZN(n323) );
  XOR2_X1 U329 ( .A(n325), .B(n326), .Z(n324) );
  AND2_X1 U330 ( .A1(n327), .A2(n282), .ZN(n322) );
  XNOR2_X1 U331 ( .A(n326), .B(n328), .ZN(n327) );
  OR2_X1 U332 ( .A1(n329), .A2(n330), .ZN(n326) );
  INV_X1 U333 ( .A(n331), .ZN(n330) );
  OR2_X1 U334 ( .A1(n332), .A2(n333), .ZN(Result_25_) );
  AND2_X1 U335 ( .A1(n334), .A2(Result_9_), .ZN(n333) );
  XOR2_X1 U336 ( .A(n335), .B(n336), .Z(n334) );
  AND2_X1 U337 ( .A1(n337), .A2(n282), .ZN(n332) );
  XNOR2_X1 U338 ( .A(n336), .B(n338), .ZN(n337) );
  OR2_X1 U339 ( .A1(n339), .A2(n340), .ZN(n336) );
  INV_X1 U340 ( .A(n341), .ZN(n340) );
  OR2_X1 U341 ( .A1(n342), .A2(n343), .ZN(Result_24_) );
  AND2_X1 U342 ( .A1(n344), .A2(Result_9_), .ZN(n343) );
  XOR2_X1 U343 ( .A(n345), .B(n346), .Z(n344) );
  AND2_X1 U344 ( .A1(n347), .A2(n282), .ZN(n342) );
  XNOR2_X1 U345 ( .A(n346), .B(n348), .ZN(n347) );
  OR2_X1 U346 ( .A1(n349), .A2(n350), .ZN(n346) );
  INV_X1 U347 ( .A(n351), .ZN(n350) );
  OR2_X1 U348 ( .A1(n352), .A2(n353), .ZN(Result_23_) );
  AND2_X1 U349 ( .A1(n354), .A2(Result_9_), .ZN(n353) );
  XOR2_X1 U350 ( .A(n355), .B(n356), .Z(n354) );
  AND2_X1 U351 ( .A1(n357), .A2(n282), .ZN(n352) );
  XNOR2_X1 U352 ( .A(n356), .B(n358), .ZN(n357) );
  OR2_X1 U353 ( .A1(n359), .A2(n360), .ZN(n356) );
  INV_X1 U354 ( .A(n361), .ZN(n360) );
  OR2_X1 U355 ( .A1(n362), .A2(n363), .ZN(Result_22_) );
  AND2_X1 U356 ( .A1(n364), .A2(Result_9_), .ZN(n363) );
  XOR2_X1 U357 ( .A(n365), .B(n366), .Z(n364) );
  AND2_X1 U358 ( .A1(n367), .A2(n282), .ZN(n362) );
  XNOR2_X1 U359 ( .A(n366), .B(n368), .ZN(n367) );
  OR2_X1 U360 ( .A1(n369), .A2(n370), .ZN(n366) );
  INV_X1 U361 ( .A(n371), .ZN(n370) );
  OR2_X1 U362 ( .A1(n372), .A2(n373), .ZN(Result_21_) );
  AND2_X1 U363 ( .A1(n374), .A2(Result_9_), .ZN(n373) );
  XOR2_X1 U364 ( .A(n375), .B(n376), .Z(n374) );
  AND2_X1 U365 ( .A1(n377), .A2(n282), .ZN(n372) );
  XNOR2_X1 U366 ( .A(n376), .B(n378), .ZN(n377) );
  OR2_X1 U367 ( .A1(n379), .A2(n380), .ZN(n376) );
  INV_X1 U368 ( .A(n381), .ZN(n380) );
  OR2_X1 U369 ( .A1(n382), .A2(n383), .ZN(Result_20_) );
  AND2_X1 U370 ( .A1(n384), .A2(Result_9_), .ZN(n383) );
  XOR2_X1 U371 ( .A(n385), .B(n386), .Z(n384) );
  AND2_X1 U372 ( .A1(n387), .A2(n282), .ZN(n382) );
  XNOR2_X1 U373 ( .A(n386), .B(n388), .ZN(n387) );
  OR2_X1 U374 ( .A1(n389), .A2(n390), .ZN(n386) );
  INV_X1 U375 ( .A(n391), .ZN(n390) );
  OR2_X1 U376 ( .A1(n392), .A2(n393), .ZN(Result_19_) );
  AND2_X1 U377 ( .A1(n394), .A2(Result_9_), .ZN(n393) );
  XOR2_X1 U378 ( .A(n395), .B(n396), .Z(n394) );
  AND2_X1 U379 ( .A1(n397), .A2(n282), .ZN(n392) );
  XNOR2_X1 U380 ( .A(n396), .B(n398), .ZN(n397) );
  OR2_X1 U381 ( .A1(n399), .A2(n400), .ZN(n396) );
  INV_X1 U382 ( .A(n401), .ZN(n400) );
  OR2_X1 U383 ( .A1(n402), .A2(n403), .ZN(Result_18_) );
  AND2_X1 U384 ( .A1(n404), .A2(Result_9_), .ZN(n403) );
  XOR2_X1 U385 ( .A(n405), .B(n406), .Z(n404) );
  AND2_X1 U386 ( .A1(n407), .A2(n282), .ZN(n402) );
  XNOR2_X1 U387 ( .A(n406), .B(n408), .ZN(n407) );
  OR2_X1 U388 ( .A1(n409), .A2(n410), .ZN(n406) );
  INV_X1 U389 ( .A(n411), .ZN(n410) );
  OR2_X1 U390 ( .A1(n412), .A2(n413), .ZN(Result_17_) );
  AND2_X1 U391 ( .A1(n414), .A2(Result_9_), .ZN(n413) );
  XOR2_X1 U392 ( .A(n415), .B(n416), .Z(n414) );
  AND2_X1 U393 ( .A1(n417), .A2(n282), .ZN(n412) );
  XOR2_X1 U394 ( .A(n416), .B(n418), .Z(n417) );
  OR2_X1 U395 ( .A1(n419), .A2(n420), .ZN(n416) );
  INV_X1 U396 ( .A(n421), .ZN(n420) );
  OR2_X1 U397 ( .A1(n422), .A2(n423), .ZN(Result_16_) );
  AND2_X1 U398 ( .A1(n424), .A2(Result_9_), .ZN(n423) );
  OR2_X1 U399 ( .A1(n425), .A2(n426), .ZN(n424) );
  INV_X1 U400 ( .A(n427), .ZN(n425) );
  OR2_X1 U401 ( .A1(n419), .A2(n428), .ZN(n427) );
  AND2_X1 U402 ( .A1(n415), .A2(n421), .ZN(n428) );
  OR2_X1 U403 ( .A1(n429), .A2(n409), .ZN(n415) );
  AND2_X1 U404 ( .A1(n405), .A2(n411), .ZN(n429) );
  OR2_X1 U405 ( .A1(n430), .A2(n399), .ZN(n405) );
  AND2_X1 U406 ( .A1(n395), .A2(n401), .ZN(n430) );
  OR2_X1 U407 ( .A1(n431), .A2(n389), .ZN(n395) );
  AND2_X1 U408 ( .A1(n385), .A2(n391), .ZN(n431) );
  OR2_X1 U409 ( .A1(n432), .A2(n379), .ZN(n385) );
  AND2_X1 U410 ( .A1(n375), .A2(n381), .ZN(n432) );
  OR2_X1 U411 ( .A1(n433), .A2(n369), .ZN(n375) );
  AND2_X1 U412 ( .A1(n365), .A2(n371), .ZN(n433) );
  OR2_X1 U413 ( .A1(n434), .A2(n359), .ZN(n365) );
  AND2_X1 U414 ( .A1(n355), .A2(n361), .ZN(n434) );
  OR2_X1 U415 ( .A1(n435), .A2(n349), .ZN(n355) );
  AND2_X1 U416 ( .A1(n345), .A2(n351), .ZN(n435) );
  OR2_X1 U417 ( .A1(n436), .A2(n339), .ZN(n345) );
  AND2_X1 U418 ( .A1(n335), .A2(n341), .ZN(n436) );
  OR2_X1 U419 ( .A1(n437), .A2(n329), .ZN(n335) );
  AND2_X1 U420 ( .A1(n325), .A2(n331), .ZN(n437) );
  OR2_X1 U421 ( .A1(n438), .A2(n319), .ZN(n325) );
  AND2_X1 U422 ( .A1(n315), .A2(n321), .ZN(n438) );
  OR2_X1 U423 ( .A1(n439), .A2(n309), .ZN(n315) );
  AND2_X1 U424 ( .A1(n305), .A2(n311), .ZN(n439) );
  OR2_X1 U425 ( .A1(n440), .A2(n299), .ZN(n305) );
  AND2_X1 U426 ( .A1(n295), .A2(n301), .ZN(n440) );
  OR2_X1 U427 ( .A1(n441), .A2(n289), .ZN(n295) );
  AND2_X1 U428 ( .A1(n442), .A2(a_14_), .ZN(n289) );
  AND2_X1 U429 ( .A1(n281), .A2(n291), .ZN(n441) );
  AND2_X1 U430 ( .A1(n443), .A2(a_1_), .ZN(n419) );
  AND2_X1 U431 ( .A1(n444), .A2(n282), .ZN(n422) );
  INV_X1 U432 ( .A(n445), .ZN(n282) );
  OR2_X1 U433 ( .A1(Result_9_), .A2(n446), .ZN(n445) );
  AND4_X1 U434 ( .A1(n447), .A2(n448), .A3(n449), .A4(n450), .ZN(n446) );
  AND4_X1 U435 ( .A1(n371), .A2(n381), .A3(n391), .A4(n401), .ZN(n450) );
  AND3_X1 U436 ( .A1(n351), .A2(n361), .A3(n341), .ZN(n449) );
  AND4_X1 U437 ( .A1(n301), .A2(n311), .A3(n321), .A4(n331), .ZN(n448) );
  AND3_X1 U438 ( .A1(n291), .A2(n273), .A3(n451), .ZN(n447) );
  OR2_X1 U439 ( .A1(a_15_), .A2(n452), .ZN(n273) );
  OR2_X1 U440 ( .A1(a_14_), .A2(n442), .ZN(n291) );
  OR3_X1 U441 ( .A1(n453), .A2(n454), .A3(n455), .ZN(Result_9_) );
  AND2_X1 U442 ( .A1(a_0_), .A2(n456), .ZN(n455) );
  AND2_X1 U443 ( .A1(n451), .A2(n457), .ZN(n454) );
  OR3_X1 U444 ( .A1(n399), .A2(n409), .A3(n458), .ZN(n457) );
  AND3_X1 U445 ( .A1(n391), .A2(n401), .A3(n459), .ZN(n458) );
  OR3_X1 U446 ( .A1(n379), .A2(n389), .A3(n460), .ZN(n459) );
  AND3_X1 U447 ( .A1(n371), .A2(n381), .A3(n461), .ZN(n460) );
  OR3_X1 U448 ( .A1(n359), .A2(n369), .A3(n462), .ZN(n461) );
  AND3_X1 U449 ( .A1(n351), .A2(n361), .A3(n463), .ZN(n462) );
  OR3_X1 U450 ( .A1(n339), .A2(n349), .A3(n464), .ZN(n463) );
  AND3_X1 U451 ( .A1(n331), .A2(n341), .A3(n465), .ZN(n464) );
  OR3_X1 U452 ( .A1(n319), .A2(n329), .A3(n466), .ZN(n465) );
  AND3_X1 U453 ( .A1(n311), .A2(n321), .A3(n467), .ZN(n466) );
  OR3_X1 U454 ( .A1(n299), .A2(n309), .A3(n468), .ZN(n467) );
  AND3_X1 U455 ( .A1(n469), .A2(n301), .A3(n470), .ZN(n468) );
  OR2_X1 U456 ( .A1(n281), .A2(a_14_), .ZN(n470) );
  OR2_X1 U457 ( .A1(a_13_), .A2(n471), .ZN(n301) );
  OR2_X1 U458 ( .A1(n472), .A2(n442), .ZN(n469) );
  INV_X1 U459 ( .A(b_14_), .ZN(n442) );
  AND2_X1 U460 ( .A1(a_14_), .A2(n281), .ZN(n472) );
  AND2_X1 U461 ( .A1(n452), .A2(a_15_), .ZN(n281) );
  INV_X1 U462 ( .A(b_15_), .ZN(n452) );
  AND2_X1 U463 ( .A1(n473), .A2(a_12_), .ZN(n309) );
  AND2_X1 U464 ( .A1(n471), .A2(a_13_), .ZN(n299) );
  OR2_X1 U465 ( .A1(a_11_), .A2(n474), .ZN(n321) );
  OR2_X1 U466 ( .A1(a_12_), .A2(n473), .ZN(n311) );
  AND2_X1 U467 ( .A1(n475), .A2(a_10_), .ZN(n329) );
  AND2_X1 U468 ( .A1(n474), .A2(a_11_), .ZN(n319) );
  OR2_X1 U469 ( .A1(a_9_), .A2(n476), .ZN(n341) );
  OR2_X1 U470 ( .A1(a_10_), .A2(n475), .ZN(n331) );
  AND2_X1 U471 ( .A1(n477), .A2(a_8_), .ZN(n349) );
  AND2_X1 U472 ( .A1(n476), .A2(a_9_), .ZN(n339) );
  OR2_X1 U473 ( .A1(a_7_), .A2(n478), .ZN(n361) );
  OR2_X1 U474 ( .A1(a_8_), .A2(n477), .ZN(n351) );
  AND2_X1 U475 ( .A1(n479), .A2(a_6_), .ZN(n369) );
  AND2_X1 U476 ( .A1(n478), .A2(a_7_), .ZN(n359) );
  OR2_X1 U477 ( .A1(a_5_), .A2(n480), .ZN(n381) );
  OR2_X1 U478 ( .A1(a_6_), .A2(n479), .ZN(n371) );
  AND2_X1 U479 ( .A1(n481), .A2(a_4_), .ZN(n389) );
  AND2_X1 U480 ( .A1(n480), .A2(a_5_), .ZN(n379) );
  OR2_X1 U481 ( .A1(a_3_), .A2(n482), .ZN(n401) );
  OR2_X1 U482 ( .A1(a_4_), .A2(n481), .ZN(n391) );
  AND2_X1 U483 ( .A1(n483), .A2(a_2_), .ZN(n409) );
  AND2_X1 U484 ( .A1(n482), .A2(a_3_), .ZN(n399) );
  AND3_X1 U485 ( .A1(n421), .A2(n484), .A3(n411), .ZN(n451) );
  OR2_X1 U486 ( .A1(a_2_), .A2(n483), .ZN(n411) );
  OR2_X1 U487 ( .A1(a_1_), .A2(n443), .ZN(n421) );
  AND3_X1 U488 ( .A1(n484), .A2(n443), .A3(a_1_), .ZN(n453) );
  INV_X1 U489 ( .A(b_1_), .ZN(n443) );
  XNOR2_X1 U490 ( .A(n426), .B(n485), .ZN(n444) );
  AND2_X1 U491 ( .A1(n486), .A2(n487), .ZN(n485) );
  OR2_X1 U492 ( .A1(b_1_), .A2(n488), .ZN(n487) );
  AND2_X1 U493 ( .A1(n418), .A2(a_1_), .ZN(n488) );
  OR2_X1 U494 ( .A1(a_1_), .A2(n418), .ZN(n486) );
  INV_X1 U495 ( .A(n489), .ZN(n418) );
  OR2_X1 U496 ( .A1(n490), .A2(n491), .ZN(n489) );
  AND2_X1 U497 ( .A1(n408), .A2(n492), .ZN(n491) );
  AND2_X1 U498 ( .A1(n493), .A2(n483), .ZN(n490) );
  INV_X1 U499 ( .A(b_2_), .ZN(n483) );
  OR2_X1 U500 ( .A1(n492), .A2(n408), .ZN(n493) );
  OR2_X1 U501 ( .A1(n494), .A2(n495), .ZN(n408) );
  AND2_X1 U502 ( .A1(n398), .A2(n496), .ZN(n495) );
  AND2_X1 U503 ( .A1(n497), .A2(n482), .ZN(n494) );
  INV_X1 U504 ( .A(b_3_), .ZN(n482) );
  OR2_X1 U505 ( .A1(n496), .A2(n398), .ZN(n497) );
  OR2_X1 U506 ( .A1(n498), .A2(n499), .ZN(n398) );
  AND2_X1 U507 ( .A1(n388), .A2(n500), .ZN(n499) );
  AND2_X1 U508 ( .A1(n501), .A2(n481), .ZN(n498) );
  INV_X1 U509 ( .A(b_4_), .ZN(n481) );
  OR2_X1 U510 ( .A1(n500), .A2(n388), .ZN(n501) );
  OR2_X1 U511 ( .A1(n502), .A2(n503), .ZN(n388) );
  AND2_X1 U512 ( .A1(n378), .A2(n504), .ZN(n503) );
  AND2_X1 U513 ( .A1(n505), .A2(n480), .ZN(n502) );
  INV_X1 U514 ( .A(b_5_), .ZN(n480) );
  OR2_X1 U515 ( .A1(n504), .A2(n378), .ZN(n505) );
  OR2_X1 U516 ( .A1(n506), .A2(n507), .ZN(n378) );
  AND2_X1 U517 ( .A1(n368), .A2(n508), .ZN(n507) );
  AND2_X1 U518 ( .A1(n509), .A2(n479), .ZN(n506) );
  INV_X1 U519 ( .A(b_6_), .ZN(n479) );
  OR2_X1 U520 ( .A1(n508), .A2(n368), .ZN(n509) );
  OR2_X1 U521 ( .A1(n510), .A2(n511), .ZN(n368) );
  AND2_X1 U522 ( .A1(n358), .A2(n512), .ZN(n511) );
  AND2_X1 U523 ( .A1(n513), .A2(n478), .ZN(n510) );
  INV_X1 U524 ( .A(b_7_), .ZN(n478) );
  OR2_X1 U525 ( .A1(n512), .A2(n358), .ZN(n513) );
  OR2_X1 U526 ( .A1(n514), .A2(n515), .ZN(n358) );
  AND2_X1 U527 ( .A1(n348), .A2(n516), .ZN(n515) );
  AND2_X1 U528 ( .A1(n517), .A2(n477), .ZN(n514) );
  INV_X1 U529 ( .A(b_8_), .ZN(n477) );
  OR2_X1 U530 ( .A1(n516), .A2(n348), .ZN(n517) );
  OR2_X1 U531 ( .A1(n518), .A2(n519), .ZN(n348) );
  AND2_X1 U532 ( .A1(n338), .A2(n520), .ZN(n519) );
  AND2_X1 U533 ( .A1(n521), .A2(n476), .ZN(n518) );
  INV_X1 U534 ( .A(b_9_), .ZN(n476) );
  OR2_X1 U535 ( .A1(n520), .A2(n338), .ZN(n521) );
  OR2_X1 U536 ( .A1(n522), .A2(n523), .ZN(n338) );
  AND2_X1 U537 ( .A1(n328), .A2(n524), .ZN(n523) );
  AND2_X1 U538 ( .A1(n525), .A2(n475), .ZN(n522) );
  INV_X1 U539 ( .A(b_10_), .ZN(n475) );
  OR2_X1 U540 ( .A1(n524), .A2(n328), .ZN(n525) );
  OR2_X1 U541 ( .A1(n526), .A2(n527), .ZN(n328) );
  AND2_X1 U542 ( .A1(n318), .A2(n528), .ZN(n527) );
  AND2_X1 U543 ( .A1(n529), .A2(n474), .ZN(n526) );
  INV_X1 U544 ( .A(b_11_), .ZN(n474) );
  OR2_X1 U545 ( .A1(n528), .A2(n318), .ZN(n529) );
  OR2_X1 U546 ( .A1(n530), .A2(n531), .ZN(n318) );
  AND2_X1 U547 ( .A1(n308), .A2(n532), .ZN(n531) );
  AND2_X1 U548 ( .A1(n533), .A2(n473), .ZN(n530) );
  INV_X1 U549 ( .A(b_12_), .ZN(n473) );
  OR2_X1 U550 ( .A1(n532), .A2(n308), .ZN(n533) );
  OR2_X1 U551 ( .A1(n534), .A2(n535), .ZN(n308) );
  AND2_X1 U552 ( .A1(n536), .A2(n537), .ZN(n535) );
  AND2_X1 U553 ( .A1(n538), .A2(n471), .ZN(n534) );
  INV_X1 U554 ( .A(b_13_), .ZN(n471) );
  OR2_X1 U555 ( .A1(n536), .A2(n537), .ZN(n538) );
  INV_X1 U556 ( .A(a_13_), .ZN(n537) );
  INV_X1 U557 ( .A(n298), .ZN(n536) );
  OR2_X1 U558 ( .A1(n539), .A2(n540), .ZN(n298) );
  AND2_X1 U559 ( .A1(b_14_), .A2(a_14_), .ZN(n540) );
  AND3_X1 U560 ( .A1(a_15_), .A2(n541), .A3(b_15_), .ZN(n539) );
  OR2_X1 U561 ( .A1(a_14_), .A2(b_14_), .ZN(n541) );
  INV_X1 U562 ( .A(a_12_), .ZN(n532) );
  INV_X1 U563 ( .A(a_11_), .ZN(n528) );
  INV_X1 U564 ( .A(a_10_), .ZN(n524) );
  INV_X1 U565 ( .A(a_9_), .ZN(n520) );
  INV_X1 U566 ( .A(a_8_), .ZN(n516) );
  INV_X1 U567 ( .A(a_7_), .ZN(n512) );
  INV_X1 U568 ( .A(a_6_), .ZN(n508) );
  INV_X1 U569 ( .A(a_5_), .ZN(n504) );
  INV_X1 U570 ( .A(a_4_), .ZN(n500) );
  INV_X1 U571 ( .A(a_3_), .ZN(n496) );
  INV_X1 U572 ( .A(a_2_), .ZN(n492) );
  AND2_X1 U573 ( .A1(n484), .A2(n542), .ZN(n426) );
  OR2_X1 U574 ( .A1(n543), .A2(b_0_), .ZN(n542) );
  INV_X1 U575 ( .A(a_0_), .ZN(n543) );
  OR2_X1 U576 ( .A1(a_0_), .A2(n456), .ZN(n484) );
  INV_X1 U577 ( .A(b_0_), .ZN(n456) );
endmodule

