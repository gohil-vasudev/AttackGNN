module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n342_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n393_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n257_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n381_, new_n388_, new_n508_, new_n194_, new_n299_, new_n142_, new_n139_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n178_, new_n295_, new_n359_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n562_, new_n525_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n598_, new_n570_, new_n143_, new_n520_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n605_, new_n182_, new_n407_, new_n480_, new_n625_, new_n151_, new_n513_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n417_, new_n591_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n550_, new_n217_, new_n269_, new_n512_, new_n412_, new_n327_, new_n561_, new_n495_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n200_, new_n422_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n138_, N1 );
xnor g001 ( new_n139_, N65, N69 );
xnor g002 ( new_n140_, new_n139_, keyIn_0_5 );
xnor g003 ( new_n141_, N73, N77 );
xnor g004 ( new_n142_, new_n141_, keyIn_0_6 );
nand g005 ( new_n143_, new_n140_, new_n142_ );
xor g006 ( new_n144_, new_n139_, keyIn_0_5 );
xor g007 ( new_n145_, new_n141_, keyIn_0_6 );
nand g008 ( new_n146_, new_n144_, new_n145_ );
nand g009 ( new_n147_, new_n146_, new_n143_ );
xnor g010 ( new_n148_, N81, N85 );
xnor g011 ( new_n149_, N89, N93 );
xnor g012 ( new_n150_, new_n148_, new_n149_ );
not g013 ( new_n151_, new_n150_ );
xnor g014 ( new_n152_, new_n147_, new_n151_ );
not g015 ( new_n153_, new_n152_ );
nand g016 ( new_n154_, N129, N137 );
nand g017 ( new_n155_, new_n153_, new_n154_ );
nand g018 ( new_n156_, new_n152_, N129, N137 );
nand g019 ( new_n157_, new_n155_, new_n156_ );
xnor g020 ( new_n158_, N1, N17 );
xnor g021 ( new_n159_, N33, N49 );
xnor g022 ( new_n160_, new_n158_, new_n159_ );
nand g023 ( new_n161_, new_n157_, new_n160_ );
not g024 ( new_n162_, new_n160_ );
nand g025 ( new_n163_, new_n155_, new_n156_, new_n162_ );
nand g026 ( new_n164_, new_n161_, new_n163_ );
not g027 ( new_n165_, new_n164_ );
xnor g028 ( new_n166_, N97, N101 );
xnor g029 ( new_n167_, N105, N109 );
xor g030 ( new_n168_, new_n166_, new_n167_ );
nand g031 ( new_n169_, new_n168_, keyIn_0_18 );
not g032 ( new_n170_, keyIn_0_18 );
xnor g033 ( new_n171_, new_n166_, new_n167_ );
nand g034 ( new_n172_, new_n171_, new_n170_ );
nand g035 ( new_n173_, new_n169_, new_n172_ );
nand g036 ( new_n174_, new_n173_, new_n147_ );
nand g037 ( new_n175_, new_n169_, new_n146_, new_n143_, new_n172_ );
nand g038 ( new_n176_, new_n174_, new_n175_ );
nand g039 ( new_n177_, new_n176_, N131, N137 );
nand g040 ( new_n178_, N131, N137 );
nand g041 ( new_n179_, new_n174_, new_n175_, new_n178_ );
nand g042 ( new_n180_, new_n177_, new_n179_ );
xnor g043 ( new_n181_, N9, N25 );
xnor g044 ( new_n182_, N41, N57 );
xnor g045 ( new_n183_, new_n181_, new_n182_ );
not g046 ( new_n184_, new_n183_ );
nand g047 ( new_n185_, new_n180_, new_n184_ );
nand g048 ( new_n186_, new_n177_, new_n179_, new_n183_ );
nand g049 ( new_n187_, new_n185_, new_n186_ );
nand g050 ( new_n188_, new_n187_, keyIn_0_24 );
not g051 ( new_n189_, keyIn_0_24 );
nand g052 ( new_n190_, new_n185_, new_n189_, new_n186_ );
nand g053 ( new_n191_, new_n188_, new_n190_ );
nand g054 ( new_n192_, new_n191_, keyIn_0_26 );
not g055 ( new_n193_, keyIn_0_26 );
nand g056 ( new_n194_, new_n188_, new_n193_, new_n190_ );
nand g057 ( new_n195_, new_n192_, new_n194_ );
not g058 ( new_n196_, keyIn_0_19 );
xnor g059 ( new_n197_, N121, N125 );
xnor g060 ( new_n198_, new_n197_, keyIn_0_7 );
xor g061 ( new_n199_, N113, N117 );
not g062 ( new_n200_, new_n199_ );
nand g063 ( new_n201_, new_n198_, new_n200_ );
not g064 ( new_n202_, keyIn_0_7 );
xnor g065 ( new_n203_, new_n197_, new_n202_ );
nand g066 ( new_n204_, new_n203_, new_n199_ );
nand g067 ( new_n205_, new_n201_, new_n204_, new_n196_ );
nand g068 ( new_n206_, new_n201_, new_n204_ );
nand g069 ( new_n207_, new_n206_, keyIn_0_19 );
nand g070 ( new_n208_, new_n207_, new_n205_ );
xnor g071 ( new_n209_, new_n208_, new_n150_ );
nand g072 ( new_n210_, N132, N137 );
xor g073 ( new_n211_, new_n210_, keyIn_0_9 );
nand g074 ( new_n212_, new_n209_, new_n211_ );
xnor g075 ( new_n213_, new_n208_, new_n151_ );
not g076 ( new_n214_, new_n211_ );
nand g077 ( new_n215_, new_n213_, new_n214_ );
nand g078 ( new_n216_, new_n212_, new_n215_, keyIn_0_23 );
not g079 ( new_n217_, keyIn_0_23 );
nand g080 ( new_n218_, new_n215_, new_n212_ );
nand g081 ( new_n219_, new_n218_, new_n217_ );
xnor g082 ( new_n220_, N13, N29 );
xnor g083 ( new_n221_, new_n220_, keyIn_0_14 );
xor g084 ( new_n222_, N45, N61 );
xnor g085 ( new_n223_, new_n221_, new_n222_ );
nand g086 ( new_n224_, new_n219_, new_n216_, new_n223_ );
nand g087 ( new_n225_, new_n219_, new_n216_ );
not g088 ( new_n226_, new_n223_ );
nand g089 ( new_n227_, new_n225_, new_n226_ );
nand g090 ( new_n228_, new_n227_, new_n224_ );
nand g091 ( new_n229_, new_n208_, new_n173_ );
nand g092 ( new_n230_, new_n207_, new_n169_, new_n172_, new_n205_ );
nand g093 ( new_n231_, new_n229_, new_n230_ );
nand g094 ( new_n232_, new_n231_, keyIn_0_22 );
not g095 ( new_n233_, keyIn_0_22 );
nand g096 ( new_n234_, new_n229_, new_n233_, new_n230_ );
nand g097 ( new_n235_, new_n232_, new_n234_ );
nand g098 ( new_n236_, N130, N137 );
xor g099 ( new_n237_, new_n236_, keyIn_0_8 );
not g100 ( new_n238_, new_n237_ );
nand g101 ( new_n239_, new_n235_, new_n238_ );
nand g102 ( new_n240_, new_n232_, new_n234_, new_n237_ );
nand g103 ( new_n241_, new_n239_, new_n240_ );
xnor g104 ( new_n242_, N5, N21 );
xnor g105 ( new_n243_, new_n242_, keyIn_0_12 );
xnor g106 ( new_n244_, N37, N53 );
xnor g107 ( new_n245_, new_n244_, keyIn_0_13 );
xnor g108 ( new_n246_, new_n243_, new_n245_ );
nand g109 ( new_n247_, new_n241_, new_n246_ );
not g110 ( new_n248_, new_n246_ );
nand g111 ( new_n249_, new_n239_, new_n240_, new_n248_ );
nand g112 ( new_n250_, new_n247_, new_n249_ );
nand g113 ( new_n251_, new_n250_, new_n165_ );
not g114 ( new_n252_, new_n251_ );
nand g115 ( new_n253_, new_n252_, keyIn_0_36, new_n195_, new_n228_ );
not g116 ( new_n254_, keyIn_0_36 );
nand g117 ( new_n255_, new_n195_, new_n228_, new_n165_, new_n250_ );
nand g118 ( new_n256_, new_n255_, new_n254_ );
nand g119 ( new_n257_, new_n256_, new_n253_ );
not g120 ( new_n258_, new_n191_ );
not g121 ( new_n259_, new_n250_ );
nand g122 ( new_n260_, new_n259_, new_n164_, new_n258_ );
not g123 ( new_n261_, keyIn_0_25 );
xnor g124 ( new_n262_, new_n164_, new_n261_ );
nand g125 ( new_n263_, new_n262_, new_n191_, new_n250_ );
nand g126 ( new_n264_, new_n260_, new_n263_ );
nand g127 ( new_n265_, new_n264_, new_n228_ );
not g128 ( new_n266_, new_n228_ );
nand g129 ( new_n267_, new_n266_, new_n164_, new_n258_, new_n250_ );
nand g130 ( new_n268_, new_n257_, new_n265_, new_n267_ );
not g131 ( new_n269_, keyIn_0_21 );
not g132 ( new_n270_, keyIn_0_17 );
not g133 ( new_n271_, keyIn_0_2 );
not g134 ( new_n272_, N33 );
not g135 ( new_n273_, N37 );
nand g136 ( new_n274_, new_n272_, new_n273_ );
nand g137 ( new_n275_, N33, N37 );
nand g138 ( new_n276_, new_n274_, new_n275_ );
nand g139 ( new_n277_, new_n276_, new_n271_ );
nand g140 ( new_n278_, new_n274_, keyIn_0_2, new_n275_ );
nand g141 ( new_n279_, new_n277_, new_n278_ );
xnor g142 ( new_n280_, N41, N45 );
nand g143 ( new_n281_, new_n280_, keyIn_0_3 );
not g144 ( new_n282_, keyIn_0_3 );
not g145 ( new_n283_, N41 );
not g146 ( new_n284_, N45 );
nand g147 ( new_n285_, new_n283_, new_n284_ );
nand g148 ( new_n286_, N41, N45 );
nand g149 ( new_n287_, new_n285_, new_n282_, new_n286_ );
nand g150 ( new_n288_, new_n281_, new_n287_ );
nand g151 ( new_n289_, new_n279_, new_n288_ );
nand g152 ( new_n290_, new_n277_, new_n281_, new_n278_, new_n287_ );
nand g153 ( new_n291_, new_n289_, new_n290_ );
nand g154 ( new_n292_, new_n291_, new_n270_ );
nand g155 ( new_n293_, new_n289_, keyIn_0_17, new_n290_ );
nand g156 ( new_n294_, new_n292_, new_n293_ );
xnor g157 ( new_n295_, N1, N5 );
xnor g158 ( new_n296_, N9, N13 );
nand g159 ( new_n297_, new_n295_, new_n296_ );
not g160 ( new_n298_, new_n295_ );
not g161 ( new_n299_, new_n296_ );
nand g162 ( new_n300_, new_n298_, new_n299_ );
nand g163 ( new_n301_, new_n300_, new_n297_ );
nand g164 ( new_n302_, new_n301_, keyIn_0_16 );
not g165 ( new_n303_, keyIn_0_16 );
nand g166 ( new_n304_, new_n300_, new_n303_, new_n297_ );
nand g167 ( new_n305_, new_n302_, new_n304_ );
nand g168 ( new_n306_, new_n294_, new_n305_ );
nand g169 ( new_n307_, new_n292_, new_n293_, new_n302_, new_n304_ );
nand g170 ( new_n308_, new_n306_, new_n307_ );
nand g171 ( new_n309_, new_n308_, new_n269_ );
nand g172 ( new_n310_, new_n306_, keyIn_0_21, new_n307_ );
nand g173 ( new_n311_, new_n309_, new_n310_ );
nand g174 ( new_n312_, N135, N137 );
xor g175 ( new_n313_, new_n312_, keyIn_0_10 );
nand g176 ( new_n314_, new_n311_, new_n313_ );
not g177 ( new_n315_, new_n313_ );
nand g178 ( new_n316_, new_n309_, new_n310_, new_n315_ );
nand g179 ( new_n317_, new_n314_, new_n316_ );
xnor g180 ( new_n318_, N73, N89 );
xnor g181 ( new_n319_, N105, N121 );
xnor g182 ( new_n320_, new_n318_, new_n319_ );
xor g183 ( new_n321_, new_n320_, keyIn_0_20 );
not g184 ( new_n322_, new_n321_ );
nand g185 ( new_n323_, new_n317_, new_n322_ );
nand g186 ( new_n324_, new_n314_, new_n316_, new_n321_ );
nand g187 ( new_n325_, new_n323_, new_n324_ );
nand g188 ( new_n326_, new_n268_, new_n325_ );
xnor g189 ( new_n327_, N57, N61 );
xnor g190 ( new_n328_, new_n327_, keyIn_0_4 );
xor g191 ( new_n329_, N49, N53 );
xnor g192 ( new_n330_, new_n328_, new_n329_ );
not g193 ( new_n331_, new_n330_ );
nand g194 ( new_n332_, new_n294_, new_n331_ );
nand g195 ( new_n333_, new_n330_, new_n292_, new_n293_ );
nand g196 ( new_n334_, new_n332_, new_n333_ );
nand g197 ( new_n335_, N134, N137 );
nand g198 ( new_n336_, new_n334_, new_n335_ );
nand g199 ( new_n337_, new_n332_, N134, N137, new_n333_ );
nand g200 ( new_n338_, new_n336_, new_n337_ );
xnor g201 ( new_n339_, N69, N85 );
xnor g202 ( new_n340_, N101, N117 );
xnor g203 ( new_n341_, new_n339_, new_n340_ );
nand g204 ( new_n342_, new_n338_, new_n341_ );
not g205 ( new_n343_, new_n341_ );
nand g206 ( new_n344_, new_n336_, new_n337_, new_n343_ );
nand g207 ( new_n345_, new_n342_, new_n344_ );
xnor g208 ( new_n346_, N17, N21 );
xnor g209 ( new_n347_, new_n346_, keyIn_0_0 );
xnor g210 ( new_n348_, N25, N29 );
xnor g211 ( new_n349_, new_n348_, keyIn_0_1 );
not g212 ( new_n350_, new_n349_ );
nand g213 ( new_n351_, new_n350_, new_n347_ );
not g214 ( new_n352_, new_n347_ );
nand g215 ( new_n353_, new_n352_, new_n349_ );
nand g216 ( new_n354_, new_n351_, new_n353_, new_n302_, new_n304_ );
nand g217 ( new_n355_, new_n351_, new_n353_ );
nand g218 ( new_n356_, new_n355_, new_n305_ );
nand g219 ( new_n357_, new_n356_, N133, N137, new_n354_ );
nand g220 ( new_n358_, new_n356_, new_n354_ );
nand g221 ( new_n359_, N133, N137 );
nand g222 ( new_n360_, new_n358_, new_n359_ );
xor g223 ( new_n361_, N97, N113 );
xnor g224 ( new_n362_, new_n361_, keyIn_0_15 );
xnor g225 ( new_n363_, N65, N81 );
xnor g226 ( new_n364_, new_n362_, new_n363_ );
nand g227 ( new_n365_, new_n360_, new_n357_, new_n364_ );
nand g228 ( new_n366_, new_n360_, new_n357_ );
not g229 ( new_n367_, new_n364_ );
nand g230 ( new_n368_, new_n366_, new_n367_ );
nand g231 ( new_n369_, new_n368_, new_n365_ );
not g232 ( new_n370_, new_n369_ );
nand g233 ( new_n371_, new_n331_, new_n355_ );
nand g234 ( new_n372_, new_n330_, new_n351_, new_n353_ );
nand g235 ( new_n373_, N136, N137 );
xnor g236 ( new_n374_, new_n373_, keyIn_0_11 );
nand g237 ( new_n375_, new_n371_, new_n372_, new_n374_ );
nand g238 ( new_n376_, new_n371_, new_n372_ );
not g239 ( new_n377_, new_n374_ );
nand g240 ( new_n378_, new_n376_, new_n377_ );
nand g241 ( new_n379_, new_n378_, new_n375_ );
xnor g242 ( new_n380_, N77, N93 );
xnor g243 ( new_n381_, N109, N125 );
xnor g244 ( new_n382_, new_n380_, new_n381_ );
nand g245 ( new_n383_, new_n379_, new_n382_ );
not g246 ( new_n384_, new_n382_ );
nand g247 ( new_n385_, new_n378_, new_n375_, new_n384_ );
nand g248 ( new_n386_, new_n383_, new_n385_ );
nand g249 ( new_n387_, new_n345_, new_n370_, new_n386_ );
nor g250 ( new_n388_, new_n326_, new_n387_ );
nand g251 ( new_n389_, new_n388_, new_n165_ );
xnor g252 ( new_n390_, new_n389_, keyIn_0_41 );
xnor g253 ( N724, new_n390_, new_n138_ );
nand g254 ( new_n392_, new_n388_, new_n259_ );
xnor g255 ( new_n393_, new_n392_, keyIn_0_42 );
xnor g256 ( N725, new_n393_, N5 );
nand g257 ( new_n395_, new_n388_, new_n191_ );
xnor g258 ( N726, new_n395_, N9 );
nand g259 ( new_n397_, new_n388_, new_n266_ );
xnor g260 ( N727, new_n397_, N13 );
not g261 ( new_n399_, keyIn_0_54 );
not g262 ( new_n400_, N17 );
nand g263 ( new_n401_, new_n370_, new_n345_ );
not g264 ( new_n402_, new_n386_ );
nand g265 ( new_n403_, new_n268_, new_n402_ );
nor g266 ( new_n404_, new_n403_, new_n325_, new_n401_ );
nand g267 ( new_n405_, new_n404_, new_n165_ );
xnor g268 ( new_n406_, new_n405_, new_n400_ );
nand g269 ( new_n407_, new_n406_, new_n399_ );
xnor g270 ( new_n408_, new_n405_, N17 );
nand g271 ( new_n409_, new_n408_, keyIn_0_54 );
nand g272 ( N728, new_n407_, new_n409_ );
not g273 ( new_n411_, keyIn_0_55 );
not g274 ( new_n412_, N21 );
nand g275 ( new_n413_, new_n404_, new_n259_ );
xnor g276 ( new_n414_, new_n413_, new_n412_ );
nand g277 ( new_n415_, new_n414_, new_n411_ );
xnor g278 ( new_n416_, new_n413_, N21 );
nand g279 ( new_n417_, new_n416_, keyIn_0_55 );
nand g280 ( N729, new_n415_, new_n417_ );
nand g281 ( new_n419_, new_n404_, new_n191_ );
xnor g282 ( N730, new_n419_, N25 );
not g283 ( new_n421_, N29 );
nand g284 ( new_n422_, new_n404_, new_n266_ );
xnor g285 ( new_n423_, new_n422_, keyIn_0_43 );
nand g286 ( new_n424_, new_n423_, new_n421_ );
not g287 ( new_n425_, keyIn_0_43 );
xnor g288 ( new_n426_, new_n422_, new_n425_ );
nand g289 ( new_n427_, new_n426_, N29 );
nand g290 ( N731, new_n424_, new_n427_ );
not g291 ( new_n429_, new_n345_ );
nand g292 ( new_n430_, new_n429_, new_n369_, new_n386_ );
nor g293 ( new_n431_, new_n326_, new_n430_ );
nand g294 ( new_n432_, new_n431_, new_n165_ );
xnor g295 ( new_n433_, new_n432_, N33 );
xnor g296 ( N732, new_n433_, keyIn_0_56 );
nand g297 ( new_n435_, new_n431_, new_n259_ );
xnor g298 ( new_n436_, new_n435_, new_n273_ );
xnor g299 ( N733, new_n436_, keyIn_0_57 );
nor g300 ( new_n438_, new_n326_, new_n258_, new_n430_ );
xnor g301 ( new_n439_, new_n438_, keyIn_0_44 );
xnor g302 ( N734, new_n439_, N41 );
not g303 ( new_n441_, new_n430_ );
nand g304 ( new_n442_, new_n268_, new_n266_, new_n325_, new_n441_ );
xnor g305 ( new_n443_, new_n442_, keyIn_0_45 );
nand g306 ( new_n444_, new_n443_, new_n284_ );
not g307 ( new_n445_, keyIn_0_45 );
xnor g308 ( new_n446_, new_n442_, new_n445_ );
nand g309 ( new_n447_, new_n446_, N45 );
nand g310 ( new_n448_, new_n444_, new_n447_ );
nand g311 ( new_n449_, new_n448_, keyIn_0_58 );
not g312 ( new_n450_, keyIn_0_58 );
nand g313 ( new_n451_, new_n444_, new_n447_, new_n450_ );
nand g314 ( N735, new_n449_, new_n451_ );
not g315 ( new_n453_, keyIn_0_59 );
not g316 ( new_n454_, N49 );
not g317 ( new_n455_, keyIn_0_39 );
not g318 ( new_n456_, keyIn_0_27 );
nand g319 ( new_n457_, new_n325_, new_n456_ );
not g320 ( new_n458_, new_n457_ );
nand g321 ( new_n459_, new_n323_, keyIn_0_27, new_n324_ );
nand g322 ( new_n460_, new_n459_, new_n429_, new_n369_ );
nor g323 ( new_n461_, new_n458_, new_n460_ );
nand g324 ( new_n462_, new_n268_, new_n402_, new_n461_ );
nand g325 ( new_n463_, new_n462_, new_n455_ );
nand g326 ( new_n464_, new_n268_, keyIn_0_39, new_n402_, new_n461_ );
nand g327 ( new_n465_, new_n463_, new_n464_ );
nand g328 ( new_n466_, new_n465_, new_n165_ );
nand g329 ( new_n467_, new_n466_, new_n454_ );
nand g330 ( new_n468_, new_n465_, N49, new_n165_ );
nand g331 ( new_n469_, new_n467_, new_n468_ );
nand g332 ( new_n470_, new_n469_, new_n453_ );
nand g333 ( new_n471_, new_n467_, keyIn_0_59, new_n468_ );
nand g334 ( N736, new_n470_, new_n471_ );
not g335 ( new_n473_, N53 );
not g336 ( new_n474_, keyIn_0_46 );
nand g337 ( new_n475_, new_n465_, new_n259_ );
nand g338 ( new_n476_, new_n475_, new_n474_ );
nand g339 ( new_n477_, new_n465_, keyIn_0_46, new_n259_ );
nand g340 ( new_n478_, new_n476_, new_n477_ );
nand g341 ( new_n479_, new_n478_, new_n473_ );
nand g342 ( new_n480_, new_n476_, N53, new_n477_ );
nand g343 ( N737, new_n479_, new_n480_ );
nand g344 ( new_n482_, new_n465_, new_n191_ );
xnor g345 ( N738, new_n482_, N57 );
nand g346 ( new_n484_, new_n465_, new_n266_ );
xnor g347 ( N739, new_n484_, N61 );
not g348 ( new_n486_, keyIn_0_47 );
not g349 ( new_n487_, keyIn_0_40 );
not g350 ( new_n488_, keyIn_0_31 );
nand g351 ( new_n489_, new_n323_, new_n488_, new_n324_ );
nand g352 ( new_n490_, new_n325_, keyIn_0_31 );
nand g353 ( new_n491_, new_n490_, new_n441_, new_n489_ );
nand g354 ( new_n492_, new_n491_, keyIn_0_37 );
not g355 ( new_n493_, keyIn_0_37 );
nand g356 ( new_n494_, new_n490_, new_n441_, new_n493_, new_n489_ );
not g357 ( new_n495_, keyIn_0_32 );
nand g358 ( new_n496_, new_n325_, new_n495_ );
nand g359 ( new_n497_, new_n323_, keyIn_0_32, new_n324_ );
nand g360 ( new_n498_, new_n496_, new_n497_ );
xnor g361 ( new_n499_, new_n386_, keyIn_0_33 );
nor g362 ( new_n500_, new_n499_, new_n401_ );
nand g363 ( new_n501_, new_n498_, new_n500_ );
not g364 ( new_n502_, keyIn_0_28 );
nand g365 ( new_n503_, new_n345_, new_n502_ );
nand g366 ( new_n504_, new_n342_, keyIn_0_28, new_n344_ );
nand g367 ( new_n505_, new_n503_, new_n504_ );
nor g368 ( new_n506_, new_n370_, new_n386_ );
nand g369 ( new_n507_, new_n505_, new_n506_, new_n323_, new_n324_ );
xnor g370 ( new_n508_, new_n386_, keyIn_0_30 );
xnor g371 ( new_n509_, new_n369_, keyIn_0_29 );
nand g372 ( new_n510_, new_n508_, new_n325_, new_n345_, new_n509_ );
nand g373 ( new_n511_, new_n510_, new_n507_ );
not g374 ( new_n512_, new_n511_ );
nand g375 ( new_n513_, new_n512_, new_n492_, new_n494_, new_n501_ );
nand g376 ( new_n514_, new_n513_, keyIn_0_38 );
not g377 ( new_n515_, keyIn_0_38 );
not g378 ( new_n516_, new_n501_ );
nor g379 ( new_n517_, new_n516_, new_n511_ );
nand g380 ( new_n518_, new_n517_, new_n515_, new_n492_, new_n494_ );
nand g381 ( new_n519_, new_n252_, new_n191_, new_n228_ );
not g382 ( new_n520_, new_n519_ );
nand g383 ( new_n521_, new_n518_, new_n487_, new_n514_, new_n520_ );
nand g384 ( new_n522_, new_n518_, new_n514_, new_n520_ );
nand g385 ( new_n523_, new_n522_, keyIn_0_40 );
nand g386 ( new_n524_, new_n523_, new_n521_ );
nand g387 ( new_n525_, new_n524_, new_n370_ );
nand g388 ( new_n526_, new_n525_, new_n486_ );
nand g389 ( new_n527_, new_n524_, keyIn_0_47, new_n370_ );
nand g390 ( new_n528_, new_n526_, new_n527_ );
nand g391 ( new_n529_, new_n528_, N65 );
not g392 ( new_n530_, N65 );
nand g393 ( new_n531_, new_n526_, new_n530_, new_n527_ );
nand g394 ( N740, new_n529_, new_n531_ );
not g395 ( new_n533_, keyIn_0_48 );
nand g396 ( new_n534_, new_n524_, new_n429_ );
nand g397 ( new_n535_, new_n534_, new_n533_ );
nand g398 ( new_n536_, new_n524_, keyIn_0_48, new_n429_ );
nand g399 ( new_n537_, new_n535_, new_n536_ );
nand g400 ( new_n538_, new_n537_, N69 );
not g401 ( new_n539_, N69 );
nand g402 ( new_n540_, new_n535_, new_n539_, new_n536_ );
nand g403 ( N741, new_n538_, new_n540_ );
nand g404 ( new_n542_, new_n524_, new_n325_ );
xnor g405 ( N742, new_n542_, N73 );
not g406 ( new_n544_, keyIn_0_60 );
not g407 ( new_n545_, N77 );
nand g408 ( new_n546_, new_n524_, new_n402_ );
nand g409 ( new_n547_, new_n546_, new_n545_ );
nand g410 ( new_n548_, new_n524_, N77, new_n402_ );
nand g411 ( new_n549_, new_n547_, new_n548_ );
nand g412 ( new_n550_, new_n549_, new_n544_ );
nand g413 ( new_n551_, new_n547_, keyIn_0_60, new_n548_ );
nand g414 ( N743, new_n550_, new_n551_ );
nand g415 ( new_n553_, new_n518_, new_n514_ );
xnor g416 ( new_n554_, new_n250_, keyIn_0_34 );
nand g417 ( new_n555_, new_n554_, new_n165_, new_n258_, new_n266_ );
nor g418 ( new_n556_, new_n553_, new_n555_ );
nand g419 ( new_n557_, new_n556_, new_n370_ );
xnor g420 ( N744, new_n557_, N81 );
not g421 ( new_n559_, N85 );
not g422 ( new_n560_, keyIn_0_49 );
nand g423 ( new_n561_, new_n556_, new_n429_ );
xnor g424 ( new_n562_, new_n561_, new_n560_ );
nand g425 ( new_n563_, new_n562_, new_n559_ );
xnor g426 ( new_n564_, new_n561_, keyIn_0_49 );
nand g427 ( new_n565_, new_n564_, N85 );
nand g428 ( N745, new_n563_, new_n565_ );
not g429 ( new_n567_, keyIn_0_61 );
not g430 ( new_n568_, N89 );
nand g431 ( new_n569_, new_n556_, new_n325_ );
xnor g432 ( new_n570_, new_n569_, new_n568_ );
nand g433 ( new_n571_, new_n570_, new_n567_ );
xnor g434 ( new_n572_, new_n569_, N89 );
nand g435 ( new_n573_, new_n572_, keyIn_0_61 );
nand g436 ( N746, new_n571_, new_n573_ );
nand g437 ( new_n575_, new_n556_, new_n402_ );
xnor g438 ( N747, new_n575_, N93 );
xor g439 ( new_n577_, new_n164_, keyIn_0_35 );
nand g440 ( new_n578_, new_n577_, new_n191_, new_n259_ );
nor g441 ( new_n579_, new_n553_, new_n266_, new_n578_ );
nand g442 ( new_n580_, new_n579_, new_n370_ );
xnor g443 ( N748, new_n580_, N97 );
nand g444 ( new_n582_, new_n579_, new_n429_ );
nand g445 ( new_n583_, new_n582_, keyIn_0_50 );
not g446 ( new_n584_, keyIn_0_50 );
nand g447 ( new_n585_, new_n579_, new_n584_, new_n429_ );
nand g448 ( new_n586_, new_n583_, new_n585_ );
nand g449 ( new_n587_, new_n586_, N101 );
not g450 ( new_n588_, N101 );
nand g451 ( new_n589_, new_n583_, new_n588_, new_n585_ );
nand g452 ( N749, new_n587_, new_n589_ );
nand g453 ( new_n591_, new_n579_, new_n325_ );
xnor g454 ( N750, new_n591_, N105 );
nand g455 ( new_n593_, new_n579_, new_n402_ );
xnor g456 ( N751, new_n593_, N109 );
nor g457 ( new_n595_, new_n260_, new_n228_ );
not g458 ( new_n596_, new_n595_ );
nor g459 ( new_n597_, new_n553_, new_n596_ );
nand g460 ( new_n598_, new_n597_, new_n370_ );
xnor g461 ( N752, new_n598_, N113 );
not g462 ( new_n600_, keyIn_0_51 );
nand g463 ( new_n601_, new_n597_, new_n429_ );
xnor g464 ( new_n602_, new_n601_, new_n600_ );
nand g465 ( new_n603_, new_n602_, N117 );
not g466 ( new_n604_, N117 );
xnor g467 ( new_n605_, new_n601_, keyIn_0_51 );
nand g468 ( new_n606_, new_n605_, new_n604_ );
nand g469 ( N753, new_n603_, new_n606_ );
nand g470 ( new_n608_, new_n518_, new_n325_, new_n514_, new_n595_ );
xnor g471 ( new_n609_, new_n608_, keyIn_0_52 );
nand g472 ( new_n610_, new_n609_, N121 );
not g473 ( new_n611_, N121 );
not g474 ( new_n612_, keyIn_0_52 );
xnor g475 ( new_n613_, new_n608_, new_n612_ );
nand g476 ( new_n614_, new_n613_, new_n611_ );
nand g477 ( new_n615_, new_n610_, new_n614_ );
nand g478 ( new_n616_, new_n615_, keyIn_0_62 );
not g479 ( new_n617_, keyIn_0_62 );
nand g480 ( new_n618_, new_n610_, new_n614_, new_n617_ );
nand g481 ( N754, new_n616_, new_n618_ );
not g482 ( new_n620_, keyIn_0_53 );
nand g483 ( new_n621_, new_n518_, new_n402_, new_n514_, new_n595_ );
xnor g484 ( new_n622_, new_n621_, new_n620_ );
nand g485 ( new_n623_, new_n622_, N125 );
not g486 ( new_n624_, N125 );
xnor g487 ( new_n625_, new_n621_, keyIn_0_53 );
nand g488 ( new_n626_, new_n625_, new_n624_ );
nand g489 ( new_n627_, new_n623_, new_n626_ );
nand g490 ( new_n628_, new_n627_, keyIn_0_63 );
not g491 ( new_n629_, keyIn_0_63 );
nand g492 ( new_n630_, new_n623_, new_n626_, new_n629_ );
nand g493 ( N755, new_n628_, new_n630_ );
endmodule