module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n1215_, new_n1249_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n1157_, new_n798_, new_n1180_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n1232_, new_n241_, new_n1025_, new_n566_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n1176_, new_n1207_, new_n1211_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1237_, new_n1172_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n1210_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n1213_, new_n840_, new_n735_, new_n1045_, new_n1132_, new_n500_, new_n898_, new_n1163_, new_n786_, new_n799_, new_n946_, new_n317_, new_n1188_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n1167_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n1238_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n1162_, new_n481_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n282_, new_n1212_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n1250_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1151_, new_n1082_, new_n849_, new_n1203_, new_n1018_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n385_, new_n1049_, new_n829_, new_n1257_, new_n988_, new_n478_, new_n694_, new_n461_, new_n1228_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n1196_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n517_, new_n325_, new_n609_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n1216_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n568_, new_n1051_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n1182_, new_n1200_, new_n650_, new_n708_, new_n750_, new_n1217_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n1222_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n1226_, new_n778_, new_n452_, new_n1198_, new_n381_, new_n1219_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1168_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n1241_, new_n882_, new_n1145_, new_n657_, new_n1150_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1159_, new_n1020_, new_n363_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n1041_, new_n917_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n1177_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n1026_, new_n1106_, new_n267_, new_n473_, new_n1147_, new_n1229_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n1247_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n1234_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n943_, new_n874_, new_n1245_, new_n402_, new_n663_, new_n579_, new_n286_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n1254_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n1218_, new_n870_, new_n945_, new_n1115_, new_n559_, new_n1201_, new_n948_, new_n1231_, new_n762_, new_n1055_, new_n1193_, new_n838_, new_n1233_, new_n923_, new_n233_, new_n1187_, new_n469_, new_n1205_, new_n391_, new_n1154_, new_n437_, new_n1085_, new_n1253_, new_n295_, new_n1256_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n1169_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n1171_, new_n688_, new_n1255_, new_n384_, new_n900_, new_n1161_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n1096_, new_n454_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n1160_, new_n809_, new_n1142_, new_n654_, new_n1166_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n328_, new_n460_, new_n1136_, new_n693_, new_n1175_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n1135_, new_n376_, new_n380_, new_n1251_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n310_, new_n1095_, new_n1252_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n1178_, new_n224_, new_n586_, new_n963_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n1191_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n1242_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1224_, new_n1137_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n1186_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n225_, new_n1040_, new_n1246_, new_n922_, new_n387_, new_n544_, new_n476_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n1179_, new_n298_, new_n499_, new_n255_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n1185_, new_n1240_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n1174_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n337_, new_n623_, new_n446_, new_n1195_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n1227_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n1248_, new_n751_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n1244_, new_n1181_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n1072_, new_n769_, new_n1190_, new_n1097_, new_n651_, new_n433_, new_n1164_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n788_, new_n841_, new_n1220_, new_n989_, new_n1204_, new_n1117_, new_n1112_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n1206_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n1258_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n1173_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1189_, new_n1153_, new_n357_, new_n1197_, new_n780_, new_n984_, new_n1183_, new_n643_, new_n474_, new_n1223_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1194_, new_n1077_, new_n1243_, new_n560_, new_n1100_, new_n1230_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n1165_, new_n1259_, new_n425_, new_n896_, new_n226_, new_n802_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n1236_, new_n709_, new_n373_, new_n866_, new_n1235_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1225_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n889_, new_n536_, new_n464_, new_n1089_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g0000 ( new_n215_, N75 );
nand g0001 ( new_n216_, N29, N42 );
nor g0002 ( N388, new_n216_, new_n215_ );
not g0003 ( new_n218_, N80 );
nand g0004 ( new_n219_, N29, N36 );
nor g0005 ( N389, new_n219_, new_n218_ );
not g0006 ( new_n221_, keyIn_0_6 );
not g0007 ( new_n222_, N42 );
nor g0008 ( new_n223_, new_n219_, new_n222_ );
nand g0009 ( new_n224_, new_n223_, new_n221_ );
not g0010 ( new_n225_, new_n223_ );
nand g0011 ( new_n226_, new_n225_, keyIn_0_6 );
nand g0012 ( N390, new_n226_, new_n224_ );
nand g0013 ( new_n228_, N85, N86 );
not g0014 ( N391, new_n228_ );
not g0015 ( new_n230_, N17 );
nand g0016 ( new_n231_, N1, N8 );
not g0017 ( new_n232_, new_n231_ );
nand g0018 ( new_n233_, new_n232_, N13 );
nor g0019 ( N418, new_n233_, new_n230_ );
nand g0020 ( new_n235_, N1, N26 );
nand g0021 ( new_n236_, N13, N17 );
nor g0022 ( new_n237_, new_n235_, new_n236_ );
not g0023 ( new_n238_, keyIn_0_0 );
nor g0024 ( new_n239_, new_n225_, new_n238_ );
nor g0025 ( new_n240_, new_n223_, keyIn_0_0 );
nor g0026 ( new_n241_, new_n239_, new_n240_ );
nand g0027 ( N419, new_n241_, new_n237_ );
nand g0028 ( new_n243_, N59, N75 );
not g0029 ( new_n244_, new_n243_ );
nand g0030 ( N420, new_n244_, N80 );
nand g0031 ( new_n246_, N36, N59 );
nor g0032 ( new_n247_, new_n246_, new_n218_ );
nor g0033 ( new_n248_, new_n247_, keyIn_0_8 );
nand g0034 ( new_n249_, new_n247_, keyIn_0_8 );
not g0035 ( new_n250_, new_n249_ );
nor g0036 ( new_n251_, new_n250_, new_n248_ );
not g0037 ( new_n252_, new_n251_ );
nand g0038 ( new_n253_, new_n252_, keyIn_0_19 );
not g0039 ( new_n254_, keyIn_0_19 );
nand g0040 ( new_n255_, new_n251_, new_n254_ );
nand g0041 ( N421, new_n253_, new_n255_ );
not g0042 ( new_n257_, keyIn_0_9 );
nor g0043 ( new_n258_, new_n246_, new_n222_ );
not g0044 ( new_n259_, new_n258_ );
nand g0045 ( new_n260_, new_n259_, new_n257_ );
nand g0046 ( new_n261_, new_n258_, keyIn_0_9 );
nand g0047 ( N422, new_n260_, new_n261_ );
nor g0048 ( new_n263_, N87, N88 );
not g0049 ( new_n264_, new_n263_ );
nand g0050 ( new_n265_, new_n264_, N90 );
nand g0051 ( new_n266_, new_n265_, keyIn_0_20 );
not g0052 ( new_n267_, keyIn_0_20 );
not g0053 ( new_n268_, new_n265_ );
nand g0054 ( new_n269_, new_n268_, new_n267_ );
nand g0055 ( N423, new_n269_, new_n266_ );
not g0056 ( new_n271_, new_n241_ );
nand g0057 ( N446, new_n271_, new_n237_ );
not g0058 ( new_n273_, keyIn_0_1 );
not g0059 ( new_n274_, new_n235_ );
nand g0060 ( new_n275_, new_n274_, N51 );
nand g0061 ( new_n276_, new_n275_, new_n273_ );
not g0062 ( new_n277_, N51 );
nor g0063 ( new_n278_, new_n235_, new_n277_ );
nand g0064 ( new_n279_, new_n278_, keyIn_0_1 );
nand g0065 ( N447, new_n276_, new_n279_ );
not g0066 ( new_n281_, keyIn_0_27 );
not g0067 ( new_n282_, keyIn_0_3 );
not g0068 ( new_n283_, N55 );
nor g0069 ( new_n284_, new_n233_, new_n283_ );
not g0070 ( new_n285_, new_n284_ );
nand g0071 ( new_n286_, new_n285_, new_n282_ );
not g0072 ( new_n287_, new_n286_ );
nor g0073 ( new_n288_, new_n285_, new_n282_ );
nor g0074 ( new_n289_, new_n287_, new_n288_ );
nand g0075 ( new_n290_, N29, N68 );
nand g0076 ( new_n291_, new_n290_, keyIn_0_4 );
not g0077 ( new_n292_, N29 );
nor g0078 ( new_n293_, new_n292_, keyIn_0_4 );
nand g0079 ( new_n294_, new_n293_, N68 );
nand g0080 ( new_n295_, new_n294_, new_n291_ );
nor g0081 ( new_n296_, new_n289_, new_n295_ );
not g0082 ( new_n297_, new_n296_ );
nand g0083 ( new_n298_, new_n297_, new_n281_ );
nand g0084 ( new_n299_, new_n296_, keyIn_0_27 );
nand g0085 ( N448, new_n298_, new_n299_ );
nand g0086 ( new_n301_, N59, N68 );
not g0087 ( new_n302_, new_n301_ );
nand g0088 ( new_n303_, new_n302_, N74 );
not g0089 ( new_n304_, new_n303_ );
nor g0090 ( new_n305_, new_n304_, keyIn_0_5 );
nand g0091 ( new_n306_, new_n304_, keyIn_0_5 );
not g0092 ( new_n307_, new_n306_ );
nor g0093 ( new_n308_, new_n307_, new_n305_ );
nor g0094 ( new_n309_, new_n289_, new_n308_ );
not g0095 ( new_n310_, new_n309_ );
nand g0096 ( new_n311_, new_n310_, keyIn_0_28 );
not g0097 ( new_n312_, keyIn_0_28 );
nand g0098 ( new_n313_, new_n309_, new_n312_ );
nand g0099 ( N449, new_n311_, new_n313_ );
nand g0100 ( new_n315_, new_n264_, N89 );
nand g0101 ( new_n316_, new_n315_, keyIn_0_29 );
not g0102 ( new_n317_, keyIn_0_29 );
not g0103 ( new_n318_, new_n315_ );
nand g0104 ( new_n319_, new_n318_, new_n317_ );
nand g0105 ( N450, new_n319_, new_n316_ );
not g0106 ( new_n321_, N130 );
not g0107 ( new_n322_, keyIn_0_22 );
not g0108 ( new_n323_, keyIn_0_11 );
nor g0109 ( new_n324_, N101, N106 );
nor g0110 ( new_n325_, new_n324_, new_n323_ );
nand g0111 ( new_n326_, new_n324_, new_n323_ );
not g0112 ( new_n327_, new_n326_ );
nor g0113 ( new_n328_, new_n327_, new_n325_ );
nand g0114 ( new_n329_, N101, N106 );
nand g0115 ( new_n330_, new_n329_, keyIn_0_10 );
not g0116 ( new_n331_, new_n330_ );
nor g0117 ( new_n332_, new_n329_, keyIn_0_10 );
nor g0118 ( new_n333_, new_n331_, new_n332_ );
nand g0119 ( new_n334_, new_n328_, new_n333_ );
not g0120 ( new_n335_, new_n334_ );
nor g0121 ( new_n336_, new_n335_, new_n322_ );
nor g0122 ( new_n337_, new_n334_, keyIn_0_22 );
nor g0123 ( new_n338_, new_n336_, new_n337_ );
not g0124 ( new_n339_, new_n338_ );
not g0125 ( new_n340_, N91 );
nor g0126 ( new_n341_, new_n340_, N96 );
not g0127 ( new_n342_, N96 );
nor g0128 ( new_n343_, new_n342_, N91 );
nor g0129 ( new_n344_, new_n341_, new_n343_ );
not g0130 ( new_n345_, new_n344_ );
nand g0131 ( new_n346_, new_n345_, keyIn_0_21 );
not g0132 ( new_n347_, new_n346_ );
nor g0133 ( new_n348_, new_n345_, keyIn_0_21 );
nor g0134 ( new_n349_, new_n347_, new_n348_ );
not g0135 ( new_n350_, new_n349_ );
nand g0136 ( new_n351_, new_n339_, new_n350_ );
nor g0137 ( new_n352_, new_n351_, keyIn_0_30 );
nand g0138 ( new_n353_, new_n351_, keyIn_0_30 );
nand g0139 ( new_n354_, new_n338_, new_n349_ );
nand g0140 ( new_n355_, new_n353_, new_n354_ );
nor g0141 ( new_n356_, new_n355_, new_n352_ );
not g0142 ( new_n357_, new_n356_ );
nor g0143 ( new_n358_, new_n357_, new_n321_ );
not g0144 ( new_n359_, new_n358_ );
nand g0145 ( new_n360_, new_n359_, keyIn_0_44 );
not g0146 ( new_n361_, new_n360_ );
nor g0147 ( new_n362_, new_n356_, N130 );
nor g0148 ( new_n363_, new_n362_, keyIn_0_45 );
nor g0149 ( new_n364_, new_n361_, new_n363_ );
nand g0150 ( new_n365_, new_n362_, keyIn_0_45 );
not g0151 ( new_n366_, new_n365_ );
nor g0152 ( new_n367_, new_n359_, keyIn_0_44 );
nor g0153 ( new_n368_, new_n367_, new_n366_ );
nand g0154 ( new_n369_, new_n364_, new_n368_ );
not g0155 ( new_n370_, new_n369_ );
nand g0156 ( new_n371_, new_n370_, keyIn_0_57 );
not g0157 ( new_n372_, keyIn_0_57 );
nand g0158 ( new_n373_, new_n369_, new_n372_ );
nand g0159 ( new_n374_, new_n371_, new_n373_ );
not g0160 ( new_n375_, keyIn_0_46 );
not g0161 ( new_n376_, keyIn_0_23 );
nor g0162 ( new_n377_, N111, N116 );
nand g0163 ( new_n378_, N111, N116 );
not g0164 ( new_n379_, new_n378_ );
nor g0165 ( new_n380_, new_n379_, new_n377_ );
nor g0166 ( new_n381_, new_n380_, new_n376_ );
nand g0167 ( new_n382_, new_n380_, new_n376_ );
not g0168 ( new_n383_, new_n382_ );
nor g0169 ( new_n384_, new_n383_, new_n381_ );
nor g0170 ( new_n385_, N121, N126 );
not g0171 ( new_n386_, new_n385_ );
nor g0172 ( new_n387_, new_n386_, keyIn_0_12 );
nand g0173 ( new_n388_, new_n386_, keyIn_0_12 );
not g0174 ( new_n389_, new_n388_ );
not g0175 ( new_n390_, keyIn_0_31 );
nand g0176 ( new_n391_, N121, N126 );
nand g0177 ( new_n392_, new_n391_, new_n390_ );
nor g0178 ( new_n393_, new_n389_, new_n392_ );
not g0179 ( new_n394_, new_n393_ );
nor g0180 ( new_n395_, new_n394_, new_n387_ );
nor g0181 ( new_n396_, new_n395_, new_n384_ );
nand g0182 ( new_n397_, new_n395_, new_n384_ );
not g0183 ( new_n398_, new_n397_ );
nor g0184 ( new_n399_, new_n398_, new_n396_ );
nor g0185 ( new_n400_, new_n399_, N135 );
not g0186 ( new_n401_, new_n400_ );
nand g0187 ( new_n402_, new_n401_, new_n375_ );
not g0188 ( new_n403_, new_n402_ );
nor g0189 ( new_n404_, new_n401_, new_n375_ );
nor g0190 ( new_n405_, new_n403_, new_n404_ );
nand g0191 ( new_n406_, new_n399_, N135 );
not g0192 ( new_n407_, new_n406_ );
nor g0193 ( new_n408_, new_n405_, new_n407_ );
not g0194 ( new_n409_, new_n408_ );
nand g0195 ( new_n410_, new_n409_, keyIn_0_53 );
not g0196 ( new_n411_, keyIn_0_53 );
nand g0197 ( new_n412_, new_n408_, new_n411_ );
nand g0198 ( new_n413_, new_n410_, new_n412_ );
nand g0199 ( new_n414_, new_n374_, new_n413_ );
nand g0200 ( new_n415_, new_n414_, keyIn_0_63 );
not g0201 ( new_n416_, new_n415_ );
nor g0202 ( new_n417_, new_n414_, keyIn_0_63 );
nor g0203 ( new_n418_, new_n416_, new_n417_ );
nor g0204 ( new_n419_, new_n370_, new_n413_ );
nor g0205 ( N767, new_n418_, new_n419_ );
not g0206 ( new_n421_, keyIn_0_64 );
not g0207 ( new_n422_, keyIn_0_62 );
not g0208 ( new_n423_, N207 );
not g0209 ( new_n424_, keyIn_0_25 );
nor g0210 ( new_n425_, N183, N189 );
nand g0211 ( new_n426_, N183, N189 );
not g0212 ( new_n427_, new_n426_ );
nor g0213 ( new_n428_, new_n427_, new_n425_ );
nor g0214 ( new_n429_, new_n428_, new_n424_ );
nand g0215 ( new_n430_, new_n428_, new_n424_ );
not g0216 ( new_n431_, new_n430_ );
nor g0217 ( new_n432_, new_n431_, new_n429_ );
not g0218 ( new_n433_, new_n432_ );
not g0219 ( new_n434_, N195 );
nor g0220 ( new_n435_, new_n434_, N201 );
not g0221 ( new_n436_, N201 );
nor g0222 ( new_n437_, new_n436_, N195 );
nor g0223 ( new_n438_, new_n435_, new_n437_ );
not g0224 ( new_n439_, new_n438_ );
nand g0225 ( new_n440_, new_n439_, keyIn_0_26 );
not g0226 ( new_n441_, new_n440_ );
nor g0227 ( new_n442_, new_n439_, keyIn_0_26 );
nor g0228 ( new_n443_, new_n441_, new_n442_ );
nor g0229 ( new_n444_, new_n443_, new_n433_ );
nand g0230 ( new_n445_, new_n443_, new_n433_ );
not g0231 ( new_n446_, new_n445_ );
nor g0232 ( new_n447_, new_n446_, new_n444_ );
nor g0233 ( new_n448_, new_n447_, new_n423_ );
not g0234 ( new_n449_, new_n448_ );
nor g0235 ( new_n450_, new_n449_, keyIn_0_51 );
nand g0236 ( new_n451_, new_n449_, keyIn_0_51 );
nand g0237 ( new_n452_, new_n447_, new_n423_ );
nand g0238 ( new_n453_, new_n451_, new_n452_ );
nor g0239 ( new_n454_, new_n453_, new_n450_ );
nand g0240 ( new_n455_, new_n454_, new_n422_ );
nor g0241 ( new_n456_, N171, N177 );
nand g0242 ( new_n457_, N171, N177 );
not g0243 ( new_n458_, new_n457_ );
nor g0244 ( new_n459_, new_n458_, new_n456_ );
not g0245 ( new_n460_, new_n459_ );
nand g0246 ( new_n461_, N159, N165 );
not g0247 ( new_n462_, new_n461_ );
nor g0248 ( new_n463_, new_n460_, new_n462_ );
nor g0249 ( new_n464_, new_n459_, new_n461_ );
nor g0250 ( new_n465_, new_n463_, new_n464_ );
nor g0251 ( new_n466_, N159, N165 );
nor g0252 ( new_n467_, new_n466_, keyIn_0_15 );
not g0253 ( new_n468_, new_n467_ );
nor g0254 ( new_n469_, new_n465_, new_n468_ );
nand g0255 ( new_n470_, new_n465_, new_n468_ );
not g0256 ( new_n471_, new_n470_ );
nor g0257 ( new_n472_, new_n471_, new_n469_ );
nor g0258 ( new_n473_, new_n472_, new_n321_ );
nand g0259 ( new_n474_, new_n472_, new_n321_ );
not g0260 ( new_n475_, new_n474_ );
nor g0261 ( new_n476_, new_n475_, new_n473_ );
not g0262 ( new_n477_, new_n476_ );
nor g0263 ( new_n478_, new_n477_, keyIn_0_61 );
not g0264 ( new_n479_, keyIn_0_61 );
nor g0265 ( new_n480_, new_n476_, new_n479_ );
nor g0266 ( new_n481_, new_n478_, new_n480_ );
nor g0267 ( new_n482_, new_n454_, new_n422_ );
nor g0268 ( new_n483_, new_n482_, new_n481_ );
nand g0269 ( new_n484_, new_n483_, new_n455_ );
nor g0270 ( new_n485_, new_n484_, new_n421_ );
not g0271 ( new_n486_, new_n454_ );
nand g0272 ( new_n487_, new_n486_, new_n476_ );
nand g0273 ( new_n488_, new_n484_, new_n421_ );
nand g0274 ( new_n489_, new_n488_, new_n487_ );
nor g0275 ( N768, new_n489_, new_n485_ );
not g0276 ( new_n491_, N261 );
not g0277 ( new_n492_, keyIn_0_82 );
not g0278 ( new_n493_, keyIn_0_56 );
not g0279 ( new_n494_, keyIn_0_50 );
not g0280 ( new_n495_, keyIn_0_36 );
not g0281 ( new_n496_, keyIn_0_2 );
nand g0282 ( new_n497_, N17, N51 );
nor g0283 ( new_n498_, new_n231_, new_n497_ );
nand g0284 ( new_n499_, new_n498_, new_n496_ );
not g0285 ( new_n500_, new_n497_ );
nand g0286 ( new_n501_, new_n232_, new_n500_ );
nand g0287 ( new_n502_, new_n501_, keyIn_0_2 );
nand g0288 ( new_n503_, new_n502_, new_n499_ );
not g0289 ( new_n504_, keyIn_0_7 );
nand g0290 ( new_n505_, new_n244_, N42 );
nand g0291 ( new_n506_, new_n505_, new_n504_ );
nor g0292 ( new_n507_, new_n243_, new_n222_ );
nand g0293 ( new_n508_, new_n507_, keyIn_0_7 );
nand g0294 ( new_n509_, new_n506_, new_n508_ );
nand g0295 ( new_n510_, new_n503_, new_n509_ );
nand g0296 ( new_n511_, N17, N42 );
not g0297 ( new_n512_, new_n511_ );
nand g0298 ( new_n513_, new_n230_, new_n222_ );
nand g0299 ( new_n514_, N59, N156 );
not g0300 ( new_n515_, new_n514_ );
nand g0301 ( new_n516_, new_n513_, new_n515_ );
nor g0302 ( new_n517_, new_n516_, new_n512_ );
nand g0303 ( new_n518_, N447, new_n517_ );
nand g0304 ( new_n519_, new_n510_, new_n518_ );
nand g0305 ( new_n520_, new_n519_, new_n495_ );
nor g0306 ( new_n521_, new_n519_, new_n495_ );
not g0307 ( new_n522_, new_n521_ );
nand g0308 ( new_n523_, new_n522_, new_n520_ );
nand g0309 ( new_n524_, new_n523_, N126 );
nand g0310 ( new_n525_, new_n524_, new_n494_ );
not g0311 ( new_n526_, N126 );
not g0312 ( new_n527_, new_n520_ );
nor g0313 ( new_n528_, new_n527_, new_n521_ );
nor g0314 ( new_n529_, new_n528_, new_n526_ );
nand g0315 ( new_n530_, new_n529_, keyIn_0_50 );
nand g0316 ( new_n531_, new_n530_, new_n525_ );
not g0317 ( new_n532_, keyIn_0_35 );
nor g0318 ( new_n533_, new_n278_, keyIn_0_1 );
nor g0319 ( new_n534_, new_n275_, new_n273_ );
nor g0320 ( new_n535_, new_n534_, new_n533_ );
not g0321 ( new_n536_, keyIn_0_14 );
nand g0322 ( new_n537_, new_n514_, new_n536_ );
not g0323 ( new_n538_, new_n537_ );
nor g0324 ( new_n539_, new_n514_, new_n536_ );
nor g0325 ( new_n540_, new_n538_, new_n539_ );
not g0326 ( new_n541_, new_n540_ );
nor g0327 ( new_n542_, new_n535_, new_n541_ );
nand g0328 ( new_n543_, new_n542_, N17 );
nand g0329 ( new_n544_, new_n543_, new_n532_ );
nand g0330 ( new_n545_, N447, new_n540_ );
nor g0331 ( new_n546_, new_n545_, new_n230_ );
nand g0332 ( new_n547_, new_n546_, keyIn_0_35 );
nand g0333 ( new_n548_, new_n544_, new_n547_ );
nand g0334 ( new_n549_, new_n548_, N1 );
nand g0335 ( new_n550_, new_n549_, N153 );
nand g0336 ( new_n551_, new_n531_, new_n550_ );
nor g0337 ( new_n552_, new_n551_, new_n493_ );
nand g0338 ( new_n553_, N29, N75 );
nor g0339 ( new_n554_, new_n553_, new_n218_ );
nand g0340 ( new_n555_, N447, new_n554_ );
nand g0341 ( new_n556_, keyIn_0_24, N268 );
not g0342 ( new_n557_, new_n556_ );
nor g0343 ( new_n558_, keyIn_0_24, N268 );
nor g0344 ( new_n559_, new_n557_, new_n558_ );
nor g0345 ( new_n560_, new_n559_, new_n283_ );
not g0346 ( new_n561_, new_n560_ );
nor g0347 ( new_n562_, new_n555_, new_n561_ );
not g0348 ( new_n563_, new_n562_ );
nand g0349 ( new_n564_, new_n551_, new_n493_ );
nand g0350 ( new_n565_, new_n564_, new_n563_ );
nor g0351 ( new_n566_, new_n565_, new_n552_ );
nor g0352 ( new_n567_, new_n566_, new_n436_ );
not g0353 ( new_n568_, new_n567_ );
nand g0354 ( new_n569_, new_n566_, new_n436_ );
nand g0355 ( new_n570_, new_n568_, new_n569_ );
not g0356 ( new_n571_, new_n570_ );
nor g0357 ( new_n572_, new_n571_, new_n492_ );
nor g0358 ( new_n573_, new_n570_, keyIn_0_82 );
nor g0359 ( new_n574_, new_n572_, new_n573_ );
nor g0360 ( new_n575_, new_n574_, new_n491_ );
nand g0361 ( new_n576_, new_n575_, keyIn_0_93 );
not g0362 ( new_n577_, keyIn_0_93 );
not g0363 ( new_n578_, new_n575_ );
nand g0364 ( new_n579_, new_n578_, new_n577_ );
not g0365 ( new_n580_, new_n579_ );
nand g0366 ( new_n581_, new_n574_, new_n491_ );
nand g0367 ( new_n582_, new_n581_, N219 );
nor g0368 ( new_n583_, new_n580_, new_n582_ );
nand g0369 ( new_n584_, new_n583_, new_n576_ );
not g0370 ( new_n585_, new_n574_ );
nand g0371 ( new_n586_, new_n585_, N228 );
not g0372 ( new_n587_, N237 );
nor g0373 ( new_n588_, new_n568_, new_n587_ );
not g0374 ( new_n589_, new_n566_ );
nand g0375 ( new_n590_, new_n589_, N246 );
not g0376 ( new_n591_, N73 );
nand g0377 ( new_n592_, N42, N72 );
nor g0378 ( new_n593_, new_n592_, new_n591_ );
nand g0379 ( new_n594_, new_n593_, new_n302_ );
nor g0380 ( new_n595_, new_n289_, new_n594_ );
nor g0381 ( new_n596_, new_n595_, keyIn_0_33 );
nand g0382 ( new_n597_, new_n595_, keyIn_0_33 );
not g0383 ( new_n598_, new_n597_ );
nor g0384 ( new_n599_, new_n598_, new_n596_ );
not g0385 ( new_n600_, new_n599_ );
nand g0386 ( new_n601_, new_n600_, N201 );
not g0387 ( new_n602_, keyIn_0_18 );
nand g0388 ( new_n603_, N255, N267 );
nor g0389 ( new_n604_, new_n603_, new_n602_ );
nand g0390 ( new_n605_, new_n603_, new_n602_ );
nand g0391 ( new_n606_, N121, N210 );
nand g0392 ( new_n607_, new_n605_, new_n606_ );
nor g0393 ( new_n608_, new_n607_, new_n604_ );
nand g0394 ( new_n609_, new_n601_, new_n608_ );
not g0395 ( new_n610_, new_n609_ );
nand g0396 ( new_n611_, new_n590_, new_n610_ );
nor g0397 ( new_n612_, new_n588_, new_n611_ );
nand g0398 ( new_n613_, new_n586_, new_n612_ );
not g0399 ( new_n614_, new_n613_ );
nand g0400 ( N850, new_n584_, new_n614_ );
not g0401 ( new_n616_, keyIn_0_120 );
not g0402 ( new_n617_, keyIn_0_106 );
not g0403 ( new_n618_, keyIn_0_103 );
not g0404 ( new_n619_, N183 );
nand g0405 ( new_n620_, new_n549_, N143 );
not g0406 ( new_n621_, new_n620_ );
nand g0407 ( new_n622_, new_n523_, N111 );
not g0408 ( new_n623_, keyIn_0_42 );
nor g0409 ( new_n624_, new_n562_, new_n623_ );
nor g0410 ( new_n625_, new_n563_, keyIn_0_42 );
nor g0411 ( new_n626_, new_n625_, new_n624_ );
nand g0412 ( new_n627_, new_n622_, new_n626_ );
nor g0413 ( new_n628_, new_n621_, new_n627_ );
nor g0414 ( new_n629_, new_n628_, new_n619_ );
not g0415 ( new_n630_, new_n628_ );
nor g0416 ( new_n631_, new_n630_, N183 );
nor g0417 ( new_n632_, new_n631_, new_n629_ );
not g0418 ( new_n633_, new_n632_ );
nand g0419 ( new_n634_, new_n633_, keyIn_0_79 );
not g0420 ( new_n635_, new_n634_ );
nor g0421 ( new_n636_, new_n633_, keyIn_0_79 );
nor g0422 ( new_n637_, new_n635_, new_n636_ );
not g0423 ( new_n638_, N189 );
nand g0424 ( new_n639_, new_n549_, N146 );
nand g0425 ( new_n640_, new_n639_, keyIn_0_48 );
nor g0426 ( new_n641_, new_n639_, keyIn_0_48 );
not g0427 ( new_n642_, new_n641_ );
nand g0428 ( new_n643_, new_n642_, new_n640_ );
nand g0429 ( new_n644_, new_n523_, N116 );
nand g0430 ( new_n645_, new_n644_, new_n563_ );
not g0431 ( new_n646_, new_n645_ );
nand g0432 ( new_n647_, new_n643_, new_n646_ );
nand g0433 ( new_n648_, new_n647_, keyIn_0_60 );
not g0434 ( new_n649_, keyIn_0_60 );
not g0435 ( new_n650_, new_n640_ );
nor g0436 ( new_n651_, new_n650_, new_n641_ );
nor g0437 ( new_n652_, new_n651_, new_n645_ );
nand g0438 ( new_n653_, new_n652_, new_n649_ );
nand g0439 ( new_n654_, new_n653_, new_n648_ );
nand g0440 ( new_n655_, new_n654_, new_n638_ );
nand g0441 ( new_n656_, new_n655_, keyIn_0_70 );
nor g0442 ( new_n657_, new_n655_, keyIn_0_70 );
not g0443 ( new_n658_, new_n657_ );
nand g0444 ( new_n659_, new_n658_, new_n656_ );
not g0445 ( new_n660_, keyIn_0_49 );
nand g0446 ( new_n661_, new_n549_, N149 );
nand g0447 ( new_n662_, new_n661_, new_n660_ );
not g0448 ( new_n663_, new_n661_ );
nand g0449 ( new_n664_, new_n663_, keyIn_0_49 );
nand g0450 ( new_n665_, new_n664_, new_n662_ );
nand g0451 ( new_n666_, new_n523_, N121 );
not g0452 ( new_n667_, new_n666_ );
nor g0453 ( new_n668_, new_n562_, keyIn_0_43 );
nand g0454 ( new_n669_, new_n562_, keyIn_0_43 );
not g0455 ( new_n670_, new_n669_ );
nor g0456 ( new_n671_, new_n670_, new_n668_ );
nor g0457 ( new_n672_, new_n667_, new_n671_ );
nand g0458 ( new_n673_, new_n665_, new_n672_ );
nor g0459 ( new_n674_, new_n673_, N195 );
nor g0460 ( new_n675_, new_n674_, keyIn_0_72 );
not g0461 ( new_n676_, new_n675_ );
nand g0462 ( new_n677_, new_n674_, keyIn_0_72 );
nand g0463 ( new_n678_, new_n676_, new_n677_ );
nand g0464 ( new_n679_, new_n678_, new_n567_ );
not g0465 ( new_n680_, new_n679_ );
nand g0466 ( new_n681_, new_n659_, new_n680_ );
nand g0467 ( new_n682_, new_n681_, keyIn_0_95 );
not g0468 ( new_n683_, keyIn_0_95 );
not g0469 ( new_n684_, new_n656_ );
nor g0470 ( new_n685_, new_n684_, new_n657_ );
nor g0471 ( new_n686_, new_n685_, new_n679_ );
nand g0472 ( new_n687_, new_n686_, new_n683_ );
nand g0473 ( new_n688_, new_n687_, new_n682_ );
not g0474 ( new_n689_, keyIn_0_71 );
nand g0475 ( new_n690_, new_n673_, N195 );
nand g0476 ( new_n691_, new_n690_, new_n689_ );
not g0477 ( new_n692_, new_n690_ );
nand g0478 ( new_n693_, new_n692_, keyIn_0_71 );
nand g0479 ( new_n694_, new_n693_, new_n691_ );
nand g0480 ( new_n695_, new_n694_, keyIn_0_80 );
not g0481 ( new_n696_, keyIn_0_80 );
not g0482 ( new_n697_, new_n691_ );
nor g0483 ( new_n698_, new_n690_, new_n689_ );
nor g0484 ( new_n699_, new_n697_, new_n698_ );
nand g0485 ( new_n700_, new_n699_, new_n696_ );
nand g0486 ( new_n701_, new_n700_, new_n695_ );
nand g0487 ( new_n702_, new_n569_, N261 );
not g0488 ( new_n703_, new_n702_ );
nand g0489 ( new_n704_, new_n703_, new_n678_ );
nand g0490 ( new_n705_, new_n701_, new_n704_ );
nand g0491 ( new_n706_, new_n705_, new_n659_ );
nor g0492 ( new_n707_, new_n654_, new_n638_ );
nand g0493 ( new_n708_, new_n707_, keyIn_0_90 );
not g0494 ( new_n709_, keyIn_0_90 );
not g0495 ( new_n710_, new_n707_ );
nand g0496 ( new_n711_, new_n710_, new_n709_ );
nand g0497 ( new_n712_, new_n711_, new_n708_ );
nand g0498 ( new_n713_, new_n706_, new_n712_ );
not g0499 ( new_n714_, new_n713_ );
nand g0500 ( new_n715_, new_n714_, new_n688_ );
nand g0501 ( new_n716_, new_n715_, new_n637_ );
not g0502 ( new_n717_, new_n716_ );
nor g0503 ( new_n718_, new_n715_, new_n637_ );
nor g0504 ( new_n719_, new_n717_, new_n718_ );
not g0505 ( new_n720_, new_n719_ );
nor g0506 ( new_n721_, new_n720_, new_n618_ );
nand g0507 ( new_n722_, new_n720_, new_n618_ );
nand g0508 ( new_n723_, new_n722_, N219 );
nor g0509 ( new_n724_, new_n723_, new_n721_ );
not g0510 ( new_n725_, new_n724_ );
nor g0511 ( new_n726_, new_n725_, new_n617_ );
nor g0512 ( new_n727_, new_n724_, keyIn_0_106 );
not g0513 ( new_n728_, N228 );
nor g0514 ( new_n729_, new_n637_, new_n728_ );
not g0515 ( new_n730_, new_n729_ );
nor g0516 ( new_n731_, new_n730_, keyIn_0_89 );
nand g0517 ( new_n732_, new_n730_, keyIn_0_89 );
nor g0518 ( new_n733_, new_n629_, keyIn_0_78 );
nand g0519 ( new_n734_, new_n629_, keyIn_0_78 );
not g0520 ( new_n735_, new_n734_ );
nor g0521 ( new_n736_, new_n735_, new_n733_ );
nand g0522 ( new_n737_, new_n736_, N237 );
nand g0523 ( new_n738_, new_n732_, new_n737_ );
nor g0524 ( new_n739_, new_n738_, new_n731_ );
not g0525 ( new_n740_, new_n739_ );
nor g0526 ( new_n741_, new_n740_, keyIn_0_98 );
nand g0527 ( new_n742_, new_n740_, keyIn_0_98 );
not g0528 ( new_n743_, N246 );
nor g0529 ( new_n744_, new_n628_, new_n743_ );
nand g0530 ( new_n745_, N106, N210 );
nand g0531 ( new_n746_, new_n600_, N183 );
nand g0532 ( new_n747_, new_n746_, new_n745_ );
nor g0533 ( new_n748_, new_n747_, new_n744_ );
nand g0534 ( new_n749_, new_n742_, new_n748_ );
nor g0535 ( new_n750_, new_n749_, new_n741_ );
not g0536 ( new_n751_, new_n750_ );
nor g0537 ( new_n752_, new_n727_, new_n751_ );
not g0538 ( new_n753_, new_n752_ );
nor g0539 ( new_n754_, new_n753_, new_n726_ );
not g0540 ( new_n755_, new_n754_ );
nand g0541 ( new_n756_, new_n755_, new_n616_ );
nand g0542 ( new_n757_, new_n754_, keyIn_0_120 );
nand g0543 ( N863, new_n756_, new_n757_ );
not g0544 ( new_n759_, keyIn_0_111 );
nor g0545 ( new_n760_, new_n685_, new_n707_ );
not g0546 ( new_n761_, new_n760_ );
not g0547 ( new_n762_, keyIn_0_99 );
not g0548 ( new_n763_, keyIn_0_83 );
not g0549 ( new_n764_, new_n704_ );
nor g0550 ( new_n765_, new_n764_, new_n763_ );
nor g0551 ( new_n766_, new_n704_, keyIn_0_83 );
nor g0552 ( new_n767_, new_n765_, new_n766_ );
nor g0553 ( new_n768_, new_n679_, keyIn_0_94 );
nand g0554 ( new_n769_, new_n679_, keyIn_0_94 );
not g0555 ( new_n770_, new_n769_ );
nor g0556 ( new_n771_, new_n770_, new_n768_ );
not g0557 ( new_n772_, keyIn_0_91 );
nor g0558 ( new_n773_, new_n701_, new_n772_ );
not g0559 ( new_n774_, new_n701_ );
nor g0560 ( new_n775_, new_n774_, keyIn_0_91 );
nor g0561 ( new_n776_, new_n775_, new_n773_ );
nor g0562 ( new_n777_, new_n776_, new_n771_ );
not g0563 ( new_n778_, new_n777_ );
nor g0564 ( new_n779_, new_n778_, new_n767_ );
not g0565 ( new_n780_, new_n779_ );
nand g0566 ( new_n781_, new_n780_, new_n762_ );
nand g0567 ( new_n782_, new_n779_, keyIn_0_99 );
nand g0568 ( new_n783_, new_n781_, new_n782_ );
nor g0569 ( new_n784_, new_n783_, new_n761_ );
nand g0570 ( new_n785_, new_n783_, new_n761_ );
nand g0571 ( new_n786_, new_n785_, N219 );
nor g0572 ( new_n787_, new_n786_, new_n784_ );
nand g0573 ( new_n788_, N111, N210 );
not g0574 ( new_n789_, new_n788_ );
nor g0575 ( new_n790_, new_n787_, new_n789_ );
nand g0576 ( new_n791_, new_n790_, new_n759_ );
nor g0577 ( new_n792_, new_n790_, new_n759_ );
nand g0578 ( new_n793_, new_n760_, N228 );
nor g0579 ( new_n794_, new_n710_, new_n587_ );
not g0580 ( new_n795_, new_n654_ );
nand g0581 ( new_n796_, new_n795_, N246 );
nand g0582 ( new_n797_, new_n600_, N189 );
nand g0583 ( new_n798_, N255, N259 );
nand g0584 ( new_n799_, new_n797_, new_n798_ );
not g0585 ( new_n800_, new_n799_ );
nand g0586 ( new_n801_, new_n796_, new_n800_ );
nor g0587 ( new_n802_, new_n794_, new_n801_ );
nand g0588 ( new_n803_, new_n793_, new_n802_ );
nor g0589 ( new_n804_, new_n792_, new_n803_ );
nand g0590 ( N864, new_n804_, new_n791_ );
not g0591 ( new_n806_, keyIn_0_117 );
not g0592 ( new_n807_, new_n678_ );
nor g0593 ( new_n808_, new_n807_, new_n694_ );
not g0594 ( new_n809_, new_n808_ );
nand g0595 ( new_n810_, new_n702_, new_n568_ );
nand g0596 ( new_n811_, new_n809_, new_n810_ );
not g0597 ( new_n812_, new_n811_ );
nor g0598 ( new_n813_, new_n809_, new_n810_ );
nor g0599 ( new_n814_, new_n812_, new_n813_ );
not g0600 ( new_n815_, new_n814_ );
nor g0601 ( new_n816_, new_n815_, keyIn_0_104 );
nand g0602 ( new_n817_, new_n815_, keyIn_0_104 );
nand g0603 ( new_n818_, new_n817_, N219 );
nor g0604 ( new_n819_, new_n818_, new_n816_ );
not g0605 ( new_n820_, keyIn_0_100 );
nor g0606 ( new_n821_, new_n809_, new_n728_ );
not g0607 ( new_n822_, new_n821_ );
nor g0608 ( new_n823_, new_n822_, keyIn_0_92 );
nor g0609 ( new_n824_, new_n701_, new_n587_ );
nand g0610 ( new_n825_, new_n822_, keyIn_0_92 );
not g0611 ( new_n826_, new_n825_ );
nor g0612 ( new_n827_, new_n826_, new_n824_ );
not g0613 ( new_n828_, new_n827_ );
nor g0614 ( new_n829_, new_n828_, new_n823_ );
not g0615 ( new_n830_, new_n829_ );
nand g0616 ( new_n831_, new_n830_, new_n820_ );
nand g0617 ( new_n832_, new_n829_, keyIn_0_100 );
nand g0618 ( new_n833_, new_n831_, new_n832_ );
nand g0619 ( new_n834_, new_n673_, N246 );
nand g0620 ( new_n835_, N255, N260 );
nand g0621 ( new_n836_, new_n834_, new_n835_ );
nand g0622 ( new_n837_, new_n836_, keyIn_0_81 );
not g0623 ( new_n838_, new_n837_ );
nor g0624 ( new_n839_, new_n836_, keyIn_0_81 );
nor g0625 ( new_n840_, new_n838_, new_n839_ );
nand g0626 ( new_n841_, new_n600_, N195 );
not g0627 ( new_n842_, keyIn_0_17 );
nand g0628 ( new_n843_, N116, N210 );
nand g0629 ( new_n844_, new_n843_, new_n842_ );
not g0630 ( new_n845_, new_n844_ );
nor g0631 ( new_n846_, new_n843_, new_n842_ );
nor g0632 ( new_n847_, new_n845_, new_n846_ );
nand g0633 ( new_n848_, new_n841_, new_n847_ );
nor g0634 ( new_n849_, new_n840_, new_n848_ );
nand g0635 ( new_n850_, new_n833_, new_n849_ );
nor g0636 ( new_n851_, new_n850_, new_n819_ );
not g0637 ( new_n852_, new_n851_ );
nand g0638 ( new_n853_, new_n852_, new_n806_ );
nand g0639 ( new_n854_, new_n851_, keyIn_0_117 );
nand g0640 ( N865, new_n853_, new_n854_ );
not g0641 ( new_n856_, keyIn_0_114 );
not g0642 ( new_n857_, keyIn_0_66 );
nor g0643 ( new_n858_, new_n545_, new_n283_ );
nor g0644 ( new_n859_, new_n858_, keyIn_0_34 );
nand g0645 ( new_n860_, new_n858_, keyIn_0_34 );
not g0646 ( new_n861_, new_n860_ );
nor g0647 ( new_n862_, new_n861_, new_n859_ );
not g0648 ( new_n863_, new_n862_ );
nand g0649 ( new_n864_, new_n863_, N146 );
nor g0650 ( new_n865_, new_n864_, keyIn_0_39 );
nand g0651 ( new_n866_, new_n864_, keyIn_0_39 );
nor g0652 ( new_n867_, new_n528_, new_n342_ );
nor g0653 ( new_n868_, new_n230_, N268 );
not g0654 ( new_n869_, new_n868_ );
nor g0655 ( new_n870_, new_n555_, new_n869_ );
nor g0656 ( new_n871_, new_n870_, keyIn_0_40 );
nand g0657 ( new_n872_, new_n870_, keyIn_0_40 );
nand g0658 ( new_n873_, N51, N138 );
nand g0659 ( new_n874_, new_n872_, new_n873_ );
nor g0660 ( new_n875_, new_n874_, new_n871_ );
not g0661 ( new_n876_, new_n875_ );
nor g0662 ( new_n877_, new_n867_, new_n876_ );
nand g0663 ( new_n878_, new_n866_, new_n877_ );
nor g0664 ( new_n879_, new_n878_, new_n865_ );
not g0665 ( new_n880_, new_n879_ );
nor g0666 ( new_n881_, new_n880_, N165 );
not g0667 ( new_n882_, new_n881_ );
nor g0668 ( new_n883_, new_n882_, new_n857_ );
nor g0669 ( new_n884_, new_n881_, keyIn_0_66 );
nor g0670 ( new_n885_, new_n883_, new_n884_ );
not g0671 ( new_n886_, keyIn_0_68 );
not g0672 ( new_n887_, keyIn_0_55 );
nand g0673 ( new_n888_, new_n523_, N101 );
nand g0674 ( new_n889_, N17, N138 );
nand g0675 ( new_n890_, new_n888_, new_n889_ );
nand g0676 ( new_n891_, new_n890_, new_n887_ );
not g0677 ( new_n892_, new_n891_ );
nor g0678 ( new_n893_, new_n890_, new_n887_ );
nor g0679 ( new_n894_, new_n892_, new_n893_ );
nand g0680 ( new_n895_, new_n863_, N149 );
nor g0681 ( new_n896_, new_n895_, keyIn_0_41 );
not g0682 ( new_n897_, new_n870_ );
nand g0683 ( new_n898_, new_n895_, keyIn_0_41 );
nand g0684 ( new_n899_, new_n898_, new_n897_ );
nor g0685 ( new_n900_, new_n899_, new_n896_ );
not g0686 ( new_n901_, new_n900_ );
nor g0687 ( new_n902_, new_n901_, new_n894_ );
not g0688 ( new_n903_, new_n902_ );
nor g0689 ( new_n904_, new_n903_, N171 );
nor g0690 ( new_n905_, new_n904_, new_n886_ );
nand g0691 ( new_n906_, new_n904_, new_n886_ );
not g0692 ( new_n907_, new_n906_ );
nor g0693 ( new_n908_, new_n907_, new_n905_ );
not g0694 ( new_n909_, new_n908_ );
not g0695 ( new_n910_, keyIn_0_69 );
not g0696 ( new_n911_, keyIn_0_59 );
nand g0697 ( new_n912_, new_n863_, N153 );
nand g0698 ( new_n913_, new_n912_, new_n897_ );
nor g0699 ( new_n914_, new_n913_, keyIn_0_47 );
nand g0700 ( new_n915_, new_n913_, keyIn_0_47 );
not g0701 ( new_n916_, N106 );
nor g0702 ( new_n917_, new_n528_, new_n916_ );
nand g0703 ( new_n918_, N138, N152 );
nand g0704 ( new_n919_, new_n918_, keyIn_0_13 );
not g0705 ( new_n920_, keyIn_0_13 );
not g0706 ( new_n921_, new_n918_ );
nand g0707 ( new_n922_, new_n921_, new_n920_ );
nand g0708 ( new_n923_, new_n922_, new_n919_ );
nor g0709 ( new_n924_, new_n917_, new_n923_ );
nand g0710 ( new_n925_, new_n915_, new_n924_ );
nor g0711 ( new_n926_, new_n925_, new_n914_ );
not g0712 ( new_n927_, new_n926_ );
nor g0713 ( new_n928_, new_n927_, new_n911_ );
nor g0714 ( new_n929_, new_n926_, keyIn_0_59 );
nor g0715 ( new_n930_, new_n928_, new_n929_ );
nor g0716 ( new_n931_, new_n930_, N177 );
not g0717 ( new_n932_, new_n931_ );
nand g0718 ( new_n933_, new_n932_, new_n910_ );
not g0719 ( new_n934_, new_n933_ );
nor g0720 ( new_n935_, new_n932_, new_n910_ );
nor g0721 ( new_n936_, new_n934_, new_n935_ );
not g0722 ( new_n937_, keyIn_0_102 );
not g0723 ( new_n938_, new_n736_ );
not g0724 ( new_n939_, keyIn_0_101 );
not g0725 ( new_n940_, new_n631_ );
nand g0726 ( new_n941_, new_n715_, new_n940_ );
nand g0727 ( new_n942_, new_n941_, new_n939_ );
nor g0728 ( new_n943_, new_n941_, new_n939_ );
not g0729 ( new_n944_, new_n943_ );
nand g0730 ( new_n945_, new_n944_, new_n942_ );
nand g0731 ( new_n946_, new_n945_, new_n938_ );
nand g0732 ( new_n947_, new_n946_, new_n937_ );
not g0733 ( new_n948_, new_n942_ );
nor g0734 ( new_n949_, new_n948_, new_n943_ );
nor g0735 ( new_n950_, new_n949_, new_n736_ );
nand g0736 ( new_n951_, new_n950_, keyIn_0_102 );
nand g0737 ( new_n952_, new_n951_, new_n947_ );
nor g0738 ( new_n953_, new_n952_, new_n936_ );
nand g0739 ( new_n954_, new_n953_, new_n909_ );
nor g0740 ( new_n955_, new_n954_, new_n885_ );
not g0741 ( new_n956_, new_n885_ );
not g0742 ( new_n957_, N177 );
not g0743 ( new_n958_, new_n930_ );
nor g0744 ( new_n959_, new_n958_, new_n957_ );
not g0745 ( new_n960_, new_n959_ );
nor g0746 ( new_n961_, new_n908_, new_n960_ );
not g0747 ( new_n962_, new_n961_ );
not g0748 ( new_n963_, keyIn_0_67 );
nand g0749 ( new_n964_, new_n903_, N171 );
nand g0750 ( new_n965_, new_n964_, new_n963_ );
not g0751 ( new_n966_, new_n965_ );
nor g0752 ( new_n967_, new_n964_, new_n963_ );
nor g0753 ( new_n968_, new_n966_, new_n967_ );
nand g0754 ( new_n969_, new_n962_, new_n968_ );
nand g0755 ( new_n970_, new_n969_, new_n956_ );
not g0756 ( new_n971_, N165 );
nor g0757 ( new_n972_, new_n879_, new_n971_ );
not g0758 ( new_n973_, new_n972_ );
nand g0759 ( new_n974_, new_n970_, new_n973_ );
nor g0760 ( new_n975_, new_n955_, new_n974_ );
not g0761 ( new_n976_, keyIn_0_58 );
not g0762 ( new_n977_, keyIn_0_54 );
nor g0763 ( new_n978_, new_n528_, new_n340_ );
nand g0764 ( new_n979_, N8, N138 );
not g0765 ( new_n980_, new_n979_ );
nor g0766 ( new_n981_, new_n978_, new_n980_ );
not g0767 ( new_n982_, new_n981_ );
nand g0768 ( new_n983_, new_n982_, new_n977_ );
not g0769 ( new_n984_, new_n983_ );
nor g0770 ( new_n985_, new_n982_, new_n977_ );
nor g0771 ( new_n986_, new_n984_, new_n985_ );
not g0772 ( new_n987_, keyIn_0_37 );
nand g0773 ( new_n988_, new_n863_, N143 );
nor g0774 ( new_n989_, new_n988_, new_n987_ );
not g0775 ( new_n990_, keyIn_0_38 );
nand g0776 ( new_n991_, new_n870_, new_n990_ );
nand g0777 ( new_n992_, new_n897_, keyIn_0_38 );
nand g0778 ( new_n993_, new_n992_, new_n991_ );
nand g0779 ( new_n994_, new_n988_, new_n987_ );
nand g0780 ( new_n995_, new_n994_, new_n993_ );
nor g0781 ( new_n996_, new_n995_, new_n989_ );
not g0782 ( new_n997_, new_n996_ );
nor g0783 ( new_n998_, new_n986_, new_n997_ );
nor g0784 ( new_n999_, new_n998_, new_n976_ );
nand g0785 ( new_n1000_, new_n998_, new_n976_ );
not g0786 ( new_n1001_, new_n1000_ );
nor g0787 ( new_n1002_, new_n1001_, new_n999_ );
nor g0788 ( new_n1003_, new_n1002_, N159 );
not g0789 ( new_n1004_, new_n1003_ );
nand g0790 ( new_n1005_, new_n1004_, keyIn_0_65 );
not g0791 ( new_n1006_, new_n1005_ );
nor g0792 ( new_n1007_, new_n1004_, keyIn_0_65 );
nor g0793 ( new_n1008_, new_n1006_, new_n1007_ );
nor g0794 ( new_n1009_, new_n975_, new_n1008_ );
not g0795 ( new_n1010_, new_n1009_ );
nor g0796 ( new_n1011_, new_n1010_, new_n856_ );
nor g0797 ( new_n1012_, new_n1009_, keyIn_0_114 );
not g0798 ( new_n1013_, N159 );
not g0799 ( new_n1014_, new_n1002_ );
nor g0800 ( new_n1015_, new_n1014_, new_n1013_ );
nor g0801 ( new_n1016_, new_n1015_, keyIn_0_73 );
nand g0802 ( new_n1017_, new_n1015_, keyIn_0_73 );
not g0803 ( new_n1018_, new_n1017_ );
nor g0804 ( new_n1019_, new_n1018_, new_n1016_ );
not g0805 ( new_n1020_, new_n1019_ );
nor g0806 ( new_n1021_, new_n1012_, new_n1020_ );
not g0807 ( new_n1022_, new_n1021_ );
nor g0808 ( new_n1023_, new_n1022_, new_n1011_ );
not g0809 ( new_n1024_, new_n1023_ );
nand g0810 ( new_n1025_, new_n1024_, keyIn_0_118 );
not g0811 ( new_n1026_, keyIn_0_118 );
nand g0812 ( new_n1027_, new_n1023_, new_n1026_ );
nand g0813 ( N866, new_n1025_, new_n1027_ );
not g0814 ( new_n1029_, keyIn_0_110 );
not g0815 ( new_n1030_, keyIn_0_105 );
not g0816 ( new_n1031_, new_n952_ );
nor g0817 ( new_n1032_, new_n936_, new_n959_ );
nor g0818 ( new_n1033_, new_n1031_, new_n1032_ );
not g0819 ( new_n1034_, new_n1033_ );
nor g0820 ( new_n1035_, new_n1034_, new_n1030_ );
nand g0821 ( new_n1036_, new_n1031_, new_n1032_ );
nand g0822 ( new_n1037_, new_n1034_, new_n1030_ );
nand g0823 ( new_n1038_, new_n1037_, new_n1036_ );
nor g0824 ( new_n1039_, new_n1038_, new_n1035_ );
not g0825 ( new_n1040_, new_n1039_ );
nor g0826 ( new_n1041_, new_n1040_, new_n1029_ );
not g0827 ( new_n1042_, N219 );
nor g0828 ( new_n1043_, new_n1039_, keyIn_0_110 );
nor g0829 ( new_n1044_, new_n1043_, new_n1042_ );
not g0830 ( new_n1045_, new_n1044_ );
nor g0831 ( new_n1046_, new_n1045_, new_n1041_ );
nand g0832 ( new_n1047_, new_n1032_, N228 );
nor g0833 ( new_n1048_, new_n960_, new_n587_ );
nor g0834 ( new_n1049_, new_n958_, new_n743_ );
nor g0835 ( new_n1050_, new_n599_, new_n957_ );
not g0836 ( new_n1051_, new_n1050_ );
nand g0837 ( new_n1052_, new_n1051_, keyIn_0_52 );
not g0838 ( new_n1053_, new_n1052_ );
nor g0839 ( new_n1054_, new_n1051_, keyIn_0_52 );
nor g0840 ( new_n1055_, new_n1053_, new_n1054_ );
nand g0841 ( new_n1056_, N101, N210 );
not g0842 ( new_n1057_, new_n1056_ );
nor g0843 ( new_n1058_, new_n1055_, new_n1057_ );
not g0844 ( new_n1059_, new_n1058_ );
nor g0845 ( new_n1060_, new_n1049_, new_n1059_ );
not g0846 ( new_n1061_, new_n1060_ );
nor g0847 ( new_n1062_, new_n1048_, new_n1061_ );
nand g0848 ( new_n1063_, new_n1047_, new_n1062_ );
nor g0849 ( new_n1064_, new_n1046_, new_n1063_ );
not g0850 ( new_n1065_, new_n1064_ );
nand g0851 ( new_n1066_, new_n1065_, keyIn_0_123 );
not g0852 ( new_n1067_, keyIn_0_123 );
nand g0853 ( new_n1068_, new_n1064_, new_n1067_ );
nand g0854 ( N874, new_n1066_, new_n1068_ );
not g0855 ( new_n1070_, keyIn_0_124 );
nor g0856 ( new_n1071_, new_n1008_, new_n1015_ );
nor g0857 ( new_n1072_, new_n1071_, keyIn_0_74 );
nand g0858 ( new_n1073_, new_n1071_, keyIn_0_74 );
not g0859 ( new_n1074_, new_n1073_ );
nor g0860 ( new_n1075_, new_n1074_, new_n1072_ );
not g0861 ( new_n1076_, new_n1075_ );
nand g0862 ( new_n1077_, new_n975_, new_n1076_ );
nor g0863 ( new_n1078_, new_n1077_, keyIn_0_112 );
nand g0864 ( new_n1079_, new_n1077_, keyIn_0_112 );
not g0865 ( new_n1080_, new_n975_ );
nand g0866 ( new_n1081_, new_n1080_, new_n1075_ );
nand g0867 ( new_n1082_, new_n1079_, new_n1081_ );
nor g0868 ( new_n1083_, new_n1082_, new_n1078_ );
nor g0869 ( new_n1084_, new_n1083_, keyIn_0_115 );
not g0870 ( new_n1085_, new_n1084_ );
nand g0871 ( new_n1086_, new_n1083_, keyIn_0_115 );
nand g0872 ( new_n1087_, new_n1086_, N219 );
not g0873 ( new_n1088_, new_n1087_ );
nand g0874 ( new_n1089_, new_n1088_, new_n1085_ );
nand g0875 ( new_n1090_, new_n559_, N210 );
not g0876 ( new_n1091_, new_n1090_ );
nor g0877 ( new_n1092_, new_n1091_, keyIn_0_32 );
nand g0878 ( new_n1093_, new_n1091_, keyIn_0_32 );
not g0879 ( new_n1094_, new_n1093_ );
nor g0880 ( new_n1095_, new_n1094_, new_n1092_ );
not g0881 ( new_n1096_, new_n1095_ );
nand g0882 ( new_n1097_, new_n1089_, new_n1096_ );
nand g0883 ( new_n1098_, new_n1097_, keyIn_0_121 );
not g0884 ( new_n1099_, keyIn_0_121 );
nor g0885 ( new_n1100_, new_n1087_, new_n1084_ );
nor g0886 ( new_n1101_, new_n1100_, new_n1095_ );
nand g0887 ( new_n1102_, new_n1101_, new_n1099_ );
nand g0888 ( new_n1103_, new_n1098_, new_n1102_ );
nor g0889 ( new_n1104_, new_n1076_, new_n728_ );
nor g0890 ( new_n1105_, new_n1019_, new_n587_ );
not g0891 ( new_n1106_, new_n1105_ );
nor g0892 ( new_n1107_, new_n1106_, keyIn_0_84 );
nand g0893 ( new_n1108_, new_n1106_, keyIn_0_84 );
nor g0894 ( new_n1109_, new_n1014_, new_n743_ );
nor g0895 ( new_n1110_, new_n599_, new_n1013_ );
nor g0896 ( new_n1111_, new_n1109_, new_n1110_ );
nand g0897 ( new_n1112_, new_n1108_, new_n1111_ );
nor g0898 ( new_n1113_, new_n1112_, new_n1107_ );
not g0899 ( new_n1114_, new_n1113_ );
nor g0900 ( new_n1115_, new_n1104_, new_n1114_ );
nand g0901 ( new_n1116_, new_n1103_, new_n1115_ );
nand g0902 ( new_n1117_, new_n1116_, new_n1070_ );
not g0903 ( new_n1118_, new_n1116_ );
nand g0904 ( new_n1119_, new_n1118_, keyIn_0_124 );
nand g0905 ( new_n1120_, new_n1119_, new_n1117_ );
nand g0906 ( new_n1121_, new_n1120_, keyIn_0_125 );
not g0907 ( new_n1122_, keyIn_0_125 );
not g0908 ( new_n1123_, new_n1117_ );
nor g0909 ( new_n1124_, new_n1116_, new_n1070_ );
nor g0910 ( new_n1125_, new_n1123_, new_n1124_ );
nand g0911 ( new_n1126_, new_n1125_, new_n1122_ );
nand g0912 ( N878, new_n1126_, new_n1121_ );
not g0913 ( new_n1128_, keyIn_0_126 );
nand g0914 ( new_n1129_, new_n956_, new_n973_ );
not g0915 ( new_n1130_, keyIn_0_108 );
not g0916 ( new_n1131_, keyIn_0_107 );
not g0917 ( new_n1132_, new_n954_ );
nor g0918 ( new_n1133_, new_n1132_, new_n1131_ );
nor g0919 ( new_n1134_, new_n954_, keyIn_0_107 );
not g0920 ( new_n1135_, keyIn_0_96 );
nor g0921 ( new_n1136_, new_n962_, new_n1135_ );
nand g0922 ( new_n1137_, new_n962_, new_n1135_ );
nor g0923 ( new_n1138_, new_n968_, keyIn_0_86 );
nand g0924 ( new_n1139_, new_n968_, keyIn_0_86 );
not g0925 ( new_n1140_, new_n1139_ );
nor g0926 ( new_n1141_, new_n1140_, new_n1138_ );
nand g0927 ( new_n1142_, new_n1137_, new_n1141_ );
nor g0928 ( new_n1143_, new_n1142_, new_n1136_ );
not g0929 ( new_n1144_, new_n1143_ );
nor g0930 ( new_n1145_, new_n1134_, new_n1144_ );
not g0931 ( new_n1146_, new_n1145_ );
nor g0932 ( new_n1147_, new_n1146_, new_n1133_ );
nor g0933 ( new_n1148_, new_n1147_, new_n1130_ );
nand g0934 ( new_n1149_, new_n1147_, new_n1130_ );
not g0935 ( new_n1150_, new_n1149_ );
nor g0936 ( new_n1151_, new_n1150_, new_n1148_ );
nor g0937 ( new_n1152_, new_n1151_, new_n1129_ );
nand g0938 ( new_n1153_, new_n1151_, new_n1129_ );
nand g0939 ( new_n1154_, new_n1153_, N219 );
nor g0940 ( new_n1155_, new_n1154_, new_n1152_ );
not g0941 ( new_n1156_, new_n1155_ );
nor g0942 ( new_n1157_, new_n1156_, keyIn_0_119 );
not g0943 ( new_n1158_, keyIn_0_119 );
nor g0944 ( new_n1159_, new_n1155_, new_n1158_ );
nor g0945 ( new_n1160_, new_n1129_, new_n728_ );
nor g0946 ( new_n1161_, new_n1160_, keyIn_0_85 );
nand g0947 ( new_n1162_, new_n1160_, keyIn_0_85 );
not g0948 ( new_n1163_, new_n1162_ );
nor g0949 ( new_n1164_, new_n1163_, new_n1161_ );
nor g0950 ( new_n1165_, new_n879_, new_n743_ );
nor g0951 ( new_n1166_, new_n599_, new_n971_ );
nor g0952 ( new_n1167_, new_n1165_, new_n1166_ );
not g0953 ( new_n1168_, new_n1167_ );
nand g0954 ( new_n1169_, new_n1168_, keyIn_0_75 );
not g0955 ( new_n1170_, new_n1169_ );
nor g0956 ( new_n1171_, new_n1168_, keyIn_0_75 );
nor g0957 ( new_n1172_, new_n1170_, new_n1171_ );
nor g0958 ( new_n1173_, new_n973_, new_n587_ );
nand g0959 ( new_n1174_, N91, N210 );
nand g0960 ( new_n1175_, new_n1174_, keyIn_0_16 );
not g0961 ( new_n1176_, new_n1175_ );
nor g0962 ( new_n1177_, new_n1174_, keyIn_0_16 );
nor g0963 ( new_n1178_, new_n1176_, new_n1177_ );
not g0964 ( new_n1179_, new_n1178_ );
nor g0965 ( new_n1180_, new_n1173_, new_n1179_ );
not g0966 ( new_n1181_, new_n1180_ );
nor g0967 ( new_n1182_, new_n1172_, new_n1181_ );
not g0968 ( new_n1183_, new_n1182_ );
nor g0969 ( new_n1184_, new_n1164_, new_n1183_ );
not g0970 ( new_n1185_, new_n1184_ );
nor g0971 ( new_n1186_, new_n1159_, new_n1185_ );
not g0972 ( new_n1187_, new_n1186_ );
nor g0973 ( new_n1188_, new_n1187_, new_n1157_ );
not g0974 ( new_n1189_, new_n1188_ );
nand g0975 ( new_n1190_, new_n1189_, new_n1128_ );
nand g0976 ( new_n1191_, new_n1188_, keyIn_0_126 );
nand g0977 ( N879, new_n1190_, new_n1191_ );
not g0978 ( new_n1193_, keyIn_0_127 );
not g0979 ( new_n1194_, keyIn_0_122 );
not g0980 ( new_n1195_, keyIn_0_116 );
not g0981 ( new_n1196_, keyIn_0_113 );
not g0982 ( new_n1197_, new_n968_ );
nor g0983 ( new_n1198_, new_n1197_, new_n908_ );
nor g0984 ( new_n1199_, new_n1198_, keyIn_0_76 );
nand g0985 ( new_n1200_, new_n1198_, keyIn_0_76 );
not g0986 ( new_n1201_, new_n1200_ );
nor g0987 ( new_n1202_, new_n1201_, new_n1199_ );
not g0988 ( new_n1203_, new_n1202_ );
not g0989 ( new_n1204_, keyIn_0_109 );
nor g0990 ( new_n1205_, new_n960_, keyIn_0_88 );
nand g0991 ( new_n1206_, new_n960_, keyIn_0_88 );
not g0992 ( new_n1207_, new_n1206_ );
nor g0993 ( new_n1208_, new_n1207_, new_n1205_ );
nor g0994 ( new_n1209_, new_n953_, new_n1208_ );
not g0995 ( new_n1210_, new_n1209_ );
nand g0996 ( new_n1211_, new_n1210_, new_n1204_ );
nand g0997 ( new_n1212_, new_n1209_, keyIn_0_109 );
nand g0998 ( new_n1213_, new_n1211_, new_n1212_ );
nand g0999 ( new_n1214_, new_n1213_, new_n1203_ );
nand g1000 ( new_n1215_, new_n1214_, new_n1196_ );
not g1001 ( new_n1216_, new_n1214_ );
nand g1002 ( new_n1217_, new_n1216_, keyIn_0_113 );
nand g1003 ( new_n1218_, new_n1217_, new_n1215_ );
nor g1004 ( new_n1219_, new_n1213_, new_n1203_ );
not g1005 ( new_n1220_, new_n1219_ );
nand g1006 ( new_n1221_, new_n1218_, new_n1220_ );
nor g1007 ( new_n1222_, new_n1221_, new_n1195_ );
nand g1008 ( new_n1223_, new_n1221_, new_n1195_ );
nand g1009 ( new_n1224_, new_n1223_, N219 );
nor g1010 ( new_n1225_, new_n1224_, new_n1222_ );
nand g1011 ( new_n1226_, N96, N210 );
not g1012 ( new_n1227_, new_n1226_ );
nor g1013 ( new_n1228_, new_n1225_, new_n1227_ );
not g1014 ( new_n1229_, new_n1228_ );
nor g1015 ( new_n1230_, new_n1229_, new_n1194_ );
not g1016 ( new_n1231_, new_n1230_ );
nor g1017 ( new_n1232_, new_n1228_, keyIn_0_122 );
not g1018 ( new_n1233_, keyIn_0_97 );
not g1019 ( new_n1234_, keyIn_0_87 );
nor g1020 ( new_n1235_, new_n1203_, new_n728_ );
nor g1021 ( new_n1236_, new_n1235_, new_n1234_ );
nand g1022 ( new_n1237_, new_n1235_, new_n1234_ );
not g1023 ( new_n1238_, new_n1237_ );
nor g1024 ( new_n1239_, new_n1238_, new_n1236_ );
nor g1025 ( new_n1240_, new_n968_, new_n587_ );
nor g1026 ( new_n1241_, new_n1239_, new_n1240_ );
not g1027 ( new_n1242_, new_n1241_ );
nand g1028 ( new_n1243_, new_n1242_, new_n1233_ );
not g1029 ( new_n1244_, new_n1243_ );
nor g1030 ( new_n1245_, new_n1242_, new_n1233_ );
nor g1031 ( new_n1246_, new_n1244_, new_n1245_ );
nand g1032 ( new_n1247_, new_n903_, N246 );
nand g1033 ( new_n1248_, new_n600_, N171 );
nand g1034 ( new_n1249_, new_n1247_, new_n1248_ );
nand g1035 ( new_n1250_, new_n1249_, keyIn_0_77 );
not g1036 ( new_n1251_, new_n1250_ );
nor g1037 ( new_n1252_, new_n1249_, keyIn_0_77 );
nor g1038 ( new_n1253_, new_n1251_, new_n1252_ );
nor g1039 ( new_n1254_, new_n1246_, new_n1253_ );
not g1040 ( new_n1255_, new_n1254_ );
nor g1041 ( new_n1256_, new_n1232_, new_n1255_ );
nand g1042 ( new_n1257_, new_n1231_, new_n1256_ );
nand g1043 ( new_n1258_, new_n1257_, new_n1193_ );
not g1044 ( new_n1259_, new_n1257_ );
nand g1045 ( new_n1260_, new_n1259_, keyIn_0_127 );
nand g1046 ( N880, new_n1260_, new_n1258_ );
endmodule