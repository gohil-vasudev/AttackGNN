module add_mul_comp_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, 
        a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, 
        a_17_, a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, 
        a_27_, a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, 
        b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, 
        b_16_, b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, 
        b_26_, b_27_, b_28_, b_29_, b_30_, b_31_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, 
        Result_32_, Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, 
        Result_38_, Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, 
        Result_44_, Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, 
        Result_50_, Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, 
        Result_56_, Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, 
        Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   Result_9_, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127;
  assign Result_8_ = Result_9_;
  assign Result_6_ = Result_9_;
  assign Result_4_ = Result_9_;
  assign Result_31_ = Result_9_;
  assign Result_2_ = Result_9_;
  assign Result_28_ = Result_9_;
  assign Result_26_ = Result_9_;
  assign Result_24_ = Result_9_;
  assign Result_22_ = Result_9_;
  assign Result_20_ = Result_9_;
  assign Result_19_ = Result_9_;
  assign Result_17_ = Result_9_;
  assign Result_15_ = Result_9_;
  assign Result_13_ = Result_9_;
  assign Result_11_ = Result_9_;
  assign Result_0_ = Result_9_;
  assign Result_10_ = Result_9_;
  assign Result_12_ = Result_9_;
  assign Result_14_ = Result_9_;
  assign Result_16_ = Result_9_;
  assign Result_18_ = Result_9_;
  assign Result_1_ = Result_9_;
  assign Result_21_ = Result_9_;
  assign Result_23_ = Result_9_;
  assign Result_25_ = Result_9_;
  assign Result_27_ = Result_9_;
  assign Result_29_ = Result_9_;
  assign Result_30_ = Result_9_;
  assign Result_3_ = Result_9_;
  assign Result_5_ = Result_9_;
  assign Result_7_ = Result_9_;

  NAND2_X2 U601 ( .A1(n988), .A2(n989), .ZN(Result_9_) );
  INV_X2 U602 ( .A(n578), .ZN(n589) );
  XOR2_X1 U603 ( .A(b_31_), .B(a_31_), .Z(Result_63_) );
  NAND2_X1 U604 ( .A1(n568), .A2(n569), .ZN(Result_62_) );
  NAND2_X1 U605 ( .A1(n570), .A2(n571), .ZN(n569) );
  AND2_X1 U606 ( .A1(n572), .A2(n573), .ZN(n571) );
  NOR2_X1 U607 ( .A1(n574), .A2(n575), .ZN(n570) );
  NAND2_X1 U608 ( .A1(n576), .A2(n577), .ZN(n575) );
  NAND2_X1 U609 ( .A1(b_31_), .A2(n578), .ZN(n577) );
  NAND2_X1 U610 ( .A1(n579), .A2(n580), .ZN(n576) );
  NAND2_X1 U611 ( .A1(n581), .A2(n582), .ZN(n568) );
  XOR2_X1 U612 ( .A(b_30_), .B(a_30_), .Z(n582) );
  NOR2_X1 U613 ( .A1(n583), .A2(n584), .ZN(n581) );
  NOR2_X1 U614 ( .A1(Result_9_), .A2(n585), .ZN(n584) );
  NOR2_X1 U615 ( .A1(n574), .A2(n586), .ZN(n583) );
  NAND2_X1 U616 ( .A1(n578), .A2(n580), .ZN(n586) );
  NAND2_X1 U617 ( .A1(n587), .A2(n588), .ZN(Result_61_) );
  NAND2_X1 U618 ( .A1(n589), .A2(n590), .ZN(n588) );
  XOR2_X1 U619 ( .A(n591), .B(n592), .Z(n590) );
  NAND2_X1 U620 ( .A1(n593), .A2(Result_9_), .ZN(n587) );
  XNOR2_X1 U621 ( .A(n594), .B(n591), .ZN(n593) );
  NAND2_X1 U622 ( .A1(n595), .A2(n596), .ZN(n591) );
  NAND2_X1 U623 ( .A1(n597), .A2(n598), .ZN(Result_60_) );
  NAND2_X1 U624 ( .A1(n589), .A2(n599), .ZN(n598) );
  XNOR2_X1 U625 ( .A(n600), .B(n601), .ZN(n599) );
  NAND2_X1 U626 ( .A1(n602), .A2(Result_9_), .ZN(n597) );
  XOR2_X1 U627 ( .A(n603), .B(n600), .Z(n602) );
  AND2_X1 U628 ( .A1(n604), .A2(n605), .ZN(n600) );
  NAND2_X1 U629 ( .A1(n606), .A2(n607), .ZN(Result_59_) );
  NAND2_X1 U630 ( .A1(n589), .A2(n608), .ZN(n607) );
  XOR2_X1 U631 ( .A(n609), .B(n610), .Z(n608) );
  NAND2_X1 U632 ( .A1(n611), .A2(Result_9_), .ZN(n606) );
  XNOR2_X1 U633 ( .A(n612), .B(n609), .ZN(n611) );
  NAND2_X1 U634 ( .A1(n613), .A2(n614), .ZN(n609) );
  NAND2_X1 U635 ( .A1(n615), .A2(n616), .ZN(Result_58_) );
  NAND2_X1 U636 ( .A1(n589), .A2(n617), .ZN(n616) );
  XNOR2_X1 U637 ( .A(n618), .B(n619), .ZN(n617) );
  NAND2_X1 U638 ( .A1(n620), .A2(Result_9_), .ZN(n615) );
  XOR2_X1 U639 ( .A(n621), .B(n618), .Z(n620) );
  AND2_X1 U640 ( .A1(n622), .A2(n623), .ZN(n618) );
  NAND2_X1 U641 ( .A1(n624), .A2(n625), .ZN(Result_57_) );
  NAND2_X1 U642 ( .A1(n589), .A2(n626), .ZN(n625) );
  XOR2_X1 U643 ( .A(n627), .B(n628), .Z(n626) );
  NAND2_X1 U644 ( .A1(n629), .A2(Result_9_), .ZN(n624) );
  XNOR2_X1 U645 ( .A(n630), .B(n627), .ZN(n629) );
  NAND2_X1 U646 ( .A1(n631), .A2(n632), .ZN(n627) );
  NAND2_X1 U647 ( .A1(n633), .A2(n634), .ZN(Result_56_) );
  NAND2_X1 U648 ( .A1(n589), .A2(n635), .ZN(n634) );
  XNOR2_X1 U649 ( .A(n636), .B(n637), .ZN(n635) );
  NAND2_X1 U650 ( .A1(n638), .A2(Result_9_), .ZN(n633) );
  XOR2_X1 U651 ( .A(n639), .B(n636), .Z(n638) );
  AND2_X1 U652 ( .A1(n640), .A2(n641), .ZN(n636) );
  NAND2_X1 U653 ( .A1(n642), .A2(n643), .ZN(Result_55_) );
  NAND2_X1 U654 ( .A1(n589), .A2(n644), .ZN(n643) );
  XOR2_X1 U655 ( .A(n645), .B(n646), .Z(n644) );
  NAND2_X1 U656 ( .A1(n647), .A2(Result_9_), .ZN(n642) );
  XNOR2_X1 U657 ( .A(n648), .B(n645), .ZN(n647) );
  NAND2_X1 U658 ( .A1(n649), .A2(n650), .ZN(n645) );
  NAND2_X1 U659 ( .A1(n651), .A2(n652), .ZN(Result_54_) );
  NAND2_X1 U660 ( .A1(n589), .A2(n653), .ZN(n652) );
  XNOR2_X1 U661 ( .A(n654), .B(n655), .ZN(n653) );
  NAND2_X1 U662 ( .A1(n656), .A2(Result_9_), .ZN(n651) );
  XOR2_X1 U663 ( .A(n657), .B(n654), .Z(n656) );
  AND2_X1 U664 ( .A1(n658), .A2(n659), .ZN(n654) );
  NAND2_X1 U665 ( .A1(n660), .A2(n661), .ZN(Result_53_) );
  NAND2_X1 U666 ( .A1(n589), .A2(n662), .ZN(n661) );
  XOR2_X1 U667 ( .A(n663), .B(n664), .Z(n662) );
  NAND2_X1 U668 ( .A1(n665), .A2(Result_9_), .ZN(n660) );
  XNOR2_X1 U669 ( .A(n666), .B(n663), .ZN(n665) );
  NAND2_X1 U670 ( .A1(n667), .A2(n668), .ZN(n663) );
  NAND2_X1 U671 ( .A1(n669), .A2(n670), .ZN(Result_52_) );
  NAND2_X1 U672 ( .A1(n589), .A2(n671), .ZN(n670) );
  XNOR2_X1 U673 ( .A(n672), .B(n673), .ZN(n671) );
  NAND2_X1 U674 ( .A1(n674), .A2(Result_9_), .ZN(n669) );
  XOR2_X1 U675 ( .A(n675), .B(n672), .Z(n674) );
  AND2_X1 U676 ( .A1(n676), .A2(n677), .ZN(n672) );
  NAND2_X1 U677 ( .A1(n678), .A2(n679), .ZN(Result_51_) );
  NAND2_X1 U678 ( .A1(n589), .A2(n680), .ZN(n679) );
  XOR2_X1 U679 ( .A(n681), .B(n682), .Z(n680) );
  NAND2_X1 U680 ( .A1(n683), .A2(Result_9_), .ZN(n678) );
  XNOR2_X1 U681 ( .A(n684), .B(n681), .ZN(n683) );
  NAND2_X1 U682 ( .A1(n685), .A2(n686), .ZN(n681) );
  NAND2_X1 U683 ( .A1(n687), .A2(n688), .ZN(Result_50_) );
  NAND2_X1 U684 ( .A1(n589), .A2(n689), .ZN(n688) );
  XNOR2_X1 U685 ( .A(n690), .B(n691), .ZN(n689) );
  NAND2_X1 U686 ( .A1(n692), .A2(Result_9_), .ZN(n687) );
  XOR2_X1 U687 ( .A(n693), .B(n690), .Z(n692) );
  AND2_X1 U688 ( .A1(n694), .A2(n695), .ZN(n690) );
  NAND2_X1 U689 ( .A1(n696), .A2(n697), .ZN(Result_49_) );
  NAND2_X1 U690 ( .A1(n589), .A2(n698), .ZN(n697) );
  XOR2_X1 U691 ( .A(n699), .B(n700), .Z(n698) );
  NAND2_X1 U692 ( .A1(n701), .A2(Result_9_), .ZN(n696) );
  XNOR2_X1 U693 ( .A(n702), .B(n699), .ZN(n701) );
  NAND2_X1 U694 ( .A1(n703), .A2(n704), .ZN(n699) );
  NAND2_X1 U695 ( .A1(n705), .A2(n706), .ZN(Result_48_) );
  NAND2_X1 U696 ( .A1(n589), .A2(n707), .ZN(n706) );
  XNOR2_X1 U697 ( .A(n708), .B(n709), .ZN(n707) );
  NAND2_X1 U698 ( .A1(n710), .A2(Result_9_), .ZN(n705) );
  XOR2_X1 U699 ( .A(n711), .B(n708), .Z(n710) );
  AND2_X1 U700 ( .A1(n712), .A2(n713), .ZN(n708) );
  NAND2_X1 U701 ( .A1(n714), .A2(n715), .ZN(Result_47_) );
  NAND2_X1 U702 ( .A1(n589), .A2(n716), .ZN(n715) );
  XOR2_X1 U703 ( .A(n717), .B(n718), .Z(n716) );
  NAND2_X1 U704 ( .A1(n719), .A2(Result_9_), .ZN(n714) );
  XNOR2_X1 U705 ( .A(n720), .B(n717), .ZN(n719) );
  NAND2_X1 U706 ( .A1(n721), .A2(n722), .ZN(n717) );
  NAND2_X1 U707 ( .A1(n723), .A2(n724), .ZN(Result_46_) );
  NAND2_X1 U708 ( .A1(n589), .A2(n725), .ZN(n724) );
  XNOR2_X1 U709 ( .A(n726), .B(n727), .ZN(n725) );
  NAND2_X1 U710 ( .A1(n728), .A2(Result_9_), .ZN(n723) );
  XOR2_X1 U711 ( .A(n729), .B(n726), .Z(n728) );
  AND2_X1 U712 ( .A1(n730), .A2(n731), .ZN(n726) );
  NAND2_X1 U713 ( .A1(n732), .A2(n733), .ZN(Result_45_) );
  NAND2_X1 U714 ( .A1(n589), .A2(n734), .ZN(n733) );
  XOR2_X1 U715 ( .A(n735), .B(n736), .Z(n734) );
  NAND2_X1 U716 ( .A1(n737), .A2(Result_9_), .ZN(n732) );
  XNOR2_X1 U717 ( .A(n738), .B(n735), .ZN(n737) );
  NAND2_X1 U718 ( .A1(n739), .A2(n740), .ZN(n735) );
  NAND2_X1 U719 ( .A1(n741), .A2(n742), .ZN(Result_44_) );
  NAND2_X1 U720 ( .A1(n589), .A2(n743), .ZN(n742) );
  XNOR2_X1 U721 ( .A(n744), .B(n745), .ZN(n743) );
  NAND2_X1 U722 ( .A1(n746), .A2(Result_9_), .ZN(n741) );
  XOR2_X1 U723 ( .A(n747), .B(n744), .Z(n746) );
  AND2_X1 U724 ( .A1(n748), .A2(n749), .ZN(n744) );
  NAND2_X1 U725 ( .A1(n750), .A2(n751), .ZN(Result_43_) );
  NAND2_X1 U726 ( .A1(n589), .A2(n752), .ZN(n751) );
  XOR2_X1 U727 ( .A(n753), .B(n754), .Z(n752) );
  NAND2_X1 U728 ( .A1(n755), .A2(Result_9_), .ZN(n750) );
  XNOR2_X1 U729 ( .A(n756), .B(n753), .ZN(n755) );
  NAND2_X1 U730 ( .A1(n757), .A2(n758), .ZN(n753) );
  NAND2_X1 U731 ( .A1(n759), .A2(n760), .ZN(Result_42_) );
  NAND2_X1 U732 ( .A1(n589), .A2(n761), .ZN(n760) );
  XNOR2_X1 U733 ( .A(n762), .B(n763), .ZN(n761) );
  NAND2_X1 U734 ( .A1(n764), .A2(Result_9_), .ZN(n759) );
  XOR2_X1 U735 ( .A(n765), .B(n762), .Z(n764) );
  AND2_X1 U736 ( .A1(n766), .A2(n767), .ZN(n762) );
  NAND2_X1 U737 ( .A1(n768), .A2(n769), .ZN(Result_41_) );
  NAND2_X1 U738 ( .A1(n589), .A2(n770), .ZN(n769) );
  XOR2_X1 U739 ( .A(n771), .B(n772), .Z(n770) );
  NAND2_X1 U740 ( .A1(n773), .A2(Result_9_), .ZN(n768) );
  XNOR2_X1 U741 ( .A(n774), .B(n771), .ZN(n773) );
  NAND2_X1 U742 ( .A1(n775), .A2(n776), .ZN(n771) );
  NAND2_X1 U743 ( .A1(n777), .A2(n778), .ZN(Result_40_) );
  NAND2_X1 U744 ( .A1(n589), .A2(n779), .ZN(n778) );
  XNOR2_X1 U745 ( .A(n780), .B(n781), .ZN(n779) );
  NAND2_X1 U746 ( .A1(n782), .A2(Result_9_), .ZN(n777) );
  XOR2_X1 U747 ( .A(n783), .B(n780), .Z(n782) );
  AND2_X1 U748 ( .A1(n784), .A2(n785), .ZN(n780) );
  NAND2_X1 U749 ( .A1(n786), .A2(n787), .ZN(Result_39_) );
  NAND2_X1 U750 ( .A1(n589), .A2(n788), .ZN(n787) );
  XOR2_X1 U751 ( .A(n789), .B(n790), .Z(n788) );
  NAND2_X1 U752 ( .A1(n791), .A2(Result_9_), .ZN(n786) );
  XNOR2_X1 U753 ( .A(n792), .B(n789), .ZN(n791) );
  NAND2_X1 U754 ( .A1(n793), .A2(n794), .ZN(n789) );
  NAND2_X1 U755 ( .A1(n795), .A2(n796), .ZN(Result_38_) );
  NAND2_X1 U756 ( .A1(n589), .A2(n797), .ZN(n796) );
  XNOR2_X1 U757 ( .A(n798), .B(n799), .ZN(n797) );
  NAND2_X1 U758 ( .A1(n800), .A2(Result_9_), .ZN(n795) );
  XOR2_X1 U759 ( .A(n801), .B(n798), .Z(n800) );
  AND2_X1 U760 ( .A1(n802), .A2(n803), .ZN(n798) );
  NAND2_X1 U761 ( .A1(n804), .A2(n805), .ZN(Result_37_) );
  NAND2_X1 U762 ( .A1(n589), .A2(n806), .ZN(n805) );
  XOR2_X1 U763 ( .A(n807), .B(n808), .Z(n806) );
  NAND2_X1 U764 ( .A1(n809), .A2(Result_9_), .ZN(n804) );
  XNOR2_X1 U765 ( .A(n810), .B(n807), .ZN(n809) );
  NAND2_X1 U766 ( .A1(n811), .A2(n812), .ZN(n807) );
  NAND2_X1 U767 ( .A1(n813), .A2(n814), .ZN(Result_36_) );
  NAND2_X1 U768 ( .A1(n589), .A2(n815), .ZN(n814) );
  XNOR2_X1 U769 ( .A(n816), .B(n817), .ZN(n815) );
  NAND2_X1 U770 ( .A1(n818), .A2(Result_9_), .ZN(n813) );
  XOR2_X1 U771 ( .A(n819), .B(n816), .Z(n818) );
  AND2_X1 U772 ( .A1(n820), .A2(n821), .ZN(n816) );
  NAND2_X1 U773 ( .A1(n822), .A2(n823), .ZN(Result_35_) );
  NAND2_X1 U774 ( .A1(n589), .A2(n824), .ZN(n823) );
  XOR2_X1 U775 ( .A(n825), .B(n826), .Z(n824) );
  NAND2_X1 U776 ( .A1(n827), .A2(Result_9_), .ZN(n822) );
  XNOR2_X1 U777 ( .A(n828), .B(n825), .ZN(n827) );
  NAND2_X1 U778 ( .A1(n829), .A2(n830), .ZN(n825) );
  NAND2_X1 U779 ( .A1(n831), .A2(n832), .ZN(Result_34_) );
  NAND2_X1 U780 ( .A1(n589), .A2(n833), .ZN(n832) );
  XNOR2_X1 U781 ( .A(n834), .B(n835), .ZN(n833) );
  NAND2_X1 U782 ( .A1(n836), .A2(Result_9_), .ZN(n831) );
  XOR2_X1 U783 ( .A(n837), .B(n834), .Z(n836) );
  AND2_X1 U784 ( .A1(n838), .A2(n839), .ZN(n834) );
  NAND2_X1 U785 ( .A1(n840), .A2(n841), .ZN(Result_33_) );
  NAND2_X1 U786 ( .A1(n589), .A2(n842), .ZN(n841) );
  XOR2_X1 U787 ( .A(n843), .B(n844), .Z(n842) );
  NAND2_X1 U788 ( .A1(n845), .A2(Result_9_), .ZN(n840) );
  XNOR2_X1 U789 ( .A(n846), .B(n843), .ZN(n845) );
  NAND2_X1 U790 ( .A1(n847), .A2(n848), .ZN(n843) );
  NAND2_X1 U791 ( .A1(n849), .A2(n850), .ZN(Result_32_) );
  NAND2_X1 U792 ( .A1(n589), .A2(n851), .ZN(n850) );
  XOR2_X1 U793 ( .A(n852), .B(n853), .Z(n851) );
  NOR2_X1 U794 ( .A1(n854), .A2(n855), .ZN(n853) );
  AND2_X1 U795 ( .A1(n844), .A2(a_1_), .ZN(n855) );
  NOR2_X1 U796 ( .A1(n856), .A2(n857), .ZN(n854) );
  NOR2_X1 U797 ( .A1(a_1_), .A2(n844), .ZN(n856) );
  NAND2_X1 U798 ( .A1(n858), .A2(n859), .ZN(n844) );
  NAND2_X1 U799 ( .A1(b_2_), .A2(n860), .ZN(n859) );
  OR2_X1 U800 ( .A1(n835), .A2(a_2_), .ZN(n860) );
  NAND2_X1 U801 ( .A1(a_2_), .A2(n835), .ZN(n858) );
  NAND2_X1 U802 ( .A1(n861), .A2(n862), .ZN(n835) );
  NAND2_X1 U803 ( .A1(b_3_), .A2(n863), .ZN(n862) );
  OR2_X1 U804 ( .A1(n826), .A2(a_3_), .ZN(n863) );
  NAND2_X1 U805 ( .A1(a_3_), .A2(n826), .ZN(n861) );
  NAND2_X1 U806 ( .A1(n864), .A2(n865), .ZN(n826) );
  NAND2_X1 U807 ( .A1(b_4_), .A2(n866), .ZN(n865) );
  OR2_X1 U808 ( .A1(n817), .A2(a_4_), .ZN(n866) );
  NAND2_X1 U809 ( .A1(a_4_), .A2(n817), .ZN(n864) );
  NAND2_X1 U810 ( .A1(n867), .A2(n868), .ZN(n817) );
  NAND2_X1 U811 ( .A1(b_5_), .A2(n869), .ZN(n868) );
  OR2_X1 U812 ( .A1(n808), .A2(a_5_), .ZN(n869) );
  NAND2_X1 U813 ( .A1(a_5_), .A2(n808), .ZN(n867) );
  NAND2_X1 U814 ( .A1(n870), .A2(n871), .ZN(n808) );
  NAND2_X1 U815 ( .A1(b_6_), .A2(n872), .ZN(n871) );
  OR2_X1 U816 ( .A1(n799), .A2(a_6_), .ZN(n872) );
  NAND2_X1 U817 ( .A1(a_6_), .A2(n799), .ZN(n870) );
  NAND2_X1 U818 ( .A1(n873), .A2(n874), .ZN(n799) );
  NAND2_X1 U819 ( .A1(b_7_), .A2(n875), .ZN(n874) );
  OR2_X1 U820 ( .A1(n790), .A2(a_7_), .ZN(n875) );
  NAND2_X1 U821 ( .A1(a_7_), .A2(n790), .ZN(n873) );
  NAND2_X1 U822 ( .A1(n876), .A2(n877), .ZN(n790) );
  NAND2_X1 U823 ( .A1(b_8_), .A2(n878), .ZN(n877) );
  OR2_X1 U824 ( .A1(n781), .A2(a_8_), .ZN(n878) );
  NAND2_X1 U825 ( .A1(a_8_), .A2(n781), .ZN(n876) );
  NAND2_X1 U826 ( .A1(n879), .A2(n880), .ZN(n781) );
  NAND2_X1 U827 ( .A1(b_9_), .A2(n881), .ZN(n880) );
  OR2_X1 U828 ( .A1(n772), .A2(a_9_), .ZN(n881) );
  NAND2_X1 U829 ( .A1(a_9_), .A2(n772), .ZN(n879) );
  NAND2_X1 U830 ( .A1(n882), .A2(n883), .ZN(n772) );
  NAND2_X1 U831 ( .A1(b_10_), .A2(n884), .ZN(n883) );
  OR2_X1 U832 ( .A1(n763), .A2(a_10_), .ZN(n884) );
  NAND2_X1 U833 ( .A1(a_10_), .A2(n763), .ZN(n882) );
  NAND2_X1 U834 ( .A1(n885), .A2(n886), .ZN(n763) );
  NAND2_X1 U835 ( .A1(b_11_), .A2(n887), .ZN(n886) );
  OR2_X1 U836 ( .A1(n754), .A2(a_11_), .ZN(n887) );
  NAND2_X1 U837 ( .A1(a_11_), .A2(n754), .ZN(n885) );
  NAND2_X1 U838 ( .A1(n888), .A2(n889), .ZN(n754) );
  NAND2_X1 U839 ( .A1(b_12_), .A2(n890), .ZN(n889) );
  OR2_X1 U840 ( .A1(n745), .A2(a_12_), .ZN(n890) );
  NAND2_X1 U841 ( .A1(a_12_), .A2(n745), .ZN(n888) );
  NAND2_X1 U842 ( .A1(n891), .A2(n892), .ZN(n745) );
  NAND2_X1 U843 ( .A1(b_13_), .A2(n893), .ZN(n892) );
  OR2_X1 U844 ( .A1(n736), .A2(a_13_), .ZN(n893) );
  NAND2_X1 U845 ( .A1(a_13_), .A2(n736), .ZN(n891) );
  NAND2_X1 U846 ( .A1(n894), .A2(n895), .ZN(n736) );
  NAND2_X1 U847 ( .A1(b_14_), .A2(n896), .ZN(n895) );
  OR2_X1 U848 ( .A1(n727), .A2(a_14_), .ZN(n896) );
  NAND2_X1 U849 ( .A1(a_14_), .A2(n727), .ZN(n894) );
  NAND2_X1 U850 ( .A1(n897), .A2(n898), .ZN(n727) );
  NAND2_X1 U851 ( .A1(b_15_), .A2(n899), .ZN(n898) );
  OR2_X1 U852 ( .A1(n718), .A2(a_15_), .ZN(n899) );
  NAND2_X1 U853 ( .A1(a_15_), .A2(n718), .ZN(n897) );
  NAND2_X1 U854 ( .A1(n900), .A2(n901), .ZN(n718) );
  NAND2_X1 U855 ( .A1(b_16_), .A2(n902), .ZN(n901) );
  OR2_X1 U856 ( .A1(n709), .A2(a_16_), .ZN(n902) );
  NAND2_X1 U857 ( .A1(a_16_), .A2(n709), .ZN(n900) );
  NAND2_X1 U858 ( .A1(n903), .A2(n904), .ZN(n709) );
  NAND2_X1 U859 ( .A1(b_17_), .A2(n905), .ZN(n904) );
  OR2_X1 U860 ( .A1(n700), .A2(a_17_), .ZN(n905) );
  NAND2_X1 U861 ( .A1(a_17_), .A2(n700), .ZN(n903) );
  NAND2_X1 U862 ( .A1(n906), .A2(n907), .ZN(n700) );
  NAND2_X1 U863 ( .A1(b_18_), .A2(n908), .ZN(n907) );
  OR2_X1 U864 ( .A1(n691), .A2(a_18_), .ZN(n908) );
  NAND2_X1 U865 ( .A1(a_18_), .A2(n691), .ZN(n906) );
  NAND2_X1 U866 ( .A1(n909), .A2(n910), .ZN(n691) );
  NAND2_X1 U867 ( .A1(b_19_), .A2(n911), .ZN(n910) );
  OR2_X1 U868 ( .A1(n682), .A2(a_19_), .ZN(n911) );
  NAND2_X1 U869 ( .A1(a_19_), .A2(n682), .ZN(n909) );
  NAND2_X1 U870 ( .A1(n912), .A2(n913), .ZN(n682) );
  NAND2_X1 U871 ( .A1(b_20_), .A2(n914), .ZN(n913) );
  OR2_X1 U872 ( .A1(n673), .A2(a_20_), .ZN(n914) );
  NAND2_X1 U873 ( .A1(a_20_), .A2(n673), .ZN(n912) );
  NAND2_X1 U874 ( .A1(n915), .A2(n916), .ZN(n673) );
  NAND2_X1 U875 ( .A1(b_21_), .A2(n917), .ZN(n916) );
  OR2_X1 U876 ( .A1(n664), .A2(a_21_), .ZN(n917) );
  NAND2_X1 U877 ( .A1(a_21_), .A2(n664), .ZN(n915) );
  NAND2_X1 U878 ( .A1(n918), .A2(n919), .ZN(n664) );
  NAND2_X1 U879 ( .A1(b_22_), .A2(n920), .ZN(n919) );
  OR2_X1 U880 ( .A1(n655), .A2(a_22_), .ZN(n920) );
  NAND2_X1 U881 ( .A1(a_22_), .A2(n655), .ZN(n918) );
  NAND2_X1 U882 ( .A1(n921), .A2(n922), .ZN(n655) );
  NAND2_X1 U883 ( .A1(b_23_), .A2(n923), .ZN(n922) );
  OR2_X1 U884 ( .A1(n646), .A2(a_23_), .ZN(n923) );
  NAND2_X1 U885 ( .A1(a_23_), .A2(n646), .ZN(n921) );
  NAND2_X1 U886 ( .A1(n924), .A2(n925), .ZN(n646) );
  NAND2_X1 U887 ( .A1(b_24_), .A2(n926), .ZN(n925) );
  OR2_X1 U888 ( .A1(n637), .A2(a_24_), .ZN(n926) );
  NAND2_X1 U889 ( .A1(a_24_), .A2(n637), .ZN(n924) );
  NAND2_X1 U890 ( .A1(n927), .A2(n928), .ZN(n637) );
  NAND2_X1 U891 ( .A1(b_25_), .A2(n929), .ZN(n928) );
  OR2_X1 U892 ( .A1(n628), .A2(a_25_), .ZN(n929) );
  NAND2_X1 U893 ( .A1(a_25_), .A2(n628), .ZN(n927) );
  NAND2_X1 U894 ( .A1(n930), .A2(n931), .ZN(n628) );
  NAND2_X1 U895 ( .A1(b_26_), .A2(n932), .ZN(n931) );
  OR2_X1 U896 ( .A1(n619), .A2(a_26_), .ZN(n932) );
  NAND2_X1 U897 ( .A1(a_26_), .A2(n619), .ZN(n930) );
  NAND2_X1 U898 ( .A1(n933), .A2(n934), .ZN(n619) );
  NAND2_X1 U899 ( .A1(b_27_), .A2(n935), .ZN(n934) );
  OR2_X1 U900 ( .A1(n610), .A2(a_27_), .ZN(n935) );
  NAND2_X1 U901 ( .A1(a_27_), .A2(n610), .ZN(n933) );
  NAND2_X1 U902 ( .A1(n936), .A2(n937), .ZN(n610) );
  NAND2_X1 U903 ( .A1(b_28_), .A2(n938), .ZN(n937) );
  OR2_X1 U904 ( .A1(n601), .A2(a_28_), .ZN(n938) );
  NAND2_X1 U905 ( .A1(a_28_), .A2(n601), .ZN(n936) );
  NAND2_X1 U906 ( .A1(n939), .A2(n940), .ZN(n601) );
  NAND2_X1 U907 ( .A1(b_29_), .A2(n941), .ZN(n940) );
  OR2_X1 U908 ( .A1(n592), .A2(a_29_), .ZN(n941) );
  NAND2_X1 U909 ( .A1(a_29_), .A2(n592), .ZN(n939) );
  NAND2_X1 U910 ( .A1(n942), .A2(n943), .ZN(n592) );
  NAND2_X1 U911 ( .A1(b_30_), .A2(n944), .ZN(n943) );
  NAND2_X1 U912 ( .A1(n945), .A2(n585), .ZN(n944) );
  OR2_X1 U913 ( .A1(n585), .A2(n945), .ZN(n942) );
  NAND2_X1 U914 ( .A1(b_31_), .A2(a_31_), .ZN(n585) );
  NAND2_X1 U915 ( .A1(n946), .A2(n579), .ZN(n578) );
  INV_X1 U916 ( .A(Result_9_), .ZN(n579) );
  NAND2_X1 U917 ( .A1(n947), .A2(n948), .ZN(n946) );
  NOR2_X1 U918 ( .A1(n949), .A2(n950), .ZN(n948) );
  NAND2_X1 U919 ( .A1(n951), .A2(n952), .ZN(n950) );
  NOR2_X1 U920 ( .A1(n953), .A2(n954), .ZN(n952) );
  NAND2_X1 U921 ( .A1(n712), .A2(n757), .ZN(n954) );
  NOR2_X1 U922 ( .A1(n955), .A2(n956), .ZN(n951) );
  NAND2_X1 U923 ( .A1(n640), .A2(n649), .ZN(n956) );
  NAND2_X1 U924 ( .A1(n957), .A2(n958), .ZN(n949) );
  NOR2_X1 U925 ( .A1(n959), .A2(n960), .ZN(n958) );
  NAND2_X1 U926 ( .A1(n572), .A2(n838), .ZN(n960) );
  NOR2_X1 U927 ( .A1(n961), .A2(n962), .ZN(n957) );
  NAND2_X1 U928 ( .A1(n848), .A2(n963), .ZN(n962) );
  NOR2_X1 U929 ( .A1(n964), .A2(n965), .ZN(n947) );
  NAND2_X1 U930 ( .A1(n966), .A2(n967), .ZN(n965) );
  NOR2_X1 U931 ( .A1(n968), .A2(n969), .ZN(n967) );
  NAND2_X1 U932 ( .A1(n970), .A2(n971), .ZN(n969) );
  INV_X1 U933 ( .A(n972), .ZN(n971) );
  NOR2_X1 U934 ( .A1(n973), .A2(n974), .ZN(n966) );
  NAND2_X1 U935 ( .A1(n975), .A2(n976), .ZN(n974) );
  INV_X1 U936 ( .A(n977), .ZN(n975) );
  NAND2_X1 U937 ( .A1(n978), .A2(n979), .ZN(n964) );
  NOR2_X1 U938 ( .A1(n980), .A2(n981), .ZN(n979) );
  NAND2_X1 U939 ( .A1(n748), .A2(n721), .ZN(n981) );
  NOR2_X1 U940 ( .A1(n982), .A2(n983), .ZN(n978) );
  NAND2_X1 U941 ( .A1(n984), .A2(n985), .ZN(n983) );
  NAND2_X1 U942 ( .A1(b_31_), .A2(n574), .ZN(n985) );
  INV_X1 U943 ( .A(a_31_), .ZN(n574) );
  INV_X1 U944 ( .A(n986), .ZN(n984) );
  NAND2_X1 U945 ( .A1(n987), .A2(Result_9_), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n990), .A2(n963), .ZN(n989) );
  NAND2_X1 U947 ( .A1(n847), .A2(n991), .ZN(n990) );
  NAND2_X1 U948 ( .A1(n992), .A2(n848), .ZN(n991) );
  INV_X1 U949 ( .A(n993), .ZN(n848) );
  NAND2_X1 U950 ( .A1(n839), .A2(n994), .ZN(n992) );
  NAND2_X1 U951 ( .A1(n995), .A2(n838), .ZN(n994) );
  NAND2_X1 U952 ( .A1(n830), .A2(n996), .ZN(n995) );
  NAND2_X1 U953 ( .A1(n997), .A2(n998), .ZN(n996) );
  NAND2_X1 U954 ( .A1(n999), .A2(n812), .ZN(n998) );
  NOR2_X1 U955 ( .A1(n1000), .A2(n1001), .ZN(n999) );
  NOR2_X1 U956 ( .A1(b_4_), .A2(n1002), .ZN(n1001) );
  NOR2_X1 U957 ( .A1(n1003), .A2(n977), .ZN(n1000) );
  NAND2_X1 U958 ( .A1(n802), .A2(n811), .ZN(n977) );
  NOR2_X1 U959 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
  NAND2_X1 U960 ( .A1(n803), .A2(n1006), .ZN(n1005) );
  NAND2_X1 U961 ( .A1(n976), .A2(n1007), .ZN(n1006) );
  NAND2_X1 U962 ( .A1(n1008), .A2(n776), .ZN(n1007) );
  NOR2_X1 U963 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
  NOR2_X1 U964 ( .A1(b_8_), .A2(n1011), .ZN(n1010) );
  NOR2_X1 U965 ( .A1(n980), .A2(n1012), .ZN(n1009) );
  NAND2_X1 U966 ( .A1(n1013), .A2(n775), .ZN(n1012) );
  NAND2_X1 U967 ( .A1(n1014), .A2(n758), .ZN(n1013) );
  NOR2_X1 U968 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
  AND2_X1 U969 ( .A1(n1017), .A2(a_10_), .ZN(n1016) );
  NOR2_X1 U970 ( .A1(n1018), .A2(n1019), .ZN(n1015) );
  NAND2_X1 U971 ( .A1(n1020), .A2(n757), .ZN(n1019) );
  NAND2_X1 U972 ( .A1(n1021), .A2(n740), .ZN(n1020) );
  NOR2_X1 U973 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
  AND2_X1 U974 ( .A1(n1024), .A2(a_12_), .ZN(n1023) );
  NOR2_X1 U975 ( .A1(n1025), .A2(n968), .ZN(n1022) );
  NAND2_X1 U976 ( .A1(n730), .A2(n739), .ZN(n968) );
  NOR2_X1 U977 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
  NAND2_X1 U978 ( .A1(n731), .A2(n1028), .ZN(n1027) );
  NAND2_X1 U979 ( .A1(n1029), .A2(n721), .ZN(n1028) );
  NOR2_X1 U980 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
  NOR2_X1 U981 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
  NAND2_X1 U982 ( .A1(n713), .A2(n1034), .ZN(n1033) );
  NAND2_X1 U983 ( .A1(n970), .A2(n1035), .ZN(n1034) );
  NAND2_X1 U984 ( .A1(n1036), .A2(n686), .ZN(n1035) );
  NOR2_X1 U985 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
  NOR2_X1 U986 ( .A1(b_18_), .A2(n1039), .ZN(n1038) );
  NOR2_X1 U987 ( .A1(n1040), .A2(n972), .ZN(n1037) );
  NAND2_X1 U988 ( .A1(n676), .A2(n685), .ZN(n972) );
  NOR2_X1 U989 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
  NAND2_X1 U990 ( .A1(n677), .A2(n1043), .ZN(n1042) );
  NAND2_X1 U991 ( .A1(n1044), .A2(n658), .ZN(n1043) );
  NOR2_X1 U992 ( .A1(n953), .A2(n1045), .ZN(n1044) );
  NOR2_X1 U993 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
  NAND2_X1 U994 ( .A1(n659), .A2(n1048), .ZN(n1047) );
  NAND2_X1 U995 ( .A1(n1049), .A2(n640), .ZN(n1048) );
  NOR2_X1 U996 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
  NOR2_X1 U997 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
  NAND2_X1 U998 ( .A1(n641), .A2(n1054), .ZN(n1053) );
  NAND2_X1 U999 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
  NAND2_X1 U1000 ( .A1(n1057), .A2(n614), .ZN(n1056) );
  NOR2_X1 U1001 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
  NOR2_X1 U1002 ( .A1(b_26_), .A2(n1060), .ZN(n1059) );
  NOR2_X1 U1003 ( .A1(n1061), .A2(n986), .ZN(n1058) );
  NAND2_X1 U1004 ( .A1(n604), .A2(n613), .ZN(n986) );
  NOR2_X1 U1005 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
  INV_X1 U1006 ( .A(n603), .ZN(n1063) );
  NOR2_X1 U1007 ( .A1(b_28_), .A2(n1064), .ZN(n1062) );
  INV_X1 U1008 ( .A(n982), .ZN(n1055) );
  NAND2_X1 U1009 ( .A1(n622), .A2(n631), .ZN(n982) );
  NOR2_X1 U1010 ( .A1(b_25_), .A2(n1065), .ZN(n1052) );
  AND2_X1 U1011 ( .A1(n1066), .A2(a_23_), .ZN(n1046) );
  AND2_X1 U1012 ( .A1(n1067), .A2(a_21_), .ZN(n1041) );
  AND2_X1 U1013 ( .A1(n694), .A2(n703), .ZN(n970) );
  NOR2_X1 U1014 ( .A1(b_17_), .A2(n1068), .ZN(n1032) );
  NOR2_X1 U1015 ( .A1(b_15_), .A2(n1069), .ZN(n1026) );
  AND2_X1 U1016 ( .A1(n784), .A2(n793), .ZN(n976) );
  NOR2_X1 U1017 ( .A1(b_7_), .A2(n1070), .ZN(n1004) );
  INV_X1 U1018 ( .A(n973), .ZN(n997) );
  NAND2_X1 U1019 ( .A1(n820), .A2(n829), .ZN(n973) );
  NAND2_X1 U1020 ( .A1(n1071), .A2(n1072), .ZN(n987) );
  NAND2_X1 U1021 ( .A1(n847), .A2(n846), .ZN(n1072) );
  NAND2_X1 U1022 ( .A1(n1073), .A2(n838), .ZN(n846) );
  NAND2_X1 U1023 ( .A1(b_2_), .A2(n1074), .ZN(n838) );
  NAND2_X1 U1024 ( .A1(n837), .A2(n839), .ZN(n1073) );
  OR2_X1 U1025 ( .A1(n1074), .A2(b_2_), .ZN(n839) );
  INV_X1 U1026 ( .A(a_2_), .ZN(n1074) );
  NAND2_X1 U1027 ( .A1(n829), .A2(n1075), .ZN(n837) );
  NAND2_X1 U1028 ( .A1(n830), .A2(n828), .ZN(n1075) );
  NAND2_X1 U1029 ( .A1(n820), .A2(n1076), .ZN(n828) );
  NAND2_X1 U1030 ( .A1(n821), .A2(n819), .ZN(n1076) );
  NAND2_X1 U1031 ( .A1(n811), .A2(n1077), .ZN(n819) );
  NAND2_X1 U1032 ( .A1(n812), .A2(n810), .ZN(n1077) );
  NAND2_X1 U1033 ( .A1(n802), .A2(n1078), .ZN(n810) );
  NAND2_X1 U1034 ( .A1(n803), .A2(n801), .ZN(n1078) );
  NAND2_X1 U1035 ( .A1(n793), .A2(n1079), .ZN(n801) );
  NAND2_X1 U1036 ( .A1(n794), .A2(n792), .ZN(n1079) );
  NAND2_X1 U1037 ( .A1(n784), .A2(n1080), .ZN(n792) );
  NAND2_X1 U1038 ( .A1(n785), .A2(n783), .ZN(n1080) );
  NAND2_X1 U1039 ( .A1(n775), .A2(n1081), .ZN(n783) );
  NAND2_X1 U1040 ( .A1(n776), .A2(n774), .ZN(n1081) );
  NAND2_X1 U1041 ( .A1(n766), .A2(n1082), .ZN(n774) );
  NAND2_X1 U1042 ( .A1(n767), .A2(n765), .ZN(n1082) );
  NAND2_X1 U1043 ( .A1(n757), .A2(n1083), .ZN(n765) );
  NAND2_X1 U1044 ( .A1(n758), .A2(n756), .ZN(n1083) );
  NAND2_X1 U1045 ( .A1(n748), .A2(n1084), .ZN(n756) );
  NAND2_X1 U1046 ( .A1(n749), .A2(n747), .ZN(n1084) );
  NAND2_X1 U1047 ( .A1(n739), .A2(n1085), .ZN(n747) );
  NAND2_X1 U1048 ( .A1(n740), .A2(n738), .ZN(n1085) );
  NAND2_X1 U1049 ( .A1(n730), .A2(n1086), .ZN(n738) );
  NAND2_X1 U1050 ( .A1(n731), .A2(n729), .ZN(n1086) );
  NAND2_X1 U1051 ( .A1(n721), .A2(n1087), .ZN(n729) );
  NAND2_X1 U1052 ( .A1(n722), .A2(n720), .ZN(n1087) );
  NAND2_X1 U1053 ( .A1(n712), .A2(n1088), .ZN(n720) );
  NAND2_X1 U1054 ( .A1(n713), .A2(n711), .ZN(n1088) );
  NAND2_X1 U1055 ( .A1(n703), .A2(n1089), .ZN(n711) );
  NAND2_X1 U1056 ( .A1(n704), .A2(n702), .ZN(n1089) );
  NAND2_X1 U1057 ( .A1(n694), .A2(n1090), .ZN(n702) );
  NAND2_X1 U1058 ( .A1(n695), .A2(n693), .ZN(n1090) );
  NAND2_X1 U1059 ( .A1(n685), .A2(n1091), .ZN(n693) );
  NAND2_X1 U1060 ( .A1(n686), .A2(n684), .ZN(n1091) );
  NAND2_X1 U1061 ( .A1(n676), .A2(n1092), .ZN(n684) );
  NAND2_X1 U1062 ( .A1(n677), .A2(n675), .ZN(n1092) );
  NAND2_X1 U1063 ( .A1(n667), .A2(n1093), .ZN(n675) );
  NAND2_X1 U1064 ( .A1(n668), .A2(n666), .ZN(n1093) );
  NAND2_X1 U1065 ( .A1(n658), .A2(n1094), .ZN(n666) );
  NAND2_X1 U1066 ( .A1(n659), .A2(n657), .ZN(n1094) );
  NAND2_X1 U1067 ( .A1(n649), .A2(n1095), .ZN(n657) );
  NAND2_X1 U1068 ( .A1(n650), .A2(n648), .ZN(n1095) );
  NAND2_X1 U1069 ( .A1(n640), .A2(n1096), .ZN(n648) );
  NAND2_X1 U1070 ( .A1(n641), .A2(n639), .ZN(n1096) );
  NAND2_X1 U1071 ( .A1(n631), .A2(n1097), .ZN(n639) );
  NAND2_X1 U1072 ( .A1(n632), .A2(n630), .ZN(n1097) );
  NAND2_X1 U1073 ( .A1(n622), .A2(n1098), .ZN(n630) );
  NAND2_X1 U1074 ( .A1(n623), .A2(n621), .ZN(n1098) );
  NAND2_X1 U1075 ( .A1(n613), .A2(n1099), .ZN(n621) );
  NAND2_X1 U1076 ( .A1(n614), .A2(n612), .ZN(n1099) );
  NAND2_X1 U1077 ( .A1(n604), .A2(n1100), .ZN(n612) );
  NAND2_X1 U1078 ( .A1(n605), .A2(n603), .ZN(n1100) );
  NAND2_X1 U1079 ( .A1(n595), .A2(n1101), .ZN(n603) );
  NAND2_X1 U1080 ( .A1(n596), .A2(n594), .ZN(n1101) );
  NAND2_X1 U1081 ( .A1(n572), .A2(n1102), .ZN(n594) );
  NAND2_X1 U1082 ( .A1(n1103), .A2(n573), .ZN(n1102) );
  OR2_X1 U1083 ( .A1(n945), .A2(b_30_), .ZN(n573) );
  NAND2_X1 U1084 ( .A1(a_31_), .A2(n580), .ZN(n1103) );
  INV_X1 U1085 ( .A(b_31_), .ZN(n580) );
  NAND2_X1 U1086 ( .A1(b_30_), .A2(n945), .ZN(n572) );
  INV_X1 U1087 ( .A(a_30_), .ZN(n945) );
  NAND2_X1 U1088 ( .A1(a_29_), .A2(n1104), .ZN(n596) );
  INV_X1 U1089 ( .A(n959), .ZN(n595) );
  NOR2_X1 U1090 ( .A1(n1104), .A2(a_29_), .ZN(n959) );
  INV_X1 U1091 ( .A(b_29_), .ZN(n1104) );
  NAND2_X1 U1092 ( .A1(a_28_), .A2(n1105), .ZN(n605) );
  INV_X1 U1093 ( .A(b_28_), .ZN(n1105) );
  NAND2_X1 U1094 ( .A1(b_28_), .A2(n1064), .ZN(n604) );
  INV_X1 U1095 ( .A(a_28_), .ZN(n1064) );
  NAND2_X1 U1096 ( .A1(a_27_), .A2(n1106), .ZN(n614) );
  OR2_X1 U1097 ( .A1(n1106), .A2(a_27_), .ZN(n613) );
  INV_X1 U1098 ( .A(b_27_), .ZN(n1106) );
  NAND2_X1 U1099 ( .A1(a_26_), .A2(n1107), .ZN(n623) );
  INV_X1 U1100 ( .A(b_26_), .ZN(n1107) );
  NAND2_X1 U1101 ( .A1(b_26_), .A2(n1060), .ZN(n622) );
  INV_X1 U1102 ( .A(a_26_), .ZN(n1060) );
  NAND2_X1 U1103 ( .A1(a_25_), .A2(n1108), .ZN(n632) );
  INV_X1 U1104 ( .A(b_25_), .ZN(n1108) );
  NAND2_X1 U1105 ( .A1(b_25_), .A2(n1065), .ZN(n631) );
  INV_X1 U1106 ( .A(a_25_), .ZN(n1065) );
  NAND2_X1 U1107 ( .A1(a_24_), .A2(n1109), .ZN(n641) );
  OR2_X1 U1108 ( .A1(n1109), .A2(a_24_), .ZN(n640) );
  INV_X1 U1109 ( .A(b_24_), .ZN(n1109) );
  NAND2_X1 U1110 ( .A1(a_23_), .A2(n1066), .ZN(n650) );
  INV_X1 U1111 ( .A(n1050), .ZN(n649) );
  NOR2_X1 U1112 ( .A1(n1066), .A2(a_23_), .ZN(n1050) );
  INV_X1 U1113 ( .A(b_23_), .ZN(n1066) );
  NAND2_X1 U1114 ( .A1(a_22_), .A2(n1110), .ZN(n659) );
  INV_X1 U1115 ( .A(n955), .ZN(n658) );
  NOR2_X1 U1116 ( .A1(n1110), .A2(a_22_), .ZN(n955) );
  INV_X1 U1117 ( .A(b_22_), .ZN(n1110) );
  NAND2_X1 U1118 ( .A1(a_21_), .A2(n1067), .ZN(n668) );
  INV_X1 U1119 ( .A(n953), .ZN(n667) );
  NOR2_X1 U1120 ( .A1(n1067), .A2(a_21_), .ZN(n953) );
  INV_X1 U1121 ( .A(b_21_), .ZN(n1067) );
  NAND2_X1 U1122 ( .A1(a_20_), .A2(n1111), .ZN(n677) );
  OR2_X1 U1123 ( .A1(n1111), .A2(a_20_), .ZN(n676) );
  INV_X1 U1124 ( .A(b_20_), .ZN(n1111) );
  NAND2_X1 U1125 ( .A1(a_19_), .A2(n1112), .ZN(n686) );
  OR2_X1 U1126 ( .A1(n1112), .A2(a_19_), .ZN(n685) );
  INV_X1 U1127 ( .A(b_19_), .ZN(n1112) );
  NAND2_X1 U1128 ( .A1(a_18_), .A2(n1113), .ZN(n695) );
  INV_X1 U1129 ( .A(b_18_), .ZN(n1113) );
  NAND2_X1 U1130 ( .A1(b_18_), .A2(n1039), .ZN(n694) );
  INV_X1 U1131 ( .A(a_18_), .ZN(n1039) );
  NAND2_X1 U1132 ( .A1(a_17_), .A2(n1114), .ZN(n704) );
  INV_X1 U1133 ( .A(b_17_), .ZN(n1114) );
  NAND2_X1 U1134 ( .A1(b_17_), .A2(n1068), .ZN(n703) );
  INV_X1 U1135 ( .A(a_17_), .ZN(n1068) );
  NAND2_X1 U1136 ( .A1(a_16_), .A2(n1115), .ZN(n713) );
  INV_X1 U1137 ( .A(n1030), .ZN(n712) );
  NOR2_X1 U1138 ( .A1(n1115), .A2(a_16_), .ZN(n1030) );
  INV_X1 U1139 ( .A(b_16_), .ZN(n1115) );
  NAND2_X1 U1140 ( .A1(a_15_), .A2(n1116), .ZN(n722) );
  INV_X1 U1141 ( .A(b_15_), .ZN(n1116) );
  NAND2_X1 U1142 ( .A1(b_15_), .A2(n1069), .ZN(n721) );
  INV_X1 U1143 ( .A(a_15_), .ZN(n1069) );
  NAND2_X1 U1144 ( .A1(a_14_), .A2(n1117), .ZN(n731) );
  OR2_X1 U1145 ( .A1(n1117), .A2(a_14_), .ZN(n730) );
  INV_X1 U1146 ( .A(b_14_), .ZN(n1117) );
  NAND2_X1 U1147 ( .A1(a_13_), .A2(n1118), .ZN(n740) );
  OR2_X1 U1148 ( .A1(n1118), .A2(a_13_), .ZN(n739) );
  INV_X1 U1149 ( .A(b_13_), .ZN(n1118) );
  NAND2_X1 U1150 ( .A1(a_12_), .A2(n1024), .ZN(n749) );
  INV_X1 U1151 ( .A(n1018), .ZN(n748) );
  NOR2_X1 U1152 ( .A1(n1024), .A2(a_12_), .ZN(n1018) );
  INV_X1 U1153 ( .A(b_12_), .ZN(n1024) );
  NAND2_X1 U1154 ( .A1(a_11_), .A2(n1119), .ZN(n758) );
  OR2_X1 U1155 ( .A1(n1119), .A2(a_11_), .ZN(n757) );
  INV_X1 U1156 ( .A(b_11_), .ZN(n1119) );
  NAND2_X1 U1157 ( .A1(a_10_), .A2(n1017), .ZN(n767) );
  INV_X1 U1158 ( .A(n980), .ZN(n766) );
  NOR2_X1 U1159 ( .A1(n1017), .A2(a_10_), .ZN(n980) );
  INV_X1 U1160 ( .A(b_10_), .ZN(n1017) );
  NAND2_X1 U1161 ( .A1(a_9_), .A2(n1120), .ZN(n776) );
  INV_X1 U1162 ( .A(n961), .ZN(n775) );
  NOR2_X1 U1163 ( .A1(n1120), .A2(a_9_), .ZN(n961) );
  INV_X1 U1164 ( .A(b_9_), .ZN(n1120) );
  NAND2_X1 U1165 ( .A1(a_8_), .A2(n1121), .ZN(n785) );
  INV_X1 U1166 ( .A(b_8_), .ZN(n1121) );
  NAND2_X1 U1167 ( .A1(b_8_), .A2(n1011), .ZN(n784) );
  INV_X1 U1168 ( .A(a_8_), .ZN(n1011) );
  NAND2_X1 U1169 ( .A1(a_7_), .A2(n1122), .ZN(n794) );
  INV_X1 U1170 ( .A(b_7_), .ZN(n1122) );
  NAND2_X1 U1171 ( .A1(b_7_), .A2(n1070), .ZN(n793) );
  INV_X1 U1172 ( .A(a_7_), .ZN(n1070) );
  NAND2_X1 U1173 ( .A1(a_6_), .A2(n1123), .ZN(n803) );
  OR2_X1 U1174 ( .A1(n1123), .A2(a_6_), .ZN(n802) );
  INV_X1 U1175 ( .A(b_6_), .ZN(n1123) );
  NAND2_X1 U1176 ( .A1(a_5_), .A2(n1124), .ZN(n812) );
  OR2_X1 U1177 ( .A1(n1124), .A2(a_5_), .ZN(n811) );
  INV_X1 U1178 ( .A(b_5_), .ZN(n1124) );
  NAND2_X1 U1179 ( .A1(a_4_), .A2(n1125), .ZN(n821) );
  INV_X1 U1180 ( .A(b_4_), .ZN(n1125) );
  NAND2_X1 U1181 ( .A1(b_4_), .A2(n1002), .ZN(n820) );
  INV_X1 U1182 ( .A(a_4_), .ZN(n1002) );
  NAND2_X1 U1183 ( .A1(a_3_), .A2(n1126), .ZN(n830) );
  OR2_X1 U1184 ( .A1(n1126), .A2(a_3_), .ZN(n829) );
  INV_X1 U1185 ( .A(b_3_), .ZN(n1126) );
  NAND2_X1 U1186 ( .A1(a_1_), .A2(n857), .ZN(n847) );
  NOR2_X1 U1187 ( .A1(n993), .A2(n852), .ZN(n1071) );
  AND2_X1 U1188 ( .A1(n963), .A2(n988), .ZN(n852) );
  NAND2_X1 U1189 ( .A1(a_0_), .A2(n1127), .ZN(n988) );
  OR2_X1 U1190 ( .A1(n1127), .A2(a_0_), .ZN(n963) );
  INV_X1 U1191 ( .A(b_0_), .ZN(n1127) );
  NOR2_X1 U1192 ( .A1(n857), .A2(a_1_), .ZN(n993) );
  INV_X1 U1193 ( .A(b_1_), .ZN(n857) );
endmodule

