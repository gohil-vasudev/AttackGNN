module locked_c2670 (  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire new_n359_, new_n368_, new_n369_, new_n370_, new_n371_, new_n375_, new_n376_, new_n378_, new_n381_, new_n382_, new_n383_, new_n384_, new_n387_, new_n388_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n487_, new_n489_, new_n491_, new_n492_, new_n493_, new_n494_, new_n498_, new_n499_, new_n500_, new_n501_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n509_, new_n510_, new_n511_, new_n512_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n525_, new_n526_, new_n528_, new_n529_, new_n530_, new_n532_, new_n533_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_;
  XOR2_X1 g000 ( .A(G44), .B(KEYINPUT3), .Z(new_n359_) );
  INV_X1 g001 ( .A(new_n359_), .ZN(G218) );
  INV_X1 g002 ( .A(G132), .ZN(G219) );
  INV_X1 g003 ( .A(G82), .ZN(G220) );
  INV_X1 g004 ( .A(G96), .ZN(G221) );
  INV_X1 g005 ( .A(G69), .ZN(G235) );
  INV_X1 g006 ( .A(G120), .ZN(G236) );
  INV_X1 g007 ( .A(G57), .ZN(G237) );
  INV_X1 g008 ( .A(G108), .ZN(G238) );
  NAND2_X1 g009 ( .A1(G2078), .A2(G2084), .ZN(new_n368_) );
  XOR2_X1 g010 ( .A(new_n368_), .B(KEYINPUT20), .Z(new_n369_) );
  NAND2_X1 g011 ( .A1(new_n369_), .A2(G2090), .ZN(new_n370_) );
  XNOR2_X1 g012 ( .A(new_n370_), .B(KEYINPUT21), .ZN(new_n371_) );
  NAND2_X1 g013 ( .A1(new_n371_), .A2(G2072), .ZN(G158) );
  NAND3_X1 g014 ( .A1(G2), .A2(G15), .A3(G661), .ZN(G259) );
  AND2_X1 g015 ( .A1(G94), .A2(G452), .ZN(G173) );
  NAND2_X1 g016 ( .A1(G7), .A2(G661), .ZN(new_n375_) );
  XOR2_X1 g017 ( .A(new_n375_), .B(KEYINPUT10), .Z(new_n376_) );
  INV_X1 g018 ( .A(new_n376_), .ZN(G223) );
  NAND2_X1 g019 ( .A1(new_n376_), .A2(G567), .ZN(new_n378_) );
  XOR2_X1 g020 ( .A(new_n378_), .B(KEYINPUT11), .Z(G234) );
  NAND2_X1 g021 ( .A1(new_n376_), .A2(G2106), .ZN(G217) );
  NAND2_X1 g022 ( .A1(G82), .A2(G132), .ZN(new_n381_) );
  XOR2_X1 g023 ( .A(new_n381_), .B(KEYINPUT22), .Z(new_n382_) );
  NAND3_X1 g024 ( .A1(new_n382_), .A2(G96), .A3(new_n359_), .ZN(new_n383_) );
  NAND4_X1 g025 ( .A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n384_) );
  NOR2_X1 g026 ( .A1(new_n383_), .A2(new_n384_), .ZN(G325) );
  INV_X1 g027 ( .A(G325), .ZN(G261) );
  NAND2_X1 g028 ( .A1(new_n383_), .A2(G2106), .ZN(new_n387_) );
  NAND2_X1 g029 ( .A1(new_n384_), .A2(G567), .ZN(new_n388_) );
  AND2_X1 g030 ( .A1(new_n387_), .A2(new_n388_), .ZN(G319) );
  INV_X1 g031 ( .A(KEYINPUT23), .ZN(new_n390_) );
  INV_X1 g032 ( .A(G2105), .ZN(new_n391_) );
  NAND3_X1 g033 ( .A1(new_n391_), .A2(G101), .A3(G2104), .ZN(new_n392_) );
  NAND2_X1 g034 ( .A1(new_n392_), .A2(new_n390_), .ZN(new_n393_) );
  NAND4_X1 g035 ( .A1(new_n391_), .A2(G101), .A3(G2104), .A4(KEYINPUT23), .ZN(new_n394_) );
  NAND2_X1 g036 ( .A1(new_n393_), .A2(new_n394_), .ZN(new_n395_) );
  INV_X1 g037 ( .A(KEYINPUT17), .ZN(new_n396_) );
  INV_X1 g038 ( .A(G2104), .ZN(new_n397_) );
  NAND2_X1 g039 ( .A1(new_n397_), .A2(new_n391_), .ZN(new_n398_) );
  NAND2_X1 g040 ( .A1(new_n398_), .A2(new_n396_), .ZN(new_n399_) );
  NAND3_X1 g041 ( .A1(new_n397_), .A2(new_n391_), .A3(KEYINPUT17), .ZN(new_n400_) );
  NAND3_X1 g042 ( .A1(new_n399_), .A2(G137), .A3(new_n400_), .ZN(new_n401_) );
  NAND2_X1 g043 ( .A1(new_n401_), .A2(new_n395_), .ZN(new_n402_) );
  NAND3_X1 g044 ( .A1(new_n397_), .A2(G125), .A3(G2105), .ZN(new_n403_) );
  NAND3_X1 g045 ( .A1(G113), .A2(G2104), .A3(G2105), .ZN(new_n404_) );
  NAND2_X1 g046 ( .A1(new_n403_), .A2(new_n404_), .ZN(new_n405_) );
  NOR2_X1 g047 ( .A1(new_n402_), .A2(new_n405_), .ZN(G160) );
  NAND2_X1 g048 ( .A1(new_n399_), .A2(new_n400_), .ZN(new_n407_) );
  INV_X1 g049 ( .A(new_n407_), .ZN(new_n408_) );
  NAND2_X1 g050 ( .A1(new_n408_), .A2(G136), .ZN(new_n409_) );
  NOR2_X1 g051 ( .A1(new_n391_), .A2(G2104), .ZN(new_n410_) );
  AND2_X1 g052 ( .A1(new_n410_), .A2(G124), .ZN(new_n411_) );
  NAND2_X1 g053 ( .A1(new_n411_), .A2(KEYINPUT44), .ZN(new_n412_) );
  OR2_X1 g054 ( .A1(new_n411_), .A2(KEYINPUT44), .ZN(new_n413_) );
  NOR2_X1 g055 ( .A1(new_n397_), .A2(G2105), .ZN(new_n414_) );
  NAND2_X1 g056 ( .A1(new_n414_), .A2(G100), .ZN(new_n415_) );
  NOR2_X1 g057 ( .A1(new_n397_), .A2(new_n391_), .ZN(new_n416_) );
  NAND2_X1 g058 ( .A1(new_n416_), .A2(G112), .ZN(new_n417_) );
  AND2_X1 g059 ( .A1(new_n417_), .A2(new_n415_), .ZN(new_n418_) );
  AND4_X1 g060 ( .A1(new_n409_), .A2(new_n412_), .A3(new_n413_), .A4(new_n418_), .ZN(G162) );
  NAND3_X1 g061 ( .A1(new_n399_), .A2(G138), .A3(new_n400_), .ZN(new_n420_) );
  NAND3_X1 g062 ( .A1(G114), .A2(G2104), .A3(G2105), .ZN(new_n421_) );
  NAND3_X1 g063 ( .A1(new_n391_), .A2(G102), .A3(G2104), .ZN(new_n422_) );
  NAND3_X1 g064 ( .A1(new_n397_), .A2(G126), .A3(G2105), .ZN(new_n423_) );
  AND3_X1 g065 ( .A1(new_n422_), .A2(new_n423_), .A3(new_n421_), .ZN(new_n424_) );
  NAND2_X1 g066 ( .A1(new_n420_), .A2(new_n424_), .ZN(new_n425_) );
  INV_X1 g067 ( .A(new_n425_), .ZN(G164) );
  INV_X1 g068 ( .A(G543), .ZN(new_n427_) );
  NAND2_X1 g069 ( .A1(new_n427_), .A2(G651), .ZN(new_n428_) );
  NAND2_X1 g070 ( .A1(new_n428_), .A2(KEYINPUT1), .ZN(new_n429_) );
  INV_X1 g071 ( .A(KEYINPUT1), .ZN(new_n430_) );
  NAND3_X1 g072 ( .A1(new_n427_), .A2(new_n430_), .A3(G651), .ZN(new_n431_) );
  NAND2_X1 g073 ( .A1(new_n429_), .A2(new_n431_), .ZN(new_n432_) );
  NAND2_X1 g074 ( .A1(new_n432_), .A2(G62), .ZN(new_n433_) );
  NOR2_X1 g075 ( .A1(G543), .A2(G651), .ZN(new_n434_) );
  NAND2_X1 g076 ( .A1(new_n434_), .A2(G88), .ZN(new_n435_) );
  INV_X1 g077 ( .A(G651), .ZN(new_n436_) );
  XOR2_X1 g078 ( .A(G543), .B(KEYINPUT0), .Z(new_n437_) );
  NOR2_X1 g079 ( .A1(new_n437_), .A2(new_n436_), .ZN(new_n438_) );
  NAND2_X1 g080 ( .A1(new_n438_), .A2(G75), .ZN(new_n439_) );
  NOR2_X1 g081 ( .A1(new_n437_), .A2(G651), .ZN(new_n440_) );
  NAND2_X1 g082 ( .A1(new_n440_), .A2(G50), .ZN(new_n441_) );
  NAND4_X1 g083 ( .A1(new_n439_), .A2(new_n441_), .A3(new_n433_), .A4(new_n435_), .ZN(G303) );
  INV_X1 g084 ( .A(G303), .ZN(G166) );
  INV_X1 g085 ( .A(KEYINPUT7), .ZN(new_n444_) );
  NAND2_X1 g086 ( .A1(new_n440_), .A2(G51), .ZN(new_n445_) );
  NAND2_X1 g087 ( .A1(new_n432_), .A2(G63), .ZN(new_n446_) );
  NAND2_X1 g088 ( .A1(new_n445_), .A2(new_n446_), .ZN(new_n447_) );
  XOR2_X1 g089 ( .A(new_n447_), .B(KEYINPUT6), .Z(new_n448_) );
  NAND2_X1 g090 ( .A1(new_n438_), .A2(G76), .ZN(new_n449_) );
  NAND2_X1 g091 ( .A1(new_n434_), .A2(G89), .ZN(new_n450_) );
  XNOR2_X1 g092 ( .A(new_n450_), .B(KEYINPUT4), .ZN(new_n451_) );
  NAND2_X1 g093 ( .A1(new_n449_), .A2(new_n451_), .ZN(new_n452_) );
  XNOR2_X1 g094 ( .A(new_n452_), .B(KEYINPUT5), .ZN(new_n453_) );
  NAND2_X1 g095 ( .A1(new_n448_), .A2(new_n453_), .ZN(new_n454_) );
  XNOR2_X1 g096 ( .A(new_n454_), .B(new_n444_), .ZN(new_n455_) );
  INV_X1 g097 ( .A(new_n455_), .ZN(G168) );
  NAND2_X1 g098 ( .A1(new_n438_), .A2(G77), .ZN(new_n457_) );
  NAND2_X1 g099 ( .A1(new_n434_), .A2(G90), .ZN(new_n458_) );
  AND2_X1 g100 ( .A1(new_n457_), .A2(new_n458_), .ZN(new_n459_) );
  NAND2_X1 g101 ( .A1(new_n459_), .A2(KEYINPUT9), .ZN(new_n460_) );
  OR2_X1 g102 ( .A1(new_n459_), .A2(KEYINPUT9), .ZN(new_n461_) );
  NAND2_X1 g103 ( .A1(new_n440_), .A2(G52), .ZN(new_n462_) );
  NAND2_X1 g104 ( .A1(new_n432_), .A2(G64), .ZN(new_n463_) );
  AND4_X1 g105 ( .A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .A4(new_n463_), .ZN(G171) );
  NAND3_X1 g106 ( .A1(new_n427_), .A2(new_n436_), .A3(G81), .ZN(new_n465_) );
  NAND2_X1 g107 ( .A1(new_n465_), .A2(KEYINPUT12), .ZN(new_n466_) );
  INV_X1 g108 ( .A(KEYINPUT12), .ZN(new_n467_) );
  NAND3_X1 g109 ( .A1(new_n434_), .A2(G81), .A3(new_n467_), .ZN(new_n468_) );
  NAND2_X1 g110 ( .A1(new_n466_), .A2(new_n468_), .ZN(new_n469_) );
  XNOR2_X1 g111 ( .A(G543), .B(KEYINPUT0), .ZN(new_n470_) );
  AND2_X1 g112 ( .A1(G68), .A2(G651), .ZN(new_n471_) );
  NAND2_X1 g113 ( .A1(new_n470_), .A2(new_n471_), .ZN(new_n472_) );
  NAND2_X1 g114 ( .A1(new_n469_), .A2(new_n472_), .ZN(new_n473_) );
  NAND2_X1 g115 ( .A1(new_n473_), .A2(KEYINPUT13), .ZN(new_n474_) );
  INV_X1 g116 ( .A(KEYINPUT13), .ZN(new_n475_) );
  NAND3_X1 g117 ( .A1(new_n469_), .A2(new_n475_), .A3(new_n472_), .ZN(new_n476_) );
  NAND2_X1 g118 ( .A1(new_n474_), .A2(new_n476_), .ZN(new_n477_) );
  NAND3_X1 g119 ( .A1(new_n470_), .A2(G43), .A3(new_n436_), .ZN(new_n478_) );
  NAND2_X1 g120 ( .A1(new_n432_), .A2(G56), .ZN(new_n479_) );
  NAND2_X1 g121 ( .A1(new_n479_), .A2(KEYINPUT14), .ZN(new_n480_) );
  INV_X1 g122 ( .A(KEYINPUT14), .ZN(new_n481_) );
  NAND3_X1 g123 ( .A1(new_n432_), .A2(G56), .A3(new_n481_), .ZN(new_n482_) );
  NAND2_X1 g124 ( .A1(new_n480_), .A2(new_n482_), .ZN(new_n483_) );
  NAND3_X1 g125 ( .A1(new_n477_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n484_) );
  INV_X1 g126 ( .A(new_n484_), .ZN(new_n485_) );
  NAND2_X1 g127 ( .A1(new_n485_), .A2(G860), .ZN(G153) );
  AND3_X1 g128 ( .A1(G319), .A2(G483), .A3(G661), .ZN(new_n487_) );
  NAND2_X1 g129 ( .A1(new_n487_), .A2(G36), .ZN(G176) );
  NAND2_X1 g130 ( .A1(G1), .A2(G3), .ZN(new_n489_) );
  NAND2_X1 g131 ( .A1(new_n487_), .A2(new_n489_), .ZN(G188) );
  NAND2_X1 g132 ( .A1(new_n432_), .A2(G65), .ZN(new_n491_) );
  NAND2_X1 g133 ( .A1(new_n434_), .A2(G91), .ZN(new_n492_) );
  NAND2_X1 g134 ( .A1(new_n440_), .A2(G53), .ZN(new_n493_) );
  NAND2_X1 g135 ( .A1(new_n438_), .A2(G78), .ZN(new_n494_) );
  NAND4_X1 g136 ( .A1(new_n493_), .A2(new_n494_), .A3(new_n491_), .A4(new_n492_), .ZN(G299) );
  INV_X1 g137 ( .A(G171), .ZN(G301) );
  XNOR2_X1 g138 ( .A(new_n455_), .B(KEYINPUT8), .ZN(G286) );
  INV_X1 g139 ( .A(new_n432_), .ZN(new_n498_) );
  NAND2_X1 g140 ( .A1(new_n440_), .A2(G49), .ZN(new_n499_) );
  NAND2_X1 g141 ( .A1(new_n437_), .A2(G87), .ZN(new_n500_) );
  NAND2_X1 g142 ( .A1(G74), .A2(G651), .ZN(new_n501_) );
  NAND4_X1 g143 ( .A1(new_n499_), .A2(new_n498_), .A3(new_n500_), .A4(new_n501_), .ZN(G288) );
  NAND2_X1 g144 ( .A1(new_n432_), .A2(G61), .ZN(new_n503_) );
  NAND2_X1 g145 ( .A1(new_n434_), .A2(G86), .ZN(new_n504_) );
  NAND2_X1 g146 ( .A1(new_n440_), .A2(G48), .ZN(new_n505_) );
  NAND2_X1 g147 ( .A1(new_n438_), .A2(G73), .ZN(new_n506_) );
  XNOR2_X1 g148 ( .A(new_n506_), .B(KEYINPUT2), .ZN(new_n507_) );
  NAND4_X1 g149 ( .A1(new_n507_), .A2(new_n503_), .A3(new_n504_), .A4(new_n505_), .ZN(G305) );
  NAND2_X1 g150 ( .A1(new_n434_), .A2(G85), .ZN(new_n509_) );
  NAND2_X1 g151 ( .A1(new_n432_), .A2(G60), .ZN(new_n510_) );
  NAND2_X1 g152 ( .A1(new_n440_), .A2(G47), .ZN(new_n511_) );
  NAND2_X1 g153 ( .A1(new_n438_), .A2(G72), .ZN(new_n512_) );
  NAND4_X1 g154 ( .A1(new_n511_), .A2(new_n512_), .A3(new_n509_), .A4(new_n510_), .ZN(G290) );
  INV_X1 g155 ( .A(G868), .ZN(new_n514_) );
  NAND2_X1 g156 ( .A1(new_n432_), .A2(G66), .ZN(new_n515_) );
  NAND2_X1 g157 ( .A1(new_n438_), .A2(G79), .ZN(new_n516_) );
  NAND3_X1 g158 ( .A1(new_n470_), .A2(G54), .A3(new_n436_), .ZN(new_n517_) );
  NAND2_X1 g159 ( .A1(new_n434_), .A2(G92), .ZN(new_n518_) );
  NAND4_X1 g160 ( .A1(new_n516_), .A2(new_n515_), .A3(new_n517_), .A4(new_n518_), .ZN(new_n519_) );
  XNOR2_X1 g161 ( .A(new_n519_), .B(KEYINPUT15), .ZN(new_n520_) );
  INV_X1 g162 ( .A(new_n520_), .ZN(new_n521_) );
  NAND2_X1 g163 ( .A1(new_n521_), .A2(new_n514_), .ZN(new_n522_) );
  NAND2_X1 g164 ( .A1(G301), .A2(G868), .ZN(new_n523_) );
  NAND2_X1 g165 ( .A1(new_n523_), .A2(new_n522_), .ZN(G284) );
  NOR2_X1 g166 ( .A1(G286), .A2(new_n514_), .ZN(new_n525_) );
  NOR2_X1 g167 ( .A1(G299), .A2(G868), .ZN(new_n526_) );
  NOR2_X1 g168 ( .A1(new_n525_), .A2(new_n526_), .ZN(G297) );
  INV_X1 g169 ( .A(G860), .ZN(new_n528_) );
  NAND2_X1 g170 ( .A1(new_n528_), .A2(G559), .ZN(new_n529_) );
  NAND2_X1 g171 ( .A1(new_n520_), .A2(new_n529_), .ZN(new_n530_) );
  XNOR2_X1 g172 ( .A(new_n530_), .B(KEYINPUT16), .ZN(G148) );
  NOR3_X1 g173 ( .A1(new_n521_), .A2(G559), .A3(new_n514_), .ZN(new_n532_) );
  NOR2_X1 g174 ( .A1(new_n484_), .A2(G868), .ZN(new_n533_) );
  NOR2_X1 g175 ( .A1(new_n532_), .A2(new_n533_), .ZN(G282) );
  NAND2_X1 g176 ( .A1(new_n410_), .A2(G123), .ZN(new_n535_) );
  XNOR2_X1 g177 ( .A(new_n535_), .B(KEYINPUT18), .ZN(new_n536_) );
  NAND2_X1 g178 ( .A1(new_n408_), .A2(G135), .ZN(new_n537_) );
  NAND2_X1 g179 ( .A1(new_n416_), .A2(G111), .ZN(new_n538_) );
  NAND2_X1 g180 ( .A1(new_n414_), .A2(G99), .ZN(new_n539_) );
  NAND4_X1 g181 ( .A1(new_n537_), .A2(new_n536_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_) );
  XNOR2_X1 g182 ( .A(new_n540_), .B(G2096), .ZN(new_n541_) );
  OR2_X1 g183 ( .A1(new_n541_), .A2(G2100), .ZN(G156) );
  XOR2_X1 g184 ( .A(G2430), .B(G2454), .Z(new_n543_) );
  XNOR2_X1 g185 ( .A(G1341), .B(G1348), .ZN(new_n544_) );
  XNOR2_X1 g186 ( .A(new_n543_), .B(new_n544_), .ZN(new_n545_) );
  XNOR2_X1 g187 ( .A(G2435), .B(G2438), .ZN(new_n546_) );
  XNOR2_X1 g188 ( .A(new_n545_), .B(new_n546_), .ZN(new_n547_) );
  XNOR2_X1 g189 ( .A(G2446), .B(G2451), .ZN(new_n548_) );
  XNOR2_X1 g190 ( .A(G2427), .B(G2443), .ZN(new_n549_) );
  XNOR2_X1 g191 ( .A(new_n548_), .B(new_n549_), .ZN(new_n550_) );
  OR2_X1 g192 ( .A1(new_n547_), .A2(new_n550_), .ZN(new_n551_) );
  NAND2_X1 g193 ( .A1(new_n547_), .A2(new_n550_), .ZN(new_n552_) );
  NAND3_X1 g194 ( .A1(new_n551_), .A2(G14), .A3(new_n552_), .ZN(new_n553_) );
  INV_X1 g195 ( .A(new_n553_), .ZN(G401) );
  XOR2_X1 g196 ( .A(G2090), .B(KEYINPUT42), .Z(new_n555_) );
  XNOR2_X1 g197 ( .A(G2067), .B(G2072), .ZN(new_n556_) );
  XNOR2_X1 g198 ( .A(new_n555_), .B(new_n556_), .ZN(new_n557_) );
  XNOR2_X1 g199 ( .A(G2096), .B(G2100), .ZN(new_n558_) );
  XNOR2_X1 g200 ( .A(G2678), .B(KEYINPUT43), .ZN(new_n559_) );
  XNOR2_X1 g201 ( .A(new_n558_), .B(new_n559_), .ZN(new_n560_) );
  XNOR2_X1 g202 ( .A(new_n557_), .B(new_n560_), .ZN(new_n561_) );
  XNOR2_X1 g203 ( .A(G2078), .B(G2084), .ZN(new_n562_) );
  XNOR2_X1 g204 ( .A(new_n561_), .B(new_n562_), .ZN(G227) );
  XOR2_X1 g205 ( .A(G1976), .B(G1981), .Z(new_n564_) );
  XNOR2_X1 g206 ( .A(G1956), .B(G1966), .ZN(new_n565_) );
  XNOR2_X1 g207 ( .A(new_n564_), .B(new_n565_), .ZN(new_n566_) );
  XNOR2_X1 g208 ( .A(new_n566_), .B(G2474), .ZN(new_n567_) );
  XOR2_X1 g209 ( .A(G1991), .B(G1996), .Z(new_n568_) );
  XNOR2_X1 g210 ( .A(new_n567_), .B(new_n568_), .ZN(new_n569_) );
  XOR2_X1 g211 ( .A(G1971), .B(KEYINPUT41), .Z(new_n570_) );
  XNOR2_X1 g212 ( .A(G1961), .B(G1986), .ZN(new_n571_) );
  XNOR2_X1 g213 ( .A(new_n570_), .B(new_n571_), .ZN(new_n572_) );
  XNOR2_X1 g214 ( .A(new_n569_), .B(new_n572_), .ZN(G229) );
  INV_X1 g215 ( .A(KEYINPUT51), .ZN(new_n574_) );
  NAND2_X1 g216 ( .A1(new_n408_), .A2(G141), .ZN(new_n575_) );
  AND2_X1 g217 ( .A1(new_n414_), .A2(G105), .ZN(new_n576_) );
  OR2_X1 g218 ( .A1(new_n576_), .A2(KEYINPUT38), .ZN(new_n577_) );
  NAND2_X1 g219 ( .A1(new_n576_), .A2(KEYINPUT38), .ZN(new_n578_) );
  NAND2_X1 g220 ( .A1(new_n410_), .A2(G129), .ZN(new_n579_) );
  NAND2_X1 g221 ( .A1(new_n416_), .A2(G117), .ZN(new_n580_) );
  AND2_X1 g222 ( .A1(new_n580_), .A2(new_n579_), .ZN(new_n581_) );
  NAND4_X1 g223 ( .A1(new_n575_), .A2(new_n577_), .A3(new_n578_), .A4(new_n581_), .ZN(new_n582_) );
  OR2_X1 g224 ( .A1(new_n582_), .A2(G1996), .ZN(new_n583_) );
  INV_X1 g225 ( .A(G2090), .ZN(new_n584_) );
  NAND2_X1 g226 ( .A1(G162), .A2(new_n584_), .ZN(new_n585_) );
  OR2_X1 g227 ( .A1(G162), .A2(new_n584_), .ZN(new_n586_) );
  NAND3_X1 g228 ( .A1(new_n586_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n587_) );
  OR2_X1 g229 ( .A1(new_n587_), .A2(new_n574_), .ZN(new_n588_) );
  NAND2_X1 g230 ( .A1(new_n408_), .A2(G139), .ZN(new_n589_) );
  NAND2_X1 g231 ( .A1(new_n414_), .A2(G103), .ZN(new_n590_) );
  NAND2_X1 g232 ( .A1(new_n410_), .A2(G127), .ZN(new_n591_) );
  NAND2_X1 g233 ( .A1(new_n416_), .A2(G115), .ZN(new_n592_) );
  NAND2_X1 g234 ( .A1(new_n592_), .A2(new_n591_), .ZN(new_n593_) );
  XNOR2_X1 g235 ( .A(new_n593_), .B(KEYINPUT47), .ZN(new_n594_) );
  NAND3_X1 g236 ( .A1(new_n594_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n595_) );
  OR2_X1 g237 ( .A1(new_n595_), .A2(G2072), .ZN(new_n596_) );
  NAND2_X1 g238 ( .A1(new_n595_), .A2(G2072), .ZN(new_n597_) );
  XOR2_X1 g239 ( .A(new_n425_), .B(G2078), .Z(new_n598_) );
  NAND3_X1 g240 ( .A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_) );
  XOR2_X1 g241 ( .A(new_n599_), .B(KEYINPUT50), .Z(new_n600_) );
  NAND2_X1 g242 ( .A1(new_n408_), .A2(G140), .ZN(new_n601_) );
  NAND2_X1 g243 ( .A1(new_n414_), .A2(G104), .ZN(new_n602_) );
  NAND2_X1 g244 ( .A1(new_n601_), .A2(new_n602_), .ZN(new_n603_) );
  OR2_X1 g245 ( .A1(new_n603_), .A2(KEYINPUT34), .ZN(new_n604_) );
  NAND2_X1 g246 ( .A1(new_n410_), .A2(G128), .ZN(new_n605_) );
  NAND2_X1 g247 ( .A1(new_n416_), .A2(G116), .ZN(new_n606_) );
  NAND2_X1 g248 ( .A1(new_n606_), .A2(new_n605_), .ZN(new_n607_) );
  XNOR2_X1 g249 ( .A(new_n607_), .B(KEYINPUT35), .ZN(new_n608_) );
  NAND2_X1 g250 ( .A1(new_n603_), .A2(KEYINPUT34), .ZN(new_n609_) );
  NAND3_X1 g251 ( .A1(new_n604_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_) );
  XNOR2_X1 g252 ( .A(new_n610_), .B(KEYINPUT36), .ZN(new_n611_) );
  XOR2_X1 g253 ( .A(G2067), .B(KEYINPUT37), .Z(new_n612_) );
  OR2_X1 g254 ( .A1(new_n611_), .A2(new_n612_), .ZN(new_n613_) );
  NAND2_X1 g255 ( .A1(new_n611_), .A2(new_n612_), .ZN(new_n614_) );
  NAND2_X1 g256 ( .A1(new_n587_), .A2(new_n574_), .ZN(new_n615_) );
  NAND2_X1 g257 ( .A1(new_n408_), .A2(G131), .ZN(new_n616_) );
  NAND2_X1 g258 ( .A1(new_n414_), .A2(G95), .ZN(new_n617_) );
  NAND2_X1 g259 ( .A1(new_n416_), .A2(G107), .ZN(new_n618_) );
  NAND2_X1 g260 ( .A1(new_n410_), .A2(G119), .ZN(new_n619_) );
  NAND4_X1 g261 ( .A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .A4(new_n619_), .ZN(new_n620_) );
  NAND2_X1 g262 ( .A1(new_n620_), .A2(G1991), .ZN(new_n621_) );
  NAND2_X1 g263 ( .A1(new_n582_), .A2(G1996), .ZN(new_n622_) );
  NAND2_X1 g264 ( .A1(new_n622_), .A2(new_n621_), .ZN(new_n623_) );
  INV_X1 g265 ( .A(G160), .ZN(new_n624_) );
  NOR2_X1 g266 ( .A1(new_n624_), .A2(G2084), .ZN(new_n625_) );
  NAND2_X1 g267 ( .A1(new_n624_), .A2(G2084), .ZN(new_n626_) );
  OR2_X1 g268 ( .A1(new_n620_), .A2(G1991), .ZN(new_n627_) );
  NAND3_X1 g269 ( .A1(new_n627_), .A2(new_n540_), .A3(new_n626_), .ZN(new_n628_) );
  NOR3_X1 g270 ( .A1(new_n628_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n629_) );
  AND3_X1 g271 ( .A1(new_n614_), .A2(new_n615_), .A3(new_n629_), .ZN(new_n630_) );
  NAND4_X1 g272 ( .A1(new_n630_), .A2(new_n588_), .A3(new_n600_), .A4(new_n613_), .ZN(new_n631_) );
  XNOR2_X1 g273 ( .A(new_n631_), .B(KEYINPUT52), .ZN(new_n632_) );
  OR2_X1 g274 ( .A1(new_n632_), .A2(KEYINPUT55), .ZN(new_n633_) );
  NAND2_X1 g275 ( .A1(new_n633_), .A2(G29), .ZN(new_n634_) );
  INV_X1 g276 ( .A(KEYINPUT57), .ZN(new_n635_) );
  NAND2_X1 g277 ( .A1(new_n455_), .A2(G1966), .ZN(new_n636_) );
  INV_X1 g278 ( .A(G1966), .ZN(new_n637_) );
  NAND2_X1 g279 ( .A1(G168), .A2(new_n637_), .ZN(new_n638_) );
  XOR2_X1 g280 ( .A(G305), .B(G1981), .Z(new_n639_) );
  NAND3_X1 g281 ( .A1(new_n638_), .A2(new_n636_), .A3(new_n639_), .ZN(new_n640_) );
  OR2_X1 g282 ( .A1(new_n640_), .A2(new_n635_), .ZN(new_n641_) );
  NAND2_X1 g283 ( .A1(new_n640_), .A2(new_n635_), .ZN(new_n642_) );
  XNOR2_X1 g284 ( .A(new_n484_), .B(G1341), .ZN(new_n643_) );
  XOR2_X1 g285 ( .A(new_n520_), .B(G1348), .Z(new_n644_) );
  XOR2_X1 g286 ( .A(G299), .B(G1956), .Z(new_n645_) );
  NAND2_X1 g287 ( .A1(G288), .A2(G1976), .ZN(new_n646_) );
  NAND2_X1 g288 ( .A1(G303), .A2(G1971), .ZN(new_n647_) );
  AND2_X1 g289 ( .A1(new_n647_), .A2(new_n646_), .ZN(new_n648_) );
  NOR2_X1 g290 ( .A1(G303), .A2(G1971), .ZN(new_n649_) );
  NOR2_X1 g291 ( .A1(G288), .A2(G1976), .ZN(new_n650_) );
  NOR2_X1 g292 ( .A1(new_n649_), .A2(new_n650_), .ZN(new_n651_) );
  XOR2_X1 g293 ( .A(G290), .B(G1986), .Z(new_n652_) );
  NAND4_X1 g294 ( .A1(new_n645_), .A2(new_n648_), .A3(new_n651_), .A4(new_n652_), .ZN(new_n653_) );
  INV_X1 g295 ( .A(G1961), .ZN(new_n654_) );
  XNOR2_X1 g296 ( .A(G171), .B(new_n654_), .ZN(new_n655_) );
  NOR4_X1 g297 ( .A1(new_n655_), .A2(new_n643_), .A3(new_n644_), .A4(new_n653_), .ZN(new_n656_) );
  NAND3_X1 g298 ( .A1(new_n641_), .A2(new_n642_), .A3(new_n656_), .ZN(new_n657_) );
  XNOR2_X1 g299 ( .A(G16), .B(KEYINPUT56), .ZN(new_n658_) );
  NAND2_X1 g300 ( .A1(new_n657_), .A2(new_n658_), .ZN(new_n659_) );
  INV_X1 g301 ( .A(G11), .ZN(new_n660_) );
  INV_X1 g302 ( .A(KEYINPUT53), .ZN(new_n661_) );
  NAND2_X1 g303 ( .A1(G33), .A2(G2072), .ZN(new_n662_) );
  AND2_X1 g304 ( .A1(G26), .A2(G2067), .ZN(new_n663_) );
  NOR2_X1 g305 ( .A1(G26), .A2(G2067), .ZN(new_n664_) );
  AND2_X1 g306 ( .A1(G32), .A2(G1996), .ZN(new_n665_) );
  NOR2_X1 g307 ( .A1(G32), .A2(G1996), .ZN(new_n666_) );
  NOR4_X1 g308 ( .A1(new_n663_), .A2(new_n665_), .A3(new_n664_), .A4(new_n666_), .ZN(new_n667_) );
  AND3_X1 g309 ( .A1(new_n667_), .A2(G28), .A3(new_n662_), .ZN(new_n668_) );
  INV_X1 g310 ( .A(G27), .ZN(new_n669_) );
  XNOR2_X1 g311 ( .A(G2078), .B(KEYINPUT25), .ZN(new_n670_) );
  NAND2_X1 g312 ( .A1(new_n670_), .A2(new_n669_), .ZN(new_n671_) );
  NOR2_X1 g313 ( .A1(new_n670_), .A2(new_n669_), .ZN(new_n672_) );
  NOR2_X1 g314 ( .A1(G25), .A2(G1991), .ZN(new_n673_) );
  NOR2_X1 g315 ( .A1(G33), .A2(G2072), .ZN(new_n674_) );
  AND2_X1 g316 ( .A1(G25), .A2(G1991), .ZN(new_n675_) );
  NOR4_X1 g317 ( .A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .A4(new_n675_), .ZN(new_n676_) );
  NAND3_X1 g318 ( .A1(new_n668_), .A2(new_n676_), .A3(new_n671_), .ZN(new_n677_) );
  NAND2_X1 g319 ( .A1(new_n677_), .A2(new_n661_), .ZN(new_n678_) );
  OR2_X1 g320 ( .A1(new_n677_), .A2(new_n661_), .ZN(new_n679_) );
  XNOR2_X1 g321 ( .A(G2084), .B(KEYINPUT54), .ZN(new_n680_) );
  NOR2_X1 g322 ( .A1(new_n680_), .A2(G34), .ZN(new_n681_) );
  XNOR2_X1 g323 ( .A(G35), .B(G2090), .ZN(new_n682_) );
  AND2_X1 g324 ( .A1(new_n680_), .A2(G34), .ZN(new_n683_) );
  NOR3_X1 g325 ( .A1(new_n683_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n684_) );
  NAND3_X1 g326 ( .A1(new_n679_), .A2(new_n678_), .A3(new_n684_), .ZN(new_n685_) );
  XNOR2_X1 g327 ( .A(new_n685_), .B(KEYINPUT55), .ZN(new_n686_) );
  NOR2_X1 g328 ( .A1(new_n686_), .A2(G29), .ZN(new_n687_) );
  XNOR2_X1 g329 ( .A(G1348), .B(KEYINPUT59), .ZN(new_n688_) );
  XNOR2_X1 g330 ( .A(new_n688_), .B(G4), .ZN(new_n689_) );
  XOR2_X1 g331 ( .A(G20), .B(G1956), .Z(new_n690_) );
  XOR2_X1 g332 ( .A(G6), .B(G1981), .Z(new_n691_) );
  XOR2_X1 g333 ( .A(G19), .B(G1341), .Z(new_n692_) );
  NAND4_X1 g334 ( .A1(new_n689_), .A2(new_n690_), .A3(new_n691_), .A4(new_n692_), .ZN(new_n693_) );
  XOR2_X1 g335 ( .A(new_n693_), .B(KEYINPUT60), .Z(new_n694_) );
  XOR2_X1 g336 ( .A(G23), .B(G1976), .Z(new_n695_) );
  XOR2_X1 g337 ( .A(G22), .B(G1971), .Z(new_n696_) );
  XOR2_X1 g338 ( .A(G24), .B(G1986), .Z(new_n697_) );
  NAND3_X1 g339 ( .A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_) );
  NOR2_X1 g340 ( .A1(new_n698_), .A2(KEYINPUT58), .ZN(new_n699_) );
  AND2_X1 g341 ( .A1(new_n698_), .A2(KEYINPUT58), .ZN(new_n700_) );
  XNOR2_X1 g342 ( .A(G21), .B(G1966), .ZN(new_n701_) );
  XNOR2_X1 g343 ( .A(G5), .B(G1961), .ZN(new_n702_) );
  NOR4_X1 g344 ( .A1(new_n700_), .A2(new_n699_), .A3(new_n701_), .A4(new_n702_), .ZN(new_n703_) );
  NAND2_X1 g345 ( .A1(new_n694_), .A2(new_n703_), .ZN(new_n704_) );
  XNOR2_X1 g346 ( .A(new_n704_), .B(KEYINPUT61), .ZN(new_n705_) );
  NOR2_X1 g347 ( .A1(new_n705_), .A2(G16), .ZN(new_n706_) );
  NOR3_X1 g348 ( .A1(new_n706_), .A2(new_n687_), .A3(new_n660_), .ZN(new_n707_) );
  NAND3_X1 g349 ( .A1(new_n634_), .A2(new_n659_), .A3(new_n707_), .ZN(new_n708_) );
  XNOR2_X1 g350 ( .A(new_n708_), .B(KEYINPUT62), .ZN(G150) );
  INV_X1 g351 ( .A(G150), .ZN(G311) );
  NAND2_X1 g352 ( .A1(new_n520_), .A2(G559), .ZN(new_n711_) );
  NAND2_X1 g353 ( .A1(new_n711_), .A2(new_n484_), .ZN(new_n712_) );
  NAND3_X1 g354 ( .A1(new_n520_), .A2(G559), .A3(new_n485_), .ZN(new_n713_) );
  NAND3_X1 g355 ( .A1(new_n712_), .A2(new_n528_), .A3(new_n713_), .ZN(new_n714_) );
  NAND2_X1 g356 ( .A1(new_n434_), .A2(G93), .ZN(new_n715_) );
  NAND2_X1 g357 ( .A1(new_n432_), .A2(G67), .ZN(new_n716_) );
  NAND2_X1 g358 ( .A1(new_n440_), .A2(G55), .ZN(new_n717_) );
  NAND2_X1 g359 ( .A1(new_n438_), .A2(G80), .ZN(new_n718_) );
  NAND4_X1 g360 ( .A1(new_n717_), .A2(new_n718_), .A3(new_n715_), .A4(new_n716_), .ZN(new_n719_) );
  XNOR2_X1 g361 ( .A(new_n714_), .B(new_n719_), .ZN(G145) );
  XNOR2_X1 g362 ( .A(new_n595_), .B(new_n624_), .ZN(new_n721_) );
  XNOR2_X1 g363 ( .A(new_n611_), .B(new_n721_), .ZN(new_n722_) );
  NAND2_X1 g364 ( .A1(new_n408_), .A2(G142), .ZN(new_n723_) );
  NAND2_X1 g365 ( .A1(new_n414_), .A2(G106), .ZN(new_n724_) );
  AND2_X1 g366 ( .A1(new_n723_), .A2(new_n724_), .ZN(new_n725_) );
  NAND2_X1 g367 ( .A1(new_n725_), .A2(KEYINPUT45), .ZN(new_n726_) );
  OR2_X1 g368 ( .A1(new_n725_), .A2(KEYINPUT45), .ZN(new_n727_) );
  NAND2_X1 g369 ( .A1(new_n410_), .A2(G130), .ZN(new_n728_) );
  NAND2_X1 g370 ( .A1(new_n416_), .A2(G118), .ZN(new_n729_) );
  NAND4_X1 g371 ( .A1(new_n727_), .A2(new_n726_), .A3(new_n728_), .A4(new_n729_), .ZN(new_n730_) );
  XNOR2_X1 g372 ( .A(new_n730_), .B(new_n582_), .ZN(new_n731_) );
  XNOR2_X1 g373 ( .A(new_n731_), .B(G162), .ZN(new_n732_) );
  XNOR2_X1 g374 ( .A(new_n732_), .B(new_n722_), .ZN(new_n733_) );
  XNOR2_X1 g375 ( .A(new_n540_), .B(new_n620_), .ZN(new_n734_) );
  XOR2_X1 g376 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(new_n735_) );
  XNOR2_X1 g377 ( .A(new_n734_), .B(new_n735_), .ZN(new_n736_) );
  XNOR2_X1 g378 ( .A(new_n736_), .B(G164), .ZN(new_n737_) );
  NOR2_X1 g379 ( .A1(new_n733_), .A2(new_n737_), .ZN(new_n738_) );
  AND2_X1 g380 ( .A1(new_n733_), .A2(new_n737_), .ZN(new_n739_) );
  NOR3_X1 g381 ( .A1(new_n739_), .A2(new_n738_), .A3(G37), .ZN(G395) );
  XOR2_X1 g382 ( .A(new_n484_), .B(G290), .Z(new_n741_) );
  XNOR2_X1 g383 ( .A(new_n741_), .B(G288), .ZN(new_n742_) );
  XNOR2_X1 g384 ( .A(G299), .B(KEYINPUT19), .ZN(new_n743_) );
  XOR2_X1 g385 ( .A(new_n743_), .B(G305), .Z(new_n744_) );
  XNOR2_X1 g386 ( .A(new_n742_), .B(new_n744_), .ZN(new_n745_) );
  XNOR2_X1 g387 ( .A(G303), .B(new_n719_), .ZN(new_n746_) );
  XNOR2_X1 g388 ( .A(new_n745_), .B(new_n746_), .ZN(new_n747_) );
  XOR2_X1 g389 ( .A(new_n747_), .B(new_n711_), .Z(new_n748_) );
  NAND2_X1 g390 ( .A1(new_n748_), .A2(G868), .ZN(new_n749_) );
  NAND2_X1 g391 ( .A1(new_n719_), .A2(new_n514_), .ZN(new_n750_) );
  NAND2_X1 g392 ( .A1(new_n749_), .A2(new_n750_), .ZN(G295) );
  INV_X1 g393 ( .A(G37), .ZN(new_n752_) );
  XNOR2_X1 g394 ( .A(G286), .B(new_n520_), .ZN(new_n753_) );
  XNOR2_X1 g395 ( .A(new_n747_), .B(new_n753_), .ZN(new_n754_) );
  OR2_X1 g396 ( .A1(new_n754_), .A2(G171), .ZN(new_n755_) );
  NAND2_X1 g397 ( .A1(new_n754_), .A2(G171), .ZN(new_n756_) );
  NAND3_X1 g398 ( .A1(new_n755_), .A2(new_n752_), .A3(new_n756_), .ZN(new_n757_) );
  INV_X1 g399 ( .A(new_n757_), .ZN(G397) );
  INV_X1 g400 ( .A(KEYINPUT33), .ZN(new_n759_) );
  INV_X1 g401 ( .A(KEYINPUT29), .ZN(new_n760_) );
  INV_X1 g402 ( .A(G1384), .ZN(new_n761_) );
  NAND2_X1 g403 ( .A1(new_n425_), .A2(new_n761_), .ZN(new_n762_) );
  INV_X1 g404 ( .A(G40), .ZN(new_n763_) );
  NOR2_X1 g405 ( .A1(new_n405_), .A2(new_n763_), .ZN(new_n764_) );
  NAND3_X1 g406 ( .A1(new_n764_), .A2(new_n401_), .A3(new_n395_), .ZN(new_n765_) );
  NOR2_X1 g407 ( .A1(new_n762_), .A2(new_n765_), .ZN(new_n766_) );
  INV_X1 g408 ( .A(new_n766_), .ZN(new_n767_) );
  NAND2_X1 g409 ( .A1(new_n767_), .A2(G1348), .ZN(new_n768_) );
  NAND2_X1 g410 ( .A1(new_n766_), .A2(G2067), .ZN(new_n769_) );
  NAND2_X1 g411 ( .A1(new_n768_), .A2(new_n769_), .ZN(new_n770_) );
  NAND3_X1 g412 ( .A1(new_n766_), .A2(G1996), .A3(KEYINPUT26), .ZN(new_n771_) );
  INV_X1 g413 ( .A(KEYINPUT26), .ZN(new_n772_) );
  NAND2_X1 g414 ( .A1(new_n766_), .A2(G1996), .ZN(new_n773_) );
  NAND2_X1 g415 ( .A1(new_n773_), .A2(new_n772_), .ZN(new_n774_) );
  INV_X1 g416 ( .A(G1341), .ZN(new_n775_) );
  NOR2_X1 g417 ( .A1(new_n766_), .A2(new_n775_), .ZN(new_n776_) );
  NOR2_X1 g418 ( .A1(new_n776_), .A2(new_n484_), .ZN(new_n777_) );
  NAND4_X1 g419 ( .A1(new_n777_), .A2(new_n520_), .A3(new_n771_), .A4(new_n774_), .ZN(new_n778_) );
  NAND2_X1 g420 ( .A1(new_n778_), .A2(new_n770_), .ZN(new_n779_) );
  NAND3_X1 g421 ( .A1(new_n777_), .A2(new_n771_), .A3(new_n774_), .ZN(new_n780_) );
  NAND2_X1 g422 ( .A1(new_n780_), .A2(new_n521_), .ZN(new_n781_) );
  NAND2_X1 g423 ( .A1(new_n779_), .A2(new_n781_), .ZN(new_n782_) );
  INV_X1 g424 ( .A(KEYINPUT27), .ZN(new_n783_) );
  NAND3_X1 g425 ( .A1(new_n766_), .A2(G2072), .A3(new_n783_), .ZN(new_n784_) );
  NAND2_X1 g426 ( .A1(new_n767_), .A2(G1956), .ZN(new_n785_) );
  NAND2_X1 g427 ( .A1(new_n766_), .A2(G2072), .ZN(new_n786_) );
  NAND2_X1 g428 ( .A1(new_n786_), .A2(KEYINPUT27), .ZN(new_n787_) );
  NAND3_X1 g429 ( .A1(new_n787_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n788_) );
  OR2_X1 g430 ( .A1(new_n788_), .A2(G299), .ZN(new_n789_) );
  NAND2_X1 g431 ( .A1(new_n782_), .A2(new_n789_), .ZN(new_n790_) );
  NAND2_X1 g432 ( .A1(new_n788_), .A2(G299), .ZN(new_n791_) );
  XNOR2_X1 g433 ( .A(new_n791_), .B(KEYINPUT28), .ZN(new_n792_) );
  NAND2_X1 g434 ( .A1(new_n790_), .A2(new_n792_), .ZN(new_n793_) );
  NAND2_X1 g435 ( .A1(new_n793_), .A2(new_n760_), .ZN(new_n794_) );
  NAND3_X1 g436 ( .A1(new_n790_), .A2(new_n792_), .A3(KEYINPUT29), .ZN(new_n795_) );
  NAND2_X1 g437 ( .A1(new_n794_), .A2(new_n795_), .ZN(new_n796_) );
  NAND2_X1 g438 ( .A1(new_n767_), .A2(new_n654_), .ZN(new_n797_) );
  NAND2_X1 g439 ( .A1(new_n766_), .A2(new_n670_), .ZN(new_n798_) );
  NAND2_X1 g440 ( .A1(new_n797_), .A2(new_n798_), .ZN(new_n799_) );
  NAND2_X1 g441 ( .A1(G171), .A2(new_n799_), .ZN(new_n800_) );
  NAND2_X1 g442 ( .A1(new_n796_), .A2(new_n800_), .ZN(new_n801_) );
  INV_X1 g443 ( .A(G8), .ZN(new_n802_) );
  NOR2_X1 g444 ( .A1(new_n766_), .A2(new_n802_), .ZN(new_n803_) );
  NAND2_X1 g445 ( .A1(new_n803_), .A2(new_n637_), .ZN(new_n804_) );
  OR2_X1 g446 ( .A1(new_n767_), .A2(G2084), .ZN(new_n805_) );
  NAND3_X1 g447 ( .A1(new_n805_), .A2(new_n804_), .A3(G8), .ZN(new_n806_) );
  OR2_X1 g448 ( .A1(new_n806_), .A2(KEYINPUT30), .ZN(new_n807_) );
  NAND2_X1 g449 ( .A1(new_n806_), .A2(KEYINPUT30), .ZN(new_n808_) );
  NAND3_X1 g450 ( .A1(new_n455_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_) );
  OR2_X1 g451 ( .A1(G171), .A2(new_n799_), .ZN(new_n810_) );
  NAND2_X1 g452 ( .A1(new_n809_), .A2(new_n810_), .ZN(new_n811_) );
  XNOR2_X1 g453 ( .A(new_n811_), .B(KEYINPUT31), .ZN(new_n812_) );
  NAND2_X1 g454 ( .A1(new_n801_), .A2(new_n812_), .ZN(new_n813_) );
  NAND2_X1 g455 ( .A1(new_n813_), .A2(G286), .ZN(new_n814_) );
  INV_X1 g456 ( .A(new_n803_), .ZN(new_n815_) );
  OR2_X1 g457 ( .A1(new_n815_), .A2(G1971), .ZN(new_n816_) );
  NAND2_X1 g458 ( .A1(new_n766_), .A2(new_n584_), .ZN(new_n817_) );
  NAND3_X1 g459 ( .A1(new_n816_), .A2(G303), .A3(new_n817_), .ZN(new_n818_) );
  NAND2_X1 g460 ( .A1(new_n814_), .A2(new_n818_), .ZN(new_n819_) );
  NAND2_X1 g461 ( .A1(new_n819_), .A2(G8), .ZN(new_n820_) );
  NAND2_X1 g462 ( .A1(new_n820_), .A2(KEYINPUT32), .ZN(new_n821_) );
  INV_X1 g463 ( .A(KEYINPUT32), .ZN(new_n822_) );
  NAND3_X1 g464 ( .A1(new_n819_), .A2(G8), .A3(new_n822_), .ZN(new_n823_) );
  NAND2_X1 g465 ( .A1(new_n821_), .A2(new_n823_), .ZN(new_n824_) );
  OR2_X1 g466 ( .A1(new_n805_), .A2(new_n802_), .ZN(new_n825_) );
  NAND3_X1 g467 ( .A1(new_n813_), .A2(new_n804_), .A3(new_n825_), .ZN(new_n826_) );
  NAND2_X1 g468 ( .A1(new_n824_), .A2(new_n826_), .ZN(new_n827_) );
  NAND2_X1 g469 ( .A1(new_n827_), .A2(new_n651_), .ZN(new_n828_) );
  AND2_X1 g470 ( .A1(new_n803_), .A2(new_n646_), .ZN(new_n829_) );
  NAND2_X1 g471 ( .A1(new_n828_), .A2(new_n829_), .ZN(new_n830_) );
  NAND2_X1 g472 ( .A1(new_n830_), .A2(new_n759_), .ZN(new_n831_) );
  NAND3_X1 g473 ( .A1(new_n803_), .A2(KEYINPUT33), .A3(new_n650_), .ZN(new_n832_) );
  AND2_X1 g474 ( .A1(new_n639_), .A2(new_n832_), .ZN(new_n833_) );
  NAND2_X1 g475 ( .A1(new_n831_), .A2(new_n833_), .ZN(new_n834_) );
  NAND3_X1 g476 ( .A1(G166), .A2(G8), .A3(new_n584_), .ZN(new_n835_) );
  NAND2_X1 g477 ( .A1(new_n827_), .A2(new_n835_), .ZN(new_n836_) );
  NAND2_X1 g478 ( .A1(new_n836_), .A2(new_n815_), .ZN(new_n837_) );
  INV_X1 g479 ( .A(KEYINPUT24), .ZN(new_n838_) );
  NOR2_X1 g480 ( .A1(G305), .A2(G1981), .ZN(new_n839_) );
  OR2_X1 g481 ( .A1(new_n839_), .A2(new_n838_), .ZN(new_n840_) );
  NAND2_X1 g482 ( .A1(new_n839_), .A2(new_n838_), .ZN(new_n841_) );
  NAND3_X1 g483 ( .A1(new_n840_), .A2(new_n803_), .A3(new_n841_), .ZN(new_n842_) );
  AND2_X1 g484 ( .A1(new_n837_), .A2(new_n842_), .ZN(new_n843_) );
  NAND2_X1 g485 ( .A1(new_n834_), .A2(new_n843_), .ZN(new_n844_) );
  INV_X1 g486 ( .A(new_n765_), .ZN(new_n845_) );
  NAND2_X1 g487 ( .A1(new_n845_), .A2(new_n762_), .ZN(new_n846_) );
  INV_X1 g488 ( .A(new_n846_), .ZN(new_n847_) );
  NAND3_X1 g489 ( .A1(new_n611_), .A2(new_n612_), .A3(new_n847_), .ZN(new_n848_) );
  OR2_X1 g490 ( .A1(new_n652_), .A2(new_n846_), .ZN(new_n849_) );
  NAND2_X1 g491 ( .A1(new_n623_), .A2(new_n847_), .ZN(new_n850_) );
  AND3_X1 g492 ( .A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_) );
  NAND2_X1 g493 ( .A1(new_n844_), .A2(new_n851_), .ZN(new_n852_) );
  OR2_X1 g494 ( .A1(G290), .A2(G1986), .ZN(new_n853_) );
  NAND2_X1 g495 ( .A1(new_n853_), .A2(new_n627_), .ZN(new_n854_) );
  NAND2_X1 g496 ( .A1(new_n850_), .A2(new_n854_), .ZN(new_n855_) );
  NAND2_X1 g497 ( .A1(new_n855_), .A2(new_n583_), .ZN(new_n856_) );
  XOR2_X1 g498 ( .A(new_n856_), .B(KEYINPUT39), .Z(new_n857_) );
  NAND2_X1 g499 ( .A1(new_n857_), .A2(new_n848_), .ZN(new_n858_) );
  NAND2_X1 g500 ( .A1(new_n858_), .A2(new_n613_), .ZN(new_n859_) );
  NAND2_X1 g501 ( .A1(new_n859_), .A2(new_n847_), .ZN(new_n860_) );
  NAND2_X1 g502 ( .A1(new_n852_), .A2(new_n860_), .ZN(new_n861_) );
  NAND2_X1 g503 ( .A1(new_n861_), .A2(KEYINPUT40), .ZN(new_n862_) );
  INV_X1 g504 ( .A(KEYINPUT40), .ZN(new_n863_) );
  NAND3_X1 g505 ( .A1(new_n852_), .A2(new_n863_), .A3(new_n860_), .ZN(new_n864_) );
  NAND2_X1 g506 ( .A1(new_n862_), .A2(new_n864_), .ZN(G329) );
  INV_X1 g507 ( .A(KEYINPUT49), .ZN(new_n867_) );
  OR2_X1 g508 ( .A1(G229), .A2(G227), .ZN(new_n868_) );
  AND2_X1 g509 ( .A1(new_n868_), .A2(new_n867_), .ZN(new_n869_) );
  NOR2_X1 g510 ( .A1(new_n868_), .A2(new_n867_), .ZN(new_n870_) );
  NAND2_X1 g511 ( .A1(new_n553_), .A2(G319), .ZN(new_n871_) );
  NOR4_X1 g512 ( .A1(G395), .A2(new_n869_), .A3(new_n870_), .A4(new_n871_), .ZN(new_n872_) );
  NAND2_X1 g513 ( .A1(new_n757_), .A2(new_n872_), .ZN(G225) );
  INV_X1 g514 ( .A(G225), .ZN(G308) );
  assign   G231 = 1'b0;
  BUF_X1 g515 ( .A(G452), .Z(G350) );
  BUF_X1 g516 ( .A(G452), .Z(G335) );
  BUF_X1 g517 ( .A(G452), .Z(G409) );
  BUF_X1 g518 ( .A(G1083), .Z(G369) );
  BUF_X1 g519 ( .A(G1083), .Z(G367) );
  BUF_X1 g520 ( .A(G2066), .Z(G411) );
  BUF_X1 g521 ( .A(G2066), .Z(G337) );
  BUF_X1 g522 ( .A(G2066), .Z(G384) );
  BUF_X1 g523 ( .A(G452), .Z(G391) );
  NAND2_X1 g524 ( .A1(new_n523_), .A2(new_n522_), .ZN(G321) );
  NOR2_X1 g525 ( .A1(new_n525_), .A2(new_n526_), .ZN(G280) );
  NOR2_X1 g526 ( .A1(new_n532_), .A2(new_n533_), .ZN(G323) );
  NAND2_X1 g527 ( .A1(new_n749_), .A2(new_n750_), .ZN(G331) );
endmodule


