module add_mul_sub_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, operation_0_, 
        operation_1_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921;

  OR3_X1 U982 ( .A1(n966), .A2(n967), .A3(n968), .ZN(Result_9_) );
  AND3_X1 U983 ( .A1(n969), .A2(n970), .A3(n971), .ZN(n968) );
  INV_X1 U984 ( .A(n972), .ZN(n970) );
  AND2_X1 U985 ( .A1(n973), .A2(n974), .ZN(n972) );
  OR2_X1 U986 ( .A1(n974), .A2(n973), .ZN(n969) );
  AND2_X1 U987 ( .A1(n975), .A2(n976), .ZN(n973) );
  INV_X1 U988 ( .A(n977), .ZN(n976) );
  AND2_X1 U989 ( .A1(n978), .A2(n979), .ZN(n977) );
  OR2_X1 U990 ( .A1(n979), .A2(n978), .ZN(n975) );
  AND2_X1 U991 ( .A1(n980), .A2(n981), .ZN(n967) );
  OR3_X1 U992 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n981) );
  AND2_X1 U993 ( .A1(n985), .A2(n986), .ZN(n984) );
  AND2_X1 U994 ( .A1(n987), .A2(n988), .ZN(n983) );
  AND2_X1 U995 ( .A1(n989), .A2(n990), .ZN(n982) );
  INV_X1 U996 ( .A(n991), .ZN(n990) );
  INV_X1 U997 ( .A(n992), .ZN(n980) );
  AND2_X1 U998 ( .A1(n992), .A2(n993), .ZN(n966) );
  OR3_X1 U999 ( .A1(n994), .A2(n995), .A3(n996), .ZN(n993) );
  AND2_X1 U1000 ( .A1(n997), .A2(n985), .ZN(n996) );
  INV_X1 U1001 ( .A(n986), .ZN(n997) );
  AND2_X1 U1002 ( .A1(n998), .A2(n987), .ZN(n995) );
  INV_X1 U1003 ( .A(n988), .ZN(n998) );
  AND2_X1 U1004 ( .A1(n989), .A2(n991), .ZN(n994) );
  OR2_X1 U1005 ( .A1(n999), .A2(n1000), .ZN(n992) );
  AND2_X1 U1006 ( .A1(a_1_), .A2(n1001), .ZN(n1000) );
  AND2_X1 U1007 ( .A1(b_1_), .A2(n1002), .ZN(n999) );
  OR4_X1 U1008 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(Result_8_) );
  AND2_X1 U1009 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
  INV_X1 U1010 ( .A(n1009), .ZN(n1008) );
  OR2_X1 U1011 ( .A1(n1010), .A2(n1011), .ZN(n1007) );
  AND2_X1 U1012 ( .A1(n1012), .A2(n985), .ZN(n1011) );
  INV_X1 U1013 ( .A(n1013), .ZN(n1012) );
  AND2_X1 U1014 ( .A1(n1014), .A2(n987), .ZN(n1010) );
  INV_X1 U1015 ( .A(n1015), .ZN(n1014) );
  AND2_X1 U1016 ( .A1(n1009), .A2(n1016), .ZN(n1005) );
  OR3_X1 U1017 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
  AND2_X1 U1018 ( .A1(n985), .A2(n1013), .ZN(n1019) );
  AND2_X1 U1019 ( .A1(n987), .A2(n1015), .ZN(n1018) );
  AND2_X1 U1020 ( .A1(n989), .A2(n1020), .ZN(n1017) );
  AND2_X1 U1021 ( .A1(n971), .A2(n1021), .ZN(n1004) );
  OR2_X1 U1022 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
  AND2_X1 U1023 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
  INV_X1 U1024 ( .A(n1026), .ZN(n1022) );
  OR2_X1 U1025 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  OR2_X1 U1026 ( .A1(n1027), .A2(n1028), .ZN(n1024) );
  AND2_X1 U1027 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
  INV_X1 U1028 ( .A(n1031), .ZN(n1029) );
  AND2_X1 U1029 ( .A1(n1032), .A2(n1031), .ZN(n1027) );
  INV_X1 U1030 ( .A(n1030), .ZN(n1032) );
  AND3_X1 U1031 ( .A1(n1033), .A2(n1020), .A3(n989), .ZN(n1003) );
  INV_X1 U1032 ( .A(n1034), .ZN(n1020) );
  AND2_X1 U1033 ( .A1(n1033), .A2(n1009), .ZN(n1034) );
  AND2_X1 U1034 ( .A1(n1035), .A2(n1036), .ZN(n1009) );
  OR2_X1 U1035 ( .A1(n1037), .A2(n1038), .ZN(n1033) );
  AND2_X1 U1036 ( .A1(n1002), .A2(n1001), .ZN(n1038) );
  AND2_X1 U1037 ( .A1(n1039), .A2(n991), .ZN(n1037) );
  OR2_X1 U1038 ( .A1(n1040), .A2(n1041), .ZN(n991) );
  AND2_X1 U1039 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
  AND2_X1 U1040 ( .A1(n1044), .A2(n1045), .ZN(n1040) );
  OR2_X1 U1041 ( .A1(n1046), .A2(n1047), .ZN(Result_7_) );
  AND3_X1 U1042 ( .A1(n1048), .A2(n1049), .A3(n971), .ZN(n1046) );
  OR2_X1 U1043 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
  INV_X1 U1044 ( .A(n1052), .ZN(n1051) );
  OR2_X1 U1045 ( .A1(n1053), .A2(n1052), .ZN(n1048) );
  OR2_X1 U1046 ( .A1(n1054), .A2(n1047), .ZN(Result_6_) );
  AND3_X1 U1047 ( .A1(n1055), .A2(n1056), .A3(n971), .ZN(n1054) );
  INV_X1 U1048 ( .A(n1057), .ZN(n1056) );
  OR2_X1 U1049 ( .A1(n1058), .A2(n1059), .ZN(n1055) );
  AND2_X1 U1050 ( .A1(n1053), .A2(n1052), .ZN(n1058) );
  OR2_X1 U1051 ( .A1(n1060), .A2(n1047), .ZN(Result_5_) );
  AND2_X1 U1052 ( .A1(n971), .A2(n1061), .ZN(n1060) );
  OR2_X1 U1053 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
  INV_X1 U1054 ( .A(n1064), .ZN(n1063) );
  OR2_X1 U1055 ( .A1(n1065), .A2(n1057), .ZN(n1064) );
  AND2_X1 U1056 ( .A1(n1057), .A2(n1065), .ZN(n1062) );
  OR2_X1 U1057 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
  AND2_X1 U1058 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
  OR2_X1 U1059 ( .A1(n1070), .A2(n1047), .ZN(Result_4_) );
  AND3_X1 U1060 ( .A1(n1071), .A2(n1072), .A3(n971), .ZN(n1070) );
  OR2_X1 U1061 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
  OR3_X1 U1062 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1071) );
  INV_X1 U1063 ( .A(n1078), .ZN(n1076) );
  OR2_X1 U1064 ( .A1(n1074), .A2(n1079), .ZN(n1078) );
  AND2_X1 U1065 ( .A1(n1079), .A2(n1074), .ZN(n1075) );
  OR2_X1 U1066 ( .A1(n1080), .A2(n1047), .ZN(Result_3_) );
  AND3_X1 U1067 ( .A1(n1081), .A2(n1082), .A3(n971), .ZN(n1080) );
  OR3_X1 U1068 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
  INV_X1 U1069 ( .A(n1086), .ZN(n1085) );
  AND2_X1 U1070 ( .A1(n1087), .A2(n1088), .ZN(n1084) );
  INV_X1 U1071 ( .A(n1089), .ZN(n1083) );
  OR2_X1 U1072 ( .A1(n1088), .A2(n1087), .ZN(n1089) );
  OR2_X1 U1073 ( .A1(n1088), .A2(n1086), .ZN(n1081) );
  OR2_X1 U1074 ( .A1(n1090), .A2(n1047), .ZN(Result_2_) );
  AND3_X1 U1075 ( .A1(n1091), .A2(n1092), .A3(n971), .ZN(n1090) );
  OR3_X1 U1076 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
  INV_X1 U1077 ( .A(n1096), .ZN(n1095) );
  INV_X1 U1078 ( .A(n1097), .ZN(n1094) );
  OR2_X1 U1079 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
  AND2_X1 U1080 ( .A1(n1099), .A2(n1098), .ZN(n1093) );
  OR2_X1 U1081 ( .A1(n1098), .A2(n1096), .ZN(n1091) );
  OR2_X1 U1082 ( .A1(n1100), .A2(n1047), .ZN(Result_1_) );
  AND3_X1 U1083 ( .A1(n1101), .A2(n1102), .A3(n971), .ZN(n1100) );
  OR3_X1 U1084 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
  AND2_X1 U1085 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
  AND2_X1 U1086 ( .A1(n1108), .A2(n1109), .ZN(n1103) );
  OR2_X1 U1087 ( .A1(n1110), .A2(n1108), .ZN(n1101) );
  OR2_X1 U1088 ( .A1(n1111), .A2(n1112), .ZN(Result_15_) );
  AND2_X1 U1089 ( .A1(n971), .A2(n1113), .ZN(n1112) );
  AND2_X1 U1090 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
  OR3_X1 U1091 ( .A1(n985), .A2(n987), .A3(n989), .ZN(n1115) );
  OR2_X1 U1092 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
  OR3_X1 U1093 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(Result_14_) );
  AND2_X1 U1094 ( .A1(n971), .A2(n1121), .ZN(n1120) );
  OR4_X1 U1095 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1121) );
  AND2_X1 U1096 ( .A1(n1116), .A2(b_6_), .ZN(n1125) );
  AND2_X1 U1097 ( .A1(n1126), .A2(a_7_), .ZN(n1124) );
  AND2_X1 U1098 ( .A1(n1117), .A2(a_6_), .ZN(n1123) );
  AND2_X1 U1099 ( .A1(n1127), .A2(b_7_), .ZN(n1122) );
  AND2_X1 U1100 ( .A1(n1128), .A2(n1129), .ZN(n1119) );
  OR3_X1 U1101 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1129) );
  AND2_X1 U1102 ( .A1(n985), .A2(n1117), .ZN(n1132) );
  AND2_X1 U1103 ( .A1(n987), .A2(n1116), .ZN(n1131) );
  AND2_X1 U1104 ( .A1(n989), .A2(n1113), .ZN(n1130) );
  INV_X1 U1105 ( .A(n1133), .ZN(n1128) );
  AND2_X1 U1106 ( .A1(n1134), .A2(n1133), .ZN(n1118) );
  OR2_X1 U1107 ( .A1(n1126), .A2(n1127), .ZN(n1133) );
  OR3_X1 U1108 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
  AND2_X1 U1109 ( .A1(n985), .A2(n1138), .ZN(n1137) );
  INV_X1 U1110 ( .A(n1117), .ZN(n1138) );
  AND2_X1 U1111 ( .A1(n987), .A2(n1139), .ZN(n1136) );
  AND2_X1 U1112 ( .A1(n989), .A2(n1140), .ZN(n1135) );
  OR3_X1 U1113 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(Result_13_) );
  AND2_X1 U1114 ( .A1(n971), .A2(n1144), .ZN(n1143) );
  OR2_X1 U1115 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
  AND2_X1 U1116 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
  INV_X1 U1117 ( .A(n1149), .ZN(n1145) );
  OR2_X1 U1118 ( .A1(n1148), .A2(n1147), .ZN(n1149) );
  OR2_X1 U1119 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
  AND2_X1 U1120 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
  INV_X1 U1121 ( .A(n1154), .ZN(n1150) );
  OR2_X1 U1122 ( .A1(n1153), .A2(n1152), .ZN(n1154) );
  INV_X1 U1123 ( .A(n1155), .ZN(n1152) );
  AND2_X1 U1124 ( .A1(n1156), .A2(n1157), .ZN(n1142) );
  OR3_X1 U1125 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1157) );
  AND2_X1 U1126 ( .A1(n985), .A2(n1161), .ZN(n1160) );
  AND2_X1 U1127 ( .A1(n987), .A2(n1162), .ZN(n1159) );
  AND2_X1 U1128 ( .A1(n989), .A2(n1163), .ZN(n1158) );
  INV_X1 U1129 ( .A(n1164), .ZN(n1156) );
  AND2_X1 U1130 ( .A1(n1164), .A2(n1165), .ZN(n1141) );
  OR3_X1 U1131 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
  AND2_X1 U1132 ( .A1(n985), .A2(n1169), .ZN(n1168) );
  INV_X1 U1133 ( .A(n1161), .ZN(n1169) );
  AND2_X1 U1134 ( .A1(n987), .A2(n1170), .ZN(n1167) );
  AND2_X1 U1135 ( .A1(n989), .A2(n1171), .ZN(n1166) );
  OR2_X1 U1136 ( .A1(n1172), .A2(n1173), .ZN(n1164) );
  AND2_X1 U1137 ( .A1(a_5_), .A2(n1174), .ZN(n1173) );
  AND2_X1 U1138 ( .A1(b_5_), .A2(n1175), .ZN(n1172) );
  OR3_X1 U1139 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(Result_12_) );
  AND2_X1 U1140 ( .A1(n971), .A2(n1179), .ZN(n1178) );
  OR2_X1 U1141 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
  AND2_X1 U1142 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
  INV_X1 U1143 ( .A(n1184), .ZN(n1180) );
  OR2_X1 U1144 ( .A1(n1183), .A2(n1182), .ZN(n1184) );
  OR2_X1 U1145 ( .A1(n1185), .A2(n1186), .ZN(n1182) );
  AND2_X1 U1146 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
  INV_X1 U1147 ( .A(n1189), .ZN(n1187) );
  AND2_X1 U1148 ( .A1(n1190), .A2(n1189), .ZN(n1185) );
  INV_X1 U1149 ( .A(n1188), .ZN(n1190) );
  AND2_X1 U1150 ( .A1(n1191), .A2(n1192), .ZN(n1177) );
  OR3_X1 U1151 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1192) );
  AND2_X1 U1152 ( .A1(n985), .A2(n1196), .ZN(n1195) );
  AND2_X1 U1153 ( .A1(n987), .A2(n1197), .ZN(n1194) );
  AND2_X1 U1154 ( .A1(n1198), .A2(n989), .ZN(n1193) );
  INV_X1 U1155 ( .A(n1199), .ZN(n1198) );
  INV_X1 U1156 ( .A(n1200), .ZN(n1191) );
  AND2_X1 U1157 ( .A1(n1200), .A2(n1201), .ZN(n1176) );
  OR3_X1 U1158 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1201) );
  AND2_X1 U1159 ( .A1(n985), .A2(n1205), .ZN(n1204) );
  INV_X1 U1160 ( .A(n1196), .ZN(n1205) );
  AND2_X1 U1161 ( .A1(n987), .A2(n1206), .ZN(n1203) );
  INV_X1 U1162 ( .A(n1197), .ZN(n1206) );
  AND2_X1 U1163 ( .A1(n989), .A2(n1199), .ZN(n1202) );
  OR2_X1 U1164 ( .A1(n1207), .A2(n1208), .ZN(n1200) );
  AND2_X1 U1165 ( .A1(a_4_), .A2(n1209), .ZN(n1208) );
  AND2_X1 U1166 ( .A1(b_4_), .A2(n1210), .ZN(n1207) );
  OR3_X1 U1167 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(Result_11_) );
  AND2_X1 U1168 ( .A1(n971), .A2(n1214), .ZN(n1213) );
  OR2_X1 U1169 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
  AND2_X1 U1170 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
  INV_X1 U1171 ( .A(n1219), .ZN(n1215) );
  OR2_X1 U1172 ( .A1(n1218), .A2(n1217), .ZN(n1219) );
  OR2_X1 U1173 ( .A1(n1220), .A2(n1221), .ZN(n1217) );
  AND2_X1 U1174 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
  INV_X1 U1175 ( .A(n1224), .ZN(n1222) );
  AND2_X1 U1176 ( .A1(n1225), .A2(n1224), .ZN(n1220) );
  INV_X1 U1177 ( .A(n1223), .ZN(n1225) );
  AND2_X1 U1178 ( .A1(n1226), .A2(n1227), .ZN(n1212) );
  OR3_X1 U1179 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1227) );
  AND2_X1 U1180 ( .A1(n985), .A2(n1231), .ZN(n1230) );
  AND2_X1 U1181 ( .A1(n987), .A2(n1232), .ZN(n1229) );
  AND2_X1 U1182 ( .A1(n1233), .A2(n989), .ZN(n1228) );
  INV_X1 U1183 ( .A(n1234), .ZN(n1233) );
  INV_X1 U1184 ( .A(n1235), .ZN(n1226) );
  AND2_X1 U1185 ( .A1(n1235), .A2(n1236), .ZN(n1211) );
  OR3_X1 U1186 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1236) );
  AND2_X1 U1187 ( .A1(n985), .A2(n1240), .ZN(n1239) );
  INV_X1 U1188 ( .A(n1231), .ZN(n1240) );
  AND2_X1 U1189 ( .A1(n987), .A2(n1241), .ZN(n1238) );
  INV_X1 U1190 ( .A(n1232), .ZN(n1241) );
  AND2_X1 U1191 ( .A1(n989), .A2(n1234), .ZN(n1237) );
  OR2_X1 U1192 ( .A1(n1242), .A2(n1243), .ZN(n1235) );
  AND2_X1 U1193 ( .A1(a_3_), .A2(n1244), .ZN(n1243) );
  AND2_X1 U1194 ( .A1(b_3_), .A2(n1245), .ZN(n1242) );
  OR3_X1 U1195 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(Result_10_) );
  AND2_X1 U1196 ( .A1(n971), .A2(n1249), .ZN(n1248) );
  OR2_X1 U1197 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
  AND2_X1 U1198 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
  INV_X1 U1199 ( .A(n1254), .ZN(n1250) );
  OR2_X1 U1200 ( .A1(n1253), .A2(n1252), .ZN(n1254) );
  OR2_X1 U1201 ( .A1(n1255), .A2(n1256), .ZN(n1252) );
  AND2_X1 U1202 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
  INV_X1 U1203 ( .A(n1259), .ZN(n1257) );
  AND2_X1 U1204 ( .A1(n1260), .A2(n1259), .ZN(n1255) );
  INV_X1 U1205 ( .A(n1258), .ZN(n1260) );
  AND2_X1 U1206 ( .A1(n1261), .A2(n1262), .ZN(n1247) );
  OR3_X1 U1207 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1262) );
  AND2_X1 U1208 ( .A1(n985), .A2(n1266), .ZN(n1265) );
  AND2_X1 U1209 ( .A1(n987), .A2(n1267), .ZN(n1264) );
  AND2_X1 U1210 ( .A1(n1268), .A2(n989), .ZN(n1263) );
  INV_X1 U1211 ( .A(n1044), .ZN(n1268) );
  INV_X1 U1212 ( .A(n1269), .ZN(n1261) );
  AND2_X1 U1213 ( .A1(n1269), .A2(n1270), .ZN(n1246) );
  OR3_X1 U1214 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1270) );
  AND2_X1 U1215 ( .A1(n985), .A2(n1274), .ZN(n1273) );
  INV_X1 U1216 ( .A(n1266), .ZN(n1274) );
  AND2_X1 U1217 ( .A1(n987), .A2(n1275), .ZN(n1272) );
  INV_X1 U1218 ( .A(n1267), .ZN(n1275) );
  AND2_X1 U1219 ( .A1(n989), .A2(n1044), .ZN(n1271) );
  OR2_X1 U1220 ( .A1(n1276), .A2(n1277), .ZN(n1044) );
  AND2_X1 U1221 ( .A1(n1245), .A2(n1244), .ZN(n1277) );
  AND2_X1 U1222 ( .A1(n1234), .A2(n1278), .ZN(n1276) );
  OR2_X1 U1223 ( .A1(n1279), .A2(n1280), .ZN(n1234) );
  AND2_X1 U1224 ( .A1(n1210), .A2(n1209), .ZN(n1280) );
  AND2_X1 U1225 ( .A1(n1199), .A2(n1281), .ZN(n1279) );
  OR2_X1 U1226 ( .A1(n1282), .A2(n1283), .ZN(n1199) );
  AND2_X1 U1227 ( .A1(n1175), .A2(n1174), .ZN(n1283) );
  AND2_X1 U1228 ( .A1(n1171), .A2(n1284), .ZN(n1282) );
  INV_X1 U1229 ( .A(n1163), .ZN(n1171) );
  OR2_X1 U1230 ( .A1(n1285), .A2(n1286), .ZN(n1163) );
  AND2_X1 U1231 ( .A1(n1113), .A2(n1287), .ZN(n1285) );
  OR2_X1 U1232 ( .A1(a_6_), .A2(b_6_), .ZN(n1287) );
  AND2_X1 U1233 ( .A1(n1288), .A2(n1289), .ZN(n989) );
  OR2_X1 U1234 ( .A1(n1290), .A2(n1291), .ZN(n1269) );
  AND2_X1 U1235 ( .A1(a_2_), .A2(n1043), .ZN(n1291) );
  AND2_X1 U1236 ( .A1(b_2_), .A2(n1042), .ZN(n1290) );
  OR2_X1 U1237 ( .A1(n1292), .A2(n1047), .ZN(Result_0_) );
  OR2_X1 U1238 ( .A1(n1293), .A2(n1294), .ZN(n1047) );
  AND2_X1 U1239 ( .A1(n985), .A2(n1295), .ZN(n1294) );
  OR2_X1 U1240 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
  AND2_X1 U1241 ( .A1(n1013), .A2(n1036), .ZN(n1296) );
  INV_X1 U1242 ( .A(n1298), .ZN(n1036) );
  OR2_X1 U1243 ( .A1(n1299), .A2(n1300), .ZN(n1013) );
  AND2_X1 U1244 ( .A1(n986), .A2(n1002), .ZN(n1300) );
  AND2_X1 U1245 ( .A1(b_1_), .A2(n1301), .ZN(n1299) );
  OR2_X1 U1246 ( .A1(n1002), .A2(n986), .ZN(n1301) );
  OR2_X1 U1247 ( .A1(n1302), .A2(n1303), .ZN(n986) );
  AND2_X1 U1248 ( .A1(n1266), .A2(n1042), .ZN(n1303) );
  AND2_X1 U1249 ( .A1(b_2_), .A2(n1304), .ZN(n1302) );
  OR2_X1 U1250 ( .A1(n1042), .A2(n1266), .ZN(n1304) );
  OR2_X1 U1251 ( .A1(n1305), .A2(n1306), .ZN(n1266) );
  AND2_X1 U1252 ( .A1(n1231), .A2(n1245), .ZN(n1306) );
  AND2_X1 U1253 ( .A1(b_3_), .A2(n1307), .ZN(n1305) );
  OR2_X1 U1254 ( .A1(n1245), .A2(n1231), .ZN(n1307) );
  OR2_X1 U1255 ( .A1(n1308), .A2(n1309), .ZN(n1231) );
  AND2_X1 U1256 ( .A1(n1196), .A2(n1210), .ZN(n1309) );
  AND2_X1 U1257 ( .A1(b_4_), .A2(n1310), .ZN(n1308) );
  OR2_X1 U1258 ( .A1(n1210), .A2(n1196), .ZN(n1310) );
  OR2_X1 U1259 ( .A1(n1311), .A2(n1312), .ZN(n1196) );
  AND2_X1 U1260 ( .A1(n1161), .A2(n1175), .ZN(n1312) );
  AND2_X1 U1261 ( .A1(b_5_), .A2(n1313), .ZN(n1311) );
  OR2_X1 U1262 ( .A1(n1175), .A2(n1161), .ZN(n1313) );
  OR2_X1 U1263 ( .A1(n1314), .A2(n1126), .ZN(n1161) );
  AND2_X1 U1264 ( .A1(n1117), .A2(n1315), .ZN(n1314) );
  AND2_X1 U1265 ( .A1(n1316), .A2(b_7_), .ZN(n1117) );
  AND2_X1 U1266 ( .A1(n1289), .A2(operation_1_), .ZN(n985) );
  INV_X1 U1267 ( .A(operation_0_), .ZN(n1289) );
  AND3_X1 U1268 ( .A1(n1317), .A2(n1035), .A3(n987), .ZN(n1293) );
  AND2_X1 U1269 ( .A1(n1288), .A2(operation_0_), .ZN(n987) );
  INV_X1 U1270 ( .A(operation_1_), .ZN(n1288) );
  INV_X1 U1271 ( .A(n1297), .ZN(n1035) );
  AND2_X1 U1272 ( .A1(n1318), .A2(b_0_), .ZN(n1297) );
  OR2_X1 U1273 ( .A1(n1298), .A2(n1015), .ZN(n1317) );
  OR2_X1 U1274 ( .A1(n1319), .A2(n1320), .ZN(n1015) );
  AND2_X1 U1275 ( .A1(a_1_), .A2(n988), .ZN(n1320) );
  AND2_X1 U1276 ( .A1(n1321), .A2(n1001), .ZN(n1319) );
  OR2_X1 U1277 ( .A1(a_1_), .A2(n988), .ZN(n1321) );
  OR2_X1 U1278 ( .A1(n1322), .A2(n1323), .ZN(n988) );
  AND2_X1 U1279 ( .A1(a_2_), .A2(n1267), .ZN(n1323) );
  AND2_X1 U1280 ( .A1(n1324), .A2(n1043), .ZN(n1322) );
  OR2_X1 U1281 ( .A1(a_2_), .A2(n1267), .ZN(n1324) );
  OR2_X1 U1282 ( .A1(n1325), .A2(n1326), .ZN(n1267) );
  AND2_X1 U1283 ( .A1(a_3_), .A2(n1232), .ZN(n1326) );
  AND2_X1 U1284 ( .A1(n1327), .A2(n1244), .ZN(n1325) );
  OR2_X1 U1285 ( .A1(a_3_), .A2(n1232), .ZN(n1327) );
  OR2_X1 U1286 ( .A1(n1328), .A2(n1329), .ZN(n1232) );
  AND2_X1 U1287 ( .A1(a_4_), .A2(n1197), .ZN(n1329) );
  AND2_X1 U1288 ( .A1(n1330), .A2(n1209), .ZN(n1328) );
  OR2_X1 U1289 ( .A1(a_4_), .A2(n1197), .ZN(n1330) );
  OR2_X1 U1290 ( .A1(n1331), .A2(n1332), .ZN(n1197) );
  AND2_X1 U1291 ( .A1(a_5_), .A2(n1162), .ZN(n1332) );
  AND2_X1 U1292 ( .A1(n1333), .A2(n1174), .ZN(n1331) );
  OR2_X1 U1293 ( .A1(a_5_), .A2(n1162), .ZN(n1333) );
  INV_X1 U1294 ( .A(n1170), .ZN(n1162) );
  AND2_X1 U1295 ( .A1(n1315), .A2(n1334), .ZN(n1170) );
  OR2_X1 U1296 ( .A1(n1139), .A2(n1126), .ZN(n1334) );
  AND2_X1 U1297 ( .A1(n1335), .A2(b_6_), .ZN(n1126) );
  INV_X1 U1298 ( .A(n1116), .ZN(n1139) );
  AND2_X1 U1299 ( .A1(n1336), .A2(a_7_), .ZN(n1116) );
  INV_X1 U1300 ( .A(n1127), .ZN(n1315) );
  AND2_X1 U1301 ( .A1(n1337), .A2(a_6_), .ZN(n1127) );
  AND2_X1 U1302 ( .A1(n1338), .A2(a_0_), .ZN(n1298) );
  AND2_X1 U1303 ( .A1(n971), .A2(n1339), .ZN(n1292) );
  OR3_X1 U1304 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1339) );
  AND2_X1 U1305 ( .A1(n1343), .A2(a_0_), .ZN(n1342) );
  INV_X1 U1306 ( .A(n1344), .ZN(n1343) );
  AND2_X1 U1307 ( .A1(n1105), .A2(n1106), .ZN(n1341) );
  INV_X1 U1308 ( .A(n1110), .ZN(n1105) );
  OR2_X1 U1309 ( .A1(n1345), .A2(n1098), .ZN(n1110) );
  OR2_X1 U1310 ( .A1(n1346), .A2(n1109), .ZN(n1098) );
  AND2_X1 U1311 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
  AND2_X1 U1312 ( .A1(n1349), .A2(n1096), .ZN(n1345) );
  OR2_X1 U1313 ( .A1(n1350), .A2(n1088), .ZN(n1096) );
  OR2_X1 U1314 ( .A1(n1099), .A2(n1351), .ZN(n1088) );
  AND3_X1 U1315 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1351) );
  INV_X1 U1316 ( .A(n1349), .ZN(n1099) );
  AND2_X1 U1317 ( .A1(n1086), .A2(n1355), .ZN(n1350) );
  OR2_X1 U1318 ( .A1(n1356), .A2(n1074), .ZN(n1086) );
  OR2_X1 U1319 ( .A1(n1357), .A2(n1087), .ZN(n1074) );
  INV_X1 U1320 ( .A(n1355), .ZN(n1087) );
  OR2_X1 U1321 ( .A1(n1358), .A2(n1359), .ZN(n1355) );
  AND2_X1 U1322 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
  OR2_X1 U1323 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
  AND2_X1 U1324 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
  AND2_X1 U1325 ( .A1(n1364), .A2(n1365), .ZN(n1360) );
  OR2_X1 U1326 ( .A1(n1363), .A2(n1362), .ZN(n1365) );
  AND2_X1 U1327 ( .A1(n1366), .A2(n1367), .ZN(n1358) );
  INV_X1 U1328 ( .A(n1368), .ZN(n1367) );
  AND2_X1 U1329 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
  OR2_X1 U1330 ( .A1(n1370), .A2(n1369), .ZN(n1366) );
  OR2_X1 U1331 ( .A1(n1371), .A2(n1372), .ZN(n1369) );
  AND2_X1 U1332 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
  INV_X1 U1333 ( .A(n1375), .ZN(n1373) );
  AND2_X1 U1334 ( .A1(n1376), .A2(n1375), .ZN(n1371) );
  AND2_X1 U1335 ( .A1(n1073), .A2(n1377), .ZN(n1356) );
  INV_X1 U1336 ( .A(n1077), .ZN(n1073) );
  OR2_X1 U1337 ( .A1(n1378), .A2(n1066), .ZN(n1077) );
  AND3_X1 U1338 ( .A1(n1379), .A2(n1380), .A3(n1381), .ZN(n1066) );
  AND2_X1 U1339 ( .A1(n1057), .A2(n1381), .ZN(n1378) );
  INV_X1 U1340 ( .A(n1068), .ZN(n1381) );
  OR2_X1 U1341 ( .A1(n1079), .A2(n1382), .ZN(n1068) );
  AND3_X1 U1342 ( .A1(n1383), .A2(n1384), .A3(n1385), .ZN(n1382) );
  INV_X1 U1343 ( .A(n1377), .ZN(n1079) );
  OR2_X1 U1344 ( .A1(n1386), .A2(n1385), .ZN(n1377) );
  OR2_X1 U1345 ( .A1(n1387), .A2(n1388), .ZN(n1385) );
  AND2_X1 U1346 ( .A1(n1389), .A2(n1390), .ZN(n1388) );
  AND2_X1 U1347 ( .A1(n1391), .A2(n1392), .ZN(n1387) );
  OR2_X1 U1348 ( .A1(n1390), .A2(n1389), .ZN(n1391) );
  INV_X1 U1349 ( .A(n1393), .ZN(n1390) );
  AND2_X1 U1350 ( .A1(n1383), .A2(n1384), .ZN(n1386) );
  OR2_X1 U1351 ( .A1(n1394), .A2(n1395), .ZN(n1384) );
  INV_X1 U1352 ( .A(n1364), .ZN(n1394) );
  OR2_X1 U1353 ( .A1(n1396), .A2(n1364), .ZN(n1383) );
  AND2_X1 U1354 ( .A1(n1397), .A2(n1398), .ZN(n1364) );
  INV_X1 U1355 ( .A(n1399), .ZN(n1398) );
  AND2_X1 U1356 ( .A1(n1400), .A2(n1401), .ZN(n1399) );
  OR2_X1 U1357 ( .A1(n1401), .A2(n1400), .ZN(n1397) );
  OR2_X1 U1358 ( .A1(n1402), .A2(n1403), .ZN(n1400) );
  AND2_X1 U1359 ( .A1(n1404), .A2(n1405), .ZN(n1403) );
  INV_X1 U1360 ( .A(n1406), .ZN(n1404) );
  AND2_X1 U1361 ( .A1(n1407), .A2(n1406), .ZN(n1402) );
  INV_X1 U1362 ( .A(n1395), .ZN(n1396) );
  AND2_X1 U1363 ( .A1(n1408), .A2(n1409), .ZN(n1395) );
  INV_X1 U1364 ( .A(n1410), .ZN(n1409) );
  AND2_X1 U1365 ( .A1(n1411), .A2(n1363), .ZN(n1410) );
  OR2_X1 U1366 ( .A1(n1363), .A2(n1411), .ZN(n1408) );
  INV_X1 U1367 ( .A(n1362), .ZN(n1411) );
  OR2_X1 U1368 ( .A1(n1209), .A2(n1318), .ZN(n1362) );
  OR2_X1 U1369 ( .A1(n1412), .A2(n1413), .ZN(n1363) );
  AND2_X1 U1370 ( .A1(n1414), .A2(n1415), .ZN(n1413) );
  AND2_X1 U1371 ( .A1(n1416), .A2(n1417), .ZN(n1412) );
  OR2_X1 U1372 ( .A1(n1415), .A2(n1414), .ZN(n1416) );
  INV_X1 U1373 ( .A(n1418), .ZN(n1415) );
  AND3_X1 U1374 ( .A1(n1053), .A2(n1052), .A3(n1059), .ZN(n1057) );
  AND2_X1 U1375 ( .A1(n1069), .A2(n1419), .ZN(n1059) );
  OR2_X1 U1376 ( .A1(n1380), .A2(n1379), .ZN(n1419) );
  INV_X1 U1377 ( .A(n1420), .ZN(n1379) );
  OR2_X1 U1378 ( .A1(n1421), .A2(n1420), .ZN(n1069) );
  OR2_X1 U1379 ( .A1(n1422), .A2(n1423), .ZN(n1420) );
  AND2_X1 U1380 ( .A1(n1424), .A2(n1425), .ZN(n1423) );
  AND2_X1 U1381 ( .A1(n1426), .A2(n1427), .ZN(n1422) );
  OR2_X1 U1382 ( .A1(n1425), .A2(n1424), .ZN(n1427) );
  INV_X1 U1383 ( .A(n1428), .ZN(n1424) );
  INV_X1 U1384 ( .A(n1380), .ZN(n1421) );
  AND2_X1 U1385 ( .A1(n1429), .A2(n1430), .ZN(n1380) );
  OR2_X1 U1386 ( .A1(n1431), .A2(n1389), .ZN(n1430) );
  INV_X1 U1387 ( .A(n1432), .ZN(n1429) );
  AND2_X1 U1388 ( .A1(n1389), .A2(n1431), .ZN(n1432) );
  AND2_X1 U1389 ( .A1(n1433), .A2(n1434), .ZN(n1431) );
  INV_X1 U1390 ( .A(n1435), .ZN(n1434) );
  AND2_X1 U1391 ( .A1(n1393), .A2(n1392), .ZN(n1435) );
  OR2_X1 U1392 ( .A1(n1392), .A2(n1393), .ZN(n1433) );
  AND2_X1 U1393 ( .A1(b_5_), .A2(a_0_), .ZN(n1393) );
  OR2_X1 U1394 ( .A1(n1436), .A2(n1437), .ZN(n1392) );
  AND2_X1 U1395 ( .A1(n1438), .A2(n1439), .ZN(n1437) );
  AND2_X1 U1396 ( .A1(n1440), .A2(n1441), .ZN(n1436) );
  OR2_X1 U1397 ( .A1(n1439), .A2(n1438), .ZN(n1441) );
  INV_X1 U1398 ( .A(n1442), .ZN(n1438) );
  OR2_X1 U1399 ( .A1(n1443), .A2(n1444), .ZN(n1389) );
  INV_X1 U1400 ( .A(n1445), .ZN(n1444) );
  OR2_X1 U1401 ( .A1(n1446), .A2(n1414), .ZN(n1445) );
  AND2_X1 U1402 ( .A1(n1414), .A2(n1446), .ZN(n1443) );
  AND2_X1 U1403 ( .A1(n1447), .A2(n1448), .ZN(n1446) );
  INV_X1 U1404 ( .A(n1449), .ZN(n1448) );
  AND2_X1 U1405 ( .A1(n1418), .A2(n1417), .ZN(n1449) );
  OR2_X1 U1406 ( .A1(n1417), .A2(n1418), .ZN(n1447) );
  AND2_X1 U1407 ( .A1(b_4_), .A2(a_1_), .ZN(n1418) );
  OR2_X1 U1408 ( .A1(n1450), .A2(n1451), .ZN(n1417) );
  AND2_X1 U1409 ( .A1(n1452), .A2(n1453), .ZN(n1451) );
  AND2_X1 U1410 ( .A1(n1454), .A2(n1455), .ZN(n1450) );
  OR2_X1 U1411 ( .A1(n1453), .A2(n1452), .ZN(n1455) );
  INV_X1 U1412 ( .A(n1456), .ZN(n1452) );
  OR2_X1 U1413 ( .A1(n1457), .A2(n1458), .ZN(n1414) );
  INV_X1 U1414 ( .A(n1459), .ZN(n1458) );
  OR2_X1 U1415 ( .A1(n1460), .A2(n1461), .ZN(n1459) );
  AND2_X1 U1416 ( .A1(n1461), .A2(n1460), .ZN(n1457) );
  AND2_X1 U1417 ( .A1(n1462), .A2(n1463), .ZN(n1460) );
  OR2_X1 U1418 ( .A1(n1464), .A2(n1465), .ZN(n1463) );
  INV_X1 U1419 ( .A(n1466), .ZN(n1462) );
  AND2_X1 U1420 ( .A1(n1465), .A2(n1464), .ZN(n1466) );
  AND2_X1 U1421 ( .A1(n1467), .A2(n1468), .ZN(n1052) );
  OR2_X1 U1422 ( .A1(n1469), .A2(n1426), .ZN(n1468) );
  INV_X1 U1423 ( .A(n1470), .ZN(n1467) );
  AND2_X1 U1424 ( .A1(n1426), .A2(n1469), .ZN(n1470) );
  AND2_X1 U1425 ( .A1(n1471), .A2(n1472), .ZN(n1469) );
  INV_X1 U1426 ( .A(n1473), .ZN(n1472) );
  AND2_X1 U1427 ( .A1(n1428), .A2(n1425), .ZN(n1473) );
  OR2_X1 U1428 ( .A1(n1425), .A2(n1428), .ZN(n1471) );
  AND2_X1 U1429 ( .A1(b_6_), .A2(a_0_), .ZN(n1428) );
  OR2_X1 U1430 ( .A1(n1474), .A2(n1475), .ZN(n1425) );
  AND2_X1 U1431 ( .A1(n1476), .A2(n1477), .ZN(n1475) );
  AND2_X1 U1432 ( .A1(n1478), .A2(n1479), .ZN(n1474) );
  OR2_X1 U1433 ( .A1(n1477), .A2(n1476), .ZN(n1479) );
  OR2_X1 U1434 ( .A1(n1480), .A2(n1481), .ZN(n1426) );
  INV_X1 U1435 ( .A(n1482), .ZN(n1481) );
  OR2_X1 U1436 ( .A1(n1483), .A2(n1440), .ZN(n1482) );
  AND2_X1 U1437 ( .A1(n1440), .A2(n1483), .ZN(n1480) );
  AND2_X1 U1438 ( .A1(n1484), .A2(n1485), .ZN(n1483) );
  INV_X1 U1439 ( .A(n1486), .ZN(n1485) );
  AND2_X1 U1440 ( .A1(n1442), .A2(n1439), .ZN(n1486) );
  OR2_X1 U1441 ( .A1(n1439), .A2(n1442), .ZN(n1484) );
  AND2_X1 U1442 ( .A1(b_5_), .A2(a_1_), .ZN(n1442) );
  OR2_X1 U1443 ( .A1(n1487), .A2(n1488), .ZN(n1439) );
  AND2_X1 U1444 ( .A1(n1489), .A2(n1490), .ZN(n1488) );
  AND2_X1 U1445 ( .A1(n1491), .A2(n1492), .ZN(n1487) );
  OR2_X1 U1446 ( .A1(n1490), .A2(n1489), .ZN(n1492) );
  OR2_X1 U1447 ( .A1(n1493), .A2(n1494), .ZN(n1440) );
  INV_X1 U1448 ( .A(n1495), .ZN(n1494) );
  OR2_X1 U1449 ( .A1(n1496), .A2(n1454), .ZN(n1495) );
  AND2_X1 U1450 ( .A1(n1454), .A2(n1496), .ZN(n1493) );
  AND2_X1 U1451 ( .A1(n1497), .A2(n1498), .ZN(n1496) );
  INV_X1 U1452 ( .A(n1499), .ZN(n1498) );
  AND2_X1 U1453 ( .A1(n1456), .A2(n1453), .ZN(n1499) );
  OR2_X1 U1454 ( .A1(n1453), .A2(n1456), .ZN(n1497) );
  AND2_X1 U1455 ( .A1(b_4_), .A2(a_2_), .ZN(n1456) );
  OR2_X1 U1456 ( .A1(n1500), .A2(n1501), .ZN(n1453) );
  AND2_X1 U1457 ( .A1(n1502), .A2(n1503), .ZN(n1501) );
  AND2_X1 U1458 ( .A1(n1504), .A2(n1505), .ZN(n1500) );
  OR2_X1 U1459 ( .A1(n1503), .A2(n1502), .ZN(n1505) );
  OR2_X1 U1460 ( .A1(n1506), .A2(n1507), .ZN(n1454) );
  INV_X1 U1461 ( .A(n1508), .ZN(n1507) );
  OR2_X1 U1462 ( .A1(n1509), .A2(n1510), .ZN(n1508) );
  AND2_X1 U1463 ( .A1(n1510), .A2(n1509), .ZN(n1506) );
  AND2_X1 U1464 ( .A1(n1511), .A2(n1512), .ZN(n1509) );
  OR2_X1 U1465 ( .A1(n1513), .A2(n1514), .ZN(n1512) );
  INV_X1 U1466 ( .A(n1515), .ZN(n1511) );
  AND2_X1 U1467 ( .A1(n1514), .A2(n1513), .ZN(n1515) );
  INV_X1 U1468 ( .A(n1050), .ZN(n1053) );
  OR2_X1 U1469 ( .A1(n1516), .A2(n1517), .ZN(n1050) );
  AND2_X1 U1470 ( .A1(n1031), .A2(n1030), .ZN(n1517) );
  AND2_X1 U1471 ( .A1(n1025), .A2(n1518), .ZN(n1516) );
  OR2_X1 U1472 ( .A1(n1030), .A2(n1031), .ZN(n1518) );
  OR2_X1 U1473 ( .A1(n1336), .A2(n1318), .ZN(n1031) );
  OR2_X1 U1474 ( .A1(n1519), .A2(n1520), .ZN(n1030) );
  AND2_X1 U1475 ( .A1(n1521), .A2(n979), .ZN(n1520) );
  AND2_X1 U1476 ( .A1(n974), .A2(n1522), .ZN(n1519) );
  OR2_X1 U1477 ( .A1(n979), .A2(n1521), .ZN(n1522) );
  INV_X1 U1478 ( .A(n978), .ZN(n1521) );
  AND2_X1 U1479 ( .A1(b_7_), .A2(a_1_), .ZN(n978) );
  OR2_X1 U1480 ( .A1(n1523), .A2(n1524), .ZN(n979) );
  AND2_X1 U1481 ( .A1(n1259), .A2(n1258), .ZN(n1524) );
  AND2_X1 U1482 ( .A1(n1253), .A2(n1525), .ZN(n1523) );
  OR2_X1 U1483 ( .A1(n1259), .A2(n1258), .ZN(n1525) );
  OR2_X1 U1484 ( .A1(n1526), .A2(n1527), .ZN(n1258) );
  AND2_X1 U1485 ( .A1(n1224), .A2(n1223), .ZN(n1527) );
  AND2_X1 U1486 ( .A1(n1218), .A2(n1528), .ZN(n1526) );
  OR2_X1 U1487 ( .A1(n1224), .A2(n1223), .ZN(n1528) );
  OR2_X1 U1488 ( .A1(n1529), .A2(n1530), .ZN(n1223) );
  AND2_X1 U1489 ( .A1(n1189), .A2(n1188), .ZN(n1530) );
  AND2_X1 U1490 ( .A1(n1183), .A2(n1531), .ZN(n1529) );
  OR2_X1 U1491 ( .A1(n1189), .A2(n1188), .ZN(n1531) );
  OR2_X1 U1492 ( .A1(n1532), .A2(n1533), .ZN(n1188) );
  AND2_X1 U1493 ( .A1(n1155), .A2(n1153), .ZN(n1533) );
  AND2_X1 U1494 ( .A1(n1148), .A2(n1534), .ZN(n1532) );
  OR2_X1 U1495 ( .A1(n1155), .A2(n1153), .ZN(n1534) );
  OR2_X1 U1496 ( .A1(n1535), .A2(n1140), .ZN(n1153) );
  INV_X1 U1497 ( .A(n1113), .ZN(n1140) );
  AND2_X1 U1498 ( .A1(a_7_), .A2(b_7_), .ZN(n1113) );
  OR2_X1 U1499 ( .A1(n1175), .A2(n1336), .ZN(n1155) );
  AND2_X1 U1500 ( .A1(n1536), .A2(n1537), .ZN(n1148) );
  OR2_X1 U1501 ( .A1(n1538), .A2(n1286), .ZN(n1537) );
  OR2_X1 U1502 ( .A1(n1535), .A2(n1539), .ZN(n1536) );
  OR2_X1 U1503 ( .A1(n1210), .A2(n1336), .ZN(n1189) );
  AND2_X1 U1504 ( .A1(n1540), .A2(n1541), .ZN(n1183) );
  INV_X1 U1505 ( .A(n1542), .ZN(n1541) );
  AND2_X1 U1506 ( .A1(n1543), .A2(n1544), .ZN(n1542) );
  OR2_X1 U1507 ( .A1(n1544), .A2(n1543), .ZN(n1540) );
  OR2_X1 U1508 ( .A1(n1545), .A2(n1546), .ZN(n1543) );
  AND2_X1 U1509 ( .A1(n1547), .A2(n1548), .ZN(n1546) );
  INV_X1 U1510 ( .A(n1549), .ZN(n1545) );
  OR2_X1 U1511 ( .A1(n1548), .A2(n1547), .ZN(n1549) );
  OR2_X1 U1512 ( .A1(n1245), .A2(n1336), .ZN(n1224) );
  AND2_X1 U1513 ( .A1(n1550), .A2(n1551), .ZN(n1218) );
  INV_X1 U1514 ( .A(n1552), .ZN(n1551) );
  AND2_X1 U1515 ( .A1(n1553), .A2(n1554), .ZN(n1552) );
  OR2_X1 U1516 ( .A1(n1554), .A2(n1553), .ZN(n1550) );
  OR2_X1 U1517 ( .A1(n1555), .A2(n1556), .ZN(n1553) );
  INV_X1 U1518 ( .A(n1557), .ZN(n1556) );
  OR2_X1 U1519 ( .A1(n1558), .A2(n1559), .ZN(n1557) );
  AND2_X1 U1520 ( .A1(n1559), .A2(n1558), .ZN(n1555) );
  INV_X1 U1521 ( .A(n1560), .ZN(n1559) );
  OR2_X1 U1522 ( .A1(n1042), .A2(n1336), .ZN(n1259) );
  INV_X1 U1523 ( .A(b_7_), .ZN(n1336) );
  AND2_X1 U1524 ( .A1(n1561), .A2(n1562), .ZN(n1253) );
  INV_X1 U1525 ( .A(n1563), .ZN(n1562) );
  AND2_X1 U1526 ( .A1(n1564), .A2(n1565), .ZN(n1563) );
  OR2_X1 U1527 ( .A1(n1565), .A2(n1564), .ZN(n1561) );
  OR2_X1 U1528 ( .A1(n1566), .A2(n1567), .ZN(n1564) );
  INV_X1 U1529 ( .A(n1568), .ZN(n1567) );
  OR2_X1 U1530 ( .A1(n1569), .A2(n1570), .ZN(n1568) );
  AND2_X1 U1531 ( .A1(n1570), .A2(n1569), .ZN(n1566) );
  INV_X1 U1532 ( .A(n1571), .ZN(n1570) );
  OR2_X1 U1533 ( .A1(n1572), .A2(n1573), .ZN(n974) );
  INV_X1 U1534 ( .A(n1574), .ZN(n1573) );
  OR2_X1 U1535 ( .A1(n1575), .A2(n1576), .ZN(n1574) );
  AND2_X1 U1536 ( .A1(n1576), .A2(n1575), .ZN(n1572) );
  AND2_X1 U1537 ( .A1(n1577), .A2(n1578), .ZN(n1575) );
  INV_X1 U1538 ( .A(n1579), .ZN(n1578) );
  AND2_X1 U1539 ( .A1(n1580), .A2(n1581), .ZN(n1579) );
  OR2_X1 U1540 ( .A1(n1581), .A2(n1580), .ZN(n1577) );
  AND2_X1 U1541 ( .A1(n1582), .A2(n1583), .ZN(n1025) );
  INV_X1 U1542 ( .A(n1584), .ZN(n1583) );
  AND2_X1 U1543 ( .A1(n1585), .A2(n1478), .ZN(n1584) );
  OR2_X1 U1544 ( .A1(n1478), .A2(n1585), .ZN(n1582) );
  OR2_X1 U1545 ( .A1(n1586), .A2(n1587), .ZN(n1585) );
  INV_X1 U1546 ( .A(n1588), .ZN(n1587) );
  OR2_X1 U1547 ( .A1(n1476), .A2(n1589), .ZN(n1588) );
  AND2_X1 U1548 ( .A1(n1589), .A2(n1476), .ZN(n1586) );
  OR2_X1 U1549 ( .A1(n1337), .A2(n1002), .ZN(n1476) );
  INV_X1 U1550 ( .A(n1477), .ZN(n1589) );
  OR2_X1 U1551 ( .A1(n1590), .A2(n1591), .ZN(n1477) );
  AND2_X1 U1552 ( .A1(n1592), .A2(n1581), .ZN(n1591) );
  AND2_X1 U1553 ( .A1(n1576), .A2(n1593), .ZN(n1590) );
  OR2_X1 U1554 ( .A1(n1581), .A2(n1592), .ZN(n1593) );
  INV_X1 U1555 ( .A(n1580), .ZN(n1592) );
  AND2_X1 U1556 ( .A1(b_6_), .A2(a_2_), .ZN(n1580) );
  OR2_X1 U1557 ( .A1(n1594), .A2(n1595), .ZN(n1581) );
  AND2_X1 U1558 ( .A1(n1569), .A2(n1571), .ZN(n1595) );
  AND2_X1 U1559 ( .A1(n1565), .A2(n1596), .ZN(n1594) );
  OR2_X1 U1560 ( .A1(n1569), .A2(n1571), .ZN(n1596) );
  OR2_X1 U1561 ( .A1(n1597), .A2(n1598), .ZN(n1571) );
  AND2_X1 U1562 ( .A1(n1558), .A2(n1560), .ZN(n1598) );
  AND2_X1 U1563 ( .A1(n1554), .A2(n1599), .ZN(n1597) );
  OR2_X1 U1564 ( .A1(n1558), .A2(n1560), .ZN(n1599) );
  OR2_X1 U1565 ( .A1(n1600), .A2(n1601), .ZN(n1560) );
  AND2_X1 U1566 ( .A1(n1602), .A2(n1548), .ZN(n1601) );
  AND2_X1 U1567 ( .A1(n1544), .A2(n1603), .ZN(n1600) );
  OR2_X1 U1568 ( .A1(n1602), .A2(n1548), .ZN(n1603) );
  OR2_X1 U1569 ( .A1(n1538), .A2(n1535), .ZN(n1548) );
  INV_X1 U1570 ( .A(n1286), .ZN(n1535) );
  AND2_X1 U1571 ( .A1(a_6_), .A2(b_6_), .ZN(n1286) );
  INV_X1 U1572 ( .A(n1539), .ZN(n1538) );
  AND2_X1 U1573 ( .A1(a_7_), .A2(b_5_), .ZN(n1539) );
  INV_X1 U1574 ( .A(n1547), .ZN(n1602) );
  AND2_X1 U1575 ( .A1(a_5_), .A2(b_6_), .ZN(n1547) );
  AND2_X1 U1576 ( .A1(n1604), .A2(n1605), .ZN(n1544) );
  OR2_X1 U1577 ( .A1(n1606), .A2(n1607), .ZN(n1605) );
  OR2_X1 U1578 ( .A1(n1608), .A2(n1609), .ZN(n1604) );
  INV_X1 U1579 ( .A(n1607), .ZN(n1608) );
  OR2_X1 U1580 ( .A1(n1210), .A2(n1337), .ZN(n1558) );
  AND2_X1 U1581 ( .A1(n1610), .A2(n1611), .ZN(n1554) );
  INV_X1 U1582 ( .A(n1612), .ZN(n1611) );
  AND2_X1 U1583 ( .A1(n1613), .A2(n1614), .ZN(n1612) );
  OR2_X1 U1584 ( .A1(n1614), .A2(n1613), .ZN(n1610) );
  OR2_X1 U1585 ( .A1(n1615), .A2(n1616), .ZN(n1613) );
  AND2_X1 U1586 ( .A1(n1617), .A2(n1618), .ZN(n1616) );
  INV_X1 U1587 ( .A(n1284), .ZN(n1617) );
  AND2_X1 U1588 ( .A1(n1619), .A2(n1284), .ZN(n1615) );
  OR2_X1 U1589 ( .A1(n1245), .A2(n1337), .ZN(n1569) );
  INV_X1 U1590 ( .A(b_6_), .ZN(n1337) );
  AND2_X1 U1591 ( .A1(n1620), .A2(n1621), .ZN(n1565) );
  INV_X1 U1592 ( .A(n1622), .ZN(n1621) );
  AND2_X1 U1593 ( .A1(n1623), .A2(n1624), .ZN(n1622) );
  OR2_X1 U1594 ( .A1(n1624), .A2(n1623), .ZN(n1620) );
  OR2_X1 U1595 ( .A1(n1625), .A2(n1626), .ZN(n1623) );
  INV_X1 U1596 ( .A(n1627), .ZN(n1626) );
  OR2_X1 U1597 ( .A1(n1628), .A2(n1629), .ZN(n1627) );
  AND2_X1 U1598 ( .A1(n1629), .A2(n1628), .ZN(n1625) );
  INV_X1 U1599 ( .A(n1630), .ZN(n1629) );
  OR2_X1 U1600 ( .A1(n1631), .A2(n1632), .ZN(n1576) );
  INV_X1 U1601 ( .A(n1633), .ZN(n1632) );
  OR2_X1 U1602 ( .A1(n1634), .A2(n1635), .ZN(n1633) );
  AND2_X1 U1603 ( .A1(n1635), .A2(n1634), .ZN(n1631) );
  AND2_X1 U1604 ( .A1(n1636), .A2(n1637), .ZN(n1634) );
  INV_X1 U1605 ( .A(n1638), .ZN(n1637) );
  AND2_X1 U1606 ( .A1(n1639), .A2(n1640), .ZN(n1638) );
  OR2_X1 U1607 ( .A1(n1640), .A2(n1639), .ZN(n1636) );
  AND2_X1 U1608 ( .A1(n1641), .A2(n1642), .ZN(n1478) );
  INV_X1 U1609 ( .A(n1643), .ZN(n1642) );
  AND2_X1 U1610 ( .A1(n1644), .A2(n1491), .ZN(n1643) );
  OR2_X1 U1611 ( .A1(n1491), .A2(n1644), .ZN(n1641) );
  OR2_X1 U1612 ( .A1(n1645), .A2(n1646), .ZN(n1644) );
  INV_X1 U1613 ( .A(n1647), .ZN(n1646) );
  OR2_X1 U1614 ( .A1(n1489), .A2(n1648), .ZN(n1647) );
  AND2_X1 U1615 ( .A1(n1648), .A2(n1489), .ZN(n1645) );
  OR2_X1 U1616 ( .A1(n1174), .A2(n1042), .ZN(n1489) );
  INV_X1 U1617 ( .A(n1490), .ZN(n1648) );
  OR2_X1 U1618 ( .A1(n1649), .A2(n1650), .ZN(n1490) );
  AND2_X1 U1619 ( .A1(n1651), .A2(n1640), .ZN(n1650) );
  AND2_X1 U1620 ( .A1(n1635), .A2(n1652), .ZN(n1649) );
  OR2_X1 U1621 ( .A1(n1640), .A2(n1651), .ZN(n1652) );
  INV_X1 U1622 ( .A(n1639), .ZN(n1651) );
  AND2_X1 U1623 ( .A1(b_5_), .A2(a_3_), .ZN(n1639) );
  OR2_X1 U1624 ( .A1(n1653), .A2(n1654), .ZN(n1640) );
  AND2_X1 U1625 ( .A1(n1628), .A2(n1630), .ZN(n1654) );
  AND2_X1 U1626 ( .A1(n1624), .A2(n1655), .ZN(n1653) );
  OR2_X1 U1627 ( .A1(n1628), .A2(n1630), .ZN(n1655) );
  OR2_X1 U1628 ( .A1(n1656), .A2(n1657), .ZN(n1630) );
  AND2_X1 U1629 ( .A1(n1284), .A2(n1618), .ZN(n1657) );
  AND2_X1 U1630 ( .A1(n1614), .A2(n1658), .ZN(n1656) );
  OR2_X1 U1631 ( .A1(n1284), .A2(n1618), .ZN(n1658) );
  INV_X1 U1632 ( .A(n1619), .ZN(n1618) );
  AND2_X1 U1633 ( .A1(n1609), .A2(n1607), .ZN(n1619) );
  AND2_X1 U1634 ( .A1(a_6_), .A2(b_5_), .ZN(n1607) );
  OR2_X1 U1635 ( .A1(n1175), .A2(n1174), .ZN(n1284) );
  AND2_X1 U1636 ( .A1(n1659), .A2(n1660), .ZN(n1614) );
  OR3_X1 U1637 ( .A1(n1209), .A2(n1335), .A3(n1661), .ZN(n1660) );
  INV_X1 U1638 ( .A(n1662), .ZN(n1659) );
  AND2_X1 U1639 ( .A1(n1661), .A2(n1663), .ZN(n1662) );
  OR2_X1 U1640 ( .A1(n1335), .A2(n1209), .ZN(n1663) );
  AND2_X1 U1641 ( .A1(b_3_), .A2(a_7_), .ZN(n1661) );
  OR2_X1 U1642 ( .A1(n1210), .A2(n1174), .ZN(n1628) );
  INV_X1 U1643 ( .A(b_5_), .ZN(n1174) );
  AND2_X1 U1644 ( .A1(n1664), .A2(n1665), .ZN(n1624) );
  INV_X1 U1645 ( .A(n1666), .ZN(n1665) );
  AND2_X1 U1646 ( .A1(n1667), .A2(n1668), .ZN(n1666) );
  OR2_X1 U1647 ( .A1(n1668), .A2(n1667), .ZN(n1664) );
  OR2_X1 U1648 ( .A1(n1669), .A2(n1670), .ZN(n1667) );
  AND2_X1 U1649 ( .A1(n1671), .A2(n1672), .ZN(n1670) );
  INV_X1 U1650 ( .A(n1673), .ZN(n1669) );
  OR2_X1 U1651 ( .A1(n1672), .A2(n1671), .ZN(n1673) );
  OR2_X1 U1652 ( .A1(n1674), .A2(n1675), .ZN(n1635) );
  INV_X1 U1653 ( .A(n1676), .ZN(n1675) );
  OR2_X1 U1654 ( .A1(n1677), .A2(n1678), .ZN(n1676) );
  AND2_X1 U1655 ( .A1(n1678), .A2(n1677), .ZN(n1674) );
  AND2_X1 U1656 ( .A1(n1679), .A2(n1680), .ZN(n1677) );
  OR2_X1 U1657 ( .A1(n1681), .A2(n1682), .ZN(n1680) );
  INV_X1 U1658 ( .A(n1683), .ZN(n1679) );
  AND2_X1 U1659 ( .A1(n1682), .A2(n1681), .ZN(n1683) );
  AND2_X1 U1660 ( .A1(n1684), .A2(n1685), .ZN(n1491) );
  INV_X1 U1661 ( .A(n1686), .ZN(n1685) );
  AND2_X1 U1662 ( .A1(n1687), .A2(n1504), .ZN(n1686) );
  OR2_X1 U1663 ( .A1(n1504), .A2(n1687), .ZN(n1684) );
  OR2_X1 U1664 ( .A1(n1688), .A2(n1689), .ZN(n1687) );
  INV_X1 U1665 ( .A(n1690), .ZN(n1689) );
  OR2_X1 U1666 ( .A1(n1502), .A2(n1691), .ZN(n1690) );
  AND2_X1 U1667 ( .A1(n1691), .A2(n1502), .ZN(n1688) );
  OR2_X1 U1668 ( .A1(n1209), .A2(n1245), .ZN(n1502) );
  INV_X1 U1669 ( .A(b_4_), .ZN(n1209) );
  INV_X1 U1670 ( .A(n1503), .ZN(n1691) );
  OR2_X1 U1671 ( .A1(n1692), .A2(n1693), .ZN(n1503) );
  AND2_X1 U1672 ( .A1(n1681), .A2(n1281), .ZN(n1693) );
  AND2_X1 U1673 ( .A1(n1678), .A2(n1694), .ZN(n1692) );
  OR2_X1 U1674 ( .A1(n1281), .A2(n1681), .ZN(n1694) );
  OR2_X1 U1675 ( .A1(n1695), .A2(n1696), .ZN(n1681) );
  AND2_X1 U1676 ( .A1(n1697), .A2(n1672), .ZN(n1696) );
  AND2_X1 U1677 ( .A1(n1668), .A2(n1698), .ZN(n1695) );
  OR2_X1 U1678 ( .A1(n1697), .A2(n1672), .ZN(n1698) );
  OR2_X1 U1679 ( .A1(n1699), .A2(n1606), .ZN(n1672) );
  INV_X1 U1680 ( .A(n1609), .ZN(n1606) );
  AND2_X1 U1681 ( .A1(a_7_), .A2(b_4_), .ZN(n1609) );
  INV_X1 U1682 ( .A(n1671), .ZN(n1697) );
  AND2_X1 U1683 ( .A1(a_5_), .A2(b_4_), .ZN(n1671) );
  AND2_X1 U1684 ( .A1(n1700), .A2(n1701), .ZN(n1668) );
  OR2_X1 U1685 ( .A1(n1702), .A2(n1703), .ZN(n1701) );
  INV_X1 U1686 ( .A(n1699), .ZN(n1703) );
  OR2_X1 U1687 ( .A1(n1699), .A2(n1704), .ZN(n1700) );
  INV_X1 U1688 ( .A(n1682), .ZN(n1281) );
  AND2_X1 U1689 ( .A1(a_4_), .A2(b_4_), .ZN(n1682) );
  OR2_X1 U1690 ( .A1(n1705), .A2(n1706), .ZN(n1678) );
  AND2_X1 U1691 ( .A1(n1707), .A2(n1708), .ZN(n1706) );
  INV_X1 U1692 ( .A(n1709), .ZN(n1705) );
  OR2_X1 U1693 ( .A1(n1707), .A2(n1708), .ZN(n1709) );
  OR2_X1 U1694 ( .A1(n1710), .A2(n1711), .ZN(n1707) );
  AND2_X1 U1695 ( .A1(n1712), .A2(n1713), .ZN(n1711) );
  AND2_X1 U1696 ( .A1(n1714), .A2(n1715), .ZN(n1710) );
  AND2_X1 U1697 ( .A1(n1716), .A2(n1717), .ZN(n1504) );
  INV_X1 U1698 ( .A(n1718), .ZN(n1717) );
  AND2_X1 U1699 ( .A1(n1719), .A2(n1720), .ZN(n1718) );
  OR2_X1 U1700 ( .A1(n1720), .A2(n1719), .ZN(n1716) );
  OR2_X1 U1701 ( .A1(n1721), .A2(n1722), .ZN(n1719) );
  AND2_X1 U1702 ( .A1(n1723), .A2(n1724), .ZN(n1722) );
  INV_X1 U1703 ( .A(n1725), .ZN(n1723) );
  AND2_X1 U1704 ( .A1(n1726), .A2(n1725), .ZN(n1721) );
  OR2_X1 U1705 ( .A1(n1727), .A2(n1354), .ZN(n1349) );
  OR2_X1 U1706 ( .A1(n1728), .A2(n1729), .ZN(n1354) );
  AND2_X1 U1707 ( .A1(n1375), .A2(n1374), .ZN(n1729) );
  AND2_X1 U1708 ( .A1(n1370), .A2(n1730), .ZN(n1728) );
  OR2_X1 U1709 ( .A1(n1374), .A2(n1375), .ZN(n1730) );
  OR2_X1 U1710 ( .A1(n1731), .A2(n1732), .ZN(n1375) );
  AND2_X1 U1711 ( .A1(n1406), .A2(n1405), .ZN(n1732) );
  AND2_X1 U1712 ( .A1(n1401), .A2(n1733), .ZN(n1731) );
  OR2_X1 U1713 ( .A1(n1405), .A2(n1406), .ZN(n1733) );
  OR2_X1 U1714 ( .A1(n1734), .A2(n1735), .ZN(n1406) );
  AND2_X1 U1715 ( .A1(n1464), .A2(n1736), .ZN(n1735) );
  AND2_X1 U1716 ( .A1(n1461), .A2(n1737), .ZN(n1734) );
  OR2_X1 U1717 ( .A1(n1736), .A2(n1464), .ZN(n1737) );
  OR2_X1 U1718 ( .A1(n1738), .A2(n1739), .ZN(n1464) );
  AND2_X1 U1719 ( .A1(n1513), .A2(n1278), .ZN(n1739) );
  AND2_X1 U1720 ( .A1(n1510), .A2(n1740), .ZN(n1738) );
  OR2_X1 U1721 ( .A1(n1278), .A2(n1513), .ZN(n1740) );
  OR2_X1 U1722 ( .A1(n1741), .A2(n1742), .ZN(n1513) );
  AND2_X1 U1723 ( .A1(n1725), .A2(n1724), .ZN(n1742) );
  AND2_X1 U1724 ( .A1(n1720), .A2(n1743), .ZN(n1741) );
  OR2_X1 U1725 ( .A1(n1724), .A2(n1725), .ZN(n1743) );
  OR2_X1 U1726 ( .A1(n1744), .A2(n1745), .ZN(n1725) );
  AND2_X1 U1727 ( .A1(n1708), .A2(n1715), .ZN(n1745) );
  AND2_X1 U1728 ( .A1(n1714), .A2(n1746), .ZN(n1744) );
  OR2_X1 U1729 ( .A1(n1715), .A2(n1708), .ZN(n1746) );
  OR2_X1 U1730 ( .A1(n1702), .A2(n1699), .ZN(n1708) );
  OR2_X1 U1731 ( .A1(n1335), .A2(n1244), .ZN(n1699) );
  INV_X1 U1732 ( .A(b_3_), .ZN(n1244) );
  INV_X1 U1733 ( .A(n1712), .ZN(n1715) );
  AND2_X1 U1734 ( .A1(b_3_), .A2(a_5_), .ZN(n1712) );
  INV_X1 U1735 ( .A(n1713), .ZN(n1714) );
  OR2_X1 U1736 ( .A1(n1747), .A2(n1748), .ZN(n1713) );
  AND3_X1 U1737 ( .A1(a_7_), .A2(n1749), .A3(b_1_), .ZN(n1748) );
  OR2_X1 U1738 ( .A1(n1335), .A2(n1043), .ZN(n1749) );
  AND3_X1 U1739 ( .A1(a_6_), .A2(n1750), .A3(b_2_), .ZN(n1747) );
  OR2_X1 U1740 ( .A1(n1316), .A2(n1001), .ZN(n1750) );
  INV_X1 U1741 ( .A(a_7_), .ZN(n1316) );
  INV_X1 U1742 ( .A(n1726), .ZN(n1724) );
  AND2_X1 U1743 ( .A1(b_3_), .A2(a_4_), .ZN(n1726) );
  AND2_X1 U1744 ( .A1(n1751), .A2(n1752), .ZN(n1720) );
  INV_X1 U1745 ( .A(n1753), .ZN(n1752) );
  AND2_X1 U1746 ( .A1(n1754), .A2(n1755), .ZN(n1753) );
  OR2_X1 U1747 ( .A1(n1755), .A2(n1754), .ZN(n1751) );
  OR2_X1 U1748 ( .A1(n1756), .A2(n1757), .ZN(n1754) );
  INV_X1 U1749 ( .A(n1758), .ZN(n1757) );
  OR2_X1 U1750 ( .A1(n1759), .A2(n1760), .ZN(n1758) );
  AND2_X1 U1751 ( .A1(n1760), .A2(n1759), .ZN(n1756) );
  INV_X1 U1752 ( .A(n1761), .ZN(n1760) );
  INV_X1 U1753 ( .A(n1514), .ZN(n1278) );
  AND2_X1 U1754 ( .A1(b_3_), .A2(a_3_), .ZN(n1514) );
  OR2_X1 U1755 ( .A1(n1762), .A2(n1763), .ZN(n1510) );
  INV_X1 U1756 ( .A(n1764), .ZN(n1763) );
  OR2_X1 U1757 ( .A1(n1765), .A2(n1766), .ZN(n1764) );
  AND2_X1 U1758 ( .A1(n1766), .A2(n1765), .ZN(n1762) );
  AND2_X1 U1759 ( .A1(n1767), .A2(n1768), .ZN(n1765) );
  INV_X1 U1760 ( .A(n1769), .ZN(n1768) );
  AND2_X1 U1761 ( .A1(n1770), .A2(n1771), .ZN(n1769) );
  OR2_X1 U1762 ( .A1(n1771), .A2(n1770), .ZN(n1767) );
  INV_X1 U1763 ( .A(n1465), .ZN(n1736) );
  AND2_X1 U1764 ( .A1(b_3_), .A2(a_2_), .ZN(n1465) );
  OR2_X1 U1765 ( .A1(n1772), .A2(n1773), .ZN(n1461) );
  INV_X1 U1766 ( .A(n1774), .ZN(n1773) );
  OR2_X1 U1767 ( .A1(n1775), .A2(n1776), .ZN(n1774) );
  AND2_X1 U1768 ( .A1(n1776), .A2(n1775), .ZN(n1772) );
  AND2_X1 U1769 ( .A1(n1777), .A2(n1778), .ZN(n1775) );
  OR2_X1 U1770 ( .A1(n1779), .A2(n1780), .ZN(n1778) );
  INV_X1 U1771 ( .A(n1781), .ZN(n1777) );
  AND2_X1 U1772 ( .A1(n1780), .A2(n1779), .ZN(n1781) );
  INV_X1 U1773 ( .A(n1407), .ZN(n1405) );
  AND2_X1 U1774 ( .A1(b_3_), .A2(a_1_), .ZN(n1407) );
  AND2_X1 U1775 ( .A1(n1782), .A2(n1783), .ZN(n1401) );
  INV_X1 U1776 ( .A(n1784), .ZN(n1783) );
  AND2_X1 U1777 ( .A1(n1785), .A2(n1786), .ZN(n1784) );
  OR2_X1 U1778 ( .A1(n1786), .A2(n1785), .ZN(n1782) );
  OR2_X1 U1779 ( .A1(n1787), .A2(n1788), .ZN(n1785) );
  AND2_X1 U1780 ( .A1(n1789), .A2(n1045), .ZN(n1788) );
  INV_X1 U1781 ( .A(n1790), .ZN(n1789) );
  AND2_X1 U1782 ( .A1(n1791), .A2(n1790), .ZN(n1787) );
  INV_X1 U1783 ( .A(n1376), .ZN(n1374) );
  AND2_X1 U1784 ( .A1(b_3_), .A2(a_0_), .ZN(n1376) );
  AND2_X1 U1785 ( .A1(n1792), .A2(n1793), .ZN(n1370) );
  INV_X1 U1786 ( .A(n1794), .ZN(n1793) );
  AND2_X1 U1787 ( .A1(n1795), .A2(n1796), .ZN(n1794) );
  OR2_X1 U1788 ( .A1(n1796), .A2(n1795), .ZN(n1792) );
  OR2_X1 U1789 ( .A1(n1797), .A2(n1798), .ZN(n1795) );
  INV_X1 U1790 ( .A(n1799), .ZN(n1798) );
  OR2_X1 U1791 ( .A1(n1800), .A2(n1801), .ZN(n1799) );
  AND2_X1 U1792 ( .A1(n1801), .A2(n1800), .ZN(n1797) );
  INV_X1 U1793 ( .A(n1802), .ZN(n1801) );
  AND2_X1 U1794 ( .A1(n1352), .A2(n1353), .ZN(n1727) );
  OR2_X1 U1795 ( .A1(n1803), .A2(n1804), .ZN(n1353) );
  OR2_X1 U1796 ( .A1(n1805), .A2(n1806), .ZN(n1352) );
  INV_X1 U1797 ( .A(n1804), .ZN(n1805) );
  AND2_X1 U1798 ( .A1(n1807), .A2(n1808), .ZN(n1804) );
  INV_X1 U1799 ( .A(n1809), .ZN(n1808) );
  AND2_X1 U1800 ( .A1(n1810), .A2(n1811), .ZN(n1809) );
  OR2_X1 U1801 ( .A1(n1811), .A2(n1810), .ZN(n1807) );
  INV_X1 U1802 ( .A(n1812), .ZN(n1810) );
  AND2_X1 U1803 ( .A1(n1109), .A2(n1106), .ZN(n1340) );
  INV_X1 U1804 ( .A(n1108), .ZN(n1106) );
  AND2_X1 U1805 ( .A1(n1813), .A2(n1814), .ZN(n1108) );
  INV_X1 U1806 ( .A(n1815), .ZN(n1814) );
  AND2_X1 U1807 ( .A1(n1816), .A2(n1344), .ZN(n1815) );
  OR2_X1 U1808 ( .A1(n1344), .A2(n1816), .ZN(n1813) );
  AND2_X1 U1809 ( .A1(b_0_), .A2(a_0_), .ZN(n1816) );
  OR2_X1 U1810 ( .A1(n1817), .A2(n1818), .ZN(n1344) );
  AND2_X1 U1811 ( .A1(n1819), .A2(n1820), .ZN(n1818) );
  AND2_X1 U1812 ( .A1(n1821), .A2(n1822), .ZN(n1817) );
  OR2_X1 U1813 ( .A1(n1820), .A2(n1819), .ZN(n1821) );
  INV_X1 U1814 ( .A(n1107), .ZN(n1109) );
  OR2_X1 U1815 ( .A1(n1347), .A2(n1348), .ZN(n1107) );
  OR2_X1 U1816 ( .A1(n1823), .A2(n1824), .ZN(n1348) );
  AND2_X1 U1817 ( .A1(n1812), .A2(n1811), .ZN(n1824) );
  AND2_X1 U1818 ( .A1(n1806), .A2(n1825), .ZN(n1823) );
  OR2_X1 U1819 ( .A1(n1811), .A2(n1812), .ZN(n1825) );
  OR2_X1 U1820 ( .A1(n1043), .A2(n1318), .ZN(n1812) );
  OR2_X1 U1821 ( .A1(n1826), .A2(n1827), .ZN(n1811) );
  AND2_X1 U1822 ( .A1(n1800), .A2(n1802), .ZN(n1827) );
  AND2_X1 U1823 ( .A1(n1796), .A2(n1828), .ZN(n1826) );
  OR2_X1 U1824 ( .A1(n1802), .A2(n1800), .ZN(n1828) );
  OR2_X1 U1825 ( .A1(n1043), .A2(n1002), .ZN(n1800) );
  OR2_X1 U1826 ( .A1(n1829), .A2(n1830), .ZN(n1802) );
  AND2_X1 U1827 ( .A1(n1790), .A2(n1045), .ZN(n1830) );
  AND2_X1 U1828 ( .A1(n1786), .A2(n1831), .ZN(n1829) );
  OR2_X1 U1829 ( .A1(n1045), .A2(n1790), .ZN(n1831) );
  OR2_X1 U1830 ( .A1(n1832), .A2(n1833), .ZN(n1790) );
  AND2_X1 U1831 ( .A1(n1779), .A2(n1834), .ZN(n1833) );
  AND2_X1 U1832 ( .A1(n1776), .A2(n1835), .ZN(n1832) );
  OR2_X1 U1833 ( .A1(n1834), .A2(n1779), .ZN(n1835) );
  OR2_X1 U1834 ( .A1(n1836), .A2(n1837), .ZN(n1779) );
  AND2_X1 U1835 ( .A1(n1838), .A2(n1771), .ZN(n1837) );
  AND2_X1 U1836 ( .A1(n1766), .A2(n1839), .ZN(n1836) );
  OR2_X1 U1837 ( .A1(n1771), .A2(n1838), .ZN(n1839) );
  INV_X1 U1838 ( .A(n1770), .ZN(n1838) );
  AND2_X1 U1839 ( .A1(b_2_), .A2(a_4_), .ZN(n1770) );
  OR2_X1 U1840 ( .A1(n1840), .A2(n1841), .ZN(n1771) );
  AND2_X1 U1841 ( .A1(n1759), .A2(n1761), .ZN(n1841) );
  AND2_X1 U1842 ( .A1(n1755), .A2(n1842), .ZN(n1840) );
  OR2_X1 U1843 ( .A1(n1761), .A2(n1759), .ZN(n1842) );
  OR2_X1 U1844 ( .A1(n1043), .A2(n1175), .ZN(n1759) );
  INV_X1 U1845 ( .A(b_2_), .ZN(n1043) );
  OR2_X1 U1846 ( .A1(n1702), .A2(n1843), .ZN(n1761) );
  INV_X1 U1847 ( .A(n1704), .ZN(n1702) );
  AND2_X1 U1848 ( .A1(a_7_), .A2(b_2_), .ZN(n1704) );
  AND2_X1 U1849 ( .A1(n1844), .A2(n1845), .ZN(n1755) );
  OR2_X1 U1850 ( .A1(n1846), .A2(n1847), .ZN(n1845) );
  INV_X1 U1851 ( .A(n1848), .ZN(n1846) );
  OR2_X1 U1852 ( .A1(n1843), .A2(n1848), .ZN(n1844) );
  OR2_X1 U1853 ( .A1(n1849), .A2(n1850), .ZN(n1766) );
  INV_X1 U1854 ( .A(n1851), .ZN(n1850) );
  OR2_X1 U1855 ( .A1(n1852), .A2(n1853), .ZN(n1851) );
  AND2_X1 U1856 ( .A1(n1853), .A2(n1852), .ZN(n1849) );
  OR2_X1 U1857 ( .A1(n1854), .A2(n1855), .ZN(n1852) );
  AND3_X1 U1858 ( .A1(a_6_), .A2(n1856), .A3(b_0_), .ZN(n1855) );
  OR2_X1 U1859 ( .A1(n1001), .A2(n1175), .ZN(n1856) );
  INV_X1 U1860 ( .A(a_5_), .ZN(n1175) );
  AND3_X1 U1861 ( .A1(b_1_), .A2(n1857), .A3(a_5_), .ZN(n1854) );
  OR2_X1 U1862 ( .A1(n1335), .A2(n1338), .ZN(n1857) );
  INV_X1 U1863 ( .A(n1780), .ZN(n1834) );
  AND2_X1 U1864 ( .A1(b_2_), .A2(a_3_), .ZN(n1780) );
  OR2_X1 U1865 ( .A1(n1858), .A2(n1859), .ZN(n1776) );
  AND2_X1 U1866 ( .A1(n1860), .A2(n1861), .ZN(n1859) );
  INV_X1 U1867 ( .A(n1862), .ZN(n1858) );
  OR2_X1 U1868 ( .A1(n1860), .A2(n1861), .ZN(n1862) );
  OR2_X1 U1869 ( .A1(n1863), .A2(n1864), .ZN(n1860) );
  AND2_X1 U1870 ( .A1(n1865), .A2(n1866), .ZN(n1864) );
  AND2_X1 U1871 ( .A1(n1867), .A2(n1868), .ZN(n1863) );
  INV_X1 U1872 ( .A(n1791), .ZN(n1045) );
  AND2_X1 U1873 ( .A1(b_2_), .A2(a_2_), .ZN(n1791) );
  AND2_X1 U1874 ( .A1(n1869), .A2(n1870), .ZN(n1786) );
  INV_X1 U1875 ( .A(n1871), .ZN(n1870) );
  AND2_X1 U1876 ( .A1(n1872), .A2(n1873), .ZN(n1871) );
  OR2_X1 U1877 ( .A1(n1872), .A2(n1873), .ZN(n1869) );
  OR2_X1 U1878 ( .A1(n1874), .A2(n1875), .ZN(n1872) );
  INV_X1 U1879 ( .A(n1876), .ZN(n1875) );
  OR2_X1 U1880 ( .A1(n1877), .A2(n1878), .ZN(n1876) );
  AND2_X1 U1881 ( .A1(n1878), .A2(n1877), .ZN(n1874) );
  INV_X1 U1882 ( .A(n1879), .ZN(n1878) );
  AND2_X1 U1883 ( .A1(n1880), .A2(n1881), .ZN(n1796) );
  INV_X1 U1884 ( .A(n1882), .ZN(n1881) );
  AND2_X1 U1885 ( .A1(n1883), .A2(n1884), .ZN(n1882) );
  OR2_X1 U1886 ( .A1(n1883), .A2(n1884), .ZN(n1880) );
  OR2_X1 U1887 ( .A1(n1885), .A2(n1886), .ZN(n1883) );
  INV_X1 U1888 ( .A(n1887), .ZN(n1886) );
  OR2_X1 U1889 ( .A1(n1888), .A2(n1889), .ZN(n1887) );
  AND2_X1 U1890 ( .A1(n1889), .A2(n1888), .ZN(n1885) );
  INV_X1 U1891 ( .A(n1890), .ZN(n1889) );
  INV_X1 U1892 ( .A(n1803), .ZN(n1806) );
  OR2_X1 U1893 ( .A1(n1891), .A2(n1892), .ZN(n1803) );
  AND2_X1 U1894 ( .A1(n1893), .A2(n1894), .ZN(n1892) );
  INV_X1 U1895 ( .A(n1895), .ZN(n1891) );
  OR2_X1 U1896 ( .A1(n1893), .A2(n1894), .ZN(n1895) );
  OR2_X1 U1897 ( .A1(n1896), .A2(n1897), .ZN(n1893) );
  AND2_X1 U1898 ( .A1(n1898), .A2(n1039), .ZN(n1897) );
  INV_X1 U1899 ( .A(n1899), .ZN(n1898) );
  AND2_X1 U1900 ( .A1(n1900), .A2(n1899), .ZN(n1896) );
  AND2_X1 U1901 ( .A1(n1901), .A2(n1902), .ZN(n1347) );
  INV_X1 U1902 ( .A(n1903), .ZN(n1902) );
  AND2_X1 U1903 ( .A1(n1904), .A2(n1819), .ZN(n1903) );
  OR2_X1 U1904 ( .A1(n1904), .A2(n1819), .ZN(n1901) );
  OR2_X1 U1905 ( .A1(n1002), .A2(n1338), .ZN(n1819) );
  INV_X1 U1906 ( .A(a_1_), .ZN(n1002) );
  OR2_X1 U1907 ( .A1(n1905), .A2(n1906), .ZN(n1904) );
  INV_X1 U1908 ( .A(n1907), .ZN(n1906) );
  OR2_X1 U1909 ( .A1(n1822), .A2(n1908), .ZN(n1907) );
  AND2_X1 U1910 ( .A1(n1908), .A2(n1822), .ZN(n1905) );
  OR2_X1 U1911 ( .A1(n1001), .A2(n1318), .ZN(n1822) );
  INV_X1 U1912 ( .A(a_0_), .ZN(n1318) );
  INV_X1 U1913 ( .A(n1820), .ZN(n1908) );
  OR2_X1 U1914 ( .A1(n1909), .A2(n1910), .ZN(n1820) );
  AND2_X1 U1915 ( .A1(n1894), .A2(n1899), .ZN(n1910) );
  AND2_X1 U1916 ( .A1(n1911), .A2(n1039), .ZN(n1909) );
  INV_X1 U1917 ( .A(n1900), .ZN(n1039) );
  AND2_X1 U1918 ( .A1(b_1_), .A2(a_1_), .ZN(n1900) );
  OR2_X1 U1919 ( .A1(n1899), .A2(n1894), .ZN(n1911) );
  OR2_X1 U1920 ( .A1(n1042), .A2(n1338), .ZN(n1894) );
  OR2_X1 U1921 ( .A1(n1912), .A2(n1913), .ZN(n1899) );
  AND2_X1 U1922 ( .A1(n1884), .A2(n1890), .ZN(n1913) );
  AND2_X1 U1923 ( .A1(n1914), .A2(n1888), .ZN(n1912) );
  OR2_X1 U1924 ( .A1(n1245), .A2(n1338), .ZN(n1888) );
  OR2_X1 U1925 ( .A1(n1890), .A2(n1884), .ZN(n1914) );
  OR2_X1 U1926 ( .A1(n1001), .A2(n1042), .ZN(n1884) );
  INV_X1 U1927 ( .A(a_2_), .ZN(n1042) );
  OR2_X1 U1928 ( .A1(n1915), .A2(n1916), .ZN(n1890) );
  AND2_X1 U1929 ( .A1(n1873), .A2(n1879), .ZN(n1916) );
  AND2_X1 U1930 ( .A1(n1917), .A2(n1877), .ZN(n1915) );
  OR2_X1 U1931 ( .A1(n1001), .A2(n1245), .ZN(n1877) );
  INV_X1 U1932 ( .A(a_3_), .ZN(n1245) );
  OR2_X1 U1933 ( .A1(n1879), .A2(n1873), .ZN(n1917) );
  OR2_X1 U1934 ( .A1(n1210), .A2(n1338), .ZN(n1873) );
  INV_X1 U1935 ( .A(b_0_), .ZN(n1338) );
  OR2_X1 U1936 ( .A1(n1918), .A2(n1919), .ZN(n1879) );
  AND2_X1 U1937 ( .A1(n1861), .A2(n1866), .ZN(n1919) );
  AND2_X1 U1938 ( .A1(n1865), .A2(n1920), .ZN(n1918) );
  OR2_X1 U1939 ( .A1(n1866), .A2(n1861), .ZN(n1920) );
  OR2_X1 U1940 ( .A1(n1001), .A2(n1210), .ZN(n1861) );
  INV_X1 U1941 ( .A(a_4_), .ZN(n1210) );
  INV_X1 U1942 ( .A(n1867), .ZN(n1866) );
  INV_X1 U1943 ( .A(n1868), .ZN(n1865) );
  OR2_X1 U1944 ( .A1(n1921), .A2(n1853), .ZN(n1868) );
  AND2_X1 U1945 ( .A1(n1847), .A2(n1848), .ZN(n1853) );
  AND2_X1 U1946 ( .A1(a_7_), .A2(b_0_), .ZN(n1848) );
  AND2_X1 U1947 ( .A1(n1867), .A2(n1847), .ZN(n1921) );
  INV_X1 U1948 ( .A(n1843), .ZN(n1847) );
  OR2_X1 U1949 ( .A1(n1335), .A2(n1001), .ZN(n1843) );
  INV_X1 U1950 ( .A(b_1_), .ZN(n1001) );
  INV_X1 U1951 ( .A(a_6_), .ZN(n1335) );
  AND2_X1 U1952 ( .A1(a_5_), .A2(b_0_), .ZN(n1867) );
  AND2_X1 U1953 ( .A1(operation_0_), .A2(operation_1_), .ZN(n971) );
endmodule

