module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX646, WX647, n3527, WX648,
         WX649, n3525, WX650, WX652, WX653, n3521, WX654, WX655, n3519, WX656,
         WX657, n3517, WX658, WX659, n3515, WX660, WX661, n3513, WX662, WX663,
         n3511, WX664, WX665, n3509, WX666, WX667, n3507, WX668, WX669, n3505,
         WX670, WX671, n3503, WX672, WX673, n3501, WX674, WX675, n3499, WX676,
         WX677, n3497, WX678, WX679, n3495, WX680, WX681, n3493, WX682, WX683,
         n3491, WX684, WX685, n3489, WX686, WX688, WX689, n3485, WX690, WX691,
         n3483, WX692, WX693, n3481, WX694, WX695, n3479, WX696, WX697, n3477,
         WX698, WX699, n3475, WX700, WX701, n3473, WX702, WX703, n3471, WX704,
         WX705, n3469, WX706, WX707, n3467, WX708, WX709, WX710, WX711, WX712,
         WX713, WX714, WX715, WX716, WX717, WX718, WX719, WX720, WX721, WX722,
         WX724, WX725, WX726, WX727, WX728, WX729, WX730, WX731, WX732, WX733,
         WX734, WX735, WX736, WX737, WX738, WX739, WX740, WX741, WX742, WX743,
         WX744, WX745, WX746, WX747, WX748, WX749, WX750, WX751, WX752, WX753,
         WX754, WX755, WX756, WX757, WX758, WX760, WX761, WX762, WX763, WX764,
         WX765, WX766, WX767, WX768, WX769, WX770, WX771, WX772, WX773, WX774,
         WX775, WX776, WX777, WX778, WX779, WX780, WX781, WX782, WX783, WX784,
         WX785, WX786, WX787, WX788, WX789, WX790, WX791, WX792, WX793, WX794,
         WX796, WX797, WX798, WX799, WX800, WX801, WX802, WX803, WX804, WX805,
         WX806, WX807, WX808, WX809, WX810, WX811, WX812, WX813, WX814, WX815,
         WX816, WX817, WX818, WX819, WX820, WX821, WX822, WX823, WX824, WX825,
         WX826, WX827, WX828, WX829, WX830, WX832, WX833, WX834, WX835, WX836,
         WX837, WX838, WX839, WX840, WX841, WX842, WX843, WX844, WX845, WX846,
         WX847, WX848, WX849, WX850, WX851, WX852, WX853, WX854, WX855, WX856,
         WX857, WX858, WX859, WX860, WX861, WX862, WX863, WX864, WX865, WX866,
         WX868, WX869, WX870, WX871, WX872, WX873, WX874, WX875, WX876, WX877,
         WX878, WX879, WX880, WX881, WX882, WX883, WX884, WX885, WX886, WX887,
         WX888, WX889, WX890, WX891, WX892, WX893, WX894, WX895, WX896, WX897,
         WX898, WX899, WX1264, DFF_160_n1, WX1266, WX1268, DFF_162_n1, WX1270,
         DFF_163_n1, WX1272, DFF_164_n1, WX1274, DFF_165_n1, WX1276,
         DFF_166_n1, WX1278, DFF_167_n1, WX1280, DFF_168_n1, WX1282,
         DFF_169_n1, WX1284, DFF_170_n1, WX1286, DFF_171_n1, WX1288,
         DFF_172_n1, WX1290, DFF_173_n1, WX1292, DFF_174_n1, WX1294,
         DFF_175_n1, WX1296, DFF_176_n1, WX1298, DFF_177_n1, WX1300,
         DFF_178_n1, WX1302, WX1304, DFF_180_n1, WX1306, DFF_181_n1, WX1308,
         DFF_182_n1, WX1310, DFF_183_n1, WX1312, DFF_184_n1, WX1314,
         DFF_185_n1, WX1316, DFF_186_n1, WX1318, DFF_187_n1, WX1320,
         DFF_188_n1, WX1322, DFF_189_n1, WX1324, DFF_190_n1, WX1326,
         DFF_191_n1, WX1778, n8702, n4033, n8701, n4032, n8700, n4031, n8699,
         n4030, n4029, n8696, n4028, n8695, n4027, n8694, n4026, n8693, n4025,
         n8692, n4024, n8691, n4023, n8690, n4022, n8689, n4021, n8688, n4020,
         n8687, n4019, n8686, n4018, n8685, n4017, n8684, n4016, n8683, n4015,
         n8682, n4014, n8681, n4013, n8680, n4012, n4011, n8677, n4010, n8676,
         n4009, n8675, n4008, n8674, n4007, n8673, n4006, n8672, n4005, n8671,
         n4004, WX1839, n8670, n4003, WX1937, n8669, WX1939, n8668, WX1941,
         n8667, WX1943, n8666, WX1945, n8665, WX1947, n8664, WX1949, n8663,
         WX1951, n8662, WX1953, n8661, WX1955, WX1957, n8658, WX1959, n8657,
         WX1961, n8656, WX1963, n8655, WX1965, n8654, WX1967, n8653, WX1969,
         WX1970, WX1971, WX1972, WX1973, WX1974, WX1975, WX1976, WX1977,
         WX1978, WX1979, WX1980, WX1981, WX1982, WX1983, WX1984, WX1985,
         WX1986, WX1987, WX1988, WX1989, WX1990, WX1991, WX1993, WX1994,
         WX1995, WX1996, WX1997, WX1998, WX1999, WX2000, WX2001, WX2002,
         WX2003, WX2004, WX2005, WX2006, WX2007, WX2008, WX2009, WX2010,
         WX2011, WX2012, WX2013, WX2014, WX2015, WX2016, WX2017, WX2018,
         WX2019, WX2020, WX2021, WX2022, WX2023, WX2024, WX2025, WX2026,
         WX2027, WX2029, WX2030, WX2031, WX2032, WX2033, WX2034, WX2035,
         WX2036, WX2037, WX2038, WX2039, WX2040, WX2041, WX2042, WX2043,
         WX2044, WX2045, WX2046, WX2047, WX2048, WX2049, WX2050, WX2051,
         WX2052, WX2053, WX2054, WX2055, WX2056, WX2057, WX2058, WX2059,
         WX2060, WX2061, WX2062, WX2063, WX2065, WX2066, WX2067, WX2068,
         WX2069, WX2070, WX2071, WX2072, WX2073, WX2074, WX2075, WX2076,
         WX2077, WX2078, WX2079, WX2080, WX2081, WX2082, WX2083, WX2084,
         WX2085, WX2086, WX2087, WX2088, WX2089, WX2090, WX2091, WX2092,
         WX2093, WX2094, WX2095, WX2096, WX2097, WX2098, WX2099, WX2101,
         WX2102, WX2103, WX2104, WX2105, WX2106, WX2107, WX2108, WX2109,
         WX2110, WX2111, WX2112, WX2113, WX2114, WX2115, WX2116, WX2117,
         WX2118, WX2119, WX2120, WX2121, WX2122, WX2123, WX2124, WX2125,
         WX2126, WX2127, WX2128, WX2129, WX2130, WX2131, WX2132, WX2133,
         WX2134, WX2135, WX2137, WX2138, WX2139, WX2140, WX2141, WX2142,
         WX2143, WX2144, WX2145, WX2146, WX2147, WX2148, WX2149, WX2150,
         WX2151, WX2152, WX2153, WX2154, WX2155, WX2156, WX2157, WX2158,
         WX2159, WX2160, WX2161, WX2162, WX2163, WX2164, WX2165, WX2166,
         WX2167, WX2168, WX2169, WX2170, WX2171, WX2173, WX2174, WX2175,
         WX2176, WX2177, WX2178, WX2179, WX2180, WX2181, WX2182, WX2183,
         WX2184, WX2185, WX2186, WX2187, WX2188, WX2189, WX2190, WX2191,
         WX2192, WX2557, DFF_352_n1, WX2559, DFF_353_n1, WX2561, DFF_354_n1,
         WX2563, DFF_355_n1, WX2565, DFF_356_n1, WX2567, DFF_357_n1, WX2569,
         DFF_358_n1, WX2571, WX2573, DFF_360_n1, WX2575, DFF_361_n1, WX2577,
         DFF_362_n1, WX2579, DFF_363_n1, WX2581, DFF_364_n1, WX2583,
         DFF_365_n1, WX2585, DFF_366_n1, WX2587, DFF_367_n1, WX2589,
         DFF_368_n1, WX2591, DFF_369_n1, WX2593, DFF_370_n1, WX2595,
         DFF_371_n1, WX2597, DFF_372_n1, WX2599, DFF_373_n1, WX2601,
         DFF_374_n1, WX2603, DFF_375_n1, WX2605, DFF_376_n1, WX2607, WX2609,
         DFF_378_n1, WX2611, DFF_379_n1, WX2613, DFF_380_n1, WX2615,
         DFF_381_n1, WX2617, DFF_382_n1, WX2619, DFF_383_n1, WX3071, n8644,
         n4002, n8643, n4001, n8642, n4000, n8641, n3999, n8640, n3998, n8639,
         n3997, n8638, n3996, n8637, n3995, n8636, n3994, n8635, n3993, n3992,
         n8632, n3991, n8631, n3990, n8630, n3989, n8629, n3988, n8628, n3987,
         n8627, n3986, n8626, n3985, n8625, n3984, n8624, n3983, n8623, n3982,
         n8622, n3981, n8621, n3980, n8620, n3979, n8619, n3978, n8618, n3977,
         n8617, n3976, n8616, n3975, n3974, n8613, n3973, WX3132, n8612, n3972,
         WX3230, n8611, WX3232, n8610, WX3234, n8609, WX3236, n8608, WX3238,
         n8607, WX3240, n8606, WX3242, n8605, WX3244, n8604, WX3246, n8603,
         WX3248, n8602, WX3250, n8601, WX3252, n8600, WX3254, n8599, WX3256,
         n8598, WX3258, n8597, WX3260, WX3262, WX3263, WX3264, WX3265, WX3266,
         WX3267, WX3268, WX3269, WX3270, WX3271, WX3272, WX3273, WX3274,
         WX3275, WX3276, WX3277, WX3278, WX3279, WX3280, WX3281, WX3282,
         WX3283, WX3284, WX3285, WX3286, WX3287, WX3288, WX3289, WX3290,
         WX3291, WX3292, WX3293, WX3294, WX3295, WX3296, WX3298, WX3299,
         WX3300, WX3301, WX3302, WX3303, WX3304, WX3305, WX3306, WX3307,
         WX3308, WX3309, WX3310, WX3311, WX3312, WX3313, WX3314, WX3315,
         WX3316, WX3317, WX3318, WX3319, WX3320, WX3321, WX3322, WX3323,
         WX3324, WX3325, WX3326, WX3327, WX3328, WX3329, WX3330, WX3331,
         WX3332, WX3334, WX3335, WX3336, WX3337, WX3338, WX3339, WX3340,
         WX3341, WX3342, WX3343, WX3344, WX3345, WX3346, WX3347, WX3348,
         WX3349, WX3350, WX3351, WX3352, WX3353, WX3354, WX3355, WX3356,
         WX3357, WX3358, WX3359, WX3360, WX3361, WX3362, WX3363, WX3364,
         WX3365, WX3366, WX3367, WX3368, WX3370, WX3371, WX3372, WX3373,
         WX3374, WX3375, WX3376, WX3377, WX3378, WX3379, WX3380, WX3381,
         WX3382, WX3383, WX3384, WX3385, WX3386, WX3387, WX3388, WX3389,
         WX3390, WX3391, WX3392, WX3393, WX3394, WX3395, WX3396, WX3397,
         WX3398, WX3399, WX3400, WX3401, WX3402, WX3403, WX3404, WX3406,
         WX3407, WX3408, WX3409, WX3410, WX3411, WX3412, WX3413, WX3414,
         WX3415, WX3416, WX3417, WX3418, WX3419, WX3420, WX3421, WX3422,
         WX3423, WX3424, WX3425, WX3426, WX3427, WX3428, WX3429, WX3430,
         WX3431, WX3432, WX3433, WX3434, WX3435, WX3436, WX3437, WX3438,
         WX3440, WX3441, WX3442, WX3443, WX3444, WX3445, WX3446, WX3447,
         WX3448, WX3449, WX3450, WX3451, WX3452, WX3453, WX3454, WX3455,
         WX3456, WX3457, WX3458, WX3459, WX3460, WX3461, WX3462, WX3463,
         WX3464, WX3465, WX3466, WX3467, WX3468, WX3469, WX3470, WX3471,
         WX3472, WX3474, WX3475, WX3476, WX3477, WX3478, WX3479, WX3480,
         WX3481, WX3482, WX3483, WX3484, WX3485, WX3850, DFF_544_n1, WX3852,
         DFF_545_n1, WX3854, DFF_546_n1, WX3856, DFF_547_n1, WX3858,
         DFF_548_n1, WX3860, DFF_549_n1, WX3862, DFF_550_n1, WX3864,
         DFF_551_n1, WX3866, DFF_552_n1, WX3868, DFF_553_n1, WX3870, WX3872,
         DFF_555_n1, WX3874, DFF_556_n1, WX3876, DFF_557_n1, WX3878,
         DFF_558_n1, WX3880, DFF_559_n1, WX3882, DFF_560_n1, WX3884,
         DFF_561_n1, WX3886, DFF_562_n1, WX3888, DFF_563_n1, WX3890,
         DFF_564_n1, WX3892, DFF_565_n1, WX3894, DFF_566_n1, WX3896,
         DFF_567_n1, WX3898, DFF_568_n1, WX3900, DFF_569_n1, WX3902,
         DFF_570_n1, WX3904, WX3906, DFF_572_n1, WX3908, DFF_573_n1, WX3910,
         DFF_574_n1, WX3912, DFF_575_n1, WX4364, n8586, n3971, n8585, n3970,
         n8584, n3969, n8583, n3968, n8582, n3967, n8581, n3966, n8580, n3965,
         n8579, n3964, n8578, n3963, n8577, n3962, n8576, n3961, n3960, n8573,
         n3959, n8572, n3958, n8571, n3957, n8570, n3956, n8569, n3955, n8568,
         n3954, n8567, n3953, n8566, n3952, n8565, n3951, n8564, n3950, n8563,
         n3949, n8562, n3948, n8561, n3947, n8560, n3946, n8559, n3945, n8558,
         n3944, n3943, n8555, n3942, WX4425, n8554, n3941, WX4523, n8553,
         WX4525, n8552, WX4527, n8551, WX4529, n8550, WX4531, n8549, WX4533,
         n8548, WX4535, n8547, WX4537, n8546, WX4539, n8545, WX4541, n8544,
         WX4543, n8543, WX4545, n8542, WX4547, n8541, WX4549, n8540, WX4551,
         WX4553, n8537, WX4555, WX4556, WX4557, WX4558, WX4559, WX4560, WX4561,
         WX4562, WX4563, WX4564, WX4565, WX4566, WX4567, WX4568, WX4569,
         WX4570, WX4571, WX4572, WX4573, WX4574, WX4575, WX4576, WX4577,
         WX4578, WX4579, WX4580, WX4581, WX4582, WX4583, WX4584, WX4585,
         WX4587, WX4588, WX4589, WX4590, WX4591, WX4592, WX4593, WX4594,
         WX4595, WX4596, WX4597, WX4598, WX4599, WX4600, WX4601, WX4602,
         WX4603, WX4604, WX4605, WX4606, WX4607, WX4608, WX4609, WX4610,
         WX4611, WX4612, WX4613, WX4614, WX4615, WX4616, WX4617, WX4618,
         WX4619, WX4621, WX4622, WX4623, WX4624, WX4625, WX4626, WX4627,
         WX4628, WX4629, WX4630, WX4631, WX4632, WX4633, WX4634, WX4635,
         WX4636, WX4637, WX4638, WX4639, WX4640, WX4641, WX4642, WX4643,
         WX4644, WX4645, WX4646, WX4647, WX4648, WX4649, WX4650, WX4651,
         WX4652, WX4653, WX4655, WX4656, WX4657, WX4658, WX4659, WX4660,
         WX4661, WX4662, WX4663, WX4664, WX4665, WX4666, WX4667, WX4668,
         WX4669, WX4670, WX4671, WX4672, WX4673, WX4674, WX4675, WX4676,
         WX4677, WX4678, WX4679, WX4680, WX4681, WX4682, WX4683, WX4684,
         WX4685, WX4686, WX4687, WX4689, WX4690, WX4691, WX4692, WX4693,
         WX4694, WX4695, WX4696, WX4697, WX4698, WX4699, WX4700, WX4701,
         WX4702, WX4703, WX4704, WX4705, WX4706, WX4707, WX4708, WX4709,
         WX4710, WX4711, WX4712, WX4713, WX4714, WX4715, WX4716, WX4717,
         WX4718, WX4719, WX4720, WX4721, WX4723, WX4724, WX4725, WX4726,
         WX4727, WX4728, WX4729, WX4730, WX4731, WX4732, WX4733, WX4734,
         WX4735, WX4736, WX4737, WX4738, WX4739, WX4740, WX4741, WX4742,
         WX4743, WX4744, WX4745, WX4746, WX4747, WX4748, WX4749, WX4750,
         WX4751, WX4752, WX4753, WX4754, WX4755, WX4757, WX4758, WX4759,
         WX4760, WX4761, WX4762, WX4763, WX4764, WX4765, WX4766, WX4767,
         WX4768, WX4769, WX4770, WX4771, WX4772, WX4773, WX4774, WX4775,
         WX4776, WX4777, WX4778, WX5143, DFF_736_n1, WX5145, DFF_737_n1,
         WX5147, DFF_738_n1, WX5149, DFF_739_n1, WX5151, DFF_740_n1, WX5153,
         WX5155, DFF_742_n1, WX5157, DFF_743_n1, WX5159, DFF_744_n1, WX5161,
         DFF_745_n1, WX5163, DFF_746_n1, WX5165, DFF_747_n1, WX5167,
         DFF_748_n1, WX5169, DFF_749_n1, WX5171, DFF_750_n1, WX5173,
         DFF_751_n1, WX5175, DFF_752_n1, WX5177, DFF_753_n1, WX5179,
         DFF_754_n1, WX5181, DFF_755_n1, WX5183, DFF_756_n1, WX5185,
         DFF_757_n1, WX5187, WX5189, DFF_759_n1, WX5191, DFF_760_n1, WX5193,
         DFF_761_n1, WX5195, DFF_762_n1, WX5197, DFF_763_n1, WX5199,
         DFF_764_n1, WX5201, DFF_765_n1, WX5203, DFF_766_n1, WX5205,
         DFF_767_n1, WX5657, n8528, n3940, n8527, n3939, n8526, n3938, n8525,
         n3937, n8524, n3936, n8523, n3935, n3934, n8520, n3933, n8519, n3932,
         n8518, n3931, n8517, n3930, n8516, n3929, n8515, n3928, n8514, n3927,
         n8513, n3926, n8512, n3925, n8511, n3924, n8510, n3923, n8509, n3922,
         n8508, n3921, n8507, n3920, n8506, n3919, n8505, n3918, n3917, n8502,
         n3916, n8501, n3915, n8500, n3914, n8499, n3913, n8498, n3912, n8497,
         n3911, WX5718, n8496, n3910, WX5816, n8495, WX5818, n8494, WX5820,
         n8493, WX5822, n8492, WX5824, n8491, WX5826, n8490, WX5828, n8489,
         WX5830, n8488, WX5832, n8487, WX5834, WX5836, n8484, WX5838, n8483,
         WX5840, n8482, WX5842, n8481, WX5844, n8480, WX5846, n8479, WX5848,
         WX5849, WX5850, WX5851, WX5852, WX5853, WX5854, WX5855, WX5856,
         WX5857, WX5858, WX5859, WX5860, WX5861, WX5862, WX5863, WX5864,
         WX5865, WX5866, WX5867, WX5868, WX5870, WX5871, WX5872, WX5873,
         WX5874, WX5875, WX5876, WX5877, WX5878, WX5879, WX5880, WX5881,
         WX5882, WX5883, WX5884, WX5885, WX5886, WX5887, WX5888, WX5889,
         WX5890, WX5891, WX5892, WX5893, WX5894, WX5895, WX5896, WX5897,
         WX5898, WX5899, WX5900, WX5901, WX5902, WX5904, WX5905, WX5906,
         WX5907, WX5908, WX5909, WX5910, WX5911, WX5912, WX5913, WX5914,
         WX5915, WX5916, WX5917, WX5918, WX5919, WX5920, WX5921, WX5922,
         WX5923, WX5924, WX5925, WX5926, WX5927, WX5928, WX5929, WX5930,
         WX5931, WX5932, WX5933, WX5934, WX5935, WX5936, WX5938, WX5939,
         WX5940, WX5941, WX5942, WX5943, WX5944, WX5945, WX5946, WX5947,
         WX5948, WX5949, WX5950, WX5951, WX5952, WX5953, WX5954, WX5955,
         WX5956, WX5957, WX5958, WX5959, WX5960, WX5961, WX5962, WX5963,
         WX5964, WX5965, WX5966, WX5967, WX5968, WX5969, WX5970, WX5972,
         WX5973, WX5974, WX5975, WX5976, WX5977, WX5978, WX5979, WX5980,
         WX5981, WX5982, WX5983, WX5984, WX5985, WX5986, WX5987, WX5988,
         WX5989, WX5990, WX5991, WX5992, WX5993, WX5994, WX5995, WX5996,
         WX5997, WX5998, WX5999, WX6000, WX6001, WX6002, WX6003, WX6004,
         WX6006, WX6007, WX6008, WX6009, WX6010, WX6011, WX6012, WX6013,
         WX6014, WX6015, WX6016, WX6017, WX6018, WX6019, WX6020, WX6021,
         WX6022, WX6023, WX6024, WX6025, WX6026, WX6027, WX6028, WX6029,
         WX6030, WX6031, WX6032, WX6033, WX6034, WX6035, WX6036, WX6037,
         WX6038, WX6040, WX6041, WX6042, WX6043, WX6044, WX6045, WX6046,
         WX6047, WX6048, WX6049, WX6050, WX6051, WX6052, WX6053, WX6054,
         WX6055, WX6056, WX6057, WX6058, WX6059, WX6060, WX6061, WX6062,
         WX6063, WX6064, WX6065, WX6066, WX6067, WX6068, WX6069, WX6070,
         WX6071, WX6436, WX6438, DFF_929_n1, WX6440, DFF_930_n1, WX6442,
         DFF_931_n1, WX6444, DFF_932_n1, WX6446, DFF_933_n1, WX6448,
         DFF_934_n1, WX6450, DFF_935_n1, WX6452, DFF_936_n1, WX6454,
         DFF_937_n1, WX6456, DFF_938_n1, WX6458, DFF_939_n1, WX6460,
         DFF_940_n1, WX6462, DFF_941_n1, WX6464, DFF_942_n1, WX6466,
         DFF_943_n1, WX6468, DFF_944_n1, WX6470, WX6472, DFF_946_n1, WX6474,
         DFF_947_n1, WX6476, DFF_948_n1, WX6478, DFF_949_n1, WX6480,
         DFF_950_n1, WX6482, DFF_951_n1, WX6484, DFF_952_n1, WX6486,
         DFF_953_n1, WX6488, DFF_954_n1, WX6490, DFF_955_n1, WX6492,
         DFF_956_n1, WX6494, DFF_957_n1, WX6496, DFF_958_n1, WX6498,
         DFF_959_n1, WX6950, n8470, n3909, n3908, n8467, n3907, n8466, n3906,
         n8465, n3905, n8464, n3904, n8463, n3903, n8462, n3902, n8461, n3901,
         n8460, n3900, n8459, n3899, n8458, n3898, n8457, n3897, n8456, n3896,
         n8455, n3895, n8454, n3894, n8453, n3893, n8452, n3892, n3891, n8449,
         n3890, n8448, n3889, n8447, n3888, n8446, n3887, n8445, n3886, n8444,
         n3885, n8443, n3884, n8442, n3883, n8441, n3882, n8440, n3881, n8439,
         n3880, WX7011, n8438, n3879, WX7109, n8437, WX7111, n8436, WX7113,
         n8435, WX7115, n8434, WX7117, WX7119, n8431, WX7121, n8430, WX7123,
         n8429, WX7125, n8428, WX7127, n8427, WX7129, n8426, WX7131, n8425,
         WX7133, n8424, WX7135, n8423, WX7137, n8422, WX7139, n8421, WX7141,
         WX7142, WX7143, WX7144, WX7145, WX7146, WX7147, WX7148, WX7149,
         WX7150, WX7151, WX7153, WX7154, WX7155, WX7156, WX7157, WX7158,
         WX7159, WX7160, WX7161, WX7162, WX7163, WX7164, WX7165, WX7166,
         WX7167, WX7168, WX7169, WX7170, WX7171, WX7172, WX7173, WX7174,
         WX7175, WX7176, WX7177, WX7178, WX7179, WX7180, WX7181, WX7182,
         WX7183, WX7184, WX7185, WX7187, WX7188, WX7189, WX7190, WX7191,
         WX7192, WX7193, WX7194, WX7195, WX7196, WX7197, WX7198, WX7199,
         WX7200, WX7201, WX7202, WX7203, WX7204, WX7205, WX7206, WX7207,
         WX7208, WX7209, WX7210, WX7211, WX7212, WX7213, WX7214, WX7215,
         WX7216, WX7217, WX7218, WX7219, WX7221, WX7222, WX7223, WX7224,
         WX7225, WX7226, WX7227, WX7228, WX7229, WX7230, WX7231, WX7232,
         WX7233, WX7234, WX7235, WX7236, WX7237, WX7238, WX7239, WX7240,
         WX7241, WX7242, WX7243, WX7244, WX7245, WX7246, WX7247, WX7248,
         WX7249, WX7250, WX7251, WX7252, WX7253, WX7255, WX7256, WX7257,
         WX7258, WX7259, WX7260, WX7261, WX7262, WX7263, WX7264, WX7265,
         WX7266, WX7267, WX7268, WX7269, WX7270, WX7271, WX7272, WX7273,
         WX7274, WX7275, WX7276, WX7277, WX7278, WX7279, WX7280, WX7281,
         WX7282, WX7283, WX7284, WX7285, WX7286, WX7287, WX7289, WX7290,
         WX7291, WX7292, WX7293, WX7294, WX7295, WX7296, WX7297, WX7298,
         WX7299, WX7300, WX7301, WX7302, WX7303, WX7304, WX7305, WX7306,
         WX7307, WX7308, WX7309, WX7310, WX7311, WX7312, WX7313, WX7314,
         WX7315, WX7316, WX7317, WX7318, WX7319, WX7320, WX7321, WX7323,
         WX7324, WX7325, WX7326, WX7327, WX7328, WX7329, WX7330, WX7331,
         WX7332, WX7333, WX7334, WX7335, WX7336, WX7337, WX7338, WX7339,
         WX7340, WX7341, WX7342, WX7343, WX7344, WX7345, WX7346, WX7347,
         WX7348, WX7349, WX7350, WX7351, WX7352, WX7353, WX7354, WX7355,
         WX7357, WX7358, WX7359, WX7360, WX7361, WX7362, WX7363, WX7364,
         WX7729, DFF_1120_n1, WX7731, DFF_1121_n1, WX7733, DFF_1122_n1, WX7735,
         DFF_1123_n1, WX7737, DFF_1124_n1, WX7739, DFF_1125_n1, WX7741,
         DFF_1126_n1, WX7743, DFF_1127_n1, WX7745, DFF_1128_n1, WX7747,
         DFF_1129_n1, WX7749, DFF_1130_n1, WX7751, DFF_1131_n1, WX7753, WX7755,
         DFF_1133_n1, WX7757, DFF_1134_n1, WX7759, DFF_1135_n1, WX7761,
         DFF_1136_n1, WX7763, DFF_1137_n1, WX7765, DFF_1138_n1, WX7767,
         DFF_1139_n1, WX7769, DFF_1140_n1, WX7771, DFF_1141_n1, WX7773,
         DFF_1142_n1, WX7775, DFF_1143_n1, WX7777, DFF_1144_n1, WX7779,
         DFF_1145_n1, WX7781, DFF_1146_n1, WX7783, DFF_1147_n1, WX7785,
         DFF_1148_n1, WX7787, WX7789, DFF_1150_n1, WX7791, DFF_1151_n1, WX8243,
         n8411, n3878, n8410, n3877, n8409, n3876, n8408, n3875, n8407, n3874,
         n8406, n3873, n8405, n3872, n8404, n3871, n8403, n3870, n8402, n3869,
         n8401, n3868, n8400, n3867, n8399, n3866, n3865, n8396, n3864, n8395,
         n3863, n8394, n3862, n8393, n3861, n8392, n3860, n8391, n3859, n8390,
         n3858, n8389, n3857, n8388, n3856, n8387, n3855, n8386, n3854, n8385,
         n3853, n8384, n3852, n8383, n3851, n8382, n3850, n8381, n3849, WX8304,
         n3848, WX8402, n8378, WX8404, n8377, WX8406, n8376, WX8408, n8375,
         WX8410, n8374, WX8412, n8373, WX8414, n8372, WX8416, n8371, WX8418,
         n8370, WX8420, n8369, WX8422, n8368, WX8424, n8367, WX8426, n8366,
         WX8428, n8365, WX8430, n8364, WX8432, n8363, WX8434, WX8436, WX8437,
         WX8438, WX8439, WX8440, WX8441, WX8442, WX8443, WX8444, WX8445,
         WX8446, WX8447, WX8448, WX8449, WX8450, WX8451, WX8452, WX8453,
         WX8454, WX8455, WX8456, WX8457, WX8458, WX8459, WX8460, WX8461,
         WX8462, WX8463, WX8464, WX8465, WX8466, WX8467, WX8468, WX8470,
         WX8471, WX8472, WX8473, WX8474, WX8475, WX8476, WX8477, WX8478,
         WX8479, WX8480, WX8481, WX8482, WX8483, WX8484, WX8485, WX8486,
         WX8487, WX8488, WX8489, WX8490, WX8491, WX8492, WX8493, WX8494,
         WX8495, WX8496, WX8497, WX8498, WX8499, WX8500, WX8501, WX8502,
         WX8504, WX8505, WX8506, WX8507, WX8508, WX8509, WX8510, WX8511,
         WX8512, WX8513, WX8514, WX8515, WX8516, WX8517, WX8518, WX8519,
         WX8520, WX8521, WX8522, WX8523, WX8524, WX8525, WX8526, WX8527,
         WX8528, WX8529, WX8530, WX8531, WX8532, WX8533, WX8534, WX8535,
         WX8536, WX8538, WX8539, WX8540, WX8541, WX8542, WX8543, WX8544,
         WX8545, WX8546, WX8547, WX8548, WX8549, WX8550, WX8551, WX8552,
         WX8553, WX8554, WX8555, WX8556, WX8557, WX8558, WX8559, WX8560,
         WX8561, WX8562, WX8563, WX8564, WX8565, WX8566, WX8567, WX8568,
         WX8569, WX8570, WX8572, WX8573, WX8574, WX8575, WX8576, WX8577,
         WX8578, WX8579, WX8580, WX8581, WX8582, WX8583, WX8584, WX8585,
         WX8586, WX8587, WX8588, WX8589, WX8590, WX8591, WX8592, WX8593,
         WX8594, WX8595, WX8596, WX8597, WX8598, WX8599, WX8600, WX8601,
         WX8602, WX8603, WX8604, WX8606, WX8607, WX8608, WX8609, WX8610,
         WX8611, WX8612, WX8613, WX8614, WX8615, WX8616, WX8617, WX8618,
         WX8619, WX8620, WX8621, WX8622, WX8623, WX8624, WX8625, WX8626,
         WX8627, WX8628, WX8629, WX8630, WX8631, WX8632, WX8633, WX8634,
         WX8635, WX8636, WX8637, WX8638, WX8640, WX8641, WX8642, WX8643,
         WX8644, WX8645, WX8646, WX8647, WX8648, WX8649, WX8650, WX8651,
         WX8652, WX8653, WX8654, WX8655, WX8656, WX8657, WX9022, DFF_1312_n1,
         WX9024, DFF_1313_n1, WX9026, DFF_1314_n1, WX9028, DFF_1315_n1, WX9030,
         DFF_1316_n1, WX9032, DFF_1317_n1, WX9034, DFF_1318_n1, WX9036, WX9038,
         DFF_1320_n1, WX9040, DFF_1321_n1, WX9042, DFF_1322_n1, WX9044,
         DFF_1323_n1, WX9046, DFF_1324_n1, WX9048, DFF_1325_n1, WX9050,
         DFF_1326_n1, WX9052, DFF_1327_n1, WX9054, DFF_1328_n1, WX9056,
         DFF_1329_n1, WX9058, DFF_1330_n1, WX9060, DFF_1331_n1, WX9062,
         DFF_1332_n1, WX9064, DFF_1333_n1, WX9066, DFF_1334_n1, WX9068,
         DFF_1335_n1, WX9070, WX9072, DFF_1337_n1, WX9074, DFF_1338_n1, WX9076,
         DFF_1339_n1, WX9078, DFF_1340_n1, WX9080, DFF_1341_n1, WX9082,
         DFF_1342_n1, WX9084, DFF_1343_n1, WX9536, n8353, n3847, n8352, n3846,
         n8351, n3845, n8350, n3844, n8349, n3843, n8348, n3842, n8347, n3841,
         n8346, n3840, n3839, n8343, n3838, n8342, n3837, n8341, n3836, n8340,
         n3835, n8339, n3834, n8338, n3833, n8337, n3832, n8336, n3831, n8335,
         n3830, n8334, n3829, n8333, n3828, n8332, n3827, n8331, n3826, n8330,
         n3825, n8329, n3824, n8328, n3823, n3822, n8325, n3821, n8324, n3820,
         n8323, n3819, n8322, n3818, WX9597, n8321, n3817, WX9695, n8320,
         WX9697, n8319, WX9699, n8318, WX9701, n8317, WX9703, n8316, WX9705,
         n8315, WX9707, n8314, WX9709, n8313, WX9711, n8312, WX9713, n8311,
         WX9715, n8310, WX9717, WX9719, n8307, WX9721, n8306, WX9723, n8305,
         WX9725, n8304, WX9727, WX9728, WX9729, WX9730, WX9731, WX9732, WX9733,
         WX9734, WX9735, WX9736, WX9737, WX9738, WX9739, WX9740, WX9741,
         WX9742, WX9743, WX9744, WX9745, WX9746, WX9747, WX9748, WX9749,
         WX9750, WX9751, WX9753, WX9754, WX9755, WX9756, WX9757, WX9758,
         WX9759, WX9760, WX9761, WX9762, WX9763, WX9764, WX9765, WX9766,
         WX9767, WX9768, WX9769, WX9770, WX9771, WX9772, WX9773, WX9774,
         WX9775, WX9776, WX9777, WX9778, WX9779, WX9780, WX9781, WX9782,
         WX9783, WX9784, WX9785, WX9787, WX9788, WX9789, WX9790, WX9791,
         WX9792, WX9793, WX9794, WX9795, WX9796, WX9797, WX9798, WX9799,
         WX9800, WX9801, WX9802, WX9803, WX9804, WX9805, WX9806, WX9807,
         WX9808, WX9809, WX9810, WX9811, WX9812, WX9813, WX9814, WX9815,
         WX9816, WX9817, WX9818, WX9819, WX9821, WX9822, WX9823, WX9824,
         WX9825, WX9826, WX9827, WX9828, WX9829, WX9830, WX9831, WX9832,
         WX9833, WX9834, WX9835, WX9836, WX9837, WX9838, WX9839, WX9840,
         WX9841, WX9842, WX9843, WX9844, WX9845, WX9846, WX9847, WX9848,
         WX9849, WX9850, WX9851, WX9852, WX9853, WX9855, WX9856, WX9857,
         WX9858, WX9859, WX9860, WX9861, WX9862, WX9863, WX9864, WX9865,
         WX9866, WX9867, WX9868, WX9869, WX9870, WX9871, WX9872, WX9873,
         WX9874, WX9875, WX9876, WX9877, WX9878, WX9879, WX9880, WX9881,
         WX9882, WX9883, WX9884, WX9885, WX9886, WX9887, WX9889, WX9890,
         WX9891, WX9892, WX9893, WX9894, WX9895, WX9896, WX9897, WX9898,
         WX9899, WX9900, WX9901, WX9902, WX9903, WX9904, WX9905, WX9906,
         WX9907, WX9908, WX9909, WX9910, WX9911, WX9912, WX9913, WX9914,
         WX9915, WX9916, WX9917, WX9918, WX9919, WX9920, WX9921, WX9923,
         WX9924, WX9925, WX9926, WX9927, WX9928, WX9929, WX9930, WX9931,
         WX9932, WX9933, WX9934, WX9935, WX9936, WX9937, WX9938, WX9939,
         WX9940, WX9941, WX9942, WX9943, WX9944, WX9945, WX9946, WX9947,
         WX9948, WX9949, WX9950, WX10315, DFF_1504_n1, WX10317, DFF_1505_n1,
         WX10319, WX10321, DFF_1507_n1, WX10323, DFF_1508_n1, WX10325,
         DFF_1509_n1, WX10327, DFF_1510_n1, WX10329, DFF_1511_n1, WX10331,
         DFF_1512_n1, WX10333, DFF_1513_n1, WX10335, DFF_1514_n1, WX10337,
         DFF_1515_n1, WX10339, DFF_1516_n1, WX10341, DFF_1517_n1, WX10343,
         DFF_1518_n1, WX10345, DFF_1519_n1, WX10347, DFF_1520_n1, WX10349,
         DFF_1521_n1, WX10351, DFF_1522_n1, WX10353, WX10355, DFF_1524_n1,
         WX10357, DFF_1525_n1, WX10359, DFF_1526_n1, WX10361, DFF_1527_n1,
         WX10363, DFF_1528_n1, WX10365, DFF_1529_n1, WX10367, DFF_1530_n1,
         WX10369, DFF_1531_n1, WX10371, DFF_1532_n1, WX10373, DFF_1533_n1,
         WX10375, DFF_1534_n1, WX10377, DFF_1535_n1, WX10829, n8295, n3816,
         n8294, n3815, n8293, n3814, n3813, n8290, n3812, n8289, n3811, n8288,
         n3810, n8287, n3809, n8286, n3808, n8285, n3807, n8284, n3806, n8283,
         n3805, n8282, n3804, n8281, n3803, n8280, n3802, n8279, n3801, n8278,
         n3800, n8277, n3799, n8276, n3798, n8275, n3797, n3796, n8272, n3795,
         n8271, n3794, n8270, n3793, n8269, n3792, n8268, n3791, n8267, n3790,
         n8266, n3789, n8265, n3788, n8264, n3787, WX10890, n8263, n3786,
         WX10988, n8262, WX10990, n8261, WX10992, n8260, WX10994, n8259,
         WX10996, n8258, WX10998, n8257, WX11000, WX11002, n8254, WX11004,
         n8253, WX11006, n8252, WX11008, n8251, WX11010, n8250, WX11012, n8249,
         WX11014, n8248, WX11016, n8247, WX11018, n8246, WX11020, WX11021,
         WX11022, WX11023, WX11024, WX11025, WX11026, WX11027, WX11028,
         WX11029, WX11030, WX11031, WX11032, WX11033, WX11034, WX11036,
         WX11037, WX11038, WX11039, WX11040, WX11041, WX11042, WX11043,
         WX11044, WX11045, WX11046, WX11047, WX11048, WX11049, WX11050,
         WX11051, WX11052, WX11053, WX11054, WX11055, WX11056, WX11057,
         WX11058, WX11059, WX11060, WX11061, WX11062, WX11063, WX11064,
         WX11065, WX11066, WX11067, WX11068, WX11070, WX11071, WX11072,
         WX11073, WX11074, WX11075, WX11076, WX11077, WX11078, WX11079,
         WX11080, WX11081, WX11082, WX11083, WX11084, WX11085, WX11086,
         WX11087, WX11088, WX11089, WX11090, WX11091, WX11092, WX11093,
         WX11094, WX11095, WX11096, WX11097, WX11098, WX11099, WX11100,
         WX11101, WX11102, WX11104, WX11105, WX11106, WX11107, WX11108,
         WX11109, WX11110, WX11111, WX11112, WX11113, WX11114, WX11115,
         WX11116, WX11117, WX11118, WX11119, WX11120, WX11121, WX11122,
         WX11123, WX11124, WX11125, WX11126, WX11127, WX11128, WX11129,
         WX11130, WX11131, WX11132, WX11133, WX11134, WX11135, WX11136,
         WX11138, WX11139, WX11140, WX11141, WX11142, WX11143, WX11144,
         WX11145, WX11146, WX11147, WX11148, WX11149, WX11150, WX11151,
         WX11152, WX11153, WX11154, WX11155, WX11156, WX11157, WX11158,
         WX11159, WX11160, WX11161, WX11162, WX11163, WX11164, WX11165,
         WX11166, WX11167, WX11168, WX11169, WX11170, WX11172, WX11173,
         WX11174, WX11175, WX11176, WX11177, WX11178, WX11179, WX11180,
         WX11181, WX11182, WX11183, WX11184, WX11185, WX11186, WX11187,
         WX11188, WX11189, WX11190, WX11191, WX11192, WX11193, WX11194,
         WX11195, WX11196, WX11197, WX11198, WX11199, WX11200, WX11201,
         WX11202, WX11203, WX11204, WX11206, WX11207, WX11208, WX11209,
         WX11210, WX11211, WX11212, WX11213, WX11214, WX11215, WX11216,
         WX11217, WX11218, WX11219, WX11220, WX11221, WX11222, WX11223,
         WX11224, WX11225, WX11226, WX11227, WX11228, WX11229, WX11230,
         WX11231, WX11232, WX11233, WX11234, WX11235, WX11236, WX11237,
         WX11238, WX11240, WX11241, WX11242, WX11243, WX11608, DFF_1696_n1,
         WX11610, DFF_1697_n1, WX11612, DFF_1698_n1, WX11614, DFF_1699_n1,
         WX11616, DFF_1700_n1, WX11618, DFF_1701_n1, WX11620, DFF_1702_n1,
         WX11622, DFF_1703_n1, WX11624, DFF_1704_n1, WX11626, DFF_1705_n1,
         WX11628, DFF_1706_n1, WX11630, DFF_1707_n1, WX11632, DFF_1708_n1,
         WX11634, DFF_1709_n1, WX11636, WX11638, DFF_1711_n1, WX11640,
         DFF_1712_n1, WX11642, DFF_1713_n1, WX11644, DFF_1714_n1, WX11646,
         DFF_1715_n1, WX11648, DFF_1716_n1, WX11650, DFF_1717_n1, WX11652,
         DFF_1718_n1, WX11654, DFF_1719_n1, WX11656, DFF_1720_n1, WX11658,
         DFF_1721_n1, WX11660, DFF_1722_n1, WX11662, DFF_1723_n1, WX11664,
         DFF_1724_n1, WX11666, DFF_1725_n1, WX11668, DFF_1726_n1, WX11670,
         n2245, n2153, n3278, n2152, n2148, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4,
         Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         Tj_Trigger, Stage4, Stage1_1, Stage1_2, Stage1_3, Stage1_4, Stage1,
         Stage2_i, Stage2_7, Stage2_8, Stage2_9, Stage2_10, Stage2, Stage3_i,
         Stage3_12, Stage3_13, Stage3_14, Stage3_15, Stage4_i, Stage4_17,
         Stage4_18, Stage4_19, Stage4_20, Stage4_21, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n2199, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8245, n8255, n8256, n8273, n8274, n8291, n8292, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8308, n8309, n8326, n8327, n8344,
         n8345, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8379, n8380, n8397, n8398, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8432, n8433, n8450, n8451, n8468, n8469, n8471,
         n8472, n8473, n8475, n8476, n8477, n8478, n8485, n8486, n8503, n8504,
         n8521, n8522, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8538, n8539, n8556, n8557, n8574, n8575, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8596, n8614, n8615, n8633, n8634, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8659, n8660, n8678, n8679,
         n8697, n8698, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, U3558_n1, U3871_n1, U3991_n1,
         U5716_n1, U5717_n1, U5718_n1, U5719_n1, U5720_n1, U5721_n1, U5722_n1,
         U5723_n1, U5724_n1, U5725_n1, U5726_n1, U5727_n1, U5728_n1, U5729_n1,
         U5730_n1, U5731_n1, U5732_n1, U5733_n1, U5734_n1, U5735_n1, U5736_n1,
         U5737_n1, U5738_n1, U5739_n1, U5740_n1, U5741_n1, U5742_n1, U5743_n1,
         U5744_n1, U5745_n1, U5746_n1, U5747_n1, U5748_n1, U5749_n1, U5750_n1,
         U5751_n1, U5752_n1, U5753_n1, U5754_n1, U5755_n1, U5756_n1, U5757_n1,
         U5758_n1, U5759_n1, U5760_n1, U5761_n1, U5762_n1, U5763_n1, U5764_n1,
         U5765_n1, U5766_n1, U5767_n1, U5768_n1, U5769_n1, U5770_n1, U5771_n1,
         U5772_n1, U5773_n1, U5774_n1, U5775_n1, U5776_n1, U5777_n1, U5778_n1,
         U5779_n1, U5780_n1, U5781_n1, U5782_n1, U5783_n1, U5784_n1, U5785_n1,
         U5786_n1, U5787_n1, U5788_n1, U5789_n1, U5790_n1, U5791_n1, U5792_n1,
         U5793_n1, U5794_n1, U5795_n1, U5796_n1, U5797_n1, U5798_n1, U5799_n1,
         U5800_n1, U5801_n1, U5802_n1, U5803_n1, U5804_n1, U5805_n1, U5806_n1,
         U5807_n1, U5808_n1, U5809_n1, U5810_n1, U5811_n1, U5812_n1, U5813_n1,
         U5814_n1, U5815_n1, U5816_n1, U5817_n1, U5818_n1, U5819_n1, U5820_n1,
         U5821_n1, U5822_n1, U5823_n1, U5824_n1, U5825_n1, U5826_n1, U5827_n1,
         U5828_n1, U5829_n1, U5830_n1, U5831_n1, U5832_n1, U5833_n1, U5834_n1,
         U5835_n1, U5836_n1, U5837_n1, U5838_n1, U5839_n1, U5840_n1, U5841_n1,
         U5842_n1, U5843_n1, U5844_n1, U5845_n1, U5846_n1, U5847_n1, U5848_n1,
         U5849_n1, U5850_n1, U5851_n1, U5852_n1, U5853_n1, U5854_n1, U5855_n1,
         U5856_n1, U5857_n1, U5858_n1, U5859_n1, U5860_n1, U5861_n1, U5862_n1,
         U5863_n1, U5864_n1, U5865_n1, U5866_n1, U5867_n1, U5868_n1, U5869_n1,
         U5870_n1, U5871_n1, U5872_n1, U5873_n1, U5874_n1, U5875_n1, U5876_n1,
         U5877_n1, U5878_n1, U5879_n1, U5880_n1, U5881_n1, U5882_n1, U5883_n1,
         U5884_n1, U5885_n1, U5886_n1, U5887_n1, U5888_n1, U5889_n1, U5890_n1,
         U5891_n1, U5892_n1, U5893_n1, U5894_n1, U5895_n1, U5896_n1, U5897_n1,
         U5898_n1, U5899_n1, U5900_n1, U5901_n1, U5902_n1, U5903_n1, U5904_n1,
         U5905_n1, U5906_n1, U5907_n1, U5908_n1, U5909_n1, U5910_n1, U5911_n1,
         U5912_n1, U5913_n1, U5914_n1, U5915_n1, U5916_n1, U5917_n1, U5918_n1,
         U5919_n1, U5920_n1, U5921_n1, U5922_n1, U5923_n1, U5924_n1, U5925_n1,
         U5926_n1, U5927_n1, U5928_n1, U5929_n1, U5930_n1, U5931_n1, U5932_n1,
         U5933_n1, U5934_n1, U5935_n1, U5936_n1, U5937_n1, U5938_n1, U5939_n1,
         U5940_n1, U5941_n1, U5942_n1, U5943_n1, U5944_n1, U5945_n1, U5946_n1,
         U5947_n1, U5948_n1, U5949_n1, U5950_n1, U5951_n1, U5952_n1, U5953_n1,
         U5954_n1, U5955_n1, U5956_n1, U5957_n1, U5958_n1, U5959_n1, U5960_n1,
         U5961_n1, U5962_n1, U5963_n1, U5964_n1, U5965_n1, U5966_n1, U5967_n1,
         U5968_n1, U5969_n1, U5970_n1, U5971_n1, U5972_n1, U5973_n1, U5974_n1,
         U5975_n1, U5976_n1, U5977_n1, U5978_n1, U5979_n1, U5980_n1, U5981_n1,
         U5982_n1, U5983_n1, U5984_n1, U5985_n1, U5986_n1, U5987_n1, U5988_n1,
         U5989_n1, U5990_n1, U5991_n1, U5992_n1, U5993_n1, U5994_n1, U5995_n1,
         U5996_n1, U5997_n1, U5998_n1, U5999_n1, U6000_n1, U6001_n1, U6002_n1,
         U6003_n1, U6004_n1, U6005_n1, U6006_n1, U6007_n1, U6008_n1, U6009_n1,
         U6010_n1, U6011_n1, U6012_n1, U6013_n1, U6014_n1, U6015_n1, U6016_n1,
         U6017_n1, U6018_n1, U6019_n1, U6020_n1, U6021_n1, U6022_n1, U6023_n1,
         U6024_n1, U6025_n1, U6026_n1, U6027_n1, U6028_n1, U6029_n1, U6030_n1,
         U6031_n1, U6032_n1, U6033_n1, U6034_n1, U6035_n1, U6036_n1, U6037_n1,
         U6038_n1, U6039_n1, U6040_n1, U6041_n1, U6042_n1, U6043_n1, U6044_n1,
         U6045_n1, U6046_n1, U6047_n1, U6048_n1, U6049_n1, U6050_n1, U6051_n1,
         U6052_n1, U6053_n1, U6054_n1, U6055_n1, U6056_n1, U6057_n1, U6058_n1,
         U6059_n1, U6060_n1, U6061_n1, U6062_n1, U6063_n1, U6064_n1, U6065_n1,
         U6066_n1, U6067_n1, U6068_n1, U6069_n1, U6070_n1, U6071_n1, U6072_n1,
         U6073_n1, U6074_n1, U6075_n1, U6076_n1, U6077_n1, U6078_n1, U6079_n1,
         U6080_n1, U6081_n1, U6082_n1, U6083_n1, U6084_n1, U6085_n1, U6086_n1,
         U6087_n1, U6088_n1, U6089_n1, U6090_n1, U6091_n1, U6092_n1, U6093_n1,
         U6094_n1, U6095_n1, U6096_n1, U6097_n1, U6098_n1, U6099_n1, U6100_n1,
         U6101_n1, U6102_n1, U6103_n1, U6104_n1, U6105_n1, U6106_n1, U6107_n1,
         U6108_n1, U6109_n1, U6110_n1, U6111_n1, U6112_n1, U6113_n1, U6114_n1,
         U6115_n1, U6116_n1, U6117_n1, U6118_n1, U6119_n1, U6120_n1, U6121_n1,
         U6122_n1, U6123_n1, U6124_n1, U6125_n1, U6126_n1, U6127_n1, U6128_n1,
         U6129_n1, U6130_n1, U6131_n1, U6132_n1, U6133_n1, U6134_n1, U6135_n1,
         U6136_n1, U6137_n1, U6138_n1, U6139_n1, U6140_n1, U6141_n1, U6142_n1,
         U6143_n1, U6144_n1, U6145_n1, U6146_n1, U6147_n1, U6148_n1, U6149_n1,
         U6150_n1, U6151_n1, U6152_n1, U6153_n1, U6154_n1, U6155_n1, U6156_n1,
         U6157_n1, U6158_n1, U6159_n1, U6160_n1, U6161_n1, U6162_n1, U6163_n1,
         U6164_n1, U6165_n1, U6166_n1, U6167_n1, U6168_n1, U6169_n1, U6170_n1,
         U6171_n1, U6172_n1, U6173_n1, U6174_n1, U6175_n1, U6176_n1, U6177_n1,
         U6178_n1, U6179_n1, U6180_n1, U6181_n1, U6182_n1, U6183_n1, U6184_n1,
         U6185_n1, U6186_n1, U6187_n1, U6188_n1, U6189_n1, U6190_n1, U6191_n1,
         U6192_n1, U6193_n1, U6194_n1, U6195_n1, U6196_n1, U6197_n1, U6198_n1,
         U6199_n1, U6200_n1, U6201_n1, U6202_n1, U6203_n1, U6204_n1, U6205_n1,
         U6206_n1, U6207_n1, U6208_n1, U6209_n1, U6210_n1, U6211_n1, U6212_n1,
         U6213_n1, U6214_n1, U6215_n1, U6216_n1, U6217_n1, U6218_n1, U6219_n1,
         U6220_n1, U6221_n1, U6222_n1, U6223_n1, U6224_n1, U6225_n1, U6226_n1,
         U6227_n1, U6228_n1, U6229_n1, U6230_n1, U6231_n1, U6232_n1, U6233_n1,
         U6234_n1, U6235_n1, U6236_n1, U6237_n1, U6238_n1, U6239_n1, U6240_n1,
         U6241_n1, U6242_n1, U6243_n1, U6244_n1, U6245_n1, U6246_n1, U6247_n1,
         U6248_n1, U6249_n1, U6250_n1, U6251_n1, U6252_n1, U6253_n1, U6254_n1,
         U6255_n1, U6256_n1, U6257_n1, U6258_n1, U6259_n1, U6260_n1, U6261_n1,
         U6262_n1, U6263_n1, U6264_n1, U6265_n1, U6266_n1, U6267_n1, U6268_n1,
         U6269_n1, U6270_n1, U6271_n1, U6272_n1, U6273_n1, U6274_n1, U6275_n1,
         U6276_n1, U6277_n1, U6278_n1, U6279_n1, U6280_n1, U6281_n1, U6282_n1,
         U6283_n1, U6284_n1, U6285_n1, U6286_n1, U6287_n1, U6288_n1, U6289_n1,
         U6290_n1, U6291_n1, U6292_n1, U6293_n1, U6294_n1, U6295_n1, U6296_n1,
         U6297_n1, U6298_n1, U6299_n1, U6300_n1, U6301_n1, U6302_n1, U6303_n1,
         U6304_n1, U6305_n1, U6306_n1, U6307_n1, U6308_n1, U6309_n1, U6310_n1,
         U6311_n1, U6312_n1, U6313_n1, U6314_n1, U6315_n1, U6316_n1, U6317_n1,
         U6318_n1, U6319_n1, U6320_n1, U6321_n1, U6322_n1, U6323_n1, U6324_n1,
         U6325_n1, U6326_n1, U6327_n1, U6328_n1, U6329_n1, U6330_n1, U6331_n1,
         U6332_n1, U6333_n1, U6334_n1, U6335_n1, U6336_n1, U6337_n1, U6338_n1,
         U6339_n1, U6340_n1, U6341_n1, U6342_n1, U6343_n1, U6344_n1, U6345_n1,
         U6346_n1, U6347_n1, U6348_n1, U6349_n1, U6350_n1, U6351_n1, U6352_n1,
         U6353_n1, U6354_n1, U6355_n1, U6356_n1, U6357_n1, U6358_n1, U6359_n1,
         U6360_n1, U6361_n1, U6362_n1, U6363_n1, U6364_n1, U6365_n1, U6366_n1,
         U6367_n1, U6368_n1, U6369_n1, U6370_n1, U6371_n1, U6372_n1, U6373_n1,
         U6374_n1, U6375_n1, U6376_n1, U6377_n1, U6378_n1, U6379_n1, U6380_n1,
         U6381_n1, U6382_n1, U6383_n1, U6384_n1, U6385_n1, U6386_n1, U6387_n1,
         U6388_n1, U6389_n1, U6390_n1, U6391_n1, U6392_n1, U6393_n1, U6394_n1,
         U6395_n1, U6396_n1, U6397_n1, U6398_n1, U6399_n1, U6400_n1, U6401_n1,
         U6402_n1, U6403_n1, U6404_n1, U6405_n1, U6406_n1, U6407_n1, U6408_n1,
         U6409_n1, U6410_n1, U6411_n1, U6412_n1, U6413_n1, U6414_n1, U6415_n1,
         U6416_n1, U6417_n1, U6418_n1, U6419_n1, U6420_n1, U6421_n1, U6422_n1,
         U6423_n1, U6424_n1, U6425_n1, U6426_n1, U6427_n1, U6428_n1, U6429_n1,
         U6430_n1, U6431_n1, U6432_n1, U6433_n1, U6434_n1, U6435_n1, U6436_n1,
         U6437_n1, U6438_n1, U6439_n1, U6440_n1, U6441_n1, U6442_n1, U6443_n1,
         U6444_n1, U6445_n1, U6446_n1, U6447_n1, U6448_n1, U6449_n1, U6450_n1,
         U6451_n1, U6452_n1, U6453_n1, U6454_n1, U6455_n1, U6456_n1, U6457_n1,
         U6458_n1, U6459_n1, U6460_n1, U6461_n1, U6462_n1, U6463_n1, U6464_n1,
         U6465_n1, U6466_n1, U6467_n1, U6468_n1, U6469_n1, U6470_n1, U6471_n1,
         U6472_n1, U6473_n1, U6474_n1, U6475_n1, U6476_n1, U6477_n1, U6478_n1,
         U6479_n1, U6480_n1, U6481_n1, U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n9289), .CLK(n9633), .Q(
        WX485), .QN(n9078) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n9316), .CLK(n9635), .Q(
        WX487), .QN(n9077) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n9417), .CLK(n9635), .Q(
        WX489), .QN(n9075) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n9297), .CLK(n9635), .Q(
        WX491), .QN(n9074) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n9396), .CLK(n9635), .Q(
        WX493), .QN(n9073) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n9384), .CLK(n9635), .Q(
        WX495), .QN(n9072) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n9381), .CLK(n9635), .Q(
        WX497), .QN(n9071) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n9369), .CLK(n9635), .Q(
        WX499), .QN(n9070) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n9374), .CLK(n9635), .Q(
        WX501), .QN(n9069) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n9288), .CLK(n9634), .Q(
        WX503), .QN(n9068) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n9285), .CLK(n9634), .Q(
        WX505), .QN(n9067) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n9286), .CLK(n9634), .Q(
        WX507), .QN(n9066) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n9289), .CLK(n9634), .Q(
        WX509), .QN(n9064) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n9290), .CLK(n9634), .Q(
        WX511), .QN(n9063) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(test_se), .CLK(n9634), .Q(
        WX513), .QN(n9062) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n9291), .CLK(n9634), .Q(
        WX515), .QN(n9061) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n9287), .CLK(n9634), .Q(
        WX517), .QN(n9060) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n9288), .CLK(n9634), .Q(
        test_so1), .QN(n9059) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n9285), .CLK(n9634), .Q(
        WX521), .QN(n9058) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n9286), .CLK(n9634), .Q(
        WX523), .QN(n9057) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n9289), .CLK(n9634), .Q(
        WX525), .QN(n9056) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(test_se), .CLK(n9633), .Q(
        WX527), .QN(n9055) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n9291), .CLK(n9633), .Q(
        WX529), .QN(n9084) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n9287), .CLK(n9633), .Q(
        WX531), .QN(n9083) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n9288), .CLK(n9633), .Q(
        WX533), .QN(n9082) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n9285), .CLK(n9633), .Q(
        WX535), .QN(n9081) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n9286), .CLK(n9633), .Q(
        WX537), .QN(n9080) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n9289), .CLK(n9633), .Q(
        WX539), .QN(n9079) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n9287), .CLK(n9633), .Q(
        WX541), .QN(n9076) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n9288), .CLK(n9633), .Q(
        WX543), .QN(n9065) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n9285), .CLK(n9633), .Q(
        WX545), .QN(n9054) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n9286), .CLK(n9633), .Q(
        WX547), .QN(n9053) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n9317), .CLK(n9635), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(n9318), .CLK(n9635), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(n9319), .CLK(n9635), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(n9320), .CLK(n9635), .Q(
        test_so2), .QN(n9166) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(n9378), .CLK(n9636), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(n9379), .CLK(n9636), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(n9296), .CLK(n9636), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n9298), .CLK(n9636), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(n9322), .CLK(n9636), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(n9324), .CLK(n9636), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(n9425), .CLK(n9637), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n9425), .CLK(n9637), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(n9425), .CLK(n9637), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(n9425), .CLK(n9637), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(n9425), .CLK(n9637), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n9424), .CLK(n9638), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(n9424), .CLK(n9638), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(n9424), .CLK(n9638), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(n9423), .CLK(n9639), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(n9423), .CLK(n9639), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(n9423), .CLK(n9639), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n9399), .CLK(n9640), .Q(
        test_so3), .QN(n9167) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(n9424), .CLK(n9640), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(n9340), .CLK(n9640), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(n9422), .CLK(n9641), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(n9422), .CLK(n9641), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(n9422), .CLK(n9641), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(n9421), .CLK(n9642), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(n9421), .CLK(n9642), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(n9421), .CLK(n9642), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(n9420), .CLK(n9643), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(n9420), .CLK(n9643), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n9420), .CLK(n9643), .Q(
        WX709), .QN(n9028) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n9419), .CLK(n9644), .Q(
        WX711), .QN(n8954) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n9419), .CLK(n9644), .Q(
        WX713), .QN(n8965) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n9321), .CLK(n9636), .Q(
        WX715), .QN(n8974) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n9397), .CLK(n9636), .Q(
        WX717), .QN(n8980) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n9385), .CLK(n9636), .Q(
        WX719), .QN(n8983) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n9422), .CLK(n9636), .Q(
        WX721), .QN(n8992) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n9423), .CLK(n9636), .Q(
        test_so4), .QN(n9148) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n9323), .CLK(n9636), .Q(
        WX725), .QN(n9003) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n9425), .CLK(n9637), .Q(
        WX727), .QN(n9015) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n9425), .CLK(n9637), .Q(
        WX729), .QN(n9021) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n9425), .CLK(n9637), .Q(
        WX731), .QN(n9027) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n9425), .CLK(n9637), .Q(
        WX733), .QN(n8962) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n9425), .CLK(n9637), .Q(
        WX735), .QN(n8977) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n9424), .CLK(n9638), .Q(
        WX737), .QN(n8989) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n9424), .CLK(n9638), .Q(
        WX739), .QN(n9004) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n9424), .CLK(n9638), .Q(
        WX741), .QN(n9018) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n9424), .CLK(n9638), .Q(
        WX743), .QN(n9033) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n9423), .CLK(n9639), .Q(
        WX745), .QN(n8968) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n9423), .CLK(n9639), .Q(
        WX747), .QN(n8995) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n9423), .CLK(n9639), .Q(
        WX749), .QN(n9041) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n9364), .CLK(n9640), .Q(
        WX751), .QN(n8986) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n9390), .CLK(n9640), .Q(
        WX753), .QN(n8996) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n9341), .CLK(n9640), .Q(
        WX755), .QN(n9008) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n9422), .CLK(n9641), .Q(
        WX757), .QN(n9036) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n9422), .CLK(n9641), .Q(
        test_so5), .QN(n9147) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n9422), .CLK(n9641), .Q(
        WX761), .QN(n9011) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n9421), .CLK(n9642), .Q(
        WX763), .QN(n9014) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n9421), .CLK(n9642), .Q(
        WX765), .QN(n8959) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n9421), .CLK(n9642), .Q(
        WX767), .QN(n9034) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n9420), .CLK(n9643), .Q(
        WX769), .QN(n8970) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n9420), .CLK(n9643), .Q(
        WX771), .QN(n9042) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n9420), .CLK(n9643), .Q(
        WX773), .QN(n9029) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n9419), .CLK(n9644), .Q(
        WX775), .QN(n8955) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n9419), .CLK(n9644), .Q(
        WX777), .QN(n8963) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n9419), .CLK(n9644), .Q(
        WX779), .QN(n8972) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n9419), .CLK(n9644), .Q(
        WX781), .QN(n8978) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n9419), .CLK(n9644), .Q(
        WX783), .QN(n8981) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n9418), .CLK(n9645), .Q(
        WX785), .QN(n8990) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n9418), .CLK(n9645), .Q(
        WX787), .QN(n8999) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n9418), .CLK(n9645), .Q(
        WX789), .QN(n9001) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n9418), .CLK(n9645), .Q(
        WX791), .QN(n9016) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n9418), .CLK(n9645), .Q(
        WX793), .QN(n9022) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n9418), .CLK(n9645), .Q(
        test_so6), .QN(n9098) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n9425), .CLK(n9637), 
        .Q(WX797), .QN(n8960) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n9425), .CLK(n9637), .Q(
        WX799), .QN(n8975) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n9424), .CLK(n9638), .Q(
        WX801), .QN(n8987) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n9424), .CLK(n9638), .Q(
        WX803), .QN(n9005) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n9424), .CLK(n9638), .Q(
        WX805), .QN(n9019) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n9424), .CLK(n9638), .Q(
        WX807), .QN(n9031) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n9423), .CLK(n9639), .Q(
        WX809), .QN(n8966) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n9423), .CLK(n9639), .Q(
        WX811), .QN(n8993) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n9423), .CLK(n9639), .Q(
        WX813), .QN(n9039) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n9370), .CLK(n9640), .Q(
        WX815), .QN(n8984) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n9418), .CLK(n9640), .Q(
        WX817), .QN(n8997) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n9342), .CLK(n9640), .Q(
        WX819), .QN(n9006) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n9422), .CLK(n9641), .Q(
        WX821), .QN(n9037) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n9422), .CLK(n9641), .Q(
        WX823), .QN(n9024) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n9422), .CLK(n9641), .Q(
        WX825), .QN(n9009) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n9421), .CLK(n9642), .Q(
        WX827), .QN(n9012) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n9421), .CLK(n9642), .Q(
        WX829), .QN(n8957) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n9421), .CLK(n9642), .Q(
        test_so7), .QN(n9149) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n9420), .CLK(n9643), 
        .Q(WX833), .QN(n8971) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n9420), .CLK(n9643), .Q(
        WX835), .QN(n9043) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n9420), .CLK(n9643), .Q(
        WX837), .QN(n9030) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n9419), .CLK(n9644), .Q(
        WX839), .QN(n8956) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n9419), .CLK(n9644), .Q(
        WX841), .QN(n8964) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n9419), .CLK(n9644), .Q(
        WX843), .QN(n8973) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n9419), .CLK(n9644), .Q(
        WX845), .QN(n8979) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n9419), .CLK(n9644), .Q(
        WX847), .QN(n8982) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n9418), .CLK(n9645), .Q(
        WX849), .QN(n8991) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n9418), .CLK(n9645), .Q(
        WX851), .QN(n9000) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n9418), .CLK(n9645), .Q(
        WX853), .QN(n9002) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n9418), .CLK(n9645), .Q(
        WX855), .QN(n9017) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n9418), .CLK(n9645), .Q(
        WX857), .QN(n9023) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n9418), .CLK(n9645), .Q(
        WX859), .QN(n9026) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n9417), .CLK(n9646), .Q(
        WX861), .QN(n8961) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n9417), .CLK(n9646), .Q(
        WX863), .QN(n8976) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n9417), .CLK(n9646), .Q(
        WX865), .QN(n8988) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n9417), .CLK(n9646), .Q(
        test_so8), .QN(n9086) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n9424), .CLK(n9638), 
        .Q(WX869), .QN(n9020) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n9423), .CLK(n9639), .Q(
        WX871), .QN(n9032) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n9423), .CLK(n9639), .Q(
        WX873), .QN(n8967) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n9423), .CLK(n9639), .Q(
        WX875), .QN(n8994) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n9368), .CLK(n9640), .Q(
        WX877), .QN(n9040) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n9294), .CLK(n9640), .Q(
        WX879), .QN(n8985) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n9410), .CLK(n9640), .Q(
        WX881), .QN(n8998) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n9422), .CLK(n9641), .Q(
        WX883), .QN(n9007) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n9422), .CLK(n9641), .Q(
        WX885), .QN(n9038) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n9422), .CLK(n9641), .Q(
        WX887), .QN(n9025) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n9421), .CLK(n9642), .Q(
        WX889), .QN(n9010) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n9421), .CLK(n9642), .Q(
        WX891), .QN(n9013) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n9421), .CLK(n9642), .Q(
        WX893), .QN(n8958) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n9420), .CLK(n9643), .Q(
        WX895), .QN(n9035) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n9420), .CLK(n9643), .Q(
        WX897), .QN(n8969) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n9420), .CLK(n9643), .Q(
        WX899), .QN(n9044) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n9293), .CLK(n9775), .Q(
        CRC_OUT_9_0), .QN(DFF_160_n1) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n9293), .CLK(n9775), 
        .Q(test_so9), .QN(n9162) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n9293), .CLK(n9775), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n9293), .CLK(n9775), 
        .Q(CRC_OUT_9_3), .QN(DFF_163_n1) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n9293), .CLK(n9775), 
        .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n9293), .CLK(n9775), 
        .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n9293), .CLK(n9775), 
        .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n9293), .CLK(n9775), 
        .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n9292), .CLK(n9776), 
        .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n9292), .CLK(n9776), 
        .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n9292), .CLK(n9776), 
        .Q(CRC_OUT_9_10), .QN(DFF_170_n1) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n9292), .CLK(n9776), .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n9292), .CLK(n9776), .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n9292), .CLK(n9776), .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n9292), .CLK(n9776), .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n9292), .CLK(n9776), .Q(CRC_OUT_9_15), .QN(DFF_175_n1) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n9292), .CLK(n9776), .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n9292), .CLK(n9776), .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n9292), .CLK(n9776), .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n9292), .CLK(n9776), .Q(test_so10), .QN(n9161) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n9417), .CLK(n9646), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n9417), .CLK(n9646), .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n9417), .CLK(n9646), .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n9417), .CLK(n9646), .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n9417), .CLK(n9646), .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n9417), .CLK(n9646), .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n9417), .CLK(n9646), .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n9417), .CLK(n9646), .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n9287), .CLK(n9647), .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n9291), .CLK(n9647), .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(test_se), .CLK(
        n9647), .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n9290), .CLK(n9647), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n267), .SI(CRC_OUT_9_31), .SE(n9289), .CLK(n9647), 
        .Q(WX1778), .QN(n9045) );
  SDFFX1 DFF_193_Q_reg ( .D(n268), .SI(WX1778), .SE(n9415), .CLK(n9649), .Q(
        n8702), .QN(n4033) );
  SDFFX1 DFF_194_Q_reg ( .D(n269), .SI(n8702), .SE(n9415), .CLK(n9649), .Q(
        n8701), .QN(n4032) );
  SDFFX1 DFF_195_Q_reg ( .D(n270), .SI(n8701), .SE(n9415), .CLK(n9649), .Q(
        n8700), .QN(n4031) );
  SDFFX1 DFF_196_Q_reg ( .D(n271), .SI(n8700), .SE(n9415), .CLK(n9649), .Q(
        n8699), .QN(n4030) );
  SDFFX1 DFF_197_Q_reg ( .D(n272), .SI(n8699), .SE(n9415), .CLK(n9649), .Q(
        test_so11), .QN(n4029) );
  SDFFX1 DFF_198_Q_reg ( .D(n273), .SI(test_si12), .SE(n9415), .CLK(n9649), 
        .Q(n8696), .QN(n4028) );
  SDFFX1 DFF_199_Q_reg ( .D(n274), .SI(n8696), .SE(n9415), .CLK(n9649), .Q(
        n8695), .QN(n4027) );
  SDFFX1 DFF_200_Q_reg ( .D(n275), .SI(n8695), .SE(n9415), .CLK(n9649), .Q(
        n8694), .QN(n4026) );
  SDFFX1 DFF_201_Q_reg ( .D(n276), .SI(n8694), .SE(n9415), .CLK(n9649), .Q(
        n8693), .QN(n4025) );
  SDFFX1 DFF_202_Q_reg ( .D(n277), .SI(n8693), .SE(n9415), .CLK(n9649), .Q(
        n8692), .QN(n4024) );
  SDFFX1 DFF_203_Q_reg ( .D(n278), .SI(n8692), .SE(n9415), .CLK(n9649), .Q(
        n8691), .QN(n4023) );
  SDFFX1 DFF_204_Q_reg ( .D(n279), .SI(n8691), .SE(n9415), .CLK(n9649), .Q(
        n8690), .QN(n4022) );
  SDFFX1 DFF_205_Q_reg ( .D(n280), .SI(n8690), .SE(n9416), .CLK(n9648), .Q(
        n8689), .QN(n4021) );
  SDFFX1 DFF_206_Q_reg ( .D(n281), .SI(n8689), .SE(n9416), .CLK(n9648), .Q(
        n8688), .QN(n4020) );
  SDFFX1 DFF_207_Q_reg ( .D(n282), .SI(n8688), .SE(n9416), .CLK(n9648), .Q(
        n8687), .QN(n4019) );
  SDFFX1 DFF_208_Q_reg ( .D(n283), .SI(n8687), .SE(n9416), .CLK(n9648), .Q(
        n8686), .QN(n4018) );
  SDFFX1 DFF_209_Q_reg ( .D(n284), .SI(n8686), .SE(n9416), .CLK(n9648), .Q(
        n8685), .QN(n4017) );
  SDFFX1 DFF_210_Q_reg ( .D(n285), .SI(n8685), .SE(n9416), .CLK(n9648), .Q(
        n8684), .QN(n4016) );
  SDFFX1 DFF_211_Q_reg ( .D(n286), .SI(n8684), .SE(n9416), .CLK(n9648), .Q(
        n8683), .QN(n4015) );
  SDFFX1 DFF_212_Q_reg ( .D(n287), .SI(n8683), .SE(n9416), .CLK(n9648), .Q(
        n8682), .QN(n4014) );
  SDFFX1 DFF_213_Q_reg ( .D(n288), .SI(n8682), .SE(n9416), .CLK(n9648), .Q(
        n8681), .QN(n4013) );
  SDFFX1 DFF_214_Q_reg ( .D(n289), .SI(n8681), .SE(n9416), .CLK(n9648), .Q(
        n8680), .QN(n4012) );
  SDFFX1 DFF_215_Q_reg ( .D(n290), .SI(n8680), .SE(n9416), .CLK(n9648), .Q(
        test_so12), .QN(n4011) );
  SDFFX1 DFF_216_Q_reg ( .D(n291), .SI(test_si13), .SE(n9416), .CLK(n9648), 
        .Q(n8677), .QN(n4010) );
  SDFFX1 DFF_217_Q_reg ( .D(n292), .SI(n8677), .SE(n9290), .CLK(n9647), .Q(
        n8676), .QN(n4009) );
  SDFFX1 DFF_218_Q_reg ( .D(n293), .SI(n8676), .SE(test_se), .CLK(n9647), .Q(
        n8675), .QN(n4008) );
  SDFFX1 DFF_219_Q_reg ( .D(n294), .SI(n8675), .SE(n9291), .CLK(n9647), .Q(
        n8674), .QN(n4007) );
  SDFFX1 DFF_220_Q_reg ( .D(n295), .SI(n8674), .SE(n9287), .CLK(n9647), .Q(
        n8673), .QN(n4006) );
  SDFFX1 DFF_221_Q_reg ( .D(n296), .SI(n8673), .SE(n9288), .CLK(n9647), .Q(
        n8672), .QN(n4005) );
  SDFFX1 DFF_222_Q_reg ( .D(n297), .SI(n8672), .SE(n9285), .CLK(n9647), .Q(
        n8671), .QN(n4004) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n9286), .CLK(n9647), .Q(
        n8670), .QN(n4003) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n9293), .CLK(n9775), .Q(
        n8669), .QN(n15982) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n9414), .CLK(n9650), .Q(
        n8668), .QN(n15979) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n9414), .CLK(n9650), .Q(
        n8667), .QN(n15977) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n9414), .CLK(n9650), .Q(
        n8666), .QN(n15975) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n9414), .CLK(n9650), .Q(
        n8665), .QN(n15973) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n9414), .CLK(n9650), .Q(
        n8664), .QN(n15971) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n9414), .CLK(n9650), .Q(
        n8663), .QN(n15969) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n9413), .CLK(n9651), .Q(
        n8662), .QN(n15967) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n9413), .CLK(n9651), .Q(
        n8661), .QN(n15965) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n9413), .CLK(n9651), .Q(
        test_so13), .QN(n9096) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n9413), .CLK(n9651), 
        .Q(n8658), .QN(n15962) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n9413), .CLK(n9651), .Q(
        n8657), .QN(n15960) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n9413), .CLK(n9651), .Q(
        n8656), .QN(n15958) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n9412), .CLK(n9652), .Q(
        n8655), .QN(n15956) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n9412), .CLK(n9652), .Q(
        n8654), .QN(n15954) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n9412), .CLK(n9652), .Q(
        n8653), .QN(n15953) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n9412), .CLK(n9652), .Q(
        WX1970), .QN(n8711) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n9411), .CLK(n9653), .Q(
        WX1972), .QN(n8710) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n9411), .CLK(n9653), .Q(
        WX1974), .QN(n8708) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n9411), .CLK(n9653), .Q(
        WX1976), .QN(n8706) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n9411), .CLK(n9653), .Q(
        WX1978), .QN(n8704) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n9410), .CLK(n9654), .Q(
        WX1980), .QN(n8698) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n9410), .CLK(n9654), .Q(
        WX1982), .QN(n8679) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n9410), .CLK(n9654), .Q(
        WX1984), .QN(n8660) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n9410), .CLK(n9654), .Q(
        WX1986), .QN(n8652) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n9409), .CLK(n9655), .Q(
        WX1988), .QN(n8650) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n9409), .CLK(n9655), .Q(
        WX1990), .QN(n8648) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n9409), .CLK(n9655), .Q(
        test_so14), .QN(n9135) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n9408), .CLK(n9656), 
        .Q(WX1994), .QN(n8645) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n9408), .CLK(n9656), .Q(
        WX1996), .QN(n8633) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n9408), .CLK(n9656), .Q(
        WX1998), .QN(n8614) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n9407), .CLK(n9657), .Q(
        WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n9407), .CLK(n9657), .Q(
        WX2002), .QN(n7890) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n9414), .CLK(n9650), .Q(
        WX2004), .QN(n8116) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n9414), .CLK(n9650), .Q(
        WX2006), .QN(n8114) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n9414), .CLK(n9650), .Q(
        WX2008), .QN(n8112) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n9414), .CLK(n9650), .Q(
        WX2010), .QN(n8110) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n9414), .CLK(n9650), .Q(
        WX2012), .QN(n8108) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n9414), .CLK(n9650), .Q(
        WX2014), .QN(n8106) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n9413), .CLK(n9651), .Q(
        WX2016), .QN(n8104) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n9413), .CLK(n9651), .Q(
        WX2018), .QN(n8102) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n9413), .CLK(n9651), .Q(
        WX2020), .QN(n8100) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n9413), .CLK(n9651), .Q(
        WX2022), .QN(n8098) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n9413), .CLK(n9651), .Q(
        WX2024), .QN(n8096) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n9413), .CLK(n9651), .Q(
        WX2026), .QN(n8094) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n9412), .CLK(n9652), .Q(
        test_so15), .QN(n9139) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n9412), .CLK(n9652), 
        .Q(WX2030), .QN(n8091) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n9412), .CLK(n9652), .Q(
        WX2032), .QN(n8089) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n9412), .CLK(n9652), .Q(
        WX2034) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n9411), .CLK(n9653), .Q(
        WX2036) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n9411), .CLK(n9653), .Q(
        WX2038) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n9411), .CLK(n9653), .Q(
        WX2040) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n9411), .CLK(n9653), .Q(
        WX2042) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n9410), .CLK(n9654), .Q(
        WX2044) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n9410), .CLK(n9654), .Q(
        WX2046) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n9410), .CLK(n9654), .Q(
        WX2048) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n9409), .CLK(n9655), .Q(
        WX2050) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n9409), .CLK(n9655), .Q(
        WX2052) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n9409), .CLK(n9655), .Q(
        WX2054) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n9408), .CLK(n9656), .Q(
        WX2056) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n9408), .CLK(n9656), .Q(
        WX2058) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n9408), .CLK(n9656), .Q(
        WX2060) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n9407), .CLK(n9657), .Q(
        WX2062) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n9407), .CLK(n9657), .Q(
        test_so16), .QN(n9134) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n9407), .CLK(n9657), 
        .Q(WX2066), .QN(n7891) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n9407), .CLK(n9657), .Q(
        WX2068), .QN(n8117) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n9289), .CLK(n9658), .Q(
        WX2070), .QN(n8115) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n9285), .CLK(n9658), .Q(
        WX2072), .QN(n8113) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n9287), .CLK(n9658), .Q(
        WX2074), .QN(n8111) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(test_se), .CLK(n9658), 
        .Q(WX2076), .QN(n8109) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n9289), .CLK(n9658), .Q(
        WX2078), .QN(n8107) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n9285), .CLK(n9658), .Q(
        WX2080), .QN(n8105) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n9406), .CLK(n9659), .Q(
        WX2082), .QN(n8103) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n9406), .CLK(n9659), .Q(
        WX2084), .QN(n8101) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n9406), .CLK(n9659), .Q(
        WX2086), .QN(n8099) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n9406), .CLK(n9659), .Q(
        WX2088), .QN(n8097) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n9406), .CLK(n9659), .Q(
        WX2090), .QN(n8095) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n9412), .CLK(n9652), .Q(
        WX2092), .QN(n8093) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n9412), .CLK(n9652), .Q(
        WX2094), .QN(n8092) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n9412), .CLK(n9652), .Q(
        WX2096), .QN(n8090) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n9412), .CLK(n9652), .Q(
        WX2098), .QN(n8712) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n9411), .CLK(n9653), .Q(
        test_so17), .QN(n9138) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n9411), .CLK(n9653), 
        .Q(WX2102), .QN(n8709) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n9411), .CLK(n9653), .Q(
        WX2104), .QN(n8707) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n9411), .CLK(n9653), .Q(
        WX2106), .QN(n8705) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n9410), .CLK(n9654), .Q(
        WX2108), .QN(n8703) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n9410), .CLK(n9654), .Q(
        WX2110), .QN(n8697) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n9410), .CLK(n9654), .Q(
        WX2112), .QN(n8678) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n9409), .CLK(n9655), .Q(
        WX2114), .QN(n8659) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n9409), .CLK(n9655), .Q(
        WX2116), .QN(n8651) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n9409), .CLK(n9655), .Q(
        WX2118), .QN(n8649) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n9408), .CLK(n9656), .Q(
        WX2120), .QN(n8647) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n9408), .CLK(n9656), .Q(
        WX2122), .QN(n8646) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n9408), .CLK(n9656), .Q(
        WX2124), .QN(n8634) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n9407), .CLK(n9657), .Q(
        WX2126), .QN(n8615) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n9407), .CLK(n9657), .Q(
        WX2128), .QN(n8596) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n9407), .CLK(n9657), .Q(
        WX2130), .QN(n8928) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n9407), .CLK(n9657), .Q(
        WX2132), .QN(n8929) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n9286), .CLK(n9658), .Q(
        WX2134), .QN(n8930) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n9288), .CLK(n9658), .Q(
        test_so18), .QN(n9108) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n9291), .CLK(n9658), 
        .Q(WX2138), .QN(n8931) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n9290), .CLK(n9658), .Q(
        WX2140), .QN(n8932) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n9286), .CLK(n9658), .Q(
        WX2142), .QN(n8933) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n9288), .CLK(n9658), .Q(
        WX2144), .QN(n8934) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n9406), .CLK(n9659), .Q(
        WX2146), .QN(n8935) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n9406), .CLK(n9659), .Q(
        WX2148), .QN(n8936) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n9406), .CLK(n9659), .Q(
        WX2150), .QN(n8937) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n9406), .CLK(n9659), .Q(
        WX2152), .QN(n8938) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n9406), .CLK(n9659), .Q(
        WX2154), .QN(n8939) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n9406), .CLK(n9659), .Q(
        WX2156), .QN(n8940) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n9406), .CLK(n9659), .Q(
        WX2158), .QN(n8941) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n9405), .CLK(n9660), .Q(
        WX2160), .QN(n8731) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n9405), .CLK(n9660), .Q(
        WX2162), .QN(n8942) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n9405), .CLK(n9660), .Q(
        WX2164), .QN(n8943) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n9405), .CLK(n9660), .Q(
        WX2166), .QN(n8944) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n9405), .CLK(n9660), .Q(
        WX2168), .QN(n8945) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n9405), .CLK(n9660), .Q(
        WX2170), .QN(n8732) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n9405), .CLK(n9660), .Q(
        test_so19), .QN(n9101) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n9410), .CLK(n9654), 
        .Q(WX2174), .QN(n8946) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n9410), .CLK(n9654), .Q(
        WX2176), .QN(n8947) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n9409), .CLK(n9655), .Q(
        WX2178), .QN(n8948) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n9409), .CLK(n9655), .Q(
        WX2180), .QN(n8949) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(n9409), .CLK(n9655), .Q(
        WX2182), .QN(n8950) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n9408), .CLK(n9656), .Q(
        WX2184), .QN(n8733) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n9408), .CLK(n9656), .Q(
        WX2186), .QN(n8951) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n9408), .CLK(n9656), .Q(
        WX2188), .QN(n8952) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n9407), .CLK(n9657), .Q(
        WX2190), .QN(n8953) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n9407), .CLK(n9657), .Q(
        WX2192), .QN(n8741) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n9295), .CLK(n9773), .Q(
        CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n9295), .CLK(n9773), 
        .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n9295), .CLK(n9773), 
        .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n9295), .CLK(n9773), 
        .Q(CRC_OUT_8_3), .QN(DFF_355_n1) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n9294), .CLK(n9774), 
        .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n9294), .CLK(n9774), 
        .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n9294), .CLK(n9774), 
        .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n9294), .CLK(n9774), 
        .Q(test_so20), .QN(n9160) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n9294), .CLK(n9774), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n9294), .CLK(n9774), 
        .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n9294), .CLK(n9774), 
        .Q(CRC_OUT_8_10), .QN(DFF_362_n1) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n9294), .CLK(n9774), .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n9294), .CLK(n9774), .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n9294), .CLK(n9774), .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n9294), .CLK(n9774), .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n9294), .CLK(n9774), .Q(CRC_OUT_8_15), .QN(DFF_367_n1) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n9293), .CLK(n9775), .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n9293), .CLK(n9775), .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n9293), .CLK(n9775), .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n9405), .CLK(n9660), .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n9405), .CLK(n9660), .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n9405), .CLK(n9660), .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n9405), .CLK(n9660), .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n9405), .CLK(n9660), .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n9404), .CLK(n9661), .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n9404), .CLK(n9661), .Q(test_so21), .QN(n9159) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n9404), .CLK(n9661), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n9404), .CLK(n9661), .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n9404), .CLK(n9661), .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n9404), .CLK(n9661), .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n9404), .CLK(n9661), .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n9404), .CLK(n9661), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n508), .SI(CRC_OUT_8_31), .SE(n9404), .CLK(n9661), 
        .Q(WX3071), .QN(n9046) );
  SDFFX1 DFF_385_Q_reg ( .D(n509), .SI(WX3071), .SE(n9401), .CLK(n9664), .Q(
        n8644), .QN(n4002) );
  SDFFX1 DFF_386_Q_reg ( .D(n510), .SI(n8644), .SE(n9401), .CLK(n9664), .Q(
        n8643), .QN(n4001) );
  SDFFX1 DFF_387_Q_reg ( .D(n511), .SI(n8643), .SE(n9401), .CLK(n9664), .Q(
        n8642), .QN(n4000) );
  SDFFX1 DFF_388_Q_reg ( .D(n512), .SI(n8642), .SE(n9401), .CLK(n9664), .Q(
        n8641), .QN(n3999) );
  SDFFX1 DFF_389_Q_reg ( .D(n513), .SI(n8641), .SE(n9402), .CLK(n9663), .Q(
        n8640), .QN(n3998) );
  SDFFX1 DFF_390_Q_reg ( .D(n514), .SI(n8640), .SE(n9402), .CLK(n9663), .Q(
        n8639), .QN(n3997) );
  SDFFX1 DFF_391_Q_reg ( .D(n515), .SI(n8639), .SE(n9402), .CLK(n9663), .Q(
        n8638), .QN(n3996) );
  SDFFX1 DFF_392_Q_reg ( .D(n516), .SI(n8638), .SE(n9402), .CLK(n9663), .Q(
        n8637), .QN(n3995) );
  SDFFX1 DFF_393_Q_reg ( .D(n517), .SI(n8637), .SE(n9402), .CLK(n9663), .Q(
        n8636), .QN(n3994) );
  SDFFX1 DFF_394_Q_reg ( .D(n518), .SI(n8636), .SE(n9402), .CLK(n9663), .Q(
        n8635), .QN(n3993) );
  SDFFX1 DFF_395_Q_reg ( .D(n519), .SI(n8635), .SE(n9402), .CLK(n9663), .Q(
        test_so22), .QN(n3992) );
  SDFFX1 DFF_396_Q_reg ( .D(n520), .SI(test_si23), .SE(n9402), .CLK(n9663), 
        .Q(n8632), .QN(n3991) );
  SDFFX1 DFF_397_Q_reg ( .D(n521), .SI(n8632), .SE(n9402), .CLK(n9663), .Q(
        n8631), .QN(n3990) );
  SDFFX1 DFF_398_Q_reg ( .D(n522), .SI(n8631), .SE(n9402), .CLK(n9663), .Q(
        n8630), .QN(n3989) );
  SDFFX1 DFF_399_Q_reg ( .D(n523), .SI(n8630), .SE(n9402), .CLK(n9663), .Q(
        n8629), .QN(n3988) );
  SDFFX1 DFF_400_Q_reg ( .D(n524), .SI(n8629), .SE(n9402), .CLK(n9663), .Q(
        n8628), .QN(n3987) );
  SDFFX1 DFF_401_Q_reg ( .D(n525), .SI(n8628), .SE(n9403), .CLK(n9662), .Q(
        n8627), .QN(n3986) );
  SDFFX1 DFF_402_Q_reg ( .D(n526), .SI(n8627), .SE(n9403), .CLK(n9662), .Q(
        n8626), .QN(n3985) );
  SDFFX1 DFF_403_Q_reg ( .D(n527), .SI(n8626), .SE(n9403), .CLK(n9662), .Q(
        n8625), .QN(n3984) );
  SDFFX1 DFF_404_Q_reg ( .D(n528), .SI(n8625), .SE(n9403), .CLK(n9662), .Q(
        n8624), .QN(n3983) );
  SDFFX1 DFF_405_Q_reg ( .D(n529), .SI(n8624), .SE(n9403), .CLK(n9662), .Q(
        n8623), .QN(n3982) );
  SDFFX1 DFF_406_Q_reg ( .D(n530), .SI(n8623), .SE(n9403), .CLK(n9662), .Q(
        n8622), .QN(n3981) );
  SDFFX1 DFF_407_Q_reg ( .D(n531), .SI(n8622), .SE(n9403), .CLK(n9662), .Q(
        n8621), .QN(n3980) );
  SDFFX1 DFF_408_Q_reg ( .D(n532), .SI(n8621), .SE(n9403), .CLK(n9662), .Q(
        n8620), .QN(n3979) );
  SDFFX1 DFF_409_Q_reg ( .D(n533), .SI(n8620), .SE(n9403), .CLK(n9662), .Q(
        n8619), .QN(n3978) );
  SDFFX1 DFF_410_Q_reg ( .D(n534), .SI(n8619), .SE(n9403), .CLK(n9662), .Q(
        n8618), .QN(n3977) );
  SDFFX1 DFF_411_Q_reg ( .D(n535), .SI(n8618), .SE(n9403), .CLK(n9662), .Q(
        n8617), .QN(n3976) );
  SDFFX1 DFF_412_Q_reg ( .D(n536), .SI(n8617), .SE(n9403), .CLK(n9662), .Q(
        n8616), .QN(n3975) );
  SDFFX1 DFF_413_Q_reg ( .D(n537), .SI(n8616), .SE(n9404), .CLK(n9661), .Q(
        test_so23), .QN(n3974) );
  SDFFX1 DFF_414_Q_reg ( .D(n538), .SI(test_si24), .SE(n9404), .CLK(n9661), 
        .Q(n8613), .QN(n3973) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n9404), .CLK(n9661), .Q(
        n8612), .QN(n3972) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n9295), .CLK(n9773), .Q(
        n8611), .QN(n15981) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n9401), .CLK(n9664), .Q(
        n8610), .QN(n15980) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n9401), .CLK(n9664), .Q(
        n8609), .QN(n15978) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n9400), .CLK(n9665), .Q(
        n8608), .QN(n15976) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n9400), .CLK(n9665), .Q(
        n8607), .QN(n15974) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n9400), .CLK(n9665), .Q(
        n8606), .QN(n15972) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n9400), .CLK(n9665), .Q(
        n8605), .QN(n15970) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n9399), .CLK(n9666), .Q(
        n8604), .QN(n15968) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n9399), .CLK(n9666), .Q(
        n8603), .QN(n15966) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n9399), .CLK(n9666), .Q(
        n8602), .QN(n15964) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n9399), .CLK(n9666), .Q(
        n8601), .QN(n15963) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n9290), .CLK(n9667), .Q(
        n8600), .QN(n15961) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n9289), .CLK(n9667), .Q(
        n8599), .QN(n15959) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n9290), .CLK(n9667), .Q(
        n8598), .QN(n15957) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n9398), .CLK(n9668), .Q(
        n8597), .QN(n15955) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n9295), .CLK(n9773), .Q(
        test_so24), .QN(n9095) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n9398), .CLK(n9668), 
        .Q(WX3263), .QN(n8593) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n9398), .CLK(n9668), .Q(
        WX3265), .QN(n8591) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n9397), .CLK(n9669), .Q(
        WX3267), .QN(n8589) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n9397), .CLK(n9669), .Q(
        WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n9397), .CLK(n9669), .Q(
        WX3271), .QN(n8574) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n9396), .CLK(n9670), .Q(
        WX3273), .QN(n8556) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n9396), .CLK(n9670), .Q(
        WX3275), .QN(n8538) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n9396), .CLK(n9670), .Q(
        WX3277), .QN(n8536) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n9288), .CLK(n9671), .Q(
        WX3279), .QN(n8534) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n9290), .CLK(n9671), .Q(
        WX3281), .QN(n8532) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n9288), .CLK(n9671), .Q(
        WX3283), .QN(n8530) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n9395), .CLK(n9672), .Q(
        WX3285), .QN(n8522) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n9395), .CLK(n9672), .Q(
        WX3287), .QN(n8504) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n9395), .CLK(n9672), .Q(
        WX3289), .QN(n8486) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n9394), .CLK(n9673), .Q(
        WX3291), .QN(n8478) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n9394), .CLK(n9673), .Q(
        WX3293), .QN(n8476) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n9394), .CLK(n9673), .Q(
        WX3295), .QN(n7888) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n9401), .CLK(n9664), .Q(
        test_so25), .QN(n9141) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n9401), .CLK(n9664), 
        .Q(WX3299), .QN(n8086) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n9401), .CLK(n9664), .Q(
        WX3301), .QN(n8084) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n9400), .CLK(n9665), .Q(
        WX3303), .QN(n8082) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n9400), .CLK(n9665), .Q(
        WX3305), .QN(n8081) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n9400), .CLK(n9665), .Q(
        WX3307), .QN(n8079) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n9400), .CLK(n9665), .Q(
        WX3309), .QN(n8077) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n9399), .CLK(n9666), .Q(
        WX3311), .QN(n8075) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n9399), .CLK(n9666), .Q(
        WX3313), .QN(n8073) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n9399), .CLK(n9666), .Q(
        WX3315), .QN(n8071) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n9287), .CLK(n9667), .Q(
        WX3317), .QN(n8069) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n9286), .CLK(n9667), .Q(
        WX3319), .QN(n8067) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n9287), .CLK(n9667), .Q(
        WX3321), .QN(n8065) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n9398), .CLK(n9668), .Q(
        WX3323), .QN(n8063) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n9398), .CLK(n9668), .Q(
        WX3325), .QN(n8061) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n9398), .CLK(n9668), .Q(
        WX3327) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n9397), .CLK(n9669), .Q(
        WX3329) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n9397), .CLK(n9669), .Q(
        WX3331) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n9397), .CLK(n9669), .Q(
        test_so26), .QN(n9137) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n9396), .CLK(n9670), 
        .Q(WX3335) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n9396), .CLK(n9670), .Q(
        WX3337) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n9396), .CLK(n9670), .Q(
        WX3339) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n9289), .CLK(n9671), .Q(
        WX3341) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n9287), .CLK(n9671), .Q(
        WX3343) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n9289), .CLK(n9671), .Q(
        WX3345) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n9395), .CLK(n9672), .Q(
        WX3347) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n9395), .CLK(n9672), .Q(
        WX3349) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n9395), .CLK(n9672), .Q(
        WX3351) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n9394), .CLK(n9673), .Q(
        WX3353) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n9394), .CLK(n9673), .Q(
        WX3355) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n9394), .CLK(n9673), .Q(
        WX3357) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n9393), .CLK(n9674), .Q(
        WX3359), .QN(n7889) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n9401), .CLK(n9664), .Q(
        WX3361), .QN(n8088) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n9401), .CLK(n9664), .Q(
        WX3363), .QN(n8087) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n9401), .CLK(n9664), .Q(
        WX3365), .QN(n8085) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n9400), .CLK(n9665), .Q(
        WX3367), .QN(n8083) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n9400), .CLK(n9665), .Q(
        test_so27), .QN(n9140) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n9400), .CLK(n9665), 
        .Q(WX3371), .QN(n8080) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n9400), .CLK(n9665), .Q(
        WX3373), .QN(n8078) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n9399), .CLK(n9666), .Q(
        WX3375), .QN(n8076) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n9399), .CLK(n9666), .Q(
        WX3377), .QN(n8074) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n9399), .CLK(n9666), .Q(
        WX3379), .QN(n8072) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n9291), .CLK(n9667), .Q(
        WX3381), .QN(n8070) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n9285), .CLK(n9667), .Q(
        WX3383), .QN(n8068) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n9291), .CLK(n9667), .Q(
        WX3385), .QN(n8066) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n9398), .CLK(n9668), .Q(
        WX3387), .QN(n8064) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(n9398), .CLK(n9668), .Q(
        WX3389), .QN(n8062) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n9398), .CLK(n9668), .Q(
        WX3391), .QN(n8594) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(n9397), .CLK(n9669), .Q(
        WX3393), .QN(n8592) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n9397), .CLK(n9669), .Q(
        WX3395), .QN(n8590) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n9397), .CLK(n9669), .Q(
        WX3397), .QN(n8588) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n9396), .CLK(n9670), .Q(
        WX3399), .QN(n8575) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n9396), .CLK(n9670), .Q(
        WX3401), .QN(n8557) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n9396), .CLK(n9670), .Q(
        WX3403), .QN(n8539) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n9286), .CLK(n9671), .Q(
        test_so28), .QN(n9136) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n9291), .CLK(n9671), 
        .Q(WX3407), .QN(n8535) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n9286), .CLK(n9671), .Q(
        WX3409), .QN(n8533) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n9395), .CLK(n9672), .Q(
        WX3411), .QN(n8531) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n9395), .CLK(n9672), .Q(
        WX3413), .QN(n8529) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n9395), .CLK(n9672), .Q(
        WX3415), .QN(n8521) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n9394), .CLK(n9673), .Q(
        WX3417), .QN(n8503) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n9394), .CLK(n9673), .Q(
        WX3419), .QN(n8485) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n9394), .CLK(n9673), .Q(
        WX3421), .QN(n8477) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n9393), .CLK(n9674), .Q(
        WX3423), .QN(n8902) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n9393), .CLK(n9674), .Q(
        WX3425), .QN(n8903) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n9393), .CLK(n9674), .Q(
        WX3427), .QN(n8904) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n9393), .CLK(n9674), .Q(
        WX3429), .QN(n8905) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n9393), .CLK(n9674), .Q(
        WX3431), .QN(n8906) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n9393), .CLK(n9674), .Q(
        WX3433), .QN(n8907) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n9393), .CLK(n9674), .Q(
        WX3435), .QN(n8908) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n9393), .CLK(n9674), .Q(
        WX3437), .QN(n8909) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n9393), .CLK(n9674), .Q(
        test_so29), .QN(n9107) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n9399), .CLK(n9666), 
        .Q(WX3441), .QN(n8910) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n9399), .CLK(n9666), .Q(
        WX3443), .QN(n8911) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(test_se), .CLK(n9667), 
        .Q(WX3445), .QN(n8912) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n9288), .CLK(n9667), .Q(
        WX3447), .QN(n8913) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(test_se), .CLK(n9667), 
        .Q(WX3449), .QN(n8914) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n9398), .CLK(n9668), .Q(
        WX3451), .QN(n8915) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n9398), .CLK(n9668), .Q(
        WX3453), .QN(n8728) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n9398), .CLK(n9668), .Q(
        WX3455), .QN(n8916) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n9397), .CLK(n9669), .Q(
        WX3457), .QN(n8917) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n9397), .CLK(n9669), .Q(
        WX3459), .QN(n8918) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n9397), .CLK(n9669), .Q(
        WX3461), .QN(n8919) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n9396), .CLK(n9670), .Q(
        WX3463), .QN(n8729) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n9396), .CLK(n9670), .Q(
        WX3465), .QN(n8920) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n9396), .CLK(n9670), .Q(
        WX3467), .QN(n8921) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n9285), .CLK(n9671), .Q(
        WX3469), .QN(n8922) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(test_se), .CLK(n9671), 
        .Q(WX3471), .QN(n8923) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n9285), .CLK(n9671), .Q(
        test_so30), .QN(n9100) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n9395), .CLK(n9672), 
        .Q(WX3475), .QN(n8924) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n9395), .CLK(n9672), .Q(
        WX3477), .QN(n8730) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n9395), .CLK(n9672), .Q(
        WX3479), .QN(n8925) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n9394), .CLK(n9673), .Q(
        WX3481), .QN(n8926) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n9394), .CLK(n9673), .Q(
        WX3483), .QN(n8927) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n9394), .CLK(n9673), .Q(
        WX3485), .QN(n8740) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n9298), .CLK(n9770), .Q(
        CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_3), .QN(DFF_547_n1) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n9297), .CLK(n9771), 
        .Q(test_so31), .QN(n9090) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n9297), .CLK(n9771), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n9297), .CLK(n9771), .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_15), .QN(DFF_559_n1) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n9296), .CLK(n9772), .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n9295), .CLK(n9773), .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n9295), .CLK(n9773), .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n9295), .CLK(n9773), .Q(test_so32), .QN(n9158) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n9295), .CLK(n9773), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n9295), .CLK(n9773), .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n9295), .CLK(n9773), .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n9393), .CLK(n9674), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n749), .SI(CRC_OUT_7_31), .SE(n9393), .CLK(n9674), 
        .Q(WX4364), .QN(n9047) );
  SDFFX1 DFF_577_Q_reg ( .D(n750), .SI(WX4364), .SE(n9390), .CLK(n9677), .Q(
        n8586), .QN(n3971) );
  SDFFX1 DFF_578_Q_reg ( .D(n751), .SI(n8586), .SE(n9390), .CLK(n9677), .Q(
        n8585), .QN(n3970) );
  SDFFX1 DFF_579_Q_reg ( .D(n752), .SI(n8585), .SE(n9390), .CLK(n9677), .Q(
        n8584), .QN(n3969) );
  SDFFX1 DFF_580_Q_reg ( .D(n753), .SI(n8584), .SE(n9390), .CLK(n9677), .Q(
        n8583), .QN(n3968) );
  SDFFX1 DFF_581_Q_reg ( .D(n754), .SI(n8583), .SE(n9390), .CLK(n9677), .Q(
        n8582), .QN(n3967) );
  SDFFX1 DFF_582_Q_reg ( .D(n755), .SI(n8582), .SE(n9390), .CLK(n9677), .Q(
        n8581), .QN(n3966) );
  SDFFX1 DFF_583_Q_reg ( .D(n756), .SI(n8581), .SE(n9390), .CLK(n9677), .Q(
        n8580), .QN(n3965) );
  SDFFX1 DFF_584_Q_reg ( .D(n757), .SI(n8580), .SE(n9391), .CLK(n9676), .Q(
        n8579), .QN(n3964) );
  SDFFX1 DFF_585_Q_reg ( .D(n758), .SI(n8579), .SE(n9391), .CLK(n9676), .Q(
        n8578), .QN(n3963) );
  SDFFX1 DFF_586_Q_reg ( .D(n759), .SI(n8578), .SE(n9391), .CLK(n9676), .Q(
        n8577), .QN(n3962) );
  SDFFX1 DFF_587_Q_reg ( .D(n760), .SI(n8577), .SE(n9391), .CLK(n9676), .Q(
        n8576), .QN(n3961) );
  SDFFX1 DFF_588_Q_reg ( .D(n761), .SI(n8576), .SE(n9391), .CLK(n9676), .Q(
        test_so33), .QN(n3960) );
  SDFFX1 DFF_589_Q_reg ( .D(n762), .SI(test_si34), .SE(n9391), .CLK(n9676), 
        .Q(n8573), .QN(n3959) );
  SDFFX1 DFF_590_Q_reg ( .D(n763), .SI(n8573), .SE(n9391), .CLK(n9676), .Q(
        n8572), .QN(n3958) );
  SDFFX1 DFF_591_Q_reg ( .D(n764), .SI(n8572), .SE(n9391), .CLK(n9676), .Q(
        n8571), .QN(n3957) );
  SDFFX1 DFF_592_Q_reg ( .D(n765), .SI(n8571), .SE(n9391), .CLK(n9676), .Q(
        n8570), .QN(n3956) );
  SDFFX1 DFF_593_Q_reg ( .D(n766), .SI(n8570), .SE(n9391), .CLK(n9676), .Q(
        n8569), .QN(n3955) );
  SDFFX1 DFF_594_Q_reg ( .D(n767), .SI(n8569), .SE(n9391), .CLK(n9676), .Q(
        n8568), .QN(n3954) );
  SDFFX1 DFF_595_Q_reg ( .D(n768), .SI(n8568), .SE(n9391), .CLK(n9676), .Q(
        n8567), .QN(n3953) );
  SDFFX1 DFF_596_Q_reg ( .D(n769), .SI(n8567), .SE(n9392), .CLK(n9675), .Q(
        n8566), .QN(n3952) );
  SDFFX1 DFF_597_Q_reg ( .D(n770), .SI(n8566), .SE(n9392), .CLK(n9675), .Q(
        n8565), .QN(n3951) );
  SDFFX1 DFF_598_Q_reg ( .D(n771), .SI(n8565), .SE(n9392), .CLK(n9675), .Q(
        n8564), .QN(n3950) );
  SDFFX1 DFF_599_Q_reg ( .D(n772), .SI(n8564), .SE(n9392), .CLK(n9675), .Q(
        n8563), .QN(n3949) );
  SDFFX1 DFF_600_Q_reg ( .D(n773), .SI(n8563), .SE(n9392), .CLK(n9675), .Q(
        n8562), .QN(n3948) );
  SDFFX1 DFF_601_Q_reg ( .D(n774), .SI(n8562), .SE(n9392), .CLK(n9675), .Q(
        n8561), .QN(n3947) );
  SDFFX1 DFF_602_Q_reg ( .D(n775), .SI(n8561), .SE(n9392), .CLK(n9675), .Q(
        n8560), .QN(n3946) );
  SDFFX1 DFF_603_Q_reg ( .D(n776), .SI(n8560), .SE(n9392), .CLK(n9675), .Q(
        n8559), .QN(n3945) );
  SDFFX1 DFF_604_Q_reg ( .D(n777), .SI(n8559), .SE(n9392), .CLK(n9675), .Q(
        n8558), .QN(n3944) );
  SDFFX1 DFF_605_Q_reg ( .D(n778), .SI(n8558), .SE(n9392), .CLK(n9675), .Q(
        test_so34), .QN(n3943) );
  SDFFX1 DFF_606_Q_reg ( .D(n779), .SI(test_si35), .SE(n9392), .CLK(n9675), 
        .Q(n8555), .QN(n3942) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n9392), .CLK(n9675), .Q(
        n8554), .QN(n3941) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n9298), .CLK(n9770), .Q(
        n8553), .QN(n15952) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n9390), .CLK(n9677), .Q(
        n8552), .QN(n15951) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n9390), .CLK(n9677), .Q(
        n8551), .QN(n15950) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n9287), .CLK(n9678), .Q(
        n8550), .QN(n15949) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n9285), .CLK(n9678), .Q(
        n8549), .QN(n15948) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n9288), .CLK(n9678), .Q(
        n8548), .QN(n15947) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n9389), .CLK(n9679), .Q(
        n8547), .QN(n15946) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n9389), .CLK(n9679), .Q(
        n8546), .QN(n15945) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n9389), .CLK(n9679), .Q(
        n8545), .QN(n15944) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n9389), .CLK(n9679), .Q(
        n8544), .QN(n15943) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n9388), .CLK(n9680), .Q(
        n8543), .QN(n15942) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n9388), .CLK(n9680), .Q(
        n8542), .QN(n15941) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n9387), .CLK(n9681), .Q(
        n8541), .QN(n15940) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n9387), .CLK(n9681), .Q(
        n8540), .QN(n15939) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n9298), .CLK(n9770), .Q(
        test_so35), .QN(n9094) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n9386), .CLK(n9682), 
        .Q(n8537), .QN(n15938) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n9386), .CLK(n9682), .Q(
        WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n9386), .CLK(n9682), .Q(
        WX4558), .QN(n8472) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n9386), .CLK(n9682), .Q(
        WX4560), .QN(n8471) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n9385), .CLK(n9683), .Q(
        WX4562), .QN(n8468) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n9385), .CLK(n9683), .Q(
        WX4564), .QN(n8450) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n9385), .CLK(n9683), .Q(
        WX4566), .QN(n8432) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n9384), .CLK(n9684), .Q(
        WX4568), .QN(n8419) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n9384), .CLK(n9684), .Q(
        WX4570), .QN(n8417) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n9384), .CLK(n9684), .Q(
        WX4572), .QN(n8415) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n9383), .CLK(n9685), .Q(
        WX4574), .QN(n8413) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n9383), .CLK(n9685), .Q(
        WX4576), .QN(n8398) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n9383), .CLK(n9685), .Q(
        WX4578), .QN(n8380) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n9382), .CLK(n9686), .Q(
        WX4580), .QN(n8362) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n9382), .CLK(n9686), .Q(
        WX4582), .QN(n8360) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n9382), .CLK(n9686), .Q(
        WX4584), .QN(n8358) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n9381), .CLK(n9687), .Q(
        test_so36), .QN(n9130) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n9298), .CLK(n9770), 
        .Q(WX4588), .QN(n7886) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n9390), .CLK(n9677), .Q(
        WX4590), .QN(n8060) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n9390), .CLK(n9677), .Q(
        WX4592), .QN(n8058) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n9291), .CLK(n9678), .Q(
        WX4594), .QN(n8056) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n9290), .CLK(n9678), .Q(
        WX4596), .QN(n8054) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n9287), .CLK(n9678), .Q(
        WX4598), .QN(n8052) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n9290), .CLK(n9678), .Q(
        WX4600), .QN(n8050) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n9389), .CLK(n9679), .Q(
        WX4602), .QN(n8048) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n9389), .CLK(n9679), .Q(
        WX4604), .QN(n8046) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n9388), .CLK(n9680), .Q(
        WX4606), .QN(n8044) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n9388), .CLK(n9680), .Q(
        WX4608), .QN(n8042) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n9388), .CLK(n9680), .Q(
        WX4610), .QN(n8040) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n9388), .CLK(n9680), .Q(
        WX4612), .QN(n8038) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n9387), .CLK(n9681), .Q(
        WX4614), .QN(n8036) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n9387), .CLK(n9681), .Q(
        WX4616), .QN(n8034) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n9387), .CLK(n9681), .Q(
        WX4618), .QN(n8032) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n9386), .CLK(n9682), .Q(
        test_so37), .QN(n9132) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n9386), .CLK(n9682), 
        .Q(WX4622) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n9386), .CLK(n9682), .Q(
        WX4624) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n9385), .CLK(n9683), .Q(
        WX4626) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n9385), .CLK(n9683), .Q(
        WX4628) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n9385), .CLK(n9683), .Q(
        WX4630) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n9384), .CLK(n9684), .Q(
        WX4632) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n9384), .CLK(n9684), .Q(
        WX4634) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n9384), .CLK(n9684), .Q(
        WX4636) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n9383), .CLK(n9685), .Q(
        WX4638) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n9383), .CLK(n9685), .Q(
        WX4640) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n9383), .CLK(n9685), .Q(
        WX4642) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n9382), .CLK(n9686), .Q(
        WX4644) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n9382), .CLK(n9686), .Q(
        WX4646) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n9382), .CLK(n9686), .Q(
        WX4648) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n9381), .CLK(n9687), .Q(
        WX4650) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n9381), .CLK(n9687), .Q(
        WX4652), .QN(n7887) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n9381), .CLK(n9687), .Q(
        test_so38), .QN(n9133) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n9390), .CLK(n9677), 
        .Q(WX4656), .QN(n8059) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(test_se), .CLK(n9678), 
        .Q(WX4658), .QN(n8057) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n9289), .CLK(n9678), .Q(
        WX4660), .QN(n8055) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n9291), .CLK(n9678), .Q(
        WX4662), .QN(n8053) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n9389), .CLK(n9679), .Q(
        WX4664), .QN(n8051) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n9389), .CLK(n9679), .Q(
        WX4666), .QN(n8049) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n9389), .CLK(n9679), .Q(
        WX4668), .QN(n8047) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n9388), .CLK(n9680), .Q(
        WX4670), .QN(n8045) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n9388), .CLK(n9680), .Q(
        WX4672), .QN(n8043) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n9388), .CLK(n9680), .Q(
        WX4674), .QN(n8041) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n9387), .CLK(n9681), .Q(
        WX4676), .QN(n8039) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n9387), .CLK(n9681), .Q(
        WX4678), .QN(n8037) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n9387), .CLK(n9681), .Q(
        WX4680), .QN(n8035) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n9387), .CLK(n9681), .Q(
        WX4682), .QN(n8033) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n9386), .CLK(n9682), .Q(
        WX4684), .QN(n8475) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n9386), .CLK(n9682), .Q(
        WX4686), .QN(n8473) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n9385), .CLK(n9683), .Q(
        test_so39), .QN(n9131) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n9385), .CLK(n9683), 
        .Q(WX4690), .QN(n8469) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n9385), .CLK(n9683), .Q(
        WX4692), .QN(n8451) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n9384), .CLK(n9684), .Q(
        WX4694), .QN(n8433) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n9384), .CLK(n9684), .Q(
        WX4696), .QN(n8420) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n9384), .CLK(n9684), .Q(
        WX4698), .QN(n8418) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n9383), .CLK(n9685), .Q(
        WX4700), .QN(n8416) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n9383), .CLK(n9685), .Q(
        WX4702), .QN(n8414) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n9383), .CLK(n9685), .Q(
        WX4704), .QN(n8412) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n9382), .CLK(n9686), .Q(
        WX4706), .QN(n8397) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n9382), .CLK(n9686), .Q(
        WX4708), .QN(n8379) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n9382), .CLK(n9686), .Q(
        WX4710), .QN(n8361) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n9381), .CLK(n9687), .Q(
        WX4712), .QN(n8359) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n9381), .CLK(n9687), .Q(
        WX4714), .QN(n8357) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n9381), .CLK(n9687), .Q(
        WX4716), .QN(n8875) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n9381), .CLK(n9687), .Q(
        WX4718), .QN(n8876) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n9381), .CLK(n9687), .Q(
        WX4720), .QN(n8877) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n9381), .CLK(n9687), .Q(
        test_so40), .QN(n9106) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n9286), .CLK(n9678), 
        .Q(WX4724), .QN(n8878) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(test_se), .CLK(n9678), 
        .Q(WX4726), .QN(n8879) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n9389), .CLK(n9679), .Q(
        WX4728), .QN(n8880) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n9389), .CLK(n9679), .Q(
        WX4730), .QN(n8881) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n9389), .CLK(n9679), .Q(
        WX4732), .QN(n8882) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n9388), .CLK(n9680), .Q(
        WX4734), .QN(n8883) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n9388), .CLK(n9680), .Q(
        WX4736), .QN(n8884) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n9388), .CLK(n9680), .Q(
        WX4738), .QN(n8885) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n9387), .CLK(n9681), .Q(
        WX4740), .QN(n8886) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n9387), .CLK(n9681), .Q(
        WX4742), .QN(n8887) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n9387), .CLK(n9681), .Q(
        WX4744), .QN(n8888) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n9386), .CLK(n9682), .Q(
        WX4746), .QN(n8726) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n9386), .CLK(n9682), .Q(
        WX4748), .QN(n8889) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n9386), .CLK(n9682), .Q(
        WX4750), .QN(n8890) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n9385), .CLK(n9683), .Q(
        WX4752), .QN(n8891) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n9385), .CLK(n9683), .Q(
        WX4754), .QN(n8892) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n9385), .CLK(n9683), .Q(
        test_so41), .QN(n9088) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n9384), .CLK(n9684), 
        .Q(WX4758), .QN(n8893) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n9384), .CLK(n9684), .Q(
        WX4760), .QN(n8894) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n9384), .CLK(n9684), .Q(
        WX4762), .QN(n8895) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n9383), .CLK(n9685), .Q(
        WX4764), .QN(n8896) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n9383), .CLK(n9685), .Q(
        WX4766), .QN(n8897) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n9383), .CLK(n9685), .Q(
        WX4768), .QN(n8898) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n9382), .CLK(n9686), .Q(
        WX4770), .QN(n8727) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n9382), .CLK(n9686), .Q(
        WX4772), .QN(n8899) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n9382), .CLK(n9686), .Q(
        WX4774), .QN(n8900) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n9381), .CLK(n9687), .Q(
        WX4776), .QN(n8901) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n9381), .CLK(n9687), .Q(
        WX4778), .QN(n8739) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n9300), .CLK(n9768), .Q(
        CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n9300), .CLK(n9768), 
        .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n9300), .CLK(n9768), 
        .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n9300), .CLK(n9768), 
        .Q(CRC_OUT_6_3), .QN(DFF_739_n1) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n9300), .CLK(n9768), 
        .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n9300), .CLK(n9768), 
        .Q(test_so42), .QN(n9157) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n9300), .CLK(n9768), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n9300), .CLK(n9768), 
        .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n9300), .CLK(n9768), 
        .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n9300), .CLK(n9768), 
        .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n9299), .CLK(n9769), 
        .Q(CRC_OUT_6_10), .QN(DFF_746_n1) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_15), .QN(DFF_751_n1) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n9299), .CLK(n9769), .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n9298), .CLK(n9770), .Q(test_so43), .QN(n9156) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n9298), .CLK(n9770), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n9298), .CLK(n9770), .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n9298), .CLK(n9770), .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n9298), .CLK(n9770), .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n9298), .CLK(n9770), .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n9298), .CLK(n9770), .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n9298), .CLK(n9770), .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n9380), .CLK(n9688), .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n9380), .CLK(n9688), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n990), .SI(CRC_OUT_6_31), .SE(n9380), .CLK(n9688), 
        .Q(WX5657), .QN(n9048) );
  SDFFX1 DFF_769_Q_reg ( .D(n991), .SI(WX5657), .SE(n9378), .CLK(n9690), .Q(
        n8528), .QN(n3940) );
  SDFFX1 DFF_770_Q_reg ( .D(n992), .SI(n8528), .SE(n9378), .CLK(n9690), .Q(
        n8527), .QN(n3939) );
  SDFFX1 DFF_771_Q_reg ( .D(n993), .SI(n8527), .SE(n9378), .CLK(n9690), .Q(
        n8526), .QN(n3938) );
  SDFFX1 DFF_772_Q_reg ( .D(n994), .SI(n8526), .SE(n9378), .CLK(n9690), .Q(
        n8525), .QN(n3937) );
  SDFFX1 DFF_773_Q_reg ( .D(n995), .SI(n8525), .SE(n9378), .CLK(n9690), .Q(
        n8524), .QN(n3936) );
  SDFFX1 DFF_774_Q_reg ( .D(n996), .SI(n8524), .SE(n9378), .CLK(n9690), .Q(
        n8523), .QN(n3935) );
  SDFFX1 DFF_775_Q_reg ( .D(n997), .SI(n8523), .SE(n9378), .CLK(n9690), .Q(
        test_so44), .QN(n3934) );
  SDFFX1 DFF_776_Q_reg ( .D(n998), .SI(test_si45), .SE(n9378), .CLK(n9690), 
        .Q(n8520), .QN(n3933) );
  SDFFX1 DFF_777_Q_reg ( .D(n999), .SI(n8520), .SE(n9378), .CLK(n9690), .Q(
        n8519), .QN(n3932) );
  SDFFX1 DFF_778_Q_reg ( .D(n1000), .SI(n8519), .SE(n9378), .CLK(n9690), .Q(
        n8518), .QN(n3931) );
  SDFFX1 DFF_779_Q_reg ( .D(n1001), .SI(n8518), .SE(n9379), .CLK(n9689), .Q(
        n8517), .QN(n3930) );
  SDFFX1 DFF_780_Q_reg ( .D(n1002), .SI(n8517), .SE(n9379), .CLK(n9689), .Q(
        n8516), .QN(n3929) );
  SDFFX1 DFF_781_Q_reg ( .D(n1003), .SI(n8516), .SE(n9379), .CLK(n9689), .Q(
        n8515), .QN(n3928) );
  SDFFX1 DFF_782_Q_reg ( .D(n1004), .SI(n8515), .SE(n9379), .CLK(n9689), .Q(
        n8514), .QN(n3927) );
  SDFFX1 DFF_783_Q_reg ( .D(n1005), .SI(n8514), .SE(n9379), .CLK(n9689), .Q(
        n8513), .QN(n3926) );
  SDFFX1 DFF_784_Q_reg ( .D(n1006), .SI(n8513), .SE(n9379), .CLK(n9689), .Q(
        n8512), .QN(n3925) );
  SDFFX1 DFF_785_Q_reg ( .D(n1007), .SI(n8512), .SE(n9379), .CLK(n9689), .Q(
        n8511), .QN(n3924) );
  SDFFX1 DFF_786_Q_reg ( .D(n1008), .SI(n8511), .SE(n9379), .CLK(n9689), .Q(
        n8510), .QN(n3923) );
  SDFFX1 DFF_787_Q_reg ( .D(n1009), .SI(n8510), .SE(n9379), .CLK(n9689), .Q(
        n8509), .QN(n3922) );
  SDFFX1 DFF_788_Q_reg ( .D(n1010), .SI(n8509), .SE(n9379), .CLK(n9689), .Q(
        n8508), .QN(n3921) );
  SDFFX1 DFF_789_Q_reg ( .D(n1011), .SI(n8508), .SE(n9379), .CLK(n9689), .Q(
        n8507), .QN(n3920) );
  SDFFX1 DFF_790_Q_reg ( .D(n1012), .SI(n8507), .SE(n9379), .CLK(n9689), .Q(
        n8506), .QN(n3919) );
  SDFFX1 DFF_791_Q_reg ( .D(n1013), .SI(n8506), .SE(n9380), .CLK(n9688), .Q(
        n8505), .QN(n3918) );
  SDFFX1 DFF_792_Q_reg ( .D(n1014), .SI(n8505), .SE(n9380), .CLK(n9688), .Q(
        test_so45), .QN(n3917) );
  SDFFX1 DFF_793_Q_reg ( .D(n1015), .SI(test_si46), .SE(n9380), .CLK(n9688), 
        .Q(n8502), .QN(n3916) );
  SDFFX1 DFF_794_Q_reg ( .D(n1016), .SI(n8502), .SE(n9380), .CLK(n9688), .Q(
        n8501), .QN(n3915) );
  SDFFX1 DFF_795_Q_reg ( .D(n1017), .SI(n8501), .SE(n9380), .CLK(n9688), .Q(
        n8500), .QN(n3914) );
  SDFFX1 DFF_796_Q_reg ( .D(n1018), .SI(n8500), .SE(n9380), .CLK(n9688), .Q(
        n8499), .QN(n3913) );
  SDFFX1 DFF_797_Q_reg ( .D(n1019), .SI(n8499), .SE(n9380), .CLK(n9688), .Q(
        n8498), .QN(n3912) );
  SDFFX1 DFF_798_Q_reg ( .D(n1020), .SI(n8498), .SE(n9380), .CLK(n9688), .Q(
        n8497), .QN(n3911) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n9380), .CLK(n9688), .Q(
        n8496), .QN(n3910) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n9300), .CLK(n9768), .Q(
        n8495), .QN(n15937) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n9378), .CLK(n9690), .Q(
        n8494), .QN(n15936) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n9377), .CLK(n9691), .Q(
        n8493), .QN(n15935) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n9377), .CLK(n9691), .Q(
        n8492), .QN(n15934) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n9377), .CLK(n9691), .Q(
        n8491), .QN(n15933) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n9377), .CLK(n9691), .Q(
        n8490), .QN(n15932) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n9377), .CLK(n9691), .Q(
        n8489), .QN(n15931) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n9377), .CLK(n9691), .Q(
        n8488), .QN(n15930) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n9376), .CLK(n9692), .Q(
        n8487), .QN(n15929) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n9376), .CLK(n9692), .Q(
        test_so46), .QN(n9093) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n9376), .CLK(n9692), 
        .Q(n8484), .QN(n15928) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n9376), .CLK(n9692), .Q(
        n8483), .QN(n15927) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n9376), .CLK(n9692), .Q(
        n8482), .QN(n15926) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n9375), .CLK(n9693), .Q(
        n8481), .QN(n15925) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n9375), .CLK(n9693), .Q(
        n8480), .QN(n15924) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n9375), .CLK(n9693), .Q(
        n8479), .QN(n15923) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n9375), .CLK(n9693), .Q(
        WX5849), .QN(n8355) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n9374), .CLK(n9694), .Q(
        WX5851), .QN(n8345) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n9374), .CLK(n9694), .Q(
        WX5853), .QN(n8327) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n9374), .CLK(n9694), .Q(
        WX5855), .QN(n8309) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n9373), .CLK(n9695), .Q(
        WX5857), .QN(n8303) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n9373), .CLK(n9695), .Q(
        WX5859), .QN(n8301) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n9373), .CLK(n9695), .Q(
        WX5861), .QN(n8299) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n9372), .CLK(n9696), .Q(
        WX5863), .QN(n8297) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n9372), .CLK(n9696), .Q(
        WX5865), .QN(n8292) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n9372), .CLK(n9696), .Q(
        WX5867), .QN(n8274) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n9371), .CLK(n9697), .Q(
        test_so47), .QN(n9127) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n9371), .CLK(n9697), 
        .Q(WX5871), .QN(n8255) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n9371), .CLK(n9697), .Q(
        WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n9370), .CLK(n9698), .Q(
        WX5875), .QN(n8242) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n9370), .CLK(n9698), .Q(
        WX5877), .QN(n8241) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n9370), .CLK(n9698), .Q(
        WX5879), .QN(n8239) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n9369), .CLK(n9699), .Q(
        WX5881), .QN(n7884) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n9378), .CLK(n9690), .Q(
        WX5883), .QN(n8030) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n9377), .CLK(n9691), .Q(
        WX5885), .QN(n8028) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n9377), .CLK(n9691), .Q(
        WX5887), .QN(n8026) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n9377), .CLK(n9691), .Q(
        WX5889), .QN(n8024) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n9377), .CLK(n9691), .Q(
        WX5891), .QN(n8022) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n9377), .CLK(n9691), .Q(
        WX5893), .QN(n8020) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n9377), .CLK(n9691), .Q(
        WX5895), .QN(n8018) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n9376), .CLK(n9692), .Q(
        WX5897), .QN(n8016) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n9376), .CLK(n9692), .Q(
        WX5899), .QN(n8014) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n9376), .CLK(n9692), .Q(
        WX5901), .QN(n8012) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n9376), .CLK(n9692), .Q(
        test_so48), .QN(n9129) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n9376), .CLK(n9692), 
        .Q(WX5905), .QN(n8009) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n9375), .CLK(n9693), .Q(
        WX5907), .QN(n8008) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n9375), .CLK(n9693), .Q(
        WX5909), .QN(n8006) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n9375), .CLK(n9693), .Q(
        WX5911), .QN(n8004) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n9375), .CLK(n9693), .Q(
        WX5913) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n9374), .CLK(n9694), .Q(
        WX5915) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n9374), .CLK(n9694), .Q(
        WX5917) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n9374), .CLK(n9694), .Q(
        WX5919) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n9373), .CLK(n9695), .Q(
        WX5921) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n9373), .CLK(n9695), .Q(
        WX5923) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n9373), .CLK(n9695), .Q(
        WX5925) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n9372), .CLK(n9696), .Q(
        WX5927) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n9372), .CLK(n9696), .Q(
        WX5929) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n9372), .CLK(n9696), .Q(
        WX5931) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n9371), .CLK(n9697), .Q(
        WX5933) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n9371), .CLK(n9697), .Q(
        WX5935) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n9371), .CLK(n9697), .Q(
        test_so49), .QN(n9126) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n9370), .CLK(n9698), 
        .Q(WX5939) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n9370), .CLK(n9698), .Q(
        WX5941) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n9370), .CLK(n9698), .Q(
        WX5943) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n9369), .CLK(n9699), .Q(
        WX5945), .QN(n7885) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n9369), .CLK(n9699), .Q(
        WX5947), .QN(n8031) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n9369), .CLK(n9699), .Q(
        WX5949), .QN(n8029) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n9369), .CLK(n9699), .Q(
        WX5951), .QN(n8027) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n9369), .CLK(n9699), .Q(
        WX5953), .QN(n8025) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n9368), .CLK(n9700), .Q(
        WX5955), .QN(n8023) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n9368), .CLK(n9700), .Q(
        WX5957), .QN(n8021) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n9368), .CLK(n9700), .Q(
        WX5959), .QN(n8019) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n9368), .CLK(n9700), .Q(
        WX5961), .QN(n8017) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n9368), .CLK(n9700), .Q(
        WX5963), .QN(n8015) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n9368), .CLK(n9700), .Q(
        WX5965), .QN(n8013) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n9376), .CLK(n9692), .Q(
        WX5967), .QN(n8011) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n9376), .CLK(n9692), .Q(
        WX5969), .QN(n8010) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n9375), .CLK(n9693), .Q(
        test_so50), .QN(n9128) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n9375), .CLK(n9693), 
        .Q(WX5973), .QN(n8007) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n9375), .CLK(n9693), .Q(
        WX5975), .QN(n8005) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n9375), .CLK(n9693), .Q(
        WX5977), .QN(n8356) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n9374), .CLK(n9694), .Q(
        WX5979), .QN(n8354) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n9374), .CLK(n9694), .Q(
        WX5981), .QN(n8344) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n9374), .CLK(n9694), .Q(
        WX5983), .QN(n8326) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n9373), .CLK(n9695), .Q(
        WX5985), .QN(n8308) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n9373), .CLK(n9695), .Q(
        WX5987), .QN(n8302) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n9373), .CLK(n9695), .Q(
        WX5989), .QN(n8300) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n9372), .CLK(n9696), .Q(
        WX5991), .QN(n8298) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n9372), .CLK(n9696), .Q(
        WX5993), .QN(n8296) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n9372), .CLK(n9696), .Q(
        WX5995), .QN(n8291) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n9371), .CLK(n9697), .Q(
        WX5997), .QN(n8273) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n9371), .CLK(n9697), .Q(
        WX5999), .QN(n8256) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n9371), .CLK(n9697), .Q(
        WX6001), .QN(n8245) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n9370), .CLK(n9698), .Q(
        WX6003), .QN(n8243) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n9370), .CLK(n9698), .Q(
        test_so51), .QN(n9125) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n9370), .CLK(n9698), 
        .Q(WX6007), .QN(n8240) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n9369), .CLK(n9699), .Q(
        WX6009), .QN(n8847) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n9369), .CLK(n9699), .Q(
        WX6011), .QN(n8848) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n9369), .CLK(n9699), .Q(
        WX6013), .QN(n8849) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n9369), .CLK(n9699), .Q(
        WX6015), .QN(n8850) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n9369), .CLK(n9699), .Q(
        WX6017), .QN(n8851) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n9368), .CLK(n9700), .Q(
        WX6019), .QN(n8852) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n9368), .CLK(n9700), .Q(
        WX6021), .QN(n8853) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n9368), .CLK(n9700), .Q(
        WX6023), .QN(n8854) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n9368), .CLK(n9700), .Q(
        WX6025), .QN(n8855) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n9368), .CLK(n9700), .Q(
        WX6027), .QN(n8856) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n9368), .CLK(n9700), .Q(
        WX6029), .QN(n8857) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n9367), .CLK(n9701), .Q(
        WX6031), .QN(n8858) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n9367), .CLK(n9701), .Q(
        WX6033), .QN(n8859) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n9367), .CLK(n9701), .Q(
        WX6035), .QN(n8860) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n9367), .CLK(n9701), .Q(
        WX6037), .QN(n8861) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n9367), .CLK(n9701), .Q(
        test_so52), .QN(n9089) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n9374), .CLK(n9694), 
        .Q(WX6041), .QN(n8862) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n9374), .CLK(n9694), .Q(
        WX6043), .QN(n8863) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n9374), .CLK(n9694), .Q(
        WX6045), .QN(n8864) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n9373), .CLK(n9695), .Q(
        WX6047), .QN(n8865) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n9373), .CLK(n9695), .Q(
        WX6049), .QN(n8724) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n9373), .CLK(n9695), .Q(
        WX6051), .QN(n8866) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n9372), .CLK(n9696), .Q(
        WX6053), .QN(n8867) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n9372), .CLK(n9696), .Q(
        WX6055), .QN(n8868) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n9372), .CLK(n9696), .Q(
        WX6057), .QN(n8869) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n9371), .CLK(n9697), .Q(
        WX6059), .QN(n8870) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n9371), .CLK(n9697), .Q(
        WX6061), .QN(n8871) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n9371), .CLK(n9697), .Q(
        WX6063), .QN(n8725) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n9370), .CLK(n9698), .Q(
        WX6065), .QN(n8872) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n9370), .CLK(n9698), .Q(
        WX6067), .QN(n8873) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n9370), .CLK(n9698), .Q(
        WX6069), .QN(n8874) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n9369), .CLK(n9699), .Q(
        WX6071), .QN(n8738) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n9302), .CLK(n9766), .Q(
        test_so53), .QN(n9155) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n9302), .CLK(n9766), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n9302), .CLK(n9766), 
        .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n9302), .CLK(n9766), 
        .Q(CRC_OUT_5_3), .QN(DFF_931_n1) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n9302), .CLK(n9766), 
        .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n9302), .CLK(n9766), 
        .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n9302), .CLK(n9766), 
        .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n9302), .CLK(n9766), 
        .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n9301), .CLK(n9767), 
        .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n9301), .CLK(n9767), 
        .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n9301), .CLK(n9767), 
        .Q(CRC_OUT_5_10), .QN(DFF_938_n1) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n9301), .CLK(n9767), .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n9301), .CLK(n9767), .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n9301), .CLK(n9767), .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n9301), .CLK(n9767), .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n9301), .CLK(n9767), .Q(CRC_OUT_5_15), .QN(DFF_943_n1) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n9301), .CLK(n9767), .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n9301), .CLK(n9767), .Q(test_so54), .QN(n9154) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n9301), .CLK(n9767), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n9301), .CLK(n9767), .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n9300), .CLK(n9768), .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n9367), .CLK(n9701), .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n9367), .CLK(n9701), .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n9367), .CLK(n9701), .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n9367), .CLK(n9701), .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n9367), .CLK(n9701), .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n9367), .CLK(n9701), .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n9367), .CLK(n9701), .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n9366), .CLK(n9702), .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n9366), .CLK(n9702), .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n9366), .CLK(n9702), .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n9366), .CLK(n9702), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n1231), .SI(CRC_OUT_5_31), .SE(n9366), .CLK(n9702), 
        .Q(WX6950), .QN(n9049) );
  SDFFX1 DFF_961_Q_reg ( .D(n1232), .SI(WX6950), .SE(n9364), .CLK(n9704), .Q(
        n8470), .QN(n3909) );
  SDFFX1 DFF_962_Q_reg ( .D(n1233), .SI(n8470), .SE(n9364), .CLK(n9704), .Q(
        test_so55), .QN(n3908) );
  SDFFX1 DFF_963_Q_reg ( .D(n1234), .SI(test_si56), .SE(n9364), .CLK(n9704), 
        .Q(n8467), .QN(n3907) );
  SDFFX1 DFF_964_Q_reg ( .D(n1235), .SI(n8467), .SE(n9364), .CLK(n9704), .Q(
        n8466), .QN(n3906) );
  SDFFX1 DFF_965_Q_reg ( .D(n1236), .SI(n8466), .SE(n9364), .CLK(n9704), .Q(
        n8465), .QN(n3905) );
  SDFFX1 DFF_966_Q_reg ( .D(n1237), .SI(n8465), .SE(n9364), .CLK(n9704), .Q(
        n8464), .QN(n3904) );
  SDFFX1 DFF_967_Q_reg ( .D(n1238), .SI(n8464), .SE(n9364), .CLK(n9704), .Q(
        n8463), .QN(n3903) );
  SDFFX1 DFF_968_Q_reg ( .D(n1239), .SI(n8463), .SE(n9364), .CLK(n9704), .Q(
        n8462), .QN(n3902) );
  SDFFX1 DFF_969_Q_reg ( .D(n1240), .SI(n8462), .SE(n9364), .CLK(n9704), .Q(
        n8461), .QN(n3901) );
  SDFFX1 DFF_970_Q_reg ( .D(n1241), .SI(n8461), .SE(n9364), .CLK(n9704), .Q(
        n8460), .QN(n3900) );
  SDFFX1 DFF_971_Q_reg ( .D(n1242), .SI(n8460), .SE(n9364), .CLK(n9704), .Q(
        n8459), .QN(n3899) );
  SDFFX1 DFF_972_Q_reg ( .D(n1243), .SI(n8459), .SE(n9364), .CLK(n9704), .Q(
        n8458), .QN(n3898) );
  SDFFX1 DFF_973_Q_reg ( .D(n1244), .SI(n8458), .SE(n9365), .CLK(n9703), .Q(
        n8457), .QN(n3897) );
  SDFFX1 DFF_974_Q_reg ( .D(n1245), .SI(n8457), .SE(n9365), .CLK(n9703), .Q(
        n8456), .QN(n3896) );
  SDFFX1 DFF_975_Q_reg ( .D(n1246), .SI(n8456), .SE(n9365), .CLK(n9703), .Q(
        n8455), .QN(n3895) );
  SDFFX1 DFF_976_Q_reg ( .D(n1247), .SI(n8455), .SE(n9365), .CLK(n9703), .Q(
        n8454), .QN(n3894) );
  SDFFX1 DFF_977_Q_reg ( .D(n1248), .SI(n8454), .SE(n9365), .CLK(n9703), .Q(
        n8453), .QN(n3893) );
  SDFFX1 DFF_978_Q_reg ( .D(n1249), .SI(n8453), .SE(n9365), .CLK(n9703), .Q(
        n8452), .QN(n3892) );
  SDFFX1 DFF_979_Q_reg ( .D(n1250), .SI(n8452), .SE(n9365), .CLK(n9703), .Q(
        test_so56), .QN(n3891) );
  SDFFX1 DFF_980_Q_reg ( .D(n1251), .SI(test_si57), .SE(n9365), .CLK(n9703), 
        .Q(n8449), .QN(n3890) );
  SDFFX1 DFF_981_Q_reg ( .D(n1252), .SI(n8449), .SE(n9365), .CLK(n9703), .Q(
        n8448), .QN(n3889) );
  SDFFX1 DFF_982_Q_reg ( .D(n1253), .SI(n8448), .SE(n9365), .CLK(n9703), .Q(
        n8447), .QN(n3888) );
  SDFFX1 DFF_983_Q_reg ( .D(n1254), .SI(n8447), .SE(n9365), .CLK(n9703), .Q(
        n8446), .QN(n3887) );
  SDFFX1 DFF_984_Q_reg ( .D(n1255), .SI(n8446), .SE(n9365), .CLK(n9703), .Q(
        n8445), .QN(n3886) );
  SDFFX1 DFF_985_Q_reg ( .D(n1256), .SI(n8445), .SE(n9366), .CLK(n9702), .Q(
        n8444), .QN(n3885) );
  SDFFX1 DFF_986_Q_reg ( .D(n1257), .SI(n8444), .SE(n9366), .CLK(n9702), .Q(
        n8443), .QN(n3884) );
  SDFFX1 DFF_987_Q_reg ( .D(n1258), .SI(n8443), .SE(n9366), .CLK(n9702), .Q(
        n8442), .QN(n3883) );
  SDFFX1 DFF_988_Q_reg ( .D(n1259), .SI(n8442), .SE(n9366), .CLK(n9702), .Q(
        n8441), .QN(n3882) );
  SDFFX1 DFF_989_Q_reg ( .D(n1260), .SI(n8441), .SE(n9366), .CLK(n9702), .Q(
        n8440), .QN(n3881) );
  SDFFX1 DFF_990_Q_reg ( .D(n1261), .SI(n8440), .SE(n9366), .CLK(n9702), .Q(
        n8439), .QN(n3880) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n9366), .CLK(n9702), .Q(
        n8438), .QN(n3879) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n9302), .CLK(n9766), .Q(
        n8437), .QN(n15922) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n9363), .CLK(n9705), .Q(
        n8436), .QN(n15921) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n9363), .CLK(n9705), .Q(
        n8435), .QN(n15920) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n9363), .CLK(n9705), .Q(
        n8434), .QN(n15919) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n9302), .CLK(n9766), .Q(
        test_so57), .QN(n9092) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n9363), .CLK(n9705), 
        .Q(n8431), .QN(n15918) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n9363), .CLK(n9705), .Q(
        n8430), .QN(n15917) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n9362), .CLK(n9706), .Q(
        n8429), .QN(n15916) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n9362), .CLK(n9706), .Q(
        n8428), .QN(n15915) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n9362), .CLK(n9706), .Q(
        n8427), .QN(n15914) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n9362), .CLK(n9706), .Q(
        n8426), .QN(n15913) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n9361), .CLK(n9707), .Q(
        n8425), .QN(n15912) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n9361), .CLK(n9707), .Q(
        n8424), .QN(n15911) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n9361), .CLK(n9707), .Q(
        n8423), .QN(n15910) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n9360), .CLK(n9708), .Q(
        n8422), .QN(n15909) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n9360), .CLK(n9708), .Q(
        n8421), .QN(n15908) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n9360), .CLK(n9708), .Q(
        WX7142), .QN(n8237) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n9359), .CLK(n9709), 
        .Q(WX7144), .QN(n8235) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n9359), .CLK(n9709), 
        .Q(WX7146), .QN(n8233) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n9359), .CLK(n9709), 
        .Q(WX7148), .QN(n8231) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n9358), .CLK(n9710), 
        .Q(WX7150), .QN(n8229) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n9358), .CLK(n9710), 
        .Q(test_so58), .QN(n9122) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n9358), .CLK(n9710), 
        .Q(WX7154), .QN(n8226) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n9357), .CLK(n9711), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n9357), .CLK(n9711), 
        .Q(WX7158), .QN(n8222) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n9357), .CLK(n9711), 
        .Q(WX7160), .QN(n8221) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n9356), .CLK(n9712), 
        .Q(WX7162), .QN(n8219) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n9356), .CLK(n9712), 
        .Q(WX7164), .QN(n8217) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n9356), .CLK(n9712), 
        .Q(WX7166), .QN(n8215) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n9355), .CLK(n9713), 
        .Q(WX7168), .QN(n8213) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n9355), .CLK(n9713), 
        .Q(WX7170), .QN(n8211) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n9355), .CLK(n9713), 
        .Q(WX7172), .QN(n8209) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n9354), .CLK(n9714), 
        .Q(WX7174), .QN(n7882) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n9363), .CLK(n9705), 
        .Q(WX7176), .QN(n8002) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n9363), .CLK(n9705), 
        .Q(WX7178), .QN(n8000) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n9363), .CLK(n9705), 
        .Q(WX7180), .QN(n7998) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n9363), .CLK(n9705), 
        .Q(WX7182), .QN(n7996) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n9363), .CLK(n9705), 
        .Q(WX7184), .QN(n7994) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n9363), .CLK(n9705), 
        .Q(test_so59), .QN(n9124) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n9362), .CLK(n9706), 
        .Q(WX7188), .QN(n7991) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n9362), .CLK(n9706), 
        .Q(WX7190), .QN(n7990) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n9362), .CLK(n9706), 
        .Q(WX7192), .QN(n7988) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n9362), .CLK(n9706), 
        .Q(WX7194), .QN(n7986) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n9361), .CLK(n9707), 
        .Q(WX7196), .QN(n7984) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n9361), .CLK(n9707), 
        .Q(WX7198), .QN(n7982) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n9361), .CLK(n9707), 
        .Q(WX7200), .QN(n7980) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n9360), .CLK(n9708), 
        .Q(WX7202), .QN(n7978) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n9360), .CLK(n9708), 
        .Q(WX7204), .QN(n7976) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n9360), .CLK(n9708), 
        .Q(WX7206) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n9359), .CLK(n9709), 
        .Q(WX7208) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n9359), .CLK(n9709), 
        .Q(WX7210) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n9359), .CLK(n9709), 
        .Q(WX7212) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n9358), .CLK(n9710), 
        .Q(WX7214) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n9358), .CLK(n9710), 
        .Q(WX7216) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n9358), .CLK(n9710), 
        .Q(WX7218) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n9357), .CLK(n9711), 
        .Q(test_so60), .QN(n9121) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n9357), .CLK(n9711), 
        .Q(WX7222) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n9357), .CLK(n9711), 
        .Q(WX7224) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n9356), .CLK(n9712), 
        .Q(WX7226) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n9356), .CLK(n9712), 
        .Q(WX7228) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n9356), .CLK(n9712), 
        .Q(WX7230) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n9355), .CLK(n9713), 
        .Q(WX7232) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n9355), .CLK(n9713), 
        .Q(WX7234) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n9355), .CLK(n9713), 
        .Q(WX7236) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n9354), .CLK(n9714), 
        .Q(WX7238), .QN(n7883) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n9354), .CLK(n9714), 
        .Q(WX7240), .QN(n8003) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n9354), .CLK(n9714), 
        .Q(WX7242), .QN(n8001) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n9354), .CLK(n9714), 
        .Q(WX7244), .QN(n7999) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n9354), .CLK(n9714), 
        .Q(WX7246), .QN(n7997) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n9354), .CLK(n9714), 
        .Q(WX7248), .QN(n7995) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n9363), .CLK(n9705), 
        .Q(WX7250), .QN(n7993) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n9362), .CLK(n9706), 
        .Q(WX7252), .QN(n7992) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n9362), .CLK(n9706), 
        .Q(test_so61), .QN(n9123) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n9362), .CLK(n9706), 
        .Q(WX7256), .QN(n7989) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n9362), .CLK(n9706), 
        .Q(WX7258), .QN(n7987) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n9361), .CLK(n9707), 
        .Q(WX7260), .QN(n7985) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n9361), .CLK(n9707), 
        .Q(WX7262), .QN(n7983) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n9361), .CLK(n9707), 
        .Q(WX7264), .QN(n7981) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n9360), .CLK(n9708), 
        .Q(WX7266), .QN(n7979) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n9360), .CLK(n9708), 
        .Q(WX7268), .QN(n7977) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n9360), .CLK(n9708), 
        .Q(WX7270), .QN(n8238) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n9359), .CLK(n9709), 
        .Q(WX7272), .QN(n8236) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n9359), .CLK(n9709), 
        .Q(WX7274), .QN(n8234) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n9359), .CLK(n9709), 
        .Q(WX7276), .QN(n8232) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n9358), .CLK(n9710), 
        .Q(WX7278), .QN(n8230) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n9358), .CLK(n9710), 
        .Q(WX7280), .QN(n8228) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n9358), .CLK(n9710), 
        .Q(WX7282), .QN(n8227) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n9357), .CLK(n9711), 
        .Q(WX7284), .QN(n8225) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n9357), .CLK(n9711), 
        .Q(WX7286), .QN(n8223) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n9357), .CLK(n9711), 
        .Q(test_so62), .QN(n9120) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n9356), .CLK(n9712), 
        .Q(WX7290), .QN(n8220) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n9356), .CLK(n9712), 
        .Q(WX7292), .QN(n8218) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n9356), .CLK(n9712), 
        .Q(WX7294), .QN(n8216) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n9355), .CLK(n9713), 
        .Q(WX7296), .QN(n8214) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n9355), .CLK(n9713), 
        .Q(WX7298), .QN(n8212) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n9355), .CLK(n9713), 
        .Q(WX7300), .QN(n8210) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n9354), .CLK(n9714), 
        .Q(WX7302), .QN(n8820) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n9354), .CLK(n9714), 
        .Q(WX7304), .QN(n8821) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n9354), .CLK(n9714), 
        .Q(WX7306), .QN(n8822) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n9354), .CLK(n9714), 
        .Q(WX7308), .QN(n8823) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n9354), .CLK(n9714), 
        .Q(WX7310), .QN(n8824) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n9353), .CLK(n9715), 
        .Q(WX7312), .QN(n8825) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n9353), .CLK(n9715), 
        .Q(WX7314), .QN(n8826) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n9353), .CLK(n9715), 
        .Q(WX7316), .QN(n8827) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n9353), .CLK(n9715), 
        .Q(WX7318), .QN(n8828) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n9353), .CLK(n9715), 
        .Q(WX7320), .QN(n8829) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n9353), .CLK(n9715), 
        .Q(test_so63), .QN(n9105) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n9361), .CLK(n9707), 
        .Q(WX7324), .QN(n8830) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n9361), .CLK(n9707), 
        .Q(WX7326), .QN(n8831) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n9361), .CLK(n9707), 
        .Q(WX7328), .QN(n8832) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n9360), .CLK(n9708), 
        .Q(WX7330), .QN(n8833) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n9360), .CLK(n9708), 
        .Q(WX7332), .QN(n8722) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n9360), .CLK(n9708), 
        .Q(WX7334), .QN(n8834) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n9359), .CLK(n9709), 
        .Q(WX7336), .QN(n8835) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n9359), .CLK(n9709), 
        .Q(WX7338), .QN(n8836) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n9359), .CLK(n9709), 
        .Q(WX7340), .QN(n8837) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n9358), .CLK(n9710), 
        .Q(WX7342), .QN(n8723) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n9358), .CLK(n9710), 
        .Q(WX7344), .QN(n8838) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n9358), .CLK(n9710), 
        .Q(WX7346), .QN(n8839) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n9357), .CLK(n9711), 
        .Q(WX7348), .QN(n8840) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n9357), .CLK(n9711), 
        .Q(WX7350), .QN(n8841) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n9357), .CLK(n9711), 
        .Q(WX7352), .QN(n8842) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n9356), .CLK(n9712), 
        .Q(WX7354), .QN(n8843) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n9356), .CLK(n9712), 
        .Q(test_so64), .QN(n9087) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n9356), .CLK(n9712), 
        .Q(WX7358), .QN(n8844) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n9355), .CLK(n9713), 
        .Q(WX7360), .QN(n8845) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n9355), .CLK(n9713), 
        .Q(WX7362), .QN(n8846) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n9355), .CLK(n9713), 
        .Q(WX7364), .QN(n8737) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n9304), .CLK(n9764), 
        .Q(CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_3), .QN(DFF_1123_n1) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n9304), .CLK(n9764), .Q(CRC_OUT_4_10), .QN(DFF_1130_n1) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n9304), .CLK(
        n9764), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n9303), .CLK(
        n9765), .Q(test_so65), .QN(n9153) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n9303), .CLK(n9765), 
        .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_15), .QN(DFF_1135_n1) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n9303), .CLK(
        n9765), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n9302), .CLK(
        n9766), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n9302), .CLK(
        n9766), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n9353), .CLK(
        n9715), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n9353), .CLK(
        n9715), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n9353), .CLK(
        n9715), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n9353), .CLK(
        n9715), .Q(test_so66), .QN(n9152) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n9353), .CLK(n9715), 
        .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n9353), .CLK(
        n9715), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n1472), .SI(CRC_OUT_4_31), .SE(n9352), .CLK(n9716), .Q(WX8243), .QN(n9050) );
  SDFFX1 DFF_1153_Q_reg ( .D(n1473), .SI(WX8243), .SE(n9350), .CLK(n9718), .Q(
        n8411), .QN(n3878) );
  SDFFX1 DFF_1154_Q_reg ( .D(n1474), .SI(n8411), .SE(n9350), .CLK(n9718), .Q(
        n8410), .QN(n3877) );
  SDFFX1 DFF_1155_Q_reg ( .D(n1475), .SI(n8410), .SE(n9350), .CLK(n9718), .Q(
        n8409), .QN(n3876) );
  SDFFX1 DFF_1156_Q_reg ( .D(n1476), .SI(n8409), .SE(n9350), .CLK(n9718), .Q(
        n8408), .QN(n3875) );
  SDFFX1 DFF_1157_Q_reg ( .D(n1477), .SI(n8408), .SE(n9350), .CLK(n9718), .Q(
        n8407), .QN(n3874) );
  SDFFX1 DFF_1158_Q_reg ( .D(n1478), .SI(n8407), .SE(n9350), .CLK(n9718), .Q(
        n8406), .QN(n3873) );
  SDFFX1 DFF_1159_Q_reg ( .D(n1479), .SI(n8406), .SE(n9350), .CLK(n9718), .Q(
        n8405), .QN(n3872) );
  SDFFX1 DFF_1160_Q_reg ( .D(n1480), .SI(n8405), .SE(n9350), .CLK(n9718), .Q(
        n8404), .QN(n3871) );
  SDFFX1 DFF_1161_Q_reg ( .D(n1481), .SI(n8404), .SE(n9351), .CLK(n9717), .Q(
        n8403), .QN(n3870) );
  SDFFX1 DFF_1162_Q_reg ( .D(n1482), .SI(n8403), .SE(n9351), .CLK(n9717), .Q(
        n8402), .QN(n3869) );
  SDFFX1 DFF_1163_Q_reg ( .D(n1483), .SI(n8402), .SE(n9351), .CLK(n9717), .Q(
        n8401), .QN(n3868) );
  SDFFX1 DFF_1164_Q_reg ( .D(n1484), .SI(n8401), .SE(n9351), .CLK(n9717), .Q(
        n8400), .QN(n3867) );
  SDFFX1 DFF_1165_Q_reg ( .D(n1485), .SI(n8400), .SE(n9351), .CLK(n9717), .Q(
        n8399), .QN(n3866) );
  SDFFX1 DFF_1166_Q_reg ( .D(n1486), .SI(n8399), .SE(n9351), .CLK(n9717), .Q(
        test_so67), .QN(n3865) );
  SDFFX1 DFF_1167_Q_reg ( .D(n1487), .SI(test_si68), .SE(n9351), .CLK(n9717), 
        .Q(n8396), .QN(n3864) );
  SDFFX1 DFF_1168_Q_reg ( .D(n1488), .SI(n8396), .SE(n9351), .CLK(n9717), .Q(
        n8395), .QN(n3863) );
  SDFFX1 DFF_1169_Q_reg ( .D(n1489), .SI(n8395), .SE(n9351), .CLK(n9717), .Q(
        n8394), .QN(n3862) );
  SDFFX1 DFF_1170_Q_reg ( .D(n1490), .SI(n8394), .SE(n9351), .CLK(n9717), .Q(
        n8393), .QN(n3861) );
  SDFFX1 DFF_1171_Q_reg ( .D(n1491), .SI(n8393), .SE(n9351), .CLK(n9717), .Q(
        n8392), .QN(n3860) );
  SDFFX1 DFF_1172_Q_reg ( .D(n1492), .SI(n8392), .SE(n9351), .CLK(n9717), .Q(
        n8391), .QN(n3859) );
  SDFFX1 DFF_1173_Q_reg ( .D(n1493), .SI(n8391), .SE(n9352), .CLK(n9716), .Q(
        n8390), .QN(n3858) );
  SDFFX1 DFF_1174_Q_reg ( .D(n1494), .SI(n8390), .SE(n9352), .CLK(n9716), .Q(
        n8389), .QN(n3857) );
  SDFFX1 DFF_1175_Q_reg ( .D(n1495), .SI(n8389), .SE(n9352), .CLK(n9716), .Q(
        n8388), .QN(n3856) );
  SDFFX1 DFF_1176_Q_reg ( .D(n1496), .SI(n8388), .SE(n9352), .CLK(n9716), .Q(
        n8387), .QN(n3855) );
  SDFFX1 DFF_1177_Q_reg ( .D(n1497), .SI(n8387), .SE(n9352), .CLK(n9716), .Q(
        n8386), .QN(n3854) );
  SDFFX1 DFF_1178_Q_reg ( .D(n1498), .SI(n8386), .SE(n9352), .CLK(n9716), .Q(
        n8385), .QN(n3853) );
  SDFFX1 DFF_1179_Q_reg ( .D(n1499), .SI(n8385), .SE(n9352), .CLK(n9716), .Q(
        n8384), .QN(n3852) );
  SDFFX1 DFF_1180_Q_reg ( .D(n1500), .SI(n8384), .SE(n9352), .CLK(n9716), .Q(
        n8383), .QN(n3851) );
  SDFFX1 DFF_1181_Q_reg ( .D(n1501), .SI(n8383), .SE(n9352), .CLK(n9716), .Q(
        n8382), .QN(n3850) );
  SDFFX1 DFF_1182_Q_reg ( .D(n1502), .SI(n8382), .SE(n9352), .CLK(n9716), .Q(
        n8381), .QN(n3849) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n9352), .CLK(n9716), .Q(
        test_so68), .QN(n3848) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n9305), .CLK(n9763), 
        .Q(n8378), .QN(n15907) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n9350), .CLK(n9718), .Q(
        n8377), .QN(n15906) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n9349), .CLK(n9719), .Q(
        n8376), .QN(n15905) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n9349), .CLK(n9719), .Q(
        n8375), .QN(n15904) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n9349), .CLK(n9719), .Q(
        n8374), .QN(n15903) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n9349), .CLK(n9719), .Q(
        n8373), .QN(n15902) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n9349), .CLK(n9719), .Q(
        n8372), .QN(n15901) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n9348), .CLK(n9720), .Q(
        n8371), .QN(n15900) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n9348), .CLK(n9720), .Q(
        n8370), .QN(n15899) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n9347), .CLK(n9721), .Q(
        n8369), .QN(n15898) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n9347), .CLK(n9721), .Q(
        n8368), .QN(n15897) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n9347), .CLK(n9721), .Q(
        n8367), .QN(n15896) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n9347), .CLK(n9721), .Q(
        n8366), .QN(n15895) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n9346), .CLK(n9722), .Q(
        n8365), .QN(n15894) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n9346), .CLK(n9722), .Q(
        n8364), .QN(n15893) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n9345), .CLK(n9723), .Q(
        n8363), .QN(n15892) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n9345), .CLK(n9723), .Q(
        test_so69), .QN(n9117) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n9345), .CLK(n9723), 
        .Q(WX8437), .QN(n8206) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n9345), .CLK(n9723), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n9344), .CLK(n9724), 
        .Q(WX8441), .QN(n8202) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n9344), .CLK(n9724), 
        .Q(WX8443), .QN(n8201) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n9344), .CLK(n9724), 
        .Q(WX8445), .QN(n8199) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n9343), .CLK(n9725), 
        .Q(WX8447), .QN(n8197) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n9343), .CLK(n9725), 
        .Q(WX8449), .QN(n8195) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n9343), .CLK(n9725), 
        .Q(WX8451), .QN(n8193) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n9342), .CLK(n9726), 
        .Q(WX8453), .QN(n8191) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n9342), .CLK(n9726), 
        .Q(WX8455), .QN(n8189) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n9342), .CLK(n9726), 
        .Q(WX8457), .QN(n8187) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n9341), .CLK(n9727), 
        .Q(WX8459), .QN(n8185) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n9341), .CLK(n9727), 
        .Q(WX8461), .QN(n8183) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n9341), .CLK(n9727), 
        .Q(WX8463), .QN(n8181) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n9340), .CLK(n9728), 
        .Q(WX8465), .QN(n8179) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n9340), .CLK(n9728), 
        .Q(WX8467), .QN(n7880) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n9350), .CLK(n9718), 
        .Q(test_so70), .QN(n9119) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n9349), .CLK(n9719), 
        .Q(WX8471), .QN(n7973) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n9349), .CLK(n9719), 
        .Q(WX8473), .QN(n7972) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n9349), .CLK(n9719), 
        .Q(WX8475), .QN(n7970) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n9349), .CLK(n9719), 
        .Q(WX8477), .QN(n7968) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n9348), .CLK(n9720), 
        .Q(WX8479), .QN(n7966) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n9348), .CLK(n9720), 
        .Q(WX8481), .QN(n7964) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n9348), .CLK(n9720), 
        .Q(WX8483), .QN(n7962) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n9348), .CLK(n9720), 
        .Q(WX8485), .QN(n7960) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n9347), .CLK(n9721), 
        .Q(WX8487), .QN(n7958) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n9347), .CLK(n9721), 
        .Q(WX8489), .QN(n7956) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n9346), .CLK(n9722), 
        .Q(WX8491), .QN(n7954) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n9346), .CLK(n9722), 
        .Q(WX8493), .QN(n7952) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n9346), .CLK(n9722), 
        .Q(WX8495), .QN(n7950) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n9346), .CLK(n9722), 
        .Q(WX8497), .QN(n7948) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n9345), .CLK(n9723), 
        .Q(WX8499) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n9345), .CLK(n9723), 
        .Q(WX8501) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n9344), .CLK(n9724), 
        .Q(test_so71), .QN(n9116) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n9344), .CLK(n9724), 
        .Q(WX8505) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n9344), .CLK(n9724), 
        .Q(WX8507) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n9343), .CLK(n9725), 
        .Q(WX8509) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n9343), .CLK(n9725), 
        .Q(WX8511) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n9343), .CLK(n9725), 
        .Q(WX8513) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n9342), .CLK(n9726), 
        .Q(WX8515) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n9342), .CLK(n9726), 
        .Q(WX8517) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n9342), .CLK(n9726), 
        .Q(WX8519) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n9341), .CLK(n9727), 
        .Q(WX8521) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n9341), .CLK(n9727), 
        .Q(WX8523) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n9341), .CLK(n9727), 
        .Q(WX8525) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n9340), .CLK(n9728), 
        .Q(WX8527) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n9340), .CLK(n9728), 
        .Q(WX8529) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n9340), .CLK(n9728), 
        .Q(WX8531), .QN(n7881) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n9350), .CLK(n9718), 
        .Q(WX8533), .QN(n7975) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n9350), .CLK(n9718), 
        .Q(WX8535), .QN(n7974) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n9349), .CLK(n9719), 
        .Q(test_so72), .QN(n9118) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n9349), .CLK(n9719), 
        .Q(WX8539), .QN(n7971) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n9349), .CLK(n9719), 
        .Q(WX8541), .QN(n7969) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n9348), .CLK(n9720), 
        .Q(WX8543), .QN(n7967) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n9348), .CLK(n9720), 
        .Q(WX8545), .QN(n7965) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n9348), .CLK(n9720), 
        .Q(WX8547), .QN(n7963) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n9347), .CLK(n9721), 
        .Q(WX8549), .QN(n7961) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n9347), .CLK(n9721), 
        .Q(WX8551), .QN(n7959) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n9347), .CLK(n9721), 
        .Q(WX8553), .QN(n7957) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n9346), .CLK(n9722), 
        .Q(WX8555), .QN(n7955) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n9346), .CLK(n9722), 
        .Q(WX8557), .QN(n7953) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n9346), .CLK(n9722), 
        .Q(WX8559), .QN(n7951) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n9345), .CLK(n9723), 
        .Q(WX8561), .QN(n7949) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n9345), .CLK(n9723), 
        .Q(WX8563), .QN(n8208) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n9345), .CLK(n9723), 
        .Q(WX8565), .QN(n8207) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n9344), .CLK(n9724), 
        .Q(WX8567), .QN(n8205) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n9344), .CLK(n9724), 
        .Q(WX8569), .QN(n8203) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n9344), .CLK(n9724), 
        .Q(test_so73), .QN(n9115) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n9343), .CLK(n9725), 
        .Q(WX8573), .QN(n8200) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n9343), .CLK(n9725), 
        .Q(WX8575), .QN(n8198) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n9343), .CLK(n9725), 
        .Q(WX8577), .QN(n8196) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n9342), .CLK(n9726), 
        .Q(WX8579), .QN(n8194) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n9342), .CLK(n9726), 
        .Q(WX8581), .QN(n8192) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n9342), .CLK(n9726), 
        .Q(WX8583), .QN(n8190) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n9341), .CLK(n9727), 
        .Q(WX8585), .QN(n8188) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n9341), .CLK(n9727), 
        .Q(WX8587), .QN(n8186) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n9341), .CLK(n9727), 
        .Q(WX8589), .QN(n8184) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n9340), .CLK(n9728), 
        .Q(WX8591), .QN(n8182) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n9340), .CLK(n9728), 
        .Q(WX8593), .QN(n8180) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n9340), .CLK(n9728), 
        .Q(WX8595), .QN(n8794) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n9340), .CLK(n9728), 
        .Q(WX8597), .QN(n8795) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n9340), .CLK(n9728), 
        .Q(WX8599), .QN(n8796) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n9339), .CLK(n9729), 
        .Q(WX8601), .QN(n8797) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n9339), .CLK(n9729), 
        .Q(WX8603), .QN(n8798) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n9339), .CLK(n9729), 
        .Q(test_so74), .QN(n9104) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n9348), .CLK(n9720), 
        .Q(WX8607), .QN(n8799) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n9348), .CLK(n9720), 
        .Q(WX8609), .QN(n8800) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n9348), .CLK(n9720), 
        .Q(WX8611), .QN(n8801) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n9347), .CLK(n9721), 
        .Q(WX8613), .QN(n8802) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n9347), .CLK(n9721), 
        .Q(WX8615), .QN(n8803) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n9347), .CLK(n9721), 
        .Q(WX8617), .QN(n8804) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n9346), .CLK(n9722), 
        .Q(WX8619), .QN(n8805) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n9346), .CLK(n9722), 
        .Q(WX8621), .QN(n8806) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n9346), .CLK(n9722), 
        .Q(WX8623), .QN(n8807) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n9345), .CLK(n9723), 
        .Q(WX8625), .QN(n8719) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n9345), .CLK(n9723), 
        .Q(WX8627), .QN(n8808) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n9345), .CLK(n9723), 
        .Q(WX8629), .QN(n8809) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n9344), .CLK(n9724), 
        .Q(WX8631), .QN(n8810) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n9344), .CLK(n9724), 
        .Q(WX8633), .QN(n8811) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n9344), .CLK(n9724), 
        .Q(WX8635), .QN(n8720) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n9343), .CLK(n9725), 
        .Q(WX8637), .QN(n8812) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n9343), .CLK(n9725), 
        .Q(test_so75), .QN(n9099) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n9343), .CLK(n9725), 
        .Q(WX8641), .QN(n8813) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n9342), .CLK(n9726), 
        .Q(WX8643), .QN(n8814) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n9342), .CLK(n9726), 
        .Q(WX8645), .QN(n8815) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n9342), .CLK(n9726), 
        .Q(WX8647), .QN(n8816) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n9341), .CLK(n9727), 
        .Q(WX8649), .QN(n8721) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n9341), .CLK(n9727), 
        .Q(WX8651), .QN(n8817) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n9341), .CLK(n9727), 
        .Q(WX8653), .QN(n8818) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n9340), .CLK(n9728), 
        .Q(WX8655), .QN(n8819) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n9340), .CLK(n9728), 
        .Q(WX8657), .QN(n8736) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n9307), .CLK(n9761), 
        .Q(CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n9307), .CLK(n9761), .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n9307), .CLK(n9761), .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n9307), .CLK(n9761), .Q(CRC_OUT_3_3), .QN(DFF_1315_n1) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n9307), .CLK(n9761), .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n9307), .CLK(n9761), .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n9307), .CLK(n9761), .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n9307), .CLK(n9761), .Q(test_so76), .QN(n9151) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n9306), .CLK(n9762), 
        .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n9306), .CLK(n9762), .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n9306), .CLK(n9762), .Q(CRC_OUT_3_10), .QN(DFF_1322_n1) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n9306), .CLK(
        n9762), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n9306), .CLK(
        n9762), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n9306), .CLK(
        n9762), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n9306), .CLK(
        n9762), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n9306), .CLK(
        n9762), .Q(CRC_OUT_3_15), .QN(DFF_1327_n1) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n9306), .CLK(
        n9762), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n9306), .CLK(
        n9762), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n9306), .CLK(
        n9762), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n9306), .CLK(
        n9762), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n9305), .CLK(
        n9763), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n9305), .CLK(
        n9763), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n9305), .CLK(
        n9763), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n9305), .CLK(
        n9763), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n9305), .CLK(
        n9763), .Q(test_so77), .QN(n9150) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n9305), .CLK(n9763), 
        .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n9305), .CLK(
        n9763), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n9305), .CLK(
        n9763), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n9305), .CLK(
        n9763), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n9305), .CLK(
        n9763), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n9305), .CLK(
        n9763), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n9339), .CLK(
        n9729), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n1714), .SI(CRC_OUT_3_31), .SE(n9339), .CLK(n9729), .Q(WX9536), .QN(n9051) );
  SDFFX1 DFF_1345_Q_reg ( .D(n1715), .SI(WX9536), .SE(n9337), .CLK(n9731), .Q(
        n8353), .QN(n3847) );
  SDFFX1 DFF_1346_Q_reg ( .D(n1716), .SI(n8353), .SE(n9337), .CLK(n9731), .Q(
        n8352), .QN(n3846) );
  SDFFX1 DFF_1347_Q_reg ( .D(n1717), .SI(n8352), .SE(n9337), .CLK(n9731), .Q(
        n8351), .QN(n3845) );
  SDFFX1 DFF_1348_Q_reg ( .D(n1718), .SI(n8351), .SE(n9337), .CLK(n9731), .Q(
        n8350), .QN(n3844) );
  SDFFX1 DFF_1349_Q_reg ( .D(n1719), .SI(n8350), .SE(n9337), .CLK(n9731), .Q(
        n8349), .QN(n3843) );
  SDFFX1 DFF_1350_Q_reg ( .D(n1720), .SI(n8349), .SE(n9337), .CLK(n9731), .Q(
        n8348), .QN(n3842) );
  SDFFX1 DFF_1351_Q_reg ( .D(n1721), .SI(n8348), .SE(n9337), .CLK(n9731), .Q(
        n8347), .QN(n3841) );
  SDFFX1 DFF_1352_Q_reg ( .D(n1722), .SI(n8347), .SE(n9337), .CLK(n9731), .Q(
        n8346), .QN(n3840) );
  SDFFX1 DFF_1353_Q_reg ( .D(n1723), .SI(n8346), .SE(n9337), .CLK(n9731), .Q(
        test_so78), .QN(n3839) );
  SDFFX1 DFF_1354_Q_reg ( .D(n1724), .SI(test_si79), .SE(n9337), .CLK(n9731), 
        .Q(n8343), .QN(n3838) );
  SDFFX1 DFF_1355_Q_reg ( .D(n1725), .SI(n8343), .SE(n9337), .CLK(n9731), .Q(
        n8342), .QN(n3837) );
  SDFFX1 DFF_1356_Q_reg ( .D(n1726), .SI(n8342), .SE(n9337), .CLK(n9731), .Q(
        n8341), .QN(n3836) );
  SDFFX1 DFF_1357_Q_reg ( .D(n1727), .SI(n8341), .SE(n9338), .CLK(n9730), .Q(
        n8340), .QN(n3835) );
  SDFFX1 DFF_1358_Q_reg ( .D(n1728), .SI(n8340), .SE(n9338), .CLK(n9730), .Q(
        n8339), .QN(n3834) );
  SDFFX1 DFF_1359_Q_reg ( .D(n1729), .SI(n8339), .SE(n9338), .CLK(n9730), .Q(
        n8338), .QN(n3833) );
  SDFFX1 DFF_1360_Q_reg ( .D(n1730), .SI(n8338), .SE(n9338), .CLK(n9730), .Q(
        n8337), .QN(n3832) );
  SDFFX1 DFF_1361_Q_reg ( .D(n1731), .SI(n8337), .SE(n9338), .CLK(n9730), .Q(
        n8336), .QN(n3831) );
  SDFFX1 DFF_1362_Q_reg ( .D(n1732), .SI(n8336), .SE(n9338), .CLK(n9730), .Q(
        n8335), .QN(n3830) );
  SDFFX1 DFF_1363_Q_reg ( .D(n1733), .SI(n8335), .SE(n9338), .CLK(n9730), .Q(
        n8334), .QN(n3829) );
  SDFFX1 DFF_1364_Q_reg ( .D(n1734), .SI(n8334), .SE(n9338), .CLK(n9730), .Q(
        n8333), .QN(n3828) );
  SDFFX1 DFF_1365_Q_reg ( .D(n1735), .SI(n8333), .SE(n9338), .CLK(n9730), .Q(
        n8332), .QN(n3827) );
  SDFFX1 DFF_1366_Q_reg ( .D(n1736), .SI(n8332), .SE(n9338), .CLK(n9730), .Q(
        n8331), .QN(n3826) );
  SDFFX1 DFF_1367_Q_reg ( .D(n1737), .SI(n8331), .SE(n9338), .CLK(n9730), .Q(
        n8330), .QN(n3825) );
  SDFFX1 DFF_1368_Q_reg ( .D(n1738), .SI(n8330), .SE(n9338), .CLK(n9730), .Q(
        n8329), .QN(n3824) );
  SDFFX1 DFF_1369_Q_reg ( .D(n1739), .SI(n8329), .SE(n9339), .CLK(n9729), .Q(
        n8328), .QN(n3823) );
  SDFFX1 DFF_1370_Q_reg ( .D(n1740), .SI(n8328), .SE(n9339), .CLK(n9729), .Q(
        test_so79), .QN(n3822) );
  SDFFX1 DFF_1371_Q_reg ( .D(n1741), .SI(test_si80), .SE(n9339), .CLK(n9729), 
        .Q(n8325), .QN(n3821) );
  SDFFX1 DFF_1372_Q_reg ( .D(n1742), .SI(n8325), .SE(n9339), .CLK(n9729), .Q(
        n8324), .QN(n3820) );
  SDFFX1 DFF_1373_Q_reg ( .D(n1743), .SI(n8324), .SE(n9339), .CLK(n9729), .Q(
        n8323), .QN(n3819) );
  SDFFX1 DFF_1374_Q_reg ( .D(n1744), .SI(n8323), .SE(n9339), .CLK(n9729), .Q(
        n8322), .QN(n3818) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n9339), .CLK(n9729), .Q(
        n8321), .QN(n3817) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n9307), .CLK(n9761), .Q(
        n8320), .QN(n15891) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n9336), .CLK(n9732), .Q(
        n8319), .QN(n15890) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n9336), .CLK(n9732), .Q(
        n8318), .QN(n15889) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n9336), .CLK(n9732), .Q(
        n8317), .QN(n15888) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n9336), .CLK(n9732), .Q(
        n8316), .QN(n15887) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n9336), .CLK(n9732), .Q(
        n8315), .QN(n15886) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n9336), .CLK(n9732), .Q(
        n8314), .QN(n15885) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n9335), .CLK(n9733), .Q(
        n8313), .QN(n15884) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n9335), .CLK(n9733), .Q(
        n8312), .QN(n15883) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n9335), .CLK(n9733), .Q(
        n8311), .QN(n15882) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n9335), .CLK(n9733), .Q(
        n8310), .QN(n15881) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n9335), .CLK(n9733), .Q(
        test_so80), .QN(n9091) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n9335), .CLK(n9733), 
        .Q(n8307), .QN(n15880) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n9334), .CLK(n9734), .Q(
        n8306), .QN(n15879) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n9334), .CLK(n9734), .Q(
        n8305), .QN(n15878) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n9334), .CLK(n9734), .Q(
        n8304), .QN(n15877) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n9334), .CLK(n9734), .Q(
        WX9728), .QN(n8177) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n9333), .CLK(n9735), 
        .Q(WX9730), .QN(n8175) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n9333), .CLK(n9735), 
        .Q(WX9732), .QN(n8173) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n9333), .CLK(n9735), 
        .Q(WX9734), .QN(n8171) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n9333), .CLK(n9735), 
        .Q(WX9736), .QN(n8169) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n9332), .CLK(n9736), 
        .Q(WX9738), .QN(n8167) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n9332), .CLK(n9736), 
        .Q(WX9740), .QN(n8165) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n9332), .CLK(n9736), 
        .Q(WX9742), .QN(n8163) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n9331), .CLK(n9737), 
        .Q(WX9744), .QN(n8161) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n9331), .CLK(n9737), 
        .Q(WX9746), .QN(n8159) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n9331), .CLK(n9737), 
        .Q(WX9748), .QN(n8157) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n9330), .CLK(n9738), 
        .Q(WX9750), .QN(n8155) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n9330), .CLK(n9738), 
        .Q(test_so81), .QN(n9112) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n9329), .CLK(n9739), 
        .Q(WX9754), .QN(n8152) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n9329), .CLK(n9739), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n9329), .CLK(n9739), 
        .Q(WX9758), .QN(n8148) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n9329), .CLK(n9739), 
        .Q(WX9760), .QN(n7878) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n9336), .CLK(n9732), 
        .Q(WX9762), .QN(n7946) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n9336), .CLK(n9732), 
        .Q(WX9764), .QN(n7944) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n9336), .CLK(n9732), 
        .Q(WX9766), .QN(n7942) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n9336), .CLK(n9732), 
        .Q(WX9768), .QN(n7940) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n9336), .CLK(n9732), 
        .Q(WX9770), .QN(n7938) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n9336), .CLK(n9732), 
        .Q(WX9772), .QN(n7936) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n9335), .CLK(n9733), 
        .Q(WX9774), .QN(n7934) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n9335), .CLK(n9733), 
        .Q(WX9776), .QN(n7932) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n9335), .CLK(n9733), 
        .Q(WX9778), .QN(n7930) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n9335), .CLK(n9733), 
        .Q(WX9780), .QN(n7928) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n9335), .CLK(n9733), 
        .Q(WX9782), .QN(n7926) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n9335), .CLK(n9733), 
        .Q(WX9784), .QN(n7924) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n9334), .CLK(n9734), 
        .Q(test_so82), .QN(n9114) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n9334), .CLK(n9734), 
        .Q(WX9788), .QN(n7921) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n9334), .CLK(n9734), 
        .Q(WX9790), .QN(n7920) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n9334), .CLK(n9734), 
        .Q(WX9792) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n9333), .CLK(n9735), 
        .Q(WX9794) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n9333), .CLK(n9735), 
        .Q(WX9796) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n9333), .CLK(n9735), 
        .Q(WX9798) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n9332), .CLK(n9736), 
        .Q(WX9800) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n9332), .CLK(n9736), 
        .Q(WX9802) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n9332), .CLK(n9736), 
        .Q(WX9804) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n9331), .CLK(n9737), 
        .Q(WX9806) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n9331), .CLK(n9737), 
        .Q(WX9808) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n9331), .CLK(n9737), 
        .Q(WX9810) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n9330), .CLK(n9738), 
        .Q(WX9812) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n9330), .CLK(n9738), 
        .Q(WX9814) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n9330), .CLK(n9738), 
        .Q(WX9816) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n9330), .CLK(n9738), 
        .Q(WX9818) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n9329), .CLK(n9739), 
        .Q(test_so83), .QN(n9111) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n9329), .CLK(n9739), 
        .Q(WX9822) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n9328), .CLK(n9740), 
        .Q(WX9824), .QN(n7879) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n9328), .CLK(n9740), 
        .Q(WX9826), .QN(n7947) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n9328), .CLK(n9740), 
        .Q(WX9828), .QN(n7945) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n9328), .CLK(n9740), 
        .Q(WX9830), .QN(n7943) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n9328), .CLK(n9740), 
        .Q(WX9832), .QN(n7941) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n9328), .CLK(n9740), 
        .Q(WX9834), .QN(n7939) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n9327), .CLK(n9741), 
        .Q(WX9836), .QN(n7937) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n9327), .CLK(n9741), 
        .Q(WX9838), .QN(n7935) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n9327), .CLK(n9741), 
        .Q(WX9840), .QN(n7933) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n9327), .CLK(n9741), 
        .Q(WX9842), .QN(n7931) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n9327), .CLK(n9741), 
        .Q(WX9844), .QN(n7929) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n9327), .CLK(n9741), 
        .Q(WX9846), .QN(n7927) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n9326), .CLK(n9742), 
        .Q(WX9848), .QN(n7925) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n9334), .CLK(n9734), 
        .Q(WX9850), .QN(n7923) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n9334), .CLK(n9734), 
        .Q(WX9852), .QN(n7922) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n9334), .CLK(n9734), 
        .Q(test_so84), .QN(n9113) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n9334), .CLK(n9734), 
        .Q(WX9856), .QN(n8178) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n9333), .CLK(n9735), 
        .Q(WX9858), .QN(n8176) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n9333), .CLK(n9735), 
        .Q(WX9860), .QN(n8174) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n9333), .CLK(n9735), 
        .Q(WX9862), .QN(n8172) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n9332), .CLK(n9736), 
        .Q(WX9864), .QN(n8170) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n9332), .CLK(n9736), 
        .Q(WX9866), .QN(n8168) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n9332), .CLK(n9736), 
        .Q(WX9868), .QN(n8166) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n9331), .CLK(n9737), 
        .Q(WX9870), .QN(n8164) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n9331), .CLK(n9737), 
        .Q(WX9872), .QN(n8162) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n9331), .CLK(n9737), 
        .Q(WX9874), .QN(n8160) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n9330), .CLK(n9738), 
        .Q(WX9876), .QN(n8158) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n9330), .CLK(n9738), 
        .Q(WX9878), .QN(n8156) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n9330), .CLK(n9738), 
        .Q(WX9880), .QN(n8154) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n9329), .CLK(n9739), 
        .Q(WX9882), .QN(n8153) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n9329), .CLK(n9739), 
        .Q(WX9884), .QN(n8151) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n9329), .CLK(n9739), 
        .Q(WX9886), .QN(n8149) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n9328), .CLK(n9740), 
        .Q(test_so85), .QN(n9110) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n9328), .CLK(n9740), 
        .Q(WX9890), .QN(n8768) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n9328), .CLK(n9740), 
        .Q(WX9892), .QN(n8769) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n9328), .CLK(n9740), 
        .Q(WX9894), .QN(n8770) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n9328), .CLK(n9740), 
        .Q(WX9896), .QN(n8771) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n9328), .CLK(n9740), 
        .Q(WX9898), .QN(n8772) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n9327), .CLK(n9741), 
        .Q(WX9900), .QN(n8773) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n9327), .CLK(n9741), 
        .Q(WX9902), .QN(n8774) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n9327), .CLK(n9741), 
        .Q(WX9904), .QN(n8775) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n9327), .CLK(n9741), 
        .Q(WX9906), .QN(n8776) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n9327), .CLK(n9741), 
        .Q(WX9908), .QN(n8777) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n9327), .CLK(n9741), 
        .Q(WX9910), .QN(n8778) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n9326), .CLK(n9742), 
        .Q(WX9912), .QN(n8779) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n9326), .CLK(n9742), 
        .Q(WX9914), .QN(n8780) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n9326), .CLK(n9742), 
        .Q(WX9916), .QN(n8781) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n9326), .CLK(n9742), 
        .Q(WX9918), .QN(n8716) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n9326), .CLK(n9742), 
        .Q(WX9920), .QN(n8782) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n9326), .CLK(n9742), 
        .Q(test_so86), .QN(n9103) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n9333), .CLK(n9735), 
        .Q(WX9924), .QN(n8783) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n9333), .CLK(n9735), 
        .Q(WX9926), .QN(n8784) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n9332), .CLK(n9736), 
        .Q(WX9928), .QN(n8717) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n9332), .CLK(n9736), 
        .Q(WX9930), .QN(n8785) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n9332), .CLK(n9736), 
        .Q(WX9932), .QN(n8786) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n9331), .CLK(n9737), 
        .Q(WX9934), .QN(n8787) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n9331), .CLK(n9737), 
        .Q(WX9936), .QN(n8788) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n9331), .CLK(n9737), 
        .Q(WX9938), .QN(n8789) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n9330), .CLK(n9738), 
        .Q(WX9940), .QN(n8790) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n9330), .CLK(n9738), 
        .Q(WX9942), .QN(n8718) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n9330), .CLK(n9738), 
        .Q(WX9944), .QN(n8791) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n9329), .CLK(n9739), 
        .Q(WX9946), .QN(n8792) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n9329), .CLK(n9739), 
        .Q(WX9948), .QN(n8793) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n9329), .CLK(n9739), 
        .Q(WX9950), .QN(n8735) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n9309), .CLK(n9759), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n9309), .CLK(
        n9759), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n9309), .CLK(
        n9759), .Q(test_so87), .QN(n9165) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n9309), .CLK(n9759), 
        .Q(CRC_OUT_2_3), .QN(DFF_1507_n1) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_10), .QN(DFF_1514_n1) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n9308), .CLK(
        n9760), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n9307), .CLK(
        n9761), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n9307), .CLK(
        n9761), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n9307), .CLK(
        n9761), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n9326), .CLK(
        n9742), .Q(test_so88), .QN(n9164) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n9326), .CLK(n9742), 
        .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n9326), .CLK(
        n9742), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n9326), .CLK(
        n9742), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n9326), .CLK(
        n9742), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n9325), .CLK(
        n9743), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n9325), .CLK(
        n9743), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n9325), .CLK(
        n9743), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n9325), .CLK(
        n9743), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n9325), .CLK(
        n9743), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n9325), .CLK(
        n9743), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n9325), .CLK(
        n9743), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n9325), .CLK(
        n9743), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(n1955), .SI(CRC_OUT_2_31), .SE(n9325), .CLK(n9743), .Q(WX10829), .QN(n9052) );
  SDFFX1 DFF_1537_Q_reg ( .D(n1956), .SI(WX10829), .SE(n9322), .CLK(n9746), 
        .Q(n8295), .QN(n3816) );
  SDFFX1 DFF_1538_Q_reg ( .D(n1957), .SI(n8295), .SE(n9322), .CLK(n9746), .Q(
        n8294), .QN(n3815) );
  SDFFX1 DFF_1539_Q_reg ( .D(n1958), .SI(n8294), .SE(n9322), .CLK(n9746), .Q(
        n8293), .QN(n3814) );
  SDFFX1 DFF_1540_Q_reg ( .D(n1959), .SI(n8293), .SE(n9322), .CLK(n9746), .Q(
        test_so89), .QN(n3813) );
  SDFFX1 DFF_1541_Q_reg ( .D(n1960), .SI(test_si90), .SE(n9323), .CLK(n9745), 
        .Q(n8290), .QN(n3812) );
  SDFFX1 DFF_1542_Q_reg ( .D(n1961), .SI(n8290), .SE(n9323), .CLK(n9745), .Q(
        n8289), .QN(n3811) );
  SDFFX1 DFF_1543_Q_reg ( .D(n1962), .SI(n8289), .SE(n9323), .CLK(n9745), .Q(
        n8288), .QN(n3810) );
  SDFFX1 DFF_1544_Q_reg ( .D(n1963), .SI(n8288), .SE(n9323), .CLK(n9745), .Q(
        n8287), .QN(n3809) );
  SDFFX1 DFF_1545_Q_reg ( .D(n1964), .SI(n8287), .SE(n9323), .CLK(n9745), .Q(
        n8286), .QN(n3808) );
  SDFFX1 DFF_1546_Q_reg ( .D(n1965), .SI(n8286), .SE(n9323), .CLK(n9745), .Q(
        n8285), .QN(n3807) );
  SDFFX1 DFF_1547_Q_reg ( .D(n1966), .SI(n8285), .SE(n9323), .CLK(n9745), .Q(
        n8284), .QN(n3806) );
  SDFFX1 DFF_1548_Q_reg ( .D(n1967), .SI(n8284), .SE(n9323), .CLK(n9745), .Q(
        n8283), .QN(n3805) );
  SDFFX1 DFF_1549_Q_reg ( .D(n1968), .SI(n8283), .SE(n9323), .CLK(n9745), .Q(
        n8282), .QN(n3804) );
  SDFFX1 DFF_1550_Q_reg ( .D(n1969), .SI(n8282), .SE(n9323), .CLK(n9745), .Q(
        n8281), .QN(n3803) );
  SDFFX1 DFF_1551_Q_reg ( .D(n1970), .SI(n8281), .SE(n9323), .CLK(n9745), .Q(
        n8280), .QN(n3802) );
  SDFFX1 DFF_1552_Q_reg ( .D(n1971), .SI(n8280), .SE(n9323), .CLK(n9745), .Q(
        n8279), .QN(n3801) );
  SDFFX1 DFF_1553_Q_reg ( .D(n1972), .SI(n8279), .SE(n9324), .CLK(n9744), .Q(
        n8278), .QN(n3800) );
  SDFFX1 DFF_1554_Q_reg ( .D(n1973), .SI(n8278), .SE(n9324), .CLK(n9744), .Q(
        n8277), .QN(n3799) );
  SDFFX1 DFF_1555_Q_reg ( .D(n1974), .SI(n8277), .SE(n9324), .CLK(n9744), .Q(
        n8276), .QN(n3798) );
  SDFFX1 DFF_1556_Q_reg ( .D(n1975), .SI(n8276), .SE(n9324), .CLK(n9744), .Q(
        n8275), .QN(n3797) );
  SDFFX1 DFF_1557_Q_reg ( .D(n1976), .SI(n8275), .SE(n9324), .CLK(n9744), .Q(
        test_so90), .QN(n3796) );
  SDFFX1 DFF_1558_Q_reg ( .D(n1977), .SI(test_si91), .SE(n9324), .CLK(n9744), 
        .Q(n8272), .QN(n3795) );
  SDFFX1 DFF_1559_Q_reg ( .D(n1978), .SI(n8272), .SE(n9324), .CLK(n9744), .Q(
        n8271), .QN(n3794) );
  SDFFX1 DFF_1560_Q_reg ( .D(n1979), .SI(n8271), .SE(n9324), .CLK(n9744), .Q(
        n8270), .QN(n3793) );
  SDFFX1 DFF_1561_Q_reg ( .D(n1980), .SI(n8270), .SE(n9324), .CLK(n9744), .Q(
        n8269), .QN(n3792) );
  SDFFX1 DFF_1562_Q_reg ( .D(n1981), .SI(n8269), .SE(n9324), .CLK(n9744), .Q(
        n8268), .QN(n3791) );
  SDFFX1 DFF_1563_Q_reg ( .D(n1982), .SI(n8268), .SE(n9324), .CLK(n9744), .Q(
        n8267), .QN(n3790) );
  SDFFX1 DFF_1564_Q_reg ( .D(n1983), .SI(n8267), .SE(n9324), .CLK(n9744), .Q(
        n8266), .QN(n3789) );
  SDFFX1 DFF_1565_Q_reg ( .D(n1984), .SI(n8266), .SE(n9325), .CLK(n9743), .Q(
        n8265), .QN(n3788) );
  SDFFX1 DFF_1566_Q_reg ( .D(n1985), .SI(n8265), .SE(n9325), .CLK(n9743), .Q(
        n8264), .QN(n3787) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n9325), .CLK(n9743), 
        .Q(n8263), .QN(n3786) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(n9309), .CLK(n9759), 
        .Q(n8262), .QN(n15997) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(n9322), .CLK(n9746), 
        .Q(n8261), .QN(n15996) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(n9322), .CLK(n9746), 
        .Q(n8260), .QN(n15995) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(n9322), .CLK(n9746), 
        .Q(n8259), .QN(n15994) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(n9322), .CLK(n9746), 
        .Q(n8258), .QN(n15993) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(n9321), .CLK(n9747), 
        .Q(n8257), .QN(n15992) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(n9309), .CLK(n9759), 
        .Q(test_so91), .QN(n9097) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(n9321), .CLK(n9747), 
        .Q(n8254), .QN(n15991) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(n9321), .CLK(n9747), 
        .Q(n8253), .QN(n15990) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(n9321), .CLK(n9747), 
        .Q(n8252), .QN(n15989) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(n9320), .CLK(n9748), 
        .Q(n8251), .QN(n15988) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(n9320), .CLK(n9748), 
        .Q(n8250), .QN(n15987) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(n9320), .CLK(n9748), 
        .Q(n8249), .QN(n15986) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(n9320), .CLK(n9748), 
        .Q(n8248), .QN(n15985) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(n9319), .CLK(n9749), 
        .Q(n8247), .QN(n15984) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(n9319), .CLK(n9749), 
        .Q(n8246), .QN(n15983) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(n9319), .CLK(n9749), 
        .Q(WX11021), .QN(n8146) );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(n9318), .CLK(n9750), 
        .Q(WX11023), .QN(n8144) );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(n9318), .CLK(n9750), 
        .Q(WX11025), .QN(n8142) );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(n9318), .CLK(n9750), 
        .Q(WX11027), .QN(n8140) );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(n9317), .CLK(n9751), 
        .Q(WX11029), .QN(n8138) );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(n9317), .CLK(n9751), 
        .Q(WX11031), .QN(n8136) );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(n9317), .CLK(n9751), 
        .Q(WX11033), .QN(n8134) );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(n9316), .CLK(n9752), 
        .Q(test_so92), .QN(n9144) );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(n9316), .CLK(n9752), 
        .Q(WX11037), .QN(n8131) );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(n9316), .CLK(n9752), 
        .Q(WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(n9315), .CLK(n9753), 
        .Q(WX11041), .QN(n8127) );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(n9315), .CLK(n9753), 
        .Q(WX11043), .QN(n8126) );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(n9315), .CLK(n9753), 
        .Q(WX11045), .QN(n8124) );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(n9314), .CLK(n9754), 
        .Q(WX11047), .QN(n8122) );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(n9314), .CLK(n9754), 
        .Q(WX11049), .QN(n8120) );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(n9314), .CLK(n9754), 
        .Q(WX11051), .QN(n8118) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n9313), .CLK(n9755), 
        .Q(WX11053), .QN(n7876) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n9322), .CLK(n9746), 
        .Q(WX11055), .QN(n7918) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n9322), .CLK(n9746), 
        .Q(WX11057), .QN(n7916) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n9322), .CLK(n9746), 
        .Q(WX11059), .QN(n7914) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n9322), .CLK(n9746), 
        .Q(WX11061), .QN(n7912) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n9321), .CLK(n9747), 
        .Q(WX11063), .QN(n7910) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n9321), .CLK(n9747), 
        .Q(WX11065), .QN(n7908) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n9321), .CLK(n9747), 
        .Q(WX11067), .QN(n7906) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n9321), .CLK(n9747), 
        .Q(test_so93), .QN(n9146) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n9321), .CLK(n9747), 
        .Q(WX11071), .QN(n7903) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n9321), .CLK(n9747), 
        .Q(WX11073), .QN(n7902) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n9320), .CLK(n9748), 
        .Q(WX11075), .QN(n7900) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n9320), .CLK(n9748), 
        .Q(WX11077), .QN(n7898) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n9320), .CLK(n9748), 
        .Q(WX11079), .QN(n7896) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n9319), .CLK(n9749), 
        .Q(WX11081), .QN(n7894) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n9319), .CLK(n9749), 
        .Q(WX11083), .QN(n7892) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n9319), .CLK(n9749), 
        .Q(WX11085) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n9318), .CLK(n9750), 
        .Q(WX11087) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n9318), .CLK(n9750), 
        .Q(WX11089) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n9318), .CLK(n9750), 
        .Q(WX11091) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n9317), .CLK(n9751), 
        .Q(WX11093) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n9317), .CLK(n9751), 
        .Q(WX11095) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n9317), .CLK(n9751), 
        .Q(WX11097) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n9316), .CLK(n9752), 
        .Q(WX11099) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n9316), .CLK(n9752), 
        .Q(WX11101) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n9316), .CLK(n9752), 
        .Q(test_so94), .QN(n9143) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n9315), .CLK(n9753), 
        .Q(WX11105) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n9315), .CLK(n9753), 
        .Q(WX11107) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n9315), .CLK(n9753), 
        .Q(WX11109) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n9314), .CLK(n9754), 
        .Q(WX11111) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n9314), .CLK(n9754), 
        .Q(WX11113) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n9314), .CLK(n9754), 
        .Q(WX11115) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n9313), .CLK(n9755), 
        .Q(WX11117), .QN(n7877) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n9313), .CLK(n9755), 
        .Q(WX11119), .QN(n7919) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n9313), .CLK(n9755), 
        .Q(WX11121), .QN(n7917) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n9313), .CLK(n9755), 
        .Q(WX11123), .QN(n7915) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n9313), .CLK(n9755), 
        .Q(WX11125), .QN(n7913) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n9313), .CLK(n9755), 
        .Q(WX11127), .QN(n7911) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n9312), .CLK(n9756), 
        .Q(WX11129), .QN(n7909) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n9312), .CLK(n9756), 
        .Q(WX11131), .QN(n7907) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n9321), .CLK(n9747), 
        .Q(WX11133), .QN(n7905) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n9321), .CLK(n9747), 
        .Q(WX11135), .QN(n7904) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n9320), .CLK(n9748), 
        .Q(test_so95), .QN(n9145) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n9320), .CLK(n9748), 
        .Q(WX11139), .QN(n7901) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n9320), .CLK(n9748), 
        .Q(WX11141), .QN(n7899) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n9320), .CLK(n9748), 
        .Q(WX11143), .QN(n7897) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n9319), .CLK(n9749), 
        .Q(WX11145), .QN(n7895) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n9319), .CLK(n9749), 
        .Q(WX11147), .QN(n7893) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n9319), .CLK(n9749), 
        .Q(WX11149), .QN(n8147) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n9318), .CLK(n9750), 
        .Q(WX11151), .QN(n8145) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n9318), .CLK(n9750), 
        .Q(WX11153), .QN(n8143) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n9318), .CLK(n9750), 
        .Q(WX11155), .QN(n8141) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155), .SE(n9317), .CLK(n9751), 
        .Q(WX11157), .QN(n8139) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(n9317), .CLK(n9751), 
        .Q(WX11159), .QN(n8137) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(n9317), .CLK(n9751), 
        .Q(WX11161), .QN(n8135) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(n9316), .CLK(n9752), 
        .Q(WX11163), .QN(n8133) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(n9316), .CLK(n9752), 
        .Q(WX11165), .QN(n8132) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(n9316), .CLK(n9752), 
        .Q(WX11167), .QN(n8130) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(n9315), .CLK(n9753), 
        .Q(WX11169), .QN(n8128) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(n9315), .CLK(n9753), 
        .Q(test_so96), .QN(n9142) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n9315), .CLK(n9753), 
        .Q(WX11173), .QN(n8125) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n9314), .CLK(n9754), 
        .Q(WX11175), .QN(n8123) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n9314), .CLK(n9754), 
        .Q(WX11177), .QN(n8121) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n9314), .CLK(n9754), 
        .Q(WX11179), .QN(n8119) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n9313), .CLK(n9755), 
        .Q(WX11181), .QN(n8742) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n9313), .CLK(n9755), 
        .Q(WX11183), .QN(n8743) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n9313), .CLK(n9755), 
        .Q(WX11185), .QN(n8744) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n9313), .CLK(n9755), 
        .Q(WX11187), .QN(n8745) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n9313), .CLK(n9755), 
        .Q(WX11189), .QN(n8746) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n9312), .CLK(n9756), 
        .Q(WX11191), .QN(n8747) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n9312), .CLK(n9756), 
        .Q(WX11193), .QN(n8748) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n9312), .CLK(n9756), 
        .Q(WX11195), .QN(n8749) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n9312), .CLK(n9756), 
        .Q(WX11197), .QN(n8750) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n9312), .CLK(n9756), 
        .Q(WX11199), .QN(n8751) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n9312), .CLK(n9756), 
        .Q(WX11201), .QN(n8752) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n9312), .CLK(n9756), 
        .Q(WX11203), .QN(n8753) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n9312), .CLK(n9756), 
        .Q(test_so97), .QN(n9109) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n9320), .CLK(n9748), 
        .Q(WX11207), .QN(n8754) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n9319), .CLK(n9749), 
        .Q(WX11209), .QN(n8755) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n9319), .CLK(n9749), 
        .Q(WX11211), .QN(n8713) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n9319), .CLK(n9749), 
        .Q(WX11213), .QN(n8756) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n9318), .CLK(n9750), 
        .Q(WX11215), .QN(n8757) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n9318), .CLK(n9750), 
        .Q(WX11217), .QN(n8758) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n9318), .CLK(n9750), 
        .Q(WX11219), .QN(n8759) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n9317), .CLK(n9751), 
        .Q(WX11221), .QN(n8714) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n9317), .CLK(n9751), 
        .Q(WX11223), .QN(n8760) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n9317), .CLK(n9751), 
        .Q(WX11225), .QN(n8761) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n9316), .CLK(n9752), 
        .Q(WX11227), .QN(n8762) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n9316), .CLK(n9752), 
        .Q(WX11229), .QN(n8763) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n9316), .CLK(n9752), 
        .Q(WX11231), .QN(n8764) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n9315), .CLK(n9753), 
        .Q(WX11233), .QN(n8765) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n9315), .CLK(n9753), 
        .Q(WX11235), .QN(n8715) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n9315), .CLK(n9753), 
        .Q(WX11237), .QN(n8766) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n9314), .CLK(n9754), 
        .Q(test_so98), .QN(n9102) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n9314), .CLK(n9754), 
        .Q(WX11241), .QN(n8767) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n9314), .CLK(n9754), 
        .Q(WX11243), .QN(n8734) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n9311), .CLK(n9757), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_1), .QN(DFF_1697_n1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_3), .QN(DFF_1699_n1) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_10), .QN(DFF_1706_n1) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n9310), .CLK(
        n9758), .Q(test_so99), .QN(n9163) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n9310), .CLK(n9758), .Q(CRC_OUT_1_15), .QN(DFF_1711_n1) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n9310), .CLK(
        n9758), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n9309), .CLK(
        n9759), .Q(CRC_OUT_1_18), .QN(DFF_1714_n1) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n9309), .CLK(
        n9759), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n9309), .CLK(
        n9759), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n9309), .CLK(
        n9759), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n9309), .CLK(
        n9759), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n9309), .CLK(
        n9759), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n9312), .CLK(
        n9756), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n9312), .CLK(
        n9756), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n9311), .CLK(
        n9757), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n9311), .CLK(
        n9757), .Q(test_so100), .QN(n9085) );
  NOR2X0 Trojan1 ( .IN1(WX3442), .IN2(WX5974), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(WX806), .IN2(WX782), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(WX11632), .IN2(n524), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(WX5964), .IN2(WX3324), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(WX8634), .IN2(WX3330), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n536), .IN2(n528), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(WX862), .IN2(WX7227), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(WX11616), .IN2(n1972), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(n9433), .Q(
        Tj_Trigger) );
  NAND3X4 TrojanPayload1 ( .IN1(WX547), .IN2(Tj_Trigger), .IN3(Stage4), .QN(
        Stage1_1) );
  INVX8 TrojanPayload2 ( .INP(Stage1_1), .ZN(Stage1_2) );
  INVX8 TrojanPayload3 ( .INP(Stage1_2), .ZN(Stage1_3) );
  INVX8 TrojanPayload4 ( .INP(Stage1_3), .ZN(Stage1_4) );
  INVX8 TrojanPayload5 ( .INP(Stage1_4), .ZN(Stage1) );
  MUX21X2 TrojanPayload6 ( .IN1(WX544), .IN2(Stage1), .S(1'b0), .Q(Stage2_i)
         );
  INVX8 TrojanPayload7 ( .INP(Stage2_i), .ZN(Stage2_7) );
  INVX8 TrojanPayload8 ( .INP(Stage2_7), .ZN(Stage2_8) );
  INVX8 TrojanPayload9 ( .INP(Stage2_8), .ZN(Stage2_9) );
  INVX8 TrojanPayload10 ( .INP(Stage2_9), .ZN(Stage2_10) );
  INVX8 TrojanPayload11 ( .INP(Stage2_10), .ZN(Stage2) );
  MUX21X2 TrojanPayload12 ( .IN1(WX706), .IN2(Stage2), .S(1'b0), .Q(Stage3_i)
         );
  INVX8 TrojanPayload13 ( .INP(Stage3_i), .ZN(Stage3_12) );
  INVX8 TrojanPayload14 ( .INP(Stage3_12), .ZN(Stage3_13) );
  INVX8 TrojanPayload15 ( .INP(Stage3_13), .ZN(Stage3_14) );
  INVX8 TrojanPayload16 ( .INP(Stage3_14), .ZN(Stage3_15) );
  INVX8 TrojanPayload17 ( .INP(Stage3_15) );
  MUX21X2 TrojanPayload18 ( .IN1(n3467), .IN2(1'b0), .S(1'b0), .Q(Stage4_i) );
  INVX8 TrojanPayload19 ( .INP(Stage4_i), .ZN(Stage4_17) );
  INVX8 TrojanPayload20 ( .INP(Stage4_17), .ZN(Stage4_18) );
  INVX8 TrojanPayload21 ( .INP(Stage4_18), .ZN(Stage4_19) );
  INVX8 TrojanPayload22 ( .INP(Stage4_19), .ZN(Stage4_20) );
  INVX8 TrojanPayload23 ( .INP(Stage4_20), .ZN(Stage4_21) );
  INVX8 TrojanPayload24 ( .INP(Stage4_21), .ZN(Stage4) );
  INVX2 U8990 ( .INP(TM0), .ZN(n2199) );
  NBUFFX2 U8991 ( .INP(n9254), .Z(n9228) );
  NBUFFX2 U8992 ( .INP(n9254), .Z(n9229) );
  NBUFFX2 U8993 ( .INP(n9252), .Z(n9237) );
  NBUFFX2 U8994 ( .INP(n9252), .Z(n9239) );
  NBUFFX2 U8995 ( .INP(n9251), .Z(n9240) );
  NBUFFX2 U8996 ( .INP(n9251), .Z(n9241) );
  NBUFFX2 U8997 ( .INP(n9251), .Z(n9242) );
  NBUFFX2 U8998 ( .INP(n9251), .Z(n9243) );
  NBUFFX2 U8999 ( .INP(n9251), .Z(n9244) );
  NBUFFX2 U9000 ( .INP(n9250), .Z(n9248) );
  NBUFFX2 U9001 ( .INP(n9253), .Z(n9230) );
  NBUFFX2 U9002 ( .INP(n9253), .Z(n9231) );
  NBUFFX2 U9003 ( .INP(n9253), .Z(n9232) );
  NBUFFX2 U9004 ( .INP(n9252), .Z(n9238) );
  NBUFFX2 U9005 ( .INP(n9253), .Z(n9233) );
  NBUFFX2 U9006 ( .INP(n9253), .Z(n9234) );
  NBUFFX2 U9007 ( .INP(n9252), .Z(n9235) );
  NBUFFX2 U9008 ( .INP(n9252), .Z(n9236) );
  NBUFFX2 U9009 ( .INP(n9250), .Z(n9245) );
  NBUFFX2 U9010 ( .INP(n9250), .Z(n9246) );
  NBUFFX2 U9011 ( .INP(n9250), .Z(n9247) );
  NBUFFX2 U9012 ( .INP(n9254), .Z(n9227) );
  NBUFFX2 U9013 ( .INP(n9805), .Z(n9636) );
  NBUFFX2 U9014 ( .INP(n9805), .Z(n9634) );
  NBUFFX2 U9015 ( .INP(n9805), .Z(n9635) );
  NBUFFX2 U9016 ( .INP(n9805), .Z(n9633) );
  NBUFFX2 U9017 ( .INP(n9780), .Z(n9758) );
  NBUFFX2 U9018 ( .INP(n9780), .Z(n9757) );
  NBUFFX2 U9019 ( .INP(n9781), .Z(n9756) );
  NBUFFX2 U9020 ( .INP(n9781), .Z(n9755) );
  NBUFFX2 U9021 ( .INP(n9781), .Z(n9754) );
  NBUFFX2 U9022 ( .INP(n9781), .Z(n9753) );
  NBUFFX2 U9023 ( .INP(n9781), .Z(n9752) );
  NBUFFX2 U9024 ( .INP(n9782), .Z(n9751) );
  NBUFFX2 U9025 ( .INP(n9782), .Z(n9750) );
  NBUFFX2 U9026 ( .INP(n9782), .Z(n9749) );
  NBUFFX2 U9027 ( .INP(n9782), .Z(n9748) );
  NBUFFX2 U9028 ( .INP(n9782), .Z(n9747) );
  NBUFFX2 U9029 ( .INP(n9783), .Z(n9744) );
  NBUFFX2 U9030 ( .INP(n9783), .Z(n9745) );
  NBUFFX2 U9031 ( .INP(n9783), .Z(n9746) );
  NBUFFX2 U9032 ( .INP(n9783), .Z(n9743) );
  NBUFFX2 U9033 ( .INP(n9780), .Z(n9760) );
  NBUFFX2 U9034 ( .INP(n9780), .Z(n9759) );
  NBUFFX2 U9035 ( .INP(n9783), .Z(n9742) );
  NBUFFX2 U9036 ( .INP(n9784), .Z(n9741) );
  NBUFFX2 U9037 ( .INP(n9784), .Z(n9740) );
  NBUFFX2 U9038 ( .INP(n9784), .Z(n9739) );
  NBUFFX2 U9039 ( .INP(n9784), .Z(n9738) );
  NBUFFX2 U9040 ( .INP(n9784), .Z(n9737) );
  NBUFFX2 U9041 ( .INP(n9785), .Z(n9736) );
  NBUFFX2 U9042 ( .INP(n9785), .Z(n9735) );
  NBUFFX2 U9043 ( .INP(n9785), .Z(n9734) );
  NBUFFX2 U9044 ( .INP(n9785), .Z(n9733) );
  NBUFFX2 U9045 ( .INP(n9785), .Z(n9732) );
  NBUFFX2 U9046 ( .INP(n9786), .Z(n9730) );
  NBUFFX2 U9047 ( .INP(n9786), .Z(n9731) );
  NBUFFX2 U9048 ( .INP(n9779), .Z(n9762) );
  NBUFFX2 U9049 ( .INP(n9780), .Z(n9761) );
  NBUFFX2 U9050 ( .INP(n9786), .Z(n9729) );
  NBUFFX2 U9051 ( .INP(n9786), .Z(n9728) );
  NBUFFX2 U9052 ( .INP(n9786), .Z(n9727) );
  NBUFFX2 U9053 ( .INP(n9787), .Z(n9726) );
  NBUFFX2 U9054 ( .INP(n9787), .Z(n9725) );
  NBUFFX2 U9055 ( .INP(n9787), .Z(n9724) );
  NBUFFX2 U9056 ( .INP(n9787), .Z(n9723) );
  NBUFFX2 U9057 ( .INP(n9787), .Z(n9722) );
  NBUFFX2 U9058 ( .INP(n9788), .Z(n9721) );
  NBUFFX2 U9059 ( .INP(n9788), .Z(n9720) );
  NBUFFX2 U9060 ( .INP(n9788), .Z(n9719) );
  NBUFFX2 U9061 ( .INP(n9779), .Z(n9763) );
  NBUFFX2 U9062 ( .INP(n9788), .Z(n9717) );
  NBUFFX2 U9063 ( .INP(n9788), .Z(n9718) );
  NBUFFX2 U9064 ( .INP(n9789), .Z(n9716) );
  NBUFFX2 U9065 ( .INP(n9779), .Z(n9765) );
  NBUFFX2 U9066 ( .INP(n9779), .Z(n9764) );
  NBUFFX2 U9067 ( .INP(n9789), .Z(n9715) );
  NBUFFX2 U9068 ( .INP(n9789), .Z(n9714) );
  NBUFFX2 U9069 ( .INP(n9789), .Z(n9713) );
  NBUFFX2 U9070 ( .INP(n9789), .Z(n9712) );
  NBUFFX2 U9071 ( .INP(n9790), .Z(n9711) );
  NBUFFX2 U9072 ( .INP(n9790), .Z(n9710) );
  NBUFFX2 U9073 ( .INP(n9790), .Z(n9709) );
  NBUFFX2 U9074 ( .INP(n9790), .Z(n9708) );
  NBUFFX2 U9075 ( .INP(n9790), .Z(n9707) );
  NBUFFX2 U9076 ( .INP(n9791), .Z(n9706) );
  NBUFFX2 U9077 ( .INP(n9791), .Z(n9705) );
  NBUFFX2 U9078 ( .INP(n9791), .Z(n9703) );
  NBUFFX2 U9079 ( .INP(n9791), .Z(n9704) );
  NBUFFX2 U9080 ( .INP(n9791), .Z(n9702) );
  NBUFFX2 U9081 ( .INP(n9778), .Z(n9767) );
  NBUFFX2 U9082 ( .INP(n9779), .Z(n9766) );
  NBUFFX2 U9083 ( .INP(n9792), .Z(n9701) );
  NBUFFX2 U9084 ( .INP(n9792), .Z(n9700) );
  NBUFFX2 U9085 ( .INP(n9792), .Z(n9699) );
  NBUFFX2 U9086 ( .INP(n9792), .Z(n9698) );
  NBUFFX2 U9087 ( .INP(n9792), .Z(n9697) );
  NBUFFX2 U9088 ( .INP(n9793), .Z(n9696) );
  NBUFFX2 U9089 ( .INP(n9793), .Z(n9695) );
  NBUFFX2 U9090 ( .INP(n9793), .Z(n9694) );
  NBUFFX2 U9091 ( .INP(n9793), .Z(n9693) );
  NBUFFX2 U9092 ( .INP(n9793), .Z(n9692) );
  NBUFFX2 U9093 ( .INP(n9794), .Z(n9691) );
  NBUFFX2 U9094 ( .INP(n9794), .Z(n9689) );
  NBUFFX2 U9095 ( .INP(n9794), .Z(n9690) );
  NBUFFX2 U9096 ( .INP(n9794), .Z(n9688) );
  NBUFFX2 U9097 ( .INP(n9778), .Z(n9769) );
  NBUFFX2 U9098 ( .INP(n9778), .Z(n9768) );
  NBUFFX2 U9099 ( .INP(n9794), .Z(n9687) );
  NBUFFX2 U9100 ( .INP(n9795), .Z(n9686) );
  NBUFFX2 U9101 ( .INP(n9795), .Z(n9685) );
  NBUFFX2 U9102 ( .INP(n9795), .Z(n9684) );
  NBUFFX2 U9103 ( .INP(n9795), .Z(n9683) );
  NBUFFX2 U9104 ( .INP(n9795), .Z(n9682) );
  NBUFFX2 U9105 ( .INP(n9796), .Z(n9681) );
  NBUFFX2 U9106 ( .INP(n9796), .Z(n9680) );
  NBUFFX2 U9107 ( .INP(n9796), .Z(n9679) );
  NBUFFX2 U9108 ( .INP(n9796), .Z(n9678) );
  NBUFFX2 U9109 ( .INP(n9797), .Z(n9675) );
  NBUFFX2 U9110 ( .INP(n9797), .Z(n9676) );
  NBUFFX2 U9111 ( .INP(n9796), .Z(n9677) );
  NBUFFX2 U9112 ( .INP(n9777), .Z(n9772) );
  NBUFFX2 U9113 ( .INP(n9778), .Z(n9771) );
  NBUFFX2 U9114 ( .INP(n9778), .Z(n9770) );
  NBUFFX2 U9115 ( .INP(n9797), .Z(n9674) );
  NBUFFX2 U9116 ( .INP(n9797), .Z(n9673) );
  NBUFFX2 U9117 ( .INP(n9797), .Z(n9672) );
  NBUFFX2 U9118 ( .INP(n9798), .Z(n9671) );
  NBUFFX2 U9119 ( .INP(n9798), .Z(n9670) );
  NBUFFX2 U9120 ( .INP(n9798), .Z(n9669) );
  NBUFFX2 U9121 ( .INP(n9798), .Z(n9668) );
  NBUFFX2 U9122 ( .INP(n9798), .Z(n9667) );
  NBUFFX2 U9123 ( .INP(n9799), .Z(n9666) );
  NBUFFX2 U9124 ( .INP(n9799), .Z(n9665) );
  NBUFFX2 U9125 ( .INP(n9799), .Z(n9662) );
  NBUFFX2 U9126 ( .INP(n9799), .Z(n9663) );
  NBUFFX2 U9127 ( .INP(n9799), .Z(n9664) );
  NBUFFX2 U9128 ( .INP(n9800), .Z(n9661) );
  NBUFFX2 U9129 ( .INP(n9777), .Z(n9774) );
  NBUFFX2 U9130 ( .INP(n9777), .Z(n9773) );
  NBUFFX2 U9131 ( .INP(n9800), .Z(n9660) );
  NBUFFX2 U9132 ( .INP(n9800), .Z(n9659) );
  NBUFFX2 U9133 ( .INP(n9800), .Z(n9658) );
  NBUFFX2 U9134 ( .INP(n9800), .Z(n9657) );
  NBUFFX2 U9135 ( .INP(n9801), .Z(n9656) );
  NBUFFX2 U9136 ( .INP(n9801), .Z(n9655) );
  NBUFFX2 U9137 ( .INP(n9801), .Z(n9654) );
  NBUFFX2 U9138 ( .INP(n9801), .Z(n9653) );
  NBUFFX2 U9139 ( .INP(n9801), .Z(n9652) );
  NBUFFX2 U9140 ( .INP(n9802), .Z(n9651) );
  NBUFFX2 U9141 ( .INP(n9802), .Z(n9650) );
  NBUFFX2 U9142 ( .INP(n9802), .Z(n9648) );
  NBUFFX2 U9143 ( .INP(n9802), .Z(n9649) );
  NBUFFX2 U9144 ( .INP(n9802), .Z(n9647) );
  NBUFFX2 U9145 ( .INP(n9777), .Z(n9776) );
  NBUFFX2 U9146 ( .INP(n9777), .Z(n9775) );
  NBUFFX2 U9147 ( .INP(n9803), .Z(n9646) );
  NBUFFX2 U9148 ( .INP(n9803), .Z(n9645) );
  NBUFFX2 U9149 ( .INP(n9803), .Z(n9644) );
  NBUFFX2 U9150 ( .INP(n9803), .Z(n9643) );
  NBUFFX2 U9151 ( .INP(n9803), .Z(n9642) );
  NBUFFX2 U9152 ( .INP(n9804), .Z(n9641) );
  NBUFFX2 U9153 ( .INP(n9804), .Z(n9640) );
  NBUFFX2 U9154 ( .INP(n9804), .Z(n9639) );
  NBUFFX2 U9155 ( .INP(n9804), .Z(n9638) );
  NBUFFX2 U9156 ( .INP(n9804), .Z(n9637) );
  NBUFFX2 U9157 ( .INP(n9250), .Z(n9249) );
  NBUFFX2 U9158 ( .INP(n9283), .Z(n9264) );
  NBUFFX2 U9159 ( .INP(n9169), .Z(n9178) );
  NBUFFX2 U9160 ( .INP(n9172), .Z(n9194) );
  NBUFFX2 U9161 ( .INP(n9172), .Z(n9193) );
  NBUFFX2 U9162 ( .INP(n9281), .Z(n9271) );
  NBUFFX2 U9163 ( .INP(n9281), .Z(n9272) );
  NBUFFX2 U9164 ( .INP(n9281), .Z(n9273) );
  NBUFFX2 U9165 ( .INP(n9281), .Z(n9274) );
  NBUFFX2 U9166 ( .INP(n9280), .Z(n9278) );
  NBUFFX2 U9167 ( .INP(n9282), .Z(n9266) );
  NBUFFX2 U9168 ( .INP(n9282), .Z(n9267) );
  NBUFFX2 U9169 ( .INP(n9282), .Z(n9268) );
  NBUFFX2 U9170 ( .INP(n9282), .Z(n9265) );
  NBUFFX2 U9171 ( .INP(n9281), .Z(n9270) );
  NBUFFX2 U9172 ( .INP(n9282), .Z(n9269) );
  NBUFFX2 U9173 ( .INP(n9280), .Z(n9275) );
  NBUFFX2 U9174 ( .INP(n9280), .Z(n9276) );
  NBUFFX2 U9175 ( .INP(n9280), .Z(n9277) );
  NBUFFX2 U9176 ( .INP(n9170), .Z(n9186) );
  NBUFFX2 U9177 ( .INP(n9170), .Z(n9185) );
  NBUFFX2 U9178 ( .INP(n9170), .Z(n9184) );
  NBUFFX2 U9179 ( .INP(n9170), .Z(n9183) );
  NBUFFX2 U9180 ( .INP(n9169), .Z(n9182) );
  NBUFFX2 U9181 ( .INP(n9171), .Z(n9192) );
  NBUFFX2 U9182 ( .INP(n9171), .Z(n9191) );
  NBUFFX2 U9183 ( .INP(n9171), .Z(n9190) );
  NBUFFX2 U9184 ( .INP(n9171), .Z(n9189) );
  NBUFFX2 U9185 ( .INP(n9171), .Z(n9188) );
  NBUFFX2 U9186 ( .INP(n9170), .Z(n9187) );
  NBUFFX2 U9187 ( .INP(n9169), .Z(n9179) );
  NBUFFX2 U9188 ( .INP(n9169), .Z(n9180) );
  NBUFFX2 U9189 ( .INP(n9169), .Z(n9181) );
  NBUFFX2 U9190 ( .INP(n9284), .Z(n9257) );
  NBUFFX2 U9191 ( .INP(n9284), .Z(n9259) );
  NBUFFX2 U9192 ( .INP(n9284), .Z(n9258) );
  NBUFFX2 U9193 ( .INP(n9283), .Z(n9263) );
  NBUFFX2 U9194 ( .INP(n9283), .Z(n9262) );
  NBUFFX2 U9195 ( .INP(n9283), .Z(n9260) );
  NBUFFX2 U9196 ( .INP(n9283), .Z(n9261) );
  NBUFFX2 U9197 ( .INP(n9168), .Z(n9177) );
  NBUFFX2 U9198 ( .INP(n9168), .Z(n9176) );
  NBUFFX2 U9199 ( .INP(n9168), .Z(n9175) );
  NBUFFX2 U9200 ( .INP(n9168), .Z(n9174) );
  NBUFFX2 U9201 ( .INP(n9168), .Z(n9173) );
  NBUFFX2 U9202 ( .INP(n9280), .Z(n9279) );
  NBUFFX2 U9203 ( .INP(n9172), .Z(n9195) );
  NBUFFX2 U9204 ( .INP(n9200), .Z(n9223) );
  NBUFFX2 U9205 ( .INP(n9200), .Z(n9221) );
  NBUFFX2 U9206 ( .INP(n9200), .Z(n9222) );
  NBUFFX2 U9207 ( .INP(n9198), .Z(n9211) );
  NBUFFX2 U9208 ( .INP(n9198), .Z(n9212) );
  NBUFFX2 U9209 ( .INP(n9198), .Z(n9213) );
  NBUFFX2 U9210 ( .INP(n9198), .Z(n9214) );
  NBUFFX2 U9211 ( .INP(n9198), .Z(n9215) );
  NBUFFX2 U9212 ( .INP(n9199), .Z(n9216) );
  NBUFFX2 U9213 ( .INP(n9199), .Z(n9217) );
  NBUFFX2 U9214 ( .INP(n9199), .Z(n9218) );
  NBUFFX2 U9215 ( .INP(n9199), .Z(n9219) );
  NBUFFX2 U9216 ( .INP(n9196), .Z(n9201) );
  NBUFFX2 U9217 ( .INP(n9196), .Z(n9202) );
  NBUFFX2 U9218 ( .INP(n9196), .Z(n9203) );
  NBUFFX2 U9219 ( .INP(n9196), .Z(n9204) );
  NBUFFX2 U9220 ( .INP(n9196), .Z(n9205) );
  NBUFFX2 U9221 ( .INP(n9197), .Z(n9206) );
  NBUFFX2 U9222 ( .INP(n9197), .Z(n9207) );
  NBUFFX2 U9223 ( .INP(n9197), .Z(n9208) );
  NBUFFX2 U9224 ( .INP(n9197), .Z(n9209) );
  NBUFFX2 U9225 ( .INP(n9197), .Z(n9210) );
  NBUFFX2 U9226 ( .INP(n9199), .Z(n9220) );
  NBUFFX2 U9227 ( .INP(n9200), .Z(n9224) );
  INVX0 U9228 ( .INP(n9289), .ZN(n9434) );
  INVX0 U9229 ( .INP(n9288), .ZN(n9433) );
  INVX0 U9230 ( .INP(n9288), .ZN(n9432) );
  INVX0 U9231 ( .INP(n9287), .ZN(n9431) );
  INVX0 U9232 ( .INP(n9287), .ZN(n9430) );
  INVX0 U9233 ( .INP(n9286), .ZN(n9429) );
  INVX0 U9234 ( .INP(n9286), .ZN(n9428) );
  INVX0 U9235 ( .INP(n9289), .ZN(n9435) );
  INVX0 U9236 ( .INP(n9285), .ZN(n9427) );
  INVX0 U9237 ( .INP(n9285), .ZN(n9426) );
  NBUFFX2 U9238 ( .INP(n9290), .Z(n9288) );
  NBUFFX2 U9239 ( .INP(n9290), .Z(n9287) );
  NBUFFX2 U9240 ( .INP(n9291), .Z(n9286) );
  NBUFFX2 U9241 ( .INP(n9290), .Z(n9289) );
  NBUFFX2 U9242 ( .INP(n9291), .Z(n9285) );
  NBUFFX2 U9243 ( .INP(n9821), .Z(n9168) );
  NBUFFX2 U9244 ( .INP(n9821), .Z(n9169) );
  NBUFFX2 U9245 ( .INP(n9821), .Z(n9170) );
  NBUFFX2 U9246 ( .INP(n9821), .Z(n9171) );
  NBUFFX2 U9247 ( .INP(n9821), .Z(n9172) );
  NBUFFX2 U9248 ( .INP(n2148), .Z(n9196) );
  NBUFFX2 U9249 ( .INP(n2148), .Z(n9197) );
  NBUFFX2 U9250 ( .INP(n2148), .Z(n9198) );
  NBUFFX2 U9251 ( .INP(n2148), .Z(n9199) );
  NBUFFX2 U9252 ( .INP(n2148), .Z(n9200) );
  NBUFFX2 U9253 ( .INP(n2152), .Z(n9225) );
  NBUFFX2 U9254 ( .INP(n2152), .Z(n9226) );
  NBUFFX2 U9255 ( .INP(n9225), .Z(n9250) );
  NBUFFX2 U9256 ( .INP(n9225), .Z(n9251) );
  NBUFFX2 U9257 ( .INP(n9225), .Z(n9252) );
  NBUFFX2 U9258 ( .INP(n9226), .Z(n9253) );
  NBUFFX2 U9259 ( .INP(n9226), .Z(n9254) );
  NBUFFX2 U9260 ( .INP(n2153), .Z(n9255) );
  NBUFFX2 U9261 ( .INP(n2153), .Z(n9256) );
  NBUFFX2 U9262 ( .INP(n9255), .Z(n9280) );
  NBUFFX2 U9263 ( .INP(n9255), .Z(n9281) );
  NBUFFX2 U9264 ( .INP(n9255), .Z(n9282) );
  NBUFFX2 U9265 ( .INP(n9256), .Z(n9283) );
  NBUFFX2 U9266 ( .INP(n9256), .Z(n9284) );
  NBUFFX2 U9267 ( .INP(test_se), .Z(n9290) );
  NBUFFX2 U9268 ( .INP(test_se), .Z(n9291) );
  INVX0 U9269 ( .INP(n9434), .ZN(n9292) );
  INVX0 U9270 ( .INP(n9434), .ZN(n9293) );
  INVX0 U9271 ( .INP(n9429), .ZN(n9294) );
  INVX0 U9272 ( .INP(n9431), .ZN(n9295) );
  INVX0 U9273 ( .INP(n9432), .ZN(n9296) );
  INVX0 U9274 ( .INP(n9433), .ZN(n9297) );
  INVX0 U9275 ( .INP(n9432), .ZN(n9298) );
  INVX0 U9276 ( .INP(n9431), .ZN(n9299) );
  INVX0 U9277 ( .INP(n9430), .ZN(n9300) );
  INVX0 U9278 ( .INP(n9434), .ZN(n9301) );
  INVX0 U9279 ( .INP(n9435), .ZN(n9302) );
  INVX0 U9280 ( .INP(n9431), .ZN(n9303) );
  INVX0 U9281 ( .INP(n9435), .ZN(n9304) );
  INVX0 U9282 ( .INP(n9435), .ZN(n9305) );
  INVX0 U9283 ( .INP(n9435), .ZN(n9306) );
  INVX0 U9284 ( .INP(n9435), .ZN(n9307) );
  INVX0 U9285 ( .INP(n9435), .ZN(n9308) );
  INVX0 U9286 ( .INP(n9435), .ZN(n9309) );
  INVX0 U9287 ( .INP(n9434), .ZN(n9310) );
  INVX0 U9288 ( .INP(n9434), .ZN(n9311) );
  INVX0 U9289 ( .INP(n9434), .ZN(n9312) );
  INVX0 U9290 ( .INP(n9434), .ZN(n9313) );
  INVX0 U9291 ( .INP(n9434), .ZN(n9314) );
  INVX0 U9292 ( .INP(n9434), .ZN(n9315) );
  INVX0 U9293 ( .INP(n9433), .ZN(n9316) );
  INVX0 U9294 ( .INP(n9433), .ZN(n9317) );
  INVX0 U9295 ( .INP(n9433), .ZN(n9318) );
  INVX0 U9296 ( .INP(n9433), .ZN(n9319) );
  INVX0 U9297 ( .INP(n9433), .ZN(n9320) );
  INVX0 U9298 ( .INP(n9433), .ZN(n9321) );
  INVX0 U9299 ( .INP(n9432), .ZN(n9322) );
  INVX0 U9300 ( .INP(n9432), .ZN(n9323) );
  INVX0 U9301 ( .INP(n9432), .ZN(n9324) );
  INVX0 U9302 ( .INP(n9432), .ZN(n9325) );
  INVX0 U9303 ( .INP(n9432), .ZN(n9326) );
  INVX0 U9304 ( .INP(n9432), .ZN(n9327) );
  INVX0 U9305 ( .INP(n9431), .ZN(n9328) );
  INVX0 U9306 ( .INP(n9431), .ZN(n9329) );
  INVX0 U9307 ( .INP(n9431), .ZN(n9330) );
  INVX0 U9308 ( .INP(n9431), .ZN(n9331) );
  INVX0 U9309 ( .INP(n9431), .ZN(n9332) );
  INVX0 U9310 ( .INP(n9431), .ZN(n9333) );
  INVX0 U9311 ( .INP(n9430), .ZN(n9334) );
  INVX0 U9312 ( .INP(n9430), .ZN(n9335) );
  INVX0 U9313 ( .INP(n9430), .ZN(n9336) );
  INVX0 U9314 ( .INP(n9430), .ZN(n9337) );
  INVX0 U9315 ( .INP(n9430), .ZN(n9338) );
  INVX0 U9316 ( .INP(n9430), .ZN(n9339) );
  INVX0 U9317 ( .INP(n9429), .ZN(n9340) );
  INVX0 U9318 ( .INP(n9429), .ZN(n9341) );
  INVX0 U9319 ( .INP(n9429), .ZN(n9342) );
  INVX0 U9320 ( .INP(n9429), .ZN(n9343) );
  INVX0 U9321 ( .INP(n9429), .ZN(n9344) );
  INVX0 U9322 ( .INP(n9429), .ZN(n9345) );
  INVX0 U9323 ( .INP(n9428), .ZN(n9346) );
  INVX0 U9324 ( .INP(n9428), .ZN(n9347) );
  INVX0 U9325 ( .INP(n9428), .ZN(n9348) );
  INVX0 U9326 ( .INP(n9428), .ZN(n9349) );
  INVX0 U9327 ( .INP(n9428), .ZN(n9350) );
  INVX0 U9328 ( .INP(n9428), .ZN(n9351) );
  INVX0 U9329 ( .INP(n9427), .ZN(n9352) );
  INVX0 U9330 ( .INP(n9427), .ZN(n9353) );
  INVX0 U9331 ( .INP(n9427), .ZN(n9354) );
  INVX0 U9332 ( .INP(n9427), .ZN(n9355) );
  INVX0 U9333 ( .INP(n9427), .ZN(n9356) );
  INVX0 U9334 ( .INP(n9427), .ZN(n9357) );
  INVX0 U9335 ( .INP(n9426), .ZN(n9358) );
  INVX0 U9336 ( .INP(n9426), .ZN(n9359) );
  INVX0 U9337 ( .INP(n9426), .ZN(n9360) );
  INVX0 U9338 ( .INP(n9426), .ZN(n9361) );
  INVX0 U9339 ( .INP(n9426), .ZN(n9362) );
  INVX0 U9340 ( .INP(n9426), .ZN(n9363) );
  INVX0 U9341 ( .INP(n9429), .ZN(n9364) );
  INVX0 U9342 ( .INP(n9428), .ZN(n9365) );
  INVX0 U9343 ( .INP(n9427), .ZN(n9366) );
  INVX0 U9344 ( .INP(n9426), .ZN(n9367) );
  INVX0 U9345 ( .INP(n9429), .ZN(n9368) );
  INVX0 U9346 ( .INP(n9433), .ZN(n9369) );
  INVX0 U9347 ( .INP(n9429), .ZN(n9370) );
  INVX0 U9348 ( .INP(n9428), .ZN(n9371) );
  INVX0 U9349 ( .INP(n9427), .ZN(n9372) );
  INVX0 U9350 ( .INP(n9426), .ZN(n9373) );
  INVX0 U9351 ( .INP(n9433), .ZN(n9374) );
  INVX0 U9352 ( .INP(n9428), .ZN(n9375) );
  INVX0 U9353 ( .INP(n9427), .ZN(n9376) );
  INVX0 U9354 ( .INP(n9426), .ZN(n9377) );
  INVX0 U9355 ( .INP(n9432), .ZN(n9378) );
  INVX0 U9356 ( .INP(n9432), .ZN(n9379) );
  INVX0 U9357 ( .INP(n9427), .ZN(n9380) );
  INVX0 U9358 ( .INP(n9433), .ZN(n9381) );
  INVX0 U9359 ( .INP(n9434), .ZN(n9382) );
  INVX0 U9360 ( .INP(n9426), .ZN(n9383) );
  INVX0 U9361 ( .INP(n9433), .ZN(n9384) );
  INVX0 U9362 ( .INP(n9432), .ZN(n9385) );
  INVX0 U9363 ( .INP(n9431), .ZN(n9386) );
  INVX0 U9364 ( .INP(n9430), .ZN(n9387) );
  INVX0 U9365 ( .INP(n9430), .ZN(n9388) );
  INVX0 U9366 ( .INP(n9434), .ZN(n9389) );
  INVX0 U9367 ( .INP(n9429), .ZN(n9390) );
  INVX0 U9368 ( .INP(n9428), .ZN(n9391) );
  INVX0 U9369 ( .INP(n9427), .ZN(n9392) );
  INVX0 U9370 ( .INP(n9431), .ZN(n9393) );
  INVX0 U9371 ( .INP(n9430), .ZN(n9394) );
  INVX0 U9372 ( .INP(n9434), .ZN(n9395) );
  INVX0 U9373 ( .INP(n9433), .ZN(n9396) );
  INVX0 U9374 ( .INP(n9432), .ZN(n9397) );
  INVX0 U9375 ( .INP(n9434), .ZN(n9398) );
  INVX0 U9376 ( .INP(n9429), .ZN(n9399) );
  INVX0 U9377 ( .INP(n9428), .ZN(n9400) );
  INVX0 U9378 ( .INP(n9427), .ZN(n9401) );
  INVX0 U9379 ( .INP(n9426), .ZN(n9402) );
  INVX0 U9380 ( .INP(n9427), .ZN(n9403) );
  INVX0 U9381 ( .INP(n9426), .ZN(n9404) );
  INVX0 U9382 ( .INP(n9430), .ZN(n9405) );
  INVX0 U9383 ( .INP(n9430), .ZN(n9406) );
  INVX0 U9384 ( .INP(n9426), .ZN(n9407) );
  INVX0 U9385 ( .INP(n9428), .ZN(n9408) );
  INVX0 U9386 ( .INP(n9430), .ZN(n9409) );
  INVX0 U9387 ( .INP(n9429), .ZN(n9410) );
  INVX0 U9388 ( .INP(n9428), .ZN(n9411) );
  INVX0 U9389 ( .INP(n9427), .ZN(n9412) );
  INVX0 U9390 ( .INP(n9426), .ZN(n9413) );
  INVX0 U9391 ( .INP(n9431), .ZN(n9414) );
  INVX0 U9392 ( .INP(n9430), .ZN(n9415) );
  INVX0 U9393 ( .INP(n9434), .ZN(n9416) );
  INVX0 U9394 ( .INP(n9433), .ZN(n9417) );
  INVX0 U9395 ( .INP(n9429), .ZN(n9418) );
  INVX0 U9396 ( .INP(n9428), .ZN(n9419) );
  INVX0 U9397 ( .INP(n9431), .ZN(n9420) );
  INVX0 U9398 ( .INP(n9431), .ZN(n9421) );
  INVX0 U9399 ( .INP(n9432), .ZN(n9422) );
  INVX0 U9400 ( .INP(n9432), .ZN(n9423) );
  INVX0 U9401 ( .INP(n9429), .ZN(n9424) );
  INVX0 U9402 ( .INP(n9428), .ZN(n9425) );
  NBUFFX2 U9403 ( .INP(TM1), .Z(n9436) );
  NBUFFX2 U9404 ( .INP(TM1), .Z(n9437) );
  NBUFFX2 U9405 ( .INP(TM1), .Z(n9438) );
  NBUFFX2 U9406 ( .INP(TM1), .Z(n9439) );
  NBUFFX2 U9407 ( .INP(TM1), .Z(n9440) );
  INVX0 U9408 ( .INP(n9455), .ZN(n9441) );
  INVX0 U9409 ( .INP(n9456), .ZN(n9442) );
  INVX0 U9410 ( .INP(n9476), .ZN(n9443) );
  INVX0 U9411 ( .INP(n9457), .ZN(n9444) );
  INVX0 U9412 ( .INP(n9459), .ZN(n9445) );
  INVX0 U9413 ( .INP(n9472), .ZN(n9446) );
  INVX0 U9414 ( .INP(n9453), .ZN(n9447) );
  INVX0 U9415 ( .INP(n9453), .ZN(n9448) );
  INVX0 U9416 ( .INP(n9477), .ZN(n9449) );
  INVX0 U9417 ( .INP(n9454), .ZN(n9450) );
  INVX0 U9418 ( .INP(n9455), .ZN(n9451) );
  INVX0 U9419 ( .INP(n9436), .ZN(n9452) );
  INVX0 U9420 ( .INP(n9436), .ZN(n9453) );
  INVX0 U9421 ( .INP(n9436), .ZN(n9454) );
  INVX0 U9422 ( .INP(n9436), .ZN(n9455) );
  INVX0 U9423 ( .INP(n9436), .ZN(n9456) );
  INVX0 U9424 ( .INP(n9436), .ZN(n9457) );
  INVX0 U9425 ( .INP(n9437), .ZN(n9458) );
  INVX0 U9426 ( .INP(n9437), .ZN(n9459) );
  INVX0 U9427 ( .INP(n9437), .ZN(n9460) );
  INVX0 U9428 ( .INP(n9437), .ZN(n9461) );
  INVX0 U9429 ( .INP(n9437), .ZN(n9462) );
  INVX0 U9430 ( .INP(n9437), .ZN(n9463) );
  INVX0 U9431 ( .INP(n9437), .ZN(n9464) );
  INVX0 U9432 ( .INP(n9437), .ZN(n9465) );
  INVX0 U9433 ( .INP(n9438), .ZN(n9466) );
  INVX0 U9434 ( .INP(n9438), .ZN(n9467) );
  INVX0 U9435 ( .INP(n9438), .ZN(n9468) );
  INVX0 U9436 ( .INP(n9438), .ZN(n9469) );
  INVX0 U9437 ( .INP(n9438), .ZN(n9470) );
  INVX0 U9438 ( .INP(n9438), .ZN(n9471) );
  INVX0 U9439 ( .INP(n9438), .ZN(n9472) );
  INVX0 U9440 ( .INP(n9439), .ZN(n9473) );
  INVX0 U9441 ( .INP(n9439), .ZN(n9474) );
  INVX0 U9442 ( .INP(n9439), .ZN(n9475) );
  INVX0 U9443 ( .INP(n9439), .ZN(n9476) );
  INVX0 U9444 ( .INP(n9439), .ZN(n9477) );
  INVX0 U9445 ( .INP(n9439), .ZN(n9478) );
  INVX0 U9446 ( .INP(n9439), .ZN(n9479) );
  INVX0 U9447 ( .INP(n9439), .ZN(n9480) );
  INVX0 U9448 ( .INP(n9440), .ZN(n9481) );
  INVX0 U9449 ( .INP(n9440), .ZN(n9482) );
  NBUFFX2 U9450 ( .INP(n9550), .Z(n9483) );
  NBUFFX2 U9451 ( .INP(n9550), .Z(n9484) );
  NBUFFX2 U9452 ( .INP(n9550), .Z(n9485) );
  NBUFFX2 U9453 ( .INP(n9549), .Z(n9486) );
  NBUFFX2 U9454 ( .INP(n9549), .Z(n9487) );
  NBUFFX2 U9455 ( .INP(n9549), .Z(n9488) );
  NBUFFX2 U9456 ( .INP(n9548), .Z(n9489) );
  NBUFFX2 U9457 ( .INP(n9548), .Z(n9490) );
  NBUFFX2 U9458 ( .INP(n9548), .Z(n9491) );
  NBUFFX2 U9459 ( .INP(n9547), .Z(n9492) );
  NBUFFX2 U9460 ( .INP(n9547), .Z(n9493) );
  NBUFFX2 U9461 ( .INP(n9547), .Z(n9494) );
  NBUFFX2 U9462 ( .INP(n9546), .Z(n9495) );
  NBUFFX2 U9463 ( .INP(n9546), .Z(n9496) );
  NBUFFX2 U9464 ( .INP(n9546), .Z(n9497) );
  NBUFFX2 U9465 ( .INP(n9545), .Z(n9498) );
  NBUFFX2 U9466 ( .INP(n9545), .Z(n9499) );
  NBUFFX2 U9467 ( .INP(n9545), .Z(n9500) );
  NBUFFX2 U9468 ( .INP(n9544), .Z(n9501) );
  NBUFFX2 U9469 ( .INP(n9544), .Z(n9502) );
  NBUFFX2 U9470 ( .INP(n9544), .Z(n9503) );
  NBUFFX2 U9471 ( .INP(n9543), .Z(n9504) );
  NBUFFX2 U9472 ( .INP(n9543), .Z(n9505) );
  NBUFFX2 U9473 ( .INP(n9543), .Z(n9506) );
  NBUFFX2 U9474 ( .INP(n9542), .Z(n9507) );
  NBUFFX2 U9475 ( .INP(n9542), .Z(n9508) );
  NBUFFX2 U9476 ( .INP(n9542), .Z(n9509) );
  NBUFFX2 U9477 ( .INP(n9541), .Z(n9510) );
  NBUFFX2 U9478 ( .INP(n9541), .Z(n9511) );
  NBUFFX2 U9479 ( .INP(n9541), .Z(n9512) );
  NBUFFX2 U9480 ( .INP(n9540), .Z(n9513) );
  NBUFFX2 U9481 ( .INP(n9540), .Z(n9514) );
  NBUFFX2 U9482 ( .INP(n9540), .Z(n9515) );
  NBUFFX2 U9483 ( .INP(n9539), .Z(n9516) );
  NBUFFX2 U9484 ( .INP(n9539), .Z(n9517) );
  NBUFFX2 U9485 ( .INP(n9539), .Z(n9518) );
  NBUFFX2 U9486 ( .INP(n9538), .Z(n9519) );
  NBUFFX2 U9487 ( .INP(n9538), .Z(n9520) );
  NBUFFX2 U9488 ( .INP(n9538), .Z(n9521) );
  NBUFFX2 U9489 ( .INP(n9537), .Z(n9522) );
  NBUFFX2 U9490 ( .INP(n9537), .Z(n9523) );
  NBUFFX2 U9491 ( .INP(n9537), .Z(n9524) );
  NBUFFX2 U9492 ( .INP(n9536), .Z(n9525) );
  NBUFFX2 U9493 ( .INP(n9536), .Z(n9526) );
  NBUFFX2 U9494 ( .INP(n9536), .Z(n9527) );
  NBUFFX2 U9495 ( .INP(n9535), .Z(n9528) );
  NBUFFX2 U9496 ( .INP(n9535), .Z(n9529) );
  NBUFFX2 U9497 ( .INP(n9535), .Z(n9530) );
  NBUFFX2 U9498 ( .INP(n9534), .Z(n9531) );
  NBUFFX2 U9499 ( .INP(n9534), .Z(n9532) );
  NBUFFX2 U9500 ( .INP(n9534), .Z(n9533) );
  NBUFFX2 U9501 ( .INP(n9556), .Z(n9534) );
  NBUFFX2 U9502 ( .INP(n9556), .Z(n9535) );
  NBUFFX2 U9503 ( .INP(n9555), .Z(n9536) );
  NBUFFX2 U9504 ( .INP(n9555), .Z(n9537) );
  NBUFFX2 U9505 ( .INP(n9555), .Z(n9538) );
  NBUFFX2 U9506 ( .INP(n9554), .Z(n9539) );
  NBUFFX2 U9507 ( .INP(n9554), .Z(n9540) );
  NBUFFX2 U9508 ( .INP(n9554), .Z(n9541) );
  NBUFFX2 U9509 ( .INP(n9553), .Z(n9542) );
  NBUFFX2 U9510 ( .INP(n9553), .Z(n9543) );
  NBUFFX2 U9511 ( .INP(n9553), .Z(n9544) );
  NBUFFX2 U9512 ( .INP(n9552), .Z(n9545) );
  NBUFFX2 U9513 ( .INP(n9552), .Z(n9546) );
  NBUFFX2 U9514 ( .INP(n9552), .Z(n9547) );
  NBUFFX2 U9515 ( .INP(n9551), .Z(n9548) );
  NBUFFX2 U9516 ( .INP(n9551), .Z(n9549) );
  NBUFFX2 U9517 ( .INP(n9551), .Z(n9550) );
  NBUFFX2 U9518 ( .INP(RESET), .Z(n9551) );
  NBUFFX2 U9519 ( .INP(RESET), .Z(n9552) );
  NBUFFX2 U9520 ( .INP(RESET), .Z(n9553) );
  NBUFFX2 U9521 ( .INP(RESET), .Z(n9554) );
  NBUFFX2 U9522 ( .INP(RESET), .Z(n9555) );
  NBUFFX2 U9523 ( .INP(RESET), .Z(n9556) );
  INVX0 U9524 ( .INP(n9483), .ZN(n9557) );
  INVX0 U9525 ( .INP(n9483), .ZN(n9558) );
  INVX0 U9526 ( .INP(n9483), .ZN(n9559) );
  INVX0 U9527 ( .INP(n9483), .ZN(n9560) );
  INVX0 U9528 ( .INP(n9483), .ZN(n9561) );
  INVX0 U9529 ( .INP(n9483), .ZN(n9562) );
  INVX0 U9530 ( .INP(n9483), .ZN(n9563) );
  INVX0 U9531 ( .INP(n9484), .ZN(n9564) );
  INVX0 U9532 ( .INP(n9484), .ZN(n9565) );
  INVX0 U9533 ( .INP(n9484), .ZN(n9566) );
  INVX0 U9534 ( .INP(n9484), .ZN(n9567) );
  INVX0 U9535 ( .INP(n9484), .ZN(n9568) );
  INVX0 U9536 ( .INP(n9484), .ZN(n9569) );
  INVX0 U9537 ( .INP(n9484), .ZN(n9570) );
  INVX0 U9538 ( .INP(n9484), .ZN(n9571) );
  INVX0 U9539 ( .INP(n9485), .ZN(n9572) );
  INVX0 U9540 ( .INP(n9485), .ZN(n9573) );
  INVX0 U9541 ( .INP(n9489), .ZN(n9574) );
  INVX0 U9542 ( .INP(n9485), .ZN(n9575) );
  INVX0 U9543 ( .INP(n9485), .ZN(n9576) );
  INVX0 U9544 ( .INP(n9485), .ZN(n9577) );
  INVX0 U9545 ( .INP(n9485), .ZN(n9578) );
  INVX0 U9546 ( .INP(n9485), .ZN(n9579) );
  INVX0 U9547 ( .INP(n9485), .ZN(n9580) );
  INVX0 U9548 ( .INP(n9486), .ZN(n9581) );
  INVX0 U9549 ( .INP(n9486), .ZN(n9582) );
  INVX0 U9550 ( .INP(n9486), .ZN(n9583) );
  INVX0 U9551 ( .INP(n9486), .ZN(n9584) );
  INVX0 U9552 ( .INP(n9486), .ZN(n9585) );
  INVX0 U9553 ( .INP(n9486), .ZN(n9586) );
  INVX0 U9554 ( .INP(n9486), .ZN(n9587) );
  INVX0 U9555 ( .INP(n9486), .ZN(n9588) );
  INVX0 U9556 ( .INP(n9487), .ZN(n9589) );
  INVX0 U9557 ( .INP(n9487), .ZN(n9590) );
  INVX0 U9558 ( .INP(n9487), .ZN(n9591) );
  INVX0 U9559 ( .INP(n9487), .ZN(n9592) );
  INVX0 U9560 ( .INP(n9487), .ZN(n9593) );
  INVX0 U9561 ( .INP(n9487), .ZN(n9594) );
  INVX0 U9562 ( .INP(n9487), .ZN(n9595) );
  INVX0 U9563 ( .INP(n9487), .ZN(n9596) );
  INVX0 U9564 ( .INP(n9488), .ZN(n9597) );
  INVX0 U9565 ( .INP(n9488), .ZN(n9598) );
  INVX0 U9566 ( .INP(n9488), .ZN(n9599) );
  INVX0 U9567 ( .INP(n9488), .ZN(n9600) );
  INVX0 U9568 ( .INP(n9488), .ZN(n9601) );
  INVX0 U9569 ( .INP(n9488), .ZN(n9602) );
  INVX0 U9570 ( .INP(n9488), .ZN(n9603) );
  INVX0 U9571 ( .INP(n9488), .ZN(n9604) );
  INVX0 U9572 ( .INP(n9489), .ZN(n9605) );
  INVX0 U9573 ( .INP(n9489), .ZN(n9606) );
  INVX0 U9574 ( .INP(n9489), .ZN(n9607) );
  INVX0 U9575 ( .INP(n9489), .ZN(n9608) );
  INVX0 U9576 ( .INP(n9490), .ZN(n9609) );
  INVX0 U9577 ( .INP(n9490), .ZN(n9610) );
  INVX0 U9578 ( .INP(n9489), .ZN(n9611) );
  INVX0 U9579 ( .INP(n9491), .ZN(n9612) );
  INVX0 U9580 ( .INP(n9490), .ZN(n9613) );
  INVX0 U9581 ( .INP(n9491), .ZN(n9614) );
  INVX0 U9582 ( .INP(n9490), .ZN(n9615) );
  INVX0 U9583 ( .INP(n9491), .ZN(n9616) );
  INVX0 U9584 ( .INP(n9491), .ZN(n9617) );
  INVX0 U9585 ( .INP(n9491), .ZN(n9618) );
  INVX0 U9586 ( .INP(n9489), .ZN(n9619) );
  INVX0 U9587 ( .INP(n9491), .ZN(n9620) );
  INVX0 U9588 ( .INP(n9489), .ZN(n9621) );
  INVX0 U9589 ( .INP(n9491), .ZN(n9622) );
  INVX0 U9590 ( .INP(n9491), .ZN(n9623) );
  INVX0 U9591 ( .INP(n9490), .ZN(n9624) );
  INVX0 U9592 ( .INP(n9490), .ZN(n9625) );
  INVX0 U9593 ( .INP(n9492), .ZN(n9626) );
  INVX0 U9594 ( .INP(n9492), .ZN(n9627) );
  INVX0 U9595 ( .INP(n9490), .ZN(n9628) );
  INVX0 U9596 ( .INP(n9492), .ZN(n9629) );
  INVX0 U9597 ( .INP(n9490), .ZN(n9630) );
  INVX0 U9598 ( .INP(n9492), .ZN(n9631) );
  INVX0 U9599 ( .INP(n9483), .ZN(n9632) );
  NBUFFX2 U9600 ( .INP(n9815), .Z(n9777) );
  NBUFFX2 U9601 ( .INP(n9815), .Z(n9778) );
  NBUFFX2 U9602 ( .INP(n9814), .Z(n9779) );
  NBUFFX2 U9603 ( .INP(n9814), .Z(n9780) );
  NBUFFX2 U9604 ( .INP(n9814), .Z(n9781) );
  NBUFFX2 U9605 ( .INP(n9813), .Z(n9782) );
  NBUFFX2 U9606 ( .INP(n9813), .Z(n9783) );
  NBUFFX2 U9607 ( .INP(n9813), .Z(n9784) );
  NBUFFX2 U9608 ( .INP(n9812), .Z(n9785) );
  NBUFFX2 U9609 ( .INP(n9812), .Z(n9786) );
  NBUFFX2 U9610 ( .INP(n9812), .Z(n9787) );
  NBUFFX2 U9611 ( .INP(n9811), .Z(n9788) );
  NBUFFX2 U9612 ( .INP(n9811), .Z(n9789) );
  NBUFFX2 U9613 ( .INP(n9811), .Z(n9790) );
  NBUFFX2 U9614 ( .INP(n9810), .Z(n9791) );
  NBUFFX2 U9615 ( .INP(n9810), .Z(n9792) );
  NBUFFX2 U9616 ( .INP(n9810), .Z(n9793) );
  NBUFFX2 U9617 ( .INP(n9809), .Z(n9794) );
  NBUFFX2 U9618 ( .INP(n9809), .Z(n9795) );
  NBUFFX2 U9619 ( .INP(n9809), .Z(n9796) );
  NBUFFX2 U9620 ( .INP(n9808), .Z(n9797) );
  NBUFFX2 U9621 ( .INP(n9808), .Z(n9798) );
  NBUFFX2 U9622 ( .INP(n9808), .Z(n9799) );
  NBUFFX2 U9623 ( .INP(n9807), .Z(n9800) );
  NBUFFX2 U9624 ( .INP(n9807), .Z(n9801) );
  NBUFFX2 U9625 ( .INP(n9807), .Z(n9802) );
  NBUFFX2 U9626 ( .INP(n9806), .Z(n9803) );
  NBUFFX2 U9627 ( .INP(n9806), .Z(n9804) );
  NBUFFX2 U9628 ( .INP(n9806), .Z(n9805) );
  NBUFFX2 U9629 ( .INP(CK), .Z(n9806) );
  NBUFFX2 U9630 ( .INP(CK), .Z(n9807) );
  NBUFFX2 U9631 ( .INP(n9815), .Z(n9808) );
  NBUFFX2 U9632 ( .INP(CK), .Z(n9809) );
  NBUFFX2 U9633 ( .INP(n9811), .Z(n9810) );
  NBUFFX2 U9634 ( .INP(CK), .Z(n9811) );
  NBUFFX2 U9635 ( .INP(n9806), .Z(n9812) );
  NBUFFX2 U9636 ( .INP(n9807), .Z(n9813) );
  NBUFFX2 U9637 ( .INP(n9809), .Z(n9814) );
  NBUFFX2 U9638 ( .INP(n9646), .Z(n9815) );
  AND2X1 U9639 ( .IN1(n9510), .IN2(n9478), .Q(n3278) );
  AND2X1 U9640 ( .IN1(n9510), .IN2(n8304), .Q(WX9789) );
  AND2X1 U9641 ( .IN1(n9510), .IN2(n8305), .Q(WX9787) );
  AND2X1 U9642 ( .IN1(n9510), .IN2(n8306), .Q(WX9785) );
  AND2X1 U9643 ( .IN1(n9508), .IN2(n8307), .Q(WX9783) );
  AND2X1 U9644 ( .IN1(test_so80), .IN2(n9497), .Q(WX9781) );
  AND2X1 U9645 ( .IN1(n9508), .IN2(n8310), .Q(WX9779) );
  AND2X1 U9646 ( .IN1(n9508), .IN2(n8311), .Q(WX9777) );
  AND2X1 U9647 ( .IN1(n9511), .IN2(n8312), .Q(WX9775) );
  AND2X1 U9648 ( .IN1(n9508), .IN2(n8313), .Q(WX9773) );
  AND2X1 U9649 ( .IN1(n9508), .IN2(n8314), .Q(WX9771) );
  AND2X1 U9650 ( .IN1(n9509), .IN2(n8315), .Q(WX9769) );
  AND2X1 U9651 ( .IN1(n9509), .IN2(n8316), .Q(WX9767) );
  AND2X1 U9652 ( .IN1(n9509), .IN2(n8317), .Q(WX9765) );
  AND2X1 U9653 ( .IN1(n9509), .IN2(n8318), .Q(WX9763) );
  AND2X1 U9654 ( .IN1(n9509), .IN2(n8319), .Q(WX9761) );
  AND2X1 U9655 ( .IN1(n9510), .IN2(n8320), .Q(WX9759) );
  OR4X1 U9656 ( .IN1(n9816), .IN2(n9817), .IN3(n9818), .IN4(n9819), .Q(WX9757)
         );
  AND2X1 U9657 ( .IN1(n9266), .IN2(n9820), .Q(n9819) );
  AND2X1 U9658 ( .IN1(n9185), .IN2(n9822), .Q(n9818) );
  AND2X1 U9659 ( .IN1(n9229), .IN2(CRC_OUT_2_0), .Q(n9817) );
  AND2X1 U9660 ( .IN1(n9224), .IN2(n1744), .Q(n9816) );
  INVX0 U9661 ( .INP(n9823), .ZN(n1744) );
  OR2X1 U9662 ( .IN1(n9577), .IN2(n3817), .Q(n9823) );
  OR4X1 U9663 ( .IN1(n9824), .IN2(n9825), .IN3(n9826), .IN4(n9827), .Q(WX9755)
         );
  AND2X1 U9664 ( .IN1(n9274), .IN2(n9828), .Q(n9827) );
  AND2X1 U9665 ( .IN1(n9829), .IN2(n9173), .Q(n9826) );
  AND2X1 U9666 ( .IN1(n9243), .IN2(CRC_OUT_2_1), .Q(n9825) );
  AND2X1 U9667 ( .IN1(n1743), .IN2(n9212), .Q(n9824) );
  INVX0 U9668 ( .INP(n9830), .ZN(n1743) );
  OR2X1 U9669 ( .IN1(n9577), .IN2(n3818), .Q(n9830) );
  OR4X1 U9670 ( .IN1(n9831), .IN2(n9832), .IN3(n9833), .IN4(n9834), .Q(WX9753)
         );
  AND2X1 U9671 ( .IN1(n9835), .IN2(n9261), .Q(n9834) );
  AND2X1 U9672 ( .IN1(n9185), .IN2(n9836), .Q(n9833) );
  AND2X1 U9673 ( .IN1(test_so87), .IN2(n9227), .Q(n9832) );
  AND2X1 U9674 ( .IN1(n1742), .IN2(n9212), .Q(n9831) );
  INVX0 U9675 ( .INP(n9837), .ZN(n1742) );
  OR2X1 U9676 ( .IN1(n9577), .IN2(n3819), .Q(n9837) );
  OR4X1 U9677 ( .IN1(n9838), .IN2(n9839), .IN3(n9840), .IN4(n9841), .Q(WX9751)
         );
  AND2X1 U9678 ( .IN1(n9270), .IN2(n9842), .Q(n9841) );
  AND2X1 U9679 ( .IN1(n9843), .IN2(n9173), .Q(n9840) );
  AND2X1 U9680 ( .IN1(n9238), .IN2(CRC_OUT_2_3), .Q(n9839) );
  AND2X1 U9681 ( .IN1(n1741), .IN2(n9212), .Q(n9838) );
  INVX0 U9682 ( .INP(n9844), .ZN(n1741) );
  OR2X1 U9683 ( .IN1(n9577), .IN2(n3820), .Q(n9844) );
  OR4X1 U9684 ( .IN1(n9845), .IN2(n9846), .IN3(n9847), .IN4(n9848), .Q(WX9749)
         );
  AND2X1 U9685 ( .IN1(n9849), .IN2(n9261), .Q(n9848) );
  AND2X1 U9686 ( .IN1(n9185), .IN2(n9850), .Q(n9847) );
  AND2X1 U9687 ( .IN1(n9238), .IN2(CRC_OUT_2_4), .Q(n9846) );
  AND2X1 U9688 ( .IN1(n1740), .IN2(n9212), .Q(n9845) );
  INVX0 U9689 ( .INP(n9851), .ZN(n1740) );
  OR2X1 U9690 ( .IN1(n9577), .IN2(n3821), .Q(n9851) );
  OR4X1 U9691 ( .IN1(n9852), .IN2(n9853), .IN3(n9854), .IN4(n9855), .Q(WX9747)
         );
  AND2X1 U9692 ( .IN1(n9270), .IN2(n9856), .Q(n9855) );
  AND2X1 U9693 ( .IN1(n9185), .IN2(n9857), .Q(n9854) );
  AND2X1 U9694 ( .IN1(n9238), .IN2(CRC_OUT_2_5), .Q(n9853) );
  AND2X1 U9695 ( .IN1(n1739), .IN2(n9213), .Q(n9852) );
  INVX0 U9696 ( .INP(n9858), .ZN(n1739) );
  OR2X1 U9697 ( .IN1(n9577), .IN2(n3822), .Q(n9858) );
  OR4X1 U9698 ( .IN1(n9859), .IN2(n9860), .IN3(n9861), .IN4(n9862), .Q(WX9745)
         );
  AND2X1 U9699 ( .IN1(n9863), .IN2(n9262), .Q(n9862) );
  AND2X1 U9700 ( .IN1(n9185), .IN2(n9864), .Q(n9861) );
  AND2X1 U9701 ( .IN1(n9238), .IN2(CRC_OUT_2_6), .Q(n9860) );
  AND2X1 U9702 ( .IN1(n1738), .IN2(n9213), .Q(n9859) );
  INVX0 U9703 ( .INP(n9865), .ZN(n1738) );
  OR2X1 U9704 ( .IN1(n9577), .IN2(n3823), .Q(n9865) );
  OR4X1 U9705 ( .IN1(n9866), .IN2(n9867), .IN3(n9868), .IN4(n9869), .Q(WX9743)
         );
  AND2X1 U9706 ( .IN1(n9270), .IN2(n9870), .Q(n9869) );
  AND2X1 U9707 ( .IN1(n9185), .IN2(n9871), .Q(n9868) );
  AND2X1 U9708 ( .IN1(n9238), .IN2(CRC_OUT_2_7), .Q(n9867) );
  AND2X1 U9709 ( .IN1(n1737), .IN2(n9213), .Q(n9866) );
  INVX0 U9710 ( .INP(n9872), .ZN(n1737) );
  OR2X1 U9711 ( .IN1(n9577), .IN2(n3824), .Q(n9872) );
  OR4X1 U9712 ( .IN1(n9873), .IN2(n9874), .IN3(n9875), .IN4(n9876), .Q(WX9741)
         );
  AND2X1 U9713 ( .IN1(n9877), .IN2(n9262), .Q(n9876) );
  AND2X1 U9714 ( .IN1(n9185), .IN2(n9878), .Q(n9875) );
  AND2X1 U9715 ( .IN1(n9239), .IN2(CRC_OUT_2_8), .Q(n9874) );
  AND2X1 U9716 ( .IN1(n1736), .IN2(n9213), .Q(n9873) );
  INVX0 U9717 ( .INP(n9879), .ZN(n1736) );
  OR2X1 U9718 ( .IN1(n9576), .IN2(n3825), .Q(n9879) );
  OR4X1 U9719 ( .IN1(n9880), .IN2(n9881), .IN3(n9882), .IN4(n9883), .Q(WX9739)
         );
  AND2X1 U9720 ( .IN1(n9270), .IN2(n9884), .Q(n9883) );
  AND2X1 U9721 ( .IN1(n9185), .IN2(n9885), .Q(n9882) );
  AND2X1 U9722 ( .IN1(n9239), .IN2(CRC_OUT_2_9), .Q(n9881) );
  AND2X1 U9723 ( .IN1(n1735), .IN2(n9213), .Q(n9880) );
  INVX0 U9724 ( .INP(n9886), .ZN(n1735) );
  OR2X1 U9725 ( .IN1(n9576), .IN2(n3826), .Q(n9886) );
  OR4X1 U9726 ( .IN1(n9887), .IN2(n9888), .IN3(n9889), .IN4(n9890), .Q(WX9737)
         );
  AND2X1 U9727 ( .IN1(n9270), .IN2(n9891), .Q(n9890) );
  AND2X1 U9728 ( .IN1(n9185), .IN2(n9892), .Q(n9889) );
  AND2X1 U9729 ( .IN1(n9239), .IN2(CRC_OUT_2_10), .Q(n9888) );
  AND2X1 U9730 ( .IN1(n1734), .IN2(n9213), .Q(n9887) );
  INVX0 U9731 ( .INP(n9893), .ZN(n1734) );
  OR2X1 U9732 ( .IN1(n9576), .IN2(n3827), .Q(n9893) );
  OR4X1 U9733 ( .IN1(n9894), .IN2(n9895), .IN3(n9896), .IN4(n9897), .Q(WX9735)
         );
  AND2X1 U9734 ( .IN1(n9270), .IN2(n9898), .Q(n9897) );
  AND2X1 U9735 ( .IN1(n9185), .IN2(n9899), .Q(n9896) );
  AND2X1 U9736 ( .IN1(n9239), .IN2(CRC_OUT_2_11), .Q(n9895) );
  AND2X1 U9737 ( .IN1(n1733), .IN2(n9213), .Q(n9894) );
  INVX0 U9738 ( .INP(n9900), .ZN(n1733) );
  OR2X1 U9739 ( .IN1(n9576), .IN2(n3828), .Q(n9900) );
  OR4X1 U9740 ( .IN1(n9901), .IN2(n9902), .IN3(n9903), .IN4(n9904), .Q(WX9733)
         );
  AND2X1 U9741 ( .IN1(n9270), .IN2(n9905), .Q(n9904) );
  AND2X1 U9742 ( .IN1(n9185), .IN2(n9906), .Q(n9903) );
  AND2X1 U9743 ( .IN1(n9239), .IN2(CRC_OUT_2_12), .Q(n9902) );
  AND2X1 U9744 ( .IN1(n1732), .IN2(n9213), .Q(n9901) );
  INVX0 U9745 ( .INP(n9907), .ZN(n1732) );
  OR2X1 U9746 ( .IN1(n9576), .IN2(n3829), .Q(n9907) );
  OR4X1 U9747 ( .IN1(n9908), .IN2(n9909), .IN3(n9910), .IN4(n9911), .Q(WX9731)
         );
  AND2X1 U9748 ( .IN1(n9270), .IN2(n9912), .Q(n9911) );
  AND2X1 U9749 ( .IN1(n9185), .IN2(n9913), .Q(n9910) );
  AND2X1 U9750 ( .IN1(n9239), .IN2(CRC_OUT_2_13), .Q(n9909) );
  AND2X1 U9751 ( .IN1(n1731), .IN2(n9213), .Q(n9908) );
  INVX0 U9752 ( .INP(n9914), .ZN(n1731) );
  OR2X1 U9753 ( .IN1(n9576), .IN2(n3830), .Q(n9914) );
  OR4X1 U9754 ( .IN1(n9915), .IN2(n9916), .IN3(n9917), .IN4(n9918), .Q(WX9729)
         );
  AND2X1 U9755 ( .IN1(n9270), .IN2(n9919), .Q(n9918) );
  AND2X1 U9756 ( .IN1(n9920), .IN2(n9174), .Q(n9917) );
  AND2X1 U9757 ( .IN1(n9239), .IN2(CRC_OUT_2_14), .Q(n9916) );
  AND2X1 U9758 ( .IN1(n1730), .IN2(n9213), .Q(n9915) );
  INVX0 U9759 ( .INP(n9921), .ZN(n1730) );
  OR2X1 U9760 ( .IN1(n9576), .IN2(n3831), .Q(n9921) );
  OR4X1 U9761 ( .IN1(n9922), .IN2(n9923), .IN3(n9924), .IN4(n9925), .Q(WX9727)
         );
  AND2X1 U9762 ( .IN1(n9270), .IN2(n9926), .Q(n9925) );
  AND2X1 U9763 ( .IN1(n9184), .IN2(n9927), .Q(n9924) );
  AND2X1 U9764 ( .IN1(n9239), .IN2(CRC_OUT_2_15), .Q(n9923) );
  AND2X1 U9765 ( .IN1(n1729), .IN2(n9213), .Q(n9922) );
  INVX0 U9766 ( .INP(n9928), .ZN(n1729) );
  OR2X1 U9767 ( .IN1(n9576), .IN2(n3832), .Q(n9928) );
  OR4X1 U9768 ( .IN1(n9929), .IN2(n9930), .IN3(n9931), .IN4(n9932), .Q(WX9725)
         );
  AND2X1 U9769 ( .IN1(n9270), .IN2(n9933), .Q(n9932) );
  AND2X1 U9770 ( .IN1(n9934), .IN2(n9174), .Q(n9931) );
  AND2X1 U9771 ( .IN1(n9239), .IN2(CRC_OUT_2_16), .Q(n9930) );
  AND2X1 U9772 ( .IN1(n1728), .IN2(n9213), .Q(n9929) );
  INVX0 U9773 ( .INP(n9935), .ZN(n1728) );
  OR2X1 U9774 ( .IN1(n9576), .IN2(n3833), .Q(n9935) );
  OR4X1 U9775 ( .IN1(n9936), .IN2(n9937), .IN3(n9938), .IN4(n9939), .Q(WX9723)
         );
  AND2X1 U9776 ( .IN1(n9271), .IN2(n9940), .Q(n9939) );
  AND2X1 U9777 ( .IN1(n9184), .IN2(n9941), .Q(n9938) );
  AND2X1 U9778 ( .IN1(n9239), .IN2(CRC_OUT_2_17), .Q(n9937) );
  AND2X1 U9779 ( .IN1(n1727), .IN2(n9214), .Q(n9936) );
  INVX0 U9780 ( .INP(n9942), .ZN(n1727) );
  OR2X1 U9781 ( .IN1(n9576), .IN2(n3834), .Q(n9942) );
  OR4X1 U9782 ( .IN1(n9943), .IN2(n9944), .IN3(n9945), .IN4(n9946), .Q(WX9721)
         );
  AND2X1 U9783 ( .IN1(n9271), .IN2(n9947), .Q(n9946) );
  AND2X1 U9784 ( .IN1(n9948), .IN2(n9174), .Q(n9945) );
  AND2X1 U9785 ( .IN1(n9239), .IN2(CRC_OUT_2_18), .Q(n9944) );
  AND2X1 U9786 ( .IN1(n1726), .IN2(n9214), .Q(n9943) );
  INVX0 U9787 ( .INP(n9949), .ZN(n1726) );
  OR2X1 U9788 ( .IN1(n9576), .IN2(n3835), .Q(n9949) );
  OR4X1 U9789 ( .IN1(n9950), .IN2(n9951), .IN3(n9952), .IN4(n9953), .Q(WX9719)
         );
  AND2X1 U9790 ( .IN1(n9954), .IN2(n9264), .Q(n9953) );
  AND2X1 U9791 ( .IN1(n9184), .IN2(n9955), .Q(n9952) );
  AND2X1 U9792 ( .IN1(test_so88), .IN2(n9227), .Q(n9951) );
  AND2X1 U9793 ( .IN1(n1725), .IN2(n9214), .Q(n9950) );
  INVX0 U9794 ( .INP(n9956), .ZN(n1725) );
  OR2X1 U9795 ( .IN1(n9576), .IN2(n3836), .Q(n9956) );
  OR4X1 U9796 ( .IN1(n9957), .IN2(n9958), .IN3(n9959), .IN4(n9960), .Q(WX9717)
         );
  AND2X1 U9797 ( .IN1(n9271), .IN2(n9961), .Q(n9960) );
  AND2X1 U9798 ( .IN1(n9962), .IN2(n9174), .Q(n9959) );
  AND2X1 U9799 ( .IN1(n9239), .IN2(CRC_OUT_2_20), .Q(n9958) );
  AND2X1 U9800 ( .IN1(n1724), .IN2(n9214), .Q(n9957) );
  INVX0 U9801 ( .INP(n9963), .ZN(n1724) );
  OR2X1 U9802 ( .IN1(n9575), .IN2(n3837), .Q(n9963) );
  OR4X1 U9803 ( .IN1(n9964), .IN2(n9965), .IN3(n9966), .IN4(n9967), .Q(WX9715)
         );
  AND2X1 U9804 ( .IN1(n9968), .IN2(n9263), .Q(n9967) );
  AND2X1 U9805 ( .IN1(n9184), .IN2(n9969), .Q(n9966) );
  AND2X1 U9806 ( .IN1(n9239), .IN2(CRC_OUT_2_21), .Q(n9965) );
  AND2X1 U9807 ( .IN1(n1723), .IN2(n9214), .Q(n9964) );
  INVX0 U9808 ( .INP(n9970), .ZN(n1723) );
  OR2X1 U9809 ( .IN1(n9575), .IN2(n3838), .Q(n9970) );
  OR4X1 U9810 ( .IN1(n9971), .IN2(n9972), .IN3(n9973), .IN4(n9974), .Q(WX9713)
         );
  AND2X1 U9811 ( .IN1(n9271), .IN2(n9975), .Q(n9974) );
  AND2X1 U9812 ( .IN1(n9184), .IN2(n9976), .Q(n9973) );
  AND2X1 U9813 ( .IN1(n9240), .IN2(CRC_OUT_2_22), .Q(n9972) );
  AND2X1 U9814 ( .IN1(n1722), .IN2(n9214), .Q(n9971) );
  INVX0 U9815 ( .INP(n9977), .ZN(n1722) );
  OR2X1 U9816 ( .IN1(n9575), .IN2(n3839), .Q(n9977) );
  OR4X1 U9817 ( .IN1(n9978), .IN2(n9979), .IN3(n9980), .IN4(n9981), .Q(WX9711)
         );
  AND2X1 U9818 ( .IN1(n9982), .IN2(n9264), .Q(n9981) );
  AND2X1 U9819 ( .IN1(n9184), .IN2(n9983), .Q(n9980) );
  AND2X1 U9820 ( .IN1(n9240), .IN2(CRC_OUT_2_23), .Q(n9979) );
  AND2X1 U9821 ( .IN1(n1721), .IN2(n9214), .Q(n9978) );
  INVX0 U9822 ( .INP(n9984), .ZN(n1721) );
  OR2X1 U9823 ( .IN1(n9575), .IN2(n3840), .Q(n9984) );
  OR4X1 U9824 ( .IN1(n9985), .IN2(n9986), .IN3(n9987), .IN4(n9988), .Q(WX9709)
         );
  AND2X1 U9825 ( .IN1(n9271), .IN2(n9989), .Q(n9988) );
  AND2X1 U9826 ( .IN1(n9184), .IN2(n9990), .Q(n9987) );
  AND2X1 U9827 ( .IN1(n9240), .IN2(CRC_OUT_2_24), .Q(n9986) );
  AND2X1 U9828 ( .IN1(n1720), .IN2(n9214), .Q(n9985) );
  INVX0 U9829 ( .INP(n9991), .ZN(n1720) );
  OR2X1 U9830 ( .IN1(n9575), .IN2(n3841), .Q(n9991) );
  OR4X1 U9831 ( .IN1(n9992), .IN2(n9993), .IN3(n9994), .IN4(n9995), .Q(WX9707)
         );
  AND2X1 U9832 ( .IN1(n9996), .IN2(n9263), .Q(n9995) );
  AND2X1 U9833 ( .IN1(n9184), .IN2(n9997), .Q(n9994) );
  AND2X1 U9834 ( .IN1(n9240), .IN2(CRC_OUT_2_25), .Q(n9993) );
  AND2X1 U9835 ( .IN1(n1719), .IN2(n9214), .Q(n9992) );
  INVX0 U9836 ( .INP(n9998), .ZN(n1719) );
  OR2X1 U9837 ( .IN1(n9575), .IN2(n3842), .Q(n9998) );
  OR4X1 U9838 ( .IN1(n9999), .IN2(n10000), .IN3(n10001), .IN4(n10002), .Q(
        WX9705) );
  AND2X1 U9839 ( .IN1(n9271), .IN2(n10003), .Q(n10002) );
  AND2X1 U9840 ( .IN1(n9184), .IN2(n10004), .Q(n10001) );
  AND2X1 U9841 ( .IN1(n9240), .IN2(CRC_OUT_2_26), .Q(n10000) );
  AND2X1 U9842 ( .IN1(n1718), .IN2(n9214), .Q(n9999) );
  INVX0 U9843 ( .INP(n10005), .ZN(n1718) );
  OR2X1 U9844 ( .IN1(n9575), .IN2(n3843), .Q(n10005) );
  OR4X1 U9845 ( .IN1(n10006), .IN2(n10007), .IN3(n10008), .IN4(n10009), .Q(
        WX9703) );
  AND2X1 U9846 ( .IN1(n9271), .IN2(n10010), .Q(n10009) );
  AND2X1 U9847 ( .IN1(n9184), .IN2(n10011), .Q(n10008) );
  AND2X1 U9848 ( .IN1(n9240), .IN2(CRC_OUT_2_27), .Q(n10007) );
  AND2X1 U9849 ( .IN1(n1717), .IN2(n9214), .Q(n10006) );
  INVX0 U9850 ( .INP(n10012), .ZN(n1717) );
  OR2X1 U9851 ( .IN1(n9575), .IN2(n3844), .Q(n10012) );
  OR4X1 U9852 ( .IN1(n10013), .IN2(n10014), .IN3(n10015), .IN4(n10016), .Q(
        WX9701) );
  AND2X1 U9853 ( .IN1(n9271), .IN2(n10017), .Q(n10016) );
  AND2X1 U9854 ( .IN1(n9184), .IN2(n10018), .Q(n10015) );
  AND2X1 U9855 ( .IN1(n9240), .IN2(CRC_OUT_2_28), .Q(n10014) );
  AND2X1 U9856 ( .IN1(n1716), .IN2(n9214), .Q(n10013) );
  INVX0 U9857 ( .INP(n10019), .ZN(n1716) );
  OR2X1 U9858 ( .IN1(n9575), .IN2(n3845), .Q(n10019) );
  OR4X1 U9859 ( .IN1(n10020), .IN2(n10021), .IN3(n10022), .IN4(n10023), .Q(
        WX9699) );
  AND2X1 U9860 ( .IN1(n9271), .IN2(n10024), .Q(n10023) );
  AND2X1 U9861 ( .IN1(n9184), .IN2(n10025), .Q(n10022) );
  AND2X1 U9862 ( .IN1(n9240), .IN2(CRC_OUT_2_29), .Q(n10021) );
  AND2X1 U9863 ( .IN1(n1715), .IN2(n9215), .Q(n10020) );
  INVX0 U9864 ( .INP(n10026), .ZN(n1715) );
  OR2X1 U9865 ( .IN1(n9575), .IN2(n3846), .Q(n10026) );
  OR4X1 U9866 ( .IN1(n10027), .IN2(n10028), .IN3(n10029), .IN4(n10030), .Q(
        WX9697) );
  AND2X1 U9867 ( .IN1(n9271), .IN2(n10031), .Q(n10030) );
  AND2X1 U9868 ( .IN1(n9184), .IN2(n10032), .Q(n10029) );
  AND2X1 U9869 ( .IN1(n9240), .IN2(CRC_OUT_2_30), .Q(n10028) );
  AND2X1 U9870 ( .IN1(n1714), .IN2(n9215), .Q(n10027) );
  INVX0 U9871 ( .INP(n10033), .ZN(n1714) );
  OR2X1 U9872 ( .IN1(n9575), .IN2(n3847), .Q(n10033) );
  OR4X1 U9873 ( .IN1(n10034), .IN2(n10035), .IN3(n10036), .IN4(n10037), .Q(
        WX9695) );
  AND2X1 U9874 ( .IN1(n9271), .IN2(n10038), .Q(n10037) );
  AND2X1 U9875 ( .IN1(n10039), .IN2(n9176), .Q(n10036) );
  AND2X1 U9876 ( .IN1(n2245), .IN2(WX9536), .Q(n10035) );
  AND2X1 U9877 ( .IN1(n9240), .IN2(CRC_OUT_2_31), .Q(n10034) );
  AND2X1 U9878 ( .IN1(n9051), .IN2(n9496), .Q(WX9597) );
  AND3X1 U9879 ( .IN1(n10040), .IN2(n10041), .IN3(n9515), .Q(WX9084) );
  OR2X1 U9880 ( .IN1(DFF_1342_n1), .IN2(WX8595), .Q(n10041) );
  OR2X1 U9881 ( .IN1(n8794), .IN2(CRC_OUT_3_30), .Q(n10040) );
  AND3X1 U9882 ( .IN1(n10042), .IN2(n10043), .IN3(n9514), .Q(WX9082) );
  OR2X1 U9883 ( .IN1(DFF_1341_n1), .IN2(WX8597), .Q(n10043) );
  OR2X1 U9884 ( .IN1(n8795), .IN2(CRC_OUT_3_29), .Q(n10042) );
  AND3X1 U9885 ( .IN1(n10044), .IN2(n10045), .IN3(n9515), .Q(WX9080) );
  OR2X1 U9886 ( .IN1(DFF_1340_n1), .IN2(WX8599), .Q(n10045) );
  OR2X1 U9887 ( .IN1(n8796), .IN2(CRC_OUT_3_28), .Q(n10044) );
  AND3X1 U9888 ( .IN1(n10046), .IN2(n10047), .IN3(n9514), .Q(WX9078) );
  OR2X1 U9889 ( .IN1(DFF_1339_n1), .IN2(WX8601), .Q(n10047) );
  OR2X1 U9890 ( .IN1(n8797), .IN2(CRC_OUT_3_27), .Q(n10046) );
  AND3X1 U9891 ( .IN1(n10048), .IN2(n10049), .IN3(n9514), .Q(WX9076) );
  OR2X1 U9892 ( .IN1(DFF_1338_n1), .IN2(WX8603), .Q(n10049) );
  OR2X1 U9893 ( .IN1(n8798), .IN2(CRC_OUT_3_26), .Q(n10048) );
  AND2X1 U9894 ( .IN1(n10050), .IN2(n9496), .Q(WX9074) );
  OR2X1 U9895 ( .IN1(n10051), .IN2(n10052), .Q(n10050) );
  AND2X1 U9896 ( .IN1(DFF_1337_n1), .IN2(n9104), .Q(n10052) );
  AND2X1 U9897 ( .IN1(test_so74), .IN2(CRC_OUT_3_25), .Q(n10051) );
  AND2X1 U9898 ( .IN1(n10053), .IN2(n9496), .Q(WX9072) );
  OR2X1 U9899 ( .IN1(n10054), .IN2(n10055), .Q(n10053) );
  AND2X1 U9900 ( .IN1(n8799), .IN2(n9150), .Q(n10055) );
  AND2X1 U9901 ( .IN1(test_so77), .IN2(WX8607), .Q(n10054) );
  AND3X1 U9902 ( .IN1(n10056), .IN2(n10057), .IN3(n9514), .Q(WX9070) );
  OR2X1 U9903 ( .IN1(DFF_1335_n1), .IN2(WX8609), .Q(n10057) );
  OR2X1 U9904 ( .IN1(n8800), .IN2(CRC_OUT_3_23), .Q(n10056) );
  AND3X1 U9905 ( .IN1(n10058), .IN2(n10059), .IN3(n9513), .Q(WX9068) );
  OR2X1 U9906 ( .IN1(DFF_1334_n1), .IN2(WX8611), .Q(n10059) );
  OR2X1 U9907 ( .IN1(n8801), .IN2(CRC_OUT_3_22), .Q(n10058) );
  AND3X1 U9908 ( .IN1(n10060), .IN2(n10061), .IN3(n9514), .Q(WX9066) );
  OR2X1 U9909 ( .IN1(DFF_1333_n1), .IN2(WX8613), .Q(n10061) );
  OR2X1 U9910 ( .IN1(n8802), .IN2(CRC_OUT_3_21), .Q(n10060) );
  AND3X1 U9911 ( .IN1(n10062), .IN2(n10063), .IN3(n9513), .Q(WX9064) );
  OR2X1 U9912 ( .IN1(DFF_1332_n1), .IN2(WX8615), .Q(n10063) );
  OR2X1 U9913 ( .IN1(n8803), .IN2(CRC_OUT_3_20), .Q(n10062) );
  AND3X1 U9914 ( .IN1(n10064), .IN2(n10065), .IN3(n9514), .Q(WX9062) );
  OR2X1 U9915 ( .IN1(DFF_1331_n1), .IN2(WX8617), .Q(n10065) );
  OR2X1 U9916 ( .IN1(n8804), .IN2(CRC_OUT_3_19), .Q(n10064) );
  AND3X1 U9917 ( .IN1(n10066), .IN2(n10067), .IN3(n9515), .Q(WX9060) );
  OR2X1 U9918 ( .IN1(DFF_1330_n1), .IN2(WX8619), .Q(n10067) );
  OR2X1 U9919 ( .IN1(n8805), .IN2(CRC_OUT_3_18), .Q(n10066) );
  AND3X1 U9920 ( .IN1(n10068), .IN2(n10069), .IN3(n9515), .Q(WX9058) );
  OR2X1 U9921 ( .IN1(DFF_1329_n1), .IN2(WX8621), .Q(n10069) );
  OR2X1 U9922 ( .IN1(n8806), .IN2(CRC_OUT_3_17), .Q(n10068) );
  AND3X1 U9923 ( .IN1(n10070), .IN2(n10071), .IN3(n9516), .Q(WX9056) );
  OR2X1 U9924 ( .IN1(DFF_1328_n1), .IN2(WX8623), .Q(n10071) );
  OR2X1 U9925 ( .IN1(n8807), .IN2(CRC_OUT_3_16), .Q(n10070) );
  AND2X1 U9926 ( .IN1(n10072), .IN2(n9494), .Q(WX9054) );
  OR2X1 U9927 ( .IN1(n10073), .IN2(n10074), .Q(n10072) );
  AND2X1 U9928 ( .IN1(n10075), .IN2(CRC_OUT_3_15), .Q(n10074) );
  AND2X1 U9929 ( .IN1(DFF_1327_n1), .IN2(n10076), .Q(n10073) );
  INVX0 U9930 ( .INP(n10075), .ZN(n10076) );
  OR2X1 U9931 ( .IN1(n10077), .IN2(n10078), .Q(n10075) );
  AND2X1 U9932 ( .IN1(DFF_1343_n1), .IN2(WX8625), .Q(n10078) );
  AND2X1 U9933 ( .IN1(n8719), .IN2(CRC_OUT_3_31), .Q(n10077) );
  AND3X1 U9934 ( .IN1(n10079), .IN2(n10080), .IN3(n9515), .Q(WX9052) );
  OR2X1 U9935 ( .IN1(DFF_1326_n1), .IN2(WX8627), .Q(n10080) );
  OR2X1 U9936 ( .IN1(n8808), .IN2(CRC_OUT_3_14), .Q(n10079) );
  AND3X1 U9937 ( .IN1(n10081), .IN2(n10082), .IN3(n9517), .Q(WX9050) );
  OR2X1 U9938 ( .IN1(DFF_1325_n1), .IN2(WX8629), .Q(n10082) );
  OR2X1 U9939 ( .IN1(n8809), .IN2(CRC_OUT_3_13), .Q(n10081) );
  AND3X1 U9940 ( .IN1(n10083), .IN2(n10084), .IN3(n9516), .Q(WX9048) );
  OR2X1 U9941 ( .IN1(DFF_1324_n1), .IN2(WX8631), .Q(n10084) );
  OR2X1 U9942 ( .IN1(n8810), .IN2(CRC_OUT_3_12), .Q(n10083) );
  AND3X1 U9943 ( .IN1(n10085), .IN2(n10086), .IN3(n9516), .Q(WX9046) );
  OR2X1 U9944 ( .IN1(DFF_1323_n1), .IN2(WX8633), .Q(n10086) );
  OR2X1 U9945 ( .IN1(n8811), .IN2(CRC_OUT_3_11), .Q(n10085) );
  AND2X1 U9946 ( .IN1(n10087), .IN2(n9493), .Q(WX9044) );
  OR2X1 U9947 ( .IN1(n10088), .IN2(n10089), .Q(n10087) );
  AND2X1 U9948 ( .IN1(n10090), .IN2(CRC_OUT_3_10), .Q(n10089) );
  AND2X1 U9949 ( .IN1(DFF_1322_n1), .IN2(n10091), .Q(n10088) );
  INVX0 U9950 ( .INP(n10090), .ZN(n10091) );
  OR2X1 U9951 ( .IN1(n10092), .IN2(n10093), .Q(n10090) );
  AND2X1 U9952 ( .IN1(DFF_1343_n1), .IN2(WX8635), .Q(n10093) );
  AND2X1 U9953 ( .IN1(n8720), .IN2(CRC_OUT_3_31), .Q(n10092) );
  AND3X1 U9954 ( .IN1(n10094), .IN2(n10095), .IN3(n9517), .Q(WX9042) );
  OR2X1 U9955 ( .IN1(DFF_1321_n1), .IN2(WX8637), .Q(n10095) );
  OR2X1 U9956 ( .IN1(n8812), .IN2(CRC_OUT_3_9), .Q(n10094) );
  AND2X1 U9957 ( .IN1(n10096), .IN2(n9493), .Q(WX9040) );
  OR2X1 U9958 ( .IN1(n10097), .IN2(n10098), .Q(n10096) );
  AND2X1 U9959 ( .IN1(DFF_1320_n1), .IN2(n9099), .Q(n10098) );
  AND2X1 U9960 ( .IN1(test_so75), .IN2(CRC_OUT_3_8), .Q(n10097) );
  AND2X1 U9961 ( .IN1(n10099), .IN2(n9493), .Q(WX9038) );
  OR2X1 U9962 ( .IN1(n10100), .IN2(n10101), .Q(n10099) );
  AND2X1 U9963 ( .IN1(n8813), .IN2(n9151), .Q(n10101) );
  AND2X1 U9964 ( .IN1(test_so76), .IN2(WX8641), .Q(n10100) );
  AND3X1 U9965 ( .IN1(n10102), .IN2(n10103), .IN3(n9516), .Q(WX9036) );
  OR2X1 U9966 ( .IN1(DFF_1318_n1), .IN2(WX8643), .Q(n10103) );
  OR2X1 U9967 ( .IN1(n8814), .IN2(CRC_OUT_3_6), .Q(n10102) );
  AND3X1 U9968 ( .IN1(n10104), .IN2(n10105), .IN3(n9517), .Q(WX9034) );
  OR2X1 U9969 ( .IN1(DFF_1317_n1), .IN2(WX8645), .Q(n10105) );
  OR2X1 U9970 ( .IN1(n8815), .IN2(CRC_OUT_3_5), .Q(n10104) );
  AND3X1 U9971 ( .IN1(n10106), .IN2(n10107), .IN3(n9516), .Q(WX9032) );
  OR2X1 U9972 ( .IN1(DFF_1316_n1), .IN2(WX8647), .Q(n10107) );
  OR2X1 U9973 ( .IN1(n8816), .IN2(CRC_OUT_3_4), .Q(n10106) );
  AND2X1 U9974 ( .IN1(n10108), .IN2(n9493), .Q(WX9030) );
  OR2X1 U9975 ( .IN1(n10109), .IN2(n10110), .Q(n10108) );
  AND2X1 U9976 ( .IN1(n10111), .IN2(CRC_OUT_3_3), .Q(n10110) );
  AND2X1 U9977 ( .IN1(DFF_1315_n1), .IN2(n10112), .Q(n10109) );
  INVX0 U9978 ( .INP(n10111), .ZN(n10112) );
  OR2X1 U9979 ( .IN1(n10113), .IN2(n10114), .Q(n10111) );
  AND2X1 U9980 ( .IN1(DFF_1343_n1), .IN2(WX8649), .Q(n10114) );
  AND2X1 U9981 ( .IN1(n8721), .IN2(CRC_OUT_3_31), .Q(n10113) );
  AND3X1 U9982 ( .IN1(n10115), .IN2(n10116), .IN3(n9517), .Q(WX9028) );
  OR2X1 U9983 ( .IN1(DFF_1314_n1), .IN2(WX8651), .Q(n10116) );
  OR2X1 U9984 ( .IN1(n8817), .IN2(CRC_OUT_3_2), .Q(n10115) );
  AND3X1 U9985 ( .IN1(n10117), .IN2(n10118), .IN3(n9517), .Q(WX9026) );
  OR2X1 U9986 ( .IN1(DFF_1313_n1), .IN2(WX8653), .Q(n10118) );
  OR2X1 U9987 ( .IN1(n8818), .IN2(CRC_OUT_3_1), .Q(n10117) );
  AND3X1 U9988 ( .IN1(n10119), .IN2(n10120), .IN3(n9517), .Q(WX9024) );
  OR2X1 U9989 ( .IN1(DFF_1312_n1), .IN2(WX8655), .Q(n10120) );
  OR2X1 U9990 ( .IN1(n8819), .IN2(CRC_OUT_3_0), .Q(n10119) );
  AND3X1 U9991 ( .IN1(n10121), .IN2(n10122), .IN3(n9517), .Q(WX9022) );
  OR2X1 U9992 ( .IN1(DFF_1343_n1), .IN2(WX8657), .Q(n10122) );
  OR2X1 U9993 ( .IN1(n8736), .IN2(CRC_OUT_3_31), .Q(n10121) );
  AND2X1 U9994 ( .IN1(n9512), .IN2(n8363), .Q(WX8496) );
  AND2X1 U9995 ( .IN1(n9512), .IN2(n8364), .Q(WX8494) );
  AND2X1 U9996 ( .IN1(n9512), .IN2(n8365), .Q(WX8492) );
  AND2X1 U9997 ( .IN1(n9511), .IN2(n8366), .Q(WX8490) );
  AND2X1 U9998 ( .IN1(n9507), .IN2(n8367), .Q(WX8488) );
  AND2X1 U9999 ( .IN1(n9507), .IN2(n8368), .Q(WX8486) );
  AND2X1 U10000 ( .IN1(n9504), .IN2(n8369), .Q(WX8484) );
  AND2X1 U10001 ( .IN1(n9505), .IN2(n8370), .Q(WX8482) );
  AND2X1 U10002 ( .IN1(n9505), .IN2(n8371), .Q(WX8480) );
  AND2X1 U10003 ( .IN1(n9504), .IN2(n8372), .Q(WX8478) );
  AND2X1 U10004 ( .IN1(n9503), .IN2(n8373), .Q(WX8476) );
  AND2X1 U10005 ( .IN1(n9505), .IN2(n8374), .Q(WX8474) );
  AND2X1 U10006 ( .IN1(n9504), .IN2(n8375), .Q(WX8472) );
  AND2X1 U10007 ( .IN1(n9504), .IN2(n8376), .Q(WX8470) );
  AND2X1 U10008 ( .IN1(n9503), .IN2(n8377), .Q(WX8468) );
  AND2X1 U10009 ( .IN1(n9503), .IN2(n8378), .Q(WX8466) );
  OR4X1 U10010 ( .IN1(n10123), .IN2(n10124), .IN3(n10125), .IN4(n10126), .Q(
        WX8464) );
  AND2X1 U10011 ( .IN1(n9183), .IN2(n10127), .Q(n10126) );
  AND2X1 U10012 ( .IN1(n9271), .IN2(n9822), .Q(n10125) );
  OR2X1 U10013 ( .IN1(n10128), .IN2(n10129), .Q(n9822) );
  INVX0 U10014 ( .INP(n10130), .ZN(n10129) );
  OR2X1 U10015 ( .IN1(n10131), .IN2(n10132), .Q(n10130) );
  AND2X1 U10016 ( .IN1(n10132), .IN2(n10131), .Q(n10128) );
  AND2X1 U10017 ( .IN1(n10133), .IN2(n10134), .Q(n10131) );
  OR2X1 U10018 ( .IN1(WX9822), .IN2(n8148), .Q(n10134) );
  INVX0 U10019 ( .INP(n10135), .ZN(n10133) );
  AND2X1 U10020 ( .IN1(n8148), .IN2(WX9822), .Q(n10135) );
  OR2X1 U10021 ( .IN1(n10136), .IN2(n10137), .Q(n10132) );
  AND2X1 U10022 ( .IN1(n8149), .IN2(WX9950), .Q(n10137) );
  AND2X1 U10023 ( .IN1(n8735), .IN2(WX9886), .Q(n10136) );
  AND2X1 U10024 ( .IN1(n9240), .IN2(CRC_OUT_3_0), .Q(n10124) );
  AND2X1 U10025 ( .IN1(n1502), .IN2(n9215), .Q(n10123) );
  INVX0 U10026 ( .INP(n10138), .ZN(n1502) );
  OR2X1 U10027 ( .IN1(n9575), .IN2(n3848), .Q(n10138) );
  OR4X1 U10028 ( .IN1(n10139), .IN2(n10140), .IN3(n10141), .IN4(n10142), .Q(
        WX8462) );
  AND2X1 U10029 ( .IN1(n9183), .IN2(n10143), .Q(n10142) );
  AND2X1 U10030 ( .IN1(n9829), .IN2(n9262), .Q(n10141) );
  AND2X1 U10031 ( .IN1(n10144), .IN2(n10145), .Q(n9829) );
  INVX0 U10032 ( .INP(n10146), .ZN(n10145) );
  AND2X1 U10033 ( .IN1(n10147), .IN2(n10148), .Q(n10146) );
  OR2X1 U10034 ( .IN1(n10148), .IN2(n10147), .Q(n10144) );
  OR2X1 U10035 ( .IN1(n10149), .IN2(n10150), .Q(n10147) );
  INVX0 U10036 ( .INP(n10151), .ZN(n10150) );
  OR2X1 U10037 ( .IN1(WX9756), .IN2(n8151), .Q(n10151) );
  AND2X1 U10038 ( .IN1(n8151), .IN2(WX9756), .Q(n10149) );
  AND2X1 U10039 ( .IN1(n10152), .IN2(n10153), .Q(n10148) );
  OR2X1 U10040 ( .IN1(WX9948), .IN2(test_so83), .Q(n10153) );
  OR2X1 U10041 ( .IN1(n9111), .IN2(n8793), .Q(n10152) );
  AND2X1 U10042 ( .IN1(n9240), .IN2(CRC_OUT_3_1), .Q(n10140) );
  AND2X1 U10043 ( .IN1(n1501), .IN2(n9215), .Q(n10139) );
  INVX0 U10044 ( .INP(n10154), .ZN(n1501) );
  OR2X1 U10045 ( .IN1(n9574), .IN2(n3849), .Q(n10154) );
  OR4X1 U10046 ( .IN1(n10155), .IN2(n10156), .IN3(n10157), .IN4(n10158), .Q(
        WX8460) );
  AND2X1 U10047 ( .IN1(n9183), .IN2(n10159), .Q(n10158) );
  AND2X1 U10048 ( .IN1(n9271), .IN2(n9836), .Q(n10157) );
  OR2X1 U10049 ( .IN1(n10160), .IN2(n10161), .Q(n9836) );
  INVX0 U10050 ( .INP(n10162), .ZN(n10161) );
  OR2X1 U10051 ( .IN1(n10163), .IN2(n10164), .Q(n10162) );
  AND2X1 U10052 ( .IN1(n10164), .IN2(n10163), .Q(n10160) );
  AND2X1 U10053 ( .IN1(n10165), .IN2(n10166), .Q(n10163) );
  OR2X1 U10054 ( .IN1(WX9818), .IN2(n8152), .Q(n10166) );
  INVX0 U10055 ( .INP(n10167), .ZN(n10165) );
  AND2X1 U10056 ( .IN1(n8152), .IN2(WX9818), .Q(n10167) );
  OR2X1 U10057 ( .IN1(n10168), .IN2(n10169), .Q(n10164) );
  AND2X1 U10058 ( .IN1(n8153), .IN2(WX9946), .Q(n10169) );
  AND2X1 U10059 ( .IN1(n8792), .IN2(WX9882), .Q(n10168) );
  AND2X1 U10060 ( .IN1(n9240), .IN2(CRC_OUT_3_2), .Q(n10156) );
  AND2X1 U10061 ( .IN1(n1500), .IN2(n9218), .Q(n10155) );
  INVX0 U10062 ( .INP(n10170), .ZN(n1500) );
  OR2X1 U10063 ( .IN1(n9574), .IN2(n3850), .Q(n10170) );
  OR4X1 U10064 ( .IN1(n10171), .IN2(n10172), .IN3(n10173), .IN4(n10174), .Q(
        WX8458) );
  AND2X1 U10065 ( .IN1(n9183), .IN2(n10175), .Q(n10174) );
  AND2X1 U10066 ( .IN1(n9843), .IN2(n9261), .Q(n10173) );
  AND2X1 U10067 ( .IN1(n10176), .IN2(n10177), .Q(n9843) );
  INVX0 U10068 ( .INP(n10178), .ZN(n10177) );
  AND2X1 U10069 ( .IN1(n10179), .IN2(n10180), .Q(n10178) );
  OR2X1 U10070 ( .IN1(n10180), .IN2(n10179), .Q(n10176) );
  OR2X1 U10071 ( .IN1(n10181), .IN2(n10182), .Q(n10179) );
  INVX0 U10072 ( .INP(n10183), .ZN(n10182) );
  OR2X1 U10073 ( .IN1(WX9816), .IN2(n8154), .Q(n10183) );
  AND2X1 U10074 ( .IN1(n8154), .IN2(WX9816), .Q(n10181) );
  AND2X1 U10075 ( .IN1(n10184), .IN2(n10185), .Q(n10180) );
  OR2X1 U10076 ( .IN1(WX9944), .IN2(test_so81), .Q(n10185) );
  OR2X1 U10077 ( .IN1(n9112), .IN2(n8791), .Q(n10184) );
  AND2X1 U10078 ( .IN1(n9241), .IN2(CRC_OUT_3_3), .Q(n10172) );
  AND2X1 U10079 ( .IN1(n1499), .IN2(n9215), .Q(n10171) );
  INVX0 U10080 ( .INP(n10186), .ZN(n1499) );
  OR2X1 U10081 ( .IN1(n9574), .IN2(n3851), .Q(n10186) );
  OR4X1 U10082 ( .IN1(n10187), .IN2(n10188), .IN3(n10189), .IN4(n10190), .Q(
        WX8456) );
  AND2X1 U10083 ( .IN1(n9183), .IN2(n10191), .Q(n10190) );
  AND2X1 U10084 ( .IN1(n9272), .IN2(n9850), .Q(n10189) );
  OR2X1 U10085 ( .IN1(n10192), .IN2(n10193), .Q(n9850) );
  INVX0 U10086 ( .INP(n10194), .ZN(n10193) );
  OR2X1 U10087 ( .IN1(n10195), .IN2(n10196), .Q(n10194) );
  AND2X1 U10088 ( .IN1(n10196), .IN2(n10195), .Q(n10192) );
  AND2X1 U10089 ( .IN1(n10197), .IN2(n10198), .Q(n10195) );
  OR2X1 U10090 ( .IN1(WX9814), .IN2(n8155), .Q(n10198) );
  INVX0 U10091 ( .INP(n10199), .ZN(n10197) );
  AND2X1 U10092 ( .IN1(n8155), .IN2(WX9814), .Q(n10199) );
  OR2X1 U10093 ( .IN1(n10200), .IN2(n10201), .Q(n10196) );
  AND2X1 U10094 ( .IN1(n8156), .IN2(WX9942), .Q(n10201) );
  AND2X1 U10095 ( .IN1(n8718), .IN2(WX9878), .Q(n10200) );
  AND2X1 U10096 ( .IN1(n9241), .IN2(CRC_OUT_3_4), .Q(n10188) );
  AND2X1 U10097 ( .IN1(n1498), .IN2(n9215), .Q(n10187) );
  INVX0 U10098 ( .INP(n10202), .ZN(n1498) );
  OR2X1 U10099 ( .IN1(n9574), .IN2(n3852), .Q(n10202) );
  OR4X1 U10100 ( .IN1(n10203), .IN2(n10204), .IN3(n10205), .IN4(n10206), .Q(
        WX8454) );
  AND2X1 U10101 ( .IN1(n9183), .IN2(n10207), .Q(n10206) );
  AND2X1 U10102 ( .IN1(n9272), .IN2(n9857), .Q(n10205) );
  OR2X1 U10103 ( .IN1(n10208), .IN2(n10209), .Q(n9857) );
  INVX0 U10104 ( .INP(n10210), .ZN(n10209) );
  OR2X1 U10105 ( .IN1(n10211), .IN2(n10212), .Q(n10210) );
  AND2X1 U10106 ( .IN1(n10212), .IN2(n10211), .Q(n10208) );
  AND2X1 U10107 ( .IN1(n10213), .IN2(n10214), .Q(n10211) );
  OR2X1 U10108 ( .IN1(WX9812), .IN2(n8157), .Q(n10214) );
  INVX0 U10109 ( .INP(n10215), .ZN(n10213) );
  AND2X1 U10110 ( .IN1(n8157), .IN2(WX9812), .Q(n10215) );
  OR2X1 U10111 ( .IN1(n10216), .IN2(n10217), .Q(n10212) );
  AND2X1 U10112 ( .IN1(n8158), .IN2(WX9940), .Q(n10217) );
  AND2X1 U10113 ( .IN1(n8790), .IN2(WX9876), .Q(n10216) );
  AND2X1 U10114 ( .IN1(n9241), .IN2(CRC_OUT_3_5), .Q(n10204) );
  AND2X1 U10115 ( .IN1(n1497), .IN2(n9215), .Q(n10203) );
  INVX0 U10116 ( .INP(n10218), .ZN(n1497) );
  OR2X1 U10117 ( .IN1(n9574), .IN2(n3853), .Q(n10218) );
  OR4X1 U10118 ( .IN1(n10219), .IN2(n10220), .IN3(n10221), .IN4(n10222), .Q(
        WX8452) );
  AND2X1 U10119 ( .IN1(n9183), .IN2(n10223), .Q(n10222) );
  AND2X1 U10120 ( .IN1(n9272), .IN2(n9864), .Q(n10221) );
  OR2X1 U10121 ( .IN1(n10224), .IN2(n10225), .Q(n9864) );
  INVX0 U10122 ( .INP(n10226), .ZN(n10225) );
  OR2X1 U10123 ( .IN1(n10227), .IN2(n10228), .Q(n10226) );
  AND2X1 U10124 ( .IN1(n10228), .IN2(n10227), .Q(n10224) );
  AND2X1 U10125 ( .IN1(n10229), .IN2(n10230), .Q(n10227) );
  OR2X1 U10126 ( .IN1(WX9810), .IN2(n8159), .Q(n10230) );
  INVX0 U10127 ( .INP(n10231), .ZN(n10229) );
  AND2X1 U10128 ( .IN1(n8159), .IN2(WX9810), .Q(n10231) );
  OR2X1 U10129 ( .IN1(n10232), .IN2(n10233), .Q(n10228) );
  AND2X1 U10130 ( .IN1(n8160), .IN2(WX9938), .Q(n10233) );
  AND2X1 U10131 ( .IN1(n8789), .IN2(WX9874), .Q(n10232) );
  AND2X1 U10132 ( .IN1(n9241), .IN2(CRC_OUT_3_6), .Q(n10220) );
  AND2X1 U10133 ( .IN1(n1496), .IN2(n9215), .Q(n10219) );
  INVX0 U10134 ( .INP(n10234), .ZN(n1496) );
  OR2X1 U10135 ( .IN1(n9574), .IN2(n3854), .Q(n10234) );
  OR4X1 U10136 ( .IN1(n10235), .IN2(n10236), .IN3(n10237), .IN4(n10238), .Q(
        WX8450) );
  AND2X1 U10137 ( .IN1(n9183), .IN2(n10239), .Q(n10238) );
  AND2X1 U10138 ( .IN1(n9272), .IN2(n9871), .Q(n10237) );
  OR2X1 U10139 ( .IN1(n10240), .IN2(n10241), .Q(n9871) );
  INVX0 U10140 ( .INP(n10242), .ZN(n10241) );
  OR2X1 U10141 ( .IN1(n10243), .IN2(n10244), .Q(n10242) );
  AND2X1 U10142 ( .IN1(n10244), .IN2(n10243), .Q(n10240) );
  AND2X1 U10143 ( .IN1(n10245), .IN2(n10246), .Q(n10243) );
  OR2X1 U10144 ( .IN1(WX9808), .IN2(n8161), .Q(n10246) );
  INVX0 U10145 ( .INP(n10247), .ZN(n10245) );
  AND2X1 U10146 ( .IN1(n8161), .IN2(WX9808), .Q(n10247) );
  OR2X1 U10147 ( .IN1(n10248), .IN2(n10249), .Q(n10244) );
  AND2X1 U10148 ( .IN1(n8162), .IN2(WX9936), .Q(n10249) );
  AND2X1 U10149 ( .IN1(n8788), .IN2(WX9872), .Q(n10248) );
  AND2X1 U10150 ( .IN1(test_so76), .IN2(n9228), .Q(n10236) );
  AND2X1 U10151 ( .IN1(n1495), .IN2(n9215), .Q(n10235) );
  INVX0 U10152 ( .INP(n10250), .ZN(n1495) );
  OR2X1 U10153 ( .IN1(n9574), .IN2(n3855), .Q(n10250) );
  OR4X1 U10154 ( .IN1(n10251), .IN2(n10252), .IN3(n10253), .IN4(n10254), .Q(
        WX8448) );
  AND2X1 U10155 ( .IN1(n9183), .IN2(n10255), .Q(n10254) );
  AND2X1 U10156 ( .IN1(n9272), .IN2(n9878), .Q(n10253) );
  OR2X1 U10157 ( .IN1(n10256), .IN2(n10257), .Q(n9878) );
  INVX0 U10158 ( .INP(n10258), .ZN(n10257) );
  OR2X1 U10159 ( .IN1(n10259), .IN2(n10260), .Q(n10258) );
  AND2X1 U10160 ( .IN1(n10260), .IN2(n10259), .Q(n10256) );
  AND2X1 U10161 ( .IN1(n10261), .IN2(n10262), .Q(n10259) );
  OR2X1 U10162 ( .IN1(WX9806), .IN2(n8163), .Q(n10262) );
  INVX0 U10163 ( .INP(n10263), .ZN(n10261) );
  AND2X1 U10164 ( .IN1(n8163), .IN2(WX9806), .Q(n10263) );
  OR2X1 U10165 ( .IN1(n10264), .IN2(n10265), .Q(n10260) );
  AND2X1 U10166 ( .IN1(n8164), .IN2(WX9934), .Q(n10265) );
  AND2X1 U10167 ( .IN1(n8787), .IN2(WX9870), .Q(n10264) );
  AND2X1 U10168 ( .IN1(n9241), .IN2(CRC_OUT_3_8), .Q(n10252) );
  AND2X1 U10169 ( .IN1(n1494), .IN2(n9215), .Q(n10251) );
  INVX0 U10170 ( .INP(n10266), .ZN(n1494) );
  OR2X1 U10171 ( .IN1(n9574), .IN2(n3856), .Q(n10266) );
  OR4X1 U10172 ( .IN1(n10267), .IN2(n10268), .IN3(n10269), .IN4(n10270), .Q(
        WX8446) );
  AND2X1 U10173 ( .IN1(n10271), .IN2(n9177), .Q(n10270) );
  AND2X1 U10174 ( .IN1(n9272), .IN2(n9885), .Q(n10269) );
  OR2X1 U10175 ( .IN1(n10272), .IN2(n10273), .Q(n9885) );
  INVX0 U10176 ( .INP(n10274), .ZN(n10273) );
  OR2X1 U10177 ( .IN1(n10275), .IN2(n10276), .Q(n10274) );
  AND2X1 U10178 ( .IN1(n10276), .IN2(n10275), .Q(n10272) );
  AND2X1 U10179 ( .IN1(n10277), .IN2(n10278), .Q(n10275) );
  OR2X1 U10180 ( .IN1(WX9804), .IN2(n8165), .Q(n10278) );
  INVX0 U10181 ( .INP(n10279), .ZN(n10277) );
  AND2X1 U10182 ( .IN1(n8165), .IN2(WX9804), .Q(n10279) );
  OR2X1 U10183 ( .IN1(n10280), .IN2(n10281), .Q(n10276) );
  AND2X1 U10184 ( .IN1(n8166), .IN2(WX9932), .Q(n10281) );
  AND2X1 U10185 ( .IN1(n8786), .IN2(WX9868), .Q(n10280) );
  AND2X1 U10186 ( .IN1(n9241), .IN2(CRC_OUT_3_9), .Q(n10268) );
  AND2X1 U10187 ( .IN1(n1493), .IN2(n9215), .Q(n10267) );
  INVX0 U10188 ( .INP(n10282), .ZN(n1493) );
  OR2X1 U10189 ( .IN1(n9574), .IN2(n3857), .Q(n10282) );
  OR4X1 U10190 ( .IN1(n10283), .IN2(n10284), .IN3(n10285), .IN4(n10286), .Q(
        WX8444) );
  AND2X1 U10191 ( .IN1(n9183), .IN2(n10287), .Q(n10286) );
  AND2X1 U10192 ( .IN1(n9272), .IN2(n9892), .Q(n10285) );
  OR2X1 U10193 ( .IN1(n10288), .IN2(n10289), .Q(n9892) );
  INVX0 U10194 ( .INP(n10290), .ZN(n10289) );
  OR2X1 U10195 ( .IN1(n10291), .IN2(n10292), .Q(n10290) );
  AND2X1 U10196 ( .IN1(n10292), .IN2(n10291), .Q(n10288) );
  AND2X1 U10197 ( .IN1(n10293), .IN2(n10294), .Q(n10291) );
  OR2X1 U10198 ( .IN1(WX9802), .IN2(n8167), .Q(n10294) );
  INVX0 U10199 ( .INP(n10295), .ZN(n10293) );
  AND2X1 U10200 ( .IN1(n8167), .IN2(WX9802), .Q(n10295) );
  OR2X1 U10201 ( .IN1(n10296), .IN2(n10297), .Q(n10292) );
  AND2X1 U10202 ( .IN1(n8168), .IN2(WX9930), .Q(n10297) );
  AND2X1 U10203 ( .IN1(n8785), .IN2(WX9866), .Q(n10296) );
  AND2X1 U10204 ( .IN1(n9241), .IN2(CRC_OUT_3_10), .Q(n10284) );
  AND2X1 U10205 ( .IN1(n1492), .IN2(n9215), .Q(n10283) );
  INVX0 U10206 ( .INP(n10298), .ZN(n1492) );
  OR2X1 U10207 ( .IN1(n9574), .IN2(n3858), .Q(n10298) );
  OR4X1 U10208 ( .IN1(n10299), .IN2(n10300), .IN3(n10301), .IN4(n10302), .Q(
        WX8442) );
  AND2X1 U10209 ( .IN1(n10303), .IN2(n9177), .Q(n10302) );
  AND2X1 U10210 ( .IN1(n9272), .IN2(n9899), .Q(n10301) );
  OR2X1 U10211 ( .IN1(n10304), .IN2(n10305), .Q(n9899) );
  INVX0 U10212 ( .INP(n10306), .ZN(n10305) );
  OR2X1 U10213 ( .IN1(n10307), .IN2(n10308), .Q(n10306) );
  AND2X1 U10214 ( .IN1(n10308), .IN2(n10307), .Q(n10304) );
  AND2X1 U10215 ( .IN1(n10309), .IN2(n10310), .Q(n10307) );
  OR2X1 U10216 ( .IN1(WX9800), .IN2(n8169), .Q(n10310) );
  INVX0 U10217 ( .INP(n10311), .ZN(n10309) );
  AND2X1 U10218 ( .IN1(n8169), .IN2(WX9800), .Q(n10311) );
  OR2X1 U10219 ( .IN1(n10312), .IN2(n10313), .Q(n10308) );
  AND2X1 U10220 ( .IN1(n8170), .IN2(WX9928), .Q(n10313) );
  AND2X1 U10221 ( .IN1(n8717), .IN2(WX9864), .Q(n10312) );
  AND2X1 U10222 ( .IN1(n9241), .IN2(CRC_OUT_3_11), .Q(n10300) );
  AND2X1 U10223 ( .IN1(n1491), .IN2(n9216), .Q(n10299) );
  INVX0 U10224 ( .INP(n10314), .ZN(n1491) );
  OR2X1 U10225 ( .IN1(n9574), .IN2(n3859), .Q(n10314) );
  OR4X1 U10226 ( .IN1(n10315), .IN2(n10316), .IN3(n10317), .IN4(n10318), .Q(
        WX8440) );
  AND2X1 U10227 ( .IN1(n9183), .IN2(n10319), .Q(n10318) );
  AND2X1 U10228 ( .IN1(n9272), .IN2(n9906), .Q(n10317) );
  OR2X1 U10229 ( .IN1(n10320), .IN2(n10321), .Q(n9906) );
  INVX0 U10230 ( .INP(n10322), .ZN(n10321) );
  OR2X1 U10231 ( .IN1(n10323), .IN2(n10324), .Q(n10322) );
  AND2X1 U10232 ( .IN1(n10324), .IN2(n10323), .Q(n10320) );
  AND2X1 U10233 ( .IN1(n10325), .IN2(n10326), .Q(n10323) );
  OR2X1 U10234 ( .IN1(WX9798), .IN2(n8171), .Q(n10326) );
  INVX0 U10235 ( .INP(n10327), .ZN(n10325) );
  AND2X1 U10236 ( .IN1(n8171), .IN2(WX9798), .Q(n10327) );
  OR2X1 U10237 ( .IN1(n10328), .IN2(n10329), .Q(n10324) );
  AND2X1 U10238 ( .IN1(n8172), .IN2(WX9926), .Q(n10329) );
  AND2X1 U10239 ( .IN1(n8784), .IN2(WX9862), .Q(n10328) );
  AND2X1 U10240 ( .IN1(n9241), .IN2(CRC_OUT_3_12), .Q(n10316) );
  AND2X1 U10241 ( .IN1(n1490), .IN2(n9216), .Q(n10315) );
  INVX0 U10242 ( .INP(n10330), .ZN(n1490) );
  OR2X1 U10243 ( .IN1(n9574), .IN2(n3860), .Q(n10330) );
  OR4X1 U10244 ( .IN1(n10331), .IN2(n10332), .IN3(n10333), .IN4(n10334), .Q(
        WX8438) );
  AND2X1 U10245 ( .IN1(n10335), .IN2(n9177), .Q(n10334) );
  AND2X1 U10246 ( .IN1(n9272), .IN2(n9913), .Q(n10333) );
  OR2X1 U10247 ( .IN1(n10336), .IN2(n10337), .Q(n9913) );
  INVX0 U10248 ( .INP(n10338), .ZN(n10337) );
  OR2X1 U10249 ( .IN1(n10339), .IN2(n10340), .Q(n10338) );
  AND2X1 U10250 ( .IN1(n10340), .IN2(n10339), .Q(n10336) );
  AND2X1 U10251 ( .IN1(n10341), .IN2(n10342), .Q(n10339) );
  OR2X1 U10252 ( .IN1(WX9796), .IN2(n8173), .Q(n10342) );
  INVX0 U10253 ( .INP(n10343), .ZN(n10341) );
  AND2X1 U10254 ( .IN1(n8173), .IN2(WX9796), .Q(n10343) );
  OR2X1 U10255 ( .IN1(n10344), .IN2(n10345), .Q(n10340) );
  AND2X1 U10256 ( .IN1(n8174), .IN2(WX9924), .Q(n10345) );
  AND2X1 U10257 ( .IN1(n8783), .IN2(WX9860), .Q(n10344) );
  AND2X1 U10258 ( .IN1(n9241), .IN2(CRC_OUT_3_13), .Q(n10332) );
  AND2X1 U10259 ( .IN1(n1489), .IN2(n9216), .Q(n10331) );
  INVX0 U10260 ( .INP(n10346), .ZN(n1489) );
  OR2X1 U10261 ( .IN1(n9573), .IN2(n3861), .Q(n10346) );
  OR4X1 U10262 ( .IN1(n10347), .IN2(n10348), .IN3(n10349), .IN4(n10350), .Q(
        WX8436) );
  AND2X1 U10263 ( .IN1(n9183), .IN2(n10351), .Q(n10350) );
  AND2X1 U10264 ( .IN1(n9920), .IN2(n9261), .Q(n10349) );
  AND2X1 U10265 ( .IN1(n10352), .IN2(n10353), .Q(n9920) );
  INVX0 U10266 ( .INP(n10354), .ZN(n10353) );
  AND2X1 U10267 ( .IN1(n10355), .IN2(n10356), .Q(n10354) );
  OR2X1 U10268 ( .IN1(n10356), .IN2(n10355), .Q(n10352) );
  OR2X1 U10269 ( .IN1(n10357), .IN2(n10358), .Q(n10355) );
  INVX0 U10270 ( .INP(n10359), .ZN(n10358) );
  OR2X1 U10271 ( .IN1(WX9794), .IN2(n8175), .Q(n10359) );
  AND2X1 U10272 ( .IN1(n8175), .IN2(WX9794), .Q(n10357) );
  AND2X1 U10273 ( .IN1(n10360), .IN2(n10361), .Q(n10356) );
  OR2X1 U10274 ( .IN1(WX9858), .IN2(test_so86), .Q(n10361) );
  OR2X1 U10275 ( .IN1(n9103), .IN2(n8176), .Q(n10360) );
  AND2X1 U10276 ( .IN1(n9241), .IN2(CRC_OUT_3_14), .Q(n10348) );
  AND2X1 U10277 ( .IN1(n1488), .IN2(n9216), .Q(n10347) );
  INVX0 U10278 ( .INP(n10362), .ZN(n1488) );
  OR2X1 U10279 ( .IN1(n9573), .IN2(n3862), .Q(n10362) );
  OR4X1 U10280 ( .IN1(n10363), .IN2(n10364), .IN3(n10365), .IN4(n10366), .Q(
        WX8434) );
  AND2X1 U10281 ( .IN1(n10367), .IN2(n9176), .Q(n10366) );
  AND2X1 U10282 ( .IN1(n9272), .IN2(n9927), .Q(n10365) );
  OR2X1 U10283 ( .IN1(n10368), .IN2(n10369), .Q(n9927) );
  INVX0 U10284 ( .INP(n10370), .ZN(n10369) );
  OR2X1 U10285 ( .IN1(n10371), .IN2(n10372), .Q(n10370) );
  AND2X1 U10286 ( .IN1(n10372), .IN2(n10371), .Q(n10368) );
  AND2X1 U10287 ( .IN1(n10373), .IN2(n10374), .Q(n10371) );
  OR2X1 U10288 ( .IN1(WX9792), .IN2(n8177), .Q(n10374) );
  INVX0 U10289 ( .INP(n10375), .ZN(n10373) );
  AND2X1 U10290 ( .IN1(n8177), .IN2(WX9792), .Q(n10375) );
  OR2X1 U10291 ( .IN1(n10376), .IN2(n10377), .Q(n10372) );
  AND2X1 U10292 ( .IN1(n8178), .IN2(WX9920), .Q(n10377) );
  AND2X1 U10293 ( .IN1(n8782), .IN2(WX9856), .Q(n10376) );
  AND2X1 U10294 ( .IN1(n9241), .IN2(CRC_OUT_3_15), .Q(n10364) );
  AND2X1 U10295 ( .IN1(n1487), .IN2(n9216), .Q(n10363) );
  INVX0 U10296 ( .INP(n10378), .ZN(n1487) );
  OR2X1 U10297 ( .IN1(n9573), .IN2(n3863), .Q(n10378) );
  OR4X1 U10298 ( .IN1(n10379), .IN2(n10380), .IN3(n10381), .IN4(n10382), .Q(
        WX8432) );
  AND2X1 U10299 ( .IN1(n9183), .IN2(n10383), .Q(n10382) );
  AND2X1 U10300 ( .IN1(n9934), .IN2(n9260), .Q(n10381) );
  AND2X1 U10301 ( .IN1(n10384), .IN2(n10385), .Q(n9934) );
  INVX0 U10302 ( .INP(n10386), .ZN(n10385) );
  AND2X1 U10303 ( .IN1(n10387), .IN2(n10388), .Q(n10386) );
  OR2X1 U10304 ( .IN1(n10388), .IN2(n10387), .Q(n10384) );
  OR2X1 U10305 ( .IN1(n10389), .IN2(n10390), .Q(n10387) );
  AND2X1 U10306 ( .IN1(n9451), .IN2(WX9790), .Q(n10390) );
  AND2X1 U10307 ( .IN1(n7920), .IN2(n9475), .Q(n10389) );
  AND2X1 U10308 ( .IN1(n10391), .IN2(n10392), .Q(n10388) );
  OR2X1 U10309 ( .IN1(n10393), .IN2(n8716), .Q(n10392) );
  OR2X1 U10310 ( .IN1(WX9918), .IN2(n10394), .Q(n10391) );
  INVX0 U10311 ( .INP(n10393), .ZN(n10394) );
  AND2X1 U10312 ( .IN1(n10395), .IN2(n10396), .Q(n10393) );
  OR2X1 U10313 ( .IN1(n8304), .IN2(test_so84), .Q(n10396) );
  OR2X1 U10314 ( .IN1(n9113), .IN2(n15877), .Q(n10395) );
  AND2X1 U10315 ( .IN1(n9241), .IN2(CRC_OUT_3_16), .Q(n10380) );
  AND2X1 U10316 ( .IN1(n1486), .IN2(n9216), .Q(n10379) );
  INVX0 U10317 ( .INP(n10397), .ZN(n1486) );
  OR2X1 U10318 ( .IN1(n9573), .IN2(n3864), .Q(n10397) );
  OR4X1 U10319 ( .IN1(n10398), .IN2(n10399), .IN3(n10400), .IN4(n10401), .Q(
        WX8430) );
  AND2X1 U10320 ( .IN1(n9182), .IN2(n10402), .Q(n10401) );
  AND2X1 U10321 ( .IN1(n9272), .IN2(n9941), .Q(n10400) );
  OR2X1 U10322 ( .IN1(n10403), .IN2(n10404), .Q(n9941) );
  INVX0 U10323 ( .INP(n10405), .ZN(n10404) );
  OR2X1 U10324 ( .IN1(n10406), .IN2(n10407), .Q(n10405) );
  AND2X1 U10325 ( .IN1(n10407), .IN2(n10406), .Q(n10403) );
  AND2X1 U10326 ( .IN1(n10408), .IN2(n10409), .Q(n10406) );
  OR2X1 U10327 ( .IN1(n9452), .IN2(n7921), .Q(n10409) );
  OR2X1 U10328 ( .IN1(WX9788), .IN2(n9450), .Q(n10408) );
  OR2X1 U10329 ( .IN1(n10410), .IN2(n10411), .Q(n10407) );
  INVX0 U10330 ( .INP(n10412), .ZN(n10411) );
  OR2X1 U10331 ( .IN1(n10413), .IN2(n7922), .Q(n10412) );
  AND2X1 U10332 ( .IN1(n7922), .IN2(n10413), .Q(n10410) );
  INVX0 U10333 ( .INP(n10414), .ZN(n10413) );
  OR2X1 U10334 ( .IN1(n10415), .IN2(n10416), .Q(n10414) );
  AND2X1 U10335 ( .IN1(n8781), .IN2(n8305), .Q(n10416) );
  AND2X1 U10336 ( .IN1(n15878), .IN2(WX9916), .Q(n10415) );
  AND2X1 U10337 ( .IN1(n9242), .IN2(CRC_OUT_3_17), .Q(n10399) );
  AND2X1 U10338 ( .IN1(n1485), .IN2(n9216), .Q(n10398) );
  INVX0 U10339 ( .INP(n10417), .ZN(n1485) );
  OR2X1 U10340 ( .IN1(n9573), .IN2(n3865), .Q(n10417) );
  OR4X1 U10341 ( .IN1(n10418), .IN2(n10419), .IN3(n10420), .IN4(n10421), .Q(
        WX8428) );
  AND2X1 U10342 ( .IN1(n9182), .IN2(n10422), .Q(n10421) );
  AND2X1 U10343 ( .IN1(n9948), .IN2(n9260), .Q(n10420) );
  AND2X1 U10344 ( .IN1(n10423), .IN2(n10424), .Q(n9948) );
  INVX0 U10345 ( .INP(n10425), .ZN(n10424) );
  AND2X1 U10346 ( .IN1(n10426), .IN2(n10427), .Q(n10425) );
  OR2X1 U10347 ( .IN1(n10427), .IN2(n10426), .Q(n10423) );
  OR2X1 U10348 ( .IN1(n10428), .IN2(n10429), .Q(n10426) );
  AND2X1 U10349 ( .IN1(n9451), .IN2(WX9850), .Q(n10429) );
  AND2X1 U10350 ( .IN1(n7923), .IN2(n9472), .Q(n10428) );
  AND2X1 U10351 ( .IN1(n10430), .IN2(n10431), .Q(n10427) );
  OR2X1 U10352 ( .IN1(n10432), .IN2(n8780), .Q(n10431) );
  OR2X1 U10353 ( .IN1(WX9914), .IN2(n10433), .Q(n10430) );
  INVX0 U10354 ( .INP(n10432), .ZN(n10433) );
  AND2X1 U10355 ( .IN1(n10434), .IN2(n10435), .Q(n10432) );
  OR2X1 U10356 ( .IN1(n8306), .IN2(test_so82), .Q(n10435) );
  OR2X1 U10357 ( .IN1(n9114), .IN2(n15879), .Q(n10434) );
  AND2X1 U10358 ( .IN1(n9242), .IN2(CRC_OUT_3_18), .Q(n10419) );
  AND2X1 U10359 ( .IN1(n1484), .IN2(n9216), .Q(n10418) );
  INVX0 U10360 ( .INP(n10436), .ZN(n1484) );
  OR2X1 U10361 ( .IN1(n9573), .IN2(n3866), .Q(n10436) );
  OR4X1 U10362 ( .IN1(n10437), .IN2(n10438), .IN3(n10439), .IN4(n10440), .Q(
        WX8426) );
  AND2X1 U10363 ( .IN1(n9182), .IN2(n10441), .Q(n10440) );
  AND2X1 U10364 ( .IN1(n9272), .IN2(n9955), .Q(n10439) );
  OR2X1 U10365 ( .IN1(n10442), .IN2(n10443), .Q(n9955) );
  INVX0 U10366 ( .INP(n10444), .ZN(n10443) );
  OR2X1 U10367 ( .IN1(n10445), .IN2(n10446), .Q(n10444) );
  AND2X1 U10368 ( .IN1(n10446), .IN2(n10445), .Q(n10442) );
  AND2X1 U10369 ( .IN1(n10447), .IN2(n10448), .Q(n10445) );
  OR2X1 U10370 ( .IN1(n9452), .IN2(n7924), .Q(n10448) );
  OR2X1 U10371 ( .IN1(WX9784), .IN2(n9448), .Q(n10447) );
  OR2X1 U10372 ( .IN1(n10449), .IN2(n10450), .Q(n10446) );
  INVX0 U10373 ( .INP(n10451), .ZN(n10450) );
  OR2X1 U10374 ( .IN1(n10452), .IN2(n7925), .Q(n10451) );
  AND2X1 U10375 ( .IN1(n7925), .IN2(n10452), .Q(n10449) );
  INVX0 U10376 ( .INP(n10453), .ZN(n10452) );
  OR2X1 U10377 ( .IN1(n10454), .IN2(n10455), .Q(n10453) );
  AND2X1 U10378 ( .IN1(n8779), .IN2(n8307), .Q(n10455) );
  AND2X1 U10379 ( .IN1(n15880), .IN2(WX9912), .Q(n10454) );
  AND2X1 U10380 ( .IN1(n9242), .IN2(CRC_OUT_3_19), .Q(n10438) );
  AND2X1 U10381 ( .IN1(n1483), .IN2(n9216), .Q(n10437) );
  INVX0 U10382 ( .INP(n10456), .ZN(n1483) );
  OR2X1 U10383 ( .IN1(n9573), .IN2(n3867), .Q(n10456) );
  OR4X1 U10384 ( .IN1(n10457), .IN2(n10458), .IN3(n10459), .IN4(n10460), .Q(
        WX8424) );
  AND2X1 U10385 ( .IN1(n9182), .IN2(n10461), .Q(n10460) );
  AND2X1 U10386 ( .IN1(n9962), .IN2(n9260), .Q(n10459) );
  AND2X1 U10387 ( .IN1(n10462), .IN2(n10463), .Q(n9962) );
  OR2X1 U10388 ( .IN1(n10464), .IN2(n10465), .Q(n10463) );
  INVX0 U10389 ( .INP(n10466), .ZN(n10462) );
  AND2X1 U10390 ( .IN1(n10465), .IN2(n10464), .Q(n10466) );
  INVX0 U10391 ( .INP(n10467), .ZN(n10464) );
  OR2X1 U10392 ( .IN1(n10468), .IN2(n10469), .Q(n10467) );
  AND2X1 U10393 ( .IN1(n9451), .IN2(WX9910), .Q(n10469) );
  AND2X1 U10394 ( .IN1(n8778), .IN2(n9458), .Q(n10468) );
  OR2X1 U10395 ( .IN1(n10470), .IN2(n10471), .Q(n10465) );
  AND3X1 U10396 ( .IN1(n10472), .IN2(n10473), .IN3(n7927), .Q(n10471) );
  OR2X1 U10397 ( .IN1(n7926), .IN2(n9091), .Q(n10473) );
  OR2X1 U10398 ( .IN1(test_so80), .IN2(WX9782), .Q(n10472) );
  AND2X1 U10399 ( .IN1(n10474), .IN2(WX9846), .Q(n10470) );
  OR2X1 U10400 ( .IN1(n10475), .IN2(n10476), .Q(n10474) );
  AND2X1 U10401 ( .IN1(n7926), .IN2(n9091), .Q(n10476) );
  AND2X1 U10402 ( .IN1(test_so80), .IN2(WX9782), .Q(n10475) );
  AND2X1 U10403 ( .IN1(n9242), .IN2(CRC_OUT_3_20), .Q(n10458) );
  AND2X1 U10404 ( .IN1(n1482), .IN2(n9216), .Q(n10457) );
  INVX0 U10405 ( .INP(n10477), .ZN(n1482) );
  OR2X1 U10406 ( .IN1(n9573), .IN2(n3868), .Q(n10477) );
  OR4X1 U10407 ( .IN1(n10478), .IN2(n10479), .IN3(n10480), .IN4(n10481), .Q(
        WX8422) );
  AND2X1 U10408 ( .IN1(n9182), .IN2(n10482), .Q(n10481) );
  AND2X1 U10409 ( .IN1(n9273), .IN2(n9969), .Q(n10480) );
  OR2X1 U10410 ( .IN1(n10483), .IN2(n10484), .Q(n9969) );
  INVX0 U10411 ( .INP(n10485), .ZN(n10484) );
  OR2X1 U10412 ( .IN1(n10486), .IN2(n10487), .Q(n10485) );
  AND2X1 U10413 ( .IN1(n10487), .IN2(n10486), .Q(n10483) );
  AND2X1 U10414 ( .IN1(n10488), .IN2(n10489), .Q(n10486) );
  OR2X1 U10415 ( .IN1(n9456), .IN2(n7928), .Q(n10489) );
  OR2X1 U10416 ( .IN1(WX9780), .IN2(n9449), .Q(n10488) );
  OR2X1 U10417 ( .IN1(n10490), .IN2(n10491), .Q(n10487) );
  INVX0 U10418 ( .INP(n10492), .ZN(n10491) );
  OR2X1 U10419 ( .IN1(n10493), .IN2(n7929), .Q(n10492) );
  AND2X1 U10420 ( .IN1(n7929), .IN2(n10493), .Q(n10490) );
  INVX0 U10421 ( .INP(n10494), .ZN(n10493) );
  OR2X1 U10422 ( .IN1(n10495), .IN2(n10496), .Q(n10494) );
  AND2X1 U10423 ( .IN1(n8777), .IN2(n8310), .Q(n10496) );
  AND2X1 U10424 ( .IN1(n15881), .IN2(WX9908), .Q(n10495) );
  AND2X1 U10425 ( .IN1(n9242), .IN2(CRC_OUT_3_21), .Q(n10479) );
  AND2X1 U10426 ( .IN1(n1481), .IN2(n9216), .Q(n10478) );
  INVX0 U10427 ( .INP(n10497), .ZN(n1481) );
  OR2X1 U10428 ( .IN1(n9573), .IN2(n3869), .Q(n10497) );
  OR4X1 U10429 ( .IN1(n10498), .IN2(n10499), .IN3(n10500), .IN4(n10501), .Q(
        WX8420) );
  AND2X1 U10430 ( .IN1(n9182), .IN2(n10502), .Q(n10501) );
  AND2X1 U10431 ( .IN1(n9273), .IN2(n9976), .Q(n10500) );
  OR2X1 U10432 ( .IN1(n10503), .IN2(n10504), .Q(n9976) );
  INVX0 U10433 ( .INP(n10505), .ZN(n10504) );
  OR2X1 U10434 ( .IN1(n10506), .IN2(n10507), .Q(n10505) );
  AND2X1 U10435 ( .IN1(n10507), .IN2(n10506), .Q(n10503) );
  AND2X1 U10436 ( .IN1(n10508), .IN2(n10509), .Q(n10506) );
  OR2X1 U10437 ( .IN1(n9454), .IN2(n7930), .Q(n10509) );
  OR2X1 U10438 ( .IN1(WX9778), .IN2(n9448), .Q(n10508) );
  OR2X1 U10439 ( .IN1(n10510), .IN2(n10511), .Q(n10507) );
  INVX0 U10440 ( .INP(n10512), .ZN(n10511) );
  OR2X1 U10441 ( .IN1(n10513), .IN2(n7931), .Q(n10512) );
  AND2X1 U10442 ( .IN1(n7931), .IN2(n10513), .Q(n10510) );
  INVX0 U10443 ( .INP(n10514), .ZN(n10513) );
  OR2X1 U10444 ( .IN1(n10515), .IN2(n10516), .Q(n10514) );
  AND2X1 U10445 ( .IN1(n8776), .IN2(n8311), .Q(n10516) );
  AND2X1 U10446 ( .IN1(n15882), .IN2(WX9906), .Q(n10515) );
  AND2X1 U10447 ( .IN1(n9242), .IN2(CRC_OUT_3_22), .Q(n10499) );
  AND2X1 U10448 ( .IN1(n1480), .IN2(n9216), .Q(n10498) );
  INVX0 U10449 ( .INP(n10517), .ZN(n1480) );
  OR2X1 U10450 ( .IN1(n9573), .IN2(n3870), .Q(n10517) );
  OR4X1 U10451 ( .IN1(n10518), .IN2(n10519), .IN3(n10520), .IN4(n10521), .Q(
        WX8418) );
  AND2X1 U10452 ( .IN1(n9182), .IN2(n10522), .Q(n10521) );
  AND2X1 U10453 ( .IN1(n9273), .IN2(n9983), .Q(n10520) );
  OR2X1 U10454 ( .IN1(n10523), .IN2(n10524), .Q(n9983) );
  INVX0 U10455 ( .INP(n10525), .ZN(n10524) );
  OR2X1 U10456 ( .IN1(n10526), .IN2(n10527), .Q(n10525) );
  AND2X1 U10457 ( .IN1(n10527), .IN2(n10526), .Q(n10523) );
  AND2X1 U10458 ( .IN1(n10528), .IN2(n10529), .Q(n10526) );
  OR2X1 U10459 ( .IN1(n9482), .IN2(n7932), .Q(n10529) );
  OR2X1 U10460 ( .IN1(WX9776), .IN2(n9449), .Q(n10528) );
  OR2X1 U10461 ( .IN1(n10530), .IN2(n10531), .Q(n10527) );
  INVX0 U10462 ( .INP(n10532), .ZN(n10531) );
  OR2X1 U10463 ( .IN1(n10533), .IN2(n7933), .Q(n10532) );
  AND2X1 U10464 ( .IN1(n7933), .IN2(n10533), .Q(n10530) );
  INVX0 U10465 ( .INP(n10534), .ZN(n10533) );
  OR2X1 U10466 ( .IN1(n10535), .IN2(n10536), .Q(n10534) );
  AND2X1 U10467 ( .IN1(n8775), .IN2(n8312), .Q(n10536) );
  AND2X1 U10468 ( .IN1(n15883), .IN2(WX9904), .Q(n10535) );
  AND2X1 U10469 ( .IN1(n9242), .IN2(CRC_OUT_3_23), .Q(n10519) );
  AND2X1 U10470 ( .IN1(n1479), .IN2(n9217), .Q(n10518) );
  INVX0 U10471 ( .INP(n10537), .ZN(n1479) );
  OR2X1 U10472 ( .IN1(n9573), .IN2(n3871), .Q(n10537) );
  OR4X1 U10473 ( .IN1(n10538), .IN2(n10539), .IN3(n10540), .IN4(n10541), .Q(
        WX8416) );
  AND2X1 U10474 ( .IN1(n9182), .IN2(n10542), .Q(n10541) );
  AND2X1 U10475 ( .IN1(n9273), .IN2(n9990), .Q(n10540) );
  OR2X1 U10476 ( .IN1(n10543), .IN2(n10544), .Q(n9990) );
  INVX0 U10477 ( .INP(n10545), .ZN(n10544) );
  OR2X1 U10478 ( .IN1(n10546), .IN2(n10547), .Q(n10545) );
  AND2X1 U10479 ( .IN1(n10547), .IN2(n10546), .Q(n10543) );
  AND2X1 U10480 ( .IN1(n10548), .IN2(n10549), .Q(n10546) );
  OR2X1 U10481 ( .IN1(n9482), .IN2(n7934), .Q(n10549) );
  OR2X1 U10482 ( .IN1(WX9774), .IN2(n9448), .Q(n10548) );
  OR2X1 U10483 ( .IN1(n10550), .IN2(n10551), .Q(n10547) );
  INVX0 U10484 ( .INP(n10552), .ZN(n10551) );
  OR2X1 U10485 ( .IN1(n10553), .IN2(n7935), .Q(n10552) );
  AND2X1 U10486 ( .IN1(n7935), .IN2(n10553), .Q(n10550) );
  INVX0 U10487 ( .INP(n10554), .ZN(n10553) );
  OR2X1 U10488 ( .IN1(n10555), .IN2(n10556), .Q(n10554) );
  AND2X1 U10489 ( .IN1(n8774), .IN2(n8313), .Q(n10556) );
  AND2X1 U10490 ( .IN1(n15884), .IN2(WX9902), .Q(n10555) );
  AND2X1 U10491 ( .IN1(test_so77), .IN2(n9227), .Q(n10539) );
  AND2X1 U10492 ( .IN1(n1478), .IN2(n9217), .Q(n10538) );
  INVX0 U10493 ( .INP(n10557), .ZN(n1478) );
  OR2X1 U10494 ( .IN1(n9573), .IN2(n3872), .Q(n10557) );
  OR4X1 U10495 ( .IN1(n10558), .IN2(n10559), .IN3(n10560), .IN4(n10561), .Q(
        WX8414) );
  AND2X1 U10496 ( .IN1(n9182), .IN2(n10562), .Q(n10561) );
  AND2X1 U10497 ( .IN1(n9273), .IN2(n9997), .Q(n10560) );
  OR2X1 U10498 ( .IN1(n10563), .IN2(n10564), .Q(n9997) );
  INVX0 U10499 ( .INP(n10565), .ZN(n10564) );
  OR2X1 U10500 ( .IN1(n10566), .IN2(n10567), .Q(n10565) );
  AND2X1 U10501 ( .IN1(n10567), .IN2(n10566), .Q(n10563) );
  AND2X1 U10502 ( .IN1(n10568), .IN2(n10569), .Q(n10566) );
  OR2X1 U10503 ( .IN1(n9481), .IN2(n7936), .Q(n10569) );
  OR2X1 U10504 ( .IN1(WX9772), .IN2(n9449), .Q(n10568) );
  OR2X1 U10505 ( .IN1(n10570), .IN2(n10571), .Q(n10567) );
  INVX0 U10506 ( .INP(n10572), .ZN(n10571) );
  OR2X1 U10507 ( .IN1(n10573), .IN2(n7937), .Q(n10572) );
  AND2X1 U10508 ( .IN1(n7937), .IN2(n10573), .Q(n10570) );
  INVX0 U10509 ( .INP(n10574), .ZN(n10573) );
  OR2X1 U10510 ( .IN1(n10575), .IN2(n10576), .Q(n10574) );
  AND2X1 U10511 ( .IN1(n8773), .IN2(n8314), .Q(n10576) );
  AND2X1 U10512 ( .IN1(n15885), .IN2(WX9900), .Q(n10575) );
  AND2X1 U10513 ( .IN1(n9242), .IN2(CRC_OUT_3_25), .Q(n10559) );
  AND2X1 U10514 ( .IN1(n1477), .IN2(n9217), .Q(n10558) );
  INVX0 U10515 ( .INP(n10577), .ZN(n1477) );
  OR2X1 U10516 ( .IN1(n9572), .IN2(n3873), .Q(n10577) );
  OR4X1 U10517 ( .IN1(n10578), .IN2(n10579), .IN3(n10580), .IN4(n10581), .Q(
        WX8412) );
  AND2X1 U10518 ( .IN1(n10582), .IN2(n9177), .Q(n10581) );
  AND2X1 U10519 ( .IN1(n9273), .IN2(n10004), .Q(n10580) );
  OR2X1 U10520 ( .IN1(n10583), .IN2(n10584), .Q(n10004) );
  INVX0 U10521 ( .INP(n10585), .ZN(n10584) );
  OR2X1 U10522 ( .IN1(n10586), .IN2(n10587), .Q(n10585) );
  AND2X1 U10523 ( .IN1(n10587), .IN2(n10586), .Q(n10583) );
  AND2X1 U10524 ( .IN1(n10588), .IN2(n10589), .Q(n10586) );
  OR2X1 U10525 ( .IN1(n9481), .IN2(n7938), .Q(n10589) );
  OR2X1 U10526 ( .IN1(WX9770), .IN2(n9449), .Q(n10588) );
  OR2X1 U10527 ( .IN1(n10590), .IN2(n10591), .Q(n10587) );
  INVX0 U10528 ( .INP(n10592), .ZN(n10591) );
  OR2X1 U10529 ( .IN1(n10593), .IN2(n7939), .Q(n10592) );
  AND2X1 U10530 ( .IN1(n7939), .IN2(n10593), .Q(n10590) );
  INVX0 U10531 ( .INP(n10594), .ZN(n10593) );
  OR2X1 U10532 ( .IN1(n10595), .IN2(n10596), .Q(n10594) );
  AND2X1 U10533 ( .IN1(n8772), .IN2(n8315), .Q(n10596) );
  AND2X1 U10534 ( .IN1(n15886), .IN2(WX9898), .Q(n10595) );
  AND2X1 U10535 ( .IN1(n9242), .IN2(CRC_OUT_3_26), .Q(n10579) );
  AND2X1 U10536 ( .IN1(n1476), .IN2(n9217), .Q(n10578) );
  INVX0 U10537 ( .INP(n10597), .ZN(n1476) );
  OR2X1 U10538 ( .IN1(n9572), .IN2(n3874), .Q(n10597) );
  OR4X1 U10539 ( .IN1(n10598), .IN2(n10599), .IN3(n10600), .IN4(n10601), .Q(
        WX8410) );
  AND2X1 U10540 ( .IN1(n9182), .IN2(n10602), .Q(n10601) );
  AND2X1 U10541 ( .IN1(n9273), .IN2(n10011), .Q(n10600) );
  OR2X1 U10542 ( .IN1(n10603), .IN2(n10604), .Q(n10011) );
  INVX0 U10543 ( .INP(n10605), .ZN(n10604) );
  OR2X1 U10544 ( .IN1(n10606), .IN2(n10607), .Q(n10605) );
  AND2X1 U10545 ( .IN1(n10607), .IN2(n10606), .Q(n10603) );
  AND2X1 U10546 ( .IN1(n10608), .IN2(n10609), .Q(n10606) );
  OR2X1 U10547 ( .IN1(n9482), .IN2(n7940), .Q(n10609) );
  OR2X1 U10548 ( .IN1(WX9768), .IN2(n9449), .Q(n10608) );
  OR2X1 U10549 ( .IN1(n10610), .IN2(n10611), .Q(n10607) );
  INVX0 U10550 ( .INP(n10612), .ZN(n10611) );
  OR2X1 U10551 ( .IN1(n10613), .IN2(n7941), .Q(n10612) );
  AND2X1 U10552 ( .IN1(n7941), .IN2(n10613), .Q(n10610) );
  INVX0 U10553 ( .INP(n10614), .ZN(n10613) );
  OR2X1 U10554 ( .IN1(n10615), .IN2(n10616), .Q(n10614) );
  AND2X1 U10555 ( .IN1(n8771), .IN2(n8316), .Q(n10616) );
  AND2X1 U10556 ( .IN1(n15887), .IN2(WX9896), .Q(n10615) );
  AND2X1 U10557 ( .IN1(n9242), .IN2(CRC_OUT_3_27), .Q(n10599) );
  AND2X1 U10558 ( .IN1(n1475), .IN2(n9217), .Q(n10598) );
  INVX0 U10559 ( .INP(n10617), .ZN(n1475) );
  OR2X1 U10560 ( .IN1(n9572), .IN2(n3875), .Q(n10617) );
  OR4X1 U10561 ( .IN1(n10618), .IN2(n10619), .IN3(n10620), .IN4(n10621), .Q(
        WX8408) );
  AND2X1 U10562 ( .IN1(n10622), .IN2(n9178), .Q(n10621) );
  AND2X1 U10563 ( .IN1(n9273), .IN2(n10018), .Q(n10620) );
  OR2X1 U10564 ( .IN1(n10623), .IN2(n10624), .Q(n10018) );
  INVX0 U10565 ( .INP(n10625), .ZN(n10624) );
  OR2X1 U10566 ( .IN1(n10626), .IN2(n10627), .Q(n10625) );
  AND2X1 U10567 ( .IN1(n10627), .IN2(n10626), .Q(n10623) );
  AND2X1 U10568 ( .IN1(n10628), .IN2(n10629), .Q(n10626) );
  OR2X1 U10569 ( .IN1(n9481), .IN2(n7942), .Q(n10629) );
  OR2X1 U10570 ( .IN1(WX9766), .IN2(n9447), .Q(n10628) );
  OR2X1 U10571 ( .IN1(n10630), .IN2(n10631), .Q(n10627) );
  INVX0 U10572 ( .INP(n10632), .ZN(n10631) );
  OR2X1 U10573 ( .IN1(n10633), .IN2(n7943), .Q(n10632) );
  AND2X1 U10574 ( .IN1(n7943), .IN2(n10633), .Q(n10630) );
  INVX0 U10575 ( .INP(n10634), .ZN(n10633) );
  OR2X1 U10576 ( .IN1(n10635), .IN2(n10636), .Q(n10634) );
  AND2X1 U10577 ( .IN1(n8770), .IN2(n8317), .Q(n10636) );
  AND2X1 U10578 ( .IN1(n15888), .IN2(WX9894), .Q(n10635) );
  AND2X1 U10579 ( .IN1(n9242), .IN2(CRC_OUT_3_28), .Q(n10619) );
  AND2X1 U10580 ( .IN1(n1474), .IN2(n9217), .Q(n10618) );
  INVX0 U10581 ( .INP(n10637), .ZN(n1474) );
  OR2X1 U10582 ( .IN1(n9572), .IN2(n3876), .Q(n10637) );
  OR4X1 U10583 ( .IN1(n10638), .IN2(n10639), .IN3(n10640), .IN4(n10641), .Q(
        WX8406) );
  AND2X1 U10584 ( .IN1(n9182), .IN2(n10642), .Q(n10641) );
  AND2X1 U10585 ( .IN1(n9273), .IN2(n10025), .Q(n10640) );
  OR2X1 U10586 ( .IN1(n10643), .IN2(n10644), .Q(n10025) );
  INVX0 U10587 ( .INP(n10645), .ZN(n10644) );
  OR2X1 U10588 ( .IN1(n10646), .IN2(n10647), .Q(n10645) );
  AND2X1 U10589 ( .IN1(n10647), .IN2(n10646), .Q(n10643) );
  AND2X1 U10590 ( .IN1(n10648), .IN2(n10649), .Q(n10646) );
  OR2X1 U10591 ( .IN1(n9481), .IN2(n7944), .Q(n10649) );
  OR2X1 U10592 ( .IN1(WX9764), .IN2(n9448), .Q(n10648) );
  OR2X1 U10593 ( .IN1(n10650), .IN2(n10651), .Q(n10647) );
  INVX0 U10594 ( .INP(n10652), .ZN(n10651) );
  OR2X1 U10595 ( .IN1(n10653), .IN2(n7945), .Q(n10652) );
  AND2X1 U10596 ( .IN1(n7945), .IN2(n10653), .Q(n10650) );
  INVX0 U10597 ( .INP(n10654), .ZN(n10653) );
  OR2X1 U10598 ( .IN1(n10655), .IN2(n10656), .Q(n10654) );
  AND2X1 U10599 ( .IN1(n8769), .IN2(n8318), .Q(n10656) );
  AND2X1 U10600 ( .IN1(n15889), .IN2(WX9892), .Q(n10655) );
  AND2X1 U10601 ( .IN1(n9242), .IN2(CRC_OUT_3_29), .Q(n10639) );
  AND2X1 U10602 ( .IN1(n1473), .IN2(n9217), .Q(n10638) );
  INVX0 U10603 ( .INP(n10657), .ZN(n1473) );
  OR2X1 U10604 ( .IN1(n9572), .IN2(n3877), .Q(n10657) );
  OR4X1 U10605 ( .IN1(n10658), .IN2(n10659), .IN3(n10660), .IN4(n10661), .Q(
        WX8404) );
  AND2X1 U10606 ( .IN1(n10662), .IN2(n9177), .Q(n10661) );
  AND2X1 U10607 ( .IN1(n9273), .IN2(n10032), .Q(n10660) );
  OR2X1 U10608 ( .IN1(n10663), .IN2(n10664), .Q(n10032) );
  INVX0 U10609 ( .INP(n10665), .ZN(n10664) );
  OR2X1 U10610 ( .IN1(n10666), .IN2(n10667), .Q(n10665) );
  AND2X1 U10611 ( .IN1(n10667), .IN2(n10666), .Q(n10663) );
  AND2X1 U10612 ( .IN1(n10668), .IN2(n10669), .Q(n10666) );
  OR2X1 U10613 ( .IN1(n9452), .IN2(n7946), .Q(n10669) );
  OR2X1 U10614 ( .IN1(WX9762), .IN2(n9449), .Q(n10668) );
  OR2X1 U10615 ( .IN1(n10670), .IN2(n10671), .Q(n10667) );
  INVX0 U10616 ( .INP(n10672), .ZN(n10671) );
  OR2X1 U10617 ( .IN1(n10673), .IN2(n7947), .Q(n10672) );
  AND2X1 U10618 ( .IN1(n7947), .IN2(n10673), .Q(n10670) );
  INVX0 U10619 ( .INP(n10674), .ZN(n10673) );
  OR2X1 U10620 ( .IN1(n10675), .IN2(n10676), .Q(n10674) );
  AND2X1 U10621 ( .IN1(n8768), .IN2(n8319), .Q(n10676) );
  AND2X1 U10622 ( .IN1(n15890), .IN2(WX9890), .Q(n10675) );
  AND2X1 U10623 ( .IN1(n9242), .IN2(CRC_OUT_3_30), .Q(n10659) );
  AND2X1 U10624 ( .IN1(n1472), .IN2(n9217), .Q(n10658) );
  INVX0 U10625 ( .INP(n10677), .ZN(n1472) );
  OR2X1 U10626 ( .IN1(n9572), .IN2(n3878), .Q(n10677) );
  OR4X1 U10627 ( .IN1(n10678), .IN2(n10679), .IN3(n10680), .IN4(n10681), .Q(
        WX8402) );
  AND2X1 U10628 ( .IN1(n9182), .IN2(n10682), .Q(n10681) );
  AND2X1 U10629 ( .IN1(n10039), .IN2(n9260), .Q(n10680) );
  AND2X1 U10630 ( .IN1(n10683), .IN2(n10684), .Q(n10039) );
  INVX0 U10631 ( .INP(n10685), .ZN(n10684) );
  AND2X1 U10632 ( .IN1(n10686), .IN2(n10687), .Q(n10685) );
  OR2X1 U10633 ( .IN1(n10687), .IN2(n10686), .Q(n10683) );
  OR2X1 U10634 ( .IN1(n10688), .IN2(n10689), .Q(n10686) );
  AND2X1 U10635 ( .IN1(n9451), .IN2(WX9760), .Q(n10689) );
  AND2X1 U10636 ( .IN1(n7878), .IN2(n9469), .Q(n10688) );
  AND2X1 U10637 ( .IN1(n10690), .IN2(n10691), .Q(n10687) );
  OR2X1 U10638 ( .IN1(n10692), .IN2(n7879), .Q(n10691) );
  INVX0 U10639 ( .INP(n10693), .ZN(n10692) );
  OR2X1 U10640 ( .IN1(WX9824), .IN2(n10693), .Q(n10690) );
  OR2X1 U10641 ( .IN1(n10694), .IN2(n10695), .Q(n10693) );
  AND2X1 U10642 ( .IN1(n15891), .IN2(n9110), .Q(n10695) );
  AND2X1 U10643 ( .IN1(test_so85), .IN2(n8320), .Q(n10694) );
  AND2X1 U10644 ( .IN1(n2245), .IN2(WX8243), .Q(n10679) );
  AND2X1 U10645 ( .IN1(n9243), .IN2(CRC_OUT_3_31), .Q(n10678) );
  AND2X1 U10646 ( .IN1(n9050), .IN2(n9492), .Q(WX8304) );
  AND3X1 U10647 ( .IN1(n10696), .IN2(n10697), .IN3(n9514), .Q(WX7791) );
  OR2X1 U10648 ( .IN1(DFF_1150_n1), .IN2(WX7302), .Q(n10697) );
  OR2X1 U10649 ( .IN1(n8820), .IN2(CRC_OUT_4_30), .Q(n10696) );
  AND2X1 U10650 ( .IN1(n10698), .IN2(n9495), .Q(WX7789) );
  OR2X1 U10651 ( .IN1(n10699), .IN2(n10700), .Q(n10698) );
  AND2X1 U10652 ( .IN1(n8821), .IN2(n9152), .Q(n10700) );
  AND2X1 U10653 ( .IN1(test_so66), .IN2(WX7304), .Q(n10699) );
  AND3X1 U10654 ( .IN1(n10701), .IN2(n10702), .IN3(n9513), .Q(WX7787) );
  OR2X1 U10655 ( .IN1(DFF_1148_n1), .IN2(WX7306), .Q(n10702) );
  OR2X1 U10656 ( .IN1(n8822), .IN2(CRC_OUT_4_28), .Q(n10701) );
  AND3X1 U10657 ( .IN1(n10703), .IN2(n10704), .IN3(n9513), .Q(WX7785) );
  OR2X1 U10658 ( .IN1(DFF_1147_n1), .IN2(WX7308), .Q(n10704) );
  OR2X1 U10659 ( .IN1(n8823), .IN2(CRC_OUT_4_27), .Q(n10703) );
  AND3X1 U10660 ( .IN1(n10705), .IN2(n10706), .IN3(n9514), .Q(WX7783) );
  OR2X1 U10661 ( .IN1(DFF_1146_n1), .IN2(WX7310), .Q(n10706) );
  OR2X1 U10662 ( .IN1(n8824), .IN2(CRC_OUT_4_26), .Q(n10705) );
  AND3X1 U10663 ( .IN1(n10707), .IN2(n10708), .IN3(n9513), .Q(WX7781) );
  OR2X1 U10664 ( .IN1(DFF_1145_n1), .IN2(WX7312), .Q(n10708) );
  OR2X1 U10665 ( .IN1(n8825), .IN2(CRC_OUT_4_25), .Q(n10707) );
  AND3X1 U10666 ( .IN1(n10709), .IN2(n10710), .IN3(n9514), .Q(WX7779) );
  OR2X1 U10667 ( .IN1(DFF_1144_n1), .IN2(WX7314), .Q(n10710) );
  OR2X1 U10668 ( .IN1(n8826), .IN2(CRC_OUT_4_24), .Q(n10709) );
  AND3X1 U10669 ( .IN1(n10711), .IN2(n10712), .IN3(n9513), .Q(WX7777) );
  OR2X1 U10670 ( .IN1(DFF_1143_n1), .IN2(WX7316), .Q(n10712) );
  OR2X1 U10671 ( .IN1(n8827), .IN2(CRC_OUT_4_23), .Q(n10711) );
  AND3X1 U10672 ( .IN1(n10713), .IN2(n10714), .IN3(n9514), .Q(WX7775) );
  OR2X1 U10673 ( .IN1(DFF_1142_n1), .IN2(WX7318), .Q(n10714) );
  OR2X1 U10674 ( .IN1(n8828), .IN2(CRC_OUT_4_22), .Q(n10713) );
  AND3X1 U10675 ( .IN1(n10715), .IN2(n10716), .IN3(n9515), .Q(WX7773) );
  OR2X1 U10676 ( .IN1(DFF_1141_n1), .IN2(WX7320), .Q(n10716) );
  OR2X1 U10677 ( .IN1(n8829), .IN2(CRC_OUT_4_21), .Q(n10715) );
  AND2X1 U10678 ( .IN1(n10717), .IN2(n9494), .Q(WX7771) );
  OR2X1 U10679 ( .IN1(n10718), .IN2(n10719), .Q(n10717) );
  AND2X1 U10680 ( .IN1(DFF_1140_n1), .IN2(n9105), .Q(n10719) );
  AND2X1 U10681 ( .IN1(test_so63), .IN2(CRC_OUT_4_20), .Q(n10718) );
  AND3X1 U10682 ( .IN1(n10720), .IN2(n10721), .IN3(n9514), .Q(WX7769) );
  OR2X1 U10683 ( .IN1(DFF_1139_n1), .IN2(WX7324), .Q(n10721) );
  OR2X1 U10684 ( .IN1(n8830), .IN2(CRC_OUT_4_19), .Q(n10720) );
  AND3X1 U10685 ( .IN1(n10722), .IN2(n10723), .IN3(n9513), .Q(WX7767) );
  OR2X1 U10686 ( .IN1(DFF_1138_n1), .IN2(WX7326), .Q(n10723) );
  OR2X1 U10687 ( .IN1(n8831), .IN2(CRC_OUT_4_18), .Q(n10722) );
  AND3X1 U10688 ( .IN1(n10724), .IN2(n10725), .IN3(n9513), .Q(WX7765) );
  OR2X1 U10689 ( .IN1(DFF_1137_n1), .IN2(WX7328), .Q(n10725) );
  OR2X1 U10690 ( .IN1(n8832), .IN2(CRC_OUT_4_17), .Q(n10724) );
  AND3X1 U10691 ( .IN1(n10726), .IN2(n10727), .IN3(n9514), .Q(WX7763) );
  OR2X1 U10692 ( .IN1(DFF_1136_n1), .IN2(WX7330), .Q(n10727) );
  OR2X1 U10693 ( .IN1(n8833), .IN2(CRC_OUT_4_16), .Q(n10726) );
  AND2X1 U10694 ( .IN1(n10728), .IN2(n9493), .Q(WX7761) );
  OR2X1 U10695 ( .IN1(n10729), .IN2(n10730), .Q(n10728) );
  AND2X1 U10696 ( .IN1(n10731), .IN2(CRC_OUT_4_15), .Q(n10730) );
  AND2X1 U10697 ( .IN1(DFF_1135_n1), .IN2(n10732), .Q(n10729) );
  INVX0 U10698 ( .INP(n10731), .ZN(n10732) );
  OR2X1 U10699 ( .IN1(n10733), .IN2(n10734), .Q(n10731) );
  AND2X1 U10700 ( .IN1(DFF_1151_n1), .IN2(WX7332), .Q(n10734) );
  AND2X1 U10701 ( .IN1(n8722), .IN2(CRC_OUT_4_31), .Q(n10733) );
  AND3X1 U10702 ( .IN1(n10735), .IN2(n10736), .IN3(n9515), .Q(WX7759) );
  OR2X1 U10703 ( .IN1(DFF_1134_n1), .IN2(WX7334), .Q(n10736) );
  OR2X1 U10704 ( .IN1(n8834), .IN2(CRC_OUT_4_14), .Q(n10735) );
  AND3X1 U10705 ( .IN1(n10737), .IN2(n10738), .IN3(n9515), .Q(WX7757) );
  OR2X1 U10706 ( .IN1(DFF_1133_n1), .IN2(WX7336), .Q(n10738) );
  OR2X1 U10707 ( .IN1(n8835), .IN2(CRC_OUT_4_13), .Q(n10737) );
  AND2X1 U10708 ( .IN1(n10739), .IN2(n9495), .Q(WX7755) );
  OR2X1 U10709 ( .IN1(n10740), .IN2(n10741), .Q(n10739) );
  AND2X1 U10710 ( .IN1(n8836), .IN2(n9153), .Q(n10741) );
  AND2X1 U10711 ( .IN1(test_so65), .IN2(WX7338), .Q(n10740) );
  AND3X1 U10712 ( .IN1(n10742), .IN2(n10743), .IN3(n9517), .Q(WX7753) );
  OR2X1 U10713 ( .IN1(DFF_1131_n1), .IN2(WX7340), .Q(n10743) );
  OR2X1 U10714 ( .IN1(n8837), .IN2(CRC_OUT_4_11), .Q(n10742) );
  AND2X1 U10715 ( .IN1(n10744), .IN2(n9495), .Q(WX7751) );
  OR2X1 U10716 ( .IN1(n10745), .IN2(n10746), .Q(n10744) );
  AND2X1 U10717 ( .IN1(n10747), .IN2(CRC_OUT_4_10), .Q(n10746) );
  AND2X1 U10718 ( .IN1(DFF_1130_n1), .IN2(n10748), .Q(n10745) );
  INVX0 U10719 ( .INP(n10747), .ZN(n10748) );
  OR2X1 U10720 ( .IN1(n10749), .IN2(n10750), .Q(n10747) );
  AND2X1 U10721 ( .IN1(DFF_1151_n1), .IN2(WX7342), .Q(n10750) );
  AND2X1 U10722 ( .IN1(n8723), .IN2(CRC_OUT_4_31), .Q(n10749) );
  AND3X1 U10723 ( .IN1(n10751), .IN2(n10752), .IN3(n9515), .Q(WX7749) );
  OR2X1 U10724 ( .IN1(DFF_1129_n1), .IN2(WX7344), .Q(n10752) );
  OR2X1 U10725 ( .IN1(n8838), .IN2(CRC_OUT_4_9), .Q(n10751) );
  AND3X1 U10726 ( .IN1(n10753), .IN2(n10754), .IN3(n9515), .Q(WX7747) );
  OR2X1 U10727 ( .IN1(DFF_1128_n1), .IN2(WX7346), .Q(n10754) );
  OR2X1 U10728 ( .IN1(n8839), .IN2(CRC_OUT_4_8), .Q(n10753) );
  AND3X1 U10729 ( .IN1(n10755), .IN2(n10756), .IN3(n9515), .Q(WX7745) );
  OR2X1 U10730 ( .IN1(DFF_1127_n1), .IN2(WX7348), .Q(n10756) );
  OR2X1 U10731 ( .IN1(n8840), .IN2(CRC_OUT_4_7), .Q(n10755) );
  AND3X1 U10732 ( .IN1(n10757), .IN2(n10758), .IN3(n9516), .Q(WX7743) );
  OR2X1 U10733 ( .IN1(DFF_1126_n1), .IN2(WX7350), .Q(n10758) );
  OR2X1 U10734 ( .IN1(n8841), .IN2(CRC_OUT_4_6), .Q(n10757) );
  AND3X1 U10735 ( .IN1(n10759), .IN2(n10760), .IN3(n9516), .Q(WX7741) );
  OR2X1 U10736 ( .IN1(DFF_1125_n1), .IN2(WX7352), .Q(n10760) );
  OR2X1 U10737 ( .IN1(n8842), .IN2(CRC_OUT_4_5), .Q(n10759) );
  AND3X1 U10738 ( .IN1(n10761), .IN2(n10762), .IN3(n9515), .Q(WX7739) );
  OR2X1 U10739 ( .IN1(DFF_1124_n1), .IN2(WX7354), .Q(n10762) );
  OR2X1 U10740 ( .IN1(n8843), .IN2(CRC_OUT_4_4), .Q(n10761) );
  AND3X1 U10741 ( .IN1(n10763), .IN2(n10764), .IN3(n9516), .Q(WX7737) );
  OR2X1 U10742 ( .IN1(DFF_1123_n1), .IN2(n10765), .Q(n10764) );
  AND2X1 U10743 ( .IN1(n10766), .IN2(n10767), .Q(n10765) );
  OR2X1 U10744 ( .IN1(DFF_1151_n1), .IN2(n9087), .Q(n10767) );
  OR2X1 U10745 ( .IN1(test_so64), .IN2(CRC_OUT_4_31), .Q(n10766) );
  OR3X1 U10746 ( .IN1(n10768), .IN2(n10769), .IN3(CRC_OUT_4_3), .Q(n10763) );
  AND2X1 U10747 ( .IN1(DFF_1151_n1), .IN2(n9087), .Q(n10769) );
  AND2X1 U10748 ( .IN1(test_so64), .IN2(CRC_OUT_4_31), .Q(n10768) );
  AND3X1 U10749 ( .IN1(n10770), .IN2(n10771), .IN3(n9516), .Q(WX7735) );
  OR2X1 U10750 ( .IN1(DFF_1122_n1), .IN2(WX7358), .Q(n10771) );
  OR2X1 U10751 ( .IN1(n8844), .IN2(CRC_OUT_4_2), .Q(n10770) );
  AND3X1 U10752 ( .IN1(n10772), .IN2(n10773), .IN3(n9516), .Q(WX7733) );
  OR2X1 U10753 ( .IN1(DFF_1121_n1), .IN2(WX7360), .Q(n10773) );
  OR2X1 U10754 ( .IN1(n8845), .IN2(CRC_OUT_4_1), .Q(n10772) );
  AND3X1 U10755 ( .IN1(n10774), .IN2(n10775), .IN3(n9516), .Q(WX7731) );
  OR2X1 U10756 ( .IN1(DFF_1120_n1), .IN2(WX7362), .Q(n10775) );
  OR2X1 U10757 ( .IN1(n8846), .IN2(CRC_OUT_4_0), .Q(n10774) );
  AND3X1 U10758 ( .IN1(n10776), .IN2(n10777), .IN3(n9516), .Q(WX7729) );
  OR2X1 U10759 ( .IN1(DFF_1151_n1), .IN2(WX7364), .Q(n10777) );
  OR2X1 U10760 ( .IN1(n8737), .IN2(CRC_OUT_4_31), .Q(n10776) );
  AND2X1 U10761 ( .IN1(n9501), .IN2(n8421), .Q(WX7203) );
  AND2X1 U10762 ( .IN1(n9500), .IN2(n8422), .Q(WX7201) );
  AND2X1 U10763 ( .IN1(n9501), .IN2(n8423), .Q(WX7199) );
  AND2X1 U10764 ( .IN1(n9500), .IN2(n8424), .Q(WX7197) );
  AND2X1 U10765 ( .IN1(n9500), .IN2(n8425), .Q(WX7195) );
  AND2X1 U10766 ( .IN1(n9501), .IN2(n8426), .Q(WX7193) );
  AND2X1 U10767 ( .IN1(n9500), .IN2(n8427), .Q(WX7191) );
  AND2X1 U10768 ( .IN1(n9500), .IN2(n8428), .Q(WX7189) );
  AND2X1 U10769 ( .IN1(n9500), .IN2(n8429), .Q(WX7187) );
  AND2X1 U10770 ( .IN1(n9499), .IN2(n8430), .Q(WX7185) );
  AND2X1 U10771 ( .IN1(n9499), .IN2(n8431), .Q(WX7183) );
  AND2X1 U10772 ( .IN1(test_so57), .IN2(n9496), .Q(WX7181) );
  AND2X1 U10773 ( .IN1(n9510), .IN2(n8434), .Q(WX7179) );
  AND2X1 U10774 ( .IN1(n9502), .IN2(n8435), .Q(WX7177) );
  AND2X1 U10775 ( .IN1(n9500), .IN2(n8436), .Q(WX7175) );
  AND2X1 U10776 ( .IN1(n9499), .IN2(n8437), .Q(WX7173) );
  OR4X1 U10777 ( .IN1(n10778), .IN2(n10779), .IN3(n10780), .IN4(n10781), .Q(
        WX7171) );
  AND2X1 U10778 ( .IN1(n9182), .IN2(n10782), .Q(n10781) );
  AND2X1 U10779 ( .IN1(n9273), .IN2(n10127), .Q(n10780) );
  OR2X1 U10780 ( .IN1(n10783), .IN2(n10784), .Q(n10127) );
  INVX0 U10781 ( .INP(n10785), .ZN(n10784) );
  OR2X1 U10782 ( .IN1(n10786), .IN2(n10787), .Q(n10785) );
  AND2X1 U10783 ( .IN1(n10787), .IN2(n10786), .Q(n10783) );
  AND2X1 U10784 ( .IN1(n10788), .IN2(n10789), .Q(n10786) );
  OR2X1 U10785 ( .IN1(WX8529), .IN2(n8179), .Q(n10789) );
  INVX0 U10786 ( .INP(n10790), .ZN(n10788) );
  AND2X1 U10787 ( .IN1(n8179), .IN2(WX8529), .Q(n10790) );
  OR2X1 U10788 ( .IN1(n10791), .IN2(n10792), .Q(n10787) );
  AND2X1 U10789 ( .IN1(n8180), .IN2(WX8657), .Q(n10792) );
  AND2X1 U10790 ( .IN1(n8736), .IN2(WX8593), .Q(n10791) );
  AND2X1 U10791 ( .IN1(n9243), .IN2(CRC_OUT_4_0), .Q(n10779) );
  AND2X1 U10792 ( .IN1(n1261), .IN2(n9217), .Q(n10778) );
  INVX0 U10793 ( .INP(n10793), .ZN(n1261) );
  OR2X1 U10794 ( .IN1(n9572), .IN2(n3879), .Q(n10793) );
  OR4X1 U10795 ( .IN1(n10794), .IN2(n10795), .IN3(n10796), .IN4(n10797), .Q(
        WX7169) );
  AND2X1 U10796 ( .IN1(n9181), .IN2(n10798), .Q(n10797) );
  AND2X1 U10797 ( .IN1(n9273), .IN2(n10143), .Q(n10796) );
  OR2X1 U10798 ( .IN1(n10799), .IN2(n10800), .Q(n10143) );
  INVX0 U10799 ( .INP(n10801), .ZN(n10800) );
  OR2X1 U10800 ( .IN1(n10802), .IN2(n10803), .Q(n10801) );
  AND2X1 U10801 ( .IN1(n10803), .IN2(n10802), .Q(n10799) );
  AND2X1 U10802 ( .IN1(n10804), .IN2(n10805), .Q(n10802) );
  OR2X1 U10803 ( .IN1(WX8527), .IN2(n8181), .Q(n10805) );
  INVX0 U10804 ( .INP(n10806), .ZN(n10804) );
  AND2X1 U10805 ( .IN1(n8181), .IN2(WX8527), .Q(n10806) );
  OR2X1 U10806 ( .IN1(n10807), .IN2(n10808), .Q(n10803) );
  AND2X1 U10807 ( .IN1(n8182), .IN2(WX8655), .Q(n10808) );
  AND2X1 U10808 ( .IN1(n8819), .IN2(WX8591), .Q(n10807) );
  AND2X1 U10809 ( .IN1(n9243), .IN2(CRC_OUT_4_1), .Q(n10795) );
  AND2X1 U10810 ( .IN1(n1260), .IN2(n9217), .Q(n10794) );
  INVX0 U10811 ( .INP(n10809), .ZN(n1260) );
  OR2X1 U10812 ( .IN1(n9572), .IN2(n3880), .Q(n10809) );
  OR4X1 U10813 ( .IN1(n10810), .IN2(n10811), .IN3(n10812), .IN4(n10813), .Q(
        WX7167) );
  AND2X1 U10814 ( .IN1(n9181), .IN2(n10814), .Q(n10813) );
  AND2X1 U10815 ( .IN1(n9273), .IN2(n10159), .Q(n10812) );
  OR2X1 U10816 ( .IN1(n10815), .IN2(n10816), .Q(n10159) );
  INVX0 U10817 ( .INP(n10817), .ZN(n10816) );
  OR2X1 U10818 ( .IN1(n10818), .IN2(n10819), .Q(n10817) );
  AND2X1 U10819 ( .IN1(n10819), .IN2(n10818), .Q(n10815) );
  AND2X1 U10820 ( .IN1(n10820), .IN2(n10821), .Q(n10818) );
  OR2X1 U10821 ( .IN1(WX8525), .IN2(n8183), .Q(n10821) );
  INVX0 U10822 ( .INP(n10822), .ZN(n10820) );
  AND2X1 U10823 ( .IN1(n8183), .IN2(WX8525), .Q(n10822) );
  OR2X1 U10824 ( .IN1(n10823), .IN2(n10824), .Q(n10819) );
  AND2X1 U10825 ( .IN1(n8184), .IN2(WX8653), .Q(n10824) );
  AND2X1 U10826 ( .IN1(n8818), .IN2(WX8589), .Q(n10823) );
  AND2X1 U10827 ( .IN1(n9243), .IN2(CRC_OUT_4_2), .Q(n10811) );
  AND2X1 U10828 ( .IN1(n1259), .IN2(n9217), .Q(n10810) );
  INVX0 U10829 ( .INP(n10825), .ZN(n1259) );
  OR2X1 U10830 ( .IN1(n9572), .IN2(n3881), .Q(n10825) );
  OR4X1 U10831 ( .IN1(n10826), .IN2(n10827), .IN3(n10828), .IN4(n10829), .Q(
        WX7165) );
  AND2X1 U10832 ( .IN1(n9181), .IN2(n10830), .Q(n10829) );
  AND2X1 U10833 ( .IN1(n9274), .IN2(n10175), .Q(n10828) );
  OR2X1 U10834 ( .IN1(n10831), .IN2(n10832), .Q(n10175) );
  INVX0 U10835 ( .INP(n10833), .ZN(n10832) );
  OR2X1 U10836 ( .IN1(n10834), .IN2(n10835), .Q(n10833) );
  AND2X1 U10837 ( .IN1(n10835), .IN2(n10834), .Q(n10831) );
  AND2X1 U10838 ( .IN1(n10836), .IN2(n10837), .Q(n10834) );
  OR2X1 U10839 ( .IN1(WX8523), .IN2(n8185), .Q(n10837) );
  INVX0 U10840 ( .INP(n10838), .ZN(n10836) );
  AND2X1 U10841 ( .IN1(n8185), .IN2(WX8523), .Q(n10838) );
  OR2X1 U10842 ( .IN1(n10839), .IN2(n10840), .Q(n10835) );
  AND2X1 U10843 ( .IN1(n8186), .IN2(WX8651), .Q(n10840) );
  AND2X1 U10844 ( .IN1(n8817), .IN2(WX8587), .Q(n10839) );
  AND2X1 U10845 ( .IN1(n9243), .IN2(CRC_OUT_4_3), .Q(n10827) );
  AND2X1 U10846 ( .IN1(n1258), .IN2(n9217), .Q(n10826) );
  INVX0 U10847 ( .INP(n10841), .ZN(n1258) );
  OR2X1 U10848 ( .IN1(n9572), .IN2(n3882), .Q(n10841) );
  OR4X1 U10849 ( .IN1(n10842), .IN2(n10843), .IN3(n10844), .IN4(n10845), .Q(
        WX7163) );
  AND2X1 U10850 ( .IN1(n10846), .IN2(n9175), .Q(n10845) );
  AND2X1 U10851 ( .IN1(n9274), .IN2(n10191), .Q(n10844) );
  OR2X1 U10852 ( .IN1(n10847), .IN2(n10848), .Q(n10191) );
  INVX0 U10853 ( .INP(n10849), .ZN(n10848) );
  OR2X1 U10854 ( .IN1(n10850), .IN2(n10851), .Q(n10849) );
  AND2X1 U10855 ( .IN1(n10851), .IN2(n10850), .Q(n10847) );
  AND2X1 U10856 ( .IN1(n10852), .IN2(n10853), .Q(n10850) );
  OR2X1 U10857 ( .IN1(WX8521), .IN2(n8187), .Q(n10853) );
  INVX0 U10858 ( .INP(n10854), .ZN(n10852) );
  AND2X1 U10859 ( .IN1(n8187), .IN2(WX8521), .Q(n10854) );
  OR2X1 U10860 ( .IN1(n10855), .IN2(n10856), .Q(n10851) );
  AND2X1 U10861 ( .IN1(n8188), .IN2(WX8649), .Q(n10856) );
  AND2X1 U10862 ( .IN1(n8721), .IN2(WX8585), .Q(n10855) );
  AND2X1 U10863 ( .IN1(n9243), .IN2(CRC_OUT_4_4), .Q(n10843) );
  AND2X1 U10864 ( .IN1(n1257), .IN2(n9218), .Q(n10842) );
  INVX0 U10865 ( .INP(n10857), .ZN(n1257) );
  OR2X1 U10866 ( .IN1(n9572), .IN2(n3883), .Q(n10857) );
  OR4X1 U10867 ( .IN1(n10858), .IN2(n10859), .IN3(n10860), .IN4(n10861), .Q(
        WX7161) );
  AND2X1 U10868 ( .IN1(n9181), .IN2(n10862), .Q(n10861) );
  AND2X1 U10869 ( .IN1(n9274), .IN2(n10207), .Q(n10860) );
  OR2X1 U10870 ( .IN1(n10863), .IN2(n10864), .Q(n10207) );
  INVX0 U10871 ( .INP(n10865), .ZN(n10864) );
  OR2X1 U10872 ( .IN1(n10866), .IN2(n10867), .Q(n10865) );
  AND2X1 U10873 ( .IN1(n10867), .IN2(n10866), .Q(n10863) );
  AND2X1 U10874 ( .IN1(n10868), .IN2(n10869), .Q(n10866) );
  OR2X1 U10875 ( .IN1(WX8519), .IN2(n8189), .Q(n10869) );
  INVX0 U10876 ( .INP(n10870), .ZN(n10868) );
  AND2X1 U10877 ( .IN1(n8189), .IN2(WX8519), .Q(n10870) );
  OR2X1 U10878 ( .IN1(n10871), .IN2(n10872), .Q(n10867) );
  AND2X1 U10879 ( .IN1(n8190), .IN2(WX8647), .Q(n10872) );
  AND2X1 U10880 ( .IN1(n8816), .IN2(WX8583), .Q(n10871) );
  AND2X1 U10881 ( .IN1(n9243), .IN2(CRC_OUT_4_5), .Q(n10859) );
  AND2X1 U10882 ( .IN1(n1256), .IN2(n9218), .Q(n10858) );
  INVX0 U10883 ( .INP(n10873), .ZN(n1256) );
  OR2X1 U10884 ( .IN1(n9572), .IN2(n3884), .Q(n10873) );
  OR4X1 U10885 ( .IN1(n10874), .IN2(n10875), .IN3(n10876), .IN4(n10877), .Q(
        WX7159) );
  AND2X1 U10886 ( .IN1(n10878), .IN2(n9175), .Q(n10877) );
  AND2X1 U10887 ( .IN1(n9274), .IN2(n10223), .Q(n10876) );
  OR2X1 U10888 ( .IN1(n10879), .IN2(n10880), .Q(n10223) );
  INVX0 U10889 ( .INP(n10881), .ZN(n10880) );
  OR2X1 U10890 ( .IN1(n10882), .IN2(n10883), .Q(n10881) );
  AND2X1 U10891 ( .IN1(n10883), .IN2(n10882), .Q(n10879) );
  AND2X1 U10892 ( .IN1(n10884), .IN2(n10885), .Q(n10882) );
  OR2X1 U10893 ( .IN1(WX8517), .IN2(n8191), .Q(n10885) );
  INVX0 U10894 ( .INP(n10886), .ZN(n10884) );
  AND2X1 U10895 ( .IN1(n8191), .IN2(WX8517), .Q(n10886) );
  OR2X1 U10896 ( .IN1(n10887), .IN2(n10888), .Q(n10883) );
  AND2X1 U10897 ( .IN1(n8192), .IN2(WX8645), .Q(n10888) );
  AND2X1 U10898 ( .IN1(n8815), .IN2(WX8581), .Q(n10887) );
  AND2X1 U10899 ( .IN1(n9243), .IN2(CRC_OUT_4_6), .Q(n10875) );
  AND2X1 U10900 ( .IN1(n1255), .IN2(n9218), .Q(n10874) );
  INVX0 U10901 ( .INP(n10889), .ZN(n1255) );
  OR2X1 U10902 ( .IN1(n9571), .IN2(n3885), .Q(n10889) );
  OR4X1 U10903 ( .IN1(n10890), .IN2(n10891), .IN3(n10892), .IN4(n10893), .Q(
        WX7157) );
  AND2X1 U10904 ( .IN1(n9181), .IN2(n10894), .Q(n10893) );
  AND2X1 U10905 ( .IN1(n9274), .IN2(n10239), .Q(n10892) );
  OR2X1 U10906 ( .IN1(n10895), .IN2(n10896), .Q(n10239) );
  INVX0 U10907 ( .INP(n10897), .ZN(n10896) );
  OR2X1 U10908 ( .IN1(n10898), .IN2(n10899), .Q(n10897) );
  AND2X1 U10909 ( .IN1(n10899), .IN2(n10898), .Q(n10895) );
  AND2X1 U10910 ( .IN1(n10900), .IN2(n10901), .Q(n10898) );
  OR2X1 U10911 ( .IN1(WX8515), .IN2(n8193), .Q(n10901) );
  INVX0 U10912 ( .INP(n10902), .ZN(n10900) );
  AND2X1 U10913 ( .IN1(n8193), .IN2(WX8515), .Q(n10902) );
  OR2X1 U10914 ( .IN1(n10903), .IN2(n10904), .Q(n10899) );
  AND2X1 U10915 ( .IN1(n8194), .IN2(WX8643), .Q(n10904) );
  AND2X1 U10916 ( .IN1(n8814), .IN2(WX8579), .Q(n10903) );
  AND2X1 U10917 ( .IN1(n9243), .IN2(CRC_OUT_4_7), .Q(n10891) );
  AND2X1 U10918 ( .IN1(n1254), .IN2(n9218), .Q(n10890) );
  INVX0 U10919 ( .INP(n10905), .ZN(n1254) );
  OR2X1 U10920 ( .IN1(n9571), .IN2(n3886), .Q(n10905) );
  OR4X1 U10921 ( .IN1(n10906), .IN2(n10907), .IN3(n10908), .IN4(n10909), .Q(
        WX7155) );
  AND2X1 U10922 ( .IN1(n10910), .IN2(n9174), .Q(n10909) );
  AND2X1 U10923 ( .IN1(n9274), .IN2(n10255), .Q(n10908) );
  OR2X1 U10924 ( .IN1(n10911), .IN2(n10912), .Q(n10255) );
  INVX0 U10925 ( .INP(n10913), .ZN(n10912) );
  OR2X1 U10926 ( .IN1(n10914), .IN2(n10915), .Q(n10913) );
  AND2X1 U10927 ( .IN1(n10915), .IN2(n10914), .Q(n10911) );
  AND2X1 U10928 ( .IN1(n10916), .IN2(n10917), .Q(n10914) );
  OR2X1 U10929 ( .IN1(WX8513), .IN2(n8195), .Q(n10917) );
  INVX0 U10930 ( .INP(n10918), .ZN(n10916) );
  AND2X1 U10931 ( .IN1(n8195), .IN2(WX8513), .Q(n10918) );
  OR2X1 U10932 ( .IN1(n10919), .IN2(n10920), .Q(n10915) );
  AND2X1 U10933 ( .IN1(n8196), .IN2(WX8641), .Q(n10920) );
  AND2X1 U10934 ( .IN1(n8813), .IN2(WX8577), .Q(n10919) );
  AND2X1 U10935 ( .IN1(n9243), .IN2(CRC_OUT_4_8), .Q(n10907) );
  AND2X1 U10936 ( .IN1(n1253), .IN2(n9218), .Q(n10906) );
  INVX0 U10937 ( .INP(n10921), .ZN(n1253) );
  OR2X1 U10938 ( .IN1(n9571), .IN2(n3887), .Q(n10921) );
  OR4X1 U10939 ( .IN1(n10922), .IN2(n10923), .IN3(n10924), .IN4(n10925), .Q(
        WX7153) );
  AND2X1 U10940 ( .IN1(n9181), .IN2(n10926), .Q(n10925) );
  AND2X1 U10941 ( .IN1(n10271), .IN2(n9259), .Q(n10924) );
  AND2X1 U10942 ( .IN1(n10927), .IN2(n10928), .Q(n10271) );
  INVX0 U10943 ( .INP(n10929), .ZN(n10928) );
  AND2X1 U10944 ( .IN1(n10930), .IN2(n10931), .Q(n10929) );
  OR2X1 U10945 ( .IN1(n10931), .IN2(n10930), .Q(n10927) );
  OR2X1 U10946 ( .IN1(n10932), .IN2(n10933), .Q(n10930) );
  INVX0 U10947 ( .INP(n10934), .ZN(n10933) );
  OR2X1 U10948 ( .IN1(WX8511), .IN2(n8197), .Q(n10934) );
  AND2X1 U10949 ( .IN1(n8197), .IN2(WX8511), .Q(n10932) );
  AND2X1 U10950 ( .IN1(n10935), .IN2(n10936), .Q(n10931) );
  OR2X1 U10951 ( .IN1(WX8575), .IN2(test_so75), .Q(n10936) );
  OR2X1 U10952 ( .IN1(n9099), .IN2(n8198), .Q(n10935) );
  AND2X1 U10953 ( .IN1(n9243), .IN2(CRC_OUT_4_9), .Q(n10923) );
  AND2X1 U10954 ( .IN1(n1252), .IN2(n9218), .Q(n10922) );
  INVX0 U10955 ( .INP(n10937), .ZN(n1252) );
  OR2X1 U10956 ( .IN1(n9571), .IN2(n3888), .Q(n10937) );
  OR4X1 U10957 ( .IN1(n10938), .IN2(n10939), .IN3(n10940), .IN4(n10941), .Q(
        WX7151) );
  AND2X1 U10958 ( .IN1(n10942), .IN2(n9174), .Q(n10941) );
  AND2X1 U10959 ( .IN1(n9274), .IN2(n10287), .Q(n10940) );
  OR2X1 U10960 ( .IN1(n10943), .IN2(n10944), .Q(n10287) );
  INVX0 U10961 ( .INP(n10945), .ZN(n10944) );
  OR2X1 U10962 ( .IN1(n10946), .IN2(n10947), .Q(n10945) );
  AND2X1 U10963 ( .IN1(n10947), .IN2(n10946), .Q(n10943) );
  AND2X1 U10964 ( .IN1(n10948), .IN2(n10949), .Q(n10946) );
  OR2X1 U10965 ( .IN1(WX8509), .IN2(n8199), .Q(n10949) );
  INVX0 U10966 ( .INP(n10950), .ZN(n10948) );
  AND2X1 U10967 ( .IN1(n8199), .IN2(WX8509), .Q(n10950) );
  OR2X1 U10968 ( .IN1(n10951), .IN2(n10952), .Q(n10947) );
  AND2X1 U10969 ( .IN1(n8200), .IN2(WX8637), .Q(n10952) );
  AND2X1 U10970 ( .IN1(n8812), .IN2(WX8573), .Q(n10951) );
  AND2X1 U10971 ( .IN1(n9243), .IN2(CRC_OUT_4_10), .Q(n10939) );
  AND2X1 U10972 ( .IN1(n1251), .IN2(n9218), .Q(n10938) );
  INVX0 U10973 ( .INP(n10953), .ZN(n1251) );
  OR2X1 U10974 ( .IN1(n9571), .IN2(n3889), .Q(n10953) );
  OR4X1 U10975 ( .IN1(n10954), .IN2(n10955), .IN3(n10956), .IN4(n10957), .Q(
        WX7149) );
  AND2X1 U10976 ( .IN1(n9181), .IN2(n10958), .Q(n10957) );
  AND2X1 U10977 ( .IN1(n10303), .IN2(n9259), .Q(n10956) );
  AND2X1 U10978 ( .IN1(n10959), .IN2(n10960), .Q(n10303) );
  INVX0 U10979 ( .INP(n10961), .ZN(n10960) );
  AND2X1 U10980 ( .IN1(n10962), .IN2(n10963), .Q(n10961) );
  OR2X1 U10981 ( .IN1(n10963), .IN2(n10962), .Q(n10959) );
  OR2X1 U10982 ( .IN1(n10964), .IN2(n10965), .Q(n10962) );
  INVX0 U10983 ( .INP(n10966), .ZN(n10965) );
  OR2X1 U10984 ( .IN1(WX8507), .IN2(n8201), .Q(n10966) );
  AND2X1 U10985 ( .IN1(n8201), .IN2(WX8507), .Q(n10964) );
  AND2X1 U10986 ( .IN1(n10967), .IN2(n10968), .Q(n10963) );
  OR2X1 U10987 ( .IN1(WX8635), .IN2(test_so73), .Q(n10968) );
  OR2X1 U10988 ( .IN1(n9115), .IN2(n8720), .Q(n10967) );
  AND2X1 U10989 ( .IN1(n9244), .IN2(CRC_OUT_4_11), .Q(n10955) );
  AND2X1 U10990 ( .IN1(n1250), .IN2(n9218), .Q(n10954) );
  INVX0 U10991 ( .INP(n10969), .ZN(n1250) );
  OR2X1 U10992 ( .IN1(n9571), .IN2(n3890), .Q(n10969) );
  OR4X1 U10993 ( .IN1(n10970), .IN2(n10971), .IN3(n10972), .IN4(n10973), .Q(
        WX7147) );
  AND2X1 U10994 ( .IN1(n9181), .IN2(n10974), .Q(n10973) );
  AND2X1 U10995 ( .IN1(n9274), .IN2(n10319), .Q(n10972) );
  OR2X1 U10996 ( .IN1(n10975), .IN2(n10976), .Q(n10319) );
  INVX0 U10997 ( .INP(n10977), .ZN(n10976) );
  OR2X1 U10998 ( .IN1(n10978), .IN2(n10979), .Q(n10977) );
  AND2X1 U10999 ( .IN1(n10979), .IN2(n10978), .Q(n10975) );
  AND2X1 U11000 ( .IN1(n10980), .IN2(n10981), .Q(n10978) );
  OR2X1 U11001 ( .IN1(WX8505), .IN2(n8202), .Q(n10981) );
  INVX0 U11002 ( .INP(n10982), .ZN(n10980) );
  AND2X1 U11003 ( .IN1(n8202), .IN2(WX8505), .Q(n10982) );
  OR2X1 U11004 ( .IN1(n10983), .IN2(n10984), .Q(n10979) );
  AND2X1 U11005 ( .IN1(n8203), .IN2(WX8633), .Q(n10984) );
  AND2X1 U11006 ( .IN1(n8811), .IN2(WX8569), .Q(n10983) );
  AND2X1 U11007 ( .IN1(test_so65), .IN2(n9227), .Q(n10971) );
  AND2X1 U11008 ( .IN1(n1249), .IN2(n9218), .Q(n10970) );
  INVX0 U11009 ( .INP(n10985), .ZN(n1249) );
  OR2X1 U11010 ( .IN1(n9571), .IN2(n3891), .Q(n10985) );
  OR4X1 U11011 ( .IN1(n10986), .IN2(n10987), .IN3(n10988), .IN4(n10989), .Q(
        WX7145) );
  AND2X1 U11012 ( .IN1(n9181), .IN2(n10990), .Q(n10989) );
  AND2X1 U11013 ( .IN1(n10335), .IN2(n9259), .Q(n10988) );
  AND2X1 U11014 ( .IN1(n10991), .IN2(n10992), .Q(n10335) );
  INVX0 U11015 ( .INP(n10993), .ZN(n10992) );
  AND2X1 U11016 ( .IN1(n10994), .IN2(n10995), .Q(n10993) );
  OR2X1 U11017 ( .IN1(n10995), .IN2(n10994), .Q(n10991) );
  OR2X1 U11018 ( .IN1(n10996), .IN2(n10997), .Q(n10994) );
  INVX0 U11019 ( .INP(n10998), .ZN(n10997) );
  OR2X1 U11020 ( .IN1(WX8439), .IN2(n8205), .Q(n10998) );
  AND2X1 U11021 ( .IN1(n8205), .IN2(WX8439), .Q(n10996) );
  AND2X1 U11022 ( .IN1(n10999), .IN2(n11000), .Q(n10995) );
  OR2X1 U11023 ( .IN1(WX8631), .IN2(test_so71), .Q(n11000) );
  OR2X1 U11024 ( .IN1(n9116), .IN2(n8810), .Q(n10999) );
  AND2X1 U11025 ( .IN1(n9244), .IN2(CRC_OUT_4_13), .Q(n10987) );
  AND2X1 U11026 ( .IN1(n1248), .IN2(n9218), .Q(n10986) );
  INVX0 U11027 ( .INP(n11001), .ZN(n1248) );
  OR2X1 U11028 ( .IN1(n9571), .IN2(n3892), .Q(n11001) );
  OR4X1 U11029 ( .IN1(n11002), .IN2(n11003), .IN3(n11004), .IN4(n11005), .Q(
        WX7143) );
  AND2X1 U11030 ( .IN1(n9178), .IN2(n11006), .Q(n11005) );
  AND2X1 U11031 ( .IN1(n9274), .IN2(n10351), .Q(n11004) );
  OR2X1 U11032 ( .IN1(n11007), .IN2(n11008), .Q(n10351) );
  INVX0 U11033 ( .INP(n11009), .ZN(n11008) );
  OR2X1 U11034 ( .IN1(n11010), .IN2(n11011), .Q(n11009) );
  AND2X1 U11035 ( .IN1(n11011), .IN2(n11010), .Q(n11007) );
  AND2X1 U11036 ( .IN1(n11012), .IN2(n11013), .Q(n11010) );
  OR2X1 U11037 ( .IN1(WX8501), .IN2(n8206), .Q(n11013) );
  INVX0 U11038 ( .INP(n11014), .ZN(n11012) );
  AND2X1 U11039 ( .IN1(n8206), .IN2(WX8501), .Q(n11014) );
  OR2X1 U11040 ( .IN1(n11015), .IN2(n11016), .Q(n11011) );
  AND2X1 U11041 ( .IN1(n8207), .IN2(WX8629), .Q(n11016) );
  AND2X1 U11042 ( .IN1(n8809), .IN2(WX8565), .Q(n11015) );
  AND2X1 U11043 ( .IN1(n9244), .IN2(CRC_OUT_4_14), .Q(n11003) );
  AND2X1 U11044 ( .IN1(n1247), .IN2(n9218), .Q(n11002) );
  INVX0 U11045 ( .INP(n11017), .ZN(n1247) );
  OR2X1 U11046 ( .IN1(n9571), .IN2(n3893), .Q(n11017) );
  OR4X1 U11047 ( .IN1(n11018), .IN2(n11019), .IN3(n11020), .IN4(n11021), .Q(
        WX7141) );
  AND2X1 U11048 ( .IN1(n9178), .IN2(n11022), .Q(n11021) );
  AND2X1 U11049 ( .IN1(n10367), .IN2(n9259), .Q(n11020) );
  AND2X1 U11050 ( .IN1(n11023), .IN2(n11024), .Q(n10367) );
  INVX0 U11051 ( .INP(n11025), .ZN(n11024) );
  AND2X1 U11052 ( .IN1(n11026), .IN2(n11027), .Q(n11025) );
  OR2X1 U11053 ( .IN1(n11027), .IN2(n11026), .Q(n11023) );
  OR2X1 U11054 ( .IN1(n11028), .IN2(n11029), .Q(n11026) );
  INVX0 U11055 ( .INP(n11030), .ZN(n11029) );
  OR2X1 U11056 ( .IN1(WX8499), .IN2(n8208), .Q(n11030) );
  AND2X1 U11057 ( .IN1(n8208), .IN2(WX8499), .Q(n11028) );
  AND2X1 U11058 ( .IN1(n11031), .IN2(n11032), .Q(n11027) );
  OR2X1 U11059 ( .IN1(WX8627), .IN2(test_so69), .Q(n11032) );
  OR2X1 U11060 ( .IN1(n9117), .IN2(n8808), .Q(n11031) );
  AND2X1 U11061 ( .IN1(n9244), .IN2(CRC_OUT_4_15), .Q(n11019) );
  AND2X1 U11062 ( .IN1(n1246), .IN2(n9219), .Q(n11018) );
  INVX0 U11063 ( .INP(n11033), .ZN(n1246) );
  OR2X1 U11064 ( .IN1(n9571), .IN2(n3894), .Q(n11033) );
  OR4X1 U11065 ( .IN1(n11034), .IN2(n11035), .IN3(n11036), .IN4(n11037), .Q(
        WX7139) );
  AND2X1 U11066 ( .IN1(n9178), .IN2(n11038), .Q(n11037) );
  AND2X1 U11067 ( .IN1(n9274), .IN2(n10383), .Q(n11036) );
  OR2X1 U11068 ( .IN1(n11039), .IN2(n11040), .Q(n10383) );
  INVX0 U11069 ( .INP(n11041), .ZN(n11040) );
  OR2X1 U11070 ( .IN1(n11042), .IN2(n11043), .Q(n11041) );
  AND2X1 U11071 ( .IN1(n11043), .IN2(n11042), .Q(n11039) );
  AND2X1 U11072 ( .IN1(n11044), .IN2(n11045), .Q(n11042) );
  OR2X1 U11073 ( .IN1(n9471), .IN2(n7948), .Q(n11045) );
  OR2X1 U11074 ( .IN1(WX8497), .IN2(n9449), .Q(n11044) );
  OR2X1 U11075 ( .IN1(n11046), .IN2(n11047), .Q(n11043) );
  INVX0 U11076 ( .INP(n11048), .ZN(n11047) );
  OR2X1 U11077 ( .IN1(n11049), .IN2(n7949), .Q(n11048) );
  AND2X1 U11078 ( .IN1(n7949), .IN2(n11049), .Q(n11046) );
  INVX0 U11079 ( .INP(n11050), .ZN(n11049) );
  OR2X1 U11080 ( .IN1(n11051), .IN2(n11052), .Q(n11050) );
  AND2X1 U11081 ( .IN1(n8719), .IN2(n8363), .Q(n11052) );
  AND2X1 U11082 ( .IN1(n15892), .IN2(WX8625), .Q(n11051) );
  AND2X1 U11083 ( .IN1(n9244), .IN2(CRC_OUT_4_16), .Q(n11035) );
  AND2X1 U11084 ( .IN1(n1245), .IN2(n9219), .Q(n11034) );
  INVX0 U11085 ( .INP(n11053), .ZN(n1245) );
  OR2X1 U11086 ( .IN1(n9571), .IN2(n3895), .Q(n11053) );
  OR4X1 U11087 ( .IN1(n11054), .IN2(n11055), .IN3(n11056), .IN4(n11057), .Q(
        WX7137) );
  AND2X1 U11088 ( .IN1(n9178), .IN2(n11058), .Q(n11057) );
  AND2X1 U11089 ( .IN1(n9274), .IN2(n10402), .Q(n11056) );
  OR2X1 U11090 ( .IN1(n11059), .IN2(n11060), .Q(n10402) );
  INVX0 U11091 ( .INP(n11061), .ZN(n11060) );
  OR2X1 U11092 ( .IN1(n11062), .IN2(n11063), .Q(n11061) );
  AND2X1 U11093 ( .IN1(n11063), .IN2(n11062), .Q(n11059) );
  AND2X1 U11094 ( .IN1(n11064), .IN2(n11065), .Q(n11062) );
  OR2X1 U11095 ( .IN1(n9466), .IN2(n7950), .Q(n11065) );
  OR2X1 U11096 ( .IN1(WX8495), .IN2(n9448), .Q(n11064) );
  OR2X1 U11097 ( .IN1(n11066), .IN2(n11067), .Q(n11063) );
  INVX0 U11098 ( .INP(n11068), .ZN(n11067) );
  OR2X1 U11099 ( .IN1(n11069), .IN2(n7951), .Q(n11068) );
  AND2X1 U11100 ( .IN1(n7951), .IN2(n11069), .Q(n11066) );
  INVX0 U11101 ( .INP(n11070), .ZN(n11069) );
  OR2X1 U11102 ( .IN1(n11071), .IN2(n11072), .Q(n11070) );
  AND2X1 U11103 ( .IN1(n8807), .IN2(n8364), .Q(n11072) );
  AND2X1 U11104 ( .IN1(n15893), .IN2(WX8623), .Q(n11071) );
  AND2X1 U11105 ( .IN1(n9244), .IN2(CRC_OUT_4_17), .Q(n11055) );
  AND2X1 U11106 ( .IN1(n1244), .IN2(n9219), .Q(n11054) );
  INVX0 U11107 ( .INP(n11073), .ZN(n1244) );
  OR2X1 U11108 ( .IN1(n9571), .IN2(n3896), .Q(n11073) );
  OR4X1 U11109 ( .IN1(n11074), .IN2(n11075), .IN3(n11076), .IN4(n11077), .Q(
        WX7135) );
  AND2X1 U11110 ( .IN1(n9178), .IN2(n11078), .Q(n11077) );
  AND2X1 U11111 ( .IN1(n9274), .IN2(n10422), .Q(n11076) );
  OR2X1 U11112 ( .IN1(n11079), .IN2(n11080), .Q(n10422) );
  INVX0 U11113 ( .INP(n11081), .ZN(n11080) );
  OR2X1 U11114 ( .IN1(n11082), .IN2(n11083), .Q(n11081) );
  AND2X1 U11115 ( .IN1(n11083), .IN2(n11082), .Q(n11079) );
  AND2X1 U11116 ( .IN1(n11084), .IN2(n11085), .Q(n11082) );
  OR2X1 U11117 ( .IN1(n9478), .IN2(n7952), .Q(n11085) );
  OR2X1 U11118 ( .IN1(WX8493), .IN2(n9449), .Q(n11084) );
  OR2X1 U11119 ( .IN1(n11086), .IN2(n11087), .Q(n11083) );
  INVX0 U11120 ( .INP(n11088), .ZN(n11087) );
  OR2X1 U11121 ( .IN1(n11089), .IN2(n7953), .Q(n11088) );
  AND2X1 U11122 ( .IN1(n7953), .IN2(n11089), .Q(n11086) );
  INVX0 U11123 ( .INP(n11090), .ZN(n11089) );
  OR2X1 U11124 ( .IN1(n11091), .IN2(n11092), .Q(n11090) );
  AND2X1 U11125 ( .IN1(n8806), .IN2(n8365), .Q(n11092) );
  AND2X1 U11126 ( .IN1(n15894), .IN2(WX8621), .Q(n11091) );
  AND2X1 U11127 ( .IN1(n9244), .IN2(CRC_OUT_4_18), .Q(n11075) );
  AND2X1 U11128 ( .IN1(n1243), .IN2(n9219), .Q(n11074) );
  INVX0 U11129 ( .INP(n11093), .ZN(n1243) );
  OR2X1 U11130 ( .IN1(n9570), .IN2(n3897), .Q(n11093) );
  OR4X1 U11131 ( .IN1(n11094), .IN2(n11095), .IN3(n11096), .IN4(n11097), .Q(
        WX7133) );
  AND2X1 U11132 ( .IN1(n9179), .IN2(n11098), .Q(n11097) );
  AND2X1 U11133 ( .IN1(n9275), .IN2(n10441), .Q(n11096) );
  OR2X1 U11134 ( .IN1(n11099), .IN2(n11100), .Q(n10441) );
  INVX0 U11135 ( .INP(n11101), .ZN(n11100) );
  OR2X1 U11136 ( .IN1(n11102), .IN2(n11103), .Q(n11101) );
  AND2X1 U11137 ( .IN1(n11103), .IN2(n11102), .Q(n11099) );
  AND2X1 U11138 ( .IN1(n11104), .IN2(n11105), .Q(n11102) );
  OR2X1 U11139 ( .IN1(n9477), .IN2(n7954), .Q(n11105) );
  OR2X1 U11140 ( .IN1(WX8491), .IN2(n9449), .Q(n11104) );
  OR2X1 U11141 ( .IN1(n11106), .IN2(n11107), .Q(n11103) );
  INVX0 U11142 ( .INP(n11108), .ZN(n11107) );
  OR2X1 U11143 ( .IN1(n11109), .IN2(n7955), .Q(n11108) );
  AND2X1 U11144 ( .IN1(n7955), .IN2(n11109), .Q(n11106) );
  INVX0 U11145 ( .INP(n11110), .ZN(n11109) );
  OR2X1 U11146 ( .IN1(n11111), .IN2(n11112), .Q(n11110) );
  AND2X1 U11147 ( .IN1(n8805), .IN2(n8366), .Q(n11112) );
  AND2X1 U11148 ( .IN1(n15895), .IN2(WX8619), .Q(n11111) );
  AND2X1 U11149 ( .IN1(n9244), .IN2(CRC_OUT_4_19), .Q(n11095) );
  AND2X1 U11150 ( .IN1(n1242), .IN2(n9219), .Q(n11094) );
  INVX0 U11151 ( .INP(n11113), .ZN(n1242) );
  OR2X1 U11152 ( .IN1(n9570), .IN2(n3898), .Q(n11113) );
  OR4X1 U11153 ( .IN1(n11114), .IN2(n11115), .IN3(n11116), .IN4(n11117), .Q(
        WX7131) );
  AND2X1 U11154 ( .IN1(n9178), .IN2(n11118), .Q(n11117) );
  AND2X1 U11155 ( .IN1(n9275), .IN2(n10461), .Q(n11116) );
  OR2X1 U11156 ( .IN1(n11119), .IN2(n11120), .Q(n10461) );
  INVX0 U11157 ( .INP(n11121), .ZN(n11120) );
  OR2X1 U11158 ( .IN1(n11122), .IN2(n11123), .Q(n11121) );
  AND2X1 U11159 ( .IN1(n11123), .IN2(n11122), .Q(n11119) );
  AND2X1 U11160 ( .IN1(n11124), .IN2(n11125), .Q(n11122) );
  OR2X1 U11161 ( .IN1(n9476), .IN2(n7956), .Q(n11125) );
  OR2X1 U11162 ( .IN1(WX8489), .IN2(n9449), .Q(n11124) );
  OR2X1 U11163 ( .IN1(n11126), .IN2(n11127), .Q(n11123) );
  INVX0 U11164 ( .INP(n11128), .ZN(n11127) );
  OR2X1 U11165 ( .IN1(n11129), .IN2(n7957), .Q(n11128) );
  AND2X1 U11166 ( .IN1(n7957), .IN2(n11129), .Q(n11126) );
  INVX0 U11167 ( .INP(n11130), .ZN(n11129) );
  OR2X1 U11168 ( .IN1(n11131), .IN2(n11132), .Q(n11130) );
  AND2X1 U11169 ( .IN1(n8804), .IN2(n8367), .Q(n11132) );
  AND2X1 U11170 ( .IN1(n15896), .IN2(WX8617), .Q(n11131) );
  AND2X1 U11171 ( .IN1(n9244), .IN2(CRC_OUT_4_20), .Q(n11115) );
  AND2X1 U11172 ( .IN1(n1241), .IN2(n9219), .Q(n11114) );
  INVX0 U11173 ( .INP(n11133), .ZN(n1241) );
  OR2X1 U11174 ( .IN1(n9570), .IN2(n3899), .Q(n11133) );
  OR4X1 U11175 ( .IN1(n11134), .IN2(n11135), .IN3(n11136), .IN4(n11137), .Q(
        WX7129) );
  AND2X1 U11176 ( .IN1(n11138), .IN2(n9176), .Q(n11137) );
  AND2X1 U11177 ( .IN1(n9275), .IN2(n10482), .Q(n11136) );
  OR2X1 U11178 ( .IN1(n11139), .IN2(n11140), .Q(n10482) );
  INVX0 U11179 ( .INP(n11141), .ZN(n11140) );
  OR2X1 U11180 ( .IN1(n11142), .IN2(n11143), .Q(n11141) );
  AND2X1 U11181 ( .IN1(n11143), .IN2(n11142), .Q(n11139) );
  AND2X1 U11182 ( .IN1(n11144), .IN2(n11145), .Q(n11142) );
  OR2X1 U11183 ( .IN1(n9475), .IN2(n7958), .Q(n11145) );
  OR2X1 U11184 ( .IN1(WX8487), .IN2(n9447), .Q(n11144) );
  OR2X1 U11185 ( .IN1(n11146), .IN2(n11147), .Q(n11143) );
  INVX0 U11186 ( .INP(n11148), .ZN(n11147) );
  OR2X1 U11187 ( .IN1(n11149), .IN2(n7959), .Q(n11148) );
  AND2X1 U11188 ( .IN1(n7959), .IN2(n11149), .Q(n11146) );
  INVX0 U11189 ( .INP(n11150), .ZN(n11149) );
  OR2X1 U11190 ( .IN1(n11151), .IN2(n11152), .Q(n11150) );
  AND2X1 U11191 ( .IN1(n8803), .IN2(n8368), .Q(n11152) );
  AND2X1 U11192 ( .IN1(n15897), .IN2(WX8615), .Q(n11151) );
  AND2X1 U11193 ( .IN1(n9244), .IN2(CRC_OUT_4_21), .Q(n11135) );
  AND2X1 U11194 ( .IN1(n1240), .IN2(n9219), .Q(n11134) );
  INVX0 U11195 ( .INP(n11153), .ZN(n1240) );
  OR2X1 U11196 ( .IN1(n9570), .IN2(n3900), .Q(n11153) );
  OR4X1 U11197 ( .IN1(n11154), .IN2(n11155), .IN3(n11156), .IN4(n11157), .Q(
        WX7127) );
  AND2X1 U11198 ( .IN1(n9178), .IN2(n11158), .Q(n11157) );
  AND2X1 U11199 ( .IN1(n9275), .IN2(n10502), .Q(n11156) );
  OR2X1 U11200 ( .IN1(n11159), .IN2(n11160), .Q(n10502) );
  INVX0 U11201 ( .INP(n11161), .ZN(n11160) );
  OR2X1 U11202 ( .IN1(n11162), .IN2(n11163), .Q(n11161) );
  AND2X1 U11203 ( .IN1(n11163), .IN2(n11162), .Q(n11159) );
  AND2X1 U11204 ( .IN1(n11164), .IN2(n11165), .Q(n11162) );
  OR2X1 U11205 ( .IN1(n9472), .IN2(n7960), .Q(n11165) );
  OR2X1 U11206 ( .IN1(WX8485), .IN2(n9449), .Q(n11164) );
  OR2X1 U11207 ( .IN1(n11166), .IN2(n11167), .Q(n11163) );
  INVX0 U11208 ( .INP(n11168), .ZN(n11167) );
  OR2X1 U11209 ( .IN1(n11169), .IN2(n7961), .Q(n11168) );
  AND2X1 U11210 ( .IN1(n7961), .IN2(n11169), .Q(n11166) );
  INVX0 U11211 ( .INP(n11170), .ZN(n11169) );
  OR2X1 U11212 ( .IN1(n11171), .IN2(n11172), .Q(n11170) );
  AND2X1 U11213 ( .IN1(n8802), .IN2(n8369), .Q(n11172) );
  AND2X1 U11214 ( .IN1(n15898), .IN2(WX8613), .Q(n11171) );
  AND2X1 U11215 ( .IN1(n9244), .IN2(CRC_OUT_4_22), .Q(n11155) );
  AND2X1 U11216 ( .IN1(n1239), .IN2(n9219), .Q(n11154) );
  INVX0 U11217 ( .INP(n11173), .ZN(n1239) );
  OR2X1 U11218 ( .IN1(n9570), .IN2(n3901), .Q(n11173) );
  OR4X1 U11219 ( .IN1(n11174), .IN2(n11175), .IN3(n11176), .IN4(n11177), .Q(
        WX7125) );
  AND2X1 U11220 ( .IN1(n11178), .IN2(n9177), .Q(n11177) );
  AND2X1 U11221 ( .IN1(n9275), .IN2(n10522), .Q(n11176) );
  OR2X1 U11222 ( .IN1(n11179), .IN2(n11180), .Q(n10522) );
  INVX0 U11223 ( .INP(n11181), .ZN(n11180) );
  OR2X1 U11224 ( .IN1(n11182), .IN2(n11183), .Q(n11181) );
  AND2X1 U11225 ( .IN1(n11183), .IN2(n11182), .Q(n11179) );
  AND2X1 U11226 ( .IN1(n11184), .IN2(n11185), .Q(n11182) );
  OR2X1 U11227 ( .IN1(n9470), .IN2(n7962), .Q(n11185) );
  OR2X1 U11228 ( .IN1(WX8483), .IN2(n9449), .Q(n11184) );
  OR2X1 U11229 ( .IN1(n11186), .IN2(n11187), .Q(n11183) );
  INVX0 U11230 ( .INP(n11188), .ZN(n11187) );
  OR2X1 U11231 ( .IN1(n11189), .IN2(n7963), .Q(n11188) );
  AND2X1 U11232 ( .IN1(n7963), .IN2(n11189), .Q(n11186) );
  INVX0 U11233 ( .INP(n11190), .ZN(n11189) );
  OR2X1 U11234 ( .IN1(n11191), .IN2(n11192), .Q(n11190) );
  AND2X1 U11235 ( .IN1(n8801), .IN2(n8370), .Q(n11192) );
  AND2X1 U11236 ( .IN1(n15899), .IN2(WX8611), .Q(n11191) );
  AND2X1 U11237 ( .IN1(n9244), .IN2(CRC_OUT_4_23), .Q(n11175) );
  AND2X1 U11238 ( .IN1(n1238), .IN2(n9219), .Q(n11174) );
  INVX0 U11239 ( .INP(n11193), .ZN(n1238) );
  OR2X1 U11240 ( .IN1(n9570), .IN2(n3902), .Q(n11193) );
  OR4X1 U11241 ( .IN1(n11194), .IN2(n11195), .IN3(n11196), .IN4(n11197), .Q(
        WX7123) );
  AND2X1 U11242 ( .IN1(n9178), .IN2(n11198), .Q(n11197) );
  AND2X1 U11243 ( .IN1(n9275), .IN2(n10542), .Q(n11196) );
  OR2X1 U11244 ( .IN1(n11199), .IN2(n11200), .Q(n10542) );
  INVX0 U11245 ( .INP(n11201), .ZN(n11200) );
  OR2X1 U11246 ( .IN1(n11202), .IN2(n11203), .Q(n11201) );
  AND2X1 U11247 ( .IN1(n11203), .IN2(n11202), .Q(n11199) );
  AND2X1 U11248 ( .IN1(n11204), .IN2(n11205), .Q(n11202) );
  OR2X1 U11249 ( .IN1(n9470), .IN2(n7964), .Q(n11205) );
  OR2X1 U11250 ( .IN1(WX8481), .IN2(n9447), .Q(n11204) );
  OR2X1 U11251 ( .IN1(n11206), .IN2(n11207), .Q(n11203) );
  INVX0 U11252 ( .INP(n11208), .ZN(n11207) );
  OR2X1 U11253 ( .IN1(n11209), .IN2(n7965), .Q(n11208) );
  AND2X1 U11254 ( .IN1(n7965), .IN2(n11209), .Q(n11206) );
  INVX0 U11255 ( .INP(n11210), .ZN(n11209) );
  OR2X1 U11256 ( .IN1(n11211), .IN2(n11212), .Q(n11210) );
  AND2X1 U11257 ( .IN1(n8800), .IN2(n8371), .Q(n11212) );
  AND2X1 U11258 ( .IN1(n15900), .IN2(WX8609), .Q(n11211) );
  AND2X1 U11259 ( .IN1(n9244), .IN2(CRC_OUT_4_24), .Q(n11195) );
  AND2X1 U11260 ( .IN1(n1237), .IN2(n9219), .Q(n11194) );
  INVX0 U11261 ( .INP(n11213), .ZN(n1237) );
  OR2X1 U11262 ( .IN1(n9570), .IN2(n3903), .Q(n11213) );
  OR4X1 U11263 ( .IN1(n11214), .IN2(n11215), .IN3(n11216), .IN4(n11217), .Q(
        WX7121) );
  AND2X1 U11264 ( .IN1(n11218), .IN2(n9177), .Q(n11217) );
  AND2X1 U11265 ( .IN1(n9275), .IN2(n10562), .Q(n11216) );
  OR2X1 U11266 ( .IN1(n11219), .IN2(n11220), .Q(n10562) );
  AND2X1 U11267 ( .IN1(n11221), .IN2(n11222), .Q(n11220) );
  INVX0 U11268 ( .INP(n11223), .ZN(n11222) );
  AND2X1 U11269 ( .IN1(n11223), .IN2(n11224), .Q(n11219) );
  INVX0 U11270 ( .INP(n11221), .ZN(n11224) );
  OR2X1 U11271 ( .IN1(n11225), .IN2(n11226), .Q(n11221) );
  AND2X1 U11272 ( .IN1(n9451), .IN2(n8372), .Q(n11226) );
  AND2X1 U11273 ( .IN1(n15901), .IN2(n9469), .Q(n11225) );
  OR2X1 U11274 ( .IN1(n11227), .IN2(n11228), .Q(n11223) );
  AND3X1 U11275 ( .IN1(n11229), .IN2(n11230), .IN3(n8799), .Q(n11228) );
  OR2X1 U11276 ( .IN1(n7966), .IN2(WX8543), .Q(n11230) );
  OR2X1 U11277 ( .IN1(n7967), .IN2(WX8479), .Q(n11229) );
  AND2X1 U11278 ( .IN1(n11231), .IN2(WX8607), .Q(n11227) );
  OR2X1 U11279 ( .IN1(n11232), .IN2(n11233), .Q(n11231) );
  AND2X1 U11280 ( .IN1(n7966), .IN2(WX8543), .Q(n11233) );
  AND2X1 U11281 ( .IN1(n7967), .IN2(WX8479), .Q(n11232) );
  AND2X1 U11282 ( .IN1(n9245), .IN2(CRC_OUT_4_25), .Q(n11215) );
  AND2X1 U11283 ( .IN1(n1236), .IN2(n9219), .Q(n11214) );
  INVX0 U11284 ( .INP(n11234), .ZN(n1236) );
  OR2X1 U11285 ( .IN1(n9570), .IN2(n3904), .Q(n11234) );
  OR4X1 U11286 ( .IN1(n11235), .IN2(n11236), .IN3(n11237), .IN4(n11238), .Q(
        WX7119) );
  AND2X1 U11287 ( .IN1(n9179), .IN2(n11239), .Q(n11238) );
  AND2X1 U11288 ( .IN1(n10582), .IN2(n9259), .Q(n11237) );
  AND2X1 U11289 ( .IN1(n11240), .IN2(n11241), .Q(n10582) );
  INVX0 U11290 ( .INP(n11242), .ZN(n11241) );
  AND2X1 U11291 ( .IN1(n11243), .IN2(n11244), .Q(n11242) );
  OR2X1 U11292 ( .IN1(n11244), .IN2(n11243), .Q(n11240) );
  OR2X1 U11293 ( .IN1(n11245), .IN2(n11246), .Q(n11243) );
  AND2X1 U11294 ( .IN1(n9450), .IN2(WX8477), .Q(n11246) );
  AND2X1 U11295 ( .IN1(n7968), .IN2(n9477), .Q(n11245) );
  AND2X1 U11296 ( .IN1(n11247), .IN2(n11248), .Q(n11244) );
  OR2X1 U11297 ( .IN1(n11249), .IN2(n7969), .Q(n11248) );
  INVX0 U11298 ( .INP(n11250), .ZN(n11249) );
  OR2X1 U11299 ( .IN1(WX8541), .IN2(n11250), .Q(n11247) );
  OR2X1 U11300 ( .IN1(n11251), .IN2(n11252), .Q(n11250) );
  AND2X1 U11301 ( .IN1(n15902), .IN2(n9104), .Q(n11252) );
  AND2X1 U11302 ( .IN1(test_so74), .IN2(n8373), .Q(n11251) );
  AND2X1 U11303 ( .IN1(n9245), .IN2(CRC_OUT_4_26), .Q(n11236) );
  AND2X1 U11304 ( .IN1(n1235), .IN2(n9219), .Q(n11235) );
  INVX0 U11305 ( .INP(n11253), .ZN(n1235) );
  OR2X1 U11306 ( .IN1(n9570), .IN2(n3905), .Q(n11253) );
  OR4X1 U11307 ( .IN1(n11254), .IN2(n11255), .IN3(n11256), .IN4(n11257), .Q(
        WX7117) );
  AND2X1 U11308 ( .IN1(n11258), .IN2(n9178), .Q(n11257) );
  AND2X1 U11309 ( .IN1(n9275), .IN2(n10602), .Q(n11256) );
  OR2X1 U11310 ( .IN1(n11259), .IN2(n11260), .Q(n10602) );
  INVX0 U11311 ( .INP(n11261), .ZN(n11260) );
  OR2X1 U11312 ( .IN1(n11262), .IN2(n11263), .Q(n11261) );
  AND2X1 U11313 ( .IN1(n11263), .IN2(n11262), .Q(n11259) );
  AND2X1 U11314 ( .IN1(n11264), .IN2(n11265), .Q(n11262) );
  OR2X1 U11315 ( .IN1(n9467), .IN2(n7970), .Q(n11265) );
  OR2X1 U11316 ( .IN1(WX8475), .IN2(n9448), .Q(n11264) );
  OR2X1 U11317 ( .IN1(n11266), .IN2(n11267), .Q(n11263) );
  INVX0 U11318 ( .INP(n11268), .ZN(n11267) );
  OR2X1 U11319 ( .IN1(n11269), .IN2(n7971), .Q(n11268) );
  AND2X1 U11320 ( .IN1(n7971), .IN2(n11269), .Q(n11266) );
  INVX0 U11321 ( .INP(n11270), .ZN(n11269) );
  OR2X1 U11322 ( .IN1(n11271), .IN2(n11272), .Q(n11270) );
  AND2X1 U11323 ( .IN1(n8798), .IN2(n8374), .Q(n11272) );
  AND2X1 U11324 ( .IN1(n15903), .IN2(WX8603), .Q(n11271) );
  AND2X1 U11325 ( .IN1(n9245), .IN2(CRC_OUT_4_27), .Q(n11255) );
  AND2X1 U11326 ( .IN1(n1234), .IN2(n9220), .Q(n11254) );
  INVX0 U11327 ( .INP(n11273), .ZN(n1234) );
  OR2X1 U11328 ( .IN1(n9570), .IN2(n3906), .Q(n11273) );
  OR4X1 U11329 ( .IN1(n11274), .IN2(n11275), .IN3(n11276), .IN4(n11277), .Q(
        WX7115) );
  AND2X1 U11330 ( .IN1(n9179), .IN2(n11278), .Q(n11277) );
  AND2X1 U11331 ( .IN1(n10622), .IN2(n9259), .Q(n11276) );
  AND2X1 U11332 ( .IN1(n11279), .IN2(n11280), .Q(n10622) );
  INVX0 U11333 ( .INP(n11281), .ZN(n11280) );
  AND2X1 U11334 ( .IN1(n11282), .IN2(n11283), .Q(n11281) );
  OR2X1 U11335 ( .IN1(n11283), .IN2(n11282), .Q(n11279) );
  OR2X1 U11336 ( .IN1(n11284), .IN2(n11285), .Q(n11282) );
  AND2X1 U11337 ( .IN1(n9451), .IN2(WX8473), .Q(n11285) );
  AND2X1 U11338 ( .IN1(n7972), .IN2(n9455), .Q(n11284) );
  AND2X1 U11339 ( .IN1(n11286), .IN2(n11287), .Q(n11283) );
  OR2X1 U11340 ( .IN1(n11288), .IN2(n8797), .Q(n11287) );
  OR2X1 U11341 ( .IN1(WX8601), .IN2(n11289), .Q(n11286) );
  INVX0 U11342 ( .INP(n11288), .ZN(n11289) );
  AND2X1 U11343 ( .IN1(n11290), .IN2(n11291), .Q(n11288) );
  OR2X1 U11344 ( .IN1(n8375), .IN2(test_so72), .Q(n11291) );
  OR2X1 U11345 ( .IN1(n9118), .IN2(n15904), .Q(n11290) );
  AND2X1 U11346 ( .IN1(n9245), .IN2(CRC_OUT_4_28), .Q(n11275) );
  AND2X1 U11347 ( .IN1(n1233), .IN2(n9220), .Q(n11274) );
  INVX0 U11348 ( .INP(n11292), .ZN(n1233) );
  OR2X1 U11349 ( .IN1(n9570), .IN2(n3907), .Q(n11292) );
  OR4X1 U11350 ( .IN1(n11293), .IN2(n11294), .IN3(n11295), .IN4(n11296), .Q(
        WX7113) );
  AND2X1 U11351 ( .IN1(n9179), .IN2(n11297), .Q(n11296) );
  AND2X1 U11352 ( .IN1(n9275), .IN2(n10642), .Q(n11295) );
  OR2X1 U11353 ( .IN1(n11298), .IN2(n11299), .Q(n10642) );
  INVX0 U11354 ( .INP(n11300), .ZN(n11299) );
  OR2X1 U11355 ( .IN1(n11301), .IN2(n11302), .Q(n11300) );
  AND2X1 U11356 ( .IN1(n11302), .IN2(n11301), .Q(n11298) );
  AND2X1 U11357 ( .IN1(n11303), .IN2(n11304), .Q(n11301) );
  OR2X1 U11358 ( .IN1(n9465), .IN2(n7973), .Q(n11304) );
  OR2X1 U11359 ( .IN1(WX8471), .IN2(n9448), .Q(n11303) );
  OR2X1 U11360 ( .IN1(n11305), .IN2(n11306), .Q(n11302) );
  INVX0 U11361 ( .INP(n11307), .ZN(n11306) );
  OR2X1 U11362 ( .IN1(n11308), .IN2(n7974), .Q(n11307) );
  AND2X1 U11363 ( .IN1(n7974), .IN2(n11308), .Q(n11305) );
  INVX0 U11364 ( .INP(n11309), .ZN(n11308) );
  OR2X1 U11365 ( .IN1(n11310), .IN2(n11311), .Q(n11309) );
  AND2X1 U11366 ( .IN1(n8796), .IN2(n8376), .Q(n11311) );
  AND2X1 U11367 ( .IN1(n15905), .IN2(WX8599), .Q(n11310) );
  AND2X1 U11368 ( .IN1(test_so66), .IN2(n9227), .Q(n11294) );
  AND2X1 U11369 ( .IN1(n1232), .IN2(n9220), .Q(n11293) );
  INVX0 U11370 ( .INP(n11312), .ZN(n1232) );
  OR2X1 U11371 ( .IN1(n9570), .IN2(n3908), .Q(n11312) );
  OR4X1 U11372 ( .IN1(n11313), .IN2(n11314), .IN3(n11315), .IN4(n11316), .Q(
        WX7111) );
  AND2X1 U11373 ( .IN1(n9179), .IN2(n11317), .Q(n11316) );
  AND2X1 U11374 ( .IN1(n10662), .IN2(n9259), .Q(n11315) );
  AND2X1 U11375 ( .IN1(n11318), .IN2(n11319), .Q(n10662) );
  INVX0 U11376 ( .INP(n11320), .ZN(n11319) );
  AND2X1 U11377 ( .IN1(n11321), .IN2(n11322), .Q(n11320) );
  OR2X1 U11378 ( .IN1(n11322), .IN2(n11321), .Q(n11318) );
  OR2X1 U11379 ( .IN1(n11323), .IN2(n11324), .Q(n11321) );
  AND2X1 U11380 ( .IN1(n9451), .IN2(WX8533), .Q(n11324) );
  AND2X1 U11381 ( .IN1(n7975), .IN2(n9465), .Q(n11323) );
  AND2X1 U11382 ( .IN1(n11325), .IN2(n11326), .Q(n11322) );
  OR2X1 U11383 ( .IN1(n11327), .IN2(n8795), .Q(n11326) );
  OR2X1 U11384 ( .IN1(WX8597), .IN2(n11328), .Q(n11325) );
  INVX0 U11385 ( .INP(n11327), .ZN(n11328) );
  AND2X1 U11386 ( .IN1(n11329), .IN2(n11330), .Q(n11327) );
  OR2X1 U11387 ( .IN1(n8377), .IN2(test_so70), .Q(n11330) );
  OR2X1 U11388 ( .IN1(n9119), .IN2(n15906), .Q(n11329) );
  AND2X1 U11389 ( .IN1(n9245), .IN2(CRC_OUT_4_30), .Q(n11314) );
  AND2X1 U11390 ( .IN1(n1231), .IN2(n9220), .Q(n11313) );
  INVX0 U11391 ( .INP(n11331), .ZN(n1231) );
  OR2X1 U11392 ( .IN1(n9569), .IN2(n3909), .Q(n11331) );
  OR4X1 U11393 ( .IN1(n11332), .IN2(n11333), .IN3(n11334), .IN4(n11335), .Q(
        WX7109) );
  AND2X1 U11394 ( .IN1(n9179), .IN2(n11336), .Q(n11335) );
  AND2X1 U11395 ( .IN1(n9275), .IN2(n10682), .Q(n11334) );
  OR2X1 U11396 ( .IN1(n11337), .IN2(n11338), .Q(n10682) );
  INVX0 U11397 ( .INP(n11339), .ZN(n11338) );
  OR2X1 U11398 ( .IN1(n11340), .IN2(n11341), .Q(n11339) );
  AND2X1 U11399 ( .IN1(n11341), .IN2(n11340), .Q(n11337) );
  AND2X1 U11400 ( .IN1(n11342), .IN2(n11343), .Q(n11340) );
  OR2X1 U11401 ( .IN1(n9465), .IN2(n7880), .Q(n11343) );
  OR2X1 U11402 ( .IN1(WX8467), .IN2(n9447), .Q(n11342) );
  OR2X1 U11403 ( .IN1(n11344), .IN2(n11345), .Q(n11341) );
  INVX0 U11404 ( .INP(n11346), .ZN(n11345) );
  OR2X1 U11405 ( .IN1(n11347), .IN2(n7881), .Q(n11346) );
  AND2X1 U11406 ( .IN1(n7881), .IN2(n11347), .Q(n11344) );
  INVX0 U11407 ( .INP(n11348), .ZN(n11347) );
  OR2X1 U11408 ( .IN1(n11349), .IN2(n11350), .Q(n11348) );
  AND2X1 U11409 ( .IN1(n8794), .IN2(n8378), .Q(n11350) );
  AND2X1 U11410 ( .IN1(n15907), .IN2(WX8595), .Q(n11349) );
  AND2X1 U11411 ( .IN1(n2245), .IN2(WX6950), .Q(n11333) );
  AND2X1 U11412 ( .IN1(n9245), .IN2(CRC_OUT_4_31), .Q(n11332) );
  OR4X1 U11413 ( .IN1(n11351), .IN2(n11352), .IN3(n11353), .IN4(n11354), .Q(
        WX706) );
  AND2X1 U11414 ( .IN1(n9179), .IN2(n11355), .Q(n11354) );
  AND2X1 U11415 ( .IN1(n11356), .IN2(n9259), .Q(n11353) );
  AND2X1 U11416 ( .IN1(n9245), .IN2(CRC_OUT_9_0), .Q(n11352) );
  AND2X1 U11417 ( .IN1(WX544), .IN2(n9220), .Q(n11351) );
  OR4X1 U11418 ( .IN1(n11357), .IN2(n11358), .IN3(n11359), .IN4(n11360), .Q(
        WX704) );
  AND2X1 U11419 ( .IN1(n9179), .IN2(n11361), .Q(n11360) );
  AND2X1 U11420 ( .IN1(n9275), .IN2(n11362), .Q(n11359) );
  AND2X1 U11421 ( .IN1(test_so9), .IN2(n9228), .Q(n11358) );
  AND2X1 U11422 ( .IN1(WX542), .IN2(n9220), .Q(n11357) );
  OR4X1 U11423 ( .IN1(n11363), .IN2(n11364), .IN3(n11365), .IN4(n11366), .Q(
        WX702) );
  AND2X1 U11424 ( .IN1(n11367), .IN2(n9176), .Q(n11366) );
  AND2X1 U11425 ( .IN1(n9275), .IN2(n11368), .Q(n11365) );
  AND2X1 U11426 ( .IN1(n9245), .IN2(CRC_OUT_9_2), .Q(n11364) );
  AND2X1 U11427 ( .IN1(WX540), .IN2(n9220), .Q(n11363) );
  AND2X1 U11428 ( .IN1(n9049), .IN2(n9497), .Q(WX7011) );
  OR4X1 U11429 ( .IN1(n11369), .IN2(n11370), .IN3(n11371), .IN4(n11372), .Q(
        WX700) );
  AND2X1 U11430 ( .IN1(n9179), .IN2(n11373), .Q(n11372) );
  AND2X1 U11431 ( .IN1(n9275), .IN2(n11374), .Q(n11371) );
  AND2X1 U11432 ( .IN1(n9245), .IN2(CRC_OUT_9_3), .Q(n11370) );
  AND2X1 U11433 ( .IN1(WX538), .IN2(n9220), .Q(n11369) );
  OR4X1 U11434 ( .IN1(n11375), .IN2(n11376), .IN3(n11377), .IN4(n11378), .Q(
        WX698) );
  AND2X1 U11435 ( .IN1(n9179), .IN2(n11379), .Q(n11378) );
  AND2X1 U11436 ( .IN1(n11380), .IN2(n9259), .Q(n11377) );
  AND2X1 U11437 ( .IN1(n9245), .IN2(CRC_OUT_9_4), .Q(n11376) );
  AND2X1 U11438 ( .IN1(WX536), .IN2(n9220), .Q(n11375) );
  OR4X1 U11439 ( .IN1(n11381), .IN2(n11382), .IN3(n11383), .IN4(n11384), .Q(
        WX696) );
  AND2X1 U11440 ( .IN1(n9179), .IN2(n11385), .Q(n11384) );
  AND2X1 U11441 ( .IN1(n9276), .IN2(n11386), .Q(n11383) );
  AND2X1 U11442 ( .IN1(n9245), .IN2(CRC_OUT_9_5), .Q(n11382) );
  AND2X1 U11443 ( .IN1(WX534), .IN2(n9220), .Q(n11381) );
  OR4X1 U11444 ( .IN1(n11387), .IN2(n11388), .IN3(n11389), .IN4(n11390), .Q(
        WX694) );
  AND2X1 U11445 ( .IN1(n11391), .IN2(n9176), .Q(n11390) );
  AND2X1 U11446 ( .IN1(n9276), .IN2(n11392), .Q(n11389) );
  AND2X1 U11447 ( .IN1(n9245), .IN2(CRC_OUT_9_6), .Q(n11388) );
  AND2X1 U11448 ( .IN1(WX532), .IN2(n9220), .Q(n11387) );
  OR4X1 U11449 ( .IN1(n11393), .IN2(n11394), .IN3(n11395), .IN4(n11396), .Q(
        WX692) );
  AND2X1 U11450 ( .IN1(n9179), .IN2(n11397), .Q(n11396) );
  AND2X1 U11451 ( .IN1(n9276), .IN2(n11398), .Q(n11395) );
  AND2X1 U11452 ( .IN1(n9245), .IN2(CRC_OUT_9_7), .Q(n11394) );
  AND2X1 U11453 ( .IN1(WX530), .IN2(n9220), .Q(n11393) );
  OR4X1 U11454 ( .IN1(n11399), .IN2(n11400), .IN3(n11401), .IN4(n11402), .Q(
        WX690) );
  AND2X1 U11455 ( .IN1(n9180), .IN2(n11403), .Q(n11402) );
  AND2X1 U11456 ( .IN1(n9276), .IN2(n11404), .Q(n11401) );
  AND2X1 U11457 ( .IN1(n9246), .IN2(CRC_OUT_9_8), .Q(n11400) );
  AND2X1 U11458 ( .IN1(WX528), .IN2(n9221), .Q(n11399) );
  OR4X1 U11459 ( .IN1(n11405), .IN2(n11406), .IN3(n11407), .IN4(n11408), .Q(
        WX688) );
  AND2X1 U11460 ( .IN1(n9180), .IN2(n11409), .Q(n11408) );
  AND2X1 U11461 ( .IN1(n9276), .IN2(n11410), .Q(n11407) );
  AND2X1 U11462 ( .IN1(n9246), .IN2(CRC_OUT_9_9), .Q(n11406) );
  AND2X1 U11463 ( .IN1(WX526), .IN2(n9221), .Q(n11405) );
  OR4X1 U11464 ( .IN1(n11411), .IN2(n11412), .IN3(n11413), .IN4(n11414), .Q(
        WX686) );
  AND2X1 U11465 ( .IN1(n11415), .IN2(n9175), .Q(n11414) );
  AND2X1 U11466 ( .IN1(n11416), .IN2(n9258), .Q(n11413) );
  AND2X1 U11467 ( .IN1(n9246), .IN2(CRC_OUT_9_10), .Q(n11412) );
  AND2X1 U11468 ( .IN1(WX524), .IN2(n9221), .Q(n11411) );
  OR4X1 U11469 ( .IN1(n11417), .IN2(n11418), .IN3(n11419), .IN4(n11420), .Q(
        WX684) );
  AND2X1 U11470 ( .IN1(n9180), .IN2(n11421), .Q(n11420) );
  AND2X1 U11471 ( .IN1(n9276), .IN2(n11422), .Q(n11419) );
  AND2X1 U11472 ( .IN1(n9246), .IN2(CRC_OUT_9_11), .Q(n11418) );
  AND2X1 U11473 ( .IN1(WX522), .IN2(n9221), .Q(n11417) );
  OR4X1 U11474 ( .IN1(n11423), .IN2(n11424), .IN3(n11425), .IN4(n11426), .Q(
        WX682) );
  AND2X1 U11475 ( .IN1(n9180), .IN2(n11427), .Q(n11426) );
  AND2X1 U11476 ( .IN1(n9276), .IN2(n11428), .Q(n11425) );
  AND2X1 U11477 ( .IN1(n9246), .IN2(CRC_OUT_9_12), .Q(n11424) );
  AND2X1 U11478 ( .IN1(WX520), .IN2(n9221), .Q(n11423) );
  OR4X1 U11479 ( .IN1(n11429), .IN2(n11430), .IN3(n11431), .IN4(n11432), .Q(
        WX680) );
  AND2X1 U11480 ( .IN1(n9180), .IN2(n11433), .Q(n11432) );
  AND2X1 U11481 ( .IN1(n9276), .IN2(n11434), .Q(n11431) );
  AND2X1 U11482 ( .IN1(n9246), .IN2(CRC_OUT_9_13), .Q(n11430) );
  AND2X1 U11483 ( .IN1(WX518), .IN2(n9221), .Q(n11429) );
  OR4X1 U11484 ( .IN1(n11435), .IN2(n11436), .IN3(n11437), .IN4(n11438), .Q(
        WX678) );
  AND2X1 U11485 ( .IN1(n9180), .IN2(n11439), .Q(n11438) );
  AND2X1 U11486 ( .IN1(n11440), .IN2(n9258), .Q(n11437) );
  AND2X1 U11487 ( .IN1(n9246), .IN2(CRC_OUT_9_14), .Q(n11436) );
  AND2X1 U11488 ( .IN1(WX516), .IN2(n9221), .Q(n11435) );
  OR4X1 U11489 ( .IN1(n11441), .IN2(n11442), .IN3(n11443), .IN4(n11444), .Q(
        WX676) );
  AND2X1 U11490 ( .IN1(n9180), .IN2(n11445), .Q(n11444) );
  AND2X1 U11491 ( .IN1(n9276), .IN2(n11446), .Q(n11443) );
  AND2X1 U11492 ( .IN1(n9246), .IN2(CRC_OUT_9_15), .Q(n11442) );
  AND2X1 U11493 ( .IN1(WX514), .IN2(n9221), .Q(n11441) );
  OR4X1 U11494 ( .IN1(n11447), .IN2(n11448), .IN3(n11449), .IN4(n11450), .Q(
        WX674) );
  AND2X1 U11495 ( .IN1(n11451), .IN2(n9175), .Q(n11450) );
  AND2X1 U11496 ( .IN1(n9276), .IN2(n11452), .Q(n11449) );
  AND2X1 U11497 ( .IN1(n9246), .IN2(CRC_OUT_9_16), .Q(n11448) );
  AND2X1 U11498 ( .IN1(WX512), .IN2(n9221), .Q(n11447) );
  OR4X1 U11499 ( .IN1(n11453), .IN2(n11454), .IN3(n11455), .IN4(n11456), .Q(
        WX672) );
  AND2X1 U11500 ( .IN1(n9180), .IN2(n11457), .Q(n11456) );
  AND2X1 U11501 ( .IN1(n9276), .IN2(n11458), .Q(n11455) );
  AND2X1 U11502 ( .IN1(n9246), .IN2(CRC_OUT_9_17), .Q(n11454) );
  AND2X1 U11503 ( .IN1(WX510), .IN2(n9221), .Q(n11453) );
  OR4X1 U11504 ( .IN1(n11459), .IN2(n11460), .IN3(n11461), .IN4(n11462), .Q(
        WX670) );
  AND2X1 U11505 ( .IN1(n9180), .IN2(n11463), .Q(n11462) );
  AND2X1 U11506 ( .IN1(n11464), .IN2(n9258), .Q(n11461) );
  AND2X1 U11507 ( .IN1(n9246), .IN2(CRC_OUT_9_18), .Q(n11460) );
  AND2X1 U11508 ( .IN1(WX508), .IN2(n9221), .Q(n11459) );
  OR4X1 U11509 ( .IN1(n11465), .IN2(n11466), .IN3(n11467), .IN4(n11468), .Q(
        WX668) );
  AND2X1 U11510 ( .IN1(n9180), .IN2(n11469), .Q(n11468) );
  AND2X1 U11511 ( .IN1(n9276), .IN2(n11470), .Q(n11467) );
  AND2X1 U11512 ( .IN1(test_so10), .IN2(n9227), .Q(n11466) );
  AND2X1 U11513 ( .IN1(WX506), .IN2(n9222), .Q(n11465) );
  OR4X1 U11514 ( .IN1(n11471), .IN2(n11472), .IN3(n11473), .IN4(n11474), .Q(
        WX666) );
  AND2X1 U11515 ( .IN1(n11475), .IN2(n9174), .Q(n11474) );
  AND2X1 U11516 ( .IN1(n9276), .IN2(n11476), .Q(n11473) );
  AND2X1 U11517 ( .IN1(n9246), .IN2(CRC_OUT_9_20), .Q(n11472) );
  AND2X1 U11518 ( .IN1(WX504), .IN2(n9221), .Q(n11471) );
  OR4X1 U11519 ( .IN1(n11477), .IN2(n11478), .IN3(n11479), .IN4(n11480), .Q(
        WX664) );
  AND2X1 U11520 ( .IN1(n9180), .IN2(n11481), .Q(n11480) );
  AND2X1 U11521 ( .IN1(n9277), .IN2(n11482), .Q(n11479) );
  AND2X1 U11522 ( .IN1(n9246), .IN2(CRC_OUT_9_21), .Q(n11478) );
  AND2X1 U11523 ( .IN1(WX502), .IN2(n9222), .Q(n11477) );
  OR4X1 U11524 ( .IN1(n11483), .IN2(n11484), .IN3(n11485), .IN4(n11486), .Q(
        WX662) );
  AND2X1 U11525 ( .IN1(n9180), .IN2(n11487), .Q(n11486) );
  AND2X1 U11526 ( .IN1(n11488), .IN2(n9258), .Q(n11485) );
  AND2X1 U11527 ( .IN1(n9247), .IN2(CRC_OUT_9_22), .Q(n11484) );
  AND2X1 U11528 ( .IN1(WX500), .IN2(n9222), .Q(n11483) );
  OR4X1 U11529 ( .IN1(n11489), .IN2(n11490), .IN3(n11491), .IN4(n11492), .Q(
        WX660) );
  AND2X1 U11530 ( .IN1(n9180), .IN2(n11493), .Q(n11492) );
  AND2X1 U11531 ( .IN1(n9277), .IN2(n11494), .Q(n11491) );
  AND2X1 U11532 ( .IN1(n9247), .IN2(CRC_OUT_9_23), .Q(n11490) );
  AND2X1 U11533 ( .IN1(WX498), .IN2(n9222), .Q(n11489) );
  OR4X1 U11534 ( .IN1(n11495), .IN2(n11496), .IN3(n11497), .IN4(n11498), .Q(
        WX658) );
  AND2X1 U11535 ( .IN1(n11499), .IN2(n9174), .Q(n11498) );
  AND2X1 U11536 ( .IN1(n9277), .IN2(n11500), .Q(n11497) );
  AND2X1 U11537 ( .IN1(n9247), .IN2(CRC_OUT_9_24), .Q(n11496) );
  AND2X1 U11538 ( .IN1(WX496), .IN2(n9222), .Q(n11495) );
  OR4X1 U11539 ( .IN1(n11501), .IN2(n11502), .IN3(n11503), .IN4(n11504), .Q(
        WX656) );
  AND2X1 U11540 ( .IN1(n9181), .IN2(n11505), .Q(n11504) );
  AND2X1 U11541 ( .IN1(n9277), .IN2(n11506), .Q(n11503) );
  AND2X1 U11542 ( .IN1(n9247), .IN2(CRC_OUT_9_25), .Q(n11502) );
  AND2X1 U11543 ( .IN1(WX494), .IN2(n9222), .Q(n11501) );
  OR4X1 U11544 ( .IN1(n11507), .IN2(n11508), .IN3(n11509), .IN4(n11510), .Q(
        WX654) );
  AND2X1 U11545 ( .IN1(n9181), .IN2(n11511), .Q(n11510) );
  AND2X1 U11546 ( .IN1(n9277), .IN2(n11512), .Q(n11509) );
  AND2X1 U11547 ( .IN1(n9247), .IN2(CRC_OUT_9_26), .Q(n11508) );
  AND2X1 U11548 ( .IN1(WX492), .IN2(n9222), .Q(n11507) );
  OR4X1 U11549 ( .IN1(n11513), .IN2(n11514), .IN3(n11515), .IN4(n11516), .Q(
        WX652) );
  AND2X1 U11550 ( .IN1(n9181), .IN2(n11517), .Q(n11516) );
  AND2X1 U11551 ( .IN1(n9277), .IN2(n11518), .Q(n11515) );
  AND2X1 U11552 ( .IN1(n9247), .IN2(CRC_OUT_9_27), .Q(n11514) );
  AND2X1 U11553 ( .IN1(WX490), .IN2(n9222), .Q(n11513) );
  OR4X1 U11554 ( .IN1(n11519), .IN2(n11520), .IN3(n11521), .IN4(n11522), .Q(
        WX650) );
  AND2X1 U11555 ( .IN1(n11523), .IN2(n9173), .Q(n11522) );
  AND2X1 U11556 ( .IN1(n11524), .IN2(n9258), .Q(n11521) );
  AND2X1 U11557 ( .IN1(n9247), .IN2(CRC_OUT_9_28), .Q(n11520) );
  AND2X1 U11558 ( .IN1(WX488), .IN2(n9222), .Q(n11519) );
  AND3X1 U11559 ( .IN1(n11525), .IN2(n11526), .IN3(n9533), .Q(WX6498) );
  OR2X1 U11560 ( .IN1(DFF_958_n1), .IN2(WX6009), .Q(n11526) );
  OR2X1 U11561 ( .IN1(n8847), .IN2(CRC_OUT_5_30), .Q(n11525) );
  AND3X1 U11562 ( .IN1(n11527), .IN2(n11528), .IN3(n9533), .Q(WX6496) );
  OR2X1 U11563 ( .IN1(DFF_957_n1), .IN2(WX6011), .Q(n11528) );
  OR2X1 U11564 ( .IN1(n8848), .IN2(CRC_OUT_5_29), .Q(n11527) );
  AND3X1 U11565 ( .IN1(n11529), .IN2(n11530), .IN3(n9533), .Q(WX6494) );
  OR2X1 U11566 ( .IN1(DFF_956_n1), .IN2(WX6013), .Q(n11530) );
  OR2X1 U11567 ( .IN1(n8849), .IN2(CRC_OUT_5_28), .Q(n11529) );
  AND3X1 U11568 ( .IN1(n11531), .IN2(n11532), .IN3(n9532), .Q(WX6492) );
  OR2X1 U11569 ( .IN1(DFF_955_n1), .IN2(WX6015), .Q(n11532) );
  OR2X1 U11570 ( .IN1(n8850), .IN2(CRC_OUT_5_27), .Q(n11531) );
  AND3X1 U11571 ( .IN1(n11533), .IN2(n11534), .IN3(n9532), .Q(WX6490) );
  OR2X1 U11572 ( .IN1(DFF_954_n1), .IN2(WX6017), .Q(n11534) );
  OR2X1 U11573 ( .IN1(n8851), .IN2(CRC_OUT_5_26), .Q(n11533) );
  AND3X1 U11574 ( .IN1(n11535), .IN2(n11536), .IN3(n9532), .Q(WX6488) );
  OR2X1 U11575 ( .IN1(DFF_953_n1), .IN2(WX6019), .Q(n11536) );
  OR2X1 U11576 ( .IN1(n8852), .IN2(CRC_OUT_5_25), .Q(n11535) );
  AND3X1 U11577 ( .IN1(n11537), .IN2(n11538), .IN3(n9532), .Q(WX6486) );
  OR2X1 U11578 ( .IN1(DFF_952_n1), .IN2(WX6021), .Q(n11538) );
  OR2X1 U11579 ( .IN1(n8853), .IN2(CRC_OUT_5_24), .Q(n11537) );
  AND3X1 U11580 ( .IN1(n11539), .IN2(n11540), .IN3(n9532), .Q(WX6484) );
  OR2X1 U11581 ( .IN1(DFF_951_n1), .IN2(WX6023), .Q(n11540) );
  OR2X1 U11582 ( .IN1(n8854), .IN2(CRC_OUT_5_23), .Q(n11539) );
  AND3X1 U11583 ( .IN1(n11541), .IN2(n11542), .IN3(n9532), .Q(WX6482) );
  OR2X1 U11584 ( .IN1(DFF_950_n1), .IN2(WX6025), .Q(n11542) );
  OR2X1 U11585 ( .IN1(n8855), .IN2(CRC_OUT_5_22), .Q(n11541) );
  AND3X1 U11586 ( .IN1(n11543), .IN2(n11544), .IN3(n9532), .Q(WX6480) );
  OR2X1 U11587 ( .IN1(DFF_949_n1), .IN2(WX6027), .Q(n11544) );
  OR2X1 U11588 ( .IN1(n8856), .IN2(CRC_OUT_5_21), .Q(n11543) );
  OR4X1 U11589 ( .IN1(n11545), .IN2(n11546), .IN3(n11547), .IN4(n11548), .Q(
        WX648) );
  AND2X1 U11590 ( .IN1(n9181), .IN2(n11549), .Q(n11548) );
  AND2X1 U11591 ( .IN1(n9277), .IN2(n11550), .Q(n11547) );
  AND2X1 U11592 ( .IN1(n9247), .IN2(CRC_OUT_9_29), .Q(n11546) );
  AND2X1 U11593 ( .IN1(WX486), .IN2(n9222), .Q(n11545) );
  AND3X1 U11594 ( .IN1(n11551), .IN2(n11552), .IN3(n9532), .Q(WX6478) );
  OR2X1 U11595 ( .IN1(DFF_948_n1), .IN2(WX6029), .Q(n11552) );
  OR2X1 U11596 ( .IN1(n8857), .IN2(CRC_OUT_5_20), .Q(n11551) );
  AND3X1 U11597 ( .IN1(n11553), .IN2(n11554), .IN3(n9532), .Q(WX6476) );
  OR2X1 U11598 ( .IN1(DFF_947_n1), .IN2(WX6031), .Q(n11554) );
  OR2X1 U11599 ( .IN1(n8858), .IN2(CRC_OUT_5_19), .Q(n11553) );
  AND3X1 U11600 ( .IN1(n11555), .IN2(n11556), .IN3(n9532), .Q(WX6474) );
  OR2X1 U11601 ( .IN1(DFF_946_n1), .IN2(WX6033), .Q(n11556) );
  OR2X1 U11602 ( .IN1(n8859), .IN2(CRC_OUT_5_18), .Q(n11555) );
  AND2X1 U11603 ( .IN1(n11557), .IN2(n9496), .Q(WX6472) );
  OR2X1 U11604 ( .IN1(n11558), .IN2(n11559), .Q(n11557) );
  AND2X1 U11605 ( .IN1(n8860), .IN2(n9154), .Q(n11559) );
  AND2X1 U11606 ( .IN1(test_so54), .IN2(WX6035), .Q(n11558) );
  AND3X1 U11607 ( .IN1(n11560), .IN2(n11561), .IN3(n9532), .Q(WX6470) );
  OR2X1 U11608 ( .IN1(DFF_944_n1), .IN2(WX6037), .Q(n11561) );
  OR2X1 U11609 ( .IN1(n8861), .IN2(CRC_OUT_5_16), .Q(n11560) );
  AND3X1 U11610 ( .IN1(n11562), .IN2(n11563), .IN3(n9532), .Q(WX6468) );
  OR2X1 U11611 ( .IN1(DFF_943_n1), .IN2(n11564), .Q(n11563) );
  AND2X1 U11612 ( .IN1(n11565), .IN2(n11566), .Q(n11564) );
  OR2X1 U11613 ( .IN1(DFF_959_n1), .IN2(n9089), .Q(n11566) );
  OR2X1 U11614 ( .IN1(test_so52), .IN2(CRC_OUT_5_31), .Q(n11565) );
  OR3X1 U11615 ( .IN1(n11567), .IN2(n11568), .IN3(CRC_OUT_5_15), .Q(n11562) );
  AND2X1 U11616 ( .IN1(DFF_959_n1), .IN2(n9089), .Q(n11568) );
  AND2X1 U11617 ( .IN1(test_so52), .IN2(CRC_OUT_5_31), .Q(n11567) );
  AND3X1 U11618 ( .IN1(n11569), .IN2(n11570), .IN3(n9531), .Q(WX6466) );
  OR2X1 U11619 ( .IN1(DFF_942_n1), .IN2(WX6041), .Q(n11570) );
  OR2X1 U11620 ( .IN1(n8862), .IN2(CRC_OUT_5_14), .Q(n11569) );
  AND3X1 U11621 ( .IN1(n11571), .IN2(n11572), .IN3(n9531), .Q(WX6464) );
  OR2X1 U11622 ( .IN1(DFF_941_n1), .IN2(WX6043), .Q(n11572) );
  OR2X1 U11623 ( .IN1(n8863), .IN2(CRC_OUT_5_13), .Q(n11571) );
  AND3X1 U11624 ( .IN1(n11573), .IN2(n11574), .IN3(n9531), .Q(WX6462) );
  OR2X1 U11625 ( .IN1(DFF_940_n1), .IN2(WX6045), .Q(n11574) );
  OR2X1 U11626 ( .IN1(n8864), .IN2(CRC_OUT_5_12), .Q(n11573) );
  AND3X1 U11627 ( .IN1(n11575), .IN2(n11576), .IN3(n9531), .Q(WX6460) );
  OR2X1 U11628 ( .IN1(DFF_939_n1), .IN2(WX6047), .Q(n11576) );
  OR2X1 U11629 ( .IN1(n8865), .IN2(CRC_OUT_5_11), .Q(n11575) );
  OR4X1 U11630 ( .IN1(n11577), .IN2(n11578), .IN3(n11579), .IN4(n11580), .Q(
        WX646) );
  AND2X1 U11631 ( .IN1(n9195), .IN2(n11581), .Q(n11580) );
  AND2X1 U11632 ( .IN1(n9277), .IN2(n11582), .Q(n11579) );
  AND2X1 U11633 ( .IN1(n9247), .IN2(CRC_OUT_9_30), .Q(n11578) );
  AND2X1 U11634 ( .IN1(WX484), .IN2(n9222), .Q(n11577) );
  AND2X1 U11635 ( .IN1(n11583), .IN2(n9495), .Q(WX6458) );
  OR2X1 U11636 ( .IN1(n11584), .IN2(n11585), .Q(n11583) );
  AND2X1 U11637 ( .IN1(n11586), .IN2(CRC_OUT_5_10), .Q(n11585) );
  AND2X1 U11638 ( .IN1(DFF_938_n1), .IN2(n11587), .Q(n11584) );
  INVX0 U11639 ( .INP(n11586), .ZN(n11587) );
  OR2X1 U11640 ( .IN1(n11588), .IN2(n11589), .Q(n11586) );
  AND2X1 U11641 ( .IN1(DFF_959_n1), .IN2(WX6049), .Q(n11589) );
  AND2X1 U11642 ( .IN1(n8724), .IN2(CRC_OUT_5_31), .Q(n11588) );
  AND3X1 U11643 ( .IN1(n11590), .IN2(n11591), .IN3(n9531), .Q(WX6456) );
  OR2X1 U11644 ( .IN1(DFF_937_n1), .IN2(WX6051), .Q(n11591) );
  OR2X1 U11645 ( .IN1(n8866), .IN2(CRC_OUT_5_9), .Q(n11590) );
  AND3X1 U11646 ( .IN1(n11592), .IN2(n11593), .IN3(n9531), .Q(WX6454) );
  OR2X1 U11647 ( .IN1(DFF_936_n1), .IN2(WX6053), .Q(n11593) );
  OR2X1 U11648 ( .IN1(n8867), .IN2(CRC_OUT_5_8), .Q(n11592) );
  AND3X1 U11649 ( .IN1(n11594), .IN2(n11595), .IN3(n9531), .Q(WX6452) );
  OR2X1 U11650 ( .IN1(DFF_935_n1), .IN2(WX6055), .Q(n11595) );
  OR2X1 U11651 ( .IN1(n8868), .IN2(CRC_OUT_5_7), .Q(n11594) );
  AND3X1 U11652 ( .IN1(n11596), .IN2(n11597), .IN3(n9531), .Q(WX6450) );
  OR2X1 U11653 ( .IN1(DFF_934_n1), .IN2(WX6057), .Q(n11597) );
  OR2X1 U11654 ( .IN1(n8869), .IN2(CRC_OUT_5_6), .Q(n11596) );
  AND3X1 U11655 ( .IN1(n11598), .IN2(n11599), .IN3(n9531), .Q(WX6448) );
  OR2X1 U11656 ( .IN1(DFF_933_n1), .IN2(WX6059), .Q(n11599) );
  OR2X1 U11657 ( .IN1(n8870), .IN2(CRC_OUT_5_5), .Q(n11598) );
  AND3X1 U11658 ( .IN1(n11600), .IN2(n11601), .IN3(n9531), .Q(WX6446) );
  OR2X1 U11659 ( .IN1(DFF_932_n1), .IN2(WX6061), .Q(n11601) );
  OR2X1 U11660 ( .IN1(n8871), .IN2(CRC_OUT_5_4), .Q(n11600) );
  AND2X1 U11661 ( .IN1(n11602), .IN2(n9495), .Q(WX6444) );
  OR2X1 U11662 ( .IN1(n11603), .IN2(n11604), .Q(n11602) );
  AND2X1 U11663 ( .IN1(n11605), .IN2(CRC_OUT_5_3), .Q(n11604) );
  AND2X1 U11664 ( .IN1(DFF_931_n1), .IN2(n11606), .Q(n11603) );
  INVX0 U11665 ( .INP(n11605), .ZN(n11606) );
  OR2X1 U11666 ( .IN1(n11607), .IN2(n11608), .Q(n11605) );
  AND2X1 U11667 ( .IN1(DFF_959_n1), .IN2(WX6063), .Q(n11608) );
  AND2X1 U11668 ( .IN1(n8725), .IN2(CRC_OUT_5_31), .Q(n11607) );
  AND3X1 U11669 ( .IN1(n11609), .IN2(n11610), .IN3(n9531), .Q(WX6442) );
  OR2X1 U11670 ( .IN1(DFF_930_n1), .IN2(WX6065), .Q(n11610) );
  OR2X1 U11671 ( .IN1(n8872), .IN2(CRC_OUT_5_2), .Q(n11609) );
  AND3X1 U11672 ( .IN1(n11611), .IN2(n11612), .IN3(n9531), .Q(WX6440) );
  OR2X1 U11673 ( .IN1(DFF_929_n1), .IN2(WX6067), .Q(n11612) );
  OR2X1 U11674 ( .IN1(n8873), .IN2(CRC_OUT_5_1), .Q(n11611) );
  OR4X1 U11675 ( .IN1(n11613), .IN2(n11614), .IN3(n11615), .IN4(n11616), .Q(
        WX644) );
  AND2X1 U11676 ( .IN1(n9195), .IN2(n11617), .Q(n11616) );
  AND2X1 U11677 ( .IN1(n9277), .IN2(n11618), .Q(n11615) );
  AND2X1 U11678 ( .IN1(n2245), .IN2(WX485), .Q(n11614) );
  AND2X1 U11679 ( .IN1(n9247), .IN2(CRC_OUT_9_31), .Q(n11613) );
  AND2X1 U11680 ( .IN1(n11619), .IN2(n9493), .Q(WX6438) );
  OR2X1 U11681 ( .IN1(n11620), .IN2(n11621), .Q(n11619) );
  AND2X1 U11682 ( .IN1(n8874), .IN2(n9155), .Q(n11621) );
  AND2X1 U11683 ( .IN1(test_so53), .IN2(WX6069), .Q(n11620) );
  AND3X1 U11684 ( .IN1(n11622), .IN2(n11623), .IN3(n9530), .Q(WX6436) );
  OR2X1 U11685 ( .IN1(DFF_959_n1), .IN2(WX6071), .Q(n11623) );
  OR2X1 U11686 ( .IN1(n8738), .IN2(CRC_OUT_5_31), .Q(n11622) );
  AND2X1 U11687 ( .IN1(n9501), .IN2(n8479), .Q(WX5910) );
  AND2X1 U11688 ( .IN1(n9500), .IN2(n8480), .Q(WX5908) );
  AND2X1 U11689 ( .IN1(n9500), .IN2(n8481), .Q(WX5906) );
  AND2X1 U11690 ( .IN1(n9501), .IN2(n8482), .Q(WX5904) );
  AND2X1 U11691 ( .IN1(n9501), .IN2(n8483), .Q(WX5902) );
  AND2X1 U11692 ( .IN1(n9502), .IN2(n8484), .Q(WX5900) );
  AND2X1 U11693 ( .IN1(test_so46), .IN2(n9494), .Q(WX5898) );
  AND2X1 U11694 ( .IN1(n9502), .IN2(n8487), .Q(WX5896) );
  AND2X1 U11695 ( .IN1(n9501), .IN2(n8488), .Q(WX5894) );
  AND2X1 U11696 ( .IN1(n9502), .IN2(n8489), .Q(WX5892) );
  AND2X1 U11697 ( .IN1(n9501), .IN2(n8490), .Q(WX5890) );
  AND2X1 U11698 ( .IN1(n9501), .IN2(n8491), .Q(WX5888) );
  AND2X1 U11699 ( .IN1(n9503), .IN2(n8492), .Q(WX5886) );
  AND2X1 U11700 ( .IN1(n9502), .IN2(n8493), .Q(WX5884) );
  AND2X1 U11701 ( .IN1(n9503), .IN2(n8494), .Q(WX5882) );
  AND2X1 U11702 ( .IN1(n9503), .IN2(n8495), .Q(WX5880) );
  OR4X1 U11703 ( .IN1(n11624), .IN2(n11625), .IN3(n11626), .IN4(n11627), .Q(
        WX5878) );
  AND2X1 U11704 ( .IN1(n9195), .IN2(n11628), .Q(n11627) );
  AND2X1 U11705 ( .IN1(n9277), .IN2(n10782), .Q(n11626) );
  OR2X1 U11706 ( .IN1(n11629), .IN2(n11630), .Q(n10782) );
  INVX0 U11707 ( .INP(n11631), .ZN(n11630) );
  OR2X1 U11708 ( .IN1(n11632), .IN2(n11633), .Q(n11631) );
  AND2X1 U11709 ( .IN1(n11633), .IN2(n11632), .Q(n11629) );
  AND2X1 U11710 ( .IN1(n11634), .IN2(n11635), .Q(n11632) );
  OR2X1 U11711 ( .IN1(WX7236), .IN2(n8209), .Q(n11635) );
  INVX0 U11712 ( .INP(n11636), .ZN(n11634) );
  AND2X1 U11713 ( .IN1(n8209), .IN2(WX7236), .Q(n11636) );
  OR2X1 U11714 ( .IN1(n11637), .IN2(n11638), .Q(n11633) );
  AND2X1 U11715 ( .IN1(n8210), .IN2(WX7364), .Q(n11638) );
  AND2X1 U11716 ( .IN1(n8737), .IN2(WX7300), .Q(n11637) );
  AND2X1 U11717 ( .IN1(test_so53), .IN2(n9228), .Q(n11625) );
  AND2X1 U11718 ( .IN1(n1020), .IN2(n9223), .Q(n11624) );
  INVX0 U11719 ( .INP(n11639), .ZN(n1020) );
  OR2X1 U11720 ( .IN1(n9569), .IN2(n3910), .Q(n11639) );
  OR4X1 U11721 ( .IN1(n11640), .IN2(n11641), .IN3(n11642), .IN4(n11643), .Q(
        WX5876) );
  AND2X1 U11722 ( .IN1(n11644), .IN2(n9173), .Q(n11643) );
  AND2X1 U11723 ( .IN1(n9277), .IN2(n10798), .Q(n11642) );
  OR2X1 U11724 ( .IN1(n11645), .IN2(n11646), .Q(n10798) );
  INVX0 U11725 ( .INP(n11647), .ZN(n11646) );
  OR2X1 U11726 ( .IN1(n11648), .IN2(n11649), .Q(n11647) );
  AND2X1 U11727 ( .IN1(n11649), .IN2(n11648), .Q(n11645) );
  AND2X1 U11728 ( .IN1(n11650), .IN2(n11651), .Q(n11648) );
  OR2X1 U11729 ( .IN1(WX7234), .IN2(n8211), .Q(n11651) );
  INVX0 U11730 ( .INP(n11652), .ZN(n11650) );
  AND2X1 U11731 ( .IN1(n8211), .IN2(WX7234), .Q(n11652) );
  OR2X1 U11732 ( .IN1(n11653), .IN2(n11654), .Q(n11649) );
  AND2X1 U11733 ( .IN1(n8212), .IN2(WX7362), .Q(n11654) );
  AND2X1 U11734 ( .IN1(n8846), .IN2(WX7298), .Q(n11653) );
  AND2X1 U11735 ( .IN1(n9247), .IN2(CRC_OUT_5_1), .Q(n11641) );
  AND2X1 U11736 ( .IN1(n1019), .IN2(n9222), .Q(n11640) );
  INVX0 U11737 ( .INP(n11655), .ZN(n1019) );
  OR2X1 U11738 ( .IN1(n9569), .IN2(n3911), .Q(n11655) );
  OR4X1 U11739 ( .IN1(n11656), .IN2(n11657), .IN3(n11658), .IN4(n11659), .Q(
        WX5874) );
  AND2X1 U11740 ( .IN1(n9195), .IN2(n11660), .Q(n11659) );
  AND2X1 U11741 ( .IN1(n9277), .IN2(n10814), .Q(n11658) );
  OR2X1 U11742 ( .IN1(n11661), .IN2(n11662), .Q(n10814) );
  INVX0 U11743 ( .INP(n11663), .ZN(n11662) );
  OR2X1 U11744 ( .IN1(n11664), .IN2(n11665), .Q(n11663) );
  AND2X1 U11745 ( .IN1(n11665), .IN2(n11664), .Q(n11661) );
  AND2X1 U11746 ( .IN1(n11666), .IN2(n11667), .Q(n11664) );
  OR2X1 U11747 ( .IN1(WX7232), .IN2(n8213), .Q(n11667) );
  INVX0 U11748 ( .INP(n11668), .ZN(n11666) );
  AND2X1 U11749 ( .IN1(n8213), .IN2(WX7232), .Q(n11668) );
  OR2X1 U11750 ( .IN1(n11669), .IN2(n11670), .Q(n11665) );
  AND2X1 U11751 ( .IN1(n8214), .IN2(WX7360), .Q(n11670) );
  AND2X1 U11752 ( .IN1(n8845), .IN2(WX7296), .Q(n11669) );
  AND2X1 U11753 ( .IN1(n9247), .IN2(CRC_OUT_5_2), .Q(n11657) );
  AND2X1 U11754 ( .IN1(n1018), .IN2(n9223), .Q(n11656) );
  INVX0 U11755 ( .INP(n11671), .ZN(n1018) );
  OR2X1 U11756 ( .IN1(n9569), .IN2(n3912), .Q(n11671) );
  OR4X1 U11757 ( .IN1(n11672), .IN2(n11673), .IN3(n11674), .IN4(n11675), .Q(
        WX5872) );
  AND2X1 U11758 ( .IN1(n11676), .IN2(n9173), .Q(n11675) );
  AND2X1 U11759 ( .IN1(n9277), .IN2(n10830), .Q(n11674) );
  OR2X1 U11760 ( .IN1(n11677), .IN2(n11678), .Q(n10830) );
  INVX0 U11761 ( .INP(n11679), .ZN(n11678) );
  OR2X1 U11762 ( .IN1(n11680), .IN2(n11681), .Q(n11679) );
  AND2X1 U11763 ( .IN1(n11681), .IN2(n11680), .Q(n11677) );
  AND2X1 U11764 ( .IN1(n11682), .IN2(n11683), .Q(n11680) );
  OR2X1 U11765 ( .IN1(WX7230), .IN2(n8215), .Q(n11683) );
  INVX0 U11766 ( .INP(n11684), .ZN(n11682) );
  AND2X1 U11767 ( .IN1(n8215), .IN2(WX7230), .Q(n11684) );
  OR2X1 U11768 ( .IN1(n11685), .IN2(n11686), .Q(n11681) );
  AND2X1 U11769 ( .IN1(n8216), .IN2(WX7358), .Q(n11686) );
  AND2X1 U11770 ( .IN1(n8844), .IN2(WX7294), .Q(n11685) );
  AND2X1 U11771 ( .IN1(n9247), .IN2(CRC_OUT_5_3), .Q(n11673) );
  AND2X1 U11772 ( .IN1(n1017), .IN2(n9223), .Q(n11672) );
  INVX0 U11773 ( .INP(n11687), .ZN(n1017) );
  OR2X1 U11774 ( .IN1(n9569), .IN2(n3913), .Q(n11687) );
  OR4X1 U11775 ( .IN1(n11688), .IN2(n11689), .IN3(n11690), .IN4(n11691), .Q(
        WX5870) );
  AND2X1 U11776 ( .IN1(n9195), .IN2(n11692), .Q(n11691) );
  AND2X1 U11777 ( .IN1(n10846), .IN2(n9258), .Q(n11690) );
  AND2X1 U11778 ( .IN1(n11693), .IN2(n11694), .Q(n10846) );
  INVX0 U11779 ( .INP(n11695), .ZN(n11694) );
  AND2X1 U11780 ( .IN1(n11696), .IN2(n11697), .Q(n11695) );
  OR2X1 U11781 ( .IN1(n11697), .IN2(n11696), .Q(n11693) );
  OR2X1 U11782 ( .IN1(n11698), .IN2(n11699), .Q(n11696) );
  INVX0 U11783 ( .INP(n11700), .ZN(n11699) );
  OR2X1 U11784 ( .IN1(WX7228), .IN2(n8217), .Q(n11700) );
  AND2X1 U11785 ( .IN1(n8217), .IN2(WX7228), .Q(n11698) );
  AND2X1 U11786 ( .IN1(n11701), .IN2(n11702), .Q(n11697) );
  OR2X1 U11787 ( .IN1(WX7292), .IN2(test_so64), .Q(n11702) );
  OR2X1 U11788 ( .IN1(n9087), .IN2(n8218), .Q(n11701) );
  AND2X1 U11789 ( .IN1(n9248), .IN2(CRC_OUT_5_4), .Q(n11689) );
  AND2X1 U11790 ( .IN1(n1016), .IN2(n9223), .Q(n11688) );
  INVX0 U11791 ( .INP(n11703), .ZN(n1016) );
  OR2X1 U11792 ( .IN1(n9569), .IN2(n3914), .Q(n11703) );
  OR4X1 U11793 ( .IN1(n11704), .IN2(n11705), .IN3(n11706), .IN4(n11707), .Q(
        WX5868) );
  AND2X1 U11794 ( .IN1(n11708), .IN2(n9173), .Q(n11707) );
  AND2X1 U11795 ( .IN1(n9278), .IN2(n10862), .Q(n11706) );
  OR2X1 U11796 ( .IN1(n11709), .IN2(n11710), .Q(n10862) );
  INVX0 U11797 ( .INP(n11711), .ZN(n11710) );
  OR2X1 U11798 ( .IN1(n11712), .IN2(n11713), .Q(n11711) );
  AND2X1 U11799 ( .IN1(n11713), .IN2(n11712), .Q(n11709) );
  AND2X1 U11800 ( .IN1(n11714), .IN2(n11715), .Q(n11712) );
  OR2X1 U11801 ( .IN1(WX7226), .IN2(n8219), .Q(n11715) );
  INVX0 U11802 ( .INP(n11716), .ZN(n11714) );
  AND2X1 U11803 ( .IN1(n8219), .IN2(WX7226), .Q(n11716) );
  OR2X1 U11804 ( .IN1(n11717), .IN2(n11718), .Q(n11713) );
  AND2X1 U11805 ( .IN1(n8220), .IN2(WX7354), .Q(n11718) );
  AND2X1 U11806 ( .IN1(n8843), .IN2(WX7290), .Q(n11717) );
  AND2X1 U11807 ( .IN1(n9248), .IN2(CRC_OUT_5_5), .Q(n11705) );
  AND2X1 U11808 ( .IN1(n1015), .IN2(n9223), .Q(n11704) );
  INVX0 U11809 ( .INP(n11719), .ZN(n1015) );
  OR2X1 U11810 ( .IN1(n9569), .IN2(n3915), .Q(n11719) );
  OR4X1 U11811 ( .IN1(n11720), .IN2(n11721), .IN3(n11722), .IN4(n11723), .Q(
        WX5866) );
  AND2X1 U11812 ( .IN1(n9195), .IN2(n11724), .Q(n11723) );
  AND2X1 U11813 ( .IN1(n10878), .IN2(n9258), .Q(n11722) );
  AND2X1 U11814 ( .IN1(n11725), .IN2(n11726), .Q(n10878) );
  INVX0 U11815 ( .INP(n11727), .ZN(n11726) );
  AND2X1 U11816 ( .IN1(n11728), .IN2(n11729), .Q(n11727) );
  OR2X1 U11817 ( .IN1(n11729), .IN2(n11728), .Q(n11725) );
  OR2X1 U11818 ( .IN1(n11730), .IN2(n11731), .Q(n11728) );
  INVX0 U11819 ( .INP(n11732), .ZN(n11731) );
  OR2X1 U11820 ( .IN1(WX7224), .IN2(n8221), .Q(n11732) );
  AND2X1 U11821 ( .IN1(n8221), .IN2(WX7224), .Q(n11730) );
  AND2X1 U11822 ( .IN1(n11733), .IN2(n11734), .Q(n11729) );
  OR2X1 U11823 ( .IN1(WX7352), .IN2(test_so62), .Q(n11734) );
  OR2X1 U11824 ( .IN1(n9120), .IN2(n8842), .Q(n11733) );
  AND2X1 U11825 ( .IN1(n9248), .IN2(CRC_OUT_5_6), .Q(n11721) );
  AND2X1 U11826 ( .IN1(n1014), .IN2(n9223), .Q(n11720) );
  INVX0 U11827 ( .INP(n11735), .ZN(n1014) );
  OR2X1 U11828 ( .IN1(n9569), .IN2(n3916), .Q(n11735) );
  OR4X1 U11829 ( .IN1(n11736), .IN2(n11737), .IN3(n11738), .IN4(n11739), .Q(
        WX5864) );
  AND2X1 U11830 ( .IN1(n9195), .IN2(n11740), .Q(n11739) );
  AND2X1 U11831 ( .IN1(n9278), .IN2(n10894), .Q(n11738) );
  OR2X1 U11832 ( .IN1(n11741), .IN2(n11742), .Q(n10894) );
  INVX0 U11833 ( .INP(n11743), .ZN(n11742) );
  OR2X1 U11834 ( .IN1(n11744), .IN2(n11745), .Q(n11743) );
  AND2X1 U11835 ( .IN1(n11745), .IN2(n11744), .Q(n11741) );
  AND2X1 U11836 ( .IN1(n11746), .IN2(n11747), .Q(n11744) );
  OR2X1 U11837 ( .IN1(WX7222), .IN2(n8222), .Q(n11747) );
  INVX0 U11838 ( .INP(n11748), .ZN(n11746) );
  AND2X1 U11839 ( .IN1(n8222), .IN2(WX7222), .Q(n11748) );
  OR2X1 U11840 ( .IN1(n11749), .IN2(n11750), .Q(n11745) );
  AND2X1 U11841 ( .IN1(n8223), .IN2(WX7350), .Q(n11750) );
  AND2X1 U11842 ( .IN1(n8841), .IN2(WX7286), .Q(n11749) );
  AND2X1 U11843 ( .IN1(n9248), .IN2(CRC_OUT_5_7), .Q(n11737) );
  AND2X1 U11844 ( .IN1(n1013), .IN2(n9223), .Q(n11736) );
  INVX0 U11845 ( .INP(n11751), .ZN(n1013) );
  OR2X1 U11846 ( .IN1(n9569), .IN2(n3917), .Q(n11751) );
  OR4X1 U11847 ( .IN1(n11752), .IN2(n11753), .IN3(n11754), .IN4(n11755), .Q(
        WX5862) );
  AND2X1 U11848 ( .IN1(n9194), .IN2(n11756), .Q(n11755) );
  AND2X1 U11849 ( .IN1(n10910), .IN2(n9257), .Q(n11754) );
  AND2X1 U11850 ( .IN1(n11757), .IN2(n11758), .Q(n10910) );
  INVX0 U11851 ( .INP(n11759), .ZN(n11758) );
  AND2X1 U11852 ( .IN1(n11760), .IN2(n11761), .Q(n11759) );
  OR2X1 U11853 ( .IN1(n11761), .IN2(n11760), .Q(n11757) );
  OR2X1 U11854 ( .IN1(n11762), .IN2(n11763), .Q(n11760) );
  INVX0 U11855 ( .INP(n11764), .ZN(n11763) );
  OR2X1 U11856 ( .IN1(WX7156), .IN2(n8225), .Q(n11764) );
  AND2X1 U11857 ( .IN1(n8225), .IN2(WX7156), .Q(n11762) );
  AND2X1 U11858 ( .IN1(n11765), .IN2(n11766), .Q(n11761) );
  OR2X1 U11859 ( .IN1(WX7348), .IN2(test_so60), .Q(n11766) );
  OR2X1 U11860 ( .IN1(n9121), .IN2(n8840), .Q(n11765) );
  AND2X1 U11861 ( .IN1(n9248), .IN2(CRC_OUT_5_8), .Q(n11753) );
  AND2X1 U11862 ( .IN1(n1012), .IN2(n9223), .Q(n11752) );
  INVX0 U11863 ( .INP(n11767), .ZN(n1012) );
  OR2X1 U11864 ( .IN1(n9569), .IN2(n3918), .Q(n11767) );
  OR4X1 U11865 ( .IN1(n11768), .IN2(n11769), .IN3(n11770), .IN4(n11771), .Q(
        WX5860) );
  AND2X1 U11866 ( .IN1(n9194), .IN2(n11772), .Q(n11771) );
  AND2X1 U11867 ( .IN1(n9278), .IN2(n10926), .Q(n11770) );
  OR2X1 U11868 ( .IN1(n11773), .IN2(n11774), .Q(n10926) );
  INVX0 U11869 ( .INP(n11775), .ZN(n11774) );
  OR2X1 U11870 ( .IN1(n11776), .IN2(n11777), .Q(n11775) );
  AND2X1 U11871 ( .IN1(n11777), .IN2(n11776), .Q(n11773) );
  AND2X1 U11872 ( .IN1(n11778), .IN2(n11779), .Q(n11776) );
  OR2X1 U11873 ( .IN1(WX7218), .IN2(n8226), .Q(n11779) );
  INVX0 U11874 ( .INP(n11780), .ZN(n11778) );
  AND2X1 U11875 ( .IN1(n8226), .IN2(WX7218), .Q(n11780) );
  OR2X1 U11876 ( .IN1(n11781), .IN2(n11782), .Q(n11777) );
  AND2X1 U11877 ( .IN1(n8227), .IN2(WX7346), .Q(n11782) );
  AND2X1 U11878 ( .IN1(n8839), .IN2(WX7282), .Q(n11781) );
  AND2X1 U11879 ( .IN1(n9248), .IN2(CRC_OUT_5_9), .Q(n11769) );
  AND2X1 U11880 ( .IN1(n1011), .IN2(n9223), .Q(n11768) );
  INVX0 U11881 ( .INP(n11783), .ZN(n1011) );
  OR2X1 U11882 ( .IN1(n9569), .IN2(n3919), .Q(n11783) );
  OR4X1 U11883 ( .IN1(n11784), .IN2(n11785), .IN3(n11786), .IN4(n11787), .Q(
        WX5858) );
  AND2X1 U11884 ( .IN1(n9194), .IN2(n11788), .Q(n11787) );
  AND2X1 U11885 ( .IN1(n10942), .IN2(n9257), .Q(n11786) );
  AND2X1 U11886 ( .IN1(n11789), .IN2(n11790), .Q(n10942) );
  INVX0 U11887 ( .INP(n11791), .ZN(n11790) );
  AND2X1 U11888 ( .IN1(n11792), .IN2(n11793), .Q(n11791) );
  OR2X1 U11889 ( .IN1(n11793), .IN2(n11792), .Q(n11789) );
  OR2X1 U11890 ( .IN1(n11794), .IN2(n11795), .Q(n11792) );
  INVX0 U11891 ( .INP(n11796), .ZN(n11795) );
  OR2X1 U11892 ( .IN1(WX7216), .IN2(n8228), .Q(n11796) );
  AND2X1 U11893 ( .IN1(n8228), .IN2(WX7216), .Q(n11794) );
  AND2X1 U11894 ( .IN1(n11797), .IN2(n11798), .Q(n11793) );
  OR2X1 U11895 ( .IN1(WX7344), .IN2(test_so58), .Q(n11798) );
  OR2X1 U11896 ( .IN1(n9122), .IN2(n8838), .Q(n11797) );
  AND2X1 U11897 ( .IN1(n9248), .IN2(CRC_OUT_5_10), .Q(n11785) );
  AND2X1 U11898 ( .IN1(n1010), .IN2(n9223), .Q(n11784) );
  INVX0 U11899 ( .INP(n11799), .ZN(n1010) );
  OR2X1 U11900 ( .IN1(n9569), .IN2(n3920), .Q(n11799) );
  OR4X1 U11901 ( .IN1(n11800), .IN2(n11801), .IN3(n11802), .IN4(n11803), .Q(
        WX5856) );
  AND2X1 U11902 ( .IN1(n9194), .IN2(n11804), .Q(n11803) );
  AND2X1 U11903 ( .IN1(n9278), .IN2(n10958), .Q(n11802) );
  OR2X1 U11904 ( .IN1(n11805), .IN2(n11806), .Q(n10958) );
  INVX0 U11905 ( .INP(n11807), .ZN(n11806) );
  OR2X1 U11906 ( .IN1(n11808), .IN2(n11809), .Q(n11807) );
  AND2X1 U11907 ( .IN1(n11809), .IN2(n11808), .Q(n11805) );
  AND2X1 U11908 ( .IN1(n11810), .IN2(n11811), .Q(n11808) );
  OR2X1 U11909 ( .IN1(WX7214), .IN2(n8229), .Q(n11811) );
  INVX0 U11910 ( .INP(n11812), .ZN(n11810) );
  AND2X1 U11911 ( .IN1(n8229), .IN2(WX7214), .Q(n11812) );
  OR2X1 U11912 ( .IN1(n11813), .IN2(n11814), .Q(n11809) );
  AND2X1 U11913 ( .IN1(n8230), .IN2(WX7342), .Q(n11814) );
  AND2X1 U11914 ( .IN1(n8723), .IN2(WX7278), .Q(n11813) );
  AND2X1 U11915 ( .IN1(n9248), .IN2(CRC_OUT_5_11), .Q(n11801) );
  AND2X1 U11916 ( .IN1(n1009), .IN2(n9223), .Q(n11800) );
  INVX0 U11917 ( .INP(n11815), .ZN(n1009) );
  OR2X1 U11918 ( .IN1(n9568), .IN2(n3921), .Q(n11815) );
  OR4X1 U11919 ( .IN1(n11816), .IN2(n11817), .IN3(n11818), .IN4(n11819), .Q(
        WX5854) );
  AND2X1 U11920 ( .IN1(n9194), .IN2(n11820), .Q(n11819) );
  AND2X1 U11921 ( .IN1(n9278), .IN2(n10974), .Q(n11818) );
  OR2X1 U11922 ( .IN1(n11821), .IN2(n11822), .Q(n10974) );
  INVX0 U11923 ( .INP(n11823), .ZN(n11822) );
  OR2X1 U11924 ( .IN1(n11824), .IN2(n11825), .Q(n11823) );
  AND2X1 U11925 ( .IN1(n11825), .IN2(n11824), .Q(n11821) );
  AND2X1 U11926 ( .IN1(n11826), .IN2(n11827), .Q(n11824) );
  OR2X1 U11927 ( .IN1(WX7212), .IN2(n8231), .Q(n11827) );
  INVX0 U11928 ( .INP(n11828), .ZN(n11826) );
  AND2X1 U11929 ( .IN1(n8231), .IN2(WX7212), .Q(n11828) );
  OR2X1 U11930 ( .IN1(n11829), .IN2(n11830), .Q(n11825) );
  AND2X1 U11931 ( .IN1(n8232), .IN2(WX7340), .Q(n11830) );
  AND2X1 U11932 ( .IN1(n8837), .IN2(WX7276), .Q(n11829) );
  AND2X1 U11933 ( .IN1(n9248), .IN2(CRC_OUT_5_12), .Q(n11817) );
  AND2X1 U11934 ( .IN1(n1008), .IN2(n9224), .Q(n11816) );
  INVX0 U11935 ( .INP(n11831), .ZN(n1008) );
  OR2X1 U11936 ( .IN1(n9568), .IN2(n3922), .Q(n11831) );
  OR4X1 U11937 ( .IN1(n11832), .IN2(n11833), .IN3(n11834), .IN4(n11835), .Q(
        WX5852) );
  AND2X1 U11938 ( .IN1(n9194), .IN2(n11836), .Q(n11835) );
  AND2X1 U11939 ( .IN1(n9278), .IN2(n10990), .Q(n11834) );
  OR2X1 U11940 ( .IN1(n11837), .IN2(n11838), .Q(n10990) );
  INVX0 U11941 ( .INP(n11839), .ZN(n11838) );
  OR2X1 U11942 ( .IN1(n11840), .IN2(n11841), .Q(n11839) );
  AND2X1 U11943 ( .IN1(n11841), .IN2(n11840), .Q(n11837) );
  AND2X1 U11944 ( .IN1(n11842), .IN2(n11843), .Q(n11840) );
  OR2X1 U11945 ( .IN1(WX7210), .IN2(n8233), .Q(n11843) );
  INVX0 U11946 ( .INP(n11844), .ZN(n11842) );
  AND2X1 U11947 ( .IN1(n8233), .IN2(WX7210), .Q(n11844) );
  OR2X1 U11948 ( .IN1(n11845), .IN2(n11846), .Q(n11841) );
  AND2X1 U11949 ( .IN1(n8234), .IN2(WX7338), .Q(n11846) );
  AND2X1 U11950 ( .IN1(n8836), .IN2(WX7274), .Q(n11845) );
  AND2X1 U11951 ( .IN1(n9248), .IN2(CRC_OUT_5_13), .Q(n11833) );
  AND2X1 U11952 ( .IN1(n1007), .IN2(n9223), .Q(n11832) );
  INVX0 U11953 ( .INP(n11847), .ZN(n1007) );
  OR2X1 U11954 ( .IN1(n9568), .IN2(n3923), .Q(n11847) );
  OR4X1 U11955 ( .IN1(n11848), .IN2(n11849), .IN3(n11850), .IN4(n11851), .Q(
        WX5850) );
  AND2X1 U11956 ( .IN1(n9194), .IN2(n11852), .Q(n11851) );
  AND2X1 U11957 ( .IN1(n9278), .IN2(n11006), .Q(n11850) );
  OR2X1 U11958 ( .IN1(n11853), .IN2(n11854), .Q(n11006) );
  INVX0 U11959 ( .INP(n11855), .ZN(n11854) );
  OR2X1 U11960 ( .IN1(n11856), .IN2(n11857), .Q(n11855) );
  AND2X1 U11961 ( .IN1(n11857), .IN2(n11856), .Q(n11853) );
  AND2X1 U11962 ( .IN1(n11858), .IN2(n11859), .Q(n11856) );
  OR2X1 U11963 ( .IN1(WX7208), .IN2(n8235), .Q(n11859) );
  INVX0 U11964 ( .INP(n11860), .ZN(n11858) );
  AND2X1 U11965 ( .IN1(n8235), .IN2(WX7208), .Q(n11860) );
  OR2X1 U11966 ( .IN1(n11861), .IN2(n11862), .Q(n11857) );
  AND2X1 U11967 ( .IN1(n8236), .IN2(WX7336), .Q(n11862) );
  AND2X1 U11968 ( .IN1(n8835), .IN2(WX7272), .Q(n11861) );
  AND2X1 U11969 ( .IN1(n9248), .IN2(CRC_OUT_5_14), .Q(n11849) );
  AND2X1 U11970 ( .IN1(n1006), .IN2(n9224), .Q(n11848) );
  INVX0 U11971 ( .INP(n11863), .ZN(n1006) );
  OR2X1 U11972 ( .IN1(n9568), .IN2(n3924), .Q(n11863) );
  OR4X1 U11973 ( .IN1(n11864), .IN2(n11865), .IN3(n11866), .IN4(n11867), .Q(
        WX5848) );
  AND2X1 U11974 ( .IN1(n9194), .IN2(n11868), .Q(n11867) );
  AND2X1 U11975 ( .IN1(n9278), .IN2(n11022), .Q(n11866) );
  OR2X1 U11976 ( .IN1(n11869), .IN2(n11870), .Q(n11022) );
  INVX0 U11977 ( .INP(n11871), .ZN(n11870) );
  OR2X1 U11978 ( .IN1(n11872), .IN2(n11873), .Q(n11871) );
  AND2X1 U11979 ( .IN1(n11873), .IN2(n11872), .Q(n11869) );
  AND2X1 U11980 ( .IN1(n11874), .IN2(n11875), .Q(n11872) );
  OR2X1 U11981 ( .IN1(WX7206), .IN2(n8237), .Q(n11875) );
  INVX0 U11982 ( .INP(n11876), .ZN(n11874) );
  AND2X1 U11983 ( .IN1(n8237), .IN2(WX7206), .Q(n11876) );
  OR2X1 U11984 ( .IN1(n11877), .IN2(n11878), .Q(n11873) );
  AND2X1 U11985 ( .IN1(n8238), .IN2(WX7334), .Q(n11878) );
  AND2X1 U11986 ( .IN1(n8834), .IN2(WX7270), .Q(n11877) );
  AND2X1 U11987 ( .IN1(n9248), .IN2(CRC_OUT_5_15), .Q(n11865) );
  AND2X1 U11988 ( .IN1(n1005), .IN2(n9206), .Q(n11864) );
  INVX0 U11989 ( .INP(n11879), .ZN(n1005) );
  OR2X1 U11990 ( .IN1(n9568), .IN2(n3925), .Q(n11879) );
  OR4X1 U11991 ( .IN1(n11880), .IN2(n11881), .IN3(n11882), .IN4(n11883), .Q(
        WX5846) );
  AND2X1 U11992 ( .IN1(n11884), .IN2(n9175), .Q(n11883) );
  AND2X1 U11993 ( .IN1(n9278), .IN2(n11038), .Q(n11882) );
  OR2X1 U11994 ( .IN1(n11885), .IN2(n11886), .Q(n11038) );
  INVX0 U11995 ( .INP(n11887), .ZN(n11886) );
  OR2X1 U11996 ( .IN1(n11888), .IN2(n11889), .Q(n11887) );
  AND2X1 U11997 ( .IN1(n11889), .IN2(n11888), .Q(n11885) );
  AND2X1 U11998 ( .IN1(n11890), .IN2(n11891), .Q(n11888) );
  OR2X1 U11999 ( .IN1(n9461), .IN2(n7976), .Q(n11891) );
  OR2X1 U12000 ( .IN1(WX7204), .IN2(n9448), .Q(n11890) );
  OR2X1 U12001 ( .IN1(n11892), .IN2(n11893), .Q(n11889) );
  INVX0 U12002 ( .INP(n11894), .ZN(n11893) );
  OR2X1 U12003 ( .IN1(n11895), .IN2(n7977), .Q(n11894) );
  AND2X1 U12004 ( .IN1(n7977), .IN2(n11895), .Q(n11892) );
  INVX0 U12005 ( .INP(n11896), .ZN(n11895) );
  OR2X1 U12006 ( .IN1(n11897), .IN2(n11898), .Q(n11896) );
  AND2X1 U12007 ( .IN1(n8722), .IN2(n8421), .Q(n11898) );
  AND2X1 U12008 ( .IN1(n15908), .IN2(WX7332), .Q(n11897) );
  AND2X1 U12009 ( .IN1(n9248), .IN2(CRC_OUT_5_16), .Q(n11881) );
  AND2X1 U12010 ( .IN1(n1004), .IN2(n9201), .Q(n11880) );
  INVX0 U12011 ( .INP(n11899), .ZN(n1004) );
  OR2X1 U12012 ( .IN1(n9568), .IN2(n3926), .Q(n11899) );
  OR4X1 U12013 ( .IN1(n11900), .IN2(n11901), .IN3(n11902), .IN4(n11903), .Q(
        WX5844) );
  AND2X1 U12014 ( .IN1(n9194), .IN2(n11904), .Q(n11903) );
  AND2X1 U12015 ( .IN1(n9278), .IN2(n11058), .Q(n11902) );
  OR2X1 U12016 ( .IN1(n11905), .IN2(n11906), .Q(n11058) );
  INVX0 U12017 ( .INP(n11907), .ZN(n11906) );
  OR2X1 U12018 ( .IN1(n11908), .IN2(n11909), .Q(n11907) );
  AND2X1 U12019 ( .IN1(n11909), .IN2(n11908), .Q(n11905) );
  AND2X1 U12020 ( .IN1(n11910), .IN2(n11911), .Q(n11908) );
  OR2X1 U12021 ( .IN1(n9458), .IN2(n7978), .Q(n11911) );
  OR2X1 U12022 ( .IN1(WX7202), .IN2(n9448), .Q(n11910) );
  OR2X1 U12023 ( .IN1(n11912), .IN2(n11913), .Q(n11909) );
  INVX0 U12024 ( .INP(n11914), .ZN(n11913) );
  OR2X1 U12025 ( .IN1(n11915), .IN2(n7979), .Q(n11914) );
  AND2X1 U12026 ( .IN1(n7979), .IN2(n11915), .Q(n11912) );
  INVX0 U12027 ( .INP(n11916), .ZN(n11915) );
  OR2X1 U12028 ( .IN1(n11917), .IN2(n11918), .Q(n11916) );
  AND2X1 U12029 ( .IN1(n8833), .IN2(n8422), .Q(n11918) );
  AND2X1 U12030 ( .IN1(n15909), .IN2(WX7330), .Q(n11917) );
  AND2X1 U12031 ( .IN1(test_so54), .IN2(n9227), .Q(n11901) );
  AND2X1 U12032 ( .IN1(n1003), .IN2(n9201), .Q(n11900) );
  INVX0 U12033 ( .INP(n11919), .ZN(n1003) );
  OR2X1 U12034 ( .IN1(n9568), .IN2(n3927), .Q(n11919) );
  OR4X1 U12035 ( .IN1(n11920), .IN2(n11921), .IN3(n11922), .IN4(n11923), .Q(
        WX5842) );
  AND2X1 U12036 ( .IN1(n11924), .IN2(n9175), .Q(n11923) );
  AND2X1 U12037 ( .IN1(n9278), .IN2(n11078), .Q(n11922) );
  OR2X1 U12038 ( .IN1(n11925), .IN2(n11926), .Q(n11078) );
  INVX0 U12039 ( .INP(n11927), .ZN(n11926) );
  OR2X1 U12040 ( .IN1(n11928), .IN2(n11929), .Q(n11927) );
  AND2X1 U12041 ( .IN1(n11929), .IN2(n11928), .Q(n11925) );
  AND2X1 U12042 ( .IN1(n11930), .IN2(n11931), .Q(n11928) );
  OR2X1 U12043 ( .IN1(n9474), .IN2(n7980), .Q(n11931) );
  OR2X1 U12044 ( .IN1(WX7200), .IN2(n9448), .Q(n11930) );
  OR2X1 U12045 ( .IN1(n11932), .IN2(n11933), .Q(n11929) );
  INVX0 U12046 ( .INP(n11934), .ZN(n11933) );
  OR2X1 U12047 ( .IN1(n11935), .IN2(n7981), .Q(n11934) );
  AND2X1 U12048 ( .IN1(n7981), .IN2(n11935), .Q(n11932) );
  INVX0 U12049 ( .INP(n11936), .ZN(n11935) );
  OR2X1 U12050 ( .IN1(n11937), .IN2(n11938), .Q(n11936) );
  AND2X1 U12051 ( .IN1(n8832), .IN2(n8423), .Q(n11938) );
  AND2X1 U12052 ( .IN1(n15910), .IN2(WX7328), .Q(n11937) );
  AND2X1 U12053 ( .IN1(n9249), .IN2(CRC_OUT_5_18), .Q(n11921) );
  AND2X1 U12054 ( .IN1(n1002), .IN2(n9201), .Q(n11920) );
  INVX0 U12055 ( .INP(n11939), .ZN(n1002) );
  OR2X1 U12056 ( .IN1(n9568), .IN2(n3928), .Q(n11939) );
  OR4X1 U12057 ( .IN1(n11940), .IN2(n11941), .IN3(n11942), .IN4(n11943), .Q(
        WX5840) );
  AND2X1 U12058 ( .IN1(n9194), .IN2(n11944), .Q(n11943) );
  AND2X1 U12059 ( .IN1(n9278), .IN2(n11098), .Q(n11942) );
  OR2X1 U12060 ( .IN1(n11945), .IN2(n11946), .Q(n11098) );
  INVX0 U12061 ( .INP(n11947), .ZN(n11946) );
  OR2X1 U12062 ( .IN1(n11948), .IN2(n11949), .Q(n11947) );
  AND2X1 U12063 ( .IN1(n11949), .IN2(n11948), .Q(n11945) );
  AND2X1 U12064 ( .IN1(n11950), .IN2(n11951), .Q(n11948) );
  OR2X1 U12065 ( .IN1(n9473), .IN2(n7982), .Q(n11951) );
  OR2X1 U12066 ( .IN1(WX7198), .IN2(n9448), .Q(n11950) );
  OR2X1 U12067 ( .IN1(n11952), .IN2(n11953), .Q(n11949) );
  INVX0 U12068 ( .INP(n11954), .ZN(n11953) );
  OR2X1 U12069 ( .IN1(n11955), .IN2(n7983), .Q(n11954) );
  AND2X1 U12070 ( .IN1(n7983), .IN2(n11955), .Q(n11952) );
  INVX0 U12071 ( .INP(n11956), .ZN(n11955) );
  OR2X1 U12072 ( .IN1(n11957), .IN2(n11958), .Q(n11956) );
  AND2X1 U12073 ( .IN1(n8831), .IN2(n8424), .Q(n11958) );
  AND2X1 U12074 ( .IN1(n15911), .IN2(WX7326), .Q(n11957) );
  AND2X1 U12075 ( .IN1(n9249), .IN2(CRC_OUT_5_19), .Q(n11941) );
  AND2X1 U12076 ( .IN1(n1001), .IN2(n9201), .Q(n11940) );
  INVX0 U12077 ( .INP(n11959), .ZN(n1001) );
  OR2X1 U12078 ( .IN1(n9568), .IN2(n3929), .Q(n11959) );
  OR4X1 U12079 ( .IN1(n11960), .IN2(n11961), .IN3(n11962), .IN4(n11963), .Q(
        WX5838) );
  AND2X1 U12080 ( .IN1(n11964), .IN2(n9175), .Q(n11963) );
  AND2X1 U12081 ( .IN1(n9278), .IN2(n11118), .Q(n11962) );
  OR2X1 U12082 ( .IN1(n11965), .IN2(n11966), .Q(n11118) );
  INVX0 U12083 ( .INP(n11967), .ZN(n11966) );
  OR2X1 U12084 ( .IN1(n11968), .IN2(n11969), .Q(n11967) );
  AND2X1 U12085 ( .IN1(n11969), .IN2(n11968), .Q(n11965) );
  AND2X1 U12086 ( .IN1(n11970), .IN2(n11971), .Q(n11968) );
  OR2X1 U12087 ( .IN1(n9475), .IN2(n7984), .Q(n11971) );
  OR2X1 U12088 ( .IN1(WX7196), .IN2(n9447), .Q(n11970) );
  OR2X1 U12089 ( .IN1(n11972), .IN2(n11973), .Q(n11969) );
  INVX0 U12090 ( .INP(n11974), .ZN(n11973) );
  OR2X1 U12091 ( .IN1(n11975), .IN2(n7985), .Q(n11974) );
  AND2X1 U12092 ( .IN1(n7985), .IN2(n11975), .Q(n11972) );
  INVX0 U12093 ( .INP(n11976), .ZN(n11975) );
  OR2X1 U12094 ( .IN1(n11977), .IN2(n11978), .Q(n11976) );
  AND2X1 U12095 ( .IN1(n8830), .IN2(n8425), .Q(n11978) );
  AND2X1 U12096 ( .IN1(n15912), .IN2(WX7324), .Q(n11977) );
  AND2X1 U12097 ( .IN1(n9249), .IN2(CRC_OUT_5_20), .Q(n11961) );
  AND2X1 U12098 ( .IN1(n1000), .IN2(n9201), .Q(n11960) );
  INVX0 U12099 ( .INP(n11979), .ZN(n1000) );
  OR2X1 U12100 ( .IN1(n9568), .IN2(n3930), .Q(n11979) );
  OR4X1 U12101 ( .IN1(n11980), .IN2(n11981), .IN3(n11982), .IN4(n11983), .Q(
        WX5836) );
  AND2X1 U12102 ( .IN1(n9194), .IN2(n11984), .Q(n11983) );
  AND2X1 U12103 ( .IN1(n11138), .IN2(n9257), .Q(n11982) );
  AND2X1 U12104 ( .IN1(n11985), .IN2(n11986), .Q(n11138) );
  INVX0 U12105 ( .INP(n11987), .ZN(n11986) );
  AND2X1 U12106 ( .IN1(n11988), .IN2(n11989), .Q(n11987) );
  OR2X1 U12107 ( .IN1(n11989), .IN2(n11988), .Q(n11985) );
  OR2X1 U12108 ( .IN1(n11990), .IN2(n11991), .Q(n11988) );
  AND2X1 U12109 ( .IN1(n9451), .IN2(WX7194), .Q(n11991) );
  AND2X1 U12110 ( .IN1(n7986), .IN2(n9459), .Q(n11990) );
  AND2X1 U12111 ( .IN1(n11992), .IN2(n11993), .Q(n11989) );
  OR2X1 U12112 ( .IN1(n11994), .IN2(n7987), .Q(n11993) );
  INVX0 U12113 ( .INP(n11995), .ZN(n11994) );
  OR2X1 U12114 ( .IN1(WX7258), .IN2(n11995), .Q(n11992) );
  OR2X1 U12115 ( .IN1(n11996), .IN2(n11997), .Q(n11995) );
  AND2X1 U12116 ( .IN1(n15913), .IN2(n9105), .Q(n11997) );
  AND2X1 U12117 ( .IN1(test_so63), .IN2(n8426), .Q(n11996) );
  AND2X1 U12118 ( .IN1(n9233), .IN2(CRC_OUT_5_21), .Q(n11981) );
  AND2X1 U12119 ( .IN1(n999), .IN2(n9201), .Q(n11980) );
  INVX0 U12120 ( .INP(n11998), .ZN(n999) );
  OR2X1 U12121 ( .IN1(n9568), .IN2(n3931), .Q(n11998) );
  OR4X1 U12122 ( .IN1(n11999), .IN2(n12000), .IN3(n12001), .IN4(n12002), .Q(
        WX5834) );
  AND2X1 U12123 ( .IN1(n12003), .IN2(n9175), .Q(n12002) );
  AND2X1 U12124 ( .IN1(n9279), .IN2(n11158), .Q(n12001) );
  OR2X1 U12125 ( .IN1(n12004), .IN2(n12005), .Q(n11158) );
  INVX0 U12126 ( .INP(n12006), .ZN(n12005) );
  OR2X1 U12127 ( .IN1(n12007), .IN2(n12008), .Q(n12006) );
  AND2X1 U12128 ( .IN1(n12008), .IN2(n12007), .Q(n12004) );
  AND2X1 U12129 ( .IN1(n12009), .IN2(n12010), .Q(n12007) );
  OR2X1 U12130 ( .IN1(n9463), .IN2(n7988), .Q(n12010) );
  OR2X1 U12131 ( .IN1(WX7192), .IN2(n9448), .Q(n12009) );
  OR2X1 U12132 ( .IN1(n12011), .IN2(n12012), .Q(n12008) );
  INVX0 U12133 ( .INP(n12013), .ZN(n12012) );
  OR2X1 U12134 ( .IN1(n12014), .IN2(n7989), .Q(n12013) );
  AND2X1 U12135 ( .IN1(n7989), .IN2(n12014), .Q(n12011) );
  INVX0 U12136 ( .INP(n12015), .ZN(n12014) );
  OR2X1 U12137 ( .IN1(n12016), .IN2(n12017), .Q(n12015) );
  AND2X1 U12138 ( .IN1(n8829), .IN2(n8427), .Q(n12017) );
  AND2X1 U12139 ( .IN1(n15914), .IN2(WX7320), .Q(n12016) );
  AND2X1 U12140 ( .IN1(n9228), .IN2(CRC_OUT_5_22), .Q(n12000) );
  AND2X1 U12141 ( .IN1(n998), .IN2(n9201), .Q(n11999) );
  INVX0 U12142 ( .INP(n12018), .ZN(n998) );
  OR2X1 U12143 ( .IN1(n9568), .IN2(n3932), .Q(n12018) );
  OR4X1 U12144 ( .IN1(n12019), .IN2(n12020), .IN3(n12021), .IN4(n12022), .Q(
        WX5832) );
  AND2X1 U12145 ( .IN1(n9194), .IN2(n12023), .Q(n12022) );
  AND2X1 U12146 ( .IN1(n11178), .IN2(n9257), .Q(n12021) );
  AND2X1 U12147 ( .IN1(n12024), .IN2(n12025), .Q(n11178) );
  INVX0 U12148 ( .INP(n12026), .ZN(n12025) );
  AND2X1 U12149 ( .IN1(n12027), .IN2(n12028), .Q(n12026) );
  OR2X1 U12150 ( .IN1(n12028), .IN2(n12027), .Q(n12024) );
  OR2X1 U12151 ( .IN1(n12029), .IN2(n12030), .Q(n12027) );
  AND2X1 U12152 ( .IN1(n9450), .IN2(WX7190), .Q(n12030) );
  AND2X1 U12153 ( .IN1(n7990), .IN2(n9467), .Q(n12029) );
  AND2X1 U12154 ( .IN1(n12031), .IN2(n12032), .Q(n12028) );
  OR2X1 U12155 ( .IN1(n12033), .IN2(n8828), .Q(n12032) );
  OR2X1 U12156 ( .IN1(WX7318), .IN2(n12034), .Q(n12031) );
  INVX0 U12157 ( .INP(n12033), .ZN(n12034) );
  AND2X1 U12158 ( .IN1(n12035), .IN2(n12036), .Q(n12033) );
  OR2X1 U12159 ( .IN1(n8428), .IN2(test_so61), .Q(n12036) );
  OR2X1 U12160 ( .IN1(n9123), .IN2(n15915), .Q(n12035) );
  AND2X1 U12161 ( .IN1(n9230), .IN2(CRC_OUT_5_23), .Q(n12020) );
  AND2X1 U12162 ( .IN1(n997), .IN2(n9201), .Q(n12019) );
  INVX0 U12163 ( .INP(n12037), .ZN(n997) );
  OR2X1 U12164 ( .IN1(n9567), .IN2(n3933), .Q(n12037) );
  OR4X1 U12165 ( .IN1(n12038), .IN2(n12039), .IN3(n12040), .IN4(n12041), .Q(
        WX5830) );
  AND2X1 U12166 ( .IN1(n9194), .IN2(n12042), .Q(n12041) );
  AND2X1 U12167 ( .IN1(n9279), .IN2(n11198), .Q(n12040) );
  OR2X1 U12168 ( .IN1(n12043), .IN2(n12044), .Q(n11198) );
  INVX0 U12169 ( .INP(n12045), .ZN(n12044) );
  OR2X1 U12170 ( .IN1(n12046), .IN2(n12047), .Q(n12045) );
  AND2X1 U12171 ( .IN1(n12047), .IN2(n12046), .Q(n12043) );
  AND2X1 U12172 ( .IN1(n12048), .IN2(n12049), .Q(n12046) );
  OR2X1 U12173 ( .IN1(n9453), .IN2(n7991), .Q(n12049) );
  OR2X1 U12174 ( .IN1(WX7188), .IN2(n9447), .Q(n12048) );
  OR2X1 U12175 ( .IN1(n12050), .IN2(n12051), .Q(n12047) );
  INVX0 U12176 ( .INP(n12052), .ZN(n12051) );
  OR2X1 U12177 ( .IN1(n12053), .IN2(n7992), .Q(n12052) );
  AND2X1 U12178 ( .IN1(n7992), .IN2(n12053), .Q(n12050) );
  INVX0 U12179 ( .INP(n12054), .ZN(n12053) );
  OR2X1 U12180 ( .IN1(n12055), .IN2(n12056), .Q(n12054) );
  AND2X1 U12181 ( .IN1(n8827), .IN2(n8429), .Q(n12056) );
  AND2X1 U12182 ( .IN1(n15916), .IN2(WX7316), .Q(n12055) );
  AND2X1 U12183 ( .IN1(n9228), .IN2(CRC_OUT_5_24), .Q(n12039) );
  AND2X1 U12184 ( .IN1(n996), .IN2(n9201), .Q(n12038) );
  INVX0 U12185 ( .INP(n12057), .ZN(n996) );
  OR2X1 U12186 ( .IN1(n9567), .IN2(n3934), .Q(n12057) );
  OR4X1 U12187 ( .IN1(n12058), .IN2(n12059), .IN3(n12060), .IN4(n12061), .Q(
        WX5828) );
  AND2X1 U12188 ( .IN1(n9193), .IN2(n12062), .Q(n12061) );
  AND2X1 U12189 ( .IN1(n11218), .IN2(n9257), .Q(n12060) );
  AND2X1 U12190 ( .IN1(n12063), .IN2(n12064), .Q(n11218) );
  INVX0 U12191 ( .INP(n12065), .ZN(n12064) );
  AND2X1 U12192 ( .IN1(n12066), .IN2(n12067), .Q(n12065) );
  OR2X1 U12193 ( .IN1(n12067), .IN2(n12066), .Q(n12063) );
  OR2X1 U12194 ( .IN1(n12068), .IN2(n12069), .Q(n12066) );
  AND2X1 U12195 ( .IN1(n9450), .IN2(WX7250), .Q(n12069) );
  AND2X1 U12196 ( .IN1(n7993), .IN2(n9470), .Q(n12068) );
  AND2X1 U12197 ( .IN1(n12070), .IN2(n12071), .Q(n12067) );
  OR2X1 U12198 ( .IN1(n12072), .IN2(n8826), .Q(n12071) );
  OR2X1 U12199 ( .IN1(WX7314), .IN2(n12073), .Q(n12070) );
  INVX0 U12200 ( .INP(n12072), .ZN(n12073) );
  AND2X1 U12201 ( .IN1(n12074), .IN2(n12075), .Q(n12072) );
  OR2X1 U12202 ( .IN1(n8430), .IN2(test_so59), .Q(n12075) );
  OR2X1 U12203 ( .IN1(n9124), .IN2(n15917), .Q(n12074) );
  AND2X1 U12204 ( .IN1(n9229), .IN2(CRC_OUT_5_25), .Q(n12059) );
  AND2X1 U12205 ( .IN1(n995), .IN2(n9201), .Q(n12058) );
  INVX0 U12206 ( .INP(n12076), .ZN(n995) );
  OR2X1 U12207 ( .IN1(n9567), .IN2(n3935), .Q(n12076) );
  OR4X1 U12208 ( .IN1(n12077), .IN2(n12078), .IN3(n12079), .IN4(n12080), .Q(
        WX5826) );
  AND2X1 U12209 ( .IN1(n9193), .IN2(n12081), .Q(n12080) );
  AND2X1 U12210 ( .IN1(n9279), .IN2(n11239), .Q(n12079) );
  OR2X1 U12211 ( .IN1(n12082), .IN2(n12083), .Q(n11239) );
  INVX0 U12212 ( .INP(n12084), .ZN(n12083) );
  OR2X1 U12213 ( .IN1(n12085), .IN2(n12086), .Q(n12084) );
  AND2X1 U12214 ( .IN1(n12086), .IN2(n12085), .Q(n12082) );
  AND2X1 U12215 ( .IN1(n12087), .IN2(n12088), .Q(n12085) );
  OR2X1 U12216 ( .IN1(n9480), .IN2(n7994), .Q(n12088) );
  OR2X1 U12217 ( .IN1(WX7184), .IN2(n9447), .Q(n12087) );
  OR2X1 U12218 ( .IN1(n12089), .IN2(n12090), .Q(n12086) );
  INVX0 U12219 ( .INP(n12091), .ZN(n12090) );
  OR2X1 U12220 ( .IN1(n12092), .IN2(n7995), .Q(n12091) );
  AND2X1 U12221 ( .IN1(n7995), .IN2(n12092), .Q(n12089) );
  INVX0 U12222 ( .INP(n12093), .ZN(n12092) );
  OR2X1 U12223 ( .IN1(n12094), .IN2(n12095), .Q(n12093) );
  AND2X1 U12224 ( .IN1(n8825), .IN2(n8431), .Q(n12095) );
  AND2X1 U12225 ( .IN1(n15918), .IN2(WX7312), .Q(n12094) );
  AND2X1 U12226 ( .IN1(n9228), .IN2(CRC_OUT_5_26), .Q(n12078) );
  AND2X1 U12227 ( .IN1(n994), .IN2(n9201), .Q(n12077) );
  INVX0 U12228 ( .INP(n12096), .ZN(n994) );
  OR2X1 U12229 ( .IN1(n9567), .IN2(n3936), .Q(n12096) );
  OR4X1 U12230 ( .IN1(n12097), .IN2(n12098), .IN3(n12099), .IN4(n12100), .Q(
        WX5824) );
  AND2X1 U12231 ( .IN1(n9193), .IN2(n12101), .Q(n12100) );
  AND2X1 U12232 ( .IN1(n11258), .IN2(n9257), .Q(n12099) );
  AND2X1 U12233 ( .IN1(n12102), .IN2(n12103), .Q(n11258) );
  OR2X1 U12234 ( .IN1(n12104), .IN2(n12105), .Q(n12103) );
  INVX0 U12235 ( .INP(n12106), .ZN(n12102) );
  AND2X1 U12236 ( .IN1(n12105), .IN2(n12104), .Q(n12106) );
  INVX0 U12237 ( .INP(n12107), .ZN(n12104) );
  OR2X1 U12238 ( .IN1(n12108), .IN2(n12109), .Q(n12107) );
  AND2X1 U12239 ( .IN1(n9450), .IN2(WX7310), .Q(n12109) );
  AND2X1 U12240 ( .IN1(n8824), .IN2(n9464), .Q(n12108) );
  OR2X1 U12241 ( .IN1(n12110), .IN2(n12111), .Q(n12105) );
  AND3X1 U12242 ( .IN1(n12112), .IN2(n12113), .IN3(n7997), .Q(n12111) );
  OR2X1 U12243 ( .IN1(n7996), .IN2(n9092), .Q(n12113) );
  OR2X1 U12244 ( .IN1(test_so57), .IN2(WX7182), .Q(n12112) );
  AND2X1 U12245 ( .IN1(n12114), .IN2(WX7246), .Q(n12110) );
  OR2X1 U12246 ( .IN1(n12115), .IN2(n12116), .Q(n12114) );
  AND2X1 U12247 ( .IN1(n7996), .IN2(n9092), .Q(n12116) );
  AND2X1 U12248 ( .IN1(test_so57), .IN2(WX7182), .Q(n12115) );
  AND2X1 U12249 ( .IN1(n9229), .IN2(CRC_OUT_5_27), .Q(n12098) );
  AND2X1 U12250 ( .IN1(n993), .IN2(n9202), .Q(n12097) );
  INVX0 U12251 ( .INP(n12117), .ZN(n993) );
  OR2X1 U12252 ( .IN1(n9567), .IN2(n3937), .Q(n12117) );
  OR4X1 U12253 ( .IN1(n12118), .IN2(n12119), .IN3(n12120), .IN4(n12121), .Q(
        WX5822) );
  AND2X1 U12254 ( .IN1(n9193), .IN2(n12122), .Q(n12121) );
  AND2X1 U12255 ( .IN1(n9279), .IN2(n11278), .Q(n12120) );
  OR2X1 U12256 ( .IN1(n12123), .IN2(n12124), .Q(n11278) );
  INVX0 U12257 ( .INP(n12125), .ZN(n12124) );
  OR2X1 U12258 ( .IN1(n12126), .IN2(n12127), .Q(n12125) );
  AND2X1 U12259 ( .IN1(n12127), .IN2(n12126), .Q(n12123) );
  AND2X1 U12260 ( .IN1(n12128), .IN2(n12129), .Q(n12126) );
  OR2X1 U12261 ( .IN1(n9481), .IN2(n7998), .Q(n12129) );
  OR2X1 U12262 ( .IN1(WX7180), .IN2(n9447), .Q(n12128) );
  OR2X1 U12263 ( .IN1(n12130), .IN2(n12131), .Q(n12127) );
  INVX0 U12264 ( .INP(n12132), .ZN(n12131) );
  OR2X1 U12265 ( .IN1(n12133), .IN2(n7999), .Q(n12132) );
  AND2X1 U12266 ( .IN1(n7999), .IN2(n12133), .Q(n12130) );
  INVX0 U12267 ( .INP(n12134), .ZN(n12133) );
  OR2X1 U12268 ( .IN1(n12135), .IN2(n12136), .Q(n12134) );
  AND2X1 U12269 ( .IN1(n8823), .IN2(n8434), .Q(n12136) );
  AND2X1 U12270 ( .IN1(n15919), .IN2(WX7308), .Q(n12135) );
  AND2X1 U12271 ( .IN1(n9228), .IN2(CRC_OUT_5_28), .Q(n12119) );
  AND2X1 U12272 ( .IN1(n992), .IN2(n9202), .Q(n12118) );
  INVX0 U12273 ( .INP(n12137), .ZN(n992) );
  OR2X1 U12274 ( .IN1(n9567), .IN2(n3938), .Q(n12137) );
  OR4X1 U12275 ( .IN1(n12138), .IN2(n12139), .IN3(n12140), .IN4(n12141), .Q(
        WX5820) );
  AND2X1 U12276 ( .IN1(n9193), .IN2(n12142), .Q(n12141) );
  AND2X1 U12277 ( .IN1(n9279), .IN2(n11297), .Q(n12140) );
  OR2X1 U12278 ( .IN1(n12143), .IN2(n12144), .Q(n11297) );
  INVX0 U12279 ( .INP(n12145), .ZN(n12144) );
  OR2X1 U12280 ( .IN1(n12146), .IN2(n12147), .Q(n12145) );
  AND2X1 U12281 ( .IN1(n12147), .IN2(n12146), .Q(n12143) );
  AND2X1 U12282 ( .IN1(n12148), .IN2(n12149), .Q(n12146) );
  OR2X1 U12283 ( .IN1(n9452), .IN2(n8000), .Q(n12149) );
  OR2X1 U12284 ( .IN1(WX7178), .IN2(n9447), .Q(n12148) );
  OR2X1 U12285 ( .IN1(n12150), .IN2(n12151), .Q(n12147) );
  INVX0 U12286 ( .INP(n12152), .ZN(n12151) );
  OR2X1 U12287 ( .IN1(n12153), .IN2(n8001), .Q(n12152) );
  AND2X1 U12288 ( .IN1(n8001), .IN2(n12153), .Q(n12150) );
  INVX0 U12289 ( .INP(n12154), .ZN(n12153) );
  OR2X1 U12290 ( .IN1(n12155), .IN2(n12156), .Q(n12154) );
  AND2X1 U12291 ( .IN1(n8822), .IN2(n8435), .Q(n12156) );
  AND2X1 U12292 ( .IN1(n15920), .IN2(WX7306), .Q(n12155) );
  AND2X1 U12293 ( .IN1(n9229), .IN2(CRC_OUT_5_29), .Q(n12139) );
  AND2X1 U12294 ( .IN1(n991), .IN2(n9202), .Q(n12138) );
  INVX0 U12295 ( .INP(n12157), .ZN(n991) );
  OR2X1 U12296 ( .IN1(n9567), .IN2(n3939), .Q(n12157) );
  OR4X1 U12297 ( .IN1(n12158), .IN2(n12159), .IN3(n12160), .IN4(n12161), .Q(
        WX5818) );
  AND2X1 U12298 ( .IN1(n9193), .IN2(n12162), .Q(n12161) );
  AND2X1 U12299 ( .IN1(n9279), .IN2(n11317), .Q(n12160) );
  OR2X1 U12300 ( .IN1(n12163), .IN2(n12164), .Q(n11317) );
  AND2X1 U12301 ( .IN1(n12165), .IN2(n12166), .Q(n12164) );
  INVX0 U12302 ( .INP(n12167), .ZN(n12166) );
  AND2X1 U12303 ( .IN1(n12167), .IN2(n12168), .Q(n12163) );
  INVX0 U12304 ( .INP(n12165), .ZN(n12168) );
  OR2X1 U12305 ( .IN1(n12169), .IN2(n12170), .Q(n12165) );
  AND2X1 U12306 ( .IN1(n9450), .IN2(n8436), .Q(n12170) );
  AND2X1 U12307 ( .IN1(n15921), .IN2(n9469), .Q(n12169) );
  OR2X1 U12308 ( .IN1(n12171), .IN2(n12172), .Q(n12167) );
  AND3X1 U12309 ( .IN1(n12173), .IN2(n12174), .IN3(n8821), .Q(n12172) );
  OR2X1 U12310 ( .IN1(n8002), .IN2(WX7240), .Q(n12174) );
  OR2X1 U12311 ( .IN1(n8003), .IN2(WX7176), .Q(n12173) );
  AND2X1 U12312 ( .IN1(n12175), .IN2(WX7304), .Q(n12171) );
  OR2X1 U12313 ( .IN1(n12176), .IN2(n12177), .Q(n12175) );
  AND2X1 U12314 ( .IN1(n8002), .IN2(WX7240), .Q(n12177) );
  AND2X1 U12315 ( .IN1(n8003), .IN2(WX7176), .Q(n12176) );
  AND2X1 U12316 ( .IN1(n9228), .IN2(CRC_OUT_5_30), .Q(n12159) );
  AND2X1 U12317 ( .IN1(n990), .IN2(n9202), .Q(n12158) );
  INVX0 U12318 ( .INP(n12178), .ZN(n990) );
  OR2X1 U12319 ( .IN1(n9567), .IN2(n3940), .Q(n12178) );
  OR4X1 U12320 ( .IN1(n12179), .IN2(n12180), .IN3(n12181), .IN4(n12182), .Q(
        WX5816) );
  AND2X1 U12321 ( .IN1(n9193), .IN2(n12183), .Q(n12182) );
  AND2X1 U12322 ( .IN1(n9279), .IN2(n11336), .Q(n12181) );
  OR2X1 U12323 ( .IN1(n12184), .IN2(n12185), .Q(n11336) );
  INVX0 U12324 ( .INP(n12186), .ZN(n12185) );
  OR2X1 U12325 ( .IN1(n12187), .IN2(n12188), .Q(n12186) );
  AND2X1 U12326 ( .IN1(n12188), .IN2(n12187), .Q(n12184) );
  AND2X1 U12327 ( .IN1(n12189), .IN2(n12190), .Q(n12187) );
  OR2X1 U12328 ( .IN1(n9468), .IN2(n7882), .Q(n12190) );
  OR2X1 U12329 ( .IN1(WX7174), .IN2(n9447), .Q(n12189) );
  OR2X1 U12330 ( .IN1(n12191), .IN2(n12192), .Q(n12188) );
  INVX0 U12331 ( .INP(n12193), .ZN(n12192) );
  OR2X1 U12332 ( .IN1(n12194), .IN2(n7883), .Q(n12193) );
  AND2X1 U12333 ( .IN1(n7883), .IN2(n12194), .Q(n12191) );
  INVX0 U12334 ( .INP(n12195), .ZN(n12194) );
  OR2X1 U12335 ( .IN1(n12196), .IN2(n12197), .Q(n12195) );
  AND2X1 U12336 ( .IN1(n8820), .IN2(n8437), .Q(n12197) );
  AND2X1 U12337 ( .IN1(n15922), .IN2(WX7302), .Q(n12196) );
  AND2X1 U12338 ( .IN1(n2245), .IN2(WX5657), .Q(n12180) );
  AND2X1 U12339 ( .IN1(n9230), .IN2(CRC_OUT_5_31), .Q(n12179) );
  AND2X1 U12340 ( .IN1(n9048), .IN2(n9493), .Q(WX5718) );
  AND2X1 U12341 ( .IN1(n9078), .IN2(n9494), .Q(WX546) );
  AND3X1 U12342 ( .IN1(n12198), .IN2(n12199), .IN3(n9530), .Q(WX5205) );
  OR2X1 U12343 ( .IN1(DFF_766_n1), .IN2(WX4716), .Q(n12199) );
  OR2X1 U12344 ( .IN1(n8875), .IN2(CRC_OUT_6_30), .Q(n12198) );
  AND3X1 U12345 ( .IN1(n12200), .IN2(n12201), .IN3(n9530), .Q(WX5203) );
  OR2X1 U12346 ( .IN1(DFF_765_n1), .IN2(WX4718), .Q(n12201) );
  OR2X1 U12347 ( .IN1(n8876), .IN2(CRC_OUT_6_29), .Q(n12200) );
  AND3X1 U12348 ( .IN1(n12202), .IN2(n12203), .IN3(n9530), .Q(WX5201) );
  OR2X1 U12349 ( .IN1(DFF_764_n1), .IN2(WX4720), .Q(n12203) );
  OR2X1 U12350 ( .IN1(n8877), .IN2(CRC_OUT_6_28), .Q(n12202) );
  AND2X1 U12351 ( .IN1(n12204), .IN2(n9494), .Q(WX5199) );
  OR2X1 U12352 ( .IN1(n12205), .IN2(n12206), .Q(n12204) );
  AND2X1 U12353 ( .IN1(DFF_763_n1), .IN2(n9106), .Q(n12206) );
  AND2X1 U12354 ( .IN1(test_so40), .IN2(CRC_OUT_6_27), .Q(n12205) );
  AND3X1 U12355 ( .IN1(n12207), .IN2(n12208), .IN3(n9530), .Q(WX5197) );
  OR2X1 U12356 ( .IN1(DFF_762_n1), .IN2(WX4724), .Q(n12208) );
  OR2X1 U12357 ( .IN1(n8878), .IN2(CRC_OUT_6_26), .Q(n12207) );
  AND3X1 U12358 ( .IN1(n12209), .IN2(n12210), .IN3(n9530), .Q(WX5195) );
  OR2X1 U12359 ( .IN1(DFF_761_n1), .IN2(WX4726), .Q(n12210) );
  OR2X1 U12360 ( .IN1(n8879), .IN2(CRC_OUT_6_25), .Q(n12209) );
  AND3X1 U12361 ( .IN1(n12211), .IN2(n12212), .IN3(n9530), .Q(WX5193) );
  OR2X1 U12362 ( .IN1(DFF_760_n1), .IN2(WX4728), .Q(n12212) );
  OR2X1 U12363 ( .IN1(n8880), .IN2(CRC_OUT_6_24), .Q(n12211) );
  AND3X1 U12364 ( .IN1(n12213), .IN2(n12214), .IN3(n9530), .Q(WX5191) );
  OR2X1 U12365 ( .IN1(DFF_759_n1), .IN2(WX4730), .Q(n12214) );
  OR2X1 U12366 ( .IN1(n8881), .IN2(CRC_OUT_6_23), .Q(n12213) );
  AND2X1 U12367 ( .IN1(n12215), .IN2(n9493), .Q(WX5189) );
  OR2X1 U12368 ( .IN1(n12216), .IN2(n12217), .Q(n12215) );
  AND2X1 U12369 ( .IN1(n8882), .IN2(n9156), .Q(n12217) );
  AND2X1 U12370 ( .IN1(test_so43), .IN2(WX4732), .Q(n12216) );
  AND3X1 U12371 ( .IN1(n12218), .IN2(n12219), .IN3(n9530), .Q(WX5187) );
  OR2X1 U12372 ( .IN1(DFF_757_n1), .IN2(WX4734), .Q(n12219) );
  OR2X1 U12373 ( .IN1(n8883), .IN2(CRC_OUT_6_21), .Q(n12218) );
  AND3X1 U12374 ( .IN1(n12220), .IN2(n12221), .IN3(n9530), .Q(WX5185) );
  OR2X1 U12375 ( .IN1(DFF_756_n1), .IN2(WX4736), .Q(n12221) );
  OR2X1 U12376 ( .IN1(n8884), .IN2(CRC_OUT_6_20), .Q(n12220) );
  AND3X1 U12377 ( .IN1(n12222), .IN2(n12223), .IN3(n9530), .Q(WX5183) );
  OR2X1 U12378 ( .IN1(DFF_755_n1), .IN2(WX4738), .Q(n12223) );
  OR2X1 U12379 ( .IN1(n8885), .IN2(CRC_OUT_6_19), .Q(n12222) );
  AND3X1 U12380 ( .IN1(n12224), .IN2(n12225), .IN3(n9530), .Q(WX5181) );
  OR2X1 U12381 ( .IN1(DFF_754_n1), .IN2(WX4740), .Q(n12225) );
  OR2X1 U12382 ( .IN1(n8886), .IN2(CRC_OUT_6_18), .Q(n12224) );
  AND3X1 U12383 ( .IN1(n12226), .IN2(n12227), .IN3(n9529), .Q(WX5179) );
  OR2X1 U12384 ( .IN1(DFF_753_n1), .IN2(WX4742), .Q(n12227) );
  OR2X1 U12385 ( .IN1(n8887), .IN2(CRC_OUT_6_17), .Q(n12226) );
  AND3X1 U12386 ( .IN1(n12228), .IN2(n12229), .IN3(n9529), .Q(WX5177) );
  OR2X1 U12387 ( .IN1(DFF_752_n1), .IN2(WX4744), .Q(n12229) );
  OR2X1 U12388 ( .IN1(n8888), .IN2(CRC_OUT_6_16), .Q(n12228) );
  AND2X1 U12389 ( .IN1(n12230), .IN2(n9494), .Q(WX5175) );
  OR2X1 U12390 ( .IN1(n12231), .IN2(n12232), .Q(n12230) );
  AND2X1 U12391 ( .IN1(n12233), .IN2(CRC_OUT_6_15), .Q(n12232) );
  AND2X1 U12392 ( .IN1(DFF_751_n1), .IN2(n12234), .Q(n12231) );
  INVX0 U12393 ( .INP(n12233), .ZN(n12234) );
  OR2X1 U12394 ( .IN1(n12235), .IN2(n12236), .Q(n12233) );
  AND2X1 U12395 ( .IN1(DFF_767_n1), .IN2(WX4746), .Q(n12236) );
  AND2X1 U12396 ( .IN1(n8726), .IN2(CRC_OUT_6_31), .Q(n12235) );
  AND3X1 U12397 ( .IN1(n12237), .IN2(n12238), .IN3(n9529), .Q(WX5173) );
  OR2X1 U12398 ( .IN1(DFF_750_n1), .IN2(WX4748), .Q(n12238) );
  OR2X1 U12399 ( .IN1(n8889), .IN2(CRC_OUT_6_14), .Q(n12237) );
  AND3X1 U12400 ( .IN1(n12239), .IN2(n12240), .IN3(n9529), .Q(WX5171) );
  OR2X1 U12401 ( .IN1(DFF_749_n1), .IN2(WX4750), .Q(n12240) );
  OR2X1 U12402 ( .IN1(n8890), .IN2(CRC_OUT_6_13), .Q(n12239) );
  AND3X1 U12403 ( .IN1(n12241), .IN2(n12242), .IN3(n9529), .Q(WX5169) );
  OR2X1 U12404 ( .IN1(DFF_748_n1), .IN2(WX4752), .Q(n12242) );
  OR2X1 U12405 ( .IN1(n8891), .IN2(CRC_OUT_6_12), .Q(n12241) );
  AND3X1 U12406 ( .IN1(n12243), .IN2(n12244), .IN3(n9529), .Q(WX5167) );
  OR2X1 U12407 ( .IN1(DFF_747_n1), .IN2(WX4754), .Q(n12244) );
  OR2X1 U12408 ( .IN1(n8892), .IN2(CRC_OUT_6_11), .Q(n12243) );
  AND3X1 U12409 ( .IN1(n12245), .IN2(n12246), .IN3(n9529), .Q(WX5165) );
  OR2X1 U12410 ( .IN1(DFF_746_n1), .IN2(n12247), .Q(n12246) );
  AND2X1 U12411 ( .IN1(n12248), .IN2(n12249), .Q(n12247) );
  OR2X1 U12412 ( .IN1(DFF_767_n1), .IN2(n9088), .Q(n12249) );
  OR2X1 U12413 ( .IN1(test_so41), .IN2(CRC_OUT_6_31), .Q(n12248) );
  OR3X1 U12414 ( .IN1(n12250), .IN2(n12251), .IN3(CRC_OUT_6_10), .Q(n12245) );
  AND2X1 U12415 ( .IN1(DFF_767_n1), .IN2(n9088), .Q(n12251) );
  AND2X1 U12416 ( .IN1(test_so41), .IN2(CRC_OUT_6_31), .Q(n12250) );
  AND3X1 U12417 ( .IN1(n12252), .IN2(n12253), .IN3(n9529), .Q(WX5163) );
  OR2X1 U12418 ( .IN1(DFF_745_n1), .IN2(WX4758), .Q(n12253) );
  OR2X1 U12419 ( .IN1(n8893), .IN2(CRC_OUT_6_9), .Q(n12252) );
  AND3X1 U12420 ( .IN1(n12254), .IN2(n12255), .IN3(n9529), .Q(WX5161) );
  OR2X1 U12421 ( .IN1(DFF_744_n1), .IN2(WX4760), .Q(n12255) );
  OR2X1 U12422 ( .IN1(n8894), .IN2(CRC_OUT_6_8), .Q(n12254) );
  AND3X1 U12423 ( .IN1(n12256), .IN2(n12257), .IN3(n9529), .Q(WX5159) );
  OR2X1 U12424 ( .IN1(DFF_743_n1), .IN2(WX4762), .Q(n12257) );
  OR2X1 U12425 ( .IN1(n8895), .IN2(CRC_OUT_6_7), .Q(n12256) );
  AND3X1 U12426 ( .IN1(n12258), .IN2(n12259), .IN3(n9529), .Q(WX5157) );
  OR2X1 U12427 ( .IN1(DFF_742_n1), .IN2(WX4764), .Q(n12259) );
  OR2X1 U12428 ( .IN1(n8896), .IN2(CRC_OUT_6_6), .Q(n12258) );
  AND2X1 U12429 ( .IN1(n12260), .IN2(n9494), .Q(WX5155) );
  OR2X1 U12430 ( .IN1(n12261), .IN2(n12262), .Q(n12260) );
  AND2X1 U12431 ( .IN1(n8897), .IN2(n9157), .Q(n12262) );
  AND2X1 U12432 ( .IN1(test_so42), .IN2(WX4766), .Q(n12261) );
  AND3X1 U12433 ( .IN1(n12263), .IN2(n12264), .IN3(n9529), .Q(WX5153) );
  OR2X1 U12434 ( .IN1(DFF_740_n1), .IN2(WX4768), .Q(n12264) );
  OR2X1 U12435 ( .IN1(n8898), .IN2(CRC_OUT_6_4), .Q(n12263) );
  AND2X1 U12436 ( .IN1(n12265), .IN2(n9492), .Q(WX5151) );
  OR2X1 U12437 ( .IN1(n12266), .IN2(n12267), .Q(n12265) );
  AND2X1 U12438 ( .IN1(n12268), .IN2(CRC_OUT_6_3), .Q(n12267) );
  AND2X1 U12439 ( .IN1(DFF_739_n1), .IN2(n12269), .Q(n12266) );
  INVX0 U12440 ( .INP(n12268), .ZN(n12269) );
  OR2X1 U12441 ( .IN1(n12270), .IN2(n12271), .Q(n12268) );
  AND2X1 U12442 ( .IN1(DFF_767_n1), .IN2(WX4770), .Q(n12271) );
  AND2X1 U12443 ( .IN1(n8727), .IN2(CRC_OUT_6_31), .Q(n12270) );
  AND3X1 U12444 ( .IN1(n12272), .IN2(n12273), .IN3(n9528), .Q(WX5149) );
  OR2X1 U12445 ( .IN1(DFF_738_n1), .IN2(WX4772), .Q(n12273) );
  OR2X1 U12446 ( .IN1(n8899), .IN2(CRC_OUT_6_2), .Q(n12272) );
  AND3X1 U12447 ( .IN1(n12274), .IN2(n12275), .IN3(n9528), .Q(WX5147) );
  OR2X1 U12448 ( .IN1(DFF_737_n1), .IN2(WX4774), .Q(n12275) );
  OR2X1 U12449 ( .IN1(n8900), .IN2(CRC_OUT_6_1), .Q(n12274) );
  AND3X1 U12450 ( .IN1(n12276), .IN2(n12277), .IN3(n9528), .Q(WX5145) );
  OR2X1 U12451 ( .IN1(DFF_736_n1), .IN2(WX4776), .Q(n12277) );
  OR2X1 U12452 ( .IN1(n8901), .IN2(CRC_OUT_6_0), .Q(n12276) );
  AND3X1 U12453 ( .IN1(n12278), .IN2(n12279), .IN3(n9528), .Q(WX5143) );
  OR2X1 U12454 ( .IN1(DFF_767_n1), .IN2(WX4778), .Q(n12279) );
  OR2X1 U12455 ( .IN1(n8739), .IN2(CRC_OUT_6_31), .Q(n12278) );
  AND2X1 U12456 ( .IN1(n9504), .IN2(n8537), .Q(WX4617) );
  AND2X1 U12457 ( .IN1(test_so35), .IN2(n9494), .Q(WX4615) );
  AND2X1 U12458 ( .IN1(n9504), .IN2(n8540), .Q(WX4613) );
  AND2X1 U12459 ( .IN1(n9505), .IN2(n8541), .Q(WX4611) );
  AND2X1 U12460 ( .IN1(n9505), .IN2(n8542), .Q(WX4609) );
  AND2X1 U12461 ( .IN1(n9505), .IN2(n8543), .Q(WX4607) );
  AND2X1 U12462 ( .IN1(n9505), .IN2(n8544), .Q(WX4605) );
  AND2X1 U12463 ( .IN1(n9505), .IN2(n8545), .Q(WX4603) );
  AND2X1 U12464 ( .IN1(n9506), .IN2(n8546), .Q(WX4601) );
  AND2X1 U12465 ( .IN1(n9506), .IN2(n8547), .Q(WX4599) );
  AND2X1 U12466 ( .IN1(n9506), .IN2(n8548), .Q(WX4597) );
  AND2X1 U12467 ( .IN1(n9506), .IN2(n8549), .Q(WX4595) );
  AND2X1 U12468 ( .IN1(n9506), .IN2(n8550), .Q(WX4593) );
  AND2X1 U12469 ( .IN1(n9506), .IN2(n8551), .Q(WX4591) );
  AND2X1 U12470 ( .IN1(n9506), .IN2(n8552), .Q(WX4589) );
  AND2X1 U12471 ( .IN1(n9506), .IN2(n8553), .Q(WX4587) );
  OR4X1 U12472 ( .IN1(n12280), .IN2(n12281), .IN3(n12282), .IN4(n12283), .Q(
        WX4585) );
  AND2X1 U12473 ( .IN1(n12284), .IN2(n9176), .Q(n12283) );
  AND2X1 U12474 ( .IN1(n9279), .IN2(n11628), .Q(n12282) );
  OR2X1 U12475 ( .IN1(n12285), .IN2(n12286), .Q(n11628) );
  INVX0 U12476 ( .INP(n12287), .ZN(n12286) );
  OR2X1 U12477 ( .IN1(n12288), .IN2(n12289), .Q(n12287) );
  AND2X1 U12478 ( .IN1(n12289), .IN2(n12288), .Q(n12285) );
  AND2X1 U12479 ( .IN1(n12290), .IN2(n12291), .Q(n12288) );
  OR2X1 U12480 ( .IN1(WX5943), .IN2(n8239), .Q(n12291) );
  INVX0 U12481 ( .INP(n12292), .ZN(n12290) );
  AND2X1 U12482 ( .IN1(n8239), .IN2(WX5943), .Q(n12292) );
  OR2X1 U12483 ( .IN1(n12293), .IN2(n12294), .Q(n12289) );
  AND2X1 U12484 ( .IN1(n8240), .IN2(WX6071), .Q(n12294) );
  AND2X1 U12485 ( .IN1(n8738), .IN2(WX6007), .Q(n12293) );
  AND2X1 U12486 ( .IN1(n9228), .IN2(CRC_OUT_6_0), .Q(n12281) );
  AND2X1 U12487 ( .IN1(n779), .IN2(n9202), .Q(n12280) );
  INVX0 U12488 ( .INP(n12295), .ZN(n779) );
  OR2X1 U12489 ( .IN1(n9567), .IN2(n3941), .Q(n12295) );
  OR4X1 U12490 ( .IN1(n12296), .IN2(n12297), .IN3(n12298), .IN4(n12299), .Q(
        WX4583) );
  AND2X1 U12491 ( .IN1(n9193), .IN2(n12300), .Q(n12299) );
  AND2X1 U12492 ( .IN1(n11644), .IN2(n9257), .Q(n12298) );
  AND2X1 U12493 ( .IN1(n12301), .IN2(n12302), .Q(n11644) );
  INVX0 U12494 ( .INP(n12303), .ZN(n12302) );
  AND2X1 U12495 ( .IN1(n12304), .IN2(n12305), .Q(n12303) );
  OR2X1 U12496 ( .IN1(n12305), .IN2(n12304), .Q(n12301) );
  OR2X1 U12497 ( .IN1(n12306), .IN2(n12307), .Q(n12304) );
  INVX0 U12498 ( .INP(n12308), .ZN(n12307) );
  OR2X1 U12499 ( .IN1(WX5941), .IN2(n8241), .Q(n12308) );
  AND2X1 U12500 ( .IN1(n8241), .IN2(WX5941), .Q(n12306) );
  AND2X1 U12501 ( .IN1(n12309), .IN2(n12310), .Q(n12305) );
  OR2X1 U12502 ( .IN1(WX6069), .IN2(test_so51), .Q(n12310) );
  OR2X1 U12503 ( .IN1(n9125), .IN2(n8874), .Q(n12309) );
  AND2X1 U12504 ( .IN1(n9229), .IN2(CRC_OUT_6_1), .Q(n12297) );
  AND2X1 U12505 ( .IN1(n778), .IN2(n9202), .Q(n12296) );
  INVX0 U12506 ( .INP(n12311), .ZN(n778) );
  OR2X1 U12507 ( .IN1(n9567), .IN2(n3942), .Q(n12311) );
  OR4X1 U12508 ( .IN1(n12312), .IN2(n12313), .IN3(n12314), .IN4(n12315), .Q(
        WX4581) );
  AND2X1 U12509 ( .IN1(n9193), .IN2(n12316), .Q(n12315) );
  AND2X1 U12510 ( .IN1(n9279), .IN2(n11660), .Q(n12314) );
  OR2X1 U12511 ( .IN1(n12317), .IN2(n12318), .Q(n11660) );
  INVX0 U12512 ( .INP(n12319), .ZN(n12318) );
  OR2X1 U12513 ( .IN1(n12320), .IN2(n12321), .Q(n12319) );
  AND2X1 U12514 ( .IN1(n12321), .IN2(n12320), .Q(n12317) );
  AND2X1 U12515 ( .IN1(n12322), .IN2(n12323), .Q(n12320) );
  OR2X1 U12516 ( .IN1(WX5939), .IN2(n8242), .Q(n12323) );
  INVX0 U12517 ( .INP(n12324), .ZN(n12322) );
  AND2X1 U12518 ( .IN1(n8242), .IN2(WX5939), .Q(n12324) );
  OR2X1 U12519 ( .IN1(n12325), .IN2(n12326), .Q(n12321) );
  AND2X1 U12520 ( .IN1(n8243), .IN2(WX6067), .Q(n12326) );
  AND2X1 U12521 ( .IN1(n8873), .IN2(WX6003), .Q(n12325) );
  AND2X1 U12522 ( .IN1(n9228), .IN2(CRC_OUT_6_2), .Q(n12313) );
  AND2X1 U12523 ( .IN1(n777), .IN2(n9202), .Q(n12312) );
  INVX0 U12524 ( .INP(n12327), .ZN(n777) );
  OR2X1 U12525 ( .IN1(n9567), .IN2(n3943), .Q(n12327) );
  OR4X1 U12526 ( .IN1(n12328), .IN2(n12329), .IN3(n12330), .IN4(n12331), .Q(
        WX4579) );
  AND2X1 U12527 ( .IN1(n9193), .IN2(n12332), .Q(n12331) );
  AND2X1 U12528 ( .IN1(n11676), .IN2(n9257), .Q(n12330) );
  AND2X1 U12529 ( .IN1(n12333), .IN2(n12334), .Q(n11676) );
  INVX0 U12530 ( .INP(n12335), .ZN(n12334) );
  AND2X1 U12531 ( .IN1(n12336), .IN2(n12337), .Q(n12335) );
  OR2X1 U12532 ( .IN1(n12337), .IN2(n12336), .Q(n12333) );
  OR2X1 U12533 ( .IN1(n12338), .IN2(n12339), .Q(n12336) );
  INVX0 U12534 ( .INP(n12340), .ZN(n12339) );
  OR2X1 U12535 ( .IN1(WX5873), .IN2(n8245), .Q(n12340) );
  AND2X1 U12536 ( .IN1(n8245), .IN2(WX5873), .Q(n12338) );
  AND2X1 U12537 ( .IN1(n12341), .IN2(n12342), .Q(n12337) );
  OR2X1 U12538 ( .IN1(WX6065), .IN2(test_so49), .Q(n12342) );
  OR2X1 U12539 ( .IN1(n9126), .IN2(n8872), .Q(n12341) );
  AND2X1 U12540 ( .IN1(n9229), .IN2(CRC_OUT_6_3), .Q(n12329) );
  AND2X1 U12541 ( .IN1(n776), .IN2(n9202), .Q(n12328) );
  INVX0 U12542 ( .INP(n12343), .ZN(n776) );
  OR2X1 U12543 ( .IN1(n9567), .IN2(n3944), .Q(n12343) );
  OR4X1 U12544 ( .IN1(n12344), .IN2(n12345), .IN3(n12346), .IN4(n12347), .Q(
        WX4577) );
  AND2X1 U12545 ( .IN1(n9193), .IN2(n12348), .Q(n12347) );
  AND2X1 U12546 ( .IN1(n9264), .IN2(n11692), .Q(n12346) );
  OR2X1 U12547 ( .IN1(n12349), .IN2(n12350), .Q(n11692) );
  INVX0 U12548 ( .INP(n12351), .ZN(n12350) );
  OR2X1 U12549 ( .IN1(n12352), .IN2(n12353), .Q(n12351) );
  AND2X1 U12550 ( .IN1(n12353), .IN2(n12352), .Q(n12349) );
  AND2X1 U12551 ( .IN1(n12354), .IN2(n12355), .Q(n12352) );
  OR2X1 U12552 ( .IN1(WX5935), .IN2(n8255), .Q(n12355) );
  INVX0 U12553 ( .INP(n12356), .ZN(n12354) );
  AND2X1 U12554 ( .IN1(n8255), .IN2(WX5935), .Q(n12356) );
  OR2X1 U12555 ( .IN1(n12357), .IN2(n12358), .Q(n12353) );
  AND2X1 U12556 ( .IN1(n8256), .IN2(WX6063), .Q(n12358) );
  AND2X1 U12557 ( .IN1(n8725), .IN2(WX5999), .Q(n12357) );
  AND2X1 U12558 ( .IN1(n9229), .IN2(CRC_OUT_6_4), .Q(n12345) );
  AND2X1 U12559 ( .IN1(n775), .IN2(n9202), .Q(n12344) );
  INVX0 U12560 ( .INP(n12359), .ZN(n775) );
  OR2X1 U12561 ( .IN1(n9566), .IN2(n3945), .Q(n12359) );
  OR4X1 U12562 ( .IN1(n12360), .IN2(n12361), .IN3(n12362), .IN4(n12363), .Q(
        WX4575) );
  AND2X1 U12563 ( .IN1(n9193), .IN2(n12364), .Q(n12363) );
  AND2X1 U12564 ( .IN1(n11708), .IN2(n9257), .Q(n12362) );
  AND2X1 U12565 ( .IN1(n12365), .IN2(n12366), .Q(n11708) );
  INVX0 U12566 ( .INP(n12367), .ZN(n12366) );
  AND2X1 U12567 ( .IN1(n12368), .IN2(n12369), .Q(n12367) );
  OR2X1 U12568 ( .IN1(n12369), .IN2(n12368), .Q(n12365) );
  OR2X1 U12569 ( .IN1(n12370), .IN2(n12371), .Q(n12368) );
  INVX0 U12570 ( .INP(n12372), .ZN(n12371) );
  OR2X1 U12571 ( .IN1(WX5933), .IN2(n8273), .Q(n12372) );
  AND2X1 U12572 ( .IN1(n8273), .IN2(WX5933), .Q(n12370) );
  AND2X1 U12573 ( .IN1(n12373), .IN2(n12374), .Q(n12369) );
  OR2X1 U12574 ( .IN1(WX6061), .IN2(test_so47), .Q(n12374) );
  OR2X1 U12575 ( .IN1(n9127), .IN2(n8871), .Q(n12373) );
  AND2X1 U12576 ( .IN1(test_so42), .IN2(n9227), .Q(n12361) );
  AND2X1 U12577 ( .IN1(n774), .IN2(n9202), .Q(n12360) );
  INVX0 U12578 ( .INP(n12375), .ZN(n774) );
  OR2X1 U12579 ( .IN1(n9566), .IN2(n3946), .Q(n12375) );
  OR4X1 U12580 ( .IN1(n12376), .IN2(n12377), .IN3(n12378), .IN4(n12379), .Q(
        WX4573) );
  AND2X1 U12581 ( .IN1(n9193), .IN2(n12380), .Q(n12379) );
  AND2X1 U12582 ( .IN1(n9266), .IN2(n11724), .Q(n12378) );
  OR2X1 U12583 ( .IN1(n12381), .IN2(n12382), .Q(n11724) );
  INVX0 U12584 ( .INP(n12383), .ZN(n12382) );
  OR2X1 U12585 ( .IN1(n12384), .IN2(n12385), .Q(n12383) );
  AND2X1 U12586 ( .IN1(n12385), .IN2(n12384), .Q(n12381) );
  AND2X1 U12587 ( .IN1(n12386), .IN2(n12387), .Q(n12384) );
  OR2X1 U12588 ( .IN1(WX5931), .IN2(n8274), .Q(n12387) );
  INVX0 U12589 ( .INP(n12388), .ZN(n12386) );
  AND2X1 U12590 ( .IN1(n8274), .IN2(WX5931), .Q(n12388) );
  OR2X1 U12591 ( .IN1(n12389), .IN2(n12390), .Q(n12385) );
  AND2X1 U12592 ( .IN1(n8291), .IN2(WX6059), .Q(n12390) );
  AND2X1 U12593 ( .IN1(n8870), .IN2(WX5995), .Q(n12389) );
  AND2X1 U12594 ( .IN1(n9229), .IN2(CRC_OUT_6_6), .Q(n12377) );
  AND2X1 U12595 ( .IN1(n773), .IN2(n9202), .Q(n12376) );
  INVX0 U12596 ( .INP(n12391), .ZN(n773) );
  OR2X1 U12597 ( .IN1(n9566), .IN2(n3947), .Q(n12391) );
  OR4X1 U12598 ( .IN1(n12392), .IN2(n12393), .IN3(n12394), .IN4(n12395), .Q(
        WX4571) );
  AND2X1 U12599 ( .IN1(n9192), .IN2(n12396), .Q(n12395) );
  AND2X1 U12600 ( .IN1(n9264), .IN2(n11740), .Q(n12394) );
  OR2X1 U12601 ( .IN1(n12397), .IN2(n12398), .Q(n11740) );
  INVX0 U12602 ( .INP(n12399), .ZN(n12398) );
  OR2X1 U12603 ( .IN1(n12400), .IN2(n12401), .Q(n12399) );
  AND2X1 U12604 ( .IN1(n12401), .IN2(n12400), .Q(n12397) );
  AND2X1 U12605 ( .IN1(n12402), .IN2(n12403), .Q(n12400) );
  OR2X1 U12606 ( .IN1(WX5929), .IN2(n8292), .Q(n12403) );
  INVX0 U12607 ( .INP(n12404), .ZN(n12402) );
  AND2X1 U12608 ( .IN1(n8292), .IN2(WX5929), .Q(n12404) );
  OR2X1 U12609 ( .IN1(n12405), .IN2(n12406), .Q(n12401) );
  AND2X1 U12610 ( .IN1(n8296), .IN2(WX6057), .Q(n12406) );
  AND2X1 U12611 ( .IN1(n8869), .IN2(WX5993), .Q(n12405) );
  AND2X1 U12612 ( .IN1(n9229), .IN2(CRC_OUT_6_7), .Q(n12393) );
  AND2X1 U12613 ( .IN1(n772), .IN2(n9202), .Q(n12392) );
  INVX0 U12614 ( .INP(n12407), .ZN(n772) );
  OR2X1 U12615 ( .IN1(n9566), .IN2(n3948), .Q(n12407) );
  OR4X1 U12616 ( .IN1(n12408), .IN2(n12409), .IN3(n12410), .IN4(n12411), .Q(
        WX4569) );
  AND2X1 U12617 ( .IN1(n9192), .IN2(n12412), .Q(n12411) );
  AND2X1 U12618 ( .IN1(n9264), .IN2(n11756), .Q(n12410) );
  OR2X1 U12619 ( .IN1(n12413), .IN2(n12414), .Q(n11756) );
  INVX0 U12620 ( .INP(n12415), .ZN(n12414) );
  OR2X1 U12621 ( .IN1(n12416), .IN2(n12417), .Q(n12415) );
  AND2X1 U12622 ( .IN1(n12417), .IN2(n12416), .Q(n12413) );
  AND2X1 U12623 ( .IN1(n12418), .IN2(n12419), .Q(n12416) );
  OR2X1 U12624 ( .IN1(WX5927), .IN2(n8297), .Q(n12419) );
  INVX0 U12625 ( .INP(n12420), .ZN(n12418) );
  AND2X1 U12626 ( .IN1(n8297), .IN2(WX5927), .Q(n12420) );
  OR2X1 U12627 ( .IN1(n12421), .IN2(n12422), .Q(n12417) );
  AND2X1 U12628 ( .IN1(n8298), .IN2(WX6055), .Q(n12422) );
  AND2X1 U12629 ( .IN1(n8868), .IN2(WX5991), .Q(n12421) );
  AND2X1 U12630 ( .IN1(n9231), .IN2(CRC_OUT_6_8), .Q(n12409) );
  AND2X1 U12631 ( .IN1(n771), .IN2(n9203), .Q(n12408) );
  INVX0 U12632 ( .INP(n12423), .ZN(n771) );
  OR2X1 U12633 ( .IN1(n9566), .IN2(n3949), .Q(n12423) );
  OR4X1 U12634 ( .IN1(n12424), .IN2(n12425), .IN3(n12426), .IN4(n12427), .Q(
        WX4567) );
  AND2X1 U12635 ( .IN1(n9192), .IN2(n12428), .Q(n12427) );
  AND2X1 U12636 ( .IN1(n9265), .IN2(n11772), .Q(n12426) );
  OR2X1 U12637 ( .IN1(n12429), .IN2(n12430), .Q(n11772) );
  INVX0 U12638 ( .INP(n12431), .ZN(n12430) );
  OR2X1 U12639 ( .IN1(n12432), .IN2(n12433), .Q(n12431) );
  AND2X1 U12640 ( .IN1(n12433), .IN2(n12432), .Q(n12429) );
  AND2X1 U12641 ( .IN1(n12434), .IN2(n12435), .Q(n12432) );
  OR2X1 U12642 ( .IN1(WX5925), .IN2(n8299), .Q(n12435) );
  INVX0 U12643 ( .INP(n12436), .ZN(n12434) );
  AND2X1 U12644 ( .IN1(n8299), .IN2(WX5925), .Q(n12436) );
  OR2X1 U12645 ( .IN1(n12437), .IN2(n12438), .Q(n12433) );
  AND2X1 U12646 ( .IN1(n8300), .IN2(WX6053), .Q(n12438) );
  AND2X1 U12647 ( .IN1(n8867), .IN2(WX5989), .Q(n12437) );
  AND2X1 U12648 ( .IN1(n9229), .IN2(CRC_OUT_6_9), .Q(n12425) );
  AND2X1 U12649 ( .IN1(n770), .IN2(n9203), .Q(n12424) );
  INVX0 U12650 ( .INP(n12439), .ZN(n770) );
  OR2X1 U12651 ( .IN1(n9566), .IN2(n3950), .Q(n12439) );
  OR4X1 U12652 ( .IN1(n12440), .IN2(n12441), .IN3(n12442), .IN4(n12443), .Q(
        WX4565) );
  AND2X1 U12653 ( .IN1(n9192), .IN2(n12444), .Q(n12443) );
  AND2X1 U12654 ( .IN1(n9265), .IN2(n11788), .Q(n12442) );
  OR2X1 U12655 ( .IN1(n12445), .IN2(n12446), .Q(n11788) );
  INVX0 U12656 ( .INP(n12447), .ZN(n12446) );
  OR2X1 U12657 ( .IN1(n12448), .IN2(n12449), .Q(n12447) );
  AND2X1 U12658 ( .IN1(n12449), .IN2(n12448), .Q(n12445) );
  AND2X1 U12659 ( .IN1(n12450), .IN2(n12451), .Q(n12448) );
  OR2X1 U12660 ( .IN1(WX5923), .IN2(n8301), .Q(n12451) );
  INVX0 U12661 ( .INP(n12452), .ZN(n12450) );
  AND2X1 U12662 ( .IN1(n8301), .IN2(WX5923), .Q(n12452) );
  OR2X1 U12663 ( .IN1(n12453), .IN2(n12454), .Q(n12449) );
  AND2X1 U12664 ( .IN1(n8302), .IN2(WX6051), .Q(n12454) );
  AND2X1 U12665 ( .IN1(n8866), .IN2(WX5987), .Q(n12453) );
  AND2X1 U12666 ( .IN1(n9230), .IN2(CRC_OUT_6_10), .Q(n12441) );
  AND2X1 U12667 ( .IN1(n769), .IN2(n9203), .Q(n12440) );
  INVX0 U12668 ( .INP(n12455), .ZN(n769) );
  OR2X1 U12669 ( .IN1(n9566), .IN2(n3951), .Q(n12455) );
  OR4X1 U12670 ( .IN1(n12456), .IN2(n12457), .IN3(n12458), .IN4(n12459), .Q(
        WX4563) );
  AND2X1 U12671 ( .IN1(n12460), .IN2(n9178), .Q(n12459) );
  AND2X1 U12672 ( .IN1(n9264), .IN2(n11804), .Q(n12458) );
  OR2X1 U12673 ( .IN1(n12461), .IN2(n12462), .Q(n11804) );
  INVX0 U12674 ( .INP(n12463), .ZN(n12462) );
  OR2X1 U12675 ( .IN1(n12464), .IN2(n12465), .Q(n12463) );
  AND2X1 U12676 ( .IN1(n12465), .IN2(n12464), .Q(n12461) );
  AND2X1 U12677 ( .IN1(n12466), .IN2(n12467), .Q(n12464) );
  OR2X1 U12678 ( .IN1(WX5921), .IN2(n8303), .Q(n12467) );
  INVX0 U12679 ( .INP(n12468), .ZN(n12466) );
  AND2X1 U12680 ( .IN1(n8303), .IN2(WX5921), .Q(n12468) );
  OR2X1 U12681 ( .IN1(n12469), .IN2(n12470), .Q(n12465) );
  AND2X1 U12682 ( .IN1(n8308), .IN2(WX6049), .Q(n12470) );
  AND2X1 U12683 ( .IN1(n8724), .IN2(WX5985), .Q(n12469) );
  AND2X1 U12684 ( .IN1(n9229), .IN2(CRC_OUT_6_11), .Q(n12457) );
  AND2X1 U12685 ( .IN1(n768), .IN2(n9203), .Q(n12456) );
  INVX0 U12686 ( .INP(n12471), .ZN(n768) );
  OR2X1 U12687 ( .IN1(n9566), .IN2(n3952), .Q(n12471) );
  OR4X1 U12688 ( .IN1(n12472), .IN2(n12473), .IN3(n12474), .IN4(n12475), .Q(
        WX4561) );
  AND2X1 U12689 ( .IN1(n9192), .IN2(n12476), .Q(n12475) );
  AND2X1 U12690 ( .IN1(n9265), .IN2(n11820), .Q(n12474) );
  OR2X1 U12691 ( .IN1(n12477), .IN2(n12478), .Q(n11820) );
  INVX0 U12692 ( .INP(n12479), .ZN(n12478) );
  OR2X1 U12693 ( .IN1(n12480), .IN2(n12481), .Q(n12479) );
  AND2X1 U12694 ( .IN1(n12481), .IN2(n12480), .Q(n12477) );
  AND2X1 U12695 ( .IN1(n12482), .IN2(n12483), .Q(n12480) );
  OR2X1 U12696 ( .IN1(WX5919), .IN2(n8309), .Q(n12483) );
  INVX0 U12697 ( .INP(n12484), .ZN(n12482) );
  AND2X1 U12698 ( .IN1(n8309), .IN2(WX5919), .Q(n12484) );
  OR2X1 U12699 ( .IN1(n12485), .IN2(n12486), .Q(n12481) );
  AND2X1 U12700 ( .IN1(n8326), .IN2(WX6047), .Q(n12486) );
  AND2X1 U12701 ( .IN1(n8865), .IN2(WX5983), .Q(n12485) );
  AND2X1 U12702 ( .IN1(n9230), .IN2(CRC_OUT_6_12), .Q(n12473) );
  AND2X1 U12703 ( .IN1(n767), .IN2(n9203), .Q(n12472) );
  INVX0 U12704 ( .INP(n12487), .ZN(n767) );
  OR2X1 U12705 ( .IN1(n9566), .IN2(n3953), .Q(n12487) );
  OR4X1 U12706 ( .IN1(n12488), .IN2(n12489), .IN3(n12490), .IN4(n12491), .Q(
        WX4559) );
  AND2X1 U12707 ( .IN1(n12492), .IN2(n9178), .Q(n12491) );
  AND2X1 U12708 ( .IN1(n9265), .IN2(n11836), .Q(n12490) );
  OR2X1 U12709 ( .IN1(n12493), .IN2(n12494), .Q(n11836) );
  INVX0 U12710 ( .INP(n12495), .ZN(n12494) );
  OR2X1 U12711 ( .IN1(n12496), .IN2(n12497), .Q(n12495) );
  AND2X1 U12712 ( .IN1(n12497), .IN2(n12496), .Q(n12493) );
  AND2X1 U12713 ( .IN1(n12498), .IN2(n12499), .Q(n12496) );
  OR2X1 U12714 ( .IN1(WX5917), .IN2(n8327), .Q(n12499) );
  INVX0 U12715 ( .INP(n12500), .ZN(n12498) );
  AND2X1 U12716 ( .IN1(n8327), .IN2(WX5917), .Q(n12500) );
  OR2X1 U12717 ( .IN1(n12501), .IN2(n12502), .Q(n12497) );
  AND2X1 U12718 ( .IN1(n8344), .IN2(WX6045), .Q(n12502) );
  AND2X1 U12719 ( .IN1(n8864), .IN2(WX5981), .Q(n12501) );
  AND2X1 U12720 ( .IN1(n9229), .IN2(CRC_OUT_6_13), .Q(n12489) );
  AND2X1 U12721 ( .IN1(n766), .IN2(n9203), .Q(n12488) );
  INVX0 U12722 ( .INP(n12503), .ZN(n766) );
  OR2X1 U12723 ( .IN1(n9566), .IN2(n3954), .Q(n12503) );
  OR4X1 U12724 ( .IN1(n12504), .IN2(n12505), .IN3(n12506), .IN4(n12507), .Q(
        WX4557) );
  AND2X1 U12725 ( .IN1(n9192), .IN2(n12508), .Q(n12507) );
  AND2X1 U12726 ( .IN1(n9264), .IN2(n11852), .Q(n12506) );
  OR2X1 U12727 ( .IN1(n12509), .IN2(n12510), .Q(n11852) );
  INVX0 U12728 ( .INP(n12511), .ZN(n12510) );
  OR2X1 U12729 ( .IN1(n12512), .IN2(n12513), .Q(n12511) );
  AND2X1 U12730 ( .IN1(n12513), .IN2(n12512), .Q(n12509) );
  AND2X1 U12731 ( .IN1(n12514), .IN2(n12515), .Q(n12512) );
  OR2X1 U12732 ( .IN1(WX5915), .IN2(n8345), .Q(n12515) );
  INVX0 U12733 ( .INP(n12516), .ZN(n12514) );
  AND2X1 U12734 ( .IN1(n8345), .IN2(WX5915), .Q(n12516) );
  OR2X1 U12735 ( .IN1(n12517), .IN2(n12518), .Q(n12513) );
  AND2X1 U12736 ( .IN1(n8354), .IN2(WX6043), .Q(n12518) );
  AND2X1 U12737 ( .IN1(n8863), .IN2(WX5979), .Q(n12517) );
  AND2X1 U12738 ( .IN1(n9231), .IN2(CRC_OUT_6_14), .Q(n12505) );
  AND2X1 U12739 ( .IN1(n765), .IN2(n9203), .Q(n12504) );
  INVX0 U12740 ( .INP(n12519), .ZN(n765) );
  OR2X1 U12741 ( .IN1(n9566), .IN2(n3955), .Q(n12519) );
  OR4X1 U12742 ( .IN1(n12520), .IN2(n12521), .IN3(n12522), .IN4(n12523), .Q(
        WX4555) );
  AND2X1 U12743 ( .IN1(n12524), .IN2(n9176), .Q(n12523) );
  AND2X1 U12744 ( .IN1(n9265), .IN2(n11868), .Q(n12522) );
  OR2X1 U12745 ( .IN1(n12525), .IN2(n12526), .Q(n11868) );
  INVX0 U12746 ( .INP(n12527), .ZN(n12526) );
  OR2X1 U12747 ( .IN1(n12528), .IN2(n12529), .Q(n12527) );
  AND2X1 U12748 ( .IN1(n12529), .IN2(n12528), .Q(n12525) );
  AND2X1 U12749 ( .IN1(n12530), .IN2(n12531), .Q(n12528) );
  OR2X1 U12750 ( .IN1(WX5913), .IN2(n8355), .Q(n12531) );
  INVX0 U12751 ( .INP(n12532), .ZN(n12530) );
  AND2X1 U12752 ( .IN1(n8355), .IN2(WX5913), .Q(n12532) );
  OR2X1 U12753 ( .IN1(n12533), .IN2(n12534), .Q(n12529) );
  AND2X1 U12754 ( .IN1(n8356), .IN2(WX6041), .Q(n12534) );
  AND2X1 U12755 ( .IN1(n8862), .IN2(WX5977), .Q(n12533) );
  AND2X1 U12756 ( .IN1(n9229), .IN2(CRC_OUT_6_15), .Q(n12521) );
  AND2X1 U12757 ( .IN1(n764), .IN2(n9203), .Q(n12520) );
  INVX0 U12758 ( .INP(n12535), .ZN(n764) );
  OR2X1 U12759 ( .IN1(n9566), .IN2(n3956), .Q(n12535) );
  OR4X1 U12760 ( .IN1(n12536), .IN2(n12537), .IN3(n12538), .IN4(n12539), .Q(
        WX4553) );
  AND2X1 U12761 ( .IN1(n9192), .IN2(n12540), .Q(n12539) );
  AND2X1 U12762 ( .IN1(n11884), .IN2(n9257), .Q(n12538) );
  AND2X1 U12763 ( .IN1(n12541), .IN2(n12542), .Q(n11884) );
  INVX0 U12764 ( .INP(n12543), .ZN(n12542) );
  AND2X1 U12765 ( .IN1(n12544), .IN2(n12545), .Q(n12543) );
  OR2X1 U12766 ( .IN1(n12545), .IN2(n12544), .Q(n12541) );
  OR2X1 U12767 ( .IN1(n12546), .IN2(n12547), .Q(n12544) );
  AND2X1 U12768 ( .IN1(n9451), .IN2(WX5911), .Q(n12547) );
  AND2X1 U12769 ( .IN1(n8004), .IN2(n9471), .Q(n12546) );
  AND2X1 U12770 ( .IN1(n12548), .IN2(n12549), .Q(n12545) );
  OR2X1 U12771 ( .IN1(n12550), .IN2(n8005), .Q(n12549) );
  INVX0 U12772 ( .INP(n12551), .ZN(n12550) );
  OR2X1 U12773 ( .IN1(WX5975), .IN2(n12551), .Q(n12548) );
  OR2X1 U12774 ( .IN1(n12552), .IN2(n12553), .Q(n12551) );
  AND2X1 U12775 ( .IN1(n15923), .IN2(n9089), .Q(n12553) );
  AND2X1 U12776 ( .IN1(test_so52), .IN2(n8479), .Q(n12552) );
  AND2X1 U12777 ( .IN1(n9230), .IN2(CRC_OUT_6_16), .Q(n12537) );
  AND2X1 U12778 ( .IN1(n763), .IN2(n9203), .Q(n12536) );
  INVX0 U12779 ( .INP(n12554), .ZN(n763) );
  OR2X1 U12780 ( .IN1(n9565), .IN2(n3957), .Q(n12554) );
  OR4X1 U12781 ( .IN1(n12555), .IN2(n12556), .IN3(n12557), .IN4(n12558), .Q(
        WX4551) );
  AND2X1 U12782 ( .IN1(n12559), .IN2(n9176), .Q(n12558) );
  AND2X1 U12783 ( .IN1(n9264), .IN2(n11904), .Q(n12557) );
  OR2X1 U12784 ( .IN1(n12560), .IN2(n12561), .Q(n11904) );
  INVX0 U12785 ( .INP(n12562), .ZN(n12561) );
  OR2X1 U12786 ( .IN1(n12563), .IN2(n12564), .Q(n12562) );
  AND2X1 U12787 ( .IN1(n12564), .IN2(n12563), .Q(n12560) );
  AND2X1 U12788 ( .IN1(n12565), .IN2(n12566), .Q(n12563) );
  OR2X1 U12789 ( .IN1(n9452), .IN2(n8006), .Q(n12566) );
  OR2X1 U12790 ( .IN1(WX5909), .IN2(n9446), .Q(n12565) );
  OR2X1 U12791 ( .IN1(n12567), .IN2(n12568), .Q(n12564) );
  INVX0 U12792 ( .INP(n12569), .ZN(n12568) );
  OR2X1 U12793 ( .IN1(n12570), .IN2(n8007), .Q(n12569) );
  AND2X1 U12794 ( .IN1(n8007), .IN2(n12570), .Q(n12567) );
  INVX0 U12795 ( .INP(n12571), .ZN(n12570) );
  OR2X1 U12796 ( .IN1(n12572), .IN2(n12573), .Q(n12571) );
  AND2X1 U12797 ( .IN1(n8861), .IN2(n8480), .Q(n12573) );
  AND2X1 U12798 ( .IN1(n15924), .IN2(WX6037), .Q(n12572) );
  AND2X1 U12799 ( .IN1(n9230), .IN2(CRC_OUT_6_17), .Q(n12556) );
  AND2X1 U12800 ( .IN1(n762), .IN2(n9203), .Q(n12555) );
  INVX0 U12801 ( .INP(n12574), .ZN(n762) );
  OR2X1 U12802 ( .IN1(n9565), .IN2(n3958), .Q(n12574) );
  OR4X1 U12803 ( .IN1(n12575), .IN2(n12576), .IN3(n12577), .IN4(n12578), .Q(
        WX4549) );
  AND2X1 U12804 ( .IN1(n9192), .IN2(n12579), .Q(n12578) );
  AND2X1 U12805 ( .IN1(n11924), .IN2(n9260), .Q(n12577) );
  AND2X1 U12806 ( .IN1(n12580), .IN2(n12581), .Q(n11924) );
  INVX0 U12807 ( .INP(n12582), .ZN(n12581) );
  AND2X1 U12808 ( .IN1(n12583), .IN2(n12584), .Q(n12582) );
  OR2X1 U12809 ( .IN1(n12584), .IN2(n12583), .Q(n12580) );
  OR2X1 U12810 ( .IN1(n12585), .IN2(n12586), .Q(n12583) );
  AND2X1 U12811 ( .IN1(n9450), .IN2(WX5907), .Q(n12586) );
  AND2X1 U12812 ( .IN1(n8008), .IN2(n9465), .Q(n12585) );
  AND2X1 U12813 ( .IN1(n12587), .IN2(n12588), .Q(n12584) );
  OR2X1 U12814 ( .IN1(n12589), .IN2(n8860), .Q(n12588) );
  OR2X1 U12815 ( .IN1(WX6035), .IN2(n12590), .Q(n12587) );
  INVX0 U12816 ( .INP(n12589), .ZN(n12590) );
  AND2X1 U12817 ( .IN1(n12591), .IN2(n12592), .Q(n12589) );
  OR2X1 U12818 ( .IN1(n8481), .IN2(test_so50), .Q(n12592) );
  OR2X1 U12819 ( .IN1(n9128), .IN2(n15925), .Q(n12591) );
  AND2X1 U12820 ( .IN1(n9230), .IN2(CRC_OUT_6_18), .Q(n12576) );
  AND2X1 U12821 ( .IN1(n761), .IN2(n9203), .Q(n12575) );
  INVX0 U12822 ( .INP(n12593), .ZN(n761) );
  OR2X1 U12823 ( .IN1(n9565), .IN2(n3959), .Q(n12593) );
  OR4X1 U12824 ( .IN1(n12594), .IN2(n12595), .IN3(n12596), .IN4(n12597), .Q(
        WX4547) );
  AND2X1 U12825 ( .IN1(n9192), .IN2(n12598), .Q(n12597) );
  AND2X1 U12826 ( .IN1(n9264), .IN2(n11944), .Q(n12596) );
  OR2X1 U12827 ( .IN1(n12599), .IN2(n12600), .Q(n11944) );
  INVX0 U12828 ( .INP(n12601), .ZN(n12600) );
  OR2X1 U12829 ( .IN1(n12602), .IN2(n12603), .Q(n12601) );
  AND2X1 U12830 ( .IN1(n12603), .IN2(n12602), .Q(n12599) );
  AND2X1 U12831 ( .IN1(n12604), .IN2(n12605), .Q(n12602) );
  OR2X1 U12832 ( .IN1(n9479), .IN2(n8009), .Q(n12605) );
  OR2X1 U12833 ( .IN1(WX5905), .IN2(n9447), .Q(n12604) );
  OR2X1 U12834 ( .IN1(n12606), .IN2(n12607), .Q(n12603) );
  INVX0 U12835 ( .INP(n12608), .ZN(n12607) );
  OR2X1 U12836 ( .IN1(n12609), .IN2(n8010), .Q(n12608) );
  AND2X1 U12837 ( .IN1(n8010), .IN2(n12609), .Q(n12606) );
  INVX0 U12838 ( .INP(n12610), .ZN(n12609) );
  OR2X1 U12839 ( .IN1(n12611), .IN2(n12612), .Q(n12610) );
  AND2X1 U12840 ( .IN1(n8859), .IN2(n8482), .Q(n12612) );
  AND2X1 U12841 ( .IN1(n15926), .IN2(WX6033), .Q(n12611) );
  AND2X1 U12842 ( .IN1(n9230), .IN2(CRC_OUT_6_19), .Q(n12595) );
  AND2X1 U12843 ( .IN1(n760), .IN2(n9203), .Q(n12594) );
  INVX0 U12844 ( .INP(n12613), .ZN(n760) );
  OR2X1 U12845 ( .IN1(n9565), .IN2(n3960), .Q(n12613) );
  OR4X1 U12846 ( .IN1(n12614), .IN2(n12615), .IN3(n12616), .IN4(n12617), .Q(
        WX4545) );
  AND2X1 U12847 ( .IN1(n9192), .IN2(n12618), .Q(n12617) );
  AND2X1 U12848 ( .IN1(n11964), .IN2(n9257), .Q(n12616) );
  AND2X1 U12849 ( .IN1(n12619), .IN2(n12620), .Q(n11964) );
  INVX0 U12850 ( .INP(n12621), .ZN(n12620) );
  AND2X1 U12851 ( .IN1(n12622), .IN2(n12623), .Q(n12621) );
  OR2X1 U12852 ( .IN1(n12623), .IN2(n12622), .Q(n12619) );
  OR2X1 U12853 ( .IN1(n12624), .IN2(n12625), .Q(n12622) );
  AND2X1 U12854 ( .IN1(n9451), .IN2(WX5967), .Q(n12625) );
  AND2X1 U12855 ( .IN1(n8011), .IN2(n9472), .Q(n12624) );
  AND2X1 U12856 ( .IN1(n12626), .IN2(n12627), .Q(n12623) );
  OR2X1 U12857 ( .IN1(n12628), .IN2(n8858), .Q(n12627) );
  OR2X1 U12858 ( .IN1(WX6031), .IN2(n12629), .Q(n12626) );
  INVX0 U12859 ( .INP(n12628), .ZN(n12629) );
  AND2X1 U12860 ( .IN1(n12630), .IN2(n12631), .Q(n12628) );
  OR2X1 U12861 ( .IN1(n8483), .IN2(test_so48), .Q(n12631) );
  OR2X1 U12862 ( .IN1(n9129), .IN2(n15927), .Q(n12630) );
  AND2X1 U12863 ( .IN1(n9230), .IN2(CRC_OUT_6_20), .Q(n12615) );
  AND2X1 U12864 ( .IN1(n759), .IN2(n9204), .Q(n12614) );
  INVX0 U12865 ( .INP(n12632), .ZN(n759) );
  OR2X1 U12866 ( .IN1(n9565), .IN2(n3961), .Q(n12632) );
  OR4X1 U12867 ( .IN1(n12633), .IN2(n12634), .IN3(n12635), .IN4(n12636), .Q(
        WX4543) );
  AND2X1 U12868 ( .IN1(n9192), .IN2(n12637), .Q(n12636) );
  AND2X1 U12869 ( .IN1(n9265), .IN2(n11984), .Q(n12635) );
  OR2X1 U12870 ( .IN1(n12638), .IN2(n12639), .Q(n11984) );
  INVX0 U12871 ( .INP(n12640), .ZN(n12639) );
  OR2X1 U12872 ( .IN1(n12641), .IN2(n12642), .Q(n12640) );
  AND2X1 U12873 ( .IN1(n12642), .IN2(n12641), .Q(n12638) );
  AND2X1 U12874 ( .IN1(n12643), .IN2(n12644), .Q(n12641) );
  OR2X1 U12875 ( .IN1(n9453), .IN2(n8012), .Q(n12644) );
  OR2X1 U12876 ( .IN1(WX5901), .IN2(n9447), .Q(n12643) );
  OR2X1 U12877 ( .IN1(n12645), .IN2(n12646), .Q(n12642) );
  INVX0 U12878 ( .INP(n12647), .ZN(n12646) );
  OR2X1 U12879 ( .IN1(n12648), .IN2(n8013), .Q(n12647) );
  AND2X1 U12880 ( .IN1(n8013), .IN2(n12648), .Q(n12645) );
  INVX0 U12881 ( .INP(n12649), .ZN(n12648) );
  OR2X1 U12882 ( .IN1(n12650), .IN2(n12651), .Q(n12649) );
  AND2X1 U12883 ( .IN1(n8857), .IN2(n8484), .Q(n12651) );
  AND2X1 U12884 ( .IN1(n15928), .IN2(WX6029), .Q(n12650) );
  AND2X1 U12885 ( .IN1(n9230), .IN2(CRC_OUT_6_21), .Q(n12634) );
  AND2X1 U12886 ( .IN1(n758), .IN2(n9204), .Q(n12633) );
  INVX0 U12887 ( .INP(n12652), .ZN(n758) );
  OR2X1 U12888 ( .IN1(n9565), .IN2(n3962), .Q(n12652) );
  OR4X1 U12889 ( .IN1(n12653), .IN2(n12654), .IN3(n12655), .IN4(n12656), .Q(
        WX4541) );
  AND2X1 U12890 ( .IN1(n9192), .IN2(n12657), .Q(n12656) );
  AND2X1 U12891 ( .IN1(n12003), .IN2(n9257), .Q(n12655) );
  AND2X1 U12892 ( .IN1(n12658), .IN2(n12659), .Q(n12003) );
  OR2X1 U12893 ( .IN1(n12660), .IN2(n12661), .Q(n12659) );
  INVX0 U12894 ( .INP(n12662), .ZN(n12658) );
  AND2X1 U12895 ( .IN1(n12661), .IN2(n12660), .Q(n12662) );
  INVX0 U12896 ( .INP(n12663), .ZN(n12660) );
  OR2X1 U12897 ( .IN1(n12664), .IN2(n12665), .Q(n12663) );
  AND2X1 U12898 ( .IN1(n9450), .IN2(WX6027), .Q(n12665) );
  AND2X1 U12899 ( .IN1(n8856), .IN2(n9458), .Q(n12664) );
  OR2X1 U12900 ( .IN1(n12666), .IN2(n12667), .Q(n12661) );
  AND3X1 U12901 ( .IN1(n12668), .IN2(n12669), .IN3(n8015), .Q(n12667) );
  OR2X1 U12902 ( .IN1(n8014), .IN2(n9093), .Q(n12669) );
  OR2X1 U12903 ( .IN1(test_so46), .IN2(WX5899), .Q(n12668) );
  AND2X1 U12904 ( .IN1(n12670), .IN2(WX5963), .Q(n12666) );
  OR2X1 U12905 ( .IN1(n12671), .IN2(n12672), .Q(n12670) );
  AND2X1 U12906 ( .IN1(n8014), .IN2(n9093), .Q(n12672) );
  AND2X1 U12907 ( .IN1(test_so46), .IN2(WX5899), .Q(n12671) );
  AND2X1 U12908 ( .IN1(test_so43), .IN2(n9227), .Q(n12654) );
  AND2X1 U12909 ( .IN1(n757), .IN2(n9204), .Q(n12653) );
  INVX0 U12910 ( .INP(n12673), .ZN(n757) );
  OR2X1 U12911 ( .IN1(n9565), .IN2(n3963), .Q(n12673) );
  OR4X1 U12912 ( .IN1(n12674), .IN2(n12675), .IN3(n12676), .IN4(n12677), .Q(
        WX4539) );
  AND2X1 U12913 ( .IN1(n9192), .IN2(n12678), .Q(n12677) );
  AND2X1 U12914 ( .IN1(n9265), .IN2(n12023), .Q(n12676) );
  OR2X1 U12915 ( .IN1(n12679), .IN2(n12680), .Q(n12023) );
  INVX0 U12916 ( .INP(n12681), .ZN(n12680) );
  OR2X1 U12917 ( .IN1(n12682), .IN2(n12683), .Q(n12681) );
  AND2X1 U12918 ( .IN1(n12683), .IN2(n12682), .Q(n12679) );
  AND2X1 U12919 ( .IN1(n12684), .IN2(n12685), .Q(n12682) );
  OR2X1 U12920 ( .IN1(n9454), .IN2(n8016), .Q(n12685) );
  OR2X1 U12921 ( .IN1(WX5897), .IN2(n9446), .Q(n12684) );
  OR2X1 U12922 ( .IN1(n12686), .IN2(n12687), .Q(n12683) );
  INVX0 U12923 ( .INP(n12688), .ZN(n12687) );
  OR2X1 U12924 ( .IN1(n12689), .IN2(n8017), .Q(n12688) );
  AND2X1 U12925 ( .IN1(n8017), .IN2(n12689), .Q(n12686) );
  INVX0 U12926 ( .INP(n12690), .ZN(n12689) );
  OR2X1 U12927 ( .IN1(n12691), .IN2(n12692), .Q(n12690) );
  AND2X1 U12928 ( .IN1(n8855), .IN2(n8487), .Q(n12692) );
  AND2X1 U12929 ( .IN1(n15929), .IN2(WX6025), .Q(n12691) );
  AND2X1 U12930 ( .IN1(n9231), .IN2(CRC_OUT_6_23), .Q(n12675) );
  AND2X1 U12931 ( .IN1(n756), .IN2(n9204), .Q(n12674) );
  INVX0 U12932 ( .INP(n12693), .ZN(n756) );
  OR2X1 U12933 ( .IN1(n9565), .IN2(n3964), .Q(n12693) );
  OR4X1 U12934 ( .IN1(n12694), .IN2(n12695), .IN3(n12696), .IN4(n12697), .Q(
        WX4537) );
  AND2X1 U12935 ( .IN1(n9191), .IN2(n12698), .Q(n12697) );
  AND2X1 U12936 ( .IN1(n9265), .IN2(n12042), .Q(n12696) );
  OR2X1 U12937 ( .IN1(n12699), .IN2(n12700), .Q(n12042) );
  INVX0 U12938 ( .INP(n12701), .ZN(n12700) );
  OR2X1 U12939 ( .IN1(n12702), .IN2(n12703), .Q(n12701) );
  AND2X1 U12940 ( .IN1(n12703), .IN2(n12702), .Q(n12699) );
  AND2X1 U12941 ( .IN1(n12704), .IN2(n12705), .Q(n12702) );
  OR2X1 U12942 ( .IN1(n9454), .IN2(n8018), .Q(n12705) );
  OR2X1 U12943 ( .IN1(WX5895), .IN2(n9446), .Q(n12704) );
  OR2X1 U12944 ( .IN1(n12706), .IN2(n12707), .Q(n12703) );
  INVX0 U12945 ( .INP(n12708), .ZN(n12707) );
  OR2X1 U12946 ( .IN1(n12709), .IN2(n8019), .Q(n12708) );
  AND2X1 U12947 ( .IN1(n8019), .IN2(n12709), .Q(n12706) );
  INVX0 U12948 ( .INP(n12710), .ZN(n12709) );
  OR2X1 U12949 ( .IN1(n12711), .IN2(n12712), .Q(n12710) );
  AND2X1 U12950 ( .IN1(n8854), .IN2(n8488), .Q(n12712) );
  AND2X1 U12951 ( .IN1(n15930), .IN2(WX6023), .Q(n12711) );
  AND2X1 U12952 ( .IN1(n9230), .IN2(CRC_OUT_6_24), .Q(n12695) );
  AND2X1 U12953 ( .IN1(n755), .IN2(n9204), .Q(n12694) );
  INVX0 U12954 ( .INP(n12713), .ZN(n755) );
  OR2X1 U12955 ( .IN1(n9565), .IN2(n3965), .Q(n12713) );
  OR4X1 U12956 ( .IN1(n12714), .IN2(n12715), .IN3(n12716), .IN4(n12717), .Q(
        WX4535) );
  AND2X1 U12957 ( .IN1(n9191), .IN2(n12718), .Q(n12717) );
  AND2X1 U12958 ( .IN1(n9265), .IN2(n12062), .Q(n12716) );
  OR2X1 U12959 ( .IN1(n12719), .IN2(n12720), .Q(n12062) );
  INVX0 U12960 ( .INP(n12721), .ZN(n12720) );
  OR2X1 U12961 ( .IN1(n12722), .IN2(n12723), .Q(n12721) );
  AND2X1 U12962 ( .IN1(n12723), .IN2(n12722), .Q(n12719) );
  AND2X1 U12963 ( .IN1(n12724), .IN2(n12725), .Q(n12722) );
  OR2X1 U12964 ( .IN1(n9455), .IN2(n8020), .Q(n12725) );
  OR2X1 U12965 ( .IN1(WX5893), .IN2(n9446), .Q(n12724) );
  OR2X1 U12966 ( .IN1(n12726), .IN2(n12727), .Q(n12723) );
  INVX0 U12967 ( .INP(n12728), .ZN(n12727) );
  OR2X1 U12968 ( .IN1(n12729), .IN2(n8021), .Q(n12728) );
  AND2X1 U12969 ( .IN1(n8021), .IN2(n12729), .Q(n12726) );
  INVX0 U12970 ( .INP(n12730), .ZN(n12729) );
  OR2X1 U12971 ( .IN1(n12731), .IN2(n12732), .Q(n12730) );
  AND2X1 U12972 ( .IN1(n8853), .IN2(n8489), .Q(n12732) );
  AND2X1 U12973 ( .IN1(n15931), .IN2(WX6021), .Q(n12731) );
  AND2X1 U12974 ( .IN1(n9231), .IN2(CRC_OUT_6_25), .Q(n12715) );
  AND2X1 U12975 ( .IN1(n754), .IN2(n9204), .Q(n12714) );
  INVX0 U12976 ( .INP(n12733), .ZN(n754) );
  OR2X1 U12977 ( .IN1(n9565), .IN2(n3966), .Q(n12733) );
  OR4X1 U12978 ( .IN1(n12734), .IN2(n12735), .IN3(n12736), .IN4(n12737), .Q(
        WX4533) );
  AND2X1 U12979 ( .IN1(n9191), .IN2(n12738), .Q(n12737) );
  AND2X1 U12980 ( .IN1(n9265), .IN2(n12081), .Q(n12736) );
  OR2X1 U12981 ( .IN1(n12739), .IN2(n12740), .Q(n12081) );
  INVX0 U12982 ( .INP(n12741), .ZN(n12740) );
  OR2X1 U12983 ( .IN1(n12742), .IN2(n12743), .Q(n12741) );
  AND2X1 U12984 ( .IN1(n12743), .IN2(n12742), .Q(n12739) );
  AND2X1 U12985 ( .IN1(n12744), .IN2(n12745), .Q(n12742) );
  OR2X1 U12986 ( .IN1(n9455), .IN2(n8022), .Q(n12745) );
  OR2X1 U12987 ( .IN1(WX5891), .IN2(n9446), .Q(n12744) );
  OR2X1 U12988 ( .IN1(n12746), .IN2(n12747), .Q(n12743) );
  INVX0 U12989 ( .INP(n12748), .ZN(n12747) );
  OR2X1 U12990 ( .IN1(n12749), .IN2(n8023), .Q(n12748) );
  AND2X1 U12991 ( .IN1(n8023), .IN2(n12749), .Q(n12746) );
  INVX0 U12992 ( .INP(n12750), .ZN(n12749) );
  OR2X1 U12993 ( .IN1(n12751), .IN2(n12752), .Q(n12750) );
  AND2X1 U12994 ( .IN1(n8852), .IN2(n8490), .Q(n12752) );
  AND2X1 U12995 ( .IN1(n15932), .IN2(WX6019), .Q(n12751) );
  AND2X1 U12996 ( .IN1(n9230), .IN2(CRC_OUT_6_26), .Q(n12735) );
  AND2X1 U12997 ( .IN1(n753), .IN2(n9204), .Q(n12734) );
  INVX0 U12998 ( .INP(n12753), .ZN(n753) );
  OR2X1 U12999 ( .IN1(n9565), .IN2(n3967), .Q(n12753) );
  OR4X1 U13000 ( .IN1(n12754), .IN2(n12755), .IN3(n12756), .IN4(n12757), .Q(
        WX4531) );
  AND2X1 U13001 ( .IN1(n9191), .IN2(n12758), .Q(n12757) );
  AND2X1 U13002 ( .IN1(n9265), .IN2(n12101), .Q(n12756) );
  OR2X1 U13003 ( .IN1(n12759), .IN2(n12760), .Q(n12101) );
  INVX0 U13004 ( .INP(n12761), .ZN(n12760) );
  OR2X1 U13005 ( .IN1(n12762), .IN2(n12763), .Q(n12761) );
  AND2X1 U13006 ( .IN1(n12763), .IN2(n12762), .Q(n12759) );
  AND2X1 U13007 ( .IN1(n12764), .IN2(n12765), .Q(n12762) );
  OR2X1 U13008 ( .IN1(n9456), .IN2(n8024), .Q(n12765) );
  OR2X1 U13009 ( .IN1(WX5889), .IN2(n9446), .Q(n12764) );
  OR2X1 U13010 ( .IN1(n12766), .IN2(n12767), .Q(n12763) );
  INVX0 U13011 ( .INP(n12768), .ZN(n12767) );
  OR2X1 U13012 ( .IN1(n12769), .IN2(n8025), .Q(n12768) );
  AND2X1 U13013 ( .IN1(n8025), .IN2(n12769), .Q(n12766) );
  INVX0 U13014 ( .INP(n12770), .ZN(n12769) );
  OR2X1 U13015 ( .IN1(n12771), .IN2(n12772), .Q(n12770) );
  AND2X1 U13016 ( .IN1(n8851), .IN2(n8491), .Q(n12772) );
  AND2X1 U13017 ( .IN1(n15933), .IN2(WX6017), .Q(n12771) );
  AND2X1 U13018 ( .IN1(n9231), .IN2(CRC_OUT_6_27), .Q(n12755) );
  AND2X1 U13019 ( .IN1(n752), .IN2(n9204), .Q(n12754) );
  INVX0 U13020 ( .INP(n12773), .ZN(n752) );
  OR2X1 U13021 ( .IN1(n9565), .IN2(n3968), .Q(n12773) );
  OR4X1 U13022 ( .IN1(n12774), .IN2(n12775), .IN3(n12776), .IN4(n12777), .Q(
        WX4529) );
  AND2X1 U13023 ( .IN1(n12778), .IN2(n9173), .Q(n12777) );
  AND2X1 U13024 ( .IN1(n9266), .IN2(n12122), .Q(n12776) );
  OR2X1 U13025 ( .IN1(n12779), .IN2(n12780), .Q(n12122) );
  INVX0 U13026 ( .INP(n12781), .ZN(n12780) );
  OR2X1 U13027 ( .IN1(n12782), .IN2(n12783), .Q(n12781) );
  AND2X1 U13028 ( .IN1(n12783), .IN2(n12782), .Q(n12779) );
  AND2X1 U13029 ( .IN1(n12784), .IN2(n12785), .Q(n12782) );
  OR2X1 U13030 ( .IN1(n9456), .IN2(n8026), .Q(n12785) );
  OR2X1 U13031 ( .IN1(WX5887), .IN2(n9446), .Q(n12784) );
  OR2X1 U13032 ( .IN1(n12786), .IN2(n12787), .Q(n12783) );
  INVX0 U13033 ( .INP(n12788), .ZN(n12787) );
  OR2X1 U13034 ( .IN1(n12789), .IN2(n8027), .Q(n12788) );
  AND2X1 U13035 ( .IN1(n8027), .IN2(n12789), .Q(n12786) );
  INVX0 U13036 ( .INP(n12790), .ZN(n12789) );
  OR2X1 U13037 ( .IN1(n12791), .IN2(n12792), .Q(n12790) );
  AND2X1 U13038 ( .IN1(n8850), .IN2(n8492), .Q(n12792) );
  AND2X1 U13039 ( .IN1(n15934), .IN2(WX6015), .Q(n12791) );
  AND2X1 U13040 ( .IN1(n9230), .IN2(CRC_OUT_6_28), .Q(n12775) );
  AND2X1 U13041 ( .IN1(n751), .IN2(n9204), .Q(n12774) );
  INVX0 U13042 ( .INP(n12793), .ZN(n751) );
  OR2X1 U13043 ( .IN1(n9564), .IN2(n3969), .Q(n12793) );
  OR4X1 U13044 ( .IN1(n12794), .IN2(n12795), .IN3(n12796), .IN4(n12797), .Q(
        WX4527) );
  AND2X1 U13045 ( .IN1(n9191), .IN2(n12798), .Q(n12797) );
  AND2X1 U13046 ( .IN1(n9265), .IN2(n12142), .Q(n12796) );
  OR2X1 U13047 ( .IN1(n12799), .IN2(n12800), .Q(n12142) );
  INVX0 U13048 ( .INP(n12801), .ZN(n12800) );
  OR2X1 U13049 ( .IN1(n12802), .IN2(n12803), .Q(n12801) );
  AND2X1 U13050 ( .IN1(n12803), .IN2(n12802), .Q(n12799) );
  AND2X1 U13051 ( .IN1(n12804), .IN2(n12805), .Q(n12802) );
  OR2X1 U13052 ( .IN1(n9457), .IN2(n8028), .Q(n12805) );
  OR2X1 U13053 ( .IN1(WX5885), .IN2(n9446), .Q(n12804) );
  OR2X1 U13054 ( .IN1(n12806), .IN2(n12807), .Q(n12803) );
  INVX0 U13055 ( .INP(n12808), .ZN(n12807) );
  OR2X1 U13056 ( .IN1(n12809), .IN2(n8029), .Q(n12808) );
  AND2X1 U13057 ( .IN1(n8029), .IN2(n12809), .Q(n12806) );
  INVX0 U13058 ( .INP(n12810), .ZN(n12809) );
  OR2X1 U13059 ( .IN1(n12811), .IN2(n12812), .Q(n12810) );
  AND2X1 U13060 ( .IN1(n8849), .IN2(n8493), .Q(n12812) );
  AND2X1 U13061 ( .IN1(n15935), .IN2(WX6013), .Q(n12811) );
  AND2X1 U13062 ( .IN1(n9232), .IN2(CRC_OUT_6_29), .Q(n12795) );
  AND2X1 U13063 ( .IN1(n750), .IN2(n9204), .Q(n12794) );
  INVX0 U13064 ( .INP(n12813), .ZN(n750) );
  OR2X1 U13065 ( .IN1(n9564), .IN2(n3970), .Q(n12813) );
  OR4X1 U13066 ( .IN1(n12814), .IN2(n12815), .IN3(n12816), .IN4(n12817), .Q(
        WX4525) );
  AND2X1 U13067 ( .IN1(n12818), .IN2(n9173), .Q(n12817) );
  AND2X1 U13068 ( .IN1(n9266), .IN2(n12162), .Q(n12816) );
  OR2X1 U13069 ( .IN1(n12819), .IN2(n12820), .Q(n12162) );
  INVX0 U13070 ( .INP(n12821), .ZN(n12820) );
  OR2X1 U13071 ( .IN1(n12822), .IN2(n12823), .Q(n12821) );
  AND2X1 U13072 ( .IN1(n12823), .IN2(n12822), .Q(n12819) );
  AND2X1 U13073 ( .IN1(n12824), .IN2(n12825), .Q(n12822) );
  OR2X1 U13074 ( .IN1(n9457), .IN2(n8030), .Q(n12825) );
  OR2X1 U13075 ( .IN1(WX5883), .IN2(n9446), .Q(n12824) );
  OR2X1 U13076 ( .IN1(n12826), .IN2(n12827), .Q(n12823) );
  INVX0 U13077 ( .INP(n12828), .ZN(n12827) );
  OR2X1 U13078 ( .IN1(n12829), .IN2(n8031), .Q(n12828) );
  AND2X1 U13079 ( .IN1(n8031), .IN2(n12829), .Q(n12826) );
  INVX0 U13080 ( .INP(n12830), .ZN(n12829) );
  OR2X1 U13081 ( .IN1(n12831), .IN2(n12832), .Q(n12830) );
  AND2X1 U13082 ( .IN1(n8848), .IN2(n8494), .Q(n12832) );
  AND2X1 U13083 ( .IN1(n15936), .IN2(WX6011), .Q(n12831) );
  AND2X1 U13084 ( .IN1(n9231), .IN2(CRC_OUT_6_30), .Q(n12815) );
  AND2X1 U13085 ( .IN1(n749), .IN2(n9204), .Q(n12814) );
  INVX0 U13086 ( .INP(n12833), .ZN(n749) );
  OR2X1 U13087 ( .IN1(n9564), .IN2(n3971), .Q(n12833) );
  OR4X1 U13088 ( .IN1(n12834), .IN2(n12835), .IN3(n12836), .IN4(n12837), .Q(
        WX4523) );
  AND2X1 U13089 ( .IN1(n9191), .IN2(n12838), .Q(n12837) );
  AND2X1 U13090 ( .IN1(n9266), .IN2(n12183), .Q(n12836) );
  OR2X1 U13091 ( .IN1(n12839), .IN2(n12840), .Q(n12183) );
  INVX0 U13092 ( .INP(n12841), .ZN(n12840) );
  OR2X1 U13093 ( .IN1(n12842), .IN2(n12843), .Q(n12841) );
  AND2X1 U13094 ( .IN1(n12843), .IN2(n12842), .Q(n12839) );
  AND2X1 U13095 ( .IN1(n12844), .IN2(n12845), .Q(n12842) );
  OR2X1 U13096 ( .IN1(n9460), .IN2(n7884), .Q(n12845) );
  OR2X1 U13097 ( .IN1(WX5881), .IN2(n9446), .Q(n12844) );
  OR2X1 U13098 ( .IN1(n12846), .IN2(n12847), .Q(n12843) );
  INVX0 U13099 ( .INP(n12848), .ZN(n12847) );
  OR2X1 U13100 ( .IN1(n12849), .IN2(n7885), .Q(n12848) );
  AND2X1 U13101 ( .IN1(n7885), .IN2(n12849), .Q(n12846) );
  INVX0 U13102 ( .INP(n12850), .ZN(n12849) );
  OR2X1 U13103 ( .IN1(n12851), .IN2(n12852), .Q(n12850) );
  AND2X1 U13104 ( .IN1(n8847), .IN2(n8495), .Q(n12852) );
  AND2X1 U13105 ( .IN1(n15937), .IN2(WX6009), .Q(n12851) );
  AND2X1 U13106 ( .IN1(n2245), .IN2(WX4364), .Q(n12835) );
  AND2X1 U13107 ( .IN1(n9231), .IN2(CRC_OUT_6_31), .Q(n12834) );
  AND2X1 U13108 ( .IN1(n9047), .IN2(n9492), .Q(WX4425) );
  AND3X1 U13109 ( .IN1(n12853), .IN2(n12854), .IN3(n9528), .Q(WX3912) );
  OR2X1 U13110 ( .IN1(DFF_574_n1), .IN2(WX3423), .Q(n12854) );
  OR2X1 U13111 ( .IN1(n8902), .IN2(CRC_OUT_7_30), .Q(n12853) );
  AND3X1 U13112 ( .IN1(n12855), .IN2(n12856), .IN3(n9528), .Q(WX3910) );
  OR2X1 U13113 ( .IN1(DFF_573_n1), .IN2(WX3425), .Q(n12856) );
  OR2X1 U13114 ( .IN1(n8903), .IN2(CRC_OUT_7_29), .Q(n12855) );
  AND3X1 U13115 ( .IN1(n12857), .IN2(n12858), .IN3(n9528), .Q(WX3908) );
  OR2X1 U13116 ( .IN1(DFF_572_n1), .IN2(WX3427), .Q(n12858) );
  OR2X1 U13117 ( .IN1(n8904), .IN2(CRC_OUT_7_28), .Q(n12857) );
  AND2X1 U13118 ( .IN1(n12859), .IN2(n9494), .Q(WX3906) );
  OR2X1 U13119 ( .IN1(n12860), .IN2(n12861), .Q(n12859) );
  AND2X1 U13120 ( .IN1(n8905), .IN2(n9158), .Q(n12861) );
  AND2X1 U13121 ( .IN1(test_so32), .IN2(WX3429), .Q(n12860) );
  AND3X1 U13122 ( .IN1(n12862), .IN2(n12863), .IN3(n9528), .Q(WX3904) );
  OR2X1 U13123 ( .IN1(DFF_570_n1), .IN2(WX3431), .Q(n12863) );
  OR2X1 U13124 ( .IN1(n8906), .IN2(CRC_OUT_7_26), .Q(n12862) );
  AND3X1 U13125 ( .IN1(n12864), .IN2(n12865), .IN3(n9528), .Q(WX3902) );
  OR2X1 U13126 ( .IN1(DFF_569_n1), .IN2(WX3433), .Q(n12865) );
  OR2X1 U13127 ( .IN1(n8907), .IN2(CRC_OUT_7_25), .Q(n12864) );
  AND3X1 U13128 ( .IN1(n12866), .IN2(n12867), .IN3(n9528), .Q(WX3900) );
  OR2X1 U13129 ( .IN1(DFF_568_n1), .IN2(WX3435), .Q(n12867) );
  OR2X1 U13130 ( .IN1(n8908), .IN2(CRC_OUT_7_24), .Q(n12866) );
  AND3X1 U13131 ( .IN1(n12868), .IN2(n12869), .IN3(n9528), .Q(WX3898) );
  OR2X1 U13132 ( .IN1(DFF_567_n1), .IN2(WX3437), .Q(n12869) );
  OR2X1 U13133 ( .IN1(n8909), .IN2(CRC_OUT_7_23), .Q(n12868) );
  AND2X1 U13134 ( .IN1(n12870), .IN2(n9492), .Q(WX3896) );
  OR2X1 U13135 ( .IN1(n12871), .IN2(n12872), .Q(n12870) );
  AND2X1 U13136 ( .IN1(DFF_566_n1), .IN2(n9107), .Q(n12872) );
  AND2X1 U13137 ( .IN1(test_so29), .IN2(CRC_OUT_7_22), .Q(n12871) );
  AND3X1 U13138 ( .IN1(n12873), .IN2(n12874), .IN3(n9528), .Q(WX3894) );
  OR2X1 U13139 ( .IN1(DFF_565_n1), .IN2(WX3441), .Q(n12874) );
  OR2X1 U13140 ( .IN1(n8910), .IN2(CRC_OUT_7_21), .Q(n12873) );
  AND3X1 U13141 ( .IN1(n12875), .IN2(n12876), .IN3(n9527), .Q(WX3892) );
  OR2X1 U13142 ( .IN1(DFF_564_n1), .IN2(WX3443), .Q(n12876) );
  OR2X1 U13143 ( .IN1(n8911), .IN2(CRC_OUT_7_20), .Q(n12875) );
  AND3X1 U13144 ( .IN1(n12877), .IN2(n12878), .IN3(n9527), .Q(WX3890) );
  OR2X1 U13145 ( .IN1(DFF_563_n1), .IN2(WX3445), .Q(n12878) );
  OR2X1 U13146 ( .IN1(n8912), .IN2(CRC_OUT_7_19), .Q(n12877) );
  AND3X1 U13147 ( .IN1(n12879), .IN2(n12880), .IN3(n9527), .Q(WX3888) );
  OR2X1 U13148 ( .IN1(DFF_562_n1), .IN2(WX3447), .Q(n12880) );
  OR2X1 U13149 ( .IN1(n8913), .IN2(CRC_OUT_7_18), .Q(n12879) );
  AND3X1 U13150 ( .IN1(n12881), .IN2(n12882), .IN3(n9527), .Q(WX3886) );
  OR2X1 U13151 ( .IN1(DFF_561_n1), .IN2(WX3449), .Q(n12882) );
  OR2X1 U13152 ( .IN1(n8914), .IN2(CRC_OUT_7_17), .Q(n12881) );
  AND3X1 U13153 ( .IN1(n12883), .IN2(n12884), .IN3(n9527), .Q(WX3884) );
  OR2X1 U13154 ( .IN1(DFF_560_n1), .IN2(WX3451), .Q(n12884) );
  OR2X1 U13155 ( .IN1(n8915), .IN2(CRC_OUT_7_16), .Q(n12883) );
  AND2X1 U13156 ( .IN1(n12885), .IN2(n9492), .Q(WX3882) );
  OR2X1 U13157 ( .IN1(n12886), .IN2(n12887), .Q(n12885) );
  AND2X1 U13158 ( .IN1(n12888), .IN2(CRC_OUT_7_15), .Q(n12887) );
  AND2X1 U13159 ( .IN1(DFF_559_n1), .IN2(n12889), .Q(n12886) );
  INVX0 U13160 ( .INP(n12888), .ZN(n12889) );
  OR2X1 U13161 ( .IN1(n12890), .IN2(n12891), .Q(n12888) );
  AND2X1 U13162 ( .IN1(DFF_575_n1), .IN2(WX3453), .Q(n12891) );
  AND2X1 U13163 ( .IN1(n8728), .IN2(CRC_OUT_7_31), .Q(n12890) );
  AND3X1 U13164 ( .IN1(n12892), .IN2(n12893), .IN3(n9527), .Q(WX3880) );
  OR2X1 U13165 ( .IN1(DFF_558_n1), .IN2(WX3455), .Q(n12893) );
  OR2X1 U13166 ( .IN1(n8916), .IN2(CRC_OUT_7_14), .Q(n12892) );
  AND3X1 U13167 ( .IN1(n12894), .IN2(n12895), .IN3(n9527), .Q(WX3878) );
  OR2X1 U13168 ( .IN1(DFF_557_n1), .IN2(WX3457), .Q(n12895) );
  OR2X1 U13169 ( .IN1(n8917), .IN2(CRC_OUT_7_13), .Q(n12894) );
  AND3X1 U13170 ( .IN1(n12896), .IN2(n12897), .IN3(n9527), .Q(WX3876) );
  OR2X1 U13171 ( .IN1(DFF_556_n1), .IN2(WX3459), .Q(n12897) );
  OR2X1 U13172 ( .IN1(n8918), .IN2(CRC_OUT_7_12), .Q(n12896) );
  AND3X1 U13173 ( .IN1(n12898), .IN2(n12899), .IN3(n9527), .Q(WX3874) );
  OR2X1 U13174 ( .IN1(DFF_555_n1), .IN2(WX3461), .Q(n12899) );
  OR2X1 U13175 ( .IN1(n8919), .IN2(CRC_OUT_7_11), .Q(n12898) );
  AND3X1 U13176 ( .IN1(n12900), .IN2(n12901), .IN3(n9527), .Q(WX3872) );
  OR2X1 U13177 ( .IN1(DFF_575_n1), .IN2(n12902), .Q(n12901) );
  AND2X1 U13178 ( .IN1(n12903), .IN2(n12904), .Q(n12902) );
  OR2X1 U13179 ( .IN1(n8729), .IN2(n9090), .Q(n12904) );
  OR2X1 U13180 ( .IN1(test_so31), .IN2(WX3463), .Q(n12903) );
  OR3X1 U13181 ( .IN1(n12905), .IN2(n12906), .IN3(CRC_OUT_7_31), .Q(n12900) );
  AND2X1 U13182 ( .IN1(n8729), .IN2(n9090), .Q(n12906) );
  AND2X1 U13183 ( .IN1(test_so31), .IN2(WX3463), .Q(n12905) );
  AND3X1 U13184 ( .IN1(n12907), .IN2(n12908), .IN3(n9527), .Q(WX3870) );
  OR2X1 U13185 ( .IN1(DFF_553_n1), .IN2(WX3465), .Q(n12908) );
  OR2X1 U13186 ( .IN1(n8920), .IN2(CRC_OUT_7_9), .Q(n12907) );
  AND3X1 U13187 ( .IN1(n12909), .IN2(n12910), .IN3(n9527), .Q(WX3868) );
  OR2X1 U13188 ( .IN1(DFF_552_n1), .IN2(WX3467), .Q(n12910) );
  OR2X1 U13189 ( .IN1(n8921), .IN2(CRC_OUT_7_8), .Q(n12909) );
  AND3X1 U13190 ( .IN1(n12911), .IN2(n12912), .IN3(n9526), .Q(WX3866) );
  OR2X1 U13191 ( .IN1(DFF_551_n1), .IN2(WX3469), .Q(n12912) );
  OR2X1 U13192 ( .IN1(n8922), .IN2(CRC_OUT_7_7), .Q(n12911) );
  AND3X1 U13193 ( .IN1(n12913), .IN2(n12914), .IN3(n9526), .Q(WX3864) );
  OR2X1 U13194 ( .IN1(DFF_550_n1), .IN2(WX3471), .Q(n12914) );
  OR2X1 U13195 ( .IN1(n8923), .IN2(CRC_OUT_7_6), .Q(n12913) );
  AND2X1 U13196 ( .IN1(n12915), .IN2(n9493), .Q(WX3862) );
  OR2X1 U13197 ( .IN1(n12916), .IN2(n12917), .Q(n12915) );
  AND2X1 U13198 ( .IN1(DFF_549_n1), .IN2(n9100), .Q(n12917) );
  AND2X1 U13199 ( .IN1(test_so30), .IN2(CRC_OUT_7_5), .Q(n12916) );
  AND3X1 U13200 ( .IN1(n12918), .IN2(n12919), .IN3(n9526), .Q(WX3860) );
  OR2X1 U13201 ( .IN1(DFF_548_n1), .IN2(WX3475), .Q(n12919) );
  OR2X1 U13202 ( .IN1(n8924), .IN2(CRC_OUT_7_4), .Q(n12918) );
  AND2X1 U13203 ( .IN1(n12920), .IN2(n9495), .Q(WX3858) );
  OR2X1 U13204 ( .IN1(n12921), .IN2(n12922), .Q(n12920) );
  AND2X1 U13205 ( .IN1(n12923), .IN2(CRC_OUT_7_3), .Q(n12922) );
  AND2X1 U13206 ( .IN1(DFF_547_n1), .IN2(n12924), .Q(n12921) );
  INVX0 U13207 ( .INP(n12923), .ZN(n12924) );
  OR2X1 U13208 ( .IN1(n12925), .IN2(n12926), .Q(n12923) );
  AND2X1 U13209 ( .IN1(DFF_575_n1), .IN2(WX3477), .Q(n12926) );
  AND2X1 U13210 ( .IN1(n8730), .IN2(CRC_OUT_7_31), .Q(n12925) );
  AND3X1 U13211 ( .IN1(n12927), .IN2(n12928), .IN3(n9526), .Q(WX3856) );
  OR2X1 U13212 ( .IN1(DFF_546_n1), .IN2(WX3479), .Q(n12928) );
  OR2X1 U13213 ( .IN1(n8925), .IN2(CRC_OUT_7_2), .Q(n12927) );
  AND3X1 U13214 ( .IN1(n12929), .IN2(n12930), .IN3(n9526), .Q(WX3854) );
  OR2X1 U13215 ( .IN1(DFF_545_n1), .IN2(WX3481), .Q(n12930) );
  OR2X1 U13216 ( .IN1(n8926), .IN2(CRC_OUT_7_1), .Q(n12929) );
  AND3X1 U13217 ( .IN1(n12931), .IN2(n12932), .IN3(n9526), .Q(WX3852) );
  OR2X1 U13218 ( .IN1(DFF_544_n1), .IN2(WX3483), .Q(n12932) );
  OR2X1 U13219 ( .IN1(n8927), .IN2(CRC_OUT_7_0), .Q(n12931) );
  AND3X1 U13220 ( .IN1(n12933), .IN2(n12934), .IN3(n9526), .Q(WX3850) );
  OR2X1 U13221 ( .IN1(DFF_575_n1), .IN2(WX3485), .Q(n12934) );
  OR2X1 U13222 ( .IN1(n8740), .IN2(CRC_OUT_7_31), .Q(n12933) );
  AND2X1 U13223 ( .IN1(test_so24), .IN2(n9495), .Q(WX3324) );
  AND2X1 U13224 ( .IN1(n9512), .IN2(n8597), .Q(WX3322) );
  AND2X1 U13225 ( .IN1(n9512), .IN2(n8598), .Q(WX3320) );
  AND2X1 U13226 ( .IN1(n9512), .IN2(n8599), .Q(WX3318) );
  AND2X1 U13227 ( .IN1(n9511), .IN2(n8600), .Q(WX3316) );
  AND2X1 U13228 ( .IN1(n9512), .IN2(n8601), .Q(WX3314) );
  AND2X1 U13229 ( .IN1(n9511), .IN2(n8602), .Q(WX3312) );
  AND2X1 U13230 ( .IN1(n9511), .IN2(n8603), .Q(WX3310) );
  AND2X1 U13231 ( .IN1(n9511), .IN2(n8604), .Q(WX3308) );
  AND2X1 U13232 ( .IN1(n9512), .IN2(n8605), .Q(WX3306) );
  AND2X1 U13233 ( .IN1(n9507), .IN2(n8606), .Q(WX3304) );
  AND2X1 U13234 ( .IN1(n9511), .IN2(n8607), .Q(WX3302) );
  AND2X1 U13235 ( .IN1(n9511), .IN2(n8608), .Q(WX3300) );
  AND2X1 U13236 ( .IN1(n9510), .IN2(n8609), .Q(WX3298) );
  AND2X1 U13237 ( .IN1(n9510), .IN2(n8610), .Q(WX3296) );
  AND2X1 U13238 ( .IN1(n9510), .IN2(n8611), .Q(WX3294) );
  OR4X1 U13239 ( .IN1(n12935), .IN2(n12936), .IN3(n12937), .IN4(n12938), .Q(
        WX3292) );
  AND2X1 U13240 ( .IN1(n9191), .IN2(n12939), .Q(n12938) );
  AND2X1 U13241 ( .IN1(n12284), .IN2(n9258), .Q(n12937) );
  AND2X1 U13242 ( .IN1(n12940), .IN2(n12941), .Q(n12284) );
  INVX0 U13243 ( .INP(n12942), .ZN(n12941) );
  AND2X1 U13244 ( .IN1(n12943), .IN2(n12944), .Q(n12942) );
  OR2X1 U13245 ( .IN1(n12944), .IN2(n12943), .Q(n12940) );
  OR2X1 U13246 ( .IN1(n12945), .IN2(n12946), .Q(n12943) );
  INVX0 U13247 ( .INP(n12947), .ZN(n12946) );
  OR2X1 U13248 ( .IN1(WX4650), .IN2(n8357), .Q(n12947) );
  AND2X1 U13249 ( .IN1(n8357), .IN2(WX4650), .Q(n12945) );
  AND2X1 U13250 ( .IN1(n12948), .IN2(n12949), .Q(n12944) );
  OR2X1 U13251 ( .IN1(WX4778), .IN2(test_so36), .Q(n12949) );
  OR2X1 U13252 ( .IN1(n9130), .IN2(n8739), .Q(n12948) );
  AND2X1 U13253 ( .IN1(n9231), .IN2(CRC_OUT_7_0), .Q(n12936) );
  AND2X1 U13254 ( .IN1(n538), .IN2(n9204), .Q(n12935) );
  INVX0 U13255 ( .INP(n12950), .ZN(n538) );
  OR2X1 U13256 ( .IN1(n9564), .IN2(n3972), .Q(n12950) );
  OR4X1 U13257 ( .IN1(n12951), .IN2(n12952), .IN3(n12953), .IN4(n12954), .Q(
        WX3290) );
  AND2X1 U13258 ( .IN1(n9191), .IN2(n12955), .Q(n12954) );
  AND2X1 U13259 ( .IN1(n9266), .IN2(n12300), .Q(n12953) );
  OR2X1 U13260 ( .IN1(n12956), .IN2(n12957), .Q(n12300) );
  INVX0 U13261 ( .INP(n12958), .ZN(n12957) );
  OR2X1 U13262 ( .IN1(n12959), .IN2(n12960), .Q(n12958) );
  AND2X1 U13263 ( .IN1(n12960), .IN2(n12959), .Q(n12956) );
  AND2X1 U13264 ( .IN1(n12961), .IN2(n12962), .Q(n12959) );
  OR2X1 U13265 ( .IN1(WX4648), .IN2(n8358), .Q(n12962) );
  INVX0 U13266 ( .INP(n12963), .ZN(n12961) );
  AND2X1 U13267 ( .IN1(n8358), .IN2(WX4648), .Q(n12963) );
  OR2X1 U13268 ( .IN1(n12964), .IN2(n12965), .Q(n12960) );
  AND2X1 U13269 ( .IN1(n8359), .IN2(WX4776), .Q(n12965) );
  AND2X1 U13270 ( .IN1(n8901), .IN2(WX4712), .Q(n12964) );
  AND2X1 U13271 ( .IN1(n9231), .IN2(CRC_OUT_7_1), .Q(n12952) );
  AND2X1 U13272 ( .IN1(n537), .IN2(n9205), .Q(n12951) );
  INVX0 U13273 ( .INP(n12966), .ZN(n537) );
  OR2X1 U13274 ( .IN1(n9564), .IN2(n3973), .Q(n12966) );
  OR4X1 U13275 ( .IN1(n12967), .IN2(n12968), .IN3(n12969), .IN4(n12970), .Q(
        WX3288) );
  AND2X1 U13276 ( .IN1(n9191), .IN2(n12971), .Q(n12970) );
  AND2X1 U13277 ( .IN1(n9266), .IN2(n12316), .Q(n12969) );
  OR2X1 U13278 ( .IN1(n12972), .IN2(n12973), .Q(n12316) );
  INVX0 U13279 ( .INP(n12974), .ZN(n12973) );
  OR2X1 U13280 ( .IN1(n12975), .IN2(n12976), .Q(n12974) );
  AND2X1 U13281 ( .IN1(n12976), .IN2(n12975), .Q(n12972) );
  AND2X1 U13282 ( .IN1(n12977), .IN2(n12978), .Q(n12975) );
  OR2X1 U13283 ( .IN1(WX4646), .IN2(n8360), .Q(n12978) );
  INVX0 U13284 ( .INP(n12979), .ZN(n12977) );
  AND2X1 U13285 ( .IN1(n8360), .IN2(WX4646), .Q(n12979) );
  OR2X1 U13286 ( .IN1(n12980), .IN2(n12981), .Q(n12976) );
  AND2X1 U13287 ( .IN1(n8361), .IN2(WX4774), .Q(n12981) );
  AND2X1 U13288 ( .IN1(n8900), .IN2(WX4710), .Q(n12980) );
  AND2X1 U13289 ( .IN1(n9231), .IN2(CRC_OUT_7_2), .Q(n12968) );
  AND2X1 U13290 ( .IN1(n536), .IN2(n9205), .Q(n12967) );
  INVX0 U13291 ( .INP(n12982), .ZN(n536) );
  OR2X1 U13292 ( .IN1(n9564), .IN2(n3974), .Q(n12982) );
  OR4X1 U13293 ( .IN1(n12983), .IN2(n12984), .IN3(n12985), .IN4(n12986), .Q(
        WX3286) );
  AND2X1 U13294 ( .IN1(n9191), .IN2(n12987), .Q(n12986) );
  AND2X1 U13295 ( .IN1(n9266), .IN2(n12332), .Q(n12985) );
  OR2X1 U13296 ( .IN1(n12988), .IN2(n12989), .Q(n12332) );
  INVX0 U13297 ( .INP(n12990), .ZN(n12989) );
  OR2X1 U13298 ( .IN1(n12991), .IN2(n12992), .Q(n12990) );
  AND2X1 U13299 ( .IN1(n12992), .IN2(n12991), .Q(n12988) );
  AND2X1 U13300 ( .IN1(n12993), .IN2(n12994), .Q(n12991) );
  OR2X1 U13301 ( .IN1(WX4644), .IN2(n8362), .Q(n12994) );
  INVX0 U13302 ( .INP(n12995), .ZN(n12993) );
  AND2X1 U13303 ( .IN1(n8362), .IN2(WX4644), .Q(n12995) );
  OR2X1 U13304 ( .IN1(n12996), .IN2(n12997), .Q(n12992) );
  AND2X1 U13305 ( .IN1(n8379), .IN2(WX4772), .Q(n12997) );
  AND2X1 U13306 ( .IN1(n8899), .IN2(WX4708), .Q(n12996) );
  AND2X1 U13307 ( .IN1(n9232), .IN2(CRC_OUT_7_3), .Q(n12984) );
  AND2X1 U13308 ( .IN1(n535), .IN2(n9205), .Q(n12983) );
  INVX0 U13309 ( .INP(n12998), .ZN(n535) );
  OR2X1 U13310 ( .IN1(n9564), .IN2(n3975), .Q(n12998) );
  OR4X1 U13311 ( .IN1(n12999), .IN2(n13000), .IN3(n13001), .IN4(n13002), .Q(
        WX3284) );
  AND2X1 U13312 ( .IN1(n9191), .IN2(n13003), .Q(n13002) );
  AND2X1 U13313 ( .IN1(n9266), .IN2(n12348), .Q(n13001) );
  OR2X1 U13314 ( .IN1(n13004), .IN2(n13005), .Q(n12348) );
  INVX0 U13315 ( .INP(n13006), .ZN(n13005) );
  OR2X1 U13316 ( .IN1(n13007), .IN2(n13008), .Q(n13006) );
  AND2X1 U13317 ( .IN1(n13008), .IN2(n13007), .Q(n13004) );
  AND2X1 U13318 ( .IN1(n13009), .IN2(n13010), .Q(n13007) );
  OR2X1 U13319 ( .IN1(WX4642), .IN2(n8380), .Q(n13010) );
  INVX0 U13320 ( .INP(n13011), .ZN(n13009) );
  AND2X1 U13321 ( .IN1(n8380), .IN2(WX4642), .Q(n13011) );
  OR2X1 U13322 ( .IN1(n13012), .IN2(n13013), .Q(n13008) );
  AND2X1 U13323 ( .IN1(n8397), .IN2(WX4770), .Q(n13013) );
  AND2X1 U13324 ( .IN1(n8727), .IN2(WX4706), .Q(n13012) );
  AND2X1 U13325 ( .IN1(n9231), .IN2(CRC_OUT_7_4), .Q(n13000) );
  AND2X1 U13326 ( .IN1(n534), .IN2(n9205), .Q(n12999) );
  INVX0 U13327 ( .INP(n13014), .ZN(n534) );
  OR2X1 U13328 ( .IN1(n9564), .IN2(n3976), .Q(n13014) );
  OR4X1 U13329 ( .IN1(n13015), .IN2(n13016), .IN3(n13017), .IN4(n13018), .Q(
        WX3282) );
  AND2X1 U13330 ( .IN1(n9191), .IN2(n13019), .Q(n13018) );
  AND2X1 U13331 ( .IN1(n9266), .IN2(n12364), .Q(n13017) );
  OR2X1 U13332 ( .IN1(n13020), .IN2(n13021), .Q(n12364) );
  INVX0 U13333 ( .INP(n13022), .ZN(n13021) );
  OR2X1 U13334 ( .IN1(n13023), .IN2(n13024), .Q(n13022) );
  AND2X1 U13335 ( .IN1(n13024), .IN2(n13023), .Q(n13020) );
  AND2X1 U13336 ( .IN1(n13025), .IN2(n13026), .Q(n13023) );
  OR2X1 U13337 ( .IN1(WX4640), .IN2(n8398), .Q(n13026) );
  INVX0 U13338 ( .INP(n13027), .ZN(n13025) );
  AND2X1 U13339 ( .IN1(n8398), .IN2(WX4640), .Q(n13027) );
  OR2X1 U13340 ( .IN1(n13028), .IN2(n13029), .Q(n13024) );
  AND2X1 U13341 ( .IN1(n8412), .IN2(WX4768), .Q(n13029) );
  AND2X1 U13342 ( .IN1(n8898), .IN2(WX4704), .Q(n13028) );
  AND2X1 U13343 ( .IN1(n9232), .IN2(CRC_OUT_7_5), .Q(n13016) );
  AND2X1 U13344 ( .IN1(n533), .IN2(n9205), .Q(n13015) );
  INVX0 U13345 ( .INP(n13030), .ZN(n533) );
  OR2X1 U13346 ( .IN1(n9564), .IN2(n3977), .Q(n13030) );
  OR4X1 U13347 ( .IN1(n13031), .IN2(n13032), .IN3(n13033), .IN4(n13034), .Q(
        WX3280) );
  AND2X1 U13348 ( .IN1(n13035), .IN2(n9175), .Q(n13034) );
  AND2X1 U13349 ( .IN1(n9266), .IN2(n12380), .Q(n13033) );
  OR2X1 U13350 ( .IN1(n13036), .IN2(n13037), .Q(n12380) );
  INVX0 U13351 ( .INP(n13038), .ZN(n13037) );
  OR2X1 U13352 ( .IN1(n13039), .IN2(n13040), .Q(n13038) );
  AND2X1 U13353 ( .IN1(n13040), .IN2(n13039), .Q(n13036) );
  AND2X1 U13354 ( .IN1(n13041), .IN2(n13042), .Q(n13039) );
  OR2X1 U13355 ( .IN1(WX4638), .IN2(n8413), .Q(n13042) );
  INVX0 U13356 ( .INP(n13043), .ZN(n13041) );
  AND2X1 U13357 ( .IN1(n8413), .IN2(WX4638), .Q(n13043) );
  OR2X1 U13358 ( .IN1(n13044), .IN2(n13045), .Q(n13040) );
  AND2X1 U13359 ( .IN1(n8414), .IN2(WX4766), .Q(n13045) );
  AND2X1 U13360 ( .IN1(n8897), .IN2(WX4702), .Q(n13044) );
  AND2X1 U13361 ( .IN1(n9231), .IN2(CRC_OUT_7_6), .Q(n13032) );
  AND2X1 U13362 ( .IN1(n532), .IN2(n9205), .Q(n13031) );
  INVX0 U13363 ( .INP(n13046), .ZN(n532) );
  OR2X1 U13364 ( .IN1(n9564), .IN2(n3978), .Q(n13046) );
  OR4X1 U13365 ( .IN1(n13047), .IN2(n13048), .IN3(n13049), .IN4(n13050), .Q(
        WX3278) );
  AND2X1 U13366 ( .IN1(n9191), .IN2(n13051), .Q(n13050) );
  AND2X1 U13367 ( .IN1(n9266), .IN2(n12396), .Q(n13049) );
  OR2X1 U13368 ( .IN1(n13052), .IN2(n13053), .Q(n12396) );
  INVX0 U13369 ( .INP(n13054), .ZN(n13053) );
  OR2X1 U13370 ( .IN1(n13055), .IN2(n13056), .Q(n13054) );
  AND2X1 U13371 ( .IN1(n13056), .IN2(n13055), .Q(n13052) );
  AND2X1 U13372 ( .IN1(n13057), .IN2(n13058), .Q(n13055) );
  OR2X1 U13373 ( .IN1(WX4636), .IN2(n8415), .Q(n13058) );
  INVX0 U13374 ( .INP(n13059), .ZN(n13057) );
  AND2X1 U13375 ( .IN1(n8415), .IN2(WX4636), .Q(n13059) );
  OR2X1 U13376 ( .IN1(n13060), .IN2(n13061), .Q(n13056) );
  AND2X1 U13377 ( .IN1(n8416), .IN2(WX4764), .Q(n13061) );
  AND2X1 U13378 ( .IN1(n8896), .IN2(WX4700), .Q(n13060) );
  AND2X1 U13379 ( .IN1(n9231), .IN2(CRC_OUT_7_7), .Q(n13048) );
  AND2X1 U13380 ( .IN1(n531), .IN2(n9205), .Q(n13047) );
  INVX0 U13381 ( .INP(n13062), .ZN(n531) );
  OR2X1 U13382 ( .IN1(n9564), .IN2(n3979), .Q(n13062) );
  OR4X1 U13383 ( .IN1(n13063), .IN2(n13064), .IN3(n13065), .IN4(n13066), .Q(
        WX3276) );
  AND2X1 U13384 ( .IN1(n13067), .IN2(n9176), .Q(n13066) );
  AND2X1 U13385 ( .IN1(n9266), .IN2(n12412), .Q(n13065) );
  OR2X1 U13386 ( .IN1(n13068), .IN2(n13069), .Q(n12412) );
  INVX0 U13387 ( .INP(n13070), .ZN(n13069) );
  OR2X1 U13388 ( .IN1(n13071), .IN2(n13072), .Q(n13070) );
  AND2X1 U13389 ( .IN1(n13072), .IN2(n13071), .Q(n13068) );
  AND2X1 U13390 ( .IN1(n13073), .IN2(n13074), .Q(n13071) );
  OR2X1 U13391 ( .IN1(WX4634), .IN2(n8417), .Q(n13074) );
  INVX0 U13392 ( .INP(n13075), .ZN(n13073) );
  AND2X1 U13393 ( .IN1(n8417), .IN2(WX4634), .Q(n13075) );
  OR2X1 U13394 ( .IN1(n13076), .IN2(n13077), .Q(n13072) );
  AND2X1 U13395 ( .IN1(n8418), .IN2(WX4762), .Q(n13077) );
  AND2X1 U13396 ( .IN1(n8895), .IN2(WX4698), .Q(n13076) );
  AND2X1 U13397 ( .IN1(n9232), .IN2(CRC_OUT_7_8), .Q(n13064) );
  AND2X1 U13398 ( .IN1(n530), .IN2(n9205), .Q(n13063) );
  INVX0 U13399 ( .INP(n13078), .ZN(n530) );
  OR2X1 U13400 ( .IN1(n9564), .IN2(n3980), .Q(n13078) );
  OR4X1 U13401 ( .IN1(n13079), .IN2(n13080), .IN3(n13081), .IN4(n13082), .Q(
        WX3274) );
  AND2X1 U13402 ( .IN1(n9190), .IN2(n13083), .Q(n13082) );
  AND2X1 U13403 ( .IN1(n9267), .IN2(n12428), .Q(n13081) );
  OR2X1 U13404 ( .IN1(n13084), .IN2(n13085), .Q(n12428) );
  INVX0 U13405 ( .INP(n13086), .ZN(n13085) );
  OR2X1 U13406 ( .IN1(n13087), .IN2(n13088), .Q(n13086) );
  AND2X1 U13407 ( .IN1(n13088), .IN2(n13087), .Q(n13084) );
  AND2X1 U13408 ( .IN1(n13089), .IN2(n13090), .Q(n13087) );
  OR2X1 U13409 ( .IN1(WX4632), .IN2(n8419), .Q(n13090) );
  INVX0 U13410 ( .INP(n13091), .ZN(n13089) );
  AND2X1 U13411 ( .IN1(n8419), .IN2(WX4632), .Q(n13091) );
  OR2X1 U13412 ( .IN1(n13092), .IN2(n13093), .Q(n13088) );
  AND2X1 U13413 ( .IN1(n8420), .IN2(WX4760), .Q(n13093) );
  AND2X1 U13414 ( .IN1(n8894), .IN2(WX4696), .Q(n13092) );
  AND2X1 U13415 ( .IN1(n9232), .IN2(CRC_OUT_7_9), .Q(n13080) );
  AND2X1 U13416 ( .IN1(n529), .IN2(n9205), .Q(n13079) );
  INVX0 U13417 ( .INP(n13094), .ZN(n529) );
  OR2X1 U13418 ( .IN1(n9563), .IN2(n3981), .Q(n13094) );
  OR4X1 U13419 ( .IN1(n13095), .IN2(n13096), .IN3(n13097), .IN4(n13098), .Q(
        WX3272) );
  AND2X1 U13420 ( .IN1(n9190), .IN2(n13099), .Q(n13098) );
  AND2X1 U13421 ( .IN1(n9267), .IN2(n12444), .Q(n13097) );
  OR2X1 U13422 ( .IN1(n13100), .IN2(n13101), .Q(n12444) );
  INVX0 U13423 ( .INP(n13102), .ZN(n13101) );
  OR2X1 U13424 ( .IN1(n13103), .IN2(n13104), .Q(n13102) );
  AND2X1 U13425 ( .IN1(n13104), .IN2(n13103), .Q(n13100) );
  AND2X1 U13426 ( .IN1(n13105), .IN2(n13106), .Q(n13103) );
  OR2X1 U13427 ( .IN1(WX4630), .IN2(n8432), .Q(n13106) );
  INVX0 U13428 ( .INP(n13107), .ZN(n13105) );
  AND2X1 U13429 ( .IN1(n8432), .IN2(WX4630), .Q(n13107) );
  OR2X1 U13430 ( .IN1(n13108), .IN2(n13109), .Q(n13104) );
  AND2X1 U13431 ( .IN1(n8433), .IN2(WX4758), .Q(n13109) );
  AND2X1 U13432 ( .IN1(n8893), .IN2(WX4694), .Q(n13108) );
  AND2X1 U13433 ( .IN1(test_so31), .IN2(n9228), .Q(n13096) );
  AND2X1 U13434 ( .IN1(n528), .IN2(n9205), .Q(n13095) );
  INVX0 U13435 ( .INP(n13110), .ZN(n528) );
  OR2X1 U13436 ( .IN1(n9563), .IN2(n3982), .Q(n13110) );
  OR4X1 U13437 ( .IN1(n13111), .IN2(n13112), .IN3(n13113), .IN4(n13114), .Q(
        WX3270) );
  AND2X1 U13438 ( .IN1(n9190), .IN2(n13115), .Q(n13114) );
  AND2X1 U13439 ( .IN1(n12460), .IN2(n9258), .Q(n13113) );
  AND2X1 U13440 ( .IN1(n13116), .IN2(n13117), .Q(n12460) );
  INVX0 U13441 ( .INP(n13118), .ZN(n13117) );
  AND2X1 U13442 ( .IN1(n13119), .IN2(n13120), .Q(n13118) );
  OR2X1 U13443 ( .IN1(n13120), .IN2(n13119), .Q(n13116) );
  OR2X1 U13444 ( .IN1(n13121), .IN2(n13122), .Q(n13119) );
  INVX0 U13445 ( .INP(n13123), .ZN(n13122) );
  OR2X1 U13446 ( .IN1(WX4628), .IN2(n8450), .Q(n13123) );
  AND2X1 U13447 ( .IN1(n8450), .IN2(WX4628), .Q(n13121) );
  AND2X1 U13448 ( .IN1(n13124), .IN2(n13125), .Q(n13120) );
  OR2X1 U13449 ( .IN1(WX4692), .IN2(test_so41), .Q(n13125) );
  OR2X1 U13450 ( .IN1(n9088), .IN2(n8451), .Q(n13124) );
  AND2X1 U13451 ( .IN1(n9232), .IN2(CRC_OUT_7_11), .Q(n13112) );
  AND2X1 U13452 ( .IN1(n527), .IN2(n9205), .Q(n13111) );
  INVX0 U13453 ( .INP(n13126), .ZN(n527) );
  OR2X1 U13454 ( .IN1(n9563), .IN2(n3983), .Q(n13126) );
  OR4X1 U13455 ( .IN1(n13127), .IN2(n13128), .IN3(n13129), .IN4(n13130), .Q(
        WX3268) );
  AND2X1 U13456 ( .IN1(n13131), .IN2(n9176), .Q(n13130) );
  AND2X1 U13457 ( .IN1(n9267), .IN2(n12476), .Q(n13129) );
  OR2X1 U13458 ( .IN1(n13132), .IN2(n13133), .Q(n12476) );
  INVX0 U13459 ( .INP(n13134), .ZN(n13133) );
  OR2X1 U13460 ( .IN1(n13135), .IN2(n13136), .Q(n13134) );
  AND2X1 U13461 ( .IN1(n13136), .IN2(n13135), .Q(n13132) );
  AND2X1 U13462 ( .IN1(n13137), .IN2(n13138), .Q(n13135) );
  OR2X1 U13463 ( .IN1(WX4626), .IN2(n8468), .Q(n13138) );
  INVX0 U13464 ( .INP(n13139), .ZN(n13137) );
  AND2X1 U13465 ( .IN1(n8468), .IN2(WX4626), .Q(n13139) );
  OR2X1 U13466 ( .IN1(n13140), .IN2(n13141), .Q(n13136) );
  AND2X1 U13467 ( .IN1(n8469), .IN2(WX4754), .Q(n13141) );
  AND2X1 U13468 ( .IN1(n8892), .IN2(WX4690), .Q(n13140) );
  AND2X1 U13469 ( .IN1(n9232), .IN2(CRC_OUT_7_12), .Q(n13128) );
  AND2X1 U13470 ( .IN1(n526), .IN2(n9205), .Q(n13127) );
  INVX0 U13471 ( .INP(n13142), .ZN(n526) );
  OR2X1 U13472 ( .IN1(n9563), .IN2(n3984), .Q(n13142) );
  OR4X1 U13473 ( .IN1(n13143), .IN2(n13144), .IN3(n13145), .IN4(n13146), .Q(
        WX3266) );
  AND2X1 U13474 ( .IN1(n9190), .IN2(n13147), .Q(n13146) );
  AND2X1 U13475 ( .IN1(n12492), .IN2(n9258), .Q(n13145) );
  AND2X1 U13476 ( .IN1(n13148), .IN2(n13149), .Q(n12492) );
  INVX0 U13477 ( .INP(n13150), .ZN(n13149) );
  AND2X1 U13478 ( .IN1(n13151), .IN2(n13152), .Q(n13150) );
  OR2X1 U13479 ( .IN1(n13152), .IN2(n13151), .Q(n13148) );
  OR2X1 U13480 ( .IN1(n13153), .IN2(n13154), .Q(n13151) );
  INVX0 U13481 ( .INP(n13155), .ZN(n13154) );
  OR2X1 U13482 ( .IN1(WX4624), .IN2(n8471), .Q(n13155) );
  AND2X1 U13483 ( .IN1(n8471), .IN2(WX4624), .Q(n13153) );
  AND2X1 U13484 ( .IN1(n13156), .IN2(n13157), .Q(n13152) );
  OR2X1 U13485 ( .IN1(WX4752), .IN2(test_so39), .Q(n13157) );
  OR2X1 U13486 ( .IN1(n9131), .IN2(n8891), .Q(n13156) );
  AND2X1 U13487 ( .IN1(n9232), .IN2(CRC_OUT_7_13), .Q(n13144) );
  AND2X1 U13488 ( .IN1(n525), .IN2(n9206), .Q(n13143) );
  INVX0 U13489 ( .INP(n13158), .ZN(n525) );
  OR2X1 U13490 ( .IN1(n9563), .IN2(n3985), .Q(n13158) );
  OR4X1 U13491 ( .IN1(n13159), .IN2(n13160), .IN3(n13161), .IN4(n13162), .Q(
        WX3264) );
  AND2X1 U13492 ( .IN1(n9190), .IN2(n13163), .Q(n13162) );
  AND2X1 U13493 ( .IN1(n9267), .IN2(n12508), .Q(n13161) );
  OR2X1 U13494 ( .IN1(n13164), .IN2(n13165), .Q(n12508) );
  INVX0 U13495 ( .INP(n13166), .ZN(n13165) );
  OR2X1 U13496 ( .IN1(n13167), .IN2(n13168), .Q(n13166) );
  AND2X1 U13497 ( .IN1(n13168), .IN2(n13167), .Q(n13164) );
  AND2X1 U13498 ( .IN1(n13169), .IN2(n13170), .Q(n13167) );
  OR2X1 U13499 ( .IN1(WX4622), .IN2(n8472), .Q(n13170) );
  INVX0 U13500 ( .INP(n13171), .ZN(n13169) );
  AND2X1 U13501 ( .IN1(n8472), .IN2(WX4622), .Q(n13171) );
  OR2X1 U13502 ( .IN1(n13172), .IN2(n13173), .Q(n13168) );
  AND2X1 U13503 ( .IN1(n8473), .IN2(WX4750), .Q(n13173) );
  AND2X1 U13504 ( .IN1(n8890), .IN2(WX4686), .Q(n13172) );
  AND2X1 U13505 ( .IN1(n9232), .IN2(CRC_OUT_7_14), .Q(n13160) );
  AND2X1 U13506 ( .IN1(n524), .IN2(n9206), .Q(n13159) );
  INVX0 U13507 ( .INP(n13174), .ZN(n524) );
  OR2X1 U13508 ( .IN1(n9563), .IN2(n3986), .Q(n13174) );
  OR4X1 U13509 ( .IN1(n13175), .IN2(n13176), .IN3(n13177), .IN4(n13178), .Q(
        WX3262) );
  AND2X1 U13510 ( .IN1(n9190), .IN2(n13179), .Q(n13178) );
  AND2X1 U13511 ( .IN1(n12524), .IN2(n9258), .Q(n13177) );
  AND2X1 U13512 ( .IN1(n13180), .IN2(n13181), .Q(n12524) );
  INVX0 U13513 ( .INP(n13182), .ZN(n13181) );
  AND2X1 U13514 ( .IN1(n13183), .IN2(n13184), .Q(n13182) );
  OR2X1 U13515 ( .IN1(n13184), .IN2(n13183), .Q(n13180) );
  OR2X1 U13516 ( .IN1(n13185), .IN2(n13186), .Q(n13183) );
  INVX0 U13517 ( .INP(n13187), .ZN(n13186) );
  OR2X1 U13518 ( .IN1(WX4556), .IN2(n8475), .Q(n13187) );
  AND2X1 U13519 ( .IN1(n8475), .IN2(WX4556), .Q(n13185) );
  AND2X1 U13520 ( .IN1(n13188), .IN2(n13189), .Q(n13184) );
  OR2X1 U13521 ( .IN1(WX4748), .IN2(test_so37), .Q(n13189) );
  OR2X1 U13522 ( .IN1(n9132), .IN2(n8889), .Q(n13188) );
  AND2X1 U13523 ( .IN1(n9232), .IN2(CRC_OUT_7_15), .Q(n13176) );
  AND2X1 U13524 ( .IN1(n523), .IN2(n9206), .Q(n13175) );
  INVX0 U13525 ( .INP(n13190), .ZN(n523) );
  OR2X1 U13526 ( .IN1(n9563), .IN2(n3987), .Q(n13190) );
  OR4X1 U13527 ( .IN1(n13191), .IN2(n13192), .IN3(n13193), .IN4(n13194), .Q(
        WX3260) );
  AND2X1 U13528 ( .IN1(n13195), .IN2(n9177), .Q(n13194) );
  AND2X1 U13529 ( .IN1(n9267), .IN2(n12540), .Q(n13193) );
  OR2X1 U13530 ( .IN1(n13196), .IN2(n13197), .Q(n12540) );
  INVX0 U13531 ( .INP(n13198), .ZN(n13197) );
  OR2X1 U13532 ( .IN1(n13199), .IN2(n13200), .Q(n13198) );
  AND2X1 U13533 ( .IN1(n13200), .IN2(n13199), .Q(n13196) );
  AND2X1 U13534 ( .IN1(n13201), .IN2(n13202), .Q(n13199) );
  OR2X1 U13535 ( .IN1(n9462), .IN2(n8032), .Q(n13202) );
  OR2X1 U13536 ( .IN1(WX4618), .IN2(n9446), .Q(n13201) );
  OR2X1 U13537 ( .IN1(n13203), .IN2(n13204), .Q(n13200) );
  INVX0 U13538 ( .INP(n13205), .ZN(n13204) );
  OR2X1 U13539 ( .IN1(n13206), .IN2(n8033), .Q(n13205) );
  AND2X1 U13540 ( .IN1(n8033), .IN2(n13206), .Q(n13203) );
  INVX0 U13541 ( .INP(n13207), .ZN(n13206) );
  OR2X1 U13542 ( .IN1(n13208), .IN2(n13209), .Q(n13207) );
  AND2X1 U13543 ( .IN1(n8726), .IN2(n8537), .Q(n13209) );
  AND2X1 U13544 ( .IN1(n15938), .IN2(WX4746), .Q(n13208) );
  AND2X1 U13545 ( .IN1(n9232), .IN2(CRC_OUT_7_16), .Q(n13192) );
  AND2X1 U13546 ( .IN1(n522), .IN2(n9206), .Q(n13191) );
  INVX0 U13547 ( .INP(n13210), .ZN(n522) );
  OR2X1 U13548 ( .IN1(n9563), .IN2(n3988), .Q(n13210) );
  OR4X1 U13549 ( .IN1(n13211), .IN2(n13212), .IN3(n13213), .IN4(n13214), .Q(
        WX3258) );
  AND2X1 U13550 ( .IN1(n9190), .IN2(n13215), .Q(n13214) );
  AND2X1 U13551 ( .IN1(n12559), .IN2(n9258), .Q(n13213) );
  AND2X1 U13552 ( .IN1(n13216), .IN2(n13217), .Q(n12559) );
  OR2X1 U13553 ( .IN1(n13218), .IN2(n13219), .Q(n13217) );
  INVX0 U13554 ( .INP(n13220), .ZN(n13216) );
  AND2X1 U13555 ( .IN1(n13219), .IN2(n13218), .Q(n13220) );
  INVX0 U13556 ( .INP(n13221), .ZN(n13218) );
  OR2X1 U13557 ( .IN1(n13222), .IN2(n13223), .Q(n13221) );
  AND2X1 U13558 ( .IN1(n9451), .IN2(WX4744), .Q(n13223) );
  AND2X1 U13559 ( .IN1(n8888), .IN2(n9460), .Q(n13222) );
  OR2X1 U13560 ( .IN1(n13224), .IN2(n13225), .Q(n13219) );
  AND3X1 U13561 ( .IN1(n13226), .IN2(n13227), .IN3(n8035), .Q(n13225) );
  OR2X1 U13562 ( .IN1(n8034), .IN2(n9094), .Q(n13227) );
  OR2X1 U13563 ( .IN1(test_so35), .IN2(WX4616), .Q(n13226) );
  AND2X1 U13564 ( .IN1(n13228), .IN2(WX4680), .Q(n13224) );
  OR2X1 U13565 ( .IN1(n13229), .IN2(n13230), .Q(n13228) );
  AND2X1 U13566 ( .IN1(n8034), .IN2(n9094), .Q(n13230) );
  AND2X1 U13567 ( .IN1(test_so35), .IN2(WX4616), .Q(n13229) );
  AND2X1 U13568 ( .IN1(n9232), .IN2(CRC_OUT_7_17), .Q(n13212) );
  AND2X1 U13569 ( .IN1(n521), .IN2(n9206), .Q(n13211) );
  INVX0 U13570 ( .INP(n13231), .ZN(n521) );
  OR2X1 U13571 ( .IN1(n9563), .IN2(n3989), .Q(n13231) );
  OR4X1 U13572 ( .IN1(n13232), .IN2(n13233), .IN3(n13234), .IN4(n13235), .Q(
        WX3256) );
  AND2X1 U13573 ( .IN1(n9190), .IN2(n13236), .Q(n13235) );
  AND2X1 U13574 ( .IN1(n9267), .IN2(n12579), .Q(n13234) );
  OR2X1 U13575 ( .IN1(n13237), .IN2(n13238), .Q(n12579) );
  INVX0 U13576 ( .INP(n13239), .ZN(n13238) );
  OR2X1 U13577 ( .IN1(n13240), .IN2(n13241), .Q(n13239) );
  AND2X1 U13578 ( .IN1(n13241), .IN2(n13240), .Q(n13237) );
  AND2X1 U13579 ( .IN1(n13242), .IN2(n13243), .Q(n13240) );
  OR2X1 U13580 ( .IN1(n9482), .IN2(n8036), .Q(n13243) );
  OR2X1 U13581 ( .IN1(WX4614), .IN2(n9445), .Q(n13242) );
  OR2X1 U13582 ( .IN1(n13244), .IN2(n13245), .Q(n13241) );
  INVX0 U13583 ( .INP(n13246), .ZN(n13245) );
  OR2X1 U13584 ( .IN1(n13247), .IN2(n8037), .Q(n13246) );
  AND2X1 U13585 ( .IN1(n8037), .IN2(n13247), .Q(n13244) );
  INVX0 U13586 ( .INP(n13248), .ZN(n13247) );
  OR2X1 U13587 ( .IN1(n13249), .IN2(n13250), .Q(n13248) );
  AND2X1 U13588 ( .IN1(n8887), .IN2(n8540), .Q(n13250) );
  AND2X1 U13589 ( .IN1(n15939), .IN2(WX4742), .Q(n13249) );
  AND2X1 U13590 ( .IN1(n9233), .IN2(CRC_OUT_7_18), .Q(n13233) );
  AND2X1 U13591 ( .IN1(n520), .IN2(n9206), .Q(n13232) );
  INVX0 U13592 ( .INP(n13251), .ZN(n520) );
  OR2X1 U13593 ( .IN1(n9563), .IN2(n3990), .Q(n13251) );
  OR4X1 U13594 ( .IN1(n13252), .IN2(n13253), .IN3(n13254), .IN4(n13255), .Q(
        WX3254) );
  AND2X1 U13595 ( .IN1(n9190), .IN2(n13256), .Q(n13255) );
  AND2X1 U13596 ( .IN1(n9267), .IN2(n12598), .Q(n13254) );
  OR2X1 U13597 ( .IN1(n13257), .IN2(n13258), .Q(n12598) );
  INVX0 U13598 ( .INP(n13259), .ZN(n13258) );
  OR2X1 U13599 ( .IN1(n13260), .IN2(n13261), .Q(n13259) );
  AND2X1 U13600 ( .IN1(n13261), .IN2(n13260), .Q(n13257) );
  AND2X1 U13601 ( .IN1(n13262), .IN2(n13263), .Q(n13260) );
  OR2X1 U13602 ( .IN1(n9453), .IN2(n8038), .Q(n13263) );
  OR2X1 U13603 ( .IN1(WX4612), .IN2(n9445), .Q(n13262) );
  OR2X1 U13604 ( .IN1(n13264), .IN2(n13265), .Q(n13261) );
  INVX0 U13605 ( .INP(n13266), .ZN(n13265) );
  OR2X1 U13606 ( .IN1(n13267), .IN2(n8039), .Q(n13266) );
  AND2X1 U13607 ( .IN1(n8039), .IN2(n13267), .Q(n13264) );
  INVX0 U13608 ( .INP(n13268), .ZN(n13267) );
  OR2X1 U13609 ( .IN1(n13269), .IN2(n13270), .Q(n13268) );
  AND2X1 U13610 ( .IN1(n8886), .IN2(n8541), .Q(n13270) );
  AND2X1 U13611 ( .IN1(n15940), .IN2(WX4740), .Q(n13269) );
  AND2X1 U13612 ( .IN1(n9232), .IN2(CRC_OUT_7_19), .Q(n13253) );
  AND2X1 U13613 ( .IN1(n519), .IN2(n9206), .Q(n13252) );
  INVX0 U13614 ( .INP(n13271), .ZN(n519) );
  OR2X1 U13615 ( .IN1(n9563), .IN2(n3991), .Q(n13271) );
  OR4X1 U13616 ( .IN1(n13272), .IN2(n13273), .IN3(n13274), .IN4(n13275), .Q(
        WX3252) );
  AND2X1 U13617 ( .IN1(n9190), .IN2(n13276), .Q(n13275) );
  AND2X1 U13618 ( .IN1(n9267), .IN2(n12618), .Q(n13274) );
  OR2X1 U13619 ( .IN1(n13277), .IN2(n13278), .Q(n12618) );
  INVX0 U13620 ( .INP(n13279), .ZN(n13278) );
  OR2X1 U13621 ( .IN1(n13280), .IN2(n13281), .Q(n13279) );
  AND2X1 U13622 ( .IN1(n13281), .IN2(n13280), .Q(n13277) );
  AND2X1 U13623 ( .IN1(n13282), .IN2(n13283), .Q(n13280) );
  OR2X1 U13624 ( .IN1(n9454), .IN2(n8040), .Q(n13283) );
  OR2X1 U13625 ( .IN1(WX4610), .IN2(n9445), .Q(n13282) );
  OR2X1 U13626 ( .IN1(n13284), .IN2(n13285), .Q(n13281) );
  INVX0 U13627 ( .INP(n13286), .ZN(n13285) );
  OR2X1 U13628 ( .IN1(n13287), .IN2(n8041), .Q(n13286) );
  AND2X1 U13629 ( .IN1(n8041), .IN2(n13287), .Q(n13284) );
  INVX0 U13630 ( .INP(n13288), .ZN(n13287) );
  OR2X1 U13631 ( .IN1(n13289), .IN2(n13290), .Q(n13288) );
  AND2X1 U13632 ( .IN1(n8885), .IN2(n8542), .Q(n13290) );
  AND2X1 U13633 ( .IN1(n15941), .IN2(WX4738), .Q(n13289) );
  AND2X1 U13634 ( .IN1(n9233), .IN2(CRC_OUT_7_20), .Q(n13273) );
  AND2X1 U13635 ( .IN1(n518), .IN2(n9206), .Q(n13272) );
  INVX0 U13636 ( .INP(n13291), .ZN(n518) );
  OR2X1 U13637 ( .IN1(n9563), .IN2(n3992), .Q(n13291) );
  OR4X1 U13638 ( .IN1(n13292), .IN2(n13293), .IN3(n13294), .IN4(n13295), .Q(
        WX3250) );
  AND2X1 U13639 ( .IN1(n9190), .IN2(n13296), .Q(n13295) );
  AND2X1 U13640 ( .IN1(n9267), .IN2(n12637), .Q(n13294) );
  OR2X1 U13641 ( .IN1(n13297), .IN2(n13298), .Q(n12637) );
  INVX0 U13642 ( .INP(n13299), .ZN(n13298) );
  OR2X1 U13643 ( .IN1(n13300), .IN2(n13301), .Q(n13299) );
  AND2X1 U13644 ( .IN1(n13301), .IN2(n13300), .Q(n13297) );
  AND2X1 U13645 ( .IN1(n13302), .IN2(n13303), .Q(n13300) );
  OR2X1 U13646 ( .IN1(n9456), .IN2(n8042), .Q(n13303) );
  OR2X1 U13647 ( .IN1(WX4608), .IN2(n9445), .Q(n13302) );
  OR2X1 U13648 ( .IN1(n13304), .IN2(n13305), .Q(n13301) );
  INVX0 U13649 ( .INP(n13306), .ZN(n13305) );
  OR2X1 U13650 ( .IN1(n13307), .IN2(n8043), .Q(n13306) );
  AND2X1 U13651 ( .IN1(n8043), .IN2(n13307), .Q(n13304) );
  INVX0 U13652 ( .INP(n13308), .ZN(n13307) );
  OR2X1 U13653 ( .IN1(n13309), .IN2(n13310), .Q(n13308) );
  AND2X1 U13654 ( .IN1(n8884), .IN2(n8543), .Q(n13310) );
  AND2X1 U13655 ( .IN1(n15942), .IN2(WX4736), .Q(n13309) );
  AND2X1 U13656 ( .IN1(n9233), .IN2(CRC_OUT_7_21), .Q(n13293) );
  AND2X1 U13657 ( .IN1(n517), .IN2(n9206), .Q(n13292) );
  INVX0 U13658 ( .INP(n13311), .ZN(n517) );
  OR2X1 U13659 ( .IN1(n9562), .IN2(n3993), .Q(n13311) );
  OR4X1 U13660 ( .IN1(n13312), .IN2(n13313), .IN3(n13314), .IN4(n13315), .Q(
        WX3248) );
  AND2X1 U13661 ( .IN1(n9190), .IN2(n13316), .Q(n13315) );
  AND2X1 U13662 ( .IN1(n9267), .IN2(n12657), .Q(n13314) );
  OR2X1 U13663 ( .IN1(n13317), .IN2(n13318), .Q(n12657) );
  INVX0 U13664 ( .INP(n13319), .ZN(n13318) );
  OR2X1 U13665 ( .IN1(n13320), .IN2(n13321), .Q(n13319) );
  AND2X1 U13666 ( .IN1(n13321), .IN2(n13320), .Q(n13317) );
  AND2X1 U13667 ( .IN1(n13322), .IN2(n13323), .Q(n13320) );
  OR2X1 U13668 ( .IN1(n9457), .IN2(n8044), .Q(n13323) );
  OR2X1 U13669 ( .IN1(WX4606), .IN2(n9445), .Q(n13322) );
  OR2X1 U13670 ( .IN1(n13324), .IN2(n13325), .Q(n13321) );
  INVX0 U13671 ( .INP(n13326), .ZN(n13325) );
  OR2X1 U13672 ( .IN1(n13327), .IN2(n8045), .Q(n13326) );
  AND2X1 U13673 ( .IN1(n8045), .IN2(n13327), .Q(n13324) );
  INVX0 U13674 ( .INP(n13328), .ZN(n13327) );
  OR2X1 U13675 ( .IN1(n13329), .IN2(n13330), .Q(n13328) );
  AND2X1 U13676 ( .IN1(n8883), .IN2(n8544), .Q(n13330) );
  AND2X1 U13677 ( .IN1(n15943), .IN2(WX4734), .Q(n13329) );
  AND2X1 U13678 ( .IN1(n9233), .IN2(CRC_OUT_7_22), .Q(n13313) );
  AND2X1 U13679 ( .IN1(n516), .IN2(n9206), .Q(n13312) );
  INVX0 U13680 ( .INP(n13331), .ZN(n516) );
  OR2X1 U13681 ( .IN1(n9562), .IN2(n3994), .Q(n13331) );
  OR4X1 U13682 ( .IN1(n13332), .IN2(n13333), .IN3(n13334), .IN4(n13335), .Q(
        WX3246) );
  AND2X1 U13683 ( .IN1(n13336), .IN2(n9178), .Q(n13335) );
  AND2X1 U13684 ( .IN1(n9270), .IN2(n12678), .Q(n13334) );
  OR2X1 U13685 ( .IN1(n13337), .IN2(n13338), .Q(n12678) );
  AND2X1 U13686 ( .IN1(n13339), .IN2(n13340), .Q(n13338) );
  INVX0 U13687 ( .INP(n13341), .ZN(n13340) );
  AND2X1 U13688 ( .IN1(n13341), .IN2(n13342), .Q(n13337) );
  INVX0 U13689 ( .INP(n13339), .ZN(n13342) );
  OR2X1 U13690 ( .IN1(n13343), .IN2(n13344), .Q(n13339) );
  AND2X1 U13691 ( .IN1(n9450), .IN2(n8545), .Q(n13344) );
  AND2X1 U13692 ( .IN1(n15944), .IN2(n9468), .Q(n13343) );
  OR2X1 U13693 ( .IN1(n13345), .IN2(n13346), .Q(n13341) );
  AND3X1 U13694 ( .IN1(n13347), .IN2(n13348), .IN3(n8882), .Q(n13346) );
  OR2X1 U13695 ( .IN1(n8046), .IN2(WX4668), .Q(n13348) );
  OR2X1 U13696 ( .IN1(n8047), .IN2(WX4604), .Q(n13347) );
  AND2X1 U13697 ( .IN1(n13349), .IN2(WX4732), .Q(n13345) );
  OR2X1 U13698 ( .IN1(n13350), .IN2(n13351), .Q(n13349) );
  AND2X1 U13699 ( .IN1(n8046), .IN2(WX4668), .Q(n13351) );
  AND2X1 U13700 ( .IN1(n8047), .IN2(WX4604), .Q(n13350) );
  AND2X1 U13701 ( .IN1(n9238), .IN2(CRC_OUT_7_23), .Q(n13333) );
  AND2X1 U13702 ( .IN1(n515), .IN2(n9206), .Q(n13332) );
  INVX0 U13703 ( .INP(n13352), .ZN(n515) );
  OR2X1 U13704 ( .IN1(n9562), .IN2(n3995), .Q(n13352) );
  OR4X1 U13705 ( .IN1(n13353), .IN2(n13354), .IN3(n13355), .IN4(n13356), .Q(
        WX3244) );
  AND2X1 U13706 ( .IN1(n9189), .IN2(n13357), .Q(n13356) );
  AND2X1 U13707 ( .IN1(n9267), .IN2(n12698), .Q(n13355) );
  OR2X1 U13708 ( .IN1(n13358), .IN2(n13359), .Q(n12698) );
  INVX0 U13709 ( .INP(n13360), .ZN(n13359) );
  OR2X1 U13710 ( .IN1(n13361), .IN2(n13362), .Q(n13360) );
  AND2X1 U13711 ( .IN1(n13362), .IN2(n13361), .Q(n13358) );
  AND2X1 U13712 ( .IN1(n13363), .IN2(n13364), .Q(n13361) );
  OR2X1 U13713 ( .IN1(n9478), .IN2(n8048), .Q(n13364) );
  OR2X1 U13714 ( .IN1(WX4602), .IN2(n9445), .Q(n13363) );
  OR2X1 U13715 ( .IN1(n13365), .IN2(n13366), .Q(n13362) );
  INVX0 U13716 ( .INP(n13367), .ZN(n13366) );
  OR2X1 U13717 ( .IN1(n13368), .IN2(n8049), .Q(n13367) );
  AND2X1 U13718 ( .IN1(n8049), .IN2(n13368), .Q(n13365) );
  INVX0 U13719 ( .INP(n13369), .ZN(n13368) );
  OR2X1 U13720 ( .IN1(n13370), .IN2(n13371), .Q(n13369) );
  AND2X1 U13721 ( .IN1(n8881), .IN2(n8546), .Q(n13371) );
  AND2X1 U13722 ( .IN1(n15945), .IN2(WX4730), .Q(n13370) );
  AND2X1 U13723 ( .IN1(n9233), .IN2(CRC_OUT_7_24), .Q(n13354) );
  AND2X1 U13724 ( .IN1(n514), .IN2(n9207), .Q(n13353) );
  INVX0 U13725 ( .INP(n13372), .ZN(n514) );
  OR2X1 U13726 ( .IN1(n9562), .IN2(n3996), .Q(n13372) );
  OR4X1 U13727 ( .IN1(n13373), .IN2(n13374), .IN3(n13375), .IN4(n13376), .Q(
        WX3242) );
  AND2X1 U13728 ( .IN1(n9189), .IN2(n13377), .Q(n13376) );
  AND2X1 U13729 ( .IN1(n9267), .IN2(n12718), .Q(n13375) );
  OR2X1 U13730 ( .IN1(n13378), .IN2(n13379), .Q(n12718) );
  INVX0 U13731 ( .INP(n13380), .ZN(n13379) );
  OR2X1 U13732 ( .IN1(n13381), .IN2(n13382), .Q(n13380) );
  AND2X1 U13733 ( .IN1(n13382), .IN2(n13381), .Q(n13378) );
  AND2X1 U13734 ( .IN1(n13383), .IN2(n13384), .Q(n13381) );
  OR2X1 U13735 ( .IN1(n9466), .IN2(n8050), .Q(n13384) );
  OR2X1 U13736 ( .IN1(WX4600), .IN2(n9445), .Q(n13383) );
  OR2X1 U13737 ( .IN1(n13385), .IN2(n13386), .Q(n13382) );
  INVX0 U13738 ( .INP(n13387), .ZN(n13386) );
  OR2X1 U13739 ( .IN1(n13388), .IN2(n8051), .Q(n13387) );
  AND2X1 U13740 ( .IN1(n8051), .IN2(n13388), .Q(n13385) );
  INVX0 U13741 ( .INP(n13389), .ZN(n13388) );
  OR2X1 U13742 ( .IN1(n13390), .IN2(n13391), .Q(n13389) );
  AND2X1 U13743 ( .IN1(n8880), .IN2(n8547), .Q(n13391) );
  AND2X1 U13744 ( .IN1(n15946), .IN2(WX4728), .Q(n13390) );
  AND2X1 U13745 ( .IN1(n9233), .IN2(CRC_OUT_7_25), .Q(n13374) );
  AND2X1 U13746 ( .IN1(n513), .IN2(n9207), .Q(n13373) );
  INVX0 U13747 ( .INP(n13392), .ZN(n513) );
  OR2X1 U13748 ( .IN1(n9562), .IN2(n3997), .Q(n13392) );
  OR4X1 U13749 ( .IN1(n13393), .IN2(n13394), .IN3(n13395), .IN4(n13396), .Q(
        WX3240) );
  AND2X1 U13750 ( .IN1(n13397), .IN2(n9177), .Q(n13396) );
  AND2X1 U13751 ( .IN1(n9267), .IN2(n12738), .Q(n13395) );
  OR2X1 U13752 ( .IN1(n13398), .IN2(n13399), .Q(n12738) );
  INVX0 U13753 ( .INP(n13400), .ZN(n13399) );
  OR2X1 U13754 ( .IN1(n13401), .IN2(n13402), .Q(n13400) );
  AND2X1 U13755 ( .IN1(n13402), .IN2(n13401), .Q(n13398) );
  AND2X1 U13756 ( .IN1(n13403), .IN2(n13404), .Q(n13401) );
  OR2X1 U13757 ( .IN1(n9467), .IN2(n8052), .Q(n13404) );
  OR2X1 U13758 ( .IN1(WX4598), .IN2(n9445), .Q(n13403) );
  OR2X1 U13759 ( .IN1(n13405), .IN2(n13406), .Q(n13402) );
  INVX0 U13760 ( .INP(n13407), .ZN(n13406) );
  OR2X1 U13761 ( .IN1(n13408), .IN2(n8053), .Q(n13407) );
  AND2X1 U13762 ( .IN1(n8053), .IN2(n13408), .Q(n13405) );
  INVX0 U13763 ( .INP(n13409), .ZN(n13408) );
  OR2X1 U13764 ( .IN1(n13410), .IN2(n13411), .Q(n13409) );
  AND2X1 U13765 ( .IN1(n8879), .IN2(n8548), .Q(n13411) );
  AND2X1 U13766 ( .IN1(n15947), .IN2(WX4726), .Q(n13410) );
  AND2X1 U13767 ( .IN1(n9233), .IN2(CRC_OUT_7_26), .Q(n13394) );
  AND2X1 U13768 ( .IN1(n512), .IN2(n9207), .Q(n13393) );
  INVX0 U13769 ( .INP(n13412), .ZN(n512) );
  OR2X1 U13770 ( .IN1(n9562), .IN2(n3998), .Q(n13412) );
  OR4X1 U13771 ( .IN1(n13413), .IN2(n13414), .IN3(n13415), .IN4(n13416), .Q(
        WX3238) );
  AND2X1 U13772 ( .IN1(n9189), .IN2(n13417), .Q(n13416) );
  AND2X1 U13773 ( .IN1(n9268), .IN2(n12758), .Q(n13415) );
  OR2X1 U13774 ( .IN1(n13418), .IN2(n13419), .Q(n12758) );
  INVX0 U13775 ( .INP(n13420), .ZN(n13419) );
  OR2X1 U13776 ( .IN1(n13421), .IN2(n13422), .Q(n13420) );
  AND2X1 U13777 ( .IN1(n13422), .IN2(n13421), .Q(n13418) );
  AND2X1 U13778 ( .IN1(n13423), .IN2(n13424), .Q(n13421) );
  OR2X1 U13779 ( .IN1(n9471), .IN2(n8054), .Q(n13424) );
  OR2X1 U13780 ( .IN1(WX4596), .IN2(n9445), .Q(n13423) );
  OR2X1 U13781 ( .IN1(n13425), .IN2(n13426), .Q(n13422) );
  INVX0 U13782 ( .INP(n13427), .ZN(n13426) );
  OR2X1 U13783 ( .IN1(n13428), .IN2(n8055), .Q(n13427) );
  AND2X1 U13784 ( .IN1(n8055), .IN2(n13428), .Q(n13425) );
  INVX0 U13785 ( .INP(n13429), .ZN(n13428) );
  OR2X1 U13786 ( .IN1(n13430), .IN2(n13431), .Q(n13429) );
  AND2X1 U13787 ( .IN1(n8878), .IN2(n8549), .Q(n13431) );
  AND2X1 U13788 ( .IN1(n15948), .IN2(WX4724), .Q(n13430) );
  AND2X1 U13789 ( .IN1(test_so32), .IN2(n9227), .Q(n13414) );
  AND2X1 U13790 ( .IN1(n511), .IN2(n9207), .Q(n13413) );
  INVX0 U13791 ( .INP(n13432), .ZN(n511) );
  OR2X1 U13792 ( .IN1(n9562), .IN2(n3999), .Q(n13432) );
  OR4X1 U13793 ( .IN1(n13433), .IN2(n13434), .IN3(n13435), .IN4(n13436), .Q(
        WX3236) );
  AND2X1 U13794 ( .IN1(n9189), .IN2(n13437), .Q(n13436) );
  AND2X1 U13795 ( .IN1(n12778), .IN2(n9259), .Q(n13435) );
  AND2X1 U13796 ( .IN1(n13438), .IN2(n13439), .Q(n12778) );
  INVX0 U13797 ( .INP(n13440), .ZN(n13439) );
  AND2X1 U13798 ( .IN1(n13441), .IN2(n13442), .Q(n13440) );
  OR2X1 U13799 ( .IN1(n13442), .IN2(n13441), .Q(n13438) );
  OR2X1 U13800 ( .IN1(n13443), .IN2(n13444), .Q(n13441) );
  AND2X1 U13801 ( .IN1(n9450), .IN2(WX4594), .Q(n13444) );
  AND2X1 U13802 ( .IN1(n8056), .IN2(n9461), .Q(n13443) );
  AND2X1 U13803 ( .IN1(n13445), .IN2(n13446), .Q(n13442) );
  OR2X1 U13804 ( .IN1(n13447), .IN2(n8057), .Q(n13446) );
  INVX0 U13805 ( .INP(n13448), .ZN(n13447) );
  OR2X1 U13806 ( .IN1(WX4658), .IN2(n13448), .Q(n13445) );
  OR2X1 U13807 ( .IN1(n13449), .IN2(n13450), .Q(n13448) );
  AND2X1 U13808 ( .IN1(n15949), .IN2(n9106), .Q(n13450) );
  AND2X1 U13809 ( .IN1(test_so40), .IN2(n8550), .Q(n13449) );
  AND2X1 U13810 ( .IN1(n9233), .IN2(CRC_OUT_7_28), .Q(n13434) );
  AND2X1 U13811 ( .IN1(n510), .IN2(n9207), .Q(n13433) );
  INVX0 U13812 ( .INP(n13451), .ZN(n510) );
  OR2X1 U13813 ( .IN1(n9562), .IN2(n4000), .Q(n13451) );
  OR4X1 U13814 ( .IN1(n13452), .IN2(n13453), .IN3(n13454), .IN4(n13455), .Q(
        WX3234) );
  AND2X1 U13815 ( .IN1(n9189), .IN2(n13456), .Q(n13455) );
  AND2X1 U13816 ( .IN1(n9268), .IN2(n12798), .Q(n13454) );
  OR2X1 U13817 ( .IN1(n13457), .IN2(n13458), .Q(n12798) );
  INVX0 U13818 ( .INP(n13459), .ZN(n13458) );
  OR2X1 U13819 ( .IN1(n13460), .IN2(n13461), .Q(n13459) );
  AND2X1 U13820 ( .IN1(n13461), .IN2(n13460), .Q(n13457) );
  AND2X1 U13821 ( .IN1(n13462), .IN2(n13463), .Q(n13460) );
  OR2X1 U13822 ( .IN1(n9468), .IN2(n8058), .Q(n13463) );
  OR2X1 U13823 ( .IN1(WX4592), .IN2(n9445), .Q(n13462) );
  OR2X1 U13824 ( .IN1(n13464), .IN2(n13465), .Q(n13461) );
  INVX0 U13825 ( .INP(n13466), .ZN(n13465) );
  OR2X1 U13826 ( .IN1(n13467), .IN2(n8059), .Q(n13466) );
  AND2X1 U13827 ( .IN1(n8059), .IN2(n13467), .Q(n13464) );
  INVX0 U13828 ( .INP(n13468), .ZN(n13467) );
  OR2X1 U13829 ( .IN1(n13469), .IN2(n13470), .Q(n13468) );
  AND2X1 U13830 ( .IN1(n8877), .IN2(n8551), .Q(n13470) );
  AND2X1 U13831 ( .IN1(n15950), .IN2(WX4720), .Q(n13469) );
  AND2X1 U13832 ( .IN1(n9233), .IN2(CRC_OUT_7_29), .Q(n13453) );
  AND2X1 U13833 ( .IN1(n509), .IN2(n9207), .Q(n13452) );
  INVX0 U13834 ( .INP(n13471), .ZN(n509) );
  OR2X1 U13835 ( .IN1(n9562), .IN2(n4001), .Q(n13471) );
  OR4X1 U13836 ( .IN1(n13472), .IN2(n13473), .IN3(n13474), .IN4(n13475), .Q(
        WX3232) );
  AND2X1 U13837 ( .IN1(n13476), .IN2(n9177), .Q(n13475) );
  AND2X1 U13838 ( .IN1(n12818), .IN2(n9259), .Q(n13474) );
  AND2X1 U13839 ( .IN1(n13477), .IN2(n13478), .Q(n12818) );
  INVX0 U13840 ( .INP(n13479), .ZN(n13478) );
  AND2X1 U13841 ( .IN1(n13480), .IN2(n13481), .Q(n13479) );
  OR2X1 U13842 ( .IN1(n13481), .IN2(n13480), .Q(n13477) );
  OR2X1 U13843 ( .IN1(n13482), .IN2(n13483), .Q(n13480) );
  AND2X1 U13844 ( .IN1(n9450), .IN2(WX4590), .Q(n13483) );
  AND2X1 U13845 ( .IN1(n8060), .IN2(n9462), .Q(n13482) );
  AND2X1 U13846 ( .IN1(n13484), .IN2(n13485), .Q(n13481) );
  OR2X1 U13847 ( .IN1(n13486), .IN2(n8876), .Q(n13485) );
  OR2X1 U13848 ( .IN1(WX4718), .IN2(n13487), .Q(n13484) );
  INVX0 U13849 ( .INP(n13486), .ZN(n13487) );
  AND2X1 U13850 ( .IN1(n13488), .IN2(n13489), .Q(n13486) );
  OR2X1 U13851 ( .IN1(n8552), .IN2(test_so38), .Q(n13489) );
  OR2X1 U13852 ( .IN1(n9133), .IN2(n15951), .Q(n13488) );
  AND2X1 U13853 ( .IN1(n9233), .IN2(CRC_OUT_7_30), .Q(n13473) );
  AND2X1 U13854 ( .IN1(n508), .IN2(n9207), .Q(n13472) );
  INVX0 U13855 ( .INP(n13490), .ZN(n508) );
  OR2X1 U13856 ( .IN1(n9562), .IN2(n4002), .Q(n13490) );
  OR4X1 U13857 ( .IN1(n13491), .IN2(n13492), .IN3(n13493), .IN4(n13494), .Q(
        WX3230) );
  AND2X1 U13858 ( .IN1(n9189), .IN2(n13495), .Q(n13494) );
  AND2X1 U13859 ( .IN1(n9268), .IN2(n12838), .Q(n13493) );
  OR2X1 U13860 ( .IN1(n13496), .IN2(n13497), .Q(n12838) );
  INVX0 U13861 ( .INP(n13498), .ZN(n13497) );
  OR2X1 U13862 ( .IN1(n13499), .IN2(n13500), .Q(n13498) );
  AND2X1 U13863 ( .IN1(n13500), .IN2(n13499), .Q(n13496) );
  AND2X1 U13864 ( .IN1(n13501), .IN2(n13502), .Q(n13499) );
  OR2X1 U13865 ( .IN1(n9458), .IN2(n7886), .Q(n13502) );
  OR2X1 U13866 ( .IN1(WX4588), .IN2(n9445), .Q(n13501) );
  OR2X1 U13867 ( .IN1(n13503), .IN2(n13504), .Q(n13500) );
  INVX0 U13868 ( .INP(n13505), .ZN(n13504) );
  OR2X1 U13869 ( .IN1(n13506), .IN2(n7887), .Q(n13505) );
  AND2X1 U13870 ( .IN1(n7887), .IN2(n13506), .Q(n13503) );
  INVX0 U13871 ( .INP(n13507), .ZN(n13506) );
  OR2X1 U13872 ( .IN1(n13508), .IN2(n13509), .Q(n13507) );
  AND2X1 U13873 ( .IN1(n8875), .IN2(n8553), .Q(n13509) );
  AND2X1 U13874 ( .IN1(n15952), .IN2(WX4716), .Q(n13508) );
  AND2X1 U13875 ( .IN1(n2245), .IN2(WX3071), .Q(n13492) );
  AND2X1 U13876 ( .IN1(n9233), .IN2(CRC_OUT_7_31), .Q(n13491) );
  AND2X1 U13877 ( .IN1(n9046), .IN2(n9495), .Q(WX3132) );
  AND3X1 U13878 ( .IN1(n13510), .IN2(n13511), .IN3(n9526), .Q(WX2619) );
  OR2X1 U13879 ( .IN1(DFF_382_n1), .IN2(WX2130), .Q(n13511) );
  OR2X1 U13880 ( .IN1(n8928), .IN2(CRC_OUT_8_30), .Q(n13510) );
  AND3X1 U13881 ( .IN1(n13512), .IN2(n13513), .IN3(n9526), .Q(WX2617) );
  OR2X1 U13882 ( .IN1(DFF_381_n1), .IN2(WX2132), .Q(n13513) );
  OR2X1 U13883 ( .IN1(n8929), .IN2(CRC_OUT_8_29), .Q(n13512) );
  AND3X1 U13884 ( .IN1(n13514), .IN2(n13515), .IN3(n9526), .Q(WX2615) );
  OR2X1 U13885 ( .IN1(DFF_380_n1), .IN2(WX2134), .Q(n13515) );
  OR2X1 U13886 ( .IN1(n8930), .IN2(CRC_OUT_8_28), .Q(n13514) );
  AND2X1 U13887 ( .IN1(n13516), .IN2(n9496), .Q(WX2613) );
  OR2X1 U13888 ( .IN1(n13517), .IN2(n13518), .Q(n13516) );
  AND2X1 U13889 ( .IN1(DFF_379_n1), .IN2(n9108), .Q(n13518) );
  AND2X1 U13890 ( .IN1(test_so18), .IN2(CRC_OUT_8_27), .Q(n13517) );
  AND3X1 U13891 ( .IN1(n13519), .IN2(n13520), .IN3(n9526), .Q(WX2611) );
  OR2X1 U13892 ( .IN1(DFF_378_n1), .IN2(WX2138), .Q(n13520) );
  OR2X1 U13893 ( .IN1(n8931), .IN2(CRC_OUT_8_26), .Q(n13519) );
  AND2X1 U13894 ( .IN1(n13521), .IN2(n9497), .Q(WX2609) );
  OR2X1 U13895 ( .IN1(n13522), .IN2(n13523), .Q(n13521) );
  AND2X1 U13896 ( .IN1(n8932), .IN2(n9159), .Q(n13523) );
  AND2X1 U13897 ( .IN1(test_so21), .IN2(WX2140), .Q(n13522) );
  AND3X1 U13898 ( .IN1(n13524), .IN2(n13525), .IN3(n9526), .Q(WX2607) );
  OR2X1 U13899 ( .IN1(DFF_376_n1), .IN2(WX2142), .Q(n13525) );
  OR2X1 U13900 ( .IN1(n8933), .IN2(CRC_OUT_8_24), .Q(n13524) );
  AND3X1 U13901 ( .IN1(n13526), .IN2(n13527), .IN3(n9525), .Q(WX2605) );
  OR2X1 U13902 ( .IN1(DFF_375_n1), .IN2(WX2144), .Q(n13527) );
  OR2X1 U13903 ( .IN1(n8934), .IN2(CRC_OUT_8_23), .Q(n13526) );
  AND3X1 U13904 ( .IN1(n13528), .IN2(n13529), .IN3(n9525), .Q(WX2603) );
  OR2X1 U13905 ( .IN1(DFF_374_n1), .IN2(WX2146), .Q(n13529) );
  OR2X1 U13906 ( .IN1(n8935), .IN2(CRC_OUT_8_22), .Q(n13528) );
  AND3X1 U13907 ( .IN1(n13530), .IN2(n13531), .IN3(n9525), .Q(WX2601) );
  OR2X1 U13908 ( .IN1(DFF_373_n1), .IN2(WX2148), .Q(n13531) );
  OR2X1 U13909 ( .IN1(n8936), .IN2(CRC_OUT_8_21), .Q(n13530) );
  AND3X1 U13910 ( .IN1(n13532), .IN2(n13533), .IN3(n9525), .Q(WX2599) );
  OR2X1 U13911 ( .IN1(DFF_372_n1), .IN2(WX2150), .Q(n13533) );
  OR2X1 U13912 ( .IN1(n8937), .IN2(CRC_OUT_8_20), .Q(n13532) );
  AND3X1 U13913 ( .IN1(n13534), .IN2(n13535), .IN3(n9525), .Q(WX2597) );
  OR2X1 U13914 ( .IN1(DFF_371_n1), .IN2(WX2152), .Q(n13535) );
  OR2X1 U13915 ( .IN1(n8938), .IN2(CRC_OUT_8_19), .Q(n13534) );
  AND3X1 U13916 ( .IN1(n13536), .IN2(n13537), .IN3(n9525), .Q(WX2595) );
  OR2X1 U13917 ( .IN1(DFF_370_n1), .IN2(WX2154), .Q(n13537) );
  OR2X1 U13918 ( .IN1(n8939), .IN2(CRC_OUT_8_18), .Q(n13536) );
  AND3X1 U13919 ( .IN1(n13538), .IN2(n13539), .IN3(n9525), .Q(WX2593) );
  OR2X1 U13920 ( .IN1(DFF_369_n1), .IN2(WX2156), .Q(n13539) );
  OR2X1 U13921 ( .IN1(n8940), .IN2(CRC_OUT_8_17), .Q(n13538) );
  AND3X1 U13922 ( .IN1(n13540), .IN2(n13541), .IN3(n9525), .Q(WX2591) );
  OR2X1 U13923 ( .IN1(DFF_368_n1), .IN2(WX2158), .Q(n13541) );
  OR2X1 U13924 ( .IN1(n8941), .IN2(CRC_OUT_8_16), .Q(n13540) );
  AND2X1 U13925 ( .IN1(n13542), .IN2(n9496), .Q(WX2589) );
  OR2X1 U13926 ( .IN1(n13543), .IN2(n13544), .Q(n13542) );
  AND2X1 U13927 ( .IN1(n13545), .IN2(CRC_OUT_8_15), .Q(n13544) );
  AND2X1 U13928 ( .IN1(DFF_367_n1), .IN2(n13546), .Q(n13543) );
  INVX0 U13929 ( .INP(n13545), .ZN(n13546) );
  OR2X1 U13930 ( .IN1(n13547), .IN2(n13548), .Q(n13545) );
  AND2X1 U13931 ( .IN1(DFF_383_n1), .IN2(WX2160), .Q(n13548) );
  AND2X1 U13932 ( .IN1(n8731), .IN2(CRC_OUT_8_31), .Q(n13547) );
  AND3X1 U13933 ( .IN1(n13549), .IN2(n13550), .IN3(n9525), .Q(WX2587) );
  OR2X1 U13934 ( .IN1(DFF_366_n1), .IN2(WX2162), .Q(n13550) );
  OR2X1 U13935 ( .IN1(n8942), .IN2(CRC_OUT_8_14), .Q(n13549) );
  AND3X1 U13936 ( .IN1(n13551), .IN2(n13552), .IN3(n9525), .Q(WX2585) );
  OR2X1 U13937 ( .IN1(DFF_365_n1), .IN2(WX2164), .Q(n13552) );
  OR2X1 U13938 ( .IN1(n8943), .IN2(CRC_OUT_8_13), .Q(n13551) );
  AND3X1 U13939 ( .IN1(n13553), .IN2(n13554), .IN3(n9525), .Q(WX2583) );
  OR2X1 U13940 ( .IN1(DFF_364_n1), .IN2(WX2166), .Q(n13554) );
  OR2X1 U13941 ( .IN1(n8944), .IN2(CRC_OUT_8_12), .Q(n13553) );
  AND3X1 U13942 ( .IN1(n13555), .IN2(n13556), .IN3(n9524), .Q(WX2581) );
  OR2X1 U13943 ( .IN1(DFF_363_n1), .IN2(WX2168), .Q(n13556) );
  OR2X1 U13944 ( .IN1(n8945), .IN2(CRC_OUT_8_11), .Q(n13555) );
  AND2X1 U13945 ( .IN1(n13557), .IN2(n9496), .Q(WX2579) );
  OR2X1 U13946 ( .IN1(n13558), .IN2(n13559), .Q(n13557) );
  AND2X1 U13947 ( .IN1(n13560), .IN2(CRC_OUT_8_10), .Q(n13559) );
  AND2X1 U13948 ( .IN1(DFF_362_n1), .IN2(n13561), .Q(n13558) );
  INVX0 U13949 ( .INP(n13560), .ZN(n13561) );
  OR2X1 U13950 ( .IN1(n13562), .IN2(n13563), .Q(n13560) );
  AND2X1 U13951 ( .IN1(DFF_383_n1), .IN2(WX2170), .Q(n13563) );
  AND2X1 U13952 ( .IN1(n8732), .IN2(CRC_OUT_8_31), .Q(n13562) );
  AND2X1 U13953 ( .IN1(n13564), .IN2(n9496), .Q(WX2577) );
  OR2X1 U13954 ( .IN1(n13565), .IN2(n13566), .Q(n13564) );
  AND2X1 U13955 ( .IN1(DFF_361_n1), .IN2(n9101), .Q(n13566) );
  AND2X1 U13956 ( .IN1(test_so19), .IN2(CRC_OUT_8_9), .Q(n13565) );
  AND3X1 U13957 ( .IN1(n13567), .IN2(n13568), .IN3(n9524), .Q(WX2575) );
  OR2X1 U13958 ( .IN1(DFF_360_n1), .IN2(WX2174), .Q(n13568) );
  OR2X1 U13959 ( .IN1(n8946), .IN2(CRC_OUT_8_8), .Q(n13567) );
  AND2X1 U13960 ( .IN1(n13569), .IN2(n9497), .Q(WX2573) );
  OR2X1 U13961 ( .IN1(n13570), .IN2(n13571), .Q(n13569) );
  AND2X1 U13962 ( .IN1(n8947), .IN2(n9160), .Q(n13571) );
  AND2X1 U13963 ( .IN1(test_so20), .IN2(WX2176), .Q(n13570) );
  AND3X1 U13964 ( .IN1(n13572), .IN2(n13573), .IN3(n9524), .Q(WX2571) );
  OR2X1 U13965 ( .IN1(DFF_358_n1), .IN2(WX2178), .Q(n13573) );
  OR2X1 U13966 ( .IN1(n8948), .IN2(CRC_OUT_8_6), .Q(n13572) );
  AND3X1 U13967 ( .IN1(n13574), .IN2(n13575), .IN3(n9524), .Q(WX2569) );
  OR2X1 U13968 ( .IN1(DFF_357_n1), .IN2(WX2180), .Q(n13575) );
  OR2X1 U13969 ( .IN1(n8949), .IN2(CRC_OUT_8_5), .Q(n13574) );
  AND3X1 U13970 ( .IN1(n13576), .IN2(n13577), .IN3(n9524), .Q(WX2567) );
  OR2X1 U13971 ( .IN1(DFF_356_n1), .IN2(WX2182), .Q(n13577) );
  OR2X1 U13972 ( .IN1(n8950), .IN2(CRC_OUT_8_4), .Q(n13576) );
  AND2X1 U13973 ( .IN1(n13578), .IN2(n9497), .Q(WX2565) );
  OR2X1 U13974 ( .IN1(n13579), .IN2(n13580), .Q(n13578) );
  AND2X1 U13975 ( .IN1(n13581), .IN2(CRC_OUT_8_3), .Q(n13580) );
  AND2X1 U13976 ( .IN1(DFF_355_n1), .IN2(n13582), .Q(n13579) );
  INVX0 U13977 ( .INP(n13581), .ZN(n13582) );
  OR2X1 U13978 ( .IN1(n13583), .IN2(n13584), .Q(n13581) );
  AND2X1 U13979 ( .IN1(DFF_383_n1), .IN2(WX2184), .Q(n13584) );
  AND2X1 U13980 ( .IN1(n8733), .IN2(CRC_OUT_8_31), .Q(n13583) );
  AND3X1 U13981 ( .IN1(n13585), .IN2(n13586), .IN3(n9524), .Q(WX2563) );
  OR2X1 U13982 ( .IN1(DFF_354_n1), .IN2(WX2186), .Q(n13586) );
  OR2X1 U13983 ( .IN1(n8951), .IN2(CRC_OUT_8_2), .Q(n13585) );
  AND3X1 U13984 ( .IN1(n13587), .IN2(n13588), .IN3(n9524), .Q(WX2561) );
  OR2X1 U13985 ( .IN1(DFF_353_n1), .IN2(WX2188), .Q(n13588) );
  OR2X1 U13986 ( .IN1(n8952), .IN2(CRC_OUT_8_1), .Q(n13587) );
  AND3X1 U13987 ( .IN1(n13589), .IN2(n13590), .IN3(n9524), .Q(WX2559) );
  OR2X1 U13988 ( .IN1(DFF_352_n1), .IN2(WX2190), .Q(n13590) );
  OR2X1 U13989 ( .IN1(n8953), .IN2(CRC_OUT_8_0), .Q(n13589) );
  AND3X1 U13990 ( .IN1(n13591), .IN2(n13592), .IN3(n9524), .Q(WX2557) );
  OR2X1 U13991 ( .IN1(DFF_383_n1), .IN2(WX2192), .Q(n13592) );
  OR2X1 U13992 ( .IN1(n8741), .IN2(CRC_OUT_8_31), .Q(n13591) );
  AND2X1 U13993 ( .IN1(n9508), .IN2(n8653), .Q(WX2031) );
  AND2X1 U13994 ( .IN1(n9507), .IN2(n8654), .Q(WX2029) );
  AND2X1 U13995 ( .IN1(n9507), .IN2(n8655), .Q(WX2027) );
  AND2X1 U13996 ( .IN1(n9507), .IN2(n8656), .Q(WX2025) );
  AND2X1 U13997 ( .IN1(n9507), .IN2(n8657), .Q(WX2023) );
  AND2X1 U13998 ( .IN1(n9507), .IN2(n8658), .Q(WX2021) );
  AND2X1 U13999 ( .IN1(test_so13), .IN2(n9495), .Q(WX2019) );
  AND2X1 U14000 ( .IN1(n9508), .IN2(n8661), .Q(WX2017) );
  AND2X1 U14001 ( .IN1(n9499), .IN2(n8662), .Q(WX2015) );
  AND2X1 U14002 ( .IN1(n9507), .IN2(n8663), .Q(WX2013) );
  AND2X1 U14003 ( .IN1(n9508), .IN2(n8664), .Q(WX2011) );
  AND2X1 U14004 ( .IN1(n9508), .IN2(n8665), .Q(WX2009) );
  AND2X1 U14005 ( .IN1(n9509), .IN2(n8666), .Q(WX2007) );
  AND2X1 U14006 ( .IN1(n9509), .IN2(n8667), .Q(WX2005) );
  AND2X1 U14007 ( .IN1(n9509), .IN2(n8668), .Q(WX2003) );
  AND2X1 U14008 ( .IN1(n9509), .IN2(n8669), .Q(WX2001) );
  OR4X1 U14009 ( .IN1(n13593), .IN2(n13594), .IN3(n13595), .IN4(n13596), .Q(
        WX1999) );
  AND2X1 U14010 ( .IN1(n9268), .IN2(n12939), .Q(n13596) );
  OR2X1 U14011 ( .IN1(n13597), .IN2(n13598), .Q(n12939) );
  INVX0 U14012 ( .INP(n13599), .ZN(n13598) );
  OR2X1 U14013 ( .IN1(n13600), .IN2(n13601), .Q(n13599) );
  AND2X1 U14014 ( .IN1(n13601), .IN2(n13600), .Q(n13597) );
  AND2X1 U14015 ( .IN1(n13602), .IN2(n13603), .Q(n13600) );
  OR2X1 U14016 ( .IN1(WX3357), .IN2(n8476), .Q(n13603) );
  INVX0 U14017 ( .INP(n13604), .ZN(n13602) );
  AND2X1 U14018 ( .IN1(n8476), .IN2(WX3357), .Q(n13604) );
  OR2X1 U14019 ( .IN1(n13605), .IN2(n13606), .Q(n13601) );
  AND2X1 U14020 ( .IN1(n8477), .IN2(WX3485), .Q(n13606) );
  AND2X1 U14021 ( .IN1(n8740), .IN2(WX3421), .Q(n13605) );
  AND2X1 U14022 ( .IN1(n11356), .IN2(n9177), .Q(n13595) );
  AND2X1 U14023 ( .IN1(n13607), .IN2(n13608), .Q(n11356) );
  INVX0 U14024 ( .INP(n13609), .ZN(n13608) );
  AND2X1 U14025 ( .IN1(n13610), .IN2(n13611), .Q(n13609) );
  OR2X1 U14026 ( .IN1(n13611), .IN2(n13610), .Q(n13607) );
  OR2X1 U14027 ( .IN1(n13612), .IN2(n13613), .Q(n13610) );
  INVX0 U14028 ( .INP(n13614), .ZN(n13613) );
  OR2X1 U14029 ( .IN1(WX2000), .IN2(n8596), .Q(n13614) );
  AND2X1 U14030 ( .IN1(n8596), .IN2(WX2000), .Q(n13612) );
  AND2X1 U14031 ( .IN1(n13615), .IN2(n13616), .Q(n13611) );
  OR2X1 U14032 ( .IN1(WX2192), .IN2(test_so16), .Q(n13616) );
  OR2X1 U14033 ( .IN1(n9134), .IN2(n8741), .Q(n13615) );
  AND2X1 U14034 ( .IN1(n9233), .IN2(CRC_OUT_8_0), .Q(n13594) );
  AND2X1 U14035 ( .IN1(n297), .IN2(n9207), .Q(n13593) );
  INVX0 U14036 ( .INP(n13617), .ZN(n297) );
  OR2X1 U14037 ( .IN1(n9562), .IN2(n4003), .Q(n13617) );
  OR4X1 U14038 ( .IN1(n13618), .IN2(n13619), .IN3(n13620), .IN4(n13621), .Q(
        WX1997) );
  AND2X1 U14039 ( .IN1(n9268), .IN2(n12955), .Q(n13621) );
  OR2X1 U14040 ( .IN1(n13622), .IN2(n13623), .Q(n12955) );
  INVX0 U14041 ( .INP(n13624), .ZN(n13623) );
  OR2X1 U14042 ( .IN1(n13625), .IN2(n13626), .Q(n13624) );
  AND2X1 U14043 ( .IN1(n13626), .IN2(n13625), .Q(n13622) );
  AND2X1 U14044 ( .IN1(n13627), .IN2(n13628), .Q(n13625) );
  OR2X1 U14045 ( .IN1(WX3355), .IN2(n8478), .Q(n13628) );
  INVX0 U14046 ( .INP(n13629), .ZN(n13627) );
  AND2X1 U14047 ( .IN1(n8478), .IN2(WX3355), .Q(n13629) );
  OR2X1 U14048 ( .IN1(n13630), .IN2(n13631), .Q(n13626) );
  AND2X1 U14049 ( .IN1(n8485), .IN2(WX3483), .Q(n13631) );
  AND2X1 U14050 ( .IN1(n8927), .IN2(WX3419), .Q(n13630) );
  AND2X1 U14051 ( .IN1(n9189), .IN2(n11362), .Q(n13620) );
  OR2X1 U14052 ( .IN1(n13632), .IN2(n13633), .Q(n11362) );
  INVX0 U14053 ( .INP(n13634), .ZN(n13633) );
  OR2X1 U14054 ( .IN1(n13635), .IN2(n13636), .Q(n13634) );
  AND2X1 U14055 ( .IN1(n13636), .IN2(n13635), .Q(n13632) );
  AND2X1 U14056 ( .IN1(n13637), .IN2(n13638), .Q(n13635) );
  OR2X1 U14057 ( .IN1(WX2062), .IN2(n8614), .Q(n13638) );
  INVX0 U14058 ( .INP(n13639), .ZN(n13637) );
  AND2X1 U14059 ( .IN1(n8614), .IN2(WX2062), .Q(n13639) );
  OR2X1 U14060 ( .IN1(n13640), .IN2(n13641), .Q(n13636) );
  AND2X1 U14061 ( .IN1(n8615), .IN2(WX2190), .Q(n13641) );
  AND2X1 U14062 ( .IN1(n8953), .IN2(WX2126), .Q(n13640) );
  AND2X1 U14063 ( .IN1(n9234), .IN2(CRC_OUT_8_1), .Q(n13619) );
  AND2X1 U14064 ( .IN1(n296), .IN2(n9207), .Q(n13618) );
  INVX0 U14065 ( .INP(n13642), .ZN(n296) );
  OR2X1 U14066 ( .IN1(n9562), .IN2(n4004), .Q(n13642) );
  OR4X1 U14067 ( .IN1(n13643), .IN2(n13644), .IN3(n13645), .IN4(n13646), .Q(
        WX1995) );
  AND2X1 U14068 ( .IN1(n9268), .IN2(n12971), .Q(n13646) );
  OR2X1 U14069 ( .IN1(n13647), .IN2(n13648), .Q(n12971) );
  INVX0 U14070 ( .INP(n13649), .ZN(n13648) );
  OR2X1 U14071 ( .IN1(n13650), .IN2(n13651), .Q(n13649) );
  AND2X1 U14072 ( .IN1(n13651), .IN2(n13650), .Q(n13647) );
  AND2X1 U14073 ( .IN1(n13652), .IN2(n13653), .Q(n13650) );
  OR2X1 U14074 ( .IN1(WX3353), .IN2(n8486), .Q(n13653) );
  INVX0 U14075 ( .INP(n13654), .ZN(n13652) );
  AND2X1 U14076 ( .IN1(n8486), .IN2(WX3353), .Q(n13654) );
  OR2X1 U14077 ( .IN1(n13655), .IN2(n13656), .Q(n13651) );
  AND2X1 U14078 ( .IN1(n8503), .IN2(WX3481), .Q(n13656) );
  AND2X1 U14079 ( .IN1(n8926), .IN2(WX3417), .Q(n13655) );
  AND2X1 U14080 ( .IN1(n9189), .IN2(n11368), .Q(n13645) );
  OR2X1 U14081 ( .IN1(n13657), .IN2(n13658), .Q(n11368) );
  INVX0 U14082 ( .INP(n13659), .ZN(n13658) );
  OR2X1 U14083 ( .IN1(n13660), .IN2(n13661), .Q(n13659) );
  AND2X1 U14084 ( .IN1(n13661), .IN2(n13660), .Q(n13657) );
  AND2X1 U14085 ( .IN1(n13662), .IN2(n13663), .Q(n13660) );
  OR2X1 U14086 ( .IN1(WX2060), .IN2(n8633), .Q(n13663) );
  INVX0 U14087 ( .INP(n13664), .ZN(n13662) );
  AND2X1 U14088 ( .IN1(n8633), .IN2(WX2060), .Q(n13664) );
  OR2X1 U14089 ( .IN1(n13665), .IN2(n13666), .Q(n13661) );
  AND2X1 U14090 ( .IN1(n8634), .IN2(WX2188), .Q(n13666) );
  AND2X1 U14091 ( .IN1(n8952), .IN2(WX2124), .Q(n13665) );
  AND2X1 U14092 ( .IN1(n9234), .IN2(CRC_OUT_8_2), .Q(n13644) );
  AND2X1 U14093 ( .IN1(n295), .IN2(n9207), .Q(n13643) );
  INVX0 U14094 ( .INP(n13667), .ZN(n295) );
  OR2X1 U14095 ( .IN1(n9561), .IN2(n4005), .Q(n13667) );
  OR4X1 U14096 ( .IN1(n13668), .IN2(n13669), .IN3(n13670), .IN4(n13671), .Q(
        WX1993) );
  AND2X1 U14097 ( .IN1(n9268), .IN2(n12987), .Q(n13671) );
  OR2X1 U14098 ( .IN1(n13672), .IN2(n13673), .Q(n12987) );
  INVX0 U14099 ( .INP(n13674), .ZN(n13673) );
  OR2X1 U14100 ( .IN1(n13675), .IN2(n13676), .Q(n13674) );
  AND2X1 U14101 ( .IN1(n13676), .IN2(n13675), .Q(n13672) );
  AND2X1 U14102 ( .IN1(n13677), .IN2(n13678), .Q(n13675) );
  OR2X1 U14103 ( .IN1(WX3351), .IN2(n8504), .Q(n13678) );
  INVX0 U14104 ( .INP(n13679), .ZN(n13677) );
  AND2X1 U14105 ( .IN1(n8504), .IN2(WX3351), .Q(n13679) );
  OR2X1 U14106 ( .IN1(n13680), .IN2(n13681), .Q(n13676) );
  AND2X1 U14107 ( .IN1(n8521), .IN2(WX3479), .Q(n13681) );
  AND2X1 U14108 ( .IN1(n8925), .IN2(WX3415), .Q(n13680) );
  AND2X1 U14109 ( .IN1(n9189), .IN2(n11374), .Q(n13670) );
  OR2X1 U14110 ( .IN1(n13682), .IN2(n13683), .Q(n11374) );
  INVX0 U14111 ( .INP(n13684), .ZN(n13683) );
  OR2X1 U14112 ( .IN1(n13685), .IN2(n13686), .Q(n13684) );
  AND2X1 U14113 ( .IN1(n13686), .IN2(n13685), .Q(n13682) );
  AND2X1 U14114 ( .IN1(n13687), .IN2(n13688), .Q(n13685) );
  OR2X1 U14115 ( .IN1(WX2058), .IN2(n8645), .Q(n13688) );
  INVX0 U14116 ( .INP(n13689), .ZN(n13687) );
  AND2X1 U14117 ( .IN1(n8645), .IN2(WX2058), .Q(n13689) );
  OR2X1 U14118 ( .IN1(n13690), .IN2(n13691), .Q(n13686) );
  AND2X1 U14119 ( .IN1(n8646), .IN2(WX2186), .Q(n13691) );
  AND2X1 U14120 ( .IN1(n8951), .IN2(WX2122), .Q(n13690) );
  AND2X1 U14121 ( .IN1(n9234), .IN2(CRC_OUT_8_3), .Q(n13669) );
  AND2X1 U14122 ( .IN1(n294), .IN2(n9207), .Q(n13668) );
  INVX0 U14123 ( .INP(n13692), .ZN(n294) );
  OR2X1 U14124 ( .IN1(n9561), .IN2(n4006), .Q(n13692) );
  OR4X1 U14125 ( .IN1(n13693), .IN2(n13694), .IN3(n13695), .IN4(n13696), .Q(
        WX1991) );
  AND2X1 U14126 ( .IN1(n9268), .IN2(n13003), .Q(n13696) );
  OR2X1 U14127 ( .IN1(n13697), .IN2(n13698), .Q(n13003) );
  INVX0 U14128 ( .INP(n13699), .ZN(n13698) );
  OR2X1 U14129 ( .IN1(n13700), .IN2(n13701), .Q(n13699) );
  AND2X1 U14130 ( .IN1(n13701), .IN2(n13700), .Q(n13697) );
  AND2X1 U14131 ( .IN1(n13702), .IN2(n13703), .Q(n13700) );
  OR2X1 U14132 ( .IN1(WX3349), .IN2(n8522), .Q(n13703) );
  INVX0 U14133 ( .INP(n13704), .ZN(n13702) );
  AND2X1 U14134 ( .IN1(n8522), .IN2(WX3349), .Q(n13704) );
  OR2X1 U14135 ( .IN1(n13705), .IN2(n13706), .Q(n13701) );
  AND2X1 U14136 ( .IN1(n8529), .IN2(WX3477), .Q(n13706) );
  AND2X1 U14137 ( .IN1(n8730), .IN2(WX3413), .Q(n13705) );
  AND2X1 U14138 ( .IN1(n11380), .IN2(n9177), .Q(n13695) );
  AND2X1 U14139 ( .IN1(n13707), .IN2(n13708), .Q(n11380) );
  INVX0 U14140 ( .INP(n13709), .ZN(n13708) );
  AND2X1 U14141 ( .IN1(n13710), .IN2(n13711), .Q(n13709) );
  OR2X1 U14142 ( .IN1(n13711), .IN2(n13710), .Q(n13707) );
  OR2X1 U14143 ( .IN1(n13712), .IN2(n13713), .Q(n13710) );
  INVX0 U14144 ( .INP(n13714), .ZN(n13713) );
  OR2X1 U14145 ( .IN1(WX2056), .IN2(n8647), .Q(n13714) );
  AND2X1 U14146 ( .IN1(n8647), .IN2(WX2056), .Q(n13712) );
  AND2X1 U14147 ( .IN1(n13715), .IN2(n13716), .Q(n13711) );
  OR2X1 U14148 ( .IN1(WX2184), .IN2(test_so14), .Q(n13716) );
  OR2X1 U14149 ( .IN1(n9135), .IN2(n8733), .Q(n13715) );
  AND2X1 U14150 ( .IN1(n9234), .IN2(CRC_OUT_8_4), .Q(n13694) );
  AND2X1 U14151 ( .IN1(n293), .IN2(n9207), .Q(n13693) );
  INVX0 U14152 ( .INP(n13717), .ZN(n293) );
  OR2X1 U14153 ( .IN1(n9561), .IN2(n4007), .Q(n13717) );
  OR4X1 U14154 ( .IN1(n13718), .IN2(n13719), .IN3(n13720), .IN4(n13721), .Q(
        WX1989) );
  AND2X1 U14155 ( .IN1(n9268), .IN2(n13019), .Q(n13721) );
  OR2X1 U14156 ( .IN1(n13722), .IN2(n13723), .Q(n13019) );
  INVX0 U14157 ( .INP(n13724), .ZN(n13723) );
  OR2X1 U14158 ( .IN1(n13725), .IN2(n13726), .Q(n13724) );
  AND2X1 U14159 ( .IN1(n13726), .IN2(n13725), .Q(n13722) );
  AND2X1 U14160 ( .IN1(n13727), .IN2(n13728), .Q(n13725) );
  OR2X1 U14161 ( .IN1(WX3347), .IN2(n8530), .Q(n13728) );
  INVX0 U14162 ( .INP(n13729), .ZN(n13727) );
  AND2X1 U14163 ( .IN1(n8530), .IN2(WX3347), .Q(n13729) );
  OR2X1 U14164 ( .IN1(n13730), .IN2(n13731), .Q(n13726) );
  AND2X1 U14165 ( .IN1(n8531), .IN2(WX3475), .Q(n13731) );
  AND2X1 U14166 ( .IN1(n8924), .IN2(WX3411), .Q(n13730) );
  AND2X1 U14167 ( .IN1(n9189), .IN2(n11386), .Q(n13720) );
  OR2X1 U14168 ( .IN1(n13732), .IN2(n13733), .Q(n11386) );
  INVX0 U14169 ( .INP(n13734), .ZN(n13733) );
  OR2X1 U14170 ( .IN1(n13735), .IN2(n13736), .Q(n13734) );
  AND2X1 U14171 ( .IN1(n13736), .IN2(n13735), .Q(n13732) );
  AND2X1 U14172 ( .IN1(n13737), .IN2(n13738), .Q(n13735) );
  OR2X1 U14173 ( .IN1(WX2054), .IN2(n8648), .Q(n13738) );
  INVX0 U14174 ( .INP(n13739), .ZN(n13737) );
  AND2X1 U14175 ( .IN1(n8648), .IN2(WX2054), .Q(n13739) );
  OR2X1 U14176 ( .IN1(n13740), .IN2(n13741), .Q(n13736) );
  AND2X1 U14177 ( .IN1(n8649), .IN2(WX2182), .Q(n13741) );
  AND2X1 U14178 ( .IN1(n8950), .IN2(WX2118), .Q(n13740) );
  AND2X1 U14179 ( .IN1(n9234), .IN2(CRC_OUT_8_5), .Q(n13719) );
  AND2X1 U14180 ( .IN1(n292), .IN2(n9208), .Q(n13718) );
  INVX0 U14181 ( .INP(n13742), .ZN(n292) );
  OR2X1 U14182 ( .IN1(n9561), .IN2(n4008), .Q(n13742) );
  OR4X1 U14183 ( .IN1(n13743), .IN2(n13744), .IN3(n13745), .IN4(n13746), .Q(
        WX1987) );
  AND2X1 U14184 ( .IN1(n13035), .IN2(n9260), .Q(n13746) );
  AND2X1 U14185 ( .IN1(n13747), .IN2(n13748), .Q(n13035) );
  INVX0 U14186 ( .INP(n13749), .ZN(n13748) );
  AND2X1 U14187 ( .IN1(n13750), .IN2(n13751), .Q(n13749) );
  OR2X1 U14188 ( .IN1(n13751), .IN2(n13750), .Q(n13747) );
  OR2X1 U14189 ( .IN1(n13752), .IN2(n13753), .Q(n13750) );
  INVX0 U14190 ( .INP(n13754), .ZN(n13753) );
  OR2X1 U14191 ( .IN1(WX3345), .IN2(n8532), .Q(n13754) );
  AND2X1 U14192 ( .IN1(n8532), .IN2(WX3345), .Q(n13752) );
  AND2X1 U14193 ( .IN1(n13755), .IN2(n13756), .Q(n13751) );
  OR2X1 U14194 ( .IN1(WX3409), .IN2(test_so30), .Q(n13756) );
  OR2X1 U14195 ( .IN1(n9100), .IN2(n8533), .Q(n13755) );
  AND2X1 U14196 ( .IN1(n9189), .IN2(n11392), .Q(n13745) );
  OR2X1 U14197 ( .IN1(n13757), .IN2(n13758), .Q(n11392) );
  INVX0 U14198 ( .INP(n13759), .ZN(n13758) );
  OR2X1 U14199 ( .IN1(n13760), .IN2(n13761), .Q(n13759) );
  AND2X1 U14200 ( .IN1(n13761), .IN2(n13760), .Q(n13757) );
  AND2X1 U14201 ( .IN1(n13762), .IN2(n13763), .Q(n13760) );
  OR2X1 U14202 ( .IN1(WX2052), .IN2(n8650), .Q(n13763) );
  INVX0 U14203 ( .INP(n13764), .ZN(n13762) );
  AND2X1 U14204 ( .IN1(n8650), .IN2(WX2052), .Q(n13764) );
  OR2X1 U14205 ( .IN1(n13765), .IN2(n13766), .Q(n13761) );
  AND2X1 U14206 ( .IN1(n8651), .IN2(WX2180), .Q(n13766) );
  AND2X1 U14207 ( .IN1(n8949), .IN2(WX2116), .Q(n13765) );
  AND2X1 U14208 ( .IN1(n9234), .IN2(CRC_OUT_8_6), .Q(n13744) );
  AND2X1 U14209 ( .IN1(n291), .IN2(n9208), .Q(n13743) );
  INVX0 U14210 ( .INP(n13767), .ZN(n291) );
  OR2X1 U14211 ( .IN1(n9561), .IN2(n4009), .Q(n13767) );
  OR4X1 U14212 ( .IN1(n13768), .IN2(n13769), .IN3(n13770), .IN4(n13771), .Q(
        WX1985) );
  AND2X1 U14213 ( .IN1(n9268), .IN2(n13051), .Q(n13771) );
  OR2X1 U14214 ( .IN1(n13772), .IN2(n13773), .Q(n13051) );
  INVX0 U14215 ( .INP(n13774), .ZN(n13773) );
  OR2X1 U14216 ( .IN1(n13775), .IN2(n13776), .Q(n13774) );
  AND2X1 U14217 ( .IN1(n13776), .IN2(n13775), .Q(n13772) );
  AND2X1 U14218 ( .IN1(n13777), .IN2(n13778), .Q(n13775) );
  OR2X1 U14219 ( .IN1(WX3343), .IN2(n8534), .Q(n13778) );
  INVX0 U14220 ( .INP(n13779), .ZN(n13777) );
  AND2X1 U14221 ( .IN1(n8534), .IN2(WX3343), .Q(n13779) );
  OR2X1 U14222 ( .IN1(n13780), .IN2(n13781), .Q(n13776) );
  AND2X1 U14223 ( .IN1(n8535), .IN2(WX3471), .Q(n13781) );
  AND2X1 U14224 ( .IN1(n8923), .IN2(WX3407), .Q(n13780) );
  AND2X1 U14225 ( .IN1(n9189), .IN2(n11398), .Q(n13770) );
  OR2X1 U14226 ( .IN1(n13782), .IN2(n13783), .Q(n11398) );
  INVX0 U14227 ( .INP(n13784), .ZN(n13783) );
  OR2X1 U14228 ( .IN1(n13785), .IN2(n13786), .Q(n13784) );
  AND2X1 U14229 ( .IN1(n13786), .IN2(n13785), .Q(n13782) );
  AND2X1 U14230 ( .IN1(n13787), .IN2(n13788), .Q(n13785) );
  OR2X1 U14231 ( .IN1(WX2050), .IN2(n8652), .Q(n13788) );
  INVX0 U14232 ( .INP(n13789), .ZN(n13787) );
  AND2X1 U14233 ( .IN1(n8652), .IN2(WX2050), .Q(n13789) );
  OR2X1 U14234 ( .IN1(n13790), .IN2(n13791), .Q(n13786) );
  AND2X1 U14235 ( .IN1(n8659), .IN2(WX2178), .Q(n13791) );
  AND2X1 U14236 ( .IN1(n8948), .IN2(WX2114), .Q(n13790) );
  AND2X1 U14237 ( .IN1(test_so20), .IN2(n9227), .Q(n13769) );
  AND2X1 U14238 ( .IN1(n290), .IN2(n9208), .Q(n13768) );
  INVX0 U14239 ( .INP(n13792), .ZN(n290) );
  OR2X1 U14240 ( .IN1(n9561), .IN2(n4010), .Q(n13792) );
  OR4X1 U14241 ( .IN1(n13793), .IN2(n13794), .IN3(n13795), .IN4(n13796), .Q(
        WX1983) );
  AND2X1 U14242 ( .IN1(n13067), .IN2(n9260), .Q(n13796) );
  AND2X1 U14243 ( .IN1(n13797), .IN2(n13798), .Q(n13067) );
  INVX0 U14244 ( .INP(n13799), .ZN(n13798) );
  AND2X1 U14245 ( .IN1(n13800), .IN2(n13801), .Q(n13799) );
  OR2X1 U14246 ( .IN1(n13801), .IN2(n13800), .Q(n13797) );
  OR2X1 U14247 ( .IN1(n13802), .IN2(n13803), .Q(n13800) );
  INVX0 U14248 ( .INP(n13804), .ZN(n13803) );
  OR2X1 U14249 ( .IN1(WX3341), .IN2(n8536), .Q(n13804) );
  AND2X1 U14250 ( .IN1(n8536), .IN2(WX3341), .Q(n13802) );
  AND2X1 U14251 ( .IN1(n13805), .IN2(n13806), .Q(n13801) );
  OR2X1 U14252 ( .IN1(WX3469), .IN2(test_so28), .Q(n13806) );
  OR2X1 U14253 ( .IN1(n9136), .IN2(n8922), .Q(n13805) );
  AND2X1 U14254 ( .IN1(n9189), .IN2(n11404), .Q(n13795) );
  OR2X1 U14255 ( .IN1(n13807), .IN2(n13808), .Q(n11404) );
  INVX0 U14256 ( .INP(n13809), .ZN(n13808) );
  OR2X1 U14257 ( .IN1(n13810), .IN2(n13811), .Q(n13809) );
  AND2X1 U14258 ( .IN1(n13811), .IN2(n13810), .Q(n13807) );
  AND2X1 U14259 ( .IN1(n13812), .IN2(n13813), .Q(n13810) );
  OR2X1 U14260 ( .IN1(WX2048), .IN2(n8660), .Q(n13813) );
  INVX0 U14261 ( .INP(n13814), .ZN(n13812) );
  AND2X1 U14262 ( .IN1(n8660), .IN2(WX2048), .Q(n13814) );
  OR2X1 U14263 ( .IN1(n13815), .IN2(n13816), .Q(n13811) );
  AND2X1 U14264 ( .IN1(n8678), .IN2(WX2176), .Q(n13816) );
  AND2X1 U14265 ( .IN1(n8947), .IN2(WX2112), .Q(n13815) );
  AND2X1 U14266 ( .IN1(n9234), .IN2(CRC_OUT_8_8), .Q(n13794) );
  AND2X1 U14267 ( .IN1(n289), .IN2(n9208), .Q(n13793) );
  INVX0 U14268 ( .INP(n13817), .ZN(n289) );
  OR2X1 U14269 ( .IN1(n9561), .IN2(n4011), .Q(n13817) );
  OR4X1 U14270 ( .IN1(n13818), .IN2(n13819), .IN3(n13820), .IN4(n13821), .Q(
        WX1981) );
  AND2X1 U14271 ( .IN1(n9268), .IN2(n13083), .Q(n13821) );
  OR2X1 U14272 ( .IN1(n13822), .IN2(n13823), .Q(n13083) );
  INVX0 U14273 ( .INP(n13824), .ZN(n13823) );
  OR2X1 U14274 ( .IN1(n13825), .IN2(n13826), .Q(n13824) );
  AND2X1 U14275 ( .IN1(n13826), .IN2(n13825), .Q(n13822) );
  AND2X1 U14276 ( .IN1(n13827), .IN2(n13828), .Q(n13825) );
  OR2X1 U14277 ( .IN1(WX3339), .IN2(n8538), .Q(n13828) );
  INVX0 U14278 ( .INP(n13829), .ZN(n13827) );
  AND2X1 U14279 ( .IN1(n8538), .IN2(WX3339), .Q(n13829) );
  OR2X1 U14280 ( .IN1(n13830), .IN2(n13831), .Q(n13826) );
  AND2X1 U14281 ( .IN1(n8539), .IN2(WX3467), .Q(n13831) );
  AND2X1 U14282 ( .IN1(n8921), .IN2(WX3403), .Q(n13830) );
  AND2X1 U14283 ( .IN1(n9188), .IN2(n11410), .Q(n13820) );
  OR2X1 U14284 ( .IN1(n13832), .IN2(n13833), .Q(n11410) );
  INVX0 U14285 ( .INP(n13834), .ZN(n13833) );
  OR2X1 U14286 ( .IN1(n13835), .IN2(n13836), .Q(n13834) );
  AND2X1 U14287 ( .IN1(n13836), .IN2(n13835), .Q(n13832) );
  AND2X1 U14288 ( .IN1(n13837), .IN2(n13838), .Q(n13835) );
  OR2X1 U14289 ( .IN1(WX2046), .IN2(n8679), .Q(n13838) );
  INVX0 U14290 ( .INP(n13839), .ZN(n13837) );
  AND2X1 U14291 ( .IN1(n8679), .IN2(WX2046), .Q(n13839) );
  OR2X1 U14292 ( .IN1(n13840), .IN2(n13841), .Q(n13836) );
  AND2X1 U14293 ( .IN1(n8697), .IN2(WX2174), .Q(n13841) );
  AND2X1 U14294 ( .IN1(n8946), .IN2(WX2110), .Q(n13840) );
  AND2X1 U14295 ( .IN1(n9234), .IN2(CRC_OUT_8_9), .Q(n13819) );
  AND2X1 U14296 ( .IN1(n288), .IN2(n9208), .Q(n13818) );
  INVX0 U14297 ( .INP(n13842), .ZN(n288) );
  OR2X1 U14298 ( .IN1(n9561), .IN2(n4012), .Q(n13842) );
  OR4X1 U14299 ( .IN1(n13843), .IN2(n13844), .IN3(n13845), .IN4(n13846), .Q(
        WX1979) );
  AND2X1 U14300 ( .IN1(n9268), .IN2(n13099), .Q(n13846) );
  OR2X1 U14301 ( .IN1(n13847), .IN2(n13848), .Q(n13099) );
  INVX0 U14302 ( .INP(n13849), .ZN(n13848) );
  OR2X1 U14303 ( .IN1(n13850), .IN2(n13851), .Q(n13849) );
  AND2X1 U14304 ( .IN1(n13851), .IN2(n13850), .Q(n13847) );
  AND2X1 U14305 ( .IN1(n13852), .IN2(n13853), .Q(n13850) );
  OR2X1 U14306 ( .IN1(WX3337), .IN2(n8556), .Q(n13853) );
  INVX0 U14307 ( .INP(n13854), .ZN(n13852) );
  AND2X1 U14308 ( .IN1(n8556), .IN2(WX3337), .Q(n13854) );
  OR2X1 U14309 ( .IN1(n13855), .IN2(n13856), .Q(n13851) );
  AND2X1 U14310 ( .IN1(n8557), .IN2(WX3465), .Q(n13856) );
  AND2X1 U14311 ( .IN1(n8920), .IN2(WX3401), .Q(n13855) );
  AND2X1 U14312 ( .IN1(n11416), .IN2(n9176), .Q(n13845) );
  AND2X1 U14313 ( .IN1(n13857), .IN2(n13858), .Q(n11416) );
  INVX0 U14314 ( .INP(n13859), .ZN(n13858) );
  AND2X1 U14315 ( .IN1(n13860), .IN2(n13861), .Q(n13859) );
  OR2X1 U14316 ( .IN1(n13861), .IN2(n13860), .Q(n13857) );
  OR2X1 U14317 ( .IN1(n13862), .IN2(n13863), .Q(n13860) );
  INVX0 U14318 ( .INP(n13864), .ZN(n13863) );
  OR2X1 U14319 ( .IN1(WX2044), .IN2(n8698), .Q(n13864) );
  AND2X1 U14320 ( .IN1(n8698), .IN2(WX2044), .Q(n13862) );
  AND2X1 U14321 ( .IN1(n13865), .IN2(n13866), .Q(n13861) );
  OR2X1 U14322 ( .IN1(WX2108), .IN2(test_so19), .Q(n13866) );
  OR2X1 U14323 ( .IN1(n9101), .IN2(n8703), .Q(n13865) );
  AND2X1 U14324 ( .IN1(n9234), .IN2(CRC_OUT_8_10), .Q(n13844) );
  AND2X1 U14325 ( .IN1(n287), .IN2(n9208), .Q(n13843) );
  INVX0 U14326 ( .INP(n13867), .ZN(n287) );
  OR2X1 U14327 ( .IN1(n9561), .IN2(n4013), .Q(n13867) );
  OR4X1 U14328 ( .IN1(n13868), .IN2(n13869), .IN3(n13870), .IN4(n13871), .Q(
        WX1977) );
  AND2X1 U14329 ( .IN1(n9268), .IN2(n13115), .Q(n13871) );
  OR2X1 U14330 ( .IN1(n13872), .IN2(n13873), .Q(n13115) );
  INVX0 U14331 ( .INP(n13874), .ZN(n13873) );
  OR2X1 U14332 ( .IN1(n13875), .IN2(n13876), .Q(n13874) );
  AND2X1 U14333 ( .IN1(n13876), .IN2(n13875), .Q(n13872) );
  AND2X1 U14334 ( .IN1(n13877), .IN2(n13878), .Q(n13875) );
  OR2X1 U14335 ( .IN1(WX3335), .IN2(n8574), .Q(n13878) );
  INVX0 U14336 ( .INP(n13879), .ZN(n13877) );
  AND2X1 U14337 ( .IN1(n8574), .IN2(WX3335), .Q(n13879) );
  OR2X1 U14338 ( .IN1(n13880), .IN2(n13881), .Q(n13876) );
  AND2X1 U14339 ( .IN1(n8575), .IN2(WX3463), .Q(n13881) );
  AND2X1 U14340 ( .IN1(n8729), .IN2(WX3399), .Q(n13880) );
  AND2X1 U14341 ( .IN1(n9188), .IN2(n11422), .Q(n13870) );
  OR2X1 U14342 ( .IN1(n13882), .IN2(n13883), .Q(n11422) );
  INVX0 U14343 ( .INP(n13884), .ZN(n13883) );
  OR2X1 U14344 ( .IN1(n13885), .IN2(n13886), .Q(n13884) );
  AND2X1 U14345 ( .IN1(n13886), .IN2(n13885), .Q(n13882) );
  AND2X1 U14346 ( .IN1(n13887), .IN2(n13888), .Q(n13885) );
  OR2X1 U14347 ( .IN1(WX2042), .IN2(n8704), .Q(n13888) );
  INVX0 U14348 ( .INP(n13889), .ZN(n13887) );
  AND2X1 U14349 ( .IN1(n8704), .IN2(WX2042), .Q(n13889) );
  OR2X1 U14350 ( .IN1(n13890), .IN2(n13891), .Q(n13886) );
  AND2X1 U14351 ( .IN1(n8705), .IN2(WX2170), .Q(n13891) );
  AND2X1 U14352 ( .IN1(n8732), .IN2(WX2106), .Q(n13890) );
  AND2X1 U14353 ( .IN1(n9234), .IN2(CRC_OUT_8_11), .Q(n13869) );
  AND2X1 U14354 ( .IN1(n286), .IN2(n9208), .Q(n13868) );
  INVX0 U14355 ( .INP(n13892), .ZN(n286) );
  OR2X1 U14356 ( .IN1(n9561), .IN2(n4014), .Q(n13892) );
  OR4X1 U14357 ( .IN1(n13893), .IN2(n13894), .IN3(n13895), .IN4(n13896), .Q(
        WX1975) );
  AND2X1 U14358 ( .IN1(n13131), .IN2(n9260), .Q(n13896) );
  AND2X1 U14359 ( .IN1(n13897), .IN2(n13898), .Q(n13131) );
  INVX0 U14360 ( .INP(n13899), .ZN(n13898) );
  AND2X1 U14361 ( .IN1(n13900), .IN2(n13901), .Q(n13899) );
  OR2X1 U14362 ( .IN1(n13901), .IN2(n13900), .Q(n13897) );
  OR2X1 U14363 ( .IN1(n13902), .IN2(n13903), .Q(n13900) );
  INVX0 U14364 ( .INP(n13904), .ZN(n13903) );
  OR2X1 U14365 ( .IN1(WX3269), .IN2(n8588), .Q(n13904) );
  AND2X1 U14366 ( .IN1(n8588), .IN2(WX3269), .Q(n13902) );
  AND2X1 U14367 ( .IN1(n13905), .IN2(n13906), .Q(n13901) );
  OR2X1 U14368 ( .IN1(WX3461), .IN2(test_so26), .Q(n13906) );
  OR2X1 U14369 ( .IN1(n9137), .IN2(n8919), .Q(n13905) );
  AND2X1 U14370 ( .IN1(n9188), .IN2(n11428), .Q(n13895) );
  OR2X1 U14371 ( .IN1(n13907), .IN2(n13908), .Q(n11428) );
  INVX0 U14372 ( .INP(n13909), .ZN(n13908) );
  OR2X1 U14373 ( .IN1(n13910), .IN2(n13911), .Q(n13909) );
  AND2X1 U14374 ( .IN1(n13911), .IN2(n13910), .Q(n13907) );
  AND2X1 U14375 ( .IN1(n13912), .IN2(n13913), .Q(n13910) );
  OR2X1 U14376 ( .IN1(WX2040), .IN2(n8706), .Q(n13913) );
  INVX0 U14377 ( .INP(n13914), .ZN(n13912) );
  AND2X1 U14378 ( .IN1(n8706), .IN2(WX2040), .Q(n13914) );
  OR2X1 U14379 ( .IN1(n13915), .IN2(n13916), .Q(n13911) );
  AND2X1 U14380 ( .IN1(n8707), .IN2(WX2168), .Q(n13916) );
  AND2X1 U14381 ( .IN1(n8945), .IN2(WX2104), .Q(n13915) );
  AND2X1 U14382 ( .IN1(n9234), .IN2(CRC_OUT_8_12), .Q(n13894) );
  AND2X1 U14383 ( .IN1(n285), .IN2(n9208), .Q(n13893) );
  INVX0 U14384 ( .INP(n13917), .ZN(n285) );
  OR2X1 U14385 ( .IN1(n9561), .IN2(n4015), .Q(n13917) );
  OR4X1 U14386 ( .IN1(n13918), .IN2(n13919), .IN3(n13920), .IN4(n13921), .Q(
        WX1973) );
  AND2X1 U14387 ( .IN1(n9269), .IN2(n13147), .Q(n13921) );
  OR2X1 U14388 ( .IN1(n13922), .IN2(n13923), .Q(n13147) );
  INVX0 U14389 ( .INP(n13924), .ZN(n13923) );
  OR2X1 U14390 ( .IN1(n13925), .IN2(n13926), .Q(n13924) );
  AND2X1 U14391 ( .IN1(n13926), .IN2(n13925), .Q(n13922) );
  AND2X1 U14392 ( .IN1(n13927), .IN2(n13928), .Q(n13925) );
  OR2X1 U14393 ( .IN1(WX3331), .IN2(n8589), .Q(n13928) );
  INVX0 U14394 ( .INP(n13929), .ZN(n13927) );
  AND2X1 U14395 ( .IN1(n8589), .IN2(WX3331), .Q(n13929) );
  OR2X1 U14396 ( .IN1(n13930), .IN2(n13931), .Q(n13926) );
  AND2X1 U14397 ( .IN1(n8590), .IN2(WX3459), .Q(n13931) );
  AND2X1 U14398 ( .IN1(n8918), .IN2(WX3395), .Q(n13930) );
  AND2X1 U14399 ( .IN1(n9188), .IN2(n11434), .Q(n13920) );
  OR2X1 U14400 ( .IN1(n13932), .IN2(n13933), .Q(n11434) );
  INVX0 U14401 ( .INP(n13934), .ZN(n13933) );
  OR2X1 U14402 ( .IN1(n13935), .IN2(n13936), .Q(n13934) );
  AND2X1 U14403 ( .IN1(n13936), .IN2(n13935), .Q(n13932) );
  AND2X1 U14404 ( .IN1(n13937), .IN2(n13938), .Q(n13935) );
  OR2X1 U14405 ( .IN1(WX2038), .IN2(n8708), .Q(n13938) );
  INVX0 U14406 ( .INP(n13939), .ZN(n13937) );
  AND2X1 U14407 ( .IN1(n8708), .IN2(WX2038), .Q(n13939) );
  OR2X1 U14408 ( .IN1(n13940), .IN2(n13941), .Q(n13936) );
  AND2X1 U14409 ( .IN1(n8709), .IN2(WX2166), .Q(n13941) );
  AND2X1 U14410 ( .IN1(n8944), .IN2(WX2102), .Q(n13940) );
  AND2X1 U14411 ( .IN1(n9234), .IN2(CRC_OUT_8_13), .Q(n13919) );
  AND2X1 U14412 ( .IN1(n284), .IN2(n9208), .Q(n13918) );
  INVX0 U14413 ( .INP(n13942), .ZN(n284) );
  OR2X1 U14414 ( .IN1(n9561), .IN2(n4016), .Q(n13942) );
  OR4X1 U14415 ( .IN1(n13943), .IN2(n13944), .IN3(n13945), .IN4(n13946), .Q(
        WX1971) );
  AND2X1 U14416 ( .IN1(n9269), .IN2(n13163), .Q(n13946) );
  OR2X1 U14417 ( .IN1(n13947), .IN2(n13948), .Q(n13163) );
  INVX0 U14418 ( .INP(n13949), .ZN(n13948) );
  OR2X1 U14419 ( .IN1(n13950), .IN2(n13951), .Q(n13949) );
  AND2X1 U14420 ( .IN1(n13951), .IN2(n13950), .Q(n13947) );
  AND2X1 U14421 ( .IN1(n13952), .IN2(n13953), .Q(n13950) );
  OR2X1 U14422 ( .IN1(WX3329), .IN2(n8591), .Q(n13953) );
  INVX0 U14423 ( .INP(n13954), .ZN(n13952) );
  AND2X1 U14424 ( .IN1(n8591), .IN2(WX3329), .Q(n13954) );
  OR2X1 U14425 ( .IN1(n13955), .IN2(n13956), .Q(n13951) );
  AND2X1 U14426 ( .IN1(n8592), .IN2(WX3457), .Q(n13956) );
  AND2X1 U14427 ( .IN1(n8917), .IN2(WX3393), .Q(n13955) );
  AND2X1 U14428 ( .IN1(n11440), .IN2(n9175), .Q(n13945) );
  AND2X1 U14429 ( .IN1(n13957), .IN2(n13958), .Q(n11440) );
  INVX0 U14430 ( .INP(n13959), .ZN(n13958) );
  AND2X1 U14431 ( .IN1(n13960), .IN2(n13961), .Q(n13959) );
  OR2X1 U14432 ( .IN1(n13961), .IN2(n13960), .Q(n13957) );
  OR2X1 U14433 ( .IN1(n13962), .IN2(n13963), .Q(n13960) );
  INVX0 U14434 ( .INP(n13964), .ZN(n13963) );
  OR2X1 U14435 ( .IN1(WX2036), .IN2(n8710), .Q(n13964) );
  AND2X1 U14436 ( .IN1(n8710), .IN2(WX2036), .Q(n13962) );
  AND2X1 U14437 ( .IN1(n13965), .IN2(n13966), .Q(n13961) );
  OR2X1 U14438 ( .IN1(WX2164), .IN2(test_so17), .Q(n13966) );
  OR2X1 U14439 ( .IN1(n9138), .IN2(n8943), .Q(n13965) );
  AND2X1 U14440 ( .IN1(n9234), .IN2(CRC_OUT_8_14), .Q(n13944) );
  AND2X1 U14441 ( .IN1(n283), .IN2(n9208), .Q(n13943) );
  INVX0 U14442 ( .INP(n13967), .ZN(n283) );
  OR2X1 U14443 ( .IN1(n9560), .IN2(n4017), .Q(n13967) );
  OR4X1 U14444 ( .IN1(n13968), .IN2(n13969), .IN3(n13970), .IN4(n13971), .Q(
        WX1969) );
  AND2X1 U14445 ( .IN1(n9269), .IN2(n13179), .Q(n13971) );
  OR2X1 U14446 ( .IN1(n13972), .IN2(n13973), .Q(n13179) );
  INVX0 U14447 ( .INP(n13974), .ZN(n13973) );
  OR2X1 U14448 ( .IN1(n13975), .IN2(n13976), .Q(n13974) );
  AND2X1 U14449 ( .IN1(n13976), .IN2(n13975), .Q(n13972) );
  AND2X1 U14450 ( .IN1(n13977), .IN2(n13978), .Q(n13975) );
  OR2X1 U14451 ( .IN1(WX3327), .IN2(n8593), .Q(n13978) );
  INVX0 U14452 ( .INP(n13979), .ZN(n13977) );
  AND2X1 U14453 ( .IN1(n8593), .IN2(WX3327), .Q(n13979) );
  OR2X1 U14454 ( .IN1(n13980), .IN2(n13981), .Q(n13976) );
  AND2X1 U14455 ( .IN1(n8594), .IN2(WX3455), .Q(n13981) );
  AND2X1 U14456 ( .IN1(n8916), .IN2(WX3391), .Q(n13980) );
  AND2X1 U14457 ( .IN1(n9188), .IN2(n11446), .Q(n13970) );
  OR2X1 U14458 ( .IN1(n13982), .IN2(n13983), .Q(n11446) );
  INVX0 U14459 ( .INP(n13984), .ZN(n13983) );
  OR2X1 U14460 ( .IN1(n13985), .IN2(n13986), .Q(n13984) );
  AND2X1 U14461 ( .IN1(n13986), .IN2(n13985), .Q(n13982) );
  AND2X1 U14462 ( .IN1(n13987), .IN2(n13988), .Q(n13985) );
  OR2X1 U14463 ( .IN1(WX2034), .IN2(n8711), .Q(n13988) );
  INVX0 U14464 ( .INP(n13989), .ZN(n13987) );
  AND2X1 U14465 ( .IN1(n8711), .IN2(WX2034), .Q(n13989) );
  OR2X1 U14466 ( .IN1(n13990), .IN2(n13991), .Q(n13986) );
  AND2X1 U14467 ( .IN1(n8712), .IN2(WX2162), .Q(n13991) );
  AND2X1 U14468 ( .IN1(n8942), .IN2(WX2098), .Q(n13990) );
  AND2X1 U14469 ( .IN1(n9235), .IN2(CRC_OUT_8_15), .Q(n13969) );
  AND2X1 U14470 ( .IN1(n282), .IN2(n9208), .Q(n13968) );
  INVX0 U14471 ( .INP(n13992), .ZN(n282) );
  OR2X1 U14472 ( .IN1(n9560), .IN2(n4018), .Q(n13992) );
  OR4X1 U14473 ( .IN1(n13993), .IN2(n13994), .IN3(n13995), .IN4(n13996), .Q(
        WX1967) );
  AND2X1 U14474 ( .IN1(n13195), .IN2(n9260), .Q(n13996) );
  AND2X1 U14475 ( .IN1(n13997), .IN2(n13998), .Q(n13195) );
  OR2X1 U14476 ( .IN1(n13999), .IN2(n14000), .Q(n13998) );
  INVX0 U14477 ( .INP(n14001), .ZN(n13997) );
  AND2X1 U14478 ( .IN1(n14000), .IN2(n13999), .Q(n14001) );
  INVX0 U14479 ( .INP(n14002), .ZN(n13999) );
  OR2X1 U14480 ( .IN1(n14003), .IN2(n14004), .Q(n14002) );
  AND2X1 U14481 ( .IN1(n9450), .IN2(WX3453), .Q(n14004) );
  AND2X1 U14482 ( .IN1(n8728), .IN2(n9463), .Q(n14003) );
  OR2X1 U14483 ( .IN1(n14005), .IN2(n14006), .Q(n14000) );
  AND3X1 U14484 ( .IN1(n14007), .IN2(n14008), .IN3(n8062), .Q(n14006) );
  OR2X1 U14485 ( .IN1(n8061), .IN2(n9095), .Q(n14008) );
  OR2X1 U14486 ( .IN1(test_so24), .IN2(WX3325), .Q(n14007) );
  AND2X1 U14487 ( .IN1(n14009), .IN2(WX3389), .Q(n14005) );
  OR2X1 U14488 ( .IN1(n14010), .IN2(n14011), .Q(n14009) );
  AND2X1 U14489 ( .IN1(n8061), .IN2(n9095), .Q(n14011) );
  AND2X1 U14490 ( .IN1(test_so24), .IN2(WX3325), .Q(n14010) );
  AND2X1 U14491 ( .IN1(n9188), .IN2(n11452), .Q(n13995) );
  OR2X1 U14492 ( .IN1(n14012), .IN2(n14013), .Q(n11452) );
  INVX0 U14493 ( .INP(n14014), .ZN(n14013) );
  OR2X1 U14494 ( .IN1(n14015), .IN2(n14016), .Q(n14014) );
  AND2X1 U14495 ( .IN1(n14016), .IN2(n14015), .Q(n14012) );
  AND2X1 U14496 ( .IN1(n14017), .IN2(n14018), .Q(n14015) );
  OR2X1 U14497 ( .IN1(n9459), .IN2(n8089), .Q(n14018) );
  OR2X1 U14498 ( .IN1(WX2032), .IN2(n9445), .Q(n14017) );
  OR2X1 U14499 ( .IN1(n14019), .IN2(n14020), .Q(n14016) );
  INVX0 U14500 ( .INP(n14021), .ZN(n14020) );
  OR2X1 U14501 ( .IN1(n14022), .IN2(n8090), .Q(n14021) );
  AND2X1 U14502 ( .IN1(n8090), .IN2(n14022), .Q(n14019) );
  INVX0 U14503 ( .INP(n14023), .ZN(n14022) );
  OR2X1 U14504 ( .IN1(n14024), .IN2(n14025), .Q(n14023) );
  AND2X1 U14505 ( .IN1(n8731), .IN2(n8653), .Q(n14025) );
  AND2X1 U14506 ( .IN1(n15953), .IN2(WX2160), .Q(n14024) );
  AND2X1 U14507 ( .IN1(n9235), .IN2(CRC_OUT_8_16), .Q(n13994) );
  AND2X1 U14508 ( .IN1(n281), .IN2(n9208), .Q(n13993) );
  INVX0 U14509 ( .INP(n14026), .ZN(n281) );
  OR2X1 U14510 ( .IN1(n9560), .IN2(n4019), .Q(n14026) );
  OR4X1 U14511 ( .IN1(n14027), .IN2(n14028), .IN3(n14029), .IN4(n14030), .Q(
        WX1965) );
  AND2X1 U14512 ( .IN1(n9269), .IN2(n13215), .Q(n14030) );
  OR2X1 U14513 ( .IN1(n14031), .IN2(n14032), .Q(n13215) );
  INVX0 U14514 ( .INP(n14033), .ZN(n14032) );
  OR2X1 U14515 ( .IN1(n14034), .IN2(n14035), .Q(n14033) );
  AND2X1 U14516 ( .IN1(n14035), .IN2(n14034), .Q(n14031) );
  AND2X1 U14517 ( .IN1(n14036), .IN2(n14037), .Q(n14034) );
  OR2X1 U14518 ( .IN1(n9459), .IN2(n8063), .Q(n14037) );
  OR2X1 U14519 ( .IN1(WX3323), .IN2(n9444), .Q(n14036) );
  OR2X1 U14520 ( .IN1(n14038), .IN2(n14039), .Q(n14035) );
  INVX0 U14521 ( .INP(n14040), .ZN(n14039) );
  OR2X1 U14522 ( .IN1(n14041), .IN2(n8064), .Q(n14040) );
  AND2X1 U14523 ( .IN1(n8064), .IN2(n14041), .Q(n14038) );
  INVX0 U14524 ( .INP(n14042), .ZN(n14041) );
  OR2X1 U14525 ( .IN1(n14043), .IN2(n14044), .Q(n14042) );
  AND2X1 U14526 ( .IN1(n8915), .IN2(n8597), .Q(n14044) );
  AND2X1 U14527 ( .IN1(n15955), .IN2(WX3451), .Q(n14043) );
  AND2X1 U14528 ( .IN1(n9188), .IN2(n11458), .Q(n14029) );
  OR2X1 U14529 ( .IN1(n14045), .IN2(n14046), .Q(n11458) );
  INVX0 U14530 ( .INP(n14047), .ZN(n14046) );
  OR2X1 U14531 ( .IN1(n14048), .IN2(n14049), .Q(n14047) );
  AND2X1 U14532 ( .IN1(n14049), .IN2(n14048), .Q(n14045) );
  AND2X1 U14533 ( .IN1(n14050), .IN2(n14051), .Q(n14048) );
  OR2X1 U14534 ( .IN1(n9460), .IN2(n8091), .Q(n14051) );
  OR2X1 U14535 ( .IN1(WX2030), .IN2(n9444), .Q(n14050) );
  OR2X1 U14536 ( .IN1(n14052), .IN2(n14053), .Q(n14049) );
  INVX0 U14537 ( .INP(n14054), .ZN(n14053) );
  OR2X1 U14538 ( .IN1(n14055), .IN2(n8092), .Q(n14054) );
  AND2X1 U14539 ( .IN1(n8092), .IN2(n14055), .Q(n14052) );
  INVX0 U14540 ( .INP(n14056), .ZN(n14055) );
  OR2X1 U14541 ( .IN1(n14057), .IN2(n14058), .Q(n14056) );
  AND2X1 U14542 ( .IN1(n8941), .IN2(n8654), .Q(n14058) );
  AND2X1 U14543 ( .IN1(n15954), .IN2(WX2158), .Q(n14057) );
  AND2X1 U14544 ( .IN1(n9235), .IN2(CRC_OUT_8_17), .Q(n14028) );
  AND2X1 U14545 ( .IN1(n280), .IN2(n9209), .Q(n14027) );
  INVX0 U14546 ( .INP(n14059), .ZN(n280) );
  OR2X1 U14547 ( .IN1(n9560), .IN2(n4020), .Q(n14059) );
  OR4X1 U14548 ( .IN1(n14060), .IN2(n14061), .IN3(n14062), .IN4(n14063), .Q(
        WX1963) );
  AND2X1 U14549 ( .IN1(n9269), .IN2(n13236), .Q(n14063) );
  OR2X1 U14550 ( .IN1(n14064), .IN2(n14065), .Q(n13236) );
  INVX0 U14551 ( .INP(n14066), .ZN(n14065) );
  OR2X1 U14552 ( .IN1(n14067), .IN2(n14068), .Q(n14066) );
  AND2X1 U14553 ( .IN1(n14068), .IN2(n14067), .Q(n14064) );
  AND2X1 U14554 ( .IN1(n14069), .IN2(n14070), .Q(n14067) );
  OR2X1 U14555 ( .IN1(n9460), .IN2(n8065), .Q(n14070) );
  OR2X1 U14556 ( .IN1(WX3321), .IN2(n9444), .Q(n14069) );
  OR2X1 U14557 ( .IN1(n14071), .IN2(n14072), .Q(n14068) );
  INVX0 U14558 ( .INP(n14073), .ZN(n14072) );
  OR2X1 U14559 ( .IN1(n14074), .IN2(n8066), .Q(n14073) );
  AND2X1 U14560 ( .IN1(n8066), .IN2(n14074), .Q(n14071) );
  INVX0 U14561 ( .INP(n14075), .ZN(n14074) );
  OR2X1 U14562 ( .IN1(n14076), .IN2(n14077), .Q(n14075) );
  AND2X1 U14563 ( .IN1(n8914), .IN2(n8598), .Q(n14077) );
  AND2X1 U14564 ( .IN1(n15957), .IN2(WX3449), .Q(n14076) );
  AND2X1 U14565 ( .IN1(n11464), .IN2(n9176), .Q(n14062) );
  AND2X1 U14566 ( .IN1(n14078), .IN2(n14079), .Q(n11464) );
  INVX0 U14567 ( .INP(n14080), .ZN(n14079) );
  AND2X1 U14568 ( .IN1(n14081), .IN2(n14082), .Q(n14080) );
  OR2X1 U14569 ( .IN1(n14082), .IN2(n14081), .Q(n14078) );
  OR2X1 U14570 ( .IN1(n14083), .IN2(n14084), .Q(n14081) );
  AND2X1 U14571 ( .IN1(n9450), .IN2(WX2092), .Q(n14084) );
  AND2X1 U14572 ( .IN1(n8093), .IN2(n9475), .Q(n14083) );
  AND2X1 U14573 ( .IN1(n14085), .IN2(n14086), .Q(n14082) );
  OR2X1 U14574 ( .IN1(n14087), .IN2(n8940), .Q(n14086) );
  OR2X1 U14575 ( .IN1(WX2156), .IN2(n14088), .Q(n14085) );
  INVX0 U14576 ( .INP(n14087), .ZN(n14088) );
  AND2X1 U14577 ( .IN1(n14089), .IN2(n14090), .Q(n14087) );
  OR2X1 U14578 ( .IN1(n8655), .IN2(test_so15), .Q(n14090) );
  OR2X1 U14579 ( .IN1(n9139), .IN2(n15956), .Q(n14089) );
  AND2X1 U14580 ( .IN1(n9235), .IN2(CRC_OUT_8_18), .Q(n14061) );
  AND2X1 U14581 ( .IN1(n279), .IN2(n9209), .Q(n14060) );
  INVX0 U14582 ( .INP(n14091), .ZN(n279) );
  OR2X1 U14583 ( .IN1(n9560), .IN2(n4021), .Q(n14091) );
  OR4X1 U14584 ( .IN1(n14092), .IN2(n14093), .IN3(n14094), .IN4(n14095), .Q(
        WX1961) );
  AND2X1 U14585 ( .IN1(n9269), .IN2(n13256), .Q(n14095) );
  OR2X1 U14586 ( .IN1(n14096), .IN2(n14097), .Q(n13256) );
  INVX0 U14587 ( .INP(n14098), .ZN(n14097) );
  OR2X1 U14588 ( .IN1(n14099), .IN2(n14100), .Q(n14098) );
  AND2X1 U14589 ( .IN1(n14100), .IN2(n14099), .Q(n14096) );
  AND2X1 U14590 ( .IN1(n14101), .IN2(n14102), .Q(n14099) );
  OR2X1 U14591 ( .IN1(n9461), .IN2(n8067), .Q(n14102) );
  OR2X1 U14592 ( .IN1(WX3319), .IN2(n9444), .Q(n14101) );
  OR2X1 U14593 ( .IN1(n14103), .IN2(n14104), .Q(n14100) );
  INVX0 U14594 ( .INP(n14105), .ZN(n14104) );
  OR2X1 U14595 ( .IN1(n14106), .IN2(n8068), .Q(n14105) );
  AND2X1 U14596 ( .IN1(n8068), .IN2(n14106), .Q(n14103) );
  INVX0 U14597 ( .INP(n14107), .ZN(n14106) );
  OR2X1 U14598 ( .IN1(n14108), .IN2(n14109), .Q(n14107) );
  AND2X1 U14599 ( .IN1(n8913), .IN2(n8599), .Q(n14109) );
  AND2X1 U14600 ( .IN1(n15959), .IN2(WX3447), .Q(n14108) );
  AND2X1 U14601 ( .IN1(n9188), .IN2(n11470), .Q(n14094) );
  OR2X1 U14602 ( .IN1(n14110), .IN2(n14111), .Q(n11470) );
  INVX0 U14603 ( .INP(n14112), .ZN(n14111) );
  OR2X1 U14604 ( .IN1(n14113), .IN2(n14114), .Q(n14112) );
  AND2X1 U14605 ( .IN1(n14114), .IN2(n14113), .Q(n14110) );
  AND2X1 U14606 ( .IN1(n14115), .IN2(n14116), .Q(n14113) );
  OR2X1 U14607 ( .IN1(n9462), .IN2(n8094), .Q(n14116) );
  OR2X1 U14608 ( .IN1(WX2026), .IN2(n9444), .Q(n14115) );
  OR2X1 U14609 ( .IN1(n14117), .IN2(n14118), .Q(n14114) );
  INVX0 U14610 ( .INP(n14119), .ZN(n14118) );
  OR2X1 U14611 ( .IN1(n14120), .IN2(n8095), .Q(n14119) );
  AND2X1 U14612 ( .IN1(n8095), .IN2(n14120), .Q(n14117) );
  INVX0 U14613 ( .INP(n14121), .ZN(n14120) );
  OR2X1 U14614 ( .IN1(n14122), .IN2(n14123), .Q(n14121) );
  AND2X1 U14615 ( .IN1(n8939), .IN2(n8656), .Q(n14123) );
  AND2X1 U14616 ( .IN1(n15958), .IN2(WX2154), .Q(n14122) );
  AND2X1 U14617 ( .IN1(n9235), .IN2(CRC_OUT_8_19), .Q(n14093) );
  AND2X1 U14618 ( .IN1(n278), .IN2(n9209), .Q(n14092) );
  INVX0 U14619 ( .INP(n14124), .ZN(n278) );
  OR2X1 U14620 ( .IN1(n9560), .IN2(n4022), .Q(n14124) );
  OR4X1 U14621 ( .IN1(n14125), .IN2(n14126), .IN3(n14127), .IN4(n14128), .Q(
        WX1959) );
  AND2X1 U14622 ( .IN1(n9269), .IN2(n13276), .Q(n14128) );
  OR2X1 U14623 ( .IN1(n14129), .IN2(n14130), .Q(n13276) );
  INVX0 U14624 ( .INP(n14131), .ZN(n14130) );
  OR2X1 U14625 ( .IN1(n14132), .IN2(n14133), .Q(n14131) );
  AND2X1 U14626 ( .IN1(n14133), .IN2(n14132), .Q(n14129) );
  AND2X1 U14627 ( .IN1(n14134), .IN2(n14135), .Q(n14132) );
  OR2X1 U14628 ( .IN1(n9462), .IN2(n8069), .Q(n14135) );
  OR2X1 U14629 ( .IN1(WX3317), .IN2(n9444), .Q(n14134) );
  OR2X1 U14630 ( .IN1(n14136), .IN2(n14137), .Q(n14133) );
  INVX0 U14631 ( .INP(n14138), .ZN(n14137) );
  OR2X1 U14632 ( .IN1(n14139), .IN2(n8070), .Q(n14138) );
  AND2X1 U14633 ( .IN1(n8070), .IN2(n14139), .Q(n14136) );
  INVX0 U14634 ( .INP(n14140), .ZN(n14139) );
  OR2X1 U14635 ( .IN1(n14141), .IN2(n14142), .Q(n14140) );
  AND2X1 U14636 ( .IN1(n8912), .IN2(n8600), .Q(n14142) );
  AND2X1 U14637 ( .IN1(n15961), .IN2(WX3445), .Q(n14141) );
  AND2X1 U14638 ( .IN1(n9188), .IN2(n11476), .Q(n14127) );
  OR2X1 U14639 ( .IN1(n14143), .IN2(n14144), .Q(n11476) );
  INVX0 U14640 ( .INP(n14145), .ZN(n14144) );
  OR2X1 U14641 ( .IN1(n14146), .IN2(n14147), .Q(n14145) );
  AND2X1 U14642 ( .IN1(n14147), .IN2(n14146), .Q(n14143) );
  AND2X1 U14643 ( .IN1(n14148), .IN2(n14149), .Q(n14146) );
  OR2X1 U14644 ( .IN1(n9463), .IN2(n8096), .Q(n14149) );
  OR2X1 U14645 ( .IN1(WX2024), .IN2(n9444), .Q(n14148) );
  OR2X1 U14646 ( .IN1(n14150), .IN2(n14151), .Q(n14147) );
  INVX0 U14647 ( .INP(n14152), .ZN(n14151) );
  OR2X1 U14648 ( .IN1(n14153), .IN2(n8097), .Q(n14152) );
  AND2X1 U14649 ( .IN1(n8097), .IN2(n14153), .Q(n14150) );
  INVX0 U14650 ( .INP(n14154), .ZN(n14153) );
  OR2X1 U14651 ( .IN1(n14155), .IN2(n14156), .Q(n14154) );
  AND2X1 U14652 ( .IN1(n8938), .IN2(n8657), .Q(n14156) );
  AND2X1 U14653 ( .IN1(n15960), .IN2(WX2152), .Q(n14155) );
  AND2X1 U14654 ( .IN1(n9235), .IN2(CRC_OUT_8_20), .Q(n14126) );
  AND2X1 U14655 ( .IN1(n277), .IN2(n9209), .Q(n14125) );
  INVX0 U14656 ( .INP(n14157), .ZN(n277) );
  OR2X1 U14657 ( .IN1(n9560), .IN2(n4023), .Q(n14157) );
  OR4X1 U14658 ( .IN1(n14158), .IN2(n14159), .IN3(n14160), .IN4(n14161), .Q(
        WX1957) );
  AND2X1 U14659 ( .IN1(n9269), .IN2(n13296), .Q(n14161) );
  OR2X1 U14660 ( .IN1(n14162), .IN2(n14163), .Q(n13296) );
  INVX0 U14661 ( .INP(n14164), .ZN(n14163) );
  OR2X1 U14662 ( .IN1(n14165), .IN2(n14166), .Q(n14164) );
  AND2X1 U14663 ( .IN1(n14166), .IN2(n14165), .Q(n14162) );
  AND2X1 U14664 ( .IN1(n14167), .IN2(n14168), .Q(n14165) );
  OR2X1 U14665 ( .IN1(n9463), .IN2(n8071), .Q(n14168) );
  OR2X1 U14666 ( .IN1(WX3315), .IN2(n9444), .Q(n14167) );
  OR2X1 U14667 ( .IN1(n14169), .IN2(n14170), .Q(n14166) );
  INVX0 U14668 ( .INP(n14171), .ZN(n14170) );
  OR2X1 U14669 ( .IN1(n14172), .IN2(n8072), .Q(n14171) );
  AND2X1 U14670 ( .IN1(n8072), .IN2(n14172), .Q(n14169) );
  INVX0 U14671 ( .INP(n14173), .ZN(n14172) );
  OR2X1 U14672 ( .IN1(n14174), .IN2(n14175), .Q(n14173) );
  AND2X1 U14673 ( .IN1(n8911), .IN2(n8601), .Q(n14175) );
  AND2X1 U14674 ( .IN1(n15963), .IN2(WX3443), .Q(n14174) );
  AND2X1 U14675 ( .IN1(n9188), .IN2(n11482), .Q(n14160) );
  OR2X1 U14676 ( .IN1(n14176), .IN2(n14177), .Q(n11482) );
  INVX0 U14677 ( .INP(n14178), .ZN(n14177) );
  OR2X1 U14678 ( .IN1(n14179), .IN2(n14180), .Q(n14178) );
  AND2X1 U14679 ( .IN1(n14180), .IN2(n14179), .Q(n14176) );
  AND2X1 U14680 ( .IN1(n14181), .IN2(n14182), .Q(n14179) );
  OR2X1 U14681 ( .IN1(n9464), .IN2(n8098), .Q(n14182) );
  OR2X1 U14682 ( .IN1(WX2022), .IN2(n9444), .Q(n14181) );
  OR2X1 U14683 ( .IN1(n14183), .IN2(n14184), .Q(n14180) );
  INVX0 U14684 ( .INP(n14185), .ZN(n14184) );
  OR2X1 U14685 ( .IN1(n14186), .IN2(n8099), .Q(n14185) );
  AND2X1 U14686 ( .IN1(n8099), .IN2(n14186), .Q(n14183) );
  INVX0 U14687 ( .INP(n14187), .ZN(n14186) );
  OR2X1 U14688 ( .IN1(n14188), .IN2(n14189), .Q(n14187) );
  AND2X1 U14689 ( .IN1(n8937), .IN2(n8658), .Q(n14189) );
  AND2X1 U14690 ( .IN1(n15962), .IN2(WX2150), .Q(n14188) );
  AND2X1 U14691 ( .IN1(n9235), .IN2(CRC_OUT_8_21), .Q(n14159) );
  AND2X1 U14692 ( .IN1(n276), .IN2(n9209), .Q(n14158) );
  INVX0 U14693 ( .INP(n14190), .ZN(n276) );
  OR2X1 U14694 ( .IN1(n9560), .IN2(n4024), .Q(n14190) );
  OR4X1 U14695 ( .IN1(n14191), .IN2(n14192), .IN3(n14193), .IN4(n14194), .Q(
        WX1955) );
  AND2X1 U14696 ( .IN1(n9269), .IN2(n13316), .Q(n14194) );
  OR2X1 U14697 ( .IN1(n14195), .IN2(n14196), .Q(n13316) );
  INVX0 U14698 ( .INP(n14197), .ZN(n14196) );
  OR2X1 U14699 ( .IN1(n14198), .IN2(n14199), .Q(n14197) );
  AND2X1 U14700 ( .IN1(n14199), .IN2(n14198), .Q(n14195) );
  AND2X1 U14701 ( .IN1(n14200), .IN2(n14201), .Q(n14198) );
  OR2X1 U14702 ( .IN1(n9464), .IN2(n8073), .Q(n14201) );
  OR2X1 U14703 ( .IN1(WX3313), .IN2(n9444), .Q(n14200) );
  OR2X1 U14704 ( .IN1(n14202), .IN2(n14203), .Q(n14199) );
  INVX0 U14705 ( .INP(n14204), .ZN(n14203) );
  OR2X1 U14706 ( .IN1(n14205), .IN2(n8074), .Q(n14204) );
  AND2X1 U14707 ( .IN1(n8074), .IN2(n14205), .Q(n14202) );
  INVX0 U14708 ( .INP(n14206), .ZN(n14205) );
  OR2X1 U14709 ( .IN1(n14207), .IN2(n14208), .Q(n14206) );
  AND2X1 U14710 ( .IN1(n8910), .IN2(n8602), .Q(n14208) );
  AND2X1 U14711 ( .IN1(n15964), .IN2(WX3441), .Q(n14207) );
  AND2X1 U14712 ( .IN1(n11488), .IN2(n9175), .Q(n14193) );
  AND2X1 U14713 ( .IN1(n14209), .IN2(n14210), .Q(n11488) );
  OR2X1 U14714 ( .IN1(n14211), .IN2(n14212), .Q(n14210) );
  INVX0 U14715 ( .INP(n14213), .ZN(n14209) );
  AND2X1 U14716 ( .IN1(n14212), .IN2(n14211), .Q(n14213) );
  INVX0 U14717 ( .INP(n14214), .ZN(n14211) );
  OR2X1 U14718 ( .IN1(n14215), .IN2(n14216), .Q(n14214) );
  AND2X1 U14719 ( .IN1(n9450), .IN2(WX2148), .Q(n14216) );
  AND2X1 U14720 ( .IN1(n8936), .IN2(n9466), .Q(n14215) );
  OR2X1 U14721 ( .IN1(n14217), .IN2(n14218), .Q(n14212) );
  AND3X1 U14722 ( .IN1(n14219), .IN2(n14220), .IN3(n8101), .Q(n14218) );
  OR2X1 U14723 ( .IN1(n8100), .IN2(n9096), .Q(n14220) );
  OR2X1 U14724 ( .IN1(test_so13), .IN2(WX2020), .Q(n14219) );
  AND2X1 U14725 ( .IN1(n14221), .IN2(WX2084), .Q(n14217) );
  OR2X1 U14726 ( .IN1(n14222), .IN2(n14223), .Q(n14221) );
  AND2X1 U14727 ( .IN1(n8100), .IN2(n9096), .Q(n14223) );
  AND2X1 U14728 ( .IN1(test_so13), .IN2(WX2020), .Q(n14222) );
  AND2X1 U14729 ( .IN1(n9235), .IN2(CRC_OUT_8_22), .Q(n14192) );
  AND2X1 U14730 ( .IN1(n275), .IN2(n9209), .Q(n14191) );
  INVX0 U14731 ( .INP(n14224), .ZN(n275) );
  OR2X1 U14732 ( .IN1(n9560), .IN2(n4025), .Q(n14224) );
  OR4X1 U14733 ( .IN1(n14225), .IN2(n14226), .IN3(n14227), .IN4(n14228), .Q(
        WX1953) );
  AND2X1 U14734 ( .IN1(n13336), .IN2(n9260), .Q(n14228) );
  AND2X1 U14735 ( .IN1(n14229), .IN2(n14230), .Q(n13336) );
  INVX0 U14736 ( .INP(n14231), .ZN(n14230) );
  AND2X1 U14737 ( .IN1(n14232), .IN2(n14233), .Q(n14231) );
  OR2X1 U14738 ( .IN1(n14233), .IN2(n14232), .Q(n14229) );
  OR2X1 U14739 ( .IN1(n14234), .IN2(n14235), .Q(n14232) );
  AND2X1 U14740 ( .IN1(n9451), .IN2(WX3311), .Q(n14235) );
  AND2X1 U14741 ( .IN1(n8075), .IN2(n9479), .Q(n14234) );
  AND2X1 U14742 ( .IN1(n14236), .IN2(n14237), .Q(n14233) );
  OR2X1 U14743 ( .IN1(n14238), .IN2(n8076), .Q(n14237) );
  INVX0 U14744 ( .INP(n14239), .ZN(n14238) );
  OR2X1 U14745 ( .IN1(WX3375), .IN2(n14239), .Q(n14236) );
  OR2X1 U14746 ( .IN1(n14240), .IN2(n14241), .Q(n14239) );
  AND2X1 U14747 ( .IN1(n15966), .IN2(n9107), .Q(n14241) );
  AND2X1 U14748 ( .IN1(test_so29), .IN2(n8603), .Q(n14240) );
  AND2X1 U14749 ( .IN1(n9188), .IN2(n11494), .Q(n14227) );
  OR2X1 U14750 ( .IN1(n14242), .IN2(n14243), .Q(n11494) );
  INVX0 U14751 ( .INP(n14244), .ZN(n14243) );
  OR2X1 U14752 ( .IN1(n14245), .IN2(n14246), .Q(n14244) );
  AND2X1 U14753 ( .IN1(n14246), .IN2(n14245), .Q(n14242) );
  AND2X1 U14754 ( .IN1(n14247), .IN2(n14248), .Q(n14245) );
  OR2X1 U14755 ( .IN1(n9466), .IN2(n8102), .Q(n14248) );
  OR2X1 U14756 ( .IN1(WX2018), .IN2(n9444), .Q(n14247) );
  OR2X1 U14757 ( .IN1(n14249), .IN2(n14250), .Q(n14246) );
  INVX0 U14758 ( .INP(n14251), .ZN(n14250) );
  OR2X1 U14759 ( .IN1(n14252), .IN2(n8103), .Q(n14251) );
  AND2X1 U14760 ( .IN1(n8103), .IN2(n14252), .Q(n14249) );
  INVX0 U14761 ( .INP(n14253), .ZN(n14252) );
  OR2X1 U14762 ( .IN1(n14254), .IN2(n14255), .Q(n14253) );
  AND2X1 U14763 ( .IN1(n8935), .IN2(n8661), .Q(n14255) );
  AND2X1 U14764 ( .IN1(n15965), .IN2(WX2146), .Q(n14254) );
  AND2X1 U14765 ( .IN1(n9235), .IN2(CRC_OUT_8_23), .Q(n14226) );
  AND2X1 U14766 ( .IN1(n274), .IN2(n9209), .Q(n14225) );
  INVX0 U14767 ( .INP(n14256), .ZN(n274) );
  OR2X1 U14768 ( .IN1(n9560), .IN2(n4026), .Q(n14256) );
  OR4X1 U14769 ( .IN1(n14257), .IN2(n14258), .IN3(n14259), .IN4(n14260), .Q(
        WX1951) );
  AND2X1 U14770 ( .IN1(n9269), .IN2(n13357), .Q(n14260) );
  OR2X1 U14771 ( .IN1(n14261), .IN2(n14262), .Q(n13357) );
  INVX0 U14772 ( .INP(n14263), .ZN(n14262) );
  OR2X1 U14773 ( .IN1(n14264), .IN2(n14265), .Q(n14263) );
  AND2X1 U14774 ( .IN1(n14265), .IN2(n14264), .Q(n14261) );
  AND2X1 U14775 ( .IN1(n14266), .IN2(n14267), .Q(n14264) );
  OR2X1 U14776 ( .IN1(n9466), .IN2(n8077), .Q(n14267) );
  OR2X1 U14777 ( .IN1(WX3309), .IN2(n9444), .Q(n14266) );
  OR2X1 U14778 ( .IN1(n14268), .IN2(n14269), .Q(n14265) );
  INVX0 U14779 ( .INP(n14270), .ZN(n14269) );
  OR2X1 U14780 ( .IN1(n14271), .IN2(n8078), .Q(n14270) );
  AND2X1 U14781 ( .IN1(n8078), .IN2(n14271), .Q(n14268) );
  INVX0 U14782 ( .INP(n14272), .ZN(n14271) );
  OR2X1 U14783 ( .IN1(n14273), .IN2(n14274), .Q(n14272) );
  AND2X1 U14784 ( .IN1(n8909), .IN2(n8604), .Q(n14274) );
  AND2X1 U14785 ( .IN1(n15968), .IN2(WX3437), .Q(n14273) );
  AND2X1 U14786 ( .IN1(n9188), .IN2(n11500), .Q(n14259) );
  OR2X1 U14787 ( .IN1(n14275), .IN2(n14276), .Q(n11500) );
  INVX0 U14788 ( .INP(n14277), .ZN(n14276) );
  OR2X1 U14789 ( .IN1(n14278), .IN2(n14279), .Q(n14277) );
  AND2X1 U14790 ( .IN1(n14279), .IN2(n14278), .Q(n14275) );
  AND2X1 U14791 ( .IN1(n14280), .IN2(n14281), .Q(n14278) );
  OR2X1 U14792 ( .IN1(n9461), .IN2(n8104), .Q(n14281) );
  OR2X1 U14793 ( .IN1(WX2016), .IN2(n9443), .Q(n14280) );
  OR2X1 U14794 ( .IN1(n14282), .IN2(n14283), .Q(n14279) );
  INVX0 U14795 ( .INP(n14284), .ZN(n14283) );
  OR2X1 U14796 ( .IN1(n14285), .IN2(n8105), .Q(n14284) );
  AND2X1 U14797 ( .IN1(n8105), .IN2(n14285), .Q(n14282) );
  INVX0 U14798 ( .INP(n14286), .ZN(n14285) );
  OR2X1 U14799 ( .IN1(n14287), .IN2(n14288), .Q(n14286) );
  AND2X1 U14800 ( .IN1(n8934), .IN2(n8662), .Q(n14288) );
  AND2X1 U14801 ( .IN1(n15967), .IN2(WX2144), .Q(n14287) );
  AND2X1 U14802 ( .IN1(n9235), .IN2(CRC_OUT_8_24), .Q(n14258) );
  AND2X1 U14803 ( .IN1(n273), .IN2(n9209), .Q(n14257) );
  INVX0 U14804 ( .INP(n14289), .ZN(n273) );
  OR2X1 U14805 ( .IN1(n9560), .IN2(n4027), .Q(n14289) );
  OR4X1 U14806 ( .IN1(n14290), .IN2(n14291), .IN3(n14292), .IN4(n14293), .Q(
        WX1949) );
  AND2X1 U14807 ( .IN1(n9269), .IN2(n13377), .Q(n14293) );
  OR2X1 U14808 ( .IN1(n14294), .IN2(n14295), .Q(n13377) );
  INVX0 U14809 ( .INP(n14296), .ZN(n14295) );
  OR2X1 U14810 ( .IN1(n14297), .IN2(n14298), .Q(n14296) );
  AND2X1 U14811 ( .IN1(n14298), .IN2(n14297), .Q(n14294) );
  AND2X1 U14812 ( .IN1(n14299), .IN2(n14300), .Q(n14297) );
  OR2X1 U14813 ( .IN1(n9464), .IN2(n8079), .Q(n14300) );
  OR2X1 U14814 ( .IN1(WX3307), .IN2(n9443), .Q(n14299) );
  OR2X1 U14815 ( .IN1(n14301), .IN2(n14302), .Q(n14298) );
  INVX0 U14816 ( .INP(n14303), .ZN(n14302) );
  OR2X1 U14817 ( .IN1(n14304), .IN2(n8080), .Q(n14303) );
  AND2X1 U14818 ( .IN1(n8080), .IN2(n14304), .Q(n14301) );
  INVX0 U14819 ( .INP(n14305), .ZN(n14304) );
  OR2X1 U14820 ( .IN1(n14306), .IN2(n14307), .Q(n14305) );
  AND2X1 U14821 ( .IN1(n8908), .IN2(n8605), .Q(n14307) );
  AND2X1 U14822 ( .IN1(n15970), .IN2(WX3435), .Q(n14306) );
  AND2X1 U14823 ( .IN1(n9188), .IN2(n11506), .Q(n14292) );
  OR2X1 U14824 ( .IN1(n14308), .IN2(n14309), .Q(n11506) );
  INVX0 U14825 ( .INP(n14310), .ZN(n14309) );
  OR2X1 U14826 ( .IN1(n14311), .IN2(n14312), .Q(n14310) );
  AND2X1 U14827 ( .IN1(n14312), .IN2(n14311), .Q(n14308) );
  AND2X1 U14828 ( .IN1(n14313), .IN2(n14314), .Q(n14311) );
  OR2X1 U14829 ( .IN1(n9467), .IN2(n8106), .Q(n14314) );
  OR2X1 U14830 ( .IN1(WX2014), .IN2(n9443), .Q(n14313) );
  OR2X1 U14831 ( .IN1(n14315), .IN2(n14316), .Q(n14312) );
  INVX0 U14832 ( .INP(n14317), .ZN(n14316) );
  OR2X1 U14833 ( .IN1(n14318), .IN2(n8107), .Q(n14317) );
  AND2X1 U14834 ( .IN1(n8107), .IN2(n14318), .Q(n14315) );
  INVX0 U14835 ( .INP(n14319), .ZN(n14318) );
  OR2X1 U14836 ( .IN1(n14320), .IN2(n14321), .Q(n14319) );
  AND2X1 U14837 ( .IN1(n8933), .IN2(n8663), .Q(n14321) );
  AND2X1 U14838 ( .IN1(n15969), .IN2(WX2142), .Q(n14320) );
  AND2X1 U14839 ( .IN1(test_so21), .IN2(n9228), .Q(n14291) );
  AND2X1 U14840 ( .IN1(n272), .IN2(n9209), .Q(n14290) );
  INVX0 U14841 ( .INP(n14322), .ZN(n272) );
  OR2X1 U14842 ( .IN1(n9560), .IN2(n4028), .Q(n14322) );
  OR4X1 U14843 ( .IN1(n14323), .IN2(n14324), .IN3(n14325), .IN4(n14326), .Q(
        WX1947) );
  AND2X1 U14844 ( .IN1(n13397), .IN2(n9260), .Q(n14326) );
  AND2X1 U14845 ( .IN1(n14327), .IN2(n14328), .Q(n13397) );
  INVX0 U14846 ( .INP(n14329), .ZN(n14328) );
  AND2X1 U14847 ( .IN1(n14330), .IN2(n14331), .Q(n14329) );
  OR2X1 U14848 ( .IN1(n14331), .IN2(n14330), .Q(n14327) );
  OR2X1 U14849 ( .IN1(n14332), .IN2(n14333), .Q(n14330) );
  AND2X1 U14850 ( .IN1(n9451), .IN2(WX3305), .Q(n14333) );
  AND2X1 U14851 ( .IN1(n8081), .IN2(n9470), .Q(n14332) );
  AND2X1 U14852 ( .IN1(n14334), .IN2(n14335), .Q(n14331) );
  OR2X1 U14853 ( .IN1(n14336), .IN2(n8907), .Q(n14335) );
  OR2X1 U14854 ( .IN1(WX3433), .IN2(n14337), .Q(n14334) );
  INVX0 U14855 ( .INP(n14336), .ZN(n14337) );
  AND2X1 U14856 ( .IN1(n14338), .IN2(n14339), .Q(n14336) );
  OR2X1 U14857 ( .IN1(n8606), .IN2(test_so27), .Q(n14339) );
  OR2X1 U14858 ( .IN1(n9140), .IN2(n15972), .Q(n14338) );
  AND2X1 U14859 ( .IN1(n9187), .IN2(n11512), .Q(n14325) );
  OR2X1 U14860 ( .IN1(n14340), .IN2(n14341), .Q(n11512) );
  INVX0 U14861 ( .INP(n14342), .ZN(n14341) );
  OR2X1 U14862 ( .IN1(n14343), .IN2(n14344), .Q(n14342) );
  AND2X1 U14863 ( .IN1(n14344), .IN2(n14343), .Q(n14340) );
  AND2X1 U14864 ( .IN1(n14345), .IN2(n14346), .Q(n14343) );
  OR2X1 U14865 ( .IN1(n9468), .IN2(n8108), .Q(n14346) );
  OR2X1 U14866 ( .IN1(WX2012), .IN2(n9443), .Q(n14345) );
  OR2X1 U14867 ( .IN1(n14347), .IN2(n14348), .Q(n14344) );
  INVX0 U14868 ( .INP(n14349), .ZN(n14348) );
  OR2X1 U14869 ( .IN1(n14350), .IN2(n8109), .Q(n14349) );
  AND2X1 U14870 ( .IN1(n8109), .IN2(n14350), .Q(n14347) );
  INVX0 U14871 ( .INP(n14351), .ZN(n14350) );
  OR2X1 U14872 ( .IN1(n14352), .IN2(n14353), .Q(n14351) );
  AND2X1 U14873 ( .IN1(n8932), .IN2(n8664), .Q(n14353) );
  AND2X1 U14874 ( .IN1(n15971), .IN2(WX2140), .Q(n14352) );
  AND2X1 U14875 ( .IN1(n9235), .IN2(CRC_OUT_8_26), .Q(n14324) );
  AND2X1 U14876 ( .IN1(n271), .IN2(n9209), .Q(n14323) );
  INVX0 U14877 ( .INP(n14354), .ZN(n271) );
  OR2X1 U14878 ( .IN1(n9559), .IN2(n4029), .Q(n14354) );
  OR4X1 U14879 ( .IN1(n14355), .IN2(n14356), .IN3(n14357), .IN4(n14358), .Q(
        WX1945) );
  AND2X1 U14880 ( .IN1(n9265), .IN2(n13417), .Q(n14358) );
  OR2X1 U14881 ( .IN1(n14359), .IN2(n14360), .Q(n13417) );
  INVX0 U14882 ( .INP(n14361), .ZN(n14360) );
  OR2X1 U14883 ( .IN1(n14362), .IN2(n14363), .Q(n14361) );
  AND2X1 U14884 ( .IN1(n14363), .IN2(n14362), .Q(n14359) );
  AND2X1 U14885 ( .IN1(n14364), .IN2(n14365), .Q(n14362) );
  OR2X1 U14886 ( .IN1(n9469), .IN2(n8082), .Q(n14365) );
  OR2X1 U14887 ( .IN1(WX3303), .IN2(n9443), .Q(n14364) );
  OR2X1 U14888 ( .IN1(n14366), .IN2(n14367), .Q(n14363) );
  INVX0 U14889 ( .INP(n14368), .ZN(n14367) );
  OR2X1 U14890 ( .IN1(n14369), .IN2(n8083), .Q(n14368) );
  AND2X1 U14891 ( .IN1(n8083), .IN2(n14369), .Q(n14366) );
  INVX0 U14892 ( .INP(n14370), .ZN(n14369) );
  OR2X1 U14893 ( .IN1(n14371), .IN2(n14372), .Q(n14370) );
  AND2X1 U14894 ( .IN1(n8906), .IN2(n8607), .Q(n14372) );
  AND2X1 U14895 ( .IN1(n15974), .IN2(WX3431), .Q(n14371) );
  AND2X1 U14896 ( .IN1(n9187), .IN2(n11518), .Q(n14357) );
  OR2X1 U14897 ( .IN1(n14373), .IN2(n14374), .Q(n11518) );
  INVX0 U14898 ( .INP(n14375), .ZN(n14374) );
  OR2X1 U14899 ( .IN1(n14376), .IN2(n14377), .Q(n14375) );
  AND2X1 U14900 ( .IN1(n14377), .IN2(n14376), .Q(n14373) );
  AND2X1 U14901 ( .IN1(n14378), .IN2(n14379), .Q(n14376) );
  OR2X1 U14902 ( .IN1(n9469), .IN2(n8110), .Q(n14379) );
  OR2X1 U14903 ( .IN1(WX2010), .IN2(n9443), .Q(n14378) );
  OR2X1 U14904 ( .IN1(n14380), .IN2(n14381), .Q(n14377) );
  INVX0 U14905 ( .INP(n14382), .ZN(n14381) );
  OR2X1 U14906 ( .IN1(n14383), .IN2(n8111), .Q(n14382) );
  AND2X1 U14907 ( .IN1(n8111), .IN2(n14383), .Q(n14380) );
  INVX0 U14908 ( .INP(n14384), .ZN(n14383) );
  OR2X1 U14909 ( .IN1(n14385), .IN2(n14386), .Q(n14384) );
  AND2X1 U14910 ( .IN1(n8931), .IN2(n8665), .Q(n14386) );
  AND2X1 U14911 ( .IN1(n15973), .IN2(WX2138), .Q(n14385) );
  AND2X1 U14912 ( .IN1(n9235), .IN2(CRC_OUT_8_27), .Q(n14356) );
  AND2X1 U14913 ( .IN1(n270), .IN2(n9209), .Q(n14355) );
  INVX0 U14914 ( .INP(n14387), .ZN(n270) );
  OR2X1 U14915 ( .IN1(n9559), .IN2(n4030), .Q(n14387) );
  OR4X1 U14916 ( .IN1(n14388), .IN2(n14389), .IN3(n14390), .IN4(n14391), .Q(
        WX1943) );
  AND2X1 U14917 ( .IN1(n9270), .IN2(n13437), .Q(n14391) );
  OR2X1 U14918 ( .IN1(n14392), .IN2(n14393), .Q(n13437) );
  AND2X1 U14919 ( .IN1(n14394), .IN2(n14395), .Q(n14393) );
  INVX0 U14920 ( .INP(n14396), .ZN(n14395) );
  AND2X1 U14921 ( .IN1(n14396), .IN2(n14397), .Q(n14392) );
  INVX0 U14922 ( .INP(n14394), .ZN(n14397) );
  OR2X1 U14923 ( .IN1(n14398), .IN2(n14399), .Q(n14394) );
  AND2X1 U14924 ( .IN1(n9450), .IN2(n8608), .Q(n14399) );
  AND2X1 U14925 ( .IN1(n15976), .IN2(n9458), .Q(n14398) );
  OR2X1 U14926 ( .IN1(n14400), .IN2(n14401), .Q(n14396) );
  AND3X1 U14927 ( .IN1(n14402), .IN2(n14403), .IN3(n8905), .Q(n14401) );
  OR2X1 U14928 ( .IN1(n8084), .IN2(WX3365), .Q(n14403) );
  OR2X1 U14929 ( .IN1(n8085), .IN2(WX3301), .Q(n14402) );
  AND2X1 U14930 ( .IN1(n14404), .IN2(WX3429), .Q(n14400) );
  OR2X1 U14931 ( .IN1(n14405), .IN2(n14406), .Q(n14404) );
  AND2X1 U14932 ( .IN1(n8084), .IN2(WX3365), .Q(n14406) );
  AND2X1 U14933 ( .IN1(n8085), .IN2(WX3301), .Q(n14405) );
  AND2X1 U14934 ( .IN1(n11524), .IN2(n9175), .Q(n14390) );
  AND2X1 U14935 ( .IN1(n14407), .IN2(n14408), .Q(n11524) );
  INVX0 U14936 ( .INP(n14409), .ZN(n14408) );
  AND2X1 U14937 ( .IN1(n14410), .IN2(n14411), .Q(n14409) );
  OR2X1 U14938 ( .IN1(n14411), .IN2(n14410), .Q(n14407) );
  OR2X1 U14939 ( .IN1(n14412), .IN2(n14413), .Q(n14410) );
  AND2X1 U14940 ( .IN1(n9450), .IN2(WX2008), .Q(n14413) );
  AND2X1 U14941 ( .IN1(n8112), .IN2(n9472), .Q(n14412) );
  AND2X1 U14942 ( .IN1(n14414), .IN2(n14415), .Q(n14411) );
  OR2X1 U14943 ( .IN1(n14416), .IN2(n8113), .Q(n14415) );
  INVX0 U14944 ( .INP(n14417), .ZN(n14416) );
  OR2X1 U14945 ( .IN1(WX2072), .IN2(n14417), .Q(n14414) );
  OR2X1 U14946 ( .IN1(n14418), .IN2(n14419), .Q(n14417) );
  AND2X1 U14947 ( .IN1(n15975), .IN2(n9108), .Q(n14419) );
  AND2X1 U14948 ( .IN1(test_so18), .IN2(n8666), .Q(n14418) );
  AND2X1 U14949 ( .IN1(n9235), .IN2(CRC_OUT_8_28), .Q(n14389) );
  AND2X1 U14950 ( .IN1(n269), .IN2(n9209), .Q(n14388) );
  INVX0 U14951 ( .INP(n14420), .ZN(n269) );
  OR2X1 U14952 ( .IN1(n9559), .IN2(n4031), .Q(n14420) );
  OR4X1 U14953 ( .IN1(n14421), .IN2(n14422), .IN3(n14423), .IN4(n14424), .Q(
        WX1941) );
  AND2X1 U14954 ( .IN1(n9269), .IN2(n13456), .Q(n14424) );
  OR2X1 U14955 ( .IN1(n14425), .IN2(n14426), .Q(n13456) );
  INVX0 U14956 ( .INP(n14427), .ZN(n14426) );
  OR2X1 U14957 ( .IN1(n14428), .IN2(n14429), .Q(n14427) );
  AND2X1 U14958 ( .IN1(n14429), .IN2(n14428), .Q(n14425) );
  AND2X1 U14959 ( .IN1(n14430), .IN2(n14431), .Q(n14428) );
  OR2X1 U14960 ( .IN1(n9471), .IN2(n8086), .Q(n14431) );
  OR2X1 U14961 ( .IN1(WX3299), .IN2(n9443), .Q(n14430) );
  OR2X1 U14962 ( .IN1(n14432), .IN2(n14433), .Q(n14429) );
  INVX0 U14963 ( .INP(n14434), .ZN(n14433) );
  OR2X1 U14964 ( .IN1(n14435), .IN2(n8087), .Q(n14434) );
  AND2X1 U14965 ( .IN1(n8087), .IN2(n14435), .Q(n14432) );
  INVX0 U14966 ( .INP(n14436), .ZN(n14435) );
  OR2X1 U14967 ( .IN1(n14437), .IN2(n14438), .Q(n14436) );
  AND2X1 U14968 ( .IN1(n8904), .IN2(n8609), .Q(n14438) );
  AND2X1 U14969 ( .IN1(n15978), .IN2(WX3427), .Q(n14437) );
  AND2X1 U14970 ( .IN1(n9187), .IN2(n11550), .Q(n14423) );
  OR2X1 U14971 ( .IN1(n14439), .IN2(n14440), .Q(n11550) );
  INVX0 U14972 ( .INP(n14441), .ZN(n14440) );
  OR2X1 U14973 ( .IN1(n14442), .IN2(n14443), .Q(n14441) );
  AND2X1 U14974 ( .IN1(n14443), .IN2(n14442), .Q(n14439) );
  AND2X1 U14975 ( .IN1(n14444), .IN2(n14445), .Q(n14442) );
  OR2X1 U14976 ( .IN1(n9471), .IN2(n8114), .Q(n14445) );
  OR2X1 U14977 ( .IN1(WX2006), .IN2(n9443), .Q(n14444) );
  OR2X1 U14978 ( .IN1(n14446), .IN2(n14447), .Q(n14443) );
  INVX0 U14979 ( .INP(n14448), .ZN(n14447) );
  OR2X1 U14980 ( .IN1(n14449), .IN2(n8115), .Q(n14448) );
  AND2X1 U14981 ( .IN1(n8115), .IN2(n14449), .Q(n14446) );
  INVX0 U14982 ( .INP(n14450), .ZN(n14449) );
  OR2X1 U14983 ( .IN1(n14451), .IN2(n14452), .Q(n14450) );
  AND2X1 U14984 ( .IN1(n8930), .IN2(n8667), .Q(n14452) );
  AND2X1 U14985 ( .IN1(n15977), .IN2(WX2134), .Q(n14451) );
  AND2X1 U14986 ( .IN1(n9236), .IN2(CRC_OUT_8_29), .Q(n14422) );
  AND2X1 U14987 ( .IN1(n268), .IN2(n9210), .Q(n14421) );
  INVX0 U14988 ( .INP(n14453), .ZN(n268) );
  OR2X1 U14989 ( .IN1(n9559), .IN2(n4032), .Q(n14453) );
  OR4X1 U14990 ( .IN1(n14454), .IN2(n14455), .IN3(n14456), .IN4(n14457), .Q(
        WX1939) );
  AND2X1 U14991 ( .IN1(n13476), .IN2(n9261), .Q(n14457) );
  AND2X1 U14992 ( .IN1(n14458), .IN2(n14459), .Q(n13476) );
  INVX0 U14993 ( .INP(n14460), .ZN(n14459) );
  AND2X1 U14994 ( .IN1(n14461), .IN2(n14462), .Q(n14460) );
  OR2X1 U14995 ( .IN1(n14462), .IN2(n14461), .Q(n14458) );
  OR2X1 U14996 ( .IN1(n14463), .IN2(n14464), .Q(n14461) );
  AND2X1 U14997 ( .IN1(n9450), .IN2(WX3361), .Q(n14464) );
  AND2X1 U14998 ( .IN1(n8088), .IN2(n9473), .Q(n14463) );
  AND2X1 U14999 ( .IN1(n14465), .IN2(n14466), .Q(n14462) );
  OR2X1 U15000 ( .IN1(n14467), .IN2(n8903), .Q(n14466) );
  OR2X1 U15001 ( .IN1(WX3425), .IN2(n14468), .Q(n14465) );
  INVX0 U15002 ( .INP(n14467), .ZN(n14468) );
  AND2X1 U15003 ( .IN1(n14469), .IN2(n14470), .Q(n14467) );
  OR2X1 U15004 ( .IN1(n8610), .IN2(test_so25), .Q(n14470) );
  OR2X1 U15005 ( .IN1(n9141), .IN2(n15980), .Q(n14469) );
  AND2X1 U15006 ( .IN1(n9187), .IN2(n11582), .Q(n14456) );
  OR2X1 U15007 ( .IN1(n14471), .IN2(n14472), .Q(n11582) );
  INVX0 U15008 ( .INP(n14473), .ZN(n14472) );
  OR2X1 U15009 ( .IN1(n14474), .IN2(n14475), .Q(n14473) );
  AND2X1 U15010 ( .IN1(n14475), .IN2(n14474), .Q(n14471) );
  AND2X1 U15011 ( .IN1(n14476), .IN2(n14477), .Q(n14474) );
  OR2X1 U15012 ( .IN1(n9472), .IN2(n8116), .Q(n14477) );
  OR2X1 U15013 ( .IN1(WX2004), .IN2(n9443), .Q(n14476) );
  OR2X1 U15014 ( .IN1(n14478), .IN2(n14479), .Q(n14475) );
  INVX0 U15015 ( .INP(n14480), .ZN(n14479) );
  OR2X1 U15016 ( .IN1(n14481), .IN2(n8117), .Q(n14480) );
  AND2X1 U15017 ( .IN1(n8117), .IN2(n14481), .Q(n14478) );
  INVX0 U15018 ( .INP(n14482), .ZN(n14481) );
  OR2X1 U15019 ( .IN1(n14483), .IN2(n14484), .Q(n14482) );
  AND2X1 U15020 ( .IN1(n8929), .IN2(n8668), .Q(n14484) );
  AND2X1 U15021 ( .IN1(n15979), .IN2(WX2132), .Q(n14483) );
  AND2X1 U15022 ( .IN1(n9236), .IN2(CRC_OUT_8_30), .Q(n14455) );
  AND2X1 U15023 ( .IN1(n267), .IN2(n9210), .Q(n14454) );
  INVX0 U15024 ( .INP(n14485), .ZN(n267) );
  OR2X1 U15025 ( .IN1(n9559), .IN2(n4033), .Q(n14485) );
  OR4X1 U15026 ( .IN1(n14486), .IN2(n14487), .IN3(n14488), .IN4(n14489), .Q(
        WX1937) );
  AND2X1 U15027 ( .IN1(n9187), .IN2(n11618), .Q(n14489) );
  OR2X1 U15028 ( .IN1(n14490), .IN2(n14491), .Q(n11618) );
  INVX0 U15029 ( .INP(n14492), .ZN(n14491) );
  OR2X1 U15030 ( .IN1(n14493), .IN2(n14494), .Q(n14492) );
  AND2X1 U15031 ( .IN1(n14494), .IN2(n14493), .Q(n14490) );
  AND2X1 U15032 ( .IN1(n14495), .IN2(n14496), .Q(n14493) );
  OR2X1 U15033 ( .IN1(n9473), .IN2(n7890), .Q(n14496) );
  OR2X1 U15034 ( .IN1(WX2002), .IN2(n9443), .Q(n14495) );
  OR2X1 U15035 ( .IN1(n14497), .IN2(n14498), .Q(n14494) );
  INVX0 U15036 ( .INP(n14499), .ZN(n14498) );
  OR2X1 U15037 ( .IN1(n14500), .IN2(n7891), .Q(n14499) );
  AND2X1 U15038 ( .IN1(n7891), .IN2(n14500), .Q(n14497) );
  INVX0 U15039 ( .INP(n14501), .ZN(n14500) );
  OR2X1 U15040 ( .IN1(n14502), .IN2(n14503), .Q(n14501) );
  AND2X1 U15041 ( .IN1(n8928), .IN2(n8669), .Q(n14503) );
  AND2X1 U15042 ( .IN1(n15982), .IN2(WX2130), .Q(n14502) );
  AND2X1 U15043 ( .IN1(n9269), .IN2(n13495), .Q(n14488) );
  OR2X1 U15044 ( .IN1(n14504), .IN2(n14505), .Q(n13495) );
  INVX0 U15045 ( .INP(n14506), .ZN(n14505) );
  OR2X1 U15046 ( .IN1(n14507), .IN2(n14508), .Q(n14506) );
  AND2X1 U15047 ( .IN1(n14508), .IN2(n14507), .Q(n14504) );
  AND2X1 U15048 ( .IN1(n14509), .IN2(n14510), .Q(n14507) );
  OR2X1 U15049 ( .IN1(n9473), .IN2(n7888), .Q(n14510) );
  OR2X1 U15050 ( .IN1(WX3295), .IN2(n9443), .Q(n14509) );
  OR2X1 U15051 ( .IN1(n14511), .IN2(n14512), .Q(n14508) );
  INVX0 U15052 ( .INP(n14513), .ZN(n14512) );
  OR2X1 U15053 ( .IN1(n14514), .IN2(n7889), .Q(n14513) );
  AND2X1 U15054 ( .IN1(n7889), .IN2(n14514), .Q(n14511) );
  INVX0 U15055 ( .INP(n14515), .ZN(n14514) );
  OR2X1 U15056 ( .IN1(n14516), .IN2(n14517), .Q(n14515) );
  AND2X1 U15057 ( .IN1(n8902), .IN2(n8611), .Q(n14517) );
  AND2X1 U15058 ( .IN1(n15981), .IN2(WX3423), .Q(n14516) );
  AND2X1 U15059 ( .IN1(n2245), .IN2(WX1778), .Q(n14487) );
  AND2X1 U15060 ( .IN1(n9236), .IN2(CRC_OUT_8_31), .Q(n14486) );
  AND2X1 U15061 ( .IN1(n9045), .IN2(n9499), .Q(WX1839) );
  AND3X1 U15062 ( .IN1(n14518), .IN2(n14519), .IN3(n9524), .Q(WX1326) );
  OR2X1 U15063 ( .IN1(DFF_190_n1), .IN2(WX837), .Q(n14519) );
  OR2X1 U15064 ( .IN1(n9030), .IN2(CRC_OUT_9_30), .Q(n14518) );
  AND3X1 U15065 ( .IN1(n14520), .IN2(n14521), .IN3(n9524), .Q(WX1324) );
  OR2X1 U15066 ( .IN1(DFF_189_n1), .IN2(WX839), .Q(n14521) );
  OR2X1 U15067 ( .IN1(n8956), .IN2(CRC_OUT_9_29), .Q(n14520) );
  AND3X1 U15068 ( .IN1(n14522), .IN2(n14523), .IN3(n9524), .Q(WX1322) );
  OR2X1 U15069 ( .IN1(DFF_188_n1), .IN2(WX841), .Q(n14523) );
  OR2X1 U15070 ( .IN1(n8964), .IN2(CRC_OUT_9_28), .Q(n14522) );
  AND3X1 U15071 ( .IN1(n14524), .IN2(n14525), .IN3(n9523), .Q(WX1320) );
  OR2X1 U15072 ( .IN1(DFF_187_n1), .IN2(WX843), .Q(n14525) );
  OR2X1 U15073 ( .IN1(n8973), .IN2(CRC_OUT_9_27), .Q(n14524) );
  AND3X1 U15074 ( .IN1(n14526), .IN2(n14527), .IN3(n9523), .Q(WX1318) );
  OR2X1 U15075 ( .IN1(DFF_186_n1), .IN2(WX845), .Q(n14527) );
  OR2X1 U15076 ( .IN1(n8979), .IN2(CRC_OUT_9_26), .Q(n14526) );
  AND3X1 U15077 ( .IN1(n14528), .IN2(n14529), .IN3(n9523), .Q(WX1316) );
  OR2X1 U15078 ( .IN1(DFF_185_n1), .IN2(WX847), .Q(n14529) );
  OR2X1 U15079 ( .IN1(n8982), .IN2(CRC_OUT_9_25), .Q(n14528) );
  AND3X1 U15080 ( .IN1(n14530), .IN2(n14531), .IN3(n9523), .Q(WX1314) );
  OR2X1 U15081 ( .IN1(DFF_184_n1), .IN2(WX849), .Q(n14531) );
  OR2X1 U15082 ( .IN1(n8991), .IN2(CRC_OUT_9_24), .Q(n14530) );
  AND3X1 U15083 ( .IN1(n14532), .IN2(n14533), .IN3(n9523), .Q(WX1312) );
  OR2X1 U15084 ( .IN1(DFF_183_n1), .IN2(WX851), .Q(n14533) );
  OR2X1 U15085 ( .IN1(n9000), .IN2(CRC_OUT_9_23), .Q(n14532) );
  AND3X1 U15086 ( .IN1(n14534), .IN2(n14535), .IN3(n9523), .Q(WX1310) );
  OR2X1 U15087 ( .IN1(DFF_182_n1), .IN2(WX853), .Q(n14535) );
  OR2X1 U15088 ( .IN1(n9002), .IN2(CRC_OUT_9_22), .Q(n14534) );
  AND3X1 U15089 ( .IN1(n14536), .IN2(n14537), .IN3(n9523), .Q(WX1308) );
  OR2X1 U15090 ( .IN1(DFF_181_n1), .IN2(WX855), .Q(n14537) );
  OR2X1 U15091 ( .IN1(n9017), .IN2(CRC_OUT_9_21), .Q(n14536) );
  AND3X1 U15092 ( .IN1(n14538), .IN2(n14539), .IN3(n9523), .Q(WX1306) );
  OR2X1 U15093 ( .IN1(DFF_180_n1), .IN2(WX857), .Q(n14539) );
  OR2X1 U15094 ( .IN1(n9023), .IN2(CRC_OUT_9_20), .Q(n14538) );
  AND2X1 U15095 ( .IN1(n14540), .IN2(n9499), .Q(WX1304) );
  OR2X1 U15096 ( .IN1(n14541), .IN2(n14542), .Q(n14540) );
  AND2X1 U15097 ( .IN1(n9026), .IN2(n9161), .Q(n14542) );
  AND2X1 U15098 ( .IN1(test_so10), .IN2(WX859), .Q(n14541) );
  AND3X1 U15099 ( .IN1(n14543), .IN2(n14544), .IN3(n9523), .Q(WX1302) );
  OR2X1 U15100 ( .IN1(DFF_178_n1), .IN2(WX861), .Q(n14544) );
  OR2X1 U15101 ( .IN1(n8961), .IN2(CRC_OUT_9_18), .Q(n14543) );
  AND3X1 U15102 ( .IN1(n14545), .IN2(n14546), .IN3(n9523), .Q(WX1300) );
  OR2X1 U15103 ( .IN1(DFF_177_n1), .IN2(WX863), .Q(n14546) );
  OR2X1 U15104 ( .IN1(n8976), .IN2(CRC_OUT_9_17), .Q(n14545) );
  AND3X1 U15105 ( .IN1(n14547), .IN2(n14548), .IN3(n9523), .Q(WX1298) );
  OR2X1 U15106 ( .IN1(DFF_176_n1), .IN2(WX865), .Q(n14548) );
  OR2X1 U15107 ( .IN1(n8988), .IN2(CRC_OUT_9_16), .Q(n14547) );
  AND3X1 U15108 ( .IN1(n14549), .IN2(n14550), .IN3(n9523), .Q(WX1296) );
  OR2X1 U15109 ( .IN1(DFF_175_n1), .IN2(n14551), .Q(n14550) );
  AND2X1 U15110 ( .IN1(n14552), .IN2(n14553), .Q(n14551) );
  OR2X1 U15111 ( .IN1(DFF_191_n1), .IN2(n9086), .Q(n14553) );
  OR2X1 U15112 ( .IN1(test_so8), .IN2(CRC_OUT_9_31), .Q(n14552) );
  OR3X1 U15113 ( .IN1(n14554), .IN2(n14555), .IN3(CRC_OUT_9_15), .Q(n14549) );
  AND2X1 U15114 ( .IN1(DFF_191_n1), .IN2(n9086), .Q(n14555) );
  AND2X1 U15115 ( .IN1(test_so8), .IN2(CRC_OUT_9_31), .Q(n14554) );
  AND3X1 U15116 ( .IN1(n14556), .IN2(n14557), .IN3(n9522), .Q(WX1294) );
  OR2X1 U15117 ( .IN1(DFF_174_n1), .IN2(WX869), .Q(n14557) );
  OR2X1 U15118 ( .IN1(n9020), .IN2(CRC_OUT_9_14), .Q(n14556) );
  AND3X1 U15119 ( .IN1(n14558), .IN2(n14559), .IN3(n9522), .Q(WX1292) );
  OR2X1 U15120 ( .IN1(DFF_173_n1), .IN2(WX871), .Q(n14559) );
  OR2X1 U15121 ( .IN1(n9032), .IN2(CRC_OUT_9_13), .Q(n14558) );
  AND3X1 U15122 ( .IN1(n14560), .IN2(n14561), .IN3(n9522), .Q(WX1290) );
  OR2X1 U15123 ( .IN1(DFF_172_n1), .IN2(WX873), .Q(n14561) );
  OR2X1 U15124 ( .IN1(n8967), .IN2(CRC_OUT_9_12), .Q(n14560) );
  AND3X1 U15125 ( .IN1(n14562), .IN2(n14563), .IN3(n9522), .Q(WX1288) );
  OR2X1 U15126 ( .IN1(DFF_171_n1), .IN2(WX875), .Q(n14563) );
  OR2X1 U15127 ( .IN1(n8994), .IN2(CRC_OUT_9_11), .Q(n14562) );
  AND2X1 U15128 ( .IN1(n14564), .IN2(n9498), .Q(WX1286) );
  OR2X1 U15129 ( .IN1(n14565), .IN2(n14566), .Q(n14564) );
  AND2X1 U15130 ( .IN1(n14567), .IN2(CRC_OUT_9_10), .Q(n14566) );
  AND2X1 U15131 ( .IN1(DFF_170_n1), .IN2(n14568), .Q(n14565) );
  INVX0 U15132 ( .INP(n14567), .ZN(n14568) );
  OR2X1 U15133 ( .IN1(n14569), .IN2(n14570), .Q(n14567) );
  AND2X1 U15134 ( .IN1(DFF_191_n1), .IN2(WX877), .Q(n14570) );
  AND2X1 U15135 ( .IN1(n9040), .IN2(CRC_OUT_9_31), .Q(n14569) );
  AND3X1 U15136 ( .IN1(n14571), .IN2(n14572), .IN3(n9522), .Q(WX1284) );
  OR2X1 U15137 ( .IN1(DFF_169_n1), .IN2(WX879), .Q(n14572) );
  OR2X1 U15138 ( .IN1(n8985), .IN2(CRC_OUT_9_9), .Q(n14571) );
  AND3X1 U15139 ( .IN1(n14573), .IN2(n14574), .IN3(n9522), .Q(WX1282) );
  OR2X1 U15140 ( .IN1(DFF_168_n1), .IN2(WX881), .Q(n14574) );
  OR2X1 U15141 ( .IN1(n8998), .IN2(CRC_OUT_9_8), .Q(n14573) );
  AND3X1 U15142 ( .IN1(n14575), .IN2(n14576), .IN3(n9522), .Q(WX1280) );
  OR2X1 U15143 ( .IN1(DFF_167_n1), .IN2(WX883), .Q(n14576) );
  OR2X1 U15144 ( .IN1(n9007), .IN2(CRC_OUT_9_7), .Q(n14575) );
  AND3X1 U15145 ( .IN1(n14577), .IN2(n14578), .IN3(n9522), .Q(WX1278) );
  OR2X1 U15146 ( .IN1(DFF_166_n1), .IN2(WX885), .Q(n14578) );
  OR2X1 U15147 ( .IN1(n9038), .IN2(CRC_OUT_9_6), .Q(n14577) );
  AND3X1 U15148 ( .IN1(n14579), .IN2(n14580), .IN3(n9522), .Q(WX1276) );
  OR2X1 U15149 ( .IN1(DFF_165_n1), .IN2(WX887), .Q(n14580) );
  OR2X1 U15150 ( .IN1(n9025), .IN2(CRC_OUT_9_5), .Q(n14579) );
  AND3X1 U15151 ( .IN1(n14581), .IN2(n14582), .IN3(n9522), .Q(WX1274) );
  OR2X1 U15152 ( .IN1(DFF_164_n1), .IN2(WX889), .Q(n14582) );
  OR2X1 U15153 ( .IN1(n9010), .IN2(CRC_OUT_9_4), .Q(n14581) );
  AND2X1 U15154 ( .IN1(n14583), .IN2(n9499), .Q(WX1272) );
  OR2X1 U15155 ( .IN1(n14584), .IN2(n14585), .Q(n14583) );
  AND2X1 U15156 ( .IN1(n14586), .IN2(CRC_OUT_9_3), .Q(n14585) );
  AND2X1 U15157 ( .IN1(DFF_163_n1), .IN2(n14587), .Q(n14584) );
  INVX0 U15158 ( .INP(n14586), .ZN(n14587) );
  OR2X1 U15159 ( .IN1(n14588), .IN2(n14589), .Q(n14586) );
  AND2X1 U15160 ( .IN1(DFF_191_n1), .IN2(WX891), .Q(n14589) );
  AND2X1 U15161 ( .IN1(n9013), .IN2(CRC_OUT_9_31), .Q(n14588) );
  AND3X1 U15162 ( .IN1(n14590), .IN2(n14591), .IN3(n9522), .Q(WX1270) );
  OR2X1 U15163 ( .IN1(DFF_162_n1), .IN2(WX893), .Q(n14591) );
  OR2X1 U15164 ( .IN1(n8958), .IN2(CRC_OUT_9_2), .Q(n14590) );
  AND2X1 U15165 ( .IN1(n14592), .IN2(n9499), .Q(WX1268) );
  OR2X1 U15166 ( .IN1(n14593), .IN2(n14594), .Q(n14592) );
  AND2X1 U15167 ( .IN1(n9035), .IN2(n9162), .Q(n14594) );
  AND2X1 U15168 ( .IN1(test_so9), .IN2(WX895), .Q(n14593) );
  AND3X1 U15169 ( .IN1(n14595), .IN2(n14596), .IN3(n9522), .Q(WX1266) );
  OR2X1 U15170 ( .IN1(DFF_160_n1), .IN2(WX897), .Q(n14596) );
  OR2X1 U15171 ( .IN1(n8969), .IN2(CRC_OUT_9_0), .Q(n14595) );
  AND3X1 U15172 ( .IN1(n14597), .IN2(n14598), .IN3(n9521), .Q(WX1264) );
  OR2X1 U15173 ( .IN1(DFF_191_n1), .IN2(WX899), .Q(n14598) );
  OR2X1 U15174 ( .IN1(n9044), .IN2(CRC_OUT_9_31), .Q(n14597) );
  AND3X1 U15175 ( .IN1(n14599), .IN2(n14600), .IN3(n9521), .Q(WX11670) );
  OR2X1 U15176 ( .IN1(DFF_1726_n1), .IN2(WX11181), .Q(n14600) );
  OR2X1 U15177 ( .IN1(n8742), .IN2(CRC_OUT_1_30), .Q(n14599) );
  AND3X1 U15178 ( .IN1(n14601), .IN2(n14602), .IN3(n9521), .Q(WX11668) );
  OR2X1 U15179 ( .IN1(DFF_1725_n1), .IN2(WX11183), .Q(n14602) );
  OR2X1 U15180 ( .IN1(n8743), .IN2(CRC_OUT_1_29), .Q(n14601) );
  AND3X1 U15181 ( .IN1(n14603), .IN2(n14604), .IN3(n9521), .Q(WX11666) );
  OR2X1 U15182 ( .IN1(DFF_1724_n1), .IN2(WX11185), .Q(n14604) );
  OR2X1 U15183 ( .IN1(n8744), .IN2(CRC_OUT_1_28), .Q(n14603) );
  AND3X1 U15184 ( .IN1(n14605), .IN2(n14606), .IN3(n9521), .Q(WX11664) );
  OR2X1 U15185 ( .IN1(DFF_1723_n1), .IN2(WX11187), .Q(n14606) );
  OR2X1 U15186 ( .IN1(n8745), .IN2(CRC_OUT_1_27), .Q(n14605) );
  AND3X1 U15187 ( .IN1(n14607), .IN2(n14608), .IN3(n9521), .Q(WX11662) );
  OR2X1 U15188 ( .IN1(DFF_1722_n1), .IN2(WX11189), .Q(n14608) );
  OR2X1 U15189 ( .IN1(n8746), .IN2(CRC_OUT_1_26), .Q(n14607) );
  AND3X1 U15190 ( .IN1(n14609), .IN2(n14610), .IN3(n9521), .Q(WX11660) );
  OR2X1 U15191 ( .IN1(DFF_1721_n1), .IN2(WX11191), .Q(n14610) );
  OR2X1 U15192 ( .IN1(n8747), .IN2(CRC_OUT_1_25), .Q(n14609) );
  AND3X1 U15193 ( .IN1(n14611), .IN2(n14612), .IN3(n9521), .Q(WX11658) );
  OR2X1 U15194 ( .IN1(DFF_1720_n1), .IN2(WX11193), .Q(n14612) );
  OR2X1 U15195 ( .IN1(n8748), .IN2(CRC_OUT_1_24), .Q(n14611) );
  AND3X1 U15196 ( .IN1(n14613), .IN2(n14614), .IN3(n9521), .Q(WX11656) );
  OR2X1 U15197 ( .IN1(DFF_1719_n1), .IN2(WX11195), .Q(n14614) );
  OR2X1 U15198 ( .IN1(n8749), .IN2(CRC_OUT_1_23), .Q(n14613) );
  AND3X1 U15199 ( .IN1(n14615), .IN2(n14616), .IN3(n9521), .Q(WX11654) );
  OR2X1 U15200 ( .IN1(DFF_1718_n1), .IN2(WX11197), .Q(n14616) );
  OR2X1 U15201 ( .IN1(n8750), .IN2(CRC_OUT_1_22), .Q(n14615) );
  AND3X1 U15202 ( .IN1(n14617), .IN2(n14618), .IN3(n9521), .Q(WX11652) );
  OR2X1 U15203 ( .IN1(DFF_1717_n1), .IN2(WX11199), .Q(n14618) );
  OR2X1 U15204 ( .IN1(n8751), .IN2(CRC_OUT_1_21), .Q(n14617) );
  AND3X1 U15205 ( .IN1(n14619), .IN2(n14620), .IN3(n9521), .Q(WX11650) );
  OR2X1 U15206 ( .IN1(DFF_1716_n1), .IN2(WX11201), .Q(n14620) );
  OR2X1 U15207 ( .IN1(n8752), .IN2(CRC_OUT_1_20), .Q(n14619) );
  AND3X1 U15208 ( .IN1(n14621), .IN2(n14622), .IN3(n9520), .Q(WX11648) );
  OR2X1 U15209 ( .IN1(DFF_1715_n1), .IN2(WX11203), .Q(n14622) );
  OR2X1 U15210 ( .IN1(n8753), .IN2(CRC_OUT_1_19), .Q(n14621) );
  AND2X1 U15211 ( .IN1(n14623), .IN2(n9498), .Q(WX11646) );
  OR2X1 U15212 ( .IN1(n14624), .IN2(n14625), .Q(n14623) );
  AND2X1 U15213 ( .IN1(DFF_1714_n1), .IN2(n9109), .Q(n14625) );
  AND2X1 U15214 ( .IN1(test_so97), .IN2(CRC_OUT_1_18), .Q(n14624) );
  AND3X1 U15215 ( .IN1(n14626), .IN2(n14627), .IN3(n9520), .Q(WX11644) );
  OR2X1 U15216 ( .IN1(DFF_1713_n1), .IN2(WX11207), .Q(n14627) );
  OR2X1 U15217 ( .IN1(n8754), .IN2(CRC_OUT_1_17), .Q(n14626) );
  AND3X1 U15218 ( .IN1(n14628), .IN2(n14629), .IN3(n9520), .Q(WX11642) );
  OR2X1 U15219 ( .IN1(DFF_1712_n1), .IN2(WX11209), .Q(n14629) );
  OR2X1 U15220 ( .IN1(n8755), .IN2(CRC_OUT_1_16), .Q(n14628) );
  AND3X1 U15221 ( .IN1(n14630), .IN2(n14631), .IN3(n9520), .Q(WX11640) );
  OR2X1 U15222 ( .IN1(DFF_1711_n1), .IN2(n14632), .Q(n14631) );
  AND2X1 U15223 ( .IN1(n14633), .IN2(n14634), .Q(n14632) );
  OR2X1 U15224 ( .IN1(n8713), .IN2(n9085), .Q(n14634) );
  OR2X1 U15225 ( .IN1(test_so100), .IN2(WX11211), .Q(n14633) );
  OR3X1 U15226 ( .IN1(n14635), .IN2(n14636), .IN3(CRC_OUT_1_15), .Q(n14630) );
  AND2X1 U15227 ( .IN1(n8713), .IN2(n9085), .Q(n14636) );
  AND2X1 U15228 ( .IN1(test_so100), .IN2(WX11211), .Q(n14635) );
  AND2X1 U15229 ( .IN1(n14637), .IN2(n9498), .Q(WX11638) );
  OR2X1 U15230 ( .IN1(n14638), .IN2(n14639), .Q(n14637) );
  AND2X1 U15231 ( .IN1(n8756), .IN2(n9163), .Q(n14639) );
  AND2X1 U15232 ( .IN1(test_so99), .IN2(WX11213), .Q(n14638) );
  AND3X1 U15233 ( .IN1(n14640), .IN2(n14641), .IN3(n9520), .Q(WX11636) );
  OR2X1 U15234 ( .IN1(DFF_1709_n1), .IN2(WX11215), .Q(n14641) );
  OR2X1 U15235 ( .IN1(n8757), .IN2(CRC_OUT_1_13), .Q(n14640) );
  AND3X1 U15236 ( .IN1(n14642), .IN2(n14643), .IN3(n9520), .Q(WX11634) );
  OR2X1 U15237 ( .IN1(DFF_1708_n1), .IN2(WX11217), .Q(n14643) );
  OR2X1 U15238 ( .IN1(n8758), .IN2(CRC_OUT_1_12), .Q(n14642) );
  AND3X1 U15239 ( .IN1(n14644), .IN2(n14645), .IN3(n9520), .Q(WX11632) );
  OR2X1 U15240 ( .IN1(DFF_1707_n1), .IN2(WX11219), .Q(n14645) );
  OR2X1 U15241 ( .IN1(n8759), .IN2(CRC_OUT_1_11), .Q(n14644) );
  AND3X1 U15242 ( .IN1(n14646), .IN2(n14647), .IN3(n9520), .Q(WX11630) );
  OR2X1 U15243 ( .IN1(DFF_1706_n1), .IN2(n14648), .Q(n14647) );
  AND2X1 U15244 ( .IN1(n14649), .IN2(n14650), .Q(n14648) );
  OR2X1 U15245 ( .IN1(n8714), .IN2(n9085), .Q(n14650) );
  OR2X1 U15246 ( .IN1(test_so100), .IN2(WX11221), .Q(n14649) );
  OR3X1 U15247 ( .IN1(n14651), .IN2(n14652), .IN3(CRC_OUT_1_10), .Q(n14646) );
  AND2X1 U15248 ( .IN1(n8714), .IN2(n9085), .Q(n14652) );
  AND2X1 U15249 ( .IN1(test_so100), .IN2(WX11221), .Q(n14651) );
  AND3X1 U15250 ( .IN1(n14653), .IN2(n14654), .IN3(n9520), .Q(WX11628) );
  OR2X1 U15251 ( .IN1(DFF_1705_n1), .IN2(WX11223), .Q(n14654) );
  OR2X1 U15252 ( .IN1(n8760), .IN2(CRC_OUT_1_9), .Q(n14653) );
  AND3X1 U15253 ( .IN1(n14655), .IN2(n14656), .IN3(n9520), .Q(WX11626) );
  OR2X1 U15254 ( .IN1(DFF_1704_n1), .IN2(WX11225), .Q(n14656) );
  OR2X1 U15255 ( .IN1(n8761), .IN2(CRC_OUT_1_8), .Q(n14655) );
  AND3X1 U15256 ( .IN1(n14657), .IN2(n14658), .IN3(n9520), .Q(WX11624) );
  OR2X1 U15257 ( .IN1(DFF_1703_n1), .IN2(WX11227), .Q(n14658) );
  OR2X1 U15258 ( .IN1(n8762), .IN2(CRC_OUT_1_7), .Q(n14657) );
  AND3X1 U15259 ( .IN1(n14659), .IN2(n14660), .IN3(n9520), .Q(WX11622) );
  OR2X1 U15260 ( .IN1(DFF_1702_n1), .IN2(WX11229), .Q(n14660) );
  OR2X1 U15261 ( .IN1(n8763), .IN2(CRC_OUT_1_6), .Q(n14659) );
  AND3X1 U15262 ( .IN1(n14661), .IN2(n14662), .IN3(n9519), .Q(WX11620) );
  OR2X1 U15263 ( .IN1(DFF_1701_n1), .IN2(WX11231), .Q(n14662) );
  OR2X1 U15264 ( .IN1(n8764), .IN2(CRC_OUT_1_5), .Q(n14661) );
  AND3X1 U15265 ( .IN1(n14663), .IN2(n14664), .IN3(n9519), .Q(WX11618) );
  OR2X1 U15266 ( .IN1(DFF_1700_n1), .IN2(WX11233), .Q(n14664) );
  OR2X1 U15267 ( .IN1(n8765), .IN2(CRC_OUT_1_4), .Q(n14663) );
  AND3X1 U15268 ( .IN1(n14665), .IN2(n14666), .IN3(n9519), .Q(WX11616) );
  OR2X1 U15269 ( .IN1(DFF_1699_n1), .IN2(n14667), .Q(n14666) );
  AND2X1 U15270 ( .IN1(n14668), .IN2(n14669), .Q(n14667) );
  OR2X1 U15271 ( .IN1(n8715), .IN2(n9085), .Q(n14669) );
  OR2X1 U15272 ( .IN1(test_so100), .IN2(WX11235), .Q(n14668) );
  OR3X1 U15273 ( .IN1(n14670), .IN2(n14671), .IN3(CRC_OUT_1_3), .Q(n14665) );
  AND2X1 U15274 ( .IN1(n8715), .IN2(n9085), .Q(n14671) );
  AND2X1 U15275 ( .IN1(test_so100), .IN2(WX11235), .Q(n14670) );
  AND3X1 U15276 ( .IN1(n14672), .IN2(n14673), .IN3(n9519), .Q(WX11614) );
  OR2X1 U15277 ( .IN1(DFF_1698_n1), .IN2(WX11237), .Q(n14673) );
  OR2X1 U15278 ( .IN1(n8766), .IN2(CRC_OUT_1_2), .Q(n14672) );
  AND2X1 U15279 ( .IN1(n14674), .IN2(n9497), .Q(WX11612) );
  OR2X1 U15280 ( .IN1(n14675), .IN2(n14676), .Q(n14674) );
  AND2X1 U15281 ( .IN1(DFF_1697_n1), .IN2(n9102), .Q(n14676) );
  AND2X1 U15282 ( .IN1(test_so98), .IN2(CRC_OUT_1_1), .Q(n14675) );
  AND3X1 U15283 ( .IN1(n14677), .IN2(n14678), .IN3(n9519), .Q(WX11610) );
  OR2X1 U15284 ( .IN1(DFF_1696_n1), .IN2(WX11241), .Q(n14678) );
  OR2X1 U15285 ( .IN1(n8767), .IN2(CRC_OUT_1_0), .Q(n14677) );
  AND2X1 U15286 ( .IN1(n14679), .IN2(n9498), .Q(WX11608) );
  OR2X1 U15287 ( .IN1(n14680), .IN2(n14681), .Q(n14679) );
  AND2X1 U15288 ( .IN1(n8734), .IN2(n9085), .Q(n14681) );
  AND2X1 U15289 ( .IN1(test_so100), .IN2(WX11243), .Q(n14680) );
  AND2X1 U15290 ( .IN1(n9512), .IN2(n8246), .Q(WX11082) );
  AND2X1 U15291 ( .IN1(n9511), .IN2(n8247), .Q(WX11080) );
  AND2X1 U15292 ( .IN1(n9513), .IN2(n8248), .Q(WX11078) );
  AND2X1 U15293 ( .IN1(n9506), .IN2(n8249), .Q(WX11076) );
  AND2X1 U15294 ( .IN1(n9505), .IN2(n8250), .Q(WX11074) );
  AND2X1 U15295 ( .IN1(n9504), .IN2(n8251), .Q(WX11072) );
  AND2X1 U15296 ( .IN1(n9504), .IN2(n8252), .Q(WX11070) );
  AND2X1 U15297 ( .IN1(n9504), .IN2(n8253), .Q(WX11068) );
  AND2X1 U15298 ( .IN1(n9503), .IN2(n8254), .Q(WX11066) );
  AND2X1 U15299 ( .IN1(test_so91), .IN2(n9499), .Q(WX11064) );
  AND2X1 U15300 ( .IN1(n9503), .IN2(n8257), .Q(WX11062) );
  AND2X1 U15301 ( .IN1(n9502), .IN2(n8258), .Q(WX11060) );
  AND2X1 U15302 ( .IN1(n9502), .IN2(n8259), .Q(WX11058) );
  AND2X1 U15303 ( .IN1(n9503), .IN2(n8260), .Q(WX11056) );
  AND2X1 U15304 ( .IN1(n9502), .IN2(n8261), .Q(WX11054) );
  AND2X1 U15305 ( .IN1(n9502), .IN2(n8262), .Q(WX11052) );
  OR4X1 U15306 ( .IN1(n14682), .IN2(n14683), .IN3(n14684), .IN4(n14685), .Q(
        WX11050) );
  AND2X1 U15307 ( .IN1(n1985), .IN2(n9210), .Q(n14685) );
  INVX0 U15308 ( .INP(n14686), .ZN(n1985) );
  OR2X1 U15309 ( .IN1(n9559), .IN2(n3786), .Q(n14686) );
  AND2X1 U15310 ( .IN1(n9187), .IN2(n9820), .Q(n14684) );
  OR2X1 U15311 ( .IN1(n14687), .IN2(n14688), .Q(n9820) );
  INVX0 U15312 ( .INP(n14689), .ZN(n14688) );
  OR2X1 U15313 ( .IN1(n14690), .IN2(n14691), .Q(n14689) );
  AND2X1 U15314 ( .IN1(n14691), .IN2(n14690), .Q(n14687) );
  AND2X1 U15315 ( .IN1(n14692), .IN2(n14693), .Q(n14690) );
  OR2X1 U15316 ( .IN1(WX11115), .IN2(n8118), .Q(n14693) );
  INVX0 U15317 ( .INP(n14694), .ZN(n14692) );
  AND2X1 U15318 ( .IN1(n8118), .IN2(WX11115), .Q(n14694) );
  OR2X1 U15319 ( .IN1(n14695), .IN2(n14696), .Q(n14691) );
  AND2X1 U15320 ( .IN1(n8119), .IN2(WX11243), .Q(n14696) );
  AND2X1 U15321 ( .IN1(n8734), .IN2(WX11179), .Q(n14695) );
  AND2X1 U15322 ( .IN1(n9236), .IN2(CRC_OUT_1_0), .Q(n14683) );
  AND2X1 U15323 ( .IN1(DATA_0_0), .IN2(n9260), .Q(n14682) );
  OR4X1 U15324 ( .IN1(n14697), .IN2(n14698), .IN3(n14699), .IN4(n14700), .Q(
        WX11048) );
  AND2X1 U15325 ( .IN1(n1984), .IN2(n9210), .Q(n14700) );
  INVX0 U15326 ( .INP(n14701), .ZN(n1984) );
  OR2X1 U15327 ( .IN1(n9559), .IN2(n3787), .Q(n14701) );
  AND2X1 U15328 ( .IN1(n9187), .IN2(n9828), .Q(n14699) );
  OR2X1 U15329 ( .IN1(n14702), .IN2(n14703), .Q(n9828) );
  INVX0 U15330 ( .INP(n14704), .ZN(n14703) );
  OR2X1 U15331 ( .IN1(n14705), .IN2(n14706), .Q(n14704) );
  AND2X1 U15332 ( .IN1(n14706), .IN2(n14705), .Q(n14702) );
  AND2X1 U15333 ( .IN1(n14707), .IN2(n14708), .Q(n14705) );
  OR2X1 U15334 ( .IN1(WX11113), .IN2(n8120), .Q(n14708) );
  INVX0 U15335 ( .INP(n14709), .ZN(n14707) );
  AND2X1 U15336 ( .IN1(n8120), .IN2(WX11113), .Q(n14709) );
  OR2X1 U15337 ( .IN1(n14710), .IN2(n14711), .Q(n14706) );
  AND2X1 U15338 ( .IN1(n8121), .IN2(WX11241), .Q(n14711) );
  AND2X1 U15339 ( .IN1(n8767), .IN2(WX11177), .Q(n14710) );
  AND2X1 U15340 ( .IN1(n9236), .IN2(CRC_OUT_1_1), .Q(n14698) );
  AND2X1 U15341 ( .IN1(DATA_0_1), .IN2(n9261), .Q(n14697) );
  OR4X1 U15342 ( .IN1(n14712), .IN2(n14713), .IN3(n14714), .IN4(n14715), .Q(
        WX11046) );
  AND2X1 U15343 ( .IN1(n1983), .IN2(n9210), .Q(n14715) );
  INVX0 U15344 ( .INP(n14716), .ZN(n1983) );
  OR2X1 U15345 ( .IN1(n9559), .IN2(n3788), .Q(n14716) );
  AND2X1 U15346 ( .IN1(n9835), .IN2(n9174), .Q(n14714) );
  AND2X1 U15347 ( .IN1(n14717), .IN2(n14718), .Q(n9835) );
  INVX0 U15348 ( .INP(n14719), .ZN(n14718) );
  AND2X1 U15349 ( .IN1(n14720), .IN2(n14721), .Q(n14719) );
  OR2X1 U15350 ( .IN1(n14721), .IN2(n14720), .Q(n14717) );
  OR2X1 U15351 ( .IN1(n14722), .IN2(n14723), .Q(n14720) );
  INVX0 U15352 ( .INP(n14724), .ZN(n14723) );
  OR2X1 U15353 ( .IN1(WX11111), .IN2(n8122), .Q(n14724) );
  AND2X1 U15354 ( .IN1(n8122), .IN2(WX11111), .Q(n14722) );
  AND2X1 U15355 ( .IN1(n14725), .IN2(n14726), .Q(n14721) );
  OR2X1 U15356 ( .IN1(WX11175), .IN2(test_so98), .Q(n14726) );
  OR2X1 U15357 ( .IN1(n9102), .IN2(n8123), .Q(n14725) );
  AND2X1 U15358 ( .IN1(n9236), .IN2(CRC_OUT_1_2), .Q(n14713) );
  AND2X1 U15359 ( .IN1(DATA_0_2), .IN2(n9262), .Q(n14712) );
  OR4X1 U15360 ( .IN1(n14727), .IN2(n14728), .IN3(n14729), .IN4(n14730), .Q(
        WX11044) );
  AND2X1 U15361 ( .IN1(n1982), .IN2(n9210), .Q(n14730) );
  INVX0 U15362 ( .INP(n14731), .ZN(n1982) );
  OR2X1 U15363 ( .IN1(n9559), .IN2(n3789), .Q(n14731) );
  AND2X1 U15364 ( .IN1(n9187), .IN2(n9842), .Q(n14729) );
  OR2X1 U15365 ( .IN1(n14732), .IN2(n14733), .Q(n9842) );
  INVX0 U15366 ( .INP(n14734), .ZN(n14733) );
  OR2X1 U15367 ( .IN1(n14735), .IN2(n14736), .Q(n14734) );
  AND2X1 U15368 ( .IN1(n14736), .IN2(n14735), .Q(n14732) );
  AND2X1 U15369 ( .IN1(n14737), .IN2(n14738), .Q(n14735) );
  OR2X1 U15370 ( .IN1(WX11109), .IN2(n8124), .Q(n14738) );
  INVX0 U15371 ( .INP(n14739), .ZN(n14737) );
  AND2X1 U15372 ( .IN1(n8124), .IN2(WX11109), .Q(n14739) );
  OR2X1 U15373 ( .IN1(n14740), .IN2(n14741), .Q(n14736) );
  AND2X1 U15374 ( .IN1(n8125), .IN2(WX11237), .Q(n14741) );
  AND2X1 U15375 ( .IN1(n8766), .IN2(WX11173), .Q(n14740) );
  AND2X1 U15376 ( .IN1(n9236), .IN2(CRC_OUT_1_3), .Q(n14728) );
  AND2X1 U15377 ( .IN1(DATA_0_3), .IN2(n9262), .Q(n14727) );
  OR4X1 U15378 ( .IN1(n14742), .IN2(n14743), .IN3(n14744), .IN4(n14745), .Q(
        WX11042) );
  AND2X1 U15379 ( .IN1(n1981), .IN2(n9210), .Q(n14745) );
  INVX0 U15380 ( .INP(n14746), .ZN(n1981) );
  OR2X1 U15381 ( .IN1(n9559), .IN2(n3790), .Q(n14746) );
  AND2X1 U15382 ( .IN1(n9849), .IN2(n9174), .Q(n14744) );
  AND2X1 U15383 ( .IN1(n14747), .IN2(n14748), .Q(n9849) );
  INVX0 U15384 ( .INP(n14749), .ZN(n14748) );
  AND2X1 U15385 ( .IN1(n14750), .IN2(n14751), .Q(n14749) );
  OR2X1 U15386 ( .IN1(n14751), .IN2(n14750), .Q(n14747) );
  OR2X1 U15387 ( .IN1(n14752), .IN2(n14753), .Q(n14750) );
  INVX0 U15388 ( .INP(n14754), .ZN(n14753) );
  OR2X1 U15389 ( .IN1(WX11107), .IN2(n8126), .Q(n14754) );
  AND2X1 U15390 ( .IN1(n8126), .IN2(WX11107), .Q(n14752) );
  AND2X1 U15391 ( .IN1(n14755), .IN2(n14756), .Q(n14751) );
  OR2X1 U15392 ( .IN1(WX11235), .IN2(test_so96), .Q(n14756) );
  OR2X1 U15393 ( .IN1(n9142), .IN2(n8715), .Q(n14755) );
  AND2X1 U15394 ( .IN1(n9236), .IN2(CRC_OUT_1_4), .Q(n14743) );
  AND2X1 U15395 ( .IN1(DATA_0_4), .IN2(n9262), .Q(n14742) );
  OR4X1 U15396 ( .IN1(n14757), .IN2(n14758), .IN3(n14759), .IN4(n14760), .Q(
        WX11040) );
  AND2X1 U15397 ( .IN1(n1980), .IN2(n9210), .Q(n14760) );
  INVX0 U15398 ( .INP(n14761), .ZN(n1980) );
  OR2X1 U15399 ( .IN1(n9559), .IN2(n3791), .Q(n14761) );
  AND2X1 U15400 ( .IN1(n9187), .IN2(n9856), .Q(n14759) );
  OR2X1 U15401 ( .IN1(n14762), .IN2(n14763), .Q(n9856) );
  INVX0 U15402 ( .INP(n14764), .ZN(n14763) );
  OR2X1 U15403 ( .IN1(n14765), .IN2(n14766), .Q(n14764) );
  AND2X1 U15404 ( .IN1(n14766), .IN2(n14765), .Q(n14762) );
  AND2X1 U15405 ( .IN1(n14767), .IN2(n14768), .Q(n14765) );
  OR2X1 U15406 ( .IN1(WX11105), .IN2(n8127), .Q(n14768) );
  INVX0 U15407 ( .INP(n14769), .ZN(n14767) );
  AND2X1 U15408 ( .IN1(n8127), .IN2(WX11105), .Q(n14769) );
  OR2X1 U15409 ( .IN1(n14770), .IN2(n14771), .Q(n14766) );
  AND2X1 U15410 ( .IN1(n8128), .IN2(WX11233), .Q(n14771) );
  AND2X1 U15411 ( .IN1(n8765), .IN2(WX11169), .Q(n14770) );
  AND2X1 U15412 ( .IN1(n9236), .IN2(CRC_OUT_1_5), .Q(n14758) );
  AND2X1 U15413 ( .IN1(DATA_0_5), .IN2(n9262), .Q(n14757) );
  OR4X1 U15414 ( .IN1(n14772), .IN2(n14773), .IN3(n14774), .IN4(n14775), .Q(
        WX11038) );
  AND2X1 U15415 ( .IN1(n1979), .IN2(n9210), .Q(n14775) );
  INVX0 U15416 ( .INP(n14776), .ZN(n1979) );
  OR2X1 U15417 ( .IN1(n9559), .IN2(n3792), .Q(n14776) );
  AND2X1 U15418 ( .IN1(n9863), .IN2(n9174), .Q(n14774) );
  AND2X1 U15419 ( .IN1(n14777), .IN2(n14778), .Q(n9863) );
  INVX0 U15420 ( .INP(n14779), .ZN(n14778) );
  AND2X1 U15421 ( .IN1(n14780), .IN2(n14781), .Q(n14779) );
  OR2X1 U15422 ( .IN1(n14781), .IN2(n14780), .Q(n14777) );
  OR2X1 U15423 ( .IN1(n14782), .IN2(n14783), .Q(n14780) );
  INVX0 U15424 ( .INP(n14784), .ZN(n14783) );
  OR2X1 U15425 ( .IN1(WX11039), .IN2(n8130), .Q(n14784) );
  AND2X1 U15426 ( .IN1(n8130), .IN2(WX11039), .Q(n14782) );
  AND2X1 U15427 ( .IN1(n14785), .IN2(n14786), .Q(n14781) );
  OR2X1 U15428 ( .IN1(WX11231), .IN2(test_so94), .Q(n14786) );
  OR2X1 U15429 ( .IN1(n9143), .IN2(n8764), .Q(n14785) );
  AND2X1 U15430 ( .IN1(n9236), .IN2(CRC_OUT_1_6), .Q(n14773) );
  AND2X1 U15431 ( .IN1(DATA_0_6), .IN2(n9262), .Q(n14772) );
  OR4X1 U15432 ( .IN1(n14787), .IN2(n14788), .IN3(n14789), .IN4(n14790), .Q(
        WX11036) );
  AND2X1 U15433 ( .IN1(n1978), .IN2(n9210), .Q(n14790) );
  INVX0 U15434 ( .INP(n14791), .ZN(n1978) );
  OR2X1 U15435 ( .IN1(n9558), .IN2(n3793), .Q(n14791) );
  AND2X1 U15436 ( .IN1(n9187), .IN2(n9870), .Q(n14789) );
  OR2X1 U15437 ( .IN1(n14792), .IN2(n14793), .Q(n9870) );
  INVX0 U15438 ( .INP(n14794), .ZN(n14793) );
  OR2X1 U15439 ( .IN1(n14795), .IN2(n14796), .Q(n14794) );
  AND2X1 U15440 ( .IN1(n14796), .IN2(n14795), .Q(n14792) );
  AND2X1 U15441 ( .IN1(n14797), .IN2(n14798), .Q(n14795) );
  OR2X1 U15442 ( .IN1(WX11101), .IN2(n8131), .Q(n14798) );
  INVX0 U15443 ( .INP(n14799), .ZN(n14797) );
  AND2X1 U15444 ( .IN1(n8131), .IN2(WX11101), .Q(n14799) );
  OR2X1 U15445 ( .IN1(n14800), .IN2(n14801), .Q(n14796) );
  AND2X1 U15446 ( .IN1(n8132), .IN2(WX11229), .Q(n14801) );
  AND2X1 U15447 ( .IN1(n8763), .IN2(WX11165), .Q(n14800) );
  AND2X1 U15448 ( .IN1(n9236), .IN2(CRC_OUT_1_7), .Q(n14788) );
  AND2X1 U15449 ( .IN1(DATA_0_7), .IN2(n9263), .Q(n14787) );
  OR4X1 U15450 ( .IN1(n14802), .IN2(n14803), .IN3(n14804), .IN4(n14805), .Q(
        WX11034) );
  AND2X1 U15451 ( .IN1(n1977), .IN2(n9210), .Q(n14805) );
  INVX0 U15452 ( .INP(n14806), .ZN(n1977) );
  OR2X1 U15453 ( .IN1(n9558), .IN2(n3794), .Q(n14806) );
  AND2X1 U15454 ( .IN1(n9877), .IN2(n9174), .Q(n14804) );
  AND2X1 U15455 ( .IN1(n14807), .IN2(n14808), .Q(n9877) );
  INVX0 U15456 ( .INP(n14809), .ZN(n14808) );
  AND2X1 U15457 ( .IN1(n14810), .IN2(n14811), .Q(n14809) );
  OR2X1 U15458 ( .IN1(n14811), .IN2(n14810), .Q(n14807) );
  OR2X1 U15459 ( .IN1(n14812), .IN2(n14813), .Q(n14810) );
  INVX0 U15460 ( .INP(n14814), .ZN(n14813) );
  OR2X1 U15461 ( .IN1(WX11099), .IN2(n8133), .Q(n14814) );
  AND2X1 U15462 ( .IN1(n8133), .IN2(WX11099), .Q(n14812) );
  AND2X1 U15463 ( .IN1(n14815), .IN2(n14816), .Q(n14811) );
  OR2X1 U15464 ( .IN1(WX11227), .IN2(test_so92), .Q(n14816) );
  OR2X1 U15465 ( .IN1(n9144), .IN2(n8762), .Q(n14815) );
  AND2X1 U15466 ( .IN1(n9236), .IN2(CRC_OUT_1_8), .Q(n14803) );
  AND2X1 U15467 ( .IN1(DATA_0_8), .IN2(n9263), .Q(n14802) );
  OR4X1 U15468 ( .IN1(n14817), .IN2(n14818), .IN3(n14819), .IN4(n14820), .Q(
        WX11032) );
  AND2X1 U15469 ( .IN1(n1976), .IN2(n9210), .Q(n14820) );
  INVX0 U15470 ( .INP(n14821), .ZN(n1976) );
  OR2X1 U15471 ( .IN1(n9558), .IN2(n3795), .Q(n14821) );
  AND2X1 U15472 ( .IN1(n9187), .IN2(n9884), .Q(n14819) );
  OR2X1 U15473 ( .IN1(n14822), .IN2(n14823), .Q(n9884) );
  INVX0 U15474 ( .INP(n14824), .ZN(n14823) );
  OR2X1 U15475 ( .IN1(n14825), .IN2(n14826), .Q(n14824) );
  AND2X1 U15476 ( .IN1(n14826), .IN2(n14825), .Q(n14822) );
  AND2X1 U15477 ( .IN1(n14827), .IN2(n14828), .Q(n14825) );
  OR2X1 U15478 ( .IN1(WX11097), .IN2(n8134), .Q(n14828) );
  INVX0 U15479 ( .INP(n14829), .ZN(n14827) );
  AND2X1 U15480 ( .IN1(n8134), .IN2(WX11097), .Q(n14829) );
  OR2X1 U15481 ( .IN1(n14830), .IN2(n14831), .Q(n14826) );
  AND2X1 U15482 ( .IN1(n8135), .IN2(WX11225), .Q(n14831) );
  AND2X1 U15483 ( .IN1(n8761), .IN2(WX11161), .Q(n14830) );
  AND2X1 U15484 ( .IN1(n9236), .IN2(CRC_OUT_1_9), .Q(n14818) );
  AND2X1 U15485 ( .IN1(DATA_0_9), .IN2(n9263), .Q(n14817) );
  OR4X1 U15486 ( .IN1(n14832), .IN2(n14833), .IN3(n14834), .IN4(n14835), .Q(
        WX11030) );
  AND2X1 U15487 ( .IN1(n1975), .IN2(n9211), .Q(n14835) );
  INVX0 U15488 ( .INP(n14836), .ZN(n1975) );
  OR2X1 U15489 ( .IN1(n9558), .IN2(n3796), .Q(n14836) );
  AND2X1 U15490 ( .IN1(n9187), .IN2(n9891), .Q(n14834) );
  OR2X1 U15491 ( .IN1(n14837), .IN2(n14838), .Q(n9891) );
  INVX0 U15492 ( .INP(n14839), .ZN(n14838) );
  OR2X1 U15493 ( .IN1(n14840), .IN2(n14841), .Q(n14839) );
  AND2X1 U15494 ( .IN1(n14841), .IN2(n14840), .Q(n14837) );
  AND2X1 U15495 ( .IN1(n14842), .IN2(n14843), .Q(n14840) );
  OR2X1 U15496 ( .IN1(WX11095), .IN2(n8136), .Q(n14843) );
  INVX0 U15497 ( .INP(n14844), .ZN(n14842) );
  AND2X1 U15498 ( .IN1(n8136), .IN2(WX11095), .Q(n14844) );
  OR2X1 U15499 ( .IN1(n14845), .IN2(n14846), .Q(n14841) );
  AND2X1 U15500 ( .IN1(n8137), .IN2(WX11223), .Q(n14846) );
  AND2X1 U15501 ( .IN1(n8760), .IN2(WX11159), .Q(n14845) );
  AND2X1 U15502 ( .IN1(n9237), .IN2(CRC_OUT_1_10), .Q(n14833) );
  AND2X1 U15503 ( .IN1(DATA_0_10), .IN2(n9263), .Q(n14832) );
  OR4X1 U15504 ( .IN1(n14847), .IN2(n14848), .IN3(n14849), .IN4(n14850), .Q(
        WX11028) );
  AND2X1 U15505 ( .IN1(n1974), .IN2(n9211), .Q(n14850) );
  INVX0 U15506 ( .INP(n14851), .ZN(n1974) );
  OR2X1 U15507 ( .IN1(n9558), .IN2(n3797), .Q(n14851) );
  AND2X1 U15508 ( .IN1(n9187), .IN2(n9898), .Q(n14849) );
  OR2X1 U15509 ( .IN1(n14852), .IN2(n14853), .Q(n9898) );
  INVX0 U15510 ( .INP(n14854), .ZN(n14853) );
  OR2X1 U15511 ( .IN1(n14855), .IN2(n14856), .Q(n14854) );
  AND2X1 U15512 ( .IN1(n14856), .IN2(n14855), .Q(n14852) );
  AND2X1 U15513 ( .IN1(n14857), .IN2(n14858), .Q(n14855) );
  OR2X1 U15514 ( .IN1(WX11093), .IN2(n8138), .Q(n14858) );
  INVX0 U15515 ( .INP(n14859), .ZN(n14857) );
  AND2X1 U15516 ( .IN1(n8138), .IN2(WX11093), .Q(n14859) );
  OR2X1 U15517 ( .IN1(n14860), .IN2(n14861), .Q(n14856) );
  AND2X1 U15518 ( .IN1(n8139), .IN2(WX11221), .Q(n14861) );
  AND2X1 U15519 ( .IN1(n8714), .IN2(WX11157), .Q(n14860) );
  AND2X1 U15520 ( .IN1(n9237), .IN2(CRC_OUT_1_11), .Q(n14848) );
  AND2X1 U15521 ( .IN1(DATA_0_11), .IN2(n9261), .Q(n14847) );
  OR4X1 U15522 ( .IN1(n14862), .IN2(n14863), .IN3(n14864), .IN4(n14865), .Q(
        WX11026) );
  AND2X1 U15523 ( .IN1(n1973), .IN2(n9211), .Q(n14865) );
  INVX0 U15524 ( .INP(n14866), .ZN(n1973) );
  OR2X1 U15525 ( .IN1(n9558), .IN2(n3798), .Q(n14866) );
  AND2X1 U15526 ( .IN1(n9186), .IN2(n9905), .Q(n14864) );
  OR2X1 U15527 ( .IN1(n14867), .IN2(n14868), .Q(n9905) );
  INVX0 U15528 ( .INP(n14869), .ZN(n14868) );
  OR2X1 U15529 ( .IN1(n14870), .IN2(n14871), .Q(n14869) );
  AND2X1 U15530 ( .IN1(n14871), .IN2(n14870), .Q(n14867) );
  AND2X1 U15531 ( .IN1(n14872), .IN2(n14873), .Q(n14870) );
  OR2X1 U15532 ( .IN1(WX11091), .IN2(n8140), .Q(n14873) );
  INVX0 U15533 ( .INP(n14874), .ZN(n14872) );
  AND2X1 U15534 ( .IN1(n8140), .IN2(WX11091), .Q(n14874) );
  OR2X1 U15535 ( .IN1(n14875), .IN2(n14876), .Q(n14871) );
  AND2X1 U15536 ( .IN1(n8141), .IN2(WX11219), .Q(n14876) );
  AND2X1 U15537 ( .IN1(n8759), .IN2(WX11155), .Q(n14875) );
  AND2X1 U15538 ( .IN1(n9237), .IN2(CRC_OUT_1_12), .Q(n14863) );
  AND2X1 U15539 ( .IN1(DATA_0_12), .IN2(n9263), .Q(n14862) );
  OR4X1 U15540 ( .IN1(n14877), .IN2(n14878), .IN3(n14879), .IN4(n14880), .Q(
        WX11024) );
  AND2X1 U15541 ( .IN1(n1972), .IN2(n9211), .Q(n14880) );
  INVX0 U15542 ( .INP(n14881), .ZN(n1972) );
  OR2X1 U15543 ( .IN1(n9558), .IN2(n3799), .Q(n14881) );
  AND2X1 U15544 ( .IN1(n9186), .IN2(n9912), .Q(n14879) );
  OR2X1 U15545 ( .IN1(n14882), .IN2(n14883), .Q(n9912) );
  INVX0 U15546 ( .INP(n14884), .ZN(n14883) );
  OR2X1 U15547 ( .IN1(n14885), .IN2(n14886), .Q(n14884) );
  AND2X1 U15548 ( .IN1(n14886), .IN2(n14885), .Q(n14882) );
  AND2X1 U15549 ( .IN1(n14887), .IN2(n14888), .Q(n14885) );
  OR2X1 U15550 ( .IN1(WX11089), .IN2(n8142), .Q(n14888) );
  INVX0 U15551 ( .INP(n14889), .ZN(n14887) );
  AND2X1 U15552 ( .IN1(n8142), .IN2(WX11089), .Q(n14889) );
  OR2X1 U15553 ( .IN1(n14890), .IN2(n14891), .Q(n14886) );
  AND2X1 U15554 ( .IN1(n8143), .IN2(WX11217), .Q(n14891) );
  AND2X1 U15555 ( .IN1(n8758), .IN2(WX11153), .Q(n14890) );
  AND2X1 U15556 ( .IN1(n9237), .IN2(CRC_OUT_1_13), .Q(n14878) );
  AND2X1 U15557 ( .IN1(DATA_0_13), .IN2(n9263), .Q(n14877) );
  OR4X1 U15558 ( .IN1(n14892), .IN2(n14893), .IN3(n14894), .IN4(n14895), .Q(
        WX11022) );
  AND2X1 U15559 ( .IN1(n1971), .IN2(n9211), .Q(n14895) );
  INVX0 U15560 ( .INP(n14896), .ZN(n1971) );
  OR2X1 U15561 ( .IN1(n9558), .IN2(n3800), .Q(n14896) );
  AND2X1 U15562 ( .IN1(n9186), .IN2(n9919), .Q(n14894) );
  OR2X1 U15563 ( .IN1(n14897), .IN2(n14898), .Q(n9919) );
  INVX0 U15564 ( .INP(n14899), .ZN(n14898) );
  OR2X1 U15565 ( .IN1(n14900), .IN2(n14901), .Q(n14899) );
  AND2X1 U15566 ( .IN1(n14901), .IN2(n14900), .Q(n14897) );
  AND2X1 U15567 ( .IN1(n14902), .IN2(n14903), .Q(n14900) );
  OR2X1 U15568 ( .IN1(WX11087), .IN2(n8144), .Q(n14903) );
  INVX0 U15569 ( .INP(n14904), .ZN(n14902) );
  AND2X1 U15570 ( .IN1(n8144), .IN2(WX11087), .Q(n14904) );
  OR2X1 U15571 ( .IN1(n14905), .IN2(n14906), .Q(n14901) );
  AND2X1 U15572 ( .IN1(n8145), .IN2(WX11215), .Q(n14906) );
  AND2X1 U15573 ( .IN1(n8757), .IN2(WX11151), .Q(n14905) );
  AND2X1 U15574 ( .IN1(test_so99), .IN2(n9227), .Q(n14893) );
  AND2X1 U15575 ( .IN1(DATA_0_14), .IN2(n9264), .Q(n14892) );
  OR4X1 U15576 ( .IN1(n14907), .IN2(n14908), .IN3(n14909), .IN4(n14910), .Q(
        WX11020) );
  AND2X1 U15577 ( .IN1(n1970), .IN2(n9211), .Q(n14910) );
  INVX0 U15578 ( .INP(n14911), .ZN(n1970) );
  OR2X1 U15579 ( .IN1(n9558), .IN2(n3801), .Q(n14911) );
  AND2X1 U15580 ( .IN1(n9186), .IN2(n9926), .Q(n14909) );
  OR2X1 U15581 ( .IN1(n14912), .IN2(n14913), .Q(n9926) );
  INVX0 U15582 ( .INP(n14914), .ZN(n14913) );
  OR2X1 U15583 ( .IN1(n14915), .IN2(n14916), .Q(n14914) );
  AND2X1 U15584 ( .IN1(n14916), .IN2(n14915), .Q(n14912) );
  AND2X1 U15585 ( .IN1(n14917), .IN2(n14918), .Q(n14915) );
  OR2X1 U15586 ( .IN1(WX11085), .IN2(n8146), .Q(n14918) );
  INVX0 U15587 ( .INP(n14919), .ZN(n14917) );
  AND2X1 U15588 ( .IN1(n8146), .IN2(WX11085), .Q(n14919) );
  OR2X1 U15589 ( .IN1(n14920), .IN2(n14921), .Q(n14916) );
  AND2X1 U15590 ( .IN1(n8147), .IN2(WX11213), .Q(n14921) );
  AND2X1 U15591 ( .IN1(n8756), .IN2(WX11149), .Q(n14920) );
  AND2X1 U15592 ( .IN1(n9237), .IN2(CRC_OUT_1_15), .Q(n14908) );
  AND2X1 U15593 ( .IN1(DATA_0_15), .IN2(n9264), .Q(n14907) );
  OR4X1 U15594 ( .IN1(n14922), .IN2(n14923), .IN3(n14924), .IN4(n14925), .Q(
        WX11018) );
  AND2X1 U15595 ( .IN1(n1969), .IN2(n9211), .Q(n14925) );
  INVX0 U15596 ( .INP(n14926), .ZN(n1969) );
  OR2X1 U15597 ( .IN1(n9558), .IN2(n3802), .Q(n14926) );
  AND2X1 U15598 ( .IN1(n9186), .IN2(n9933), .Q(n14924) );
  OR2X1 U15599 ( .IN1(n14927), .IN2(n14928), .Q(n9933) );
  INVX0 U15600 ( .INP(n14929), .ZN(n14928) );
  OR2X1 U15601 ( .IN1(n14930), .IN2(n14931), .Q(n14929) );
  AND2X1 U15602 ( .IN1(n14931), .IN2(n14930), .Q(n14927) );
  AND2X1 U15603 ( .IN1(n14932), .IN2(n14933), .Q(n14930) );
  OR2X1 U15604 ( .IN1(n9474), .IN2(n7892), .Q(n14933) );
  OR2X1 U15605 ( .IN1(WX11083), .IN2(n9443), .Q(n14932) );
  OR2X1 U15606 ( .IN1(n14934), .IN2(n14935), .Q(n14931) );
  INVX0 U15607 ( .INP(n14936), .ZN(n14935) );
  OR2X1 U15608 ( .IN1(n14937), .IN2(n7893), .Q(n14936) );
  AND2X1 U15609 ( .IN1(n7893), .IN2(n14937), .Q(n14934) );
  INVX0 U15610 ( .INP(n14938), .ZN(n14937) );
  OR2X1 U15611 ( .IN1(n14939), .IN2(n14940), .Q(n14938) );
  AND2X1 U15612 ( .IN1(n8713), .IN2(n8246), .Q(n14940) );
  AND2X1 U15613 ( .IN1(n15983), .IN2(WX11211), .Q(n14939) );
  AND2X1 U15614 ( .IN1(n9237), .IN2(CRC_OUT_1_16), .Q(n14923) );
  AND2X1 U15615 ( .IN1(DATA_0_16), .IN2(n9263), .Q(n14922) );
  OR4X1 U15616 ( .IN1(n14941), .IN2(n14942), .IN3(n14943), .IN4(n14944), .Q(
        WX11016) );
  AND2X1 U15617 ( .IN1(n1968), .IN2(n9211), .Q(n14944) );
  INVX0 U15618 ( .INP(n14945), .ZN(n1968) );
  OR2X1 U15619 ( .IN1(n9558), .IN2(n3803), .Q(n14945) );
  AND2X1 U15620 ( .IN1(n9186), .IN2(n9940), .Q(n14943) );
  OR2X1 U15621 ( .IN1(n14946), .IN2(n14947), .Q(n9940) );
  INVX0 U15622 ( .INP(n14948), .ZN(n14947) );
  OR2X1 U15623 ( .IN1(n14949), .IN2(n14950), .Q(n14948) );
  AND2X1 U15624 ( .IN1(n14950), .IN2(n14949), .Q(n14946) );
  AND2X1 U15625 ( .IN1(n14951), .IN2(n14952), .Q(n14949) );
  OR2X1 U15626 ( .IN1(n9474), .IN2(n7894), .Q(n14952) );
  OR2X1 U15627 ( .IN1(WX11081), .IN2(n9442), .Q(n14951) );
  OR2X1 U15628 ( .IN1(n14953), .IN2(n14954), .Q(n14950) );
  INVX0 U15629 ( .INP(n14955), .ZN(n14954) );
  OR2X1 U15630 ( .IN1(n14956), .IN2(n7895), .Q(n14955) );
  AND2X1 U15631 ( .IN1(n7895), .IN2(n14956), .Q(n14953) );
  INVX0 U15632 ( .INP(n14957), .ZN(n14956) );
  OR2X1 U15633 ( .IN1(n14958), .IN2(n14959), .Q(n14957) );
  AND2X1 U15634 ( .IN1(n8755), .IN2(n8247), .Q(n14959) );
  AND2X1 U15635 ( .IN1(n15984), .IN2(WX11209), .Q(n14958) );
  AND2X1 U15636 ( .IN1(n9237), .IN2(CRC_OUT_1_17), .Q(n14942) );
  AND2X1 U15637 ( .IN1(DATA_0_17), .IN2(n9264), .Q(n14941) );
  OR4X1 U15638 ( .IN1(n14960), .IN2(n14961), .IN3(n14962), .IN4(n14963), .Q(
        WX11014) );
  AND2X1 U15639 ( .IN1(n1967), .IN2(n9211), .Q(n14963) );
  INVX0 U15640 ( .INP(n14964), .ZN(n1967) );
  OR2X1 U15641 ( .IN1(n9558), .IN2(n3804), .Q(n14964) );
  AND2X1 U15642 ( .IN1(n9186), .IN2(n9947), .Q(n14962) );
  OR2X1 U15643 ( .IN1(n14965), .IN2(n14966), .Q(n9947) );
  INVX0 U15644 ( .INP(n14967), .ZN(n14966) );
  OR2X1 U15645 ( .IN1(n14968), .IN2(n14969), .Q(n14967) );
  AND2X1 U15646 ( .IN1(n14969), .IN2(n14968), .Q(n14965) );
  AND2X1 U15647 ( .IN1(n14970), .IN2(n14971), .Q(n14968) );
  OR2X1 U15648 ( .IN1(n9475), .IN2(n7896), .Q(n14971) );
  OR2X1 U15649 ( .IN1(WX11079), .IN2(n9442), .Q(n14970) );
  OR2X1 U15650 ( .IN1(n14972), .IN2(n14973), .Q(n14969) );
  INVX0 U15651 ( .INP(n14974), .ZN(n14973) );
  OR2X1 U15652 ( .IN1(n14975), .IN2(n7897), .Q(n14974) );
  AND2X1 U15653 ( .IN1(n7897), .IN2(n14975), .Q(n14972) );
  INVX0 U15654 ( .INP(n14976), .ZN(n14975) );
  OR2X1 U15655 ( .IN1(n14977), .IN2(n14978), .Q(n14976) );
  AND2X1 U15656 ( .IN1(n8754), .IN2(n8248), .Q(n14978) );
  AND2X1 U15657 ( .IN1(n15985), .IN2(WX11207), .Q(n14977) );
  AND2X1 U15658 ( .IN1(n9237), .IN2(CRC_OUT_1_18), .Q(n14961) );
  AND2X1 U15659 ( .IN1(DATA_0_18), .IN2(n9262), .Q(n14960) );
  OR4X1 U15660 ( .IN1(n14979), .IN2(n14980), .IN3(n14981), .IN4(n14982), .Q(
        WX11012) );
  AND2X1 U15661 ( .IN1(n1966), .IN2(n9211), .Q(n14982) );
  INVX0 U15662 ( .INP(n14983), .ZN(n1966) );
  OR2X1 U15663 ( .IN1(n9557), .IN2(n3805), .Q(n14983) );
  AND2X1 U15664 ( .IN1(n9954), .IN2(n9173), .Q(n14981) );
  AND2X1 U15665 ( .IN1(n14984), .IN2(n14985), .Q(n9954) );
  INVX0 U15666 ( .INP(n14986), .ZN(n14985) );
  AND2X1 U15667 ( .IN1(n14987), .IN2(n14988), .Q(n14986) );
  OR2X1 U15668 ( .IN1(n14988), .IN2(n14987), .Q(n14984) );
  OR2X1 U15669 ( .IN1(n14989), .IN2(n14990), .Q(n14987) );
  AND2X1 U15670 ( .IN1(n9451), .IN2(WX11077), .Q(n14990) );
  AND2X1 U15671 ( .IN1(n7898), .IN2(n9474), .Q(n14989) );
  AND2X1 U15672 ( .IN1(n14991), .IN2(n14992), .Q(n14988) );
  OR2X1 U15673 ( .IN1(n14993), .IN2(n7899), .Q(n14992) );
  INVX0 U15674 ( .INP(n14994), .ZN(n14993) );
  OR2X1 U15675 ( .IN1(WX11141), .IN2(n14994), .Q(n14991) );
  OR2X1 U15676 ( .IN1(n14995), .IN2(n14996), .Q(n14994) );
  AND2X1 U15677 ( .IN1(n15986), .IN2(n9109), .Q(n14996) );
  AND2X1 U15678 ( .IN1(test_so97), .IN2(n8249), .Q(n14995) );
  AND2X1 U15679 ( .IN1(n9237), .IN2(CRC_OUT_1_19), .Q(n14980) );
  AND2X1 U15680 ( .IN1(DATA_0_19), .IN2(n9261), .Q(n14979) );
  OR4X1 U15681 ( .IN1(n14997), .IN2(n14998), .IN3(n14999), .IN4(n15000), .Q(
        WX11010) );
  AND2X1 U15682 ( .IN1(n1965), .IN2(n9211), .Q(n15000) );
  INVX0 U15683 ( .INP(n15001), .ZN(n1965) );
  OR2X1 U15684 ( .IN1(n9557), .IN2(n3806), .Q(n15001) );
  AND2X1 U15685 ( .IN1(n9186), .IN2(n9961), .Q(n14999) );
  OR2X1 U15686 ( .IN1(n15002), .IN2(n15003), .Q(n9961) );
  INVX0 U15687 ( .INP(n15004), .ZN(n15003) );
  OR2X1 U15688 ( .IN1(n15005), .IN2(n15006), .Q(n15004) );
  AND2X1 U15689 ( .IN1(n15006), .IN2(n15005), .Q(n15002) );
  AND2X1 U15690 ( .IN1(n15007), .IN2(n15008), .Q(n15005) );
  OR2X1 U15691 ( .IN1(n9476), .IN2(n7900), .Q(n15008) );
  OR2X1 U15692 ( .IN1(WX11075), .IN2(n9442), .Q(n15007) );
  OR2X1 U15693 ( .IN1(n15009), .IN2(n15010), .Q(n15006) );
  INVX0 U15694 ( .INP(n15011), .ZN(n15010) );
  OR2X1 U15695 ( .IN1(n15012), .IN2(n7901), .Q(n15011) );
  AND2X1 U15696 ( .IN1(n7901), .IN2(n15012), .Q(n15009) );
  INVX0 U15697 ( .INP(n15013), .ZN(n15012) );
  OR2X1 U15698 ( .IN1(n15014), .IN2(n15015), .Q(n15013) );
  AND2X1 U15699 ( .IN1(n8753), .IN2(n8250), .Q(n15015) );
  AND2X1 U15700 ( .IN1(n15987), .IN2(WX11203), .Q(n15014) );
  AND2X1 U15701 ( .IN1(n9237), .IN2(CRC_OUT_1_20), .Q(n14998) );
  AND2X1 U15702 ( .IN1(DATA_0_20), .IN2(n9264), .Q(n14997) );
  OR4X1 U15703 ( .IN1(n15016), .IN2(n15017), .IN3(n15018), .IN4(n15019), .Q(
        WX11008) );
  AND2X1 U15704 ( .IN1(n1964), .IN2(n9211), .Q(n15019) );
  INVX0 U15705 ( .INP(n15020), .ZN(n1964) );
  OR2X1 U15706 ( .IN1(n9557), .IN2(n3807), .Q(n15020) );
  AND2X1 U15707 ( .IN1(n9968), .IN2(n9173), .Q(n15018) );
  AND2X1 U15708 ( .IN1(n15021), .IN2(n15022), .Q(n9968) );
  INVX0 U15709 ( .INP(n15023), .ZN(n15022) );
  AND2X1 U15710 ( .IN1(n15024), .IN2(n15025), .Q(n15023) );
  OR2X1 U15711 ( .IN1(n15025), .IN2(n15024), .Q(n15021) );
  OR2X1 U15712 ( .IN1(n15026), .IN2(n15027), .Q(n15024) );
  AND2X1 U15713 ( .IN1(n9451), .IN2(WX11073), .Q(n15027) );
  AND2X1 U15714 ( .IN1(n7902), .IN2(n9464), .Q(n15026) );
  AND2X1 U15715 ( .IN1(n15028), .IN2(n15029), .Q(n15025) );
  OR2X1 U15716 ( .IN1(n15030), .IN2(n8752), .Q(n15029) );
  OR2X1 U15717 ( .IN1(WX11201), .IN2(n15031), .Q(n15028) );
  INVX0 U15718 ( .INP(n15030), .ZN(n15031) );
  AND2X1 U15719 ( .IN1(n15032), .IN2(n15033), .Q(n15030) );
  OR2X1 U15720 ( .IN1(n8251), .IN2(test_so95), .Q(n15033) );
  OR2X1 U15721 ( .IN1(n9145), .IN2(n15988), .Q(n15032) );
  AND2X1 U15722 ( .IN1(n9237), .IN2(CRC_OUT_1_21), .Q(n15017) );
  AND2X1 U15723 ( .IN1(DATA_0_21), .IN2(n9262), .Q(n15016) );
  OR4X1 U15724 ( .IN1(n15034), .IN2(n15035), .IN3(n15036), .IN4(n15037), .Q(
        WX11006) );
  AND2X1 U15725 ( .IN1(n1963), .IN2(n9212), .Q(n15037) );
  INVX0 U15726 ( .INP(n15038), .ZN(n1963) );
  OR2X1 U15727 ( .IN1(n9557), .IN2(n3808), .Q(n15038) );
  AND2X1 U15728 ( .IN1(n9186), .IN2(n9975), .Q(n15036) );
  OR2X1 U15729 ( .IN1(n15039), .IN2(n15040), .Q(n9975) );
  INVX0 U15730 ( .INP(n15041), .ZN(n15040) );
  OR2X1 U15731 ( .IN1(n15042), .IN2(n15043), .Q(n15041) );
  AND2X1 U15732 ( .IN1(n15043), .IN2(n15042), .Q(n15039) );
  AND2X1 U15733 ( .IN1(n15044), .IN2(n15045), .Q(n15042) );
  OR2X1 U15734 ( .IN1(n9477), .IN2(n7903), .Q(n15045) );
  OR2X1 U15735 ( .IN1(WX11071), .IN2(n9442), .Q(n15044) );
  OR2X1 U15736 ( .IN1(n15046), .IN2(n15047), .Q(n15043) );
  INVX0 U15737 ( .INP(n15048), .ZN(n15047) );
  OR2X1 U15738 ( .IN1(n15049), .IN2(n7904), .Q(n15048) );
  AND2X1 U15739 ( .IN1(n7904), .IN2(n15049), .Q(n15046) );
  INVX0 U15740 ( .INP(n15050), .ZN(n15049) );
  OR2X1 U15741 ( .IN1(n15051), .IN2(n15052), .Q(n15050) );
  AND2X1 U15742 ( .IN1(n8751), .IN2(n8252), .Q(n15052) );
  AND2X1 U15743 ( .IN1(n15989), .IN2(WX11199), .Q(n15051) );
  AND2X1 U15744 ( .IN1(n9237), .IN2(CRC_OUT_1_22), .Q(n15035) );
  AND2X1 U15745 ( .IN1(DATA_0_22), .IN2(n9263), .Q(n15034) );
  OR4X1 U15746 ( .IN1(n15053), .IN2(n15054), .IN3(n15055), .IN4(n15056), .Q(
        WX11004) );
  AND2X1 U15747 ( .IN1(n1962), .IN2(n9212), .Q(n15056) );
  INVX0 U15748 ( .INP(n15057), .ZN(n1962) );
  OR2X1 U15749 ( .IN1(n9557), .IN2(n3809), .Q(n15057) );
  AND2X1 U15750 ( .IN1(n9982), .IN2(n9173), .Q(n15055) );
  AND2X1 U15751 ( .IN1(n15058), .IN2(n15059), .Q(n9982) );
  INVX0 U15752 ( .INP(n15060), .ZN(n15059) );
  AND2X1 U15753 ( .IN1(n15061), .IN2(n15062), .Q(n15060) );
  OR2X1 U15754 ( .IN1(n15062), .IN2(n15061), .Q(n15058) );
  OR2X1 U15755 ( .IN1(n15063), .IN2(n15064), .Q(n15061) );
  AND2X1 U15756 ( .IN1(n9451), .IN2(WX11133), .Q(n15064) );
  AND2X1 U15757 ( .IN1(n7905), .IN2(n9476), .Q(n15063) );
  AND2X1 U15758 ( .IN1(n15065), .IN2(n15066), .Q(n15062) );
  OR2X1 U15759 ( .IN1(n15067), .IN2(n8750), .Q(n15066) );
  OR2X1 U15760 ( .IN1(WX11197), .IN2(n15068), .Q(n15065) );
  INVX0 U15761 ( .INP(n15067), .ZN(n15068) );
  AND2X1 U15762 ( .IN1(n15069), .IN2(n15070), .Q(n15067) );
  OR2X1 U15763 ( .IN1(n8253), .IN2(test_so93), .Q(n15070) );
  OR2X1 U15764 ( .IN1(n9146), .IN2(n15990), .Q(n15069) );
  AND2X1 U15765 ( .IN1(n9237), .IN2(CRC_OUT_1_23), .Q(n15054) );
  AND2X1 U15766 ( .IN1(DATA_0_23), .IN2(n9261), .Q(n15053) );
  OR4X1 U15767 ( .IN1(n15071), .IN2(n15072), .IN3(n15073), .IN4(n15074), .Q(
        WX11002) );
  AND2X1 U15768 ( .IN1(n1961), .IN2(n9212), .Q(n15074) );
  INVX0 U15769 ( .INP(n15075), .ZN(n1961) );
  OR2X1 U15770 ( .IN1(n9557), .IN2(n3810), .Q(n15075) );
  AND2X1 U15771 ( .IN1(n9186), .IN2(n9989), .Q(n15073) );
  OR2X1 U15772 ( .IN1(n15076), .IN2(n15077), .Q(n9989) );
  INVX0 U15773 ( .INP(n15078), .ZN(n15077) );
  OR2X1 U15774 ( .IN1(n15079), .IN2(n15080), .Q(n15078) );
  AND2X1 U15775 ( .IN1(n15080), .IN2(n15079), .Q(n15076) );
  AND2X1 U15776 ( .IN1(n15081), .IN2(n15082), .Q(n15079) );
  OR2X1 U15777 ( .IN1(n9478), .IN2(n7906), .Q(n15082) );
  OR2X1 U15778 ( .IN1(WX11067), .IN2(n9442), .Q(n15081) );
  OR2X1 U15779 ( .IN1(n15083), .IN2(n15084), .Q(n15080) );
  INVX0 U15780 ( .INP(n15085), .ZN(n15084) );
  OR2X1 U15781 ( .IN1(n15086), .IN2(n7907), .Q(n15085) );
  AND2X1 U15782 ( .IN1(n7907), .IN2(n15086), .Q(n15083) );
  INVX0 U15783 ( .INP(n15087), .ZN(n15086) );
  OR2X1 U15784 ( .IN1(n15088), .IN2(n15089), .Q(n15087) );
  AND2X1 U15785 ( .IN1(n8749), .IN2(n8254), .Q(n15089) );
  AND2X1 U15786 ( .IN1(n15991), .IN2(WX11195), .Q(n15088) );
  AND2X1 U15787 ( .IN1(n9238), .IN2(CRC_OUT_1_24), .Q(n15072) );
  AND2X1 U15788 ( .IN1(DATA_0_24), .IN2(n9262), .Q(n15071) );
  OR4X1 U15789 ( .IN1(n15090), .IN2(n15091), .IN3(n15092), .IN4(n15093), .Q(
        WX11000) );
  AND2X1 U15790 ( .IN1(n1960), .IN2(n9212), .Q(n15093) );
  INVX0 U15791 ( .INP(n15094), .ZN(n1960) );
  OR2X1 U15792 ( .IN1(n9557), .IN2(n3811), .Q(n15094) );
  AND2X1 U15793 ( .IN1(n9996), .IN2(n9173), .Q(n15092) );
  AND2X1 U15794 ( .IN1(n15095), .IN2(n15096), .Q(n9996) );
  OR2X1 U15795 ( .IN1(n15097), .IN2(n15098), .Q(n15096) );
  INVX0 U15796 ( .INP(n15099), .ZN(n15095) );
  AND2X1 U15797 ( .IN1(n15098), .IN2(n15097), .Q(n15099) );
  INVX0 U15798 ( .INP(n15100), .ZN(n15097) );
  OR2X1 U15799 ( .IN1(n15101), .IN2(n15102), .Q(n15100) );
  AND2X1 U15800 ( .IN1(n9451), .IN2(WX11193), .Q(n15102) );
  AND2X1 U15801 ( .IN1(n8748), .IN2(n9461), .Q(n15101) );
  OR2X1 U15802 ( .IN1(n15103), .IN2(n15104), .Q(n15098) );
  AND3X1 U15803 ( .IN1(n15105), .IN2(n15106), .IN3(n7909), .Q(n15104) );
  OR2X1 U15804 ( .IN1(n7908), .IN2(n9097), .Q(n15106) );
  OR2X1 U15805 ( .IN1(test_so91), .IN2(WX11065), .Q(n15105) );
  AND2X1 U15806 ( .IN1(n15107), .IN2(WX11129), .Q(n15103) );
  OR2X1 U15807 ( .IN1(n15108), .IN2(n15109), .Q(n15107) );
  AND2X1 U15808 ( .IN1(n7908), .IN2(n9097), .Q(n15109) );
  AND2X1 U15809 ( .IN1(test_so91), .IN2(WX11065), .Q(n15108) );
  AND2X1 U15810 ( .IN1(n9238), .IN2(CRC_OUT_1_25), .Q(n15091) );
  AND2X1 U15811 ( .IN1(DATA_0_25), .IN2(n9263), .Q(n15090) );
  OR4X1 U15812 ( .IN1(n15110), .IN2(n15111), .IN3(n15112), .IN4(n15113), .Q(
        WX10998) );
  AND2X1 U15813 ( .IN1(n1959), .IN2(n9212), .Q(n15113) );
  INVX0 U15814 ( .INP(n15114), .ZN(n1959) );
  OR2X1 U15815 ( .IN1(n9557), .IN2(n3812), .Q(n15114) );
  AND2X1 U15816 ( .IN1(n9186), .IN2(n10003), .Q(n15112) );
  OR2X1 U15817 ( .IN1(n15115), .IN2(n15116), .Q(n10003) );
  INVX0 U15818 ( .INP(n15117), .ZN(n15116) );
  OR2X1 U15819 ( .IN1(n15118), .IN2(n15119), .Q(n15117) );
  AND2X1 U15820 ( .IN1(n15119), .IN2(n15118), .Q(n15115) );
  AND2X1 U15821 ( .IN1(n15120), .IN2(n15121), .Q(n15118) );
  OR2X1 U15822 ( .IN1(n9479), .IN2(n7910), .Q(n15121) );
  OR2X1 U15823 ( .IN1(WX11063), .IN2(n9442), .Q(n15120) );
  OR2X1 U15824 ( .IN1(n15122), .IN2(n15123), .Q(n15119) );
  INVX0 U15825 ( .INP(n15124), .ZN(n15123) );
  OR2X1 U15826 ( .IN1(n15125), .IN2(n7911), .Q(n15124) );
  AND2X1 U15827 ( .IN1(n7911), .IN2(n15125), .Q(n15122) );
  INVX0 U15828 ( .INP(n15126), .ZN(n15125) );
  OR2X1 U15829 ( .IN1(n15127), .IN2(n15128), .Q(n15126) );
  AND2X1 U15830 ( .IN1(n8747), .IN2(n8257), .Q(n15128) );
  AND2X1 U15831 ( .IN1(n15992), .IN2(WX11191), .Q(n15127) );
  AND2X1 U15832 ( .IN1(n9238), .IN2(CRC_OUT_1_26), .Q(n15111) );
  AND2X1 U15833 ( .IN1(DATA_0_26), .IN2(n9263), .Q(n15110) );
  OR4X1 U15834 ( .IN1(n15129), .IN2(n15130), .IN3(n15131), .IN4(n15132), .Q(
        WX10996) );
  AND2X1 U15835 ( .IN1(n1958), .IN2(n9212), .Q(n15132) );
  INVX0 U15836 ( .INP(n15133), .ZN(n1958) );
  OR2X1 U15837 ( .IN1(n9557), .IN2(n3813), .Q(n15133) );
  AND2X1 U15838 ( .IN1(n9186), .IN2(n10010), .Q(n15131) );
  OR2X1 U15839 ( .IN1(n15134), .IN2(n15135), .Q(n10010) );
  INVX0 U15840 ( .INP(n15136), .ZN(n15135) );
  OR2X1 U15841 ( .IN1(n15137), .IN2(n15138), .Q(n15136) );
  AND2X1 U15842 ( .IN1(n15138), .IN2(n15137), .Q(n15134) );
  AND2X1 U15843 ( .IN1(n15139), .IN2(n15140), .Q(n15137) );
  OR2X1 U15844 ( .IN1(n9479), .IN2(n7912), .Q(n15140) );
  OR2X1 U15845 ( .IN1(WX11061), .IN2(n9442), .Q(n15139) );
  OR2X1 U15846 ( .IN1(n15141), .IN2(n15142), .Q(n15138) );
  INVX0 U15847 ( .INP(n15143), .ZN(n15142) );
  OR2X1 U15848 ( .IN1(n15144), .IN2(n7913), .Q(n15143) );
  AND2X1 U15849 ( .IN1(n7913), .IN2(n15144), .Q(n15141) );
  INVX0 U15850 ( .INP(n15145), .ZN(n15144) );
  OR2X1 U15851 ( .IN1(n15146), .IN2(n15147), .Q(n15145) );
  AND2X1 U15852 ( .IN1(n8746), .IN2(n8258), .Q(n15147) );
  AND2X1 U15853 ( .IN1(n15993), .IN2(WX11189), .Q(n15146) );
  AND2X1 U15854 ( .IN1(n9238), .IN2(CRC_OUT_1_27), .Q(n15130) );
  AND2X1 U15855 ( .IN1(DATA_0_27), .IN2(n9262), .Q(n15129) );
  OR4X1 U15856 ( .IN1(n15148), .IN2(n15149), .IN3(n15150), .IN4(n15151), .Q(
        WX10994) );
  AND2X1 U15857 ( .IN1(n1957), .IN2(n9212), .Q(n15151) );
  INVX0 U15858 ( .INP(n15152), .ZN(n1957) );
  OR2X1 U15859 ( .IN1(n9557), .IN2(n3814), .Q(n15152) );
  AND2X1 U15860 ( .IN1(n9186), .IN2(n10017), .Q(n15150) );
  OR2X1 U15861 ( .IN1(n15153), .IN2(n15154), .Q(n10017) );
  INVX0 U15862 ( .INP(n15155), .ZN(n15154) );
  OR2X1 U15863 ( .IN1(n15156), .IN2(n15157), .Q(n15155) );
  AND2X1 U15864 ( .IN1(n15157), .IN2(n15156), .Q(n15153) );
  AND2X1 U15865 ( .IN1(n15158), .IN2(n15159), .Q(n15156) );
  OR2X1 U15866 ( .IN1(n9480), .IN2(n7914), .Q(n15159) );
  OR2X1 U15867 ( .IN1(WX11059), .IN2(n9442), .Q(n15158) );
  OR2X1 U15868 ( .IN1(n15160), .IN2(n15161), .Q(n15157) );
  INVX0 U15869 ( .INP(n15162), .ZN(n15161) );
  OR2X1 U15870 ( .IN1(n15163), .IN2(n7915), .Q(n15162) );
  AND2X1 U15871 ( .IN1(n7915), .IN2(n15163), .Q(n15160) );
  INVX0 U15872 ( .INP(n15164), .ZN(n15163) );
  OR2X1 U15873 ( .IN1(n15165), .IN2(n15166), .Q(n15164) );
  AND2X1 U15874 ( .IN1(n8745), .IN2(n8259), .Q(n15166) );
  AND2X1 U15875 ( .IN1(n15994), .IN2(WX11187), .Q(n15165) );
  AND2X1 U15876 ( .IN1(n9238), .IN2(CRC_OUT_1_28), .Q(n15149) );
  AND2X1 U15877 ( .IN1(DATA_0_28), .IN2(n9261), .Q(n15148) );
  OR4X1 U15878 ( .IN1(n15167), .IN2(n15168), .IN3(n15169), .IN4(n15170), .Q(
        WX10992) );
  AND2X1 U15879 ( .IN1(n1956), .IN2(n9201), .Q(n15170) );
  INVX0 U15880 ( .INP(n15171), .ZN(n1956) );
  OR2X1 U15881 ( .IN1(n9557), .IN2(n3815), .Q(n15171) );
  AND2X1 U15882 ( .IN1(n9185), .IN2(n10024), .Q(n15169) );
  OR2X1 U15883 ( .IN1(n15172), .IN2(n15173), .Q(n10024) );
  INVX0 U15884 ( .INP(n15174), .ZN(n15173) );
  OR2X1 U15885 ( .IN1(n15175), .IN2(n15176), .Q(n15174) );
  AND2X1 U15886 ( .IN1(n15176), .IN2(n15175), .Q(n15172) );
  AND2X1 U15887 ( .IN1(n15177), .IN2(n15178), .Q(n15175) );
  OR2X1 U15888 ( .IN1(n9480), .IN2(n7916), .Q(n15178) );
  OR2X1 U15889 ( .IN1(WX11057), .IN2(n9442), .Q(n15177) );
  OR2X1 U15890 ( .IN1(n15179), .IN2(n15180), .Q(n15176) );
  INVX0 U15891 ( .INP(n15181), .ZN(n15180) );
  OR2X1 U15892 ( .IN1(n15182), .IN2(n7917), .Q(n15181) );
  AND2X1 U15893 ( .IN1(n7917), .IN2(n15182), .Q(n15179) );
  INVX0 U15894 ( .INP(n15183), .ZN(n15182) );
  OR2X1 U15895 ( .IN1(n15184), .IN2(n15185), .Q(n15183) );
  AND2X1 U15896 ( .IN1(n8744), .IN2(n8260), .Q(n15185) );
  AND2X1 U15897 ( .IN1(n15995), .IN2(WX11185), .Q(n15184) );
  AND2X1 U15898 ( .IN1(n9238), .IN2(CRC_OUT_1_29), .Q(n15168) );
  AND2X1 U15899 ( .IN1(DATA_0_29), .IN2(n9261), .Q(n15167) );
  OR4X1 U15900 ( .IN1(n15186), .IN2(n15187), .IN3(n15188), .IN4(n15189), .Q(
        WX10990) );
  AND2X1 U15901 ( .IN1(n1955), .IN2(n9212), .Q(n15189) );
  AND2X1 U15902 ( .IN1(TM0), .IN2(n9450), .Q(n2148) );
  INVX0 U15903 ( .INP(n15190), .ZN(n1955) );
  OR2X1 U15904 ( .IN1(n9557), .IN2(n3816), .Q(n15190) );
  AND2X1 U15905 ( .IN1(n9190), .IN2(n10031), .Q(n15188) );
  OR2X1 U15906 ( .IN1(n15191), .IN2(n15192), .Q(n10031) );
  INVX0 U15907 ( .INP(n15193), .ZN(n15192) );
  OR2X1 U15908 ( .IN1(n15194), .IN2(n15195), .Q(n15193) );
  AND2X1 U15909 ( .IN1(n15195), .IN2(n15194), .Q(n15191) );
  AND2X1 U15910 ( .IN1(n15196), .IN2(n15197), .Q(n15194) );
  OR2X1 U15911 ( .IN1(n9459), .IN2(n7918), .Q(n15197) );
  OR2X1 U15912 ( .IN1(WX11055), .IN2(n9442), .Q(n15196) );
  OR2X1 U15913 ( .IN1(n15198), .IN2(n15199), .Q(n15195) );
  INVX0 U15914 ( .INP(n15200), .ZN(n15199) );
  OR2X1 U15915 ( .IN1(n15201), .IN2(n7919), .Q(n15200) );
  AND2X1 U15916 ( .IN1(n7919), .IN2(n15201), .Q(n15198) );
  INVX0 U15917 ( .INP(n15202), .ZN(n15201) );
  OR2X1 U15918 ( .IN1(n15203), .IN2(n15204), .Q(n15202) );
  AND2X1 U15919 ( .IN1(n8743), .IN2(n8261), .Q(n15204) );
  AND2X1 U15920 ( .IN1(n15996), .IN2(WX11183), .Q(n15203) );
  AND2X1 U15921 ( .IN1(n9238), .IN2(CRC_OUT_1_30), .Q(n15187) );
  AND2X1 U15922 ( .IN1(DATA_0_30), .IN2(n9261), .Q(n15186) );
  OR4X1 U15923 ( .IN1(n15205), .IN2(n15206), .IN3(n15207), .IN4(n15208), .Q(
        WX10988) );
  AND2X1 U15924 ( .IN1(DATA_0_31), .IN2(n9259), .Q(n15208) );
  AND2X1 U15925 ( .IN1(n9179), .IN2(n10038), .Q(n15207) );
  OR2X1 U15926 ( .IN1(n15209), .IN2(n15210), .Q(n10038) );
  INVX0 U15927 ( .INP(n15211), .ZN(n15210) );
  OR2X1 U15928 ( .IN1(n15212), .IN2(n15213), .Q(n15211) );
  AND2X1 U15929 ( .IN1(n15213), .IN2(n15212), .Q(n15209) );
  AND2X1 U15930 ( .IN1(n15214), .IN2(n15215), .Q(n15212) );
  OR2X1 U15931 ( .IN1(n9460), .IN2(n7876), .Q(n15215) );
  OR2X1 U15932 ( .IN1(WX11053), .IN2(n9442), .Q(n15214) );
  OR2X1 U15933 ( .IN1(n15216), .IN2(n15217), .Q(n15213) );
  INVX0 U15934 ( .INP(n15218), .ZN(n15217) );
  OR2X1 U15935 ( .IN1(n15219), .IN2(n7877), .Q(n15218) );
  AND2X1 U15936 ( .IN1(n7877), .IN2(n15219), .Q(n15216) );
  INVX0 U15937 ( .INP(n15220), .ZN(n15219) );
  OR2X1 U15938 ( .IN1(n15221), .IN2(n15222), .Q(n15220) );
  AND2X1 U15939 ( .IN1(n8742), .IN2(n8262), .Q(n15222) );
  AND2X1 U15940 ( .IN1(n15997), .IN2(WX11181), .Q(n15221) );
  AND3X1 U15941 ( .IN1(n2199), .IN2(n9513), .IN3(n9440), .Q(n9821) );
  AND2X1 U15942 ( .IN1(n2245), .IN2(WX10829), .Q(n15206) );
  AND2X1 U15943 ( .IN1(test_so100), .IN2(n9228), .Q(n15205) );
  AND2X1 U15944 ( .IN1(n9052), .IN2(n9498), .Q(WX10890) );
  AND2X1 U15945 ( .IN1(n15223), .IN2(n9498), .Q(WX10377) );
  OR2X1 U15946 ( .IN1(n15224), .IN2(n15225), .Q(n15223) );
  AND2X1 U15947 ( .IN1(DFF_1534_n1), .IN2(n9110), .Q(n15225) );
  AND2X1 U15948 ( .IN1(test_so85), .IN2(CRC_OUT_2_30), .Q(n15224) );
  AND3X1 U15949 ( .IN1(n15226), .IN2(n15227), .IN3(n9519), .Q(WX10375) );
  OR2X1 U15950 ( .IN1(DFF_1533_n1), .IN2(WX9890), .Q(n15227) );
  OR2X1 U15951 ( .IN1(n8768), .IN2(CRC_OUT_2_29), .Q(n15226) );
  AND3X1 U15952 ( .IN1(n15228), .IN2(n15229), .IN3(n9519), .Q(WX10373) );
  OR2X1 U15953 ( .IN1(DFF_1532_n1), .IN2(WX9892), .Q(n15229) );
  OR2X1 U15954 ( .IN1(n8769), .IN2(CRC_OUT_2_28), .Q(n15228) );
  AND3X1 U15955 ( .IN1(n15230), .IN2(n15231), .IN3(n9519), .Q(WX10371) );
  OR2X1 U15956 ( .IN1(DFF_1531_n1), .IN2(WX9894), .Q(n15231) );
  OR2X1 U15957 ( .IN1(n8770), .IN2(CRC_OUT_2_27), .Q(n15230) );
  AND3X1 U15958 ( .IN1(n15232), .IN2(n15233), .IN3(n9519), .Q(WX10369) );
  OR2X1 U15959 ( .IN1(DFF_1530_n1), .IN2(WX9896), .Q(n15233) );
  OR2X1 U15960 ( .IN1(n8771), .IN2(CRC_OUT_2_26), .Q(n15232) );
  AND3X1 U15961 ( .IN1(n15234), .IN2(n15235), .IN3(n9519), .Q(WX10367) );
  OR2X1 U15962 ( .IN1(DFF_1529_n1), .IN2(WX9898), .Q(n15235) );
  OR2X1 U15963 ( .IN1(n8772), .IN2(CRC_OUT_2_25), .Q(n15234) );
  AND3X1 U15964 ( .IN1(n15236), .IN2(n15237), .IN3(n9519), .Q(WX10365) );
  OR2X1 U15965 ( .IN1(DFF_1528_n1), .IN2(WX9900), .Q(n15237) );
  OR2X1 U15966 ( .IN1(n8773), .IN2(CRC_OUT_2_24), .Q(n15236) );
  AND3X1 U15967 ( .IN1(n15238), .IN2(n15239), .IN3(n9519), .Q(WX10363) );
  OR2X1 U15968 ( .IN1(DFF_1527_n1), .IN2(WX9902), .Q(n15239) );
  OR2X1 U15969 ( .IN1(n8774), .IN2(CRC_OUT_2_23), .Q(n15238) );
  AND3X1 U15970 ( .IN1(n15240), .IN2(n15241), .IN3(n9518), .Q(WX10361) );
  OR2X1 U15971 ( .IN1(DFF_1526_n1), .IN2(WX9904), .Q(n15241) );
  OR2X1 U15972 ( .IN1(n8775), .IN2(CRC_OUT_2_22), .Q(n15240) );
  AND3X1 U15973 ( .IN1(n15242), .IN2(n15243), .IN3(n9518), .Q(WX10359) );
  OR2X1 U15974 ( .IN1(DFF_1525_n1), .IN2(WX9906), .Q(n15243) );
  OR2X1 U15975 ( .IN1(n8776), .IN2(CRC_OUT_2_21), .Q(n15242) );
  AND3X1 U15976 ( .IN1(n15244), .IN2(n15245), .IN3(n9518), .Q(WX10357) );
  OR2X1 U15977 ( .IN1(DFF_1524_n1), .IN2(WX9908), .Q(n15245) );
  OR2X1 U15978 ( .IN1(n8777), .IN2(CRC_OUT_2_20), .Q(n15244) );
  AND2X1 U15979 ( .IN1(n15246), .IN2(n9498), .Q(WX10355) );
  OR2X1 U15980 ( .IN1(n15247), .IN2(n15248), .Q(n15246) );
  AND2X1 U15981 ( .IN1(n8778), .IN2(n9164), .Q(n15248) );
  AND2X1 U15982 ( .IN1(test_so88), .IN2(WX9910), .Q(n15247) );
  AND3X1 U15983 ( .IN1(n15249), .IN2(n15250), .IN3(n9518), .Q(WX10353) );
  OR2X1 U15984 ( .IN1(DFF_1522_n1), .IN2(WX9912), .Q(n15250) );
  OR2X1 U15985 ( .IN1(n8779), .IN2(CRC_OUT_2_18), .Q(n15249) );
  AND3X1 U15986 ( .IN1(n15251), .IN2(n15252), .IN3(n9518), .Q(WX10351) );
  OR2X1 U15987 ( .IN1(DFF_1521_n1), .IN2(WX9914), .Q(n15252) );
  OR2X1 U15988 ( .IN1(n8780), .IN2(CRC_OUT_2_17), .Q(n15251) );
  AND3X1 U15989 ( .IN1(n15253), .IN2(n15254), .IN3(n9518), .Q(WX10349) );
  OR2X1 U15990 ( .IN1(DFF_1520_n1), .IN2(WX9916), .Q(n15254) );
  OR2X1 U15991 ( .IN1(n8781), .IN2(CRC_OUT_2_16), .Q(n15253) );
  AND2X1 U15992 ( .IN1(n15255), .IN2(n9498), .Q(WX10347) );
  OR2X1 U15993 ( .IN1(n15256), .IN2(n15257), .Q(n15255) );
  AND2X1 U15994 ( .IN1(n15258), .IN2(CRC_OUT_2_15), .Q(n15257) );
  INVX0 U15995 ( .INP(n15259), .ZN(n15258) );
  AND2X1 U15996 ( .IN1(DFF_1519_n1), .IN2(n15259), .Q(n15256) );
  AND2X1 U15997 ( .IN1(n15260), .IN2(n15261), .Q(n15259) );
  OR2X1 U15998 ( .IN1(CRC_OUT_2_31), .IN2(n8716), .Q(n15261) );
  OR2X1 U15999 ( .IN1(WX9918), .IN2(DFF_1535_n1), .Q(n15260) );
  AND3X1 U16000 ( .IN1(n15262), .IN2(n15263), .IN3(n9518), .Q(WX10345) );
  OR2X1 U16001 ( .IN1(DFF_1518_n1), .IN2(WX9920), .Q(n15263) );
  OR2X1 U16002 ( .IN1(n8782), .IN2(CRC_OUT_2_14), .Q(n15262) );
  AND2X1 U16003 ( .IN1(n15264), .IN2(n9497), .Q(WX10343) );
  OR2X1 U16004 ( .IN1(n15265), .IN2(n15266), .Q(n15264) );
  AND2X1 U16005 ( .IN1(DFF_1517_n1), .IN2(n9103), .Q(n15266) );
  AND2X1 U16006 ( .IN1(test_so86), .IN2(CRC_OUT_2_13), .Q(n15265) );
  AND3X1 U16007 ( .IN1(n15267), .IN2(n15268), .IN3(n9518), .Q(WX10341) );
  OR2X1 U16008 ( .IN1(DFF_1516_n1), .IN2(WX9924), .Q(n15268) );
  OR2X1 U16009 ( .IN1(n8783), .IN2(CRC_OUT_2_12), .Q(n15267) );
  AND3X1 U16010 ( .IN1(n15269), .IN2(n15270), .IN3(n9518), .Q(WX10339) );
  OR2X1 U16011 ( .IN1(DFF_1515_n1), .IN2(WX9926), .Q(n15270) );
  OR2X1 U16012 ( .IN1(n8784), .IN2(CRC_OUT_2_11), .Q(n15269) );
  AND2X1 U16013 ( .IN1(n15271), .IN2(n9498), .Q(WX10337) );
  OR2X1 U16014 ( .IN1(n15272), .IN2(n15273), .Q(n15271) );
  AND2X1 U16015 ( .IN1(n15274), .IN2(CRC_OUT_2_10), .Q(n15273) );
  AND2X1 U16016 ( .IN1(DFF_1514_n1), .IN2(n15275), .Q(n15272) );
  INVX0 U16017 ( .INP(n15274), .ZN(n15275) );
  OR2X1 U16018 ( .IN1(n15276), .IN2(n15277), .Q(n15274) );
  AND2X1 U16019 ( .IN1(DFF_1535_n1), .IN2(WX9928), .Q(n15277) );
  AND2X1 U16020 ( .IN1(n8717), .IN2(CRC_OUT_2_31), .Q(n15276) );
  AND3X1 U16021 ( .IN1(n15278), .IN2(n15279), .IN3(n9518), .Q(WX10335) );
  OR2X1 U16022 ( .IN1(DFF_1513_n1), .IN2(WX9930), .Q(n15279) );
  OR2X1 U16023 ( .IN1(n8785), .IN2(CRC_OUT_2_9), .Q(n15278) );
  AND3X1 U16024 ( .IN1(n15280), .IN2(n15281), .IN3(n9518), .Q(WX10333) );
  OR2X1 U16025 ( .IN1(DFF_1512_n1), .IN2(WX9932), .Q(n15281) );
  OR2X1 U16026 ( .IN1(n8786), .IN2(CRC_OUT_2_8), .Q(n15280) );
  AND3X1 U16027 ( .IN1(n15282), .IN2(n15283), .IN3(n9518), .Q(WX10331) );
  OR2X1 U16028 ( .IN1(DFF_1511_n1), .IN2(WX9934), .Q(n15283) );
  OR2X1 U16029 ( .IN1(n8787), .IN2(CRC_OUT_2_7), .Q(n15282) );
  AND3X1 U16030 ( .IN1(n15284), .IN2(n15285), .IN3(n9517), .Q(WX10329) );
  OR2X1 U16031 ( .IN1(DFF_1510_n1), .IN2(WX9936), .Q(n15285) );
  OR2X1 U16032 ( .IN1(n8788), .IN2(CRC_OUT_2_6), .Q(n15284) );
  AND3X1 U16033 ( .IN1(n15286), .IN2(n15287), .IN3(n9517), .Q(WX10327) );
  OR2X1 U16034 ( .IN1(DFF_1509_n1), .IN2(WX9938), .Q(n15287) );
  OR2X1 U16035 ( .IN1(n8789), .IN2(CRC_OUT_2_5), .Q(n15286) );
  AND3X1 U16036 ( .IN1(n15288), .IN2(n15289), .IN3(n9517), .Q(WX10325) );
  OR2X1 U16037 ( .IN1(DFF_1508_n1), .IN2(WX9940), .Q(n15289) );
  OR2X1 U16038 ( .IN1(n8790), .IN2(CRC_OUT_2_4), .Q(n15288) );
  AND2X1 U16039 ( .IN1(n15290), .IN2(n9497), .Q(WX10323) );
  OR2X1 U16040 ( .IN1(n15291), .IN2(n15292), .Q(n15290) );
  AND2X1 U16041 ( .IN1(n15293), .IN2(CRC_OUT_2_3), .Q(n15292) );
  AND2X1 U16042 ( .IN1(DFF_1507_n1), .IN2(n15294), .Q(n15291) );
  INVX0 U16043 ( .INP(n15293), .ZN(n15294) );
  OR2X1 U16044 ( .IN1(n15295), .IN2(n15296), .Q(n15293) );
  AND2X1 U16045 ( .IN1(DFF_1535_n1), .IN2(WX9942), .Q(n15296) );
  AND2X1 U16046 ( .IN1(n8718), .IN2(CRC_OUT_2_31), .Q(n15295) );
  AND2X1 U16047 ( .IN1(n15297), .IN2(n9497), .Q(WX10321) );
  OR2X1 U16048 ( .IN1(n15298), .IN2(n15299), .Q(n15297) );
  AND2X1 U16049 ( .IN1(n8791), .IN2(n9165), .Q(n15299) );
  AND2X1 U16050 ( .IN1(test_so87), .IN2(WX9944), .Q(n15298) );
  AND3X1 U16051 ( .IN1(n15300), .IN2(n15301), .IN3(n9525), .Q(WX10319) );
  OR2X1 U16052 ( .IN1(DFF_1505_n1), .IN2(WX9946), .Q(n15301) );
  OR2X1 U16053 ( .IN1(n8792), .IN2(CRC_OUT_2_1), .Q(n15300) );
  AND3X1 U16054 ( .IN1(n15302), .IN2(n15303), .IN3(n9513), .Q(WX10317) );
  OR2X1 U16055 ( .IN1(DFF_1504_n1), .IN2(WX9948), .Q(n15303) );
  OR2X1 U16056 ( .IN1(n8793), .IN2(CRC_OUT_2_0), .Q(n15302) );
  AND3X1 U16057 ( .IN1(n15304), .IN2(n15305), .IN3(n9517), .Q(WX10315) );
  OR2X1 U16058 ( .IN1(DFF_1535_n1), .IN2(WX9950), .Q(n15305) );
  OR2X1 U16059 ( .IN1(n8735), .IN2(CRC_OUT_2_31), .Q(n15304) );
  OR2X1 U16060 ( .IN1(n15306), .IN2(n15307), .Q(DATA_9_9) );
  AND2X1 U16061 ( .IN1(n11409), .IN2(n15308), .Q(n15307) );
  INVX0 U16062 ( .INP(n15309), .ZN(n15306) );
  OR2X1 U16063 ( .IN1(n15308), .IN2(n11409), .Q(n15309) );
  OR2X1 U16064 ( .IN1(n15310), .IN2(n15311), .Q(n11409) );
  INVX0 U16065 ( .INP(n15312), .ZN(n15311) );
  OR2X1 U16066 ( .IN1(n15313), .IN2(n15314), .Q(n15312) );
  AND2X1 U16067 ( .IN1(n15314), .IN2(n15313), .Q(n15310) );
  AND2X1 U16068 ( .IN1(n15315), .IN2(n15316), .Q(n15313) );
  OR2X1 U16069 ( .IN1(n2199), .IN2(n3485), .Q(n15316) );
  OR2X1 U16070 ( .IN1(WX689), .IN2(TM0), .Q(n15315) );
  INVX0 U16071 ( .INP(n15317), .ZN(n15314) );
  AND2X1 U16072 ( .IN1(n15318), .IN2(n15319), .Q(n15317) );
  OR2X1 U16073 ( .IN1(n15320), .IN2(n8996), .Q(n15319) );
  INVX0 U16074 ( .INP(n15321), .ZN(n15318) );
  AND2X1 U16075 ( .IN1(n8996), .IN2(n15320), .Q(n15321) );
  AND2X1 U16076 ( .IN1(n15322), .IN2(n15323), .Q(n15320) );
  OR2X1 U16077 ( .IN1(WX817), .IN2(n8998), .Q(n15323) );
  OR2X1 U16078 ( .IN1(WX881), .IN2(n8997), .Q(n15322) );
  OR2X1 U16079 ( .IN1(n9084), .IN2(n2199), .Q(n15308) );
  OR2X1 U16080 ( .IN1(n15324), .IN2(n15325), .Q(DATA_9_8) );
  AND2X1 U16081 ( .IN1(n11403), .IN2(n15326), .Q(n15325) );
  INVX0 U16082 ( .INP(n15327), .ZN(n15324) );
  OR2X1 U16083 ( .IN1(n15326), .IN2(n11403), .Q(n15327) );
  OR2X1 U16084 ( .IN1(n15328), .IN2(n15329), .Q(n11403) );
  INVX0 U16085 ( .INP(n15330), .ZN(n15329) );
  OR2X1 U16086 ( .IN1(n15331), .IN2(n15332), .Q(n15330) );
  AND2X1 U16087 ( .IN1(n15332), .IN2(n15331), .Q(n15328) );
  AND2X1 U16088 ( .IN1(n15333), .IN2(n15334), .Q(n15331) );
  OR2X1 U16089 ( .IN1(n2199), .IN2(n3483), .Q(n15334) );
  OR2X1 U16090 ( .IN1(WX691), .IN2(TM0), .Q(n15333) );
  OR2X1 U16091 ( .IN1(n15335), .IN2(n15336), .Q(n15332) );
  AND3X1 U16092 ( .IN1(n15337), .IN2(n15338), .IN3(n9008), .Q(n15336) );
  OR2X1 U16093 ( .IN1(n9006), .IN2(WX883), .Q(n15338) );
  OR2X1 U16094 ( .IN1(n9007), .IN2(WX819), .Q(n15337) );
  AND2X1 U16095 ( .IN1(n15339), .IN2(WX755), .Q(n15335) );
  OR2X1 U16096 ( .IN1(n15340), .IN2(n15341), .Q(n15339) );
  AND2X1 U16097 ( .IN1(n9006), .IN2(WX883), .Q(n15341) );
  AND2X1 U16098 ( .IN1(n9007), .IN2(WX819), .Q(n15340) );
  OR2X1 U16099 ( .IN1(n9083), .IN2(n2199), .Q(n15326) );
  OR2X1 U16100 ( .IN1(n15342), .IN2(n15343), .Q(DATA_9_7) );
  AND2X1 U16101 ( .IN1(n11397), .IN2(n15344), .Q(n15343) );
  INVX0 U16102 ( .INP(n15345), .ZN(n15342) );
  OR2X1 U16103 ( .IN1(n15344), .IN2(n11397), .Q(n15345) );
  OR2X1 U16104 ( .IN1(n15346), .IN2(n15347), .Q(n11397) );
  INVX0 U16105 ( .INP(n15348), .ZN(n15347) );
  OR2X1 U16106 ( .IN1(n15349), .IN2(n15350), .Q(n15348) );
  AND2X1 U16107 ( .IN1(n15350), .IN2(n15349), .Q(n15346) );
  AND2X1 U16108 ( .IN1(n15351), .IN2(n15352), .Q(n15349) );
  OR2X1 U16109 ( .IN1(n2199), .IN2(n3481), .Q(n15352) );
  OR2X1 U16110 ( .IN1(WX693), .IN2(TM0), .Q(n15351) );
  INVX0 U16111 ( .INP(n15353), .ZN(n15350) );
  AND2X1 U16112 ( .IN1(n15354), .IN2(n15355), .Q(n15353) );
  OR2X1 U16113 ( .IN1(n15356), .IN2(n9036), .Q(n15355) );
  INVX0 U16114 ( .INP(n15357), .ZN(n15354) );
  AND2X1 U16115 ( .IN1(n9036), .IN2(n15356), .Q(n15357) );
  AND2X1 U16116 ( .IN1(n15358), .IN2(n15359), .Q(n15356) );
  OR2X1 U16117 ( .IN1(WX821), .IN2(n9038), .Q(n15359) );
  OR2X1 U16118 ( .IN1(WX885), .IN2(n9037), .Q(n15358) );
  OR2X1 U16119 ( .IN1(n9082), .IN2(n2199), .Q(n15344) );
  OR2X1 U16120 ( .IN1(n15360), .IN2(n15361), .Q(DATA_9_6) );
  INVX0 U16121 ( .INP(n15362), .ZN(n15361) );
  OR3X1 U16122 ( .IN1(n2199), .IN2(n9081), .IN3(n11391), .Q(n15362) );
  AND2X1 U16123 ( .IN1(n11391), .IN2(n15363), .Q(n15360) );
  OR2X1 U16124 ( .IN1(n9081), .IN2(n2199), .Q(n15363) );
  AND2X1 U16125 ( .IN1(n15364), .IN2(n15365), .Q(n11391) );
  INVX0 U16126 ( .INP(n15366), .ZN(n15365) );
  AND2X1 U16127 ( .IN1(n15367), .IN2(n15368), .Q(n15366) );
  OR2X1 U16128 ( .IN1(n15368), .IN2(n15367), .Q(n15364) );
  OR2X1 U16129 ( .IN1(n15369), .IN2(n15370), .Q(n15367) );
  AND2X1 U16130 ( .IN1(TM0), .IN2(WX695), .Q(n15370) );
  AND2X1 U16131 ( .IN1(n3479), .IN2(n2199), .Q(n15369) );
  AND2X1 U16132 ( .IN1(n15371), .IN2(n15372), .Q(n15368) );
  OR2X1 U16133 ( .IN1(n15373), .IN2(n9024), .Q(n15372) );
  INVX0 U16134 ( .INP(n15374), .ZN(n15371) );
  AND2X1 U16135 ( .IN1(n9024), .IN2(n15373), .Q(n15374) );
  AND2X1 U16136 ( .IN1(n15375), .IN2(n15376), .Q(n15373) );
  OR2X1 U16137 ( .IN1(WX887), .IN2(test_so5), .Q(n15376) );
  OR2X1 U16138 ( .IN1(n9147), .IN2(n9025), .Q(n15375) );
  OR2X1 U16139 ( .IN1(n15377), .IN2(n15378), .Q(DATA_9_5) );
  AND2X1 U16140 ( .IN1(n11385), .IN2(n15379), .Q(n15378) );
  INVX0 U16141 ( .INP(n15380), .ZN(n15377) );
  OR2X1 U16142 ( .IN1(n15379), .IN2(n11385), .Q(n15380) );
  OR2X1 U16143 ( .IN1(n15381), .IN2(n15382), .Q(n11385) );
  INVX0 U16144 ( .INP(n15383), .ZN(n15382) );
  OR2X1 U16145 ( .IN1(n15384), .IN2(n15385), .Q(n15383) );
  AND2X1 U16146 ( .IN1(n15385), .IN2(n15384), .Q(n15381) );
  AND2X1 U16147 ( .IN1(n15386), .IN2(n15387), .Q(n15384) );
  OR2X1 U16148 ( .IN1(n2199), .IN2(n3477), .Q(n15387) );
  OR2X1 U16149 ( .IN1(WX697), .IN2(TM0), .Q(n15386) );
  OR2X1 U16150 ( .IN1(n15388), .IN2(n15389), .Q(n15385) );
  AND3X1 U16151 ( .IN1(n15390), .IN2(n15391), .IN3(n9011), .Q(n15389) );
  OR2X1 U16152 ( .IN1(n9009), .IN2(WX889), .Q(n15391) );
  OR2X1 U16153 ( .IN1(n9010), .IN2(WX825), .Q(n15390) );
  AND2X1 U16154 ( .IN1(n15392), .IN2(WX761), .Q(n15388) );
  OR2X1 U16155 ( .IN1(n15393), .IN2(n15394), .Q(n15392) );
  AND2X1 U16156 ( .IN1(n9009), .IN2(WX889), .Q(n15394) );
  AND2X1 U16157 ( .IN1(n9010), .IN2(WX825), .Q(n15393) );
  OR2X1 U16158 ( .IN1(n9080), .IN2(n2199), .Q(n15379) );
  OR2X1 U16159 ( .IN1(n15395), .IN2(n15396), .Q(DATA_9_4) );
  AND2X1 U16160 ( .IN1(n11379), .IN2(n15397), .Q(n15396) );
  INVX0 U16161 ( .INP(n15398), .ZN(n15395) );
  OR2X1 U16162 ( .IN1(n15397), .IN2(n11379), .Q(n15398) );
  OR2X1 U16163 ( .IN1(n15399), .IN2(n15400), .Q(n11379) );
  INVX0 U16164 ( .INP(n15401), .ZN(n15400) );
  OR2X1 U16165 ( .IN1(n15402), .IN2(n15403), .Q(n15401) );
  AND2X1 U16166 ( .IN1(n15403), .IN2(n15402), .Q(n15399) );
  AND2X1 U16167 ( .IN1(n15404), .IN2(n15405), .Q(n15402) );
  OR2X1 U16168 ( .IN1(n2199), .IN2(n3475), .Q(n15405) );
  OR2X1 U16169 ( .IN1(WX699), .IN2(TM0), .Q(n15404) );
  OR2X1 U16170 ( .IN1(n15406), .IN2(n15407), .Q(n15403) );
  AND3X1 U16171 ( .IN1(n15408), .IN2(n15409), .IN3(n9014), .Q(n15407) );
  OR2X1 U16172 ( .IN1(n9012), .IN2(WX891), .Q(n15409) );
  OR2X1 U16173 ( .IN1(n9013), .IN2(WX827), .Q(n15408) );
  AND2X1 U16174 ( .IN1(n15410), .IN2(WX763), .Q(n15406) );
  OR2X1 U16175 ( .IN1(n15411), .IN2(n15412), .Q(n15410) );
  AND2X1 U16176 ( .IN1(n9012), .IN2(WX891), .Q(n15412) );
  AND2X1 U16177 ( .IN1(n9013), .IN2(WX827), .Q(n15411) );
  OR2X1 U16178 ( .IN1(n9079), .IN2(n2199), .Q(n15397) );
  OR2X1 U16179 ( .IN1(n15413), .IN2(n15414), .Q(DATA_9_31) );
  AND2X1 U16180 ( .IN1(n11617), .IN2(n15415), .Q(n15414) );
  INVX0 U16181 ( .INP(n15416), .ZN(n15413) );
  OR2X1 U16182 ( .IN1(n15415), .IN2(n11617), .Q(n15416) );
  OR2X1 U16183 ( .IN1(n15417), .IN2(n15418), .Q(n11617) );
  INVX0 U16184 ( .INP(n15419), .ZN(n15418) );
  OR2X1 U16185 ( .IN1(n15420), .IN2(n15421), .Q(n15419) );
  AND2X1 U16186 ( .IN1(n15421), .IN2(n15420), .Q(n15417) );
  AND2X1 U16187 ( .IN1(n15422), .IN2(n15423), .Q(n15420) );
  OR2X1 U16188 ( .IN1(n9462), .IN2(n3529), .Q(n15423) );
  OR2X1 U16189 ( .IN1(WX645), .IN2(n9442), .Q(n15422) );
  INVX0 U16190 ( .INP(n15424), .ZN(n15421) );
  AND2X1 U16191 ( .IN1(n15425), .IN2(n15426), .Q(n15424) );
  OR2X1 U16192 ( .IN1(n15427), .IN2(n9028), .Q(n15426) );
  INVX0 U16193 ( .INP(n15428), .ZN(n15425) );
  AND2X1 U16194 ( .IN1(n9028), .IN2(n15427), .Q(n15428) );
  AND2X1 U16195 ( .IN1(n15429), .IN2(n15430), .Q(n15427) );
  OR2X1 U16196 ( .IN1(WX773), .IN2(n9030), .Q(n15430) );
  OR2X1 U16197 ( .IN1(WX837), .IN2(n9029), .Q(n15429) );
  OR2X1 U16198 ( .IN1(n9078), .IN2(n2199), .Q(n15415) );
  OR2X1 U16199 ( .IN1(n15431), .IN2(n15432), .Q(DATA_9_30) );
  AND2X1 U16200 ( .IN1(n11581), .IN2(n15433), .Q(n15432) );
  INVX0 U16201 ( .INP(n15434), .ZN(n15431) );
  OR2X1 U16202 ( .IN1(n15433), .IN2(n11581), .Q(n15434) );
  OR2X1 U16203 ( .IN1(n15435), .IN2(n15436), .Q(n11581) );
  INVX0 U16204 ( .INP(n15437), .ZN(n15436) );
  OR2X1 U16205 ( .IN1(n15438), .IN2(n15439), .Q(n15437) );
  AND2X1 U16206 ( .IN1(n15439), .IN2(n15438), .Q(n15435) );
  AND2X1 U16207 ( .IN1(n15440), .IN2(n15441), .Q(n15438) );
  OR2X1 U16208 ( .IN1(n9463), .IN2(n3527), .Q(n15441) );
  OR2X1 U16209 ( .IN1(WX647), .IN2(n9441), .Q(n15440) );
  INVX0 U16210 ( .INP(n15442), .ZN(n15439) );
  AND2X1 U16211 ( .IN1(n15443), .IN2(n15444), .Q(n15442) );
  OR2X1 U16212 ( .IN1(n15445), .IN2(n8954), .Q(n15444) );
  INVX0 U16213 ( .INP(n15446), .ZN(n15443) );
  AND2X1 U16214 ( .IN1(n8954), .IN2(n15445), .Q(n15446) );
  AND2X1 U16215 ( .IN1(n15447), .IN2(n15448), .Q(n15445) );
  OR2X1 U16216 ( .IN1(WX775), .IN2(n8956), .Q(n15448) );
  OR2X1 U16217 ( .IN1(WX839), .IN2(n8955), .Q(n15447) );
  OR2X1 U16218 ( .IN1(n9077), .IN2(n2199), .Q(n15433) );
  OR2X1 U16219 ( .IN1(n15449), .IN2(n15450), .Q(DATA_9_3) );
  AND2X1 U16220 ( .IN1(n11373), .IN2(n15451), .Q(n15450) );
  INVX0 U16221 ( .INP(n15452), .ZN(n15449) );
  OR2X1 U16222 ( .IN1(n15451), .IN2(n11373), .Q(n15452) );
  OR2X1 U16223 ( .IN1(n15453), .IN2(n15454), .Q(n11373) );
  INVX0 U16224 ( .INP(n15455), .ZN(n15454) );
  OR2X1 U16225 ( .IN1(n15456), .IN2(n15457), .Q(n15455) );
  AND2X1 U16226 ( .IN1(n15457), .IN2(n15456), .Q(n15453) );
  AND2X1 U16227 ( .IN1(n15458), .IN2(n15459), .Q(n15456) );
  OR2X1 U16228 ( .IN1(n2199), .IN2(n3473), .Q(n15459) );
  OR2X1 U16229 ( .IN1(WX701), .IN2(TM0), .Q(n15458) );
  OR2X1 U16230 ( .IN1(n15460), .IN2(n15461), .Q(n15457) );
  AND3X1 U16231 ( .IN1(n15462), .IN2(n15463), .IN3(n8959), .Q(n15461) );
  OR2X1 U16232 ( .IN1(n8957), .IN2(WX893), .Q(n15463) );
  OR2X1 U16233 ( .IN1(n8958), .IN2(WX829), .Q(n15462) );
  AND2X1 U16234 ( .IN1(n15464), .IN2(WX765), .Q(n15460) );
  OR2X1 U16235 ( .IN1(n15465), .IN2(n15466), .Q(n15464) );
  AND2X1 U16236 ( .IN1(n8957), .IN2(WX893), .Q(n15466) );
  AND2X1 U16237 ( .IN1(n8958), .IN2(WX829), .Q(n15465) );
  OR2X1 U16238 ( .IN1(n9076), .IN2(n2199), .Q(n15451) );
  OR2X1 U16239 ( .IN1(n15467), .IN2(n15468), .Q(DATA_9_29) );
  AND2X1 U16240 ( .IN1(n11549), .IN2(n15469), .Q(n15468) );
  INVX0 U16241 ( .INP(n15470), .ZN(n15467) );
  OR2X1 U16242 ( .IN1(n15469), .IN2(n11549), .Q(n15470) );
  OR2X1 U16243 ( .IN1(n15471), .IN2(n15472), .Q(n11549) );
  INVX0 U16244 ( .INP(n15473), .ZN(n15472) );
  OR2X1 U16245 ( .IN1(n15474), .IN2(n15475), .Q(n15473) );
  AND2X1 U16246 ( .IN1(n15475), .IN2(n15474), .Q(n15471) );
  AND2X1 U16247 ( .IN1(n15476), .IN2(n15477), .Q(n15474) );
  OR2X1 U16248 ( .IN1(n9465), .IN2(n3525), .Q(n15477) );
  OR2X1 U16249 ( .IN1(WX649), .IN2(n9441), .Q(n15476) );
  OR2X1 U16250 ( .IN1(n15478), .IN2(n15479), .Q(n15475) );
  AND3X1 U16251 ( .IN1(n15480), .IN2(n15481), .IN3(n8965), .Q(n15479) );
  OR2X1 U16252 ( .IN1(n8963), .IN2(WX841), .Q(n15481) );
  OR2X1 U16253 ( .IN1(n8964), .IN2(WX777), .Q(n15480) );
  AND2X1 U16254 ( .IN1(n15482), .IN2(WX713), .Q(n15478) );
  OR2X1 U16255 ( .IN1(n15483), .IN2(n15484), .Q(n15482) );
  AND2X1 U16256 ( .IN1(n8963), .IN2(WX841), .Q(n15484) );
  AND2X1 U16257 ( .IN1(n8964), .IN2(WX777), .Q(n15483) );
  OR2X1 U16258 ( .IN1(n9075), .IN2(n2199), .Q(n15469) );
  OR2X1 U16259 ( .IN1(n15485), .IN2(n15486), .Q(DATA_9_28) );
  INVX0 U16260 ( .INP(n15487), .ZN(n15486) );
  OR3X1 U16261 ( .IN1(n2199), .IN2(n9074), .IN3(n11523), .Q(n15487) );
  AND2X1 U16262 ( .IN1(n11523), .IN2(n15488), .Q(n15485) );
  OR2X1 U16263 ( .IN1(n9074), .IN2(n2199), .Q(n15488) );
  AND2X1 U16264 ( .IN1(n15489), .IN2(n15490), .Q(n11523) );
  INVX0 U16265 ( .INP(n15491), .ZN(n15490) );
  AND2X1 U16266 ( .IN1(n15492), .IN2(n15493), .Q(n15491) );
  OR2X1 U16267 ( .IN1(n15493), .IN2(n15492), .Q(n15489) );
  OR2X1 U16268 ( .IN1(n15494), .IN2(n15495), .Q(n15492) );
  AND2X1 U16269 ( .IN1(n9451), .IN2(WX779), .Q(n15495) );
  AND2X1 U16270 ( .IN1(n8972), .IN2(n9478), .Q(n15494) );
  AND2X1 U16271 ( .IN1(n15496), .IN2(n15497), .Q(n15493) );
  INVX0 U16272 ( .INP(n15498), .ZN(n15497) );
  AND2X1 U16273 ( .IN1(n15499), .IN2(WX843), .Q(n15498) );
  OR2X1 U16274 ( .IN1(WX843), .IN2(n15499), .Q(n15496) );
  OR2X1 U16275 ( .IN1(n15500), .IN2(n15501), .Q(n15499) );
  AND2X1 U16276 ( .IN1(n8974), .IN2(n9166), .Q(n15501) );
  AND2X1 U16277 ( .IN1(test_so2), .IN2(WX715), .Q(n15500) );
  OR2X1 U16278 ( .IN1(n15502), .IN2(n15503), .Q(DATA_9_27) );
  AND2X1 U16279 ( .IN1(n11517), .IN2(n15504), .Q(n15503) );
  INVX0 U16280 ( .INP(n15505), .ZN(n15502) );
  OR2X1 U16281 ( .IN1(n15504), .IN2(n11517), .Q(n15505) );
  OR2X1 U16282 ( .IN1(n15506), .IN2(n15507), .Q(n11517) );
  INVX0 U16283 ( .INP(n15508), .ZN(n15507) );
  OR2X1 U16284 ( .IN1(n15509), .IN2(n15510), .Q(n15508) );
  AND2X1 U16285 ( .IN1(n15510), .IN2(n15509), .Q(n15506) );
  AND2X1 U16286 ( .IN1(n15511), .IN2(n15512), .Q(n15509) );
  OR2X1 U16287 ( .IN1(n9467), .IN2(n3521), .Q(n15512) );
  OR2X1 U16288 ( .IN1(WX653), .IN2(n9441), .Q(n15511) );
  OR2X1 U16289 ( .IN1(n15513), .IN2(n15514), .Q(n15510) );
  AND3X1 U16290 ( .IN1(n15515), .IN2(n15516), .IN3(n8980), .Q(n15514) );
  OR2X1 U16291 ( .IN1(n8978), .IN2(WX845), .Q(n15516) );
  OR2X1 U16292 ( .IN1(n8979), .IN2(WX781), .Q(n15515) );
  AND2X1 U16293 ( .IN1(n15517), .IN2(WX717), .Q(n15513) );
  OR2X1 U16294 ( .IN1(n15518), .IN2(n15519), .Q(n15517) );
  AND2X1 U16295 ( .IN1(n8978), .IN2(WX845), .Q(n15519) );
  AND2X1 U16296 ( .IN1(n8979), .IN2(WX781), .Q(n15518) );
  OR2X1 U16297 ( .IN1(n9073), .IN2(n2199), .Q(n15504) );
  OR2X1 U16298 ( .IN1(n15520), .IN2(n15521), .Q(DATA_9_26) );
  AND2X1 U16299 ( .IN1(n11511), .IN2(n15522), .Q(n15521) );
  INVX0 U16300 ( .INP(n15523), .ZN(n15520) );
  OR2X1 U16301 ( .IN1(n15522), .IN2(n11511), .Q(n15523) );
  OR2X1 U16302 ( .IN1(n15524), .IN2(n15525), .Q(n11511) );
  INVX0 U16303 ( .INP(n15526), .ZN(n15525) );
  OR2X1 U16304 ( .IN1(n15527), .IN2(n15528), .Q(n15526) );
  AND2X1 U16305 ( .IN1(n15528), .IN2(n15527), .Q(n15524) );
  AND2X1 U16306 ( .IN1(n15529), .IN2(n15530), .Q(n15527) );
  OR2X1 U16307 ( .IN1(n9468), .IN2(n3519), .Q(n15530) );
  OR2X1 U16308 ( .IN1(WX655), .IN2(n9441), .Q(n15529) );
  OR2X1 U16309 ( .IN1(n15531), .IN2(n15532), .Q(n15528) );
  AND3X1 U16310 ( .IN1(n15533), .IN2(n15534), .IN3(n8983), .Q(n15532) );
  OR2X1 U16311 ( .IN1(n8981), .IN2(WX847), .Q(n15534) );
  OR2X1 U16312 ( .IN1(n8982), .IN2(WX783), .Q(n15533) );
  AND2X1 U16313 ( .IN1(n15535), .IN2(WX719), .Q(n15531) );
  OR2X1 U16314 ( .IN1(n15536), .IN2(n15537), .Q(n15535) );
  AND2X1 U16315 ( .IN1(n8981), .IN2(WX847), .Q(n15537) );
  AND2X1 U16316 ( .IN1(n8982), .IN2(WX783), .Q(n15536) );
  OR2X1 U16317 ( .IN1(n9072), .IN2(n2199), .Q(n15522) );
  OR2X1 U16318 ( .IN1(n15538), .IN2(n15539), .Q(DATA_9_25) );
  AND2X1 U16319 ( .IN1(n11505), .IN2(n15540), .Q(n15539) );
  INVX0 U16320 ( .INP(n15541), .ZN(n15538) );
  OR2X1 U16321 ( .IN1(n15540), .IN2(n11505), .Q(n15541) );
  OR2X1 U16322 ( .IN1(n15542), .IN2(n15543), .Q(n11505) );
  INVX0 U16323 ( .INP(n15544), .ZN(n15543) );
  OR2X1 U16324 ( .IN1(n15545), .IN2(n15546), .Q(n15544) );
  AND2X1 U16325 ( .IN1(n15546), .IN2(n15545), .Q(n15542) );
  AND2X1 U16326 ( .IN1(n15547), .IN2(n15548), .Q(n15545) );
  OR2X1 U16327 ( .IN1(n9470), .IN2(n3517), .Q(n15548) );
  OR2X1 U16328 ( .IN1(WX657), .IN2(n9441), .Q(n15547) );
  OR2X1 U16329 ( .IN1(n15549), .IN2(n15550), .Q(n15546) );
  AND3X1 U16330 ( .IN1(n15551), .IN2(n15552), .IN3(n8992), .Q(n15550) );
  OR2X1 U16331 ( .IN1(n8990), .IN2(WX849), .Q(n15552) );
  OR2X1 U16332 ( .IN1(n8991), .IN2(WX785), .Q(n15551) );
  AND2X1 U16333 ( .IN1(n15553), .IN2(WX721), .Q(n15549) );
  OR2X1 U16334 ( .IN1(n15554), .IN2(n15555), .Q(n15553) );
  AND2X1 U16335 ( .IN1(n8990), .IN2(WX849), .Q(n15555) );
  AND2X1 U16336 ( .IN1(n8991), .IN2(WX785), .Q(n15554) );
  OR2X1 U16337 ( .IN1(n9071), .IN2(n2199), .Q(n15540) );
  OR2X1 U16338 ( .IN1(n15556), .IN2(n15557), .Q(DATA_9_24) );
  INVX0 U16339 ( .INP(n15558), .ZN(n15557) );
  OR3X1 U16340 ( .IN1(n2199), .IN2(n9070), .IN3(n11499), .Q(n15558) );
  AND2X1 U16341 ( .IN1(n11499), .IN2(n15559), .Q(n15556) );
  OR2X1 U16342 ( .IN1(n9070), .IN2(n2199), .Q(n15559) );
  AND2X1 U16343 ( .IN1(n15560), .IN2(n15561), .Q(n11499) );
  INVX0 U16344 ( .INP(n15562), .ZN(n15561) );
  AND2X1 U16345 ( .IN1(n15563), .IN2(n15564), .Q(n15562) );
  OR2X1 U16346 ( .IN1(n15564), .IN2(n15563), .Q(n15560) );
  OR2X1 U16347 ( .IN1(n15565), .IN2(n15566), .Q(n15563) );
  AND2X1 U16348 ( .IN1(n9451), .IN2(WX659), .Q(n15566) );
  AND2X1 U16349 ( .IN1(n3515), .IN2(n9480), .Q(n15565) );
  AND2X1 U16350 ( .IN1(n15567), .IN2(n15568), .Q(n15564) );
  OR2X1 U16351 ( .IN1(n15569), .IN2(n8999), .Q(n15568) );
  INVX0 U16352 ( .INP(n15570), .ZN(n15567) );
  AND2X1 U16353 ( .IN1(n8999), .IN2(n15569), .Q(n15570) );
  AND2X1 U16354 ( .IN1(n15571), .IN2(n15572), .Q(n15569) );
  OR2X1 U16355 ( .IN1(WX851), .IN2(test_so4), .Q(n15572) );
  OR2X1 U16356 ( .IN1(n9148), .IN2(n9000), .Q(n15571) );
  OR2X1 U16357 ( .IN1(n15573), .IN2(n15574), .Q(DATA_9_23) );
  AND2X1 U16358 ( .IN1(n11493), .IN2(n15575), .Q(n15574) );
  INVX0 U16359 ( .INP(n15576), .ZN(n15573) );
  OR2X1 U16360 ( .IN1(n15575), .IN2(n11493), .Q(n15576) );
  OR2X1 U16361 ( .IN1(n15577), .IN2(n15578), .Q(n11493) );
  INVX0 U16362 ( .INP(n15579), .ZN(n15578) );
  OR2X1 U16363 ( .IN1(n15580), .IN2(n15581), .Q(n15579) );
  AND2X1 U16364 ( .IN1(n15581), .IN2(n15580), .Q(n15577) );
  AND2X1 U16365 ( .IN1(n15582), .IN2(n15583), .Q(n15580) );
  OR2X1 U16366 ( .IN1(n9473), .IN2(n3513), .Q(n15583) );
  OR2X1 U16367 ( .IN1(WX661), .IN2(n9441), .Q(n15582) );
  OR2X1 U16368 ( .IN1(n15584), .IN2(n15585), .Q(n15581) );
  AND3X1 U16369 ( .IN1(n15586), .IN2(n15587), .IN3(n9003), .Q(n15585) );
  OR2X1 U16370 ( .IN1(n9001), .IN2(WX853), .Q(n15587) );
  OR2X1 U16371 ( .IN1(n9002), .IN2(WX789), .Q(n15586) );
  AND2X1 U16372 ( .IN1(n15588), .IN2(WX725), .Q(n15584) );
  OR2X1 U16373 ( .IN1(n15589), .IN2(n15590), .Q(n15588) );
  AND2X1 U16374 ( .IN1(n9001), .IN2(WX853), .Q(n15590) );
  AND2X1 U16375 ( .IN1(n9002), .IN2(WX789), .Q(n15589) );
  OR2X1 U16376 ( .IN1(n9069), .IN2(n2199), .Q(n15575) );
  OR2X1 U16377 ( .IN1(n15591), .IN2(n15592), .Q(DATA_9_22) );
  AND2X1 U16378 ( .IN1(n11487), .IN2(n15593), .Q(n15592) );
  INVX0 U16379 ( .INP(n15594), .ZN(n15591) );
  OR2X1 U16380 ( .IN1(n15593), .IN2(n11487), .Q(n15594) );
  OR2X1 U16381 ( .IN1(n15595), .IN2(n15596), .Q(n11487) );
  INVX0 U16382 ( .INP(n15597), .ZN(n15596) );
  OR2X1 U16383 ( .IN1(n15598), .IN2(n15599), .Q(n15597) );
  AND2X1 U16384 ( .IN1(n15599), .IN2(n15598), .Q(n15595) );
  AND2X1 U16385 ( .IN1(n15600), .IN2(n15601), .Q(n15598) );
  OR2X1 U16386 ( .IN1(n9474), .IN2(n3511), .Q(n15601) );
  OR2X1 U16387 ( .IN1(WX663), .IN2(n9441), .Q(n15600) );
  INVX0 U16388 ( .INP(n15602), .ZN(n15599) );
  AND2X1 U16389 ( .IN1(n15603), .IN2(n15604), .Q(n15602) );
  OR2X1 U16390 ( .IN1(n15605), .IN2(n9015), .Q(n15604) );
  INVX0 U16391 ( .INP(n15606), .ZN(n15603) );
  AND2X1 U16392 ( .IN1(n9015), .IN2(n15605), .Q(n15606) );
  AND2X1 U16393 ( .IN1(n15607), .IN2(n15608), .Q(n15605) );
  OR2X1 U16394 ( .IN1(WX791), .IN2(n9017), .Q(n15608) );
  OR2X1 U16395 ( .IN1(WX855), .IN2(n9016), .Q(n15607) );
  OR2X1 U16396 ( .IN1(n9068), .IN2(n2199), .Q(n15593) );
  OR2X1 U16397 ( .IN1(n15609), .IN2(n15610), .Q(DATA_9_21) );
  AND2X1 U16398 ( .IN1(n11481), .IN2(n15611), .Q(n15610) );
  INVX0 U16399 ( .INP(n15612), .ZN(n15609) );
  OR2X1 U16400 ( .IN1(n15611), .IN2(n11481), .Q(n15612) );
  OR2X1 U16401 ( .IN1(n15613), .IN2(n15614), .Q(n11481) );
  INVX0 U16402 ( .INP(n15615), .ZN(n15614) );
  OR2X1 U16403 ( .IN1(n15616), .IN2(n15617), .Q(n15615) );
  AND2X1 U16404 ( .IN1(n15617), .IN2(n15616), .Q(n15613) );
  AND2X1 U16405 ( .IN1(n15618), .IN2(n15619), .Q(n15616) );
  OR2X1 U16406 ( .IN1(n9476), .IN2(n3509), .Q(n15619) );
  OR2X1 U16407 ( .IN1(WX665), .IN2(n9441), .Q(n15618) );
  INVX0 U16408 ( .INP(n15620), .ZN(n15617) );
  AND2X1 U16409 ( .IN1(n15621), .IN2(n15622), .Q(n15620) );
  OR2X1 U16410 ( .IN1(n15623), .IN2(n9021), .Q(n15622) );
  INVX0 U16411 ( .INP(n15624), .ZN(n15621) );
  AND2X1 U16412 ( .IN1(n9021), .IN2(n15623), .Q(n15624) );
  AND2X1 U16413 ( .IN1(n15625), .IN2(n15626), .Q(n15623) );
  OR2X1 U16414 ( .IN1(WX793), .IN2(n9023), .Q(n15626) );
  OR2X1 U16415 ( .IN1(WX857), .IN2(n9022), .Q(n15625) );
  OR2X1 U16416 ( .IN1(n9067), .IN2(n2199), .Q(n15611) );
  OR2X1 U16417 ( .IN1(n15627), .IN2(n15628), .Q(DATA_9_20) );
  AND2X1 U16418 ( .IN1(n11475), .IN2(n15629), .Q(n15628) );
  OR2X1 U16419 ( .IN1(n9066), .IN2(n2199), .Q(n15629) );
  INVX0 U16420 ( .INP(n15630), .ZN(n15627) );
  OR3X1 U16421 ( .IN1(n2199), .IN2(n9066), .IN3(n11475), .Q(n15630) );
  AND2X1 U16422 ( .IN1(n15631), .IN2(n15632), .Q(n11475) );
  OR2X1 U16423 ( .IN1(n15633), .IN2(n15634), .Q(n15632) );
  INVX0 U16424 ( .INP(n15635), .ZN(n15631) );
  AND2X1 U16425 ( .IN1(n15634), .IN2(n15633), .Q(n15635) );
  AND2X1 U16426 ( .IN1(n15636), .IN2(n15637), .Q(n15633) );
  OR2X1 U16427 ( .IN1(n9477), .IN2(n3507), .Q(n15637) );
  OR2X1 U16428 ( .IN1(WX667), .IN2(n9441), .Q(n15636) );
  OR2X1 U16429 ( .IN1(n15638), .IN2(n15639), .Q(n15634) );
  AND3X1 U16430 ( .IN1(n15640), .IN2(n15641), .IN3(n9027), .Q(n15639) );
  OR2X1 U16431 ( .IN1(n9026), .IN2(n9098), .Q(n15641) );
  OR2X1 U16432 ( .IN1(test_so6), .IN2(WX859), .Q(n15640) );
  AND2X1 U16433 ( .IN1(n15642), .IN2(WX731), .Q(n15638) );
  OR2X1 U16434 ( .IN1(n15643), .IN2(n15644), .Q(n15642) );
  AND2X1 U16435 ( .IN1(n9026), .IN2(n9098), .Q(n15644) );
  AND2X1 U16436 ( .IN1(test_so6), .IN2(WX859), .Q(n15643) );
  OR2X1 U16437 ( .IN1(n15645), .IN2(n15646), .Q(DATA_9_2) );
  INVX0 U16438 ( .INP(n15647), .ZN(n15646) );
  OR3X1 U16439 ( .IN1(n2199), .IN2(n9065), .IN3(n11367), .Q(n15647) );
  AND2X1 U16440 ( .IN1(n11367), .IN2(n15648), .Q(n15645) );
  OR2X1 U16441 ( .IN1(n9065), .IN2(n2199), .Q(n15648) );
  AND2X1 U16442 ( .IN1(n15649), .IN2(n15650), .Q(n11367) );
  INVX0 U16443 ( .INP(n15651), .ZN(n15650) );
  AND2X1 U16444 ( .IN1(n15652), .IN2(n15653), .Q(n15651) );
  OR2X1 U16445 ( .IN1(n15653), .IN2(n15652), .Q(n15649) );
  OR2X1 U16446 ( .IN1(n15654), .IN2(n15655), .Q(n15652) );
  AND2X1 U16447 ( .IN1(TM0), .IN2(WX703), .Q(n15655) );
  AND2X1 U16448 ( .IN1(n3471), .IN2(n2199), .Q(n15654) );
  AND2X1 U16449 ( .IN1(n15656), .IN2(n15657), .Q(n15653) );
  OR2X1 U16450 ( .IN1(n15658), .IN2(n9034), .Q(n15657) );
  INVX0 U16451 ( .INP(n15659), .ZN(n15656) );
  AND2X1 U16452 ( .IN1(n9034), .IN2(n15658), .Q(n15659) );
  AND2X1 U16453 ( .IN1(n15660), .IN2(n15661), .Q(n15658) );
  OR2X1 U16454 ( .IN1(WX895), .IN2(test_so7), .Q(n15661) );
  OR2X1 U16455 ( .IN1(n9149), .IN2(n9035), .Q(n15660) );
  OR2X1 U16456 ( .IN1(n15662), .IN2(n15663), .Q(DATA_9_19) );
  AND2X1 U16457 ( .IN1(n11469), .IN2(n15664), .Q(n15663) );
  INVX0 U16458 ( .INP(n15665), .ZN(n15662) );
  OR2X1 U16459 ( .IN1(n15664), .IN2(n11469), .Q(n15665) );
  OR2X1 U16460 ( .IN1(n15666), .IN2(n15667), .Q(n11469) );
  INVX0 U16461 ( .INP(n15668), .ZN(n15667) );
  OR2X1 U16462 ( .IN1(n15669), .IN2(n15670), .Q(n15668) );
  AND2X1 U16463 ( .IN1(n15670), .IN2(n15669), .Q(n15666) );
  AND2X1 U16464 ( .IN1(n15671), .IN2(n15672), .Q(n15669) );
  OR2X1 U16465 ( .IN1(n9479), .IN2(n3505), .Q(n15672) );
  OR2X1 U16466 ( .IN1(WX669), .IN2(n9441), .Q(n15671) );
  OR2X1 U16467 ( .IN1(n15673), .IN2(n15674), .Q(n15670) );
  AND3X1 U16468 ( .IN1(n15675), .IN2(n15676), .IN3(n8962), .Q(n15674) );
  OR2X1 U16469 ( .IN1(n8960), .IN2(WX861), .Q(n15676) );
  OR2X1 U16470 ( .IN1(n8961), .IN2(WX797), .Q(n15675) );
  AND2X1 U16471 ( .IN1(n15677), .IN2(WX733), .Q(n15673) );
  OR2X1 U16472 ( .IN1(n15678), .IN2(n15679), .Q(n15677) );
  AND2X1 U16473 ( .IN1(n8960), .IN2(WX861), .Q(n15679) );
  AND2X1 U16474 ( .IN1(n8961), .IN2(WX797), .Q(n15678) );
  OR2X1 U16475 ( .IN1(n9064), .IN2(n2199), .Q(n15664) );
  OR2X1 U16476 ( .IN1(n15680), .IN2(n15681), .Q(DATA_9_18) );
  AND2X1 U16477 ( .IN1(n11463), .IN2(n15682), .Q(n15681) );
  INVX0 U16478 ( .INP(n15683), .ZN(n15680) );
  OR2X1 U16479 ( .IN1(n15682), .IN2(n11463), .Q(n15683) );
  OR2X1 U16480 ( .IN1(n15684), .IN2(n15685), .Q(n11463) );
  INVX0 U16481 ( .INP(n15686), .ZN(n15685) );
  OR2X1 U16482 ( .IN1(n15687), .IN2(n15688), .Q(n15686) );
  AND2X1 U16483 ( .IN1(n15688), .IN2(n15687), .Q(n15684) );
  AND2X1 U16484 ( .IN1(n15689), .IN2(n15690), .Q(n15687) );
  OR2X1 U16485 ( .IN1(n9480), .IN2(n3503), .Q(n15690) );
  OR2X1 U16486 ( .IN1(WX671), .IN2(n9441), .Q(n15689) );
  OR2X1 U16487 ( .IN1(n15691), .IN2(n15692), .Q(n15688) );
  AND3X1 U16488 ( .IN1(n15693), .IN2(n15694), .IN3(n8977), .Q(n15692) );
  OR2X1 U16489 ( .IN1(n8975), .IN2(WX863), .Q(n15694) );
  OR2X1 U16490 ( .IN1(n8976), .IN2(WX799), .Q(n15693) );
  AND2X1 U16491 ( .IN1(n15695), .IN2(WX735), .Q(n15691) );
  OR2X1 U16492 ( .IN1(n15696), .IN2(n15697), .Q(n15695) );
  AND2X1 U16493 ( .IN1(n8975), .IN2(WX863), .Q(n15697) );
  AND2X1 U16494 ( .IN1(n8976), .IN2(WX799), .Q(n15696) );
  OR2X1 U16495 ( .IN1(n9063), .IN2(n2199), .Q(n15682) );
  OR2X1 U16496 ( .IN1(n15698), .IN2(n15699), .Q(DATA_9_17) );
  AND2X1 U16497 ( .IN1(n11457), .IN2(n15700), .Q(n15699) );
  INVX0 U16498 ( .INP(n15701), .ZN(n15698) );
  OR2X1 U16499 ( .IN1(n15700), .IN2(n11457), .Q(n15701) );
  OR2X1 U16500 ( .IN1(n15702), .IN2(n15703), .Q(n11457) );
  INVX0 U16501 ( .INP(n15704), .ZN(n15703) );
  OR2X1 U16502 ( .IN1(n15705), .IN2(n15706), .Q(n15704) );
  AND2X1 U16503 ( .IN1(n15706), .IN2(n15705), .Q(n15702) );
  AND2X1 U16504 ( .IN1(n15707), .IN2(n15708), .Q(n15705) );
  OR2X1 U16505 ( .IN1(n9482), .IN2(n3501), .Q(n15708) );
  OR2X1 U16506 ( .IN1(WX673), .IN2(n9441), .Q(n15707) );
  OR2X1 U16507 ( .IN1(n15709), .IN2(n15710), .Q(n15706) );
  AND3X1 U16508 ( .IN1(n15711), .IN2(n15712), .IN3(n8989), .Q(n15710) );
  OR2X1 U16509 ( .IN1(n8987), .IN2(WX865), .Q(n15712) );
  OR2X1 U16510 ( .IN1(n8988), .IN2(WX801), .Q(n15711) );
  AND2X1 U16511 ( .IN1(n15713), .IN2(WX737), .Q(n15709) );
  OR2X1 U16512 ( .IN1(n15714), .IN2(n15715), .Q(n15713) );
  AND2X1 U16513 ( .IN1(n8987), .IN2(WX865), .Q(n15715) );
  AND2X1 U16514 ( .IN1(n8988), .IN2(WX801), .Q(n15714) );
  OR2X1 U16515 ( .IN1(n9062), .IN2(n2199), .Q(n15700) );
  OR2X1 U16516 ( .IN1(n15716), .IN2(n15717), .Q(DATA_9_16) );
  AND2X1 U16517 ( .IN1(n11451), .IN2(n15718), .Q(n15717) );
  OR2X1 U16518 ( .IN1(n9061), .IN2(n2199), .Q(n15718) );
  INVX0 U16519 ( .INP(n15719), .ZN(n15716) );
  OR3X1 U16520 ( .IN1(n2199), .IN2(n9061), .IN3(n11451), .Q(n15719) );
  AND2X1 U16521 ( .IN1(n15720), .IN2(n15721), .Q(n11451) );
  OR2X1 U16522 ( .IN1(n15722), .IN2(n15723), .Q(n15721) );
  INVX0 U16523 ( .INP(n15724), .ZN(n15720) );
  AND2X1 U16524 ( .IN1(n15723), .IN2(n15722), .Q(n15724) );
  AND2X1 U16525 ( .IN1(n15725), .IN2(n15726), .Q(n15722) );
  OR2X1 U16526 ( .IN1(n9457), .IN2(n3499), .Q(n15726) );
  OR2X1 U16527 ( .IN1(WX675), .IN2(n9446), .Q(n15725) );
  OR2X1 U16528 ( .IN1(n15727), .IN2(n15728), .Q(n15723) );
  AND3X1 U16529 ( .IN1(n15729), .IN2(n15730), .IN3(n9005), .Q(n15728) );
  OR2X1 U16530 ( .IN1(n9004), .IN2(n9086), .Q(n15730) );
  OR2X1 U16531 ( .IN1(test_so8), .IN2(WX739), .Q(n15729) );
  AND2X1 U16532 ( .IN1(n15731), .IN2(WX803), .Q(n15727) );
  OR2X1 U16533 ( .IN1(n15732), .IN2(n15733), .Q(n15731) );
  AND2X1 U16534 ( .IN1(n9004), .IN2(n9086), .Q(n15733) );
  AND2X1 U16535 ( .IN1(test_so8), .IN2(WX739), .Q(n15732) );
  OR2X1 U16536 ( .IN1(n15734), .IN2(n15735), .Q(DATA_9_15) );
  AND2X1 U16537 ( .IN1(n11445), .IN2(n15736), .Q(n15735) );
  INVX0 U16538 ( .INP(n15737), .ZN(n15734) );
  OR2X1 U16539 ( .IN1(n15736), .IN2(n11445), .Q(n15737) );
  OR2X1 U16540 ( .IN1(n15738), .IN2(n15739), .Q(n11445) );
  INVX0 U16541 ( .INP(n15740), .ZN(n15739) );
  OR2X1 U16542 ( .IN1(n15741), .IN2(n15742), .Q(n15740) );
  AND2X1 U16543 ( .IN1(n15742), .IN2(n15741), .Q(n15738) );
  AND2X1 U16544 ( .IN1(n15743), .IN2(n15744), .Q(n15741) );
  OR2X1 U16545 ( .IN1(n2199), .IN2(n3497), .Q(n15744) );
  OR2X1 U16546 ( .IN1(WX677), .IN2(TM0), .Q(n15743) );
  INVX0 U16547 ( .INP(n15745), .ZN(n15742) );
  AND2X1 U16548 ( .IN1(n15746), .IN2(n15747), .Q(n15745) );
  OR2X1 U16549 ( .IN1(n15748), .IN2(n9018), .Q(n15747) );
  INVX0 U16550 ( .INP(n15749), .ZN(n15746) );
  AND2X1 U16551 ( .IN1(n9018), .IN2(n15748), .Q(n15749) );
  AND2X1 U16552 ( .IN1(n15750), .IN2(n15751), .Q(n15748) );
  OR2X1 U16553 ( .IN1(WX805), .IN2(n9020), .Q(n15751) );
  OR2X1 U16554 ( .IN1(WX869), .IN2(n9019), .Q(n15750) );
  OR2X1 U16555 ( .IN1(n9060), .IN2(n2199), .Q(n15736) );
  OR2X1 U16556 ( .IN1(n15752), .IN2(n15753), .Q(DATA_9_14) );
  AND2X1 U16557 ( .IN1(n11439), .IN2(n15754), .Q(n15753) );
  INVX0 U16558 ( .INP(n15755), .ZN(n15752) );
  OR2X1 U16559 ( .IN1(n15754), .IN2(n11439), .Q(n15755) );
  OR2X1 U16560 ( .IN1(n15756), .IN2(n15757), .Q(n11439) );
  INVX0 U16561 ( .INP(n15758), .ZN(n15757) );
  OR2X1 U16562 ( .IN1(n15759), .IN2(n15760), .Q(n15758) );
  AND2X1 U16563 ( .IN1(n15760), .IN2(n15759), .Q(n15756) );
  AND2X1 U16564 ( .IN1(n15761), .IN2(n15762), .Q(n15759) );
  OR2X1 U16565 ( .IN1(n2199), .IN2(n3495), .Q(n15762) );
  OR2X1 U16566 ( .IN1(WX679), .IN2(TM0), .Q(n15761) );
  OR2X1 U16567 ( .IN1(n15763), .IN2(n15764), .Q(n15760) );
  AND3X1 U16568 ( .IN1(n15765), .IN2(n15766), .IN3(n9033), .Q(n15764) );
  OR2X1 U16569 ( .IN1(n9031), .IN2(WX871), .Q(n15766) );
  OR2X1 U16570 ( .IN1(n9032), .IN2(WX807), .Q(n15765) );
  AND2X1 U16571 ( .IN1(n15767), .IN2(WX743), .Q(n15763) );
  OR2X1 U16572 ( .IN1(n15768), .IN2(n15769), .Q(n15767) );
  AND2X1 U16573 ( .IN1(n9031), .IN2(WX871), .Q(n15769) );
  AND2X1 U16574 ( .IN1(n9032), .IN2(WX807), .Q(n15768) );
  OR2X1 U16575 ( .IN1(n2199), .IN2(n9059), .Q(n15754) );
  OR2X1 U16576 ( .IN1(n15770), .IN2(n15771), .Q(DATA_9_13) );
  AND2X1 U16577 ( .IN1(n11433), .IN2(n15772), .Q(n15771) );
  INVX0 U16578 ( .INP(n15773), .ZN(n15770) );
  OR2X1 U16579 ( .IN1(n15772), .IN2(n11433), .Q(n15773) );
  OR2X1 U16580 ( .IN1(n15774), .IN2(n15775), .Q(n11433) );
  INVX0 U16581 ( .INP(n15776), .ZN(n15775) );
  OR2X1 U16582 ( .IN1(n15777), .IN2(n15778), .Q(n15776) );
  AND2X1 U16583 ( .IN1(n15778), .IN2(n15777), .Q(n15774) );
  AND2X1 U16584 ( .IN1(n15779), .IN2(n15780), .Q(n15777) );
  OR2X1 U16585 ( .IN1(n2199), .IN2(n3493), .Q(n15780) );
  OR2X1 U16586 ( .IN1(WX681), .IN2(TM0), .Q(n15779) );
  OR2X1 U16587 ( .IN1(n15781), .IN2(n15782), .Q(n15778) );
  AND3X1 U16588 ( .IN1(n15783), .IN2(n15784), .IN3(n8968), .Q(n15782) );
  OR2X1 U16589 ( .IN1(n8966), .IN2(WX873), .Q(n15784) );
  OR2X1 U16590 ( .IN1(n8967), .IN2(WX809), .Q(n15783) );
  AND2X1 U16591 ( .IN1(n15785), .IN2(WX745), .Q(n15781) );
  OR2X1 U16592 ( .IN1(n15786), .IN2(n15787), .Q(n15785) );
  AND2X1 U16593 ( .IN1(n8966), .IN2(WX873), .Q(n15787) );
  AND2X1 U16594 ( .IN1(n8967), .IN2(WX809), .Q(n15786) );
  OR2X1 U16595 ( .IN1(n9058), .IN2(n2199), .Q(n15772) );
  OR2X1 U16596 ( .IN1(n15788), .IN2(n15789), .Q(DATA_9_12) );
  AND2X1 U16597 ( .IN1(n11427), .IN2(n15790), .Q(n15789) );
  INVX0 U16598 ( .INP(n15791), .ZN(n15788) );
  OR2X1 U16599 ( .IN1(n15790), .IN2(n11427), .Q(n15791) );
  OR2X1 U16600 ( .IN1(n15792), .IN2(n15793), .Q(n11427) );
  INVX0 U16601 ( .INP(n15794), .ZN(n15793) );
  OR2X1 U16602 ( .IN1(n15795), .IN2(n15796), .Q(n15794) );
  AND2X1 U16603 ( .IN1(n15796), .IN2(n15795), .Q(n15792) );
  AND2X1 U16604 ( .IN1(n15797), .IN2(n15798), .Q(n15795) );
  OR2X1 U16605 ( .IN1(n2199), .IN2(n3491), .Q(n15798) );
  OR2X1 U16606 ( .IN1(WX683), .IN2(TM0), .Q(n15797) );
  OR2X1 U16607 ( .IN1(n15799), .IN2(n15800), .Q(n15796) );
  AND3X1 U16608 ( .IN1(n15801), .IN2(n15802), .IN3(n8995), .Q(n15800) );
  OR2X1 U16609 ( .IN1(n8993), .IN2(WX875), .Q(n15802) );
  OR2X1 U16610 ( .IN1(n8994), .IN2(WX811), .Q(n15801) );
  AND2X1 U16611 ( .IN1(n15803), .IN2(WX747), .Q(n15799) );
  OR2X1 U16612 ( .IN1(n15804), .IN2(n15805), .Q(n15803) );
  AND2X1 U16613 ( .IN1(n8993), .IN2(WX875), .Q(n15805) );
  AND2X1 U16614 ( .IN1(n8994), .IN2(WX811), .Q(n15804) );
  OR2X1 U16615 ( .IN1(n9057), .IN2(n2199), .Q(n15790) );
  OR2X1 U16616 ( .IN1(n15806), .IN2(n15807), .Q(DATA_9_11) );
  AND2X1 U16617 ( .IN1(n11421), .IN2(n15808), .Q(n15807) );
  INVX0 U16618 ( .INP(n15809), .ZN(n15806) );
  OR2X1 U16619 ( .IN1(n15808), .IN2(n11421), .Q(n15809) );
  OR2X1 U16620 ( .IN1(n15810), .IN2(n15811), .Q(n11421) );
  INVX0 U16621 ( .INP(n15812), .ZN(n15811) );
  OR2X1 U16622 ( .IN1(n15813), .IN2(n15814), .Q(n15812) );
  AND2X1 U16623 ( .IN1(n15814), .IN2(n15813), .Q(n15810) );
  AND2X1 U16624 ( .IN1(n15815), .IN2(n15816), .Q(n15813) );
  OR2X1 U16625 ( .IN1(n2199), .IN2(n3489), .Q(n15816) );
  OR2X1 U16626 ( .IN1(WX685), .IN2(TM0), .Q(n15815) );
  OR2X1 U16627 ( .IN1(n15817), .IN2(n15818), .Q(n15814) );
  AND3X1 U16628 ( .IN1(n15819), .IN2(n15820), .IN3(n9041), .Q(n15818) );
  OR2X1 U16629 ( .IN1(n9039), .IN2(WX877), .Q(n15820) );
  OR2X1 U16630 ( .IN1(n9040), .IN2(WX813), .Q(n15819) );
  AND2X1 U16631 ( .IN1(n15821), .IN2(WX749), .Q(n15817) );
  OR2X1 U16632 ( .IN1(n15822), .IN2(n15823), .Q(n15821) );
  AND2X1 U16633 ( .IN1(n9039), .IN2(WX877), .Q(n15823) );
  AND2X1 U16634 ( .IN1(n9040), .IN2(WX813), .Q(n15822) );
  OR2X1 U16635 ( .IN1(n9056), .IN2(n2199), .Q(n15808) );
  OR2X1 U16636 ( .IN1(n15824), .IN2(n15825), .Q(DATA_9_10) );
  INVX0 U16637 ( .INP(n15826), .ZN(n15825) );
  OR3X1 U16638 ( .IN1(n2199), .IN2(n9055), .IN3(n11415), .Q(n15826) );
  AND2X1 U16639 ( .IN1(n11415), .IN2(n15827), .Q(n15824) );
  OR2X1 U16640 ( .IN1(n9055), .IN2(n2199), .Q(n15827) );
  AND2X1 U16641 ( .IN1(n15828), .IN2(n15829), .Q(n11415) );
  INVX0 U16642 ( .INP(n15830), .ZN(n15829) );
  AND2X1 U16643 ( .IN1(n15831), .IN2(n15832), .Q(n15830) );
  OR2X1 U16644 ( .IN1(n15832), .IN2(n15831), .Q(n15828) );
  OR2X1 U16645 ( .IN1(n15833), .IN2(n15834), .Q(n15831) );
  AND2X1 U16646 ( .IN1(TM0), .IN2(WX815), .Q(n15834) );
  AND2X1 U16647 ( .IN1(n8984), .IN2(n2199), .Q(n15833) );
  AND2X1 U16648 ( .IN1(n15835), .IN2(n15836), .Q(n15832) );
  INVX0 U16649 ( .INP(n15837), .ZN(n15836) );
  AND2X1 U16650 ( .IN1(n15838), .IN2(WX879), .Q(n15837) );
  OR2X1 U16651 ( .IN1(WX879), .IN2(n15838), .Q(n15835) );
  OR2X1 U16652 ( .IN1(n15839), .IN2(n15840), .Q(n15838) );
  AND2X1 U16653 ( .IN1(n8986), .IN2(n9167), .Q(n15840) );
  AND2X1 U16654 ( .IN1(test_so3), .IN2(WX751), .Q(n15839) );
  OR2X1 U16655 ( .IN1(n15841), .IN2(n15842), .Q(DATA_9_1) );
  AND2X1 U16656 ( .IN1(n11361), .IN2(n15843), .Q(n15842) );
  INVX0 U16657 ( .INP(n15844), .ZN(n15841) );
  OR2X1 U16658 ( .IN1(n15843), .IN2(n11361), .Q(n15844) );
  OR2X1 U16659 ( .IN1(n15845), .IN2(n15846), .Q(n11361) );
  INVX0 U16660 ( .INP(n15847), .ZN(n15846) );
  OR2X1 U16661 ( .IN1(n15848), .IN2(n15849), .Q(n15847) );
  AND2X1 U16662 ( .IN1(n15849), .IN2(n15848), .Q(n15845) );
  AND2X1 U16663 ( .IN1(n15850), .IN2(n15851), .Q(n15848) );
  OR2X1 U16664 ( .IN1(n2199), .IN2(n3469), .Q(n15851) );
  OR2X1 U16665 ( .IN1(WX705), .IN2(TM0), .Q(n15850) );
  OR2X1 U16666 ( .IN1(n15852), .IN2(n15853), .Q(n15849) );
  AND3X1 U16667 ( .IN1(n15854), .IN2(n15855), .IN3(n8971), .Q(n15853) );
  OR2X1 U16668 ( .IN1(n8969), .IN2(WX769), .Q(n15855) );
  OR2X1 U16669 ( .IN1(n8970), .IN2(WX897), .Q(n15854) );
  AND2X1 U16670 ( .IN1(n15856), .IN2(WX833), .Q(n15852) );
  OR2X1 U16671 ( .IN1(n15857), .IN2(n15858), .Q(n15856) );
  AND2X1 U16672 ( .IN1(n8969), .IN2(WX769), .Q(n15858) );
  AND2X1 U16673 ( .IN1(n8970), .IN2(WX897), .Q(n15857) );
  OR2X1 U16674 ( .IN1(n9054), .IN2(n2199), .Q(n15843) );
  OR2X1 U16675 ( .IN1(n15859), .IN2(n15860), .Q(DATA_9_0) );
  AND2X1 U16676 ( .IN1(n11355), .IN2(n15861), .Q(n15860) );
  INVX0 U16677 ( .INP(n15862), .ZN(n15859) );
  OR2X1 U16678 ( .IN1(n15861), .IN2(n11355), .Q(n15862) );
  OR2X1 U16679 ( .IN1(n15863), .IN2(n15864), .Q(n11355) );
  INVX0 U16680 ( .INP(n15865), .ZN(n15864) );
  OR2X1 U16681 ( .IN1(n15866), .IN2(n15867), .Q(n15865) );
  AND2X1 U16682 ( .IN1(n15867), .IN2(n15866), .Q(n15863) );
  AND2X1 U16683 ( .IN1(n15868), .IN2(n15869), .Q(n15866) );
  OR2X1 U16684 ( .IN1(n2199), .IN2(n3467), .Q(n15869) );
  OR2X1 U16685 ( .IN1(WX707), .IN2(TM0), .Q(n15868) );
  INVX0 U16686 ( .INP(n15870), .ZN(n15867) );
  AND2X1 U16687 ( .IN1(n15871), .IN2(n15872), .Q(n15870) );
  OR2X1 U16688 ( .IN1(n15873), .IN2(n9042), .Q(n15872) );
  INVX0 U16689 ( .INP(n15874), .ZN(n15871) );
  AND2X1 U16690 ( .IN1(n9042), .IN2(n15873), .Q(n15874) );
  AND2X1 U16691 ( .IN1(n15875), .IN2(n15876), .Q(n15873) );
  OR2X1 U16692 ( .IN1(WX835), .IN2(n9044), .Q(n15876) );
  OR2X1 U16693 ( .IN1(WX899), .IN2(n9043), .Q(n15875) );
  OR2X1 U16694 ( .IN1(n9053), .IN2(n2199), .Q(n15861) );
  AND2X1 U3558_U2 ( .IN1(n9224), .IN2(U3558_n1), .Q(n2245) );
  INVX0 U3558_U1 ( .INP(n9577), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(TM0), .ZN(U3871_n1) );
  AND2X1 U3871_U1 ( .IN1(n3278), .IN2(U3871_n1), .Q(n2153) );
  INVX0 U3991_U2 ( .INP(n2199), .ZN(U3991_n1) );
  AND2X1 U3991_U1 ( .IN1(n3278), .IN2(U3991_n1), .Q(n2152) );
  AND2X1 U5716_U2 ( .IN1(WX547), .IN2(U5716_n1), .Q(WX544) );
  INVX0 U5716_U1 ( .INP(n9632), .ZN(U5716_n1) );
  AND2X1 U5717_U2 ( .IN1(WX545), .IN2(U5717_n1), .Q(WX542) );
  INVX0 U5717_U1 ( .INP(n9632), .ZN(U5717_n1) );
  AND2X1 U5718_U2 ( .IN1(WX543), .IN2(U5718_n1), .Q(WX540) );
  INVX0 U5718_U1 ( .INP(n9632), .ZN(U5718_n1) );
  AND2X1 U5719_U2 ( .IN1(WX541), .IN2(U5719_n1), .Q(WX538) );
  INVX0 U5719_U1 ( .INP(n9632), .ZN(U5719_n1) );
  AND2X1 U5720_U2 ( .IN1(WX539), .IN2(U5720_n1), .Q(WX536) );
  INVX0 U5720_U1 ( .INP(n9632), .ZN(U5720_n1) );
  AND2X1 U5721_U2 ( .IN1(WX537), .IN2(U5721_n1), .Q(WX534) );
  INVX0 U5721_U1 ( .INP(n9632), .ZN(U5721_n1) );
  AND2X1 U5722_U2 ( .IN1(WX535), .IN2(U5722_n1), .Q(WX532) );
  INVX0 U5722_U1 ( .INP(n9632), .ZN(U5722_n1) );
  AND2X1 U5723_U2 ( .IN1(WX533), .IN2(U5723_n1), .Q(WX530) );
  INVX0 U5723_U1 ( .INP(n9632), .ZN(U5723_n1) );
  AND2X1 U5724_U2 ( .IN1(WX531), .IN2(U5724_n1), .Q(WX528) );
  INVX0 U5724_U1 ( .INP(n9631), .ZN(U5724_n1) );
  AND2X1 U5725_U2 ( .IN1(WX529), .IN2(U5725_n1), .Q(WX526) );
  INVX0 U5725_U1 ( .INP(n9631), .ZN(U5725_n1) );
  AND2X1 U5726_U2 ( .IN1(WX527), .IN2(U5726_n1), .Q(WX524) );
  INVX0 U5726_U1 ( .INP(n9631), .ZN(U5726_n1) );
  AND2X1 U5727_U2 ( .IN1(WX525), .IN2(U5727_n1), .Q(WX522) );
  INVX0 U5727_U1 ( .INP(n9631), .ZN(U5727_n1) );
  AND2X1 U5728_U2 ( .IN1(WX523), .IN2(U5728_n1), .Q(WX520) );
  INVX0 U5728_U1 ( .INP(n9631), .ZN(U5728_n1) );
  AND2X1 U5729_U2 ( .IN1(WX521), .IN2(U5729_n1), .Q(WX518) );
  INVX0 U5729_U1 ( .INP(n9631), .ZN(U5729_n1) );
  AND2X1 U5730_U2 ( .IN1(test_so1), .IN2(U5730_n1), .Q(WX516) );
  INVX0 U5730_U1 ( .INP(n9631), .ZN(U5730_n1) );
  AND2X1 U5731_U2 ( .IN1(WX517), .IN2(U5731_n1), .Q(WX514) );
  INVX0 U5731_U1 ( .INP(n9631), .ZN(U5731_n1) );
  AND2X1 U5732_U2 ( .IN1(WX515), .IN2(U5732_n1), .Q(WX512) );
  INVX0 U5732_U1 ( .INP(n9631), .ZN(U5732_n1) );
  AND2X1 U5733_U2 ( .IN1(WX513), .IN2(U5733_n1), .Q(WX510) );
  INVX0 U5733_U1 ( .INP(n9631), .ZN(U5733_n1) );
  AND2X1 U5734_U2 ( .IN1(WX511), .IN2(U5734_n1), .Q(WX508) );
  INVX0 U5734_U1 ( .INP(n9631), .ZN(U5734_n1) );
  AND2X1 U5735_U2 ( .IN1(WX509), .IN2(U5735_n1), .Q(WX506) );
  INVX0 U5735_U1 ( .INP(n9631), .ZN(U5735_n1) );
  AND2X1 U5736_U2 ( .IN1(WX507), .IN2(U5736_n1), .Q(WX504) );
  INVX0 U5736_U1 ( .INP(n9631), .ZN(U5736_n1) );
  AND2X1 U5737_U2 ( .IN1(WX505), .IN2(U5737_n1), .Q(WX502) );
  INVX0 U5737_U1 ( .INP(n9631), .ZN(U5737_n1) );
  AND2X1 U5738_U2 ( .IN1(WX503), .IN2(U5738_n1), .Q(WX500) );
  INVX0 U5738_U1 ( .INP(n9630), .ZN(U5738_n1) );
  AND2X1 U5739_U2 ( .IN1(WX501), .IN2(U5739_n1), .Q(WX498) );
  INVX0 U5739_U1 ( .INP(n9630), .ZN(U5739_n1) );
  AND2X1 U5740_U2 ( .IN1(WX499), .IN2(U5740_n1), .Q(WX496) );
  INVX0 U5740_U1 ( .INP(n9630), .ZN(U5740_n1) );
  AND2X1 U5741_U2 ( .IN1(WX497), .IN2(U5741_n1), .Q(WX494) );
  INVX0 U5741_U1 ( .INP(n9630), .ZN(U5741_n1) );
  AND2X1 U5742_U2 ( .IN1(WX495), .IN2(U5742_n1), .Q(WX492) );
  INVX0 U5742_U1 ( .INP(n9630), .ZN(U5742_n1) );
  AND2X1 U5743_U2 ( .IN1(WX493), .IN2(U5743_n1), .Q(WX490) );
  INVX0 U5743_U1 ( .INP(n9630), .ZN(U5743_n1) );
  AND2X1 U5744_U2 ( .IN1(WX491), .IN2(U5744_n1), .Q(WX488) );
  INVX0 U5744_U1 ( .INP(n9630), .ZN(U5744_n1) );
  AND2X1 U5745_U2 ( .IN1(WX489), .IN2(U5745_n1), .Q(WX486) );
  INVX0 U5745_U1 ( .INP(n9630), .ZN(U5745_n1) );
  AND2X1 U5746_U2 ( .IN1(WX487), .IN2(U5746_n1), .Q(WX484) );
  INVX0 U5746_U1 ( .INP(n9630), .ZN(U5746_n1) );
  AND2X1 U5747_U2 ( .IN1(WX5939), .IN2(U5747_n1), .Q(WX6002) );
  INVX0 U5747_U1 ( .INP(n9630), .ZN(U5747_n1) );
  AND2X1 U5748_U2 ( .IN1(test_so49), .IN2(U5748_n1), .Q(WX6000) );
  INVX0 U5748_U1 ( .INP(n9630), .ZN(U5748_n1) );
  AND2X1 U5749_U2 ( .IN1(WX5935), .IN2(U5749_n1), .Q(WX5998) );
  INVX0 U5749_U1 ( .INP(n9630), .ZN(U5749_n1) );
  AND2X1 U5750_U2 ( .IN1(WX5933), .IN2(U5750_n1), .Q(WX5996) );
  INVX0 U5750_U1 ( .INP(n9630), .ZN(U5750_n1) );
  AND2X1 U5751_U2 ( .IN1(WX5931), .IN2(U5751_n1), .Q(WX5994) );
  INVX0 U5751_U1 ( .INP(n9630), .ZN(U5751_n1) );
  AND2X1 U5752_U2 ( .IN1(WX3269), .IN2(U5752_n1), .Q(WX3332) );
  INVX0 U5752_U1 ( .INP(n9629), .ZN(U5752_n1) );
  AND2X1 U5753_U2 ( .IN1(WX3265), .IN2(U5753_n1), .Q(WX3328) );
  INVX0 U5753_U1 ( .INP(n9629), .ZN(U5753_n1) );
  AND2X1 U5754_U2 ( .IN1(WX3263), .IN2(U5754_n1), .Q(WX3326) );
  INVX0 U5754_U1 ( .INP(n9629), .ZN(U5754_n1) );
  AND2X1 U5755_U2 ( .IN1(WX11179), .IN2(U5755_n1), .Q(WX11242) );
  INVX0 U5755_U1 ( .INP(n9629), .ZN(U5755_n1) );
  AND2X1 U5756_U2 ( .IN1(WX11177), .IN2(U5756_n1), .Q(WX11240) );
  INVX0 U5756_U1 ( .INP(n9629), .ZN(U5756_n1) );
  AND2X1 U5757_U2 ( .IN1(WX11175), .IN2(U5757_n1), .Q(WX11238) );
  INVX0 U5757_U1 ( .INP(n9629), .ZN(U5757_n1) );
  AND2X1 U5758_U2 ( .IN1(WX11173), .IN2(U5758_n1), .Q(WX11236) );
  INVX0 U5758_U1 ( .INP(n9629), .ZN(U5758_n1) );
  AND2X1 U5759_U2 ( .IN1(test_so96), .IN2(U5759_n1), .Q(WX11234) );
  INVX0 U5759_U1 ( .INP(n9629), .ZN(U5759_n1) );
  AND2X1 U5760_U2 ( .IN1(WX11169), .IN2(U5760_n1), .Q(WX11232) );
  INVX0 U5760_U1 ( .INP(n9629), .ZN(U5760_n1) );
  AND2X1 U5761_U2 ( .IN1(WX11167), .IN2(U5761_n1), .Q(WX11230) );
  INVX0 U5761_U1 ( .INP(n9629), .ZN(U5761_n1) );
  AND2X1 U5762_U2 ( .IN1(WX11165), .IN2(U5762_n1), .Q(WX11228) );
  INVX0 U5762_U1 ( .INP(n9629), .ZN(U5762_n1) );
  AND2X1 U5763_U2 ( .IN1(WX11163), .IN2(U5763_n1), .Q(WX11226) );
  INVX0 U5763_U1 ( .INP(n9629), .ZN(U5763_n1) );
  AND2X1 U5764_U2 ( .IN1(WX11161), .IN2(U5764_n1), .Q(WX11224) );
  INVX0 U5764_U1 ( .INP(n9629), .ZN(U5764_n1) );
  AND2X1 U5765_U2 ( .IN1(WX11159), .IN2(U5765_n1), .Q(WX11222) );
  INVX0 U5765_U1 ( .INP(n9629), .ZN(U5765_n1) );
  AND2X1 U5766_U2 ( .IN1(WX11157), .IN2(U5766_n1), .Q(WX11220) );
  INVX0 U5766_U1 ( .INP(n9628), .ZN(U5766_n1) );
  AND2X1 U5767_U2 ( .IN1(WX11155), .IN2(U5767_n1), .Q(WX11218) );
  INVX0 U5767_U1 ( .INP(n9628), .ZN(U5767_n1) );
  AND2X1 U5768_U2 ( .IN1(WX11153), .IN2(U5768_n1), .Q(WX11216) );
  INVX0 U5768_U1 ( .INP(n9628), .ZN(U5768_n1) );
  AND2X1 U5769_U2 ( .IN1(WX11151), .IN2(U5769_n1), .Q(WX11214) );
  INVX0 U5769_U1 ( .INP(n9628), .ZN(U5769_n1) );
  AND2X1 U5770_U2 ( .IN1(WX11149), .IN2(U5770_n1), .Q(WX11212) );
  INVX0 U5770_U1 ( .INP(n9628), .ZN(U5770_n1) );
  AND2X1 U5771_U2 ( .IN1(WX11147), .IN2(U5771_n1), .Q(WX11210) );
  INVX0 U5771_U1 ( .INP(n9628), .ZN(U5771_n1) );
  AND2X1 U5772_U2 ( .IN1(WX11145), .IN2(U5772_n1), .Q(WX11208) );
  INVX0 U5772_U1 ( .INP(n9628), .ZN(U5772_n1) );
  AND2X1 U5773_U2 ( .IN1(WX11143), .IN2(U5773_n1), .Q(WX11206) );
  INVX0 U5773_U1 ( .INP(n9628), .ZN(U5773_n1) );
  AND2X1 U5774_U2 ( .IN1(WX11141), .IN2(U5774_n1), .Q(WX11204) );
  INVX0 U5774_U1 ( .INP(n9628), .ZN(U5774_n1) );
  AND2X1 U5775_U2 ( .IN1(WX11139), .IN2(U5775_n1), .Q(WX11202) );
  INVX0 U5775_U1 ( .INP(n9628), .ZN(U5775_n1) );
  AND2X1 U5776_U2 ( .IN1(test_so95), .IN2(U5776_n1), .Q(WX11200) );
  INVX0 U5776_U1 ( .INP(n9628), .ZN(U5776_n1) );
  AND2X1 U5777_U2 ( .IN1(WX11135), .IN2(U5777_n1), .Q(WX11198) );
  INVX0 U5777_U1 ( .INP(n9628), .ZN(U5777_n1) );
  AND2X1 U5778_U2 ( .IN1(WX11133), .IN2(U5778_n1), .Q(WX11196) );
  INVX0 U5778_U1 ( .INP(n9628), .ZN(U5778_n1) );
  AND2X1 U5779_U2 ( .IN1(WX11131), .IN2(U5779_n1), .Q(WX11194) );
  INVX0 U5779_U1 ( .INP(n9628), .ZN(U5779_n1) );
  AND2X1 U5780_U2 ( .IN1(WX11129), .IN2(U5780_n1), .Q(WX11192) );
  INVX0 U5780_U1 ( .INP(n9627), .ZN(U5780_n1) );
  AND2X1 U5781_U2 ( .IN1(WX11127), .IN2(U5781_n1), .Q(WX11190) );
  INVX0 U5781_U1 ( .INP(n9627), .ZN(U5781_n1) );
  AND2X1 U5782_U2 ( .IN1(WX11125), .IN2(U5782_n1), .Q(WX11188) );
  INVX0 U5782_U1 ( .INP(n9627), .ZN(U5782_n1) );
  AND2X1 U5783_U2 ( .IN1(WX11123), .IN2(U5783_n1), .Q(WX11186) );
  INVX0 U5783_U1 ( .INP(n9627), .ZN(U5783_n1) );
  AND2X1 U5784_U2 ( .IN1(WX11121), .IN2(U5784_n1), .Q(WX11184) );
  INVX0 U5784_U1 ( .INP(n9627), .ZN(U5784_n1) );
  AND2X1 U5785_U2 ( .IN1(WX11119), .IN2(U5785_n1), .Q(WX11182) );
  INVX0 U5785_U1 ( .INP(n9627), .ZN(U5785_n1) );
  AND2X1 U5786_U2 ( .IN1(WX11117), .IN2(U5786_n1), .Q(WX11180) );
  INVX0 U5786_U1 ( .INP(n9627), .ZN(U5786_n1) );
  AND2X1 U5787_U2 ( .IN1(WX11115), .IN2(U5787_n1), .Q(WX11178) );
  INVX0 U5787_U1 ( .INP(n9627), .ZN(U5787_n1) );
  AND2X1 U5788_U2 ( .IN1(WX11113), .IN2(U5788_n1), .Q(WX11176) );
  INVX0 U5788_U1 ( .INP(n9627), .ZN(U5788_n1) );
  AND2X1 U5789_U2 ( .IN1(WX11111), .IN2(U5789_n1), .Q(WX11174) );
  INVX0 U5789_U1 ( .INP(n9627), .ZN(U5789_n1) );
  AND2X1 U5790_U2 ( .IN1(WX11109), .IN2(U5790_n1), .Q(WX11172) );
  INVX0 U5790_U1 ( .INP(n9627), .ZN(U5790_n1) );
  AND2X1 U5791_U2 ( .IN1(WX11107), .IN2(U5791_n1), .Q(WX11170) );
  INVX0 U5791_U1 ( .INP(n9627), .ZN(U5791_n1) );
  AND2X1 U5792_U2 ( .IN1(WX11105), .IN2(U5792_n1), .Q(WX11168) );
  INVX0 U5792_U1 ( .INP(n9627), .ZN(U5792_n1) );
  AND2X1 U5793_U2 ( .IN1(test_so94), .IN2(U5793_n1), .Q(WX11166) );
  INVX0 U5793_U1 ( .INP(n9627), .ZN(U5793_n1) );
  AND2X1 U5794_U2 ( .IN1(WX11101), .IN2(U5794_n1), .Q(WX11164) );
  INVX0 U5794_U1 ( .INP(n9626), .ZN(U5794_n1) );
  AND2X1 U5795_U2 ( .IN1(WX11099), .IN2(U5795_n1), .Q(WX11162) );
  INVX0 U5795_U1 ( .INP(n9626), .ZN(U5795_n1) );
  AND2X1 U5796_U2 ( .IN1(WX11097), .IN2(U5796_n1), .Q(WX11160) );
  INVX0 U5796_U1 ( .INP(n9626), .ZN(U5796_n1) );
  AND2X1 U5797_U2 ( .IN1(WX11095), .IN2(U5797_n1), .Q(WX11158) );
  INVX0 U5797_U1 ( .INP(n9626), .ZN(U5797_n1) );
  AND2X1 U5798_U2 ( .IN1(WX11093), .IN2(U5798_n1), .Q(WX11156) );
  INVX0 U5798_U1 ( .INP(n9626), .ZN(U5798_n1) );
  AND2X1 U5799_U2 ( .IN1(WX11091), .IN2(U5799_n1), .Q(WX11154) );
  INVX0 U5799_U1 ( .INP(n9626), .ZN(U5799_n1) );
  AND2X1 U5800_U2 ( .IN1(WX11089), .IN2(U5800_n1), .Q(WX11152) );
  INVX0 U5800_U1 ( .INP(n9626), .ZN(U5800_n1) );
  AND2X1 U5801_U2 ( .IN1(WX11087), .IN2(U5801_n1), .Q(WX11150) );
  INVX0 U5801_U1 ( .INP(n9626), .ZN(U5801_n1) );
  AND2X1 U5802_U2 ( .IN1(WX11085), .IN2(U5802_n1), .Q(WX11148) );
  INVX0 U5802_U1 ( .INP(n9626), .ZN(U5802_n1) );
  AND2X1 U5803_U2 ( .IN1(WX11083), .IN2(U5803_n1), .Q(WX11146) );
  INVX0 U5803_U1 ( .INP(n9626), .ZN(U5803_n1) );
  AND2X1 U5804_U2 ( .IN1(WX11081), .IN2(U5804_n1), .Q(WX11144) );
  INVX0 U5804_U1 ( .INP(n9626), .ZN(U5804_n1) );
  AND2X1 U5805_U2 ( .IN1(WX11079), .IN2(U5805_n1), .Q(WX11142) );
  INVX0 U5805_U1 ( .INP(n9626), .ZN(U5805_n1) );
  AND2X1 U5806_U2 ( .IN1(WX11077), .IN2(U5806_n1), .Q(WX11140) );
  INVX0 U5806_U1 ( .INP(n9626), .ZN(U5806_n1) );
  AND2X1 U5807_U2 ( .IN1(WX11075), .IN2(U5807_n1), .Q(WX11138) );
  INVX0 U5807_U1 ( .INP(n9626), .ZN(U5807_n1) );
  AND2X1 U5808_U2 ( .IN1(WX11073), .IN2(U5808_n1), .Q(WX11136) );
  INVX0 U5808_U1 ( .INP(n9625), .ZN(U5808_n1) );
  AND2X1 U5809_U2 ( .IN1(WX11071), .IN2(U5809_n1), .Q(WX11134) );
  INVX0 U5809_U1 ( .INP(n9625), .ZN(U5809_n1) );
  AND2X1 U5810_U2 ( .IN1(test_so93), .IN2(U5810_n1), .Q(WX11132) );
  INVX0 U5810_U1 ( .INP(n9625), .ZN(U5810_n1) );
  AND2X1 U5811_U2 ( .IN1(WX11067), .IN2(U5811_n1), .Q(WX11130) );
  INVX0 U5811_U1 ( .INP(n9625), .ZN(U5811_n1) );
  AND2X1 U5812_U2 ( .IN1(WX11065), .IN2(U5812_n1), .Q(WX11128) );
  INVX0 U5812_U1 ( .INP(n9625), .ZN(U5812_n1) );
  AND2X1 U5813_U2 ( .IN1(WX11063), .IN2(U5813_n1), .Q(WX11126) );
  INVX0 U5813_U1 ( .INP(n9625), .ZN(U5813_n1) );
  AND2X1 U5814_U2 ( .IN1(WX11061), .IN2(U5814_n1), .Q(WX11124) );
  INVX0 U5814_U1 ( .INP(n9625), .ZN(U5814_n1) );
  AND2X1 U5815_U2 ( .IN1(WX11059), .IN2(U5815_n1), .Q(WX11122) );
  INVX0 U5815_U1 ( .INP(n9625), .ZN(U5815_n1) );
  AND2X1 U5816_U2 ( .IN1(WX11057), .IN2(U5816_n1), .Q(WX11120) );
  INVX0 U5816_U1 ( .INP(n9625), .ZN(U5816_n1) );
  AND2X1 U5817_U2 ( .IN1(WX11055), .IN2(U5817_n1), .Q(WX11118) );
  INVX0 U5817_U1 ( .INP(n9625), .ZN(U5817_n1) );
  AND2X1 U5818_U2 ( .IN1(WX11053), .IN2(U5818_n1), .Q(WX11116) );
  INVX0 U5818_U1 ( .INP(n9625), .ZN(U5818_n1) );
  AND2X1 U5819_U2 ( .IN1(WX11051), .IN2(U5819_n1), .Q(WX11114) );
  INVX0 U5819_U1 ( .INP(n9625), .ZN(U5819_n1) );
  AND2X1 U5820_U2 ( .IN1(WX11049), .IN2(U5820_n1), .Q(WX11112) );
  INVX0 U5820_U1 ( .INP(n9625), .ZN(U5820_n1) );
  AND2X1 U5821_U2 ( .IN1(WX11047), .IN2(U5821_n1), .Q(WX11110) );
  INVX0 U5821_U1 ( .INP(n9625), .ZN(U5821_n1) );
  AND2X1 U5822_U2 ( .IN1(WX11045), .IN2(U5822_n1), .Q(WX11108) );
  INVX0 U5822_U1 ( .INP(n9624), .ZN(U5822_n1) );
  AND2X1 U5823_U2 ( .IN1(WX11043), .IN2(U5823_n1), .Q(WX11106) );
  INVX0 U5823_U1 ( .INP(n9624), .ZN(U5823_n1) );
  AND2X1 U5824_U2 ( .IN1(WX11041), .IN2(U5824_n1), .Q(WX11104) );
  INVX0 U5824_U1 ( .INP(n9624), .ZN(U5824_n1) );
  AND2X1 U5825_U2 ( .IN1(WX11039), .IN2(U5825_n1), .Q(WX11102) );
  INVX0 U5825_U1 ( .INP(n9624), .ZN(U5825_n1) );
  AND2X1 U5826_U2 ( .IN1(WX11037), .IN2(U5826_n1), .Q(WX11100) );
  INVX0 U5826_U1 ( .INP(n9624), .ZN(U5826_n1) );
  AND2X1 U5827_U2 ( .IN1(test_so92), .IN2(U5827_n1), .Q(WX11098) );
  INVX0 U5827_U1 ( .INP(n9624), .ZN(U5827_n1) );
  AND2X1 U5828_U2 ( .IN1(WX11033), .IN2(U5828_n1), .Q(WX11096) );
  INVX0 U5828_U1 ( .INP(n9624), .ZN(U5828_n1) );
  AND2X1 U5829_U2 ( .IN1(WX11031), .IN2(U5829_n1), .Q(WX11094) );
  INVX0 U5829_U1 ( .INP(n9624), .ZN(U5829_n1) );
  AND2X1 U5830_U2 ( .IN1(WX11029), .IN2(U5830_n1), .Q(WX11092) );
  INVX0 U5830_U1 ( .INP(n9624), .ZN(U5830_n1) );
  AND2X1 U5831_U2 ( .IN1(WX11027), .IN2(U5831_n1), .Q(WX11090) );
  INVX0 U5831_U1 ( .INP(n9624), .ZN(U5831_n1) );
  AND2X1 U5832_U2 ( .IN1(WX11025), .IN2(U5832_n1), .Q(WX11088) );
  INVX0 U5832_U1 ( .INP(n9624), .ZN(U5832_n1) );
  AND2X1 U5833_U2 ( .IN1(WX11023), .IN2(U5833_n1), .Q(WX11086) );
  INVX0 U5833_U1 ( .INP(n9624), .ZN(U5833_n1) );
  AND2X1 U5834_U2 ( .IN1(WX11021), .IN2(U5834_n1), .Q(WX11084) );
  INVX0 U5834_U1 ( .INP(n9624), .ZN(U5834_n1) );
  AND2X1 U5835_U2 ( .IN1(WX9886), .IN2(U5835_n1), .Q(WX9949) );
  INVX0 U5835_U1 ( .INP(n9624), .ZN(U5835_n1) );
  AND2X1 U5836_U2 ( .IN1(WX9884), .IN2(U5836_n1), .Q(WX9947) );
  INVX0 U5836_U1 ( .INP(n9623), .ZN(U5836_n1) );
  AND2X1 U5837_U2 ( .IN1(WX9882), .IN2(U5837_n1), .Q(WX9945) );
  INVX0 U5837_U1 ( .INP(n9623), .ZN(U5837_n1) );
  AND2X1 U5838_U2 ( .IN1(WX9880), .IN2(U5838_n1), .Q(WX9943) );
  INVX0 U5838_U1 ( .INP(n9623), .ZN(U5838_n1) );
  AND2X1 U5839_U2 ( .IN1(WX9878), .IN2(U5839_n1), .Q(WX9941) );
  INVX0 U5839_U1 ( .INP(n9623), .ZN(U5839_n1) );
  AND2X1 U5840_U2 ( .IN1(WX9876), .IN2(U5840_n1), .Q(WX9939) );
  INVX0 U5840_U1 ( .INP(n9623), .ZN(U5840_n1) );
  AND2X1 U5841_U2 ( .IN1(WX9874), .IN2(U5841_n1), .Q(WX9937) );
  INVX0 U5841_U1 ( .INP(n9623), .ZN(U5841_n1) );
  AND2X1 U5842_U2 ( .IN1(WX9872), .IN2(U5842_n1), .Q(WX9935) );
  INVX0 U5842_U1 ( .INP(n9623), .ZN(U5842_n1) );
  AND2X1 U5843_U2 ( .IN1(WX9870), .IN2(U5843_n1), .Q(WX9933) );
  INVX0 U5843_U1 ( .INP(n9623), .ZN(U5843_n1) );
  AND2X1 U5844_U2 ( .IN1(WX9868), .IN2(U5844_n1), .Q(WX9931) );
  INVX0 U5844_U1 ( .INP(n9623), .ZN(U5844_n1) );
  AND2X1 U5845_U2 ( .IN1(WX9866), .IN2(U5845_n1), .Q(WX9929) );
  INVX0 U5845_U1 ( .INP(n9623), .ZN(U5845_n1) );
  AND2X1 U5846_U2 ( .IN1(WX9864), .IN2(U5846_n1), .Q(WX9927) );
  INVX0 U5846_U1 ( .INP(n9623), .ZN(U5846_n1) );
  AND2X1 U5847_U2 ( .IN1(WX9862), .IN2(U5847_n1), .Q(WX9925) );
  INVX0 U5847_U1 ( .INP(n9623), .ZN(U5847_n1) );
  AND2X1 U5848_U2 ( .IN1(WX9860), .IN2(U5848_n1), .Q(WX9923) );
  INVX0 U5848_U1 ( .INP(n9623), .ZN(U5848_n1) );
  AND2X1 U5849_U2 ( .IN1(WX9858), .IN2(U5849_n1), .Q(WX9921) );
  INVX0 U5849_U1 ( .INP(n9623), .ZN(U5849_n1) );
  AND2X1 U5850_U2 ( .IN1(WX9856), .IN2(U5850_n1), .Q(WX9919) );
  INVX0 U5850_U1 ( .INP(n9622), .ZN(U5850_n1) );
  AND2X1 U5851_U2 ( .IN1(test_so84), .IN2(U5851_n1), .Q(WX9917) );
  INVX0 U5851_U1 ( .INP(n9622), .ZN(U5851_n1) );
  AND2X1 U5852_U2 ( .IN1(WX9852), .IN2(U5852_n1), .Q(WX9915) );
  INVX0 U5852_U1 ( .INP(n9622), .ZN(U5852_n1) );
  AND2X1 U5853_U2 ( .IN1(WX9850), .IN2(U5853_n1), .Q(WX9913) );
  INVX0 U5853_U1 ( .INP(n9622), .ZN(U5853_n1) );
  AND2X1 U5854_U2 ( .IN1(WX9848), .IN2(U5854_n1), .Q(WX9911) );
  INVX0 U5854_U1 ( .INP(n9622), .ZN(U5854_n1) );
  AND2X1 U5855_U2 ( .IN1(WX9846), .IN2(U5855_n1), .Q(WX9909) );
  INVX0 U5855_U1 ( .INP(n9622), .ZN(U5855_n1) );
  AND2X1 U5856_U2 ( .IN1(WX9844), .IN2(U5856_n1), .Q(WX9907) );
  INVX0 U5856_U1 ( .INP(n9622), .ZN(U5856_n1) );
  AND2X1 U5857_U2 ( .IN1(WX9842), .IN2(U5857_n1), .Q(WX9905) );
  INVX0 U5857_U1 ( .INP(n9622), .ZN(U5857_n1) );
  AND2X1 U5858_U2 ( .IN1(WX9840), .IN2(U5858_n1), .Q(WX9903) );
  INVX0 U5858_U1 ( .INP(n9622), .ZN(U5858_n1) );
  AND2X1 U5859_U2 ( .IN1(WX9838), .IN2(U5859_n1), .Q(WX9901) );
  INVX0 U5859_U1 ( .INP(n9622), .ZN(U5859_n1) );
  AND2X1 U5860_U2 ( .IN1(WX9836), .IN2(U5860_n1), .Q(WX9899) );
  INVX0 U5860_U1 ( .INP(n9622), .ZN(U5860_n1) );
  AND2X1 U5861_U2 ( .IN1(WX9834), .IN2(U5861_n1), .Q(WX9897) );
  INVX0 U5861_U1 ( .INP(n9622), .ZN(U5861_n1) );
  AND2X1 U5862_U2 ( .IN1(WX9832), .IN2(U5862_n1), .Q(WX9895) );
  INVX0 U5862_U1 ( .INP(n9622), .ZN(U5862_n1) );
  AND2X1 U5863_U2 ( .IN1(WX9830), .IN2(U5863_n1), .Q(WX9893) );
  INVX0 U5863_U1 ( .INP(n9622), .ZN(U5863_n1) );
  AND2X1 U5864_U2 ( .IN1(WX9828), .IN2(U5864_n1), .Q(WX9891) );
  INVX0 U5864_U1 ( .INP(n9621), .ZN(U5864_n1) );
  AND2X1 U5865_U2 ( .IN1(WX9826), .IN2(U5865_n1), .Q(WX9889) );
  INVX0 U5865_U1 ( .INP(n9621), .ZN(U5865_n1) );
  AND2X1 U5866_U2 ( .IN1(WX9824), .IN2(U5866_n1), .Q(WX9887) );
  INVX0 U5866_U1 ( .INP(n9621), .ZN(U5866_n1) );
  AND2X1 U5867_U2 ( .IN1(WX9822), .IN2(U5867_n1), .Q(WX9885) );
  INVX0 U5867_U1 ( .INP(n9621), .ZN(U5867_n1) );
  AND2X1 U5868_U2 ( .IN1(test_so83), .IN2(U5868_n1), .Q(WX9883) );
  INVX0 U5868_U1 ( .INP(n9621), .ZN(U5868_n1) );
  AND2X1 U5869_U2 ( .IN1(WX9818), .IN2(U5869_n1), .Q(WX9881) );
  INVX0 U5869_U1 ( .INP(n9621), .ZN(U5869_n1) );
  AND2X1 U5870_U2 ( .IN1(WX9816), .IN2(U5870_n1), .Q(WX9879) );
  INVX0 U5870_U1 ( .INP(n9621), .ZN(U5870_n1) );
  AND2X1 U5871_U2 ( .IN1(WX9814), .IN2(U5871_n1), .Q(WX9877) );
  INVX0 U5871_U1 ( .INP(n9621), .ZN(U5871_n1) );
  AND2X1 U5872_U2 ( .IN1(WX9812), .IN2(U5872_n1), .Q(WX9875) );
  INVX0 U5872_U1 ( .INP(n9621), .ZN(U5872_n1) );
  AND2X1 U5873_U2 ( .IN1(WX9810), .IN2(U5873_n1), .Q(WX9873) );
  INVX0 U5873_U1 ( .INP(n9621), .ZN(U5873_n1) );
  AND2X1 U5874_U2 ( .IN1(WX9808), .IN2(U5874_n1), .Q(WX9871) );
  INVX0 U5874_U1 ( .INP(n9621), .ZN(U5874_n1) );
  AND2X1 U5875_U2 ( .IN1(WX9806), .IN2(U5875_n1), .Q(WX9869) );
  INVX0 U5875_U1 ( .INP(n9621), .ZN(U5875_n1) );
  AND2X1 U5876_U2 ( .IN1(WX9804), .IN2(U5876_n1), .Q(WX9867) );
  INVX0 U5876_U1 ( .INP(n9621), .ZN(U5876_n1) );
  AND2X1 U5877_U2 ( .IN1(WX9802), .IN2(U5877_n1), .Q(WX9865) );
  INVX0 U5877_U1 ( .INP(n9621), .ZN(U5877_n1) );
  AND2X1 U5878_U2 ( .IN1(WX9800), .IN2(U5878_n1), .Q(WX9863) );
  INVX0 U5878_U1 ( .INP(n9620), .ZN(U5878_n1) );
  AND2X1 U5879_U2 ( .IN1(WX9798), .IN2(U5879_n1), .Q(WX9861) );
  INVX0 U5879_U1 ( .INP(n9620), .ZN(U5879_n1) );
  AND2X1 U5880_U2 ( .IN1(WX9796), .IN2(U5880_n1), .Q(WX9859) );
  INVX0 U5880_U1 ( .INP(n9620), .ZN(U5880_n1) );
  AND2X1 U5881_U2 ( .IN1(WX9794), .IN2(U5881_n1), .Q(WX9857) );
  INVX0 U5881_U1 ( .INP(n9620), .ZN(U5881_n1) );
  AND2X1 U5882_U2 ( .IN1(WX9792), .IN2(U5882_n1), .Q(WX9855) );
  INVX0 U5882_U1 ( .INP(n9620), .ZN(U5882_n1) );
  AND2X1 U5883_U2 ( .IN1(WX9790), .IN2(U5883_n1), .Q(WX9853) );
  INVX0 U5883_U1 ( .INP(n9620), .ZN(U5883_n1) );
  AND2X1 U5884_U2 ( .IN1(WX9788), .IN2(U5884_n1), .Q(WX9851) );
  INVX0 U5884_U1 ( .INP(n9620), .ZN(U5884_n1) );
  AND2X1 U5885_U2 ( .IN1(test_so82), .IN2(U5885_n1), .Q(WX9849) );
  INVX0 U5885_U1 ( .INP(n9620), .ZN(U5885_n1) );
  AND2X1 U5886_U2 ( .IN1(WX9784), .IN2(U5886_n1), .Q(WX9847) );
  INVX0 U5886_U1 ( .INP(n9620), .ZN(U5886_n1) );
  AND2X1 U5887_U2 ( .IN1(WX9782), .IN2(U5887_n1), .Q(WX9845) );
  INVX0 U5887_U1 ( .INP(n9620), .ZN(U5887_n1) );
  AND2X1 U5888_U2 ( .IN1(WX9780), .IN2(U5888_n1), .Q(WX9843) );
  INVX0 U5888_U1 ( .INP(n9620), .ZN(U5888_n1) );
  AND2X1 U5889_U2 ( .IN1(WX9778), .IN2(U5889_n1), .Q(WX9841) );
  INVX0 U5889_U1 ( .INP(n9620), .ZN(U5889_n1) );
  AND2X1 U5890_U2 ( .IN1(WX9776), .IN2(U5890_n1), .Q(WX9839) );
  INVX0 U5890_U1 ( .INP(n9620), .ZN(U5890_n1) );
  AND2X1 U5891_U2 ( .IN1(WX9774), .IN2(U5891_n1), .Q(WX9837) );
  INVX0 U5891_U1 ( .INP(n9620), .ZN(U5891_n1) );
  AND2X1 U5892_U2 ( .IN1(WX9772), .IN2(U5892_n1), .Q(WX9835) );
  INVX0 U5892_U1 ( .INP(n9619), .ZN(U5892_n1) );
  AND2X1 U5893_U2 ( .IN1(WX9770), .IN2(U5893_n1), .Q(WX9833) );
  INVX0 U5893_U1 ( .INP(n9619), .ZN(U5893_n1) );
  AND2X1 U5894_U2 ( .IN1(WX9768), .IN2(U5894_n1), .Q(WX9831) );
  INVX0 U5894_U1 ( .INP(n9619), .ZN(U5894_n1) );
  AND2X1 U5895_U2 ( .IN1(WX9766), .IN2(U5895_n1), .Q(WX9829) );
  INVX0 U5895_U1 ( .INP(n9619), .ZN(U5895_n1) );
  AND2X1 U5896_U2 ( .IN1(WX9764), .IN2(U5896_n1), .Q(WX9827) );
  INVX0 U5896_U1 ( .INP(n9619), .ZN(U5896_n1) );
  AND2X1 U5897_U2 ( .IN1(WX9762), .IN2(U5897_n1), .Q(WX9825) );
  INVX0 U5897_U1 ( .INP(n9619), .ZN(U5897_n1) );
  AND2X1 U5898_U2 ( .IN1(WX9760), .IN2(U5898_n1), .Q(WX9823) );
  INVX0 U5898_U1 ( .INP(n9619), .ZN(U5898_n1) );
  AND2X1 U5899_U2 ( .IN1(WX9758), .IN2(U5899_n1), .Q(WX9821) );
  INVX0 U5899_U1 ( .INP(n9619), .ZN(U5899_n1) );
  AND2X1 U5900_U2 ( .IN1(WX9756), .IN2(U5900_n1), .Q(WX9819) );
  INVX0 U5900_U1 ( .INP(n9619), .ZN(U5900_n1) );
  AND2X1 U5901_U2 ( .IN1(WX9754), .IN2(U5901_n1), .Q(WX9817) );
  INVX0 U5901_U1 ( .INP(n9619), .ZN(U5901_n1) );
  AND2X1 U5902_U2 ( .IN1(test_so81), .IN2(U5902_n1), .Q(WX9815) );
  INVX0 U5902_U1 ( .INP(n9619), .ZN(U5902_n1) );
  AND2X1 U5903_U2 ( .IN1(WX9750), .IN2(U5903_n1), .Q(WX9813) );
  INVX0 U5903_U1 ( .INP(n9619), .ZN(U5903_n1) );
  AND2X1 U5904_U2 ( .IN1(WX9748), .IN2(U5904_n1), .Q(WX9811) );
  INVX0 U5904_U1 ( .INP(n9619), .ZN(U5904_n1) );
  AND2X1 U5905_U2 ( .IN1(WX9746), .IN2(U5905_n1), .Q(WX9809) );
  INVX0 U5905_U1 ( .INP(n9619), .ZN(U5905_n1) );
  AND2X1 U5906_U2 ( .IN1(WX9744), .IN2(U5906_n1), .Q(WX9807) );
  INVX0 U5906_U1 ( .INP(n9618), .ZN(U5906_n1) );
  AND2X1 U5907_U2 ( .IN1(WX9742), .IN2(U5907_n1), .Q(WX9805) );
  INVX0 U5907_U1 ( .INP(n9618), .ZN(U5907_n1) );
  AND2X1 U5908_U2 ( .IN1(WX9740), .IN2(U5908_n1), .Q(WX9803) );
  INVX0 U5908_U1 ( .INP(n9618), .ZN(U5908_n1) );
  AND2X1 U5909_U2 ( .IN1(WX9738), .IN2(U5909_n1), .Q(WX9801) );
  INVX0 U5909_U1 ( .INP(n9618), .ZN(U5909_n1) );
  AND2X1 U5910_U2 ( .IN1(WX9736), .IN2(U5910_n1), .Q(WX9799) );
  INVX0 U5910_U1 ( .INP(n9618), .ZN(U5910_n1) );
  AND2X1 U5911_U2 ( .IN1(WX9734), .IN2(U5911_n1), .Q(WX9797) );
  INVX0 U5911_U1 ( .INP(n9618), .ZN(U5911_n1) );
  AND2X1 U5912_U2 ( .IN1(WX9732), .IN2(U5912_n1), .Q(WX9795) );
  INVX0 U5912_U1 ( .INP(n9618), .ZN(U5912_n1) );
  AND2X1 U5913_U2 ( .IN1(WX9730), .IN2(U5913_n1), .Q(WX9793) );
  INVX0 U5913_U1 ( .INP(n9618), .ZN(U5913_n1) );
  AND2X1 U5914_U2 ( .IN1(WX9728), .IN2(U5914_n1), .Q(WX9791) );
  INVX0 U5914_U1 ( .INP(n9618), .ZN(U5914_n1) );
  AND2X1 U5915_U2 ( .IN1(WX8593), .IN2(U5915_n1), .Q(WX8656) );
  INVX0 U5915_U1 ( .INP(n9618), .ZN(U5915_n1) );
  AND2X1 U5916_U2 ( .IN1(WX8591), .IN2(U5916_n1), .Q(WX8654) );
  INVX0 U5916_U1 ( .INP(n9618), .ZN(U5916_n1) );
  AND2X1 U5917_U2 ( .IN1(WX8589), .IN2(U5917_n1), .Q(WX8652) );
  INVX0 U5917_U1 ( .INP(n9618), .ZN(U5917_n1) );
  AND2X1 U5918_U2 ( .IN1(WX8587), .IN2(U5918_n1), .Q(WX8650) );
  INVX0 U5918_U1 ( .INP(n9618), .ZN(U5918_n1) );
  AND2X1 U5919_U2 ( .IN1(WX8585), .IN2(U5919_n1), .Q(WX8648) );
  INVX0 U5919_U1 ( .INP(n9618), .ZN(U5919_n1) );
  AND2X1 U5920_U2 ( .IN1(WX8583), .IN2(U5920_n1), .Q(WX8646) );
  INVX0 U5920_U1 ( .INP(n9617), .ZN(U5920_n1) );
  AND2X1 U5921_U2 ( .IN1(WX8581), .IN2(U5921_n1), .Q(WX8644) );
  INVX0 U5921_U1 ( .INP(n9617), .ZN(U5921_n1) );
  AND2X1 U5922_U2 ( .IN1(WX8579), .IN2(U5922_n1), .Q(WX8642) );
  INVX0 U5922_U1 ( .INP(n9617), .ZN(U5922_n1) );
  AND2X1 U5923_U2 ( .IN1(WX8577), .IN2(U5923_n1), .Q(WX8640) );
  INVX0 U5923_U1 ( .INP(n9617), .ZN(U5923_n1) );
  AND2X1 U5924_U2 ( .IN1(WX8575), .IN2(U5924_n1), .Q(WX8638) );
  INVX0 U5924_U1 ( .INP(n9617), .ZN(U5924_n1) );
  AND2X1 U5925_U2 ( .IN1(WX8573), .IN2(U5925_n1), .Q(WX8636) );
  INVX0 U5925_U1 ( .INP(n9617), .ZN(U5925_n1) );
  AND2X1 U5926_U2 ( .IN1(test_so73), .IN2(U5926_n1), .Q(WX8634) );
  INVX0 U5926_U1 ( .INP(n9617), .ZN(U5926_n1) );
  AND2X1 U5927_U2 ( .IN1(WX8569), .IN2(U5927_n1), .Q(WX8632) );
  INVX0 U5927_U1 ( .INP(n9617), .ZN(U5927_n1) );
  AND2X1 U5928_U2 ( .IN1(WX8567), .IN2(U5928_n1), .Q(WX8630) );
  INVX0 U5928_U1 ( .INP(n9617), .ZN(U5928_n1) );
  AND2X1 U5929_U2 ( .IN1(WX8565), .IN2(U5929_n1), .Q(WX8628) );
  INVX0 U5929_U1 ( .INP(n9617), .ZN(U5929_n1) );
  AND2X1 U5930_U2 ( .IN1(WX8563), .IN2(U5930_n1), .Q(WX8626) );
  INVX0 U5930_U1 ( .INP(n9617), .ZN(U5930_n1) );
  AND2X1 U5931_U2 ( .IN1(WX8561), .IN2(U5931_n1), .Q(WX8624) );
  INVX0 U5931_U1 ( .INP(n9617), .ZN(U5931_n1) );
  AND2X1 U5932_U2 ( .IN1(WX8559), .IN2(U5932_n1), .Q(WX8622) );
  INVX0 U5932_U1 ( .INP(n9617), .ZN(U5932_n1) );
  AND2X1 U5933_U2 ( .IN1(WX8557), .IN2(U5933_n1), .Q(WX8620) );
  INVX0 U5933_U1 ( .INP(n9617), .ZN(U5933_n1) );
  AND2X1 U5934_U2 ( .IN1(WX8555), .IN2(U5934_n1), .Q(WX8618) );
  INVX0 U5934_U1 ( .INP(n9616), .ZN(U5934_n1) );
  AND2X1 U5935_U2 ( .IN1(WX8553), .IN2(U5935_n1), .Q(WX8616) );
  INVX0 U5935_U1 ( .INP(n9616), .ZN(U5935_n1) );
  AND2X1 U5936_U2 ( .IN1(WX8551), .IN2(U5936_n1), .Q(WX8614) );
  INVX0 U5936_U1 ( .INP(n9616), .ZN(U5936_n1) );
  AND2X1 U5937_U2 ( .IN1(WX8549), .IN2(U5937_n1), .Q(WX8612) );
  INVX0 U5937_U1 ( .INP(n9616), .ZN(U5937_n1) );
  AND2X1 U5938_U2 ( .IN1(WX8547), .IN2(U5938_n1), .Q(WX8610) );
  INVX0 U5938_U1 ( .INP(n9616), .ZN(U5938_n1) );
  AND2X1 U5939_U2 ( .IN1(WX8545), .IN2(U5939_n1), .Q(WX8608) );
  INVX0 U5939_U1 ( .INP(n9616), .ZN(U5939_n1) );
  AND2X1 U5940_U2 ( .IN1(WX8543), .IN2(U5940_n1), .Q(WX8606) );
  INVX0 U5940_U1 ( .INP(n9616), .ZN(U5940_n1) );
  AND2X1 U5941_U2 ( .IN1(WX8541), .IN2(U5941_n1), .Q(WX8604) );
  INVX0 U5941_U1 ( .INP(n9616), .ZN(U5941_n1) );
  AND2X1 U5942_U2 ( .IN1(WX8539), .IN2(U5942_n1), .Q(WX8602) );
  INVX0 U5942_U1 ( .INP(n9616), .ZN(U5942_n1) );
  AND2X1 U5943_U2 ( .IN1(test_so72), .IN2(U5943_n1), .Q(WX8600) );
  INVX0 U5943_U1 ( .INP(n9616), .ZN(U5943_n1) );
  AND2X1 U5944_U2 ( .IN1(WX8535), .IN2(U5944_n1), .Q(WX8598) );
  INVX0 U5944_U1 ( .INP(n9616), .ZN(U5944_n1) );
  AND2X1 U5945_U2 ( .IN1(WX8533), .IN2(U5945_n1), .Q(WX8596) );
  INVX0 U5945_U1 ( .INP(n9616), .ZN(U5945_n1) );
  AND2X1 U5946_U2 ( .IN1(WX8531), .IN2(U5946_n1), .Q(WX8594) );
  INVX0 U5946_U1 ( .INP(n9616), .ZN(U5946_n1) );
  AND2X1 U5947_U2 ( .IN1(WX8529), .IN2(U5947_n1), .Q(WX8592) );
  INVX0 U5947_U1 ( .INP(n9616), .ZN(U5947_n1) );
  AND2X1 U5948_U2 ( .IN1(WX8527), .IN2(U5948_n1), .Q(WX8590) );
  INVX0 U5948_U1 ( .INP(n9615), .ZN(U5948_n1) );
  AND2X1 U5949_U2 ( .IN1(WX8525), .IN2(U5949_n1), .Q(WX8588) );
  INVX0 U5949_U1 ( .INP(n9615), .ZN(U5949_n1) );
  AND2X1 U5950_U2 ( .IN1(WX8523), .IN2(U5950_n1), .Q(WX8586) );
  INVX0 U5950_U1 ( .INP(n9615), .ZN(U5950_n1) );
  AND2X1 U5951_U2 ( .IN1(WX8521), .IN2(U5951_n1), .Q(WX8584) );
  INVX0 U5951_U1 ( .INP(n9615), .ZN(U5951_n1) );
  AND2X1 U5952_U2 ( .IN1(WX8519), .IN2(U5952_n1), .Q(WX8582) );
  INVX0 U5952_U1 ( .INP(n9615), .ZN(U5952_n1) );
  AND2X1 U5953_U2 ( .IN1(WX8517), .IN2(U5953_n1), .Q(WX8580) );
  INVX0 U5953_U1 ( .INP(n9615), .ZN(U5953_n1) );
  AND2X1 U5954_U2 ( .IN1(WX8515), .IN2(U5954_n1), .Q(WX8578) );
  INVX0 U5954_U1 ( .INP(n9615), .ZN(U5954_n1) );
  AND2X1 U5955_U2 ( .IN1(WX8513), .IN2(U5955_n1), .Q(WX8576) );
  INVX0 U5955_U1 ( .INP(n9615), .ZN(U5955_n1) );
  AND2X1 U5956_U2 ( .IN1(WX8511), .IN2(U5956_n1), .Q(WX8574) );
  INVX0 U5956_U1 ( .INP(n9615), .ZN(U5956_n1) );
  AND2X1 U5957_U2 ( .IN1(WX8509), .IN2(U5957_n1), .Q(WX8572) );
  INVX0 U5957_U1 ( .INP(n9615), .ZN(U5957_n1) );
  AND2X1 U5958_U2 ( .IN1(WX8507), .IN2(U5958_n1), .Q(WX8570) );
  INVX0 U5958_U1 ( .INP(n9615), .ZN(U5958_n1) );
  AND2X1 U5959_U2 ( .IN1(WX8505), .IN2(U5959_n1), .Q(WX8568) );
  INVX0 U5959_U1 ( .INP(n9615), .ZN(U5959_n1) );
  AND2X1 U5960_U2 ( .IN1(test_so71), .IN2(U5960_n1), .Q(WX8566) );
  INVX0 U5960_U1 ( .INP(n9615), .ZN(U5960_n1) );
  AND2X1 U5961_U2 ( .IN1(WX8501), .IN2(U5961_n1), .Q(WX8564) );
  INVX0 U5961_U1 ( .INP(n9615), .ZN(U5961_n1) );
  AND2X1 U5962_U2 ( .IN1(WX8499), .IN2(U5962_n1), .Q(WX8562) );
  INVX0 U5962_U1 ( .INP(n9614), .ZN(U5962_n1) );
  AND2X1 U5963_U2 ( .IN1(WX8497), .IN2(U5963_n1), .Q(WX8560) );
  INVX0 U5963_U1 ( .INP(n9614), .ZN(U5963_n1) );
  AND2X1 U5964_U2 ( .IN1(WX8495), .IN2(U5964_n1), .Q(WX8558) );
  INVX0 U5964_U1 ( .INP(n9614), .ZN(U5964_n1) );
  AND2X1 U5965_U2 ( .IN1(WX8493), .IN2(U5965_n1), .Q(WX8556) );
  INVX0 U5965_U1 ( .INP(n9614), .ZN(U5965_n1) );
  AND2X1 U5966_U2 ( .IN1(WX8491), .IN2(U5966_n1), .Q(WX8554) );
  INVX0 U5966_U1 ( .INP(n9614), .ZN(U5966_n1) );
  AND2X1 U5967_U2 ( .IN1(WX8489), .IN2(U5967_n1), .Q(WX8552) );
  INVX0 U5967_U1 ( .INP(n9614), .ZN(U5967_n1) );
  AND2X1 U5968_U2 ( .IN1(WX8487), .IN2(U5968_n1), .Q(WX8550) );
  INVX0 U5968_U1 ( .INP(n9614), .ZN(U5968_n1) );
  AND2X1 U5969_U2 ( .IN1(WX8485), .IN2(U5969_n1), .Q(WX8548) );
  INVX0 U5969_U1 ( .INP(n9614), .ZN(U5969_n1) );
  AND2X1 U5970_U2 ( .IN1(WX8483), .IN2(U5970_n1), .Q(WX8546) );
  INVX0 U5970_U1 ( .INP(n9614), .ZN(U5970_n1) );
  AND2X1 U5971_U2 ( .IN1(WX8481), .IN2(U5971_n1), .Q(WX8544) );
  INVX0 U5971_U1 ( .INP(n9614), .ZN(U5971_n1) );
  AND2X1 U5972_U2 ( .IN1(WX8479), .IN2(U5972_n1), .Q(WX8542) );
  INVX0 U5972_U1 ( .INP(n9614), .ZN(U5972_n1) );
  AND2X1 U5973_U2 ( .IN1(WX8477), .IN2(U5973_n1), .Q(WX8540) );
  INVX0 U5973_U1 ( .INP(n9614), .ZN(U5973_n1) );
  AND2X1 U5974_U2 ( .IN1(WX8475), .IN2(U5974_n1), .Q(WX8538) );
  INVX0 U5974_U1 ( .INP(n9614), .ZN(U5974_n1) );
  AND2X1 U5975_U2 ( .IN1(WX8473), .IN2(U5975_n1), .Q(WX8536) );
  INVX0 U5975_U1 ( .INP(n9614), .ZN(U5975_n1) );
  AND2X1 U5976_U2 ( .IN1(WX8471), .IN2(U5976_n1), .Q(WX8534) );
  INVX0 U5976_U1 ( .INP(n9613), .ZN(U5976_n1) );
  AND2X1 U5977_U2 ( .IN1(test_so70), .IN2(U5977_n1), .Q(WX8532) );
  INVX0 U5977_U1 ( .INP(n9613), .ZN(U5977_n1) );
  AND2X1 U5978_U2 ( .IN1(WX8467), .IN2(U5978_n1), .Q(WX8530) );
  INVX0 U5978_U1 ( .INP(n9613), .ZN(U5978_n1) );
  AND2X1 U5979_U2 ( .IN1(WX8465), .IN2(U5979_n1), .Q(WX8528) );
  INVX0 U5979_U1 ( .INP(n9613), .ZN(U5979_n1) );
  AND2X1 U5980_U2 ( .IN1(WX8463), .IN2(U5980_n1), .Q(WX8526) );
  INVX0 U5980_U1 ( .INP(n9613), .ZN(U5980_n1) );
  AND2X1 U5981_U2 ( .IN1(WX8461), .IN2(U5981_n1), .Q(WX8524) );
  INVX0 U5981_U1 ( .INP(n9613), .ZN(U5981_n1) );
  AND2X1 U5982_U2 ( .IN1(WX8459), .IN2(U5982_n1), .Q(WX8522) );
  INVX0 U5982_U1 ( .INP(n9613), .ZN(U5982_n1) );
  AND2X1 U5983_U2 ( .IN1(WX8457), .IN2(U5983_n1), .Q(WX8520) );
  INVX0 U5983_U1 ( .INP(n9613), .ZN(U5983_n1) );
  AND2X1 U5984_U2 ( .IN1(WX8455), .IN2(U5984_n1), .Q(WX8518) );
  INVX0 U5984_U1 ( .INP(n9613), .ZN(U5984_n1) );
  AND2X1 U5985_U2 ( .IN1(WX8453), .IN2(U5985_n1), .Q(WX8516) );
  INVX0 U5985_U1 ( .INP(n9613), .ZN(U5985_n1) );
  AND2X1 U5986_U2 ( .IN1(WX8451), .IN2(U5986_n1), .Q(WX8514) );
  INVX0 U5986_U1 ( .INP(n9613), .ZN(U5986_n1) );
  AND2X1 U5987_U2 ( .IN1(WX8449), .IN2(U5987_n1), .Q(WX8512) );
  INVX0 U5987_U1 ( .INP(n9613), .ZN(U5987_n1) );
  AND2X1 U5988_U2 ( .IN1(WX8447), .IN2(U5988_n1), .Q(WX8510) );
  INVX0 U5988_U1 ( .INP(n9613), .ZN(U5988_n1) );
  AND2X1 U5989_U2 ( .IN1(WX8445), .IN2(U5989_n1), .Q(WX8508) );
  INVX0 U5989_U1 ( .INP(n9613), .ZN(U5989_n1) );
  AND2X1 U5990_U2 ( .IN1(WX8443), .IN2(U5990_n1), .Q(WX8506) );
  INVX0 U5990_U1 ( .INP(n9612), .ZN(U5990_n1) );
  AND2X1 U5991_U2 ( .IN1(WX8441), .IN2(U5991_n1), .Q(WX8504) );
  INVX0 U5991_U1 ( .INP(n9612), .ZN(U5991_n1) );
  AND2X1 U5992_U2 ( .IN1(WX8439), .IN2(U5992_n1), .Q(WX8502) );
  INVX0 U5992_U1 ( .INP(n9612), .ZN(U5992_n1) );
  AND2X1 U5993_U2 ( .IN1(WX8437), .IN2(U5993_n1), .Q(WX8500) );
  INVX0 U5993_U1 ( .INP(n9612), .ZN(U5993_n1) );
  AND2X1 U5994_U2 ( .IN1(test_so69), .IN2(U5994_n1), .Q(WX8498) );
  INVX0 U5994_U1 ( .INP(n9612), .ZN(U5994_n1) );
  AND2X1 U5995_U2 ( .IN1(WX7300), .IN2(U5995_n1), .Q(WX7363) );
  INVX0 U5995_U1 ( .INP(n9612), .ZN(U5995_n1) );
  AND2X1 U5996_U2 ( .IN1(WX7298), .IN2(U5996_n1), .Q(WX7361) );
  INVX0 U5996_U1 ( .INP(n9612), .ZN(U5996_n1) );
  AND2X1 U5997_U2 ( .IN1(WX7296), .IN2(U5997_n1), .Q(WX7359) );
  INVX0 U5997_U1 ( .INP(n9612), .ZN(U5997_n1) );
  AND2X1 U5998_U2 ( .IN1(WX7294), .IN2(U5998_n1), .Q(WX7357) );
  INVX0 U5998_U1 ( .INP(n9612), .ZN(U5998_n1) );
  AND2X1 U5999_U2 ( .IN1(WX7292), .IN2(U5999_n1), .Q(WX7355) );
  INVX0 U5999_U1 ( .INP(n9612), .ZN(U5999_n1) );
  AND2X1 U6000_U2 ( .IN1(WX7290), .IN2(U6000_n1), .Q(WX7353) );
  INVX0 U6000_U1 ( .INP(n9612), .ZN(U6000_n1) );
  AND2X1 U6001_U2 ( .IN1(test_so62), .IN2(U6001_n1), .Q(WX7351) );
  INVX0 U6001_U1 ( .INP(n9612), .ZN(U6001_n1) );
  AND2X1 U6002_U2 ( .IN1(WX7286), .IN2(U6002_n1), .Q(WX7349) );
  INVX0 U6002_U1 ( .INP(n9612), .ZN(U6002_n1) );
  AND2X1 U6003_U2 ( .IN1(WX7284), .IN2(U6003_n1), .Q(WX7347) );
  INVX0 U6003_U1 ( .INP(n9612), .ZN(U6003_n1) );
  AND2X1 U6004_U2 ( .IN1(WX7282), .IN2(U6004_n1), .Q(WX7345) );
  INVX0 U6004_U1 ( .INP(n9611), .ZN(U6004_n1) );
  AND2X1 U6005_U2 ( .IN1(WX7280), .IN2(U6005_n1), .Q(WX7343) );
  INVX0 U6005_U1 ( .INP(n9611), .ZN(U6005_n1) );
  AND2X1 U6006_U2 ( .IN1(WX7278), .IN2(U6006_n1), .Q(WX7341) );
  INVX0 U6006_U1 ( .INP(n9611), .ZN(U6006_n1) );
  AND2X1 U6007_U2 ( .IN1(WX7276), .IN2(U6007_n1), .Q(WX7339) );
  INVX0 U6007_U1 ( .INP(n9611), .ZN(U6007_n1) );
  AND2X1 U6008_U2 ( .IN1(WX7274), .IN2(U6008_n1), .Q(WX7337) );
  INVX0 U6008_U1 ( .INP(n9611), .ZN(U6008_n1) );
  AND2X1 U6009_U2 ( .IN1(WX7272), .IN2(U6009_n1), .Q(WX7335) );
  INVX0 U6009_U1 ( .INP(n9611), .ZN(U6009_n1) );
  AND2X1 U6010_U2 ( .IN1(WX7270), .IN2(U6010_n1), .Q(WX7333) );
  INVX0 U6010_U1 ( .INP(n9611), .ZN(U6010_n1) );
  AND2X1 U6011_U2 ( .IN1(WX7268), .IN2(U6011_n1), .Q(WX7331) );
  INVX0 U6011_U1 ( .INP(n9611), .ZN(U6011_n1) );
  AND2X1 U6012_U2 ( .IN1(WX7266), .IN2(U6012_n1), .Q(WX7329) );
  INVX0 U6012_U1 ( .INP(n9611), .ZN(U6012_n1) );
  AND2X1 U6013_U2 ( .IN1(WX7264), .IN2(U6013_n1), .Q(WX7327) );
  INVX0 U6013_U1 ( .INP(n9611), .ZN(U6013_n1) );
  AND2X1 U6014_U2 ( .IN1(WX7262), .IN2(U6014_n1), .Q(WX7325) );
  INVX0 U6014_U1 ( .INP(n9611), .ZN(U6014_n1) );
  AND2X1 U6015_U2 ( .IN1(WX7260), .IN2(U6015_n1), .Q(WX7323) );
  INVX0 U6015_U1 ( .INP(n9611), .ZN(U6015_n1) );
  AND2X1 U6016_U2 ( .IN1(WX7258), .IN2(U6016_n1), .Q(WX7321) );
  INVX0 U6016_U1 ( .INP(n9611), .ZN(U6016_n1) );
  AND2X1 U6017_U2 ( .IN1(WX7256), .IN2(U6017_n1), .Q(WX7319) );
  INVX0 U6017_U1 ( .INP(n9611), .ZN(U6017_n1) );
  AND2X1 U6018_U2 ( .IN1(test_so61), .IN2(U6018_n1), .Q(WX7317) );
  INVX0 U6018_U1 ( .INP(n9610), .ZN(U6018_n1) );
  AND2X1 U6019_U2 ( .IN1(WX7252), .IN2(U6019_n1), .Q(WX7315) );
  INVX0 U6019_U1 ( .INP(n9610), .ZN(U6019_n1) );
  AND2X1 U6020_U2 ( .IN1(WX7250), .IN2(U6020_n1), .Q(WX7313) );
  INVX0 U6020_U1 ( .INP(n9610), .ZN(U6020_n1) );
  AND2X1 U6021_U2 ( .IN1(WX7248), .IN2(U6021_n1), .Q(WX7311) );
  INVX0 U6021_U1 ( .INP(n9610), .ZN(U6021_n1) );
  AND2X1 U6022_U2 ( .IN1(WX7246), .IN2(U6022_n1), .Q(WX7309) );
  INVX0 U6022_U1 ( .INP(n9610), .ZN(U6022_n1) );
  AND2X1 U6023_U2 ( .IN1(WX7244), .IN2(U6023_n1), .Q(WX7307) );
  INVX0 U6023_U1 ( .INP(n9610), .ZN(U6023_n1) );
  AND2X1 U6024_U2 ( .IN1(WX7242), .IN2(U6024_n1), .Q(WX7305) );
  INVX0 U6024_U1 ( .INP(n9610), .ZN(U6024_n1) );
  AND2X1 U6025_U2 ( .IN1(WX7240), .IN2(U6025_n1), .Q(WX7303) );
  INVX0 U6025_U1 ( .INP(n9610), .ZN(U6025_n1) );
  AND2X1 U6026_U2 ( .IN1(WX7238), .IN2(U6026_n1), .Q(WX7301) );
  INVX0 U6026_U1 ( .INP(n9610), .ZN(U6026_n1) );
  AND2X1 U6027_U2 ( .IN1(WX7236), .IN2(U6027_n1), .Q(WX7299) );
  INVX0 U6027_U1 ( .INP(n9610), .ZN(U6027_n1) );
  AND2X1 U6028_U2 ( .IN1(WX7234), .IN2(U6028_n1), .Q(WX7297) );
  INVX0 U6028_U1 ( .INP(n9610), .ZN(U6028_n1) );
  AND2X1 U6029_U2 ( .IN1(WX7232), .IN2(U6029_n1), .Q(WX7295) );
  INVX0 U6029_U1 ( .INP(n9610), .ZN(U6029_n1) );
  AND2X1 U6030_U2 ( .IN1(WX7230), .IN2(U6030_n1), .Q(WX7293) );
  INVX0 U6030_U1 ( .INP(n9610), .ZN(U6030_n1) );
  AND2X1 U6031_U2 ( .IN1(WX7228), .IN2(U6031_n1), .Q(WX7291) );
  INVX0 U6031_U1 ( .INP(n9610), .ZN(U6031_n1) );
  AND2X1 U6032_U2 ( .IN1(WX7226), .IN2(U6032_n1), .Q(WX7289) );
  INVX0 U6032_U1 ( .INP(n9609), .ZN(U6032_n1) );
  AND2X1 U6033_U2 ( .IN1(WX7224), .IN2(U6033_n1), .Q(WX7287) );
  INVX0 U6033_U1 ( .INP(n9609), .ZN(U6033_n1) );
  AND2X1 U6034_U2 ( .IN1(WX7222), .IN2(U6034_n1), .Q(WX7285) );
  INVX0 U6034_U1 ( .INP(n9609), .ZN(U6034_n1) );
  AND2X1 U6035_U2 ( .IN1(test_so60), .IN2(U6035_n1), .Q(WX7283) );
  INVX0 U6035_U1 ( .INP(n9609), .ZN(U6035_n1) );
  AND2X1 U6036_U2 ( .IN1(WX7218), .IN2(U6036_n1), .Q(WX7281) );
  INVX0 U6036_U1 ( .INP(n9609), .ZN(U6036_n1) );
  AND2X1 U6037_U2 ( .IN1(WX7216), .IN2(U6037_n1), .Q(WX7279) );
  INVX0 U6037_U1 ( .INP(n9609), .ZN(U6037_n1) );
  AND2X1 U6038_U2 ( .IN1(WX7214), .IN2(U6038_n1), .Q(WX7277) );
  INVX0 U6038_U1 ( .INP(n9609), .ZN(U6038_n1) );
  AND2X1 U6039_U2 ( .IN1(WX7212), .IN2(U6039_n1), .Q(WX7275) );
  INVX0 U6039_U1 ( .INP(n9609), .ZN(U6039_n1) );
  AND2X1 U6040_U2 ( .IN1(WX7210), .IN2(U6040_n1), .Q(WX7273) );
  INVX0 U6040_U1 ( .INP(n9609), .ZN(U6040_n1) );
  AND2X1 U6041_U2 ( .IN1(WX7208), .IN2(U6041_n1), .Q(WX7271) );
  INVX0 U6041_U1 ( .INP(n9609), .ZN(U6041_n1) );
  AND2X1 U6042_U2 ( .IN1(WX7206), .IN2(U6042_n1), .Q(WX7269) );
  INVX0 U6042_U1 ( .INP(n9609), .ZN(U6042_n1) );
  AND2X1 U6043_U2 ( .IN1(WX7204), .IN2(U6043_n1), .Q(WX7267) );
  INVX0 U6043_U1 ( .INP(n9609), .ZN(U6043_n1) );
  AND2X1 U6044_U2 ( .IN1(WX7202), .IN2(U6044_n1), .Q(WX7265) );
  INVX0 U6044_U1 ( .INP(n9609), .ZN(U6044_n1) );
  AND2X1 U6045_U2 ( .IN1(WX7200), .IN2(U6045_n1), .Q(WX7263) );
  INVX0 U6045_U1 ( .INP(n9609), .ZN(U6045_n1) );
  AND2X1 U6046_U2 ( .IN1(WX7198), .IN2(U6046_n1), .Q(WX7261) );
  INVX0 U6046_U1 ( .INP(n9608), .ZN(U6046_n1) );
  AND2X1 U6047_U2 ( .IN1(WX7196), .IN2(U6047_n1), .Q(WX7259) );
  INVX0 U6047_U1 ( .INP(n9608), .ZN(U6047_n1) );
  AND2X1 U6048_U2 ( .IN1(WX7194), .IN2(U6048_n1), .Q(WX7257) );
  INVX0 U6048_U1 ( .INP(n9608), .ZN(U6048_n1) );
  AND2X1 U6049_U2 ( .IN1(WX7192), .IN2(U6049_n1), .Q(WX7255) );
  INVX0 U6049_U1 ( .INP(n9608), .ZN(U6049_n1) );
  AND2X1 U6050_U2 ( .IN1(WX7190), .IN2(U6050_n1), .Q(WX7253) );
  INVX0 U6050_U1 ( .INP(n9608), .ZN(U6050_n1) );
  AND2X1 U6051_U2 ( .IN1(WX7188), .IN2(U6051_n1), .Q(WX7251) );
  INVX0 U6051_U1 ( .INP(n9608), .ZN(U6051_n1) );
  AND2X1 U6052_U2 ( .IN1(test_so59), .IN2(U6052_n1), .Q(WX7249) );
  INVX0 U6052_U1 ( .INP(n9608), .ZN(U6052_n1) );
  AND2X1 U6053_U2 ( .IN1(WX7184), .IN2(U6053_n1), .Q(WX7247) );
  INVX0 U6053_U1 ( .INP(n9608), .ZN(U6053_n1) );
  AND2X1 U6054_U2 ( .IN1(WX7182), .IN2(U6054_n1), .Q(WX7245) );
  INVX0 U6054_U1 ( .INP(n9608), .ZN(U6054_n1) );
  AND2X1 U6055_U2 ( .IN1(WX7180), .IN2(U6055_n1), .Q(WX7243) );
  INVX0 U6055_U1 ( .INP(n9608), .ZN(U6055_n1) );
  AND2X1 U6056_U2 ( .IN1(WX7178), .IN2(U6056_n1), .Q(WX7241) );
  INVX0 U6056_U1 ( .INP(n9608), .ZN(U6056_n1) );
  AND2X1 U6057_U2 ( .IN1(WX7176), .IN2(U6057_n1), .Q(WX7239) );
  INVX0 U6057_U1 ( .INP(n9608), .ZN(U6057_n1) );
  AND2X1 U6058_U2 ( .IN1(WX7174), .IN2(U6058_n1), .Q(WX7237) );
  INVX0 U6058_U1 ( .INP(n9608), .ZN(U6058_n1) );
  AND2X1 U6059_U2 ( .IN1(WX7172), .IN2(U6059_n1), .Q(WX7235) );
  INVX0 U6059_U1 ( .INP(n9608), .ZN(U6059_n1) );
  AND2X1 U6060_U2 ( .IN1(WX7170), .IN2(U6060_n1), .Q(WX7233) );
  INVX0 U6060_U1 ( .INP(n9607), .ZN(U6060_n1) );
  AND2X1 U6061_U2 ( .IN1(WX7168), .IN2(U6061_n1), .Q(WX7231) );
  INVX0 U6061_U1 ( .INP(n9607), .ZN(U6061_n1) );
  AND2X1 U6062_U2 ( .IN1(WX7166), .IN2(U6062_n1), .Q(WX7229) );
  INVX0 U6062_U1 ( .INP(n9607), .ZN(U6062_n1) );
  AND2X1 U6063_U2 ( .IN1(WX7164), .IN2(U6063_n1), .Q(WX7227) );
  INVX0 U6063_U1 ( .INP(n9607), .ZN(U6063_n1) );
  AND2X1 U6064_U2 ( .IN1(WX7162), .IN2(U6064_n1), .Q(WX7225) );
  INVX0 U6064_U1 ( .INP(n9607), .ZN(U6064_n1) );
  AND2X1 U6065_U2 ( .IN1(WX7160), .IN2(U6065_n1), .Q(WX7223) );
  INVX0 U6065_U1 ( .INP(n9607), .ZN(U6065_n1) );
  AND2X1 U6066_U2 ( .IN1(WX7158), .IN2(U6066_n1), .Q(WX7221) );
  INVX0 U6066_U1 ( .INP(n9607), .ZN(U6066_n1) );
  AND2X1 U6067_U2 ( .IN1(WX7156), .IN2(U6067_n1), .Q(WX7219) );
  INVX0 U6067_U1 ( .INP(n9607), .ZN(U6067_n1) );
  AND2X1 U6068_U2 ( .IN1(WX7154), .IN2(U6068_n1), .Q(WX7217) );
  INVX0 U6068_U1 ( .INP(n9607), .ZN(U6068_n1) );
  AND2X1 U6069_U2 ( .IN1(test_so58), .IN2(U6069_n1), .Q(WX7215) );
  INVX0 U6069_U1 ( .INP(n9607), .ZN(U6069_n1) );
  AND2X1 U6070_U2 ( .IN1(WX7150), .IN2(U6070_n1), .Q(WX7213) );
  INVX0 U6070_U1 ( .INP(n9607), .ZN(U6070_n1) );
  AND2X1 U6071_U2 ( .IN1(WX7148), .IN2(U6071_n1), .Q(WX7211) );
  INVX0 U6071_U1 ( .INP(n9607), .ZN(U6071_n1) );
  AND2X1 U6072_U2 ( .IN1(WX7146), .IN2(U6072_n1), .Q(WX7209) );
  INVX0 U6072_U1 ( .INP(n9607), .ZN(U6072_n1) );
  AND2X1 U6073_U2 ( .IN1(WX7144), .IN2(U6073_n1), .Q(WX7207) );
  INVX0 U6073_U1 ( .INP(n9607), .ZN(U6073_n1) );
  AND2X1 U6074_U2 ( .IN1(WX7142), .IN2(U6074_n1), .Q(WX7205) );
  INVX0 U6074_U1 ( .INP(n9606), .ZN(U6074_n1) );
  AND2X1 U6075_U2 ( .IN1(WX6007), .IN2(U6075_n1), .Q(WX6070) );
  INVX0 U6075_U1 ( .INP(n9606), .ZN(U6075_n1) );
  AND2X1 U6076_U2 ( .IN1(test_so51), .IN2(U6076_n1), .Q(WX6068) );
  INVX0 U6076_U1 ( .INP(n9606), .ZN(U6076_n1) );
  AND2X1 U6077_U2 ( .IN1(WX6003), .IN2(U6077_n1), .Q(WX6066) );
  INVX0 U6077_U1 ( .INP(n9606), .ZN(U6077_n1) );
  AND2X1 U6078_U2 ( .IN1(WX6001), .IN2(U6078_n1), .Q(WX6064) );
  INVX0 U6078_U1 ( .INP(n9606), .ZN(U6078_n1) );
  AND2X1 U6079_U2 ( .IN1(WX5999), .IN2(U6079_n1), .Q(WX6062) );
  INVX0 U6079_U1 ( .INP(n9606), .ZN(U6079_n1) );
  AND2X1 U6080_U2 ( .IN1(WX5997), .IN2(U6080_n1), .Q(WX6060) );
  INVX0 U6080_U1 ( .INP(n9606), .ZN(U6080_n1) );
  AND2X1 U6081_U2 ( .IN1(WX5995), .IN2(U6081_n1), .Q(WX6058) );
  INVX0 U6081_U1 ( .INP(n9606), .ZN(U6081_n1) );
  AND2X1 U6082_U2 ( .IN1(WX5993), .IN2(U6082_n1), .Q(WX6056) );
  INVX0 U6082_U1 ( .INP(n9606), .ZN(U6082_n1) );
  AND2X1 U6083_U2 ( .IN1(WX5991), .IN2(U6083_n1), .Q(WX6054) );
  INVX0 U6083_U1 ( .INP(n9606), .ZN(U6083_n1) );
  AND2X1 U6084_U2 ( .IN1(WX5989), .IN2(U6084_n1), .Q(WX6052) );
  INVX0 U6084_U1 ( .INP(n9606), .ZN(U6084_n1) );
  AND2X1 U6085_U2 ( .IN1(WX5987), .IN2(U6085_n1), .Q(WX6050) );
  INVX0 U6085_U1 ( .INP(n9606), .ZN(U6085_n1) );
  AND2X1 U6086_U2 ( .IN1(WX5985), .IN2(U6086_n1), .Q(WX6048) );
  INVX0 U6086_U1 ( .INP(n9606), .ZN(U6086_n1) );
  AND2X1 U6087_U2 ( .IN1(WX5983), .IN2(U6087_n1), .Q(WX6046) );
  INVX0 U6087_U1 ( .INP(n9606), .ZN(U6087_n1) );
  AND2X1 U6088_U2 ( .IN1(WX5981), .IN2(U6088_n1), .Q(WX6044) );
  INVX0 U6088_U1 ( .INP(n9605), .ZN(U6088_n1) );
  AND2X1 U6089_U2 ( .IN1(WX5979), .IN2(U6089_n1), .Q(WX6042) );
  INVX0 U6089_U1 ( .INP(n9605), .ZN(U6089_n1) );
  AND2X1 U6090_U2 ( .IN1(WX5977), .IN2(U6090_n1), .Q(WX6040) );
  INVX0 U6090_U1 ( .INP(n9605), .ZN(U6090_n1) );
  AND2X1 U6091_U2 ( .IN1(WX5975), .IN2(U6091_n1), .Q(WX6038) );
  INVX0 U6091_U1 ( .INP(n9605), .ZN(U6091_n1) );
  AND2X1 U6092_U2 ( .IN1(WX5973), .IN2(U6092_n1), .Q(WX6036) );
  INVX0 U6092_U1 ( .INP(n9605), .ZN(U6092_n1) );
  AND2X1 U6093_U2 ( .IN1(test_so50), .IN2(U6093_n1), .Q(WX6034) );
  INVX0 U6093_U1 ( .INP(n9605), .ZN(U6093_n1) );
  AND2X1 U6094_U2 ( .IN1(WX5969), .IN2(U6094_n1), .Q(WX6032) );
  INVX0 U6094_U1 ( .INP(n9605), .ZN(U6094_n1) );
  AND2X1 U6095_U2 ( .IN1(WX5967), .IN2(U6095_n1), .Q(WX6030) );
  INVX0 U6095_U1 ( .INP(n9605), .ZN(U6095_n1) );
  AND2X1 U6096_U2 ( .IN1(WX5965), .IN2(U6096_n1), .Q(WX6028) );
  INVX0 U6096_U1 ( .INP(n9605), .ZN(U6096_n1) );
  AND2X1 U6097_U2 ( .IN1(WX5963), .IN2(U6097_n1), .Q(WX6026) );
  INVX0 U6097_U1 ( .INP(n9605), .ZN(U6097_n1) );
  AND2X1 U6098_U2 ( .IN1(WX5961), .IN2(U6098_n1), .Q(WX6024) );
  INVX0 U6098_U1 ( .INP(n9605), .ZN(U6098_n1) );
  AND2X1 U6099_U2 ( .IN1(WX5959), .IN2(U6099_n1), .Q(WX6022) );
  INVX0 U6099_U1 ( .INP(n9605), .ZN(U6099_n1) );
  AND2X1 U6100_U2 ( .IN1(WX5957), .IN2(U6100_n1), .Q(WX6020) );
  INVX0 U6100_U1 ( .INP(n9605), .ZN(U6100_n1) );
  AND2X1 U6101_U2 ( .IN1(WX5955), .IN2(U6101_n1), .Q(WX6018) );
  INVX0 U6101_U1 ( .INP(n9605), .ZN(U6101_n1) );
  AND2X1 U6102_U2 ( .IN1(WX5953), .IN2(U6102_n1), .Q(WX6016) );
  INVX0 U6102_U1 ( .INP(n9604), .ZN(U6102_n1) );
  AND2X1 U6103_U2 ( .IN1(WX5951), .IN2(U6103_n1), .Q(WX6014) );
  INVX0 U6103_U1 ( .INP(n9604), .ZN(U6103_n1) );
  AND2X1 U6104_U2 ( .IN1(WX5949), .IN2(U6104_n1), .Q(WX6012) );
  INVX0 U6104_U1 ( .INP(n9604), .ZN(U6104_n1) );
  AND2X1 U6105_U2 ( .IN1(WX5947), .IN2(U6105_n1), .Q(WX6010) );
  INVX0 U6105_U1 ( .INP(n9604), .ZN(U6105_n1) );
  AND2X1 U6106_U2 ( .IN1(WX5945), .IN2(U6106_n1), .Q(WX6008) );
  INVX0 U6106_U1 ( .INP(n9604), .ZN(U6106_n1) );
  AND2X1 U6107_U2 ( .IN1(WX5943), .IN2(U6107_n1), .Q(WX6006) );
  INVX0 U6107_U1 ( .INP(n9604), .ZN(U6107_n1) );
  AND2X1 U6108_U2 ( .IN1(WX5941), .IN2(U6108_n1), .Q(WX6004) );
  INVX0 U6108_U1 ( .INP(n9604), .ZN(U6108_n1) );
  AND2X1 U6109_U2 ( .IN1(WX5929), .IN2(U6109_n1), .Q(WX5992) );
  INVX0 U6109_U1 ( .INP(n9604), .ZN(U6109_n1) );
  AND2X1 U6110_U2 ( .IN1(WX5927), .IN2(U6110_n1), .Q(WX5990) );
  INVX0 U6110_U1 ( .INP(n9604), .ZN(U6110_n1) );
  AND2X1 U6111_U2 ( .IN1(WX5925), .IN2(U6111_n1), .Q(WX5988) );
  INVX0 U6111_U1 ( .INP(n9604), .ZN(U6111_n1) );
  AND2X1 U6112_U2 ( .IN1(WX5923), .IN2(U6112_n1), .Q(WX5986) );
  INVX0 U6112_U1 ( .INP(n9604), .ZN(U6112_n1) );
  AND2X1 U6113_U2 ( .IN1(WX5921), .IN2(U6113_n1), .Q(WX5984) );
  INVX0 U6113_U1 ( .INP(n9604), .ZN(U6113_n1) );
  AND2X1 U6114_U2 ( .IN1(WX5919), .IN2(U6114_n1), .Q(WX5982) );
  INVX0 U6114_U1 ( .INP(n9604), .ZN(U6114_n1) );
  AND2X1 U6115_U2 ( .IN1(WX5917), .IN2(U6115_n1), .Q(WX5980) );
  INVX0 U6115_U1 ( .INP(n9604), .ZN(U6115_n1) );
  AND2X1 U6116_U2 ( .IN1(WX5915), .IN2(U6116_n1), .Q(WX5978) );
  INVX0 U6116_U1 ( .INP(n9603), .ZN(U6116_n1) );
  AND2X1 U6117_U2 ( .IN1(WX5913), .IN2(U6117_n1), .Q(WX5976) );
  INVX0 U6117_U1 ( .INP(n9603), .ZN(U6117_n1) );
  AND2X1 U6118_U2 ( .IN1(WX5911), .IN2(U6118_n1), .Q(WX5974) );
  INVX0 U6118_U1 ( .INP(n9603), .ZN(U6118_n1) );
  AND2X1 U6119_U2 ( .IN1(WX5909), .IN2(U6119_n1), .Q(WX5972) );
  INVX0 U6119_U1 ( .INP(n9603), .ZN(U6119_n1) );
  AND2X1 U6120_U2 ( .IN1(WX5907), .IN2(U6120_n1), .Q(WX5970) );
  INVX0 U6120_U1 ( .INP(n9603), .ZN(U6120_n1) );
  AND2X1 U6121_U2 ( .IN1(WX5905), .IN2(U6121_n1), .Q(WX5968) );
  INVX0 U6121_U1 ( .INP(n9603), .ZN(U6121_n1) );
  AND2X1 U6122_U2 ( .IN1(test_so48), .IN2(U6122_n1), .Q(WX5966) );
  INVX0 U6122_U1 ( .INP(n9603), .ZN(U6122_n1) );
  AND2X1 U6123_U2 ( .IN1(WX5901), .IN2(U6123_n1), .Q(WX5964) );
  INVX0 U6123_U1 ( .INP(n9603), .ZN(U6123_n1) );
  AND2X1 U6124_U2 ( .IN1(WX5899), .IN2(U6124_n1), .Q(WX5962) );
  INVX0 U6124_U1 ( .INP(n9603), .ZN(U6124_n1) );
  AND2X1 U6125_U2 ( .IN1(WX5897), .IN2(U6125_n1), .Q(WX5960) );
  INVX0 U6125_U1 ( .INP(n9603), .ZN(U6125_n1) );
  AND2X1 U6126_U2 ( .IN1(WX5895), .IN2(U6126_n1), .Q(WX5958) );
  INVX0 U6126_U1 ( .INP(n9603), .ZN(U6126_n1) );
  AND2X1 U6127_U2 ( .IN1(WX5893), .IN2(U6127_n1), .Q(WX5956) );
  INVX0 U6127_U1 ( .INP(n9603), .ZN(U6127_n1) );
  AND2X1 U6128_U2 ( .IN1(WX5891), .IN2(U6128_n1), .Q(WX5954) );
  INVX0 U6128_U1 ( .INP(n9603), .ZN(U6128_n1) );
  AND2X1 U6129_U2 ( .IN1(WX5889), .IN2(U6129_n1), .Q(WX5952) );
  INVX0 U6129_U1 ( .INP(n9603), .ZN(U6129_n1) );
  AND2X1 U6130_U2 ( .IN1(WX5887), .IN2(U6130_n1), .Q(WX5950) );
  INVX0 U6130_U1 ( .INP(n9602), .ZN(U6130_n1) );
  AND2X1 U6131_U2 ( .IN1(WX5885), .IN2(U6131_n1), .Q(WX5948) );
  INVX0 U6131_U1 ( .INP(n9602), .ZN(U6131_n1) );
  AND2X1 U6132_U2 ( .IN1(WX5883), .IN2(U6132_n1), .Q(WX5946) );
  INVX0 U6132_U1 ( .INP(n9602), .ZN(U6132_n1) );
  AND2X1 U6133_U2 ( .IN1(WX5881), .IN2(U6133_n1), .Q(WX5944) );
  INVX0 U6133_U1 ( .INP(n9602), .ZN(U6133_n1) );
  AND2X1 U6134_U2 ( .IN1(WX5879), .IN2(U6134_n1), .Q(WX5942) );
  INVX0 U6134_U1 ( .INP(n9602), .ZN(U6134_n1) );
  AND2X1 U6135_U2 ( .IN1(WX5877), .IN2(U6135_n1), .Q(WX5940) );
  INVX0 U6135_U1 ( .INP(n9602), .ZN(U6135_n1) );
  AND2X1 U6136_U2 ( .IN1(WX5875), .IN2(U6136_n1), .Q(WX5938) );
  INVX0 U6136_U1 ( .INP(n9602), .ZN(U6136_n1) );
  AND2X1 U6137_U2 ( .IN1(WX5873), .IN2(U6137_n1), .Q(WX5936) );
  INVX0 U6137_U1 ( .INP(n9602), .ZN(U6137_n1) );
  AND2X1 U6138_U2 ( .IN1(WX5871), .IN2(U6138_n1), .Q(WX5934) );
  INVX0 U6138_U1 ( .INP(n9602), .ZN(U6138_n1) );
  AND2X1 U6139_U2 ( .IN1(test_so47), .IN2(U6139_n1), .Q(WX5932) );
  INVX0 U6139_U1 ( .INP(n9602), .ZN(U6139_n1) );
  AND2X1 U6140_U2 ( .IN1(WX5867), .IN2(U6140_n1), .Q(WX5930) );
  INVX0 U6140_U1 ( .INP(n9602), .ZN(U6140_n1) );
  AND2X1 U6141_U2 ( .IN1(WX5865), .IN2(U6141_n1), .Q(WX5928) );
  INVX0 U6141_U1 ( .INP(n9602), .ZN(U6141_n1) );
  AND2X1 U6142_U2 ( .IN1(WX5863), .IN2(U6142_n1), .Q(WX5926) );
  INVX0 U6142_U1 ( .INP(n9602), .ZN(U6142_n1) );
  AND2X1 U6143_U2 ( .IN1(WX5861), .IN2(U6143_n1), .Q(WX5924) );
  INVX0 U6143_U1 ( .INP(n9602), .ZN(U6143_n1) );
  AND2X1 U6144_U2 ( .IN1(WX5859), .IN2(U6144_n1), .Q(WX5922) );
  INVX0 U6144_U1 ( .INP(n9601), .ZN(U6144_n1) );
  AND2X1 U6145_U2 ( .IN1(WX5857), .IN2(U6145_n1), .Q(WX5920) );
  INVX0 U6145_U1 ( .INP(n9601), .ZN(U6145_n1) );
  AND2X1 U6146_U2 ( .IN1(WX5855), .IN2(U6146_n1), .Q(WX5918) );
  INVX0 U6146_U1 ( .INP(n9601), .ZN(U6146_n1) );
  AND2X1 U6147_U2 ( .IN1(WX5853), .IN2(U6147_n1), .Q(WX5916) );
  INVX0 U6147_U1 ( .INP(n9601), .ZN(U6147_n1) );
  AND2X1 U6148_U2 ( .IN1(WX5851), .IN2(U6148_n1), .Q(WX5914) );
  INVX0 U6148_U1 ( .INP(n9601), .ZN(U6148_n1) );
  AND2X1 U6149_U2 ( .IN1(WX5849), .IN2(U6149_n1), .Q(WX5912) );
  INVX0 U6149_U1 ( .INP(n9601), .ZN(U6149_n1) );
  AND2X1 U6150_U2 ( .IN1(WX4714), .IN2(U6150_n1), .Q(WX4777) );
  INVX0 U6150_U1 ( .INP(n9601), .ZN(U6150_n1) );
  AND2X1 U6151_U2 ( .IN1(WX4712), .IN2(U6151_n1), .Q(WX4775) );
  INVX0 U6151_U1 ( .INP(n9601), .ZN(U6151_n1) );
  AND2X1 U6152_U2 ( .IN1(WX4710), .IN2(U6152_n1), .Q(WX4773) );
  INVX0 U6152_U1 ( .INP(n9601), .ZN(U6152_n1) );
  AND2X1 U6153_U2 ( .IN1(WX4708), .IN2(U6153_n1), .Q(WX4771) );
  INVX0 U6153_U1 ( .INP(n9601), .ZN(U6153_n1) );
  AND2X1 U6154_U2 ( .IN1(WX4706), .IN2(U6154_n1), .Q(WX4769) );
  INVX0 U6154_U1 ( .INP(n9601), .ZN(U6154_n1) );
  AND2X1 U6155_U2 ( .IN1(WX4704), .IN2(U6155_n1), .Q(WX4767) );
  INVX0 U6155_U1 ( .INP(n9601), .ZN(U6155_n1) );
  AND2X1 U6156_U2 ( .IN1(WX4702), .IN2(U6156_n1), .Q(WX4765) );
  INVX0 U6156_U1 ( .INP(n9601), .ZN(U6156_n1) );
  AND2X1 U6157_U2 ( .IN1(WX4700), .IN2(U6157_n1), .Q(WX4763) );
  INVX0 U6157_U1 ( .INP(n9601), .ZN(U6157_n1) );
  AND2X1 U6158_U2 ( .IN1(WX4698), .IN2(U6158_n1), .Q(WX4761) );
  INVX0 U6158_U1 ( .INP(n9600), .ZN(U6158_n1) );
  AND2X1 U6159_U2 ( .IN1(WX4696), .IN2(U6159_n1), .Q(WX4759) );
  INVX0 U6159_U1 ( .INP(n9600), .ZN(U6159_n1) );
  AND2X1 U6160_U2 ( .IN1(WX4694), .IN2(U6160_n1), .Q(WX4757) );
  INVX0 U6160_U1 ( .INP(n9600), .ZN(U6160_n1) );
  AND2X1 U6161_U2 ( .IN1(WX4692), .IN2(U6161_n1), .Q(WX4755) );
  INVX0 U6161_U1 ( .INP(n9600), .ZN(U6161_n1) );
  AND2X1 U6162_U2 ( .IN1(WX4690), .IN2(U6162_n1), .Q(WX4753) );
  INVX0 U6162_U1 ( .INP(n9600), .ZN(U6162_n1) );
  AND2X1 U6163_U2 ( .IN1(test_so39), .IN2(U6163_n1), .Q(WX4751) );
  INVX0 U6163_U1 ( .INP(n9600), .ZN(U6163_n1) );
  AND2X1 U6164_U2 ( .IN1(WX4686), .IN2(U6164_n1), .Q(WX4749) );
  INVX0 U6164_U1 ( .INP(n9600), .ZN(U6164_n1) );
  AND2X1 U6165_U2 ( .IN1(WX4684), .IN2(U6165_n1), .Q(WX4747) );
  INVX0 U6165_U1 ( .INP(n9600), .ZN(U6165_n1) );
  AND2X1 U6166_U2 ( .IN1(WX4682), .IN2(U6166_n1), .Q(WX4745) );
  INVX0 U6166_U1 ( .INP(n9600), .ZN(U6166_n1) );
  AND2X1 U6167_U2 ( .IN1(WX4680), .IN2(U6167_n1), .Q(WX4743) );
  INVX0 U6167_U1 ( .INP(n9600), .ZN(U6167_n1) );
  AND2X1 U6168_U2 ( .IN1(WX4678), .IN2(U6168_n1), .Q(WX4741) );
  INVX0 U6168_U1 ( .INP(n9600), .ZN(U6168_n1) );
  AND2X1 U6169_U2 ( .IN1(WX4676), .IN2(U6169_n1), .Q(WX4739) );
  INVX0 U6169_U1 ( .INP(n9600), .ZN(U6169_n1) );
  AND2X1 U6170_U2 ( .IN1(WX4674), .IN2(U6170_n1), .Q(WX4737) );
  INVX0 U6170_U1 ( .INP(n9600), .ZN(U6170_n1) );
  AND2X1 U6171_U2 ( .IN1(WX4672), .IN2(U6171_n1), .Q(WX4735) );
  INVX0 U6171_U1 ( .INP(n9600), .ZN(U6171_n1) );
  AND2X1 U6172_U2 ( .IN1(WX4670), .IN2(U6172_n1), .Q(WX4733) );
  INVX0 U6172_U1 ( .INP(n9599), .ZN(U6172_n1) );
  AND2X1 U6173_U2 ( .IN1(WX4668), .IN2(U6173_n1), .Q(WX4731) );
  INVX0 U6173_U1 ( .INP(n9599), .ZN(U6173_n1) );
  AND2X1 U6174_U2 ( .IN1(WX4666), .IN2(U6174_n1), .Q(WX4729) );
  INVX0 U6174_U1 ( .INP(n9599), .ZN(U6174_n1) );
  AND2X1 U6175_U2 ( .IN1(WX4664), .IN2(U6175_n1), .Q(WX4727) );
  INVX0 U6175_U1 ( .INP(n9599), .ZN(U6175_n1) );
  AND2X1 U6176_U2 ( .IN1(WX4662), .IN2(U6176_n1), .Q(WX4725) );
  INVX0 U6176_U1 ( .INP(n9599), .ZN(U6176_n1) );
  AND2X1 U6177_U2 ( .IN1(WX4660), .IN2(U6177_n1), .Q(WX4723) );
  INVX0 U6177_U1 ( .INP(n9599), .ZN(U6177_n1) );
  AND2X1 U6178_U2 ( .IN1(WX4658), .IN2(U6178_n1), .Q(WX4721) );
  INVX0 U6178_U1 ( .INP(n9599), .ZN(U6178_n1) );
  AND2X1 U6179_U2 ( .IN1(WX4656), .IN2(U6179_n1), .Q(WX4719) );
  INVX0 U6179_U1 ( .INP(n9599), .ZN(U6179_n1) );
  AND2X1 U6180_U2 ( .IN1(test_so38), .IN2(U6180_n1), .Q(WX4717) );
  INVX0 U6180_U1 ( .INP(n9599), .ZN(U6180_n1) );
  AND2X1 U6181_U2 ( .IN1(WX4652), .IN2(U6181_n1), .Q(WX4715) );
  INVX0 U6181_U1 ( .INP(n9599), .ZN(U6181_n1) );
  AND2X1 U6182_U2 ( .IN1(WX4650), .IN2(U6182_n1), .Q(WX4713) );
  INVX0 U6182_U1 ( .INP(n9599), .ZN(U6182_n1) );
  AND2X1 U6183_U2 ( .IN1(WX4648), .IN2(U6183_n1), .Q(WX4711) );
  INVX0 U6183_U1 ( .INP(n9599), .ZN(U6183_n1) );
  AND2X1 U6184_U2 ( .IN1(WX4646), .IN2(U6184_n1), .Q(WX4709) );
  INVX0 U6184_U1 ( .INP(n9599), .ZN(U6184_n1) );
  AND2X1 U6185_U2 ( .IN1(WX4644), .IN2(U6185_n1), .Q(WX4707) );
  INVX0 U6185_U1 ( .INP(n9599), .ZN(U6185_n1) );
  AND2X1 U6186_U2 ( .IN1(WX4642), .IN2(U6186_n1), .Q(WX4705) );
  INVX0 U6186_U1 ( .INP(n9598), .ZN(U6186_n1) );
  AND2X1 U6187_U2 ( .IN1(WX4640), .IN2(U6187_n1), .Q(WX4703) );
  INVX0 U6187_U1 ( .INP(n9598), .ZN(U6187_n1) );
  AND2X1 U6188_U2 ( .IN1(WX4638), .IN2(U6188_n1), .Q(WX4701) );
  INVX0 U6188_U1 ( .INP(n9598), .ZN(U6188_n1) );
  AND2X1 U6189_U2 ( .IN1(WX4636), .IN2(U6189_n1), .Q(WX4699) );
  INVX0 U6189_U1 ( .INP(n9598), .ZN(U6189_n1) );
  AND2X1 U6190_U2 ( .IN1(WX4634), .IN2(U6190_n1), .Q(WX4697) );
  INVX0 U6190_U1 ( .INP(n9598), .ZN(U6190_n1) );
  AND2X1 U6191_U2 ( .IN1(WX4632), .IN2(U6191_n1), .Q(WX4695) );
  INVX0 U6191_U1 ( .INP(n9598), .ZN(U6191_n1) );
  AND2X1 U6192_U2 ( .IN1(WX4630), .IN2(U6192_n1), .Q(WX4693) );
  INVX0 U6192_U1 ( .INP(n9598), .ZN(U6192_n1) );
  AND2X1 U6193_U2 ( .IN1(WX4628), .IN2(U6193_n1), .Q(WX4691) );
  INVX0 U6193_U1 ( .INP(n9598), .ZN(U6193_n1) );
  AND2X1 U6194_U2 ( .IN1(WX4626), .IN2(U6194_n1), .Q(WX4689) );
  INVX0 U6194_U1 ( .INP(n9598), .ZN(U6194_n1) );
  AND2X1 U6195_U2 ( .IN1(WX4624), .IN2(U6195_n1), .Q(WX4687) );
  INVX0 U6195_U1 ( .INP(n9598), .ZN(U6195_n1) );
  AND2X1 U6196_U2 ( .IN1(WX4622), .IN2(U6196_n1), .Q(WX4685) );
  INVX0 U6196_U1 ( .INP(n9598), .ZN(U6196_n1) );
  AND2X1 U6197_U2 ( .IN1(test_so37), .IN2(U6197_n1), .Q(WX4683) );
  INVX0 U6197_U1 ( .INP(n9598), .ZN(U6197_n1) );
  AND2X1 U6198_U2 ( .IN1(WX4618), .IN2(U6198_n1), .Q(WX4681) );
  INVX0 U6198_U1 ( .INP(n9598), .ZN(U6198_n1) );
  AND2X1 U6199_U2 ( .IN1(WX4616), .IN2(U6199_n1), .Q(WX4679) );
  INVX0 U6199_U1 ( .INP(n9598), .ZN(U6199_n1) );
  AND2X1 U6200_U2 ( .IN1(WX4614), .IN2(U6200_n1), .Q(WX4677) );
  INVX0 U6200_U1 ( .INP(n9597), .ZN(U6200_n1) );
  AND2X1 U6201_U2 ( .IN1(WX4612), .IN2(U6201_n1), .Q(WX4675) );
  INVX0 U6201_U1 ( .INP(n9597), .ZN(U6201_n1) );
  AND2X1 U6202_U2 ( .IN1(WX4610), .IN2(U6202_n1), .Q(WX4673) );
  INVX0 U6202_U1 ( .INP(n9597), .ZN(U6202_n1) );
  AND2X1 U6203_U2 ( .IN1(WX4608), .IN2(U6203_n1), .Q(WX4671) );
  INVX0 U6203_U1 ( .INP(n9597), .ZN(U6203_n1) );
  AND2X1 U6204_U2 ( .IN1(WX4606), .IN2(U6204_n1), .Q(WX4669) );
  INVX0 U6204_U1 ( .INP(n9597), .ZN(U6204_n1) );
  AND2X1 U6205_U2 ( .IN1(WX4604), .IN2(U6205_n1), .Q(WX4667) );
  INVX0 U6205_U1 ( .INP(n9597), .ZN(U6205_n1) );
  AND2X1 U6206_U2 ( .IN1(WX4602), .IN2(U6206_n1), .Q(WX4665) );
  INVX0 U6206_U1 ( .INP(n9597), .ZN(U6206_n1) );
  AND2X1 U6207_U2 ( .IN1(WX4600), .IN2(U6207_n1), .Q(WX4663) );
  INVX0 U6207_U1 ( .INP(n9597), .ZN(U6207_n1) );
  AND2X1 U6208_U2 ( .IN1(WX4598), .IN2(U6208_n1), .Q(WX4661) );
  INVX0 U6208_U1 ( .INP(n9597), .ZN(U6208_n1) );
  AND2X1 U6209_U2 ( .IN1(WX4596), .IN2(U6209_n1), .Q(WX4659) );
  INVX0 U6209_U1 ( .INP(n9597), .ZN(U6209_n1) );
  AND2X1 U6210_U2 ( .IN1(WX4594), .IN2(U6210_n1), .Q(WX4657) );
  INVX0 U6210_U1 ( .INP(n9597), .ZN(U6210_n1) );
  AND2X1 U6211_U2 ( .IN1(WX4592), .IN2(U6211_n1), .Q(WX4655) );
  INVX0 U6211_U1 ( .INP(n9597), .ZN(U6211_n1) );
  AND2X1 U6212_U2 ( .IN1(WX4590), .IN2(U6212_n1), .Q(WX4653) );
  INVX0 U6212_U1 ( .INP(n9597), .ZN(U6212_n1) );
  AND2X1 U6213_U2 ( .IN1(WX4588), .IN2(U6213_n1), .Q(WX4651) );
  INVX0 U6213_U1 ( .INP(n9597), .ZN(U6213_n1) );
  AND2X1 U6214_U2 ( .IN1(test_so36), .IN2(U6214_n1), .Q(WX4649) );
  INVX0 U6214_U1 ( .INP(n9596), .ZN(U6214_n1) );
  AND2X1 U6215_U2 ( .IN1(WX4584), .IN2(U6215_n1), .Q(WX4647) );
  INVX0 U6215_U1 ( .INP(n9596), .ZN(U6215_n1) );
  AND2X1 U6216_U2 ( .IN1(WX4582), .IN2(U6216_n1), .Q(WX4645) );
  INVX0 U6216_U1 ( .INP(n9596), .ZN(U6216_n1) );
  AND2X1 U6217_U2 ( .IN1(WX4580), .IN2(U6217_n1), .Q(WX4643) );
  INVX0 U6217_U1 ( .INP(n9596), .ZN(U6217_n1) );
  AND2X1 U6218_U2 ( .IN1(WX4578), .IN2(U6218_n1), .Q(WX4641) );
  INVX0 U6218_U1 ( .INP(n9596), .ZN(U6218_n1) );
  AND2X1 U6219_U2 ( .IN1(WX4576), .IN2(U6219_n1), .Q(WX4639) );
  INVX0 U6219_U1 ( .INP(n9596), .ZN(U6219_n1) );
  AND2X1 U6220_U2 ( .IN1(WX4574), .IN2(U6220_n1), .Q(WX4637) );
  INVX0 U6220_U1 ( .INP(n9596), .ZN(U6220_n1) );
  AND2X1 U6221_U2 ( .IN1(WX4572), .IN2(U6221_n1), .Q(WX4635) );
  INVX0 U6221_U1 ( .INP(n9596), .ZN(U6221_n1) );
  AND2X1 U6222_U2 ( .IN1(WX4570), .IN2(U6222_n1), .Q(WX4633) );
  INVX0 U6222_U1 ( .INP(n9596), .ZN(U6222_n1) );
  AND2X1 U6223_U2 ( .IN1(WX4568), .IN2(U6223_n1), .Q(WX4631) );
  INVX0 U6223_U1 ( .INP(n9596), .ZN(U6223_n1) );
  AND2X1 U6224_U2 ( .IN1(WX4566), .IN2(U6224_n1), .Q(WX4629) );
  INVX0 U6224_U1 ( .INP(n9596), .ZN(U6224_n1) );
  AND2X1 U6225_U2 ( .IN1(WX4564), .IN2(U6225_n1), .Q(WX4627) );
  INVX0 U6225_U1 ( .INP(n9596), .ZN(U6225_n1) );
  AND2X1 U6226_U2 ( .IN1(WX4562), .IN2(U6226_n1), .Q(WX4625) );
  INVX0 U6226_U1 ( .INP(n9596), .ZN(U6226_n1) );
  AND2X1 U6227_U2 ( .IN1(WX4560), .IN2(U6227_n1), .Q(WX4623) );
  INVX0 U6227_U1 ( .INP(n9596), .ZN(U6227_n1) );
  AND2X1 U6228_U2 ( .IN1(WX4558), .IN2(U6228_n1), .Q(WX4621) );
  INVX0 U6228_U1 ( .INP(n9595), .ZN(U6228_n1) );
  AND2X1 U6229_U2 ( .IN1(WX4556), .IN2(U6229_n1), .Q(WX4619) );
  INVX0 U6229_U1 ( .INP(n9595), .ZN(U6229_n1) );
  AND2X1 U6230_U2 ( .IN1(WX3421), .IN2(U6230_n1), .Q(WX3484) );
  INVX0 U6230_U1 ( .INP(n9595), .ZN(U6230_n1) );
  AND2X1 U6231_U2 ( .IN1(WX3419), .IN2(U6231_n1), .Q(WX3482) );
  INVX0 U6231_U1 ( .INP(n9595), .ZN(U6231_n1) );
  AND2X1 U6232_U2 ( .IN1(WX3417), .IN2(U6232_n1), .Q(WX3480) );
  INVX0 U6232_U1 ( .INP(n9595), .ZN(U6232_n1) );
  AND2X1 U6233_U2 ( .IN1(WX3415), .IN2(U6233_n1), .Q(WX3478) );
  INVX0 U6233_U1 ( .INP(n9595), .ZN(U6233_n1) );
  AND2X1 U6234_U2 ( .IN1(WX3413), .IN2(U6234_n1), .Q(WX3476) );
  INVX0 U6234_U1 ( .INP(n9595), .ZN(U6234_n1) );
  AND2X1 U6235_U2 ( .IN1(WX3411), .IN2(U6235_n1), .Q(WX3474) );
  INVX0 U6235_U1 ( .INP(n9595), .ZN(U6235_n1) );
  AND2X1 U6236_U2 ( .IN1(WX3409), .IN2(U6236_n1), .Q(WX3472) );
  INVX0 U6236_U1 ( .INP(n9595), .ZN(U6236_n1) );
  AND2X1 U6237_U2 ( .IN1(WX3407), .IN2(U6237_n1), .Q(WX3470) );
  INVX0 U6237_U1 ( .INP(n9595), .ZN(U6237_n1) );
  AND2X1 U6238_U2 ( .IN1(test_so28), .IN2(U6238_n1), .Q(WX3468) );
  INVX0 U6238_U1 ( .INP(n9595), .ZN(U6238_n1) );
  AND2X1 U6239_U2 ( .IN1(WX3403), .IN2(U6239_n1), .Q(WX3466) );
  INVX0 U6239_U1 ( .INP(n9595), .ZN(U6239_n1) );
  AND2X1 U6240_U2 ( .IN1(WX3401), .IN2(U6240_n1), .Q(WX3464) );
  INVX0 U6240_U1 ( .INP(n9595), .ZN(U6240_n1) );
  AND2X1 U6241_U2 ( .IN1(WX3399), .IN2(U6241_n1), .Q(WX3462) );
  INVX0 U6241_U1 ( .INP(n9595), .ZN(U6241_n1) );
  AND2X1 U6242_U2 ( .IN1(WX3397), .IN2(U6242_n1), .Q(WX3460) );
  INVX0 U6242_U1 ( .INP(n9594), .ZN(U6242_n1) );
  AND2X1 U6243_U2 ( .IN1(WX3395), .IN2(U6243_n1), .Q(WX3458) );
  INVX0 U6243_U1 ( .INP(n9594), .ZN(U6243_n1) );
  AND2X1 U6244_U2 ( .IN1(WX3393), .IN2(U6244_n1), .Q(WX3456) );
  INVX0 U6244_U1 ( .INP(n9594), .ZN(U6244_n1) );
  AND2X1 U6245_U2 ( .IN1(WX3391), .IN2(U6245_n1), .Q(WX3454) );
  INVX0 U6245_U1 ( .INP(n9594), .ZN(U6245_n1) );
  AND2X1 U6246_U2 ( .IN1(WX3389), .IN2(U6246_n1), .Q(WX3452) );
  INVX0 U6246_U1 ( .INP(n9594), .ZN(U6246_n1) );
  AND2X1 U6247_U2 ( .IN1(WX3387), .IN2(U6247_n1), .Q(WX3450) );
  INVX0 U6247_U1 ( .INP(n9594), .ZN(U6247_n1) );
  AND2X1 U6248_U2 ( .IN1(WX3385), .IN2(U6248_n1), .Q(WX3448) );
  INVX0 U6248_U1 ( .INP(n9594), .ZN(U6248_n1) );
  AND2X1 U6249_U2 ( .IN1(WX3383), .IN2(U6249_n1), .Q(WX3446) );
  INVX0 U6249_U1 ( .INP(n9594), .ZN(U6249_n1) );
  AND2X1 U6250_U2 ( .IN1(WX3381), .IN2(U6250_n1), .Q(WX3444) );
  INVX0 U6250_U1 ( .INP(n9594), .ZN(U6250_n1) );
  AND2X1 U6251_U2 ( .IN1(WX3379), .IN2(U6251_n1), .Q(WX3442) );
  INVX0 U6251_U1 ( .INP(n9594), .ZN(U6251_n1) );
  AND2X1 U6252_U2 ( .IN1(WX3377), .IN2(U6252_n1), .Q(WX3440) );
  INVX0 U6252_U1 ( .INP(n9594), .ZN(U6252_n1) );
  AND2X1 U6253_U2 ( .IN1(WX3375), .IN2(U6253_n1), .Q(WX3438) );
  INVX0 U6253_U1 ( .INP(n9594), .ZN(U6253_n1) );
  AND2X1 U6254_U2 ( .IN1(WX3373), .IN2(U6254_n1), .Q(WX3436) );
  INVX0 U6254_U1 ( .INP(n9594), .ZN(U6254_n1) );
  AND2X1 U6255_U2 ( .IN1(WX3371), .IN2(U6255_n1), .Q(WX3434) );
  INVX0 U6255_U1 ( .INP(n9594), .ZN(U6255_n1) );
  AND2X1 U6256_U2 ( .IN1(test_so27), .IN2(U6256_n1), .Q(WX3432) );
  INVX0 U6256_U1 ( .INP(n9593), .ZN(U6256_n1) );
  AND2X1 U6257_U2 ( .IN1(WX3367), .IN2(U6257_n1), .Q(WX3430) );
  INVX0 U6257_U1 ( .INP(n9593), .ZN(U6257_n1) );
  AND2X1 U6258_U2 ( .IN1(WX3365), .IN2(U6258_n1), .Q(WX3428) );
  INVX0 U6258_U1 ( .INP(n9593), .ZN(U6258_n1) );
  AND2X1 U6259_U2 ( .IN1(WX3363), .IN2(U6259_n1), .Q(WX3426) );
  INVX0 U6259_U1 ( .INP(n9593), .ZN(U6259_n1) );
  AND2X1 U6260_U2 ( .IN1(WX3361), .IN2(U6260_n1), .Q(WX3424) );
  INVX0 U6260_U1 ( .INP(n9593), .ZN(U6260_n1) );
  AND2X1 U6261_U2 ( .IN1(WX3359), .IN2(U6261_n1), .Q(WX3422) );
  INVX0 U6261_U1 ( .INP(n9593), .ZN(U6261_n1) );
  AND2X1 U6262_U2 ( .IN1(WX3357), .IN2(U6262_n1), .Q(WX3420) );
  INVX0 U6262_U1 ( .INP(n9593), .ZN(U6262_n1) );
  AND2X1 U6263_U2 ( .IN1(WX3355), .IN2(U6263_n1), .Q(WX3418) );
  INVX0 U6263_U1 ( .INP(n9593), .ZN(U6263_n1) );
  AND2X1 U6264_U2 ( .IN1(WX3353), .IN2(U6264_n1), .Q(WX3416) );
  INVX0 U6264_U1 ( .INP(n9593), .ZN(U6264_n1) );
  AND2X1 U6265_U2 ( .IN1(WX3351), .IN2(U6265_n1), .Q(WX3414) );
  INVX0 U6265_U1 ( .INP(n9593), .ZN(U6265_n1) );
  AND2X1 U6266_U2 ( .IN1(WX3349), .IN2(U6266_n1), .Q(WX3412) );
  INVX0 U6266_U1 ( .INP(n9593), .ZN(U6266_n1) );
  AND2X1 U6267_U2 ( .IN1(WX3347), .IN2(U6267_n1), .Q(WX3410) );
  INVX0 U6267_U1 ( .INP(n9593), .ZN(U6267_n1) );
  AND2X1 U6268_U2 ( .IN1(WX3345), .IN2(U6268_n1), .Q(WX3408) );
  INVX0 U6268_U1 ( .INP(n9593), .ZN(U6268_n1) );
  AND2X1 U6269_U2 ( .IN1(WX3343), .IN2(U6269_n1), .Q(WX3406) );
  INVX0 U6269_U1 ( .INP(n9593), .ZN(U6269_n1) );
  AND2X1 U6270_U2 ( .IN1(WX3341), .IN2(U6270_n1), .Q(WX3404) );
  INVX0 U6270_U1 ( .INP(n9592), .ZN(U6270_n1) );
  AND2X1 U6271_U2 ( .IN1(WX3339), .IN2(U6271_n1), .Q(WX3402) );
  INVX0 U6271_U1 ( .INP(n9592), .ZN(U6271_n1) );
  AND2X1 U6272_U2 ( .IN1(WX3337), .IN2(U6272_n1), .Q(WX3400) );
  INVX0 U6272_U1 ( .INP(n9592), .ZN(U6272_n1) );
  AND2X1 U6273_U2 ( .IN1(WX3335), .IN2(U6273_n1), .Q(WX3398) );
  INVX0 U6273_U1 ( .INP(n9592), .ZN(U6273_n1) );
  AND2X1 U6274_U2 ( .IN1(test_so26), .IN2(U6274_n1), .Q(WX3396) );
  INVX0 U6274_U1 ( .INP(n9592), .ZN(U6274_n1) );
  AND2X1 U6275_U2 ( .IN1(WX3331), .IN2(U6275_n1), .Q(WX3394) );
  INVX0 U6275_U1 ( .INP(n9592), .ZN(U6275_n1) );
  AND2X1 U6276_U2 ( .IN1(WX3329), .IN2(U6276_n1), .Q(WX3392) );
  INVX0 U6276_U1 ( .INP(n9592), .ZN(U6276_n1) );
  AND2X1 U6277_U2 ( .IN1(WX3327), .IN2(U6277_n1), .Q(WX3390) );
  INVX0 U6277_U1 ( .INP(n9592), .ZN(U6277_n1) );
  AND2X1 U6278_U2 ( .IN1(WX3325), .IN2(U6278_n1), .Q(WX3388) );
  INVX0 U6278_U1 ( .INP(n9592), .ZN(U6278_n1) );
  AND2X1 U6279_U2 ( .IN1(WX3323), .IN2(U6279_n1), .Q(WX3386) );
  INVX0 U6279_U1 ( .INP(n9592), .ZN(U6279_n1) );
  AND2X1 U6280_U2 ( .IN1(WX3321), .IN2(U6280_n1), .Q(WX3384) );
  INVX0 U6280_U1 ( .INP(n9592), .ZN(U6280_n1) );
  AND2X1 U6281_U2 ( .IN1(WX3319), .IN2(U6281_n1), .Q(WX3382) );
  INVX0 U6281_U1 ( .INP(n9592), .ZN(U6281_n1) );
  AND2X1 U6282_U2 ( .IN1(WX3317), .IN2(U6282_n1), .Q(WX3380) );
  INVX0 U6282_U1 ( .INP(n9592), .ZN(U6282_n1) );
  AND2X1 U6283_U2 ( .IN1(WX3315), .IN2(U6283_n1), .Q(WX3378) );
  INVX0 U6283_U1 ( .INP(n9592), .ZN(U6283_n1) );
  AND2X1 U6284_U2 ( .IN1(WX3313), .IN2(U6284_n1), .Q(WX3376) );
  INVX0 U6284_U1 ( .INP(n9591), .ZN(U6284_n1) );
  AND2X1 U6285_U2 ( .IN1(WX3311), .IN2(U6285_n1), .Q(WX3374) );
  INVX0 U6285_U1 ( .INP(n9591), .ZN(U6285_n1) );
  AND2X1 U6286_U2 ( .IN1(WX3309), .IN2(U6286_n1), .Q(WX3372) );
  INVX0 U6286_U1 ( .INP(n9591), .ZN(U6286_n1) );
  AND2X1 U6287_U2 ( .IN1(WX3307), .IN2(U6287_n1), .Q(WX3370) );
  INVX0 U6287_U1 ( .INP(n9591), .ZN(U6287_n1) );
  AND2X1 U6288_U2 ( .IN1(WX3305), .IN2(U6288_n1), .Q(WX3368) );
  INVX0 U6288_U1 ( .INP(n9591), .ZN(U6288_n1) );
  AND2X1 U6289_U2 ( .IN1(WX3303), .IN2(U6289_n1), .Q(WX3366) );
  INVX0 U6289_U1 ( .INP(n9591), .ZN(U6289_n1) );
  AND2X1 U6290_U2 ( .IN1(WX3301), .IN2(U6290_n1), .Q(WX3364) );
  INVX0 U6290_U1 ( .INP(n9591), .ZN(U6290_n1) );
  AND2X1 U6291_U2 ( .IN1(WX3299), .IN2(U6291_n1), .Q(WX3362) );
  INVX0 U6291_U1 ( .INP(n9591), .ZN(U6291_n1) );
  AND2X1 U6292_U2 ( .IN1(test_so25), .IN2(U6292_n1), .Q(WX3360) );
  INVX0 U6292_U1 ( .INP(n9591), .ZN(U6292_n1) );
  AND2X1 U6293_U2 ( .IN1(WX3295), .IN2(U6293_n1), .Q(WX3358) );
  INVX0 U6293_U1 ( .INP(n9591), .ZN(U6293_n1) );
  AND2X1 U6294_U2 ( .IN1(WX3293), .IN2(U6294_n1), .Q(WX3356) );
  INVX0 U6294_U1 ( .INP(n9591), .ZN(U6294_n1) );
  AND2X1 U6295_U2 ( .IN1(WX3291), .IN2(U6295_n1), .Q(WX3354) );
  INVX0 U6295_U1 ( .INP(n9591), .ZN(U6295_n1) );
  AND2X1 U6296_U2 ( .IN1(WX3289), .IN2(U6296_n1), .Q(WX3352) );
  INVX0 U6296_U1 ( .INP(n9591), .ZN(U6296_n1) );
  AND2X1 U6297_U2 ( .IN1(WX3287), .IN2(U6297_n1), .Q(WX3350) );
  INVX0 U6297_U1 ( .INP(n9591), .ZN(U6297_n1) );
  AND2X1 U6298_U2 ( .IN1(WX3285), .IN2(U6298_n1), .Q(WX3348) );
  INVX0 U6298_U1 ( .INP(n9590), .ZN(U6298_n1) );
  AND2X1 U6299_U2 ( .IN1(WX3283), .IN2(U6299_n1), .Q(WX3346) );
  INVX0 U6299_U1 ( .INP(n9590), .ZN(U6299_n1) );
  AND2X1 U6300_U2 ( .IN1(WX3281), .IN2(U6300_n1), .Q(WX3344) );
  INVX0 U6300_U1 ( .INP(n9590), .ZN(U6300_n1) );
  AND2X1 U6301_U2 ( .IN1(WX3279), .IN2(U6301_n1), .Q(WX3342) );
  INVX0 U6301_U1 ( .INP(n9590), .ZN(U6301_n1) );
  AND2X1 U6302_U2 ( .IN1(WX3277), .IN2(U6302_n1), .Q(WX3340) );
  INVX0 U6302_U1 ( .INP(n9590), .ZN(U6302_n1) );
  AND2X1 U6303_U2 ( .IN1(WX3275), .IN2(U6303_n1), .Q(WX3338) );
  INVX0 U6303_U1 ( .INP(n9590), .ZN(U6303_n1) );
  AND2X1 U6304_U2 ( .IN1(WX3273), .IN2(U6304_n1), .Q(WX3336) );
  INVX0 U6304_U1 ( .INP(n9590), .ZN(U6304_n1) );
  AND2X1 U6305_U2 ( .IN1(WX3271), .IN2(U6305_n1), .Q(WX3334) );
  INVX0 U6305_U1 ( .INP(n9590), .ZN(U6305_n1) );
  AND2X1 U6306_U2 ( .IN1(WX3267), .IN2(U6306_n1), .Q(WX3330) );
  INVX0 U6306_U1 ( .INP(n9590), .ZN(U6306_n1) );
  AND2X1 U6307_U2 ( .IN1(WX2128), .IN2(U6307_n1), .Q(WX2191) );
  INVX0 U6307_U1 ( .INP(n9590), .ZN(U6307_n1) );
  AND2X1 U6308_U2 ( .IN1(WX2126), .IN2(U6308_n1), .Q(WX2189) );
  INVX0 U6308_U1 ( .INP(n9590), .ZN(U6308_n1) );
  AND2X1 U6309_U2 ( .IN1(WX2124), .IN2(U6309_n1), .Q(WX2187) );
  INVX0 U6309_U1 ( .INP(n9590), .ZN(U6309_n1) );
  AND2X1 U6310_U2 ( .IN1(WX2122), .IN2(U6310_n1), .Q(WX2185) );
  INVX0 U6310_U1 ( .INP(n9590), .ZN(U6310_n1) );
  AND2X1 U6311_U2 ( .IN1(WX2120), .IN2(U6311_n1), .Q(WX2183) );
  INVX0 U6311_U1 ( .INP(n9590), .ZN(U6311_n1) );
  AND2X1 U6312_U2 ( .IN1(WX2118), .IN2(U6312_n1), .Q(WX2181) );
  INVX0 U6312_U1 ( .INP(n9589), .ZN(U6312_n1) );
  AND2X1 U6313_U2 ( .IN1(WX2116), .IN2(U6313_n1), .Q(WX2179) );
  INVX0 U6313_U1 ( .INP(n9589), .ZN(U6313_n1) );
  AND2X1 U6314_U2 ( .IN1(WX2114), .IN2(U6314_n1), .Q(WX2177) );
  INVX0 U6314_U1 ( .INP(n9589), .ZN(U6314_n1) );
  AND2X1 U6315_U2 ( .IN1(WX2112), .IN2(U6315_n1), .Q(WX2175) );
  INVX0 U6315_U1 ( .INP(n9589), .ZN(U6315_n1) );
  AND2X1 U6316_U2 ( .IN1(WX2110), .IN2(U6316_n1), .Q(WX2173) );
  INVX0 U6316_U1 ( .INP(n9589), .ZN(U6316_n1) );
  AND2X1 U6317_U2 ( .IN1(WX2108), .IN2(U6317_n1), .Q(WX2171) );
  INVX0 U6317_U1 ( .INP(n9589), .ZN(U6317_n1) );
  AND2X1 U6318_U2 ( .IN1(WX2106), .IN2(U6318_n1), .Q(WX2169) );
  INVX0 U6318_U1 ( .INP(n9589), .ZN(U6318_n1) );
  AND2X1 U6319_U2 ( .IN1(WX2104), .IN2(U6319_n1), .Q(WX2167) );
  INVX0 U6319_U1 ( .INP(n9589), .ZN(U6319_n1) );
  AND2X1 U6320_U2 ( .IN1(WX2102), .IN2(U6320_n1), .Q(WX2165) );
  INVX0 U6320_U1 ( .INP(n9589), .ZN(U6320_n1) );
  AND2X1 U6321_U2 ( .IN1(test_so17), .IN2(U6321_n1), .Q(WX2163) );
  INVX0 U6321_U1 ( .INP(n9589), .ZN(U6321_n1) );
  AND2X1 U6322_U2 ( .IN1(WX2098), .IN2(U6322_n1), .Q(WX2161) );
  INVX0 U6322_U1 ( .INP(n9589), .ZN(U6322_n1) );
  AND2X1 U6323_U2 ( .IN1(WX2096), .IN2(U6323_n1), .Q(WX2159) );
  INVX0 U6323_U1 ( .INP(n9589), .ZN(U6323_n1) );
  AND2X1 U6324_U2 ( .IN1(WX2094), .IN2(U6324_n1), .Q(WX2157) );
  INVX0 U6324_U1 ( .INP(n9589), .ZN(U6324_n1) );
  AND2X1 U6325_U2 ( .IN1(WX2092), .IN2(U6325_n1), .Q(WX2155) );
  INVX0 U6325_U1 ( .INP(n9589), .ZN(U6325_n1) );
  AND2X1 U6326_U2 ( .IN1(WX2090), .IN2(U6326_n1), .Q(WX2153) );
  INVX0 U6326_U1 ( .INP(n9588), .ZN(U6326_n1) );
  AND2X1 U6327_U2 ( .IN1(WX2088), .IN2(U6327_n1), .Q(WX2151) );
  INVX0 U6327_U1 ( .INP(n9588), .ZN(U6327_n1) );
  AND2X1 U6328_U2 ( .IN1(WX2086), .IN2(U6328_n1), .Q(WX2149) );
  INVX0 U6328_U1 ( .INP(n9588), .ZN(U6328_n1) );
  AND2X1 U6329_U2 ( .IN1(WX2084), .IN2(U6329_n1), .Q(WX2147) );
  INVX0 U6329_U1 ( .INP(n9588), .ZN(U6329_n1) );
  AND2X1 U6330_U2 ( .IN1(WX2082), .IN2(U6330_n1), .Q(WX2145) );
  INVX0 U6330_U1 ( .INP(n9588), .ZN(U6330_n1) );
  AND2X1 U6331_U2 ( .IN1(WX2080), .IN2(U6331_n1), .Q(WX2143) );
  INVX0 U6331_U1 ( .INP(n9588), .ZN(U6331_n1) );
  AND2X1 U6332_U2 ( .IN1(WX2078), .IN2(U6332_n1), .Q(WX2141) );
  INVX0 U6332_U1 ( .INP(n9588), .ZN(U6332_n1) );
  AND2X1 U6333_U2 ( .IN1(WX2076), .IN2(U6333_n1), .Q(WX2139) );
  INVX0 U6333_U1 ( .INP(n9588), .ZN(U6333_n1) );
  AND2X1 U6334_U2 ( .IN1(WX2074), .IN2(U6334_n1), .Q(WX2137) );
  INVX0 U6334_U1 ( .INP(n9588), .ZN(U6334_n1) );
  AND2X1 U6335_U2 ( .IN1(WX2072), .IN2(U6335_n1), .Q(WX2135) );
  INVX0 U6335_U1 ( .INP(n9588), .ZN(U6335_n1) );
  AND2X1 U6336_U2 ( .IN1(WX2070), .IN2(U6336_n1), .Q(WX2133) );
  INVX0 U6336_U1 ( .INP(n9588), .ZN(U6336_n1) );
  AND2X1 U6337_U2 ( .IN1(WX2068), .IN2(U6337_n1), .Q(WX2131) );
  INVX0 U6337_U1 ( .INP(n9588), .ZN(U6337_n1) );
  AND2X1 U6338_U2 ( .IN1(WX2066), .IN2(U6338_n1), .Q(WX2129) );
  INVX0 U6338_U1 ( .INP(n9588), .ZN(U6338_n1) );
  AND2X1 U6339_U2 ( .IN1(test_so16), .IN2(U6339_n1), .Q(WX2127) );
  INVX0 U6339_U1 ( .INP(n9588), .ZN(U6339_n1) );
  AND2X1 U6340_U2 ( .IN1(WX2062), .IN2(U6340_n1), .Q(WX2125) );
  INVX0 U6340_U1 ( .INP(n9587), .ZN(U6340_n1) );
  AND2X1 U6341_U2 ( .IN1(WX2060), .IN2(U6341_n1), .Q(WX2123) );
  INVX0 U6341_U1 ( .INP(n9587), .ZN(U6341_n1) );
  AND2X1 U6342_U2 ( .IN1(WX2058), .IN2(U6342_n1), .Q(WX2121) );
  INVX0 U6342_U1 ( .INP(n9587), .ZN(U6342_n1) );
  AND2X1 U6343_U2 ( .IN1(WX2056), .IN2(U6343_n1), .Q(WX2119) );
  INVX0 U6343_U1 ( .INP(n9587), .ZN(U6343_n1) );
  AND2X1 U6344_U2 ( .IN1(WX2054), .IN2(U6344_n1), .Q(WX2117) );
  INVX0 U6344_U1 ( .INP(n9587), .ZN(U6344_n1) );
  AND2X1 U6345_U2 ( .IN1(WX2052), .IN2(U6345_n1), .Q(WX2115) );
  INVX0 U6345_U1 ( .INP(n9587), .ZN(U6345_n1) );
  AND2X1 U6346_U2 ( .IN1(WX2050), .IN2(U6346_n1), .Q(WX2113) );
  INVX0 U6346_U1 ( .INP(n9587), .ZN(U6346_n1) );
  AND2X1 U6347_U2 ( .IN1(WX2048), .IN2(U6347_n1), .Q(WX2111) );
  INVX0 U6347_U1 ( .INP(n9587), .ZN(U6347_n1) );
  AND2X1 U6348_U2 ( .IN1(WX2046), .IN2(U6348_n1), .Q(WX2109) );
  INVX0 U6348_U1 ( .INP(n9587), .ZN(U6348_n1) );
  AND2X1 U6349_U2 ( .IN1(WX2044), .IN2(U6349_n1), .Q(WX2107) );
  INVX0 U6349_U1 ( .INP(n9587), .ZN(U6349_n1) );
  AND2X1 U6350_U2 ( .IN1(WX2042), .IN2(U6350_n1), .Q(WX2105) );
  INVX0 U6350_U1 ( .INP(n9587), .ZN(U6350_n1) );
  AND2X1 U6351_U2 ( .IN1(WX2040), .IN2(U6351_n1), .Q(WX2103) );
  INVX0 U6351_U1 ( .INP(n9587), .ZN(U6351_n1) );
  AND2X1 U6352_U2 ( .IN1(WX2038), .IN2(U6352_n1), .Q(WX2101) );
  INVX0 U6352_U1 ( .INP(n9587), .ZN(U6352_n1) );
  AND2X1 U6353_U2 ( .IN1(WX2036), .IN2(U6353_n1), .Q(WX2099) );
  INVX0 U6353_U1 ( .INP(n9587), .ZN(U6353_n1) );
  AND2X1 U6354_U2 ( .IN1(WX2034), .IN2(U6354_n1), .Q(WX2097) );
  INVX0 U6354_U1 ( .INP(n9586), .ZN(U6354_n1) );
  AND2X1 U6355_U2 ( .IN1(WX2032), .IN2(U6355_n1), .Q(WX2095) );
  INVX0 U6355_U1 ( .INP(n9586), .ZN(U6355_n1) );
  AND2X1 U6356_U2 ( .IN1(WX2030), .IN2(U6356_n1), .Q(WX2093) );
  INVX0 U6356_U1 ( .INP(n9586), .ZN(U6356_n1) );
  AND2X1 U6357_U2 ( .IN1(test_so15), .IN2(U6357_n1), .Q(WX2091) );
  INVX0 U6357_U1 ( .INP(n9586), .ZN(U6357_n1) );
  AND2X1 U6358_U2 ( .IN1(WX2026), .IN2(U6358_n1), .Q(WX2089) );
  INVX0 U6358_U1 ( .INP(n9586), .ZN(U6358_n1) );
  AND2X1 U6359_U2 ( .IN1(WX2024), .IN2(U6359_n1), .Q(WX2087) );
  INVX0 U6359_U1 ( .INP(n9586), .ZN(U6359_n1) );
  AND2X1 U6360_U2 ( .IN1(WX2022), .IN2(U6360_n1), .Q(WX2085) );
  INVX0 U6360_U1 ( .INP(n9586), .ZN(U6360_n1) );
  AND2X1 U6361_U2 ( .IN1(WX2020), .IN2(U6361_n1), .Q(WX2083) );
  INVX0 U6361_U1 ( .INP(n9586), .ZN(U6361_n1) );
  AND2X1 U6362_U2 ( .IN1(WX2018), .IN2(U6362_n1), .Q(WX2081) );
  INVX0 U6362_U1 ( .INP(n9586), .ZN(U6362_n1) );
  AND2X1 U6363_U2 ( .IN1(WX2016), .IN2(U6363_n1), .Q(WX2079) );
  INVX0 U6363_U1 ( .INP(n9586), .ZN(U6363_n1) );
  AND2X1 U6364_U2 ( .IN1(WX2014), .IN2(U6364_n1), .Q(WX2077) );
  INVX0 U6364_U1 ( .INP(n9586), .ZN(U6364_n1) );
  AND2X1 U6365_U2 ( .IN1(WX2012), .IN2(U6365_n1), .Q(WX2075) );
  INVX0 U6365_U1 ( .INP(n9586), .ZN(U6365_n1) );
  AND2X1 U6366_U2 ( .IN1(WX2010), .IN2(U6366_n1), .Q(WX2073) );
  INVX0 U6366_U1 ( .INP(n9586), .ZN(U6366_n1) );
  AND2X1 U6367_U2 ( .IN1(WX2008), .IN2(U6367_n1), .Q(WX2071) );
  INVX0 U6367_U1 ( .INP(n9586), .ZN(U6367_n1) );
  AND2X1 U6368_U2 ( .IN1(WX2006), .IN2(U6368_n1), .Q(WX2069) );
  INVX0 U6368_U1 ( .INP(n9585), .ZN(U6368_n1) );
  AND2X1 U6369_U2 ( .IN1(WX2004), .IN2(U6369_n1), .Q(WX2067) );
  INVX0 U6369_U1 ( .INP(n9585), .ZN(U6369_n1) );
  AND2X1 U6370_U2 ( .IN1(WX2002), .IN2(U6370_n1), .Q(WX2065) );
  INVX0 U6370_U1 ( .INP(n9585), .ZN(U6370_n1) );
  AND2X1 U6371_U2 ( .IN1(WX2000), .IN2(U6371_n1), .Q(WX2063) );
  INVX0 U6371_U1 ( .INP(n9585), .ZN(U6371_n1) );
  AND2X1 U6372_U2 ( .IN1(WX1998), .IN2(U6372_n1), .Q(WX2061) );
  INVX0 U6372_U1 ( .INP(n9585), .ZN(U6372_n1) );
  AND2X1 U6373_U2 ( .IN1(WX1996), .IN2(U6373_n1), .Q(WX2059) );
  INVX0 U6373_U1 ( .INP(n9585), .ZN(U6373_n1) );
  AND2X1 U6374_U2 ( .IN1(WX1994), .IN2(U6374_n1), .Q(WX2057) );
  INVX0 U6374_U1 ( .INP(n9585), .ZN(U6374_n1) );
  AND2X1 U6375_U2 ( .IN1(test_so14), .IN2(U6375_n1), .Q(WX2055) );
  INVX0 U6375_U1 ( .INP(n9585), .ZN(U6375_n1) );
  AND2X1 U6376_U2 ( .IN1(WX1990), .IN2(U6376_n1), .Q(WX2053) );
  INVX0 U6376_U1 ( .INP(n9585), .ZN(U6376_n1) );
  AND2X1 U6377_U2 ( .IN1(WX1988), .IN2(U6377_n1), .Q(WX2051) );
  INVX0 U6377_U1 ( .INP(n9585), .ZN(U6377_n1) );
  AND2X1 U6378_U2 ( .IN1(WX1986), .IN2(U6378_n1), .Q(WX2049) );
  INVX0 U6378_U1 ( .INP(n9585), .ZN(U6378_n1) );
  AND2X1 U6379_U2 ( .IN1(WX1984), .IN2(U6379_n1), .Q(WX2047) );
  INVX0 U6379_U1 ( .INP(n9585), .ZN(U6379_n1) );
  AND2X1 U6380_U2 ( .IN1(WX1982), .IN2(U6380_n1), .Q(WX2045) );
  INVX0 U6380_U1 ( .INP(n9585), .ZN(U6380_n1) );
  AND2X1 U6381_U2 ( .IN1(WX1980), .IN2(U6381_n1), .Q(WX2043) );
  INVX0 U6381_U1 ( .INP(n9585), .ZN(U6381_n1) );
  AND2X1 U6382_U2 ( .IN1(WX1978), .IN2(U6382_n1), .Q(WX2041) );
  INVX0 U6382_U1 ( .INP(n9584), .ZN(U6382_n1) );
  AND2X1 U6383_U2 ( .IN1(WX1976), .IN2(U6383_n1), .Q(WX2039) );
  INVX0 U6383_U1 ( .INP(n9584), .ZN(U6383_n1) );
  AND2X1 U6384_U2 ( .IN1(WX1974), .IN2(U6384_n1), .Q(WX2037) );
  INVX0 U6384_U1 ( .INP(n9584), .ZN(U6384_n1) );
  AND2X1 U6385_U2 ( .IN1(WX1972), .IN2(U6385_n1), .Q(WX2035) );
  INVX0 U6385_U1 ( .INP(n9584), .ZN(U6385_n1) );
  AND2X1 U6386_U2 ( .IN1(WX1970), .IN2(U6386_n1), .Q(WX2033) );
  INVX0 U6386_U1 ( .INP(n9584), .ZN(U6386_n1) );
  AND2X1 U6387_U2 ( .IN1(WX835), .IN2(U6387_n1), .Q(WX898) );
  INVX0 U6387_U1 ( .INP(n9584), .ZN(U6387_n1) );
  AND2X1 U6388_U2 ( .IN1(WX833), .IN2(U6388_n1), .Q(WX896) );
  INVX0 U6388_U1 ( .INP(n9584), .ZN(U6388_n1) );
  AND2X1 U6389_U2 ( .IN1(test_so7), .IN2(U6389_n1), .Q(WX894) );
  INVX0 U6389_U1 ( .INP(n9584), .ZN(U6389_n1) );
  AND2X1 U6390_U2 ( .IN1(WX829), .IN2(U6390_n1), .Q(WX892) );
  INVX0 U6390_U1 ( .INP(n9584), .ZN(U6390_n1) );
  AND2X1 U6391_U2 ( .IN1(WX827), .IN2(U6391_n1), .Q(WX890) );
  INVX0 U6391_U1 ( .INP(n9584), .ZN(U6391_n1) );
  AND2X1 U6392_U2 ( .IN1(WX825), .IN2(U6392_n1), .Q(WX888) );
  INVX0 U6392_U1 ( .INP(n9584), .ZN(U6392_n1) );
  AND2X1 U6393_U2 ( .IN1(WX823), .IN2(U6393_n1), .Q(WX886) );
  INVX0 U6393_U1 ( .INP(n9584), .ZN(U6393_n1) );
  AND2X1 U6394_U2 ( .IN1(WX821), .IN2(U6394_n1), .Q(WX884) );
  INVX0 U6394_U1 ( .INP(n9584), .ZN(U6394_n1) );
  AND2X1 U6395_U2 ( .IN1(WX819), .IN2(U6395_n1), .Q(WX882) );
  INVX0 U6395_U1 ( .INP(n9584), .ZN(U6395_n1) );
  AND2X1 U6396_U2 ( .IN1(WX817), .IN2(U6396_n1), .Q(WX880) );
  INVX0 U6396_U1 ( .INP(n9583), .ZN(U6396_n1) );
  AND2X1 U6397_U2 ( .IN1(WX815), .IN2(U6397_n1), .Q(WX878) );
  INVX0 U6397_U1 ( .INP(n9583), .ZN(U6397_n1) );
  AND2X1 U6398_U2 ( .IN1(WX813), .IN2(U6398_n1), .Q(WX876) );
  INVX0 U6398_U1 ( .INP(n9583), .ZN(U6398_n1) );
  AND2X1 U6399_U2 ( .IN1(WX811), .IN2(U6399_n1), .Q(WX874) );
  INVX0 U6399_U1 ( .INP(n9583), .ZN(U6399_n1) );
  AND2X1 U6400_U2 ( .IN1(WX809), .IN2(U6400_n1), .Q(WX872) );
  INVX0 U6400_U1 ( .INP(n9583), .ZN(U6400_n1) );
  AND2X1 U6401_U2 ( .IN1(WX807), .IN2(U6401_n1), .Q(WX870) );
  INVX0 U6401_U1 ( .INP(n9583), .ZN(U6401_n1) );
  AND2X1 U6402_U2 ( .IN1(WX805), .IN2(U6402_n1), .Q(WX868) );
  INVX0 U6402_U1 ( .INP(n9583), .ZN(U6402_n1) );
  AND2X1 U6403_U2 ( .IN1(WX803), .IN2(U6403_n1), .Q(WX866) );
  INVX0 U6403_U1 ( .INP(n9583), .ZN(U6403_n1) );
  AND2X1 U6404_U2 ( .IN1(WX801), .IN2(U6404_n1), .Q(WX864) );
  INVX0 U6404_U1 ( .INP(n9583), .ZN(U6404_n1) );
  AND2X1 U6405_U2 ( .IN1(WX799), .IN2(U6405_n1), .Q(WX862) );
  INVX0 U6405_U1 ( .INP(n9583), .ZN(U6405_n1) );
  AND2X1 U6406_U2 ( .IN1(WX797), .IN2(U6406_n1), .Q(WX860) );
  INVX0 U6406_U1 ( .INP(n9583), .ZN(U6406_n1) );
  AND2X1 U6407_U2 ( .IN1(test_so6), .IN2(U6407_n1), .Q(WX858) );
  INVX0 U6407_U1 ( .INP(n9583), .ZN(U6407_n1) );
  AND2X1 U6408_U2 ( .IN1(WX793), .IN2(U6408_n1), .Q(WX856) );
  INVX0 U6408_U1 ( .INP(n9583), .ZN(U6408_n1) );
  AND2X1 U6409_U2 ( .IN1(WX791), .IN2(U6409_n1), .Q(WX854) );
  INVX0 U6409_U1 ( .INP(n9583), .ZN(U6409_n1) );
  AND2X1 U6410_U2 ( .IN1(WX789), .IN2(U6410_n1), .Q(WX852) );
  INVX0 U6410_U1 ( .INP(n9582), .ZN(U6410_n1) );
  AND2X1 U6411_U2 ( .IN1(WX787), .IN2(U6411_n1), .Q(WX850) );
  INVX0 U6411_U1 ( .INP(n9582), .ZN(U6411_n1) );
  AND2X1 U6412_U2 ( .IN1(WX785), .IN2(U6412_n1), .Q(WX848) );
  INVX0 U6412_U1 ( .INP(n9582), .ZN(U6412_n1) );
  AND2X1 U6413_U2 ( .IN1(WX783), .IN2(U6413_n1), .Q(WX846) );
  INVX0 U6413_U1 ( .INP(n9582), .ZN(U6413_n1) );
  AND2X1 U6414_U2 ( .IN1(WX781), .IN2(U6414_n1), .Q(WX844) );
  INVX0 U6414_U1 ( .INP(n9582), .ZN(U6414_n1) );
  AND2X1 U6415_U2 ( .IN1(WX779), .IN2(U6415_n1), .Q(WX842) );
  INVX0 U6415_U1 ( .INP(n9582), .ZN(U6415_n1) );
  AND2X1 U6416_U2 ( .IN1(WX777), .IN2(U6416_n1), .Q(WX840) );
  INVX0 U6416_U1 ( .INP(n9582), .ZN(U6416_n1) );
  AND2X1 U6417_U2 ( .IN1(WX775), .IN2(U6417_n1), .Q(WX838) );
  INVX0 U6417_U1 ( .INP(n9582), .ZN(U6417_n1) );
  AND2X1 U6418_U2 ( .IN1(WX773), .IN2(U6418_n1), .Q(WX836) );
  INVX0 U6418_U1 ( .INP(n9582), .ZN(U6418_n1) );
  AND2X1 U6419_U2 ( .IN1(WX771), .IN2(U6419_n1), .Q(WX834) );
  INVX0 U6419_U1 ( .INP(n9582), .ZN(U6419_n1) );
  AND2X1 U6420_U2 ( .IN1(WX769), .IN2(U6420_n1), .Q(WX832) );
  INVX0 U6420_U1 ( .INP(n9582), .ZN(U6420_n1) );
  AND2X1 U6421_U2 ( .IN1(WX767), .IN2(U6421_n1), .Q(WX830) );
  INVX0 U6421_U1 ( .INP(n9582), .ZN(U6421_n1) );
  AND2X1 U6422_U2 ( .IN1(WX765), .IN2(U6422_n1), .Q(WX828) );
  INVX0 U6422_U1 ( .INP(n9582), .ZN(U6422_n1) );
  AND2X1 U6423_U2 ( .IN1(WX763), .IN2(U6423_n1), .Q(WX826) );
  INVX0 U6423_U1 ( .INP(n9582), .ZN(U6423_n1) );
  AND2X1 U6424_U2 ( .IN1(WX761), .IN2(U6424_n1), .Q(WX824) );
  INVX0 U6424_U1 ( .INP(n9581), .ZN(U6424_n1) );
  AND2X1 U6425_U2 ( .IN1(test_so5), .IN2(U6425_n1), .Q(WX822) );
  INVX0 U6425_U1 ( .INP(n9581), .ZN(U6425_n1) );
  AND2X1 U6426_U2 ( .IN1(WX757), .IN2(U6426_n1), .Q(WX820) );
  INVX0 U6426_U1 ( .INP(n9581), .ZN(U6426_n1) );
  AND2X1 U6427_U2 ( .IN1(WX755), .IN2(U6427_n1), .Q(WX818) );
  INVX0 U6427_U1 ( .INP(n9581), .ZN(U6427_n1) );
  AND2X1 U6428_U2 ( .IN1(WX753), .IN2(U6428_n1), .Q(WX816) );
  INVX0 U6428_U1 ( .INP(n9581), .ZN(U6428_n1) );
  AND2X1 U6429_U2 ( .IN1(WX751), .IN2(U6429_n1), .Q(WX814) );
  INVX0 U6429_U1 ( .INP(n9581), .ZN(U6429_n1) );
  AND2X1 U6430_U2 ( .IN1(WX749), .IN2(U6430_n1), .Q(WX812) );
  INVX0 U6430_U1 ( .INP(n9581), .ZN(U6430_n1) );
  AND2X1 U6431_U2 ( .IN1(WX747), .IN2(U6431_n1), .Q(WX810) );
  INVX0 U6431_U1 ( .INP(n9581), .ZN(U6431_n1) );
  AND2X1 U6432_U2 ( .IN1(WX745), .IN2(U6432_n1), .Q(WX808) );
  INVX0 U6432_U1 ( .INP(n9581), .ZN(U6432_n1) );
  AND2X1 U6433_U2 ( .IN1(WX743), .IN2(U6433_n1), .Q(WX806) );
  INVX0 U6433_U1 ( .INP(n9581), .ZN(U6433_n1) );
  AND2X1 U6434_U2 ( .IN1(WX741), .IN2(U6434_n1), .Q(WX804) );
  INVX0 U6434_U1 ( .INP(n9581), .ZN(U6434_n1) );
  AND2X1 U6435_U2 ( .IN1(WX739), .IN2(U6435_n1), .Q(WX802) );
  INVX0 U6435_U1 ( .INP(n9581), .ZN(U6435_n1) );
  AND2X1 U6436_U2 ( .IN1(WX737), .IN2(U6436_n1), .Q(WX800) );
  INVX0 U6436_U1 ( .INP(n9581), .ZN(U6436_n1) );
  AND2X1 U6437_U2 ( .IN1(WX735), .IN2(U6437_n1), .Q(WX798) );
  INVX0 U6437_U1 ( .INP(n9581), .ZN(U6437_n1) );
  AND2X1 U6438_U2 ( .IN1(WX733), .IN2(U6438_n1), .Q(WX796) );
  INVX0 U6438_U1 ( .INP(n9580), .ZN(U6438_n1) );
  AND2X1 U6439_U2 ( .IN1(WX731), .IN2(U6439_n1), .Q(WX794) );
  INVX0 U6439_U1 ( .INP(n9580), .ZN(U6439_n1) );
  AND2X1 U6440_U2 ( .IN1(WX729), .IN2(U6440_n1), .Q(WX792) );
  INVX0 U6440_U1 ( .INP(n9580), .ZN(U6440_n1) );
  AND2X1 U6441_U2 ( .IN1(WX727), .IN2(U6441_n1), .Q(WX790) );
  INVX0 U6441_U1 ( .INP(n9580), .ZN(U6441_n1) );
  AND2X1 U6442_U2 ( .IN1(WX725), .IN2(U6442_n1), .Q(WX788) );
  INVX0 U6442_U1 ( .INP(n9580), .ZN(U6442_n1) );
  AND2X1 U6443_U2 ( .IN1(test_so4), .IN2(U6443_n1), .Q(WX786) );
  INVX0 U6443_U1 ( .INP(n9580), .ZN(U6443_n1) );
  AND2X1 U6444_U2 ( .IN1(WX721), .IN2(U6444_n1), .Q(WX784) );
  INVX0 U6444_U1 ( .INP(n9580), .ZN(U6444_n1) );
  AND2X1 U6445_U2 ( .IN1(WX719), .IN2(U6445_n1), .Q(WX782) );
  INVX0 U6445_U1 ( .INP(n9580), .ZN(U6445_n1) );
  AND2X1 U6446_U2 ( .IN1(WX717), .IN2(U6446_n1), .Q(WX780) );
  INVX0 U6446_U1 ( .INP(n9580), .ZN(U6446_n1) );
  AND2X1 U6447_U2 ( .IN1(WX715), .IN2(U6447_n1), .Q(WX778) );
  INVX0 U6447_U1 ( .INP(n9580), .ZN(U6447_n1) );
  AND2X1 U6448_U2 ( .IN1(WX713), .IN2(U6448_n1), .Q(WX776) );
  INVX0 U6448_U1 ( .INP(n9580), .ZN(U6448_n1) );
  AND2X1 U6449_U2 ( .IN1(WX711), .IN2(U6449_n1), .Q(WX774) );
  INVX0 U6449_U1 ( .INP(n9580), .ZN(U6449_n1) );
  AND2X1 U6450_U2 ( .IN1(WX709), .IN2(U6450_n1), .Q(WX772) );
  INVX0 U6450_U1 ( .INP(n9580), .ZN(U6450_n1) );
  AND2X1 U6451_U2 ( .IN1(WX707), .IN2(U6451_n1), .Q(WX770) );
  INVX0 U6451_U1 ( .INP(n9580), .ZN(U6451_n1) );
  AND2X1 U6452_U2 ( .IN1(WX705), .IN2(U6452_n1), .Q(WX768) );
  INVX0 U6452_U1 ( .INP(n9579), .ZN(U6452_n1) );
  AND2X1 U6453_U2 ( .IN1(WX703), .IN2(U6453_n1), .Q(WX766) );
  INVX0 U6453_U1 ( .INP(n9579), .ZN(U6453_n1) );
  AND2X1 U6454_U2 ( .IN1(WX701), .IN2(U6454_n1), .Q(WX764) );
  INVX0 U6454_U1 ( .INP(n9579), .ZN(U6454_n1) );
  AND2X1 U6455_U2 ( .IN1(WX699), .IN2(U6455_n1), .Q(WX762) );
  INVX0 U6455_U1 ( .INP(n9579), .ZN(U6455_n1) );
  AND2X1 U6456_U2 ( .IN1(WX697), .IN2(U6456_n1), .Q(WX760) );
  INVX0 U6456_U1 ( .INP(n9579), .ZN(U6456_n1) );
  AND2X1 U6457_U2 ( .IN1(WX695), .IN2(U6457_n1), .Q(WX758) );
  INVX0 U6457_U1 ( .INP(n9579), .ZN(U6457_n1) );
  AND2X1 U6458_U2 ( .IN1(WX693), .IN2(U6458_n1), .Q(WX756) );
  INVX0 U6458_U1 ( .INP(n9579), .ZN(U6458_n1) );
  AND2X1 U6459_U2 ( .IN1(WX691), .IN2(U6459_n1), .Q(WX754) );
  INVX0 U6459_U1 ( .INP(n9579), .ZN(U6459_n1) );
  AND2X1 U6460_U2 ( .IN1(WX689), .IN2(U6460_n1), .Q(WX752) );
  INVX0 U6460_U1 ( .INP(n9579), .ZN(U6460_n1) );
  AND2X1 U6461_U2 ( .IN1(test_so3), .IN2(U6461_n1), .Q(WX750) );
  INVX0 U6461_U1 ( .INP(n9579), .ZN(U6461_n1) );
  AND2X1 U6462_U2 ( .IN1(WX685), .IN2(U6462_n1), .Q(WX748) );
  INVX0 U6462_U1 ( .INP(n9579), .ZN(U6462_n1) );
  AND2X1 U6463_U2 ( .IN1(WX683), .IN2(U6463_n1), .Q(WX746) );
  INVX0 U6463_U1 ( .INP(n9579), .ZN(U6463_n1) );
  AND2X1 U6464_U2 ( .IN1(WX681), .IN2(U6464_n1), .Q(WX744) );
  INVX0 U6464_U1 ( .INP(n9579), .ZN(U6464_n1) );
  AND2X1 U6465_U2 ( .IN1(WX679), .IN2(U6465_n1), .Q(WX742) );
  INVX0 U6465_U1 ( .INP(n9579), .ZN(U6465_n1) );
  AND2X1 U6466_U2 ( .IN1(WX677), .IN2(U6466_n1), .Q(WX740) );
  INVX0 U6466_U1 ( .INP(n9578), .ZN(U6466_n1) );
  AND2X1 U6467_U2 ( .IN1(WX675), .IN2(U6467_n1), .Q(WX738) );
  INVX0 U6467_U1 ( .INP(n9578), .ZN(U6467_n1) );
  AND2X1 U6468_U2 ( .IN1(WX673), .IN2(U6468_n1), .Q(WX736) );
  INVX0 U6468_U1 ( .INP(n9578), .ZN(U6468_n1) );
  AND2X1 U6469_U2 ( .IN1(WX671), .IN2(U6469_n1), .Q(WX734) );
  INVX0 U6469_U1 ( .INP(n9578), .ZN(U6469_n1) );
  AND2X1 U6470_U2 ( .IN1(WX669), .IN2(U6470_n1), .Q(WX732) );
  INVX0 U6470_U1 ( .INP(n9578), .ZN(U6470_n1) );
  AND2X1 U6471_U2 ( .IN1(WX667), .IN2(U6471_n1), .Q(WX730) );
  INVX0 U6471_U1 ( .INP(n9578), .ZN(U6471_n1) );
  AND2X1 U6472_U2 ( .IN1(WX665), .IN2(U6472_n1), .Q(WX728) );
  INVX0 U6472_U1 ( .INP(n9578), .ZN(U6472_n1) );
  AND2X1 U6473_U2 ( .IN1(WX663), .IN2(U6473_n1), .Q(WX726) );
  INVX0 U6473_U1 ( .INP(n9578), .ZN(U6473_n1) );
  AND2X1 U6474_U2 ( .IN1(WX661), .IN2(U6474_n1), .Q(WX724) );
  INVX0 U6474_U1 ( .INP(n9578), .ZN(U6474_n1) );
  AND2X1 U6475_U2 ( .IN1(WX659), .IN2(U6475_n1), .Q(WX722) );
  INVX0 U6475_U1 ( .INP(n9578), .ZN(U6475_n1) );
  AND2X1 U6476_U2 ( .IN1(WX657), .IN2(U6476_n1), .Q(WX720) );
  INVX0 U6476_U1 ( .INP(n9578), .ZN(U6476_n1) );
  AND2X1 U6477_U2 ( .IN1(WX655), .IN2(U6477_n1), .Q(WX718) );
  INVX0 U6477_U1 ( .INP(n9578), .ZN(U6477_n1) );
  AND2X1 U6478_U2 ( .IN1(WX653), .IN2(U6478_n1), .Q(WX716) );
  INVX0 U6478_U1 ( .INP(n9578), .ZN(U6478_n1) );
  AND2X1 U6479_U2 ( .IN1(test_so2), .IN2(U6479_n1), .Q(WX714) );
  INVX0 U6479_U1 ( .INP(n9578), .ZN(U6479_n1) );
  AND2X1 U6480_U2 ( .IN1(WX649), .IN2(U6480_n1), .Q(WX712) );
  INVX0 U6480_U1 ( .INP(n9577), .ZN(U6480_n1) );
  AND2X1 U6481_U2 ( .IN1(WX647), .IN2(U6481_n1), .Q(WX710) );
  INVX0 U6481_U1 ( .INP(n9577), .ZN(U6481_n1) );
  AND2X1 U6482_U2 ( .IN1(WX645), .IN2(U6482_n1), .Q(WX708) );
  INVX0 U6482_U1 ( .INP(n9577), .ZN(U6482_n1) );
endmodule

