module s38584 ( CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, 
        g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, 
        g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, 
        g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, 
        g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, 
        g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, 
        g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, 
        g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, 
        g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, 
        g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, 
        g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, 
        g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, 
        g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, 
        g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, 
        g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, 
        g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, 
        g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, 
        g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, 
        g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, 
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
        g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, 
        g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, 
        g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, 
        g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, 
        g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, 
        g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, 
        g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, 
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, 
        g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, 
        g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, 
        g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, 
        g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, 
        g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, 
        g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, 
        g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g99, test_se, test_si1, 
        test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, 
        test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, 
        test_so8, test_si9, test_so9, test_si10, test_so10, test_si11, 
        test_so11, test_si12, test_so12, test_si13, test_so13, test_si14, 
        test_so14, test_si15, test_so15, test_si16, test_so16, test_si17, 
        test_so17, test_si18, test_so18, test_si19, test_so19, test_si20, 
        test_so20, test_si21, test_so21, test_si22, test_so22, test_si23, 
        test_so23, test_si24, test_so24, test_si25, test_so25, test_si26, 
        test_so26, test_si27, test_so27, test_si28, test_so28, test_si29, 
        test_so29, test_si30, test_so30, test_si31, test_so31, test_si32, 
        test_so32, test_si33, test_so33, test_si34, test_so34, test_si35, 
        test_so35, test_si36, test_so36, test_si37, test_so37, test_si38, 
        test_so38, test_si39, test_so39, test_si40, test_so40, test_si41, 
        test_so41, test_si42, test_so42, test_si43, test_so43, test_si44, 
        test_so44, test_si45, test_so45, test_si46, test_so46, test_si47, 
        test_so47, test_si48, test_so48, test_si49, test_so49, test_si50, 
        test_so50, test_si51, test_so51, test_si52, test_so52, test_si53, 
        test_so53, test_si54, test_so54, test_si55, test_so55, test_si56, 
        test_so56, test_si57, test_so57, test_si58, test_so58, test_si59, 
        test_so59, test_si60, test_so60, test_si61, test_so61, test_si62, 
        test_so62, test_si63, test_so63, test_si64, test_so64, test_si65, 
        test_so65, test_si66, test_so66, test_si67, test_so67, test_si68, 
        test_so68, test_si69, test_so69, test_si70, test_so70, test_si71, 
        test_so71, test_si72, test_so72, test_si73, test_so73, test_si74, 
        test_so74, test_si75, test_so75, test_si76, test_so76, test_si77, 
        test_so77, test_si78, test_so78, test_si79, test_so79, test_si80, 
        test_so80, test_si81, test_so81, test_si82, test_so82, test_si83, 
        test_so83, test_si84, test_so84, test_si85, test_so85, test_si86, 
        test_so86, test_si87, test_so87, test_si88, test_so88, test_si89, 
        test_so89, test_si90, test_so90, test_si91, test_so91, test_si92, 
        test_so92, test_si93, test_so93, test_si94, test_so94, test_si95, 
        test_so95, test_si96, test_so96, test_si97, test_so97, test_si98, 
        test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746,
         g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90,
         g91, g92, g99, test_se, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_si6, test_si7, test_si8, test_si9, test_si10,
         test_si11, test_si12, test_si13, test_si14, test_si15, test_si16,
         test_si17, test_si18, test_si19, test_si20, test_si21, test_si22,
         test_si23, test_si24, test_si25, test_si26, test_si27, test_si28,
         test_si29, test_si30, test_si31, test_si32, test_si33, test_si34,
         test_si35, test_si36, test_si37, test_si38, test_si39, test_si40,
         test_si41, test_si42, test_si43, test_si44, test_si45, test_si46,
         test_si47, test_si48, test_si49, test_si50, test_si51, test_si52,
         test_si53, test_si54, test_si55, test_si56, test_si57, test_si58,
         test_si59, test_si60, test_si61, test_si62, test_si63, test_si64,
         test_si65, test_si66, test_si67, test_si68, test_si69, test_si70,
         test_si71, test_si72, test_si73, test_si74, test_si75, test_si76,
         test_si77, test_si78, test_si79, test_si80, test_si81, test_si82,
         test_si83, test_si84, test_si85, test_si86, test_si87, test_si88,
         test_si89, test_si90, test_si91, test_si92, test_si93, test_si94,
         test_si95, test_si96, test_si97, test_si98, test_si99, test_si100;
  output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g18881, g23612, g23652, g73, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29219, g29220, g29221, g30327, g30331,
         g30332, g31656, g31665, g33533, g34435, g34788, g34839, g36, g44, g53,
         g54, g56, g57, g64, g6744, g6745, g6746, g6747, g6748, g6749, g6750,
         g6751, g6753, g84, g90, g91, g92, g99, test_so10, test_so26,
         test_so35, test_so39, test_so42, test_so44, test_so46, test_so80,
         test_so86, test_so92, test_so100, g34783, n2730, n4836, n4896, n4895,
         n4837, n4921, n4920, n4411, n5045, g559, n4959, g33046, g5057, n5615,
         g34441, g2771, n5544, g33982, g1882, g34007, g2299, g24276, g4040,
         n5530, g30381, g2547, n5782, g30405, g3243, g25604, g452, g30416,
         g3542, g30466, g5232, g25736, g5813, g34617, g33974, g1744, g30505,
         g5909, g33554, g1802, n5536, g30432, g3554, g33064, g6219, n5385,
         g34881, g807, n5479, g6031, g24216, g847, n5709, g24232, n9367,
         DFF_24_n1, g34733, g4172, n5493, g34882, g4372, g33026, g3512, g31867,
         n5471, g25668, g3490, n5454, g24344, n5432, g4235, g33966, g1600,
         g33550, g1714, n5460, g30393, g3155, n5366, g29248, g2236, g4571,
         g4555, g24274, g3698, g33973, g1736, n5817, g30360, g1968, n5664,
         g34460, g30494, g5607, g30384, g2657, n5316, g24340, n5439, g29223,
         g490, n5708, g26881, g311, n5317, g34252, g772, n5334, g30489, g5587,
         g29301, g6177, n5874, g6377, g33022, g3167, n5652, g30496, g5615,
         g33043, g4567, g29263, g30533, g6287, g24256, n5302, g34015, g2563,
         n5816, g34031, g4776, n5707, g34452, g4593, n5303, g34646, g6199,
         n5644, g34001, g2295, n5815, g25633, g1384, g24259, g1339, g33049,
         g5180, n5384, g34609, g2844, g31869, g1024, g30490, g30427, g3598,
         g21894, g4264, g33965, g767, n5333, g34645, g5853, n5499, g33571,
         g2089, g34267, g4933, g26971, g4521, n5752, g34644, g5507, n5643,
         g30534, g6291, g33535, g294, n5680, g30498, g25728, g25743, g25684,
         g3813, g25613, g562, g34438, g608, n5475, g24244, g1205, n5547,
         g30439, g3909, g30541, g6259, g30519, g5905, g25621, g921, g34807,
         g2955, g25599, g203, g24235, g34036, g4878, n5283, g30476, g5204,
         g30429, g3606, g32997, g1926, n5510, g33063, g6215, n5651, g30424,
         g3586, g32977, g291, n5679, g34026, g4674, n5440, g30420, g3570,
         g33560, g29226, g676, n5751, g25619, g843, g34455, g4332, n5540,
         g30457, g4153, g33625, g6336, n5592, g34790, g622, n5672, g30414,
         g3506, n5576, g26966, g4558, g25656, g3111, g30390, g25688, g34727,
         g939, n5415, g25594, g278, n5627, g26963, g4492, g34034, g4864, n5318,
         g33541, g1036, g28093, g24236, g1178, g30404, g3239, g28051, g718,
         g29303, g6195, g26917, g1135, n5328, g33624, g6395, n5396, g24337,
         g34911, g554, g33963, g496, g34627, g3853, n5641, g29282, g5134,
         n5807, g25676, g33013, g2485, n5509, g32981, g925, n5725, g34976,
         n9357, DFF_150_n1, g30483, g5555, g32994, g1798, n5833, g28070,
         g34806, g2941, g30453, g3905, g33539, g763, n5332, g30526, g6255,
         g26951, g4375, g34035, g4871, n5443, g34636, g4722, n5345, g32978,
         g590, n5472, g30348, g1632, n5836, g24336, n5438, g3100, g24250,
         g29236, g1437, g29298, g6154, n5747, g1579, g30499, g5567, g33976,
         g1752, g32996, g1917, g30335, g744, n5470, g34637, g4737, n5867,
         g25694, DFF_178_n1, g30528, g6267, g24251, g1442, g30521, g26960,
         g4477, n5849, g24239, g34259, g4643, n5382, g30474, g5264, n5703,
         g33016, g2610, g34643, g5160, n5498, g30510, g5933, g29239, g1454,
         g26897, g753, g34729, g1296, g34625, g3151, n5495, g34800, g24353,
         g6727, n5531, g33029, g3530, n5569, g33615, g4104, g24253, g1532,
         g24281, g33997, n9352, g34971, n9351, DFF_206_n1, g34263, g4754,
         n5877, g24237, g1189, n5642, g33584, g2287, n5353, g24280, g4273,
         n5764, g26920, g1389, g33548, g29296, g5835, n5663, g30338, g1171,
         n5363, g21895, g4269, n5763, g33588, g2399, n5762, g34041, g4983,
         n5367, g30495, g5611, g29279, g4572, g25655, g3143, n5882, g34795,
         g2898, g24269, g3343, g30403, g3235, g33042, g30419, g3566, g34023,
         n9348, DFF_228_n1, g28090, g4961, n5770, g34642, g4927, n5879, g30370,
         g2259, n5419, g34448, g2819, n5609, g26946, g5802, g34610, g2852,
         g24209, g417, n5358, g28047, g681, g24206, g437, g26891, g30504,
         g5901, g34798, g2886, g25669, g3494, n5889, g30480, g5511, n5575,
         g33027, g3518, n5645, g33972, g1604, g25697, g5092, g28099, g4831,
         g26947, g4382, n5714, g24350, g6386, g24210, g479, g30455, g3965,
         g28084, g33993, g2008, g736, g30444, g3933, g33537, g222, g25650,
         g3050, n5998, g25625, g1052, g30366, g2122, n5784, g33593, g2465,
         n5523, g30502, g5889, g33036, g4495, g25595, g34462, g33024, g3179,
         n5390, g33552, g1728, n5352, g34014, g2433, g29273, g3835, n5662,
         g25748, g6187, n5453, g34638, g4917, n5408, g30341, g1070, g26899,
         g822, n5422, g30336, g914, n5560, g5339, g26940, g4164, g25622,
         g34447, g2807, n5379, g33613, g4054, n5395, g25749, g6191, n5888,
         g25704, g5077, n5455, g33053, g5523, n5647, g3680, g30555, g6637,
         g25601, g174, n5402, g33971, g1682, g26892, g355, g1087, g26915,
         g1105, n5478, g33008, g30538, g6307, g3802, g25750, g6159, g30369,
         g2255, n5414, g34446, g2815, g29230, g911, n5559, g43, g33975, g1748,
         g30497, g5551, g30418, g3558, g25721, g5499, n5885, g34622, g30438,
         g3901, g34266, g4888, n5863, g30540, g6251, g32986, g1373, g25648,
         g33960, g157, n5678, g34442, g2783, g4281, g30421, g3574, g33573,
         g2112, g34730, g1283, n5635, g24205, g10122_Tj, g4297, n5698, g32979,
         g758, n5331, g4639, n5727, g25763, g6537, n5884, g30481, g5543,
         g30517, g5961, g30539, g6243, g34880, n9340, g24242, n5654, g30436,
         g29265, g3476, n5786, g32990, g1664, g24245, g1246, n5756, g30553,
         g6629, g26907, g246, n6008, g24278, g4049, g26955, g24282, g2932,
         g29276, g4575, g31894, g4098, n5350, g33037, g4498, g26894, g528,
         n5327, g34977, n5477, g25654, g3139, n5447, g33962, g34451, g4584,
         n5539, g34250, g142, n5724, g29295, g5831, n5873, g26905, g239,
         g25629, g1216, n5442, g34792, g2848, g25703, g5022, g32983, g1030,
         g30402, g3231, g25757, g1430, n9336, g33999, g2241, g24262, g1564,
         g25729, g6148, g30558, g6649, g110, g26901, g225, n5597, g26961,
         g33039, g4504, g33059, g5873, n5388, g31899, g5037, n5611, g33007,
         g2319, n5375, g25720, g5495, n5446, g21891, g30462, g5208, g30487,
         g5579, g33058, g5869, n5649, g24261, g1589, n5755, g25730, g5752,
         n5996, g30531, g6279, g30506, g34804, g2975, n5750, g25747, g6167,
         n5430, n5701, g33601, g2599, n5524, g26922, g1448, n5343, g29250,
         g2370, g30459, g5164, n5570, g1333, n5616, g33534, g153, n5677,
         g30543, g6549, n5571, g29275, g4087, n5480, g34030, g34980, g2984,
         n5842, g30451, g3961, g25627, g962, n5630, g34657, g101, g30552,
         g6625, g34979, n9332, DFF_420_n1, g30337, g1018, g24254, g24277,
         g4045, g29237, g1467, g30378, g2461, n5840, g33019, n5300, g33623,
         g5990, n5589, g29235, g1256, n5558, g31902, g5029, n5601, g29306,
         g6519, n5806, g25689, g4169, n5729, g33978, g1816, g26970, g4369,
         g29278, g4578, g34253, g4459, n5765, g29272, g3831, n5872, g33595,
         g2514, g33610, g3288, n5400, g33589, g34605, g2145, n5307, g30350,
         g1700, n5417, g25611, g513, n5548, g2841, n5963, g33619, g5297, n5588,
         g34022, g2763, g34033, g4793, n5368, g34726, g952, g31870, g1263,
         n5674, g33985, g1950, g29283, g5138, n5871, g34003, g2307, g25677,
         g34463, g4664, g33006, g2223, g29292, g5808, n5749, g30557, g6645,
         g33989, g2016, g33033, g3873, n5387, n5699, g34005, g2315, n5802,
         g26932, g2811, g30516, g5957, g33575, g2047, g33032, g30486, g5575,
         g34974, n9327, DFF_477_n1, g25678, g3752, n5994, g30440, g3917, g1585,
         n5757, g26949, g4388, g30530, g6275, g30542, g6311, g25624, g1041,
         g30383, g33597, g2537, g34598, g26957, g4430, g26967, n9325, g28102,
         g4826, g30524, g6239, g26903, g232, g30475, g5268, g34647, g6545,
         n5497, g30377, n9324, g33553, g1772, n5504, g31903, g5052, n5607,
         g25715, g33984, g1890, n5799, g33602, g2629, n5521, g28045, g572,
         n5337, g34603, g2130, n5487, g33035, g4108, n5715, g4308, g24208,
         g475, g990, n5622, g31, n5469, g34970, n9322, DFF_514_n1, g24213,
         g33614, g3990, n5594, g33060, g30362, g1992, g33023, g3171, n5603,
         g26898, g812, n5733, g25618, g832, g30518, g5897, g4570, n5702,
         g26959, g4455, g34801, g2902, g26884, g333, g25600, g168, n5606,
         g26933, g28066, g3684, g33612, g3639, n5591, g24268, g3338, n5527,
         g25716, g5406, n5992, g26906, g269, g24203, g401, g24346, g6040,
         g24207, g441, g25701, n5690, g29269, g3808, n5745, g9, n5468, g34255,
         g30450, g3957, g30456, g4093, n5340, g32991, g1760, n5602, g24348,
         n5437, g34249, g160, n5843, g30371, g2279, n5778, g29268, g3498,
         g29224, g586, n5336, g33017, g2619, n5508, g30339, g1183, n5599,
         g33967, g1608, g33559, g1779, g29255, g2652, g30368, g2193, n5839,
         g30375, g2393, n5421, g28052, g661, g28089, g4950, n5772, g33055,
         g5535, n5566, g30392, g2834, g30343, g1361, g30523, g6235, g24233,
         g1146, n5851, g33018, g32976, g150, n5676, g30349, g1696, n5628,
         g33067, g6555, g26900, g33034, g3881, n5564, g30551, g6621, g25667,
         g3470, n5424, g30452, g3897, g34719, g518, g538, g33607, g2606,
         g26923, g1472, g24211, g33050, g5188, n5567, g24341, g5689, n5529,
         g24201, g405, g30463, g5216, g6494, g34464, g4669, g24243, g996,
         g24335, g4531, g34611, g2860, g34262, g4743, g30546, g6593, g25591,
         g4411, g30347, g1413, g30556, g6641, g6, g33562, g1936, n5534, g55,
         g25610, g504, n5519, g33015, g2587, n5372, g31896, g4480, g34004,
         n9314, g30428, g30485, g5571, g30422, g3578, g25714, g29294, g5827,
         n5809, g30423, g3582, g30529, g6271, g34028, g4688, n5656, g33587,
         g2380, g30460, g5196, g30401, g3227, g33990, n9312, g29309, g6541,
         n5739, g30411, g3203, g33546, g1668, n5598, g28085, g4760, n5775,
         g26904, g262, g33556, g1840, n5451, g25722, g5467, g25605, g460,
         g33062, g6209, g26893, n5704, g28050, g655, g34626, g33583, g2204,
         n5620, g30472, g5256, g34454, g4608, n5274, g34850, g794, n5291,
         g4423, g24272, g3689, n5532, g5685, g24214, g703, n5821, g26909, g862,
         n5682, g30406, g3247, g33569, g2040, n5505, DFF_672_n1, g34628, g4146,
         n5981, g34458, g4633, n5844, g24240, n5304, g34634, g4732, n5296,
         g25700, n5689, g29293, g5817, g33009, g2351, n5511, g33603, g2648,
         g24355, g6736, g34268, g4944, n5875, g25691, g4072, g26890, g29264,
         g3466, g28072, g4116, g31900, g5041, n5605, g26956, g4434, g29271,
         g3827, n5808, g29304, g6500, n5748, g29261, g3133, n5661, g28063,
         g3333, g979, n5320, g34027, g4681, g33961, g298, n5675, g33604,
         g32995, g1894, n5374, g34624, g2988, g30415, g3538, g33536, g301,
         g26888, n9306, DFF_709_n1, g28055, g827, n5728, g24238, g33600, g2555,
         n5351, g28105, g5011, g34721, g199, g29307, g6523, n5870, g30345,
         g34453, g4601, n5365, g32980, g854, n5754, g29238, g1484, n5865,
         g34639, g4922, n5346, g25695, g5080, n5893, g33057, g5863, g26969,
         g4581, n5670, g29253, g2518, g34021, g2567, g26895, g568, n5335,
         g30413, g3263, g30549, g6613, g24347, g25758, g6444, n5990, g34808,
         g2965, g30501, g5857, n5573, g33969, n9303, g34440, g890, n5305,
         g30433, g3562, g21900, g26921, g1404, g29270, g3817, n9302, n6010,
         g33038, g4501, g31865, g26926, g2724, n5301, g28083, g4704, n5771,
         g34797, g22, g2878, g30478, g5220, g34724, g617, n5339, g24212,
         g26883, g316, g32985, g1277, g25761, g6513, n5426, g26886, g336,
         n5824, g34796, g2882, g32982, g33561, g1906, n5503, g26880, g305,
         n5282, g8, g26931, g2799, g34641, g4912, n5297, g34629, g4157, n5983,
         g33598, g2541, n5461, g33576, g2153, n5356, g34720, g550, g26902,
         g255, g29244, g30468, g5240, g26924, g1478, n5289, g33031, g3863,
         g29245, g1959, g29266, g3480, n5868, g30559, g6653, g34794, g2864,
         g28087, g4894, n5774, g30435, g3857, n5572, g25609, g28057, g1002,
         g34439, g776, n5330, g28, n5324, g1236, g34260, g4646, n5712, g33012,
         g2476, g32989, g1657, n5525, g34006, g2375, g63, g358, g26910, g896,
         n5431, g28043, g33021, g3161, g29251, g2384, n5700, g34456, g4616,
         n5608, g26968, g4561, g33991, g2024, n5801, g3451, g26930, g2795,
         g34599, g613, n5474, g28082, g4527, g33557, g1844, g30511, g5937,
         g33045, g30379, g2523, n5281, g24267, n5436, g34020, g2643, g24249,
         g1489, n5850, g25592, g30382, n9295, g29285, g5156, n5734, n5526,
         n9294, g25662, g21896, g33563, g1955, g33622, g33582, g2273, n5458,
         g28086, g4771, n5769, g25744, g6098, n5988, g29262, g3147, n5738,
         g24270, g3347, g33581, g2269, g191, g24266, g2712, g34849, g626,
         n5288, g33618, g2729, g5357, n5393, g34038, g34032, g4709, n5518,
         g34803, g2927, g34459, g4340, n5653, g30509, g5929, g34640, g4907,
         n5295, g28069, g4035, g21899, g2946, g31868, g918, n5673, g26938,
         g4082, g25756, g30363, g30334, g577, n5294, g33970, g1620, g30391,
         g2831, g25615, g667, g33540, g930, n5731, g30445, g3937, g25617, g817,
         n5822, g24247, g1249, g24215, g837, n5562, g33964, g599, n5550,
         g25719, g5475, n5425, g29228, g30514, g5949, g33627, g6682, n5590,
         g24231, g904, g34615, g2873, g30356, g1854, n5785, g25696, g5084,
         n5681, g30493, g5603, n5726, g33594, g2495, n5522, g34009, g2437,
         g30365, g2102, n5666, g33004, g2208, g34018, g25685, g4064, n5416,
         g34040, g4899, n5517, g25639, g2719, n5465, g34029, g4785, n5361,
         g30488, g5583, g34600, g781, n5551, g29300, g6173, n5810, g34802,
         g2917, g25614, g686, g28058, g1252, n5554, g29225, g671, g33580,
         g30532, g6283, g33054, g5527, n5389, g26962, g4489, g33564, g1974,
         n5450, g32984, g1270, n5716, g34039, g4966, n5706, g33065, g6227,
         n5568, g30443, g3929, g29291, g5503, n5737, g24279, g30508, g5925,
         g29232, g1124, g34269, g4955, n5614, g30464, g5224, g33988, g2012,
         g30522, g6203, n5574, g25708, g5120, g30374, g2389, n5631, g26953,
         g4438, g34008, g2429, g34444, g2787, n5610, g34731, g33606, g2675,
         n5457, g24334, n5541, g34265, g4836, n5713, g30340, g1199, g24257,
         n5401, g30482, g5547, g34604, g2138, n5275, g33591, g2338, g30525,
         g6247, g26929, g2791, g30448, g34602, g1291, n2549, g30513, g5945,
         g30469, g5244, g33608, g2759, g33626, g6741, n5398, g34725, g785,
         n5293, g30342, g1259, n5553, g29267, g3484, n5668, g25593, g209,
         n5595, g30548, g6609, g33052, g5517, g34012, g2449, g34017, n9281,
         g24263, g2715, n5299, g26912, g936, n5557, g30364, g2098, n5280,
         g34254, g4462, n5671, g34251, g604, n5473, g30560, g6589, g33983,
         n9280, g24204, g429, g33980, g1870, g34631, g29243, g1825, g25623,
         g1008, n5321, g26950, g4392, n5710, g30431, g3546, g30467, g5236,
         g30353, g1768, n5834, g34467, g4854, g30442, g3925, g29305, g6509,
         g25616, g732, n5732, g29252, g2504, g4519, g4520, g33003, g2185,
         n5376, g34613, g37, g4031, g33570, g2070, n5535, g34734, g4176, n5494,
         g24275, n5435, g4405, g872, g29302, g6181, n5667, g24349, g34264,
         g4765, n5613, g30484, g5563, g25634, g1395, g33567, g1913, g33585,
         g2331, n5513, g30527, g6263, g34978, n9276, DFF_1012_n1, g30447,
         g3945, g347, n5860, g34256, g4473, g25630, g1266, g29290, g5489,
         n5660, g29227, g31872, g2748, n5516, g29287, g5471, g31897, g4540,
         g6723, g30562, g6605, g34011, n9274, g33996, g2173, g21898, g33014,
         g2491, g34465, g4849, g33995, g2169, g30372, n9273, g30545, g30389,
         g33590, g2407, n5459, g34616, g2868, g26927, g2767, g32992, g1783,
         n5596, g25631, g1312, n5466, g30477, g5212, g34632, g4245, n5640,
         g28046, g645, g4291, g26896, g25602, g26916, g1129, n5329, g33578,
         g2227, n5538, g33579, g2246, g30354, g1830, n5413, g30425, g3590,
         g24200, g392, g33544, g1592, n5362, g25764, g6505, g24246, g1221,
         g30507, g5921, g26889, g30333, g218, g32998, g1932, g32987, g1624,
         n5370, g25702, g5062, g29286, g5462, n5744, g34606, g2689, n5347,
         g33070, g6573, n5563, g29240, g1677, g32999, g2028, n5371, g33605,
         g2671, g24255, g26945, g33558, g1848, n5464, g25699, n5669, g29289,
         g5485, n5869, g30388, g2741, n5349, n5482, g29254, g2638, g28074,
         g4122, g34450, g4322, n5506, g30512, g5941, g33572, g2108, n5452, g25,
         g33551, g33538, g595, n5476, g33005, g2217, n5512, g24248, n9267,
         DFF_1092_n1, g33002, g2066, n5832, g24234, g1152, n5618, g30471,
         g5252, g34000, g2165, g34016, g2571, g33048, g5176, n5650, g25628,
         g26934, g2827, g34468, g4859, g24202, g424, g33542, g1274, n5730,
         n9265, g34445, g2803, n5545, g33555, g1821, g34013, g2509, g28091,
         g5073, g26919, n5556, g30554, g6633, g29281, g5124, g30537, g6303,
         g28092, g5069, g34732, g2994, n5634, g28049, g650, g33545, g1636,
         n5549, g30441, g3921, g29247, g24354, g6732, g25636, g1306, n5796,
         g26914, g1061, g25670, g3462, g33998, g2181, n5803, g25626, g956,
         n5341, g33977, g1756, n5804, g29297, g5849, g28071, g4112, g30387,
         n9262, g33577, g2197, n5514, g33592, g26913, g1046, g28044, g482,
         n5820, g26948, g4401, g30344, g1514, n5364, g26885, g329, n5766,
         g33069, g6565, n5386, g34621, g2950, g28059, g1345, g25762, g6533,
         n5445, g34633, g4727, n5312, g24352, g26925, g1536, g30446, g3941,
         g25597, g370, g24342, g5694, g30357, g1858, n5892, g26908, g446,
         g30399, g3219, g29242, g1811, g30547, g6601, g34010, g2441, g33986,
         g1874, g34257, g30544, g6581, g30561, g6597, g5008, n5637, g30430,
         g3610, g34799, g2890, g33565, g1978, g33968, g1612, g34843, g112,
         g34793, g2856, g33566, g1982, n5462, g30465, g28073, g4119, g24351,
         g6390, g30346, g1542, g21893, g4258, g4818, n5636, g31904, g5033,
         g34635, g4717, n5344, g25637, g1554, n5768, g29274, g3849, g30396,
         g3199, g25735, g34037, g4975, n5360, g34791, g790, n5292, g30520,
         g5913, g30358, g1902, n5837, g29299, g6163, g25690, g4125, g28096,
         g4821, g28088, g4939, n5776, g24241, n5392, g30397, g3207, g4483,
         g30409, g29284, g5142, n5658, g30470, g5248, g30367, g2126, g24273,
         g3694, g29288, g5481, n5805, g30359, g1964, n5315, g25698, g5097,
         n5753, g30398, g3215, n9255, g26952, g4427, g26928, g2779, n5694,
         g26954, DFF_1225_n1, g30351, g1720, n5780, g31871, g1367, g5112, g19,
         g26939, g4145, g33994, g2161, n5812, g25596, g376, n5633, g33586,
         g2361, n5537, g21901, g31866, g582, n5552, g33000, g2051, g26918,
         g1193, g30373, g2327, n5841, g28056, g907, n5555, g34601, g947, n5286,
         g30355, g1834, n5665, g30426, g3594, g34805, g2999, g34002, g2303,
         g28053, g29229, g723, n5826, g33620, g5703, n5397, g34722, g546,
         n5492, g33599, g2472, n5619, g30515, g5953, g25649, g33979, g1740,
         g30417, g3550, g25683, g3845, n5886, g33574, g2116, n5463, g30410,
         g30454, g3913, g34024, g33547, g1687, g30386, g2681, n5777, g33596,
         g2533, n5761, g26887, g324, n5827, g34607, g2697, n5308, g31895,
         g4417, g33068, g6561, n5646, g29233, g1141, n5691, g24258, n5655,
         g30376, g33549, g1710, g29308, g6527, n5659, g30408, g3255, g29241,
         g1691, g34620, g2936, g33621, g5644, n5593, g25707, g5152, n5883,
         g24339, g5352, g34443, g2775, n5378, g34619, g2922, g29234, g30503,
         g5893, g30550, g6617, g33001, g2060, n5507, g33040, g4512, g30492,
         g5599, g25664, g3401, n5986, g26944, g4366, g34614, g29260, g3129,
         n5861, g33047, g5170, g24298, g25733, g5821, n5429, g30536, g6299,
         g29246, g2079, g34261, g4698, n5862, g33611, g3703, n5399, g25638,
         g1559, n5441, g34728, n9247, g29222, g411, n5629, g25742, g30449,
         g3953, g34608, g2704, n5377, g24345, g6035, n5528, n9245, g25635,
         g1300, n5483, g25686, g4057, n5711, g30461, g5200, g34466, g4843,
         g31901, g5046, n5578, g29249, g2250, g26882, n5456, g33041, g33011,
         g2453, n5373, g25734, g5841, n5449, n5705, g34618, g2912, g33010,
         g2357, g31864, g164, n5561, g34630, g4253, n5484, g31898, g5016,
         n5369, g25653, g3119, n5423, g25632, g1351, n5322, g32988, g33616,
         g29280, g5115, n5743, g33609, g3352, n5604, g30563, g6657, g33044,
         g4552, g30437, g3893, g30412, g3211, g30491, g5595, g30434, g3614,
         g34612, g29259, g3125, n5781, g25681, g3821, n5428, g25687, g4141,
         n5612, g33617, g30479, g5272, g29256, g2735, n5600, g28054, g728,
         g30535, g6295, g30385, g2661, n5418, g30361, g1988, n5783, g25705,
         g24260, g1548, n5546, g29257, g3106, n5742, g34461, g4659, g34258,
         g4358, n5348, g32993, g1792, n5359, g33992, g2084, g30394, g3187,
         g34449, g4311, n5323, g34019, g2583, n5800, g18597, n9240,
         DFF_1381_n1, g29231, g1094, g25682, g21897, g4284, g30395, g3191,
         g21892, g4239, g4180, n5380, g28048, g691, n5520, g34723, g534, n5490,
         g25598, g385, n5632, g33987, g2004, n5818, g30380, g2527, n5420,
         g5456, g26965, n6007, g25706, g30458, g4507, n5846, g24338, g5348,
         g30400, g3223, g34623, g2970, g24343, g5698, g30473, g5260, g24252,
         g1521, g33028, g3522, n5383, g29258, g3115, g30407, g3251, g26958,
         g34457, g33568, g1996, n5355, g25663, g26964, g4515, g34735, g4300,
         n5639, g30352, n9236, g33543, g1379, g24271, n5433, g33981, g1878,
         g30500, g5619, g34649, g71, g29277, g25612, n5287, g28060, n2505,
         n2499, n2461, n2396, n2668, n3160, n3141, n3122, n3102, g72, n5960,
         n4689, n5961, n4708, n3593, n3589, n3595, n3574, n3570, n3576, n3517,
         n3513, n3519, n3628, n3624, n3630, n3555, n3551, n3557, n3646, n3642,
         n3648, n3536, n3532, n3538, n3611, n3607, n3613, n3006, n3765, n3505,
         n3525, n3635, n4888, n3550, n2595, n2527, n3524, n3005, n3623, n3549,
         n3003, n3007, n3569, n3606, n3588, n3165, n3799, n3033, n3622, n3587,
         n3586, n3605, n3604, n3568, n3567, n3548, n3512, n3511, n3531, n3530,
         n3641, n3640, n3131, n3111, n3907, n3773, n3807, n3950, n3841, n3983,
         n3874, n4014, n4537, n4201, n3745, n3684, n3274, n2982, n2706, n2649,
         n2556, n2509, n2487, n2427, n2423, n2421, n4172, n4173, n4190, n4191,
         n4388, n4210, n3479, n3951, n3404, n3774, n3424, n3842, n3414, n3808,
         n3444, n3908, n3489, n3984, n3434, n3875, n3500, n4015, n3446, n3914,
         n3406, n3780, n3481, n3957, n3426, n3848, n3491, n3990, n3416, n3814,
         n3436, n3881, n3502, n4022, n3501, n4027, n3407, n3785, n3482, n3962,
         n3427, n3853, n3437, n3886, n3417, n3819, n3492, n3995, n3447, n3919,
         n3682, n3272, n2980, n2704, n2647, n2554, n2507, n2485, n2425, n2419,
         n2405, n2760, n2552, n4946, n4198, n2404, n3653, n3581, n4962, n4948,
         n2726, n2727, n3195, n2774, n3116, n4945, n4525, n4518, n3281, n3277,
         n3276, n2989, n2991, n2710, n2707, n3174, n3362, n3676, n2644, n3146,
         n3115, n3833, n3023, n3933, n3729, n4723, n2601, n3664, n3662, n3673,
         n3671, n2607, n3506, n2790, n4490, n4178, n4514, n4196, n3736, n3741,
         n2598, n4814, n4519, n2594, n3084, n2590, n4722, n3125, n3105, n3145,
         n3164, n3910, n3776, n3877, n3810, n4017, n3953, n3986, n3844, n3770,
         n3904, n3804, n3947, n3838, n3871, n3980, n4020, n3495, n3945, n3836,
         n3768, n3869, n3978, n3802, n3902, n2422, n4037, n4034, n4039, n3972,
         n3969, n3929, n3926, n3863, n3860, n4003, n4002, n4032, n4035, n3797,
         n3792, n3790, n3795, n3891, n3893, n3827, n3826, n3896, n4007, n3931,
         n3793, n3924, n3831, n3829, n3927, n3974, n3898, n3970, n4000, n3865,
         n3861, n3824, n3894, n3967, n3858, n4005, n3395, n4956, n5026, n3941,
         n3733, n4798, n4805, n4175, n4193, n3738, n4721, n4523, n4524, n4526,
         n2573, n2577, n2563, n2567, n4938, n4940, n4913, n4915, n4714, n4516,
         n4517, n5111, n4819, n3730, n3121, n3180, n4305, n4283, n2608, n4447,
         n4448, n4402, n4403, n4425, n4426, n4436, n4437, n4391, n4392, n4379,
         n4380, n4414, n4415, n4458, n4459, n5016, n5014, n3064, n3065, n4535,
         n5112, n3675, counter_31, counter_30, counter_29, counter_28,
         counter_27, counter_26, counter_25, counter_24, counter_23,
         counter_22, counter_21, counter_20, counter_19, counter_18,
         counter_17, counter_16, counter_15, counter_14, counter_13,
         counter_12, counter_11, counter_10, counter_9, counter_8, counter_7,
         counter_6, counter_5, counter_4, counter_3, counter_2, counter_1,
         counter_0, carry_31, carry_30, carry_29, carry_28, carry_27, carry_26,
         carry_25, carry_24, carry_23, carry_22, carry_21, carry_20, carry_19,
         carry_18, carry_17, carry_16, carry_15, carry_14, carry_13, carry_12,
         carry_11, carry_10, carry_9, carry_8, carry_7, carry_6, carry_5,
         carry_4, carry_3, carry_2, N31, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N23, N24, N25, N26, N2, N3, N4, N16, N17, N18, N19,
         N20, N21, N22, N27, N28, N29, N30, N1, N32, n37, n87, n73, n86, n85,
         n84, n83, n82, n81, n80, n79, n78, n77, n76, n75, n74, n58, n59, n60,
         n61, n62, n63, n64, Trigger_out, n65, n66, n67, n68, n69, n70, n71,
         n72, n5, n42, n43, n45, g33959, n155, n156, g26801, n171, n220, n233,
         n314, n322, n326, n435, n436, n456, n616, n628, n709, n911, n917,
         n965, n982, n1123, n1136, n1413, n1430, n7671, n7672, n7675, n7677,
         n7680, n7681, n7684, n7685, n7686, n7689, n7691, n7692, n7693, n7696,
         n7708, n7709, n7710, n7712, n7713, n7718, n7722, n7723, n7724, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7738,
         n7739, n7740, n7742, n7743, n7744, n7746, n7747, n7749, n7750, n7751,
         n7752, n7753, n7757, n7758, n7765, n7766, n7768, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7791, n7792, n7793, n7794,
         n7796, n7797, n7804, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7822, n7826, n7827, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7854,
         n7856, n7857, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7876, n7880, n7884,
         n7891, n7895, n7899, n7901, n7904, n7905, n7906, n7907, n7908, n7909,
         n7911, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7954,
         n7956, n7958, n7960, n7962, n7964, n7966, n7967, n7969, n7971, n7973,
         n7975, n7976, n7978, n7980, n7982, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7999,
         n8000, n8001, n8002, n8003, n8004, n8007, n8010, n8013, n8016, n8019,
         n8022, n8025, n8028, n8038, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8059, n8069, n8074, n8078, n8083, n8088, n8093, n8095, n8097, n8099,
         n8101, n8103, n8105, n8107, n8109, n8111, n8113, n8115, n8117, n8119,
         n8121, n8122, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8159, n8160, n8161, n8164, n8167, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, g31860, g31862, g31863,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9237, n9238, n9239, n9241, n9242, n9243,
         n9244, n9246, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9256,
         n9257, n9258, n9259, n9260, n9261, n9263, n9264, n9266, n9268, n9269,
         n9270, n9271, n9272, n9275, n9277, n9278, n9279, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9296,
         n9297, n9298, n9299, n9300, n9301, n9304, n9305, n9307, n9308, n9309,
         n9310, n9311, n9313, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9323, n9326, n9328, n9329, n9330, n9331, n9333, n9334, n9335, n9337,
         n9338, n9339, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9349,
         n9350, n9353, n9354, n9355, n9356, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, U5353_n1, U5355_n1, U5961_n1,
         U5962_n1, U5963_n1, U5964_n1, U5965_n1, U5966_n1, U5967_n1, U5968_n1,
         U6100_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1, U6216_n1,
         U6217_n1, U6218_n1, U6279_n1, U6280_n1, U6281_n1, U6282_n1, U6283_n1,
         U6284_n1, U6285_n1, U6286_n1, U6287_n1, U6288_n1, U6289_n1, U6290_n1,
         U6291_n1, U6292_n1, U6338_n1, U6341_n1, U6342_n1, U6343_n1, U6344_n1,
         U6345_n1, U6346_n1, U6347_n1, U6348_n1, U6349_n1, U6350_n1, U6351_n1,
         U6352_n1, U6353_n1, U6354_n1, U6355_n1, U6356_n1, U6357_n1, U6358_n1,
         U6359_n1, U6360_n1, U6361_n1, U6362_n1, U6363_n1, U6364_n1, U6365_n1,
         U6366_n1, U6367_n1, U6368_n1, U6369_n1, U6370_n1, U6371_n1, U6372_n1,
         U6373_n1, U6374_n1, U6375_n1, U6417_n1, U6446_n1, U6465_n1, U6497_n1,
         U6523_n1, U6542_n1, U6552_n1, U6553_n1, U6554_n1, U6555_n1, U6556_n1,
         U6559_n1, U6560_n1, U6561_n1, U6570_n1, U6911_n1, U6912_n1, U6917_n1,
         U6926_n1, U6927_n1, U6929_n1, U6931_n1, U6932_n1, U6933_n1, U6934_n1,
         U6935_n1, U6936_n1, U6937_n1, U6938_n1, U6939_n1, U6940_n1, U6941_n1,
         U6944_n1, U6950_n1, U6954_n1, U6955_n1, U6956_n1, U6957_n1, U7174_n1,
         U7248_n1, U7249_n1, U7402_n1, U7405_n1, U7413_n1, U7416_n1, U7427_n1,
         U7438_n1, U7449_n1, U7455_n1, U7464_n1, U7467_n1, U7482_n1, U7492_n1,
         U7513_n1, U7516_n1, U7549_n1, U7561_n1, U7574_n1, U7577_n1, U7585_n1,
         U7595_n1, U7614_n1, U7621_n1, U7629_n1, U7636_n1, U7639_n1, U7649_n1,
         U7652_n1, U7668_n1, U7673_n1, U7690_n1, U7707_n1, U7712_n1, U7792_n1,
         U7794_n1, U7895_n1, U7897_n1, U7977_n1, U8034_n1, U8036_n1, U8050_n1,
         U8055_n1, U8060_n1, U8070_n1, U8074_n1, U8088_n1, U8112_n1, U8113_n1,
         U8147_n1, U8165_n1, U8185_n1, U8192_n1, U8210_n1, U8223_n1, U8224_n1,
         U8281_n1, U8307_n1, U8974_n1, U8975_n1, U9065_n1, U9070_n1, U9075_n1,
         U9076_n1, U9080_n1, U9084_n1, U9085_n1, U9086_n1, U9090_n1, U9098_n1,
         U9099_n1, U9101_n1, U9107_n1, U9111_n1, U9116_n1, U9120_n1, U9124_n1,
         U9128_n1, U9132_n1, U9136_n1, U9315_n1, U9453_n1, U9825_n1, U9886_n1,
         U9927_n1, U9953_n1, U9957_n1, U9958_n1, U9968_n1, U9972_n1, U9992_n1,
         U10314_n1, U10318_n1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g34597 = 1'b0;
  assign g24173 = g100;
  assign g24174 = g113;
  assign g24175 = g114;
  assign g24176 = g115;
  assign g24177 = g116;
  assign g24178 = g120;
  assign g24179 = g124;
  assign g24180 = g125;
  assign g24181 = g126;
  assign g24182 = g127;
  assign g24183 = g134;
  assign g24184 = g135;
  assign g29218 = g18881;
  assign g30329 = g23612;
  assign g30330 = g23652;
  assign g24167 = g73;
  assign g20763 = g29211;
  assign g20899 = g29212;
  assign g20557 = g29213;
  assign g20652 = g29214;
  assign g20901 = g29215;
  assign g21176 = g29216;
  assign g21270 = g29217;
  assign g20654 = g29219;
  assign g21245 = g29220;
  assign g21292 = g29221;
  assign g23002 = g30327;
  assign g23759 = g30331;
  assign g23683 = g30332;
  assign g34436 = g31656;
  assign g34437 = g31665;
  assign g27831 = g33533;
  assign g31521 = g34435;
  assign g33894 = g34788;
  assign g34956 = g34839;
  assign g21698 = g36;
  assign g24185 = g44;
  assign g24161 = g53;
  assign g24162 = g54;
  assign g24163 = g56;
  assign g24164 = g57;
  assign g24165 = g64;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18101 = g6746;
  assign g18097 = g6747;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18100 = g6751;
  assign g18092 = g6753;
  assign g24168 = g84;
  assign g24169 = g90;
  assign g24170 = g91;
  assign g24171 = g92;
  assign g24172 = g99;
  assign g31861 = test_so10;
  assign g25219 = test_so10;
  assign g13881 = test_so26;
  assign g9615 = test_so35;
  assign g8785 = test_so39;
  assign g8291 = test_so42;
  assign g17316 = test_so44;
  assign g8178 = test_so46;
  assign g12470 = test_so80;
  assign g11447 = test_so86;
  assign g9682 = test_so92;
  assign g29210 = test_so100;
  assign g20049 = test_so100;
  assign g24166 = g72;
  assign g28753 = g33959;
  assign g32975 = g26801;
  assign g25114 = g31860;
  assign g25259 = g31862;
  assign g25167 = g31863;

  SDFFX1 DFF_0_Q_reg ( .D(g33046), .SI(test_si1), .SE(n8248), .CLK(n8662), .Q(
        g5057), .QN(n5615) );
  SDFFX1 DFF_1_Q_reg ( .D(g34441), .SI(g5057), .SE(n8263), .CLK(n8677), .Q(
        g2771), .QN(n5544) );
  SDFFX1 DFF_2_Q_reg ( .D(g33982), .SI(g2771), .SE(n8287), .CLK(n8701), .Q(
        g1882) );
  SDFFX1 DFF_4_Q_reg ( .D(g34007), .SI(g1882), .SE(n8287), .CLK(n8701), .Q(
        g2299) );
  SDFFX1 DFF_5_Q_reg ( .D(g24276), .SI(g2299), .SE(n8334), .CLK(n8748), .Q(
        g4040), .QN(n5530) );
  SDFFX1 DFF_6_Q_reg ( .D(g30381), .SI(g4040), .SE(n8268), .CLK(n8682), .Q(
        g2547), .QN(n5782) );
  SDFFX1 DFF_7_Q_reg ( .D(g9048), .SI(g2547), .SE(n8305), .CLK(n8719), .Q(g559) );
  SDFFX1 DFF_9_Q_reg ( .D(g30405), .SI(g559), .SE(n8320), .CLK(n8734), .Q(
        g3243) );
  SDFFX1 DFF_10_Q_reg ( .D(g25604), .SI(g3243), .SE(n8257), .CLK(n8671), .Q(
        g452), .QN(n8002) );
  SDFFX1 DFF_12_Q_reg ( .D(g30416), .SI(g452), .SE(n8305), .CLK(n8719), .Q(
        g3542), .QN(n7891) );
  SDFFX1 DFF_13_Q_reg ( .D(g30466), .SI(g3542), .SE(n8253), .CLK(n8667), .Q(
        g5232) );
  SDFFX1 DFF_14_Q_reg ( .D(g25736), .SI(g5232), .SE(n8335), .CLK(n8749), .Q(
        g5813), .QN(n7793) );
  SDFFX1 DFF_15_Q_reg ( .D(g34617), .SI(g5813), .SE(n8270), .CLK(n8684), .Q(
        test_so1) );
  SDFFX1 DFF_16_Q_reg ( .D(g33974), .SI(test_si2), .SE(n8272), .CLK(n8686), 
        .Q(g1744) );
  SDFFX1 DFF_17_Q_reg ( .D(g30505), .SI(g1744), .SE(n8288), .CLK(n8702), .Q(
        g5909), .QN(n8013) );
  SDFFX1 DFF_18_Q_reg ( .D(g33554), .SI(g5909), .SE(n8273), .CLK(n8687), .Q(
        g1802), .QN(n5536) );
  SDFFX1 DFF_19_Q_reg ( .D(g30432), .SI(g1802), .SE(n8306), .CLK(n8720), .Q(
        g3554) );
  SDFFX1 DFF_20_Q_reg ( .D(g33064), .SI(g3554), .SE(n8336), .CLK(n8750), .Q(
        g6219), .QN(n5385) );
  SDFFX1 DFF_21_Q_reg ( .D(g34881), .SI(g6219), .SE(n8299), .CLK(n8713), .Q(
        g807), .QN(n5479) );
  SDFFX1 DFF_22_Q_reg ( .D(g17715), .SI(g807), .SE(n8324), .CLK(n8738), .Q(
        g6031) );
  SDFFX1 DFF_23_Q_reg ( .D(g24216), .SI(g6031), .SE(n8257), .CLK(n8671), .Q(
        g847), .QN(n5709) );
  SDFFX1 DFF_24_Q_reg ( .D(g24232), .SI(g847), .SE(n8352), .CLK(n8766), .Q(
        n9367), .QN(DFF_24_n1) );
  SDFFX1 DFF_25_Q_reg ( .D(g34733), .SI(n9367), .SE(n8268), .CLK(n8682), .Q(
        g4172), .QN(n5493) );
  SDFFX1 DFF_26_Q_reg ( .D(g34882), .SI(g4172), .SE(n8304), .CLK(n8718), .Q(
        g4372) );
  SDFFX1 DFF_27_Q_reg ( .D(g33026), .SI(g4372), .SE(n8304), .CLK(n8718), .Q(
        g3512), .QN(n8146) );
  SDFFX1 DFF_28_Q_reg ( .D(g31867), .SI(g3512), .SE(n8316), .CLK(n8730), .Q(
        test_so2), .QN(n5471) );
  SDFFX1 DFF_29_Q_reg ( .D(g25668), .SI(test_si3), .SE(n8315), .CLK(n8729), 
        .Q(g3490), .QN(n5454) );
  SDFFX1 DFF_30_Q_reg ( .D(g24344), .SI(g3490), .SE(n8315), .CLK(n8729), .Q(
        g12350), .QN(n5432) );
  SDFFX1 DFF_31_Q_reg ( .D(g8920), .SI(g12350), .SE(n8315), .CLK(n8729), .Q(
        g4235), .QN(n7920) );
  SDFFX1 DFF_32_Q_reg ( .D(g33966), .SI(g4235), .SE(n8315), .CLK(n8729), .Q(
        g1600) );
  SDFFX1 DFF_33_Q_reg ( .D(g33550), .SI(g1600), .SE(n8296), .CLK(n8710), .Q(
        g1714), .QN(n5460) );
  SDFFX1 DFF_34_Q_reg ( .D(g16656), .SI(g1714), .SE(n8296), .CLK(n8710), .Q(
        g14451) );
  SDFFX1 DFF_35_Q_reg ( .D(g30393), .SI(g14451), .SE(n8326), .CLK(n8740), .Q(
        g3155), .QN(n5366) );
  SDFFX1 DFF_37_Q_reg ( .D(g29248), .SI(g3155), .SE(n8312), .CLK(n8726), .Q(
        g2236), .QN(n7908) );
  SDFFX1 DFF_38_Q_reg ( .D(g4571), .SI(g2236), .SE(n8339), .CLK(n8753), .Q(
        g4555) );
  SDFFX1 DFF_39_Q_reg ( .D(g24274), .SI(g4555), .SE(n8279), .CLK(n8693), .Q(
        g3698), .QN(n7989) );
  SDFFX1 DFF_41_Q_reg ( .D(g33973), .SI(g3698), .SE(n8272), .CLK(n8686), .Q(
        g1736), .QN(n5817) );
  SDFFX1 DFF_42_Q_reg ( .D(g30360), .SI(g1736), .SE(n8271), .CLK(n8685), .Q(
        g1968), .QN(n5664) );
  SDFFX1 DFF_43_Q_reg ( .D(g34460), .SI(g1968), .SE(n8331), .CLK(n8745), .Q(
        test_so3), .QN(n8226) );
  SDFFX1 DFF_44_Q_reg ( .D(g30494), .SI(test_si4), .SE(n8260), .CLK(n8674), 
        .Q(g5607) );
  SDFFX1 DFF_45_Q_reg ( .D(g30384), .SI(g5607), .SE(n8260), .CLK(n8674), .Q(
        g2657), .QN(n5316) );
  SDFFX1 DFF_46_Q_reg ( .D(g24340), .SI(g2657), .SE(n8320), .CLK(n8734), .Q(
        g12300), .QN(n5439) );
  SDFFX1 DFF_47_Q_reg ( .D(g29223), .SI(g12300), .SE(n8323), .CLK(n8737), .Q(
        g490), .QN(n5708) );
  SDFFX1 DFF_48_Q_reg ( .D(g26881), .SI(g490), .SE(n8345), .CLK(n8759), .Q(
        g311), .QN(n5317) );
  SDFFX1 DFF_50_Q_reg ( .D(g34252), .SI(g311), .SE(n8316), .CLK(n8730), .Q(
        g772), .QN(n5334) );
  SDFFX1 DFF_51_Q_reg ( .D(g30489), .SI(g772), .SE(n8259), .CLK(n8673), .Q(
        g5587) );
  SDFFX1 DFF_52_Q_reg ( .D(g29301), .SI(g5587), .SE(n8256), .CLK(n8670), .Q(
        g6177), .QN(n5874) );
  SDFFX1 DFF_53_Q_reg ( .D(g17743), .SI(g6177), .SE(n8317), .CLK(n8731), .Q(
        g6377) );
  SDFFX1 DFF_54_Q_reg ( .D(g33022), .SI(g6377), .SE(n8326), .CLK(n8740), .Q(
        g3167), .QN(n5652) );
  SDFFX1 DFF_55_Q_reg ( .D(g30496), .SI(g3167), .SE(n8250), .CLK(n8664), .Q(
        g5615) );
  SDFFX1 DFF_56_Q_reg ( .D(g33043), .SI(g5615), .SE(n8321), .CLK(n8735), .Q(
        g4567) );
  SDFFX1 DFF_58_Q_reg ( .D(g29263), .SI(g4567), .SE(n8352), .CLK(n8766), .Q(
        test_so4), .QN(n8224) );
  SDFFX1 DFF_59_Q_reg ( .D(g30533), .SI(test_si5), .SE(n8351), .CLK(n8765), 
        .Q(g6287) );
  SDFFX1 DFF_60_Q_reg ( .D(g24256), .SI(g6287), .SE(n8262), .CLK(n8676), .Q(
        g7946), .QN(n5302) );
  SDFFX1 DFF_61_Q_reg ( .D(g34015), .SI(g7946), .SE(n8303), .CLK(n8717), .Q(
        g2563), .QN(n5816) );
  SDFFX1 DFF_62_Q_reg ( .D(g34031), .SI(g2563), .SE(n8327), .CLK(n8741), .Q(
        g4776), .QN(n5707) );
  SDFFX1 DFF_63_Q_reg ( .D(g34452), .SI(g4776), .SE(n8327), .CLK(n8741), .Q(
        g4593), .QN(n5303) );
  SDFFX1 DFF_64_Q_reg ( .D(g34646), .SI(g4593), .SE(n8327), .CLK(n8741), .Q(
        g6199), .QN(n5644) );
  SDFFX1 DFF_65_Q_reg ( .D(g34001), .SI(g6199), .SE(n8287), .CLK(n8701), .Q(
        g2295), .QN(n5815) );
  SDFFX1 DFF_66_Q_reg ( .D(g25633), .SI(g2295), .SE(n8261), .CLK(n8675), .Q(
        g1384), .QN(n7693) );
  SDFFX1 DFF_67_Q_reg ( .D(g24259), .SI(g1384), .SE(n8314), .CLK(n8728), .Q(
        g1339) );
  SDFFX1 DFF_68_Q_reg ( .D(g33049), .SI(g1339), .SE(n8304), .CLK(n8718), .Q(
        g5180), .QN(n5384) );
  SDFFX1 DFF_69_Q_reg ( .D(g34609), .SI(g5180), .SE(n8289), .CLK(n8703), .Q(
        g2844) );
  SDFFX1 DFF_70_Q_reg ( .D(g31869), .SI(g2844), .SE(n8262), .CLK(n8676), .Q(
        g1024), .QN(n7815) );
  SDFFX1 DFF_71_Q_reg ( .D(g30490), .SI(g1024), .SE(n8260), .CLK(n8674), .Q(
        test_so5) );
  SDFFX1 DFF_72_Q_reg ( .D(g30427), .SI(test_si6), .SE(n8305), .CLK(n8719), 
        .Q(g3598) );
  SDFFX1 DFF_73_Q_reg ( .D(g21894), .SI(g3598), .SE(n8305), .CLK(n8719), .Q(
        g4264) );
  SDFFX1 DFF_74_Q_reg ( .D(g33965), .SI(g4264), .SE(n8316), .CLK(n8730), .Q(
        g767), .QN(n5333) );
  SDFFX1 DFF_75_Q_reg ( .D(g34645), .SI(g767), .SE(n8316), .CLK(n8730), .Q(
        g5853), .QN(n5499) );
  SDFFX1 DFF_76_Q_reg ( .D(g16874), .SI(g5853), .SE(n8343), .CLK(n8757), .Q(
        g13865) );
  SDFFX1 DFF_77_Q_reg ( .D(g33571), .SI(g13865), .SE(n8291), .CLK(n8705), .Q(
        g2089) );
  SDFFX1 DFF_78_Q_reg ( .D(g34267), .SI(g2089), .SE(n8295), .CLK(n8709), .Q(
        g4933) );
  SDFFX1 DFF_79_Q_reg ( .D(g26971), .SI(g4933), .SE(n8350), .CLK(n8764), .Q(
        g4521), .QN(n5752) );
  SDFFX1 DFF_80_Q_reg ( .D(g34644), .SI(g4521), .SE(n8350), .CLK(n8764), .Q(
        g5507), .QN(n5643) );
  SDFFX1 DFF_81_Q_reg ( .D(g16627), .SI(g5507), .SE(n8297), .CLK(n8711), .Q(
        g16656), .QN(n8088) );
  SDFFX1 DFF_82_Q_reg ( .D(g30534), .SI(g16656), .SE(n8297), .CLK(n8711), .Q(
        g6291) );
  SDFFX1 DFF_83_Q_reg ( .D(g33535), .SI(g6291), .SE(n8276), .CLK(n8690), .Q(
        g294), .QN(n5680) );
  SDFFX1 DFF_84_Q_reg ( .D(g30498), .SI(g294), .SE(n8354), .CLK(n8768), .Q(
        test_so6) );
  SDFFX1 DFF_85_Q_reg ( .D(g25728), .SI(test_si7), .SE(n8335), .CLK(n8749), 
        .Q(g9617) );
  SDFFX1 DFF_86_Q_reg ( .D(g25743), .SI(g9617), .SE(n8278), .CLK(n8692), .Q(
        g9741), .QN(n7723) );
  SDFFX1 DFF_87_Q_reg ( .D(g25684), .SI(g9741), .SE(n8278), .CLK(n8692), .Q(
        g3813), .QN(n7776) );
  SDFFX1 DFF_88_Q_reg ( .D(g25613), .SI(g3813), .SE(n8282), .CLK(n8696), .Q(
        g562), .QN(n7686) );
  SDFFX1 DFF_89_Q_reg ( .D(g34438), .SI(g562), .SE(n8283), .CLK(n8697), .Q(
        g608), .QN(n5475) );
  SDFFX1 DFF_90_Q_reg ( .D(g24244), .SI(g608), .SE(n8284), .CLK(n8698), .Q(
        g1205), .QN(n5547) );
  SDFFX1 DFF_91_Q_reg ( .D(g30439), .SI(g1205), .SE(n8265), .CLK(n8679), .Q(
        g3909), .QN(n8019) );
  SDFFX1 DFF_92_Q_reg ( .D(g30541), .SI(g3909), .SE(n8351), .CLK(n8765), .Q(
        g6259), .QN(n8119) );
  SDFFX1 DFF_93_Q_reg ( .D(g30519), .SI(g6259), .SE(n8351), .CLK(n8765), .Q(
        g5905) );
  SDFFX1 DFF_94_Q_reg ( .D(g25621), .SI(g5905), .SE(n8351), .CLK(n8765), .Q(
        g921), .QN(n7827) );
  SDFFX1 DFF_95_Q_reg ( .D(g34807), .SI(g921), .SE(n8248), .CLK(n8662), .Q(
        g2955), .QN(n7820) );
  SDFFX1 DFF_96_Q_reg ( .D(g25599), .SI(g2955), .SE(n8291), .CLK(n8705), .Q(
        g203) );
  SDFFX1 DFF_98_Q_reg ( .D(g24235), .SI(g203), .SE(n8291), .CLK(n8705), .Q(
        test_so7), .QN(n8207) );
  SDFFX1 DFF_99_Q_reg ( .D(g34036), .SI(test_si8), .SE(n8302), .CLK(n8716), 
        .Q(g4878), .QN(n5283) );
  SDFFX1 DFF_100_Q_reg ( .D(g30476), .SI(g4878), .SE(n8302), .CLK(n8716), .Q(
        g5204), .QN(n8040) );
  SDFFX1 DFF_101_Q_reg ( .D(g17580), .SI(g5204), .SE(n8302), .CLK(n8716), .Q(
        g17604), .QN(n8074) );
  SDFFX1 DFF_102_Q_reg ( .D(g30429), .SI(g17604), .SE(n8306), .CLK(n8720), .Q(
        g3606) );
  SDFFX1 DFF_103_Q_reg ( .D(g32997), .SI(g3606), .SE(n8281), .CLK(n8695), .Q(
        g1926), .QN(n5510) );
  SDFFX1 DFF_104_Q_reg ( .D(g33063), .SI(g1926), .SE(n8336), .CLK(n8750), .Q(
        g6215), .QN(n5651) );
  SDFFX1 DFF_105_Q_reg ( .D(g30424), .SI(g6215), .SE(n8305), .CLK(n8719), .Q(
        g3586) );
  SDFFX1 DFF_106_Q_reg ( .D(g32977), .SI(g3586), .SE(n8276), .CLK(n8690), .Q(
        g291), .QN(n5679) );
  SDFFX1 DFF_107_Q_reg ( .D(g34026), .SI(g291), .SE(n8331), .CLK(n8745), .Q(
        g4674), .QN(n5440) );
  SDFFX1 DFF_108_Q_reg ( .D(g30420), .SI(g4674), .SE(n8305), .CLK(n8719), .Q(
        g3570) );
  SDFFX1 DFF_109_Q_reg ( .D(g12368), .SI(g3570), .SE(n8305), .CLK(n8719), .Q(
        g9048), .QN(n7672) );
  SDFFX1 DFF_110_Q_reg ( .D(g17739), .SI(g9048), .SE(n8307), .CLK(n8721), .Q(
        g17607), .QN(n7958) );
  SDFFX1 DFF_111_Q_reg ( .D(g33560), .SI(g17607), .SE(n8345), .CLK(n8759), .Q(
        test_so8), .QN(n8205) );
  SDFFX1 DFF_112_Q_reg ( .D(g29226), .SI(test_si9), .SE(n8264), .CLK(n8678), 
        .Q(g676), .QN(n5751) );
  SDFFX1 DFF_113_Q_reg ( .D(g25619), .SI(g676), .SE(n8325), .CLK(n8739), .Q(
        g843), .QN(n7804) );
  SDFFX1 DFF_115_Q_reg ( .D(g34455), .SI(g843), .SE(n8327), .CLK(n8741), .Q(
        g4332), .QN(n5540) );
  SDFFX1 DFF_116_Q_reg ( .D(g30457), .SI(g4332), .SE(n8267), .CLK(n8681), .Q(
        g4153), .QN(n8182) );
  SDFFX1 DFF_117_Q_reg ( .D(g14694), .SI(g4153), .SE(n8286), .CLK(n8700), .Q(
        g17711), .QN(n7975) );
  SDFFX1 DFF_118_Q_reg ( .D(g33625), .SI(g17711), .SE(n8256), .CLK(n8670), .Q(
        g6336), .QN(n5592) );
  SDFFX1 DFF_119_Q_reg ( .D(g34790), .SI(g6336), .SE(n8282), .CLK(n8696), .Q(
        g622), .QN(n5672) );
  SDFFX1 DFF_120_Q_reg ( .D(g30414), .SI(g622), .SE(n8330), .CLK(n8744), .Q(
        g3506), .QN(n5576) );
  SDFFX1 DFF_121_Q_reg ( .D(g26966), .SI(g3506), .SE(n8339), .CLK(n8753), .Q(
        g4558) );
  SDFFX1 DFF_123_Q_reg ( .D(g17649), .SI(g4558), .SE(n8339), .CLK(n8753), .Q(
        g17685), .QN(n8093) );
  SDFFX1 DFF_124_Q_reg ( .D(g25656), .SI(g17685), .SE(n8342), .CLK(n8756), .Q(
        g3111), .QN(n7773) );
  SDFFX1 DFF_125_Q_reg ( .D(g30390), .SI(g3111), .SE(n8280), .CLK(n8694), .Q(
        g29217) );
  SDFFX1 DFF_126_Q_reg ( .D(g25688), .SI(g29217), .SE(n8280), .CLK(n8694), .Q(
        test_so9) );
  SDFFX1 DFF_127_Q_reg ( .D(g34727), .SI(test_si10), .SE(n8276), .CLK(n8690), 
        .Q(g939), .QN(n5415) );
  SDFFX1 DFF_128_Q_reg ( .D(g25594), .SI(g939), .SE(n8276), .CLK(n8690), .Q(
        g278), .QN(n5627) );
  SDFFX1 DFF_129_Q_reg ( .D(g26963), .SI(g278), .SE(n8341), .CLK(n8755), .Q(
        g4492) );
  SDFFX1 DFF_130_Q_reg ( .D(g34034), .SI(g4492), .SE(n8302), .CLK(n8716), .Q(
        g4864), .QN(n5318) );
  SDFFX1 DFF_131_Q_reg ( .D(g33541), .SI(g4864), .SE(n8263), .CLK(n8677), .Q(
        g1036), .QN(n7779) );
  SDFFX1 DFF_132_Q_reg ( .D(g28093), .SI(g1036), .SE(n8254), .CLK(n8668), .Q(
        g29220) );
  SDFFX1 DFF_133_Q_reg ( .D(g24236), .SI(g29220), .SE(n8254), .CLK(n8668), .Q(
        g1178) );
  SDFFX1 DFF_134_Q_reg ( .D(g30404), .SI(g1178), .SE(n8319), .CLK(n8733), .Q(
        g3239) );
  SDFFX1 DFF_135_Q_reg ( .D(g28051), .SI(g3239), .SE(n8322), .CLK(n8736), .Q(
        g718), .QN(n7905) );
  SDFFX1 DFF_136_Q_reg ( .D(g29303), .SI(g718), .SE(n8336), .CLK(n8750), .Q(
        g6195) );
  SDFFX1 DFF_137_Q_reg ( .D(g26917), .SI(g6195), .SE(n8249), .CLK(n8663), .Q(
        g1135), .QN(n5328) );
  SDFFX1 DFF_139_Q_reg ( .D(g33624), .SI(g1135), .SE(n8317), .CLK(n8731), .Q(
        g6395), .QN(n5396) );
  SDFFX1 DFF_141_Q_reg ( .D(g24337), .SI(g6395), .SE(n8317), .CLK(n8731), .Q(
        test_so10), .QN(n8236) );
  SDFFX1 DFF_142_Q_reg ( .D(g34911), .SI(test_si11), .SE(n8299), .CLK(n8713), 
        .Q(g554) );
  SDFFX1 DFF_143_Q_reg ( .D(g33963), .SI(g554), .SE(n8251), .CLK(n8665), .Q(
        g496) );
  SDFFX1 DFF_144_Q_reg ( .D(g34627), .SI(g496), .SE(n8251), .CLK(n8665), .Q(
        g3853), .QN(n5641) );
  SDFFX1 DFF_145_Q_reg ( .D(g29282), .SI(g3853), .SE(n8342), .CLK(n8756), .Q(
        g5134), .QN(n5807) );
  SDFFX1 DFF_146_Q_reg ( .D(g17320), .SI(g5134), .SE(n8347), .CLK(n8761), .Q(
        g17404) );
  SDFFX1 DFF_147_Q_reg ( .D(g25676), .SI(g17404), .SE(n8292), .CLK(n8706), .Q(
        g8344) );
  SDFFX1 DFF_148_Q_reg ( .D(g33013), .SI(g8344), .SE(n8292), .CLK(n8706), .Q(
        g2485), .QN(n5509) );
  SDFFX1 DFF_149_Q_reg ( .D(g32981), .SI(g2485), .SE(n8275), .CLK(n8689), .Q(
        g925), .QN(n5725) );
  SDFFX1 DFF_150_Q_reg ( .D(g34976), .SI(g925), .SE(n8249), .CLK(n8663), .Q(
        n9357), .QN(DFF_150_n1) );
  SDFFX1 DFF_151_Q_reg ( .D(g30483), .SI(n9357), .SE(n8249), .CLK(n8663), .Q(
        g5555), .QN(n8105) );
  SDFFX1 DFF_152_Q_reg ( .D(g14217), .SI(g5555), .SE(n8300), .CLK(n8714), .Q(
        g14096) );
  SDFFX1 DFF_153_Q_reg ( .D(g32994), .SI(g14096), .SE(n8300), .CLK(n8714), .Q(
        g1798), .QN(n5833) );
  SDFFX1 DFF_154_Q_reg ( .D(g28070), .SI(g1798), .SE(n8325), .CLK(n8739), .Q(
        test_so11), .QN(n8220) );
  SDFFX1 DFF_155_Q_reg ( .D(g34806), .SI(test_si12), .SE(n8264), .CLK(n8678), 
        .Q(g2941), .QN(n8172) );
  SDFFX1 DFF_156_Q_reg ( .D(g30453), .SI(g2941), .SE(n8264), .CLK(n8678), .Q(
        g3905) );
  SDFFX1 DFF_157_Q_reg ( .D(g33539), .SI(g3905), .SE(n8316), .CLK(n8730), .Q(
        g763), .QN(n5332) );
  SDFFX1 DFF_158_Q_reg ( .D(g30526), .SI(g763), .SE(n8352), .CLK(n8766), .Q(
        g6255), .QN(n8028) );
  SDFFX1 DFF_159_Q_reg ( .D(g26951), .SI(g6255), .SE(n8277), .CLK(n8691), .Q(
        g4375), .QN(n7680) );
  SDFFX1 DFF_160_Q_reg ( .D(g34035), .SI(g4375), .SE(n8302), .CLK(n8716), .Q(
        g4871), .QN(n5443) );
  SDFFX1 DFF_161_Q_reg ( .D(g34636), .SI(g4871), .SE(n8338), .CLK(n8752), .Q(
        g4722), .QN(n5345) );
  SDFFX1 DFF_162_Q_reg ( .D(g32978), .SI(g4722), .SE(n8283), .CLK(n8697), .Q(
        g590), .QN(n5472) );
  SDFFX1 DFF_163_Q_reg ( .D(g17722), .SI(g590), .SE(n8319), .CLK(n8733), .Q(
        g13099) );
  SDFFX1 DFF_164_Q_reg ( .D(g30348), .SI(g13099), .SE(n8263), .CLK(n8677), .Q(
        g1632), .QN(n5836) );
  SDFFX1 DFF_165_Q_reg ( .D(g24336), .SI(g1632), .SE(n8346), .CLK(n8760), .Q(
        g12238), .QN(n5438) );
  SDFFX1 DFF_166_Q_reg ( .D(g8215), .SI(g12238), .SE(n8272), .CLK(n8686), .Q(
        g3100), .QN(n7743) );
  SDFFX1 DFF_167_Q_reg ( .D(g24250), .SI(g3100), .SE(n8323), .CLK(n8737), .Q(
        test_so12) );
  SDFFX1 DFF_169_Q_reg ( .D(g29236), .SI(test_si13), .SE(n8323), .CLK(n8737), 
        .Q(g1437) );
  SDFFX1 DFF_170_Q_reg ( .D(g29298), .SI(g1437), .SE(n8256), .CLK(n8670), .Q(
        g6154), .QN(n5747) );
  SDFFX1 DFF_171_Q_reg ( .D(g10527), .SI(g6154), .SE(n8314), .CLK(n8728), .Q(
        g1579), .QN(n7809) );
  SDFFX1 DFF_172_Q_reg ( .D(g30499), .SI(g1579), .SE(n8249), .CLK(n8663), .Q(
        g5567), .QN(n8103) );
  SDFFX1 DFF_173_Q_reg ( .D(g33976), .SI(g5567), .SE(n8273), .CLK(n8687), .Q(
        g1752) );
  SDFFX1 DFF_174_Q_reg ( .D(g32996), .SI(g1752), .SE(n8316), .CLK(n8730), .Q(
        g1917), .QN(n8132) );
  SDFFX1 DFF_175_Q_reg ( .D(g30335), .SI(g1917), .SE(n8316), .CLK(n8730), .Q(
        g744), .QN(n5470) );
  SDFFX1 DFF_177_Q_reg ( .D(g34637), .SI(g744), .SE(n8338), .CLK(n8752), .Q(
        g4737), .QN(n5867) );
  SDFFX1 DFF_178_Q_reg ( .D(g25694), .SI(g4737), .SE(n8338), .CLK(n8752), .Q(
        g8132), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(g30528), .SI(g8132), .SE(n8297), .CLK(n8711), .Q(
        g6267) );
  SDFFX1 DFF_181_Q_reg ( .D(g16775), .SI(g6267), .SE(n8334), .CLK(n8748), .Q(
        g16659), .QN(n7962) );
  SDFFX1 DFF_182_Q_reg ( .D(g24251), .SI(g16659), .SE(n8323), .CLK(n8737), .Q(
        g1442), .QN(n8137) );
  SDFFX1 DFF_183_Q_reg ( .D(g30521), .SI(g1442), .SE(n8288), .CLK(n8702), .Q(
        test_so13) );
  SDFFX1 DFF_184_Q_reg ( .D(g26960), .SI(test_si14), .SE(n8290), .CLK(n8704), 
        .Q(g4477), .QN(n5849) );
  SDFFX1 DFF_185_Q_reg ( .D(g24239), .SI(g4477), .SE(n8330), .CLK(n8744), .Q(
        g10500) );
  SDFFX1 DFF_186_Q_reg ( .D(g34259), .SI(g10500), .SE(n8331), .CLK(n8745), .Q(
        g4643), .QN(n5382) );
  SDFFX1 DFF_187_Q_reg ( .D(g30474), .SI(g4643), .SE(n8253), .CLK(n8667), .Q(
        g5264) );
  SDFFX1 DFF_188_Q_reg ( .D(g12422), .SI(g5264), .SE(n8342), .CLK(n8756), .Q(
        g14779), .QN(n5703) );
  SDFFX1 DFF_189_Q_reg ( .D(g33016), .SI(g14779), .SE(n8293), .CLK(n8707), .Q(
        g2610), .QN(n8130) );
  SDFFX1 DFF_190_Q_reg ( .D(g34643), .SI(g2610), .SE(n8293), .CLK(n8707), .Q(
        g5160), .QN(n5498) );
  SDFFX1 DFF_192_Q_reg ( .D(g30510), .SI(g5160), .SE(n8337), .CLK(n8751), .Q(
        g5933) );
  SDFFX1 DFF_193_Q_reg ( .D(g29239), .SI(g5933), .SE(n8255), .CLK(n8669), .Q(
        g1454) );
  SDFFX1 DFF_194_Q_reg ( .D(g26897), .SI(g1454), .SE(n8343), .CLK(n8757), .Q(
        g753), .QN(n7771) );
  SDFFX1 DFF_195_Q_reg ( .D(g34729), .SI(g753), .SE(n8347), .CLK(n8761), .Q(
        g1296) );
  SDFFX1 DFF_196_Q_reg ( .D(g34625), .SI(g1296), .SE(n8347), .CLK(n8761), .Q(
        g3151), .QN(n5495) );
  SDFFX1 DFF_197_Q_reg ( .D(g34800), .SI(g3151), .SE(n8270), .CLK(n8684), .Q(
        test_so14) );
  SDFFX1 DFF_198_Q_reg ( .D(g24353), .SI(test_si15), .SE(n8266), .CLK(n8680), 
        .Q(g6727), .QN(n5531) );
  SDFFX1 DFF_199_Q_reg ( .D(g33029), .SI(g6727), .SE(n8315), .CLK(n8729), .Q(
        g3530), .QN(n5569) );
  SDFFX1 DFF_201_Q_reg ( .D(g33615), .SI(g3530), .SE(n8293), .CLK(n8707), .Q(
        g4104), .QN(n8001) );
  SDFFX1 DFF_202_Q_reg ( .D(g24253), .SI(g4104), .SE(n8293), .CLK(n8707), .Q(
        g1532), .QN(n7995) );
  SDFFX1 DFF_203_Q_reg ( .D(g24281), .SI(g1532), .SE(n8293), .CLK(n8707), .Q(
        g9251) );
  SDFFX1 DFF_204_Q_reg ( .D(g33997), .SI(g9251), .SE(n8312), .CLK(n8726), .Q(
        n9352) );
  SDFFX1 DFF_206_Q_reg ( .D(g34971), .SI(n9352), .SE(n8354), .CLK(n8768), .Q(
        n9351), .QN(DFF_206_n1) );
  SDFFX1 DFF_207_Q_reg ( .D(g34263), .SI(n9351), .SE(n8258), .CLK(n8672), .Q(
        g4754), .QN(n5877) );
  SDFFX1 DFF_208_Q_reg ( .D(g24237), .SI(g4754), .SE(n8332), .CLK(n8746), .Q(
        g1189), .QN(n5642) );
  SDFFX1 DFF_209_Q_reg ( .D(g33584), .SI(g1189), .SE(n8311), .CLK(n8725), .Q(
        g2287), .QN(n5353) );
  SDFFX1 DFF_210_Q_reg ( .D(g24280), .SI(g2287), .SE(n8311), .CLK(n8725), .Q(
        g4273), .QN(n5764) );
  SDFFX1 DFF_211_Q_reg ( .D(g26920), .SI(g4273), .SE(n8261), .CLK(n8675), .Q(
        g1389), .QN(n7845) );
  SDFFX1 DFF_212_Q_reg ( .D(g33548), .SI(g1389), .SE(n8322), .CLK(n8736), .Q(
        test_so15) );
  SDFFX1 DFF_213_Q_reg ( .D(g29296), .SI(test_si16), .SE(n8286), .CLK(n8700), 
        .Q(g5835), .QN(n5663) );
  SDFFX1 DFF_214_Q_reg ( .D(g30338), .SI(g5835), .SE(n8332), .CLK(n8746), .Q(
        g1171), .QN(n5363) );
  SDFFX1 DFF_215_Q_reg ( .D(g21895), .SI(g1171), .SE(n8332), .CLK(n8746), .Q(
        g4269), .QN(n5763) );
  SDFFX1 DFF_216_Q_reg ( .D(g33588), .SI(g4269), .SE(n8294), .CLK(n8708), .Q(
        g2399), .QN(n5762) );
  SDFFX1 DFF_218_Q_reg ( .D(g34041), .SI(g2399), .SE(n8294), .CLK(n8708), .Q(
        g4983), .QN(n5367) );
  SDFFX1 DFF_219_Q_reg ( .D(g30495), .SI(g4983), .SE(n8249), .CLK(n8663), .Q(
        g5611) );
  SDFFX1 DFF_220_Q_reg ( .D(g16744), .SI(g5611), .SE(n8297), .CLK(n8711), .Q(
        g16627), .QN(n7966) );
  SDFFX1 DFF_221_Q_reg ( .D(g29279), .SI(g16627), .SE(n8265), .CLK(n8679), .Q(
        g4572), .QN(n7770) );
  SDFFX1 DFF_222_Q_reg ( .D(g25655), .SI(g4572), .SE(n8270), .CLK(n8684), .Q(
        g3143), .QN(n5882) );
  SDFFX1 DFF_223_Q_reg ( .D(g34795), .SI(g3143), .SE(n8270), .CLK(n8684), .Q(
        g2898) );
  SDFFX1 DFF_224_Q_reg ( .D(g24269), .SI(g2898), .SE(n8321), .CLK(n8735), .Q(
        g3343), .QN(n7985) );
  SDFFX1 DFF_225_Q_reg ( .D(g30403), .SI(g3343), .SE(n8321), .CLK(n8735), .Q(
        g3235) );
  SDFFX1 DFF_226_Q_reg ( .D(g33042), .SI(g3235), .SE(n8321), .CLK(n8735), .Q(
        test_so16) );
  SDFFX1 DFF_227_Q_reg ( .D(g30419), .SI(test_si17), .SE(n8346), .CLK(n8760), 
        .Q(g3566) );
  SDFFX1 DFF_228_Q_reg ( .D(g34023), .SI(g3566), .SE(n8346), .CLK(n8760), .Q(
        n9348), .QN(DFF_228_n1) );
  SDFFX1 DFF_229_Q_reg ( .D(g28090), .SI(n9348), .SE(n8267), .CLK(n8681), .Q(
        g4961), .QN(n5770) );
  SDFFX1 DFF_231_Q_reg ( .D(g34642), .SI(g4961), .SE(n8267), .CLK(n8681), .Q(
        g4927), .QN(n5879) );
  SDFFX1 DFF_232_Q_reg ( .D(g30370), .SI(g4927), .SE(n8309), .CLK(n8723), .Q(
        g2259), .QN(n5419) );
  SDFFX1 DFF_233_Q_reg ( .D(g34448), .SI(g2259), .SE(n8280), .CLK(n8694), .Q(
        g2819), .QN(n5609) );
  SDFFX1 DFF_234_Q_reg ( .D(g26946), .SI(g2819), .SE(n8277), .CLK(n8691), .Q(
        g7257) );
  SDFFX1 DFF_235_Q_reg ( .D(g9617), .SI(g7257), .SE(n8277), .CLK(n8691), .Q(
        g5802), .QN(n7740) );
  SDFFX1 DFF_236_Q_reg ( .D(g34610), .SI(g5802), .SE(n8289), .CLK(n8703), .Q(
        g2852) );
  SDFFX1 DFF_237_Q_reg ( .D(g24209), .SI(g2852), .SE(n8312), .CLK(n8726), .Q(
        g417), .QN(n5358) );
  SDFFX1 DFF_238_Q_reg ( .D(g28047), .SI(g417), .SE(n8344), .CLK(n8758), .Q(
        g681) );
  SDFFX1 DFF_239_Q_reg ( .D(g24206), .SI(g681), .SE(n8257), .CLK(n8671), .Q(
        g437), .QN(n7834) );
  SDFFX1 DFF_240_Q_reg ( .D(g26891), .SI(g437), .SE(n8309), .CLK(n8723), .Q(
        test_so17), .QN(n8229) );
  SDFFX1 DFF_241_Q_reg ( .D(g30504), .SI(test_si18), .SE(n8351), .CLK(n8765), 
        .Q(g5901), .QN(n8101) );
  SDFFX1 DFF_242_Q_reg ( .D(g34798), .SI(g5901), .SE(n8270), .CLK(n8684), .Q(
        g2886), .QN(n8174) );
  SDFFX1 DFF_243_Q_reg ( .D(g25669), .SI(g2886), .SE(n8279), .CLK(n8693), .Q(
        g3494), .QN(n5889) );
  SDFFX1 DFF_244_Q_reg ( .D(g30480), .SI(g3494), .SE(n8279), .CLK(n8693), .Q(
        g5511), .QN(n5575) );
  SDFFX1 DFF_245_Q_reg ( .D(g33027), .SI(g5511), .SE(n8330), .CLK(n8744), .Q(
        g3518), .QN(n5645) );
  SDFFX1 DFF_246_Q_reg ( .D(g33972), .SI(g3518), .SE(n8346), .CLK(n8760), .Q(
        g1604) );
  SDFFX1 DFF_248_Q_reg ( .D(g25697), .SI(g1604), .SE(n8248), .CLK(n8662), .Q(
        g5092) );
  SDFFX1 DFF_249_Q_reg ( .D(g28099), .SI(g5092), .SE(n8288), .CLK(n8702), .Q(
        g4831) );
  SDFFX1 DFF_250_Q_reg ( .D(g26947), .SI(g4831), .SE(n8288), .CLK(n8702), .Q(
        g4382), .QN(n5714) );
  SDFFX1 DFF_251_Q_reg ( .D(g24350), .SI(g4382), .SE(n8346), .CLK(n8760), .Q(
        g6386), .QN(n7987) );
  SDFFX1 DFF_252_Q_reg ( .D(g24210), .SI(g6386), .SE(n8346), .CLK(n8760), .Q(
        g479) );
  SDFFX1 DFF_253_Q_reg ( .D(g30455), .SI(g479), .SE(n8265), .CLK(n8679), .Q(
        g3965) );
  SDFFX1 DFF_254_Q_reg ( .D(g28084), .SI(g3965), .SE(n8271), .CLK(n8685), .Q(
        test_so18), .QN(n8242) );
  SDFFX1 DFF_255_Q_reg ( .D(g33993), .SI(test_si19), .SE(n8291), .CLK(n8705), 
        .Q(g2008) );
  SDFFX1 DFF_256_Q_reg ( .D(g11678), .SI(g2008), .SE(n8291), .CLK(n8705), .Q(
        g736) );
  SDFFX1 DFF_257_Q_reg ( .D(g30444), .SI(g736), .SE(n8334), .CLK(n8748), .Q(
        g3933) );
  SDFFX1 DFF_258_Q_reg ( .D(g33537), .SI(g3933), .SE(n8276), .CLK(n8690), .Q(
        g222), .QN(n8187) );
  SDFFX1 DFF_259_Q_reg ( .D(g25650), .SI(g222), .SE(n8272), .CLK(n8686), .Q(
        g3050), .QN(n5998) );
  SDFFX1 DFF_261_Q_reg ( .D(g25625), .SI(g3050), .SE(n8295), .CLK(n8709), .Q(
        g1052), .QN(n8055) );
  SDFFX1 DFF_263_Q_reg ( .D(g17711), .SI(g1052), .SE(n8295), .CLK(n8709), .Q(
        g17580), .QN(n7960) );
  SDFFX1 DFF_264_Q_reg ( .D(g30366), .SI(g17580), .SE(n8279), .CLK(n8693), .Q(
        g2122), .QN(n5784) );
  SDFFX1 DFF_265_Q_reg ( .D(g33593), .SI(g2122), .SE(n8311), .CLK(n8725), .Q(
        g2465), .QN(n5523) );
  SDFFX1 DFF_267_Q_reg ( .D(g30502), .SI(g2465), .SE(n8335), .CLK(n8749), .Q(
        g5889), .QN(n8044) );
  SDFFX1 DFF_268_Q_reg ( .D(g33036), .SI(g5889), .SE(n8290), .CLK(n8704), .Q(
        g4495) );
  SDFFX1 DFF_269_Q_reg ( .D(g25595), .SI(g4495), .SE(n8290), .CLK(n8704), .Q(
        g8719), .QN(n7873) );
  SDFFX1 DFF_270_Q_reg ( .D(g34462), .SI(g8719), .SE(n8298), .CLK(n8712), .Q(
        test_so19), .QN(n8239) );
  SDFFX1 DFF_271_Q_reg ( .D(g33024), .SI(test_si20), .SE(n8272), .CLK(n8686), 
        .Q(g3179), .QN(n5390) );
  SDFFX1 DFF_272_Q_reg ( .D(g33552), .SI(g3179), .SE(n8274), .CLK(n8688), .Q(
        g1728), .QN(n5352) );
  SDFFX1 DFF_273_Q_reg ( .D(g34014), .SI(g1728), .SE(n8348), .CLK(n8762), .Q(
        g2433) );
  SDFFX1 DFF_274_Q_reg ( .D(g29273), .SI(g2433), .SE(n8278), .CLK(n8692), .Q(
        g3835), .QN(n5662) );
  SDFFX1 DFF_275_Q_reg ( .D(g25748), .SI(g3835), .SE(n8336), .CLK(n8750), .Q(
        g6187), .QN(n5453) );
  SDFFX1 DFF_276_Q_reg ( .D(g34638), .SI(g6187), .SE(n8336), .CLK(n8750), .Q(
        g4917), .QN(n5408) );
  SDFFX1 DFF_277_Q_reg ( .D(g30341), .SI(g4917), .SE(n8254), .CLK(n8668), .Q(
        g1070) );
  SDFFX1 DFF_278_Q_reg ( .D(g26899), .SI(g1070), .SE(n8324), .CLK(n8738), .Q(
        g822), .QN(n5422) );
  SDFFX1 DFF_279_Q_reg ( .D(g14673), .SI(g822), .SE(n8324), .CLK(n8738), .Q(
        g17715) );
  SDFFX1 DFF_280_Q_reg ( .D(g30336), .SI(g17715), .SE(n8275), .CLK(n8689), .Q(
        g914), .QN(n5560) );
  SDFFX1 DFF_281_Q_reg ( .D(g17639), .SI(g914), .SE(n8342), .CLK(n8756), .Q(
        g5339) );
  SDFFX1 DFF_282_Q_reg ( .D(g26940), .SI(g5339), .SE(n8353), .CLK(n8767), .Q(
        g4164), .QN(n8161) );
  SDFFX1 DFF_283_Q_reg ( .D(g25622), .SI(g4164), .SE(n8263), .CLK(n8677), .Q(
        test_so20), .QN(n8223) );
  SDFFX1 DFF_284_Q_reg ( .D(g34447), .SI(test_si21), .SE(n8280), .CLK(n8694), 
        .Q(g2807), .QN(n5379) );
  SDFFX1 DFF_286_Q_reg ( .D(g33613), .SI(g2807), .SE(n8267), .CLK(n8681), .Q(
        g4054), .QN(n5395) );
  SDFFX1 DFF_287_Q_reg ( .D(g25749), .SI(g4054), .SE(n8256), .CLK(n8670), .Q(
        g6191), .QN(n5888) );
  SDFFX1 DFF_288_Q_reg ( .D(g25704), .SI(g6191), .SE(n8256), .CLK(n8670), .Q(
        g5077), .QN(n5455) );
  SDFFX1 DFF_289_Q_reg ( .D(g33053), .SI(g5077), .SE(n8256), .CLK(n8670), .Q(
        g5523), .QN(n5647) );
  SDFFX1 DFF_290_Q_reg ( .D(g16722), .SI(g5523), .SE(n8332), .CLK(n8746), .Q(
        g3680) );
  SDFFX1 DFF_291_Q_reg ( .D(g30555), .SI(g3680), .SE(n8340), .CLK(n8754), .Q(
        g6637) );
  SDFFX1 DFF_292_Q_reg ( .D(g25601), .SI(g6637), .SE(n8344), .CLK(n8758), .Q(
        g174), .QN(n5402) );
  SDFFX1 DFF_293_Q_reg ( .D(g33971), .SI(g174), .SE(n8322), .CLK(n8736), .Q(
        g1682), .QN(n7789) );
  SDFFX1 DFF_294_Q_reg ( .D(g26892), .SI(g1682), .SE(n8322), .CLK(n8736), .Q(
        g355), .QN(n8136) );
  SDFFX1 DFF_295_Q_reg ( .D(g17400), .SI(g355), .SE(n8330), .CLK(n8744), .Q(
        g1087), .QN(n8157) );
  SDFFX1 DFF_296_Q_reg ( .D(g26915), .SI(g1087), .SE(n8294), .CLK(n8708), .Q(
        g1105), .QN(n5478) );
  SDFFX1 DFF_297_Q_reg ( .D(g33008), .SI(g1105), .SE(n8294), .CLK(n8708), .Q(
        test_so21), .QN(n8213) );
  SDFFX1 DFF_298_Q_reg ( .D(g30538), .SI(test_si22), .SE(n8297), .CLK(n8711), 
        .Q(g6307) );
  SDFFX1 DFF_299_Q_reg ( .D(g8344), .SI(g6307), .SE(n8297), .CLK(n8711), .Q(
        g3802), .QN(n7735) );
  SDFFX1 DFF_300_Q_reg ( .D(g25750), .SI(g3802), .SE(n8336), .CLK(n8750), .Q(
        g6159), .QN(n7791) );
  SDFFX1 DFF_301_Q_reg ( .D(g30369), .SI(g6159), .SE(n8309), .CLK(n8723), .Q(
        g2255), .QN(n5414) );
  SDFFX1 DFF_302_Q_reg ( .D(g34446), .SI(g2255), .SE(n8280), .CLK(n8694), .Q(
        g2815) );
  SDFFX1 DFF_303_Q_reg ( .D(g29230), .SI(g2815), .SE(n8275), .CLK(n8689), .Q(
        g911), .QN(n5559) );
  SDFFX1 DFF_304_Q_reg ( .D(n8193), .SI(g911), .SE(n8250), .CLK(n8664), .Q(g43), .QN(n7841) );
  SDFFX1 DFF_305_Q_reg ( .D(g13966), .SI(g43), .SE(n8334), .CLK(n8748), .Q(
        g16775), .QN(n7976) );
  SDFFX1 DFF_306_Q_reg ( .D(g33975), .SI(g16775), .SE(n8273), .CLK(n8687), .Q(
        g1748) );
  SDFFX1 DFF_307_Q_reg ( .D(g30497), .SI(g1748), .SE(n8259), .CLK(n8673), .Q(
        g5551), .QN(n8045) );
  SDFFX1 DFF_309_Q_reg ( .D(g30418), .SI(g5551), .SE(n8350), .CLK(n8764), .Q(
        g3558), .QN(n8025) );
  SDFFX1 DFF_310_Q_reg ( .D(g25721), .SI(g3558), .SE(n8353), .CLK(n8767), .Q(
        g5499), .QN(n5885) );
  SDFFX1 DFF_311_Q_reg ( .D(g34622), .SI(g5499), .SE(n8271), .CLK(n8685), .Q(
        test_so22), .QN(n8235) );
  SDFFX1 DFF_312_Q_reg ( .D(g30438), .SI(test_si23), .SE(n8264), .CLK(n8678), 
        .Q(g3901), .QN(n8109) );
  SDFFX1 DFF_313_Q_reg ( .D(g34266), .SI(g3901), .SE(n8266), .CLK(n8680), .Q(
        g4888), .QN(n5863) );
  SDFFX1 DFF_314_Q_reg ( .D(g30540), .SI(g4888), .SE(n8298), .CLK(n8712), .Q(
        g6251) );
  SDFFX1 DFF_315_Q_reg ( .D(g17760), .SI(g6251), .SE(n8342), .CLK(n8756), .Q(
        g17649), .QN(n7967) );
  SDFFX1 DFF_316_Q_reg ( .D(g32986), .SI(g17649), .SE(n8261), .CLK(n8675), .Q(
        g1373), .QN(n7849) );
  SDFFX1 DFF_317_Q_reg ( .D(g25648), .SI(g1373), .SE(n8272), .CLK(n8686), .Q(
        g8215) );
  SDFFX1 DFF_318_Q_reg ( .D(g33960), .SI(g8215), .SE(n8299), .CLK(n8713), .Q(
        g157), .QN(n5678) );
  SDFFX1 DFF_319_Q_reg ( .D(g34442), .SI(g157), .SE(n8281), .CLK(n8695), .Q(
        g2783) );
  SDFFX1 DFF_320_Q_reg ( .D(g8839), .SI(g2783), .SE(n8303), .CLK(n8717), .Q(
        g4281), .QN(n8190) );
  SDFFX1 DFF_321_Q_reg ( .D(g30421), .SI(g4281), .SE(n8306), .CLK(n8720), .Q(
        g3574) );
  SDFFX1 DFF_322_Q_reg ( .D(g33573), .SI(g3574), .SE(n8353), .CLK(n8767), .Q(
        g2112) );
  SDFFX1 DFF_323_Q_reg ( .D(g34730), .SI(g2112), .SE(n8353), .CLK(n8767), .Q(
        g1283), .QN(n5635) );
  SDFFX1 DFF_324_Q_reg ( .D(g24205), .SI(g1283), .SE(n8257), .CLK(n8671), .Q(
        test_so23) );
  SDFFX1 DFF_325_Q_reg ( .D(g10122_Tj), .SI(test_si24), .SE(n8306), .CLK(n8720), .Q(g4297), .QN(n7727) );
  SDFFX1 DFF_326_Q_reg ( .D(g12350), .SI(g4297), .SE(n8306), .CLK(n8720), .Q(
        g14738), .QN(n5698) );
  SDFFX1 DFF_327_Q_reg ( .D(g19357), .SI(g14738), .SE(n8307), .CLK(n8721), .Q(
        g13272), .QN(n7832) );
  SDFFX1 DFF_328_Q_reg ( .D(g32979), .SI(g13272), .SE(n8316), .CLK(n8730), .Q(
        g758), .QN(n5331) );
  SDFFX1 DFF_331_Q_reg ( .D(n322), .SI(g758), .SE(n8331), .CLK(n8745), .Q(
        g4639), .QN(n5727) );
  SDFFX1 DFF_332_Q_reg ( .D(g25763), .SI(g4639), .SE(n8259), .CLK(n8673), .Q(
        g6537), .QN(n5884) );
  SDFFX1 DFF_333_Q_reg ( .D(g30481), .SI(g6537), .SE(n8259), .CLK(n8673), .Q(
        g5543), .QN(n8046) );
  SDFFX1 DFF_334_Q_reg ( .D(g7946), .SI(g5543), .SE(n8262), .CLK(n8676), .Q(
        g8475), .QN(n7744) );
  SDFFX1 DFF_336_Q_reg ( .D(g30517), .SI(g8475), .SE(n8288), .CLK(n8702), .Q(
        g5961) );
  SDFFX1 DFF_337_Q_reg ( .D(g30539), .SI(g5961), .SE(n8344), .CLK(n8758), .Q(
        g6243), .QN(n8052) );
  SDFFX1 DFF_338_Q_reg ( .D(g34880), .SI(g6243), .SE(n8282), .CLK(n8696), .Q(
        n9340), .QN(n14519) );
  SDFFX1 DFF_339_Q_reg ( .D(g24242), .SI(n9340), .SE(n8275), .CLK(n8689), .Q(
        g12919), .QN(n5654) );
  SDFFX1 DFF_340_Q_reg ( .D(g30436), .SI(g12919), .SE(n8334), .CLK(n8748), .Q(
        test_so24) );
  SDFFX1 DFF_341_Q_reg ( .D(g29265), .SI(test_si25), .SE(n8295), .CLK(n8709), 
        .Q(g3476), .QN(n5786) );
  SDFFX1 DFF_342_Q_reg ( .D(g32990), .SI(g3476), .SE(n8296), .CLK(n8710), .Q(
        g1664) );
  SDFFX1 DFF_343_Q_reg ( .D(g24245), .SI(g1664), .SE(n8296), .CLK(n8710), .Q(
        g1246), .QN(n5756) );
  SDFFX1 DFF_345_Q_reg ( .D(g30553), .SI(g1246), .SE(n8329), .CLK(n8743), .Q(
        g6629) );
  SDFFX1 DFF_346_Q_reg ( .D(g26907), .SI(g6629), .SE(n8275), .CLK(n8689), .Q(
        g246), .QN(n6008) );
  SDFFX1 DFF_347_Q_reg ( .D(g24278), .SI(g246), .SE(n8347), .CLK(n8761), .Q(
        g4049), .QN(n7993) );
  SDFFX1 DFF_348_Q_reg ( .D(g26955), .SI(g4049), .SE(n8288), .CLK(n8702), .Q(
        g7260) );
  SDFFX1 DFF_349_Q_reg ( .D(g24282), .SI(g7260), .SE(n8289), .CLK(n8703), .Q(
        g2932), .QN(n8179) );
  SDFFX1 DFF_350_Q_reg ( .D(g29276), .SI(g2932), .SE(n8250), .CLK(n8664), .Q(
        g4575) );
  SDFFX1 DFF_351_Q_reg ( .D(g31894), .SI(g4575), .SE(n8250), .CLK(n8664), .Q(
        g4098), .QN(n5350) );
  SDFFX1 DFF_352_Q_reg ( .D(g33037), .SI(g4098), .SE(n8290), .CLK(n8704), .Q(
        g4498) );
  SDFFX1 DFF_353_Q_reg ( .D(g26894), .SI(g4498), .SE(n8323), .CLK(n8737), .Q(
        g528), .QN(n5327) );
  SDFFX1 DFF_355_Q_reg ( .D(g34977), .SI(g528), .SE(n8267), .CLK(n8681), .Q(
        test_so25), .QN(n5477) );
  SDFFX1 DFF_356_Q_reg ( .D(g25654), .SI(test_si26), .SE(n8327), .CLK(n8741), 
        .Q(g3139), .QN(n5447) );
  SDFFX1 DFF_357_Q_reg ( .D(g33962), .SI(g3139), .SE(n8275), .CLK(n8689), .Q(
        g29215) );
  SDFFX1 DFF_358_Q_reg ( .D(g34451), .SI(g29215), .SE(n8327), .CLK(n8741), .Q(
        g4584), .QN(n5539) );
  SDFFX1 DFF_359_Q_reg ( .D(g34250), .SI(g4584), .SE(n8276), .CLK(n8690), .Q(
        g142), .QN(n5724) );
  SDFFX1 DFF_360_Q_reg ( .D(g14597), .SI(g142), .SE(n8342), .CLK(n8756), .Q(
        g17639) );
  SDFFX1 DFF_361_Q_reg ( .D(g29295), .SI(g17639), .SE(n8285), .CLK(n8699), .Q(
        g5831), .QN(n5873) );
  SDFFX1 DFF_362_Q_reg ( .D(g26905), .SI(g5831), .SE(n8334), .CLK(n8748), .Q(
        g239), .QN(n7997) );
  SDFFX1 DFF_363_Q_reg ( .D(g25629), .SI(g239), .SE(n8284), .CLK(n8698), .Q(
        g1216), .QN(n5442) );
  SDFFX1 DFF_364_Q_reg ( .D(g34792), .SI(g1216), .SE(n8255), .CLK(n8669), .Q(
        g2848) );
  SDFFX1 DFF_366_Q_reg ( .D(g25703), .SI(g2848), .SE(n8317), .CLK(n8731), .Q(
        g5022), .QN(n7871) );
  SDFFX1 DFF_367_Q_reg ( .D(g14518), .SI(g5022), .SE(n8333), .CLK(n8747), .Q(
        g16955) );
  SDFFX1 DFF_368_Q_reg ( .D(g32983), .SI(g16955), .SE(n8263), .CLK(n8677), .Q(
        g1030), .QN(n7851) );
  SDFFX1 DFF_369_Q_reg ( .D(g16924), .SI(g1030), .SE(n8324), .CLK(n8738), .Q(
        test_so26) );
  SDFFX1 DFF_370_Q_reg ( .D(g30402), .SI(test_si27), .SE(n8328), .CLK(n8742), 
        .Q(g3231) );
  SDFFX1 DFF_371_Q_reg ( .D(g25757), .SI(g3231), .SE(n8313), .CLK(n8727), .Q(
        g9817), .QN(n7728) );
  SDFFX1 DFF_372_Q_reg ( .D(g17423), .SI(g9817), .SE(n8313), .CLK(n8727), .Q(
        g1430), .QN(n8155) );
  SDFFX1 DFF_373_Q_reg ( .D(g7245), .SI(g1430), .SE(n8309), .CLK(n8723), .Q(
        n9336), .QN(n14518) );
  SDFFX1 DFF_374_Q_reg ( .D(g33999), .SI(n9336), .SE(n8309), .CLK(n8723), .Q(
        g2241), .QN(n7788) );
  SDFFX1 DFF_375_Q_reg ( .D(g24262), .SI(g2241), .SE(n8313), .CLK(n8727), .Q(
        g1564), .QN(n8154) );
  SDFFX1 DFF_376_Q_reg ( .D(g25729), .SI(g1564), .SE(n8278), .CLK(n8692), .Q(
        g9680), .QN(n7739) );
  SDFFX1 DFF_377_Q_reg ( .D(test_so92), .SI(g9680), .SE(n8278), .CLK(n8692), 
        .Q(g6148), .QN(n7724) );
  SDFFX1 DFF_378_Q_reg ( .D(g30558), .SI(g6148), .SE(n8340), .CLK(n8754), .Q(
        g6649) );
  SDFFX1 DFF_379_Q_reg ( .D(n233), .SI(g6649), .SE(n8293), .CLK(n8707), .Q(
        g110) );
  SDFFX1 DFF_380_Q_reg ( .D(g14125), .SI(g110), .SE(n8300), .CLK(n8714), .Q(
        g14147) );
  SDFFX1 DFF_382_Q_reg ( .D(g26901), .SI(g14147), .SE(n8333), .CLK(n8747), .Q(
        g225), .QN(n5597) );
  SDFFX1 DFF_383_Q_reg ( .D(g26961), .SI(g225), .SE(n8333), .CLK(n8747), .Q(
        test_so27) );
  SDFFX1 DFF_384_Q_reg ( .D(g33039), .SI(test_si28), .SE(n8290), .CLK(n8704), 
        .Q(g4504) );
  SDFFX1 DFF_385_Q_reg ( .D(g33059), .SI(g4504), .SE(n8335), .CLK(n8749), .Q(
        g5873), .QN(n5388) );
  SDFFX1 DFF_386_Q_reg ( .D(g31899), .SI(g5873), .SE(n8317), .CLK(n8731), .Q(
        g5037), .QN(n5611) );
  SDFFX1 DFF_387_Q_reg ( .D(g33007), .SI(g5037), .SE(n8318), .CLK(n8732), .Q(
        g2319), .QN(n5375) );
  SDFFX1 DFF_388_Q_reg ( .D(g25720), .SI(g2319), .SE(n8353), .CLK(n8767), .Q(
        g5495), .QN(n5446) );
  SDFFX1 DFF_389_Q_reg ( .D(g21891), .SI(g5495), .SE(n8253), .CLK(n8667), .Q(
        g11770) );
  SDFFX1 DFF_390_Q_reg ( .D(g30462), .SI(g11770), .SE(n8253), .CLK(n8667), .Q(
        g5208), .QN(n8004) );
  SDFFX1 DFF_392_Q_reg ( .D(g30487), .SI(g5208), .SE(n8249), .CLK(n8663), .Q(
        g5579) );
  SDFFX1 DFF_393_Q_reg ( .D(g33058), .SI(g5579), .SE(n8335), .CLK(n8749), .Q(
        g5869), .QN(n5649) );
  SDFFX1 DFF_395_Q_reg ( .D(g24261), .SI(g5869), .SE(n8335), .CLK(n8749), .Q(
        g1589), .QN(n5755) );
  SDFFX1 DFF_396_Q_reg ( .D(g25730), .SI(g1589), .SE(n8278), .CLK(n8692), .Q(
        g5752), .QN(n5996) );
  SDFFX1 DFF_397_Q_reg ( .D(g30531), .SI(g5752), .SE(n8336), .CLK(n8750), .Q(
        g6279) );
  SDFFX1 DFF_398_Q_reg ( .D(g30506), .SI(g6279), .SE(n8337), .CLK(n8751), .Q(
        test_so28) );
  SDFFX1 DFF_399_Q_reg ( .D(g34804), .SI(test_si29), .SE(n8248), .CLK(n8662), 
        .Q(g2975), .QN(n5750) );
  SDFFX1 DFF_400_Q_reg ( .D(g25747), .SI(g2975), .SE(n8256), .CLK(n8670), .Q(
        g6167), .QN(n5430) );
  SDFFX1 DFF_401_Q_reg ( .D(g11418), .SI(g6167), .SE(n8334), .CLK(n8748), .Q(
        g13966), .QN(n5701) );
  SDFFX1 DFF_402_Q_reg ( .D(g33601), .SI(g13966), .SE(n8348), .CLK(n8762), .Q(
        g2599), .QN(n5524) );
  SDFFX1 DFF_403_Q_reg ( .D(g26922), .SI(g2599), .SE(n8255), .CLK(n8669), .Q(
        g1448), .QN(n5343) );
  SDFFX1 DFF_404_Q_reg ( .D(g14096), .SI(g1448), .SE(n8300), .CLK(n8714), .Q(
        g14125) );
  SDFFX1 DFF_406_Q_reg ( .D(g29250), .SI(g14125), .SE(n8318), .CLK(n8732), .Q(
        g2370) );
  SDFFX1 DFF_407_Q_reg ( .D(g30459), .SI(g2370), .SE(n8318), .CLK(n8732), .Q(
        g5164), .QN(n5570) );
  SDFFX1 DFF_408_Q_reg ( .D(g8475), .SI(g5164), .SE(n8318), .CLK(n8732), .Q(
        g1333), .QN(n5616) );
  SDFFX1 DFF_409_Q_reg ( .D(g33534), .SI(g1333), .SE(n8299), .CLK(n8713), .Q(
        g153), .QN(n5677) );
  SDFFX1 DFF_410_Q_reg ( .D(g30543), .SI(g153), .SE(n8326), .CLK(n8740), .Q(
        g6549), .QN(n5571) );
  SDFFX1 DFF_411_Q_reg ( .D(g29275), .SI(g6549), .SE(n8326), .CLK(n8740), .Q(
        g4087), .QN(n5480) );
  SDFFX1 DFF_412_Q_reg ( .D(g34030), .SI(g4087), .SE(n8298), .CLK(n8712), .Q(
        test_so29), .QN(n8215) );
  SDFFX1 DFF_413_Q_reg ( .D(g34980), .SI(test_si30), .SE(n8270), .CLK(n8684), 
        .Q(g2984), .QN(n5842) );
  SDFFX1 DFF_414_Q_reg ( .D(g30451), .SI(g2984), .SE(n8265), .CLK(n8679), .Q(
        g3961) );
  SDFFX1 DFF_416_Q_reg ( .D(g25627), .SI(g3961), .SE(n8332), .CLK(n8746), .Q(
        g962), .QN(n5630) );
  SDFFX1 DFF_417_Q_reg ( .D(g34657), .SI(g962), .SE(n8258), .CLK(n8672), .Q(
        g101) );
  SDFFX1 DFF_418_Q_reg ( .D(g8870), .SI(g101), .SE(n8258), .CLK(n8672), .Q(
        g8918), .QN(n14524) );
  SDFFX1 DFF_419_Q_reg ( .D(g30552), .SI(g8918), .SE(n8258), .CLK(n8672), .Q(
        g6625) );
  SDFFX1 DFF_420_Q_reg ( .D(g34979), .SI(g6625), .SE(n8262), .CLK(n8676), .Q(
        n9332), .QN(DFF_420_n1) );
  SDFFX1 DFF_421_Q_reg ( .D(g30337), .SI(n9332), .SE(n8262), .CLK(n8676), .Q(
        g1018), .QN(n7850) );
  SDFFX1 DFF_422_Q_reg ( .D(g24254), .SI(g1018), .SE(n8347), .CLK(n8761), .Q(
        g17320) );
  SDFFX1 DFF_423_Q_reg ( .D(g24277), .SI(g17320), .SE(n8347), .CLK(n8761), .Q(
        g4045), .QN(n7994) );
  SDFFX1 DFF_424_Q_reg ( .D(g29237), .SI(g4045), .SE(n8307), .CLK(n8721), .Q(
        g1467) );
  SDFFX1 DFF_425_Q_reg ( .D(g30378), .SI(g1467), .SE(n8280), .CLK(n8694), .Q(
        g2461), .QN(n5840) );
  SDFFX1 DFF_428_Q_reg ( .D(g33019), .SI(g2461), .SE(n8281), .CLK(n8695), .Q(
        test_so30), .QN(n5300) );
  SDFFX1 DFF_429_Q_reg ( .D(g33623), .SI(test_si31), .SE(n8331), .CLK(n8745), 
        .Q(g5990), .QN(n5589) );
  SDFFX1 DFF_431_Q_reg ( .D(g29235), .SI(g5990), .SE(n8314), .CLK(n8728), .Q(
        g1256), .QN(n5558) );
  SDFFX1 DFF_432_Q_reg ( .D(g31902), .SI(g1256), .SE(n8250), .CLK(n8664), .Q(
        g5029), .QN(n5601) );
  SDFFX1 DFF_433_Q_reg ( .D(g29306), .SI(g5029), .SE(n8292), .CLK(n8706), .Q(
        g6519), .QN(n5806) );
  SDFFX1 DFF_434_Q_reg ( .D(g25689), .SI(g6519), .SE(n8292), .CLK(n8706), .Q(
        g4169), .QN(n5729) );
  SDFFX1 DFF_435_Q_reg ( .D(g33978), .SI(g4169), .SE(n8274), .CLK(n8688), .Q(
        g1816), .QN(n7708) );
  SDFFX1 DFF_436_Q_reg ( .D(g26970), .SI(g1816), .SE(n8274), .CLK(n8688), .Q(
        g4369), .QN(n7999) );
  SDFFX1 DFF_439_Q_reg ( .D(g29278), .SI(g4369), .SE(n8265), .CLK(n8679), .Q(
        g4578) );
  SDFFX1 DFF_440_Q_reg ( .D(g34253), .SI(g4578), .SE(n8266), .CLK(n8680), .Q(
        g4459), .QN(n5765) );
  SDFFX1 DFF_441_Q_reg ( .D(g29272), .SI(g4459), .SE(n8278), .CLK(n8692), .Q(
        g3831), .QN(n5872) );
  SDFFX1 DFF_442_Q_reg ( .D(g33595), .SI(g3831), .SE(n8308), .CLK(n8722), .Q(
        g2514), .QN(n7750) );
  SDFFX1 DFF_443_Q_reg ( .D(g33610), .SI(g2514), .SE(n8295), .CLK(n8709), .Q(
        g3288), .QN(n5400) );
  SDFFX1 DFF_444_Q_reg ( .D(g33589), .SI(g3288), .SE(n8352), .CLK(n8766), .Q(
        test_so31) );
  SDFFX1 DFF_445_Q_reg ( .D(g34605), .SI(test_si32), .SE(n8283), .CLK(n8697), 
        .Q(g2145), .QN(n5307) );
  SDFFX1 DFF_446_Q_reg ( .D(g30350), .SI(g2145), .SE(n8296), .CLK(n8710), .Q(
        g1700), .QN(n5417) );
  SDFFX1 DFF_447_Q_reg ( .D(g25611), .SI(g1700), .SE(n8323), .CLK(n8737), .Q(
        g513), .QN(n5548) );
  SDFFX1 DFF_448_Q_reg ( .D(test_so9), .SI(g513), .SE(n8280), .CLK(n8694), .Q(
        g2841), .QN(n5963) );
  SDFFX1 DFF_449_Q_reg ( .D(g33619), .SI(g2841), .SE(n8269), .CLK(n8683), .Q(
        g5297), .QN(n5588) );
  SDFFX1 DFF_451_Q_reg ( .D(g34022), .SI(g5297), .SE(n8302), .CLK(n8716), .Q(
        g2763), .QN(n7689) );
  SDFFX1 DFF_452_Q_reg ( .D(g34033), .SI(g2763), .SE(n8298), .CLK(n8712), .Q(
        g4793), .QN(n5368) );
  SDFFX1 DFF_453_Q_reg ( .D(g34726), .SI(g4793), .SE(n8332), .CLK(n8746), .Q(
        g952) );
  SDFFX1 DFF_454_Q_reg ( .D(g31870), .SI(g952), .SE(n8314), .CLK(n8728), .Q(
        g1263), .QN(n5674) );
  SDFFX1 DFF_455_Q_reg ( .D(g33985), .SI(g1263), .SE(n8286), .CLK(n8700), .Q(
        g1950), .QN(n7787) );
  SDFFX1 DFF_456_Q_reg ( .D(g29283), .SI(g1950), .SE(n8268), .CLK(n8682), .Q(
        g5138), .QN(n5871) );
  SDFFX1 DFF_457_Q_reg ( .D(g34003), .SI(g5138), .SE(n8287), .CLK(n8701), .Q(
        g2307) );
  SDFFX1 DFF_458_Q_reg ( .D(g9497), .SI(g2307), .SE(n8287), .CLK(n8701), .Q(
        test_so32) );
  SDFFX1 DFF_460_Q_reg ( .D(g25677), .SI(test_si33), .SE(n8255), .CLK(n8669), 
        .Q(g8398), .QN(n7734) );
  SDFFX1 DFF_461_Q_reg ( .D(g34463), .SI(g8398), .SE(n8255), .CLK(n8669), .Q(
        g4664) );
  SDFFX1 DFF_462_Q_reg ( .D(g33006), .SI(g4664), .SE(n8310), .CLK(n8724), .Q(
        g2223) );
  SDFFX1 DFF_463_Q_reg ( .D(g29292), .SI(g2223), .SE(n8285), .CLK(n8699), .Q(
        g5808), .QN(n5749) );
  SDFFX1 DFF_464_Q_reg ( .D(g30557), .SI(g5808), .SE(n8329), .CLK(n8743), .Q(
        g6645) );
  SDFFX1 DFF_465_Q_reg ( .D(g33989), .SI(g6645), .SE(n8292), .CLK(n8706), .Q(
        g2016) );
  SDFFX1 DFF_467_Q_reg ( .D(g33033), .SI(g2016), .SE(n8292), .CLK(n8706), .Q(
        g3873), .QN(n5387) );
  SDFFX1 DFF_468_Q_reg ( .D(g11388), .SI(g3873), .SE(n8296), .CLK(n8710), .Q(
        g13926), .QN(n5699) );
  SDFFX1 DFF_469_Q_reg ( .D(g34005), .SI(g13926), .SE(n8287), .CLK(n8701), .Q(
        g2315), .QN(n5802) );
  SDFFX1 DFF_470_Q_reg ( .D(g26932), .SI(g2315), .SE(n8288), .CLK(n8702), .Q(
        g2811) );
  SDFFX1 DFF_471_Q_reg ( .D(g30516), .SI(g2811), .SE(n8288), .CLK(n8702), .Q(
        g5957) );
  SDFFX1 DFF_472_Q_reg ( .D(g33575), .SI(g5957), .SE(n8284), .CLK(n8698), .Q(
        g2047) );
  SDFFX1 DFF_473_Q_reg ( .D(g33032), .SI(g2047), .SE(n8330), .CLK(n8744), .Q(
        test_so33), .QN(n8209) );
  SDFFX1 DFF_474_Q_reg ( .D(g14779), .SI(test_si34), .SE(n8342), .CLK(n8756), 
        .Q(g17760), .QN(n7982) );
  SDFFX1 DFF_476_Q_reg ( .D(g30486), .SI(g17760), .SE(n8260), .CLK(n8674), .Q(
        g5575) );
  SDFFX1 DFF_477_Q_reg ( .D(g34974), .SI(g5575), .SE(n8255), .CLK(n8669), .Q(
        n9327), .QN(DFF_477_n1) );
  SDFFX1 DFF_478_Q_reg ( .D(g25678), .SI(n9327), .SE(n8255), .CLK(n8669), .Q(
        g3752), .QN(n5994) );
  SDFFX1 DFF_479_Q_reg ( .D(g30440), .SI(g3752), .SE(n8334), .CLK(n8748), .Q(
        g3917) );
  SDFFX1 DFF_480_Q_reg ( .D(test_so86), .SI(g3917), .SE(n8303), .CLK(n8717), 
        .Q(g8783), .QN(n14526) );
  SDFFX1 DFF_481_Q_reg ( .D(g12923), .SI(g8783), .SE(n8303), .CLK(n8717), .Q(
        g1585), .QN(n5757) );
  SDFFX1 DFF_482_Q_reg ( .D(g26949), .SI(g1585), .SE(n8343), .CLK(n8757), .Q(
        g4388) );
  SDFFX1 DFF_483_Q_reg ( .D(g30530), .SI(g4388), .SE(n8352), .CLK(n8766), .Q(
        g6275) );
  SDFFX1 DFF_484_Q_reg ( .D(g30542), .SI(g6275), .SE(n8297), .CLK(n8711), .Q(
        g6311) );
  SDFFX1 DFF_485_Q_reg ( .D(g8915), .SI(g6311), .SE(n8297), .CLK(n8711), .Q(
        g8916) );
  SDFFX1 DFF_486_Q_reg ( .D(g25624), .SI(g8916), .SE(n8263), .CLK(n8677), .Q(
        g1041), .QN(n7692) );
  SDFFX1 DFF_487_Q_reg ( .D(g30383), .SI(g1041), .SE(n8293), .CLK(n8707), .Q(
        test_so34), .QN(n8243) );
  SDFFX1 DFF_488_Q_reg ( .D(g33597), .SI(test_si35), .SE(n8349), .CLK(n8763), 
        .Q(g2537) );
  SDFFX1 DFF_489_Q_reg ( .D(g34598), .SI(g2537), .SE(n8277), .CLK(n8691), .Q(
        g29221), .QN(g23612) );
  SDFFX1 DFF_490_Q_reg ( .D(g26957), .SI(g29221), .SE(n8277), .CLK(n8691), .Q(
        g4430), .QN(n7772) );
  SDFFX1 DFF_491_Q_reg ( .D(g26967), .SI(g4430), .SE(n8342), .CLK(n8756), .Q(
        n9325) );
  SDFFX1 DFF_493_Q_reg ( .D(g28102), .SI(n9325), .SE(n8297), .CLK(n8711), .Q(
        g4826) );
  SDFFX1 DFF_494_Q_reg ( .D(g30524), .SI(g4826), .SE(n8297), .CLK(n8711), .Q(
        g6239), .QN(n7895) );
  SDFFX1 DFF_496_Q_reg ( .D(g26903), .SI(g6239), .SE(n8333), .CLK(n8747), .Q(
        g232), .QN(n7996) );
  SDFFX1 DFF_497_Q_reg ( .D(g30475), .SI(g232), .SE(n8254), .CLK(n8668), .Q(
        g5268) );
  SDFFX1 DFF_498_Q_reg ( .D(g34647), .SI(g5268), .SE(n8254), .CLK(n8668), .Q(
        g6545), .QN(n5497) );
  SDFFX1 DFF_499_Q_reg ( .D(g30377), .SI(g6545), .SE(n8273), .CLK(n8687), .Q(
        n9324) );
  SDFFX1 DFF_500_Q_reg ( .D(g33553), .SI(n9324), .SE(n8273), .CLK(n8687), .Q(
        g1772), .QN(n5504) );
  SDFFX1 DFF_502_Q_reg ( .D(g31903), .SI(g1772), .SE(n8251), .CLK(n8665), .Q(
        g5052), .QN(n5607) );
  SDFFX1 DFF_503_Q_reg ( .D(g25715), .SI(g5052), .SE(n8251), .CLK(n8665), .Q(
        test_so35), .QN(n7732) );
  SDFFX1 DFF_504_Q_reg ( .D(g33984), .SI(test_si36), .SE(n8287), .CLK(n8701), 
        .Q(g1890), .QN(n5799) );
  SDFFX1 DFF_505_Q_reg ( .D(g33602), .SI(g1890), .SE(n8348), .CLK(n8762), .Q(
        g2629), .QN(n5521) );
  SDFFX1 DFF_506_Q_reg ( .D(g28045), .SI(g2629), .SE(n8282), .CLK(n8696), .Q(
        g572), .QN(n5337) );
  SDFFX1 DFF_507_Q_reg ( .D(g34603), .SI(g572), .SE(n8283), .CLK(n8697), .Q(
        g2130), .QN(n5487) );
  SDFFX1 DFF_508_Q_reg ( .D(g33035), .SI(g2130), .SE(n8292), .CLK(n8706), .Q(
        g4108), .QN(n5715) );
  SDFFX1 DFF_509_Q_reg ( .D(g9251), .SI(g4108), .SE(n8293), .CLK(n8707), .Q(
        g4308) );
  SDFFX1 DFF_510_Q_reg ( .D(g24208), .SI(g4308), .SE(n8257), .CLK(n8671), .Q(
        g475) );
  SDFFX1 DFF_511_Q_reg ( .D(g8416), .SI(g475), .SE(n8332), .CLK(n8746), .Q(
        g990), .QN(n5622) );
  SDFFX1 DFF_512_Q_reg ( .D(g34971), .SI(g990), .SE(n8262), .CLK(n8676), .Q(
        g31), .QN(n5469) );
  SDFFX1 DFF_514_Q_reg ( .D(g34970), .SI(g31), .SE(n8251), .CLK(n8665), .Q(
        n9322), .QN(DFF_514_n1) );
  SDFFX1 DFF_515_Q_reg ( .D(g24213), .SI(n9322), .SE(n8251), .CLK(n8665), .Q(
        g12184) );
  SDFFX1 DFF_517_Q_reg ( .D(g33614), .SI(g12184), .SE(n8251), .CLK(n8665), .Q(
        g3990), .QN(n5594) );
  SDFFX1 DFF_519_Q_reg ( .D(g33060), .SI(g3990), .SE(n8335), .CLK(n8749), .Q(
        test_so36), .QN(n8217) );
  SDFFX1 DFF_520_Q_reg ( .D(g30362), .SI(test_si37), .SE(n8272), .CLK(n8686), 
        .Q(g1992) );
  SDFFX1 DFF_522_Q_reg ( .D(g33023), .SI(g1992), .SE(n8272), .CLK(n8686), .Q(
        g3171), .QN(n5603) );
  SDFFX1 DFF_524_Q_reg ( .D(g26898), .SI(g3171), .SE(n8325), .CLK(n8739), .Q(
        g812), .QN(n5733) );
  SDFFX1 DFF_525_Q_reg ( .D(g25618), .SI(g812), .SE(n8325), .CLK(n8739), .Q(
        g832), .QN(n8153) );
  SDFFX1 DFF_526_Q_reg ( .D(g30518), .SI(g832), .SE(n8325), .CLK(n8739), .Q(
        g5897), .QN(n8043) );
  SDFFX1 DFF_527_Q_reg ( .D(g25688), .SI(g5897), .SE(n8325), .CLK(n8739), .Q(
        g25689) );
  SDFFX1 DFF_528_Q_reg ( .D(g4570), .SI(g25689), .SE(n8338), .CLK(n8752), .Q(
        g4571) );
  SDFFX1 DFF_529_Q_reg ( .D(g11349), .SI(g4571), .SE(n8338), .CLK(n8752), .Q(
        g13895), .QN(n5702) );
  SDFFX1 DFF_530_Q_reg ( .D(g26959), .SI(g13895), .SE(n8301), .CLK(n8715), .Q(
        g4455) );
  SDFFX1 DFF_531_Q_reg ( .D(g34801), .SI(g4455), .SE(n8264), .CLK(n8678), .Q(
        g2902), .QN(n7818) );
  SDFFX1 DFF_532_Q_reg ( .D(g26884), .SI(g2902), .SE(n8309), .CLK(n8723), .Q(
        g333), .QN(n8135) );
  SDFFX1 DFF_533_Q_reg ( .D(g25600), .SI(g333), .SE(n8344), .CLK(n8758), .Q(
        g168), .QN(n5606) );
  SDFFX1 DFF_534_Q_reg ( .D(g26933), .SI(g168), .SE(n8280), .CLK(n8694), .Q(
        test_so37) );
  SDFFX1 DFF_535_Q_reg ( .D(g28066), .SI(test_si38), .SE(n8352), .CLK(n8766), 
        .Q(g3684) );
  SDFFX1 DFF_536_Q_reg ( .D(g33612), .SI(g3684), .SE(n8279), .CLK(n8693), .Q(
        g3639), .QN(n5591) );
  SDFFX1 DFF_537_Q_reg ( .D(g17787), .SI(g3639), .SE(n8342), .CLK(n8756), .Q(
        g14597) );
  SDFFX1 DFF_538_Q_reg ( .D(g24268), .SI(g14597), .SE(n8321), .CLK(n8735), .Q(
        g3338), .QN(n5527) );
  SDFFX1 DFF_539_Q_reg ( .D(g25716), .SI(g3338), .SE(n8251), .CLK(n8665), .Q(
        g5406), .QN(n5992) );
  SDFFX1 DFF_541_Q_reg ( .D(g26906), .SI(g5406), .SE(n8251), .CLK(n8665), .Q(
        g269), .QN(n7870) );
  SDFFX1 DFF_542_Q_reg ( .D(g24203), .SI(g269), .SE(n8258), .CLK(n8672), .Q(
        g401), .QN(n7813) );
  SDFFX1 DFF_543_Q_reg ( .D(g24346), .SI(g401), .SE(n8258), .CLK(n8672), .Q(
        g6040), .QN(n7988) );
  SDFFX1 DFF_544_Q_reg ( .D(g24207), .SI(g6040), .SE(n8257), .CLK(n8671), .Q(
        g441), .QN(n7864) );
  SDFFX1 DFF_545_Q_reg ( .D(g25701), .SI(g441), .SE(n8317), .CLK(n8731), .Q(
        g9553), .QN(n5690) );
  SDFFX1 DFF_546_Q_reg ( .D(g29269), .SI(g9553), .SE(n8290), .CLK(n8704), .Q(
        g3808), .QN(n5745) );
  SDFFX1 DFF_547_Q_reg ( .D(g34976), .SI(g3808), .SE(n8290), .CLK(n8704), .Q(
        g9), .QN(n5468) );
  SDFFX1 DFF_549_Q_reg ( .D(g34255), .SI(g9), .SE(n8290), .CLK(n8704), .Q(
        test_so38), .QN(n8222) );
  SDFFX1 DFF_550_Q_reg ( .D(g30450), .SI(test_si39), .SE(n8265), .CLK(n8679), 
        .Q(g3957) );
  SDFFX1 DFF_551_Q_reg ( .D(g30456), .SI(g3957), .SE(n8326), .CLK(n8740), .Q(
        g4093), .QN(n5340) );
  SDFFX1 DFF_552_Q_reg ( .D(g32991), .SI(g4093), .SE(n8326), .CLK(n8740), .Q(
        g1760), .QN(n5602) );
  SDFFX1 DFF_554_Q_reg ( .D(g24348), .SI(g1760), .SE(n8342), .CLK(n8756), .Q(
        g12422), .QN(n5437) );
  SDFFX1 DFF_555_Q_reg ( .D(g34249), .SI(g12422), .SE(n8299), .CLK(n8713), .Q(
        g160), .QN(n5843) );
  SDFFX1 DFF_558_Q_reg ( .D(g30371), .SI(g160), .SE(n8349), .CLK(n8763), .Q(
        g2279), .QN(n5778) );
  SDFFX1 DFF_559_Q_reg ( .D(g29268), .SI(g2279), .SE(n8349), .CLK(n8763), .Q(
        g3498) );
  SDFFX1 DFF_560_Q_reg ( .D(g29224), .SI(g3498), .SE(n8283), .CLK(n8697), .Q(
        g586), .QN(n5336) );
  SDFFX1 DFF_561_Q_reg ( .D(g14189), .SI(g586), .SE(n8300), .CLK(n8714), .Q(
        g14201) );
  SDFFX1 DFF_562_Q_reg ( .D(g33017), .SI(g14201), .SE(n8294), .CLK(n8708), .Q(
        g2619), .QN(n5508) );
  SDFFX1 DFF_563_Q_reg ( .D(g30339), .SI(g2619), .SE(n8294), .CLK(n8708), .Q(
        g1183), .QN(n5599) );
  SDFFX1 DFF_564_Q_reg ( .D(g33967), .SI(g1183), .SE(n8315), .CLK(n8729), .Q(
        g1608) );
  SDFFX1 DFF_565_Q_reg ( .D(g8784), .SI(g1608), .SE(n8315), .CLK(n8729), .Q(
        test_so39) );
  SDFFX1 DFF_566_Q_reg ( .D(g17519), .SI(test_si40), .SE(n8341), .CLK(n8755), 
        .Q(g17577) );
  SDFFX1 DFF_567_Q_reg ( .D(g33559), .SI(g17577), .SE(n8345), .CLK(n8759), .Q(
        g1779) );
  SDFFX1 DFF_568_Q_reg ( .D(g29255), .SI(g1779), .SE(n8353), .CLK(n8767), .Q(
        g2652), .QN(n7919) );
  SDFFX1 DFF_570_Q_reg ( .D(g30368), .SI(g2652), .SE(n8261), .CLK(n8675), .Q(
        g2193), .QN(n5839) );
  SDFFX1 DFF_571_Q_reg ( .D(g30375), .SI(g2193), .SE(n8294), .CLK(n8708), .Q(
        g2393), .QN(n5421) );
  SDFFX1 DFF_573_Q_reg ( .D(g28052), .SI(g2393), .SE(n8344), .CLK(n8758), .Q(
        g661) );
  SDFFX1 DFF_574_Q_reg ( .D(g28089), .SI(g661), .SE(n8279), .CLK(n8693), .Q(
        g4950), .QN(n5772) );
  SDFFX1 DFF_575_Q_reg ( .D(g33055), .SI(g4950), .SE(n8341), .CLK(n8755), .Q(
        g5535), .QN(n5566) );
  SDFFX1 DFF_576_Q_reg ( .D(g30392), .SI(g5535), .SE(n8261), .CLK(n8675), .Q(
        g2834), .QN(g23652) );
  SDFFX1 DFF_577_Q_reg ( .D(g30343), .SI(g2834), .SE(n8261), .CLK(n8675), .Q(
        g1361), .QN(n7848) );
  SDFFX1 DFF_579_Q_reg ( .D(g30523), .SI(g1361), .SE(n8336), .CLK(n8750), .Q(
        g6235), .QN(n8053) );
  SDFFX1 DFF_580_Q_reg ( .D(g24233), .SI(g6235), .SE(n8294), .CLK(n8708), .Q(
        g1146), .QN(n5851) );
  SDFFX1 DFF_581_Q_reg ( .D(g33018), .SI(g1146), .SE(n8294), .CLK(n8708), .Q(
        test_so40) );
  SDFFX1 DFF_582_Q_reg ( .D(g32976), .SI(test_si41), .SE(n8299), .CLK(n8713), 
        .Q(g150), .QN(n5676) );
  SDFFX1 DFF_583_Q_reg ( .D(g30349), .SI(g150), .SE(n8296), .CLK(n8710), .Q(
        g1696), .QN(n5628) );
  SDFFX1 DFF_584_Q_reg ( .D(g33067), .SI(g1696), .SE(n8328), .CLK(n8742), .Q(
        g6555), .QN(n8141) );
  SDFFX1 DFF_585_Q_reg ( .D(g26900), .SI(g6555), .SE(n8300), .CLK(n8714), .Q(
        g14189) );
  SDFFX1 DFF_587_Q_reg ( .D(g33034), .SI(g14189), .SE(n8292), .CLK(n8706), .Q(
        g3881), .QN(n5564) );
  SDFFX1 DFF_588_Q_reg ( .D(g30551), .SI(g3881), .SE(n8340), .CLK(n8754), .Q(
        g6621) );
  SDFFX1 DFF_589_Q_reg ( .D(g25667), .SI(g6621), .SE(n8295), .CLK(n8709), .Q(
        g3470), .QN(n5424) );
  SDFFX1 DFF_590_Q_reg ( .D(g30452), .SI(g3470), .SE(n8334), .CLK(n8748), .Q(
        g3897), .QN(n8047) );
  SDFFX1 DFF_593_Q_reg ( .D(g34719), .SI(g518), .SE(n8276), .CLK(n8690), .Q(
        g538) );
  SDFFX1 DFF_594_Q_reg ( .D(g33607), .SI(g538), .SE(n8348), .CLK(n8762), .Q(
        g2606) );
  SDFFX1 DFF_595_Q_reg ( .D(g26923), .SI(g2606), .SE(n8308), .CLK(n8722), .Q(
        g1472) );
  SDFFX1 DFF_597_Q_reg ( .D(g24211), .SI(g1472), .SE(n8277), .CLK(n8691), .Q(
        test_so41), .QN(n8232) );
  SDFFX1 DFF_598_Q_reg ( .D(g33050), .SI(test_si42), .SE(n8250), .CLK(n8664), 
        .Q(g5188), .QN(n5567) );
  SDFFX1 DFF_599_Q_reg ( .D(g24341), .SI(g5188), .SE(n8286), .CLK(n8700), .Q(
        g5689), .QN(n5529) );
  SDFFX1 DFF_600_Q_reg ( .D(g19334), .SI(g5689), .SE(n8286), .CLK(n8700), .Q(
        g13259), .QN(n7831) );
  SDFFX1 DFF_601_Q_reg ( .D(g24201), .SI(g13259), .SE(n8312), .CLK(n8726), .Q(
        g405), .QN(n7835) );
  SDFFX1 DFF_602_Q_reg ( .D(g30463), .SI(g405), .SE(n8253), .CLK(n8667), .Q(
        g5216), .QN(n8010) );
  SDFFX1 DFF_603_Q_reg ( .D(g9743), .SI(g5216), .SE(n8313), .CLK(n8727), .Q(
        g6494), .QN(n7729) );
  SDFFX1 DFF_604_Q_reg ( .D(g34464), .SI(g6494), .SE(n8255), .CLK(n8669), .Q(
        g4669), .QN(n7691) );
  SDFFX1 DFF_606_Q_reg ( .D(g24243), .SI(g4669), .SE(n8331), .CLK(n8745), .Q(
        g996) );
  SDFFX1 DFF_607_Q_reg ( .D(g24335), .SI(g996), .SE(n8350), .CLK(n8764), .Q(
        g4531), .QN(n14516) );
  SDFFX1 DFF_608_Q_reg ( .D(g34611), .SI(g4531), .SE(n8289), .CLK(n8703), .Q(
        g2860), .QN(n8164) );
  SDFFX1 DFF_609_Q_reg ( .D(g34262), .SI(g2860), .SE(n8271), .CLK(n8685), .Q(
        g4743) );
  SDFFX1 DFF_610_Q_reg ( .D(g30546), .SI(g4743), .SE(n8329), .CLK(n8743), .Q(
        g6593), .QN(n8113) );
  SDFFX1 DFF_612_Q_reg ( .D(g25591), .SI(g6593), .SE(n8329), .CLK(n8743), .Q(
        test_so42) );
  SDFFX1 DFF_613_Q_reg ( .D(g7257), .SI(test_si43), .SE(n8277), .CLK(n8691), 
        .Q(g4411), .QN(n7681) );
  SDFFX1 DFF_614_Q_reg ( .D(g30347), .SI(g4411), .SE(n8262), .CLK(n8676), .Q(
        g1413) );
  SDFFX1 DFF_615_Q_reg ( .D(test_so38), .SI(g1413), .SE(n8290), .CLK(n8704), 
        .Q(g26960) );
  SDFFX1 DFF_616_Q_reg ( .D(g17577), .SI(g26960), .SE(n8341), .CLK(n8755), .Q(
        g13039), .QN(n8041) );
  SDFFX1 DFF_617_Q_reg ( .D(g30556), .SI(g13039), .SE(n8258), .CLK(n8672), .Q(
        g6641) );
  SDFFX1 DFF_619_Q_reg ( .D(g34970), .SI(g6641), .SE(n8258), .CLK(n8672), .Q(
        g6), .QN(n7765) );
  SDFFX1 DFF_620_Q_reg ( .D(g33562), .SI(g6), .SE(n8345), .CLK(n8759), .Q(
        g1936), .QN(n5534) );
  SDFFX1 DFF_621_Q_reg ( .D(n8192), .SI(g1936), .SE(n8345), .CLK(n8759), .Q(
        g55) );
  SDFFX1 DFF_622_Q_reg ( .D(g25610), .SI(g55), .SE(n8322), .CLK(n8736), .Q(
        g504), .QN(n5519) );
  SDFFX1 DFF_623_Q_reg ( .D(g33015), .SI(g504), .SE(n8293), .CLK(n8707), .Q(
        g2587), .QN(n5372) );
  SDFFX1 DFF_624_Q_reg ( .D(g31896), .SI(g2587), .SE(n8290), .CLK(n8704), .Q(
        g4480) );
  SDFFX1 DFF_625_Q_reg ( .D(g34004), .SI(g4480), .SE(n8287), .CLK(n8701), .Q(
        n9314) );
  SDFFX1 DFF_626_Q_reg ( .D(g30428), .SI(n9314), .SE(n8305), .CLK(n8719), .Q(
        test_so43) );
  SDFFX1 DFF_627_Q_reg ( .D(g30485), .SI(test_si44), .SE(n8259), .CLK(n8673), 
        .Q(g5571) );
  SDFFX1 DFF_628_Q_reg ( .D(g30422), .SI(g5571), .SE(n8304), .CLK(n8718), .Q(
        g3578) );
  SDFFX1 DFF_630_Q_reg ( .D(g25714), .SI(g3578), .SE(n8305), .CLK(n8719), .Q(
        g9555) );
  SDFFX1 DFF_632_Q_reg ( .D(g29294), .SI(g9555), .SE(n8305), .CLK(n8719), .Q(
        g5827), .QN(n5809) );
  SDFFX1 DFF_633_Q_reg ( .D(g30423), .SI(g5827), .SE(n8305), .CLK(n8719), .Q(
        g3582) );
  SDFFX1 DFF_634_Q_reg ( .D(g30529), .SI(g3582), .SE(n8298), .CLK(n8712), .Q(
        g6271) );
  SDFFX1 DFF_635_Q_reg ( .D(g34028), .SI(g6271), .SE(n8298), .CLK(n8712), .Q(
        g4688), .QN(n5656) );
  SDFFX1 DFF_637_Q_reg ( .D(g33587), .SI(g4688), .SE(n8255), .CLK(n8669), .Q(
        g2380), .QN(n7749) );
  SDFFX1 DFF_638_Q_reg ( .D(g30460), .SI(g2380), .SE(n8318), .CLK(n8732), .Q(
        g5196), .QN(n8042) );
  SDFFX1 DFF_640_Q_reg ( .D(g30401), .SI(g5196), .SE(n8320), .CLK(n8734), .Q(
        g3227) );
  SDFFX1 DFF_641_Q_reg ( .D(g33990), .SI(g3227), .SE(n8291), .CLK(n8705), .Q(
        n9312) );
  SDFFX1 DFF_642_Q_reg ( .D(g16693), .SI(n9312), .SE(n8330), .CLK(n8744), .Q(
        g14518) );
  SDFFX1 DFF_643_Q_reg ( .D(g17291), .SI(g14518), .SE(n8330), .CLK(n8744), .Q(
        test_so44) );
  SDFFX1 DFF_644_Q_reg ( .D(g29309), .SI(test_si45), .SE(n8329), .CLK(n8743), 
        .Q(g6541), .QN(n5739) );
  SDFFX1 DFF_645_Q_reg ( .D(g30411), .SI(g6541), .SE(n8321), .CLK(n8735), .Q(
        g3203) );
  SDFFX1 DFF_646_Q_reg ( .D(g33546), .SI(g3203), .SE(n8321), .CLK(n8735), .Q(
        g1668), .QN(n5598) );
  SDFFX1 DFF_647_Q_reg ( .D(g28085), .SI(g1668), .SE(n8258), .CLK(n8672), .Q(
        g4760), .QN(n5775) );
  SDFFX1 DFF_648_Q_reg ( .D(g26904), .SI(g4760), .SE(n8333), .CLK(n8747), .Q(
        g262), .QN(n7869) );
  SDFFX1 DFF_649_Q_reg ( .D(g33556), .SI(g262), .SE(n8352), .CLK(n8766), .Q(
        g1840), .QN(n5451) );
  SDFFX1 DFF_651_Q_reg ( .D(g25722), .SI(g1840), .SE(n8256), .CLK(n8670), .Q(
        g5467), .QN(n7775) );
  SDFFX1 DFF_652_Q_reg ( .D(g25605), .SI(g5467), .SE(n8256), .CLK(n8670), .Q(
        g460) );
  SDFFX1 DFF_653_Q_reg ( .D(g33062), .SI(g460), .SE(n8336), .CLK(n8750), .Q(
        g6209), .QN(n8144) );
  SDFFX1 DFF_654_Q_reg ( .D(g26893), .SI(g6209), .SE(n8322), .CLK(n8736), .Q(
        g29211) );
  SDFFX1 DFF_655_Q_reg ( .D(g12238), .SI(g29211), .SE(n8322), .CLK(n8736), .Q(
        g14662), .QN(n5704) );
  SDFFX1 DFF_656_Q_reg ( .D(g28050), .SI(g14662), .SE(n8322), .CLK(n8736), .Q(
        g655), .QN(n7906) );
  SDFFX1 DFF_657_Q_reg ( .D(g34626), .SI(g655), .SE(n8322), .CLK(n8736), .Q(
        test_so45), .QN(n8227) );
  SDFFX1 DFF_658_Q_reg ( .D(g33583), .SI(test_si46), .SE(n8347), .CLK(n8761), 
        .Q(g2204), .QN(n5620) );
  SDFFX1 DFF_659_Q_reg ( .D(g30472), .SI(g2204), .SE(n8304), .CLK(n8718), .Q(
        g5256) );
  SDFFX1 DFF_660_Q_reg ( .D(g34454), .SI(g5256), .SE(n8304), .CLK(n8718), .Q(
        g4608), .QN(n5274) );
  SDFFX1 DFF_661_Q_reg ( .D(g34850), .SI(g4608), .SE(n8299), .CLK(n8713), .Q(
        g794), .QN(n5291) );
  SDFFX1 DFF_662_Q_reg ( .D(g16955), .SI(g794), .SE(n8333), .CLK(n8747), .Q(
        g13906) );
  SDFFX1 DFF_663_Q_reg ( .D(g10306), .SI(g13906), .SE(n8341), .CLK(n8755), .Q(
        g4423) );
  SDFFX1 DFF_664_Q_reg ( .D(g24272), .SI(g4423), .SE(n8352), .CLK(n8766), .Q(
        g3689), .QN(n5532) );
  SDFFX1 DFF_666_Q_reg ( .D(g17678), .SI(g3689), .SE(n8352), .CLK(n8766), .Q(
        g5685) );
  SDFFX1 DFF_667_Q_reg ( .D(g24214), .SI(g5685), .SE(n8257), .CLK(n8671), .Q(
        g703), .QN(n5821) );
  SDFFX1 DFF_669_Q_reg ( .D(g26909), .SI(g703), .SE(n8275), .CLK(n8689), .Q(
        g862), .QN(n5682) );
  SDFFX1 DFF_670_Q_reg ( .D(g30406), .SI(g862), .SE(n8328), .CLK(n8742), .Q(
        g3247) );
  SDFFX1 DFF_671_Q_reg ( .D(g33569), .SI(g3247), .SE(n8284), .CLK(n8698), .Q(
        g2040), .QN(n5505) );
  SDFFX1 DFF_672_Q_reg ( .D(g25694), .SI(g2040), .SE(n8284), .CLK(n8698), .Q(
        test_so46), .QN(DFF_672_n1) );
  SDFFX1 DFF_673_Q_reg ( .D(g34628), .SI(test_si47), .SE(n8268), .CLK(n8682), 
        .Q(g4146), .QN(n5981) );
  SDFFX1 DFF_674_Q_reg ( .D(g34458), .SI(g4146), .SE(n8331), .CLK(n8745), .Q(
        g4633), .QN(n5844) );
  SDFFX1 DFF_675_Q_reg ( .D(g24240), .SI(g4633), .SE(n8331), .CLK(n8745), .Q(
        g7916), .QN(n5304) );
  SDFFX1 DFF_677_Q_reg ( .D(g34634), .SI(g7916), .SE(n8338), .CLK(n8752), .Q(
        g4732), .QN(n5296) );
  SDFFX1 DFF_678_Q_reg ( .D(g25700), .SI(g4732), .SE(n8250), .CLK(n8664), .Q(
        g9497), .QN(n5689) );
  SDFFX1 DFF_679_Q_reg ( .D(g29293), .SI(g9497), .SE(n8285), .CLK(n8699), .Q(
        g5817) );
  SDFFX1 DFF_681_Q_reg ( .D(g33009), .SI(g5817), .SE(n8294), .CLK(n8708), .Q(
        g2351), .QN(n5511) );
  SDFFX1 DFF_682_Q_reg ( .D(g33603), .SI(g2351), .SE(n8349), .CLK(n8763), .Q(
        g2648), .QN(n7753) );
  SDFFX1 DFF_683_Q_reg ( .D(g24355), .SI(g2648), .SE(n8266), .CLK(n8680), .Q(
        g6736), .QN(n8124) );
  SDFFX1 DFF_684_Q_reg ( .D(g34268), .SI(g6736), .SE(n8279), .CLK(n8693), .Q(
        g4944), .QN(n5875) );
  SDFFX1 DFF_685_Q_reg ( .D(g25691), .SI(g4944), .SE(n8325), .CLK(n8739), .Q(
        g4072), .QN(n8181) );
  SDFFX1 DFF_686_Q_reg ( .D(g26890), .SI(g4072), .SE(n8309), .CLK(n8723), .Q(
        g7540) );
  SDFFX1 DFF_687_Q_reg ( .D(g7260), .SI(g7540), .SE(n8309), .CLK(n8723), .Q(
        test_so47) );
  SDFFX1 DFF_688_Q_reg ( .D(g29264), .SI(test_si48), .SE(n8295), .CLK(n8709), 
        .Q(g3466), .QN(n7731) );
  SDFFX1 DFF_689_Q_reg ( .D(g28072), .SI(g3466), .SE(n8267), .CLK(n8681), .Q(
        g4116) );
  SDFFX1 DFF_690_Q_reg ( .D(g31900), .SI(g4116), .SE(n8251), .CLK(n8665), .Q(
        g5041), .QN(n5605) );
  SDFFX1 DFF_692_Q_reg ( .D(g26956), .SI(g5041), .SE(n8349), .CLK(n8763), .Q(
        g4434), .QN(n7768) );
  SDFFX1 DFF_693_Q_reg ( .D(g29271), .SI(g4434), .SE(n8349), .CLK(n8763), .Q(
        g3827), .QN(n5808) );
  SDFFX1 DFF_694_Q_reg ( .D(g29304), .SI(g3827), .SE(n8259), .CLK(n8673), .Q(
        g6500), .QN(n5748) );
  SDFFX1 DFF_695_Q_reg ( .D(g13049), .SI(g6500), .SE(n8319), .CLK(n8733), .Q(
        g17813) );
  SDFFX1 DFF_696_Q_reg ( .D(g29261), .SI(g17813), .SE(n8270), .CLK(n8684), .Q(
        g3133), .QN(n5661) );
  SDFFX1 DFF_697_Q_reg ( .D(g28063), .SI(g3133), .SE(n8328), .CLK(n8742), .Q(
        g3333) );
  SDFFX1 DFF_698_Q_reg ( .D(g13259), .SI(g3333), .SE(n8328), .CLK(n8742), .Q(
        g979), .QN(n5320) );
  SDFFX1 DFF_699_Q_reg ( .D(g34027), .SI(g979), .SE(n8331), .CLK(n8745), .Q(
        g4681), .QN(n8128) );
  SDFFX1 DFF_700_Q_reg ( .D(g33961), .SI(g4681), .SE(n8276), .CLK(n8690), .Q(
        g298), .QN(n5675) );
  SDFFX1 DFF_702_Q_reg ( .D(g33604), .SI(g298), .SE(n8348), .CLK(n8762), .Q(
        test_so48) );
  SDFFX1 DFF_704_Q_reg ( .D(g8788), .SI(test_si49), .SE(n8315), .CLK(n8729), 
        .Q(g8789), .QN(n7854) );
  SDFFX1 DFF_705_Q_reg ( .D(g32995), .SI(g8789), .SE(n8316), .CLK(n8730), .Q(
        g1894), .QN(n5374) );
  SDFFX1 DFF_706_Q_reg ( .D(g34624), .SI(g1894), .SE(n8289), .CLK(n8703), .Q(
        g2988) );
  SDFFX1 DFF_707_Q_reg ( .D(g30415), .SI(g2988), .SE(n8346), .CLK(n8760), .Q(
        g3538), .QN(n8051) );
  SDFFX1 DFF_708_Q_reg ( .D(g33536), .SI(g3538), .SE(n8299), .CLK(n8713), .Q(
        g301), .QN(n8184) );
  SDFFX1 DFF_709_Q_reg ( .D(g26888), .SI(g301), .SE(n8299), .CLK(n8713), .Q(
        n9306), .QN(DFF_709_n1) );
  SDFFX1 DFF_710_Q_reg ( .D(g28055), .SI(n9306), .SE(n8324), .CLK(n8738), .Q(
        g827), .QN(n5728) );
  SDFFX1 DFF_711_Q_reg ( .D(g24238), .SI(g827), .SE(n8263), .CLK(n8677), .Q(
        g17291) );
  SDFFX1 DFF_713_Q_reg ( .D(g33600), .SI(g17291), .SE(n8348), .CLK(n8762), .Q(
        g2555), .QN(n5351) );
  SDFFX1 DFF_714_Q_reg ( .D(g28105), .SI(g2555), .SE(n8348), .CLK(n8762), .Q(
        g5011) );
  SDFFX1 DFF_715_Q_reg ( .D(g34721), .SI(g5011), .SE(n8348), .CLK(n8762), .Q(
        g199), .QN(n8186) );
  SDFFX1 DFF_716_Q_reg ( .D(g29307), .SI(g199), .SE(n8259), .CLK(n8673), .Q(
        g6523), .QN(n5870) );
  SDFFX1 DFF_717_Q_reg ( .D(g30345), .SI(g6523), .SE(n8293), .CLK(n8707), .Q(
        test_so49), .QN(n8206) );
  SDFFX1 DFF_718_Q_reg ( .D(g34453), .SI(test_si50), .SE(n8304), .CLK(n8718), 
        .Q(g4601), .QN(n5365) );
  SDFFX1 DFF_719_Q_reg ( .D(g32980), .SI(g4601), .SE(n8257), .CLK(n8671), .Q(
        g854), .QN(n5754) );
  SDFFX1 DFF_720_Q_reg ( .D(g29238), .SI(g854), .SE(n8343), .CLK(n8757), .Q(
        g1484), .QN(n5865) );
  SDFFX1 DFF_721_Q_reg ( .D(g34639), .SI(g1484), .SE(n8343), .CLK(n8757), .Q(
        g4922), .QN(n5346) );
  SDFFX1 DFF_722_Q_reg ( .D(g25695), .SI(g4922), .SE(n8248), .CLK(n8662), .Q(
        g5080), .QN(n5893) );
  SDFFX1 DFF_723_Q_reg ( .D(g33057), .SI(g5080), .SE(n8335), .CLK(n8749), .Q(
        g5863), .QN(n8143) );
  SDFFX1 DFF_724_Q_reg ( .D(g26969), .SI(g5863), .SE(n8266), .CLK(n8680), .Q(
        g4581), .QN(n5670) );
  SDFFX1 DFF_726_Q_reg ( .D(g29253), .SI(g4581), .SE(n8349), .CLK(n8763), .Q(
        g2518), .QN(n7917) );
  SDFFX1 DFF_727_Q_reg ( .D(g34021), .SI(g2518), .SE(n8303), .CLK(n8717), .Q(
        g2567) );
  SDFFX1 DFF_728_Q_reg ( .D(g26895), .SI(g2567), .SE(n8282), .CLK(n8696), .Q(
        g568), .QN(n5335) );
  SDFFX1 DFF_729_Q_reg ( .D(g30413), .SI(g568), .SE(n8328), .CLK(n8742), .Q(
        g3263) );
  SDFFX1 DFF_730_Q_reg ( .D(g30549), .SI(g3263), .SE(n8329), .CLK(n8743), .Q(
        g6613) );
  SDFFX1 DFF_731_Q_reg ( .D(g24347), .SI(g6613), .SE(n8258), .CLK(n8672), .Q(
        test_so50), .QN(n8230) );
  SDFFX1 DFF_732_Q_reg ( .D(g25758), .SI(test_si51), .SE(n8313), .CLK(n8727), 
        .Q(g6444), .QN(n5990) );
  SDFFX1 DFF_733_Q_reg ( .D(g34808), .SI(g6444), .SE(n8248), .CLK(n8662), .Q(
        g2965), .QN(n7819) );
  SDFFX1 DFF_734_Q_reg ( .D(g30501), .SI(g2965), .SE(n8335), .CLK(n8749), .Q(
        g5857), .QN(n5573) );
  SDFFX1 DFF_735_Q_reg ( .D(g33969), .SI(g5857), .SE(n8263), .CLK(n8677), .Q(
        n9303) );
  SDFFX1 DFF_736_Q_reg ( .D(g34440), .SI(n9303), .SE(n8274), .CLK(n8688), .Q(
        g890), .QN(n5305) );
  SDFFX1 DFF_737_Q_reg ( .D(g17607), .SI(g890), .SE(n8307), .CLK(n8721), .Q(
        g17646), .QN(n8069) );
  SDFFX1 DFF_738_Q_reg ( .D(g30433), .SI(g17646), .SE(n8306), .CLK(n8720), .Q(
        g3562), .QN(n8115) );
  SDFFX1 DFF_739_Q_reg ( .D(g21900), .SI(g3562), .SE(n8306), .CLK(n8720), .Q(
        g10122_Tj), .QN(n7726) );
  SDFFX1 DFF_740_Q_reg ( .D(g26921), .SI(g10122_Tj), .SE(n8318), .CLK(n8732), 
        .Q(g1404), .QN(n7839) );
  SDFFX1 DFF_742_Q_reg ( .D(g29270), .SI(g1404), .SE(n8278), .CLK(n8692), .Q(
        g3817), .QN(n7710) );
  SDFFX1 DFF_743_Q_reg ( .D(n8197), .SI(g3817), .SE(n8251), .CLK(n8665), .Q(
        n9302), .QN(n6010) );
  SDFFX1 DFF_744_Q_reg ( .D(g33038), .SI(n9302), .SE(n8290), .CLK(n8704), .Q(
        g4501) );
  SDFFX1 DFF_745_Q_reg ( .D(g31865), .SI(g4501), .SE(n8307), .CLK(n8721), .Q(
        test_so51), .QN(n8241) );
  SDFFX1 DFF_746_Q_reg ( .D(g26926), .SI(test_si52), .SE(n8281), .CLK(n8695), 
        .Q(g2724), .QN(n5301) );
  SDFFX1 DFF_747_Q_reg ( .D(g28083), .SI(g2724), .SE(n8269), .CLK(n8683), .Q(
        g4704), .QN(n5771) );
  SDFFX1 DFF_749_Q_reg ( .D(g34797), .SI(g22), .SE(n8270), .CLK(n8684), .Q(
        g2878), .QN(n8173) );
  SDFFX1 DFF_750_Q_reg ( .D(g30478), .SI(g2878), .SE(n8253), .CLK(n8667), .Q(
        g5220), .QN(n8003) );
  SDFFX1 DFF_751_Q_reg ( .D(g34724), .SI(g5220), .SE(n8282), .CLK(n8696), .Q(
        g617), .QN(n5339) );
  SDFFX1 DFF_752_Q_reg ( .D(g24212), .SI(g617), .SE(n8282), .CLK(n8696), .Q(
        g12368) );
  SDFFX1 DFF_753_Q_reg ( .D(g26883), .SI(g12368), .SE(n8308), .CLK(n8722), .Q(
        g316) );
  SDFFX1 DFF_754_Q_reg ( .D(g32985), .SI(g316), .SE(n8348), .CLK(n8762), .Q(
        g1277), .QN(n8183) );
  SDFFX1 DFF_755_Q_reg ( .D(g25761), .SI(g1277), .SE(n8259), .CLK(n8673), .Q(
        g6513), .QN(n5426) );
  SDFFX1 DFF_756_Q_reg ( .D(g26886), .SI(g6513), .SE(n8309), .CLK(n8723), .Q(
        g336), .QN(n5824) );
  SDFFX1 DFF_757_Q_reg ( .D(g34796), .SI(g336), .SE(n8270), .CLK(n8684), .Q(
        g2882), .QN(n7677) );
  SDFFX1 DFF_758_Q_reg ( .D(g32982), .SI(g2882), .SE(n8276), .CLK(n8690), .Q(
        test_so52), .QN(n8188) );
  SDFFX1 DFF_759_Q_reg ( .D(g33561), .SI(test_si53), .SE(n8345), .CLK(n8759), 
        .Q(g1906), .QN(n5503) );
  SDFFX1 DFF_760_Q_reg ( .D(g26880), .SI(g1906), .SE(n8345), .CLK(n8759), .Q(
        g305), .QN(n5282) );
  SDFFX1 DFF_761_Q_reg ( .D(n171), .SI(g305), .SE(n8345), .CLK(n8759), .Q(g8), 
        .QN(n7766) );
  SDFFX1 DFF_763_Q_reg ( .D(g26931), .SI(g8), .SE(n8261), .CLK(n8675), .Q(
        g2799) );
  SDFFX1 DFF_764_Q_reg ( .D(g14147), .SI(g2799), .SE(n8300), .CLK(n8714), .Q(
        g14167) );
  SDFFX1 DFF_765_Q_reg ( .D(g13039), .SI(g14167), .SE(n8341), .CLK(n8755), .Q(
        g17787) );
  SDFFX1 DFF_766_Q_reg ( .D(g34641), .SI(g17787), .SE(n8343), .CLK(n8757), .Q(
        g4912), .QN(n5297) );
  SDFFX1 DFF_767_Q_reg ( .D(g34629), .SI(g4912), .SE(n8268), .CLK(n8682), .Q(
        g4157), .QN(n5983) );
  SDFFX1 DFF_768_Q_reg ( .D(g33598), .SI(g4157), .SE(n8268), .CLK(n8682), .Q(
        g2541), .QN(n5461) );
  SDFFX1 DFF_769_Q_reg ( .D(g33576), .SI(g2541), .SE(n8261), .CLK(n8675), .Q(
        g2153), .QN(n5356) );
  SDFFX1 DFF_770_Q_reg ( .D(g34720), .SI(g2153), .SE(n8277), .CLK(n8691), .Q(
        g550), .QN(n8185) );
  SDFFX1 DFF_771_Q_reg ( .D(g26902), .SI(g550), .SE(n8333), .CLK(n8747), .Q(
        g255), .QN(n7868) );
  SDFFX1 DFF_772_Q_reg ( .D(g29244), .SI(g255), .SE(n8353), .CLK(n8767), .Q(
        test_so53) );
  SDFFX1 DFF_773_Q_reg ( .D(g30468), .SI(test_si54), .SE(n8318), .CLK(n8732), 
        .Q(g5240) );
  SDFFX1 DFF_774_Q_reg ( .D(g26924), .SI(g5240), .SE(n8323), .CLK(n8737), .Q(
        g1478), .QN(n5289) );
  SDFFX1 DFF_776_Q_reg ( .D(g33031), .SI(g1478), .SE(n8323), .CLK(n8737), .Q(
        g3863), .QN(n8142) );
  SDFFX1 DFF_777_Q_reg ( .D(g29245), .SI(g3863), .SE(n8353), .CLK(n8767), .Q(
        g1959), .QN(n7916) );
  SDFFX1 DFF_778_Q_reg ( .D(g29266), .SI(g1959), .SE(n8279), .CLK(n8693), .Q(
        g3480), .QN(n5868) );
  SDFFX1 DFF_779_Q_reg ( .D(g30559), .SI(g3480), .SE(n8340), .CLK(n8754), .Q(
        g6653) );
  SDFFX1 DFF_780_Q_reg ( .D(g14749), .SI(g6653), .SE(n8349), .CLK(n8763), .Q(
        g17764) );
  SDFFX1 DFF_781_Q_reg ( .D(g34794), .SI(g17764), .SE(n8252), .CLK(n8666), .Q(
        g2864) );
  SDFFX1 DFF_782_Q_reg ( .D(g28087), .SI(g2864), .SE(n8266), .CLK(n8680), .Q(
        g4894), .QN(n5774) );
  SDFFX1 DFF_783_Q_reg ( .D(g14635), .SI(g4894), .SE(n8320), .CLK(n8734), .Q(
        g17678) );
  SDFFX1 DFF_784_Q_reg ( .D(g30435), .SI(g17678), .SE(n8330), .CLK(n8744), .Q(
        g3857), .QN(n5572) );
  SDFFX1 DFF_785_Q_reg ( .D(g16659), .SI(g3857), .SE(n8330), .CLK(n8744), .Q(
        g16693), .QN(n8078) );
  SDFFX1 DFF_786_Q_reg ( .D(g25609), .SI(g16693), .SE(n8343), .CLK(n8757), .Q(
        test_so54), .QN(n8221) );
  SDFFX1 DFF_788_Q_reg ( .D(g28057), .SI(test_si55), .SE(n8263), .CLK(n8677), 
        .Q(g1002), .QN(n7837) );
  SDFFX1 DFF_789_Q_reg ( .D(g34439), .SI(g1002), .SE(n8316), .CLK(n8730), .Q(
        g776), .QN(n5330) );
  SDFFX1 DFF_790_Q_reg ( .D(g34979), .SI(g776), .SE(n8316), .CLK(n8730), .Q(
        g28), .QN(n5324) );
  SDFFX1 DFF_791_Q_reg ( .D(g10500), .SI(g28), .SE(n8330), .CLK(n8744), .Q(
        g1236), .QN(n7808) );
  SDFFX1 DFF_792_Q_reg ( .D(g34260), .SI(g1236), .SE(n8330), .CLK(n8744), .Q(
        g4646), .QN(n5712) );
  SDFFX1 DFF_793_Q_reg ( .D(g33012), .SI(g4646), .SE(n8331), .CLK(n8745), .Q(
        g2476), .QN(n8131) );
  SDFFX1 DFF_794_Q_reg ( .D(g32989), .SI(g2476), .SE(n8296), .CLK(n8710), .Q(
        g1657), .QN(n5525) );
  SDFFX1 DFF_795_Q_reg ( .D(g34006), .SI(g1657), .SE(n8255), .CLK(n8669), .Q(
        g2375), .QN(n7786) );
  SDFFX1 DFF_796_Q_reg ( .D(g34783), .SI(g2375), .SE(n8298), .CLK(n8712), .Q(
        g63) );
  SDFFX1 DFF_797_Q_reg ( .D(g14738), .SI(g63), .SE(n8306), .CLK(n8720), .Q(
        g17739), .QN(n7973) );
  SDFFX1 DFF_798_Q_reg ( .D(g8719), .SI(g17739), .SE(n8306), .CLK(n8720), .Q(
        g358), .QN(n7872) );
  SDFFX1 DFF_799_Q_reg ( .D(g26910), .SI(g358), .SE(n8306), .CLK(n8720), .Q(
        g896), .QN(n5431) );
  SDFFX1 DFF_802_Q_reg ( .D(g28043), .SI(g896), .SE(n8307), .CLK(n8721), .Q(
        test_so55), .QN(n8228) );
  SDFFX1 DFF_803_Q_reg ( .D(g33021), .SI(test_si56), .SE(n8326), .CLK(n8740), 
        .Q(g3161), .QN(n8150) );
  SDFFX1 DFF_804_Q_reg ( .D(g29251), .SI(g3161), .SE(n8318), .CLK(n8732), .Q(
        g2384), .QN(n7911) );
  SDFFX1 DFF_806_Q_reg ( .D(test_so80), .SI(g2384), .SE(n8318), .CLK(n8732), 
        .Q(g14828), .QN(n5700) );
  SDFFX1 DFF_807_Q_reg ( .D(g34456), .SI(g14828), .SE(n8304), .CLK(n8718), .Q(
        g4616), .QN(n5608) );
  SDFFX1 DFF_808_Q_reg ( .D(g26968), .SI(g4616), .SE(n8342), .CLK(n8756), .Q(
        g4561) );
  SDFFX1 DFF_809_Q_reg ( .D(g33991), .SI(g4561), .SE(n8291), .CLK(n8705), .Q(
        g2024), .QN(n5801) );
  SDFFX1 DFF_810_Q_reg ( .D(g8279), .SI(g2024), .SE(n8252), .CLK(n8666), .Q(
        g3451), .QN(n7713) );
  SDFFX1 DFF_811_Q_reg ( .D(g26930), .SI(g3451), .SE(n8282), .CLK(n8696), .Q(
        g2795) );
  SDFFX1 DFF_812_Q_reg ( .D(g34599), .SI(g2795), .SE(n8282), .CLK(n8696), .Q(
        g613), .QN(n5474) );
  SDFFX1 DFF_813_Q_reg ( .D(g28082), .SI(g613), .SE(n8350), .CLK(n8764), .Q(
        g4527), .QN(n8159) );
  SDFFX1 DFF_814_Q_reg ( .D(g33557), .SI(g4527), .SE(n8274), .CLK(n8688), .Q(
        g1844) );
  SDFFX1 DFF_815_Q_reg ( .D(g30511), .SI(g1844), .SE(n8337), .CLK(n8751), .Q(
        g5937) );
  SDFFX1 DFF_816_Q_reg ( .D(g33045), .SI(g5937), .SE(n8337), .CLK(n8751), .Q(
        test_so56) );
  SDFFX1 DFF_818_Q_reg ( .D(g30379), .SI(test_si57), .SE(n8308), .CLK(n8722), 
        .Q(g2523), .QN(n5281) );
  SDFFX1 DFF_819_Q_reg ( .D(g24267), .SI(g2523), .SE(n8339), .CLK(n8753), .Q(
        g11349), .QN(n5436) );
  SDFFX1 DFF_820_Q_reg ( .D(g34020), .SI(g11349), .SE(n8307), .CLK(n8721), .Q(
        g2643), .QN(n7785) );
  SDFFX1 DFF_822_Q_reg ( .D(g24249), .SI(g2643), .SE(n8307), .CLK(n8721), .Q(
        g1489), .QN(n5850) );
  SDFFX1 DFF_824_Q_reg ( .D(g25592), .SI(g1489), .SE(n8276), .CLK(n8690), .Q(
        g8358), .QN(n7846) );
  SDFFX1 DFF_825_Q_reg ( .D(g30382), .SI(g8358), .SE(n8268), .CLK(n8682), .Q(
        n9295) );
  SDFFX1 DFF_826_Q_reg ( .D(g29285), .SI(n9295), .SE(n8268), .CLK(n8682), .Q(
        g5156), .QN(n5734) );
  SDFFX1 DFF_828_Q_reg ( .D(g12919), .SI(g5156), .SE(n8275), .CLK(n8689), .Q(
        g30332), .QN(n5526) );
  SDFFX1 DFF_829_Q_reg ( .D(n171), .SI(g30332), .SE(n8252), .CLK(n8666), .Q(
        n9294), .QN(n14515) );
  SDFFX1 DFF_830_Q_reg ( .D(g25662), .SI(n9294), .SE(n8252), .CLK(n8666), .Q(
        g8279) );
  SDFFX1 DFF_831_Q_reg ( .D(g21896), .SI(g8279), .SE(n8303), .CLK(n8717), .Q(
        g8839) );
  SDFFX1 DFF_832_Q_reg ( .D(g33563), .SI(g8839), .SE(n8286), .CLK(n8700), .Q(
        g1955), .QN(n7746) );
  SDFFX1 DFF_833_Q_reg ( .D(g33622), .SI(g1955), .SE(n8331), .CLK(n8745), .Q(
        test_so57), .QN(n8216) );
  SDFFX1 DFF_835_Q_reg ( .D(g33582), .SI(test_si58), .SE(n8349), .CLK(n8763), 
        .Q(g2273), .QN(n5458) );
  SDFFX1 DFF_836_Q_reg ( .D(g17871), .SI(g2273), .SE(n8349), .CLK(n8763), .Q(
        g14749) );
  SDFFX1 DFF_837_Q_reg ( .D(g28086), .SI(g14749), .SE(n8351), .CLK(n8765), .Q(
        g4771), .QN(n5769) );
  SDFFX1 DFF_838_Q_reg ( .D(g25744), .SI(g4771), .SE(n8278), .CLK(n8692), .Q(
        g6098), .QN(n5988) );
  SDFFX1 DFF_839_Q_reg ( .D(g29262), .SI(g6098), .SE(n8328), .CLK(n8742), .Q(
        g3147), .QN(n5738) );
  SDFFX1 DFF_840_Q_reg ( .D(g24270), .SI(g3147), .SE(n8321), .CLK(n8735), .Q(
        g3347), .QN(n7984) );
  SDFFX1 DFF_841_Q_reg ( .D(g33581), .SI(g3347), .SE(n8310), .CLK(n8724), .Q(
        g2269) );
  SDFFX1 DFF_842_Q_reg ( .D(g8358), .SI(g2269), .SE(n8310), .CLK(n8724), .Q(
        g191), .QN(n7847) );
  SDFFX1 DFF_843_Q_reg ( .D(g24266), .SI(g191), .SE(n8310), .CLK(n8724), .Q(
        g2712), .QN(n7722) );
  SDFFX1 DFF_844_Q_reg ( .D(g34849), .SI(g2712), .SE(n8282), .CLK(n8696), .Q(
        g626), .QN(n5288) );
  SDFFX1 DFF_846_Q_reg ( .D(g33618), .SI(g2729), .SE(n8269), .CLK(n8683), .Q(
        g5357), .QN(n5393) );
  SDFFX1 DFF_847_Q_reg ( .D(g34038), .SI(g5357), .SE(n8295), .CLK(n8709), .Q(
        test_so58), .QN(n8214) );
  SDFFX1 DFF_848_Q_reg ( .D(g13068), .SI(test_si59), .SE(n8285), .CLK(n8699), 
        .Q(g17819) );
  SDFFX1 DFF_849_Q_reg ( .D(g34032), .SI(g17819), .SE(n8327), .CLK(n8741), .Q(
        g4709), .QN(n5518) );
  SDFFX1 DFF_852_Q_reg ( .D(g34803), .SI(g4709), .SE(n8264), .CLK(n8678), .Q(
        g2927), .QN(n7816) );
  SDFFX1 DFF_853_Q_reg ( .D(g34459), .SI(g2927), .SE(n8301), .CLK(n8715), .Q(
        g4340), .QN(n5653) );
  SDFFX1 DFF_854_Q_reg ( .D(g30509), .SI(g4340), .SE(n8288), .CLK(n8702), .Q(
        g5929) );
  SDFFX1 DFF_855_Q_reg ( .D(g34640), .SI(g5929), .SE(n8343), .CLK(n8757), .Q(
        g4907), .QN(n5295) );
  SDFFX1 DFF_856_Q_reg ( .D(g14421), .SI(g4907), .SE(n8343), .CLK(n8757), .Q(
        g16874) );
  SDFFX1 DFF_857_Q_reg ( .D(g28069), .SI(g16874), .SE(n8265), .CLK(n8679), .Q(
        g4035) );
  SDFFX1 DFF_858_Q_reg ( .D(g21899), .SI(g4035), .SE(n8303), .CLK(n8717), .Q(
        g2946), .QN(n8175) );
  SDFFX1 DFF_859_Q_reg ( .D(g31868), .SI(g2946), .SE(n8275), .CLK(n8689), .Q(
        g918), .QN(n5673) );
  SDFFX1 DFF_860_Q_reg ( .D(g26938), .SI(g918), .SE(n8325), .CLK(n8739), .Q(
        g4082), .QN(n7826) );
  SDFFX1 DFF_861_Q_reg ( .D(g25756), .SI(g4082), .SE(n8313), .CLK(n8727), .Q(
        g9743) );
  SDFFX1 DFF_862_Q_reg ( .D(g30363), .SI(g9743), .SE(n8284), .CLK(n8698), .Q(
        test_so59), .QN(n8244) );
  SDFFX1 DFF_863_Q_reg ( .D(g30334), .SI(test_si60), .SE(n8283), .CLK(n8697), 
        .Q(g577), .QN(n5294) );
  SDFFX1 DFF_864_Q_reg ( .D(g33970), .SI(g577), .SE(n8346), .CLK(n8760), .Q(
        g1620) );
  SDFFX1 DFF_865_Q_reg ( .D(g30391), .SI(g1620), .SE(n8264), .CLK(n8678), .Q(
        g2831), .QN(g30331) );
  SDFFX1 DFF_866_Q_reg ( .D(g25615), .SI(g2831), .SE(n8264), .CLK(n8678), .Q(
        g667) );
  SDFFX1 DFF_867_Q_reg ( .D(g33540), .SI(g667), .SE(n8276), .CLK(n8690), .Q(
        g930), .QN(n5731) );
  SDFFX1 DFF_868_Q_reg ( .D(g30445), .SI(g930), .SE(n8324), .CLK(n8738), .Q(
        g3937) );
  SDFFX1 DFF_870_Q_reg ( .D(g25617), .SI(g3937), .SE(n8324), .CLK(n8738), .Q(
        g817), .QN(n5822) );
  SDFFX1 DFF_871_Q_reg ( .D(g24247), .SI(g817), .SE(n8324), .CLK(n8738), .Q(
        g1249) );
  SDFFX1 DFF_872_Q_reg ( .D(g24215), .SI(g1249), .SE(n8324), .CLK(n8738), .Q(
        g837), .QN(n5562) );
  SDFFX1 DFF_873_Q_reg ( .D(g14451), .SI(g837), .SE(n8324), .CLK(n8738), .Q(
        g16924) );
  SDFFX1 DFF_874_Q_reg ( .D(g33964), .SI(g16924), .SE(n8283), .CLK(n8697), .Q(
        g599), .QN(n5550) );
  SDFFX1 DFF_875_Q_reg ( .D(g25719), .SI(g599), .SE(n8283), .CLK(n8697), .Q(
        g5475), .QN(n5425) );
  SDFFX1 DFF_876_Q_reg ( .D(g29228), .SI(g5475), .SE(n8299), .CLK(n8713), .Q(
        test_so60) );
  SDFFX1 DFF_877_Q_reg ( .D(g30514), .SI(test_si61), .SE(n8337), .CLK(n8751), 
        .Q(g5949) );
  SDFFX1 DFF_878_Q_reg ( .D(g33627), .SI(g5949), .SE(n8292), .CLK(n8706), .Q(
        g6682), .QN(n5590) );
  SDFFX1 DFF_880_Q_reg ( .D(g24231), .SI(g6682), .SE(n8292), .CLK(n8706), .Q(
        g904) );
  SDFFX1 DFF_881_Q_reg ( .D(g34615), .SI(g904), .SE(n8289), .CLK(n8703), .Q(
        g2873) );
  SDFFX1 DFF_882_Q_reg ( .D(g30356), .SI(g2873), .SE(n8274), .CLK(n8688), .Q(
        g1854), .QN(n5785) );
  SDFFX1 DFF_883_Q_reg ( .D(g25696), .SI(g1854), .SE(n8248), .CLK(n8662), .Q(
        g5084), .QN(n5681) );
  SDFFX1 DFF_884_Q_reg ( .D(g30493), .SI(g5084), .SE(n8259), .CLK(n8673), .Q(
        g5603) );
  SDFFX1 DFF_885_Q_reg ( .D(g8917), .SI(g5603), .SE(n8259), .CLK(n8673), .Q(
        g8870), .QN(n5726) );
  SDFFX1 DFF_886_Q_reg ( .D(g33594), .SI(g8870), .SE(n8310), .CLK(n8724), .Q(
        g2495), .QN(n5522) );
  SDFFX1 DFF_887_Q_reg ( .D(g34009), .SI(g2495), .SE(n8349), .CLK(n8763), .Q(
        g2437) );
  SDFFX1 DFF_888_Q_reg ( .D(g30365), .SI(g2437), .SE(n8285), .CLK(n8699), .Q(
        g2102), .QN(n5666) );
  SDFFX1 DFF_889_Q_reg ( .D(g33004), .SI(g2102), .SE(n8310), .CLK(n8724), .Q(
        g2208), .QN(n8133) );
  SDFFX1 DFF_890_Q_reg ( .D(g34018), .SI(g2208), .SE(n8293), .CLK(n8707), .Q(
        test_so61) );
  SDFFX1 DFF_891_Q_reg ( .D(g25685), .SI(test_si62), .SE(n8325), .CLK(n8739), 
        .Q(g4064), .QN(n5416) );
  SDFFX1 DFF_892_Q_reg ( .D(g34040), .SI(g4064), .SE(n8351), .CLK(n8765), .Q(
        g4899), .QN(n5517) );
  SDFFX1 DFF_893_Q_reg ( .D(g25639), .SI(g4899), .SE(n8281), .CLK(n8695), .Q(
        g2719), .QN(n5465) );
  SDFFX1 DFF_894_Q_reg ( .D(g34029), .SI(g2719), .SE(n8327), .CLK(n8741), .Q(
        g4785), .QN(n5361) );
  SDFFX1 DFF_895_Q_reg ( .D(g30488), .SI(g4785), .SE(n8249), .CLK(n8663), .Q(
        g5583) );
  SDFFX1 DFF_896_Q_reg ( .D(g34600), .SI(g5583), .SE(n8316), .CLK(n8730), .Q(
        g781), .QN(n5551) );
  SDFFX1 DFF_897_Q_reg ( .D(g29300), .SI(g781), .SE(n8317), .CLK(n8731), .Q(
        g6173), .QN(n5810) );
  SDFFX1 DFF_898_Q_reg ( .D(g14705), .SI(g6173), .SE(n8317), .CLK(n8731), .Q(
        g17743) );
  SDFFX1 DFF_899_Q_reg ( .D(g34802), .SI(g17743), .SE(n8264), .CLK(n8678), .Q(
        g2917), .QN(n7817) );
  SDFFX1 DFF_900_Q_reg ( .D(g25614), .SI(g2917), .SE(n8322), .CLK(n8736), .Q(
        g686) );
  SDFFX1 DFF_901_Q_reg ( .D(g28058), .SI(g686), .SE(n8314), .CLK(n8728), .Q(
        g1252), .QN(n5554) );
  SDFFX1 DFF_902_Q_reg ( .D(g29225), .SI(g1252), .SE(n8264), .CLK(n8678), .Q(
        g671), .QN(n7718) );
  SDFFX1 DFF_903_Q_reg ( .D(g33580), .SI(g671), .SE(n8347), .CLK(n8761), .Q(
        test_so62) );
  SDFFX1 DFF_904_Q_reg ( .D(g30532), .SI(test_si63), .SE(n8297), .CLK(n8711), 
        .Q(g6283) );
  SDFFX1 DFF_905_Q_reg ( .D(g17845), .SI(g6283), .SE(n8340), .CLK(n8754), .Q(
        g14705) );
  SDFFX1 DFF_906_Q_reg ( .D(g17674), .SI(g14705), .SE(n8341), .CLK(n8755), .Q(
        g17519), .QN(n7956) );
  SDFFX1 DFF_909_Q_reg ( .D(g8783), .SI(g17519), .SE(n8341), .CLK(n8755), .Q(
        g8784), .QN(n14527) );
  SDFFX1 DFF_910_Q_reg ( .D(g33054), .SI(g8784), .SE(n8341), .CLK(n8755), .Q(
        g5527), .QN(n5389) );
  SDFFX1 DFF_911_Q_reg ( .D(g26962), .SI(g5527), .SE(n8341), .CLK(n8755), .Q(
        g4489) );
  SDFFX1 DFF_912_Q_reg ( .D(g33564), .SI(g4489), .SE(n8345), .CLK(n8759), .Q(
        g1974), .QN(n5450) );
  SDFFX1 DFF_913_Q_reg ( .D(g32984), .SI(g1974), .SE(n8314), .CLK(n8728), .Q(
        g1270), .QN(n5716) );
  SDFFX1 DFF_914_Q_reg ( .D(g34039), .SI(g1270), .SE(n8298), .CLK(n8712), .Q(
        g4966), .QN(n5706) );
  SDFFX1 DFF_916_Q_reg ( .D(g33065), .SI(g4966), .SE(n8336), .CLK(n8750), .Q(
        g6227), .QN(n5568) );
  SDFFX1 DFF_917_Q_reg ( .D(g30443), .SI(g6227), .SE(n8265), .CLK(n8679), .Q(
        g3929) );
  SDFFX1 DFF_918_Q_reg ( .D(g29291), .SI(g3929), .SE(n8256), .CLK(n8670), .Q(
        g5503), .QN(n5737) );
  SDFFX1 DFF_919_Q_reg ( .D(g24279), .SI(g5503), .SE(n8253), .CLK(n8667), .Q(
        test_so63), .QN(n8177) );
  SDFFX1 DFF_920_Q_reg ( .D(g30508), .SI(test_si64), .SE(n8351), .CLK(n8765), 
        .Q(g5925) );
  SDFFX1 DFF_921_Q_reg ( .D(g29232), .SI(g5925), .SE(n8286), .CLK(n8700), .Q(
        g1124) );
  SDFFX1 DFF_922_Q_reg ( .D(g34269), .SI(g1124), .SE(n8267), .CLK(n8681), .Q(
        g4955), .QN(n5614) );
  SDFFX1 DFF_923_Q_reg ( .D(g30464), .SI(g4955), .SE(n8318), .CLK(n8732), .Q(
        g5224) );
  SDFFX1 DFF_924_Q_reg ( .D(g33988), .SI(g5224), .SE(n8291), .CLK(n8705), .Q(
        g2012) );
  SDFFX1 DFF_925_Q_reg ( .D(g30522), .SI(g2012), .SE(n8336), .CLK(n8750), .Q(
        g6203), .QN(n5574) );
  SDFFX1 DFF_926_Q_reg ( .D(g25708), .SI(g6203), .SE(n8268), .CLK(n8682), .Q(
        g5120), .QN(n7774) );
  SDFFX1 DFF_927_Q_reg ( .D(g14662), .SI(g5120), .SE(n8322), .CLK(n8736), .Q(
        g17674), .QN(n7971) );
  SDFFX1 DFF_928_Q_reg ( .D(g30374), .SI(g17674), .SE(n8255), .CLK(n8669), .Q(
        g2389), .QN(n5631) );
  SDFFX1 DFF_929_Q_reg ( .D(g26953), .SI(g2389), .SE(n8341), .CLK(n8755), .Q(
        g4438), .QN(n8139) );
  SDFFX1 DFF_930_Q_reg ( .D(g34008), .SI(g4438), .SE(n8348), .CLK(n8762), .Q(
        g2429) );
  SDFFX1 DFF_931_Q_reg ( .D(g34444), .SI(g2429), .SE(n8281), .CLK(n8695), .Q(
        g2787), .QN(n5610) );
  SDFFX1 DFF_932_Q_reg ( .D(g34731), .SI(g2787), .SE(n8262), .CLK(n8676), .Q(
        test_so64) );
  SDFFX1 DFF_933_Q_reg ( .D(g33606), .SI(test_si65), .SE(n8260), .CLK(n8674), 
        .Q(g2675), .QN(n5457) );
  SDFFX1 DFF_934_Q_reg ( .D(g24334), .SI(g2675), .SE(n8301), .CLK(n8715), .Q(
        g18881), .QN(n5541) );
  SDFFX1 DFF_935_Q_reg ( .D(g34265), .SI(g18881), .SE(n8301), .CLK(n8715), .Q(
        g4836), .QN(n5713) );
  SDFFX1 DFF_936_Q_reg ( .D(g30340), .SI(g4836), .SE(n8254), .CLK(n8668), .Q(
        g1199), .QN(n7863) );
  SDFFX1 DFF_937_Q_reg ( .D(g24257), .SI(g1199), .SE(n8254), .CLK(n8668), .Q(
        g19357), .QN(n5401) );
  SDFFX1 DFF_938_Q_reg ( .D(g30482), .SI(g19357), .SE(n8260), .CLK(n8674), .Q(
        g5547), .QN(n7884) );
  SDFFX1 DFF_941_Q_reg ( .D(g34604), .SI(g5547), .SE(n8283), .CLK(n8697), .Q(
        g2138), .QN(n5275) );
  SDFFX1 DFF_942_Q_reg ( .D(g13926), .SI(g2138), .SE(n8297), .CLK(n8711), .Q(
        g16744), .QN(n7980) );
  SDFFX1 DFF_943_Q_reg ( .D(g33591), .SI(g16744), .SE(n8311), .CLK(n8725), .Q(
        g2338) );
  SDFFX1 DFF_944_Q_reg ( .D(g8918), .SI(g2338), .SE(n8311), .CLK(n8725), .Q(
        g8919), .QN(n14525) );
  SDFFX1 DFF_945_Q_reg ( .D(g30525), .SI(g8919), .SE(n8298), .CLK(n8712), .Q(
        g6247), .QN(n8121) );
  SDFFX1 DFF_946_Q_reg ( .D(g26929), .SI(g6247), .SE(n8282), .CLK(n8696), .Q(
        g2791) );
  SDFFX1 DFF_947_Q_reg ( .D(g30448), .SI(g2791), .SE(n8334), .CLK(n8748), .Q(
        test_so65) );
  SDFFX1 DFF_948_Q_reg ( .D(g34602), .SI(test_si66), .SE(n8248), .CLK(n8662), 
        .Q(g1291), .QN(n2549) );
  SDFFX1 DFF_949_Q_reg ( .D(g30513), .SI(g1291), .SE(n8288), .CLK(n8702), .Q(
        g5945) );
  SDFFX1 DFF_950_Q_reg ( .D(g30469), .SI(g5945), .SE(n8302), .CLK(n8716), .Q(
        g5244) );
  SDFFX1 DFF_951_Q_reg ( .D(g33608), .SI(g5244), .SE(n8302), .CLK(n8716), .Q(
        g2759), .QN(n7684) );
  SDFFX1 DFF_952_Q_reg ( .D(g33626), .SI(g2759), .SE(n8327), .CLK(n8741), .Q(
        g6741), .QN(n5398) );
  SDFFX1 DFF_953_Q_reg ( .D(g34725), .SI(g6741), .SE(n8346), .CLK(n8760), .Q(
        g785), .QN(n5293) );
  SDFFX1 DFF_954_Q_reg ( .D(g30342), .SI(g785), .SE(n8314), .CLK(n8728), .Q(
        g1259), .QN(n5553) );
  SDFFX1 DFF_955_Q_reg ( .D(g29267), .SI(g1259), .SE(n8279), .CLK(n8693), .Q(
        g3484), .QN(n5668) );
  SDFFX1 DFF_956_Q_reg ( .D(g25593), .SI(g3484), .SE(n8276), .CLK(n8690), .Q(
        g209), .QN(n5595) );
  SDFFX1 DFF_957_Q_reg ( .D(g30548), .SI(g209), .SE(n8329), .CLK(n8743), .Q(
        g6609) );
  SDFFX1 DFF_958_Q_reg ( .D(g33052), .SI(g6609), .SE(n8279), .CLK(n8693), .Q(
        g5517), .QN(n8145) );
  SDFFX1 DFF_959_Q_reg ( .D(g34012), .SI(g5517), .SE(n8280), .CLK(n8694), .Q(
        g2449) );
  SDFFX1 DFF_960_Q_reg ( .D(g34017), .SI(g2449), .SE(n8293), .CLK(n8707), .Q(
        test_so66) );
  SDFFX1 DFF_961_Q_reg ( .D(g18881), .SI(test_si67), .SE(n8301), .CLK(n8715), 
        .Q(n9281) );
  SDFFX1 DFF_962_Q_reg ( .D(g24263), .SI(n9281), .SE(n8310), .CLK(n8724), .Q(
        g2715), .QN(n5299) );
  SDFFX1 DFF_963_Q_reg ( .D(g26912), .SI(g2715), .SE(n8275), .CLK(n8689), .Q(
        g936), .QN(n5557) );
  SDFFX1 DFF_964_Q_reg ( .D(g30364), .SI(g936), .SE(n8285), .CLK(n8699), .Q(
        g2098), .QN(n5280) );
  SDFFX1 DFF_965_Q_reg ( .D(g34254), .SI(g2098), .SE(n8332), .CLK(n8746), .Q(
        g4462), .QN(n5671) );
  SDFFX1 DFF_966_Q_reg ( .D(g34251), .SI(g4462), .SE(n8283), .CLK(n8697), .Q(
        g604), .QN(n5473) );
  SDFFX1 DFF_967_Q_reg ( .D(g30560), .SI(g604), .SE(n8258), .CLK(n8672), .Q(
        g6589), .QN(n8048) );
  SDFFX1 DFF_968_Q_reg ( .D(g33983), .SI(g6589), .SE(n8287), .CLK(n8701), .Q(
        n9280) );
  SDFFX1 DFF_970_Q_reg ( .D(g13085), .SI(n9280), .SE(n8340), .CLK(n8754), .Q(
        g17845) );
  SDFFX1 DFF_971_Q_reg ( .D(g13099), .SI(g17845), .SE(n8340), .CLK(n8754), .Q(
        g17871) );
  SDFFX1 DFF_972_Q_reg ( .D(g24204), .SI(g17871), .SE(n8257), .CLK(n8671), .Q(
        g429) );
  SDFFX1 DFF_973_Q_reg ( .D(g33980), .SI(g429), .SE(n8286), .CLK(n8700), .Q(
        g1870) );
  SDFFX1 DFF_974_Q_reg ( .D(g34631), .SI(g1870), .SE(n8287), .CLK(n8701), .Q(
        test_so67), .QN(n8240) );
  SDFFX1 DFF_977_Q_reg ( .D(g29243), .SI(test_si68), .SE(n8300), .CLK(n8714), 
        .Q(g1825), .QN(n7909) );
  SDFFX1 DFF_979_Q_reg ( .D(g25623), .SI(g1825), .SE(n8301), .CLK(n8715), .Q(
        g1008), .QN(n5321) );
  SDFFX1 DFF_980_Q_reg ( .D(g26950), .SI(g1008), .SE(n8301), .CLK(n8715), .Q(
        g4392), .QN(n5710) );
  SDFFX1 DFF_981_Q_reg ( .D(test_so46), .SI(g4392), .SE(n8301), .CLK(n8715), 
        .Q(g8283) );
  SDFFX1 DFF_982_Q_reg ( .D(g30431), .SI(g8283), .SE(n8305), .CLK(n8719), .Q(
        g3546), .QN(n8050) );
  SDFFX1 DFF_983_Q_reg ( .D(g30467), .SI(g3546), .SE(n8254), .CLK(n8668), .Q(
        g5236) );
  SDFFX1 DFF_984_Q_reg ( .D(g30353), .SI(g5236), .SE(n8273), .CLK(n8687), .Q(
        g1768), .QN(n5834) );
  SDFFX1 DFF_985_Q_reg ( .D(g34467), .SI(g1768), .SE(n8350), .CLK(n8764), .Q(
        g4854) );
  SDFFX1 DFF_986_Q_reg ( .D(g30442), .SI(g4854), .SE(n8265), .CLK(n8679), .Q(
        g3925) );
  SDFFX1 DFF_987_Q_reg ( .D(g29305), .SI(g3925), .SE(n8259), .CLK(n8673), .Q(
        g6509), .QN(n7758) );
  SDFFX1 DFF_988_Q_reg ( .D(g25616), .SI(g6509), .SE(n8343), .CLK(n8757), .Q(
        g732), .QN(n5732) );
  SDFFX1 DFF_989_Q_reg ( .D(g29252), .SI(g732), .SE(n8310), .CLK(n8724), .Q(
        g2504) );
  SDFFX1 DFF_990_Q_reg ( .D(g13272), .SI(g2504), .SE(n8310), .CLK(n8724), .Q(
        test_so68), .QN(n8203) );
  SDFFX1 DFF_991_Q_reg ( .D(g4519), .SI(test_si69), .SE(n8253), .CLK(n8667), 
        .Q(g4520) );
  SDFFX1 DFF_992_Q_reg ( .D(g8916), .SI(g4520), .SE(n8253), .CLK(n8667), .Q(
        g8917), .QN(n14523) );
  SDFFX1 DFF_993_Q_reg ( .D(g33003), .SI(g8917), .SE(n8310), .CLK(n8724), .Q(
        g2185), .QN(n5376) );
  SDFFX1 DFF_994_Q_reg ( .D(g34613), .SI(g2185), .SE(n8289), .CLK(n8703), .Q(
        g37), .QN(g30327) );
  SDFFX1 DFF_995_Q_reg ( .D(g16748), .SI(g37), .SE(n8290), .CLK(n8704), .Q(
        g4031) );
  SDFFX1 DFF_996_Q_reg ( .D(g33570), .SI(g4031), .SE(n8284), .CLK(n8698), .Q(
        g2070), .QN(n5535) );
  SDFFX1 DFF_997_Q_reg ( .D(g8132), .SI(g2070), .SE(n8339), .CLK(n8753), .Q(
        g8235) );
  SDFFX1 DFF_1000_Q_reg ( .D(g34734), .SI(g8235), .SE(n8268), .CLK(n8682), .Q(
        g4176), .QN(n5494) );
  SDFFX1 DFF_1001_Q_reg ( .D(g24275), .SI(g4176), .SE(n8333), .CLK(n8747), .Q(
        g11418), .QN(n5435) );
  SDFFX1 DFF_1002_Q_reg ( .D(g7243), .SI(g11418), .SE(n8333), .CLK(n8747), .Q(
        g4405), .QN(n7671) );
  SDFFX1 DFF_1003_Q_reg ( .D(g14167), .SI(g4405), .SE(n8333), .CLK(n8747), .Q(
        g872) );
  SDFFX1 DFF_1004_Q_reg ( .D(g29302), .SI(g872), .SE(n8256), .CLK(n8670), .Q(
        g6181), .QN(n5667) );
  SDFFX1 DFF_1005_Q_reg ( .D(g24349), .SI(g6181), .SE(n8317), .CLK(n8731), .Q(
        test_so69), .QN(n8237) );
  SDFFX1 DFF_1006_Q_reg ( .D(g34264), .SI(test_si70), .SE(n8351), .CLK(n8765), 
        .Q(g4765), .QN(n5613) );
  SDFFX1 DFF_1007_Q_reg ( .D(g30484), .SI(g4765), .SE(n8249), .CLK(n8663), .Q(
        g5563), .QN(n8016) );
  SDFFX1 DFF_1008_Q_reg ( .D(g25634), .SI(g5563), .SE(n8318), .CLK(n8732), .Q(
        g1395), .QN(n8054) );
  SDFFX1 DFF_1009_Q_reg ( .D(g33567), .SI(g1395), .SE(n8345), .CLK(n8759), .Q(
        g1913) );
  SDFFX1 DFF_1010_Q_reg ( .D(g33585), .SI(g1913), .SE(n8311), .CLK(n8725), .Q(
        g2331), .QN(n5513) );
  SDFFX1 DFF_1011_Q_reg ( .D(g30527), .SI(g2331), .SE(n8336), .CLK(n8750), .Q(
        g6263) );
  SDFFX1 DFF_1012_Q_reg ( .D(g34978), .SI(g6263), .SE(n8354), .CLK(n8768), .Q(
        n9276), .QN(DFF_1012_n1) );
  SDFFX1 DFF_1013_Q_reg ( .D(g30447), .SI(n9276), .SE(n8265), .CLK(n8679), .Q(
        g3945) );
  SDFFX1 DFF_1014_Q_reg ( .D(g7540), .SI(g3945), .SE(n8309), .CLK(n8723), .Q(
        g347), .QN(n5860) );
  SDFFX1 DFF_1016_Q_reg ( .D(g34256), .SI(g347), .SE(n8266), .CLK(n8680), .Q(
        g4473), .QN(n7794) );
  SDFFX1 DFF_1017_Q_reg ( .D(g25630), .SI(g4473), .SE(n8324), .CLK(n8738), .Q(
        g1266), .QN(n7830) );
  SDFFX1 DFF_1018_Q_reg ( .D(g29290), .SI(g1266), .SE(n8353), .CLK(n8767), .Q(
        g5489), .QN(n5660) );
  SDFFX1 DFF_1019_Q_reg ( .D(g29227), .SI(g5489), .SE(n8264), .CLK(n8678), .Q(
        test_so70), .QN(n8225) );
  SDFFX1 DFF_1020_Q_reg ( .D(g31872), .SI(test_si71), .SE(n8281), .CLK(n8695), 
        .Q(g2748), .QN(n5516) );
  SDFFX1 DFF_1021_Q_reg ( .D(g29287), .SI(g2748), .SE(n8252), .CLK(n8666), .Q(
        g5471) );
  SDFFX1 DFF_1022_Q_reg ( .D(g31897), .SI(g5471), .SE(n8266), .CLK(n8680), .Q(
        g4540) );
  SDFFX1 DFF_1023_Q_reg ( .D(g17764), .SI(g4540), .SE(n8266), .CLK(n8680), .Q(
        g6723) );
  SDFFX1 DFF_1024_Q_reg ( .D(g30562), .SI(g6723), .SE(n8340), .CLK(n8754), .Q(
        g6605), .QN(n8111) );
  SDFFX1 DFF_1025_Q_reg ( .D(g34011), .SI(g6605), .SE(n8280), .CLK(n8694), .Q(
        n9274) );
  SDFFX1 DFF_1026_Q_reg ( .D(g33996), .SI(n9274), .SE(n8312), .CLK(n8726), .Q(
        g2173) );
  SDFFX1 DFF_1027_Q_reg ( .D(g21898), .SI(g2173), .SE(n8303), .CLK(n8717), .Q(
        g9019) );
  SDFFX1 DFF_1028_Q_reg ( .D(g33014), .SI(g9019), .SE(n8292), .CLK(n8706), .Q(
        g2491) );
  SDFFX1 DFF_1029_Q_reg ( .D(g34465), .SI(g2491), .SE(n8292), .CLK(n8706), .Q(
        g4849), .QN(n8151) );
  SDFFX1 DFF_1030_Q_reg ( .D(g33995), .SI(g4849), .SE(n8312), .CLK(n8726), .Q(
        g2169) );
  SDFFX1 DFF_1031_Q_reg ( .D(g30372), .SI(g2169), .SE(n8349), .CLK(n8763), .Q(
        n9273), .QN(n14522) );
  SDFFX1 DFF_1032_Q_reg ( .D(g30545), .SI(n9273), .SE(n8258), .CLK(n8672), .Q(
        test_so71) );
  SDFFX1 DFF_1033_Q_reg ( .D(g30389), .SI(test_si72), .SE(n8273), .CLK(n8687), 
        .Q(g29219) );
  SDFFX1 DFF_1034_Q_reg ( .D(g33590), .SI(g29219), .SE(n8273), .CLK(n8687), 
        .Q(g2407), .QN(n5459) );
  SDFFX1 DFF_1035_Q_reg ( .D(g34616), .SI(g2407), .SE(n8289), .CLK(n8703), .Q(
        g2868) );
  SDFFX1 DFF_1036_Q_reg ( .D(g26927), .SI(g2868), .SE(n8263), .CLK(n8677), .Q(
        g2767) );
  SDFFX1 DFF_1037_Q_reg ( .D(g32992), .SI(g2767), .SE(n8326), .CLK(n8740), .Q(
        g1783), .QN(n5596) );
  SDFFX1 DFF_1038_Q_reg ( .D(g13895), .SI(g1783), .SE(n8338), .CLK(n8752), .Q(
        g16718), .QN(n7969) );
  SDFFX1 DFF_1039_Q_reg ( .D(g25631), .SI(g16718), .SE(n8262), .CLK(n8676), 
        .Q(g1312), .QN(n5466) );
  SDFFX1 DFF_1040_Q_reg ( .D(g30477), .SI(g1312), .SE(n8302), .CLK(n8716), .Q(
        g5212) );
  SDFFX1 DFF_1041_Q_reg ( .D(g34632), .SI(g5212), .SE(n8303), .CLK(n8717), .Q(
        g4245), .QN(n5640) );
  SDFFX1 DFF_1042_Q_reg ( .D(g28046), .SI(g4245), .SE(n8344), .CLK(n8758), .Q(
        g645), .QN(n7860) );
  SDFFX1 DFF_1043_Q_reg ( .D(g9019), .SI(g645), .SE(n8303), .CLK(n8717), .Q(
        g4291), .QN(n8189) );
  SDFFX1 DFF_1044_Q_reg ( .D(g26896), .SI(g4291), .SE(n8344), .CLK(n8758), .Q(
        g29212) );
  SDFFX1 DFF_1045_Q_reg ( .D(g25602), .SI(g29212), .SE(n8344), .CLK(n8758), 
        .Q(test_so72) );
  SDFFX1 DFF_1046_Q_reg ( .D(g26916), .SI(test_si73), .SE(n8286), .CLK(n8700), 
        .Q(g1129), .QN(n5329) );
  SDFFX1 DFF_1047_Q_reg ( .D(g33578), .SI(g1129), .SE(n8260), .CLK(n8674), .Q(
        g2227), .QN(n5538) );
  SDFFX1 DFF_1049_Q_reg ( .D(g8787), .SI(g2227), .SE(n8315), .CLK(n8729), .Q(
        g8788) );
  SDFFX1 DFF_1050_Q_reg ( .D(g33579), .SI(g8788), .SE(n8309), .CLK(n8723), .Q(
        g2246), .QN(n7752) );
  SDFFX1 DFF_1051_Q_reg ( .D(g30354), .SI(g2246), .SE(n8274), .CLK(n8688), .Q(
        g1830), .QN(n5413) );
  SDFFX1 DFF_1052_Q_reg ( .D(g30425), .SI(g1830), .SE(n8306), .CLK(n8720), .Q(
        g3590) );
  SDFFX1 DFF_1053_Q_reg ( .D(g24200), .SI(g3590), .SE(n8257), .CLK(n8671), .Q(
        g392), .QN(n7865) );
  SDFFX1 DFF_1054_Q_reg ( .D(g33544), .SI(g392), .SE(n8322), .CLK(n8736), .Q(
        g1592), .QN(n5362) );
  SDFFX1 DFF_1055_Q_reg ( .D(g25764), .SI(g1592), .SE(n8329), .CLK(n8743), .Q(
        g6505), .QN(n7792) );
  SDFFX1 DFF_1057_Q_reg ( .D(g24246), .SI(g6505), .SE(n8284), .CLK(n8698), .Q(
        g1221), .QN(n8156) );
  SDFFX1 DFF_1058_Q_reg ( .D(g30507), .SI(g1221), .SE(n8337), .CLK(n8751), .Q(
        g5921) );
  SDFFX1 DFF_1059_Q_reg ( .D(g26889), .SI(g5921), .SE(n8300), .CLK(n8714), .Q(
        g29216) );
  SDFFX1 DFF_1060_Q_reg ( .D(g30333), .SI(g29216), .SE(n8351), .CLK(n8765), 
        .Q(test_so73) );
  SDFFX1 DFF_1061_Q_reg ( .D(test_so42), .SI(test_si74), .SE(n8329), .CLK(
        n8743), .Q(g218), .QN(n8138) );
  SDFFX1 DFF_1063_Q_reg ( .D(g32998), .SI(g218), .SE(n8281), .CLK(n8695), .Q(
        g1932) );
  SDFFX1 DFF_1064_Q_reg ( .D(g32987), .SI(g1932), .SE(n8347), .CLK(n8761), .Q(
        g1624), .QN(n5370) );
  SDFFX1 DFF_1065_Q_reg ( .D(g25702), .SI(g1624), .SE(n8250), .CLK(n8664), .Q(
        g5062), .QN(n7842) );
  SDFFX1 DFF_1066_Q_reg ( .D(g29286), .SI(g5062), .SE(n8252), .CLK(n8666), .Q(
        g5462), .QN(n5744) );
  SDFFX1 DFF_1067_Q_reg ( .D(g34606), .SI(g5462), .SE(n8252), .CLK(n8666), .Q(
        g2689), .QN(n5347) );
  SDFFX1 DFF_1068_Q_reg ( .D(g33070), .SI(g2689), .SE(n8313), .CLK(n8727), .Q(
        g6573), .QN(n5563) );
  SDFFX1 DFF_1069_Q_reg ( .D(g29240), .SI(g6573), .SE(n8296), .CLK(n8710), .Q(
        g1677), .QN(n7914) );
  SDFFX1 DFF_1070_Q_reg ( .D(g32999), .SI(g1677), .SE(n8284), .CLK(n8698), .Q(
        g2028), .QN(n5371) );
  SDFFX1 DFF_1071_Q_reg ( .D(g33605), .SI(g2028), .SE(n8260), .CLK(n8674), .Q(
        g2671) );
  SDFFX1 DFF_1072_Q_reg ( .D(g24255), .SI(g2671), .SE(n8314), .CLK(n8728), .Q(
        g10527) );
  SDFFX1 DFF_1073_Q_reg ( .D(g26945), .SI(g10527), .SE(n8334), .CLK(n8748), 
        .Q(g7243) );
  SDFFX1 DFF_1074_Q_reg ( .D(n8192), .SI(g7243), .SE(n8345), .CLK(n8759), .Q(
        test_so74) );
  SDFFX1 DFF_1075_Q_reg ( .D(g33558), .SI(test_si75), .SE(n8274), .CLK(n8688), 
        .Q(g1848), .QN(n5464) );
  SDFFX1 DFF_1078_Q_reg ( .D(g25699), .SI(g1848), .SE(n8248), .CLK(n8662), .Q(
        g29213), .QN(n5669) );
  SDFFX1 DFF_1079_Q_reg ( .D(g29289), .SI(g29213), .SE(n8248), .CLK(n8662), 
        .Q(g5485), .QN(n5869) );
  SDFFX1 DFF_1080_Q_reg ( .D(g30388), .SI(g5485), .SE(n8281), .CLK(n8695), .Q(
        g2741), .QN(n5349) );
  SDFFX1 DFF_1081_Q_reg ( .D(g12184), .SI(g2741), .SE(n8281), .CLK(n8695), .Q(
        g11678), .QN(n5482) );
  SDFFX1 DFF_1082_Q_reg ( .D(g29254), .SI(g11678), .SE(n8352), .CLK(n8766), 
        .Q(g2638), .QN(n7918) );
  SDFFX1 DFF_1083_Q_reg ( .D(g28074), .SI(g2638), .SE(n8267), .CLK(n8681), .Q(
        g4122), .QN(n7696) );
  SDFFX1 DFF_1084_Q_reg ( .D(g34450), .SI(g4122), .SE(n8326), .CLK(n8740), .Q(
        g4322), .QN(n5506) );
  SDFFX1 DFF_1085_Q_reg ( .D(g30512), .SI(g4322), .SE(n8351), .CLK(n8765), .Q(
        g5941) );
  SDFFX1 DFF_1086_Q_reg ( .D(g33572), .SI(g5941), .SE(n8285), .CLK(n8699), .Q(
        g2108), .QN(n5452) );
  SDFFX1 DFF_1087_Q_reg ( .D(g17646), .SI(g2108), .SE(n8285), .CLK(n8699), .Q(
        g13068) );
  SDFFX1 DFF_1088_Q_reg ( .D(g25), .SI(g13068), .SE(n8285), .CLK(n8699), .Q(
        g25) );
  SDFFX1 DFF_1089_Q_reg ( .D(g33551), .SI(g25), .SE(n8321), .CLK(n8735), .Q(
        test_so75) );
  SDFFX1 DFF_1090_Q_reg ( .D(g33538), .SI(test_si76), .SE(n8283), .CLK(n8697), 
        .Q(g595), .QN(n5476) );
  SDFFX1 DFF_1091_Q_reg ( .D(g33005), .SI(g595), .SE(n8310), .CLK(n8724), .Q(
        g2217), .QN(n5512) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24248), .SI(g2217), .SE(n8254), .CLK(n8668), .Q(
        n9267), .QN(DFF_1092_n1) );
  SDFFX1 DFF_1093_Q_reg ( .D(g33002), .SI(n9267), .SE(n8339), .CLK(n8753), .Q(
        g2066), .QN(n5832) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24234), .SI(g2066), .SE(n8339), .CLK(n8753), .Q(
        g1152), .QN(n5618) );
  SDFFX1 DFF_1095_Q_reg ( .D(g30471), .SI(g1152), .SE(n8254), .CLK(n8668), .Q(
        g5252) );
  SDFFX1 DFF_1096_Q_reg ( .D(g34000), .SI(g5252), .SE(n8311), .CLK(n8725), .Q(
        g2165) );
  SDFFX1 DFF_1097_Q_reg ( .D(g34016), .SI(g2165), .SE(n8304), .CLK(n8718), .Q(
        g2571) );
  SDFFX1 DFF_1098_Q_reg ( .D(g33048), .SI(g2571), .SE(n8304), .CLK(n8718), .Q(
        g5176), .QN(n5650) );
  SDFFX1 DFF_1100_Q_reg ( .D(g8283), .SI(g5176), .SE(n8304), .CLK(n8718), .Q(
        g8403) );
  SDFFX1 DFF_1102_Q_reg ( .D(g17819), .SI(g8403), .SE(n8304), .CLK(n8718), .Q(
        g14673) );
  SDFFX1 DFF_1103_Q_reg ( .D(g25628), .SI(g14673), .SE(n8284), .CLK(n8698), 
        .Q(test_so76), .QN(n8212) );
  SDFFX1 DFF_1104_Q_reg ( .D(g26934), .SI(test_si77), .SE(n8280), .CLK(n8694), 
        .Q(g2827) );
  SDFFX1 DFF_1106_Q_reg ( .D(g14201), .SI(g2827), .SE(n8300), .CLK(n8714), .Q(
        g14217) );
  SDFFX1 DFF_1107_Q_reg ( .D(g34468), .SI(g14217), .SE(n8298), .CLK(n8712), 
        .Q(g4859) );
  SDFFX1 DFF_1108_Q_reg ( .D(g24202), .SI(g4859), .SE(n8257), .CLK(n8671), .Q(
        g424), .QN(n7833) );
  SDFFX1 DFF_1109_Q_reg ( .D(g33542), .SI(g424), .SE(n8314), .CLK(n8728), .Q(
        g1274), .QN(n5730) );
  SDFFX1 DFF_1110_Q_reg ( .D(g17404), .SI(g1274), .SE(n8314), .CLK(n8728), .Q(
        g17423), .QN(n7822) );
  SDFFX1 DFF_1111_Q_reg ( .D(g33435), .SI(g17423), .SE(n8353), .CLK(n8767), 
        .Q(n9265) );
  SDFFX1 DFF_1112_Q_reg ( .D(g34445), .SI(n9265), .SE(n8261), .CLK(n8675), .Q(
        g2803), .QN(n5545) );
  SDFFX1 DFF_1114_Q_reg ( .D(g33555), .SI(g2803), .SE(n8274), .CLK(n8688), .Q(
        g1821), .QN(n7747) );
  SDFFX1 DFF_1115_Q_reg ( .D(g34013), .SI(g1821), .SE(n8308), .CLK(n8722), .Q(
        g2509), .QN(n7784) );
  SDFFX1 DFF_1116_Q_reg ( .D(g28091), .SI(g2509), .SE(n8308), .CLK(n8722), .Q(
        g5073), .QN(n7781) );
  SDFFX1 DFF_1117_Q_reg ( .D(g26919), .SI(g5073), .SE(n8324), .CLK(n8738), .Q(
        test_so77), .QN(n5556) );
  SDFFX1 DFF_1118_Q_reg ( .D(g8235), .SI(test_si78), .SE(n8339), .CLK(n8753), 
        .Q(g8353) );
  SDFFX1 DFF_1119_Q_reg ( .D(g17685), .SI(g8353), .SE(n8340), .CLK(n8754), .Q(
        g13085) );
  SDFFX1 DFF_1120_Q_reg ( .D(g30554), .SI(g13085), .SE(n8340), .CLK(n8754), 
        .Q(g6633) );
  SDFFX1 DFF_1121_Q_reg ( .D(g29281), .SI(g6633), .SE(n8268), .CLK(n8682), .Q(
        g5124), .QN(n7709) );
  SDFFX1 DFF_1122_Q_reg ( .D(test_so44), .SI(g5124), .SE(n8330), .CLK(n8744), 
        .Q(g17400), .QN(n7811) );
  SDFFX1 DFF_1123_Q_reg ( .D(g30537), .SI(g17400), .SE(n8351), .CLK(n8765), 
        .Q(g6303) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28092), .SI(g6303), .SE(n8248), .CLK(n8662), .Q(
        g5069), .QN(n7780) );
  SDFFX1 DFF_1125_Q_reg ( .D(g34732), .SI(g5069), .SE(n8289), .CLK(n8703), .Q(
        g2994), .QN(n5634) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28049), .SI(g2994), .SE(n8344), .CLK(n8758), .Q(
        g650), .QN(n7861) );
  SDFFX1 DFF_1127_Q_reg ( .D(g33545), .SI(g650), .SE(n8321), .CLK(n8735), .Q(
        g1636), .QN(n5549) );
  SDFFX1 DFF_1128_Q_reg ( .D(g30441), .SI(g1636), .SE(n8323), .CLK(n8737), .Q(
        g3921) );
  SDFFX1 DFF_1129_Q_reg ( .D(g29247), .SI(g3921), .SE(n8285), .CLK(n8699), .Q(
        test_so78) );
  SDFFX1 DFF_1130_Q_reg ( .D(g24354), .SI(test_si79), .SE(n8266), .CLK(n8680), 
        .Q(g6732), .QN(n8125) );
  SDFFX1 DFF_1131_Q_reg ( .D(g25636), .SI(g6732), .SE(n8347), .CLK(n8761), .Q(
        g1306), .QN(n5796) );
  SDFFX1 DFF_1133_Q_reg ( .D(g26914), .SI(g1306), .SE(n8295), .CLK(n8709), .Q(
        g1061), .QN(n7840) );
  SDFFX1 DFF_1134_Q_reg ( .D(g25670), .SI(g1061), .SE(n8295), .CLK(n8709), .Q(
        g3462), .QN(n7777) );
  SDFFX1 DFF_1135_Q_reg ( .D(g33998), .SI(g3462), .SE(n8312), .CLK(n8726), .Q(
        g2181), .QN(n5803) );
  SDFFX1 DFF_1136_Q_reg ( .D(g25626), .SI(g2181), .SE(n8291), .CLK(n8705), .Q(
        g956), .QN(n5341) );
  SDFFX1 DFF_1137_Q_reg ( .D(g33977), .SI(g956), .SE(n8273), .CLK(n8687), .Q(
        g1756), .QN(n5804) );
  SDFFX1 DFF_1138_Q_reg ( .D(g29297), .SI(g1756), .SE(n8335), .CLK(n8749), .Q(
        g5849) );
  SDFFX1 DFF_1139_Q_reg ( .D(g28071), .SI(g5849), .SE(n8267), .CLK(n8681), .Q(
        g4112) );
  SDFFX1 DFF_1140_Q_reg ( .D(g30387), .SI(g4112), .SE(n8260), .CLK(n8674), .Q(
        n9262), .QN(n14517) );
  SDFFX1 DFF_1141_Q_reg ( .D(g33577), .SI(n9262), .SE(n8260), .CLK(n8674), .Q(
        g2197), .QN(n5514) );
  SDFFX1 DFF_1143_Q_reg ( .D(g33592), .SI(g2197), .SE(n8310), .CLK(n8724), .Q(
        test_so79), .QN(n8204) );
  SDFFX1 DFF_1144_Q_reg ( .D(g26913), .SI(test_si80), .SE(n8263), .CLK(n8677), 
        .Q(g1046) );
  SDFFX1 DFF_1145_Q_reg ( .D(g28044), .SI(g1046), .SE(n8323), .CLK(n8737), .Q(
        g482), .QN(n5820) );
  SDFFX1 DFF_1146_Q_reg ( .D(g26948), .SI(g482), .SE(n8323), .CLK(n8737), .Q(
        g4401) );
  SDFFX1 DFF_1148_Q_reg ( .D(g30344), .SI(g4401), .SE(n8323), .CLK(n8737), .Q(
        g1514), .QN(n5364) );
  SDFFX1 DFF_1149_Q_reg ( .D(g26885), .SI(g1514), .SE(n8313), .CLK(n8727), .Q(
        g329), .QN(n5766) );
  SDFFX1 DFF_1150_Q_reg ( .D(g33069), .SI(g329), .SE(n8313), .CLK(n8727), .Q(
        g6565), .QN(n5386) );
  SDFFX1 DFF_1151_Q_reg ( .D(g34621), .SI(g6565), .SE(n8271), .CLK(n8685), .Q(
        g2950), .QN(n8170) );
  SDFFX1 DFF_1153_Q_reg ( .D(g28059), .SI(g2950), .SE(n8261), .CLK(n8675), .Q(
        g1345), .QN(n7836) );
  SDFFX1 DFF_1154_Q_reg ( .D(g25762), .SI(g1345), .SE(n8329), .CLK(n8743), .Q(
        g6533), .QN(n5445) );
  SDFFX1 DFF_1155_Q_reg ( .D(g16624), .SI(g6533), .SE(n8338), .CLK(n8752), .Q(
        g14421) );
  SDFFX1 DFF_1157_Q_reg ( .D(g34633), .SI(g14421), .SE(n8338), .CLK(n8752), 
        .Q(g4727), .QN(n5312) );
  SDFFX1 DFF_1158_Q_reg ( .D(g24352), .SI(g4727), .SE(n8346), .CLK(n8760), .Q(
        test_so80), .QN(n8231) );
  SDFFX1 DFF_1159_Q_reg ( .D(g26925), .SI(test_si81), .SE(n8262), .CLK(n8676), 
        .Q(g1536) );
  SDFFX1 DFF_1160_Q_reg ( .D(g30446), .SI(g1536), .SE(n8265), .CLK(n8679), .Q(
        g3941) );
  SDFFX1 DFF_1161_Q_reg ( .D(g25597), .SI(g3941), .SE(n8307), .CLK(n8721), .Q(
        g370), .QN(n7874) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24342), .SI(g370), .SE(n8271), .CLK(n8685), .Q(
        g5694), .QN(n7992) );
  SDFFX1 DFF_1163_Q_reg ( .D(g30357), .SI(g5694), .SE(n8274), .CLK(n8688), .Q(
        g1858), .QN(n5892) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26908), .SI(g1858), .SE(n8274), .CLK(n8688), .Q(
        g446) );
  SDFFX1 DFF_1166_Q_reg ( .D(g30399), .SI(g446), .SE(n8328), .CLK(n8742), .Q(
        g3219) );
  SDFFX1 DFF_1167_Q_reg ( .D(g29242), .SI(g3219), .SE(n8300), .CLK(n8714), .Q(
        g1811) );
  SDFFX1 DFF_1169_Q_reg ( .D(g30547), .SI(g1811), .SE(n8340), .CLK(n8754), .Q(
        g6601), .QN(n8022) );
  SDFFX1 DFF_1171_Q_reg ( .D(g34010), .SI(g6601), .SE(n8280), .CLK(n8694), .Q(
        g2441) );
  SDFFX1 DFF_1172_Q_reg ( .D(g33986), .SI(g2441), .SE(n8286), .CLK(n8700), .Q(
        g1874) );
  SDFFX1 DFF_1173_Q_reg ( .D(g34257), .SI(g1874), .SE(n8301), .CLK(n8715), .Q(
        test_so81), .QN(n8208) );
  SDFFX1 DFF_1174_Q_reg ( .D(g30544), .SI(test_si82), .SE(n8328), .CLK(n8742), 
        .Q(g6581), .QN(n8049) );
  SDFFX1 DFF_1175_Q_reg ( .D(g30561), .SI(g6581), .SE(n8329), .CLK(n8743), .Q(
        g6597) );
  SDFFX1 DFF_1176_Q_reg ( .D(g8403), .SI(g6597), .SE(n8329), .CLK(n8743), .Q(
        g5008), .QN(n5637) );
  SDFFX1 DFF_1177_Q_reg ( .D(g30430), .SI(g5008), .SE(n8350), .CLK(n8764), .Q(
        g3610) );
  SDFFX1 DFF_1178_Q_reg ( .D(g34799), .SI(g3610), .SE(n8289), .CLK(n8703), .Q(
        g2890), .QN(n8178) );
  SDFFX1 DFF_1179_Q_reg ( .D(g33565), .SI(g2890), .SE(n8271), .CLK(n8685), .Q(
        g1978) );
  SDFFX1 DFF_1180_Q_reg ( .D(g33968), .SI(g1978), .SE(n8263), .CLK(n8677), .Q(
        g1612) );
  SDFFX1 DFF_1181_Q_reg ( .D(g34843), .SI(g1612), .SE(n8311), .CLK(n8725), .Q(
        g112), .QN(n7866) );
  SDFFX1 DFF_1182_Q_reg ( .D(g34793), .SI(g112), .SE(n8255), .CLK(n8669), .Q(
        g2856) );
  SDFFX1 DFF_1184_Q_reg ( .D(g33566), .SI(g2856), .SE(n8272), .CLK(n8686), .Q(
        g1982), .QN(n5462) );
  SDFFX1 DFF_1185_Q_reg ( .D(g17688), .SI(g1982), .SE(n8319), .CLK(n8733), .Q(
        g17722), .QN(n8083) );
  SDFFX1 DFF_1186_Q_reg ( .D(g30465), .SI(g17722), .SE(n8302), .CLK(n8716), 
        .Q(test_so82) );
  SDFFX1 DFF_1187_Q_reg ( .D(g28073), .SI(test_si83), .SE(n8267), .CLK(n8681), 
        .Q(g4119) );
  SDFFX1 DFF_1188_Q_reg ( .D(g24351), .SI(g4119), .SE(n8317), .CLK(n8731), .Q(
        g6390), .QN(n7986) );
  SDFFX1 DFF_1189_Q_reg ( .D(g30346), .SI(g6390), .SE(n8262), .CLK(n8676), .Q(
        g1542), .QN(n7862) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21893), .SI(g1542), .SE(n8262), .CLK(n8676), .Q(
        g4258) );
  SDFFX1 DFF_1191_Q_reg ( .D(g8353), .SI(g4258), .SE(n8339), .CLK(n8753), .Q(
        g4818), .QN(n5636) );
  SDFFX1 DFF_1192_Q_reg ( .D(g31904), .SI(g4818), .SE(n8250), .CLK(n8664), .Q(
        g5033), .QN(n7838) );
  SDFFX1 DFF_1193_Q_reg ( .D(g34635), .SI(g5033), .SE(n8338), .CLK(n8752), .Q(
        g4717), .QN(n5344) );
  SDFFX1 DFF_1194_Q_reg ( .D(g25637), .SI(g4717), .SE(n8313), .CLK(n8727), .Q(
        g1554), .QN(n5768) );
  SDFFX1 DFF_1195_Q_reg ( .D(g29274), .SI(g1554), .SE(n8335), .CLK(n8749), .Q(
        g3849) );
  SDFFX1 DFF_1196_Q_reg ( .D(g14828), .SI(g3849), .SE(n8319), .CLK(n8733), .Q(
        g17778), .QN(n7978) );
  SDFFX1 DFF_1197_Q_reg ( .D(g30396), .SI(g17778), .SE(n8319), .CLK(n8733), 
        .Q(g3199), .QN(n8097) );
  SDFFX1 DFF_1198_Q_reg ( .D(g25735), .SI(g3199), .SE(n8353), .CLK(n8767), .Q(
        test_so83), .QN(n8233) );
  SDFFX1 DFF_1199_Q_reg ( .D(g34037), .SI(test_si84), .SE(n8298), .CLK(n8712), 
        .Q(g4975), .QN(n5360) );
  SDFFX1 DFF_1200_Q_reg ( .D(g34791), .SI(g4975), .SE(n8299), .CLK(n8713), .Q(
        g790), .QN(n5292) );
  SDFFX1 DFF_1201_Q_reg ( .D(g30520), .SI(g790), .SE(n8288), .CLK(n8702), .Q(
        g5913), .QN(n8099) );
  SDFFX1 DFF_1202_Q_reg ( .D(g30358), .SI(g5913), .SE(n8282), .CLK(n8696), .Q(
        g1902), .QN(n5837) );
  SDFFX1 DFF_1203_Q_reg ( .D(g29299), .SI(g1902), .SE(n8256), .CLK(n8670), .Q(
        g6163), .QN(n7738) );
  SDFFX1 DFF_1204_Q_reg ( .D(g25690), .SI(g6163), .SE(n8325), .CLK(n8739), .Q(
        g4125), .QN(n8122) );
  SDFFX1 DFF_1205_Q_reg ( .D(g28096), .SI(g4125), .SE(n8250), .CLK(n8664), .Q(
        g4821) );
  SDFFX1 DFF_1206_Q_reg ( .D(g28088), .SI(g4821), .SE(n8295), .CLK(n8709), .Q(
        g4939), .QN(n5776) );
  SDFFX1 DFF_1207_Q_reg ( .D(g24241), .SI(g4939), .SE(n8295), .CLK(n8709), .Q(
        g19334), .QN(n5392) );
  SDFFX1 DFF_1208_Q_reg ( .D(g30397), .SI(g19334), .SE(n8320), .CLK(n8734), 
        .Q(g3207), .QN(n8007) );
  SDFFX1 DFF_1209_Q_reg ( .D(g4520), .SI(g3207), .SE(n8320), .CLK(n8734), .Q(
        g4483) );
  SDFFX1 DFF_1210_Q_reg ( .D(g30409), .SI(g4483), .SE(n8320), .CLK(n8734), .Q(
        test_so84) );
  SDFFX1 DFF_1211_Q_reg ( .D(g29284), .SI(test_si85), .SE(n8269), .CLK(n8683), 
        .Q(g5142), .QN(n5658) );
  SDFFX1 DFF_1212_Q_reg ( .D(g30470), .SI(g5142), .SE(n8253), .CLK(n8667), .Q(
        g5248) );
  SDFFX1 DFF_1213_Q_reg ( .D(g30367), .SI(g5248), .SE(n8279), .CLK(n8693), .Q(
        g2126) );
  SDFFX1 DFF_1214_Q_reg ( .D(g24273), .SI(g2126), .SE(n8279), .CLK(n8693), .Q(
        g3694), .QN(n7990) );
  SDFFX1 DFF_1215_Q_reg ( .D(g29288), .SI(g3694), .SE(n8271), .CLK(n8685), .Q(
        g5481), .QN(n5805) );
  SDFFX1 DFF_1216_Q_reg ( .D(g30359), .SI(g5481), .SE(n8271), .CLK(n8685), .Q(
        g1964), .QN(n5315) );
  SDFFX1 DFF_1217_Q_reg ( .D(g25698), .SI(g1964), .SE(n8248), .CLK(n8662), .Q(
        g5097), .QN(n5753) );
  SDFFX1 DFF_1218_Q_reg ( .D(g30398), .SI(g5097), .SE(n8328), .CLK(n8742), .Q(
        g3215) );
  SDFFX1 DFF_1219_Q_reg ( .D(g13906), .SI(g3215), .SE(n8333), .CLK(n8747), .Q(
        g16748) );
  SDFFX1 DFF_1220_Q_reg ( .D(g33079), .SI(g16748), .SE(n8333), .CLK(n8747), 
        .Q(n9255) );
  SDFFX1 DFF_1221_Q_reg ( .D(g26952), .SI(n9255), .SE(n8277), .CLK(n8691), .Q(
        g4427), .QN(n7856) );
  SDFFX1 DFF_1222_Q_reg ( .D(g34974), .SI(g4427), .SE(n8277), .CLK(n8691), .Q(
        test_so85), .QN(n8219) );
  SDFFX1 DFF_1223_Q_reg ( .D(g26928), .SI(test_si86), .SE(n8273), .CLK(n8687), 
        .Q(g2779) );
  SDFFX1 DFF_1224_Q_reg ( .D(test_so39), .SI(g2779), .SE(n8315), .CLK(n8729), 
        .Q(g8786), .QN(n5694) );
  SDFFX1 DFF_1225_Q_reg ( .D(g26954), .SI(g8786), .SE(n8309), .CLK(n8723), .Q(
        g7245), .QN(DFF_1225_n1) );
  SDFFX1 DFF_1226_Q_reg ( .D(g30351), .SI(g7245), .SE(n8352), .CLK(n8766), .Q(
        g1720), .QN(n5780) );
  SDFFX1 DFF_1227_Q_reg ( .D(g31871), .SI(g1720), .SE(n8261), .CLK(n8675), .Q(
        g1367), .QN(n7814) );
  SDFFX1 DFF_1228_Q_reg ( .D(g9553), .SI(g1367), .SE(n8317), .CLK(n8731), .Q(
        g5112) );
  SDFFX1 DFF_1229_Q_reg ( .D(g34978), .SI(g5112), .SE(n8267), .CLK(n8681), .Q(
        g19), .QN(n7685) );
  SDFFX1 DFF_1230_Q_reg ( .D(g26939), .SI(g19), .SE(n8267), .CLK(n8681), .Q(
        g4145), .QN(n8160) );
  SDFFX1 DFF_1231_Q_reg ( .D(g33994), .SI(g4145), .SE(n8312), .CLK(n8726), .Q(
        g2161), .QN(n5812) );
  SDFFX1 DFF_1232_Q_reg ( .D(g25596), .SI(g2161), .SE(n8312), .CLK(n8726), .Q(
        g376), .QN(n5633) );
  SDFFX1 DFF_1233_Q_reg ( .D(g33586), .SI(g376), .SE(n8311), .CLK(n8725), .Q(
        g2361), .QN(n5537) );
  SDFFX1 DFF_1234_Q_reg ( .D(g21901), .SI(g2361), .SE(n8303), .CLK(n8717), .Q(
        test_so86) );
  SDFFX1 DFF_1235_Q_reg ( .D(g31866), .SI(test_si87), .SE(n8283), .CLK(n8697), 
        .Q(g582), .QN(n5552) );
  SDFFX1 DFF_1236_Q_reg ( .D(g33000), .SI(g582), .SE(n8284), .CLK(n8698), .Q(
        g2051), .QN(n8129) );
  SDFFX1 DFF_1237_Q_reg ( .D(g26918), .SI(g2051), .SE(n8254), .CLK(n8668), .Q(
        g1193) );
  SDFFX1 DFF_1240_Q_reg ( .D(g30373), .SI(g1193), .SE(n8288), .CLK(n8702), .Q(
        g2327), .QN(n5841) );
  SDFFX1 DFF_1241_Q_reg ( .D(g28056), .SI(g2327), .SE(n8275), .CLK(n8689), .Q(
        g907), .QN(n5555) );
  SDFFX1 DFF_1242_Q_reg ( .D(g34601), .SI(g907), .SE(n8275), .CLK(n8689), .Q(
        g947), .QN(n5286) );
  SDFFX1 DFF_1243_Q_reg ( .D(g30355), .SI(g947), .SE(n8274), .CLK(n8688), .Q(
        g1834), .QN(n5665) );
  SDFFX1 DFF_1244_Q_reg ( .D(g30426), .SI(g1834), .SE(n8350), .CLK(n8764), .Q(
        g3594) );
  SDFFX1 DFF_1245_Q_reg ( .D(g34805), .SI(g3594), .SE(n8289), .CLK(n8703), .Q(
        g2999), .QN(n8180) );
  SDFFX1 DFF_1247_Q_reg ( .D(g34002), .SI(g2999), .SE(n8287), .CLK(n8701), .Q(
        g2303) );
  SDFFX1 DFF_1248_Q_reg ( .D(g17778), .SI(g2303), .SE(n8319), .CLK(n8733), .Q(
        g17688), .QN(n7964) );
  SDFFX1 DFF_1250_Q_reg ( .D(g28053), .SI(g17688), .SE(n8344), .CLK(n8758), 
        .Q(test_so87) );
  SDFFX1 DFF_1251_Q_reg ( .D(g29229), .SI(test_si88), .SE(n8342), .CLK(n8756), 
        .Q(g723), .QN(n5826) );
  SDFFX1 DFF_1252_Q_reg ( .D(g33620), .SI(g723), .SE(n8271), .CLK(n8685), .Q(
        g5703), .QN(n5397) );
  SDFFX1 DFF_1253_Q_reg ( .D(g34722), .SI(g5703), .SE(n8277), .CLK(n8691), .Q(
        g546), .QN(n5492) );
  SDFFX1 DFF_1254_Q_reg ( .D(g33599), .SI(g546), .SE(n8348), .CLK(n8762), .Q(
        g2472), .QN(n5619) );
  SDFFX1 DFF_1255_Q_reg ( .D(g30515), .SI(g2472), .SE(n8348), .CLK(n8762), .Q(
        g5953) );
  SDFFX1 DFF_1256_Q_reg ( .D(g25649), .SI(g5953), .SE(n8272), .CLK(n8686), .Q(
        g8277), .QN(n7742) );
  SDFFX1 DFF_1258_Q_reg ( .D(g33979), .SI(g8277), .SE(n8272), .CLK(n8686), .Q(
        g1740) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30417), .SI(g1740), .SE(n8306), .CLK(n8720), .Q(
        g3550), .QN(n8117) );
  SDFFX1 DFF_1260_Q_reg ( .D(g25683), .SI(g3550), .SE(n8278), .CLK(n8692), .Q(
        g3845), .QN(n5886) );
  SDFFX1 DFF_1261_Q_reg ( .D(g33574), .SI(g3845), .SE(n8278), .CLK(n8692), .Q(
        g2116), .QN(n5463) );
  SDFFX1 DFF_1262_Q_reg ( .D(g17813), .SI(g2116), .SE(n8319), .CLK(n8733), .Q(
        g14635) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30410), .SI(g14635), .SE(n8328), .CLK(n8742), 
        .Q(test_so88) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30454), .SI(test_si89), .SE(n8265), .CLK(n8679), 
        .Q(g3913), .QN(n8107) );
  SDFFX1 DFF_1265_Q_reg ( .D(g34024), .SI(g3913), .SE(n8341), .CLK(n8755), .Q(
        g10306) );
  SDFFX1 DFF_1266_Q_reg ( .D(g33547), .SI(g10306), .SE(n8346), .CLK(n8760), 
        .Q(g1687), .QN(n7751) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30386), .SI(g1687), .SE(n8260), .CLK(n8674), .Q(
        g2681), .QN(n5777) );
  SDFFX1 DFF_1268_Q_reg ( .D(g33596), .SI(g2681), .SE(n8308), .CLK(n8722), .Q(
        g2533), .QN(n5761) );
  SDFFX1 DFF_1269_Q_reg ( .D(g26887), .SI(g2533), .SE(n8308), .CLK(n8722), .Q(
        g324), .QN(n5827) );
  SDFFX1 DFF_1270_Q_reg ( .D(g34607), .SI(g324), .SE(n8308), .CLK(n8722), .Q(
        g2697), .QN(n5308) );
  SDFFX1 DFF_1272_Q_reg ( .D(g31895), .SI(g2697), .SE(n8308), .CLK(n8722), .Q(
        g4417), .QN(n7675) );
  SDFFX1 DFF_1273_Q_reg ( .D(g33068), .SI(g4417), .SE(n8326), .CLK(n8740), .Q(
        g6561), .QN(n5646) );
  SDFFX1 DFF_1274_Q_reg ( .D(g29233), .SI(g6561), .SE(n8291), .CLK(n8705), .Q(
        g1141), .QN(n5691) );
  SDFFX1 DFF_1275_Q_reg ( .D(g24258), .SI(g1141), .SE(n8314), .CLK(n8728), .Q(
        g12923), .QN(n5655) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30376), .SI(g12923), .SE(n8273), .CLK(n8687), 
        .Q(test_so89), .QN(n8234) );
  SDFFX1 DFF_1277_Q_reg ( .D(g33549), .SI(test_si90), .SE(n8296), .CLK(n8710), 
        .Q(g1710) );
  SDFFX1 DFF_1278_Q_reg ( .D(g29308), .SI(g1710), .SE(n8259), .CLK(n8673), .Q(
        g6527), .QN(n5659) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30408), .SI(g6527), .SE(n8319), .CLK(n8733), .Q(
        g3255) );
  SDFFX1 DFF_1281_Q_reg ( .D(g29241), .SI(g3255), .SE(n8296), .CLK(n8710), .Q(
        g1691), .QN(n7913) );
  SDFFX1 DFF_1282_Q_reg ( .D(g34620), .SI(g1691), .SE(n8270), .CLK(n8684), .Q(
        g2936), .QN(n8171) );
  SDFFX1 DFF_1283_Q_reg ( .D(g33621), .SI(g2936), .SE(n8252), .CLK(n8666), .Q(
        g5644), .QN(n5593) );
  SDFFX1 DFF_1284_Q_reg ( .D(g25707), .SI(g5644), .SE(n8269), .CLK(n8683), .Q(
        g5152), .QN(n5883) );
  SDFFX1 DFF_1285_Q_reg ( .D(g24339), .SI(g5152), .SE(n8269), .CLK(n8683), .Q(
        g5352), .QN(n8126) );
  SDFFX1 DFF_1286_Q_reg ( .D(g11770), .SI(g5352), .SE(n8269), .CLK(n8683), .Q(
        g8915) );
  SDFFX1 DFF_1288_Q_reg ( .D(g34443), .SI(g8915), .SE(n8273), .CLK(n8687), .Q(
        g2775), .QN(n5378) );
  SDFFX1 DFF_1289_Q_reg ( .D(g34619), .SI(g2775), .SE(n8270), .CLK(n8684), .Q(
        g2922), .QN(n8169) );
  SDFFX1 DFF_1290_Q_reg ( .D(g29234), .SI(g2922), .SE(n8294), .CLK(n8708), .Q(
        test_so90) );
  SDFFX1 DFF_1291_Q_reg ( .D(g30503), .SI(test_si91), .SE(n8337), .CLK(n8751), 
        .Q(g5893), .QN(n7901) );
  SDFFX1 DFF_1293_Q_reg ( .D(g16718), .SI(g5893), .SE(n8338), .CLK(n8752), .Q(
        g16603), .QN(n7954) );
  SDFFX1 DFF_1294_Q_reg ( .D(g30550), .SI(g16603), .SE(n8339), .CLK(n8753), 
        .Q(g6617) );
  SDFFX1 DFF_1295_Q_reg ( .D(g33001), .SI(g6617), .SE(n8339), .CLK(n8753), .Q(
        g2060), .QN(n5507) );
  SDFFX1 DFF_1296_Q_reg ( .D(g33040), .SI(g2060), .SE(n8339), .CLK(n8753), .Q(
        g4512) );
  SDFFX1 DFF_1297_Q_reg ( .D(g30492), .SI(g4512), .SE(n8249), .CLK(n8663), .Q(
        g5599) );
  SDFFX1 DFF_1298_Q_reg ( .D(g25664), .SI(g5599), .SE(n8252), .CLK(n8666), .Q(
        g3401), .QN(n5986) );
  SDFFX1 DFF_1299_Q_reg ( .D(g26944), .SI(g3401), .SE(n8332), .CLK(n8746), .Q(
        g4366), .QN(n8000) );
  SDFFX1 DFF_1300_Q_reg ( .D(test_so26), .SI(g4366), .SE(n8332), .CLK(n8746), 
        .Q(g16722) );
  SDFFX1 DFF_1301_Q_reg ( .D(g34614), .SI(g16722), .SE(n8332), .CLK(n8746), 
        .Q(g29214) );
  SDFFX1 DFF_1302_Q_reg ( .D(g29260), .SI(g29214), .SE(n8269), .CLK(n8683), 
        .Q(g3129), .QN(n5861) );
  SDFFX1 DFF_1303_Q_reg ( .D(g16686), .SI(g3129), .SE(n8321), .CLK(n8735), .Q(
        test_so91) );
  SDFFX1 DFF_1304_Q_reg ( .D(g33047), .SI(test_si92), .SE(n8318), .CLK(n8732), 
        .Q(g5170), .QN(n8140) );
  SDFFX1 DFF_1305_Q_reg ( .D(g24298), .SI(g5170), .SE(n8301), .CLK(n8715), .Q(
        g26959) );
  SDFFX1 DFF_1306_Q_reg ( .D(g25733), .SI(g26959), .SE(n8285), .CLK(n8699), 
        .Q(g5821), .QN(n5429) );
  SDFFX1 DFF_1307_Q_reg ( .D(g30536), .SI(g5821), .SE(n8298), .CLK(n8712), .Q(
        g6299) );
  SDFFX1 DFF_1308_Q_reg ( .D(g7916), .SI(g6299), .SE(n8332), .CLK(n8746), .Q(
        g8416), .QN(n7730) );
  SDFFX1 DFF_1310_Q_reg ( .D(g29246), .SI(g8416), .SE(n8285), .CLK(n8699), .Q(
        g2079), .QN(n7915) );
  SDFFX1 DFF_1311_Q_reg ( .D(g34261), .SI(g2079), .SE(n8269), .CLK(n8683), .Q(
        g4698), .QN(n5862) );
  SDFFX1 DFF_1312_Q_reg ( .D(g33611), .SI(g4698), .SE(n8327), .CLK(n8741), .Q(
        g3703), .QN(n5399) );
  SDFFX1 DFF_1313_Q_reg ( .D(g25638), .SI(g3703), .SE(n8313), .CLK(n8727), .Q(
        g1559), .QN(n5441) );
  SDFFX1 DFF_1314_Q_reg ( .D(g34728), .SI(g1559), .SE(n8353), .CLK(n8767), .Q(
        n9247), .QN(n14520) );
  SDFFX1 DFF_1315_Q_reg ( .D(g29222), .SI(n9247), .SE(n8257), .CLK(n8671), .Q(
        g411), .QN(n5629) );
  SDFFX1 DFF_1316_Q_reg ( .D(g25742), .SI(g411), .SE(n8337), .CLK(n8751), .Q(
        test_so92) );
  SDFFX1 DFF_1317_Q_reg ( .D(g30449), .SI(test_si93), .SE(n8343), .CLK(n8757), 
        .Q(g3953) );
  SDFFX1 DFF_1319_Q_reg ( .D(g34608), .SI(g3953), .SE(n8343), .CLK(n8757), .Q(
        g2704), .QN(n5377) );
  SDFFX1 DFF_1320_Q_reg ( .D(g24345), .SI(g2704), .SE(n8307), .CLK(n8721), .Q(
        g6035), .QN(n5528) );
  SDFFX1 DFF_1322_Q_reg ( .D(g34977), .SI(g6035), .SE(n8307), .CLK(n8721), .Q(
        n9245) );
  SDFFX1 DFF_1323_Q_reg ( .D(g25635), .SI(n9245), .SE(n8307), .CLK(n8721), .Q(
        g1300), .QN(n5483) );
  SDFFX1 DFF_1324_Q_reg ( .D(g25686), .SI(g1300), .SE(n8325), .CLK(n8739), .Q(
        g4057), .QN(n5711) );
  SDFFX1 DFF_1325_Q_reg ( .D(g30461), .SI(g4057), .SE(n8302), .CLK(n8716), .Q(
        g5200), .QN(n7899) );
  SDFFX1 DFF_1326_Q_reg ( .D(g34466), .SI(g5200), .SE(n8350), .CLK(n8764), .Q(
        g4843), .QN(n7796) );
  SDFFX1 DFF_1327_Q_reg ( .D(g31901), .SI(g4843), .SE(n8251), .CLK(n8665), .Q(
        g5046), .QN(n5578) );
  SDFFX1 DFF_1328_Q_reg ( .D(g29249), .SI(g5046), .SE(n8312), .CLK(n8726), .Q(
        g2250), .QN(n7907) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26882), .SI(g2250), .SE(n8312), .CLK(n8726), .Q(
        g26885), .QN(n5456) );
  SDFFX1 DFF_1330_Q_reg ( .D(g33041), .SI(g26885), .SE(n8337), .CLK(n8751), 
        .Q(test_so93) );
  SDFFX1 DFF_1331_Q_reg ( .D(g33011), .SI(test_si94), .SE(n8331), .CLK(n8745), 
        .Q(g2453), .QN(n5373) );
  SDFFX1 DFF_1332_Q_reg ( .D(g25734), .SI(g2453), .SE(n8286), .CLK(n8700), .Q(
        g5841), .QN(n5449) );
  SDFFX1 DFF_1335_Q_reg ( .D(g12300), .SI(g5841), .SE(n8286), .CLK(n8700), .Q(
        g14694), .QN(n5705) );
  SDFFX1 DFF_1336_Q_reg ( .D(g34618), .SI(g14694), .SE(n8270), .CLK(n8684), 
        .Q(g2912) );
  SDFFX1 DFF_1337_Q_reg ( .D(g33010), .SI(g2912), .SE(n8294), .CLK(n8708), .Q(
        g2357) );
  SDFFX1 DFF_1338_Q_reg ( .D(g8919), .SI(g2357), .SE(n8311), .CLK(n8725), .Q(
        g8920) );
  SDFFX1 DFF_1339_Q_reg ( .D(g31864), .SI(g8920), .SE(n8299), .CLK(n8713), .Q(
        g164), .QN(n5561) );
  SDFFX1 DFF_1340_Q_reg ( .D(g34630), .SI(g164), .SE(n8253), .CLK(n8667), .Q(
        g4253), .QN(n5484) );
  SDFFX1 DFF_1341_Q_reg ( .D(g31898), .SI(g4253), .SE(n8317), .CLK(n8731), .Q(
        g5016), .QN(n5369) );
  SDFFX1 DFF_1342_Q_reg ( .D(g25653), .SI(g5016), .SE(n8320), .CLK(n8734), .Q(
        g3119), .QN(n5423) );
  SDFFX1 DFF_1343_Q_reg ( .D(g25632), .SI(g3119), .SE(n8347), .CLK(n8761), .Q(
        g1351), .QN(n5322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g32988), .SI(g1351), .SE(n8347), .CLK(n8761), .Q(
        test_so94), .QN(n8210) );
  SDFFX1 DFF_1345_Q_reg ( .D(g33616), .SI(test_si95), .SE(n8252), .CLK(n8666), 
        .Q(g4519) );
  SDFFX1 DFF_1346_Q_reg ( .D(g29280), .SI(g4519), .SE(n8269), .CLK(n8683), .Q(
        g5115), .QN(n5743) );
  SDFFX1 DFF_1347_Q_reg ( .D(g33609), .SI(g5115), .SE(n8269), .CLK(n8683), .Q(
        g3352), .QN(n5604) );
  SDFFX1 DFF_1348_Q_reg ( .D(g30563), .SI(g3352), .SE(n8340), .CLK(n8754), .Q(
        g6657) );
  SDFFX1 DFF_1349_Q_reg ( .D(g33044), .SI(g6657), .SE(n8337), .CLK(n8751), .Q(
        g4552) );
  SDFFX1 DFF_1350_Q_reg ( .D(g30437), .SI(g4552), .SE(n8337), .CLK(n8751), .Q(
        g3893), .QN(n7904) );
  SDFFX1 DFF_1351_Q_reg ( .D(g30412), .SI(g3893), .SE(n8319), .CLK(n8733), .Q(
        g3211), .QN(n8095) );
  SDFFX1 DFF_1352_Q_reg ( .D(g17604), .SI(g3211), .SE(n8319), .CLK(n8733), .Q(
        g13049) );
  SDFFX1 DFF_1354_Q_reg ( .D(g16603), .SI(g13049), .SE(n8338), .CLK(n8752), 
        .Q(g16624), .QN(n8059) );
  SDFFX1 DFF_1355_Q_reg ( .D(g30491), .SI(g16624), .SE(n8249), .CLK(n8663), 
        .Q(g5595) );
  SDFFX1 DFF_1356_Q_reg ( .D(g30434), .SI(g5595), .SE(n8350), .CLK(n8764), .Q(
        g3614) );
  SDFFX1 DFF_1357_Q_reg ( .D(g34612), .SI(g3614), .SE(n8289), .CLK(n8703), .Q(
        test_so95) );
  SDFFX1 DFF_1358_Q_reg ( .D(g29259), .SI(test_si96), .SE(n8320), .CLK(n8734), 
        .Q(g3125), .QN(n5781) );
  SDFFX1 DFF_1359_Q_reg ( .D(g13865), .SI(g3125), .SE(n8320), .CLK(n8734), .Q(
        g16686) );
  SDFFX1 DFF_1360_Q_reg ( .D(g25681), .SI(g16686), .SE(n8278), .CLK(n8692), 
        .Q(g3821), .QN(n5428) );
  SDFFX1 DFF_1361_Q_reg ( .D(g25687), .SI(g3821), .SE(n8325), .CLK(n8739), .Q(
        g4141), .QN(n5612) );
  SDFFX1 DFF_1362_Q_reg ( .D(g33617), .SI(g4141), .SE(n8337), .CLK(n8751), .Q(
        g4570) );
  SDFFX1 DFF_1363_Q_reg ( .D(g30479), .SI(g4570), .SE(n8254), .CLK(n8668), .Q(
        g5272) );
  SDFFX1 DFF_1364_Q_reg ( .D(g29256), .SI(g5272), .SE(n8281), .CLK(n8695), .Q(
        g2735), .QN(n5600) );
  SDFFX1 DFF_1365_Q_reg ( .D(g28054), .SI(g2735), .SE(n8344), .CLK(n8758), .Q(
        g728), .QN(n7876) );
  SDFFX1 DFF_1366_Q_reg ( .D(g30535), .SI(g728), .SE(n8344), .CLK(n8758), .Q(
        g6295) );
  SDFFX1 DFF_1368_Q_reg ( .D(g30385), .SI(g6295), .SE(n8260), .CLK(n8674), .Q(
        g2661), .QN(n5418) );
  SDFFX1 DFF_1369_Q_reg ( .D(g30361), .SI(g2661), .SE(n8272), .CLK(n8686), .Q(
        g1988), .QN(n5783) );
  SDFFX1 DFF_1370_Q_reg ( .D(g25705), .SI(g1988), .SE(n8268), .CLK(n8682), .Q(
        test_so96), .QN(n8211) );
  SDFFX1 DFF_1371_Q_reg ( .D(g24260), .SI(test_si97), .SE(n8313), .CLK(n8727), 
        .Q(g1548), .QN(n5546) );
  SDFFX1 DFF_1372_Q_reg ( .D(g29257), .SI(g1548), .SE(n8320), .CLK(n8734), .Q(
        g3106), .QN(n5742) );
  SDFFX1 DFF_1373_Q_reg ( .D(g34461), .SI(g3106), .SE(n8327), .CLK(n8741), .Q(
        g4659), .QN(n8152) );
  SDFFX1 DFF_1374_Q_reg ( .D(g34258), .SI(g4659), .SE(n8327), .CLK(n8741), .Q(
        g4358), .QN(n5348) );
  SDFFX1 DFF_1375_Q_reg ( .D(g32993), .SI(g4358), .SE(n8300), .CLK(n8714), .Q(
        g1792), .QN(n5359) );
  SDFFX1 DFF_1376_Q_reg ( .D(g33992), .SI(g1792), .SE(n8291), .CLK(n8705), .Q(
        g2084), .QN(n7783) );
  SDFFX1 DFF_1378_Q_reg ( .D(g30394), .SI(g2084), .SE(n8326), .CLK(n8740), .Q(
        g3187), .QN(n8038) );
  SDFFX1 DFF_1379_Q_reg ( .D(g34449), .SI(g3187), .SE(n8326), .CLK(n8740), .Q(
        g4311), .QN(n5323) );
  SDFFX1 DFF_1380_Q_reg ( .D(g34019), .SI(g4311), .SE(n8350), .CLK(n8764), .Q(
        g2583), .QN(n5800) );
  SDFFX1 DFF_1381_Q_reg ( .D(g18597), .SI(g2583), .SE(n8249), .CLK(n8663), .Q(
        n9240), .QN(DFF_1381_n1) );
  SDFFX1 DFF_1382_Q_reg ( .D(g29231), .SI(n9240), .SE(n8249), .CLK(n8663), .Q(
        g1094) );
  SDFFX1 DFF_1383_Q_reg ( .D(g25682), .SI(g1094), .SE(n8335), .CLK(n8749), .Q(
        test_so97) );
  SDFFX1 DFF_1384_Q_reg ( .D(g21897), .SI(test_si98), .SE(n8303), .CLK(n8717), 
        .Q(g4284), .QN(n7812) );
  SDFFX1 DFF_1386_Q_reg ( .D(g30395), .SI(g4284), .SE(n8328), .CLK(n8742), .Q(
        g3191), .QN(n7880) );
  SDFFX1 DFF_1387_Q_reg ( .D(g21892), .SI(g3191), .SE(n8311), .CLK(n8725), .Q(
        g4239), .QN(n7797) );
  SDFFX1 DFF_1389_Q_reg ( .D(g8789), .SI(g4239), .SE(n8311), .CLK(n8725), .Q(
        g4180), .QN(n5380) );
  SDFFX1 DFF_1390_Q_reg ( .D(g28048), .SI(g4180), .SE(n8264), .CLK(n8678), .Q(
        g691), .QN(n5520) );
  SDFFX1 DFF_1391_Q_reg ( .D(g34723), .SI(g691), .SE(n8277), .CLK(n8691), .Q(
        g534), .QN(n5490) );
  SDFFX1 DFF_1393_Q_reg ( .D(g25598), .SI(g534), .SE(n8312), .CLK(n8726), .Q(
        g385), .QN(n5632) );
  SDFFX1 DFF_1394_Q_reg ( .D(g33987), .SI(g385), .SE(n8291), .CLK(n8705), .Q(
        g2004), .QN(n5818) );
  SDFFX1 DFF_1395_Q_reg ( .D(g30380), .SI(g2004), .SE(n8308), .CLK(n8722), .Q(
        g2527), .QN(n5420) );
  SDFFX1 DFF_1396_Q_reg ( .D(g9555), .SI(g2527), .SE(n8308), .CLK(n8722), .Q(
        g5456), .QN(n7733) );
  SDFFX1 DFF_1397_Q_reg ( .D(g26965), .SI(g5456), .SE(n8346), .CLK(n8760), .Q(
        n6007), .QN(n7857) );
  SDFFX1 DFF_1398_Q_reg ( .D(g25706), .SI(n6007), .SE(n8350), .CLK(n8764), .Q(
        test_so98), .QN(n8238) );
  SDFFX1 DFF_1399_Q_reg ( .D(g30458), .SI(test_si99), .SE(n8266), .CLK(n8680), 
        .Q(g4507), .QN(n5846) );
  SDFFX1 DFF_1400_Q_reg ( .D(g24338), .SI(g4507), .SE(n8269), .CLK(n8683), .Q(
        g5348), .QN(n8127) );
  SDFFX1 DFF_1401_Q_reg ( .D(g30400), .SI(g5348), .SE(n8319), .CLK(n8733), .Q(
        g3223) );
  SDFFX1 DFF_1403_Q_reg ( .D(g34623), .SI(g3223), .SE(n8271), .CLK(n8685), .Q(
        g2970), .QN(n8167) );
  SDFFX1 DFF_1404_Q_reg ( .D(g24343), .SI(g2970), .SE(n8271), .CLK(n8685), .Q(
        g5698), .QN(n7991) );
  SDFFX1 DFF_1406_Q_reg ( .D(g30473), .SI(g5698), .SE(n8302), .CLK(n8716), .Q(
        g5260) );
  SDFFX1 DFF_1407_Q_reg ( .D(g24252), .SI(g5260), .SE(n8314), .CLK(n8728), .Q(
        g1521) );
  SDFFX1 DFF_1408_Q_reg ( .D(g33028), .SI(g1521), .SE(n8315), .CLK(n8729), .Q(
        g3522), .QN(n5383) );
  SDFFX1 DFF_1409_Q_reg ( .D(g29258), .SI(g3522), .SE(n8320), .CLK(n8734), .Q(
        g3115), .QN(n7757) );
  SDFFX1 DFF_1410_Q_reg ( .D(g30407), .SI(g3115), .SE(n8321), .CLK(n8735), .Q(
        g3251) );
  SDFFX1 DFF_1411_Q_reg ( .D(g26958), .SI(g3251), .SE(n8301), .CLK(n8715), .Q(
        g12832) );
  SDFFX1 DFF_1412_Q_reg ( .D(g34457), .SI(g12832), .SE(n8301), .CLK(n8715), 
        .Q(test_so99), .QN(n8218) );
  SDFFX1 DFF_1413_Q_reg ( .D(g33568), .SI(test_si100), .SE(n8284), .CLK(n8698), 
        .Q(g1996), .QN(n5355) );
  SDFFX1 DFF_1414_Q_reg ( .D(g25663), .SI(g1996), .SE(n8252), .CLK(n8666), .Q(
        g8342), .QN(n7712) );
  SDFFX1 DFF_1415_Q_reg ( .D(g26964), .SI(g8342), .SE(n8252), .CLK(n8666), .Q(
        g4515), .QN(n8134) );
  SDFFX1 DFF_1416_Q_reg ( .D(g8786), .SI(g4515), .SE(n8315), .CLK(n8729), .Q(
        g8787) );
  SDFFX1 DFF_1417_Q_reg ( .D(g34735), .SI(g8787), .SE(n8253), .CLK(n8667), .Q(
        g4300), .QN(n5639) );
  SDFFX1 DFF_1418_Q_reg ( .D(g30352), .SI(g4300), .SE(n8352), .CLK(n8766), .Q(
        n9236), .QN(n14521) );
  SDFFX1 DFF_1419_Q_reg ( .D(g33543), .SI(n9236), .SE(n8261), .CLK(n8675), .Q(
        g1379), .QN(n7778) );
  SDFFX1 DFF_1420_Q_reg ( .D(g24271), .SI(g1379), .SE(n8296), .CLK(n8710), .Q(
        g11388), .QN(n5433) );
  SDFFX1 DFF_1422_Q_reg ( .D(g33981), .SI(g11388), .SE(n8287), .CLK(n8701), 
        .Q(g1878) );
  SDFFX1 DFF_1423_Q_reg ( .D(g30500), .SI(g1878), .SE(n8250), .CLK(n8664), .Q(
        g5619) );
  SDFFX1 DFF_1424_Q_reg ( .D(g34649), .SI(g5619), .SE(n8266), .CLK(n8680), .Q(
        g71) );
  SDFFX1 DFF_1425_Q_reg ( .D(g29277), .SI(g71), .SE(n8250), .CLK(n8664), .Q(
        test_so100) );
  SDFFX1 DFF_748_Q_reg ( .D(n8202), .SI(g4704), .SE(n8345), .CLK(n8759), .Q(
        g22), .QN(n7810) );
  SDFFX1 DFF_591_Q_reg ( .D(g25612), .SI(g3897), .SE(n8334), .CLK(n8748), .Q(
        g518), .QN(n5287) );
  SDFFX1 DFF_845_Q_reg ( .D(g28060), .SI(g626), .SE(n8281), .CLK(n8695), .Q(
        g2729), .QN(n7867) );
  HADDX1 Trojan_U1_1_30 ( .A0(counter_30), .B0(carry_30), .C1(carry_31), .SO(
        N31) );
  HADDX1 Trojan_U1_1_4 ( .A0(counter_4), .B0(carry_4), .C1(carry_5), .SO(N5)
         );
  HADDX1 Trojan_U1_1_5 ( .A0(counter_5), .B0(carry_5), .C1(carry_6), .SO(N6)
         );
  HADDX1 Trojan_U1_1_6 ( .A0(counter_6), .B0(carry_6), .C1(carry_7), .SO(N7)
         );
  HADDX1 Trojan_U1_1_7 ( .A0(counter_7), .B0(carry_7), .C1(carry_8), .SO(N8)
         );
  HADDX1 Trojan_U1_1_8 ( .A0(counter_8), .B0(carry_8), .C1(carry_9), .SO(N9)
         );
  HADDX1 Trojan_U1_1_9 ( .A0(counter_9), .B0(carry_9), .C1(carry_10), .SO(N10)
         );
  HADDX1 Trojan_U1_1_10 ( .A0(counter_10), .B0(carry_10), .C1(carry_11), .SO(
        N11) );
  HADDX1 Trojan_U1_1_11 ( .A0(counter_11), .B0(carry_11), .C1(carry_12), .SO(
        N12) );
  HADDX1 Trojan_U1_1_12 ( .A0(counter_12), .B0(carry_12), .C1(carry_13), .SO(
        N13) );
  HADDX1 Trojan_U1_1_13 ( .A0(counter_13), .B0(carry_13), .C1(carry_14), .SO(
        N14) );
  HADDX1 Trojan_U1_1_14 ( .A0(counter_14), .B0(carry_14), .C1(carry_15), .SO(
        N15) );
  HADDX1 Trojan_U1_1_22 ( .A0(counter_22), .B0(carry_22), .C1(carry_23), .SO(
        N23) );
  HADDX1 Trojan_U1_1_23 ( .A0(counter_23), .B0(carry_23), .C1(carry_24), .SO(
        N24) );
  HADDX1 Trojan_U1_1_24 ( .A0(counter_24), .B0(carry_24), .C1(carry_25), .SO(
        N25) );
  HADDX1 Trojan_U1_1_25 ( .A0(counter_25), .B0(carry_25), .C1(carry_26), .SO(
        N26) );
  HADDX1 Trojan_U1_1_1 ( .A0(counter_1), .B0(counter_0), .C1(carry_2), .SO(N2)
         );
  HADDX1 Trojan_U1_1_2 ( .A0(counter_2), .B0(carry_2), .C1(carry_3), .SO(N3)
         );
  HADDX1 Trojan_U1_1_3 ( .A0(counter_3), .B0(carry_3), .C1(carry_4), .SO(N4)
         );
  HADDX1 Trojan_U1_1_15 ( .A0(counter_15), .B0(carry_15), .C1(carry_16), .SO(
        N16) );
  HADDX1 Trojan_U1_1_16 ( .A0(counter_16), .B0(carry_16), .C1(carry_17), .SO(
        N17) );
  HADDX1 Trojan_U1_1_17 ( .A0(counter_17), .B0(carry_17), .C1(carry_18), .SO(
        N18) );
  HADDX1 Trojan_U1_1_18 ( .A0(counter_18), .B0(carry_18), .C1(carry_19), .SO(
        N19) );
  HADDX1 Trojan_U1_1_19 ( .A0(counter_19), .B0(carry_19), .C1(carry_20), .SO(
        N20) );
  HADDX1 Trojan_U1_1_20 ( .A0(counter_20), .B0(carry_20), .C1(carry_21), .SO(
        N21) );
  HADDX1 Trojan_U1_1_21 ( .A0(counter_21), .B0(carry_21), .C1(carry_22), .SO(
        N22) );
  HADDX1 Trojan_U1_1_26 ( .A0(counter_26), .B0(carry_26), .C1(carry_27), .SO(
        N27) );
  HADDX1 Trojan_U1_1_27 ( .A0(counter_27), .B0(carry_27), .C1(carry_28), .SO(
        N28) );
  HADDX1 Trojan_U1_1_28 ( .A0(counter_28), .B0(carry_28), .C1(carry_29), .SO(
        N29) );
  HADDX1 Trojan_U1_1_29 ( .A0(counter_29), .B0(carry_29), .C1(carry_30), .SO(
        N30) );
  INVX0 Trojan_U1 ( .INP(counter_0), .ZN(N1) );
  XOR2X1 Trojan_U2 ( .IN1(carry_31), .IN2(counter_31), .Q(N32) );
  DFFARX1 Trojan_counter_reg_31_ ( .D(N32), .CLK(n37), .RSTB(n8247), .Q(
        counter_31), .QN(n73) );
  DFFARX1 Trojan_counter_reg_1_ ( .D(N2), .CLK(n37), .RSTB(n8246), .Q(
        counter_1) );
  DFFARX1 Trojan_counter_reg_2_ ( .D(N3), .CLK(n37), .RSTB(n87), .Q(counter_2)
         );
  DFFARX1 Trojan_counter_reg_3_ ( .D(N4), .CLK(n37), .RSTB(n8247), .Q(
        counter_3), .QN(n86) );
  DFFARX1 Trojan_counter_reg_15_ ( .D(N16), .CLK(n37), .RSTB(n8246), .Q(
        counter_15), .QN(n85) );
  DFFARX1 Trojan_counter_reg_16_ ( .D(N17), .CLK(n37), .RSTB(n87), .Q(
        counter_16), .QN(n84) );
  DFFARX1 Trojan_counter_reg_17_ ( .D(N18), .CLK(n37), .RSTB(n8247), .Q(
        counter_17), .QN(n83) );
  DFFARX1 Trojan_counter_reg_18_ ( .D(N19), .CLK(n37), .RSTB(n8246), .Q(
        counter_18), .QN(n82) );
  DFFARX1 Trojan_counter_reg_19_ ( .D(N20), .CLK(n37), .RSTB(n87), .Q(
        counter_19), .QN(n81) );
  DFFARX1 Trojan_counter_reg_20_ ( .D(N21), .CLK(n37), .RSTB(n8247), .Q(
        counter_20), .QN(n80) );
  DFFARX1 Trojan_counter_reg_21_ ( .D(N22), .CLK(n37), .RSTB(n8246), .Q(
        counter_21), .QN(n79) );
  DFFARX1 Trojan_counter_reg_26_ ( .D(N27), .CLK(n37), .RSTB(n87), .Q(
        counter_26), .QN(n78) );
  DFFARX1 Trojan_counter_reg_27_ ( .D(N28), .CLK(n37), .RSTB(n8247), .Q(
        counter_27), .QN(n77) );
  DFFARX1 Trojan_counter_reg_28_ ( .D(N29), .CLK(n37), .RSTB(n8246), .Q(
        counter_28), .QN(n76) );
  DFFARX1 Trojan_counter_reg_29_ ( .D(N30), .CLK(n37), .RSTB(n87), .Q(
        counter_29), .QN(n75) );
  DFFARX1 Trojan_counter_reg_30_ ( .D(N31), .CLK(n37), .RSTB(n8247), .Q(
        counter_30), .QN(n74) );
  DFFARX1 Trojan_counter_reg_7_ ( .D(N8), .CLK(n37), .RSTB(n8246), .Q(
        counter_7) );
  DFFARX1 Trojan_counter_reg_11_ ( .D(N12), .CLK(n37), .RSTB(n87), .Q(
        counter_11) );
  DFFARX1 Trojan_counter_reg_25_ ( .D(N26), .CLK(n37), .RSTB(n8247), .Q(
        counter_25) );
  DFFARX1 Trojan_counter_reg_6_ ( .D(N7), .CLK(n37), .RSTB(n8246), .Q(
        counter_6) );
  DFFARX1 Trojan_counter_reg_10_ ( .D(N11), .CLK(n37), .RSTB(n87), .Q(
        counter_10) );
  DFFARX1 Trojan_counter_reg_12_ ( .D(N13), .CLK(n37), .RSTB(n8247), .Q(
        counter_12) );
  DFFARX1 Trojan_counter_reg_24_ ( .D(N25), .CLK(n37), .RSTB(n8246), .Q(
        counter_24) );
  DFFARX1 Trojan_counter_reg_4_ ( .D(N5), .CLK(n37), .RSTB(n87), .Q(counter_4)
         );
  DFFARX1 Trojan_counter_reg_5_ ( .D(N6), .CLK(n37), .RSTB(n8247), .Q(
        counter_5) );
  DFFARX1 Trojan_counter_reg_9_ ( .D(N10), .CLK(n37), .RSTB(n8246), .Q(
        counter_9) );
  DFFARX1 Trojan_counter_reg_14_ ( .D(N15), .CLK(n37), .RSTB(n87), .Q(
        counter_14) );
  DFFARX1 Trojan_counter_reg_23_ ( .D(N24), .CLK(n37), .RSTB(n8247), .Q(
        counter_23) );
  DFFARX1 Trojan_counter_reg_8_ ( .D(N9), .CLK(n37), .RSTB(n8246), .Q(
        counter_8) );
  DFFARX1 Trojan_counter_reg_13_ ( .D(N14), .CLK(n37), .RSTB(n87), .Q(
        counter_13) );
  DFFARX1 Trojan_counter_reg_22_ ( .D(N23), .CLK(n37), .RSTB(n8247), .Q(
        counter_22) );
  DFFARX1 Trojan_counter_reg_0_ ( .D(N1), .CLK(n37), .RSTB(n8246), .Q(
        counter_0) );
  NAND4X0 Trojan_U14 ( .IN1(n3180), .IN2(n3121), .IN3(n2461), .IN4(n58), .QN(
        n87) );
  INVX0 Trojan_U15 ( .INP(n59), .ZN(n58) );
  NOR4X0 Trojan_U16 ( .IN1(n3180), .IN2(n3121), .IN3(n2461), .IN4(n59), .QN(
        n37) );
  NAND3X0 Trojan_U17 ( .IN1(n2601), .IN2(n5111), .IN3(n60), .QN(n59) );
  AND3X1 Trojan_U18 ( .IN1(n2396), .IN2(n42), .IN3(n8194), .Q(n60) );
  NOR4X0 Trojan_U19 ( .IN1(n61), .IN2(n62), .IN3(n63), .IN4(n64), .QN(
        Trigger_out) );
  NAND4X0 Trojan_U20 ( .IN1(n78), .IN2(n77), .IN3(n76), .IN4(n75), .QN(n64) );
  NAND4X0 Trojan_U21 ( .IN1(n74), .IN2(n73), .IN3(counter_6), .IN4(counter_5), 
        .QN(n63) );
  NAND4X0 Trojan_U22 ( .IN1(n80), .IN2(n79), .IN3(n81), .IN4(n65), .QN(n62) );
  NOR4X0 Trojan_U23 ( .IN1(counter_25), .IN2(counter_24), .IN3(counter_23), 
        .IN4(counter_22), .QN(n65) );
  NAND4X0 Trojan_U24 ( .IN1(n66), .IN2(n67), .IN3(n68), .IN4(n69), .QN(n61) );
  NOR4X0 Trojan_U25 ( .IN1(n70), .IN2(counter_12), .IN3(counter_14), .IN4(
        counter_13), .QN(n69) );
  NAND4X0 Trojan_U26 ( .IN1(n85), .IN2(n84), .IN3(n83), .IN4(n82), .QN(n70) );
  NOR4X0 Trojan_U27 ( .IN1(counter_11), .IN2(counter_10), .IN3(counter_9), 
        .IN4(counter_8), .QN(n68) );
  MUX21X1 Trojan_U28 ( .IN1(n71), .IN2(n72), .S(n86), .Q(n67) );
  OA21X1 Trojan_U29 ( .IN1(counter_1), .IN2(counter_0), .IN3(counter_2), .Q(
        n72) );
  NAND2X0 Trojan_U30 ( .IN1(counter_2), .IN2(counter_1), .QN(n71) );
  NOR2X0 Trojan_U31 ( .IN1(counter_7), .IN2(counter_4), .QN(n66) );
  MUX21X1 Trojan_Paylod ( .IN1(g10122_Tj), .IN2(g25715), .S(Trigger_out), .Q(
        g10122) );
  INVX0 U8183 ( .INP(n87), .ZN(n8245) );
  INVX0 U8184 ( .INP(n8245), .ZN(n8246) );
  INVX0 U8186 ( .INP(n8245), .ZN(n8247) );
  NBUFFX2 U8187 ( .INP(n8376), .Z(n8249) );
  NBUFFX2 U8188 ( .INP(n8376), .Z(n8248) );
  NBUFFX2 U8189 ( .INP(n8375), .Z(n8252) );
  NBUFFX2 U8190 ( .INP(n8365), .Z(n8301) );
  NBUFFX2 U8191 ( .INP(n8356), .Z(n8349) );
  NBUFFX2 U8193 ( .INP(n8363), .Z(n8310) );
  NBUFFX2 U8194 ( .INP(n8372), .Z(n8269) );
  NBUFFX2 U8195 ( .INP(n8364), .Z(n8308) );
  NBUFFX2 U8196 ( .INP(n8362), .Z(n8318) );
  NBUFFX2 U8197 ( .INP(n8363), .Z(n8313) );
  NBUFFX2 U8198 ( .INP(n8360), .Z(n8328) );
  NBUFFX2 U8199 ( .INP(n8359), .Z(n8333) );
  NBUFFX2 U8200 ( .INP(n8368), .Z(n8285) );
  NBUFFX2 U8201 ( .INP(n8360), .Z(n8329) );
  NBUFFX2 U8202 ( .INP(n8357), .Z(n8340) );
  NBUFFX2 U8203 ( .INP(n8356), .Z(n8348) );
  NBUFFX2 U8204 ( .INP(n8371), .Z(n8274) );
  NBUFFX2 U8205 ( .INP(n8366), .Z(n8298) );
  NBUFFX2 U8206 ( .INP(n8357), .Z(n8344) );
  NBUFFX2 U8207 ( .INP(n8364), .Z(n8309) );
  NBUFFX2 U8208 ( .INP(n8367), .Z(n8294) );
  NBUFFX2 U8209 ( .INP(n8363), .Z(n8311) );
  NBUFFX2 U8211 ( .INP(n8359), .Z(n8332) );
  NBUFFX2 U8212 ( .INP(n8374), .Z(n8258) );
  NBUFFX2 U8213 ( .INP(n8372), .Z(n8266) );
  NBUFFX2 U8214 ( .INP(n8374), .Z(n8255) );
  NBUFFX2 U8215 ( .INP(n8358), .Z(n8337) );
  NBUFFX2 U8216 ( .INP(n8367), .Z(n8293) );
  NBUFFX2 U8217 ( .INP(n8367), .Z(n8290) );
  NBUFFX2 U8218 ( .INP(n8356), .Z(n8346) );
  NBUFFX2 U8219 ( .INP(n8358), .Z(n8338) );
  NBUFFX2 U8220 ( .INP(n8370), .Z(n8277) );
  NBUFFX2 U8221 ( .INP(n8365), .Z(n8300) );
  NBUFFX2 U8222 ( .INP(n8370), .Z(n8275) );
  NBUFFX2 U8225 ( .INP(n8367), .Z(n8292) );
  NBUFFX2 U8226 ( .INP(n8356), .Z(n8347) );
  NBUFFX2 U8227 ( .INP(n8375), .Z(n8251) );
  NBUFFX2 U8228 ( .INP(n8361), .Z(n8322) );
  NBUFFX2 U8229 ( .INP(n8362), .Z(n8319) );
  NBUFFX2 U8230 ( .INP(n8375), .Z(n8254) );
  NBUFFX2 U8231 ( .INP(n8357), .Z(n8341) );
  NBUFFX2 U8232 ( .INP(n8369), .Z(n8280) );
  NBUFFX2 U8233 ( .INP(n8357), .Z(n8342) );
  NBUFFX2 U8234 ( .INP(n8359), .Z(n8330) );
  NBUFFX2 U8235 ( .INP(n8368), .Z(n8286) );
  NBUFFX2 U8236 ( .INP(n8372), .Z(n8267) );
  NBUFFX2 U8237 ( .INP(n8360), .Z(n8325) );
  NBUFFX2 U8238 ( .INP(n8373), .Z(n8264) );
  NBUFFX2 U8239 ( .INP(n8364), .Z(n8307) );
  NBUFFX2 U8240 ( .INP(n8369), .Z(n8281) );
  NBUFFX2 U8241 ( .INP(n8365), .Z(n8302) );
  NBUFFX2 U8242 ( .INP(n8372), .Z(n8265) );
  NBUFFX2 U8243 ( .INP(n8369), .Z(n8284) );
  NBUFFX2 U8244 ( .INP(n8369), .Z(n8283) );
  NBUFFX2 U8245 ( .INP(n8369), .Z(n8282) );
  NBUFFX2 U8246 ( .INP(n8370), .Z(n8278) );
  NBUFFX2 U8247 ( .INP(n8370), .Z(n8276) );
  NBUFFX2 U8248 ( .INP(n8366), .Z(n8297) );
  NBUFFX2 U8249 ( .INP(n8366), .Z(n8295) );
  NBUFFX2 U8250 ( .INP(n8367), .Z(n8291) );
  NBUFFX2 U8251 ( .INP(n8357), .Z(n8343) );
  NBUFFX2 U8252 ( .INP(n8368), .Z(n8289) );
  NBUFFX2 U8253 ( .INP(n8363), .Z(n8314) );
  NBUFFX2 U8254 ( .INP(n8373), .Z(n8261) );
  NBUFFX2 U8255 ( .INP(n8360), .Z(n8327) );
  NBUFFX2 U8256 ( .INP(n8365), .Z(n8303) );
  NBUFFX2 U8257 ( .INP(n8373), .Z(n8262) );
  NBUFFX2 U8258 ( .INP(n8361), .Z(n8321) );
  NBUFFX2 U8259 ( .INP(n8375), .Z(n8250) );
  NBUFFX2 U8260 ( .INP(n8362), .Z(n8317) );
  NBUFFX2 U8261 ( .INP(n8374), .Z(n8256) );
  NBUFFX2 U8262 ( .INP(n8374), .Z(n8259) );
  NBUFFX2 U8263 ( .INP(n8356), .Z(n8345) );
  NBUFFX2 U8264 ( .INP(n8361), .Z(n8323) );
  NBUFFX2 U8265 ( .INP(n8373), .Z(n8260) );
  NBUFFX2 U8266 ( .INP(n8359), .Z(n8331) );
  NBUFFX2 U8267 ( .INP(n8371), .Z(n8271) );
  NBUFFX2 U8268 ( .INP(n8370), .Z(n8279) );
  NBUFFX2 U8269 ( .INP(n8358), .Z(n8339) );
  NBUFFX2 U8270 ( .INP(n8363), .Z(n8312) );
  NBUFFX2 U8271 ( .INP(n8360), .Z(n8326) );
  NBUFFX2 U8272 ( .INP(n8366), .Z(n8296) );
  NBUFFX2 U8273 ( .INP(n8362), .Z(n8315) );
  NBUFFX2 U8274 ( .INP(n8362), .Z(n8316) );
  NBUFFX2 U8275 ( .INP(n8365), .Z(n8304) );
  NBUFFX2 U8276 ( .INP(n8361), .Z(n8324) );
  NBUFFX2 U8277 ( .INP(n8366), .Z(n8299) );
  NBUFFX2 U8278 ( .INP(n8358), .Z(n8336) );
  NBUFFX2 U8279 ( .INP(n8364), .Z(n8306) );
  NBUFFX2 U8280 ( .INP(n8371), .Z(n8273) );
  NBUFFX2 U8282 ( .INP(n8368), .Z(n8288) );
  NBUFFX2 U8283 ( .INP(n8371), .Z(n8272) );
  NBUFFX2 U8284 ( .INP(n8371), .Z(n8270) );
  NBUFFX2 U8285 ( .INP(n8358), .Z(n8335) );
  NBUFFX2 U8286 ( .INP(n8375), .Z(n8253) );
  NBUFFX2 U8287 ( .INP(n8374), .Z(n8257) );
  NBUFFX2 U8288 ( .INP(n8361), .Z(n8320) );
  NBUFFX2 U8289 ( .INP(n8364), .Z(n8305) );
  NBUFFX2 U8290 ( .INP(n8372), .Z(n8268) );
  NBUFFX2 U8291 ( .INP(n8359), .Z(n8334) );
  NBUFFX2 U8292 ( .INP(n8368), .Z(n8287) );
  NBUFFX2 U8293 ( .INP(n8373), .Z(n8263) );
  NBUFFX2 U8294 ( .INP(n8790), .Z(n8663) );
  NBUFFX2 U8295 ( .INP(n8790), .Z(n8662) );
  NBUFFX2 U8296 ( .INP(n8789), .Z(n8666) );
  NBUFFX2 U8297 ( .INP(n8779), .Z(n8715) );
  NBUFFX2 U8298 ( .INP(n8770), .Z(n8763) );
  NBUFFX2 U8299 ( .INP(n8777), .Z(n8724) );
  NBUFFX2 U8300 ( .INP(n8786), .Z(n8683) );
  NBUFFX2 U8301 ( .INP(n8778), .Z(n8722) );
  NBUFFX2 U8302 ( .INP(n8776), .Z(n8732) );
  NBUFFX2 U8303 ( .INP(n8777), .Z(n8727) );
  NBUFFX2 U8304 ( .INP(n8774), .Z(n8742) );
  NBUFFX2 U8305 ( .INP(n8773), .Z(n8747) );
  NBUFFX2 U8306 ( .INP(n8782), .Z(n8699) );
  NBUFFX2 U8308 ( .INP(n8774), .Z(n8743) );
  NBUFFX2 U8309 ( .INP(n8771), .Z(n8754) );
  NBUFFX2 U8310 ( .INP(n8770), .Z(n8762) );
  NBUFFX2 U8311 ( .INP(n8785), .Z(n8688) );
  NBUFFX2 U8312 ( .INP(n8780), .Z(n8712) );
  NBUFFX2 U8313 ( .INP(n8771), .Z(n8758) );
  NBUFFX2 U8314 ( .INP(n8778), .Z(n8723) );
  NBUFFX2 U8315 ( .INP(n8781), .Z(n8708) );
  NBUFFX2 U8316 ( .INP(n8777), .Z(n8725) );
  NBUFFX2 U8317 ( .INP(n8773), .Z(n8746) );
  NBUFFX2 U8318 ( .INP(n8788), .Z(n8672) );
  NBUFFX2 U8319 ( .INP(n8786), .Z(n8680) );
  NBUFFX2 U8320 ( .INP(n8788), .Z(n8669) );
  NBUFFX2 U8321 ( .INP(n8772), .Z(n8751) );
  NBUFFX2 U8322 ( .INP(n8781), .Z(n8707) );
  NBUFFX2 U8323 ( .INP(n8781), .Z(n8704) );
  NBUFFX2 U8324 ( .INP(n8770), .Z(n8760) );
  NBUFFX2 U8325 ( .INP(n8772), .Z(n8752) );
  NBUFFX2 U8326 ( .INP(n8784), .Z(n8691) );
  NBUFFX2 U8327 ( .INP(n8779), .Z(n8714) );
  NBUFFX2 U8328 ( .INP(n8784), .Z(n8689) );
  NBUFFX2 U8329 ( .INP(n8781), .Z(n8706) );
  NBUFFX2 U8330 ( .INP(n8770), .Z(n8761) );
  NBUFFX2 U8331 ( .INP(n8789), .Z(n8665) );
  NBUFFX2 U8332 ( .INP(n8775), .Z(n8736) );
  NBUFFX2 U8333 ( .INP(n8776), .Z(n8733) );
  NBUFFX2 U8334 ( .INP(n8789), .Z(n8668) );
  NBUFFX2 U8335 ( .INP(n8771), .Z(n8755) );
  NBUFFX2 U8336 ( .INP(n8783), .Z(n8694) );
  NBUFFX2 U8337 ( .INP(n8771), .Z(n8756) );
  NBUFFX2 U8338 ( .INP(n8773), .Z(n8744) );
  NBUFFX2 U8339 ( .INP(n8782), .Z(n8700) );
  NBUFFX2 U8340 ( .INP(n8786), .Z(n8681) );
  NBUFFX2 U8341 ( .INP(n8774), .Z(n8739) );
  NBUFFX2 U8342 ( .INP(n8787), .Z(n8678) );
  NBUFFX2 U8343 ( .INP(n8778), .Z(n8721) );
  NBUFFX2 U8344 ( .INP(n8783), .Z(n8695) );
  NBUFFX2 U8345 ( .INP(n8779), .Z(n8716) );
  NBUFFX2 U8346 ( .INP(n8786), .Z(n8679) );
  NBUFFX2 U8347 ( .INP(n8783), .Z(n8698) );
  NBUFFX2 U8348 ( .INP(n8783), .Z(n8697) );
  NBUFFX2 U8349 ( .INP(n8783), .Z(n8696) );
  NBUFFX2 U8350 ( .INP(n8784), .Z(n8692) );
  NBUFFX2 U8351 ( .INP(n8784), .Z(n8690) );
  NBUFFX2 U8352 ( .INP(n8780), .Z(n8711) );
  NBUFFX2 U8353 ( .INP(n8780), .Z(n8709) );
  NBUFFX2 U8354 ( .INP(n8781), .Z(n8705) );
  NBUFFX2 U8355 ( .INP(n8771), .Z(n8757) );
  NBUFFX2 U8356 ( .INP(n8782), .Z(n8703) );
  NBUFFX2 U8357 ( .INP(n8777), .Z(n8728) );
  NBUFFX2 U8358 ( .INP(n8787), .Z(n8675) );
  NBUFFX2 U8359 ( .INP(n8774), .Z(n8741) );
  NBUFFX2 U8360 ( .INP(n8779), .Z(n8717) );
  NBUFFX2 U8361 ( .INP(n8787), .Z(n8676) );
  NBUFFX2 U8362 ( .INP(n8775), .Z(n8735) );
  NBUFFX2 U8363 ( .INP(n8789), .Z(n8664) );
  NBUFFX2 U8364 ( .INP(n8776), .Z(n8731) );
  NBUFFX2 U8365 ( .INP(n8788), .Z(n8670) );
  NBUFFX2 U8366 ( .INP(n8788), .Z(n8673) );
  NBUFFX2 U8367 ( .INP(n8770), .Z(n8759) );
  NBUFFX2 U8368 ( .INP(n8775), .Z(n8737) );
  NBUFFX2 U8369 ( .INP(n8787), .Z(n8674) );
  NBUFFX2 U8370 ( .INP(n8773), .Z(n8745) );
  NBUFFX2 U8371 ( .INP(n8785), .Z(n8685) );
  NBUFFX2 U8372 ( .INP(n8784), .Z(n8693) );
  NBUFFX2 U8373 ( .INP(n8772), .Z(n8753) );
  NBUFFX2 U8374 ( .INP(n8777), .Z(n8726) );
  NBUFFX2 U8375 ( .INP(n8774), .Z(n8740) );
  NBUFFX2 U8376 ( .INP(n8780), .Z(n8710) );
  NBUFFX2 U8377 ( .INP(n8776), .Z(n8729) );
  NBUFFX2 U8378 ( .INP(n8776), .Z(n8730) );
  NBUFFX2 U8379 ( .INP(n8779), .Z(n8718) );
  NBUFFX2 U8380 ( .INP(n8775), .Z(n8738) );
  NBUFFX2 U8381 ( .INP(n8780), .Z(n8713) );
  NBUFFX2 U8382 ( .INP(n8772), .Z(n8750) );
  NBUFFX2 U8383 ( .INP(n8778), .Z(n8720) );
  NBUFFX2 U8384 ( .INP(n8785), .Z(n8687) );
  NBUFFX2 U8385 ( .INP(n8782), .Z(n8702) );
  NBUFFX2 U8386 ( .INP(n8785), .Z(n8686) );
  NBUFFX2 U8387 ( .INP(n8785), .Z(n8684) );
  NBUFFX2 U8388 ( .INP(n8772), .Z(n8749) );
  NBUFFX2 U8389 ( .INP(n8789), .Z(n8667) );
  NBUFFX2 U8390 ( .INP(n8788), .Z(n8671) );
  NBUFFX2 U8391 ( .INP(n8775), .Z(n8734) );
  NBUFFX2 U8392 ( .INP(n8778), .Z(n8719) );
  NBUFFX2 U8393 ( .INP(n8786), .Z(n8682) );
  NBUFFX2 U8394 ( .INP(n8773), .Z(n8748) );
  NBUFFX2 U8395 ( .INP(n8782), .Z(n8701) );
  NBUFFX2 U8396 ( .INP(n8787), .Z(n8677) );
  INVX0 U8397 ( .INP(n8396), .ZN(n8544) );
  INVX0 U8398 ( .INP(n8408), .ZN(n8568) );
  INVX0 U8399 ( .INP(n8411), .ZN(n8575) );
  INVX0 U8400 ( .INP(n8409), .ZN(n8570) );
  INVX0 U8401 ( .INP(n8410), .ZN(n8573) );
  INVX0 U8402 ( .INP(n8409), .ZN(n8571) );
  INVX0 U8403 ( .INP(n8411), .ZN(n8574) );
  INVX0 U8404 ( .INP(n8408), .ZN(n8569) );
  INVX0 U8405 ( .INP(n8410), .ZN(n8572) );
  INVX0 U8406 ( .INP(n8412), .ZN(n8576) );
  INVX0 U8407 ( .INP(n8396), .ZN(n8545) );
  INVX0 U8408 ( .INP(n8397), .ZN(n8546) );
  INVX0 U8409 ( .INP(n8392), .ZN(n8537) );
  INVX0 U8410 ( .INP(n8412), .ZN(n8577) );
  INVX0 U8411 ( .INP(n8415), .ZN(n8582) );
  INVX0 U8412 ( .INP(n8413), .ZN(n8579) );
  INVX0 U8413 ( .INP(n8413), .ZN(n8578) );
  INVX0 U8414 ( .INP(n8416), .ZN(n8584) );
  INVX0 U8415 ( .INP(n8414), .ZN(n8581) );
  INVX0 U8416 ( .INP(n8414), .ZN(n8580) );
  INVX0 U8417 ( .INP(n8415), .ZN(n8583) );
  INVX0 U8418 ( .INP(n8404), .ZN(n8560) );
  INVX0 U8419 ( .INP(n8400), .ZN(n8553) );
  INVX0 U8420 ( .INP(n8405), .ZN(n8562) );
  INVX0 U8421 ( .INP(n8398), .ZN(n8549) );
  INVX0 U8422 ( .INP(n8404), .ZN(n8561) );
  INVX0 U8423 ( .INP(n8402), .ZN(n8556) );
  INVX0 U8424 ( .INP(n8399), .ZN(n8550) );
  INVX0 U8425 ( .INP(n8403), .ZN(n8559) );
  INVX0 U8426 ( .INP(n8398), .ZN(n8548) );
  INVX0 U8427 ( .INP(n8399), .ZN(n8551) );
  INVX0 U8428 ( .INP(n8405), .ZN(n8563) );
  INVX0 U8429 ( .INP(n8400), .ZN(n8552) );
  INVX0 U8430 ( .INP(n8402), .ZN(n8557) );
  INVX0 U8431 ( .INP(n8401), .ZN(n8555) );
  INVX0 U8432 ( .INP(n8401), .ZN(n8554) );
  INVX0 U8433 ( .INP(n8403), .ZN(n8558) );
  INVX0 U8434 ( .INP(n8454), .ZN(n8659) );
  INVX0 U8435 ( .INP(n8388), .ZN(n8529) );
  INVX0 U8436 ( .INP(n8388), .ZN(n8530) );
  INVX0 U8437 ( .INP(n8390), .ZN(n8533) );
  INVX0 U8438 ( .INP(n8391), .ZN(n8536) );
  INVX0 U8439 ( .INP(n8389), .ZN(n8532) );
  INVX0 U8440 ( .INP(n8389), .ZN(n8531) );
  INVX0 U8441 ( .INP(n8390), .ZN(n8534) );
  INVX0 U8442 ( .INP(n8391), .ZN(n8535) );
  INVX0 U8443 ( .INP(n8416), .ZN(n8585) );
  INVX0 U8444 ( .INP(n8455), .ZN(n8661) );
  INVX0 U8445 ( .INP(n8455), .ZN(n8660) );
  INVX0 U8446 ( .INP(n8397), .ZN(n8547) );
  INVX0 U8447 ( .INP(n8407), .ZN(n8567) );
  INVX0 U8448 ( .INP(n8407), .ZN(n8566) );
  INVX0 U8449 ( .INP(n8406), .ZN(n8565) );
  INVX0 U8450 ( .INP(n8395), .ZN(n8543) );
  INVX0 U8451 ( .INP(n8393), .ZN(n8539) );
  INVX0 U8452 ( .INP(n8394), .ZN(n8540) );
  INVX0 U8453 ( .INP(n8395), .ZN(n8542) );
  INVX0 U8454 ( .INP(n8394), .ZN(n8541) );
  INVX0 U8455 ( .INP(n8393), .ZN(n8538) );
  INVX0 U8456 ( .INP(n8406), .ZN(n8564) );
  INVX0 U8457 ( .INP(n8419), .ZN(n8590) );
  INVX0 U8458 ( .INP(n8427), .ZN(n8607) );
  INVX0 U8459 ( .INP(n8418), .ZN(n8588) );
  INVX0 U8460 ( .INP(n8429), .ZN(n8610) );
  INVX0 U8461 ( .INP(n8448), .ZN(n8647) );
  INVX0 U8462 ( .INP(n8431), .ZN(n8614) );
  INVX0 U8463 ( .INP(n8424), .ZN(n8600) );
  INVX0 U8464 ( .INP(n8452), .ZN(n8656) );
  INVX0 U8465 ( .INP(n8438), .ZN(n8628) );
  INVX0 U8466 ( .INP(n8423), .ZN(n8599) );
  INVX0 U8467 ( .INP(n8432), .ZN(n8616) );
  INVX0 U8468 ( .INP(n8426), .ZN(n8605) );
  INVX0 U8469 ( .INP(n8452), .ZN(n8655) );
  INVX0 U8470 ( .INP(n8449), .ZN(n8649) );
  INVX0 U8471 ( .INP(n8444), .ZN(n8639) );
  INVX0 U8472 ( .INP(n8451), .ZN(n8653) );
  INVX0 U8473 ( .INP(n8420), .ZN(n8593) );
  INVX0 U8474 ( .INP(n8439), .ZN(n8630) );
  INVX0 U8475 ( .INP(n8448), .ZN(n8648) );
  INVX0 U8476 ( .INP(n8432), .ZN(n8617) );
  INVX0 U8477 ( .INP(n8422), .ZN(n8597) );
  INVX0 U8478 ( .INP(n8431), .ZN(n8615) );
  INVX0 U8479 ( .INP(n8435), .ZN(n8621) );
  INVX0 U8480 ( .INP(n8422), .ZN(n8596) );
  INVX0 U8481 ( .INP(n8424), .ZN(n8601) );
  INVX0 U8482 ( .INP(n8417), .ZN(n8586) );
  INVX0 U8483 ( .INP(n8430), .ZN(n8613) );
  INVX0 U8484 ( .INP(n8441), .ZN(n8634) );
  INVX0 U8485 ( .INP(n8430), .ZN(n8612) );
  INVX0 U8486 ( .INP(n8440), .ZN(n8631) );
  INVX0 U8487 ( .INP(n8446), .ZN(n8644) );
  INVX0 U8488 ( .INP(n8450), .ZN(n8651) );
  INVX0 U8489 ( .INP(n8421), .ZN(n8595) );
  INVX0 U8490 ( .INP(n8442), .ZN(n8635) );
  INVX0 U8491 ( .INP(n8427), .ZN(n8606) );
  INVX0 U8492 ( .INP(n8423), .ZN(n8598) );
  INVX0 U8493 ( .INP(n8440), .ZN(n8632) );
  INVX0 U8494 ( .INP(n8425), .ZN(n8602) );
  INVX0 U8495 ( .INP(n8441), .ZN(n8633) );
  INVX0 U8496 ( .INP(n8451), .ZN(n8654) );
  INVX0 U8497 ( .INP(n8443), .ZN(n8638) );
  INVX0 U8498 ( .INP(n8429), .ZN(n8611) );
  INVX0 U8499 ( .INP(n8446), .ZN(n8643) );
  INVX0 U8500 ( .INP(n8447), .ZN(n8646) );
  INVX0 U8501 ( .INP(n8421), .ZN(n8594) );
  INVX0 U8502 ( .INP(n8437), .ZN(n8625) );
  INVX0 U8503 ( .INP(n8450), .ZN(n8652) );
  INVX0 U8504 ( .INP(n8425), .ZN(n8603) );
  INVX0 U8505 ( .INP(n8420), .ZN(n8592) );
  INVX0 U8506 ( .INP(n8439), .ZN(n8629) );
  INVX0 U8507 ( .INP(n8428), .ZN(n8608) );
  INVX0 U8508 ( .INP(n8435), .ZN(n8622) );
  INVX0 U8509 ( .INP(n8438), .ZN(n8627) );
  INVX0 U8510 ( .INP(n8436), .ZN(n8624) );
  INVX0 U8511 ( .INP(n8447), .ZN(n8645) );
  INVX0 U8512 ( .INP(n8445), .ZN(n8641) );
  INVX0 U8513 ( .INP(n8453), .ZN(n8658) );
  INVX0 U8514 ( .INP(n8444), .ZN(n8640) );
  INVX0 U8515 ( .INP(n8426), .ZN(n8604) );
  INVX0 U8516 ( .INP(n8428), .ZN(n8609) );
  INVX0 U8517 ( .INP(n8417), .ZN(n8587) );
  INVX0 U8518 ( .INP(n8433), .ZN(n8618) );
  INVX0 U8519 ( .INP(n8449), .ZN(n8650) );
  INVX0 U8520 ( .INP(n8442), .ZN(n8636) );
  INVX0 U8521 ( .INP(n8445), .ZN(n8642) );
  INVX0 U8522 ( .INP(n8434), .ZN(n8619) );
  INVX0 U8523 ( .INP(n8443), .ZN(n8637) );
  INVX0 U8524 ( .INP(n8419), .ZN(n8591) );
  INVX0 U8525 ( .INP(n8418), .ZN(n8589) );
  INVX0 U8526 ( .INP(n8436), .ZN(n8623) );
  INVX0 U8527 ( .INP(n8434), .ZN(n8620) );
  INVX0 U8528 ( .INP(n8437), .ZN(n8626) );
  INVX0 U8529 ( .INP(n8453), .ZN(n8657) );
  NBUFFX2 U8530 ( .INP(n8355), .Z(n8353) );
  NBUFFX2 U8531 ( .INP(n8355), .Z(n8350) );
  NBUFFX2 U8532 ( .INP(n8355), .Z(n8351) );
  NBUFFX2 U8533 ( .INP(n8355), .Z(n8352) );
  NBUFFX2 U8534 ( .INP(n8769), .Z(n8767) );
  NBUFFX2 U8535 ( .INP(n8769), .Z(n8764) );
  NBUFFX2 U8536 ( .INP(n8769), .Z(n8765) );
  NBUFFX2 U8537 ( .INP(n8769), .Z(n8766) );
  NBUFFX2 U8538 ( .INP(n8355), .Z(n8354) );
  NBUFFX2 U8539 ( .INP(n8470), .Z(n8388) );
  NBUFFX2 U8540 ( .INP(n8470), .Z(n8389) );
  NBUFFX2 U8541 ( .INP(n8470), .Z(n8390) );
  NBUFFX2 U8542 ( .INP(n8470), .Z(n8391) );
  NBUFFX2 U8543 ( .INP(n8468), .Z(n8397) );
  NBUFFX2 U8544 ( .INP(n8465), .Z(n8412) );
  NBUFFX2 U8545 ( .INP(n8467), .Z(n8406) );
  NBUFFX2 U8546 ( .INP(n8467), .Z(n8404) );
  NBUFFX2 U8547 ( .INP(n8468), .Z(n8400) );
  NBUFFX2 U8548 ( .INP(n8467), .Z(n8405) );
  NBUFFX2 U8549 ( .INP(n8465), .Z(n8415) );
  NBUFFX2 U8550 ( .INP(n8466), .Z(n8407) );
  NBUFFX2 U8551 ( .INP(n8467), .Z(n8402) );
  NBUFFX2 U8552 ( .INP(n8465), .Z(n8413) );
  NBUFFX2 U8553 ( .INP(n8465), .Z(n8416) );
  NBUFFX2 U8554 ( .INP(n8467), .Z(n8403) );
  NBUFFX2 U8555 ( .INP(n8465), .Z(n8414) );
  NBUFFX2 U8556 ( .INP(n8456), .Z(n8452) );
  NBUFFX2 U8557 ( .INP(n8466), .Z(n8411) );
  NBUFFX2 U8558 ( .INP(n8457), .Z(n8448) );
  NBUFFX2 U8559 ( .INP(n8466), .Z(n8409) );
  NBUFFX2 U8560 ( .INP(n8461), .Z(n8432) );
  NBUFFX2 U8561 ( .INP(n8461), .Z(n8431) );
  NBUFFX2 U8562 ( .INP(n8463), .Z(n8422) );
  NBUFFX2 U8563 ( .INP(n8463), .Z(n8424) );
  NBUFFX2 U8564 ( .INP(n8462), .Z(n8430) );
  NBUFFX2 U8565 ( .INP(n8456), .Z(n8455) );
  NBUFFX2 U8566 ( .INP(n8469), .Z(n8396) );
  NBUFFX2 U8567 ( .INP(n8469), .Z(n8395) );
  NBUFFX2 U8568 ( .INP(n8462), .Z(n8427) );
  NBUFFX2 U8569 ( .INP(n8463), .Z(n8423) );
  NBUFFX2 U8570 ( .INP(n8459), .Z(n8440) );
  NBUFFX2 U8571 ( .INP(n8459), .Z(n8441) );
  NBUFFX2 U8572 ( .INP(n8466), .Z(n8410) );
  NBUFFX2 U8573 ( .INP(n8468), .Z(n8398) );
  NBUFFX2 U8574 ( .INP(n8457), .Z(n8451) );
  NBUFFX2 U8575 ( .INP(n8468), .Z(n8399) );
  NBUFFX2 U8576 ( .INP(n8462), .Z(n8429) );
  NBUFFX2 U8577 ( .INP(n8458), .Z(n8446) );
  NBUFFX2 U8578 ( .INP(n8469), .Z(n8394) );
  NBUFFX2 U8579 ( .INP(n8463), .Z(n8421) );
  NBUFFX2 U8580 ( .INP(n8457), .Z(n8450) );
  NBUFFX2 U8581 ( .INP(n8463), .Z(n8425) );
  NBUFFX2 U8582 ( .INP(n8464), .Z(n8420) );
  NBUFFX2 U8583 ( .INP(n8459), .Z(n8439) );
  NBUFFX2 U8584 ( .INP(n8460), .Z(n8435) );
  NBUFFX2 U8585 ( .INP(n8459), .Z(n8438) );
  NBUFFX2 U8586 ( .INP(n8469), .Z(n8392) );
  NBUFFX2 U8587 ( .INP(n8457), .Z(n8447) );
  NBUFFX2 U8588 ( .INP(n8458), .Z(n8444) );
  NBUFFX2 U8589 ( .INP(n8462), .Z(n8426) );
  NBUFFX2 U8590 ( .INP(n8462), .Z(n8428) );
  NBUFFX2 U8591 ( .INP(n8464), .Z(n8417) );
  NBUFFX2 U8592 ( .INP(n8469), .Z(n8393) );
  NBUFFX2 U8593 ( .INP(n8460), .Z(n8433) );
  NBUFFX2 U8594 ( .INP(n8457), .Z(n8449) );
  NBUFFX2 U8595 ( .INP(n8456), .Z(n8454) );
  NBUFFX2 U8596 ( .INP(n8458), .Z(n8442) );
  NBUFFX2 U8597 ( .INP(n8458), .Z(n8445) );
  NBUFFX2 U8598 ( .INP(n8458), .Z(n8443) );
  NBUFFX2 U8599 ( .INP(n8464), .Z(n8419) );
  NBUFFX2 U8600 ( .INP(n8464), .Z(n8418) );
  NBUFFX2 U8601 ( .INP(n8460), .Z(n8436) );
  NBUFFX2 U8602 ( .INP(n8460), .Z(n8434) );
  NBUFFX2 U8603 ( .INP(n8459), .Z(n8437) );
  NBUFFX2 U8604 ( .INP(n8456), .Z(n8453) );
  NBUFFX2 U8605 ( .INP(n8468), .Z(n8401) );
  NBUFFX2 U8606 ( .INP(n8466), .Z(n8408) );
  NBUFFX2 U8607 ( .INP(n8769), .Z(n8768) );
  NBUFFX2 U8608 ( .INP(n8384), .Z(n8355) );
  NBUFFX2 U8609 ( .INP(n8383), .Z(n8356) );
  NBUFFX2 U8610 ( .INP(n8383), .Z(n8357) );
  NBUFFX2 U8611 ( .INP(n8383), .Z(n8358) );
  NBUFFX2 U8612 ( .INP(n8382), .Z(n8359) );
  NBUFFX2 U8613 ( .INP(n8382), .Z(n8360) );
  NBUFFX2 U8614 ( .INP(n8382), .Z(n8361) );
  NBUFFX2 U8615 ( .INP(n8381), .Z(n8362) );
  NBUFFX2 U8616 ( .INP(n8381), .Z(n8363) );
  NBUFFX2 U8617 ( .INP(n8381), .Z(n8364) );
  NBUFFX2 U8618 ( .INP(n8380), .Z(n8365) );
  NBUFFX2 U8619 ( .INP(n8380), .Z(n8366) );
  NBUFFX2 U8620 ( .INP(n8380), .Z(n8367) );
  NBUFFX2 U8621 ( .INP(n8379), .Z(n8368) );
  NBUFFX2 U8622 ( .INP(n8379), .Z(n8369) );
  NBUFFX2 U8623 ( .INP(n8379), .Z(n8370) );
  NBUFFX2 U8624 ( .INP(n8378), .Z(n8371) );
  NBUFFX2 U8625 ( .INP(n8378), .Z(n8372) );
  NBUFFX2 U8626 ( .INP(n8378), .Z(n8373) );
  NBUFFX2 U8627 ( .INP(n8377), .Z(n8374) );
  NBUFFX2 U8628 ( .INP(n8377), .Z(n8375) );
  NBUFFX2 U8629 ( .INP(n8377), .Z(n8376) );
  NBUFFX2 U8630 ( .INP(n8387), .Z(n8377) );
  NBUFFX2 U8631 ( .INP(n8387), .Z(n8378) );
  NBUFFX2 U8632 ( .INP(n8386), .Z(n8379) );
  NBUFFX2 U8633 ( .INP(n8386), .Z(n8380) );
  NBUFFX2 U8634 ( .INP(n8386), .Z(n8381) );
  NBUFFX2 U8635 ( .INP(n8385), .Z(n8382) );
  NBUFFX2 U8636 ( .INP(n8385), .Z(n8383) );
  NBUFFX2 U8637 ( .INP(n8385), .Z(n8384) );
  NBUFFX2 U8638 ( .INP(test_se), .Z(n8385) );
  NBUFFX2 U8639 ( .INP(test_se), .Z(n8386) );
  NBUFFX2 U8640 ( .INP(test_se), .Z(n8387) );
  NBUFFX2 U8641 ( .INP(n8475), .Z(n8456) );
  NBUFFX2 U8642 ( .INP(n8475), .Z(n8457) );
  NBUFFX2 U8643 ( .INP(n8475), .Z(n8458) );
  NBUFFX2 U8644 ( .INP(n8474), .Z(n8459) );
  NBUFFX2 U8645 ( .INP(n8474), .Z(n8460) );
  NBUFFX2 U8646 ( .INP(n8474), .Z(n8461) );
  NBUFFX2 U8647 ( .INP(n8473), .Z(n8462) );
  NBUFFX2 U8648 ( .INP(n8473), .Z(n8463) );
  NBUFFX2 U8649 ( .INP(n8473), .Z(n8464) );
  NBUFFX2 U8650 ( .INP(n8472), .Z(n8465) );
  NBUFFX2 U8651 ( .INP(n8472), .Z(n8466) );
  NBUFFX2 U8652 ( .INP(n8472), .Z(n8467) );
  NBUFFX2 U8653 ( .INP(n8471), .Z(n8468) );
  NBUFFX2 U8654 ( .INP(n8471), .Z(n8469) );
  NBUFFX2 U8655 ( .INP(n8471), .Z(n8470) );
  NBUFFX2 U8656 ( .INP(g35), .Z(n8471) );
  NBUFFX2 U8657 ( .INP(g35), .Z(n8472) );
  NBUFFX2 U8658 ( .INP(g35), .Z(n8473) );
  NBUFFX2 U8659 ( .INP(g35), .Z(n8474) );
  NBUFFX2 U8660 ( .INP(g35), .Z(n8475) );
  INVX0 U8661 ( .INP(n8579), .ZN(n8476) );
  INVX0 U8662 ( .INP(n8580), .ZN(n8477) );
  INVX0 U8663 ( .INP(n8581), .ZN(n8478) );
  INVX0 U8664 ( .INP(n8581), .ZN(n8479) );
  INVX0 U8665 ( .INP(n8578), .ZN(n8480) );
  INVX0 U8666 ( .INP(n8582), .ZN(n8481) );
  INVX0 U8667 ( .INP(n8580), .ZN(n8482) );
  INVX0 U8668 ( .INP(n8583), .ZN(n8483) );
  INVX0 U8669 ( .INP(n8578), .ZN(n8484) );
  INVX0 U8670 ( .INP(n8584), .ZN(n8485) );
  INVX0 U8671 ( .INP(n8582), .ZN(n8486) );
  INVX0 U8672 ( .INP(n8581), .ZN(n8487) );
  INVX0 U8673 ( .INP(n8583), .ZN(n8488) );
  INVX0 U8674 ( .INP(n8580), .ZN(n8489) );
  INVX0 U8675 ( .INP(n8585), .ZN(n8490) );
  INVX0 U8676 ( .INP(n8585), .ZN(n8491) );
  INVX0 U8677 ( .INP(n8585), .ZN(n8492) );
  INVX0 U8678 ( .INP(n8582), .ZN(n8493) );
  INVX0 U8679 ( .INP(n8585), .ZN(n8494) );
  INVX0 U8680 ( .INP(n8582), .ZN(n8495) );
  INVX0 U8681 ( .INP(n8580), .ZN(n8496) );
  INVX0 U8682 ( .INP(n8584), .ZN(n8497) );
  INVX0 U8683 ( .INP(n8584), .ZN(n8498) );
  INVX0 U8684 ( .INP(n8584), .ZN(n8499) );
  INVX0 U8685 ( .INP(n8581), .ZN(n8500) );
  INVX0 U8686 ( .INP(n8584), .ZN(n8501) );
  INVX0 U8687 ( .INP(n8584), .ZN(n8502) );
  INVX0 U8688 ( .INP(n8583), .ZN(n8503) );
  INVX0 U8689 ( .INP(n8583), .ZN(n8504) );
  INVX0 U8690 ( .INP(n8583), .ZN(n8505) );
  INVX0 U8691 ( .INP(n8583), .ZN(n8506) );
  INVX0 U8692 ( .INP(n8578), .ZN(n8507) );
  INVX0 U8693 ( .INP(n8582), .ZN(n8508) );
  INVX0 U8694 ( .INP(n8582), .ZN(n8509) );
  INVX0 U8695 ( .INP(n8579), .ZN(n8510) );
  INVX0 U8696 ( .INP(n8578), .ZN(n8511) );
  INVX0 U8697 ( .INP(n8581), .ZN(n8512) );
  INVX0 U8698 ( .INP(n8580), .ZN(n8513) );
  INVX0 U8699 ( .INP(n8580), .ZN(n8514) );
  INVX0 U8700 ( .INP(n8578), .ZN(n8515) );
  INVX0 U8701 ( .INP(n8579), .ZN(n8516) );
  INVX0 U8702 ( .INP(n8579), .ZN(n8517) );
  INVX0 U8703 ( .INP(n8577), .ZN(n8518) );
  INVX0 U8704 ( .INP(n8579), .ZN(n8519) );
  INVX0 U8705 ( .INP(n8579), .ZN(n8520) );
  INVX0 U8706 ( .INP(n8578), .ZN(n8521) );
  INVX0 U8707 ( .INP(n8577), .ZN(n8522) );
  INVX0 U8708 ( .INP(n8577), .ZN(n8523) );
  INVX0 U8709 ( .INP(n8577), .ZN(n8524) );
  INVX0 U8710 ( .INP(n8577), .ZN(n8525) );
  INVX0 U8711 ( .INP(n8577), .ZN(n8526) );
  INVX0 U8712 ( .INP(n8581), .ZN(n8527) );
  INVX0 U8713 ( .INP(n8576), .ZN(n8528) );
  NBUFFX2 U8714 ( .INP(n8798), .Z(n8769) );
  NBUFFX2 U8715 ( .INP(n8797), .Z(n8770) );
  NBUFFX2 U8716 ( .INP(n8797), .Z(n8771) );
  NBUFFX2 U8717 ( .INP(n8797), .Z(n8772) );
  NBUFFX2 U8718 ( .INP(n8796), .Z(n8773) );
  NBUFFX2 U8719 ( .INP(n8796), .Z(n8774) );
  NBUFFX2 U8720 ( .INP(n8796), .Z(n8775) );
  NBUFFX2 U8721 ( .INP(n8795), .Z(n8776) );
  NBUFFX2 U8722 ( .INP(n8795), .Z(n8777) );
  NBUFFX2 U8723 ( .INP(n8795), .Z(n8778) );
  NBUFFX2 U8724 ( .INP(n8794), .Z(n8779) );
  NBUFFX2 U8725 ( .INP(n8794), .Z(n8780) );
  NBUFFX2 U8726 ( .INP(n8794), .Z(n8781) );
  NBUFFX2 U8727 ( .INP(n8793), .Z(n8782) );
  NBUFFX2 U8728 ( .INP(n8793), .Z(n8783) );
  NBUFFX2 U8729 ( .INP(n8793), .Z(n8784) );
  NBUFFX2 U8730 ( .INP(n8792), .Z(n8785) );
  NBUFFX2 U8731 ( .INP(n8792), .Z(n8786) );
  NBUFFX2 U8732 ( .INP(n8792), .Z(n8787) );
  NBUFFX2 U8733 ( .INP(n8791), .Z(n8788) );
  NBUFFX2 U8734 ( .INP(n8791), .Z(n8789) );
  NBUFFX2 U8735 ( .INP(n8791), .Z(n8790) );
  NBUFFX2 U8736 ( .INP(n8801), .Z(n8791) );
  NBUFFX2 U8737 ( .INP(n8801), .Z(n8792) );
  NBUFFX2 U8738 ( .INP(n8800), .Z(n8793) );
  NBUFFX2 U8739 ( .INP(n8800), .Z(n8794) );
  NBUFFX2 U8740 ( .INP(n8800), .Z(n8795) );
  NBUFFX2 U8741 ( .INP(n8799), .Z(n8796) );
  NBUFFX2 U8742 ( .INP(n8799), .Z(n8797) );
  NBUFFX2 U8743 ( .INP(n8799), .Z(n8798) );
  NBUFFX2 U8744 ( .INP(CK), .Z(n8799) );
  NBUFFX2 U8745 ( .INP(CK), .Z(n8800) );
  NBUFFX2 U8746 ( .INP(CK), .Z(n8801) );
  INVX0 U8747 ( .INP(n8802), .ZN(n965) );
  NOR3X0 U8748 ( .IN1(n8803), .IN2(n8804), .IN3(n8805), .QN(n8193) );
  INVX0 U8749 ( .INP(n8806), .ZN(n8192) );
  INVX0 U8750 ( .INP(n8807), .ZN(n628) );
  NAND4X0 U8751 ( .IN1(n8808), .IN2(n8809), .IN3(n8810), .IN4(n8811), .QN(
        n5961) );
  NAND2X0 U8752 ( .IN1(n8812), .IN2(g5348), .QN(n8811) );
  NAND2X0 U8753 ( .IN1(n8127), .IN2(n8813), .QN(n8810) );
  NAND2X0 U8754 ( .IN1(g31860), .IN2(g5352), .QN(n8809) );
  NAND2X0 U8755 ( .IN1(n8126), .IN2(n8814), .QN(n8808) );
  NAND4X0 U8756 ( .IN1(n8815), .IN2(n8816), .IN3(n8817), .IN4(n8818), .QN(
        n5960) );
  NAND2X0 U8757 ( .IN1(n8819), .IN2(g6732), .QN(n8818) );
  NAND2X0 U8758 ( .IN1(n8125), .IN2(n8820), .QN(n8817) );
  NAND2X0 U8759 ( .IN1(n8821), .IN2(g6736), .QN(n8816) );
  NAND2X0 U8760 ( .IN1(n8124), .IN2(n8822), .QN(n8815) );
  INVX0 U8761 ( .INP(n8823), .ZN(n4940) );
  NAND2X0 U8762 ( .IN1(n8824), .IN2(g1677), .QN(n4459) );
  NAND2X0 U8763 ( .IN1(n8825), .IN2(g1811), .QN(n4448) );
  NAND2X0 U8764 ( .IN1(test_so53), .IN2(n8826), .QN(n4437) );
  OR2X1 U8765 ( .IN1(n8827), .IN2(n7915), .Q(n4426) );
  NAND2X0 U8766 ( .IN1(n8828), .IN2(g2236), .QN(n4415) );
  NAND2X0 U8767 ( .IN1(n8829), .IN2(g2370), .QN(n4403) );
  NAND2X0 U8768 ( .IN1(n8830), .IN2(g2504), .QN(n4392) );
  NAND2X0 U8769 ( .IN1(n8831), .IN2(g2638), .QN(n4380) );
  NAND4X0 U8770 ( .IN1(n8832), .IN2(n8833), .IN3(n8834), .IN4(n8835), .QN(
        n4305) );
  NOR2X0 U8771 ( .IN1(n8836), .IN2(n8837), .QN(n8835) );
  NOR2X0 U8772 ( .IN1(n5656), .IN2(g4826), .QN(n8837) );
  NOR2X0 U8773 ( .IN1(n5440), .IN2(g4821), .QN(n8836) );
  NAND2X0 U8774 ( .IN1(g4646), .IN2(g29220), .QN(n8834) );
  NAND4X0 U8775 ( .IN1(n5440), .IN2(n8838), .IN3(n8839), .IN4(n8128), .QN(
        n8833) );
  NOR2X0 U8776 ( .IN1(g4688), .IN2(g4646), .QN(n8839) );
  NAND2X0 U8777 ( .IN1(n8840), .IN2(n8841), .QN(n8838) );
  NAND3X0 U8778 ( .IN1(n8842), .IN2(n8843), .IN3(n8844), .QN(n8840) );
  NAND2X0 U8779 ( .IN1(n8845), .IN2(g4776), .QN(n8844) );
  NAND2X0 U8780 ( .IN1(n5368), .IN2(n8846), .QN(n8845) );
  XOR2X1 U8781 ( .IN1(g34657), .IN2(n8847), .Q(n8846) );
  NAND4X0 U8782 ( .IN1(n8848), .IN2(n8849), .IN3(n8850), .IN4(n8851), .QN(
        n8847) );
  NAND2X0 U8783 ( .IN1(n8852), .IN2(g4732), .QN(n8851) );
  NAND2X0 U8784 ( .IN1(n8853), .IN2(g4717), .QN(n8850) );
  NAND2X0 U8785 ( .IN1(n8854), .IN2(g4727), .QN(n8849) );
  NAND2X0 U8786 ( .IN1(n8855), .IN2(g4722), .QN(n8848) );
  NAND2X0 U8787 ( .IN1(n8856), .IN2(g4793), .QN(n8843) );
  NAND2X0 U8788 ( .IN1(n5368), .IN2(n8857), .QN(n8842) );
  NAND2X0 U8789 ( .IN1(n8215), .IN2(n8858), .QN(n8857) );
  OR4X1 U8790 ( .IN1(g4776), .IN2(n8859), .IN3(n8852), .IN4(n8853), .Q(n8858)
         );
  AND2X1 U8791 ( .IN1(n8854), .IN2(n5867), .Q(n8859) );
  NAND2X0 U8792 ( .IN1(g4831), .IN2(g4681), .QN(n8832) );
  NAND4X0 U8793 ( .IN1(n8860), .IN2(n8861), .IN3(n8862), .IN4(n8863), .QN(
        n4283) );
  NOR2X0 U8794 ( .IN1(n8864), .IN2(n8865), .QN(n8863) );
  NOR2X0 U8795 ( .IN1(n5318), .IN2(g3333), .QN(n8865) );
  NOR2X0 U8796 ( .IN1(n5283), .IN2(g4035), .QN(n8864) );
  NAND2X0 U8797 ( .IN1(g4871), .IN2(g3684), .QN(n8862) );
  NAND4X0 U8798 ( .IN1(n5283), .IN2(n8866), .IN3(n8867), .IN4(n5713), .QN(
        n8861) );
  NOR2X0 U8799 ( .IN1(g4864), .IN2(g4871), .QN(n8867) );
  NAND2X0 U8800 ( .IN1(n8868), .IN2(n8869), .QN(n8866) );
  NAND3X0 U8801 ( .IN1(n8870), .IN2(n8871), .IN3(n8872), .QN(n8868) );
  NAND2X0 U8802 ( .IN1(n8873), .IN2(g4966), .QN(n8872) );
  NAND2X0 U8803 ( .IN1(n5367), .IN2(n8874), .QN(n8873) );
  XOR2X1 U8804 ( .IN1(g34649), .IN2(n8875), .Q(n8874) );
  NAND4X0 U8805 ( .IN1(n8876), .IN2(n8877), .IN3(n8878), .IN4(n8879), .QN(
        n8875) );
  NAND2X0 U8806 ( .IN1(n8880), .IN2(g4912), .QN(n8879) );
  NAND2X0 U8807 ( .IN1(n8881), .IN2(g4917), .QN(n8878) );
  NAND2X0 U8808 ( .IN1(n8882), .IN2(g4922), .QN(n8877) );
  NAND2X0 U8809 ( .IN1(n8883), .IN2(g4907), .QN(n8876) );
  NAND2X0 U8810 ( .IN1(n8884), .IN2(g4983), .QN(n8871) );
  NAND2X0 U8811 ( .IN1(n5367), .IN2(n8885), .QN(n8870) );
  NAND2X0 U8812 ( .IN1(n8214), .IN2(n8886), .QN(n8885) );
  OR4X1 U8813 ( .IN1(g4966), .IN2(n8887), .IN3(n8882), .IN4(n8883), .Q(n8886)
         );
  AND2X1 U8814 ( .IN1(n8881), .IN2(n5879), .Q(n8887) );
  NAND2X0 U8815 ( .IN1(g4836), .IN2(g5011), .QN(n8860) );
  AND3X1 U8816 ( .IN1(n5652), .IN2(n5366), .IN3(n8150), .Q(n4034) );
  AND3X1 U8817 ( .IN1(n5645), .IN2(n5576), .IN3(n8146), .Q(n4002) );
  NOR3X0 U8818 ( .IN1(g3863), .IN2(test_so33), .IN3(g3857), .QN(n3969) );
  NOR4X0 U8819 ( .IN1(n7841), .IN2(n1430), .IN3(n8805), .IN4(n8803), .QN(n3933) );
  INVX0 U8820 ( .INP(n8888), .ZN(n8803) );
  INVX0 U8821 ( .INP(n8889), .ZN(n8805) );
  AND3X1 U8822 ( .IN1(n5650), .IN2(n5570), .IN3(n8140), .Q(n3926) );
  AND3X1 U8823 ( .IN1(n5647), .IN2(n5575), .IN3(n8145), .Q(n3893) );
  AND3X1 U8824 ( .IN1(n5649), .IN2(n5573), .IN3(n8143), .Q(n3860) );
  AND3X1 U8825 ( .IN1(n5651), .IN2(n5574), .IN3(n8144), .Q(n3826) );
  AND3X1 U8826 ( .IN1(n5646), .IN2(n5571), .IN3(n8141), .Q(n3792) );
  NAND4X0 U8827 ( .IN1(n5358), .IN2(n5520), .IN3(n8890), .IN4(n8891), .QN(
        n3675) );
  NAND2X0 U8828 ( .IN1(n7865), .IN2(n8892), .QN(n8891) );
  NAND2X0 U8829 ( .IN1(n8893), .IN2(n5629), .QN(n8892) );
  XOR2X1 U8830 ( .IN1(g174), .IN2(test_so72), .Q(n8893) );
  NAND2X0 U8831 ( .IN1(n8894), .IN2(g392), .QN(n8890) );
  NAND2X0 U8832 ( .IN1(n8895), .IN2(n7864), .QN(n8894) );
  XNOR2X1 U8833 ( .IN1(n8002), .IN2(test_so72), .Q(n8895) );
  OR2X1 U8834 ( .IN1(n8896), .IN2(n5349), .Q(n3635) );
  INVX0 U8835 ( .INP(n8897), .ZN(n3506) );
  NOR2X0 U8836 ( .IN1(n8898), .IN2(n8899), .QN(n3174) );
  XOR2X1 U8837 ( .IN1(g482), .IN2(g72), .Q(n8899) );
  XOR2X1 U8838 ( .IN1(g490), .IN2(g73), .Q(n8898) );
  NOR2X0 U8839 ( .IN1(n1430), .IN2(n6010), .QN(n3084) );
  NAND3X0 U8840 ( .IN1(n8503), .IN2(g4104), .IN3(n8900), .QN(n3065) );
  NAND2X0 U8841 ( .IN1(n8901), .IN2(g4108), .QN(n8900) );
  XOR2X1 U8842 ( .IN1(n5323), .IN2(n2607), .Q(n2608) );
  NAND2X0 U8843 ( .IN1(n8902), .IN2(g34979), .QN(n2461) );
  NOR2X0 U8844 ( .IN1(n8903), .IN2(n8904), .QN(n2396) );
  INVX0 U8845 ( .INP(n8905), .ZN(n233) );
  NAND2X0 U8846 ( .IN1(n8906), .IN2(n8907), .QN(g34980) );
  NAND2X0 U8847 ( .IN1(test_so14), .IN2(n8536), .QN(n8907) );
  NAND2X0 U8848 ( .IN1(n8908), .IN2(n8513), .QN(n8906) );
  NAND2X0 U8849 ( .IN1(n5842), .IN2(n8909), .QN(n8908) );
  OR4X1 U8850 ( .IN1(n8806), .IN2(g53), .IN3(g54), .IN4(g56), .Q(n8909) );
  NAND2X0 U8851 ( .IN1(n8806), .IN2(g22), .QN(g34972) );
  XOR3X1 U8852 ( .IN1(g34979), .IN2(n8903), .IN3(n8910), .Q(n8806) );
  XNOR3X1 U8853 ( .IN1(n8911), .IN2(g34974), .IN3(n8912), .Q(n8910) );
  XOR3X1 U8854 ( .IN1(n8913), .IN2(n171), .IN3(g34978), .Q(n8912) );
  NAND2X0 U8855 ( .IN1(n8914), .IN2(g55), .QN(n8913) );
  NAND2X0 U8856 ( .IN1(g54), .IN2(n8915), .QN(n8914) );
  XNOR3X1 U8857 ( .IN1(g34970), .IN2(g34977), .IN3(g34976), .Q(n8911) );
  OR2X1 U8858 ( .IN1(g34979), .IN2(n7810), .Q(g34927) );
  NAND4X0 U8859 ( .IN1(n8916), .IN2(n8917), .IN3(n8918), .IN4(n8919), .QN(
        g34979) );
  NOR4X0 U8860 ( .IN1(n8920), .IN2(n8921), .IN3(n8922), .IN4(n8923), .QN(n8919) );
  NOR2X0 U8861 ( .IN1(n5415), .IN2(n8924), .QN(n8923) );
  NOR2X0 U8862 ( .IN1(n5635), .IN2(n8925), .QN(n8922) );
  NOR2X0 U8863 ( .IN1(n5308), .IN2(n8926), .QN(n8921) );
  NOR2X0 U8864 ( .IN1(n8927), .IN2(DFF_420_n1), .QN(n8920) );
  NOR2X0 U8865 ( .IN1(n8928), .IN2(n8929), .QN(n8918) );
  NOR2X0 U8866 ( .IN1(n8930), .IN2(n8240), .QN(n8929) );
  NAND2X0 U8867 ( .IN1(n8202), .IN2(n8931), .QN(n8917) );
  NAND4X0 U8868 ( .IN1(n8932), .IN2(n8933), .IN3(n8934), .IN4(n8935), .QN(
        n8931) );
  NOR4X0 U8869 ( .IN1(n8936), .IN2(n8937), .IN3(n8938), .IN4(n8939), .QN(n8935) );
  AND2X1 U8870 ( .IN1(n8940), .IN2(g29221), .Q(n8939) );
  NOR2X0 U8871 ( .IN1(n5293), .IN2(n8941), .QN(n8938) );
  NOR2X0 U8872 ( .IN1(n5470), .IN2(n8942), .QN(n8937) );
  NAND3X0 U8873 ( .IN1(n8943), .IN2(n8944), .IN3(n8945), .QN(n8936) );
  NAND2X0 U8874 ( .IN1(g127), .IN2(n8946), .QN(n8945) );
  NAND2X0 U8875 ( .IN1(test_so14), .IN2(n8902), .QN(n8944) );
  INVX0 U8876 ( .INP(n8904), .ZN(n8902) );
  NAND2X0 U8877 ( .IN1(g92), .IN2(n8947), .QN(n8943) );
  NOR3X0 U8878 ( .IN1(n8948), .IN2(n8949), .IN3(n8950), .QN(n8934) );
  NOR2X0 U8879 ( .IN1(n5473), .IN2(n8951), .QN(n8950) );
  NOR2X0 U8880 ( .IN1(n5335), .IN2(n8952), .QN(n8949) );
  NOR2X0 U8881 ( .IN1(n5750), .IN2(n8953), .QN(n8948) );
  NAND2X0 U8882 ( .IN1(n8954), .IN2(g2886), .QN(n8933) );
  NOR2X0 U8883 ( .IN1(n8955), .IN2(n8956), .QN(n8932) );
  NOR2X0 U8884 ( .IN1(n8167), .IN2(n8957), .QN(n8956) );
  NOR2X0 U8885 ( .IN1(n5981), .IN2(n8958), .QN(n8955) );
  NAND2X0 U8886 ( .IN1(n8959), .IN2(g2138), .QN(n8916) );
  OR2X1 U8887 ( .IN1(g34978), .IN2(n7810), .Q(g34925) );
  NAND4X0 U8888 ( .IN1(n8960), .IN2(n8961), .IN3(n8962), .IN4(n8963), .QN(
        g34978) );
  NOR4X0 U8889 ( .IN1(n8964), .IN2(n8965), .IN3(n8966), .IN4(n8967), .QN(n8963) );
  NOR2X0 U8890 ( .IN1(n8924), .IN2(g952), .QN(n8967) );
  NOR2X0 U8891 ( .IN1(n8925), .IN2(g1296), .QN(n8966) );
  NOR2X0 U8892 ( .IN1(n5347), .IN2(n8926), .QN(n8965) );
  NOR2X0 U8893 ( .IN1(n8927), .IN2(DFF_1012_n1), .QN(n8964) );
  NOR2X0 U8894 ( .IN1(n8928), .IN2(n8968), .QN(n8962) );
  NOR2X0 U8895 ( .IN1(n5484), .IN2(n8930), .QN(n8968) );
  NAND2X0 U8896 ( .IN1(n8202), .IN2(n8969), .QN(n8961) );
  NAND4X0 U8897 ( .IN1(n8970), .IN2(n8971), .IN3(n8972), .IN4(n8973), .QN(
        n8969) );
  NOR4X0 U8898 ( .IN1(n8974), .IN2(n8975), .IN3(n8976), .IN4(n8977), .QN(n8973) );
  NOR2X0 U8899 ( .IN1(n8942), .IN2(n5471), .QN(n8977) );
  NOR2X0 U8900 ( .IN1(n8978), .IN2(g550), .QN(n8976) );
  NOR2X0 U8901 ( .IN1(n5337), .IN2(n8952), .QN(n8975) );
  NAND3X0 U8902 ( .IN1(n8979), .IN2(n8980), .IN3(n8981), .QN(n8974) );
  NAND2X0 U8903 ( .IN1(n8982), .IN2(g790), .QN(n8981) );
  NAND2X0 U8904 ( .IN1(n8947), .IN2(g29214), .QN(n8980) );
  NAND2X0 U8905 ( .IN1(n8946), .IN2(g2873), .QN(n8979) );
  NOR3X0 U8906 ( .IN1(n8983), .IN2(n8984), .IN3(n8985), .QN(n8972) );
  NOR2X0 U8907 ( .IN1(n7819), .IN2(n8953), .QN(n8985) );
  NOR2X0 U8908 ( .IN1(n5475), .IN2(n8951), .QN(n8984) );
  NOR2X0 U8909 ( .IN1(n5494), .IN2(n8958), .QN(n8983) );
  NAND2X0 U8910 ( .IN1(test_so22), .IN2(n8986), .QN(n8971) );
  NAND2X0 U8911 ( .IN1(n8954), .IN2(g2878), .QN(n8970) );
  NAND2X0 U8912 ( .IN1(n8959), .IN2(g2130), .QN(n8960) );
  INVX0 U8913 ( .INP(n8987), .ZN(n8959) );
  OR2X1 U8914 ( .IN1(g34977), .IN2(n7810), .Q(g34923) );
  NAND4X0 U8915 ( .IN1(n8988), .IN2(n8989), .IN3(n8990), .IN4(n8991), .QN(
        g34977) );
  NOR4X0 U8916 ( .IN1(n8992), .IN2(n8993), .IN3(n8994), .IN4(n8995), .QN(n8991) );
  NOR2X0 U8917 ( .IN1(n5286), .IN2(n8924), .QN(n8995) );
  NOR2X0 U8918 ( .IN1(n2549), .IN2(n8925), .QN(n8994) );
  NOR2X0 U8919 ( .IN1(n8996), .IN2(g4927), .QN(n8993) );
  NOR2X0 U8920 ( .IN1(n8997), .IN2(g4737), .QN(n8992) );
  NOR2X0 U8921 ( .IN1(n8928), .IN2(n8998), .QN(n8990) );
  NOR2X0 U8922 ( .IN1(n5639), .IN2(n8930), .QN(n8998) );
  NAND2X0 U8923 ( .IN1(n8202), .IN2(n8999), .QN(n8989) );
  NAND4X0 U8924 ( .IN1(n9000), .IN2(n9001), .IN3(n9002), .IN4(n9003), .QN(
        n8999) );
  NOR4X0 U8925 ( .IN1(n9004), .IN2(n9005), .IN3(n9006), .IN4(n9007), .QN(n9003) );
  NOR2X0 U8926 ( .IN1(n5490), .IN2(n8978), .QN(n9007) );
  NOR2X0 U8927 ( .IN1(n5291), .IN2(n8941), .QN(n9006) );
  NOR2X0 U8928 ( .IN1(n5331), .IN2(n8942), .QN(n9005) );
  NAND3X0 U8929 ( .IN1(n9008), .IN2(n9009), .IN3(n9010), .QN(n9004) );
  NAND2X0 U8930 ( .IN1(n8946), .IN2(g2868), .QN(n9010) );
  NAND2X0 U8931 ( .IN1(g37), .IN2(n8947), .QN(n9008) );
  NOR3X0 U8932 ( .IN1(n9011), .IN2(n9012), .IN3(n9013), .QN(n9002) );
  NOR2X0 U8933 ( .IN1(n5474), .IN2(n8951), .QN(n9013) );
  NOR2X0 U8934 ( .IN1(n5336), .IN2(n8952), .QN(n9012) );
  NOR2X0 U8935 ( .IN1(n7820), .IN2(n8953), .QN(n9011) );
  NAND2X0 U8936 ( .IN1(n8954), .IN2(g2882), .QN(n9001) );
  NOR2X0 U8937 ( .IN1(n9014), .IN2(n9015), .QN(n9000) );
  NOR2X0 U8938 ( .IN1(n8170), .IN2(n8957), .QN(n9015) );
  NOR2X0 U8939 ( .IN1(n5493), .IN2(n8958), .QN(n9014) );
  NAND2X0 U8940 ( .IN1(n9245), .IN2(n9016), .QN(n8988) );
  INVX0 U8941 ( .INP(n8927), .ZN(n9016) );
  OR2X1 U8942 ( .IN1(g34976), .IN2(n7810), .Q(g34921) );
  NAND4X0 U8943 ( .IN1(n9017), .IN2(n9018), .IN3(n9019), .IN4(n9020), .QN(
        g34976) );
  NOR4X0 U8944 ( .IN1(n9021), .IN2(n9022), .IN3(n9023), .IN4(n9024), .QN(n9020) );
  NOR2X0 U8945 ( .IN1(n5297), .IN2(n8996), .QN(n9024) );
  NOR2X0 U8946 ( .IN1(n5345), .IN2(n8997), .QN(n9023) );
  NOR2X0 U8947 ( .IN1(n5497), .IN2(n8926), .QN(n9022) );
  NOR2X0 U8948 ( .IN1(n8927), .IN2(DFF_150_n1), .QN(n9021) );
  NOR3X0 U8949 ( .IN1(n9025), .IN2(n8928), .IN3(n9026), .QN(n9019) );
  NOR2X0 U8950 ( .IN1(n5289), .IN2(n9027), .QN(n9026) );
  AND2X1 U8951 ( .IN1(g1135), .IN2(n9028), .Q(n9025) );
  NAND2X0 U8952 ( .IN1(n8202), .IN2(n9029), .QN(n9018) );
  NAND4X0 U8953 ( .IN1(n9030), .IN2(n9031), .IN3(n9032), .IN4(n9033), .QN(
        n9029) );
  NOR4X0 U8954 ( .IN1(n9034), .IN2(n9035), .IN3(n9036), .IN4(n9037), .QN(n9033) );
  NOR2X0 U8955 ( .IN1(n5332), .IN2(n8942), .QN(n9037) );
  NOR2X0 U8956 ( .IN1(n8978), .IN2(n8232), .QN(n9036) );
  NOR2X0 U8957 ( .IN1(n5294), .IN2(n8952), .QN(n9035) );
  NAND3X0 U8958 ( .IN1(n9038), .IN2(n9009), .IN3(n9039), .QN(n9034) );
  NAND2X0 U8959 ( .IN1(n8982), .IN2(g807), .QN(n9039) );
  NAND2X0 U8960 ( .IN1(n8946), .IN2(g2988), .QN(n9038) );
  NOR3X0 U8961 ( .IN1(n9040), .IN2(n9041), .IN3(n9042), .QN(n9032) );
  NOR2X0 U8962 ( .IN1(n8172), .IN2(n8953), .QN(n9042) );
  NOR2X0 U8963 ( .IN1(n5339), .IN2(n8951), .QN(n9041) );
  AND2X1 U8964 ( .IN1(n9043), .IN2(test_so95), .Q(n9040) );
  NAND2X0 U8965 ( .IN1(n8986), .IN2(g2936), .QN(n9031) );
  NAND2X0 U8966 ( .IN1(n8954), .IN2(g2898), .QN(n9030) );
  OR2X1 U8967 ( .IN1(n8987), .IN2(n5498), .Q(n9017) );
  OR2X1 U8968 ( .IN1(n171), .IN2(n7810), .Q(g34919) );
  NAND4X0 U8969 ( .IN1(n9044), .IN2(n9045), .IN3(n9046), .IN4(n9047), .QN(n171) );
  NOR4X0 U8970 ( .IN1(n9048), .IN2(n9049), .IN3(n9050), .IN4(n9051), .QN(n9047) );
  NOR2X0 U8971 ( .IN1(n9052), .IN2(n9053), .QN(n9051) );
  NOR4X0 U8972 ( .IN1(n9054), .IN2(n9055), .IN3(n9056), .IN4(n9057), .QN(n9052) );
  NOR2X0 U8973 ( .IN1(n5552), .IN2(n8952), .QN(n9057) );
  NOR2X0 U8976 ( .IN1(n5672), .IN2(n8951), .QN(n9056) );
  NAND3X0 U8977 ( .IN1(n9058), .IN2(n9059), .IN3(n9060), .QN(n9055) );
  NAND2X0 U8978 ( .IN1(n8982), .IN2(g554), .QN(n9060) );
  NAND2X0 U8979 ( .IN1(n8954), .IN2(g2864), .QN(n9059) );
  NAND2X0 U8980 ( .IN1(n5634), .IN2(n8946), .QN(n9058) );
  NAND4X0 U8981 ( .IN1(n9061), .IN2(n9062), .IN3(n9063), .IN4(n9064), .QN(
        n9054) );
  NOR2X0 U8982 ( .IN1(n9065), .IN2(n9066), .QN(n9064) );
  NOR2X0 U8983 ( .IN1(n8169), .IN2(n8957), .QN(n9066) );
  NOR2X0 U8984 ( .IN1(n8164), .IN2(n8958), .QN(n9065) );
  NAND2X0 U8985 ( .IN1(n9067), .IN2(g2927), .QN(n9063) );
  NAND2X0 U8986 ( .IN1(n9068), .IN2(g767), .QN(n9062) );
  NAND2X0 U8987 ( .IN1(n8940), .IN2(g546), .QN(n9061) );
  NOR2X0 U8988 ( .IN1(n5344), .IN2(n8997), .QN(n9050) );
  NOR2X0 U8989 ( .IN1(n5495), .IN2(n8926), .QN(n9049) );
  NOR2X0 U8990 ( .IN1(n14515), .IN2(n8927), .QN(n9048) );
  NOR3X0 U8991 ( .IN1(n9069), .IN2(n9070), .IN3(n8928), .QN(n9046) );
  NOR2X0 U8992 ( .IN1(n5295), .IN2(n8996), .QN(n9070) );
  NOR2X0 U8993 ( .IN1(n5343), .IN2(n9027), .QN(n9069) );
  NAND2X0 U8994 ( .IN1(n9028), .IN2(g1105), .QN(n9045) );
  OR2X1 U8995 ( .IN1(n8987), .IN2(n5643), .Q(n9044) );
  OR2X1 U8996 ( .IN1(g34974), .IN2(n7810), .Q(g34917) );
  NAND4X0 U8997 ( .IN1(n9071), .IN2(n9072), .IN3(n9073), .IN4(n9074), .QN(
        g34974) );
  NOR4X0 U8998 ( .IN1(n9075), .IN2(n9076), .IN3(n9077), .IN4(n9078), .QN(n9074) );
  NOR2X0 U8999 ( .IN1(n5346), .IN2(n8996), .QN(n9078) );
  NOR2X0 U9000 ( .IN1(n5296), .IN2(n8997), .QN(n9077) );
  NOR2X0 U9001 ( .IN1(n8926), .IN2(n8227), .QN(n9076) );
  NOR2X0 U9002 ( .IN1(n8927), .IN2(DFF_477_n1), .QN(n9075) );
  NOR2X0 U9003 ( .IN1(n9079), .IN2(n9080), .QN(n9073) );
  NOR2X0 U9004 ( .IN1(n5499), .IN2(n8987), .QN(n9080) );
  NOR2X0 U9005 ( .IN1(n9081), .IN2(n9053), .QN(n9079) );
  NOR4X0 U9006 ( .IN1(n9082), .IN2(n9083), .IN3(n9084), .IN4(n9085), .QN(n9081) );
  NOR2X0 U9007 ( .IN1(n5288), .IN2(n8951), .QN(n9085) );
  NOR2X0 U9008 ( .IN1(n5472), .IN2(n8952), .QN(n9084) );
  NAND3X0 U9009 ( .IN1(n9086), .IN2(n9087), .IN3(n9088), .QN(n9083) );
  NAND2X0 U9010 ( .IN1(n9068), .IN2(g772), .QN(n9088) );
  NAND2X0 U9011 ( .IN1(n8946), .IN2(g2999), .QN(n9086) );
  NAND4X0 U9012 ( .IN1(n9089), .IN2(n9090), .IN3(n9091), .IN4(n9092), .QN(
        n9082) );
  NAND2X0 U9013 ( .IN1(n9067), .IN2(g2917), .QN(n9092) );
  NAND2X0 U9014 ( .IN1(n9043), .IN2(g2852), .QN(n9091) );
  NAND2X0 U9015 ( .IN1(n8986), .IN2(g2912), .QN(n9090) );
  NAND2X0 U9016 ( .IN1(n8954), .IN2(g2856), .QN(n9089) );
  NAND2X0 U9017 ( .IN1(n9093), .IN2(g1472), .QN(n9072) );
  NAND2X0 U9018 ( .IN1(n9028), .IN2(g1129), .QN(n9071) );
  NAND2X0 U9019 ( .IN1(n8903), .IN2(g22), .QN(g34915) );
  INVX0 U9020 ( .INP(g34971), .ZN(n8903) );
  NAND4X0 U9021 ( .IN1(n9094), .IN2(n9095), .IN3(n9096), .IN4(n9097), .QN(
        g34971) );
  NOR4X0 U9022 ( .IN1(n8928), .IN2(n9098), .IN3(n9099), .IN4(n9100), .QN(n9097) );
  NOR2X0 U9023 ( .IN1(n5307), .IN2(n8987), .QN(n9100) );
  NOR2X0 U9024 ( .IN1(n9101), .IN2(n9053), .QN(n9099) );
  NOR4X0 U9025 ( .IN1(n9102), .IN2(n9103), .IN3(n9104), .IN4(n9105), .QN(n9101) );
  NOR2X0 U9026 ( .IN1(n5983), .IN2(n8958), .QN(n9105) );
  NOR2X0 U9027 ( .IN1(n5550), .IN2(n8951), .QN(n9104) );
  NAND3X0 U9028 ( .IN1(n9106), .IN2(n9107), .IN3(n9108), .QN(n9103) );
  OR2X1 U9029 ( .IN1(n8952), .IN2(n7686), .Q(n9108) );
  OR2X1 U9030 ( .IN1(n8978), .IN2(n8186), .Q(n9107) );
  NAND2X0 U9031 ( .IN1(test_so60), .IN2(n9068), .QN(n9106) );
  NAND4X0 U9032 ( .IN1(n9109), .IN2(n9110), .IN3(n9111), .IN4(n9112), .QN(
        n9102) );
  NAND2X0 U9033 ( .IN1(g100), .IN2(n8947), .QN(n9112) );
  AND3X1 U9034 ( .IN1(n9113), .IN2(g28), .IN3(n9114), .Q(n8947) );
  NOR2X0 U9035 ( .IN1(n9115), .IN2(n9116), .QN(n9111) );
  NOR2X0 U9036 ( .IN1(n5842), .IN2(n8904), .QN(n9116) );
  NAND4X0 U9037 ( .IN1(n9117), .IN2(test_so25), .IN3(n7685), .IN4(n5324), .QN(
        n8904) );
  INVX0 U9038 ( .INP(n9009), .ZN(n9115) );
  NAND4X0 U9039 ( .IN1(n9117), .IN2(g28), .IN3(g19), .IN4(n5477), .QN(n9009)
         );
  NAND2X0 U9040 ( .IN1(n8946), .IN2(g2890), .QN(n9110) );
  AND2X1 U9041 ( .IN1(n9118), .IN2(n9113), .Q(n8946) );
  NAND2X0 U9042 ( .IN1(n8982), .IN2(g781), .QN(n9109) );
  INVX0 U9043 ( .INP(n8941), .ZN(n8982) );
  NOR2X0 U9044 ( .IN1(n5640), .IN2(n8930), .QN(n9098) );
  NAND2X0 U9045 ( .IN1(n9119), .IN2(n9118), .QN(n8930) );
  AND3X1 U9046 ( .IN1(n9120), .IN2(n8537), .IN3(n8202), .Q(n8928) );
  NAND4X0 U9047 ( .IN1(n8941), .IN2(n8942), .IN3(n8952), .IN4(n8951), .QN(
        n9120) );
  NAND2X0 U9048 ( .IN1(n9121), .IN2(n9118), .QN(n8941) );
  NOR2X0 U9049 ( .IN1(n9122), .IN2(n9123), .QN(n9096) );
  NOR2X0 U9050 ( .IN1(n5377), .IN2(n8926), .QN(n9123) );
  NOR2X0 U9051 ( .IN1(n8927), .IN2(DFF_206_n1), .QN(n9122) );
  NAND2X0 U9052 ( .IN1(test_so64), .IN2(n9124), .QN(n9095) );
  OR2X1 U9053 ( .IN1(n8924), .IN2(n14520), .Q(n9094) );
  OR2X1 U9054 ( .IN1(g34970), .IN2(n7810), .Q(g34913) );
  NAND4X0 U9055 ( .IN1(n9125), .IN2(n9126), .IN3(n9127), .IN4(n9128), .QN(
        g34970) );
  NOR4X0 U9056 ( .IN1(n9129), .IN2(n9130), .IN3(n9131), .IN4(n9132), .QN(n9128) );
  NOR2X0 U9057 ( .IN1(n5408), .IN2(n8996), .QN(n9132) );
  NAND3X0 U9058 ( .IN1(n9118), .IN2(n8202), .IN3(n2527), .QN(n8996) );
  NOR2X0 U9059 ( .IN1(n5312), .IN2(n8997), .QN(n9131) );
  NAND3X0 U9060 ( .IN1(n8202), .IN2(n9133), .IN3(n2527), .QN(n8997) );
  NOR2X0 U9061 ( .IN1(n5641), .IN2(n8926), .QN(n9130) );
  NAND3X0 U9062 ( .IN1(n9114), .IN2(n5324), .IN3(n9119), .QN(n8926) );
  NOR2X0 U9063 ( .IN1(n8927), .IN2(DFF_514_n1), .QN(n9129) );
  NAND2X0 U9064 ( .IN1(n9053), .IN2(n9134), .QN(n8927) );
  NOR2X0 U9066 ( .IN1(n9135), .IN2(n9136), .QN(n9127) );
  NOR2X0 U9067 ( .IN1(n5644), .IN2(n8987), .QN(n9136) );
  NAND2X0 U9068 ( .IN1(n9119), .IN2(n9133), .QN(n8987) );
  NOR4X0 U9069 ( .IN1(n9053), .IN2(n5468), .IN3(n7685), .IN4(test_so25), .QN(
        n9119) );
  NOR2X0 U9071 ( .IN1(n9137), .IN2(n9053), .QN(n9135) );
  NOR4X0 U9072 ( .IN1(n9138), .IN2(n9139), .IN3(n9140), .IN4(n9141), .QN(n9137) );
  NOR2X0 U9073 ( .IN1(n14519), .IN2(n8951), .QN(n9141) );
  NOR2X0 U9074 ( .IN1(n5476), .IN2(n8952), .QN(n9140) );
  NAND3X0 U9077 ( .IN1(n9142), .IN2(n9087), .IN3(n9143), .QN(n9139) );
  NAND2X0 U9078 ( .IN1(n9068), .IN2(g776), .QN(n9143) );
  INVX0 U9079 ( .INP(n8942), .ZN(n9068) );
  NAND2X0 U9081 ( .IN1(n8636), .IN2(n9144), .QN(n9087) );
  NAND3X0 U9082 ( .IN1(n8952), .IN2(n8951), .IN3(n8942), .QN(n9144) );
  NAND3X0 U9083 ( .IN1(n9114), .IN2(g28), .IN3(n9121), .QN(n8942) );
  NAND2X0 U9087 ( .IN1(n2552), .IN2(n9133), .QN(n8951) );
  NAND3X0 U9088 ( .IN1(n2552), .IN2(n5324), .IN3(n9114), .QN(n8952) );
  NOR2X0 U9089 ( .IN1(n9145), .IN2(n5469), .QN(n9114) );
  NAND2X0 U9091 ( .IN1(n8940), .IN2(g538), .QN(n9142) );
  INVX0 U9092 ( .INP(n8978), .ZN(n8940) );
  NAND2X0 U9093 ( .IN1(n9121), .IN2(n9133), .QN(n8978) );
  AND2X1 U9094 ( .IN1(n9146), .IN2(n5468), .Q(n9121) );
  NAND4X0 U9095 ( .IN1(n9147), .IN2(n9148), .IN3(n9149), .IN4(n9150), .QN(
        n9138) );
  NAND2X0 U9096 ( .IN1(n9067), .IN2(g2902), .QN(n9150) );
  INVX0 U9097 ( .INP(n8953), .ZN(n9067) );
  NAND3X0 U9100 ( .IN1(n9146), .IN2(n5324), .IN3(n9117), .QN(n8953) );
  NAND2X0 U9102 ( .IN1(n9043), .IN2(g2844), .QN(n9149) );
  INVX0 U9103 ( .INP(n8958), .ZN(n9043) );
  NAND3X0 U9104 ( .IN1(n9133), .IN2(g9), .IN3(n9146), .QN(n8958) );
  NAND2X0 U9105 ( .IN1(test_so1), .IN2(n8986), .QN(n9148) );
  INVX0 U9106 ( .INP(n8957), .ZN(n8986) );
  NAND3X0 U9108 ( .IN1(n9146), .IN2(g28), .IN3(n9117), .QN(n8957) );
  NOR4X0 U9109 ( .IN1(n8219), .IN2(n9151), .IN3(n5468), .IN4(n7766), .QN(n9117) );
  INVX0 U9110 ( .INP(n3395), .ZN(n9151) );
  NAND2X0 U9112 ( .IN1(n8954), .IN2(g2848), .QN(n9147) );
  AND3X1 U9113 ( .IN1(n9118), .IN2(g9), .IN3(n9146), .Q(n8954) );
  NOR2X0 U9114 ( .IN1(g19), .IN2(test_so25), .QN(n9146) );
  NAND2X0 U9115 ( .IN1(n9093), .IN2(g1300), .QN(n9126) );
  INVX0 U9117 ( .INP(n9027), .ZN(n9093) );
  NAND2X0 U9118 ( .IN1(n2549), .IN2(n9124), .QN(n9027) );
  INVX0 U9119 ( .INP(n8925), .ZN(n9124) );
  NAND3X0 U9121 ( .IN1(n9133), .IN2(n9113), .IN3(n8202), .QN(n8925) );
  NOR3X0 U9122 ( .IN1(g19), .IN2(g9), .IN3(n5477), .QN(n9113) );
  AND3X1 U9123 ( .IN1(n5324), .IN2(n9152), .IN3(n5469), .Q(n9133) );
  NAND2X0 U9125 ( .IN1(n9028), .IN2(g956), .QN(n9125) );
  NOR2X0 U9126 ( .IN1(g947), .IN2(n8924), .QN(n9028) );
  NAND3X0 U9127 ( .IN1(n9118), .IN2(n8202), .IN3(n2552), .QN(n8924) );
  INVX0 U9129 ( .INP(n9053), .ZN(n8202) );
  NAND4X0 U9130 ( .IN1(g54), .IN2(n9134), .IN3(n9153), .IN4(n8915), .QN(n9053)
         );
  INVX0 U9131 ( .INP(g56), .ZN(n8915) );
  NOR2X0 U9133 ( .IN1(test_so74), .IN2(g57), .QN(n9153) );
  INVX0 U9134 ( .INP(g53), .ZN(n9134) );
  AND3X1 U9135 ( .IN1(n9152), .IN2(g28), .IN3(n5469), .Q(n9118) );
  INVX0 U9137 ( .INP(n9145), .ZN(n9152) );
  NAND3X0 U9138 ( .IN1(n7765), .IN2(n8219), .IN3(n7766), .QN(n9145) );
  NAND2X0 U9139 ( .IN1(n9154), .IN2(n9155), .QN(g34911) );
  NAND2X0 U9140 ( .IN1(n9156), .IN2(g807), .QN(n9155) );
  NAND2X0 U9141 ( .IN1(n8511), .IN2(n9157), .QN(n9156) );
  NAND2X0 U9142 ( .IN1(n2404), .IN2(g554), .QN(n9154) );
  NAND2X0 U9143 ( .IN1(n9158), .IN2(n9159), .QN(g34882) );
  OR2X1 U9144 ( .IN1(n8480), .IN2(n8000), .Q(n9159) );
  NAND2X0 U9145 ( .IN1(n9160), .IN2(n8521), .QN(n9158) );
  NAND3X0 U9146 ( .IN1(n9161), .IN2(n9162), .IN3(n9163), .QN(n9160) );
  NAND3X0 U9147 ( .IN1(n5653), .IN2(n9164), .IN3(n9165), .QN(n9163) );
  OR2X1 U9148 ( .IN1(n9166), .IN2(g4358), .Q(n9164) );
  NAND3X0 U9149 ( .IN1(test_so81), .IN2(g4340), .IN3(g4358), .QN(n9162) );
  NAND3X0 U9150 ( .IN1(n9166), .IN2(n8208), .IN3(n5348), .QN(n9161) );
  NAND4X0 U9151 ( .IN1(n5653), .IN2(n8208), .IN3(n9167), .IN4(n9168), .QN(
        n9166) );
  NAND2X0 U9152 ( .IN1(n5540), .IN2(n9169), .QN(n9168) );
  NAND3X0 U9153 ( .IN1(n9170), .IN2(n9171), .IN3(n9172), .QN(n9169) );
  NAND2X0 U9154 ( .IN1(n8134), .IN2(g4322), .QN(n9171) );
  NAND3X0 U9155 ( .IN1(g90), .IN2(n5634), .IN3(n5506), .QN(n9170) );
  NAND3X0 U9156 ( .IN1(n5506), .IN2(g4311), .IN3(g4332), .QN(n9167) );
  NAND3X0 U9157 ( .IN1(n9173), .IN2(n9174), .IN3(n9175), .QN(g34881) );
  NAND2X0 U9158 ( .IN1(n8636), .IN2(g794), .QN(n9175) );
  NAND3X0 U9159 ( .IN1(n2404), .IN2(n9157), .IN3(g807), .QN(n9174) );
  INVX0 U9160 ( .INP(n2405), .ZN(n9157) );
  NAND2X0 U9161 ( .IN1(n2405), .IN2(n5479), .QN(n9173) );
  NAND3X0 U9162 ( .IN1(n9176), .IN2(n9177), .IN3(n9178), .QN(g34880) );
  NAND2X0 U9163 ( .IN1(n8636), .IN2(g626), .QN(n9178) );
  NAND3X0 U9164 ( .IN1(n2421), .IN2(n9179), .IN3(n9340), .QN(n9177) );
  INVX0 U9165 ( .INP(n2422), .ZN(n9179) );
  NAND2X0 U9166 ( .IN1(n2422), .IN2(n14519), .QN(n9176) );
  NAND3X0 U9167 ( .IN1(n9180), .IN2(n9181), .IN3(n9182), .QN(g34850) );
  NAND2X0 U9168 ( .IN1(n8635), .IN2(g790), .QN(n9182) );
  NAND3X0 U9169 ( .IN1(n2404), .IN2(n9183), .IN3(g794), .QN(n9181) );
  INVX0 U9170 ( .INP(n2419), .ZN(n9183) );
  NAND2X0 U9171 ( .IN1(n2419), .IN2(n5291), .QN(n9180) );
  NAND3X0 U9172 ( .IN1(n9184), .IN2(n9185), .IN3(n9186), .QN(g34849) );
  NAND2X0 U9173 ( .IN1(n8635), .IN2(g622), .QN(n9186) );
  NAND3X0 U9174 ( .IN1(n2421), .IN2(n9187), .IN3(g626), .QN(n9185) );
  INVX0 U9175 ( .INP(n2423), .ZN(n9187) );
  NAND2X0 U9176 ( .IN1(n2423), .IN2(n5288), .QN(n9184) );
  INVX0 U9177 ( .INP(n9188), .ZN(g34843) );
  NOR2X0 U9178 ( .IN1(n7999), .IN2(n9189), .QN(g34839) );
  AND3X1 U9179 ( .IN1(n9190), .IN2(n9191), .IN3(n8000), .Q(n9189) );
  NAND2X0 U9180 ( .IN1(n5540), .IN2(n9192), .QN(n9191) );
  NAND3X0 U9181 ( .IN1(n9193), .IN2(n9194), .IN3(n5323), .QN(n9192) );
  NAND2X0 U9182 ( .IN1(n9195), .IN2(g4332), .QN(n9190) );
  NAND3X0 U9183 ( .IN1(n5323), .IN2(n9193), .IN3(g73), .QN(n9195) );
  NAND2X0 U9184 ( .IN1(n9196), .IN2(n9197), .QN(g34808) );
  NAND2X0 U9185 ( .IN1(n8635), .IN2(g2955), .QN(n9197) );
  NAND2X0 U9186 ( .IN1(n9198), .IN2(n8523), .QN(n9196) );
  NAND3X0 U9187 ( .IN1(g91), .IN2(n9199), .IN3(n7819), .QN(n9198) );
  NAND2X0 U9188 ( .IN1(n9200), .IN2(n9201), .QN(g34807) );
  OR2X1 U9189 ( .IN1(n8480), .IN2(n8172), .Q(n9201) );
  NAND2X0 U9190 ( .IN1(n9202), .IN2(n8523), .QN(n9200) );
  NAND4X0 U9191 ( .IN1(n9203), .IN2(n9204), .IN3(n9205), .IN4(n9206), .QN(
        n9202) );
  NOR4X0 U9192 ( .IN1(n9207), .IN2(n9208), .IN3(g2955), .IN4(g2946), .QN(n9206) );
  NOR2X0 U9193 ( .IN1(n9209), .IN2(n9210), .QN(n9205) );
  NAND2X0 U9194 ( .IN1(n9211), .IN2(n9212), .QN(g34806) );
  NAND2X0 U9195 ( .IN1(n8635), .IN2(g2927), .QN(n9212) );
  NAND2X0 U9196 ( .IN1(n9213), .IN2(n8523), .QN(n9211) );
  NAND3X0 U9197 ( .IN1(n8181), .IN2(n8172), .IN3(n8182), .QN(n9213) );
  NOR2X0 U9198 ( .IN1(n8569), .IN2(n9214), .QN(g34805) );
  AND2X1 U9199 ( .IN1(n8179), .IN2(n8180), .Q(n9214) );
  NAND2X0 U9200 ( .IN1(n9215), .IN2(n9216), .QN(g34804) );
  OR2X1 U9201 ( .IN1(n8481), .IN2(n7819), .Q(n9216) );
  NAND2X0 U9202 ( .IN1(n9217), .IN2(n8522), .QN(n9215) );
  NAND3X0 U9203 ( .IN1(g962), .IN2(g1306), .IN3(n5750), .QN(n9217) );
  NAND2X0 U9204 ( .IN1(n9218), .IN2(n9219), .QN(g34803) );
  NAND2X0 U9205 ( .IN1(n8635), .IN2(g2917), .QN(n9219) );
  NAND2X0 U9206 ( .IN1(n9220), .IN2(n8522), .QN(n9218) );
  NAND3X0 U9207 ( .IN1(g44), .IN2(n8179), .IN3(n7816), .QN(n9220) );
  NAND2X0 U9208 ( .IN1(n9221), .IN2(n9222), .QN(g34802) );
  NAND2X0 U9209 ( .IN1(n8635), .IN2(g2902), .QN(n9222) );
  NAND2X0 U9210 ( .IN1(n9223), .IN2(n8522), .QN(n9221) );
  NAND3X0 U9211 ( .IN1(n9224), .IN2(n9225), .IN3(n7817), .QN(n9223) );
  NAND2X0 U9212 ( .IN1(n9226), .IN2(n9227), .QN(g34801) );
  NAND2X0 U9213 ( .IN1(n8635), .IN2(g2970), .QN(n9227) );
  NAND2X0 U9214 ( .IN1(n9228), .IN2(n8522), .QN(n9226) );
  NAND4X0 U9215 ( .IN1(n8184), .IN2(n7818), .IN3(n5595), .IN4(g691), .QN(n9228) );
  NAND2X0 U9216 ( .IN1(n9229), .IN2(n9230), .QN(g34800) );
  NAND2X0 U9217 ( .IN1(n8634), .IN2(g2886), .QN(n9230) );
  NAND2X0 U9218 ( .IN1(n9231), .IN2(n8522), .QN(n9229) );
  OR2X1 U9219 ( .IN1(test_so74), .IN2(test_so14), .Q(n9231) );
  NAND2X0 U9220 ( .IN1(n9232), .IN2(n9233), .QN(g34799) );
  NAND2X0 U9221 ( .IN1(n8634), .IN2(g2873), .QN(n9233) );
  NAND2X0 U9222 ( .IN1(n9234), .IN2(n8522), .QN(n9232) );
  NAND2X0 U9223 ( .IN1(n8178), .IN2(g44), .QN(n9234) );
  NAND2X0 U9224 ( .IN1(n9235), .IN2(n9237), .QN(g34798) );
  NAND2X0 U9225 ( .IN1(n8634), .IN2(g2878), .QN(n9237) );
  NAND2X0 U9226 ( .IN1(n9238), .IN2(n8522), .QN(n9235) );
  NAND2X0 U9227 ( .IN1(n8174), .IN2(n8175), .QN(n9238) );
  NAND2X0 U9228 ( .IN1(n9239), .IN2(n9241), .QN(g34797) );
  NAND2X0 U9229 ( .IN1(n8634), .IN2(g2882), .QN(n9241) );
  NAND2X0 U9230 ( .IN1(n9242), .IN2(n8522), .QN(n9239) );
  NAND2X0 U9231 ( .IN1(n8173), .IN2(g91), .QN(n9242) );
  NAND2X0 U9232 ( .IN1(n9243), .IN2(n9244), .QN(g34796) );
  NAND2X0 U9233 ( .IN1(n8634), .IN2(g2898), .QN(n9244) );
  NAND2X0 U9234 ( .IN1(n9246), .IN2(n8522), .QN(n9243) );
  NAND2X0 U9235 ( .IN1(n7677), .IN2(n9199), .QN(n9246) );
  NOR2X0 U9236 ( .IN1(n9248), .IN2(n9249), .QN(n9199) );
  NAND2X0 U9237 ( .IN1(n9250), .IN2(n9251), .QN(g34795) );
  NAND2X0 U9238 ( .IN1(n8634), .IN2(g2864), .QN(n9251) );
  NAND2X0 U9239 ( .IN1(n9252), .IN2(n8522), .QN(n9250) );
  OR2X1 U9240 ( .IN1(g2898), .IN2(n9209), .Q(n9252) );
  NAND4X0 U9241 ( .IN1(n5882), .IN2(n5861), .IN3(n9253), .IN4(n9254), .QN(
        n9209) );
  NAND2X0 U9242 ( .IN1(n9256), .IN2(n9257), .QN(g34794) );
  NAND2X0 U9243 ( .IN1(n8634), .IN2(g2856), .QN(n9257) );
  NAND2X0 U9244 ( .IN1(n9258), .IN2(n8522), .QN(n9256) );
  OR2X1 U9245 ( .IN1(g2864), .IN2(n9210), .Q(n9258) );
  NAND2X0 U9246 ( .IN1(n9259), .IN2(n9260), .QN(n9210) );
  NAND2X0 U9247 ( .IN1(n9261), .IN2(n9263), .QN(g34793) );
  NAND2X0 U9248 ( .IN1(n8633), .IN2(g2848), .QN(n9263) );
  NAND2X0 U9249 ( .IN1(n9264), .IN2(n8522), .QN(n9261) );
  OR3X1 U9250 ( .IN1(n9207), .IN2(n9266), .IN3(g2856), .Q(n9264) );
  NAND2X0 U9251 ( .IN1(n9268), .IN2(n9269), .QN(g34792) );
  NAND2X0 U9252 ( .IN1(n8633), .IN2(g29214), .QN(n9269) );
  NAND2X0 U9253 ( .IN1(n9270), .IN2(n8522), .QN(n9268) );
  OR3X1 U9254 ( .IN1(n9208), .IN2(n9271), .IN3(g2848), .Q(n9270) );
  NAND3X0 U9255 ( .IN1(n9272), .IN2(n9275), .IN3(n9277), .QN(g34791) );
  NAND2X0 U9256 ( .IN1(n8633), .IN2(g785), .QN(n9277) );
  NAND3X0 U9257 ( .IN1(n2404), .IN2(n9278), .IN3(g790), .QN(n9275) );
  INVX0 U9258 ( .INP(n2425), .ZN(n9278) );
  NAND2X0 U9259 ( .IN1(n2425), .IN2(n5292), .QN(n9272) );
  NAND3X0 U9260 ( .IN1(n9279), .IN2(n9282), .IN3(n9283), .QN(g34790) );
  NAND2X0 U9261 ( .IN1(n8633), .IN2(g617), .QN(n9283) );
  NAND3X0 U9262 ( .IN1(n2421), .IN2(n9284), .IN3(g622), .QN(n9282) );
  INVX0 U9263 ( .INP(n2427), .ZN(n9284) );
  NAND2X0 U9264 ( .IN1(n2427), .IN2(n5672), .QN(n9279) );
  NOR2X0 U9265 ( .IN1(n5305), .IN2(n9285), .QN(g34788) );
  AND2X1 U9266 ( .IN1(g479), .IN2(n3195), .Q(n9285) );
  NAND2X0 U9267 ( .IN1(n9286), .IN2(n9287), .QN(g34783) );
  NAND3X0 U9268 ( .IN1(n9288), .IN2(n9289), .IN3(n9290), .QN(n9287) );
  NAND3X0 U9269 ( .IN1(n9291), .IN2(n9292), .IN3(n9293), .QN(n9286) );
  NAND2X0 U9270 ( .IN1(n9296), .IN2(n9297), .QN(g34735) );
  OR2X1 U9271 ( .IN1(n8481), .IN2(n7727), .Q(n9297) );
  NAND2X0 U9272 ( .IN1(n9298), .IN2(n8522), .QN(n9296) );
  NAND2X0 U9273 ( .IN1(n5639), .IN2(n8177), .QN(n9298) );
  NAND2X0 U9274 ( .IN1(n9299), .IN2(n9300), .QN(g34734) );
  NAND2X0 U9275 ( .IN1(n8633), .IN2(g4172), .QN(n9300) );
  NAND2X0 U9276 ( .IN1(n9301), .IN2(n8522), .QN(n9299) );
  NAND2X0 U9277 ( .IN1(n5494), .IN2(n8181), .QN(n9301) );
  NOR2X0 U9278 ( .IN1(n8572), .IN2(n9304), .QN(g34733) );
  NOR2X0 U9279 ( .IN1(g4153), .IN2(g4172), .QN(n9304) );
  NAND2X0 U9280 ( .IN1(n9305), .IN2(n9307), .QN(g34732) );
  NAND2X0 U9281 ( .IN1(n8510), .IN2(g2994), .QN(n9307) );
  NAND2X0 U9282 ( .IN1(n8633), .IN2(g2999), .QN(n9305) );
  NAND2X0 U9283 ( .IN1(n9308), .IN2(n9309), .QN(g34731) );
  OR2X1 U9284 ( .IN1(n8480), .IN2(n5635), .Q(n9309) );
  NAND2X0 U9285 ( .IN1(n9310), .IN2(n8522), .QN(n9308) );
  OR2X1 U9286 ( .IN1(n9311), .IN2(test_so64), .Q(n9310) );
  NAND2X0 U9287 ( .IN1(n9313), .IN2(n9315), .QN(g34730) );
  NAND2X0 U9288 ( .IN1(n8633), .IN2(g1296), .QN(n9315) );
  NAND2X0 U9289 ( .IN1(n9316), .IN2(n8522), .QN(n9313) );
  NAND2X0 U9290 ( .IN1(n8183), .IN2(n5635), .QN(n9316) );
  OR3X1 U9291 ( .IN1(n9317), .IN2(n9318), .IN3(n2499), .Q(g34729) );
  NOR2X0 U9292 ( .IN1(n2549), .IN2(n8504), .QN(n9318) );
  NOR2X0 U9293 ( .IN1(n8573), .IN2(g1306), .QN(n9317) );
  NAND2X0 U9294 ( .IN1(n9319), .IN2(n9320), .QN(g34728) );
  OR2X1 U9295 ( .IN1(n8481), .IN2(n5415), .Q(n9320) );
  NAND2X0 U9296 ( .IN1(n9321), .IN2(n8522), .QN(n9319) );
  NAND2X0 U9297 ( .IN1(n14520), .IN2(n9224), .QN(n9321) );
  NAND2X0 U9298 ( .IN1(n9323), .IN2(n9326), .QN(g34727) );
  NAND2X0 U9299 ( .IN1(n8632), .IN2(g952), .QN(n9326) );
  NAND2X0 U9300 ( .IN1(n9328), .IN2(n8522), .QN(n9323) );
  NAND2X0 U9301 ( .IN1(n5415), .IN2(n8188), .QN(n9328) );
  OR3X1 U9302 ( .IN1(n9329), .IN2(n9330), .IN3(n2505), .Q(g34726) );
  NOR2X0 U9303 ( .IN1(n5286), .IN2(n8505), .QN(n9330) );
  NOR2X0 U9304 ( .IN1(n8573), .IN2(g962), .QN(n9329) );
  NAND3X0 U9305 ( .IN1(n9331), .IN2(n9333), .IN3(n9334), .QN(g34725) );
  NAND2X0 U9306 ( .IN1(n8632), .IN2(g781), .QN(n9334) );
  NAND3X0 U9307 ( .IN1(n2404), .IN2(n9335), .IN3(g785), .QN(n9333) );
  INVX0 U9308 ( .INP(n2485), .ZN(n9335) );
  NAND2X0 U9309 ( .IN1(n2485), .IN2(n5293), .QN(n9331) );
  NAND3X0 U9310 ( .IN1(n9337), .IN2(n9338), .IN3(n9339), .QN(g34724) );
  NAND2X0 U9311 ( .IN1(n8632), .IN2(g613), .QN(n9339) );
  NAND3X0 U9312 ( .IN1(n2421), .IN2(n9341), .IN3(g617), .QN(n9338) );
  INVX0 U9313 ( .INP(n2487), .ZN(n9341) );
  NAND2X0 U9314 ( .IN1(n2487), .IN2(n5339), .QN(n9337) );
  NAND2X0 U9316 ( .IN1(n9342), .IN2(n9343), .QN(g34723) );
  NAND2X0 U9317 ( .IN1(test_so41), .IN2(n8562), .QN(n9343) );
  NAND2X0 U9318 ( .IN1(n9344), .IN2(n8522), .QN(n9342) );
  NAND2X0 U9319 ( .IN1(n5490), .IN2(n8184), .QN(n9344) );
  NAND2X0 U9320 ( .IN1(n9345), .IN2(n9346), .QN(g34722) );
  NAND2X0 U9321 ( .IN1(n8632), .IN2(g538), .QN(n9346) );
  NAND2X0 U9322 ( .IN1(n9347), .IN2(n8522), .QN(n9345) );
  NAND2X0 U9323 ( .IN1(n5492), .IN2(g691), .QN(n9347) );
  NAND2X0 U9324 ( .IN1(n9349), .IN2(n9350), .QN(g34721) );
  NAND2X0 U9325 ( .IN1(g29221), .IN2(n8557), .QN(n9350) );
  NAND2X0 U9326 ( .IN1(n9353), .IN2(n8521), .QN(n9349) );
  NAND2X0 U9327 ( .IN1(n8187), .IN2(n8186), .QN(n9353) );
  NAND2X0 U9328 ( .IN1(n9354), .IN2(n9355), .QN(g34720) );
  OR2X1 U9329 ( .IN1(n8480), .IN2(n5490), .Q(n9355) );
  NAND2X0 U9330 ( .IN1(n9356), .IN2(n8521), .QN(n9354) );
  NAND2X0 U9331 ( .IN1(n8185), .IN2(g29212), .QN(n9356) );
  NOR2X0 U9332 ( .IN1(n8574), .IN2(n9358), .QN(g34719) );
  NOR2X0 U9333 ( .IN1(g209), .IN2(g538), .QN(n9358) );
  NOR2X0 U9334 ( .IN1(n5497), .IN2(n8560), .QN(g34647) );
  NOR2X0 U9335 ( .IN1(n5644), .IN2(n8559), .QN(g34646) );
  NOR2X0 U9336 ( .IN1(n5499), .IN2(n8560), .QN(g34645) );
  NOR2X0 U9337 ( .IN1(n5643), .IN2(n8559), .QN(g34644) );
  NOR2X0 U9338 ( .IN1(n5498), .IN2(n8559), .QN(g34643) );
  NAND2X0 U9339 ( .IN1(n9359), .IN2(n9360), .QN(g34642) );
  NAND2X0 U9340 ( .IN1(n8510), .IN2(g4927), .QN(n9360) );
  NAND2X0 U9341 ( .IN1(n8632), .IN2(g4912), .QN(n9359) );
  NAND2X0 U9342 ( .IN1(n9361), .IN2(n9362), .QN(g34641) );
  NAND2X0 U9343 ( .IN1(n8511), .IN2(g4912), .QN(n9362) );
  NAND2X0 U9344 ( .IN1(n8632), .IN2(g4907), .QN(n9361) );
  NAND2X0 U9345 ( .IN1(n9363), .IN2(n9364), .QN(g34640) );
  NAND2X0 U9346 ( .IN1(n8510), .IN2(g4907), .QN(n9364) );
  NAND2X0 U9347 ( .IN1(n8632), .IN2(g4922), .QN(n9363) );
  NAND2X0 U9348 ( .IN1(n9365), .IN2(n9366), .QN(g34639) );
  NAND2X0 U9349 ( .IN1(n8510), .IN2(g4922), .QN(n9366) );
  NAND2X0 U9350 ( .IN1(n8631), .IN2(g4917), .QN(n9365) );
  NOR2X0 U9351 ( .IN1(n5408), .IN2(n8558), .QN(g34638) );
  NAND2X0 U9352 ( .IN1(n9368), .IN2(n9369), .QN(g34637) );
  NAND2X0 U9353 ( .IN1(n8509), .IN2(g4737), .QN(n9369) );
  NAND2X0 U9354 ( .IN1(n8631), .IN2(g4722), .QN(n9368) );
  NAND2X0 U9355 ( .IN1(n9370), .IN2(n9371), .QN(g34636) );
  NAND2X0 U9356 ( .IN1(n8511), .IN2(g4722), .QN(n9371) );
  NAND2X0 U9357 ( .IN1(n8631), .IN2(g4717), .QN(n9370) );
  NAND2X0 U9358 ( .IN1(n9372), .IN2(n9373), .QN(g34635) );
  NAND2X0 U9359 ( .IN1(n8509), .IN2(g4717), .QN(n9373) );
  NAND2X0 U9360 ( .IN1(n8631), .IN2(g4732), .QN(n9372) );
  NAND2X0 U9361 ( .IN1(n9374), .IN2(n9375), .QN(g34634) );
  NAND2X0 U9362 ( .IN1(n8509), .IN2(g4732), .QN(n9375) );
  NAND2X0 U9363 ( .IN1(n8631), .IN2(g4727), .QN(n9374) );
  NOR2X0 U9364 ( .IN1(n5312), .IN2(n8557), .QN(g34633) );
  NAND2X0 U9365 ( .IN1(n9376), .IN2(n9377), .QN(g34632) );
  NAND2X0 U9366 ( .IN1(n8509), .IN2(g4245), .QN(n9377) );
  NAND2X0 U9367 ( .IN1(test_so67), .IN2(n8659), .QN(n9376) );
  NAND2X0 U9368 ( .IN1(n9378), .IN2(n9379), .QN(g34631) );
  NAND2X0 U9369 ( .IN1(test_so67), .IN2(n8521), .QN(n9379) );
  NAND2X0 U9370 ( .IN1(n8631), .IN2(g4253), .QN(n9378) );
  NAND2X0 U9371 ( .IN1(n9380), .IN2(n9381), .QN(g34630) );
  NAND2X0 U9372 ( .IN1(n8509), .IN2(g4253), .QN(n9381) );
  OR2X1 U9373 ( .IN1(n8479), .IN2(n5639), .Q(n9380) );
  NAND2X0 U9374 ( .IN1(n9382), .IN2(n9383), .QN(g34629) );
  NAND2X0 U9375 ( .IN1(n8510), .IN2(g4157), .QN(n9383) );
  NAND2X0 U9376 ( .IN1(n8631), .IN2(g4146), .QN(n9382) );
  NAND2X0 U9377 ( .IN1(n9384), .IN2(n9385), .QN(g34628) );
  NAND2X0 U9378 ( .IN1(n8509), .IN2(g4146), .QN(n9385) );
  OR2X1 U9379 ( .IN1(n8480), .IN2(n5494), .Q(n9384) );
  NOR2X0 U9380 ( .IN1(n5641), .IN2(n8556), .QN(g34627) );
  NOR2X0 U9381 ( .IN1(n8576), .IN2(n8227), .QN(g34626) );
  NOR2X0 U9382 ( .IN1(n5495), .IN2(n8556), .QN(g34625) );
  NAND2X0 U9383 ( .IN1(n9386), .IN2(n9387), .QN(g34624) );
  NAND2X0 U9384 ( .IN1(n8509), .IN2(g2988), .QN(n9387) );
  NAND2X0 U9385 ( .IN1(n8630), .IN2(g2994), .QN(n9386) );
  NAND2X0 U9386 ( .IN1(n9388), .IN2(n9389), .QN(g34623) );
  NAND2X0 U9387 ( .IN1(n8509), .IN2(g2970), .QN(n9389) );
  NAND2X0 U9388 ( .IN1(test_so22), .IN2(n8545), .QN(n9388) );
  NAND2X0 U9389 ( .IN1(n9390), .IN2(n9391), .QN(g34622) );
  NAND2X0 U9390 ( .IN1(test_so22), .IN2(n8521), .QN(n9391) );
  NAND2X0 U9391 ( .IN1(n8630), .IN2(g2950), .QN(n9390) );
  NAND2X0 U9392 ( .IN1(n9392), .IN2(n9393), .QN(g34621) );
  NAND2X0 U9393 ( .IN1(n8510), .IN2(g2950), .QN(n9393) );
  NAND2X0 U9394 ( .IN1(n8630), .IN2(g2936), .QN(n9392) );
  NAND2X0 U9395 ( .IN1(n9394), .IN2(n9395), .QN(g34620) );
  NAND2X0 U9396 ( .IN1(n8509), .IN2(g2936), .QN(n9395) );
  NAND2X0 U9397 ( .IN1(n8630), .IN2(g2922), .QN(n9394) );
  NAND2X0 U9398 ( .IN1(n9396), .IN2(n9397), .QN(g34619) );
  NAND2X0 U9399 ( .IN1(n8509), .IN2(g2922), .QN(n9397) );
  NAND2X0 U9400 ( .IN1(n8630), .IN2(g2912), .QN(n9396) );
  NAND2X0 U9401 ( .IN1(n9398), .IN2(n9399), .QN(g34618) );
  NAND2X0 U9402 ( .IN1(n8509), .IN2(g2912), .QN(n9399) );
  NAND2X0 U9403 ( .IN1(test_so1), .IN2(n8585), .QN(n9398) );
  NAND2X0 U9404 ( .IN1(n9400), .IN2(n9401), .QN(g34617) );
  NAND2X0 U9405 ( .IN1(test_so1), .IN2(n8523), .QN(n9401) );
  OR2X1 U9406 ( .IN1(n8479), .IN2(n5842), .Q(n9400) );
  NAND2X0 U9407 ( .IN1(n9402), .IN2(n9403), .QN(g34616) );
  NAND2X0 U9408 ( .IN1(n8509), .IN2(g2868), .QN(n9403) );
  NAND2X0 U9409 ( .IN1(n8630), .IN2(g2988), .QN(n9402) );
  NAND2X0 U9410 ( .IN1(n9404), .IN2(n9405), .QN(g34615) );
  NAND2X0 U9411 ( .IN1(n8509), .IN2(g2873), .QN(n9405) );
  NAND2X0 U9412 ( .IN1(n8630), .IN2(g2868), .QN(n9404) );
  NAND2X0 U9413 ( .IN1(n9406), .IN2(n9407), .QN(g34614) );
  NAND2X0 U9414 ( .IN1(n8509), .IN2(g29214), .QN(n9407) );
  NAND2X0 U9415 ( .IN1(g37), .IN2(n8576), .QN(n9406) );
  NAND2X0 U9416 ( .IN1(n9408), .IN2(n9409), .QN(g34613) );
  NAND2X0 U9417 ( .IN1(test_so95), .IN2(n8660), .QN(n9409) );
  NAND2X0 U9418 ( .IN1(g37), .IN2(n8521), .QN(n9408) );
  NAND2X0 U9419 ( .IN1(n9410), .IN2(n9411), .QN(g34612) );
  NAND2X0 U9420 ( .IN1(test_so95), .IN2(n8521), .QN(n9411) );
  NAND2X0 U9421 ( .IN1(n8629), .IN2(g2860), .QN(n9410) );
  NAND2X0 U9422 ( .IN1(n9412), .IN2(n9413), .QN(g34611) );
  NAND2X0 U9423 ( .IN1(n8510), .IN2(g2860), .QN(n9413) );
  NAND2X0 U9424 ( .IN1(n8629), .IN2(g2852), .QN(n9412) );
  NAND2X0 U9425 ( .IN1(n9414), .IN2(n9415), .QN(g34610) );
  NAND2X0 U9426 ( .IN1(n8510), .IN2(g2852), .QN(n9415) );
  NAND2X0 U9427 ( .IN1(n8629), .IN2(g2844), .QN(n9414) );
  NAND2X0 U9428 ( .IN1(n9416), .IN2(n9417), .QN(g34609) );
  NAND2X0 U9429 ( .IN1(n8510), .IN2(g2844), .QN(n9417) );
  NAND2X0 U9430 ( .IN1(n8629), .IN2(g2890), .QN(n9416) );
  NAND2X0 U9431 ( .IN1(n9418), .IN2(n9419), .QN(g34608) );
  NAND2X0 U9432 ( .IN1(n8509), .IN2(g2704), .QN(n9419) );
  NAND2X0 U9433 ( .IN1(n8629), .IN2(g2697), .QN(n9418) );
  NAND2X0 U9434 ( .IN1(n9420), .IN2(n9421), .QN(g34607) );
  NAND2X0 U9435 ( .IN1(n8510), .IN2(g2697), .QN(n9421) );
  NAND2X0 U9436 ( .IN1(n8629), .IN2(g2689), .QN(n9420) );
  NOR2X0 U9437 ( .IN1(n5347), .IN2(n8555), .QN(g34606) );
  NAND2X0 U9438 ( .IN1(n9422), .IN2(n9423), .QN(g34605) );
  NAND2X0 U9439 ( .IN1(n8509), .IN2(g2145), .QN(n9423) );
  NAND2X0 U9440 ( .IN1(n8629), .IN2(g2138), .QN(n9422) );
  NAND2X0 U9441 ( .IN1(n9424), .IN2(n9425), .QN(g34604) );
  NAND2X0 U9442 ( .IN1(n8510), .IN2(g2138), .QN(n9425) );
  NAND2X0 U9443 ( .IN1(n8628), .IN2(g2130), .QN(n9424) );
  NOR2X0 U9444 ( .IN1(n5487), .IN2(n8554), .QN(g34603) );
  NOR2X0 U9445 ( .IN1(n2549), .IN2(n8552), .QN(g34602) );
  NOR2X0 U9446 ( .IN1(n5286), .IN2(n8552), .QN(g34601) );
  NAND3X0 U9447 ( .IN1(n9426), .IN2(n9427), .IN3(n9428), .QN(g34600) );
  NAND2X0 U9448 ( .IN1(n8628), .IN2(g776), .QN(n9428) );
  NAND3X0 U9449 ( .IN1(n2404), .IN2(n9429), .IN3(g781), .QN(n9427) );
  INVX0 U9450 ( .INP(n2507), .ZN(n9429) );
  NAND2X0 U9451 ( .IN1(n2507), .IN2(n5551), .QN(n9426) );
  NAND3X0 U9452 ( .IN1(n9430), .IN2(n9431), .IN3(n9432), .QN(g34599) );
  NAND2X0 U9454 ( .IN1(n8628), .IN2(g608), .QN(n9432) );
  NAND3X0 U9455 ( .IN1(n2421), .IN2(n9433), .IN3(g613), .QN(n9431) );
  INVX0 U9456 ( .INP(n2509), .ZN(n9433) );
  NAND2X0 U9457 ( .IN1(n2509), .IN2(n5474), .QN(n9430) );
  NAND2X0 U9458 ( .IN1(n9434), .IN2(n9435), .QN(g34598) );
  NAND2X0 U9459 ( .IN1(n8628), .IN2(g550), .QN(n9435) );
  NAND2X0 U9460 ( .IN1(g29221), .IN2(n8521), .QN(n9434) );
  NAND2X0 U9461 ( .IN1(n9436), .IN2(n9437), .QN(g34468) );
  NAND2X0 U9462 ( .IN1(n9438), .IN2(g4854), .QN(n9437) );
  NAND2X0 U9463 ( .IN1(n9439), .IN2(n8521), .QN(n9438) );
  NAND2X0 U9464 ( .IN1(n9440), .IN2(n9441), .QN(n9439) );
  NAND2X0 U9465 ( .IN1(n9442), .IN2(g4859), .QN(n9436) );
  NAND2X0 U9466 ( .IN1(n9443), .IN2(n9444), .QN(g34467) );
  NAND2X0 U9467 ( .IN1(n9445), .IN2(n9442), .QN(n9444) );
  XOR2X1 U9468 ( .IN1(g4854), .IN2(n9441), .Q(n9445) );
  AND2X1 U9469 ( .IN1(n2563), .IN2(g4849), .Q(n9441) );
  NAND2X0 U9470 ( .IN1(n8628), .IN2(g4849), .QN(n9443) );
  NAND2X0 U9471 ( .IN1(n9446), .IN2(n9447), .QN(g34466) );
  NAND2X0 U9472 ( .IN1(n9448), .IN2(g4878), .QN(n9447) );
  NAND2X0 U9473 ( .IN1(n9449), .IN2(n8521), .QN(n9448) );
  NAND2X0 U9474 ( .IN1(n7796), .IN2(n9440), .QN(n9449) );
  NAND3X0 U9475 ( .IN1(n9442), .IN2(g4843), .IN3(n5283), .QN(n9446) );
  NAND3X0 U9476 ( .IN1(n9450), .IN2(n9451), .IN3(n9452), .QN(g34465) );
  NAND2X0 U9477 ( .IN1(n8628), .IN2(g4843), .QN(n9452) );
  NAND3X0 U9478 ( .IN1(n9440), .IN2(n2563), .IN3(n8151), .QN(n9451) );
  NAND2X0 U9479 ( .IN1(n2567), .IN2(n9442), .QN(n9450) );
  INVX0 U9480 ( .INP(n9453), .ZN(n9442) );
  NAND2X0 U9481 ( .IN1(n9454), .IN2(n9455), .QN(g34464) );
  NAND2X0 U9482 ( .IN1(n9456), .IN2(g4664), .QN(n9455) );
  NAND2X0 U9483 ( .IN1(n9457), .IN2(n8521), .QN(n9456) );
  NAND2X0 U9484 ( .IN1(n9458), .IN2(n9459), .QN(n9457) );
  NAND2X0 U9485 ( .IN1(n9460), .IN2(g4669), .QN(n9454) );
  NAND2X0 U9486 ( .IN1(n9461), .IN2(n9462), .QN(g34463) );
  NAND2X0 U9487 ( .IN1(n9463), .IN2(n9460), .QN(n9462) );
  XOR2X1 U9488 ( .IN1(g4664), .IN2(n9459), .Q(n9463) );
  AND2X1 U9489 ( .IN1(n2573), .IN2(g4659), .Q(n9459) );
  NAND2X0 U9490 ( .IN1(n8628), .IN2(g4659), .QN(n9461) );
  NAND2X0 U9491 ( .IN1(n9464), .IN2(n9465), .QN(g34462) );
  NAND2X0 U9492 ( .IN1(n9466), .IN2(g4688), .QN(n9465) );
  NAND2X0 U9493 ( .IN1(n9467), .IN2(n8521), .QN(n9466) );
  NAND2X0 U9494 ( .IN1(n9458), .IN2(n8239), .QN(n9467) );
  NAND3X0 U9495 ( .IN1(n9460), .IN2(test_so19), .IN3(n5656), .QN(n9464) );
  NAND3X0 U9496 ( .IN1(n9468), .IN2(n9469), .IN3(n9470), .QN(g34461) );
  NAND2X0 U9497 ( .IN1(test_so19), .IN2(n8661), .QN(n9470) );
  NAND3X0 U9498 ( .IN1(n9458), .IN2(n2573), .IN3(n8152), .QN(n9469) );
  NAND2X0 U9499 ( .IN1(n2577), .IN2(n9460), .QN(n9468) );
  INVX0 U9500 ( .INP(n9471), .ZN(n9460) );
  NAND2X0 U9501 ( .IN1(n9472), .IN2(n9473), .QN(g34460) );
  NAND2X0 U9502 ( .IN1(n9474), .IN2(g4639), .QN(n9473) );
  NAND2X0 U9503 ( .IN1(n9475), .IN2(n8521), .QN(n9474) );
  NAND2X0 U9504 ( .IN1(n9476), .IN2(n8226), .QN(n9475) );
  NAND2X0 U9505 ( .IN1(n322), .IN2(test_so3), .QN(n9472) );
  INVX0 U9506 ( .INP(n9477), .ZN(n322) );
  NAND2X0 U9507 ( .IN1(n9478), .IN2(n9479), .QN(g34459) );
  NAND2X0 U9508 ( .IN1(n8627), .IN2(g4643), .QN(n9479) );
  NAND2X0 U9509 ( .IN1(n9480), .IN2(n8521), .QN(n9478) );
  NAND2X0 U9510 ( .IN1(n9481), .IN2(n9482), .QN(n9480) );
  NAND2X0 U9511 ( .IN1(n9483), .IN2(n9484), .QN(n9482) );
  NAND2X0 U9512 ( .IN1(n5653), .IN2(n9485), .QN(n9483) );
  NAND2X0 U9513 ( .IN1(test_so99), .IN2(n9486), .QN(n9485) );
  NAND2X0 U9514 ( .IN1(n9487), .IN2(n9488), .QN(g34458) );
  NAND2X0 U9515 ( .IN1(n9489), .IN2(g4633), .QN(n9488) );
  NAND2X0 U9516 ( .IN1(n9490), .IN2(n9491), .QN(n9489) );
  NAND3X0 U9517 ( .IN1(n8504), .IN2(n8218), .IN3(n9476), .QN(n9491) );
  INVX0 U9518 ( .INP(n9492), .ZN(n9490) );
  NAND2X0 U9519 ( .IN1(test_so99), .IN2(n9493), .QN(n9487) );
  NAND2X0 U9520 ( .IN1(n9494), .IN2(n8521), .QN(n9493) );
  NAND4X0 U9521 ( .IN1(n5844), .IN2(n9476), .IN3(test_so3), .IN4(g4639), .QN(
        n9494) );
  NAND2X0 U9522 ( .IN1(n9495), .IN2(n9496), .QN(g34457) );
  NAND2X0 U9523 ( .IN1(test_so3), .IN2(n9497), .QN(n9496) );
  NAND2X0 U9524 ( .IN1(n9498), .IN2(n8521), .QN(n9497) );
  NAND3X0 U9525 ( .IN1(g4639), .IN2(n8218), .IN3(n9476), .QN(n9498) );
  NAND2X0 U9526 ( .IN1(test_so99), .IN2(n9492), .QN(n9495) );
  NAND2X0 U9527 ( .IN1(n9477), .IN2(n9499), .QN(n9492) );
  NAND3X0 U9528 ( .IN1(n8503), .IN2(n8226), .IN3(n9476), .QN(n9499) );
  INVX0 U9529 ( .INP(n9500), .ZN(n9476) );
  NAND3X0 U9530 ( .IN1(n5382), .IN2(n9501), .IN3(n5727), .QN(n9477) );
  NAND2X0 U9531 ( .IN1(n9502), .IN2(n9503), .QN(g34456) );
  NAND2X0 U9532 ( .IN1(n9504), .IN2(g4608), .QN(n9503) );
  NAND2X0 U9533 ( .IN1(n9505), .IN2(n8521), .QN(n9504) );
  NAND2X0 U9534 ( .IN1(n2590), .IN2(n9506), .QN(n9505) );
  NAND2X0 U9535 ( .IN1(n9507), .IN2(g4616), .QN(n9502) );
  NAND2X0 U9536 ( .IN1(n9508), .IN2(n9509), .QN(g34455) );
  NAND2X0 U9537 ( .IN1(n9510), .IN2(g4322), .QN(n9509) );
  NAND2X0 U9538 ( .IN1(n9511), .IN2(n8521), .QN(n9510) );
  NAND3X0 U9539 ( .IN1(n9512), .IN2(n9481), .IN3(n2594), .QN(n9511) );
  NAND2X0 U9540 ( .IN1(n2595), .IN2(g4332), .QN(n9508) );
  NAND2X0 U9541 ( .IN1(n9513), .IN2(n9514), .QN(g34454) );
  NAND2X0 U9542 ( .IN1(n9515), .IN2(n9507), .QN(n9514) );
  XOR2X1 U9543 ( .IN1(n2590), .IN2(g4608), .Q(n9515) );
  NAND2X0 U9544 ( .IN1(n8627), .IN2(g4601), .QN(n9513) );
  NAND3X0 U9545 ( .IN1(n9516), .IN2(n9517), .IN3(n9518), .QN(g34453) );
  NAND2X0 U9546 ( .IN1(n8627), .IN2(g4593), .QN(n9518) );
  NAND3X0 U9547 ( .IN1(n9507), .IN2(n9519), .IN3(g4601), .QN(n9517) );
  INVX0 U9548 ( .INP(n2598), .ZN(n9519) );
  NAND3X0 U9549 ( .IN1(n2598), .IN2(n9506), .IN3(n5365), .QN(n9516) );
  NAND2X0 U9550 ( .IN1(n9520), .IN2(n9521), .QN(g34452) );
  NAND2X0 U9551 ( .IN1(n9522), .IN2(n9507), .QN(n9521) );
  XOR2X1 U9552 ( .IN1(g4593), .IN2(n2601), .Q(n9522) );
  NAND2X0 U9553 ( .IN1(n8627), .IN2(g4584), .QN(n9520) );
  NAND2X0 U9554 ( .IN1(n9523), .IN2(n9524), .QN(g34451) );
  NAND2X0 U9555 ( .IN1(n9525), .IN2(n9507), .QN(n9524) );
  AND2X1 U9556 ( .IN1(n9506), .IN2(n8508), .Q(n9507) );
  AND2X1 U9557 ( .IN1(n9526), .IN2(n9481), .Q(n9506) );
  NAND2X0 U9558 ( .IN1(n2601), .IN2(g4616), .QN(n9526) );
  NOR2X0 U9559 ( .IN1(n9512), .IN2(n5539), .QN(n2601) );
  XOR2X1 U9560 ( .IN1(n9512), .IN2(n5539), .Q(n9525) );
  NAND2X0 U9561 ( .IN1(n8627), .IN2(g4332), .QN(n9523) );
  NAND3X0 U9562 ( .IN1(n9527), .IN2(n9528), .IN3(n9529), .QN(g34450) );
  NAND2X0 U9563 ( .IN1(n8627), .IN2(g4311), .QN(n9529) );
  NAND3X0 U9564 ( .IN1(n2595), .IN2(n9530), .IN3(g4322), .QN(n9528) );
  INVX0 U9565 ( .INP(n2594), .ZN(n9530) );
  AND2X1 U9566 ( .IN1(n9501), .IN2(n9512), .Q(n2595) );
  NAND3X0 U9567 ( .IN1(g4322), .IN2(g4332), .IN3(n2607), .QN(n9512) );
  NOR2X0 U9568 ( .IN1(n9531), .IN2(n5348), .QN(n2607) );
  NAND3X0 U9569 ( .IN1(n2594), .IN2(n9481), .IN3(n5506), .QN(n9527) );
  NAND3X0 U9570 ( .IN1(n9532), .IN2(n9533), .IN3(n9534), .QN(g34448) );
  NAND2X0 U9571 ( .IN1(n8627), .IN2(g2827), .QN(n9534) );
  NAND3X0 U9572 ( .IN1(n8504), .IN2(g2819), .IN3(n9535), .QN(n9533) );
  NAND3X0 U9573 ( .IN1(n9536), .IN2(n9537), .IN3(n9538), .QN(n9532) );
  NAND2X0 U9574 ( .IN1(n9539), .IN2(g2827), .QN(n9537) );
  NAND3X0 U9575 ( .IN1(n9540), .IN2(n9541), .IN3(n9542), .QN(g34447) );
  NAND2X0 U9576 ( .IN1(n8626), .IN2(g2815), .QN(n9542) );
  NAND3X0 U9577 ( .IN1(n8503), .IN2(g2807), .IN3(n9543), .QN(n9541) );
  NAND3X0 U9578 ( .IN1(n9536), .IN2(n9544), .IN3(n9545), .QN(n9540) );
  NAND2X0 U9579 ( .IN1(n9539), .IN2(g2811), .QN(n9544) );
  NAND3X0 U9580 ( .IN1(n9546), .IN2(n9547), .IN3(n9548), .QN(g34446) );
  NAND2X0 U9581 ( .IN1(n8626), .IN2(g2819), .QN(n9548) );
  NAND3X0 U9582 ( .IN1(n8503), .IN2(g2815), .IN3(n9549), .QN(n9547) );
  NAND3X0 U9583 ( .IN1(n9536), .IN2(n9550), .IN3(n9551), .QN(n9546) );
  NAND2X0 U9584 ( .IN1(test_so37), .IN2(n9539), .QN(n9550) );
  NAND3X0 U9585 ( .IN1(n9552), .IN2(n9553), .IN3(n9554), .QN(g34445) );
  NAND2X0 U9586 ( .IN1(n8626), .IN2(g2807), .QN(n9554) );
  NAND3X0 U9587 ( .IN1(n8503), .IN2(g2803), .IN3(n9555), .QN(n9553) );
  NAND3X0 U9588 ( .IN1(n9536), .IN2(n9556), .IN3(n9557), .QN(n9552) );
  NAND2X0 U9589 ( .IN1(n9539), .IN2(g2799), .QN(n9556) );
  AND2X1 U9590 ( .IN1(n9558), .IN2(n8508), .Q(n9536) );
  NAND2X0 U9591 ( .IN1(n2760), .IN2(n9255), .QN(n9558) );
  NAND3X0 U9592 ( .IN1(n9559), .IN2(n9560), .IN3(n9561), .QN(g34444) );
  NAND2X0 U9593 ( .IN1(n8626), .IN2(g2795), .QN(n9561) );
  NAND3X0 U9594 ( .IN1(n8503), .IN2(g2787), .IN3(n9535), .QN(n9560) );
  NAND3X0 U9595 ( .IN1(n9562), .IN2(n9563), .IN3(n9538), .QN(n9559) );
  INVX0 U9596 ( .INP(n9535), .ZN(n9538) );
  NAND2X0 U9597 ( .IN1(n9564), .IN2(n9565), .QN(n9535) );
  NAND2X0 U9598 ( .IN1(n9539), .IN2(g2795), .QN(n9563) );
  NAND3X0 U9599 ( .IN1(n9566), .IN2(n9567), .IN3(n9568), .QN(g34443) );
  NAND2X0 U9600 ( .IN1(n8626), .IN2(g2783), .QN(n9568) );
  NAND3X0 U9601 ( .IN1(n8503), .IN2(g2775), .IN3(n9543), .QN(n9567) );
  NAND3X0 U9602 ( .IN1(n9562), .IN2(n9569), .IN3(n9545), .QN(n9566) );
  INVX0 U9603 ( .INP(n9543), .ZN(n9545) );
  NAND3X0 U9604 ( .IN1(n7867), .IN2(g2724), .IN3(n9564), .QN(n9543) );
  NAND2X0 U9605 ( .IN1(n9539), .IN2(g2779), .QN(n9569) );
  NAND3X0 U9606 ( .IN1(n9570), .IN2(n9571), .IN3(n9572), .QN(g34442) );
  NAND2X0 U9607 ( .IN1(n8626), .IN2(g2787), .QN(n9572) );
  NAND3X0 U9608 ( .IN1(n8503), .IN2(g2783), .IN3(n9549), .QN(n9571) );
  NAND3X0 U9609 ( .IN1(n9562), .IN2(n9573), .IN3(n9551), .QN(n9570) );
  INVX0 U9610 ( .INP(n9549), .ZN(n9551) );
  NAND2X0 U9611 ( .IN1(n9574), .IN2(n9564), .QN(n9549) );
  NAND2X0 U9612 ( .IN1(n9539), .IN2(g2791), .QN(n9573) );
  NAND3X0 U9613 ( .IN1(n9575), .IN2(n9576), .IN3(n9577), .QN(g34441) );
  NAND2X0 U9614 ( .IN1(n8626), .IN2(g2775), .QN(n9577) );
  NAND3X0 U9615 ( .IN1(n8504), .IN2(g2771), .IN3(n9555), .QN(n9576) );
  NAND3X0 U9616 ( .IN1(n9562), .IN2(n9578), .IN3(n9557), .QN(n9575) );
  INVX0 U9617 ( .INP(n9555), .ZN(n9557) );
  NAND2X0 U9618 ( .IN1(n9564), .IN2(n9579), .QN(n9555) );
  INVX0 U9619 ( .INP(n9580), .ZN(n9564) );
  NAND2X0 U9620 ( .IN1(n9539), .IN2(g2767), .QN(n9578) );
  AND2X1 U9621 ( .IN1(n9581), .IN2(n8509), .Q(n9562) );
  NAND2X0 U9622 ( .IN1(n2760), .IN2(n9265), .QN(n9581) );
  NAND2X0 U9623 ( .IN1(n9582), .IN2(n9583), .QN(g34440) );
  NAND2X0 U9624 ( .IN1(n8625), .IN2(g446), .QN(n9583) );
  NAND2X0 U9625 ( .IN1(n9584), .IN2(n8521), .QN(n9582) );
  NAND2X0 U9626 ( .IN1(n9585), .IN2(n9586), .QN(n9584) );
  NAND2X0 U9627 ( .IN1(n9587), .IN2(g862), .QN(n9586) );
  NAND2X0 U9628 ( .IN1(g896), .IN2(n9588), .QN(n9587) );
  NAND2X0 U9629 ( .IN1(n9589), .IN2(n9590), .QN(n9588) );
  OR3X1 U9630 ( .IN1(n9591), .IN2(n2644), .IN3(g703), .Q(n9589) );
  NAND2X0 U9631 ( .IN1(g890), .IN2(g896), .QN(n9585) );
  NAND3X0 U9632 ( .IN1(n9592), .IN2(n9593), .IN3(n9594), .QN(g34439) );
  NAND2X0 U9633 ( .IN1(n8625), .IN2(g772), .QN(n9594) );
  NAND3X0 U9634 ( .IN1(n2404), .IN2(n9595), .IN3(g776), .QN(n9593) );
  INVX0 U9635 ( .INP(n2554), .ZN(n9595) );
  NAND2X0 U9636 ( .IN1(n2554), .IN2(n5330), .QN(n9592) );
  NAND3X0 U9637 ( .IN1(n9596), .IN2(n9597), .IN3(n9598), .QN(g34438) );
  NAND2X0 U9638 ( .IN1(n8625), .IN2(g604), .QN(n9598) );
  NAND3X0 U9639 ( .IN1(n2421), .IN2(n9599), .IN3(g608), .QN(n9597) );
  INVX0 U9640 ( .INP(n2556), .ZN(n9599) );
  NAND2X0 U9641 ( .IN1(n2556), .IN2(n5475), .QN(n9596) );
  NOR4X0 U9642 ( .IN1(n9600), .IN2(g4064), .IN3(g4057), .IN4(g4125), .QN(
        g34435) );
  AND3X1 U9643 ( .IN1(n5612), .IN2(n9601), .IN3(n7826), .Q(n9600) );
  NAND4X0 U9644 ( .IN1(test_so11), .IN2(n5350), .IN3(n9602), .IN4(g4112), .QN(
        n9601) );
  NAND2X0 U9645 ( .IN1(n2730), .IN2(n9603), .QN(g34425) );
  INVX0 U9646 ( .INP(n8197), .ZN(n9603) );
  NAND2X0 U9647 ( .IN1(n9604), .IN2(n9605), .QN(n8197) );
  NAND2X0 U9648 ( .IN1(n9606), .IN2(g4358), .QN(n9605) );
  NAND2X0 U9649 ( .IN1(n9607), .IN2(n9608), .QN(n9606) );
  NAND2X0 U9650 ( .IN1(test_so81), .IN2(n9609), .QN(n9608) );
  NAND2X0 U9651 ( .IN1(n9610), .IN2(n9611), .QN(n9609) );
  NAND2X0 U9652 ( .IN1(n9612), .IN2(n9292), .QN(n9611) );
  NAND2X0 U9653 ( .IN1(n9613), .IN2(n9289), .QN(n9610) );
  NAND2X0 U9654 ( .IN1(n9614), .IN2(n8208), .QN(n9607) );
  NAND2X0 U9655 ( .IN1(n9615), .IN2(n9616), .QN(n9614) );
  NAND2X0 U9656 ( .IN1(n9617), .IN2(n9292), .QN(n9616) );
  NAND2X0 U9657 ( .IN1(n9618), .IN2(n9289), .QN(n9615) );
  NAND2X0 U9658 ( .IN1(n9619), .IN2(n5348), .QN(n9604) );
  NAND2X0 U9659 ( .IN1(n9620), .IN2(n9621), .QN(n9619) );
  NAND2X0 U9660 ( .IN1(test_so81), .IN2(n9622), .QN(n9621) );
  NAND2X0 U9661 ( .IN1(n9623), .IN2(n9624), .QN(n9622) );
  NAND2X0 U9662 ( .IN1(n9625), .IN2(n9292), .QN(n9624) );
  NAND2X0 U9663 ( .IN1(n9626), .IN2(n9289), .QN(n9623) );
  NAND2X0 U9664 ( .IN1(n9627), .IN2(n8208), .QN(n9620) );
  NAND2X0 U9665 ( .IN1(n9628), .IN2(n9629), .QN(n9627) );
  NAND2X0 U9666 ( .IN1(g31860), .IN2(n9292), .QN(n9629) );
  NAND2X0 U9667 ( .IN1(n8821), .IN2(n9289), .QN(n9628) );
  AND2X1 U9668 ( .IN1(n9630), .IN2(n9631), .Q(n2730) );
  NAND2X0 U9669 ( .IN1(n9632), .IN2(n9633), .QN(n9631) );
  NAND3X0 U9670 ( .IN1(n9634), .IN2(n9188), .IN3(n9630), .QN(g34383) );
  NOR2X0 U9671 ( .IN1(n9635), .IN2(n9636), .QN(n9188) );
  NAND4X0 U9672 ( .IN1(n9637), .IN2(n9638), .IN3(n9639), .IN4(n9640), .QN(
        n9636) );
  NAND3X0 U9673 ( .IN1(n9641), .IN2(g2227), .IN3(n5514), .QN(n9640) );
  NAND2X0 U9674 ( .IN1(n9642), .IN2(n9643), .QN(n9639) );
  NAND2X0 U9675 ( .IN1(n9644), .IN2(n9645), .QN(n9638) );
  NAND2X0 U9676 ( .IN1(g31862), .IN2(n9646), .QN(n9637) );
  NAND4X0 U9677 ( .IN1(n9647), .IN2(n9648), .IN3(n9649), .IN4(n9650), .QN(
        n9635) );
  NAND3X0 U9678 ( .IN1(n9651), .IN2(g2070), .IN3(n5505), .QN(n9650) );
  NAND3X0 U9679 ( .IN1(n9652), .IN2(g1802), .IN3(n5504), .QN(n9649) );
  NAND3X0 U9680 ( .IN1(n9653), .IN2(g2629), .IN3(n5524), .QN(n9648) );
  NAND3X0 U9681 ( .IN1(n9654), .IN2(g2361), .IN3(n5513), .QN(n9647) );
  NAND4X0 U9682 ( .IN1(n9655), .IN2(n9656), .IN3(n9657), .IN4(n9658), .QN(
        n9634) );
  NOR4X0 U9683 ( .IN1(n9659), .IN2(n9651), .IN3(n9641), .IN4(n9654), .QN(n9658) );
  NAND2X0 U9684 ( .IN1(n9660), .IN2(n9661), .QN(g34269) );
  NAND2X0 U9685 ( .IN1(n8625), .IN2(g4961), .QN(n9661) );
  NAND3X0 U9686 ( .IN1(n9662), .IN2(n9663), .IN3(n9664), .QN(n9660) );
  NAND3X0 U9687 ( .IN1(n5614), .IN2(n9665), .IN3(n9666), .QN(n9663) );
  NAND3X0 U9688 ( .IN1(n5770), .IN2(n9667), .IN3(n9668), .QN(n9662) );
  NAND2X0 U9689 ( .IN1(n9669), .IN2(n9670), .QN(g34268) );
  NAND2X0 U9690 ( .IN1(n8625), .IN2(g4950), .QN(n9670) );
  NAND3X0 U9691 ( .IN1(n9671), .IN2(n9672), .IN3(n9664), .QN(n9669) );
  NAND3X0 U9692 ( .IN1(n5875), .IN2(n9665), .IN3(n9673), .QN(n9672) );
  NAND3X0 U9693 ( .IN1(n5772), .IN2(n9667), .IN3(n9674), .QN(n9671) );
  NAND2X0 U9694 ( .IN1(n9675), .IN2(n9676), .QN(g34267) );
  NAND2X0 U9695 ( .IN1(n9677), .IN2(n8521), .QN(n9676) );
  NAND2X0 U9696 ( .IN1(n9667), .IN2(n9678), .QN(n9677) );
  NAND3X0 U9697 ( .IN1(n9665), .IN2(g4933), .IN3(n9679), .QN(n9678) );
  NAND2X0 U9698 ( .IN1(n9680), .IN2(g4939), .QN(n9675) );
  NAND2X0 U9699 ( .IN1(n9681), .IN2(n8521), .QN(n9680) );
  NAND2X0 U9700 ( .IN1(n9682), .IN2(n9665), .QN(n9681) );
  NAND2X0 U9701 ( .IN1(n9683), .IN2(n9684), .QN(g34266) );
  NAND2X0 U9702 ( .IN1(n8625), .IN2(g4894), .QN(n9684) );
  NAND3X0 U9703 ( .IN1(n9685), .IN2(n9686), .IN3(n9664), .QN(n9683) );
  AND2X1 U9704 ( .IN1(n9687), .IN2(n8508), .Q(n9664) );
  NAND2X0 U9705 ( .IN1(n9688), .IN2(n9667), .QN(n9687) );
  NAND3X0 U9706 ( .IN1(n5863), .IN2(n9665), .IN3(n9689), .QN(n9686) );
  NAND3X0 U9707 ( .IN1(n5774), .IN2(n9667), .IN3(n9288), .QN(n9685) );
  NAND2X0 U9708 ( .IN1(n9688), .IN2(g71), .QN(n9667) );
  INVX0 U9709 ( .INP(n9665), .ZN(n9688) );
  NAND3X0 U9710 ( .IN1(n2668), .IN2(DFF_672_n1), .IN3(n5637), .QN(n9665) );
  NOR4X0 U9711 ( .IN1(g4864), .IN2(g4871), .IN3(g4836), .IN4(n9453), .QN(
        g34265) );
  NAND2X0 U9712 ( .IN1(n9440), .IN2(n8520), .QN(n9453) );
  NOR2X0 U9713 ( .IN1(n9690), .IN2(n9290), .QN(n9440) );
  NAND2X0 U9714 ( .IN1(n9691), .IN2(n9692), .QN(g34264) );
  NAND2X0 U9715 ( .IN1(n8625), .IN2(g4771), .QN(n9692) );
  NAND3X0 U9716 ( .IN1(n9693), .IN2(n9694), .IN3(n9695), .QN(n9691) );
  NAND3X0 U9717 ( .IN1(n5613), .IN2(n9696), .IN3(n9697), .QN(n9694) );
  NAND3X0 U9718 ( .IN1(n5769), .IN2(n9698), .IN3(n9699), .QN(n9693) );
  NAND2X0 U9719 ( .IN1(n9700), .IN2(n9701), .QN(g34263) );
  NAND2X0 U9720 ( .IN1(n8627), .IN2(g4760), .QN(n9701) );
  NAND3X0 U9721 ( .IN1(n9702), .IN2(n9703), .IN3(n9695), .QN(n9700) );
  NAND3X0 U9722 ( .IN1(n5877), .IN2(n9696), .IN3(n9704), .QN(n9703) );
  NAND3X0 U9723 ( .IN1(n5775), .IN2(n9698), .IN3(n9705), .QN(n9702) );
  NAND2X0 U9724 ( .IN1(n9706), .IN2(n9707), .QN(g34262) );
  NAND2X0 U9725 ( .IN1(n9708), .IN2(n8520), .QN(n9707) );
  NAND2X0 U9726 ( .IN1(n9698), .IN2(n9709), .QN(n9708) );
  NAND3X0 U9727 ( .IN1(n9696), .IN2(g4743), .IN3(n9710), .QN(n9709) );
  NAND2X0 U9728 ( .IN1(test_so18), .IN2(n9711), .QN(n9706) );
  NAND2X0 U9729 ( .IN1(n9712), .IN2(n8520), .QN(n9711) );
  NAND2X0 U9730 ( .IN1(n9713), .IN2(n9696), .QN(n9712) );
  NAND2X0 U9731 ( .IN1(n9714), .IN2(n9715), .QN(g34261) );
  NAND2X0 U9732 ( .IN1(n8625), .IN2(g4704), .QN(n9715) );
  NAND3X0 U9733 ( .IN1(n9716), .IN2(n9717), .IN3(n9695), .QN(n9714) );
  AND2X1 U9734 ( .IN1(n9718), .IN2(n8508), .Q(n9695) );
  NAND2X0 U9735 ( .IN1(n9719), .IN2(n9698), .QN(n9718) );
  NAND3X0 U9736 ( .IN1(n5862), .IN2(n9696), .IN3(n9720), .QN(n9717) );
  NAND3X0 U9737 ( .IN1(n5771), .IN2(n9698), .IN3(n9291), .QN(n9716) );
  NAND2X0 U9738 ( .IN1(n9719), .IN2(g101), .QN(n9698) );
  INVX0 U9739 ( .INP(n9696), .ZN(n9719) );
  NAND3X0 U9740 ( .IN1(n2668), .IN2(DFF_178_n1), .IN3(n5636), .QN(n9696) );
  NOR4X0 U9741 ( .IN1(g4674), .IN2(g4646), .IN3(g4681), .IN4(n9471), .QN(
        g34260) );
  NAND2X0 U9742 ( .IN1(n9458), .IN2(n8520), .QN(n9471) );
  NOR2X0 U9743 ( .IN1(n9293), .IN2(n9721), .QN(n9458) );
  NOR2X0 U9744 ( .IN1(n5844), .IN2(n9722), .QN(g34259) );
  NOR2X0 U9745 ( .IN1(n8545), .IN2(n9723), .QN(n9722) );
  NOR2X0 U9746 ( .IN1(n9724), .IN2(n9500), .QN(n9723) );
  NAND2X0 U9747 ( .IN1(n5382), .IN2(n9481), .QN(n9500) );
  NAND3X0 U9748 ( .IN1(n9725), .IN2(n9726), .IN3(n9727), .QN(g34258) );
  NAND2X0 U9749 ( .IN1(test_so81), .IN2(n8547), .QN(n9727) );
  NAND3X0 U9750 ( .IN1(n9501), .IN2(n9531), .IN3(g4358), .QN(n9726) );
  NAND3X0 U9751 ( .IN1(n9728), .IN2(n9481), .IN3(n5348), .QN(n9725) );
  INVX0 U9752 ( .INP(n9531), .ZN(n9728) );
  NAND2X0 U9753 ( .IN1(n9729), .IN2(test_so81), .QN(n9531) );
  NAND3X0 U9754 ( .IN1(n9730), .IN2(n9731), .IN3(n9732), .QN(g34257) );
  NAND2X0 U9755 ( .IN1(n8626), .IN2(g4340), .QN(n9732) );
  NAND3X0 U9756 ( .IN1(n9501), .IN2(test_so81), .IN3(n9484), .QN(n9731) );
  AND2X1 U9757 ( .IN1(n9481), .IN2(n8508), .Q(n9501) );
  NAND3X0 U9758 ( .IN1(n9481), .IN2(n8208), .IN3(n9729), .QN(n9730) );
  INVX0 U9759 ( .INP(n9484), .ZN(n9729) );
  NAND3X0 U9760 ( .IN1(n9486), .IN2(g4340), .IN3(test_so99), .QN(n9484) );
  INVX0 U9761 ( .INP(n9724), .ZN(n9486) );
  NAND2X0 U9762 ( .IN1(n9281), .IN2(n9733), .QN(n9481) );
  NAND2X0 U9763 ( .IN1(n9172), .IN2(n1430), .QN(n9733) );
  NAND2X0 U9764 ( .IN1(n9734), .IN2(n9735), .QN(g34256) );
  OR2X1 U9765 ( .IN1(n8477), .IN2(n7999), .Q(n9735) );
  NAND2X0 U9766 ( .IN1(n9736), .IN2(n8520), .QN(n9734) );
  NAND3X0 U9767 ( .IN1(n9737), .IN2(n9738), .IN3(n5765), .QN(n9736) );
  NAND2X0 U9768 ( .IN1(n5671), .IN2(g4473), .QN(n9737) );
  NAND4X0 U9769 ( .IN1(n5671), .IN2(n9739), .IN3(n9738), .IN4(n8506), .QN(
        g34255) );
  NAND2X0 U9770 ( .IN1(test_so38), .IN2(g4473), .QN(n9739) );
  NAND2X0 U9771 ( .IN1(n9740), .IN2(n9741), .QN(g34254) );
  NAND2X0 U9772 ( .IN1(n9742), .IN2(g4473), .QN(n9741) );
  NAND4X0 U9773 ( .IN1(n8508), .IN2(g4643), .IN3(g4462), .IN4(n8222), .QN(
        n9742) );
  OR2X1 U9774 ( .IN1(n9738), .IN2(n8545), .Q(n9740) );
  NOR2X0 U9775 ( .IN1(n8569), .IN2(n9743), .QN(g34253) );
  AND3X1 U9776 ( .IN1(test_so38), .IN2(g4462), .IN3(n9738), .Q(n9743) );
  NAND3X0 U9777 ( .IN1(n9744), .IN2(g26960), .IN3(n5849), .QN(n9738) );
  NAND2X0 U9778 ( .IN1(n9172), .IN2(n9745), .QN(n9744) );
  NAND2X0 U9779 ( .IN1(n5846), .IN2(n2668), .QN(n9745) );
  NAND3X0 U9780 ( .IN1(n9746), .IN2(n9747), .IN3(n9748), .QN(g34252) );
  NAND2X0 U9781 ( .IN1(n8616), .IN2(g767), .QN(n9748) );
  NAND3X0 U9782 ( .IN1(n2404), .IN2(n9749), .IN3(g772), .QN(n9747) );
  INVX0 U9783 ( .INP(n2647), .ZN(n9749) );
  NAND2X0 U9784 ( .IN1(n2647), .IN2(n5334), .QN(n9746) );
  NAND3X0 U9785 ( .IN1(n9750), .IN2(n9751), .IN3(n9752), .QN(g34251) );
  NAND2X0 U9786 ( .IN1(n8617), .IN2(g599), .QN(n9752) );
  NAND3X0 U9787 ( .IN1(n2421), .IN2(n9753), .IN3(g604), .QN(n9751) );
  INVX0 U9788 ( .INP(n2649), .ZN(n9753) );
  NAND2X0 U9789 ( .IN1(n2649), .IN2(n5473), .QN(n9750) );
  NAND3X0 U9790 ( .IN1(n9754), .IN2(n9755), .IN3(n9756), .QN(g34250) );
  NAND2X0 U9791 ( .IN1(n8649), .IN2(g298), .QN(n9756) );
  NAND3X0 U9792 ( .IN1(n8194), .IN2(n9757), .IN3(g142), .QN(n9755) );
  INVX0 U9793 ( .INP(n2707), .ZN(n9757) );
  NAND2X0 U9794 ( .IN1(n5724), .IN2(n2707), .QN(n9754) );
  NAND3X0 U9795 ( .IN1(n9758), .IN2(n9759), .IN3(n9760), .QN(g34249) );
  OR2X1 U9796 ( .IN1(n8477), .IN2(n5678), .Q(n9760) );
  OR3X1 U9797 ( .IN1(n9761), .IN2(n2710), .IN3(n5843), .Q(n9759) );
  NAND2X0 U9798 ( .IN1(n2710), .IN2(n5843), .QN(n9758) );
  NAND3X0 U9799 ( .IN1(n9762), .IN2(n8905), .IN3(n9630), .QN(g34201) );
  NOR2X0 U9800 ( .IN1(n9763), .IN2(n9764), .QN(n8905) );
  NAND4X0 U9801 ( .IN1(n9765), .IN2(n9766), .IN3(n9767), .IN4(n9768), .QN(
        n9764) );
  NAND3X0 U9802 ( .IN1(n9769), .IN2(g2051), .IN3(n5507), .QN(n9768) );
  NAND3X0 U9803 ( .IN1(n9770), .IN2(g1917), .IN3(n5510), .QN(n9767) );
  NAND3X0 U9804 ( .IN1(n3005), .IN2(g1783), .IN3(n5359), .QN(n9766) );
  NAND2X0 U9805 ( .IN1(g31863), .IN2(n9771), .QN(n9765) );
  NAND4X0 U9806 ( .IN1(n9772), .IN2(n9773), .IN3(n9774), .IN4(n9775), .QN(
        n9763) );
  NAND3X0 U9807 ( .IN1(n9776), .IN2(g2610), .IN3(n5508), .QN(n9775) );
  NAND3X0 U9808 ( .IN1(n9777), .IN2(g2476), .IN3(n5509), .QN(n9774) );
  NAND3X0 U9809 ( .IN1(test_so21), .IN2(n9778), .IN3(n5511), .QN(n9773) );
  NAND3X0 U9810 ( .IN1(n9779), .IN2(g2208), .IN3(n5512), .QN(n9772) );
  NAND4X0 U9811 ( .IN1(n3588), .IN2(n3606), .IN3(n9780), .IN4(n9781), .QN(
        n9762) );
  NOR4X0 U9812 ( .IN1(n9779), .IN2(n9778), .IN3(n9777), .IN4(n9776), .QN(n9781) );
  NOR2X0 U9813 ( .IN1(n3005), .IN2(n9771), .QN(n9780) );
  NAND2X0 U9814 ( .IN1(n9782), .IN2(n9783), .QN(g34041) );
  NAND2X0 U9815 ( .IN1(n9784), .IN2(n9785), .QN(n9783) );
  XOR2X1 U9816 ( .IN1(n9786), .IN2(n5367), .Q(n9784) );
  OR2X1 U9817 ( .IN1(n8476), .IN2(n5637), .Q(n9782) );
  NAND3X0 U9818 ( .IN1(n9787), .IN2(n9788), .IN3(n9789), .QN(g34040) );
  NAND2X0 U9819 ( .IN1(n8614), .IN2(g4975), .QN(n9789) );
  NAND2X0 U9820 ( .IN1(n9790), .IN2(n9791), .QN(n9788) );
  NAND2X0 U9821 ( .IN1(n9792), .IN2(n9793), .QN(n9790) );
  NAND2X0 U9822 ( .IN1(n9794), .IN2(n8883), .QN(n9793) );
  NAND2X0 U9823 ( .IN1(n8882), .IN2(n8520), .QN(n9792) );
  NAND2X0 U9824 ( .IN1(n9785), .IN2(g4899), .QN(n9787) );
  NAND2X0 U9826 ( .IN1(n9795), .IN2(n9796), .QN(g34039) );
  NAND2X0 U9827 ( .IN1(test_so58), .IN2(n9797), .QN(n9796) );
  NAND2X0 U9828 ( .IN1(n9798), .IN2(n8520), .QN(n9797) );
  NAND2X0 U9829 ( .IN1(n9799), .IN2(n9800), .QN(n9798) );
  NAND2X0 U9830 ( .IN1(n9785), .IN2(g4966), .QN(n9795) );
  NAND3X0 U9831 ( .IN1(n9801), .IN2(n9802), .IN3(n9803), .QN(g34038) );
  NAND2X0 U9832 ( .IN1(n8615), .IN2(g4983), .QN(n9803) );
  NAND3X0 U9833 ( .IN1(n9799), .IN2(n9800), .IN3(n8214), .QN(n9802) );
  INVX0 U9834 ( .INP(n9804), .ZN(n9800) );
  NAND3X0 U9835 ( .IN1(n9785), .IN2(n9804), .IN3(test_so58), .QN(n9801) );
  NAND3X0 U9836 ( .IN1(n9805), .IN2(n9806), .IN3(n9807), .QN(g34037) );
  NAND2X0 U9837 ( .IN1(n8631), .IN2(g4966), .QN(n9807) );
  NAND2X0 U9838 ( .IN1(n9785), .IN2(g4975), .QN(n9806) );
  AND2X1 U9839 ( .IN1(n9799), .IN2(n8508), .Q(n9785) );
  NOR2X0 U9840 ( .IN1(n9794), .IN2(n9690), .QN(n9799) );
  INVX0 U9841 ( .INP(n9791), .ZN(n9690) );
  NAND3X0 U9842 ( .IN1(n9794), .IN2(n9791), .IN3(n5360), .QN(n9805) );
  NOR2X0 U9843 ( .IN1(n9804), .IN2(n5706), .QN(n9794) );
  NAND2X0 U9844 ( .IN1(n9290), .IN2(g4983), .QN(n9804) );
  INVX0 U9845 ( .INP(n9786), .ZN(n9290) );
  NAND4X0 U9846 ( .IN1(g4878), .IN2(g4859), .IN3(g4843), .IN4(g4849), .QN(
        n9786) );
  NOR2X0 U9847 ( .IN1(n5443), .IN2(n9808), .QN(g34036) );
  NOR2X0 U9848 ( .IN1(n5318), .IN2(n9808), .QN(g34035) );
  NOR2X0 U9849 ( .IN1(n5713), .IN2(n9808), .QN(g34034) );
  NOR2X0 U9850 ( .IN1(n9791), .IN2(n8551), .QN(n9808) );
  NAND3X0 U9851 ( .IN1(n2760), .IN2(g63), .IN3(n9289), .QN(n9791) );
  NAND2X0 U9852 ( .IN1(n9809), .IN2(n9810), .QN(g34033) );
  NAND2X0 U9853 ( .IN1(n9811), .IN2(n9812), .QN(n9810) );
  XOR2X1 U9854 ( .IN1(n9813), .IN2(n5368), .Q(n9811) );
  OR2X1 U9855 ( .IN1(n8476), .IN2(n5636), .Q(n9809) );
  NAND3X0 U9856 ( .IN1(n9814), .IN2(n9815), .IN3(n9816), .QN(g34032) );
  NAND2X0 U9857 ( .IN1(n8632), .IN2(g4785), .QN(n9816) );
  NAND2X0 U9858 ( .IN1(n9817), .IN2(n9818), .QN(n9815) );
  NAND2X0 U9859 ( .IN1(n9819), .IN2(n9820), .QN(n9817) );
  NAND2X0 U9860 ( .IN1(n9821), .IN2(n8853), .QN(n9820) );
  NAND2X0 U9861 ( .IN1(n8852), .IN2(n8520), .QN(n9819) );
  NAND2X0 U9862 ( .IN1(n9812), .IN2(g4709), .QN(n9814) );
  NAND2X0 U9863 ( .IN1(n9822), .IN2(n9823), .QN(g34031) );
  NAND2X0 U9864 ( .IN1(test_so29), .IN2(n9824), .QN(n9823) );
  NAND2X0 U9865 ( .IN1(n9825), .IN2(n8520), .QN(n9824) );
  NAND2X0 U9866 ( .IN1(n9826), .IN2(n9827), .QN(n9825) );
  NAND2X0 U9867 ( .IN1(n9812), .IN2(g4776), .QN(n9822) );
  NAND3X0 U9868 ( .IN1(n9828), .IN2(n9829), .IN3(n9830), .QN(g34030) );
  NAND2X0 U9869 ( .IN1(n8634), .IN2(g4793), .QN(n9830) );
  NAND3X0 U9870 ( .IN1(n9826), .IN2(n9827), .IN3(n8215), .QN(n9829) );
  INVX0 U9871 ( .INP(n9831), .ZN(n9827) );
  NAND3X0 U9872 ( .IN1(n9812), .IN2(n9831), .IN3(test_so29), .QN(n9828) );
  NAND3X0 U9873 ( .IN1(n9832), .IN2(n9833), .IN3(n9834), .QN(g34029) );
  NAND2X0 U9874 ( .IN1(n8633), .IN2(g4776), .QN(n9834) );
  NAND2X0 U9875 ( .IN1(n9812), .IN2(g4785), .QN(n9833) );
  AND2X1 U9876 ( .IN1(n9826), .IN2(n8508), .Q(n9812) );
  NOR2X0 U9877 ( .IN1(n9821), .IN2(n9721), .QN(n9826) );
  INVX0 U9878 ( .INP(n9818), .ZN(n9721) );
  NAND3X0 U9879 ( .IN1(n9821), .IN2(n9818), .IN3(n5361), .QN(n9832) );
  NOR2X0 U9880 ( .IN1(n9831), .IN2(n5707), .QN(n9821) );
  NAND2X0 U9881 ( .IN1(n9293), .IN2(g4793), .QN(n9831) );
  INVX0 U9882 ( .INP(n9813), .ZN(n9293) );
  NAND4X0 U9883 ( .IN1(test_so19), .IN2(g4688), .IN3(g4669), .IN4(g4659), .QN(
        n9813) );
  NOR2X0 U9884 ( .IN1(n5440), .IN2(n2774), .QN(g34027) );
  NOR2X0 U9885 ( .IN1(n5712), .IN2(n2774), .QN(g34026) );
  NOR2X0 U9887 ( .IN1(n9818), .IN2(n8548), .QN(n2774) );
  NAND3X0 U9888 ( .IN1(n2760), .IN2(g63), .IN3(n9292), .QN(n9818) );
  NAND4X0 U9889 ( .IN1(n9835), .IN2(n9836), .IN3(n9837), .IN4(n9838), .QN(
        g34024) );
  NAND2X0 U9890 ( .IN1(n8630), .IN2(g4492), .QN(n9838) );
  NAND2X0 U9891 ( .IN1(n9839), .IN2(n8520), .QN(n9837) );
  NAND2X0 U9892 ( .IN1(n9840), .IN2(n9841), .QN(n9839) );
  NAND2X0 U9893 ( .IN1(n9842), .IN2(g4512), .QN(n9841) );
  NAND2X0 U9894 ( .IN1(n9843), .IN2(n9172), .QN(n9840) );
  NAND4X0 U9895 ( .IN1(n9844), .IN2(n9845), .IN3(n9835), .IN4(n9836), .QN(
        g34023) );
  NAND3X0 U9896 ( .IN1(n8503), .IN2(g2988), .IN3(n9172), .QN(n9835) );
  NAND3X0 U9897 ( .IN1(n8503), .IN2(g4552), .IN3(n9842), .QN(n9845) );
  NAND2X0 U9898 ( .IN1(n9846), .IN2(n9325), .QN(n9844) );
  NAND2X0 U9899 ( .IN1(n9847), .IN2(n8520), .QN(n9846) );
  NAND4X0 U9900 ( .IN1(n9172), .IN2(g4555), .IN3(g4558), .IN4(g4561), .QN(
        n9847) );
  NAND4X0 U9901 ( .IN1(n9848), .IN2(n8807), .IN3(n9849), .IN4(n9850), .QN(
        g34022) );
  OR3X1 U9902 ( .IN1(n9851), .IN2(n7689), .IN3(n8537), .Q(n9850) );
  NAND2X0 U9903 ( .IN1(n8629), .IN2(g2759), .QN(n9849) );
  NAND2X0 U9904 ( .IN1(n9851), .IN2(n7689), .QN(n9848) );
  NOR2X0 U9905 ( .IN1(n9852), .IN2(n7684), .QN(n9851) );
  NAND3X0 U9906 ( .IN1(n9853), .IN2(n9854), .IN3(n9855), .QN(g34021) );
  NAND2X0 U9907 ( .IN1(n8624), .IN2(g2648), .QN(n9855) );
  NAND2X0 U9908 ( .IN1(n9856), .IN2(n9857), .QN(n9854) );
  NAND2X0 U9909 ( .IN1(n9858), .IN2(g2567), .QN(n9853) );
  NAND2X0 U9910 ( .IN1(n9859), .IN2(n9860), .QN(g34020) );
  NAND2X0 U9911 ( .IN1(n9861), .IN2(g2629), .QN(n9860) );
  NAND2X0 U9912 ( .IN1(n9862), .IN2(n8520), .QN(n9861) );
  NAND2X0 U9913 ( .IN1(n9863), .IN2(g2643), .QN(n9862) );
  NAND2X0 U9914 ( .IN1(n9864), .IN2(n8520), .QN(n9859) );
  NAND2X0 U9915 ( .IN1(n9865), .IN2(n9866), .QN(n9864) );
  NAND2X0 U9916 ( .IN1(n9867), .IN2(n9868), .QN(n9866) );
  NAND2X0 U9917 ( .IN1(n9869), .IN2(n9870), .QN(n9868) );
  NAND2X0 U9918 ( .IN1(n7785), .IN2(n9871), .QN(n9870) );
  NAND2X0 U9919 ( .IN1(n9872), .IN2(g2643), .QN(n9865) );
  NAND2X0 U9920 ( .IN1(n9871), .IN2(n9873), .QN(n9872) );
  NAND2X0 U9921 ( .IN1(n9863), .IN2(g2555), .QN(n9873) );
  INVX0 U9922 ( .INP(n9867), .ZN(n9863) );
  NAND2X0 U9923 ( .IN1(n9874), .IN2(n9875), .QN(n9867) );
  NAND2X0 U9924 ( .IN1(n5755), .IN2(n9876), .QN(n9875) );
  NAND2X0 U9925 ( .IN1(n9877), .IN2(n9878), .QN(n9874) );
  NAND3X0 U9926 ( .IN1(n9879), .IN2(n9880), .IN3(n9881), .QN(g34019) );
  NAND2X0 U9928 ( .IN1(n9882), .IN2(n9856), .QN(n9881) );
  OR3X1 U9929 ( .IN1(n9882), .IN2(n5800), .IN3(n8537), .Q(n9880) );
  NOR2X0 U9930 ( .IN1(n9883), .IN2(n5521), .QN(n9882) );
  NAND2X0 U9931 ( .IN1(n8624), .IN2(g2571), .QN(n9879) );
  NAND3X0 U9932 ( .IN1(n9884), .IN2(n9885), .IN3(n9886), .QN(g34018) );
  NAND2X0 U9933 ( .IN1(n9887), .IN2(n9856), .QN(n9886) );
  INVX0 U9934 ( .INP(n9888), .ZN(n9887) );
  NAND3X0 U9935 ( .IN1(test_so61), .IN2(n9888), .IN3(n8497), .QN(n9885) );
  NAND2X0 U9936 ( .IN1(n9889), .IN2(n5351), .QN(n9888) );
  NAND2X0 U9937 ( .IN1(n8624), .IN2(g2583), .QN(n9884) );
  NAND3X0 U9938 ( .IN1(n9890), .IN2(n9891), .IN3(n9892), .QN(g34017) );
  NAND2X0 U9939 ( .IN1(n9893), .IN2(n9856), .QN(n9892) );
  INVX0 U9940 ( .INP(n9894), .ZN(n9893) );
  NAND3X0 U9941 ( .IN1(test_so66), .IN2(n9894), .IN3(n8497), .QN(n9891) );
  NAND3X0 U9942 ( .IN1(g2555), .IN2(g2629), .IN3(n9871), .QN(n9894) );
  NAND2X0 U9943 ( .IN1(test_so61), .IN2(n8566), .QN(n9890) );
  NAND3X0 U9944 ( .IN1(n9895), .IN2(n9896), .IN3(n9897), .QN(g34016) );
  NAND2X0 U9945 ( .IN1(n9898), .IN2(n9856), .QN(n9897) );
  INVX0 U9946 ( .INP(n9899), .ZN(n9898) );
  NAND3X0 U9947 ( .IN1(n9899), .IN2(g2571), .IN3(n8497), .QN(n9896) );
  NAND2X0 U9948 ( .IN1(n9889), .IN2(n5521), .QN(n9899) );
  NAND2X0 U9949 ( .IN1(n8624), .IN2(g2563), .QN(n9895) );
  NAND3X0 U9950 ( .IN1(n9900), .IN2(n9901), .IN3(n9902), .QN(g34015) );
  NAND2X0 U9951 ( .IN1(n9903), .IN2(n9856), .QN(n9902) );
  AND3X1 U9952 ( .IN1(n9904), .IN2(n9905), .IN3(n8528), .Q(n9856) );
  NAND2X0 U9954 ( .IN1(n9876), .IN2(g1585), .QN(n9905) );
  OR2X1 U9955 ( .IN1(n9877), .IN2(n9876), .Q(n9904) );
  INVX0 U9956 ( .INP(n9878), .ZN(n9876) );
  NAND2X0 U9959 ( .IN1(n9906), .IN2(n9907), .QN(n9877) );
  OR3X1 U9960 ( .IN1(n9903), .IN2(n5816), .IN3(n8530), .Q(n9901) );
  NOR2X0 U9961 ( .IN1(n9883), .IN2(n5351), .QN(n9903) );
  NAND2X0 U9962 ( .IN1(n8624), .IN2(g2567), .QN(n9900) );
  NAND3X0 U9963 ( .IN1(n9908), .IN2(n9909), .IN3(n9910), .QN(g34014) );
  NAND2X0 U9964 ( .IN1(n8624), .IN2(g2514), .QN(n9910) );
  NAND2X0 U9965 ( .IN1(n9911), .IN2(n9912), .QN(n9909) );
  NAND2X0 U9966 ( .IN1(n9913), .IN2(g2433), .QN(n9908) );
  NAND2X0 U9967 ( .IN1(n9914), .IN2(n9915), .QN(g34013) );
  NAND2X0 U9969 ( .IN1(n9916), .IN2(g2495), .QN(n9915) );
  NAND2X0 U9970 ( .IN1(n9917), .IN2(n8520), .QN(n9916) );
  NAND2X0 U9971 ( .IN1(n9918), .IN2(g2509), .QN(n9917) );
  NAND2X0 U9973 ( .IN1(n9919), .IN2(n8520), .QN(n9914) );
  NAND2X0 U9974 ( .IN1(n9920), .IN2(n9921), .QN(n9919) );
  NAND2X0 U9975 ( .IN1(n9922), .IN2(n9923), .QN(n9921) );
  NAND2X0 U9976 ( .IN1(n9924), .IN2(n9925), .QN(n9923) );
  NAND2X0 U9977 ( .IN1(n7784), .IN2(n9926), .QN(n9925) );
  NAND2X0 U9978 ( .IN1(n9927), .IN2(g2509), .QN(n9920) );
  NAND2X0 U9979 ( .IN1(n9926), .IN2(n9928), .QN(n9927) );
  NAND2X0 U9980 ( .IN1(test_so79), .IN2(n9918), .QN(n9928) );
  INVX0 U9981 ( .INP(n9922), .ZN(n9918) );
  NAND2X0 U9982 ( .IN1(n9929), .IN2(n9930), .QN(n9922) );
  NAND2X0 U9983 ( .IN1(n9931), .IN2(g1589), .QN(n9930) );
  NAND2X0 U9984 ( .IN1(n9932), .IN2(n9933), .QN(n9929) );
  NAND3X0 U9985 ( .IN1(n9934), .IN2(n9935), .IN3(n9936), .QN(g34012) );
  NAND2X0 U9986 ( .IN1(n9937), .IN2(n9911), .QN(n9936) );
  INVX0 U9987 ( .INP(n9938), .ZN(n9937) );
  NAND3X0 U9988 ( .IN1(n9938), .IN2(g2449), .IN3(n8498), .QN(n9935) );
  NAND2X0 U9989 ( .IN1(n9644), .IN2(n9926), .QN(n9938) );
  NAND2X0 U9990 ( .IN1(n8624), .IN2(g2437), .QN(n9934) );
  NAND3X0 U9991 ( .IN1(n9939), .IN2(n9940), .IN3(n9941), .QN(g34011) );
  NAND2X0 U9993 ( .IN1(n9942), .IN2(n9911), .QN(n9941) );
  INVX0 U9994 ( .INP(n9943), .ZN(n9942) );
  NAND3X0 U9995 ( .IN1(n9943), .IN2(n9274), .IN3(n8498), .QN(n9940) );
  NAND2X0 U9996 ( .IN1(n9944), .IN2(n8204), .QN(n9943) );
  NAND2X0 U9997 ( .IN1(n8623), .IN2(g2449), .QN(n9939) );
  NAND3X0 U9998 ( .IN1(n9945), .IN2(n9946), .IN3(n9947), .QN(g34010) );
  NAND2X0 U9999 ( .IN1(n9948), .IN2(n9911), .QN(n9947) );
  INVX0 U10000 ( .INP(n9949), .ZN(n9948) );
  NAND3X0 U10001 ( .IN1(n9949), .IN2(g2441), .IN3(n8498), .QN(n9946) );
  NAND2X0 U10002 ( .IN1(n9950), .IN2(g2495), .QN(n9949) );
  NAND2X0 U10003 ( .IN1(n8623), .IN2(n9274), .QN(n9945) );
  NAND3X0 U10004 ( .IN1(n9951), .IN2(n9952), .IN3(n9953), .QN(g34009) );
  NAND2X0 U10005 ( .IN1(n9954), .IN2(n9911), .QN(n9953) );
  INVX0 U10006 ( .INP(n9955), .ZN(n9954) );
  NAND3X0 U10007 ( .IN1(n9955), .IN2(g2437), .IN3(n8498), .QN(n9952) );
  NAND2X0 U10008 ( .IN1(n9944), .IN2(n5522), .QN(n9955) );
  NAND2X0 U10009 ( .IN1(n8623), .IN2(g2429), .QN(n9951) );
  NAND3X0 U10010 ( .IN1(n9956), .IN2(n9957), .IN3(n9958), .QN(g34008) );
  NAND2X0 U10011 ( .IN1(n9959), .IN2(n9911), .QN(n9958) );
  AND3X1 U10012 ( .IN1(n9960), .IN2(n9961), .IN3(n8528), .Q(n9911) );
  OR2X1 U10013 ( .IN1(n9932), .IN2(n9931), .Q(n9961) );
  NAND2X0 U10014 ( .IN1(n9906), .IN2(n9962), .QN(n9932) );
  NAND2X0 U10015 ( .IN1(n5757), .IN2(n9931), .QN(n9960) );
  INVX0 U10016 ( .INP(n9933), .ZN(n9931) );
  INVX0 U10017 ( .INP(n9963), .ZN(n9959) );
  NAND3X0 U10018 ( .IN1(n9963), .IN2(g2429), .IN3(n8498), .QN(n9957) );
  NAND2X0 U10019 ( .IN1(n9950), .IN2(n5523), .QN(n9963) );
  NAND2X0 U10020 ( .IN1(n8623), .IN2(g2433), .QN(n9956) );
  NAND3X0 U10021 ( .IN1(n9964), .IN2(n9965), .IN3(n9966), .QN(g34007) );
  NAND2X0 U10022 ( .IN1(n8623), .IN2(g2380), .QN(n9966) );
  NAND2X0 U10023 ( .IN1(n9967), .IN2(n9968), .QN(n9965) );
  NAND2X0 U10024 ( .IN1(n9969), .IN2(g2299), .QN(n9964) );
  NAND2X0 U10025 ( .IN1(n9970), .IN2(n9971), .QN(g34006) );
  NAND2X0 U10026 ( .IN1(n9972), .IN2(g2361), .QN(n9971) );
  NAND2X0 U10027 ( .IN1(n9973), .IN2(n8520), .QN(n9972) );
  NAND2X0 U10028 ( .IN1(n9974), .IN2(g2375), .QN(n9973) );
  NAND2X0 U10029 ( .IN1(n9975), .IN2(n8520), .QN(n9970) );
  NAND2X0 U10030 ( .IN1(n9976), .IN2(n9977), .QN(n9975) );
  NAND2X0 U10031 ( .IN1(n9978), .IN2(n9979), .QN(n9977) );
  NAND2X0 U10032 ( .IN1(n9980), .IN2(n9981), .QN(n9979) );
  NAND2X0 U10033 ( .IN1(n7786), .IN2(n9982), .QN(n9981) );
  NAND2X0 U10034 ( .IN1(n9983), .IN2(g2375), .QN(n9976) );
  NAND2X0 U10035 ( .IN1(n9982), .IN2(n9984), .QN(n9983) );
  NAND2X0 U10036 ( .IN1(n9974), .IN2(g2287), .QN(n9984) );
  INVX0 U10037 ( .INP(n9978), .ZN(n9974) );
  NAND2X0 U10038 ( .IN1(n9985), .IN2(n9986), .QN(n9978) );
  NAND2X0 U10039 ( .IN1(n9987), .IN2(n5755), .QN(n9986) );
  NAND2X0 U10040 ( .IN1(n9988), .IN2(n9989), .QN(n9985) );
  NAND3X0 U10041 ( .IN1(n9990), .IN2(n9991), .IN3(n9992), .QN(g34005) );
  NAND2X0 U10042 ( .IN1(n9993), .IN2(n9967), .QN(n9992) );
  OR3X1 U10043 ( .IN1(n9993), .IN2(n5802), .IN3(n8539), .Q(n9991) );
  NOR2X0 U10044 ( .IN1(n9994), .IN2(n5537), .QN(n9993) );
  NAND2X0 U10045 ( .IN1(n8623), .IN2(g2303), .QN(n9990) );
  NAND3X0 U10046 ( .IN1(n9995), .IN2(n9996), .IN3(n9997), .QN(g34004) );
  NAND2X0 U10047 ( .IN1(n9998), .IN2(n9967), .QN(n9997) );
  INVX0 U10048 ( .INP(n9999), .ZN(n9998) );
  NAND3X0 U10049 ( .IN1(n9999), .IN2(n9314), .IN3(n8498), .QN(n9996) );
  NAND2X0 U10050 ( .IN1(n10000), .IN2(n5353), .QN(n9999) );
  NAND2X0 U10051 ( .IN1(n8623), .IN2(g2315), .QN(n9995) );
  NAND3X0 U10052 ( .IN1(n10001), .IN2(n10002), .IN3(n10003), .QN(g34003) );
  NAND2X0 U10053 ( .IN1(n10004), .IN2(n9967), .QN(n10003) );
  INVX0 U10054 ( .INP(n10005), .ZN(n10004) );
  NAND3X0 U10055 ( .IN1(n10005), .IN2(g2307), .IN3(n8498), .QN(n10002) );
  NAND3X0 U10056 ( .IN1(g2287), .IN2(g2361), .IN3(n9982), .QN(n10005) );
  NAND2X0 U10057 ( .IN1(n8622), .IN2(n9314), .QN(n10001) );
  NAND3X0 U10058 ( .IN1(n10006), .IN2(n10007), .IN3(n10008), .QN(g34002) );
  NAND2X0 U10059 ( .IN1(n10009), .IN2(n9967), .QN(n10008) );
  INVX0 U10060 ( .INP(n10010), .ZN(n10009) );
  NAND3X0 U10061 ( .IN1(n10010), .IN2(g2303), .IN3(n8498), .QN(n10007) );
  NAND2X0 U10062 ( .IN1(n10000), .IN2(n5537), .QN(n10010) );
  NAND2X0 U10063 ( .IN1(n8622), .IN2(g2295), .QN(n10006) );
  NAND3X0 U10064 ( .IN1(n10011), .IN2(n10012), .IN3(n10013), .QN(g34001) );
  NAND2X0 U10065 ( .IN1(n10014), .IN2(n9967), .QN(n10013) );
  AND3X1 U10066 ( .IN1(n10015), .IN2(n10016), .IN3(n8528), .Q(n9967) );
  NAND2X0 U10067 ( .IN1(n9987), .IN2(g1585), .QN(n10016) );
  OR2X1 U10068 ( .IN1(n9988), .IN2(n9987), .Q(n10015) );
  INVX0 U10069 ( .INP(n9989), .ZN(n9987) );
  NAND2X0 U10070 ( .IN1(n9906), .IN2(n10017), .QN(n9988) );
  OR3X1 U10071 ( .IN1(n10014), .IN2(n5815), .IN3(n8537), .Q(n10012) );
  NOR2X0 U10072 ( .IN1(n9994), .IN2(n5353), .QN(n10014) );
  NAND2X0 U10073 ( .IN1(n8622), .IN2(g2299), .QN(n10011) );
  NAND3X0 U10074 ( .IN1(n10018), .IN2(n10019), .IN3(n10020), .QN(g34000) );
  NAND2X0 U10075 ( .IN1(n8622), .IN2(g2246), .QN(n10020) );
  NAND2X0 U10076 ( .IN1(n10021), .IN2(n10022), .QN(n10019) );
  NAND2X0 U10077 ( .IN1(n10023), .IN2(g2165), .QN(n10018) );
  NAND2X0 U10078 ( .IN1(n10024), .IN2(n10025), .QN(g33999) );
  NAND2X0 U10079 ( .IN1(n10026), .IN2(g2227), .QN(n10025) );
  NAND2X0 U10080 ( .IN1(n10027), .IN2(n8520), .QN(n10026) );
  NAND2X0 U10081 ( .IN1(n10028), .IN2(g2241), .QN(n10027) );
  NAND2X0 U10082 ( .IN1(n10029), .IN2(n8520), .QN(n10024) );
  NAND2X0 U10083 ( .IN1(n10030), .IN2(n10031), .QN(n10029) );
  NAND2X0 U10084 ( .IN1(n10032), .IN2(n10033), .QN(n10031) );
  NAND2X0 U10085 ( .IN1(n10034), .IN2(n10035), .QN(n10033) );
  NAND2X0 U10086 ( .IN1(n7788), .IN2(n10036), .QN(n10035) );
  NAND2X0 U10087 ( .IN1(n10037), .IN2(g2241), .QN(n10030) );
  NAND2X0 U10088 ( .IN1(n10036), .IN2(n10038), .QN(n10037) );
  NAND2X0 U10089 ( .IN1(n10028), .IN2(g2153), .QN(n10038) );
  INVX0 U10090 ( .INP(n10032), .ZN(n10028) );
  NAND2X0 U10091 ( .IN1(n10039), .IN2(n10040), .QN(n10032) );
  NAND2X0 U10092 ( .IN1(n10041), .IN2(g1589), .QN(n10040) );
  NAND2X0 U10093 ( .IN1(n10042), .IN2(n10043), .QN(n10039) );
  NAND3X0 U10094 ( .IN1(n10044), .IN2(n10045), .IN3(n10046), .QN(g33998) );
  NAND2X0 U10095 ( .IN1(n10047), .IN2(n10021), .QN(n10046) );
  OR3X1 U10096 ( .IN1(n10047), .IN2(n5803), .IN3(n8531), .Q(n10045) );
  NOR2X0 U10097 ( .IN1(n10048), .IN2(n5538), .QN(n10047) );
  NAND2X0 U10098 ( .IN1(n8622), .IN2(g2169), .QN(n10044) );
  NAND3X0 U10099 ( .IN1(n10049), .IN2(n10050), .IN3(n10051), .QN(g33997) );
  NAND2X0 U10100 ( .IN1(n10052), .IN2(n10021), .QN(n10051) );
  INVX0 U10101 ( .INP(n10053), .ZN(n10052) );
  NAND3X0 U10102 ( .IN1(n10053), .IN2(n9352), .IN3(n8498), .QN(n10050) );
  NAND2X0 U10103 ( .IN1(n10054), .IN2(n5356), .QN(n10053) );
  NAND2X0 U10104 ( .IN1(n8622), .IN2(g2181), .QN(n10049) );
  NAND3X0 U10105 ( .IN1(n10055), .IN2(n10056), .IN3(n10057), .QN(g33996) );
  NAND2X0 U10106 ( .IN1(n10058), .IN2(n10021), .QN(n10057) );
  INVX0 U10107 ( .INP(n10059), .ZN(n10058) );
  NAND3X0 U10108 ( .IN1(n10059), .IN2(g2173), .IN3(n8498), .QN(n10056) );
  NAND3X0 U10109 ( .IN1(g2153), .IN2(g2227), .IN3(n10036), .QN(n10059) );
  NAND2X0 U10110 ( .IN1(n8622), .IN2(n9352), .QN(n10055) );
  NAND3X0 U10111 ( .IN1(n10060), .IN2(n10061), .IN3(n10062), .QN(g33995) );
  NAND2X0 U10112 ( .IN1(n10063), .IN2(n10021), .QN(n10062) );
  INVX0 U10113 ( .INP(n10064), .ZN(n10063) );
  NAND3X0 U10114 ( .IN1(n10064), .IN2(g2169), .IN3(n8498), .QN(n10061) );
  NAND2X0 U10115 ( .IN1(n10054), .IN2(n5538), .QN(n10064) );
  NAND2X0 U10116 ( .IN1(n8621), .IN2(g2161), .QN(n10060) );
  NAND3X0 U10117 ( .IN1(n10065), .IN2(n10066), .IN3(n10067), .QN(g33994) );
  NAND2X0 U10118 ( .IN1(n10068), .IN2(n10021), .QN(n10067) );
  AND3X1 U10119 ( .IN1(n10069), .IN2(n10070), .IN3(n8528), .Q(n10021) );
  OR2X1 U10120 ( .IN1(n10042), .IN2(n10041), .Q(n10070) );
  NAND2X0 U10121 ( .IN1(n9906), .IN2(n10071), .QN(n10042) );
  AND2X1 U10122 ( .IN1(n10072), .IN2(g4180), .Q(n9906) );
  NAND2X0 U10123 ( .IN1(n10041), .IN2(n5757), .QN(n10069) );
  INVX0 U10124 ( .INP(n10043), .ZN(n10041) );
  OR3X1 U10125 ( .IN1(n10068), .IN2(n5812), .IN3(n8540), .Q(n10066) );
  NOR2X0 U10126 ( .IN1(n10048), .IN2(n5356), .QN(n10068) );
  NAND2X0 U10127 ( .IN1(n8621), .IN2(g2165), .QN(n10065) );
  NAND3X0 U10128 ( .IN1(n10073), .IN2(n10074), .IN3(n10075), .QN(g33993) );
  NAND2X0 U10129 ( .IN1(n8621), .IN2(g2089), .QN(n10075) );
  NAND2X0 U10130 ( .IN1(n10076), .IN2(n10077), .QN(n10074) );
  NAND2X0 U10131 ( .IN1(n10078), .IN2(g2008), .QN(n10073) );
  NAND2X0 U10132 ( .IN1(n10079), .IN2(n10080), .QN(g33992) );
  NAND2X0 U10133 ( .IN1(n10081), .IN2(g2070), .QN(n10080) );
  NAND2X0 U10134 ( .IN1(n10082), .IN2(n8520), .QN(n10081) );
  NAND2X0 U10135 ( .IN1(n10083), .IN2(g2084), .QN(n10082) );
  NAND2X0 U10136 ( .IN1(n10084), .IN2(n8519), .QN(n10079) );
  NAND2X0 U10137 ( .IN1(n10085), .IN2(n10086), .QN(n10084) );
  NAND2X0 U10138 ( .IN1(n10087), .IN2(n10088), .QN(n10086) );
  NAND2X0 U10139 ( .IN1(n10089), .IN2(n10090), .QN(n10088) );
  NAND2X0 U10140 ( .IN1(n7783), .IN2(n10091), .QN(n10090) );
  NAND2X0 U10141 ( .IN1(n10092), .IN2(g2084), .QN(n10085) );
  NAND2X0 U10142 ( .IN1(n10091), .IN2(n10093), .QN(n10092) );
  NAND2X0 U10143 ( .IN1(n10083), .IN2(g1996), .QN(n10093) );
  INVX0 U10144 ( .INP(n10087), .ZN(n10083) );
  NAND2X0 U10145 ( .IN1(n10094), .IN2(n10095), .QN(n10087) );
  NAND2X0 U10146 ( .IN1(n5756), .IN2(n10096), .QN(n10095) );
  NAND2X0 U10147 ( .IN1(n10097), .IN2(n10098), .QN(n10094) );
  NAND3X0 U10148 ( .IN1(n10099), .IN2(n10100), .IN3(n10101), .QN(g33991) );
  NAND2X0 U10149 ( .IN1(n10102), .IN2(n10076), .QN(n10101) );
  OR3X1 U10150 ( .IN1(n10102), .IN2(n5801), .IN3(n8539), .Q(n10100) );
  NOR2X0 U10151 ( .IN1(n10103), .IN2(n5535), .QN(n10102) );
  NAND2X0 U10152 ( .IN1(n8621), .IN2(g2012), .QN(n10099) );
  NAND3X0 U10153 ( .IN1(n10104), .IN2(n10105), .IN3(n10106), .QN(g33990) );
  NAND2X0 U10154 ( .IN1(n10107), .IN2(n10076), .QN(n10106) );
  INVX0 U10155 ( .INP(n10108), .ZN(n10107) );
  NAND3X0 U10156 ( .IN1(n10108), .IN2(n9312), .IN3(n8499), .QN(n10105) );
  NAND2X0 U10157 ( .IN1(n10109), .IN2(n5355), .QN(n10108) );
  NAND2X0 U10158 ( .IN1(n8621), .IN2(g2024), .QN(n10104) );
  NAND3X0 U10159 ( .IN1(n10110), .IN2(n10111), .IN3(n10112), .QN(g33989) );
  NAND2X0 U10160 ( .IN1(n10113), .IN2(n10076), .QN(n10112) );
  INVX0 U10161 ( .INP(n10114), .ZN(n10113) );
  NAND3X0 U10162 ( .IN1(n10114), .IN2(g2016), .IN3(n8499), .QN(n10111) );
  NAND3X0 U10163 ( .IN1(g1996), .IN2(g2070), .IN3(n10091), .QN(n10114) );
  NAND2X0 U10164 ( .IN1(n8621), .IN2(n9312), .QN(n10110) );
  NAND3X0 U10165 ( .IN1(n10115), .IN2(n10116), .IN3(n10117), .QN(g33988) );
  NAND2X0 U10166 ( .IN1(n10118), .IN2(n10076), .QN(n10117) );
  INVX0 U10167 ( .INP(n10119), .ZN(n10118) );
  NAND3X0 U10168 ( .IN1(n10119), .IN2(g2012), .IN3(n8499), .QN(n10116) );
  NAND2X0 U10169 ( .IN1(n10109), .IN2(n5535), .QN(n10119) );
  NAND2X0 U10170 ( .IN1(n8621), .IN2(g2004), .QN(n10115) );
  NAND3X0 U10171 ( .IN1(n10120), .IN2(n10121), .IN3(n10122), .QN(g33987) );
  NAND2X0 U10172 ( .IN1(n10123), .IN2(n10076), .QN(n10122) );
  AND3X1 U10173 ( .IN1(n10124), .IN2(n10125), .IN3(n8528), .Q(n10076) );
  NAND2X0 U10174 ( .IN1(n10096), .IN2(g30332), .QN(n10125) );
  OR2X1 U10175 ( .IN1(n10097), .IN2(n10096), .Q(n10124) );
  INVX0 U10176 ( .INP(n10098), .ZN(n10096) );
  NAND2X0 U10177 ( .IN1(n10126), .IN2(n10127), .QN(n10097) );
  OR3X1 U10178 ( .IN1(n10123), .IN2(n5818), .IN3(n8539), .Q(n10121) );
  NOR2X0 U10179 ( .IN1(n10103), .IN2(n5355), .QN(n10123) );
  NAND2X0 U10180 ( .IN1(n8620), .IN2(g2008), .QN(n10120) );
  NAND3X0 U10181 ( .IN1(n10128), .IN2(n10129), .IN3(n10130), .QN(g33986) );
  NAND2X0 U10182 ( .IN1(n8620), .IN2(g1955), .QN(n10130) );
  NAND2X0 U10183 ( .IN1(n10131), .IN2(n10132), .QN(n10129) );
  NAND2X0 U10184 ( .IN1(n10133), .IN2(g1874), .QN(n10128) );
  NAND2X0 U10185 ( .IN1(n10134), .IN2(n10135), .QN(g33985) );
  NAND2X0 U10186 ( .IN1(n10136), .IN2(g1936), .QN(n10135) );
  NAND2X0 U10187 ( .IN1(n10137), .IN2(n8519), .QN(n10136) );
  NAND2X0 U10188 ( .IN1(n10138), .IN2(g1950), .QN(n10137) );
  NAND2X0 U10189 ( .IN1(n10139), .IN2(n8519), .QN(n10134) );
  NAND2X0 U10190 ( .IN1(n10140), .IN2(n10141), .QN(n10139) );
  NAND2X0 U10191 ( .IN1(n10142), .IN2(n10143), .QN(n10141) );
  NAND2X0 U10192 ( .IN1(n10144), .IN2(n10145), .QN(n10143) );
  NAND2X0 U10193 ( .IN1(n7787), .IN2(n10146), .QN(n10145) );
  NAND2X0 U10194 ( .IN1(n10147), .IN2(g1950), .QN(n10140) );
  NAND2X0 U10195 ( .IN1(n10146), .IN2(n10148), .QN(n10147) );
  NAND2X0 U10196 ( .IN1(test_so8), .IN2(n10138), .QN(n10148) );
  INVX0 U10197 ( .INP(n10142), .ZN(n10138) );
  NAND2X0 U10198 ( .IN1(n10149), .IN2(n10150), .QN(n10142) );
  NAND2X0 U10199 ( .IN1(n10151), .IN2(g1246), .QN(n10150) );
  NAND2X0 U10200 ( .IN1(n10152), .IN2(n10153), .QN(n10149) );
  NAND3X0 U10201 ( .IN1(n10154), .IN2(n10155), .IN3(n10156), .QN(g33984) );
  NAND2X0 U10202 ( .IN1(n10157), .IN2(n10131), .QN(n10156) );
  OR3X1 U10203 ( .IN1(n10157), .IN2(n5799), .IN3(n8538), .Q(n10155) );
  NOR2X0 U10204 ( .IN1(n10158), .IN2(n10159), .QN(n10157) );
  NAND2X0 U10205 ( .IN1(n8620), .IN2(g1878), .QN(n10154) );
  NAND3X0 U10206 ( .IN1(n10160), .IN2(n10161), .IN3(n10162), .QN(g33983) );
  NAND2X0 U10207 ( .IN1(n10163), .IN2(n10131), .QN(n10162) );
  INVX0 U10208 ( .INP(n10164), .ZN(n10163) );
  NAND3X0 U10209 ( .IN1(n10164), .IN2(n9280), .IN3(n8499), .QN(n10161) );
  NAND2X0 U10210 ( .IN1(n10165), .IN2(n8205), .QN(n10164) );
  NAND2X0 U10211 ( .IN1(n8620), .IN2(g1890), .QN(n10160) );
  NAND3X0 U10212 ( .IN1(n10166), .IN2(n10167), .IN3(n10168), .QN(g33982) );
  NAND2X0 U10213 ( .IN1(n10169), .IN2(n10131), .QN(n10168) );
  INVX0 U10214 ( .INP(n10170), .ZN(n10169) );
  NAND3X0 U10215 ( .IN1(n10170), .IN2(g1882), .IN3(n8499), .QN(n10167) );
  NAND2X0 U10216 ( .IN1(n10171), .IN2(g1936), .QN(n10170) );
  NAND2X0 U10217 ( .IN1(n8620), .IN2(n9280), .QN(n10166) );
  NAND3X0 U10218 ( .IN1(n10172), .IN2(n10173), .IN3(n10174), .QN(g33981) );
  NAND2X0 U10219 ( .IN1(n10175), .IN2(n10131), .QN(n10174) );
  INVX0 U10220 ( .INP(n10176), .ZN(n10175) );
  NAND3X0 U10221 ( .IN1(n10176), .IN2(g1878), .IN3(n8499), .QN(n10173) );
  NAND2X0 U10222 ( .IN1(n10165), .IN2(n5534), .QN(n10176) );
  NAND2X0 U10223 ( .IN1(n8620), .IN2(g1870), .QN(n10172) );
  NAND3X0 U10224 ( .IN1(n10177), .IN2(n10178), .IN3(n10179), .QN(g33980) );
  NAND2X0 U10225 ( .IN1(n10180), .IN2(n10131), .QN(n10179) );
  AND3X1 U10226 ( .IN1(n10181), .IN2(n10182), .IN3(n8528), .Q(n10131) );
  OR2X1 U10227 ( .IN1(n10152), .IN2(n10151), .Q(n10182) );
  NAND2X0 U10228 ( .IN1(n10126), .IN2(n10183), .QN(n10152) );
  NAND2X0 U10229 ( .IN1(n5526), .IN2(n10151), .QN(n10181) );
  INVX0 U10230 ( .INP(n10153), .ZN(n10151) );
  INVX0 U10231 ( .INP(n10184), .ZN(n10180) );
  NAND3X0 U10232 ( .IN1(n10184), .IN2(g1870), .IN3(n8499), .QN(n10178) );
  NAND2X0 U10233 ( .IN1(n10171), .IN2(n5503), .QN(n10184) );
  NAND2X0 U10234 ( .IN1(n8620), .IN2(g1874), .QN(n10177) );
  NAND3X0 U10235 ( .IN1(n10185), .IN2(n10186), .IN3(n10187), .QN(g33979) );
  NAND2X0 U10236 ( .IN1(n8619), .IN2(g1821), .QN(n10187) );
  NAND2X0 U10237 ( .IN1(n10188), .IN2(n10189), .QN(n10186) );
  NAND2X0 U10238 ( .IN1(n10190), .IN2(g1740), .QN(n10185) );
  NAND2X0 U10239 ( .IN1(n10191), .IN2(n10192), .QN(g33978) );
  NAND2X0 U10240 ( .IN1(n10193), .IN2(g1802), .QN(n10192) );
  NAND2X0 U10241 ( .IN1(n10194), .IN2(n8519), .QN(n10193) );
  NAND2X0 U10242 ( .IN1(n10195), .IN2(g1816), .QN(n10194) );
  NAND2X0 U10243 ( .IN1(n10196), .IN2(n8519), .QN(n10191) );
  NAND2X0 U10244 ( .IN1(n10197), .IN2(n10198), .QN(n10196) );
  NAND2X0 U10245 ( .IN1(n10199), .IN2(n10200), .QN(n10198) );
  NAND2X0 U10246 ( .IN1(n10201), .IN2(n10202), .QN(n10200) );
  NAND2X0 U10247 ( .IN1(n7708), .IN2(n10203), .QN(n10202) );
  NAND2X0 U10248 ( .IN1(n10204), .IN2(g1816), .QN(n10197) );
  NAND2X0 U10249 ( .IN1(n10203), .IN2(n10205), .QN(n10204) );
  NAND2X0 U10250 ( .IN1(n10195), .IN2(g1728), .QN(n10205) );
  INVX0 U10251 ( .INP(n10199), .ZN(n10195) );
  NAND2X0 U10252 ( .IN1(n10206), .IN2(n10207), .QN(n10199) );
  NAND2X0 U10253 ( .IN1(n10208), .IN2(n5756), .QN(n10207) );
  NAND2X0 U10254 ( .IN1(n10209), .IN2(n10210), .QN(n10206) );
  NAND3X0 U10255 ( .IN1(n10211), .IN2(n10212), .IN3(n10213), .QN(g33977) );
  NAND2X0 U10256 ( .IN1(n10214), .IN2(n10188), .QN(n10213) );
  OR3X1 U10257 ( .IN1(n10214), .IN2(n5804), .IN3(n8537), .Q(n10212) );
  NOR2X0 U10258 ( .IN1(n10215), .IN2(n5536), .QN(n10214) );
  NAND2X0 U10259 ( .IN1(n8619), .IN2(g1744), .QN(n10211) );
  NAND3X0 U10260 ( .IN1(n10216), .IN2(n10217), .IN3(n10218), .QN(g33976) );
  NAND2X0 U10261 ( .IN1(n10219), .IN2(n10188), .QN(n10218) );
  INVX0 U10262 ( .INP(n10220), .ZN(n10219) );
  NAND3X0 U10263 ( .IN1(n10220), .IN2(g1752), .IN3(n8499), .QN(n10217) );
  NAND2X0 U10264 ( .IN1(n10221), .IN2(n5352), .QN(n10220) );
  NAND2X0 U10265 ( .IN1(n8619), .IN2(g1756), .QN(n10216) );
  NAND3X0 U10266 ( .IN1(n10222), .IN2(n10223), .IN3(n10224), .QN(g33975) );
  NAND2X0 U10267 ( .IN1(n10225), .IN2(n10188), .QN(n10224) );
  INVX0 U10268 ( .INP(n10226), .ZN(n10225) );
  NAND3X0 U10269 ( .IN1(n10226), .IN2(g1748), .IN3(n8500), .QN(n10223) );
  NAND3X0 U10270 ( .IN1(g1728), .IN2(g1802), .IN3(n10203), .QN(n10226) );
  NAND2X0 U10271 ( .IN1(n8619), .IN2(g1752), .QN(n10222) );
  NAND3X0 U10272 ( .IN1(n10227), .IN2(n10228), .IN3(n10229), .QN(g33974) );
  NAND2X0 U10273 ( .IN1(n10230), .IN2(n10188), .QN(n10229) );
  INVX0 U10274 ( .INP(n10231), .ZN(n10230) );
  NAND3X0 U10275 ( .IN1(n10231), .IN2(g1744), .IN3(n8500), .QN(n10228) );
  NAND2X0 U10276 ( .IN1(n10221), .IN2(n5536), .QN(n10231) );
  NAND2X0 U10277 ( .IN1(n8619), .IN2(g1736), .QN(n10227) );
  NAND3X0 U10278 ( .IN1(n10232), .IN2(n10233), .IN3(n10234), .QN(g33973) );
  NAND2X0 U10279 ( .IN1(n10235), .IN2(n10188), .QN(n10234) );
  AND3X1 U10280 ( .IN1(n10236), .IN2(n10237), .IN3(n8455), .Q(n10188) );
  NAND2X0 U10281 ( .IN1(n10208), .IN2(g30332), .QN(n10237) );
  OR2X1 U10282 ( .IN1(n10209), .IN2(n10208), .Q(n10236) );
  NAND2X0 U10283 ( .IN1(n10126), .IN2(n10238), .QN(n10209) );
  OR3X1 U10284 ( .IN1(n10235), .IN2(n5817), .IN3(n8538), .Q(n10233) );
  NOR2X0 U10285 ( .IN1(n10215), .IN2(n5352), .QN(n10235) );
  NAND2X0 U10286 ( .IN1(n8619), .IN2(g1740), .QN(n10232) );
  NAND3X0 U10287 ( .IN1(n10239), .IN2(n10240), .IN3(n10241), .QN(g33972) );
  NAND2X0 U10288 ( .IN1(n8619), .IN2(g1687), .QN(n10241) );
  NAND2X0 U10289 ( .IN1(n10242), .IN2(n10243), .QN(n10240) );
  NAND2X0 U10290 ( .IN1(n10244), .IN2(g1604), .QN(n10239) );
  NAND2X0 U10291 ( .IN1(n10245), .IN2(n10246), .QN(g33971) );
  NAND2X0 U10292 ( .IN1(n10247), .IN2(g1668), .QN(n10246) );
  NAND2X0 U10293 ( .IN1(n10248), .IN2(n8519), .QN(n10247) );
  NAND2X0 U10294 ( .IN1(n10249), .IN2(g1682), .QN(n10248) );
  NAND2X0 U10295 ( .IN1(n10250), .IN2(n8519), .QN(n10245) );
  NAND2X0 U10296 ( .IN1(n10251), .IN2(n10252), .QN(n10250) );
  NAND2X0 U10297 ( .IN1(n10253), .IN2(n10254), .QN(n10252) );
  NAND2X0 U10298 ( .IN1(n10255), .IN2(n10256), .QN(n10254) );
  NAND2X0 U10299 ( .IN1(n7789), .IN2(n10257), .QN(n10256) );
  NAND2X0 U10300 ( .IN1(n10258), .IN2(g1682), .QN(n10251) );
  NAND2X0 U10301 ( .IN1(n10257), .IN2(n10259), .QN(n10258) );
  NAND2X0 U10302 ( .IN1(n10249), .IN2(g1592), .QN(n10259) );
  INVX0 U10303 ( .INP(n10253), .ZN(n10249) );
  NAND2X0 U10304 ( .IN1(n10260), .IN2(n10261), .QN(n10253) );
  NAND2X0 U10305 ( .IN1(n10262), .IN2(g1246), .QN(n10261) );
  NAND2X0 U10306 ( .IN1(n10263), .IN2(n10264), .QN(n10260) );
  NAND3X0 U10307 ( .IN1(n10265), .IN2(n10266), .IN3(n10267), .QN(g33970) );
  NAND2X0 U10308 ( .IN1(n10268), .IN2(n10242), .QN(n10267) );
  INVX0 U10309 ( .INP(n10269), .ZN(n10268) );
  NAND3X0 U10310 ( .IN1(n10269), .IN2(g1620), .IN3(n8500), .QN(n10266) );
  NAND2X0 U10311 ( .IN1(g31862), .IN2(n10257), .QN(n10269) );
  NAND2X0 U10312 ( .IN1(n8618), .IN2(g1608), .QN(n10265) );
  NAND3X0 U10313 ( .IN1(n10270), .IN2(n10271), .IN3(n10272), .QN(g33969) );
  NAND2X0 U10315 ( .IN1(n10273), .IN2(n10242), .QN(n10272) );
  INVX0 U10316 ( .INP(n10274), .ZN(n10273) );
  NAND3X0 U10317 ( .IN1(n10274), .IN2(n9303), .IN3(n8500), .QN(n10271) );
  NAND2X0 U10319 ( .IN1(n10275), .IN2(n5362), .QN(n10274) );
  NAND2X0 U10320 ( .IN1(n8618), .IN2(g1620), .QN(n10270) );
  NAND3X0 U10321 ( .IN1(n10276), .IN2(n10277), .IN3(n10278), .QN(g33968) );
  NAND2X0 U10322 ( .IN1(n10279), .IN2(n10242), .QN(n10278) );
  INVX0 U10323 ( .INP(n10280), .ZN(n10279) );
  NAND3X0 U10324 ( .IN1(n10280), .IN2(g1612), .IN3(n8500), .QN(n10277) );
  NAND2X0 U10325 ( .IN1(n10281), .IN2(g1668), .QN(n10280) );
  NAND2X0 U10326 ( .IN1(n8618), .IN2(n9303), .QN(n10276) );
  NAND3X0 U10327 ( .IN1(n10282), .IN2(n10283), .IN3(n10284), .QN(g33967) );
  NAND2X0 U10328 ( .IN1(n10285), .IN2(n10242), .QN(n10284) );
  INVX0 U10329 ( .INP(n10286), .ZN(n10285) );
  NAND3X0 U10330 ( .IN1(n10286), .IN2(g1608), .IN3(n8500), .QN(n10283) );
  NAND2X0 U10331 ( .IN1(n10275), .IN2(n5598), .QN(n10286) );
  NAND2X0 U10332 ( .IN1(n8618), .IN2(g1600), .QN(n10282) );
  NAND3X0 U10333 ( .IN1(n10287), .IN2(n10288), .IN3(n10289), .QN(g33966) );
  NAND2X0 U10334 ( .IN1(n10290), .IN2(n10242), .QN(n10289) );
  AND3X1 U10335 ( .IN1(n10291), .IN2(n10292), .IN3(n8412), .Q(n10242) );
  OR2X1 U10336 ( .IN1(n10263), .IN2(n10262), .Q(n10292) );
  NAND2X0 U10337 ( .IN1(n10126), .IN2(n10293), .QN(n10263) );
  AND2X1 U10338 ( .IN1(n10294), .IN2(g4180), .Q(n10126) );
  NAND2X0 U10339 ( .IN1(n10262), .IN2(n5526), .QN(n10291) );
  INVX0 U10340 ( .INP(n10264), .ZN(n10262) );
  INVX0 U10341 ( .INP(n10295), .ZN(n10290) );
  NAND3X0 U10342 ( .IN1(n10295), .IN2(g1600), .IN3(n8501), .QN(n10288) );
  NAND2X0 U10343 ( .IN1(n10281), .IN2(n5549), .QN(n10295) );
  NAND2X0 U10344 ( .IN1(n8618), .IN2(g1604), .QN(n10287) );
  NAND3X0 U10345 ( .IN1(n10296), .IN2(n10297), .IN3(n10298), .QN(g33965) );
  NAND2X0 U10346 ( .IN1(n8618), .IN2(g763), .QN(n10298) );
  NAND3X0 U10347 ( .IN1(n2404), .IN2(n10299), .IN3(g767), .QN(n10297) );
  INVX0 U10348 ( .INP(n2704), .ZN(n10299) );
  NAND2X0 U10349 ( .IN1(n2704), .IN2(n5333), .QN(n10296) );
  NAND3X0 U10350 ( .IN1(n10300), .IN2(n10301), .IN3(n10302), .QN(g33964) );
  NAND2X0 U10351 ( .IN1(n8618), .IN2(g595), .QN(n10302) );
  NAND3X0 U10352 ( .IN1(n2421), .IN2(n10303), .IN3(g599), .QN(n10301) );
  INVX0 U10353 ( .INP(n2706), .ZN(n10303) );
  NAND2X0 U10354 ( .IN1(n2706), .IN2(n5550), .QN(n10300) );
  NAND2X0 U10355 ( .IN1(n10304), .IN2(n10305), .QN(g33963) );
  NAND2X0 U10356 ( .IN1(n8621), .IN2(g29215), .QN(n10305) );
  NAND3X0 U10357 ( .IN1(n10306), .IN2(n10307), .IN3(n8500), .QN(n10304) );
  NAND3X0 U10358 ( .IN1(n10308), .IN2(n9194), .IN3(n10309), .QN(n10307) );
  NAND2X0 U10359 ( .IN1(g72), .IN2(g262), .QN(n10309) );
  NAND2X0 U10360 ( .IN1(n10310), .IN2(g269), .QN(n10308) );
  NAND2X0 U10361 ( .IN1(g73), .IN2(n10311), .QN(n10306) );
  NAND2X0 U10362 ( .IN1(n10310), .IN2(g255), .QN(n10311) );
  NAND2X0 U10363 ( .IN1(n10312), .IN2(n10313), .QN(g33962) );
  NAND2X0 U10364 ( .IN1(n8622), .IN2(g479), .QN(n10313) );
  NAND3X0 U10365 ( .IN1(n10314), .IN2(n10315), .IN3(n8501), .QN(n10312) );
  NAND3X0 U10366 ( .IN1(n10316), .IN2(n9194), .IN3(n10317), .QN(n10315) );
  NAND2X0 U10367 ( .IN1(g72), .IN2(g239), .QN(n10317) );
  INVX0 U10368 ( .INP(g73), .ZN(n9194) );
  NAND2X0 U10369 ( .IN1(n10310), .IN2(g246), .QN(n10316) );
  NAND2X0 U10370 ( .IN1(g73), .IN2(n10318), .QN(n10314) );
  NAND2X0 U10371 ( .IN1(n10319), .IN2(n10320), .QN(n10318) );
  NAND2X0 U10372 ( .IN1(n5597), .IN2(g72), .QN(n10320) );
  NAND2X0 U10373 ( .IN1(n7996), .IN2(n10321), .QN(n10319) );
  NAND3X0 U10374 ( .IN1(n10322), .IN2(n10323), .IN3(n10324), .QN(g33961) );
  NAND2X0 U10375 ( .IN1(n8624), .IN2(g294), .QN(n10324) );
  NAND3X0 U10376 ( .IN1(n8194), .IN2(n10325), .IN3(g298), .QN(n10323) );
  INVX0 U10377 ( .INP(n2989), .ZN(n10325) );
  NAND2X0 U10378 ( .IN1(n2989), .IN2(n5675), .QN(n10322) );
  NAND3X0 U10379 ( .IN1(n10326), .IN2(n10327), .IN3(n10328), .QN(g33960) );
  OR2X1 U10380 ( .IN1(n8478), .IN2(n5677), .Q(n10328) );
  OR3X1 U10381 ( .IN1(n9761), .IN2(n2991), .IN3(n5678), .Q(n10327) );
  NAND2X0 U10382 ( .IN1(n2991), .IN2(n5678), .QN(n10326) );
  NAND4X0 U10383 ( .IN1(n2668), .IN2(n8884), .IN3(g8403), .IN4(g8283), .QN(
        g33935) );
  INVX0 U10384 ( .INP(g34649), .ZN(n8884) );
  NAND4X0 U10385 ( .IN1(n10329), .IN2(n10330), .IN3(n10331), .IN4(n10332), 
        .QN(g34649) );
  NAND2X0 U10386 ( .IN1(n8880), .IN2(g4888), .QN(n10332) );
  NAND2X0 U10387 ( .IN1(n8881), .IN2(g4955), .QN(n10331) );
  NAND2X0 U10388 ( .IN1(n8882), .IN2(g4944), .QN(n10330) );
  NAND2X0 U10389 ( .IN1(n8883), .IN2(g4933), .QN(n10329) );
  NAND3X0 U10390 ( .IN1(n2668), .IN2(g4507), .IN3(n5541), .QN(g33874) );
  NAND4X0 U10391 ( .IN1(n8804), .IN2(n9630), .IN3(n8888), .IN4(n8889), .QN(
        g33659) );
  XNOR2X1 U10392 ( .IN1(g4104), .IN2(g73), .Q(n8889) );
  XNOR2X1 U10393 ( .IN1(g4108), .IN2(g72), .Q(n8888) );
  AND2X1 U10394 ( .IN1(g113), .IN2(n2668), .Q(n9630) );
  AND2X1 U10395 ( .IN1(n10333), .IN2(n10334), .Q(n8804) );
  NAND2X0 U10396 ( .IN1(n5350), .IN2(n10335), .QN(n10334) );
  NAND3X0 U10397 ( .IN1(n10336), .IN2(n10337), .IN3(n10338), .QN(n10335) );
  NAND2X0 U10398 ( .IN1(n10339), .IN2(n10340), .QN(n10338) );
  NAND3X0 U10399 ( .IN1(n10341), .IN2(n10342), .IN3(g4093), .QN(n10337) );
  NAND2X0 U10400 ( .IN1(n5480), .IN2(n10343), .QN(n10342) );
  NAND2X0 U10401 ( .IN1(n10344), .IN2(g4087), .QN(n10341) );
  NAND2X0 U10402 ( .IN1(g26801), .IN2(n9602), .QN(n10336) );
  NAND2X0 U10403 ( .IN1(n10345), .IN2(g4098), .QN(n10333) );
  NAND3X0 U10404 ( .IN1(n10346), .IN2(n10347), .IN3(n10348), .QN(n10345) );
  NAND2X0 U10405 ( .IN1(n10340), .IN2(n10349), .QN(n10348) );
  NAND3X0 U10406 ( .IN1(n10350), .IN2(n10351), .IN3(g4093), .QN(n10347) );
  NAND2X0 U10407 ( .IN1(n5480), .IN2(n10352), .QN(n10351) );
  NAND2X0 U10408 ( .IN1(n10353), .IN2(g4087), .QN(n10350) );
  NAND2X0 U10409 ( .IN1(n9602), .IN2(n10354), .QN(n10346) );
  NAND4X0 U10410 ( .IN1(n2668), .IN2(n8856), .IN3(g8353), .IN4(g8235), .QN(
        g33636) );
  INVX0 U10411 ( .INP(g34657), .ZN(n8856) );
  NAND4X0 U10412 ( .IN1(n10355), .IN2(n10356), .IN3(n10357), .IN4(n10358), 
        .QN(g34657) );
  NAND2X0 U10413 ( .IN1(n8852), .IN2(g4754), .QN(n10358) );
  NAND2X0 U10414 ( .IN1(n8853), .IN2(g4743), .QN(n10357) );
  NAND2X0 U10415 ( .IN1(n8854), .IN2(g4765), .QN(n10356) );
  NAND2X0 U10416 ( .IN1(n8855), .IN2(g4698), .QN(n10355) );
  NAND2X0 U10417 ( .IN1(n10359), .IN2(n10360), .QN(n2668) );
  NAND2X0 U10418 ( .IN1(g99), .IN2(g37), .QN(n10360) );
  NAND3X0 U10419 ( .IN1(n10361), .IN2(n10362), .IN3(n10363), .QN(g33627) );
  NAND3X0 U10420 ( .IN1(n10364), .IN2(n10365), .IN3(n8822), .QN(n10363) );
  NAND2X0 U10421 ( .IN1(n8623), .IN2(g6741), .QN(n10362) );
  NAND2X0 U10422 ( .IN1(n10366), .IN2(n8519), .QN(n10361) );
  NAND2X0 U10423 ( .IN1(n10367), .IN2(n10368), .QN(n10366) );
  NAND2X0 U10424 ( .IN1(n8198), .IN2(g6682), .QN(n10368) );
  NAND2X0 U10425 ( .IN1(n8819), .IN2(n10364), .QN(n10367) );
  NAND3X0 U10426 ( .IN1(n10369), .IN2(n10370), .IN3(n10371), .QN(g33626) );
  NAND2X0 U10427 ( .IN1(n10372), .IN2(g6741), .QN(n10371) );
  NAND4X0 U10428 ( .IN1(n10364), .IN2(n10365), .IN3(n5398), .IN4(n8506), .QN(
        n10370) );
  NAND2X0 U10429 ( .IN1(n10373), .IN2(n9289), .QN(n10364) );
  NAND2X0 U10430 ( .IN1(n8619), .IN2(g6736), .QN(n10369) );
  NAND3X0 U10431 ( .IN1(n10374), .IN2(n10375), .IN3(n10376), .QN(g33625) );
  NAND3X0 U10432 ( .IN1(n10377), .IN2(n10378), .IN3(n10379), .QN(n10376) );
  NAND2X0 U10433 ( .IN1(n8620), .IN2(g6395), .QN(n10375) );
  NAND2X0 U10434 ( .IN1(n10380), .IN2(n8519), .QN(n10374) );
  NAND2X0 U10435 ( .IN1(n10381), .IN2(n10382), .QN(n10380) );
  OR2X1 U10436 ( .IN1(n10377), .IN2(n5592), .Q(n10382) );
  NAND2X0 U10437 ( .IN1(n10383), .IN2(n10378), .QN(n10381) );
  NAND3X0 U10438 ( .IN1(n10384), .IN2(n10385), .IN3(n10386), .QN(g33624) );
  NAND2X0 U10439 ( .IN1(n10387), .IN2(g6395), .QN(n10386) );
  NAND4X0 U10440 ( .IN1(n10377), .IN2(n10378), .IN3(n5396), .IN4(n8506), .QN(
        n10385) );
  NAND2X0 U10441 ( .IN1(n10388), .IN2(n9292), .QN(n10378) );
  NAND2X0 U10442 ( .IN1(n8618), .IN2(g6390), .QN(n10384) );
  NAND3X0 U10443 ( .IN1(n10389), .IN2(n10390), .IN3(n10391), .QN(g33623) );
  NAND3X0 U10444 ( .IN1(n10392), .IN2(n10393), .IN3(n10394), .QN(n10391) );
  NAND2X0 U10445 ( .IN1(test_so57), .IN2(n8660), .QN(n10390) );
  NAND2X0 U10446 ( .IN1(n10395), .IN2(n8519), .QN(n10389) );
  NAND2X0 U10447 ( .IN1(n10396), .IN2(n10397), .QN(n10395) );
  OR2X1 U10448 ( .IN1(n10392), .IN2(n5589), .Q(n10397) );
  NAND2X0 U10449 ( .IN1(n10398), .IN2(n10393), .QN(n10396) );
  NAND3X0 U10450 ( .IN1(n10399), .IN2(n10400), .IN3(n10401), .QN(g33622) );
  NAND2X0 U10451 ( .IN1(n10402), .IN2(test_so57), .QN(n10401) );
  NAND4X0 U10452 ( .IN1(n10393), .IN2(n8216), .IN3(n10392), .IN4(n8506), .QN(
        n10400) );
  NAND2X0 U10453 ( .IN1(n10403), .IN2(n9292), .QN(n10393) );
  NAND2X0 U10454 ( .IN1(test_so50), .IN2(n8660), .QN(n10399) );
  NAND3X0 U10455 ( .IN1(n10404), .IN2(n10405), .IN3(n10406), .QN(g33621) );
  NAND3X0 U10456 ( .IN1(n10407), .IN2(n10408), .IN3(n10409), .QN(n10406) );
  NAND2X0 U10457 ( .IN1(n8617), .IN2(g5703), .QN(n10405) );
  NAND2X0 U10458 ( .IN1(n10410), .IN2(n8519), .QN(n10404) );
  NAND2X0 U10459 ( .IN1(n10411), .IN2(n10412), .QN(n10410) );
  OR2X1 U10460 ( .IN1(n10407), .IN2(n5593), .Q(n10412) );
  NAND2X0 U10461 ( .IN1(n10413), .IN2(n10408), .QN(n10411) );
  NAND3X0 U10462 ( .IN1(n10414), .IN2(n10415), .IN3(n10416), .QN(g33620) );
  NAND2X0 U10463 ( .IN1(n10417), .IN2(g5703), .QN(n10416) );
  NAND4X0 U10464 ( .IN1(n10407), .IN2(n10408), .IN3(n5397), .IN4(n8507), .QN(
        n10415) );
  NAND2X0 U10465 ( .IN1(n10418), .IN2(n9292), .QN(n10408) );
  NAND2X0 U10466 ( .IN1(n8617), .IN2(g5698), .QN(n10414) );
  NAND3X0 U10467 ( .IN1(n10419), .IN2(n10420), .IN3(n10421), .QN(g33619) );
  NAND3X0 U10468 ( .IN1(n10422), .IN2(g33959), .IN3(n8814), .QN(n10421) );
  NAND2X0 U10469 ( .IN1(n8617), .IN2(g5357), .QN(n10420) );
  NAND2X0 U10470 ( .IN1(n10423), .IN2(n8519), .QN(n10419) );
  NAND2X0 U10471 ( .IN1(n10424), .IN2(n10425), .QN(n10423) );
  NAND2X0 U10472 ( .IN1(n8196), .IN2(g5297), .QN(n10425) );
  NAND2X0 U10473 ( .IN1(n8812), .IN2(n10422), .QN(n10424) );
  NAND3X0 U10474 ( .IN1(n10426), .IN2(n10427), .IN3(n10428), .QN(g33618) );
  NAND2X0 U10475 ( .IN1(n10429), .IN2(g5357), .QN(n10428) );
  NAND4X0 U10476 ( .IN1(n10422), .IN2(g33959), .IN3(n5393), .IN4(n8506), .QN(
        n10427) );
  NAND2X0 U10477 ( .IN1(n10373), .IN2(n9292), .QN(n10422) );
  INVX0 U10478 ( .INP(n9633), .ZN(n9292) );
  NAND2X0 U10479 ( .IN1(n5323), .IN2(n10430), .QN(n9633) );
  AND2X1 U10480 ( .IN1(n3023), .IN2(n8208), .Q(n10373) );
  NAND2X0 U10481 ( .IN1(n8617), .IN2(g5352), .QN(n10426) );
  NAND3X0 U10482 ( .IN1(n10431), .IN2(n9836), .IN3(n10432), .QN(g33617) );
  NAND2X0 U10483 ( .IN1(n10433), .IN2(g4552), .QN(n10432) );
  NAND4X0 U10484 ( .IN1(n10434), .IN2(n10435), .IN3(n10436), .IN4(n9836), .QN(
        g33616) );
  NAND2X0 U10485 ( .IN1(n10437), .IN2(g4512), .QN(n10435) );
  OR2X1 U10486 ( .IN1(n8480), .IN2(n8134), .Q(n10434) );
  NAND2X0 U10487 ( .IN1(n3064), .IN2(n10438), .QN(g33615) );
  NAND2X0 U10488 ( .IN1(n10439), .IN2(g4108), .QN(n10438) );
  NAND2X0 U10489 ( .IN1(n10440), .IN2(n8519), .QN(n10439) );
  NAND2X0 U10490 ( .IN1(n8901), .IN2(n8001), .QN(n10440) );
  NAND3X0 U10491 ( .IN1(n10441), .IN2(n10442), .IN3(n10443), .QN(g33614) );
  NAND3X0 U10492 ( .IN1(n10444), .IN2(n10445), .IN3(n10446), .QN(n10443) );
  NAND2X0 U10493 ( .IN1(n8617), .IN2(g4054), .QN(n10442) );
  NAND2X0 U10494 ( .IN1(n10447), .IN2(n8519), .QN(n10441) );
  NAND2X0 U10495 ( .IN1(n10448), .IN2(n10449), .QN(n10447) );
  OR2X1 U10496 ( .IN1(n10444), .IN2(n5594), .Q(n10449) );
  NAND2X0 U10497 ( .IN1(n10450), .IN2(n10445), .QN(n10448) );
  NAND3X0 U10498 ( .IN1(n10451), .IN2(n10452), .IN3(n10453), .QN(g33613) );
  NAND2X0 U10499 ( .IN1(n10454), .IN2(g4054), .QN(n10453) );
  NAND4X0 U10500 ( .IN1(n10444), .IN2(n10445), .IN3(n5395), .IN4(n8506), .QN(
        n10452) );
  NAND2X0 U10501 ( .IN1(n10388), .IN2(n9289), .QN(n10445) );
  AND2X1 U10502 ( .IN1(n3033), .IN2(test_so81), .Q(n10388) );
  NAND2X0 U10503 ( .IN1(n8617), .IN2(g4049), .QN(n10451) );
  NAND3X0 U10504 ( .IN1(n10455), .IN2(n10456), .IN3(n10457), .QN(g33612) );
  NAND3X0 U10505 ( .IN1(n10458), .IN2(n10459), .IN3(n10460), .QN(n10457) );
  NAND2X0 U10506 ( .IN1(n8617), .IN2(g3703), .QN(n10456) );
  NAND2X0 U10507 ( .IN1(n10461), .IN2(n8519), .QN(n10455) );
  NAND2X0 U10508 ( .IN1(n10462), .IN2(n10463), .QN(n10461) );
  OR2X1 U10509 ( .IN1(n10458), .IN2(n5591), .Q(n10463) );
  NAND2X0 U10510 ( .IN1(n10464), .IN2(n10459), .QN(n10462) );
  NAND3X0 U10511 ( .IN1(n10465), .IN2(n10466), .IN3(n10467), .QN(g33611) );
  NAND2X0 U10512 ( .IN1(n10468), .IN2(g3703), .QN(n10467) );
  NAND4X0 U10513 ( .IN1(n10458), .IN2(n10459), .IN3(n5399), .IN4(n8507), .QN(
        n10466) );
  NAND2X0 U10514 ( .IN1(n10403), .IN2(n9289), .QN(n10459) );
  AND2X1 U10515 ( .IN1(n3033), .IN2(n8208), .Q(n10403) );
  NAND2X0 U10516 ( .IN1(n8616), .IN2(g3698), .QN(n10465) );
  NAND2X0 U10517 ( .IN1(n10469), .IN2(n10470), .QN(g33610) );
  NAND2X0 U10518 ( .IN1(n8616), .IN2(g3352), .QN(n10470) );
  NAND2X0 U10519 ( .IN1(n10471), .IN2(n8519), .QN(n10469) );
  NAND2X0 U10520 ( .IN1(n10472), .IN2(n10473), .QN(n10471) );
  NAND2X0 U10521 ( .IN1(n10474), .IN2(g3288), .QN(n10473) );
  NAND3X0 U10522 ( .IN1(n10475), .IN2(n10476), .IN3(n10477), .QN(n10472) );
  OR2X1 U10523 ( .IN1(n10478), .IN2(n10479), .Q(n10475) );
  NAND3X0 U10524 ( .IN1(n10480), .IN2(n10481), .IN3(n10482), .QN(g33609) );
  NAND2X0 U10525 ( .IN1(n10483), .IN2(g3352), .QN(n10482) );
  NAND4X0 U10526 ( .IN1(n5604), .IN2(n10476), .IN3(n10477), .IN4(n8506), .QN(
        n10481) );
  NAND2X0 U10527 ( .IN1(n10418), .IN2(n9289), .QN(n10476) );
  INVX0 U10528 ( .INP(n9632), .ZN(n9289) );
  NAND2X0 U10529 ( .IN1(n10430), .IN2(g4311), .QN(n9632) );
  AND2X1 U10530 ( .IN1(n10484), .IN2(n9193), .Q(n10430) );
  XOR2X1 U10531 ( .IN1(g72), .IN2(n5506), .Q(n9193) );
  XOR2X1 U10532 ( .IN1(n5540), .IN2(g73), .Q(n10484) );
  AND2X1 U10533 ( .IN1(n3023), .IN2(test_so81), .Q(n10418) );
  NAND2X0 U10534 ( .IN1(n8616), .IN2(g3347), .QN(n10480) );
  NAND4X0 U10535 ( .IN1(n10485), .IN2(n8807), .IN3(n10486), .IN4(n10487), .QN(
        g33608) );
  NAND3X0 U10536 ( .IN1(n9852), .IN2(g2759), .IN3(n8502), .QN(n10487) );
  NAND2X0 U10537 ( .IN1(test_so30), .IN2(n8564), .QN(n10486) );
  OR2X1 U10538 ( .IN1(n9852), .IN2(g2759), .Q(n10485) );
  NAND2X0 U10539 ( .IN1(n2790), .IN2(test_so30), .QN(n9852) );
  NAND3X0 U10540 ( .IN1(n10488), .IN2(n10489), .IN3(n10490), .QN(g33607) );
  NAND2X0 U10541 ( .IN1(n8616), .IN2(g2555), .QN(n10490) );
  NAND3X0 U10542 ( .IN1(n10491), .IN2(n10492), .IN3(n3102), .QN(n10489) );
  NAND2X0 U10543 ( .IN1(n10493), .IN2(n10494), .QN(n10492) );
  NAND4X0 U10544 ( .IN1(n5524), .IN2(n10495), .IN3(n9653), .IN4(g2629), .QN(
        n10494) );
  INVX0 U10545 ( .INP(n2726), .ZN(n9653) );
  NAND2X0 U10546 ( .IN1(n9659), .IN2(n5519), .QN(n2726) );
  NAND2X0 U10547 ( .IN1(n3111), .IN2(n8519), .QN(n10493) );
  NAND3X0 U10548 ( .IN1(g2629), .IN2(g112), .IN3(n5524), .QN(n10491) );
  NAND2X0 U10549 ( .IN1(n10496), .IN2(g2606), .QN(n10488) );
  OR2X1 U10550 ( .IN1(n10497), .IN2(n10498), .Q(n10496) );
  NOR2X0 U10551 ( .IN1(n3105), .IN2(n8548), .QN(n10497) );
  NAND3X0 U10552 ( .IN1(n10499), .IN2(n10500), .IN3(n10501), .QN(g33606) );
  NAND2X0 U10553 ( .IN1(n9858), .IN2(g2675), .QN(n10501) );
  NAND3X0 U10554 ( .IN1(n5457), .IN2(n9857), .IN3(n8502), .QN(n10500) );
  NAND2X0 U10555 ( .IN1(n8616), .IN2(g2671), .QN(n10499) );
  NAND3X0 U10556 ( .IN1(n10502), .IN2(n10503), .IN3(n10504), .QN(g33605) );
  NAND2X0 U10557 ( .IN1(n9858), .IN2(g2671), .QN(n10504) );
  NAND2X0 U10558 ( .IN1(test_so48), .IN2(n10505), .QN(n10503) );
  NAND2X0 U10559 ( .IN1(n10506), .IN2(n8519), .QN(n10505) );
  NAND2X0 U10560 ( .IN1(n9857), .IN2(g2661), .QN(n10506) );
  INVX0 U10561 ( .INP(n9869), .ZN(n9857) );
  OR4X1 U10562 ( .IN1(n9869), .IN2(n8544), .IN3(g2661), .IN4(test_so48), .Q(
        n10502) );
  NAND2X0 U10563 ( .IN1(n10507), .IN2(n10508), .QN(g33604) );
  NAND2X0 U10564 ( .IN1(test_so48), .IN2(n9858), .QN(n10508) );
  NAND2X0 U10565 ( .IN1(n10509), .IN2(g2661), .QN(n10507) );
  NAND2X0 U10566 ( .IN1(n10510), .IN2(n10511), .QN(g33603) );
  NAND2X0 U10567 ( .IN1(n9858), .IN2(g2648), .QN(n10511) );
  INVX0 U10568 ( .INP(n10509), .ZN(n9858) );
  NAND2X0 U10569 ( .IN1(n10509), .IN2(g2643), .QN(n10510) );
  NAND2X0 U10570 ( .IN1(n9869), .IN2(n8519), .QN(n10509) );
  NAND3X0 U10571 ( .IN1(n5351), .IN2(n9871), .IN3(n5521), .QN(n9869) );
  NAND3X0 U10572 ( .IN1(n10512), .IN2(n10513), .IN3(n10514), .QN(g33602) );
  NAND2X0 U10573 ( .IN1(n8616), .IN2(g2599), .QN(n10514) );
  NAND2X0 U10574 ( .IN1(n10515), .IN2(g2629), .QN(n10513) );
  NAND2X0 U10575 ( .IN1(n9889), .IN2(n10516), .QN(n10512) );
  NOR2X0 U10576 ( .IN1(n5524), .IN2(n10517), .QN(n9889) );
  NAND3X0 U10577 ( .IN1(n10518), .IN2(n10519), .IN3(n10520), .QN(g33601) );
  NAND2X0 U10578 ( .IN1(n10515), .IN2(g2599), .QN(n10520) );
  NAND2X0 U10579 ( .IN1(n8616), .IN2(g2606), .QN(n10519) );
  NAND4X0 U10580 ( .IN1(n10516), .IN2(g2555), .IN3(n9871), .IN4(n8507), .QN(
        n10518) );
  NAND2X0 U10581 ( .IN1(n10521), .IN2(n10522), .QN(g33600) );
  NAND4X0 U10582 ( .IN1(n5521), .IN2(n10523), .IN3(n8505), .IN4(n10516), .QN(
        n10522) );
  INVX0 U10583 ( .INP(n3111), .ZN(n10516) );
  NAND2X0 U10584 ( .IN1(n5351), .IN2(n9883), .QN(n10523) );
  NAND2X0 U10585 ( .IN1(n5524), .IN2(n9871), .QN(n9883) );
  NAND2X0 U10586 ( .IN1(n10515), .IN2(g2555), .QN(n10521) );
  NOR2X0 U10587 ( .IN1(n9871), .IN2(n8550), .QN(n10515) );
  INVX0 U10588 ( .INP(n10517), .ZN(n9871) );
  NOR2X0 U10589 ( .IN1(n9878), .IN2(n3102), .QN(n10517) );
  AND2X1 U10590 ( .IN1(n10524), .IN2(g1430), .Q(n3102) );
  NAND3X0 U10591 ( .IN1(n10525), .IN2(n8206), .IN3(n5364), .QN(n10524) );
  NAND3X0 U10592 ( .IN1(n10526), .IN2(n10072), .IN3(n9907), .QN(n9878) );
  NAND2X0 U10593 ( .IN1(n2549), .IN2(g1300), .QN(n9907) );
  NAND3X0 U10594 ( .IN1(g2689), .IN2(g2704), .IN3(g2697), .QN(n10526) );
  NAND4X0 U10595 ( .IN1(n10527), .IN2(n3121), .IN3(n10528), .IN4(n10529), .QN(
        g33599) );
  NAND2X0 U10596 ( .IN1(test_so79), .IN2(n8561), .QN(n10529) );
  NAND4X0 U10597 ( .IN1(n3122), .IN2(n10530), .IN3(n3131), .IN4(n8507), .QN(
        n10528) );
  NAND2X0 U10598 ( .IN1(n9644), .IN2(g112), .QN(n10530) );
  NAND4X0 U10599 ( .IN1(n3122), .IN2(n9644), .IN3(n10531), .IN4(n9645), .QN(
        n3121) );
  INVX0 U10600 ( .INP(n2727), .ZN(n9645) );
  NAND2X0 U10601 ( .IN1(n9659), .IN2(g504), .QN(n2727) );
  AND2X1 U10602 ( .IN1(n3116), .IN2(g518), .Q(n9659) );
  NOR2X0 U10603 ( .IN1(g2465), .IN2(n5522), .QN(n9644) );
  NAND2X0 U10604 ( .IN1(n10532), .IN2(g2472), .QN(n10527) );
  OR2X1 U10605 ( .IN1(n10533), .IN2(n10498), .Q(n10532) );
  NOR2X0 U10606 ( .IN1(n3125), .IN2(n8548), .QN(n10533) );
  NAND3X0 U10607 ( .IN1(n10534), .IN2(n10535), .IN3(n10536), .QN(g33598) );
  NAND2X0 U10608 ( .IN1(n9913), .IN2(g2541), .QN(n10536) );
  NAND3X0 U10609 ( .IN1(n5461), .IN2(n9912), .IN3(n8501), .QN(n10535) );
  NAND2X0 U10610 ( .IN1(n8615), .IN2(g2537), .QN(n10534) );
  NAND3X0 U10611 ( .IN1(n10537), .IN2(n10538), .IN3(n10539), .QN(g33597) );
  NAND2X0 U10612 ( .IN1(n9913), .IN2(g2537), .QN(n10539) );
  NAND2X0 U10613 ( .IN1(n10540), .IN2(g2533), .QN(n10538) );
  NAND2X0 U10614 ( .IN1(n10541), .IN2(n8519), .QN(n10540) );
  NAND2X0 U10615 ( .IN1(n9912), .IN2(g2527), .QN(n10541) );
  NAND4X0 U10616 ( .IN1(n9912), .IN2(n8506), .IN3(n5420), .IN4(n5761), .QN(
        n10537) );
  INVX0 U10617 ( .INP(n9924), .ZN(n9912) );
  NAND2X0 U10618 ( .IN1(n10542), .IN2(n10543), .QN(g33596) );
  NAND2X0 U10619 ( .IN1(n9913), .IN2(g2533), .QN(n10543) );
  NAND2X0 U10620 ( .IN1(n10544), .IN2(g2527), .QN(n10542) );
  NAND2X0 U10621 ( .IN1(n10545), .IN2(n10546), .QN(g33595) );
  NAND2X0 U10622 ( .IN1(n9913), .IN2(g2514), .QN(n10546) );
  INVX0 U10623 ( .INP(n10544), .ZN(n9913) );
  NAND2X0 U10624 ( .IN1(n10544), .IN2(g2509), .QN(n10545) );
  NAND2X0 U10625 ( .IN1(n9924), .IN2(n8519), .QN(n10544) );
  NAND3X0 U10626 ( .IN1(n9926), .IN2(n8204), .IN3(n5522), .QN(n9924) );
  NAND3X0 U10627 ( .IN1(n10547), .IN2(n10548), .IN3(n10549), .QN(g33594) );
  NAND2X0 U10628 ( .IN1(n8615), .IN2(g2465), .QN(n10549) );
  NAND2X0 U10629 ( .IN1(n10550), .IN2(g2495), .QN(n10548) );
  NAND2X0 U10630 ( .IN1(n9944), .IN2(n10551), .QN(n10547) );
  NOR2X0 U10631 ( .IN1(n5523), .IN2(n10552), .QN(n9944) );
  NAND3X0 U10632 ( .IN1(n10553), .IN2(n10554), .IN3(n10555), .QN(g33593) );
  NAND2X0 U10633 ( .IN1(n10550), .IN2(g2465), .QN(n10555) );
  NAND2X0 U10634 ( .IN1(n8615), .IN2(g2472), .QN(n10554) );
  NAND3X0 U10635 ( .IN1(n9950), .IN2(n10551), .IN3(n8486), .QN(n10553) );
  NOR2X0 U10636 ( .IN1(n8204), .IN2(n10552), .QN(n9950) );
  NAND2X0 U10637 ( .IN1(n10556), .IN2(n10557), .QN(g33592) );
  NAND4X0 U10638 ( .IN1(n5522), .IN2(n10558), .IN3(n8505), .IN4(n10551), .QN(
        n10557) );
  INVX0 U10639 ( .INP(n3131), .ZN(n10551) );
  NAND2X0 U10640 ( .IN1(n8204), .IN2(n10559), .QN(n10558) );
  NAND2X0 U10641 ( .IN1(n5523), .IN2(n9926), .QN(n10559) );
  NAND2X0 U10642 ( .IN1(n10550), .IN2(test_so79), .QN(n10556) );
  NOR2X0 U10643 ( .IN1(n9926), .IN2(n8549), .QN(n10550) );
  INVX0 U10644 ( .INP(n10552), .ZN(n9926) );
  NOR2X0 U10645 ( .IN1(n9933), .IN2(n3122), .QN(n10552) );
  AND2X1 U10646 ( .IN1(n10560), .IN2(g17423), .Q(n3122) );
  NAND2X0 U10647 ( .IN1(n10561), .IN2(n10525), .QN(n10560) );
  NAND3X0 U10648 ( .IN1(n10562), .IN2(n10072), .IN3(n9962), .QN(n9933) );
  NAND2X0 U10649 ( .IN1(n2549), .IN2(g1472), .QN(n9962) );
  NAND3X0 U10650 ( .IN1(g2697), .IN2(g2689), .IN3(n5377), .QN(n10562) );
  NAND3X0 U10651 ( .IN1(n10563), .IN2(n10564), .IN3(n10565), .QN(g33591) );
  NAND2X0 U10652 ( .IN1(n8615), .IN2(g2287), .QN(n10565) );
  NAND3X0 U10653 ( .IN1(n10566), .IN2(n10567), .IN3(n3141), .QN(n10564) );
  NAND2X0 U10654 ( .IN1(n10568), .IN2(n10569), .QN(n10567) );
  NAND4X0 U10655 ( .IN1(n5513), .IN2(n10495), .IN3(n9654), .IN4(g2361), .QN(
        n10569) );
  OR2X1 U10656 ( .IN1(n10570), .IN2(n8546), .Q(n10568) );
  NAND3X0 U10657 ( .IN1(g2361), .IN2(g112), .IN3(n5513), .QN(n10566) );
  NAND2X0 U10658 ( .IN1(n10571), .IN2(g2338), .QN(n10563) );
  OR2X1 U10659 ( .IN1(n10572), .IN2(n10498), .Q(n10571) );
  NOR2X0 U10660 ( .IN1(n3145), .IN2(n8549), .QN(n10572) );
  NAND3X0 U10661 ( .IN1(n10573), .IN2(n10574), .IN3(n10575), .QN(g33590) );
  NAND2X0 U10662 ( .IN1(n9969), .IN2(g2407), .QN(n10575) );
  NAND3X0 U10663 ( .IN1(n5459), .IN2(n9968), .IN3(n8486), .QN(n10574) );
  NAND2X0 U10664 ( .IN1(test_so31), .IN2(n8556), .QN(n10573) );
  NAND3X0 U10665 ( .IN1(n10576), .IN2(n10577), .IN3(n10578), .QN(g33589) );
  NAND2X0 U10666 ( .IN1(test_so31), .IN2(n9969), .QN(n10578) );
  NAND2X0 U10667 ( .IN1(n10579), .IN2(g2399), .QN(n10577) );
  NAND2X0 U10668 ( .IN1(n10580), .IN2(n8518), .QN(n10579) );
  NAND2X0 U10669 ( .IN1(n9968), .IN2(g2393), .QN(n10580) );
  NAND4X0 U10670 ( .IN1(n9968), .IN2(n8506), .IN3(n5421), .IN4(n5762), .QN(
        n10576) );
  INVX0 U10671 ( .INP(n9980), .ZN(n9968) );
  NAND2X0 U10672 ( .IN1(n10581), .IN2(n10582), .QN(g33588) );
  NAND2X0 U10673 ( .IN1(n9969), .IN2(g2399), .QN(n10582) );
  NAND2X0 U10674 ( .IN1(n10583), .IN2(g2393), .QN(n10581) );
  NAND2X0 U10675 ( .IN1(n10584), .IN2(n10585), .QN(g33587) );
  NAND2X0 U10676 ( .IN1(n9969), .IN2(g2380), .QN(n10585) );
  INVX0 U10677 ( .INP(n10583), .ZN(n9969) );
  NAND2X0 U10678 ( .IN1(n10583), .IN2(g2375), .QN(n10584) );
  NAND2X0 U10679 ( .IN1(n9980), .IN2(n8518), .QN(n10583) );
  NAND3X0 U10680 ( .IN1(n5353), .IN2(n9982), .IN3(n5537), .QN(n9980) );
  NAND3X0 U10681 ( .IN1(n10586), .IN2(n10587), .IN3(n10588), .QN(g33586) );
  NAND2X0 U10682 ( .IN1(n8615), .IN2(g2331), .QN(n10588) );
  NAND2X0 U10683 ( .IN1(n10589), .IN2(g2361), .QN(n10587) );
  NAND2X0 U10684 ( .IN1(n10000), .IN2(n10570), .QN(n10586) );
  NOR2X0 U10685 ( .IN1(n5513), .IN2(n10590), .QN(n10000) );
  NAND3X0 U10686 ( .IN1(n10591), .IN2(n10592), .IN3(n10593), .QN(g33585) );
  NAND2X0 U10687 ( .IN1(n10589), .IN2(g2331), .QN(n10593) );
  NAND2X0 U10688 ( .IN1(n8615), .IN2(g2338), .QN(n10592) );
  NAND4X0 U10689 ( .IN1(n9982), .IN2(g2287), .IN3(n10570), .IN4(n8507), .QN(
        n10591) );
  NAND2X0 U10690 ( .IN1(n10594), .IN2(n10595), .QN(g33584) );
  NAND2X0 U10691 ( .IN1(n10589), .IN2(g2287), .QN(n10595) );
  NOR2X0 U10692 ( .IN1(n9982), .IN2(n8550), .QN(n10589) );
  NAND4X0 U10693 ( .IN1(n5537), .IN2(n10596), .IN3(n10570), .IN4(n8507), .QN(
        n10594) );
  NAND2X0 U10694 ( .IN1(n3115), .IN2(n9654), .QN(n10570) );
  INVX0 U10695 ( .INP(n3146), .ZN(n9654) );
  NAND3X0 U10696 ( .IN1(n5287), .IN2(g504), .IN3(n3116), .QN(n3146) );
  NAND2X0 U10697 ( .IN1(n5353), .IN2(n9994), .QN(n10596) );
  NAND2X0 U10698 ( .IN1(n5513), .IN2(n9982), .QN(n9994) );
  INVX0 U10699 ( .INP(n10590), .ZN(n9982) );
  NOR2X0 U10700 ( .IN1(n9989), .IN2(n3141), .QN(n10590) );
  AND2X1 U10701 ( .IN1(n10597), .IN2(g17404), .Q(n3141) );
  NAND2X0 U10702 ( .IN1(n10598), .IN2(n10525), .QN(n10597) );
  NAND3X0 U10703 ( .IN1(n10599), .IN2(n10072), .IN3(n10017), .QN(n9989) );
  NAND2X0 U10704 ( .IN1(n2549), .IN2(g1448), .QN(n10017) );
  NAND3X0 U10705 ( .IN1(g2689), .IN2(g2704), .IN3(n5308), .QN(n10599) );
  NAND3X0 U10706 ( .IN1(n10600), .IN2(n10601), .IN3(n10602), .QN(g33583) );
  NAND2X0 U10707 ( .IN1(n8615), .IN2(g2153), .QN(n10602) );
  NAND3X0 U10708 ( .IN1(n10603), .IN2(n9641), .IN3(n3160), .QN(n10601) );
  NAND2X0 U10709 ( .IN1(n10604), .IN2(n10605), .QN(n10603) );
  NAND3X0 U10710 ( .IN1(n10531), .IN2(g2227), .IN3(n5514), .QN(n10605) );
  NAND3X0 U10711 ( .IN1(n10606), .IN2(n8481), .IN3(n3115), .QN(n10604) );
  NAND3X0 U10712 ( .IN1(g2227), .IN2(g112), .IN3(n5514), .QN(n10606) );
  NAND2X0 U10713 ( .IN1(n10607), .IN2(g2204), .QN(n10600) );
  OR2X1 U10714 ( .IN1(n10608), .IN2(n10498), .Q(n10607) );
  INVX0 U10715 ( .INP(n10609), .ZN(n10498) );
  NOR2X0 U10716 ( .IN1(n3164), .IN2(n8550), .QN(n10608) );
  NAND3X0 U10717 ( .IN1(n10610), .IN2(n10611), .IN3(n10612), .QN(g33582) );
  NAND2X0 U10718 ( .IN1(n10023), .IN2(g2273), .QN(n10612) );
  NAND3X0 U10719 ( .IN1(n5458), .IN2(n10022), .IN3(n8484), .QN(n10611) );
  NAND2X0 U10720 ( .IN1(n8614), .IN2(g2269), .QN(n10610) );
  NAND3X0 U10721 ( .IN1(n10613), .IN2(n10614), .IN3(n10615), .QN(g33581) );
  NAND2X0 U10722 ( .IN1(n10023), .IN2(g2269), .QN(n10615) );
  NAND2X0 U10723 ( .IN1(test_so62), .IN2(n10616), .QN(n10614) );
  NAND2X0 U10724 ( .IN1(n10617), .IN2(n8518), .QN(n10616) );
  NAND2X0 U10725 ( .IN1(n10022), .IN2(g2259), .QN(n10617) );
  INVX0 U10726 ( .INP(n10034), .ZN(n10022) );
  OR4X1 U10727 ( .IN1(n10034), .IN2(n8543), .IN3(g2259), .IN4(test_so62), .Q(
        n10613) );
  NAND2X0 U10728 ( .IN1(n10618), .IN2(n10619), .QN(g33580) );
  NAND2X0 U10729 ( .IN1(test_so62), .IN2(n10023), .QN(n10619) );
  NAND2X0 U10730 ( .IN1(n10620), .IN2(g2259), .QN(n10618) );
  NAND2X0 U10731 ( .IN1(n10621), .IN2(n10622), .QN(g33579) );
  NAND2X0 U10732 ( .IN1(n10023), .IN2(g2246), .QN(n10622) );
  INVX0 U10733 ( .INP(n10620), .ZN(n10023) );
  NAND2X0 U10734 ( .IN1(n10620), .IN2(g2241), .QN(n10621) );
  NAND2X0 U10735 ( .IN1(n10034), .IN2(n8518), .QN(n10620) );
  NAND3X0 U10736 ( .IN1(n5356), .IN2(n10036), .IN3(n5538), .QN(n10034) );
  NAND3X0 U10737 ( .IN1(n10623), .IN2(n10624), .IN3(n10625), .QN(g33578) );
  NAND2X0 U10738 ( .IN1(n8614), .IN2(g2197), .QN(n10625) );
  NAND2X0 U10739 ( .IN1(n10626), .IN2(g2227), .QN(n10624) );
  NAND2X0 U10740 ( .IN1(n10054), .IN2(n10627), .QN(n10623) );
  NOR2X0 U10741 ( .IN1(n5514), .IN2(n10628), .QN(n10054) );
  NAND3X0 U10742 ( .IN1(n10629), .IN2(n10630), .IN3(n10631), .QN(g33577) );
  NAND2X0 U10743 ( .IN1(n10626), .IN2(g2197), .QN(n10631) );
  NAND2X0 U10744 ( .IN1(n8614), .IN2(g2204), .QN(n10630) );
  NAND4X0 U10745 ( .IN1(n10036), .IN2(g2153), .IN3(n10627), .IN4(n8507), .QN(
        n10629) );
  NAND2X0 U10746 ( .IN1(n10632), .IN2(n10633), .QN(g33576) );
  NAND2X0 U10747 ( .IN1(n10626), .IN2(g2153), .QN(n10633) );
  NOR2X0 U10748 ( .IN1(n10036), .IN2(n8553), .QN(n10626) );
  NAND4X0 U10749 ( .IN1(n5538), .IN2(n10634), .IN3(n10627), .IN4(n8507), .QN(
        n10632) );
  NAND2X0 U10750 ( .IN1(n3115), .IN2(n9641), .QN(n10627) );
  INVX0 U10751 ( .INP(n3165), .ZN(n9641) );
  NAND3X0 U10752 ( .IN1(n5287), .IN2(n5519), .IN3(n3116), .QN(n3165) );
  NAND2X0 U10753 ( .IN1(n5356), .IN2(n10048), .QN(n10634) );
  NAND2X0 U10754 ( .IN1(n5514), .IN2(n10036), .QN(n10048) );
  INVX0 U10755 ( .INP(n10628), .ZN(n10036) );
  NOR2X0 U10756 ( .IN1(n10043), .IN2(n3160), .QN(n10628) );
  AND2X1 U10757 ( .IN1(n10635), .IN2(g17320), .Q(n3160) );
  NAND2X0 U10758 ( .IN1(n10525), .IN2(n10636), .QN(n10635) );
  NOR4X0 U10759 ( .IN1(n8203), .IN2(n7839), .IN3(g1559), .IN4(n10637), .QN(
        n10525) );
  NAND3X0 U10760 ( .IN1(n5768), .IN2(n5546), .IN3(n8154), .QN(n10637) );
  NAND3X0 U10761 ( .IN1(n10638), .IN2(n10072), .IN3(n10071), .QN(n10043) );
  NAND2X0 U10762 ( .IN1(n2549), .IN2(g1478), .QN(n10071) );
  NAND2X0 U10763 ( .IN1(n10359), .IN2(n10639), .QN(n10072) );
  NAND3X0 U10764 ( .IN1(n9225), .IN2(g691), .IN3(n5595), .QN(n10639) );
  NAND3X0 U10765 ( .IN1(n5377), .IN2(g2689), .IN3(n5308), .QN(n10638) );
  NAND4X0 U10766 ( .IN1(n10640), .IN2(n3180), .IN3(n10641), .IN4(n10642), .QN(
        g33575) );
  NAND2X0 U10767 ( .IN1(n8614), .IN2(g1996), .QN(n10642) );
  NAND4X0 U10768 ( .IN1(n10643), .IN2(n10644), .IN3(n10645), .IN4(n8507), .QN(
        n10641) );
  INVX0 U10769 ( .INP(n10646), .ZN(n10645) );
  NAND3X0 U10770 ( .IN1(g2070), .IN2(g112), .IN3(n5505), .QN(n10644) );
  NAND4X0 U10771 ( .IN1(n5505), .IN2(n10647), .IN3(n10531), .IN4(g2070), .QN(
        n3180) );
  INVX0 U10772 ( .INP(n10648), .ZN(n10647) );
  NAND2X0 U10773 ( .IN1(n10649), .IN2(g2047), .QN(n10640) );
  NAND2X0 U10774 ( .IN1(n10609), .IN2(n10650), .QN(n10649) );
  NAND2X0 U10775 ( .IN1(n10648), .IN2(n8518), .QN(n10650) );
  NAND2X0 U10776 ( .IN1(n10643), .IN2(n9651), .QN(n10648) );
  NAND3X0 U10777 ( .IN1(n10651), .IN2(n10652), .IN3(n10653), .QN(g33574) );
  NAND2X0 U10778 ( .IN1(n10078), .IN2(g2116), .QN(n10653) );
  NAND3X0 U10779 ( .IN1(n5463), .IN2(n10077), .IN3(n8484), .QN(n10652) );
  NAND2X0 U10780 ( .IN1(n8614), .IN2(g2112), .QN(n10651) );
  NAND3X0 U10781 ( .IN1(n10654), .IN2(n10655), .IN3(n10656), .QN(g33573) );
  NAND2X0 U10782 ( .IN1(n10078), .IN2(g2112), .QN(n10656) );
  NAND2X0 U10783 ( .IN1(n10657), .IN2(g2108), .QN(n10655) );
  NAND2X0 U10784 ( .IN1(n10658), .IN2(n8518), .QN(n10657) );
  NAND2X0 U10785 ( .IN1(n10077), .IN2(g2102), .QN(n10658) );
  NAND4X0 U10786 ( .IN1(n10077), .IN2(n8506), .IN3(n5666), .IN4(n5452), .QN(
        n10654) );
  INVX0 U10787 ( .INP(n10089), .ZN(n10077) );
  NAND2X0 U10788 ( .IN1(n10659), .IN2(n10660), .QN(g33572) );
  NAND2X0 U10789 ( .IN1(n10078), .IN2(g2108), .QN(n10660) );
  NAND2X0 U10790 ( .IN1(n10661), .IN2(g2102), .QN(n10659) );
  NAND2X0 U10791 ( .IN1(n10662), .IN2(n10663), .QN(g33571) );
  NAND2X0 U10792 ( .IN1(n10078), .IN2(g2089), .QN(n10663) );
  INVX0 U10793 ( .INP(n10661), .ZN(n10078) );
  NAND2X0 U10794 ( .IN1(n10661), .IN2(g2084), .QN(n10662) );
  NAND2X0 U10795 ( .IN1(n10089), .IN2(n8518), .QN(n10661) );
  NAND3X0 U10796 ( .IN1(n5355), .IN2(n10091), .IN3(n5535), .QN(n10089) );
  NAND3X0 U10797 ( .IN1(n10664), .IN2(n10665), .IN3(n10666), .QN(g33570) );
  NAND2X0 U10798 ( .IN1(n8614), .IN2(g2040), .QN(n10666) );
  NAND2X0 U10799 ( .IN1(n10667), .IN2(g2070), .QN(n10665) );
  NAND2X0 U10800 ( .IN1(n10109), .IN2(n10646), .QN(n10664) );
  NOR2X0 U10801 ( .IN1(n5505), .IN2(n10668), .QN(n10109) );
  NAND3X0 U10802 ( .IN1(n10669), .IN2(n10670), .IN3(n10671), .QN(g33569) );
  NAND2X0 U10803 ( .IN1(n10667), .IN2(g2040), .QN(n10671) );
  NAND2X0 U10804 ( .IN1(n8614), .IN2(g2047), .QN(n10670) );
  NAND4X0 U10805 ( .IN1(n10091), .IN2(g1996), .IN3(n10646), .IN4(n8507), .QN(
        n10669) );
  NAND2X0 U10806 ( .IN1(n10672), .IN2(n10673), .QN(g33568) );
  NAND2X0 U10807 ( .IN1(n10667), .IN2(g1996), .QN(n10673) );
  NOR2X0 U10808 ( .IN1(n10091), .IN2(n8553), .QN(n10667) );
  NAND4X0 U10809 ( .IN1(n5535), .IN2(n10674), .IN3(n10646), .IN4(n8507), .QN(
        n10672) );
  NAND2X0 U10810 ( .IN1(n3115), .IN2(n9651), .QN(n10646) );
  AND3X1 U10811 ( .IN1(n5519), .IN2(g518), .IN3(n3195), .Q(n9651) );
  NAND2X0 U10812 ( .IN1(n5355), .IN2(n10103), .QN(n10674) );
  NAND2X0 U10813 ( .IN1(n5505), .IN2(n10091), .QN(n10103) );
  INVX0 U10814 ( .INP(n10668), .ZN(n10091) );
  NOR2X0 U10815 ( .IN1(n10098), .IN2(n10643), .QN(n10668) );
  AND2X1 U10816 ( .IN1(g1087), .IN2(n10675), .Q(n10643) );
  NAND3X0 U10817 ( .IN1(n5363), .IN2(n10676), .IN3(n5599), .QN(n10675) );
  NAND3X0 U10818 ( .IN1(n10677), .IN2(n10294), .IN3(n10127), .QN(n10098) );
  NAND2X0 U10819 ( .IN1(n5286), .IN2(g956), .QN(n10127) );
  NAND3X0 U10820 ( .IN1(g2145), .IN2(g2130), .IN3(g2138), .QN(n10677) );
  NAND3X0 U10821 ( .IN1(n10678), .IN2(n10679), .IN3(n10680), .QN(g33567) );
  NAND2X0 U10822 ( .IN1(test_so8), .IN2(n8552), .QN(n10680) );
  NAND2X0 U10823 ( .IN1(n10681), .IN2(n10682), .QN(n10679) );
  NAND2X0 U10824 ( .IN1(n10683), .IN2(n10684), .QN(n10682) );
  NAND3X0 U10825 ( .IN1(n10158), .IN2(n8481), .IN3(n10685), .QN(n10684) );
  NAND2X0 U10826 ( .IN1(n7866), .IN2(n10686), .QN(n10683) );
  NAND2X0 U10827 ( .IN1(n10687), .IN2(n10688), .QN(n10686) );
  NAND3X0 U10828 ( .IN1(n9643), .IN2(n10495), .IN3(n9642), .QN(n10688) );
  INVX0 U10829 ( .INP(n10158), .ZN(n9643) );
  NAND2X0 U10830 ( .IN1(n5503), .IN2(g1936), .QN(n10158) );
  NAND2X0 U10831 ( .IN1(n10685), .IN2(n8518), .QN(n10687) );
  INVX0 U10832 ( .INP(n10689), .ZN(n10685) );
  NAND2X0 U10833 ( .IN1(n10690), .IN2(g1913), .QN(n10678) );
  NAND2X0 U10834 ( .IN1(n10609), .IN2(n10691), .QN(n10690) );
  NAND2X0 U10835 ( .IN1(n10692), .IN2(n8518), .QN(n10691) );
  NAND2X0 U10836 ( .IN1(n10681), .IN2(n9642), .QN(n10692) );
  NAND3X0 U10837 ( .IN1(n10693), .IN2(n10694), .IN3(n10695), .QN(g33566) );
  NAND2X0 U10838 ( .IN1(n10133), .IN2(g1982), .QN(n10695) );
  NAND3X0 U10839 ( .IN1(n5462), .IN2(n10132), .IN3(n8485), .QN(n10694) );
  NAND2X0 U10840 ( .IN1(n8657), .IN2(g1978), .QN(n10693) );
  NAND3X0 U10841 ( .IN1(n10696), .IN2(n10697), .IN3(n10698), .QN(g33565) );
  NAND2X0 U10842 ( .IN1(n10133), .IN2(g1978), .QN(n10698) );
  NAND2X0 U10843 ( .IN1(n10699), .IN2(g1974), .QN(n10697) );
  NAND2X0 U10844 ( .IN1(n10700), .IN2(n8518), .QN(n10699) );
  NAND2X0 U10845 ( .IN1(n10132), .IN2(g1968), .QN(n10700) );
  NAND4X0 U10846 ( .IN1(n10132), .IN2(n8506), .IN3(n5664), .IN4(n5450), .QN(
        n10696) );
  INVX0 U10847 ( .INP(n10144), .ZN(n10132) );
  NAND2X0 U10848 ( .IN1(n10701), .IN2(n10702), .QN(g33564) );
  NAND2X0 U10849 ( .IN1(n10133), .IN2(g1974), .QN(n10702) );
  NAND2X0 U10850 ( .IN1(n10703), .IN2(g1968), .QN(n10701) );
  NAND2X0 U10851 ( .IN1(n10704), .IN2(n10705), .QN(g33563) );
  NAND2X0 U10852 ( .IN1(n10133), .IN2(g1955), .QN(n10705) );
  INVX0 U10853 ( .INP(n10703), .ZN(n10133) );
  NAND2X0 U10854 ( .IN1(n10703), .IN2(g1950), .QN(n10704) );
  NAND2X0 U10855 ( .IN1(n10144), .IN2(n8518), .QN(n10703) );
  NAND3X0 U10856 ( .IN1(n10146), .IN2(n8205), .IN3(n5534), .QN(n10144) );
  NAND3X0 U10857 ( .IN1(n10706), .IN2(n10707), .IN3(n10708), .QN(g33562) );
  NAND2X0 U10858 ( .IN1(n8647), .IN2(g1906), .QN(n10708) );
  NAND2X0 U10859 ( .IN1(n10709), .IN2(g1936), .QN(n10707) );
  NAND2X0 U10860 ( .IN1(n10165), .IN2(n10689), .QN(n10706) );
  NOR2X0 U10861 ( .IN1(n5503), .IN2(n10159), .QN(n10165) );
  NAND3X0 U10862 ( .IN1(n10710), .IN2(n10711), .IN3(n10712), .QN(g33561) );
  NAND2X0 U10863 ( .IN1(n10709), .IN2(g1906), .QN(n10712) );
  NAND2X0 U10864 ( .IN1(n8648), .IN2(g1913), .QN(n10711) );
  NAND3X0 U10865 ( .IN1(n10171), .IN2(n10689), .IN3(n8484), .QN(n10710) );
  NOR2X0 U10866 ( .IN1(n8205), .IN2(n10159), .QN(n10171) );
  NAND2X0 U10867 ( .IN1(n10713), .IN2(n10714), .QN(g33560) );
  NAND4X0 U10868 ( .IN1(n5534), .IN2(n10715), .IN3(n10689), .IN4(n8507), .QN(
        n10714) );
  NAND2X0 U10869 ( .IN1(n3115), .IN2(n9642), .QN(n10689) );
  INVX0 U10870 ( .INP(n9657), .ZN(n9642) );
  NAND3X0 U10871 ( .IN1(g518), .IN2(g504), .IN3(n3195), .QN(n9657) );
  NAND2X0 U10872 ( .IN1(n8205), .IN2(n10716), .QN(n10715) );
  NAND2X0 U10873 ( .IN1(n5503), .IN2(n10146), .QN(n10716) );
  NAND2X0 U10874 ( .IN1(n10709), .IN2(test_so8), .QN(n10713) );
  NOR2X0 U10875 ( .IN1(n10146), .IN2(n8553), .QN(n10709) );
  INVX0 U10876 ( .INP(n10159), .ZN(n10146) );
  NOR2X0 U10877 ( .IN1(n10153), .IN2(n10681), .QN(n10159) );
  AND2X1 U10878 ( .IN1(n10717), .IN2(g17400), .Q(n10681) );
  NAND2X0 U10879 ( .IN1(n10718), .IN2(n10676), .QN(n10717) );
  NAND3X0 U10880 ( .IN1(n10719), .IN2(n10294), .IN3(n10183), .QN(n10153) );
  NAND2X0 U10881 ( .IN1(n5286), .IN2(g1129), .QN(n10183) );
  NAND3X0 U10882 ( .IN1(g2138), .IN2(g2130), .IN3(n5307), .QN(n10719) );
  NAND3X0 U10883 ( .IN1(n10720), .IN2(n10721), .IN3(n10722), .QN(g33559) );
  NAND2X0 U10884 ( .IN1(n8653), .IN2(g1728), .QN(n10722) );
  NAND3X0 U10885 ( .IN1(n10723), .IN2(n10724), .IN3(n10725), .QN(n10721) );
  NAND3X0 U10886 ( .IN1(g1802), .IN2(g112), .IN3(n5504), .QN(n10724) );
  NAND2X0 U10887 ( .IN1(n10726), .IN2(n10727), .QN(n10723) );
  NAND3X0 U10888 ( .IN1(n10495), .IN2(g1802), .IN3(n5504), .QN(n10727) );
  NAND2X0 U10889 ( .IN1(n3115), .IN2(n8518), .QN(n10726) );
  NAND2X0 U10890 ( .IN1(n10728), .IN2(g1779), .QN(n10720) );
  NAND2X0 U10891 ( .IN1(n10609), .IN2(n10729), .QN(n10728) );
  OR2X1 U10892 ( .IN1(n10725), .IN2(n8546), .Q(n10729) );
  NOR2X0 U10893 ( .IN1(n10730), .IN2(n9655), .QN(n10725) );
  NAND3X0 U10894 ( .IN1(n10731), .IN2(n10732), .IN3(n10733), .QN(g33558) );
  NAND2X0 U10895 ( .IN1(n10190), .IN2(g1848), .QN(n10733) );
  NAND3X0 U10896 ( .IN1(n5464), .IN2(n10189), .IN3(n8484), .QN(n10732) );
  NAND2X0 U10897 ( .IN1(n8654), .IN2(g1844), .QN(n10731) );
  NAND3X0 U10898 ( .IN1(n10734), .IN2(n10735), .IN3(n10736), .QN(g33557) );
  NAND2X0 U10899 ( .IN1(n10190), .IN2(g1844), .QN(n10736) );
  NAND2X0 U10900 ( .IN1(n10737), .IN2(g1840), .QN(n10735) );
  NAND2X0 U10901 ( .IN1(n10738), .IN2(n8518), .QN(n10737) );
  NAND2X0 U10902 ( .IN1(n10189), .IN2(g1834), .QN(n10738) );
  NAND4X0 U10903 ( .IN1(n10189), .IN2(n8506), .IN3(n5665), .IN4(n5451), .QN(
        n10734) );
  INVX0 U10904 ( .INP(n10201), .ZN(n10189) );
  NAND2X0 U10905 ( .IN1(n10739), .IN2(n10740), .QN(g33556) );
  NAND2X0 U10906 ( .IN1(n10190), .IN2(g1840), .QN(n10740) );
  NAND2X0 U10907 ( .IN1(n10741), .IN2(g1834), .QN(n10739) );
  NAND2X0 U10908 ( .IN1(n10742), .IN2(n10743), .QN(g33555) );
  NAND2X0 U10909 ( .IN1(n10190), .IN2(g1821), .QN(n10743) );
  INVX0 U10910 ( .INP(n10741), .ZN(n10190) );
  NAND2X0 U10911 ( .IN1(n10741), .IN2(g1816), .QN(n10742) );
  NAND2X0 U10912 ( .IN1(n10201), .IN2(n8518), .QN(n10741) );
  NAND3X0 U10913 ( .IN1(n5352), .IN2(n10203), .IN3(n5536), .QN(n10201) );
  NAND3X0 U10914 ( .IN1(n10744), .IN2(n10745), .IN3(n10746), .QN(g33554) );
  NAND2X0 U10915 ( .IN1(n8651), .IN2(g1772), .QN(n10746) );
  NAND2X0 U10916 ( .IN1(n10747), .IN2(g1802), .QN(n10745) );
  NAND2X0 U10917 ( .IN1(n10221), .IN2(n10748), .QN(n10744) );
  AND2X1 U10918 ( .IN1(g1772), .IN2(n10203), .Q(n10221) );
  NAND3X0 U10919 ( .IN1(n10749), .IN2(n10750), .IN3(n10751), .QN(g33553) );
  NAND2X0 U10920 ( .IN1(n10747), .IN2(g1772), .QN(n10751) );
  NAND2X0 U10921 ( .IN1(n8652), .IN2(g1779), .QN(n10750) );
  NAND4X0 U10922 ( .IN1(n10203), .IN2(g1728), .IN3(n10748), .IN4(n8508), .QN(
        n10749) );
  NAND2X0 U10923 ( .IN1(n10752), .IN2(n10753), .QN(g33552) );
  NAND2X0 U10924 ( .IN1(n10747), .IN2(g1728), .QN(n10753) );
  NOR2X0 U10925 ( .IN1(n10203), .IN2(n8555), .QN(n10747) );
  NAND4X0 U10926 ( .IN1(n5536), .IN2(n10754), .IN3(n10748), .IN4(n8507), .QN(
        n10752) );
  NAND2X0 U10927 ( .IN1(n3115), .IN2(n9652), .QN(n10748) );
  INVX0 U10928 ( .INP(n9655), .ZN(n9652) );
  NAND3X0 U10929 ( .IN1(n5287), .IN2(g504), .IN3(n3195), .QN(n9655) );
  NAND2X0 U10930 ( .IN1(n5352), .IN2(n10215), .QN(n10754) );
  NAND2X0 U10931 ( .IN1(n5504), .IN2(n10203), .QN(n10215) );
  NAND2X0 U10932 ( .IN1(n10208), .IN2(n10730), .QN(n10203) );
  NAND2X0 U10933 ( .IN1(test_so44), .IN2(n10755), .QN(n10730) );
  NAND2X0 U10934 ( .IN1(n10756), .IN2(n10676), .QN(n10755) );
  INVX0 U10935 ( .INP(n10210), .ZN(n10208) );
  NAND3X0 U10936 ( .IN1(n10757), .IN2(n10294), .IN3(n10238), .QN(n10210) );
  NAND2X0 U10937 ( .IN1(n5286), .IN2(g1105), .QN(n10238) );
  NAND3X0 U10938 ( .IN1(g2145), .IN2(g2130), .IN3(n5275), .QN(n10757) );
  NAND3X0 U10939 ( .IN1(n10758), .IN2(n10759), .IN3(n10760), .QN(g33551) );
  NAND2X0 U10940 ( .IN1(n8540), .IN2(g1592), .QN(n10760) );
  NAND3X0 U10941 ( .IN1(n9646), .IN2(n10761), .IN3(g33533), .QN(n10759) );
  NAND2X0 U10942 ( .IN1(n10762), .IN2(n10763), .QN(n10761) );
  NAND3X0 U10943 ( .IN1(n10764), .IN2(n8483), .IN3(n3115), .QN(n10763) );
  NAND2X0 U10944 ( .IN1(g31862), .IN2(g112), .QN(n10764) );
  NAND2X0 U10945 ( .IN1(g31862), .IN2(n10531), .QN(n10762) );
  NOR2X0 U10946 ( .IN1(g112), .IN2(n9539), .QN(n10531) );
  NAND2X0 U10947 ( .IN1(test_so75), .IN2(n10765), .QN(n10758) );
  NAND2X0 U10948 ( .IN1(n10609), .IN2(n10766), .QN(n10765) );
  NAND2X0 U10949 ( .IN1(n10767), .IN2(n8518), .QN(n10766) );
  NAND2X0 U10950 ( .IN1(g33533), .IN2(n9646), .QN(n10767) );
  NAND3X0 U10951 ( .IN1(n10768), .IN2(n10769), .IN3(n10770), .QN(g33550) );
  NAND2X0 U10952 ( .IN1(n10244), .IN2(g1714), .QN(n10770) );
  NAND3X0 U10953 ( .IN1(n5460), .IN2(n10243), .IN3(n8486), .QN(n10769) );
  NAND2X0 U10954 ( .IN1(n8541), .IN2(g1710), .QN(n10768) );
  NAND3X0 U10955 ( .IN1(n10771), .IN2(n10772), .IN3(n10773), .QN(g33549) );
  NAND2X0 U10956 ( .IN1(n10244), .IN2(g1710), .QN(n10773) );
  NAND2X0 U10957 ( .IN1(test_so15), .IN2(n10774), .QN(n10772) );
  NAND2X0 U10958 ( .IN1(n10775), .IN2(n8518), .QN(n10774) );
  NAND2X0 U10959 ( .IN1(n10243), .IN2(g1700), .QN(n10775) );
  INVX0 U10960 ( .INP(n10255), .ZN(n10243) );
  OR4X1 U10961 ( .IN1(n10255), .IN2(n8544), .IN3(g1700), .IN4(test_so15), .Q(
        n10771) );
  NAND2X0 U10962 ( .IN1(n10776), .IN2(n10777), .QN(g33548) );
  NAND2X0 U10963 ( .IN1(test_so15), .IN2(n10244), .QN(n10777) );
  NAND2X0 U10964 ( .IN1(n10778), .IN2(g1700), .QN(n10776) );
  NAND2X0 U10965 ( .IN1(n10779), .IN2(n10780), .QN(g33547) );
  NAND2X0 U10966 ( .IN1(n10244), .IN2(g1687), .QN(n10780) );
  INVX0 U10967 ( .INP(n10778), .ZN(n10244) );
  NAND2X0 U10968 ( .IN1(n10778), .IN2(g1682), .QN(n10779) );
  NAND2X0 U10969 ( .IN1(n10255), .IN2(n8518), .QN(n10778) );
  NAND3X0 U10970 ( .IN1(n5362), .IN2(n10257), .IN3(n5598), .QN(n10255) );
  NAND3X0 U10971 ( .IN1(n10781), .IN2(n10782), .IN3(n10783), .QN(g33546) );
  NAND2X0 U10972 ( .IN1(n8628), .IN2(g1636), .QN(n10783) );
  NAND2X0 U10973 ( .IN1(n10784), .IN2(g1668), .QN(n10782) );
  NAND2X0 U10974 ( .IN1(n10275), .IN2(n10785), .QN(n10781) );
  NOR2X0 U10975 ( .IN1(n5549), .IN2(n10786), .QN(n10275) );
  NAND3X0 U10976 ( .IN1(n10787), .IN2(n10788), .IN3(n10789), .QN(g33545) );
  NAND2X0 U10977 ( .IN1(n10784), .IN2(g1636), .QN(n10789) );
  NAND2X0 U10978 ( .IN1(test_so75), .IN2(n8659), .QN(n10788) );
  NAND3X0 U10979 ( .IN1(n10281), .IN2(n10785), .IN3(n8486), .QN(n10787) );
  NOR2X0 U10980 ( .IN1(n5362), .IN2(n10786), .QN(n10281) );
  NAND2X0 U10981 ( .IN1(n10790), .IN2(n10791), .QN(g33544) );
  NAND2X0 U10982 ( .IN1(n10784), .IN2(g1592), .QN(n10791) );
  NOR2X0 U10983 ( .IN1(n10257), .IN2(n8554), .QN(n10784) );
  NAND4X0 U10984 ( .IN1(n10257), .IN2(n8505), .IN3(n10785), .IN4(n10792), .QN(
        n10790) );
  AND2X1 U10985 ( .IN1(n10793), .IN2(n5598), .Q(n10792) );
  NAND2X0 U10986 ( .IN1(n3115), .IN2(n9646), .QN(n10785) );
  INVX0 U10987 ( .INP(n9656), .ZN(n9646) );
  NAND3X0 U10988 ( .IN1(n5287), .IN2(n5519), .IN3(n3195), .QN(n9656) );
  INVX0 U10989 ( .INP(n10786), .ZN(n10257) );
  NOR2X0 U10990 ( .IN1(n10264), .IN2(g33533), .QN(n10786) );
  NAND3X0 U10991 ( .IN1(n10794), .IN2(n10294), .IN3(n10293), .QN(n10264) );
  NAND2X0 U10992 ( .IN1(n5286), .IN2(g1135), .QN(n10293) );
  NAND2X0 U10993 ( .IN1(n10359), .IN2(n10795), .QN(n10294) );
  NAND3X0 U10994 ( .IN1(n9224), .IN2(g691), .IN3(n5595), .QN(n10795) );
  INVX0 U10995 ( .INP(g134), .ZN(n10359) );
  NAND3X0 U10996 ( .IN1(n5307), .IN2(g2130), .IN3(n5275), .QN(n10794) );
  NAND2X0 U10997 ( .IN1(n10796), .IN2(n10797), .QN(g33543) );
  NAND3X0 U10998 ( .IN1(n8504), .IN2(g1379), .IN3(n10798), .QN(n10797) );
  NAND2X0 U10999 ( .IN1(n10799), .IN2(n10800), .QN(n10798) );
  NAND2X0 U11000 ( .IN1(n7849), .IN2(n10801), .QN(n10800) );
  NAND2X0 U11001 ( .IN1(n10802), .IN2(g1373), .QN(n10796) );
  NAND2X0 U11002 ( .IN1(n10803), .IN2(n8518), .QN(n10802) );
  NAND3X0 U11003 ( .IN1(n10799), .IN2(n10801), .IN3(n7778), .QN(n10803) );
  NAND3X0 U11004 ( .IN1(n10804), .IN2(n10805), .IN3(n10806), .QN(g33542) );
  NAND2X0 U11005 ( .IN1(n8650), .IN2(g1270), .QN(n10806) );
  OR3X1 U11006 ( .IN1(n10807), .IN2(n10808), .IN3(n5730), .Q(n10805) );
  NAND2X0 U11007 ( .IN1(n5730), .IN2(n10808), .QN(n10804) );
  NAND2X0 U11008 ( .IN1(n10809), .IN2(n10810), .QN(g33541) );
  NAND3X0 U11009 ( .IN1(n8504), .IN2(g1036), .IN3(n10811), .QN(n10810) );
  NAND2X0 U11010 ( .IN1(n10812), .IN2(n10813), .QN(n10811) );
  NAND2X0 U11011 ( .IN1(n7851), .IN2(n10814), .QN(n10813) );
  NAND2X0 U11012 ( .IN1(n10815), .IN2(g1030), .QN(n10809) );
  NAND2X0 U11013 ( .IN1(n10816), .IN2(n8518), .QN(n10815) );
  NAND3X0 U11014 ( .IN1(n10812), .IN2(n10814), .IN3(n7779), .QN(n10816) );
  NAND3X0 U11015 ( .IN1(n10817), .IN2(n10818), .IN3(n10819), .QN(g33540) );
  NAND2X0 U11016 ( .IN1(n8651), .IN2(g925), .QN(n10819) );
  OR3X1 U11017 ( .IN1(n10820), .IN2(n10821), .IN3(n5731), .Q(n10818) );
  NAND2X0 U11018 ( .IN1(n5731), .IN2(n10821), .QN(n10817) );
  NAND3X0 U11019 ( .IN1(n10822), .IN2(n10823), .IN3(n10824), .QN(g33539) );
  NAND2X0 U11020 ( .IN1(n8651), .IN2(g758), .QN(n10824) );
  NAND3X0 U11021 ( .IN1(n2404), .IN2(n10825), .IN3(g763), .QN(n10823) );
  INVX0 U11022 ( .INP(n2980), .ZN(n10825) );
  NAND2X0 U11023 ( .IN1(n2980), .IN2(n5332), .QN(n10822) );
  NAND3X0 U11024 ( .IN1(n10826), .IN2(n10827), .IN3(n10828), .QN(g33538) );
  NAND2X0 U11025 ( .IN1(n8651), .IN2(g590), .QN(n10828) );
  NAND3X0 U11026 ( .IN1(n2421), .IN2(n10829), .IN3(g595), .QN(n10827) );
  INVX0 U11027 ( .INP(n2982), .ZN(n10829) );
  NAND2X0 U11028 ( .IN1(n2982), .IN2(n5476), .QN(n10826) );
  NAND2X0 U11029 ( .IN1(n10830), .IN2(n10831), .QN(g33537) );
  OR2X1 U11030 ( .IN1(n8476), .IN2(n8184), .Q(n10831) );
  NAND3X0 U11031 ( .IN1(n2707), .IN2(g142), .IN3(n8487), .QN(n10830) );
  NOR2X0 U11032 ( .IN1(n5843), .IN2(n10832), .QN(g33536) );
  NOR2X0 U11033 ( .IN1(n2710), .IN2(n8554), .QN(n10832) );
  NAND3X0 U11034 ( .IN1(n10833), .IN2(n10834), .IN3(n10835), .QN(g33535) );
  NAND2X0 U11035 ( .IN1(n8652), .IN2(g291), .QN(n10835) );
  NAND3X0 U11036 ( .IN1(n8194), .IN2(n10836), .IN3(g294), .QN(n10834) );
  INVX0 U11037 ( .INP(n3276), .ZN(n10836) );
  NAND2X0 U11038 ( .IN1(n3276), .IN2(n5680), .QN(n10833) );
  NAND3X0 U11039 ( .IN1(n10837), .IN2(n10838), .IN3(n10839), .QN(g33534) );
  OR2X1 U11040 ( .IN1(n8479), .IN2(n5676), .Q(n10839) );
  OR3X1 U11041 ( .IN1(n9761), .IN2(n3277), .IN3(n5677), .Q(n10838) );
  NAND2X0 U11042 ( .IN1(n3277), .IN2(n5677), .QN(n10837) );
  AND2X1 U11043 ( .IN1(n10840), .IN2(g17291), .Q(g33533) );
  NAND2X0 U11044 ( .IN1(n10841), .IN2(n10676), .QN(n10840) );
  AND4X1 U11045 ( .IN1(n5547), .IN2(n5442), .IN3(n8156), .IN4(n10842), .Q(
        n10676) );
  NOR3X0 U11046 ( .IN1(n5320), .IN2(test_so76), .IN3(n7840), .QN(n10842) );
  AND3X1 U11047 ( .IN1(n10843), .IN2(n10844), .IN3(n10845), .Q(g33435) );
  NAND2X0 U11048 ( .IN1(n9565), .IN2(g2787), .QN(n10845) );
  NAND3X0 U11049 ( .IN1(n10846), .IN2(n10847), .IN3(n7867), .QN(n10844) );
  NAND2X0 U11050 ( .IN1(n5378), .IN2(g2724), .QN(n10847) );
  NAND2X0 U11051 ( .IN1(n5544), .IN2(n5301), .QN(n10846) );
  NAND2X0 U11052 ( .IN1(n9574), .IN2(g2783), .QN(n10843) );
  AND3X1 U11053 ( .IN1(n10848), .IN2(n10849), .IN3(n10850), .Q(g33079) );
  NAND2X0 U11054 ( .IN1(n9565), .IN2(g2819), .QN(n10850) );
  NAND3X0 U11055 ( .IN1(n10851), .IN2(n10852), .IN3(n7867), .QN(n10849) );
  NAND2X0 U11056 ( .IN1(n5379), .IN2(g2724), .QN(n10852) );
  NAND2X0 U11057 ( .IN1(n5545), .IN2(n5301), .QN(n10851) );
  NAND2X0 U11058 ( .IN1(n9574), .IN2(g2815), .QN(n10848) );
  NOR2X0 U11059 ( .IN1(g2724), .IN2(n7867), .QN(n9574) );
  NAND2X0 U11060 ( .IN1(n10853), .IN2(n10854), .QN(g33070) );
  NAND2X0 U11061 ( .IN1(n10855), .IN2(n10856), .QN(n10854) );
  NAND3X0 U11062 ( .IN1(n10857), .IN2(n10858), .IN3(n10859), .QN(n10855) );
  NAND2X0 U11063 ( .IN1(n8512), .IN2(n10860), .QN(n10859) );
  NAND2X0 U11064 ( .IN1(g25756), .IN2(n5646), .QN(n10857) );
  NAND2X0 U11065 ( .IN1(n8652), .IN2(g6565), .QN(n10853) );
  NAND2X0 U11066 ( .IN1(n10861), .IN2(n10862), .QN(g33069) );
  NAND2X0 U11067 ( .IN1(n10863), .IN2(g6561), .QN(n10862) );
  NAND2X0 U11068 ( .IN1(n10864), .IN2(n8518), .QN(n10863) );
  NAND2X0 U11069 ( .IN1(n5386), .IN2(n10856), .QN(n10864) );
  OR2X1 U11070 ( .IN1(n10865), .IN2(n5386), .Q(n10861) );
  NAND2X0 U11071 ( .IN1(n10866), .IN2(n10867), .QN(g33068) );
  NAND3X0 U11072 ( .IN1(n10856), .IN2(n10868), .IN3(n5646), .QN(n10867) );
  NAND2X0 U11073 ( .IN1(n8652), .IN2(g6555), .QN(n10866) );
  NAND2X0 U11074 ( .IN1(n10869), .IN2(n10870), .QN(g33067) );
  NAND2X0 U11075 ( .IN1(n10871), .IN2(n10856), .QN(n10870) );
  NAND2X0 U11076 ( .IN1(n3407), .IN2(n10872), .QN(n10871) );
  NAND2X0 U11077 ( .IN1(n8512), .IN2(n10873), .QN(n10872) );
  NAND2X0 U11078 ( .IN1(n8653), .IN2(g6549), .QN(n10869) );
  NAND2X0 U11079 ( .IN1(n10874), .IN2(n10875), .QN(g33065) );
  NAND2X0 U11080 ( .IN1(n10876), .IN2(n10877), .QN(n10875) );
  NAND3X0 U11081 ( .IN1(n10878), .IN2(n10879), .IN3(n10880), .QN(n10876) );
  NAND2X0 U11082 ( .IN1(n8512), .IN2(n10881), .QN(n10880) );
  NAND2X0 U11083 ( .IN1(g25742), .IN2(n5651), .QN(n10878) );
  NAND2X0 U11084 ( .IN1(n8653), .IN2(g6219), .QN(n10874) );
  NAND2X0 U11085 ( .IN1(n10882), .IN2(n10883), .QN(g33064) );
  NAND2X0 U11086 ( .IN1(n10884), .IN2(g6215), .QN(n10883) );
  NAND2X0 U11087 ( .IN1(n10885), .IN2(n8518), .QN(n10884) );
  NAND2X0 U11088 ( .IN1(n5385), .IN2(n10877), .QN(n10885) );
  OR2X1 U11089 ( .IN1(n10886), .IN2(n5385), .Q(n10882) );
  NAND2X0 U11090 ( .IN1(n10887), .IN2(n10888), .QN(g33063) );
  NAND3X0 U11091 ( .IN1(n10877), .IN2(n10889), .IN3(n5651), .QN(n10888) );
  NAND2X0 U11092 ( .IN1(n8654), .IN2(g6209), .QN(n10887) );
  NAND2X0 U11093 ( .IN1(n10890), .IN2(n10891), .QN(g33062) );
  NAND2X0 U11094 ( .IN1(n10892), .IN2(n10877), .QN(n10891) );
  NAND2X0 U11095 ( .IN1(n3417), .IN2(n10893), .QN(n10892) );
  NAND2X0 U11096 ( .IN1(n8512), .IN2(n10894), .QN(n10893) );
  NAND2X0 U11097 ( .IN1(n8654), .IN2(g6203), .QN(n10890) );
  NAND2X0 U11098 ( .IN1(n10895), .IN2(n10896), .QN(g33060) );
  NAND2X0 U11099 ( .IN1(n10897), .IN2(n10898), .QN(n10896) );
  NAND3X0 U11100 ( .IN1(n10899), .IN2(n10900), .IN3(n10901), .QN(n10897) );
  NAND2X0 U11101 ( .IN1(n8512), .IN2(n10902), .QN(n10901) );
  NAND2X0 U11102 ( .IN1(g25728), .IN2(n5649), .QN(n10899) );
  NAND2X0 U11103 ( .IN1(n8655), .IN2(g5873), .QN(n10895) );
  NAND2X0 U11104 ( .IN1(n10903), .IN2(n10904), .QN(g33059) );
  NAND2X0 U11105 ( .IN1(n10905), .IN2(g5869), .QN(n10904) );
  NAND2X0 U11106 ( .IN1(n10906), .IN2(n8517), .QN(n10905) );
  NAND2X0 U11107 ( .IN1(n5388), .IN2(n10898), .QN(n10906) );
  OR2X1 U11108 ( .IN1(n10907), .IN2(n5388), .Q(n10903) );
  NAND2X0 U11109 ( .IN1(n10908), .IN2(n10909), .QN(g33058) );
  NAND3X0 U11110 ( .IN1(n10898), .IN2(n10910), .IN3(n5649), .QN(n10909) );
  NAND2X0 U11111 ( .IN1(n8655), .IN2(g5863), .QN(n10908) );
  NAND2X0 U11112 ( .IN1(n10911), .IN2(n10912), .QN(g33057) );
  NAND2X0 U11113 ( .IN1(n10913), .IN2(n10898), .QN(n10912) );
  NAND2X0 U11114 ( .IN1(n3427), .IN2(n10914), .QN(n10913) );
  NAND2X0 U11115 ( .IN1(n8512), .IN2(n10915), .QN(n10914) );
  NAND2X0 U11116 ( .IN1(n8656), .IN2(g5857), .QN(n10911) );
  NAND2X0 U11117 ( .IN1(n10916), .IN2(n10917), .QN(g33055) );
  NAND2X0 U11118 ( .IN1(n10918), .IN2(n10919), .QN(n10917) );
  NAND3X0 U11119 ( .IN1(n10920), .IN2(n10921), .IN3(n10922), .QN(n10918) );
  NAND2X0 U11120 ( .IN1(n8512), .IN2(n10923), .QN(n10922) );
  NAND2X0 U11121 ( .IN1(g25714), .IN2(n5647), .QN(n10920) );
  NAND2X0 U11122 ( .IN1(n8656), .IN2(g5527), .QN(n10916) );
  NAND2X0 U11123 ( .IN1(n10924), .IN2(n10925), .QN(g33054) );
  NAND2X0 U11124 ( .IN1(n10926), .IN2(g5523), .QN(n10925) );
  NAND2X0 U11125 ( .IN1(n10927), .IN2(n8517), .QN(n10926) );
  NAND2X0 U11126 ( .IN1(n5389), .IN2(n10919), .QN(n10927) );
  OR2X1 U11127 ( .IN1(n10928), .IN2(n5389), .Q(n10924) );
  NAND2X0 U11128 ( .IN1(n10929), .IN2(n10930), .QN(g33053) );
  NAND3X0 U11129 ( .IN1(n10919), .IN2(n10931), .IN3(n5647), .QN(n10930) );
  NAND2X0 U11130 ( .IN1(n8657), .IN2(g5517), .QN(n10929) );
  NAND2X0 U11131 ( .IN1(n10932), .IN2(n10933), .QN(g33052) );
  NAND2X0 U11132 ( .IN1(n10934), .IN2(n10919), .QN(n10933) );
  NAND2X0 U11133 ( .IN1(n3437), .IN2(n10935), .QN(n10934) );
  NAND2X0 U11134 ( .IN1(n8512), .IN2(n10936), .QN(n10935) );
  NAND2X0 U11135 ( .IN1(n8656), .IN2(g5511), .QN(n10932) );
  NAND2X0 U11136 ( .IN1(n10937), .IN2(n10938), .QN(g33050) );
  NAND2X0 U11137 ( .IN1(n10939), .IN2(n10940), .QN(n10938) );
  NAND3X0 U11138 ( .IN1(n10941), .IN2(n10942), .IN3(n10943), .QN(n10939) );
  NAND2X0 U11139 ( .IN1(n8512), .IN2(n10944), .QN(n10943) );
  NAND2X0 U11140 ( .IN1(g25700), .IN2(n5650), .QN(n10941) );
  NAND2X0 U11141 ( .IN1(n8656), .IN2(g5180), .QN(n10937) );
  NAND2X0 U11142 ( .IN1(n10945), .IN2(n10946), .QN(g33049) );
  NAND2X0 U11143 ( .IN1(n10947), .IN2(g5176), .QN(n10946) );
  NAND2X0 U11144 ( .IN1(n10948), .IN2(n8517), .QN(n10947) );
  NAND2X0 U11145 ( .IN1(n5384), .IN2(n10940), .QN(n10948) );
  OR2X1 U11146 ( .IN1(n10949), .IN2(n5384), .Q(n10945) );
  NAND2X0 U11147 ( .IN1(n10950), .IN2(n10951), .QN(g33048) );
  NAND3X0 U11148 ( .IN1(n10940), .IN2(n10952), .IN3(n5650), .QN(n10951) );
  NAND2X0 U11149 ( .IN1(n8657), .IN2(g5170), .QN(n10950) );
  NAND2X0 U11150 ( .IN1(n10953), .IN2(n10954), .QN(g33047) );
  NAND2X0 U11151 ( .IN1(n10955), .IN2(n10940), .QN(n10954) );
  NAND2X0 U11152 ( .IN1(n3447), .IN2(n10956), .QN(n10955) );
  NAND2X0 U11153 ( .IN1(n8512), .IN2(n10957), .QN(n10956) );
  NAND2X0 U11154 ( .IN1(n8658), .IN2(g5164), .QN(n10953) );
  NAND3X0 U11155 ( .IN1(n10958), .IN2(n10959), .IN3(n10960), .QN(g33046) );
  NAND2X0 U11156 ( .IN1(n8657), .IN2(g5052), .QN(n10960) );
  NAND2X0 U11157 ( .IN1(n5615), .IN2(n10961), .QN(n10959) );
  NAND2X0 U11158 ( .IN1(n10962), .IN2(n10963), .QN(n10961) );
  NAND3X0 U11159 ( .IN1(n10964), .IN2(n10963), .IN3(g5057), .QN(n10958) );
  NAND2X0 U11160 ( .IN1(n10965), .IN2(g5052), .QN(n10963) );
  NAND3X0 U11161 ( .IN1(n10966), .IN2(n10967), .IN3(n10968), .QN(g33045) );
  NAND2X0 U11162 ( .IN1(n10433), .IN2(g4567), .QN(n10968) );
  NAND3X0 U11163 ( .IN1(n10967), .IN2(n9836), .IN3(n10969), .QN(g33044) );
  NAND2X0 U11164 ( .IN1(test_so93), .IN2(n10433), .QN(n10969) );
  NAND3X0 U11165 ( .IN1(n10970), .IN2(n10431), .IN3(n10971), .QN(g33043) );
  NAND2X0 U11166 ( .IN1(test_so16), .IN2(n10433), .QN(n10971) );
  NAND3X0 U11167 ( .IN1(n10970), .IN2(n10967), .IN3(n10972), .QN(g33042) );
  NAND2X0 U11168 ( .IN1(n10433), .IN2(g4540), .QN(n10972) );
  NAND2X0 U11169 ( .IN1(n10973), .IN2(g4578), .QN(n10967) );
  NAND3X0 U11170 ( .IN1(n10966), .IN2(n10431), .IN3(n10974), .QN(g33041) );
  NAND2X0 U11171 ( .IN1(test_so56), .IN2(n10433), .QN(n10974) );
  NAND3X0 U11172 ( .IN1(n10975), .IN2(n9836), .IN3(n10976), .QN(g33040) );
  NAND2X0 U11173 ( .IN1(n10433), .IN2(g4504), .QN(n10976) );
  NAND2X0 U11174 ( .IN1(n10973), .IN2(n9842), .QN(n9836) );
  INVX0 U11175 ( .INP(n9172), .ZN(n9842) );
  NOR2X0 U11176 ( .IN1(g73), .IN2(g72), .QN(n9172) );
  NAND3X0 U11177 ( .IN1(n10966), .IN2(n10436), .IN3(n10977), .QN(g33039) );
  NAND2X0 U11178 ( .IN1(n10433), .IN2(g4501), .QN(n10977) );
  NAND3X0 U11179 ( .IN1(n10966), .IN2(n10975), .IN3(n10978), .QN(g33038) );
  NAND2X0 U11180 ( .IN1(n10433), .IN2(g4498), .QN(n10978) );
  NAND2X0 U11181 ( .IN1(n10973), .IN2(n10979), .QN(n10966) );
  OR2X1 U11182 ( .IN1(n10321), .IN2(g73), .Q(n10979) );
  INVX0 U11183 ( .INP(g72), .ZN(n10321) );
  NAND3X0 U11184 ( .IN1(n10970), .IN2(n10436), .IN3(n10980), .QN(g33037) );
  NAND2X0 U11185 ( .IN1(n10433), .IN2(g4495), .QN(n10980) );
  NAND3X0 U11186 ( .IN1(n10970), .IN2(n10975), .IN3(n10981), .QN(g33036) );
  NAND2X0 U11187 ( .IN1(n10433), .IN2(g4480), .QN(n10981) );
  OR2X1 U11188 ( .IN1(n10433), .IN2(n7770), .Q(n10975) );
  INVX0 U11189 ( .INP(n10973), .ZN(n10433) );
  NAND2X0 U11190 ( .IN1(n10973), .IN2(n10982), .QN(n10970) );
  NAND2X0 U11191 ( .IN1(g73), .IN2(n10310), .QN(n10982) );
  INVX0 U11192 ( .INP(g72), .ZN(n10310) );
  NAND4X0 U11193 ( .IN1(n10983), .IN2(n10984), .IN3(n10985), .IN4(n10986), 
        .QN(g33035) );
  OR3X1 U11194 ( .IN1(n8901), .IN2(n5715), .IN3(n8538), .Q(n10986) );
  NAND2X0 U11195 ( .IN1(n8659), .IN2(g4098), .QN(n10985) );
  NAND2X0 U11196 ( .IN1(n8901), .IN2(n5715), .QN(n10983) );
  AND2X1 U11197 ( .IN1(n10987), .IN2(g4098), .Q(n8901) );
  NAND2X0 U11198 ( .IN1(n10988), .IN2(n10989), .QN(g33034) );
  NAND2X0 U11199 ( .IN1(n10990), .IN2(n10991), .QN(n10989) );
  NAND3X0 U11200 ( .IN1(n10992), .IN2(n10993), .IN3(n10994), .QN(n10990) );
  NAND2X0 U11201 ( .IN1(n8512), .IN2(n10995), .QN(n10994) );
  NAND2X0 U11202 ( .IN1(g25676), .IN2(n8209), .QN(n10992) );
  NAND2X0 U11203 ( .IN1(n8659), .IN2(g3873), .QN(n10988) );
  NAND2X0 U11204 ( .IN1(n10996), .IN2(n10997), .QN(g33033) );
  NAND2X0 U11205 ( .IN1(test_so33), .IN2(n10998), .QN(n10997) );
  NAND2X0 U11206 ( .IN1(n10999), .IN2(n8517), .QN(n10998) );
  NAND2X0 U11207 ( .IN1(n5387), .IN2(n10991), .QN(n10999) );
  OR2X1 U11208 ( .IN1(n11000), .IN2(n5387), .Q(n10996) );
  NAND2X0 U11209 ( .IN1(n11001), .IN2(n11002), .QN(g33032) );
  NAND3X0 U11210 ( .IN1(n11003), .IN2(n8209), .IN3(n10991), .QN(n11002) );
  NAND2X0 U11211 ( .IN1(n8659), .IN2(g3863), .QN(n11001) );
  NAND2X0 U11212 ( .IN1(n11004), .IN2(n11005), .QN(g33031) );
  NAND2X0 U11213 ( .IN1(n11006), .IN2(n10991), .QN(n11005) );
  NAND2X0 U11214 ( .IN1(n3482), .IN2(n11007), .QN(n11006) );
  NAND2X0 U11215 ( .IN1(n8511), .IN2(n11008), .QN(n11007) );
  NAND2X0 U11216 ( .IN1(n8658), .IN2(g3857), .QN(n11004) );
  NAND2X0 U11217 ( .IN1(n11009), .IN2(n11010), .QN(g33029) );
  NAND2X0 U11218 ( .IN1(n11011), .IN2(n11012), .QN(n11010) );
  NAND3X0 U11219 ( .IN1(n11013), .IN2(n11014), .IN3(n11015), .QN(n11011) );
  NAND2X0 U11220 ( .IN1(n8512), .IN2(n11016), .QN(n11015) );
  NAND2X0 U11221 ( .IN1(g25662), .IN2(n5645), .QN(n11013) );
  NAND2X0 U11222 ( .IN1(n8658), .IN2(g3522), .QN(n11009) );
  NAND2X0 U11223 ( .IN1(n11017), .IN2(n11018), .QN(g33028) );
  NAND2X0 U11224 ( .IN1(n11019), .IN2(g3518), .QN(n11018) );
  NAND2X0 U11225 ( .IN1(n11020), .IN2(n8517), .QN(n11019) );
  NAND2X0 U11226 ( .IN1(n5383), .IN2(n11012), .QN(n11020) );
  OR2X1 U11227 ( .IN1(n11021), .IN2(n5383), .Q(n11017) );
  NAND2X0 U11228 ( .IN1(n11022), .IN2(n11023), .QN(g33027) );
  NAND3X0 U11229 ( .IN1(n11012), .IN2(n11024), .IN3(n5645), .QN(n11023) );
  NAND2X0 U11230 ( .IN1(n8658), .IN2(g3512), .QN(n11022) );
  NAND2X0 U11231 ( .IN1(n11025), .IN2(n11026), .QN(g33026) );
  NAND2X0 U11232 ( .IN1(n11027), .IN2(n11012), .QN(n11026) );
  NAND2X0 U11233 ( .IN1(n3492), .IN2(n11028), .QN(n11027) );
  NAND2X0 U11234 ( .IN1(n8512), .IN2(n11029), .QN(n11028) );
  NAND2X0 U11235 ( .IN1(n8659), .IN2(g3506), .QN(n11025) );
  NAND3X0 U11236 ( .IN1(n11030), .IN2(n11031), .IN3(n11032), .QN(g33024) );
  NAND2X0 U11237 ( .IN1(g25648), .IN2(n11033), .QN(n11032) );
  NAND2X0 U11238 ( .IN1(n8657), .IN2(g3171), .QN(n11031) );
  NAND3X0 U11239 ( .IN1(n11034), .IN2(n11035), .IN3(n8489), .QN(n11030) );
  NAND2X0 U11240 ( .IN1(n11036), .IN2(n3495), .QN(n11034) );
  NAND2X0 U11241 ( .IN1(n11037), .IN2(n11038), .QN(g33023) );
  NAND3X0 U11242 ( .IN1(n8504), .IN2(g3171), .IN3(n11033), .QN(n11038) );
  NAND2X0 U11243 ( .IN1(n11039), .IN2(g3167), .QN(n11037) );
  NAND2X0 U11244 ( .IN1(n11040), .IN2(n8517), .QN(n11039) );
  NAND2X0 U11245 ( .IN1(n5603), .IN2(n11035), .QN(n11040) );
  NAND2X0 U11246 ( .IN1(n11041), .IN2(n11042), .QN(g33022) );
  NAND2X0 U11247 ( .IN1(n11033), .IN2(n11043), .QN(n11042) );
  NAND2X0 U11248 ( .IN1(n8658), .IN2(g3161), .QN(n11041) );
  NAND2X0 U11249 ( .IN1(n11044), .IN2(n11045), .QN(g33021) );
  NAND2X0 U11250 ( .IN1(n11046), .IN2(n11035), .QN(n11045) );
  NAND2X0 U11251 ( .IN1(n3501), .IN2(n11047), .QN(n11046) );
  NAND2X0 U11252 ( .IN1(n8512), .IN2(n11048), .QN(n11047) );
  NAND2X0 U11253 ( .IN1(n8658), .IN2(g3155), .QN(n11044) );
  NAND3X0 U11254 ( .IN1(n11049), .IN2(n11050), .IN3(n8807), .QN(g33019) );
  NAND2X0 U11255 ( .IN1(n8658), .IN2(g2748), .QN(n11050) );
  NAND2X0 U11256 ( .IN1(n11051), .IN2(n8517), .QN(n11049) );
  XOR2X1 U11257 ( .IN1(test_so30), .IN2(n2790), .Q(n11051) );
  NAND4X0 U11258 ( .IN1(n11052), .IN2(n11053), .IN3(n11054), .IN4(n11055), 
        .QN(g33018) );
  NAND2X0 U11259 ( .IN1(n8657), .IN2(g2610), .QN(n11055) );
  NAND4X0 U11260 ( .IN1(n3511), .IN2(n10495), .IN3(n11056), .IN4(n8130), .QN(
        n11054) );
  NOR2X0 U11261 ( .IN1(n5508), .IN2(n11057), .QN(n11056) );
  NAND3X0 U11262 ( .IN1(n3512), .IN2(n11058), .IN3(n3517), .QN(n11053) );
  INVX0 U11263 ( .INP(n3513), .ZN(n11058) );
  NAND2X0 U11264 ( .IN1(n3524), .IN2(n9776), .QN(n3513) );
  INVX0 U11265 ( .INP(n3006), .ZN(n9776) );
  NAND3X0 U11266 ( .IN1(g2619), .IN2(g110), .IN3(n8130), .QN(n3512) );
  NAND2X0 U11267 ( .IN1(test_so40), .IN2(n11059), .QN(n11052) );
  NAND3X0 U11268 ( .IN1(n11060), .IN2(n10609), .IN3(n11061), .QN(n11059) );
  NAND2X0 U11269 ( .IN1(n3006), .IN2(n8520), .QN(n11061) );
  NAND2X0 U11270 ( .IN1(n3525), .IN2(n3505), .QN(n3006) );
  NAND4X0 U11271 ( .IN1(n11062), .IN2(n11063), .IN3(n11064), .IN4(n11065), 
        .QN(g33017) );
  NAND2X0 U11272 ( .IN1(n11066), .IN2(g2619), .QN(n11064) );
  NAND2X0 U11273 ( .IN1(n3517), .IN2(g2610), .QN(n11063) );
  NAND2X0 U11274 ( .IN1(test_so40), .IN2(n8660), .QN(n11062) );
  NAND3X0 U11275 ( .IN1(n11067), .IN2(n11068), .IN3(n11065), .QN(g33016) );
  NAND2X0 U11276 ( .IN1(n11066), .IN2(g2610), .QN(n11068) );
  NAND2X0 U11277 ( .IN1(n11060), .IN2(g2587), .QN(n11067) );
  NAND4X0 U11278 ( .IN1(n11069), .IN2(n11070), .IN3(n11071), .IN4(n11065), 
        .QN(g33015) );
  INVX0 U11279 ( .INP(n3519), .ZN(n11065) );
  NAND3X0 U11280 ( .IN1(n5508), .IN2(n11072), .IN3(n3517), .QN(n11071) );
  NAND2X0 U11281 ( .IN1(n11066), .IN2(g2587), .QN(n11070) );
  NAND2X0 U11282 ( .IN1(test_so34), .IN2(n8660), .QN(n11069) );
  NAND4X0 U11283 ( .IN1(n11073), .IN2(n11074), .IN3(n11075), .IN4(n11076), 
        .QN(g33014) );
  NAND2X0 U11284 ( .IN1(n8657), .IN2(g2476), .QN(n11076) );
  NAND4X0 U11285 ( .IN1(n3530), .IN2(n10495), .IN3(n11077), .IN4(n8131), .QN(
        n11075) );
  NOR2X0 U11286 ( .IN1(n5509), .IN2(n11078), .QN(n11077) );
  NAND3X0 U11287 ( .IN1(n3531), .IN2(n11079), .IN3(n3536), .QN(n11074) );
  INVX0 U11288 ( .INP(n3532), .ZN(n11079) );
  NAND2X0 U11289 ( .IN1(n3524), .IN2(n9777), .QN(n3532) );
  INVX0 U11290 ( .INP(n3007), .ZN(n9777) );
  NAND3X0 U11291 ( .IN1(g2485), .IN2(g110), .IN3(n8131), .QN(n3531) );
  NAND2X0 U11292 ( .IN1(n11080), .IN2(g2491), .QN(n11073) );
  NAND3X0 U11293 ( .IN1(n11081), .IN2(n10609), .IN3(n11082), .QN(n11080) );
  NAND2X0 U11294 ( .IN1(n3007), .IN2(n8527), .QN(n11082) );
  NAND3X0 U11295 ( .IN1(n5349), .IN2(g2748), .IN3(n3525), .QN(n3007) );
  NAND4X0 U11296 ( .IN1(n11083), .IN2(n11084), .IN3(n11085), .IN4(n11086), 
        .QN(g33013) );
  NAND2X0 U11297 ( .IN1(n11087), .IN2(g2485), .QN(n11085) );
  NAND2X0 U11298 ( .IN1(n3536), .IN2(g2476), .QN(n11084) );
  NAND2X0 U11299 ( .IN1(n8657), .IN2(g2491), .QN(n11083) );
  NAND3X0 U11300 ( .IN1(n11088), .IN2(n11089), .IN3(n11086), .QN(g33012) );
  NAND2X0 U11301 ( .IN1(n11087), .IN2(g2476), .QN(n11089) );
  NAND2X0 U11302 ( .IN1(n11081), .IN2(g2453), .QN(n11088) );
  NAND4X0 U11303 ( .IN1(n11090), .IN2(n11091), .IN3(n11092), .IN4(n11086), 
        .QN(g33011) );
  INVX0 U11304 ( .INP(n3538), .ZN(n11086) );
  NAND3X0 U11305 ( .IN1(n5509), .IN2(n11093), .IN3(n3536), .QN(n11092) );
  NAND2X0 U11306 ( .IN1(n11087), .IN2(g2453), .QN(n11091) );
  NAND2X0 U11307 ( .IN1(n8656), .IN2(g2461), .QN(n11090) );
  NAND4X0 U11308 ( .IN1(n11094), .IN2(n11095), .IN3(n11096), .IN4(n11097), 
        .QN(g33010) );
  NAND2X0 U11309 ( .IN1(test_so21), .IN2(n8661), .QN(n11097) );
  NAND4X0 U11310 ( .IN1(n3548), .IN2(n10495), .IN3(n11098), .IN4(n8213), .QN(
        n11096) );
  NOR2X0 U11311 ( .IN1(n5511), .IN2(n11099), .QN(n11098) );
  NAND3X0 U11312 ( .IN1(n3549), .IN2(n11100), .IN3(n3555), .QN(n11095) );
  INVX0 U11313 ( .INP(n3551), .ZN(n11100) );
  NAND2X0 U11314 ( .IN1(n3524), .IN2(n9778), .QN(n3551) );
  INVX0 U11315 ( .INP(n3550), .ZN(n9778) );
  NAND3X0 U11316 ( .IN1(g110), .IN2(n8213), .IN3(g2351), .QN(n3549) );
  NAND2X0 U11317 ( .IN1(n11101), .IN2(g2357), .QN(n11094) );
  NAND3X0 U11318 ( .IN1(n11102), .IN2(n10609), .IN3(n11103), .QN(n11101) );
  NAND2X0 U11319 ( .IN1(n3550), .IN2(n8528), .QN(n11103) );
  NAND3X0 U11320 ( .IN1(n5516), .IN2(g2741), .IN3(n3525), .QN(n3550) );
  NAND4X0 U11321 ( .IN1(n11104), .IN2(n11105), .IN3(n11106), .IN4(n11107), 
        .QN(g33009) );
  NAND2X0 U11322 ( .IN1(n11108), .IN2(g2351), .QN(n11106) );
  NAND2X0 U11323 ( .IN1(n3555), .IN2(test_so21), .QN(n11105) );
  NAND2X0 U11324 ( .IN1(n8656), .IN2(g2357), .QN(n11104) );
  NAND3X0 U11325 ( .IN1(n11109), .IN2(n11110), .IN3(n11107), .QN(g33008) );
  NAND2X0 U11326 ( .IN1(n11108), .IN2(test_so21), .QN(n11110) );
  NAND2X0 U11327 ( .IN1(n11102), .IN2(g2319), .QN(n11109) );
  NAND4X0 U11328 ( .IN1(n11111), .IN2(n11112), .IN3(n11113), .IN4(n11107), 
        .QN(g33007) );
  INVX0 U11329 ( .INP(n3557), .ZN(n11107) );
  NAND3X0 U11330 ( .IN1(n5511), .IN2(n11114), .IN3(n3555), .QN(n11113) );
  NAND2X0 U11331 ( .IN1(n11108), .IN2(g2319), .QN(n11112) );
  NAND2X0 U11332 ( .IN1(n8655), .IN2(g2327), .QN(n11111) );
  NAND4X0 U11333 ( .IN1(n11115), .IN2(n11116), .IN3(n11117), .IN4(n11118), 
        .QN(g33006) );
  NAND2X0 U11334 ( .IN1(n8656), .IN2(g2208), .QN(n11118) );
  NAND4X0 U11335 ( .IN1(n3567), .IN2(n10495), .IN3(n11119), .IN4(n8133), .QN(
        n11117) );
  NOR2X0 U11336 ( .IN1(n5512), .IN2(n11120), .QN(n11119) );
  NAND3X0 U11337 ( .IN1(n3568), .IN2(n11121), .IN3(n3574), .QN(n11116) );
  INVX0 U11338 ( .INP(n3570), .ZN(n11121) );
  NAND2X0 U11339 ( .IN1(n3524), .IN2(n9779), .QN(n3570) );
  INVX0 U11340 ( .INP(n3569), .ZN(n9779) );
  NAND3X0 U11341 ( .IN1(g2217), .IN2(g110), .IN3(n8133), .QN(n3568) );
  NAND2X0 U11342 ( .IN1(n11122), .IN2(g2223), .QN(n11115) );
  NAND3X0 U11343 ( .IN1(n11123), .IN2(n10609), .IN3(n11124), .QN(n11122) );
  NAND2X0 U11344 ( .IN1(n3569), .IN2(n8528), .QN(n11124) );
  NAND3X0 U11345 ( .IN1(n5349), .IN2(n5516), .IN3(n3525), .QN(n3569) );
  NAND4X0 U11346 ( .IN1(n11125), .IN2(n11126), .IN3(n11127), .IN4(n11128), 
        .QN(g33005) );
  NAND2X0 U11347 ( .IN1(n11129), .IN2(g2217), .QN(n11127) );
  NAND2X0 U11348 ( .IN1(n3574), .IN2(g2208), .QN(n11126) );
  NAND2X0 U11349 ( .IN1(n8655), .IN2(g2223), .QN(n11125) );
  NAND3X0 U11350 ( .IN1(n11130), .IN2(n11131), .IN3(n11128), .QN(g33004) );
  NAND2X0 U11351 ( .IN1(n11129), .IN2(g2208), .QN(n11131) );
  NAND2X0 U11352 ( .IN1(n11123), .IN2(g2185), .QN(n11130) );
  NAND4X0 U11353 ( .IN1(n11132), .IN2(n11133), .IN3(n11134), .IN4(n11128), 
        .QN(g33003) );
  INVX0 U11354 ( .INP(n3576), .ZN(n11128) );
  NAND3X0 U11355 ( .IN1(n5512), .IN2(n11135), .IN3(n3574), .QN(n11134) );
  NAND2X0 U11356 ( .IN1(n11129), .IN2(g2185), .QN(n11133) );
  NAND2X0 U11357 ( .IN1(n8655), .IN2(g2193), .QN(n11132) );
  NAND4X0 U11358 ( .IN1(n11136), .IN2(n11137), .IN3(n11138), .IN4(n11139), 
        .QN(g33002) );
  NAND2X0 U11359 ( .IN1(n8655), .IN2(g2051), .QN(n11139) );
  NAND4X0 U11360 ( .IN1(n3586), .IN2(n10495), .IN3(n11140), .IN4(n8129), .QN(
        n11138) );
  NOR2X0 U11361 ( .IN1(n5507), .IN2(n11141), .QN(n11140) );
  NAND3X0 U11362 ( .IN1(n3587), .IN2(n11142), .IN3(n3593), .QN(n11137) );
  INVX0 U11363 ( .INP(n3589), .ZN(n11142) );
  NAND2X0 U11364 ( .IN1(n3524), .IN2(n9769), .QN(n3589) );
  INVX0 U11365 ( .INP(n3588), .ZN(n9769) );
  NAND3X0 U11366 ( .IN1(g2060), .IN2(g110), .IN3(n8129), .QN(n3587) );
  NAND2X0 U11367 ( .IN1(n11143), .IN2(g2066), .QN(n11136) );
  NAND3X0 U11368 ( .IN1(n11144), .IN2(n10609), .IN3(n11145), .QN(n11143) );
  NAND2X0 U11369 ( .IN1(n3588), .IN2(n8528), .QN(n11145) );
  NAND3X0 U11370 ( .IN1(n3581), .IN2(n5300), .IN3(n3505), .QN(n3588) );
  NAND4X0 U11371 ( .IN1(n11146), .IN2(n11147), .IN3(n11148), .IN4(n11149), 
        .QN(g33001) );
  NAND2X0 U11372 ( .IN1(n11150), .IN2(g2060), .QN(n11148) );
  NAND2X0 U11373 ( .IN1(n3593), .IN2(g2051), .QN(n11147) );
  NAND2X0 U11374 ( .IN1(n8655), .IN2(g2066), .QN(n11146) );
  NAND3X0 U11375 ( .IN1(n11151), .IN2(n11152), .IN3(n11149), .QN(g33000) );
  NAND2X0 U11376 ( .IN1(n11150), .IN2(g2051), .QN(n11152) );
  NAND2X0 U11377 ( .IN1(n11144), .IN2(g2028), .QN(n11151) );
  NAND4X0 U11378 ( .IN1(n11153), .IN2(n11154), .IN3(n11155), .IN4(n11149), 
        .QN(g32999) );
  INVX0 U11379 ( .INP(n3595), .ZN(n11149) );
  NAND3X0 U11380 ( .IN1(n5507), .IN2(n11156), .IN3(n3593), .QN(n11155) );
  NAND2X0 U11381 ( .IN1(n11150), .IN2(g2028), .QN(n11154) );
  NAND2X0 U11382 ( .IN1(test_so59), .IN2(n8661), .QN(n11153) );
  NAND4X0 U11383 ( .IN1(n11157), .IN2(n11158), .IN3(n11159), .IN4(n11160), 
        .QN(g32998) );
  NAND2X0 U11384 ( .IN1(n8654), .IN2(g1917), .QN(n11160) );
  NAND4X0 U11385 ( .IN1(n3604), .IN2(n10495), .IN3(n11161), .IN4(n8132), .QN(
        n11159) );
  NOR2X0 U11386 ( .IN1(n5510), .IN2(n11162), .QN(n11161) );
  NAND3X0 U11387 ( .IN1(n3605), .IN2(n11163), .IN3(n3611), .QN(n11158) );
  INVX0 U11388 ( .INP(n3607), .ZN(n11163) );
  NAND2X0 U11389 ( .IN1(n3524), .IN2(n9770), .QN(n3607) );
  INVX0 U11390 ( .INP(n3606), .ZN(n9770) );
  NAND3X0 U11391 ( .IN1(g1926), .IN2(g110), .IN3(n8132), .QN(n3605) );
  NAND2X0 U11392 ( .IN1(n11164), .IN2(g1932), .QN(n11157) );
  NAND3X0 U11393 ( .IN1(n11165), .IN2(n10609), .IN3(n11166), .QN(n11164) );
  NAND2X0 U11394 ( .IN1(n3606), .IN2(n8528), .QN(n11166) );
  NAND4X0 U11395 ( .IN1(n3581), .IN2(n5349), .IN3(g2748), .IN4(n5300), .QN(
        n3606) );
  NAND4X0 U11396 ( .IN1(n11167), .IN2(n11168), .IN3(n11169), .IN4(n11170), 
        .QN(g32997) );
  NAND2X0 U11397 ( .IN1(n11171), .IN2(g1926), .QN(n11169) );
  NAND2X0 U11398 ( .IN1(n3611), .IN2(g1917), .QN(n11168) );
  NAND2X0 U11399 ( .IN1(n8654), .IN2(g1932), .QN(n11167) );
  NAND3X0 U11400 ( .IN1(n11172), .IN2(n11173), .IN3(n11170), .QN(g32996) );
  NAND2X0 U11401 ( .IN1(n11171), .IN2(g1917), .QN(n11173) );
  NAND2X0 U11402 ( .IN1(n11165), .IN2(g1894), .QN(n11172) );
  NAND4X0 U11403 ( .IN1(n11174), .IN2(n11175), .IN3(n11176), .IN4(n11170), 
        .QN(g32995) );
  INVX0 U11404 ( .INP(n3613), .ZN(n11170) );
  NAND3X0 U11405 ( .IN1(n5510), .IN2(n11177), .IN3(n3611), .QN(n11176) );
  NAND2X0 U11406 ( .IN1(n11171), .IN2(g1894), .QN(n11175) );
  NAND2X0 U11407 ( .IN1(n8654), .IN2(g1902), .QN(n11174) );
  NAND4X0 U11408 ( .IN1(n11178), .IN2(n11179), .IN3(n11180), .IN4(n11181), 
        .QN(g32994) );
  NAND2X0 U11409 ( .IN1(n8654), .IN2(g1783), .QN(n11181) );
  NAND4X0 U11410 ( .IN1(n3622), .IN2(n10495), .IN3(n11182), .IN4(n5596), .QN(
        n11180) );
  NOR2X0 U11411 ( .IN1(n5359), .IN2(n11183), .QN(n11182) );
  NAND3X0 U11412 ( .IN1(n3623), .IN2(n11184), .IN3(n3628), .QN(n11179) );
  INVX0 U11413 ( .INP(n3624), .ZN(n11184) );
  NAND2X0 U11414 ( .IN1(n3524), .IN2(n3005), .QN(n3624) );
  NAND3X0 U11415 ( .IN1(g1792), .IN2(g110), .IN3(n5596), .QN(n3623) );
  NAND2X0 U11416 ( .IN1(n11185), .IN2(g1798), .QN(n11178) );
  NAND3X0 U11417 ( .IN1(n11186), .IN2(n10609), .IN3(n11187), .QN(n11185) );
  NAND2X0 U11418 ( .IN1(n8511), .IN2(n1413), .QN(n11187) );
  INVX0 U11419 ( .INP(n3005), .ZN(n1413) );
  NAND4X0 U11420 ( .IN1(n11188), .IN2(n11189), .IN3(n11190), .IN4(n11191), 
        .QN(g32993) );
  NAND2X0 U11421 ( .IN1(n11192), .IN2(g1792), .QN(n11190) );
  NAND2X0 U11422 ( .IN1(n3628), .IN2(g1783), .QN(n11189) );
  NAND2X0 U11423 ( .IN1(n8654), .IN2(g1798), .QN(n11188) );
  NAND3X0 U11424 ( .IN1(n11193), .IN2(n11194), .IN3(n11191), .QN(g32992) );
  NAND2X0 U11425 ( .IN1(n11192), .IN2(g1783), .QN(n11194) );
  NAND2X0 U11426 ( .IN1(n11186), .IN2(g1760), .QN(n11193) );
  NAND4X0 U11427 ( .IN1(n11195), .IN2(n11196), .IN3(n11197), .IN4(n11191), 
        .QN(g32991) );
  INVX0 U11428 ( .INP(n3630), .ZN(n11191) );
  NAND3X0 U11429 ( .IN1(n5359), .IN2(n11198), .IN3(n3628), .QN(n11197) );
  NAND2X0 U11430 ( .IN1(n11192), .IN2(g1760), .QN(n11196) );
  NAND2X0 U11431 ( .IN1(n8653), .IN2(g1768), .QN(n11195) );
  NAND4X0 U11432 ( .IN1(n11199), .IN2(n11200), .IN3(n11201), .IN4(n11202), 
        .QN(g32990) );
  NAND2X0 U11433 ( .IN1(test_so94), .IN2(n8661), .QN(n11202) );
  NAND4X0 U11434 ( .IN1(n3640), .IN2(n10495), .IN3(n11203), .IN4(n8210), .QN(
        n11201) );
  NOR2X0 U11435 ( .IN1(n5525), .IN2(n11204), .QN(n11203) );
  INVX0 U11436 ( .INP(n9539), .ZN(n10495) );
  NAND3X0 U11437 ( .IN1(n3641), .IN2(n11205), .IN3(n3646), .QN(n11200) );
  INVX0 U11438 ( .INP(n3642), .ZN(n11205) );
  NAND2X0 U11439 ( .IN1(n3524), .IN2(n9771), .QN(n3642) );
  INVX0 U11440 ( .INP(n3003), .ZN(n9771) );
  NAND3X0 U11441 ( .IN1(g110), .IN2(n8210), .IN3(g1657), .QN(n3641) );
  NAND2X0 U11442 ( .IN1(n11206), .IN2(g1664), .QN(n11199) );
  NAND3X0 U11443 ( .IN1(n11207), .IN2(n10609), .IN3(n11208), .QN(n11206) );
  NAND2X0 U11444 ( .IN1(n3003), .IN2(n8528), .QN(n11208) );
  NAND2X0 U11445 ( .IN1(n3653), .IN2(n3581), .QN(n3003) );
  AND2X1 U11446 ( .IN1(n11209), .IN2(n11210), .Q(n3581) );
  XOR2X1 U11447 ( .IN1(n7684), .IN2(g72), .Q(n11210) );
  XOR2X1 U11448 ( .IN1(n7689), .IN2(g73), .Q(n11209) );
  NAND2X0 U11449 ( .IN1(n8511), .IN2(n1430), .QN(n10609) );
  INVX0 U11450 ( .INP(n2760), .ZN(n1430) );
  NAND4X0 U11451 ( .IN1(n11211), .IN2(n11212), .IN3(n11213), .IN4(n11214), 
        .QN(g32989) );
  NAND2X0 U11452 ( .IN1(n11215), .IN2(g1657), .QN(n11213) );
  NAND2X0 U11453 ( .IN1(n3646), .IN2(test_so94), .QN(n11212) );
  NAND2X0 U11454 ( .IN1(n8653), .IN2(g1664), .QN(n11211) );
  NAND3X0 U11455 ( .IN1(n11216), .IN2(n11217), .IN3(n11214), .QN(g32988) );
  NAND2X0 U11456 ( .IN1(n11215), .IN2(test_so94), .QN(n11217) );
  NAND2X0 U11457 ( .IN1(n11207), .IN2(g1624), .QN(n11216) );
  NAND4X0 U11458 ( .IN1(n11218), .IN2(n11219), .IN3(n11220), .IN4(n11214), 
        .QN(g32987) );
  INVX0 U11459 ( .INP(n3648), .ZN(n11214) );
  NAND3X0 U11460 ( .IN1(n5525), .IN2(n11221), .IN3(n3646), .QN(n11220) );
  NAND2X0 U11461 ( .IN1(n11215), .IN2(g1624), .QN(n11219) );
  NAND2X0 U11462 ( .IN1(n8653), .IN2(g1632), .QN(n11218) );
  NAND3X0 U11463 ( .IN1(n11222), .IN2(n11223), .IN3(n11224), .QN(g32986) );
  NAND3X0 U11464 ( .IN1(n10799), .IN2(n7849), .IN3(n11225), .QN(n11224) );
  INVX0 U11465 ( .INP(n11226), .ZN(n10799) );
  NAND3X0 U11466 ( .IN1(n11226), .IN2(g1373), .IN3(n8490), .QN(n11223) );
  NAND2X0 U11467 ( .IN1(n155), .IN2(n11227), .QN(n11226) );
  NAND2X0 U11468 ( .IN1(n7814), .IN2(n10801), .QN(n11227) );
  INVX0 U11469 ( .INP(n11228), .ZN(n155) );
  NAND2X0 U11470 ( .IN1(n8653), .IN2(g1367), .QN(n11222) );
  NOR2X0 U11471 ( .IN1(n5730), .IN2(n11229), .QN(g32985) );
  NOR2X0 U11472 ( .IN1(n8568), .IN2(n11230), .QN(n11229) );
  AND2X1 U11473 ( .IN1(n9311), .IN2(n10808), .Q(n11230) );
  NOR2X0 U11474 ( .IN1(n11231), .IN2(n5716), .QN(n10808) );
  NAND3X0 U11475 ( .IN1(n11232), .IN2(n11233), .IN3(n11234), .QN(g32984) );
  OR2X1 U11476 ( .IN1(n8478), .IN2(n5674), .Q(n11234) );
  NAND3X0 U11477 ( .IN1(n11235), .IN2(n11231), .IN3(g1270), .QN(n11233) );
  INVX0 U11478 ( .INP(n3662), .ZN(n11231) );
  NAND2X0 U11479 ( .IN1(n5716), .IN2(n3662), .QN(n11232) );
  NAND3X0 U11480 ( .IN1(n11236), .IN2(n11237), .IN3(n11238), .QN(g32983) );
  NAND3X0 U11481 ( .IN1(n10812), .IN2(n7851), .IN3(n11239), .QN(n11238) );
  INVX0 U11482 ( .INP(n11240), .ZN(n10812) );
  NAND3X0 U11483 ( .IN1(n11240), .IN2(g1030), .IN3(n8490), .QN(n11237) );
  NAND2X0 U11484 ( .IN1(n435), .IN2(n11241), .QN(n11240) );
  NAND2X0 U11485 ( .IN1(n7815), .IN2(n10814), .QN(n11241) );
  INVX0 U11486 ( .INP(n11242), .ZN(n435) );
  NAND2X0 U11487 ( .IN1(n8653), .IN2(g1024), .QN(n11236) );
  NOR2X0 U11488 ( .IN1(n5731), .IN2(n11243), .QN(g32982) );
  NOR2X0 U11489 ( .IN1(n8569), .IN2(n11244), .QN(n11243) );
  AND2X1 U11490 ( .IN1(n11245), .IN2(n10821), .Q(n11244) );
  NOR2X0 U11491 ( .IN1(n11246), .IN2(n5725), .QN(n10821) );
  NAND3X0 U11492 ( .IN1(n11247), .IN2(n11248), .IN3(n11249), .QN(g32981) );
  OR2X1 U11493 ( .IN1(n8478), .IN2(n5673), .Q(n11249) );
  NAND3X0 U11494 ( .IN1(n11250), .IN2(n11246), .IN3(g925), .QN(n11248) );
  INVX0 U11495 ( .INP(n3671), .ZN(n11246) );
  NAND2X0 U11496 ( .IN1(n5725), .IN2(n3671), .QN(n11247) );
  AND3X1 U11497 ( .IN1(n11251), .IN2(n11252), .IN3(n8452), .Q(g32980) );
  NAND2X0 U11498 ( .IN1(n5754), .IN2(n9591), .QN(n11252) );
  NAND2X0 U11499 ( .IN1(n2644), .IN2(n11253), .QN(n11251) );
  INVX0 U11500 ( .INP(n9591), .ZN(n11253) );
  NAND4X0 U11501 ( .IN1(n5632), .IN2(g376), .IN3(g8719), .IN4(g370), .QN(n9591) );
  NAND3X0 U11502 ( .IN1(n11254), .IN2(n11255), .IN3(n11256), .QN(g32979) );
  NAND2X0 U11503 ( .IN1(test_so2), .IN2(n8534), .QN(n11256) );
  NAND3X0 U11504 ( .IN1(n2404), .IN2(n11257), .IN3(g758), .QN(n11255) );
  INVX0 U11505 ( .INP(n3272), .ZN(n11257) );
  NAND2X0 U11506 ( .IN1(n3272), .IN2(n5331), .QN(n11254) );
  NAND3X0 U11507 ( .IN1(n11258), .IN2(n11259), .IN3(n11260), .QN(g32978) );
  NAND2X0 U11508 ( .IN1(n8652), .IN2(g582), .QN(n11260) );
  NAND3X0 U11509 ( .IN1(n2421), .IN2(n11261), .IN3(g590), .QN(n11259) );
  INVX0 U11510 ( .INP(n3274), .ZN(n11261) );
  NAND2X0 U11511 ( .IN1(n3274), .IN2(n5472), .QN(n11258) );
  NAND3X0 U11512 ( .IN1(n11262), .IN2(n11263), .IN3(n11264), .QN(g32977) );
  NAND2X0 U11513 ( .IN1(test_so51), .IN2(n8533), .QN(n11264) );
  NAND3X0 U11514 ( .IN1(n8194), .IN2(n11265), .IN3(g291), .QN(n11263) );
  NAND2X0 U11515 ( .IN1(n42), .IN2(n5679), .QN(n11262) );
  INVX0 U11516 ( .INP(n11265), .ZN(n42) );
  NAND3X0 U11517 ( .IN1(test_so51), .IN2(n11266), .IN3(test_so55), .QN(n11265)
         );
  NAND3X0 U11518 ( .IN1(n11267), .IN2(n11268), .IN3(n11269), .QN(g32976) );
  NAND2X0 U11519 ( .IN1(n8652), .IN2(g164), .QN(n11269) );
  OR3X1 U11520 ( .IN1(n9761), .IN2(n3281), .IN3(n5676), .Q(n11268) );
  NAND2X0 U11521 ( .IN1(n3281), .IN2(n5676), .QN(n11267) );
  NOR4X0 U11522 ( .IN1(n11270), .IN2(n11271), .IN3(n11272), .IN4(n11273), .QN(
        g32185) );
  NOR2X0 U11523 ( .IN1(n8172), .IN2(n8171), .QN(n11273) );
  AND2X1 U11524 ( .IN1(g2902), .IN2(test_so1), .Q(n11272) );
  NOR2X0 U11525 ( .IN1(n7819), .IN2(n8235), .QN(n11271) );
  NAND4X0 U11526 ( .IN1(n11274), .IN2(n11275), .IN3(n11276), .IN4(n11277), 
        .QN(n11270) );
  OR2X1 U11527 ( .IN1(n5750), .IN2(n8167), .Q(n11277) );
  NAND2X0 U11528 ( .IN1(g2955), .IN2(g2950), .QN(n11276) );
  NAND2X0 U11529 ( .IN1(g2927), .IN2(g2922), .QN(n11275) );
  NAND2X0 U11530 ( .IN1(g2917), .IN2(g2912), .QN(n11274) );
  NAND4X0 U11531 ( .IN1(n11278), .IN2(n11279), .IN3(n11280), .IN4(n11281), 
        .QN(g31904) );
  NAND4X0 U11532 ( .IN1(n11282), .IN2(n11283), .IN3(n10964), .IN4(g5033), .QN(
        n11281) );
  OR2X1 U11533 ( .IN1(g5033), .IN2(n11282), .Q(n11280) );
  NAND2X0 U11534 ( .IN1(n8652), .IN2(g5029), .QN(n11279) );
  NAND2X0 U11535 ( .IN1(n11284), .IN2(n8528), .QN(n11278) );
  NAND4X0 U11536 ( .IN1(n11285), .IN2(n10962), .IN3(n11286), .IN4(n11287), 
        .QN(g31903) );
  OR4X1 U11537 ( .IN1(n10965), .IN2(n11288), .IN3(n11289), .IN4(n5607), .Q(
        n11287) );
  NAND2X0 U11538 ( .IN1(n5607), .IN2(n10965), .QN(n11286) );
  NOR2X0 U11539 ( .IN1(n11290), .IN2(n5578), .QN(n10965) );
  NAND3X0 U11540 ( .IN1(n11288), .IN2(n8481), .IN3(n5607), .QN(n10962) );
  NAND2X0 U11541 ( .IN1(n8652), .IN2(g5046), .QN(n11285) );
  NAND3X0 U11542 ( .IN1(n11291), .IN2(n11292), .IN3(n11293), .QN(g31902) );
  OR2X1 U11543 ( .IN1(n11283), .IN2(n8545), .Q(n11293) );
  NAND4X0 U11544 ( .IN1(n10964), .IN2(g5029), .IN3(n11294), .IN4(n11295), .QN(
        n11292) );
  NAND2X0 U11545 ( .IN1(n5369), .IN2(g5022), .QN(n11295) );
  NAND2X0 U11546 ( .IN1(g5016), .IN2(g5062), .QN(n11294) );
  NAND2X0 U11547 ( .IN1(n11296), .IN2(g5016), .QN(n11291) );
  NAND2X0 U11548 ( .IN1(n11297), .IN2(n8528), .QN(n11296) );
  NAND2X0 U11549 ( .IN1(n5601), .IN2(g5062), .QN(n11297) );
  NAND4X0 U11550 ( .IN1(n11298), .IN2(n11299), .IN3(n11300), .IN4(n11301), 
        .QN(g31901) );
  NAND4X0 U11551 ( .IN1(n11302), .IN2(n11290), .IN3(n10964), .IN4(g5046), .QN(
        n11301) );
  OR2X1 U11552 ( .IN1(n11290), .IN2(g5046), .Q(n11300) );
  NAND3X0 U11553 ( .IN1(g5041), .IN2(g5037), .IN3(n11303), .QN(n11290) );
  NAND2X0 U11554 ( .IN1(n8651), .IN2(g5041), .QN(n11299) );
  NAND2X0 U11555 ( .IN1(n11288), .IN2(n8528), .QN(n11298) );
  NOR2X0 U11556 ( .IN1(n11302), .IN2(g5046), .QN(n11288) );
  NAND3X0 U11557 ( .IN1(n5605), .IN2(n11284), .IN3(n5611), .QN(n11302) );
  NAND3X0 U11558 ( .IN1(n11304), .IN2(n11305), .IN3(n11306), .QN(g31900) );
  OR2X1 U11559 ( .IN1(n11307), .IN2(g5041), .Q(n11306) );
  NAND4X0 U11560 ( .IN1(n11308), .IN2(g5041), .IN3(n10964), .IN4(n5611), .QN(
        n11305) );
  NAND2X0 U11561 ( .IN1(n11309), .IN2(g5037), .QN(n11304) );
  NAND3X0 U11562 ( .IN1(n11310), .IN2(n11311), .IN3(n8490), .QN(n11309) );
  NAND3X0 U11563 ( .IN1(n11312), .IN2(n11313), .IN3(g5041), .QN(n11311) );
  NAND2X0 U11564 ( .IN1(n5605), .IN2(n11303), .QN(n11310) );
  NAND4X0 U11565 ( .IN1(n11314), .IN2(n11307), .IN3(n11315), .IN4(n11316), 
        .QN(g31899) );
  NAND4X0 U11566 ( .IN1(n11308), .IN2(n11313), .IN3(n10964), .IN4(g5037), .QN(
        n11316) );
  INVX0 U11567 ( .INP(n11289), .ZN(n10964) );
  INVX0 U11568 ( .INP(n11303), .ZN(n11313) );
  INVX0 U11569 ( .INP(n11284), .ZN(n11308) );
  NAND2X0 U11570 ( .IN1(n5611), .IN2(n11303), .QN(n11315) );
  NOR2X0 U11571 ( .IN1(n11282), .IN2(n7838), .QN(n11303) );
  NAND3X0 U11572 ( .IN1(g5029), .IN2(g5062), .IN3(g5016), .QN(n11282) );
  NAND3X0 U11573 ( .IN1(n11284), .IN2(n8481), .IN3(n5611), .QN(n11307) );
  NOR2X0 U11574 ( .IN1(g5033), .IN2(n11283), .QN(n11284) );
  NAND3X0 U11575 ( .IN1(n5369), .IN2(g5022), .IN3(n5601), .QN(n11283) );
  NAND2X0 U11576 ( .IN1(n8651), .IN2(g5033), .QN(n11314) );
  NAND3X0 U11577 ( .IN1(n11317), .IN2(n11318), .IN3(n11319), .QN(g31898) );
  OR3X1 U11578 ( .IN1(n11289), .IN2(n11320), .IN3(g5016), .Q(n11319) );
  NAND2X0 U11579 ( .IN1(n11312), .IN2(n8527), .QN(n11289) );
  AND2X1 U11580 ( .IN1(n11321), .IN2(n11322), .Q(n11312) );
  NAND3X0 U11581 ( .IN1(n11320), .IN2(g5016), .IN3(n8490), .QN(n11318) );
  NOR2X0 U11582 ( .IN1(g5022), .IN2(g5062), .QN(n11320) );
  NAND2X0 U11583 ( .IN1(n8651), .IN2(g5022), .QN(n11317) );
  NAND3X0 U11584 ( .IN1(n11323), .IN2(n10431), .IN3(n11324), .QN(g31897) );
  NAND2X0 U11585 ( .IN1(n10973), .IN2(g4575), .QN(n10431) );
  NAND2X0 U11586 ( .IN1(n8651), .IN2(g4423), .QN(n11323) );
  NAND3X0 U11587 ( .IN1(n11325), .IN2(n10436), .IN3(n11324), .QN(g31896) );
  AND2X1 U11588 ( .IN1(n11326), .IN2(n11327), .Q(n11324) );
  NAND2X0 U11589 ( .IN1(n10973), .IN2(n11328), .QN(n11327) );
  NAND2X0 U11590 ( .IN1(g72), .IN2(g73), .QN(n11328) );
  NAND2X0 U11591 ( .IN1(n10437), .IN2(g4372), .QN(n11326) );
  INVX0 U11592 ( .INP(n11329), .ZN(n10437) );
  NAND2X0 U11593 ( .IN1(test_so100), .IN2(n10973), .QN(n10436) );
  NOR2X0 U11594 ( .IN1(n8575), .IN2(n5670), .QN(n10973) );
  OR2X1 U11595 ( .IN1(n8479), .IN2(n5849), .Q(n11325) );
  NAND2X0 U11596 ( .IN1(n9539), .IN2(n11330), .QN(g31895) );
  OR2X1 U11597 ( .IN1(n8479), .IN2(n5714), .Q(n11330) );
  NAND2X0 U11598 ( .IN1(n2760), .IN2(n8528), .QN(n9539) );
  NAND3X0 U11599 ( .IN1(n11331), .IN2(n11332), .IN3(n10984), .QN(g31894) );
  NAND2X0 U11600 ( .IN1(n8650), .IN2(g4093), .QN(n11332) );
  NAND2X0 U11601 ( .IN1(n11333), .IN2(n8527), .QN(n11331) );
  XOR2X1 U11602 ( .IN1(n10987), .IN2(g4098), .Q(n11333) );
  NOR2X0 U11603 ( .IN1(n3729), .IN2(n5340), .QN(n10987) );
  NAND2X0 U11604 ( .IN1(n11334), .IN2(g4087), .QN(n3729) );
  NAND2X0 U11605 ( .IN1(n11335), .IN2(n11336), .QN(g31872) );
  NAND2X0 U11606 ( .IN1(n11337), .IN2(n3730), .QN(n11336) );
  XOR2X1 U11607 ( .IN1(n11338), .IN2(n5516), .Q(n11337) );
  NAND2X0 U11608 ( .IN1(n8897), .IN2(g2741), .QN(n11338) );
  NAND2X0 U11609 ( .IN1(n8650), .IN2(g2741), .QN(n11335) );
  NAND3X0 U11610 ( .IN1(n11339), .IN2(n11340), .IN3(n11341), .QN(g31871) );
  NAND2X0 U11611 ( .IN1(n3733), .IN2(n11225), .QN(n11341) );
  NAND2X0 U11612 ( .IN1(n8650), .IN2(g1361), .QN(n11340) );
  NAND3X0 U11613 ( .IN1(n11228), .IN2(g1367), .IN3(n8490), .QN(n11339) );
  NAND2X0 U11614 ( .IN1(n156), .IN2(n11342), .QN(n11228) );
  NAND2X0 U11615 ( .IN1(n7848), .IN2(n10801), .QN(n11342) );
  INVX0 U11616 ( .INP(n11343), .ZN(n156) );
  NAND3X0 U11617 ( .IN1(n11344), .IN2(n11345), .IN3(n11346), .QN(g31870) );
  OR2X1 U11618 ( .IN1(n8479), .IN2(n5553), .Q(n11346) );
  OR3X1 U11619 ( .IN1(n10807), .IN2(n3664), .IN3(n5674), .Q(n11345) );
  NAND2X0 U11620 ( .IN1(n3664), .IN2(n5674), .QN(n11344) );
  NAND3X0 U11621 ( .IN1(n11347), .IN2(n11348), .IN3(n11349), .QN(g31869) );
  NAND2X0 U11622 ( .IN1(n3738), .IN2(n11239), .QN(n11349) );
  NAND2X0 U11623 ( .IN1(n8650), .IN2(g1018), .QN(n11348) );
  NAND3X0 U11624 ( .IN1(n11242), .IN2(g1024), .IN3(n8490), .QN(n11347) );
  NAND2X0 U11625 ( .IN1(n436), .IN2(n11350), .QN(n11242) );
  NAND2X0 U11626 ( .IN1(n7850), .IN2(n10814), .QN(n11350) );
  INVX0 U11627 ( .INP(n11351), .ZN(n436) );
  NAND3X0 U11628 ( .IN1(n11352), .IN2(n11353), .IN3(n11354), .QN(g31868) );
  OR2X1 U11629 ( .IN1(n8479), .IN2(n5560), .Q(n11354) );
  OR3X1 U11630 ( .IN1(n10820), .IN2(n3673), .IN3(n5673), .Q(n11353) );
  NAND2X0 U11631 ( .IN1(n3673), .IN2(n5673), .QN(n11352) );
  NAND3X0 U11632 ( .IN1(n11355), .IN2(n11356), .IN3(n11357), .QN(g31867) );
  NAND2X0 U11633 ( .IN1(n8650), .IN2(g744), .QN(n11357) );
  NAND3X0 U11634 ( .IN1(n2404), .IN2(test_so2), .IN3(n11358), .QN(n11356) );
  INVX0 U11635 ( .INP(n3682), .ZN(n11358) );
  NAND2X0 U11636 ( .IN1(n3682), .IN2(n5471), .QN(n11355) );
  NAND3X0 U11637 ( .IN1(n11359), .IN2(n11360), .IN3(n11361), .QN(g31866) );
  NAND2X0 U11638 ( .IN1(n8650), .IN2(g577), .QN(n11361) );
  NAND3X0 U11639 ( .IN1(n2421), .IN2(n11362), .IN3(g582), .QN(n11360) );
  INVX0 U11640 ( .INP(n3684), .ZN(n11362) );
  NAND2X0 U11641 ( .IN1(n3684), .IN2(n5552), .QN(n11359) );
  NAND2X0 U11642 ( .IN1(n11363), .IN2(n11364), .QN(g31865) );
  NAND2X0 U11643 ( .IN1(test_so55), .IN2(n11365), .QN(n11364) );
  NAND2X0 U11644 ( .IN1(n11366), .IN2(n8528), .QN(n11365) );
  NAND2X0 U11645 ( .IN1(n11266), .IN2(n8241), .QN(n11366) );
  NAND3X0 U11646 ( .IN1(n8194), .IN2(test_so51), .IN3(n8228), .QN(n11363) );
  NAND3X0 U11647 ( .IN1(n11367), .IN2(n11368), .IN3(n11369), .QN(g31864) );
  NAND2X0 U11648 ( .IN1(test_so73), .IN2(n8548), .QN(n11369) );
  NAND3X0 U11649 ( .IN1(n11370), .IN2(n11371), .IN3(g164), .QN(n11368) );
  NAND2X0 U11650 ( .IN1(n45), .IN2(n5561), .QN(n11367) );
  INVX0 U11651 ( .INP(n11371), .ZN(n45) );
  NAND3X0 U11652 ( .IN1(n11372), .IN2(n11373), .IN3(test_so73), .QN(n11371) );
  NOR2X0 U11653 ( .IN1(g1636), .IN2(n5598), .QN(g31862) );
  NAND2X0 U11654 ( .IN1(n11374), .IN2(n11375), .QN(g31793) );
  NAND3X0 U11655 ( .IN1(n11376), .IN2(n11377), .IN3(n9260), .QN(n11375) );
  NOR2X0 U11656 ( .IN1(n11378), .IN2(n11379), .QN(n9260) );
  AND2X1 U11657 ( .IN1(n11380), .IN2(n8508), .Q(n11379) );
  NAND2X0 U11658 ( .IN1(n11381), .IN2(n8527), .QN(n11377) );
  NAND2X0 U11659 ( .IN1(n11382), .IN2(n11383), .QN(n11381) );
  NAND2X0 U11660 ( .IN1(n11384), .IN2(g6509), .QN(n11383) );
  NAND2X0 U11661 ( .IN1(n11385), .IN2(n11386), .QN(n11382) );
  NAND4X0 U11662 ( .IN1(n7758), .IN2(n11387), .IN3(n11388), .IN4(n11389), .QN(
        n11385) );
  NAND2X0 U11663 ( .IN1(n11390), .IN2(g6163), .QN(n11389) );
  NAND2X0 U11664 ( .IN1(n11391), .IN2(n11392), .QN(n11390) );
  OR2X1 U11665 ( .IN1(n11392), .IN2(n11391), .Q(n11388) );
  NAND2X0 U11666 ( .IN1(g5817), .IN2(g5471), .QN(n11387) );
  NAND2X0 U11667 ( .IN1(n11384), .IN2(n11386), .QN(n11376) );
  NAND3X0 U11668 ( .IN1(n11393), .IN2(n11394), .IN3(n9259), .QN(n11374) );
  NOR3X0 U11669 ( .IN1(n11386), .IN2(n11384), .IN3(g6509), .QN(n9259) );
  NAND2X0 U11670 ( .IN1(n7857), .IN2(n7856), .QN(n11384) );
  NAND2X0 U11671 ( .IN1(n11395), .IN2(n11392), .QN(n11386) );
  INVX0 U11672 ( .INP(n11396), .ZN(n11392) );
  NAND2X0 U11673 ( .IN1(n11397), .IN2(n8527), .QN(n11395) );
  NAND2X0 U11674 ( .IN1(n7738), .IN2(n11391), .QN(n11397) );
  NOR2X0 U11675 ( .IN1(g5471), .IN2(g5817), .QN(n11391) );
  NAND2X0 U11676 ( .IN1(n11378), .IN2(n11380), .QN(n11394) );
  NAND2X0 U11677 ( .IN1(n7757), .IN2(n7731), .QN(n11380) );
  NAND2X0 U11678 ( .IN1(g3466), .IN2(g3115), .QN(n11393) );
  NAND2X0 U11679 ( .IN1(g113), .IN2(g2868), .QN(g31665) );
  NAND2X0 U11680 ( .IN1(g113), .IN2(g2873), .QN(g31656) );
  NAND3X0 U11681 ( .IN1(n11398), .IN2(n11399), .IN3(n11400), .QN(g30563) );
  NAND2X0 U11682 ( .IN1(n8649), .IN2(g6653), .QN(n11400) );
  NAND2X0 U11683 ( .IN1(n11401), .IN2(g6657), .QN(n11399) );
  NAND2X0 U11684 ( .IN1(n3765), .IN2(n10354), .QN(n11398) );
  NAND3X0 U11685 ( .IN1(n11402), .IN2(n11403), .IN3(n11404), .QN(g30562) );
  NAND2X0 U11686 ( .IN1(n11405), .IN2(n3765), .QN(n11404) );
  OR3X1 U11687 ( .IN1(n11405), .IN2(n8111), .IN3(n8539), .Q(n11403) );
  NOR2X0 U11688 ( .IN1(n3768), .IN2(n5646), .QN(n11405) );
  NAND2X0 U11689 ( .IN1(n8649), .IN2(g6649), .QN(n11402) );
  NAND3X0 U11690 ( .IN1(n11406), .IN2(n11407), .IN3(n11408), .QN(g30561) );
  NAND2X0 U11691 ( .IN1(n11409), .IN2(n3765), .QN(n11408) );
  INVX0 U11692 ( .INP(n10858), .ZN(n11409) );
  NAND3X0 U11693 ( .IN1(n10858), .IN2(g6597), .IN3(n8491), .QN(n11407) );
  NAND2X0 U11694 ( .IN1(n11410), .IN2(g6561), .QN(n10858) );
  NAND2X0 U11695 ( .IN1(n8649), .IN2(g6645), .QN(n11406) );
  NAND3X0 U11696 ( .IN1(n11411), .IN2(n11412), .IN3(n11413), .QN(g30560) );
  NAND2X0 U11697 ( .IN1(n11414), .IN2(n3765), .QN(n11413) );
  OR3X1 U11698 ( .IN1(n11414), .IN2(n8048), .IN3(n8540), .Q(n11412) );
  NOR2X0 U11699 ( .IN1(n3773), .IN2(n5646), .QN(n11414) );
  NAND2X0 U11700 ( .IN1(n8649), .IN2(g6641), .QN(n11411) );
  NAND3X0 U11701 ( .IN1(n11415), .IN2(n11416), .IN3(n11417), .QN(g30559) );
  NAND2X0 U11702 ( .IN1(n3774), .IN2(n11418), .QN(n11417) );
  NAND2X0 U11703 ( .IN1(n8649), .IN2(g6637), .QN(n11416) );
  NAND3X0 U11704 ( .IN1(n11419), .IN2(g6653), .IN3(n8491), .QN(n11415) );
  NAND2X0 U11705 ( .IN1(n10868), .IN2(n11418), .QN(n11419) );
  NAND3X0 U11706 ( .IN1(n11420), .IN2(n11421), .IN3(n11422), .QN(g30558) );
  NAND2X0 U11707 ( .IN1(n3774), .IN2(n10860), .QN(n11422) );
  NAND2X0 U11708 ( .IN1(n8649), .IN2(g6633), .QN(n11421) );
  NAND3X0 U11709 ( .IN1(n11423), .IN2(g6649), .IN3(n8491), .QN(n11420) );
  NAND2X0 U11710 ( .IN1(n10868), .IN2(n10860), .QN(n11423) );
  NAND3X0 U11711 ( .IN1(n11424), .IN2(n11425), .IN3(n11426), .QN(g30557) );
  NAND2X0 U11712 ( .IN1(n3774), .IN2(n11410), .QN(n11426) );
  NAND2X0 U11713 ( .IN1(n8648), .IN2(g6629), .QN(n11425) );
  NAND3X0 U11714 ( .IN1(n11427), .IN2(g6645), .IN3(n8491), .QN(n11424) );
  NAND2X0 U11715 ( .IN1(n10868), .IN2(n11410), .QN(n11427) );
  NAND3X0 U11716 ( .IN1(n11428), .IN2(n11429), .IN3(n11430), .QN(g30556) );
  NAND2X0 U11717 ( .IN1(n3774), .IN2(n11431), .QN(n11430) );
  NAND2X0 U11718 ( .IN1(n8648), .IN2(g6625), .QN(n11429) );
  NAND3X0 U11719 ( .IN1(n11432), .IN2(g6641), .IN3(n8491), .QN(n11428) );
  NAND2X0 U11720 ( .IN1(n10868), .IN2(n11431), .QN(n11432) );
  INVX0 U11721 ( .INP(n3404), .ZN(n10868) );
  NAND2X0 U11722 ( .IN1(g6555), .IN2(g6549), .QN(n3404) );
  NAND3X0 U11723 ( .IN1(n11433), .IN2(n11434), .IN3(n11435), .QN(g30555) );
  NAND2X0 U11724 ( .IN1(n3780), .IN2(n11418), .QN(n11435) );
  NAND2X0 U11725 ( .IN1(n8648), .IN2(g6621), .QN(n11434) );
  NAND3X0 U11726 ( .IN1(n11436), .IN2(g6637), .IN3(n8491), .QN(n11433) );
  NAND2X0 U11727 ( .IN1(n10873), .IN2(n11418), .QN(n11436) );
  NAND3X0 U11728 ( .IN1(n11437), .IN2(n11438), .IN3(n11439), .QN(g30554) );
  NAND2X0 U11729 ( .IN1(n3780), .IN2(n10860), .QN(n11439) );
  NAND2X0 U11730 ( .IN1(n8648), .IN2(g6617), .QN(n11438) );
  NAND3X0 U11731 ( .IN1(n11440), .IN2(g6633), .IN3(n8491), .QN(n11437) );
  NAND2X0 U11732 ( .IN1(n10873), .IN2(n10860), .QN(n11440) );
  NAND3X0 U11733 ( .IN1(n11441), .IN2(n11442), .IN3(n11443), .QN(g30553) );
  NAND2X0 U11734 ( .IN1(n3780), .IN2(n11410), .QN(n11443) );
  NAND2X0 U11735 ( .IN1(n8648), .IN2(g6613), .QN(n11442) );
  NAND3X0 U11736 ( .IN1(n11444), .IN2(g6629), .IN3(n8491), .QN(n11441) );
  NAND2X0 U11737 ( .IN1(n10873), .IN2(n11410), .QN(n11444) );
  NAND3X0 U11738 ( .IN1(n11445), .IN2(n11446), .IN3(n11447), .QN(g30552) );
  NAND2X0 U11739 ( .IN1(n3780), .IN2(n11431), .QN(n11447) );
  NAND2X0 U11740 ( .IN1(n8648), .IN2(g6609), .QN(n11446) );
  NAND3X0 U11741 ( .IN1(n11448), .IN2(g6625), .IN3(n8491), .QN(n11445) );
  NAND2X0 U11742 ( .IN1(n10873), .IN2(n11431), .QN(n11448) );
  INVX0 U11743 ( .INP(n3406), .ZN(n10873) );
  NAND2X0 U11744 ( .IN1(n5571), .IN2(g6555), .QN(n3406) );
  NAND3X0 U11745 ( .IN1(n11449), .IN2(n11450), .IN3(n11451), .QN(g30551) );
  NAND2X0 U11746 ( .IN1(n3785), .IN2(n11418), .QN(n11451) );
  NAND2X0 U11747 ( .IN1(n8648), .IN2(g6601), .QN(n11450) );
  NAND3X0 U11748 ( .IN1(n11452), .IN2(g6621), .IN3(n8491), .QN(n11449) );
  NAND2X0 U11749 ( .IN1(n11453), .IN2(n11418), .QN(n11452) );
  INVX0 U11750 ( .INP(n3776), .ZN(n11418) );
  NAND3X0 U11751 ( .IN1(n11454), .IN2(n11455), .IN3(n11456), .QN(g30550) );
  NAND2X0 U11752 ( .IN1(n3785), .IN2(n10860), .QN(n11456) );
  NAND2X0 U11753 ( .IN1(n8647), .IN2(g6593), .QN(n11455) );
  NAND3X0 U11754 ( .IN1(n11457), .IN2(g6617), .IN3(n8491), .QN(n11454) );
  NAND2X0 U11755 ( .IN1(n11453), .IN2(n10860), .QN(n11457) );
  INVX0 U11756 ( .INP(n3768), .ZN(n10860) );
  NAND2X0 U11757 ( .IN1(n5386), .IN2(g6573), .QN(n3768) );
  NAND3X0 U11758 ( .IN1(n11458), .IN2(n11459), .IN3(n11460), .QN(g30549) );
  NAND2X0 U11759 ( .IN1(n3785), .IN2(n11410), .QN(n11460) );
  NAND2X0 U11760 ( .IN1(test_so71), .IN2(n8543), .QN(n11459) );
  NAND3X0 U11761 ( .IN1(n11461), .IN2(g6613), .IN3(n8491), .QN(n11458) );
  NAND2X0 U11762 ( .IN1(n11453), .IN2(n11410), .QN(n11461) );
  INVX0 U11763 ( .INP(n3770), .ZN(n11410) );
  NAND2X0 U11764 ( .IN1(n5563), .IN2(g6565), .QN(n3770) );
  NAND3X0 U11765 ( .IN1(n11462), .IN2(n11463), .IN3(n11464), .QN(g30548) );
  NAND2X0 U11766 ( .IN1(n3785), .IN2(n11431), .QN(n11464) );
  NAND2X0 U11767 ( .IN1(n8647), .IN2(g6581), .QN(n11463) );
  NAND3X0 U11768 ( .IN1(n11465), .IN2(g6609), .IN3(n8491), .QN(n11462) );
  NAND2X0 U11769 ( .IN1(n11453), .IN2(n11431), .QN(n11465) );
  INVX0 U11770 ( .INP(n3773), .ZN(n11431) );
  NAND2X0 U11771 ( .IN1(n5563), .IN2(n5386), .QN(n3773) );
  INVX0 U11772 ( .INP(n3407), .ZN(n11453) );
  NAND2X0 U11773 ( .IN1(n8141), .IN2(g6549), .QN(n3407) );
  NAND3X0 U11774 ( .IN1(n11466), .IN2(n11467), .IN3(n11468), .QN(g30547) );
  NAND2X0 U11775 ( .IN1(n8647), .IN2(g6605), .QN(n11468) );
  OR3X1 U11776 ( .IN1(n8529), .IN2(n8022), .IN3(n3790), .Q(n11467) );
  NAND2X0 U11777 ( .IN1(n3790), .IN2(n3765), .QN(n11466) );
  NAND3X0 U11778 ( .IN1(n11469), .IN2(n11470), .IN3(n11471), .QN(g30546) );
  NAND2X0 U11779 ( .IN1(n8647), .IN2(g6597), .QN(n11471) );
  OR3X1 U11780 ( .IN1(n8536), .IN2(n8113), .IN3(n3793), .Q(n11470) );
  NAND2X0 U11781 ( .IN1(n3793), .IN2(n3765), .QN(n11469) );
  NAND3X0 U11782 ( .IN1(n11472), .IN2(n11473), .IN3(n11474), .QN(g30545) );
  NAND2X0 U11783 ( .IN1(n8647), .IN2(g6589), .QN(n11474) );
  NAND3X0 U11784 ( .IN1(test_so71), .IN2(n8482), .IN3(n11475), .QN(n11473) );
  INVX0 U11785 ( .INP(n3795), .ZN(n11475) );
  NAND2X0 U11786 ( .IN1(n3795), .IN2(n3765), .QN(n11472) );
  NAND3X0 U11787 ( .IN1(n11476), .IN2(n11477), .IN3(n11478), .QN(g30544) );
  NAND2X0 U11788 ( .IN1(n8647), .IN2(g6573), .QN(n11478) );
  OR3X1 U11789 ( .IN1(n8534), .IN2(n8049), .IN3(n3797), .Q(n11477) );
  NAND2X0 U11790 ( .IN1(n3797), .IN2(n3765), .QN(n11476) );
  NOR2X0 U11791 ( .IN1(g6549), .IN2(n10865), .QN(g30543) );
  NAND3X0 U11792 ( .IN1(n10856), .IN2(n8483), .IN3(n5646), .QN(n10865) );
  NAND2X0 U11793 ( .IN1(n3799), .IN2(n9602), .QN(n10856) );
  NAND3X0 U11794 ( .IN1(n11479), .IN2(n11480), .IN3(n11481), .QN(g30542) );
  NAND2X0 U11795 ( .IN1(n8647), .IN2(g6307), .QN(n11481) );
  NAND2X0 U11796 ( .IN1(n11482), .IN2(g6311), .QN(n11480) );
  NAND2X0 U11797 ( .IN1(n11483), .IN2(n3765), .QN(n11479) );
  NAND3X0 U11798 ( .IN1(n11484), .IN2(n11485), .IN3(n11486), .QN(g30541) );
  NAND2X0 U11799 ( .IN1(n11487), .IN2(n3765), .QN(n11486) );
  OR3X1 U11800 ( .IN1(n11487), .IN2(n8119), .IN3(n8541), .Q(n11485) );
  NOR2X0 U11801 ( .IN1(n3802), .IN2(n5651), .QN(n11487) );
  NAND2X0 U11802 ( .IN1(n8646), .IN2(g6303), .QN(n11484) );
  NAND3X0 U11803 ( .IN1(n11488), .IN2(n11489), .IN3(n11490), .QN(g30540) );
  NAND2X0 U11804 ( .IN1(n11491), .IN2(n3765), .QN(n11490) );
  INVX0 U11805 ( .INP(n10879), .ZN(n11491) );
  NAND3X0 U11806 ( .IN1(n10879), .IN2(g6251), .IN3(n8492), .QN(n11489) );
  NAND2X0 U11807 ( .IN1(n11492), .IN2(g6215), .QN(n10879) );
  NAND2X0 U11808 ( .IN1(n8646), .IN2(g6299), .QN(n11488) );
  NAND3X0 U11809 ( .IN1(n11493), .IN2(n11494), .IN3(n11495), .QN(g30539) );
  NAND2X0 U11810 ( .IN1(n11496), .IN2(n3765), .QN(n11495) );
  OR3X1 U11811 ( .IN1(n11496), .IN2(n8052), .IN3(n8540), .Q(n11494) );
  NOR2X0 U11812 ( .IN1(n3807), .IN2(n5651), .QN(n11496) );
  NAND2X0 U11813 ( .IN1(n8646), .IN2(g6295), .QN(n11493) );
  NAND3X0 U11814 ( .IN1(n11497), .IN2(n11498), .IN3(n11499), .QN(g30538) );
  NAND2X0 U11815 ( .IN1(n3808), .IN2(n11500), .QN(n11499) );
  NAND2X0 U11816 ( .IN1(n8646), .IN2(g6291), .QN(n11498) );
  NAND3X0 U11817 ( .IN1(n11501), .IN2(g6307), .IN3(n8492), .QN(n11497) );
  NAND2X0 U11818 ( .IN1(n10889), .IN2(n11500), .QN(n11501) );
  NAND3X0 U11819 ( .IN1(n11502), .IN2(n11503), .IN3(n11504), .QN(g30537) );
  NAND2X0 U11820 ( .IN1(n3808), .IN2(n10881), .QN(n11504) );
  NAND2X0 U11821 ( .IN1(n8646), .IN2(g6287), .QN(n11503) );
  NAND3X0 U11822 ( .IN1(n11505), .IN2(g6303), .IN3(n8492), .QN(n11502) );
  NAND2X0 U11823 ( .IN1(n10889), .IN2(n10881), .QN(n11505) );
  NAND3X0 U11824 ( .IN1(n11506), .IN2(n11507), .IN3(n11508), .QN(g30536) );
  NAND2X0 U11825 ( .IN1(n3808), .IN2(n11492), .QN(n11508) );
  NAND2X0 U11826 ( .IN1(n8646), .IN2(g6283), .QN(n11507) );
  NAND3X0 U11827 ( .IN1(n11509), .IN2(g6299), .IN3(n8492), .QN(n11506) );
  NAND2X0 U11828 ( .IN1(n10889), .IN2(n11492), .QN(n11509) );
  NAND3X0 U11829 ( .IN1(n11510), .IN2(n11511), .IN3(n11512), .QN(g30535) );
  NAND2X0 U11830 ( .IN1(n3808), .IN2(n11513), .QN(n11512) );
  NAND2X0 U11831 ( .IN1(n8646), .IN2(g6279), .QN(n11511) );
  NAND3X0 U11832 ( .IN1(n11514), .IN2(g6295), .IN3(n8492), .QN(n11510) );
  NAND2X0 U11833 ( .IN1(n10889), .IN2(n11513), .QN(n11514) );
  INVX0 U11834 ( .INP(n3414), .ZN(n10889) );
  NAND2X0 U11835 ( .IN1(g6209), .IN2(g6203), .QN(n3414) );
  NAND3X0 U11836 ( .IN1(n11515), .IN2(n11516), .IN3(n11517), .QN(g30534) );
  NAND2X0 U11837 ( .IN1(n3814), .IN2(n11500), .QN(n11517) );
  NAND2X0 U11838 ( .IN1(n8645), .IN2(g6275), .QN(n11516) );
  NAND3X0 U11839 ( .IN1(n11518), .IN2(g6291), .IN3(n8492), .QN(n11515) );
  NAND2X0 U11840 ( .IN1(n10894), .IN2(n11500), .QN(n11518) );
  NAND3X0 U11841 ( .IN1(n11519), .IN2(n11520), .IN3(n11521), .QN(g30533) );
  NAND2X0 U11842 ( .IN1(n3814), .IN2(n10881), .QN(n11521) );
  NAND2X0 U11843 ( .IN1(n8645), .IN2(g6271), .QN(n11520) );
  NAND3X0 U11844 ( .IN1(n11522), .IN2(g6287), .IN3(n8492), .QN(n11519) );
  NAND2X0 U11845 ( .IN1(n10894), .IN2(n10881), .QN(n11522) );
  NAND3X0 U11846 ( .IN1(n11523), .IN2(n11524), .IN3(n11525), .QN(g30532) );
  NAND2X0 U11847 ( .IN1(n3814), .IN2(n11492), .QN(n11525) );
  NAND2X0 U11848 ( .IN1(n8645), .IN2(g6267), .QN(n11524) );
  NAND3X0 U11849 ( .IN1(n11526), .IN2(g6283), .IN3(n8487), .QN(n11523) );
  NAND2X0 U11850 ( .IN1(n10894), .IN2(n11492), .QN(n11526) );
  NAND3X0 U11851 ( .IN1(n11527), .IN2(n11528), .IN3(n11529), .QN(g30531) );
  NAND2X0 U11852 ( .IN1(n3814), .IN2(n11513), .QN(n11529) );
  NAND2X0 U11853 ( .IN1(n8645), .IN2(g6263), .QN(n11528) );
  NAND3X0 U11854 ( .IN1(n11530), .IN2(g6279), .IN3(n8496), .QN(n11527) );
  NAND2X0 U11855 ( .IN1(n10894), .IN2(n11513), .QN(n11530) );
  INVX0 U11856 ( .INP(n3416), .ZN(n10894) );
  NAND2X0 U11857 ( .IN1(n5574), .IN2(g6209), .QN(n3416) );
  NAND3X0 U11858 ( .IN1(n11531), .IN2(n11532), .IN3(n11533), .QN(g30530) );
  NAND2X0 U11859 ( .IN1(n3819), .IN2(n11500), .QN(n11533) );
  NAND2X0 U11860 ( .IN1(n8645), .IN2(g6255), .QN(n11532) );
  NAND3X0 U11861 ( .IN1(n11534), .IN2(g6275), .IN3(n8490), .QN(n11531) );
  NAND2X0 U11862 ( .IN1(n11535), .IN2(n11500), .QN(n11534) );
  NAND3X0 U11863 ( .IN1(n11536), .IN2(n11537), .IN3(n11538), .QN(g30529) );
  NAND2X0 U11864 ( .IN1(n3819), .IN2(n10881), .QN(n11538) );
  NAND2X0 U11865 ( .IN1(n8645), .IN2(g6247), .QN(n11537) );
  NAND3X0 U11866 ( .IN1(n11539), .IN2(g6271), .IN3(n8490), .QN(n11536) );
  NAND2X0 U11867 ( .IN1(n11535), .IN2(n10881), .QN(n11539) );
  INVX0 U11868 ( .INP(n3802), .ZN(n10881) );
  NAND2X0 U11869 ( .IN1(n5385), .IN2(g6227), .QN(n3802) );
  NAND3X0 U11870 ( .IN1(n11540), .IN2(n11541), .IN3(n11542), .QN(g30528) );
  NAND2X0 U11871 ( .IN1(n3819), .IN2(n11492), .QN(n11542) );
  NAND2X0 U11872 ( .IN1(n8645), .IN2(g6239), .QN(n11541) );
  NAND3X0 U11873 ( .IN1(n11543), .IN2(g6267), .IN3(n8490), .QN(n11540) );
  NAND2X0 U11874 ( .IN1(n11535), .IN2(n11492), .QN(n11543) );
  INVX0 U11875 ( .INP(n3804), .ZN(n11492) );
  NAND2X0 U11876 ( .IN1(n5568), .IN2(g6219), .QN(n3804) );
  NAND3X0 U11877 ( .IN1(n11544), .IN2(n11545), .IN3(n11546), .QN(g30527) );
  NAND2X0 U11878 ( .IN1(n3819), .IN2(n11513), .QN(n11546) );
  NAND2X0 U11879 ( .IN1(n8644), .IN2(g6235), .QN(n11545) );
  NAND3X0 U11880 ( .IN1(n11547), .IN2(g6263), .IN3(n8490), .QN(n11544) );
  NAND2X0 U11881 ( .IN1(n11535), .IN2(n11513), .QN(n11547) );
  INVX0 U11882 ( .INP(n3807), .ZN(n11513) );
  NAND2X0 U11883 ( .IN1(n5568), .IN2(n5385), .QN(n3807) );
  INVX0 U11884 ( .INP(n3417), .ZN(n11535) );
  NAND2X0 U11885 ( .IN1(n8144), .IN2(g6203), .QN(n3417) );
  NAND3X0 U11886 ( .IN1(n11548), .IN2(n11549), .IN3(n11550), .QN(g30526) );
  NAND2X0 U11887 ( .IN1(n8644), .IN2(g6259), .QN(n11550) );
  OR3X1 U11888 ( .IN1(n8536), .IN2(n8028), .IN3(n3824), .Q(n11549) );
  NAND2X0 U11889 ( .IN1(n3824), .IN2(n3765), .QN(n11548) );
  NAND3X0 U11890 ( .IN1(n11551), .IN2(n11552), .IN3(n11553), .QN(g30525) );
  NAND2X0 U11891 ( .IN1(n8644), .IN2(g6251), .QN(n11553) );
  OR3X1 U11892 ( .IN1(n8533), .IN2(n8121), .IN3(n3827), .Q(n11552) );
  NAND2X0 U11893 ( .IN1(n3827), .IN2(n3765), .QN(n11551) );
  NAND3X0 U11894 ( .IN1(n11554), .IN2(n11555), .IN3(n11556), .QN(g30524) );
  NAND2X0 U11895 ( .IN1(n8644), .IN2(g6243), .QN(n11556) );
  OR3X1 U11896 ( .IN1(n8535), .IN2(n7895), .IN3(n3829), .Q(n11555) );
  NAND2X0 U11897 ( .IN1(n3829), .IN2(n3765), .QN(n11554) );
  NAND3X0 U11898 ( .IN1(n11557), .IN2(n11558), .IN3(n11559), .QN(g30523) );
  NAND2X0 U11899 ( .IN1(n8644), .IN2(g6227), .QN(n11559) );
  OR3X1 U11900 ( .IN1(n8535), .IN2(n8053), .IN3(n3831), .Q(n11558) );
  NAND2X0 U11901 ( .IN1(n3831), .IN2(n3765), .QN(n11557) );
  NOR2X0 U11902 ( .IN1(g6203), .IN2(n10886), .QN(g30522) );
  NAND3X0 U11903 ( .IN1(n10877), .IN2(n8482), .IN3(n5651), .QN(n10886) );
  NAND3X0 U11904 ( .IN1(g4093), .IN2(g4087), .IN3(n3833), .QN(n10877) );
  NAND3X0 U11905 ( .IN1(n11560), .IN2(n11561), .IN3(n11562), .QN(g30521) );
  NAND2X0 U11906 ( .IN1(n8644), .IN2(g5961), .QN(n11562) );
  NAND2X0 U11907 ( .IN1(test_so13), .IN2(n11563), .QN(n11561) );
  NAND2X0 U11908 ( .IN1(n11564), .IN2(n3765), .QN(n11560) );
  NAND3X0 U11909 ( .IN1(n11565), .IN2(n11566), .IN3(n11567), .QN(g30520) );
  NAND2X0 U11910 ( .IN1(n11568), .IN2(n3765), .QN(n11567) );
  OR3X1 U11911 ( .IN1(n11568), .IN2(n8099), .IN3(n8540), .Q(n11566) );
  NOR2X0 U11912 ( .IN1(n3836), .IN2(n5649), .QN(n11568) );
  NAND2X0 U11913 ( .IN1(n8644), .IN2(g5957), .QN(n11565) );
  NAND3X0 U11914 ( .IN1(n11569), .IN2(n11570), .IN3(n11571), .QN(g30519) );
  NAND2X0 U11915 ( .IN1(n11572), .IN2(n3765), .QN(n11571) );
  INVX0 U11916 ( .INP(n10900), .ZN(n11572) );
  NAND3X0 U11917 ( .IN1(n10900), .IN2(g5905), .IN3(n8490), .QN(n11570) );
  NAND2X0 U11918 ( .IN1(n11573), .IN2(g5869), .QN(n10900) );
  NAND2X0 U11919 ( .IN1(n8643), .IN2(g5953), .QN(n11569) );
  NAND3X0 U11920 ( .IN1(n11574), .IN2(n11575), .IN3(n11576), .QN(g30518) );
  NAND2X0 U11921 ( .IN1(n11577), .IN2(n3765), .QN(n11576) );
  OR3X1 U11922 ( .IN1(n11577), .IN2(n8043), .IN3(n8541), .Q(n11575) );
  NOR2X0 U11923 ( .IN1(n3841), .IN2(n5649), .QN(n11577) );
  NAND2X0 U11924 ( .IN1(n8643), .IN2(g5949), .QN(n11574) );
  NAND3X0 U11925 ( .IN1(n11578), .IN2(n11579), .IN3(n11580), .QN(g30517) );
  NAND2X0 U11926 ( .IN1(n3842), .IN2(n11581), .QN(n11580) );
  NAND2X0 U11927 ( .IN1(n8643), .IN2(g5945), .QN(n11579) );
  NAND3X0 U11928 ( .IN1(n11582), .IN2(g5961), .IN3(n8489), .QN(n11578) );
  NAND2X0 U11929 ( .IN1(n10910), .IN2(n11581), .QN(n11582) );
  NAND3X0 U11930 ( .IN1(n11583), .IN2(n11584), .IN3(n11585), .QN(g30516) );
  NAND2X0 U11931 ( .IN1(n3842), .IN2(n10902), .QN(n11585) );
  NAND2X0 U11932 ( .IN1(n8643), .IN2(g5941), .QN(n11584) );
  NAND3X0 U11933 ( .IN1(n11586), .IN2(g5957), .IN3(n8489), .QN(n11583) );
  NAND2X0 U11934 ( .IN1(n10910), .IN2(n10902), .QN(n11586) );
  NAND3X0 U11935 ( .IN1(n11587), .IN2(n11588), .IN3(n11589), .QN(g30515) );
  NAND2X0 U11936 ( .IN1(n3842), .IN2(n11573), .QN(n11589) );
  NAND2X0 U11937 ( .IN1(n8643), .IN2(g5937), .QN(n11588) );
  NAND3X0 U11938 ( .IN1(n11590), .IN2(g5953), .IN3(n8489), .QN(n11587) );
  NAND2X0 U11939 ( .IN1(n10910), .IN2(n11573), .QN(n11590) );
  NAND3X0 U11940 ( .IN1(n11591), .IN2(n11592), .IN3(n11593), .QN(g30514) );
  NAND2X0 U11941 ( .IN1(n3842), .IN2(n11594), .QN(n11593) );
  NAND2X0 U11942 ( .IN1(n8643), .IN2(g5933), .QN(n11592) );
  NAND3X0 U11943 ( .IN1(n11595), .IN2(g5949), .IN3(n8489), .QN(n11591) );
  NAND2X0 U11944 ( .IN1(n10910), .IN2(n11594), .QN(n11595) );
  INVX0 U11945 ( .INP(n3424), .ZN(n10910) );
  NAND2X0 U11946 ( .IN1(g5863), .IN2(g5857), .QN(n3424) );
  NAND3X0 U11947 ( .IN1(n11596), .IN2(n11597), .IN3(n11598), .QN(g30513) );
  NAND2X0 U11948 ( .IN1(n3848), .IN2(n11581), .QN(n11598) );
  NAND2X0 U11949 ( .IN1(n8643), .IN2(g5929), .QN(n11597) );
  NAND3X0 U11950 ( .IN1(n11599), .IN2(g5945), .IN3(n8489), .QN(n11596) );
  NAND2X0 U11951 ( .IN1(n10915), .IN2(n11581), .QN(n11599) );
  NAND3X0 U11952 ( .IN1(n11600), .IN2(n11601), .IN3(n11602), .QN(g30512) );
  NAND2X0 U11953 ( .IN1(n3848), .IN2(n10902), .QN(n11602) );
  NAND2X0 U11954 ( .IN1(n8642), .IN2(g5925), .QN(n11601) );
  NAND3X0 U11955 ( .IN1(n11603), .IN2(g5941), .IN3(n8489), .QN(n11600) );
  NAND2X0 U11956 ( .IN1(n10915), .IN2(n10902), .QN(n11603) );
  NAND3X0 U11957 ( .IN1(n11604), .IN2(n11605), .IN3(n11606), .QN(g30511) );
  NAND2X0 U11958 ( .IN1(n3848), .IN2(n11573), .QN(n11606) );
  NAND2X0 U11959 ( .IN1(n8642), .IN2(g5921), .QN(n11605) );
  NAND3X0 U11960 ( .IN1(n11607), .IN2(g5937), .IN3(n8489), .QN(n11604) );
  NAND2X0 U11961 ( .IN1(n10915), .IN2(n11573), .QN(n11607) );
  NAND3X0 U11962 ( .IN1(n11608), .IN2(n11609), .IN3(n11610), .QN(g30510) );
  NAND2X0 U11963 ( .IN1(n3848), .IN2(n11594), .QN(n11610) );
  NAND2X0 U11964 ( .IN1(test_so28), .IN2(n8660), .QN(n11609) );
  NAND3X0 U11965 ( .IN1(n11611), .IN2(g5933), .IN3(n8489), .QN(n11608) );
  NAND2X0 U11966 ( .IN1(n10915), .IN2(n11594), .QN(n11611) );
  INVX0 U11967 ( .INP(n3426), .ZN(n10915) );
  NAND2X0 U11968 ( .IN1(n5573), .IN2(g5863), .QN(n3426) );
  NAND3X0 U11969 ( .IN1(n11612), .IN2(n11613), .IN3(n11614), .QN(g30509) );
  NAND2X0 U11970 ( .IN1(n3853), .IN2(n11581), .QN(n11614) );
  NAND2X0 U11971 ( .IN1(n8642), .IN2(g5909), .QN(n11613) );
  NAND3X0 U11972 ( .IN1(n11615), .IN2(g5929), .IN3(n8489), .QN(n11612) );
  NAND2X0 U11973 ( .IN1(n11616), .IN2(n11581), .QN(n11615) );
  NAND3X0 U11974 ( .IN1(n11617), .IN2(n11618), .IN3(n11619), .QN(g30508) );
  NAND2X0 U11975 ( .IN1(n3853), .IN2(n10902), .QN(n11619) );
  NAND2X0 U11976 ( .IN1(n8642), .IN2(g5901), .QN(n11618) );
  NAND3X0 U11977 ( .IN1(n11620), .IN2(g5925), .IN3(n8488), .QN(n11617) );
  NAND2X0 U11978 ( .IN1(n11616), .IN2(n10902), .QN(n11620) );
  INVX0 U11979 ( .INP(n3836), .ZN(n10902) );
  NAND2X0 U11980 ( .IN1(n5388), .IN2(test_so36), .QN(n3836) );
  NAND3X0 U11981 ( .IN1(n11621), .IN2(n11622), .IN3(n11623), .QN(g30507) );
  NAND2X0 U11982 ( .IN1(n3853), .IN2(n11573), .QN(n11623) );
  NAND2X0 U11983 ( .IN1(n8642), .IN2(g5893), .QN(n11622) );
  NAND3X0 U11984 ( .IN1(n11624), .IN2(g5921), .IN3(n8488), .QN(n11621) );
  NAND2X0 U11985 ( .IN1(n11616), .IN2(n11573), .QN(n11624) );
  INVX0 U11986 ( .INP(n3838), .ZN(n11573) );
  NAND2X0 U11987 ( .IN1(n8217), .IN2(g5873), .QN(n3838) );
  NAND3X0 U11988 ( .IN1(n11625), .IN2(n11626), .IN3(n11627), .QN(g30506) );
  NAND2X0 U11989 ( .IN1(n3853), .IN2(n11594), .QN(n11627) );
  NAND2X0 U11990 ( .IN1(n8642), .IN2(g5889), .QN(n11626) );
  NAND3X0 U11991 ( .IN1(test_so28), .IN2(n11628), .IN3(n8488), .QN(n11625) );
  NAND2X0 U11992 ( .IN1(n11616), .IN2(n11594), .QN(n11628) );
  INVX0 U11993 ( .INP(n3841), .ZN(n11594) );
  NAND2X0 U11994 ( .IN1(n5388), .IN2(n8217), .QN(n3841) );
  INVX0 U11995 ( .INP(n3427), .ZN(n11616) );
  NAND2X0 U11996 ( .IN1(n8143), .IN2(g5857), .QN(n3427) );
  NAND3X0 U11997 ( .IN1(n11629), .IN2(n11630), .IN3(n11631), .QN(g30505) );
  NAND2X0 U11998 ( .IN1(n8642), .IN2(g5913), .QN(n11631) );
  OR3X1 U11999 ( .IN1(n8534), .IN2(n8013), .IN3(n3858), .Q(n11630) );
  NAND2X0 U12000 ( .IN1(n3858), .IN2(n3765), .QN(n11629) );
  NAND3X0 U12001 ( .IN1(n11632), .IN2(n11633), .IN3(n11634), .QN(g30504) );
  NAND2X0 U12002 ( .IN1(n8641), .IN2(g5905), .QN(n11634) );
  OR3X1 U12003 ( .IN1(n8534), .IN2(n8101), .IN3(n3861), .Q(n11633) );
  NAND2X0 U12004 ( .IN1(n3861), .IN2(n3765), .QN(n11632) );
  NAND3X0 U12005 ( .IN1(n11635), .IN2(n11636), .IN3(n11637), .QN(g30503) );
  NAND2X0 U12006 ( .IN1(n8641), .IN2(g5897), .QN(n11637) );
  OR3X1 U12007 ( .IN1(n8532), .IN2(n7901), .IN3(n3863), .Q(n11636) );
  NAND2X0 U12008 ( .IN1(n3863), .IN2(n3765), .QN(n11635) );
  NAND3X0 U12009 ( .IN1(n11638), .IN2(n11639), .IN3(n11640), .QN(g30502) );
  NAND2X0 U12010 ( .IN1(test_so36), .IN2(n8567), .QN(n11640) );
  OR3X1 U12011 ( .IN1(n8533), .IN2(n8044), .IN3(n3865), .Q(n11639) );
  NAND2X0 U12012 ( .IN1(n3865), .IN2(n3765), .QN(n11638) );
  NOR2X0 U12013 ( .IN1(g5857), .IN2(n10907), .QN(g30501) );
  NAND3X0 U12014 ( .IN1(n10898), .IN2(n8484), .IN3(n5649), .QN(n10907) );
  NAND3X0 U12015 ( .IN1(n5480), .IN2(g4093), .IN3(n3833), .QN(n10898) );
  NAND3X0 U12016 ( .IN1(n11641), .IN2(n11642), .IN3(n11643), .QN(g30500) );
  NAND2X0 U12017 ( .IN1(n8641), .IN2(g5615), .QN(n11643) );
  NAND2X0 U12018 ( .IN1(n11644), .IN2(g5619), .QN(n11642) );
  NAND2X0 U12019 ( .IN1(n3765), .IN2(n10339), .QN(n11641) );
  NAND3X0 U12020 ( .IN1(n11645), .IN2(n11646), .IN3(n11647), .QN(g30499) );
  NAND2X0 U12021 ( .IN1(n11648), .IN2(n3765), .QN(n11647) );
  OR3X1 U12022 ( .IN1(n11648), .IN2(n8103), .IN3(n8542), .Q(n11646) );
  NOR2X0 U12023 ( .IN1(n3869), .IN2(n5647), .QN(n11648) );
  NAND2X0 U12024 ( .IN1(n8641), .IN2(g5611), .QN(n11645) );
  NAND3X0 U12025 ( .IN1(n11649), .IN2(n11650), .IN3(n11651), .QN(g30498) );
  NAND2X0 U12026 ( .IN1(n11652), .IN2(n3765), .QN(n11651) );
  INVX0 U12027 ( .INP(n10921), .ZN(n11652) );
  NAND3X0 U12028 ( .IN1(test_so6), .IN2(n10921), .IN3(n8488), .QN(n11650) );
  NAND2X0 U12029 ( .IN1(n11653), .IN2(g5523), .QN(n10921) );
  NAND2X0 U12030 ( .IN1(n8641), .IN2(g5607), .QN(n11649) );
  NAND3X0 U12031 ( .IN1(n11654), .IN2(n11655), .IN3(n11656), .QN(g30497) );
  NAND2X0 U12032 ( .IN1(n11657), .IN2(n3765), .QN(n11656) );
  OR3X1 U12033 ( .IN1(n11657), .IN2(n8045), .IN3(n8543), .Q(n11655) );
  NOR2X0 U12034 ( .IN1(n3874), .IN2(n5647), .QN(n11657) );
  NAND2X0 U12035 ( .IN1(n8641), .IN2(g5603), .QN(n11654) );
  NAND3X0 U12036 ( .IN1(n11658), .IN2(n11659), .IN3(n11660), .QN(g30496) );
  NAND2X0 U12037 ( .IN1(n3875), .IN2(n11661), .QN(n11660) );
  NAND2X0 U12038 ( .IN1(n8641), .IN2(g5599), .QN(n11659) );
  NAND3X0 U12039 ( .IN1(n11662), .IN2(g5615), .IN3(n8488), .QN(n11658) );
  NAND2X0 U12040 ( .IN1(n10931), .IN2(n11661), .QN(n11662) );
  NAND3X0 U12041 ( .IN1(n11663), .IN2(n11664), .IN3(n11665), .QN(g30495) );
  NAND2X0 U12042 ( .IN1(n3875), .IN2(n10923), .QN(n11665) );
  NAND2X0 U12043 ( .IN1(n8640), .IN2(g5595), .QN(n11664) );
  NAND3X0 U12044 ( .IN1(n11666), .IN2(g5611), .IN3(n8488), .QN(n11663) );
  NAND2X0 U12045 ( .IN1(n10931), .IN2(n10923), .QN(n11666) );
  NAND3X0 U12046 ( .IN1(n11667), .IN2(n11668), .IN3(n11669), .QN(g30494) );
  NAND2X0 U12047 ( .IN1(n3875), .IN2(n11653), .QN(n11669) );
  NAND2X0 U12048 ( .IN1(test_so5), .IN2(n8659), .QN(n11668) );
  NAND3X0 U12049 ( .IN1(n11670), .IN2(g5607), .IN3(n8488), .QN(n11667) );
  NAND2X0 U12050 ( .IN1(n10931), .IN2(n11653), .QN(n11670) );
  NAND3X0 U12051 ( .IN1(n11671), .IN2(n11672), .IN3(n11673), .QN(g30493) );
  NAND2X0 U12052 ( .IN1(n3875), .IN2(n11674), .QN(n11673) );
  NAND2X0 U12053 ( .IN1(n8640), .IN2(g5587), .QN(n11672) );
  NAND3X0 U12054 ( .IN1(n11675), .IN2(g5603), .IN3(n8488), .QN(n11671) );
  NAND2X0 U12055 ( .IN1(n10931), .IN2(n11674), .QN(n11675) );
  INVX0 U12056 ( .INP(n3434), .ZN(n10931) );
  NAND2X0 U12057 ( .IN1(g5517), .IN2(g5511), .QN(n3434) );
  NAND3X0 U12058 ( .IN1(n11676), .IN2(n11677), .IN3(n11678), .QN(g30492) );
  NAND2X0 U12059 ( .IN1(n3881), .IN2(n11661), .QN(n11678) );
  NAND2X0 U12060 ( .IN1(n8640), .IN2(g5583), .QN(n11677) );
  NAND3X0 U12061 ( .IN1(n11679), .IN2(g5599), .IN3(n8488), .QN(n11676) );
  NAND2X0 U12062 ( .IN1(n10936), .IN2(n11661), .QN(n11679) );
  NAND3X0 U12063 ( .IN1(n11680), .IN2(n11681), .IN3(n11682), .QN(g30491) );
  NAND2X0 U12064 ( .IN1(n3881), .IN2(n10923), .QN(n11682) );
  NAND2X0 U12065 ( .IN1(n8640), .IN2(g5579), .QN(n11681) );
  NAND3X0 U12066 ( .IN1(n11683), .IN2(g5595), .IN3(n8488), .QN(n11680) );
  NAND2X0 U12067 ( .IN1(n10936), .IN2(n10923), .QN(n11683) );
  NAND3X0 U12068 ( .IN1(n11684), .IN2(n11685), .IN3(n11686), .QN(g30490) );
  NAND2X0 U12069 ( .IN1(n3881), .IN2(n11653), .QN(n11686) );
  NAND2X0 U12070 ( .IN1(n8640), .IN2(g5575), .QN(n11685) );
  NAND3X0 U12071 ( .IN1(test_so5), .IN2(n11687), .IN3(n8488), .QN(n11684) );
  NAND2X0 U12072 ( .IN1(n10936), .IN2(n11653), .QN(n11687) );
  NAND3X0 U12073 ( .IN1(n11688), .IN2(n11689), .IN3(n11690), .QN(g30489) );
  NAND2X0 U12074 ( .IN1(n3881), .IN2(n11674), .QN(n11690) );
  NAND2X0 U12075 ( .IN1(n8640), .IN2(g5571), .QN(n11689) );
  NAND3X0 U12076 ( .IN1(n11691), .IN2(g5587), .IN3(n8488), .QN(n11688) );
  NAND2X0 U12077 ( .IN1(n10936), .IN2(n11674), .QN(n11691) );
  INVX0 U12078 ( .INP(n3436), .ZN(n10936) );
  NAND2X0 U12079 ( .IN1(n5575), .IN2(g5517), .QN(n3436) );
  NAND3X0 U12080 ( .IN1(n11692), .IN2(n11693), .IN3(n11694), .QN(g30488) );
  NAND2X0 U12081 ( .IN1(n3886), .IN2(n11661), .QN(n11694) );
  NAND2X0 U12082 ( .IN1(n8640), .IN2(g5563), .QN(n11693) );
  NAND3X0 U12083 ( .IN1(n11695), .IN2(g5583), .IN3(n8487), .QN(n11692) );
  NAND2X0 U12084 ( .IN1(n11696), .IN2(n11661), .QN(n11695) );
  INVX0 U12085 ( .INP(n3877), .ZN(n11661) );
  NAND3X0 U12086 ( .IN1(n11697), .IN2(n11698), .IN3(n11699), .QN(g30487) );
  NAND2X0 U12087 ( .IN1(n3886), .IN2(n10923), .QN(n11699) );
  NAND2X0 U12088 ( .IN1(n8639), .IN2(g5555), .QN(n11698) );
  NAND3X0 U12089 ( .IN1(n11700), .IN2(g5579), .IN3(n8487), .QN(n11697) );
  NAND2X0 U12090 ( .IN1(n11696), .IN2(n10923), .QN(n11700) );
  INVX0 U12091 ( .INP(n3869), .ZN(n10923) );
  NAND2X0 U12092 ( .IN1(n5389), .IN2(g5535), .QN(n3869) );
  NAND3X0 U12093 ( .IN1(n11701), .IN2(n11702), .IN3(n11703), .QN(g30486) );
  NAND2X0 U12094 ( .IN1(n3886), .IN2(n11653), .QN(n11703) );
  NAND2X0 U12095 ( .IN1(n8639), .IN2(g5547), .QN(n11702) );
  NAND3X0 U12096 ( .IN1(n11704), .IN2(g5575), .IN3(n8487), .QN(n11701) );
  NAND2X0 U12097 ( .IN1(n11696), .IN2(n11653), .QN(n11704) );
  INVX0 U12098 ( .INP(n3871), .ZN(n11653) );
  NAND2X0 U12099 ( .IN1(n5566), .IN2(g5527), .QN(n3871) );
  NAND3X0 U12100 ( .IN1(n11705), .IN2(n11706), .IN3(n11707), .QN(g30485) );
  NAND2X0 U12101 ( .IN1(n3886), .IN2(n11674), .QN(n11707) );
  NAND2X0 U12102 ( .IN1(n8639), .IN2(g5543), .QN(n11706) );
  NAND3X0 U12103 ( .IN1(n11708), .IN2(g5571), .IN3(n8487), .QN(n11705) );
  NAND2X0 U12104 ( .IN1(n11696), .IN2(n11674), .QN(n11708) );
  INVX0 U12105 ( .INP(n3874), .ZN(n11674) );
  NAND2X0 U12106 ( .IN1(n5566), .IN2(n5389), .QN(n3874) );
  INVX0 U12107 ( .INP(n3437), .ZN(n11696) );
  NAND2X0 U12108 ( .IN1(n8145), .IN2(g5511), .QN(n3437) );
  NAND3X0 U12109 ( .IN1(n11709), .IN2(n11710), .IN3(n11711), .QN(g30484) );
  NAND2X0 U12110 ( .IN1(n8639), .IN2(g5567), .QN(n11711) );
  OR3X1 U12111 ( .IN1(n8532), .IN2(n8016), .IN3(n3891), .Q(n11710) );
  NAND2X0 U12112 ( .IN1(n3891), .IN2(n3765), .QN(n11709) );
  NAND3X0 U12113 ( .IN1(n11712), .IN2(n11713), .IN3(n11714), .QN(g30483) );
  NAND2X0 U12114 ( .IN1(test_so6), .IN2(n8555), .QN(n11714) );
  OR3X1 U12115 ( .IN1(n8532), .IN2(n8105), .IN3(n3894), .Q(n11713) );
  NAND2X0 U12116 ( .IN1(n3894), .IN2(n3765), .QN(n11712) );
  NAND3X0 U12117 ( .IN1(n11715), .IN2(n11716), .IN3(n11717), .QN(g30482) );
  NAND2X0 U12118 ( .IN1(n8639), .IN2(g5551), .QN(n11717) );
  OR3X1 U12119 ( .IN1(n8531), .IN2(n7884), .IN3(n3896), .Q(n11716) );
  NAND2X0 U12120 ( .IN1(n3896), .IN2(n3765), .QN(n11715) );
  NAND3X0 U12121 ( .IN1(n11718), .IN2(n11719), .IN3(n11720), .QN(g30481) );
  NAND2X0 U12122 ( .IN1(n8639), .IN2(g5535), .QN(n11720) );
  OR3X1 U12123 ( .IN1(n8530), .IN2(n8046), .IN3(n3898), .Q(n11719) );
  NAND2X0 U12124 ( .IN1(n3898), .IN2(n3765), .QN(n11718) );
  NOR2X0 U12125 ( .IN1(g5511), .IN2(n10928), .QN(g30480) );
  NAND3X0 U12126 ( .IN1(n10919), .IN2(n8484), .IN3(n5647), .QN(n10928) );
  NAND2X0 U12127 ( .IN1(n3833), .IN2(n10340), .QN(n10919) );
  NAND3X0 U12128 ( .IN1(n11721), .IN2(n11722), .IN3(n11723), .QN(g30479) );
  NAND2X0 U12129 ( .IN1(n8639), .IN2(g5268), .QN(n11723) );
  NAND2X0 U12130 ( .IN1(n11724), .IN2(g5272), .QN(n11722) );
  NAND2X0 U12131 ( .IN1(n3765), .IN2(g26801), .QN(n11721) );
  NAND3X0 U12132 ( .IN1(n11725), .IN2(n11726), .IN3(n11727), .QN(g30478) );
  NAND2X0 U12133 ( .IN1(n11728), .IN2(n3765), .QN(n11727) );
  OR3X1 U12134 ( .IN1(n11728), .IN2(n8003), .IN3(n8543), .Q(n11726) );
  NOR2X0 U12135 ( .IN1(n3902), .IN2(n5650), .QN(n11728) );
  NAND2X0 U12136 ( .IN1(n8638), .IN2(g5264), .QN(n11725) );
  NAND3X0 U12137 ( .IN1(n11729), .IN2(n11730), .IN3(n11731), .QN(g30477) );
  NAND2X0 U12138 ( .IN1(n11732), .IN2(n3765), .QN(n11731) );
  INVX0 U12139 ( .INP(n10942), .ZN(n11732) );
  NAND3X0 U12140 ( .IN1(n10942), .IN2(g5212), .IN3(n8487), .QN(n11730) );
  NAND2X0 U12141 ( .IN1(n11733), .IN2(g5176), .QN(n10942) );
  NAND2X0 U12142 ( .IN1(n8638), .IN2(g5260), .QN(n11729) );
  NAND3X0 U12143 ( .IN1(n11734), .IN2(n11735), .IN3(n11736), .QN(g30476) );
  NAND2X0 U12144 ( .IN1(n11737), .IN2(n3765), .QN(n11736) );
  OR3X1 U12145 ( .IN1(n11737), .IN2(n8040), .IN3(n8541), .Q(n11735) );
  NOR2X0 U12146 ( .IN1(n3907), .IN2(n5650), .QN(n11737) );
  NAND2X0 U12147 ( .IN1(n8638), .IN2(g5256), .QN(n11734) );
  NAND3X0 U12148 ( .IN1(n11738), .IN2(n11739), .IN3(n11740), .QN(g30475) );
  NAND2X0 U12149 ( .IN1(n3908), .IN2(n11741), .QN(n11740) );
  NAND2X0 U12150 ( .IN1(n8638), .IN2(g5252), .QN(n11739) );
  NAND3X0 U12151 ( .IN1(n11742), .IN2(g5268), .IN3(n8487), .QN(n11738) );
  NAND2X0 U12152 ( .IN1(n10952), .IN2(n11741), .QN(n11742) );
  NAND3X0 U12153 ( .IN1(n11743), .IN2(n11744), .IN3(n11745), .QN(g30474) );
  NAND2X0 U12154 ( .IN1(n3908), .IN2(n10944), .QN(n11745) );
  NAND2X0 U12155 ( .IN1(n8638), .IN2(g5248), .QN(n11744) );
  NAND3X0 U12156 ( .IN1(n11746), .IN2(g5264), .IN3(n8487), .QN(n11743) );
  NAND2X0 U12157 ( .IN1(n10952), .IN2(n10944), .QN(n11746) );
  NAND3X0 U12158 ( .IN1(n11747), .IN2(n11748), .IN3(n11749), .QN(g30473) );
  NAND2X0 U12159 ( .IN1(n3908), .IN2(n11733), .QN(n11749) );
  NAND2X0 U12160 ( .IN1(n8638), .IN2(g5244), .QN(n11748) );
  NAND3X0 U12161 ( .IN1(n11750), .IN2(g5260), .IN3(n8486), .QN(n11747) );
  NAND2X0 U12162 ( .IN1(n10952), .IN2(n11733), .QN(n11750) );
  NAND3X0 U12163 ( .IN1(n11751), .IN2(n11752), .IN3(n11753), .QN(g30472) );
  NAND2X0 U12164 ( .IN1(n3908), .IN2(n11754), .QN(n11753) );
  NAND2X0 U12165 ( .IN1(n8638), .IN2(g5240), .QN(n11752) );
  NAND3X0 U12166 ( .IN1(n11755), .IN2(g5256), .IN3(n8487), .QN(n11751) );
  NAND2X0 U12167 ( .IN1(n10952), .IN2(n11754), .QN(n11755) );
  INVX0 U12168 ( .INP(n3444), .ZN(n10952) );
  NAND2X0 U12169 ( .IN1(g5170), .IN2(g5164), .QN(n3444) );
  NAND3X0 U12170 ( .IN1(n11756), .IN2(n11757), .IN3(n11758), .QN(g30471) );
  NAND2X0 U12171 ( .IN1(n3914), .IN2(n11741), .QN(n11758) );
  NAND2X0 U12172 ( .IN1(n8637), .IN2(g5236), .QN(n11757) );
  NAND3X0 U12173 ( .IN1(n11759), .IN2(g5252), .IN3(n8486), .QN(n11756) );
  NAND2X0 U12174 ( .IN1(n10957), .IN2(n11741), .QN(n11759) );
  NAND3X0 U12175 ( .IN1(n11760), .IN2(n11761), .IN3(n11762), .QN(g30470) );
  NAND2X0 U12176 ( .IN1(n3914), .IN2(n10944), .QN(n11762) );
  NAND2X0 U12177 ( .IN1(n8637), .IN2(g5232), .QN(n11761) );
  NAND3X0 U12178 ( .IN1(n11763), .IN2(g5248), .IN3(n8486), .QN(n11760) );
  NAND2X0 U12179 ( .IN1(n10957), .IN2(n10944), .QN(n11763) );
  NAND3X0 U12180 ( .IN1(n11764), .IN2(n11765), .IN3(n11766), .QN(g30469) );
  NAND2X0 U12181 ( .IN1(n3914), .IN2(n11733), .QN(n11766) );
  NAND2X0 U12182 ( .IN1(test_so82), .IN2(n8551), .QN(n11765) );
  NAND3X0 U12183 ( .IN1(n11767), .IN2(g5244), .IN3(n8486), .QN(n11764) );
  NAND2X0 U12184 ( .IN1(n10957), .IN2(n11733), .QN(n11767) );
  NAND3X0 U12185 ( .IN1(n11768), .IN2(n11769), .IN3(n11770), .QN(g30468) );
  NAND2X0 U12186 ( .IN1(n3914), .IN2(n11754), .QN(n11770) );
  NAND2X0 U12187 ( .IN1(n8637), .IN2(g5224), .QN(n11769) );
  NAND3X0 U12188 ( .IN1(n11771), .IN2(g5240), .IN3(n8486), .QN(n11768) );
  NAND2X0 U12189 ( .IN1(n10957), .IN2(n11754), .QN(n11771) );
  INVX0 U12190 ( .INP(n3446), .ZN(n10957) );
  NAND2X0 U12191 ( .IN1(n5570), .IN2(g5170), .QN(n3446) );
  NAND3X0 U12192 ( .IN1(n11772), .IN2(n11773), .IN3(n11774), .QN(g30467) );
  NAND2X0 U12193 ( .IN1(n3919), .IN2(n11741), .QN(n11774) );
  NAND2X0 U12194 ( .IN1(n8637), .IN2(g5216), .QN(n11773) );
  NAND3X0 U12195 ( .IN1(n11775), .IN2(g5236), .IN3(n8485), .QN(n11772) );
  NAND2X0 U12196 ( .IN1(n11776), .IN2(n11741), .QN(n11775) );
  INVX0 U12197 ( .INP(n3910), .ZN(n11741) );
  NAND3X0 U12198 ( .IN1(n11777), .IN2(n11778), .IN3(n11779), .QN(g30466) );
  NAND2X0 U12199 ( .IN1(n3919), .IN2(n10944), .QN(n11779) );
  NAND2X0 U12200 ( .IN1(n8637), .IN2(g5208), .QN(n11778) );
  NAND3X0 U12201 ( .IN1(n11780), .IN2(g5232), .IN3(n8485), .QN(n11777) );
  NAND2X0 U12202 ( .IN1(n11776), .IN2(n10944), .QN(n11780) );
  INVX0 U12203 ( .INP(n3902), .ZN(n10944) );
  NAND2X0 U12204 ( .IN1(n5384), .IN2(g5188), .QN(n3902) );
  NAND3X0 U12205 ( .IN1(n11781), .IN2(n11782), .IN3(n11783), .QN(g30465) );
  NAND2X0 U12206 ( .IN1(n3919), .IN2(n11733), .QN(n11783) );
  NAND2X0 U12207 ( .IN1(n8637), .IN2(g5200), .QN(n11782) );
  NAND3X0 U12208 ( .IN1(test_so82), .IN2(n11784), .IN3(n8485), .QN(n11781) );
  NAND2X0 U12209 ( .IN1(n11776), .IN2(n11733), .QN(n11784) );
  INVX0 U12210 ( .INP(n3904), .ZN(n11733) );
  NAND2X0 U12211 ( .IN1(n5567), .IN2(g5180), .QN(n3904) );
  NAND3X0 U12212 ( .IN1(n11785), .IN2(n11786), .IN3(n11787), .QN(g30464) );
  NAND2X0 U12213 ( .IN1(n3919), .IN2(n11754), .QN(n11787) );
  NAND2X0 U12214 ( .IN1(n8637), .IN2(g5196), .QN(n11786) );
  NAND3X0 U12215 ( .IN1(n11788), .IN2(g5224), .IN3(n8485), .QN(n11785) );
  NAND2X0 U12216 ( .IN1(n11776), .IN2(n11754), .QN(n11788) );
  INVX0 U12217 ( .INP(n3907), .ZN(n11754) );
  NAND2X0 U12218 ( .IN1(n5567), .IN2(n5384), .QN(n3907) );
  INVX0 U12219 ( .INP(n3447), .ZN(n11776) );
  NAND2X0 U12220 ( .IN1(n8140), .IN2(g5164), .QN(n3447) );
  NAND3X0 U12221 ( .IN1(n11789), .IN2(n11790), .IN3(n11791), .QN(g30463) );
  NAND2X0 U12222 ( .IN1(n8636), .IN2(g5220), .QN(n11791) );
  OR3X1 U12223 ( .IN1(n8530), .IN2(n8010), .IN3(n3924), .Q(n11790) );
  NAND2X0 U12224 ( .IN1(n3924), .IN2(n3765), .QN(n11789) );
  NAND3X0 U12225 ( .IN1(n11792), .IN2(n11793), .IN3(n11794), .QN(g30462) );
  NAND2X0 U12226 ( .IN1(n8636), .IN2(g5212), .QN(n11794) );
  OR3X1 U12227 ( .IN1(n8529), .IN2(n8004), .IN3(n3927), .Q(n11793) );
  NAND2X0 U12228 ( .IN1(n3927), .IN2(n3765), .QN(n11792) );
  NAND3X0 U12229 ( .IN1(n11795), .IN2(n11796), .IN3(n11797), .QN(g30461) );
  NAND2X0 U12230 ( .IN1(n8636), .IN2(g5204), .QN(n11797) );
  OR3X1 U12231 ( .IN1(n8529), .IN2(n7899), .IN3(n3929), .Q(n11796) );
  NAND2X0 U12232 ( .IN1(n3929), .IN2(n3765), .QN(n11795) );
  NAND3X0 U12233 ( .IN1(n11798), .IN2(n11799), .IN3(n11800), .QN(g30460) );
  NAND2X0 U12234 ( .IN1(n8636), .IN2(g5188), .QN(n11800) );
  OR3X1 U12235 ( .IN1(n8529), .IN2(n8042), .IN3(n3931), .Q(n11799) );
  NAND2X0 U12236 ( .IN1(n3931), .IN2(n3765), .QN(n11798) );
  NOR2X0 U12237 ( .IN1(g5164), .IN2(n10949), .QN(g30459) );
  NAND3X0 U12238 ( .IN1(n10940), .IN2(n8482), .IN3(n5650), .QN(n10949) );
  NAND2X0 U12239 ( .IN1(n3833), .IN2(n9602), .QN(n10940) );
  NAND3X0 U12240 ( .IN1(n11801), .IN2(n11802), .IN3(n8484), .QN(g30458) );
  NAND2X0 U12241 ( .IN1(n11803), .IN2(g113), .QN(n11802) );
  OR2X1 U12242 ( .IN1(n11803), .IN2(n5846), .Q(n11801) );
  NOR2X0 U12243 ( .IN1(g4459), .IN2(n7794), .QN(n11803) );
  NAND2X0 U12244 ( .IN1(n11804), .IN2(n11805), .QN(g30457) );
  OR2X1 U12245 ( .IN1(n8478), .IN2(n7696), .Q(n11805) );
  NAND2X0 U12246 ( .IN1(n11806), .IN2(n8528), .QN(n11804) );
  NAND2X0 U12247 ( .IN1(n11807), .IN2(n11808), .QN(n11806) );
  NAND2X0 U12248 ( .IN1(n11809), .IN2(n5981), .QN(n11808) );
  XNOR2X1 U12249 ( .IN1(g126), .IN2(n11810), .Q(n11809) );
  NAND2X0 U12250 ( .IN1(n11811), .IN2(n5983), .QN(n11807) );
  XNOR2X1 U12251 ( .IN1(g115), .IN2(n11812), .Q(n11811) );
  NAND3X0 U12252 ( .IN1(n11813), .IN2(n11814), .IN3(n11815), .QN(g30456) );
  NAND2X0 U12253 ( .IN1(n8596), .IN2(g4087), .QN(n11815) );
  NAND3X0 U12254 ( .IN1(n10340), .IN2(g4169), .IN3(n11334), .QN(n11814) );
  NAND2X0 U12255 ( .IN1(n3941), .IN2(n11816), .QN(n11813) );
  NAND3X0 U12256 ( .IN1(n11817), .IN2(n11818), .IN3(n11819), .QN(g30455) );
  NAND2X0 U12257 ( .IN1(n8596), .IN2(g3961), .QN(n11819) );
  NAND2X0 U12258 ( .IN1(n11820), .IN2(g3965), .QN(n11818) );
  NAND2X0 U12259 ( .IN1(n11821), .IN2(n3765), .QN(n11817) );
  NAND3X0 U12260 ( .IN1(n11822), .IN2(n11823), .IN3(n11824), .QN(g30454) );
  NAND2X0 U12261 ( .IN1(n11825), .IN2(n3765), .QN(n11824) );
  OR3X1 U12262 ( .IN1(n11825), .IN2(n8107), .IN3(n8542), .Q(n11823) );
  NOR2X0 U12263 ( .IN1(n8209), .IN2(n3945), .QN(n11825) );
  NAND2X0 U12264 ( .IN1(n8595), .IN2(g3957), .QN(n11822) );
  NAND3X0 U12265 ( .IN1(n11826), .IN2(n11827), .IN3(n11828), .QN(g30453) );
  NAND2X0 U12266 ( .IN1(n11829), .IN2(n3765), .QN(n11828) );
  INVX0 U12267 ( .INP(n10993), .ZN(n11829) );
  NAND3X0 U12268 ( .IN1(n10993), .IN2(g3905), .IN3(n8486), .QN(n11827) );
  NAND2X0 U12269 ( .IN1(test_so33), .IN2(n11830), .QN(n10993) );
  NAND2X0 U12270 ( .IN1(n8595), .IN2(g3953), .QN(n11826) );
  NAND3X0 U12271 ( .IN1(n11831), .IN2(n11832), .IN3(n11833), .QN(g30452) );
  NAND2X0 U12272 ( .IN1(n11834), .IN2(n3765), .QN(n11833) );
  OR3X1 U12273 ( .IN1(n11834), .IN2(n8047), .IN3(n8543), .Q(n11832) );
  NOR2X0 U12274 ( .IN1(n8209), .IN2(n3950), .QN(n11834) );
  NAND2X0 U12275 ( .IN1(test_so65), .IN2(n8550), .QN(n11831) );
  NAND3X0 U12276 ( .IN1(n11835), .IN2(n11836), .IN3(n11837), .QN(g30451) );
  NAND2X0 U12277 ( .IN1(n3951), .IN2(n11838), .QN(n11837) );
  NAND2X0 U12278 ( .IN1(n8595), .IN2(g3945), .QN(n11836) );
  NAND3X0 U12279 ( .IN1(n11839), .IN2(g3961), .IN3(n8484), .QN(n11835) );
  NAND2X0 U12280 ( .IN1(n11003), .IN2(n11838), .QN(n11839) );
  NAND3X0 U12281 ( .IN1(n11840), .IN2(n11841), .IN3(n11842), .QN(g30450) );
  NAND2X0 U12282 ( .IN1(n3951), .IN2(n10995), .QN(n11842) );
  NAND2X0 U12283 ( .IN1(n8595), .IN2(g3941), .QN(n11841) );
  NAND3X0 U12284 ( .IN1(n11843), .IN2(g3957), .IN3(n8485), .QN(n11840) );
  NAND2X0 U12285 ( .IN1(n11003), .IN2(n10995), .QN(n11843) );
  NAND3X0 U12286 ( .IN1(n11844), .IN2(n11845), .IN3(n11846), .QN(g30449) );
  NAND2X0 U12287 ( .IN1(n3951), .IN2(n11830), .QN(n11846) );
  NAND2X0 U12288 ( .IN1(n8595), .IN2(g3937), .QN(n11845) );
  NAND3X0 U12289 ( .IN1(n11847), .IN2(g3953), .IN3(n8484), .QN(n11844) );
  NAND2X0 U12290 ( .IN1(n11003), .IN2(n11830), .QN(n11847) );
  NAND3X0 U12291 ( .IN1(n11848), .IN2(n11849), .IN3(n11850), .QN(g30448) );
  NAND2X0 U12292 ( .IN1(n3951), .IN2(n11851), .QN(n11850) );
  NAND2X0 U12293 ( .IN1(n8595), .IN2(g3933), .QN(n11849) );
  NAND3X0 U12294 ( .IN1(test_so65), .IN2(n11852), .IN3(n8485), .QN(n11848) );
  NAND2X0 U12295 ( .IN1(n11003), .IN2(n11851), .QN(n11852) );
  INVX0 U12296 ( .INP(n3479), .ZN(n11003) );
  NAND2X0 U12297 ( .IN1(g3863), .IN2(g3857), .QN(n3479) );
  NAND3X0 U12298 ( .IN1(n11853), .IN2(n11854), .IN3(n11855), .QN(g30447) );
  NAND2X0 U12299 ( .IN1(n3957), .IN2(n11838), .QN(n11855) );
  NAND2X0 U12300 ( .IN1(n8595), .IN2(g3929), .QN(n11854) );
  NAND3X0 U12301 ( .IN1(n11856), .IN2(g3945), .IN3(n8485), .QN(n11853) );
  NAND2X0 U12302 ( .IN1(n11008), .IN2(n11838), .QN(n11856) );
  NAND3X0 U12303 ( .IN1(n11857), .IN2(n11858), .IN3(n11859), .QN(g30446) );
  NAND2X0 U12304 ( .IN1(n3957), .IN2(n10995), .QN(n11859) );
  NAND2X0 U12305 ( .IN1(n8594), .IN2(g3925), .QN(n11858) );
  NAND3X0 U12306 ( .IN1(n11860), .IN2(g3941), .IN3(n8484), .QN(n11857) );
  NAND2X0 U12307 ( .IN1(n11008), .IN2(n10995), .QN(n11860) );
  NAND3X0 U12308 ( .IN1(n11861), .IN2(n11862), .IN3(n11863), .QN(g30445) );
  NAND2X0 U12309 ( .IN1(n3957), .IN2(n11830), .QN(n11863) );
  NAND2X0 U12310 ( .IN1(n8594), .IN2(g3921), .QN(n11862) );
  NAND3X0 U12311 ( .IN1(n11864), .IN2(g3937), .IN3(n8484), .QN(n11861) );
  NAND2X0 U12312 ( .IN1(n11008), .IN2(n11830), .QN(n11864) );
  NAND3X0 U12313 ( .IN1(n11865), .IN2(n11866), .IN3(n11867), .QN(g30444) );
  NAND2X0 U12314 ( .IN1(n3957), .IN2(n11851), .QN(n11867) );
  NAND2X0 U12315 ( .IN1(n8594), .IN2(g3917), .QN(n11866) );
  NAND3X0 U12316 ( .IN1(n11868), .IN2(g3933), .IN3(n8486), .QN(n11865) );
  NAND2X0 U12317 ( .IN1(n11008), .IN2(n11851), .QN(n11868) );
  INVX0 U12318 ( .INP(n3481), .ZN(n11008) );
  NAND2X0 U12319 ( .IN1(n5572), .IN2(g3863), .QN(n3481) );
  NAND3X0 U12320 ( .IN1(n11869), .IN2(n11870), .IN3(n11871), .QN(g30443) );
  NAND2X0 U12321 ( .IN1(n3962), .IN2(n11838), .QN(n11871) );
  NAND2X0 U12322 ( .IN1(n8594), .IN2(g3909), .QN(n11870) );
  NAND3X0 U12323 ( .IN1(n11872), .IN2(g3929), .IN3(n8485), .QN(n11869) );
  NAND2X0 U12324 ( .IN1(n11873), .IN2(n11838), .QN(n11872) );
  NAND3X0 U12325 ( .IN1(n11874), .IN2(n11875), .IN3(n11876), .QN(g30442) );
  NAND2X0 U12326 ( .IN1(n3962), .IN2(n10995), .QN(n11876) );
  NAND2X0 U12327 ( .IN1(n8594), .IN2(g3901), .QN(n11875) );
  NAND3X0 U12328 ( .IN1(n11877), .IN2(g3925), .IN3(n8486), .QN(n11874) );
  NAND2X0 U12329 ( .IN1(n11873), .IN2(n10995), .QN(n11877) );
  INVX0 U12330 ( .INP(n3945), .ZN(n10995) );
  NAND2X0 U12331 ( .IN1(n5387), .IN2(g3881), .QN(n3945) );
  NAND3X0 U12332 ( .IN1(n11878), .IN2(n11879), .IN3(n11880), .QN(g30441) );
  NAND2X0 U12333 ( .IN1(n3962), .IN2(n11830), .QN(n11880) );
  NAND2X0 U12334 ( .IN1(n8594), .IN2(g3893), .QN(n11879) );
  NAND3X0 U12335 ( .IN1(n11881), .IN2(g3921), .IN3(n8485), .QN(n11878) );
  NAND2X0 U12336 ( .IN1(n11873), .IN2(n11830), .QN(n11881) );
  INVX0 U12337 ( .INP(n3947), .ZN(n11830) );
  NAND2X0 U12338 ( .IN1(n5564), .IN2(g3873), .QN(n3947) );
  NAND3X0 U12339 ( .IN1(n11882), .IN2(n11883), .IN3(n11884), .QN(g30440) );
  NAND2X0 U12340 ( .IN1(n3962), .IN2(n11851), .QN(n11884) );
  NAND2X0 U12341 ( .IN1(test_so24), .IN2(n8554), .QN(n11883) );
  NAND3X0 U12342 ( .IN1(n11885), .IN2(g3917), .IN3(n8485), .QN(n11882) );
  NAND2X0 U12343 ( .IN1(n11873), .IN2(n11851), .QN(n11885) );
  INVX0 U12344 ( .INP(n3950), .ZN(n11851) );
  NAND2X0 U12345 ( .IN1(n5564), .IN2(n5387), .QN(n3950) );
  INVX0 U12346 ( .INP(n3482), .ZN(n11873) );
  NAND2X0 U12347 ( .IN1(n8142), .IN2(g3857), .QN(n3482) );
  NAND3X0 U12348 ( .IN1(n11886), .IN2(n11887), .IN3(n11888), .QN(g30439) );
  NAND2X0 U12349 ( .IN1(n8594), .IN2(g3913), .QN(n11888) );
  OR3X1 U12350 ( .IN1(n8531), .IN2(n8019), .IN3(n3967), .Q(n11887) );
  NAND2X0 U12351 ( .IN1(n3967), .IN2(n3765), .QN(n11886) );
  NAND3X0 U12352 ( .IN1(n11889), .IN2(n11890), .IN3(n11891), .QN(g30438) );
  NAND2X0 U12353 ( .IN1(n8593), .IN2(g3905), .QN(n11891) );
  OR3X1 U12354 ( .IN1(n8531), .IN2(n8109), .IN3(n3970), .Q(n11890) );
  NAND2X0 U12355 ( .IN1(n3970), .IN2(n3765), .QN(n11889) );
  NAND3X0 U12356 ( .IN1(n11892), .IN2(n11893), .IN3(n11894), .QN(g30437) );
  NAND2X0 U12357 ( .IN1(n8593), .IN2(g3897), .QN(n11894) );
  OR3X1 U12358 ( .IN1(n8532), .IN2(n7904), .IN3(n3972), .Q(n11893) );
  NAND2X0 U12359 ( .IN1(n3972), .IN2(n3765), .QN(n11892) );
  NAND3X0 U12360 ( .IN1(n11895), .IN2(n11896), .IN3(n11897), .QN(g30436) );
  NAND2X0 U12361 ( .IN1(n8593), .IN2(g3881), .QN(n11897) );
  NAND3X0 U12362 ( .IN1(test_so24), .IN2(n8483), .IN3(n11898), .QN(n11896) );
  INVX0 U12363 ( .INP(n3974), .ZN(n11898) );
  NAND2X0 U12364 ( .IN1(n3974), .IN2(n3765), .QN(n11895) );
  NOR2X0 U12365 ( .IN1(g3857), .IN2(n11000), .QN(g30435) );
  NAND3X0 U12366 ( .IN1(n8503), .IN2(n8209), .IN3(n10991), .QN(n11000) );
  NAND3X0 U12367 ( .IN1(g4093), .IN2(g4087), .IN3(n3799), .QN(n10991) );
  NAND3X0 U12368 ( .IN1(n11899), .IN2(n11900), .IN3(n11901), .QN(g30434) );
  NAND2X0 U12369 ( .IN1(n8593), .IN2(g3610), .QN(n11901) );
  NAND2X0 U12370 ( .IN1(n11902), .IN2(g3614), .QN(n11900) );
  NAND2X0 U12371 ( .IN1(n11903), .IN2(n3765), .QN(n11899) );
  NAND3X0 U12372 ( .IN1(n11904), .IN2(n11905), .IN3(n11906), .QN(g30433) );
  NAND2X0 U12373 ( .IN1(n11907), .IN2(n3765), .QN(n11906) );
  OR3X1 U12374 ( .IN1(n11907), .IN2(n8115), .IN3(n8542), .Q(n11905) );
  NOR2X0 U12375 ( .IN1(n3978), .IN2(n5645), .QN(n11907) );
  NAND2X0 U12376 ( .IN1(n8593), .IN2(g3606), .QN(n11904) );
  NAND3X0 U12377 ( .IN1(n11908), .IN2(n11909), .IN3(n11910), .QN(g30432) );
  NAND2X0 U12378 ( .IN1(n11911), .IN2(n3765), .QN(n11910) );
  INVX0 U12379 ( .INP(n11014), .ZN(n11911) );
  NAND3X0 U12380 ( .IN1(n11014), .IN2(g3554), .IN3(n8485), .QN(n11909) );
  NAND2X0 U12381 ( .IN1(n11912), .IN2(g3518), .QN(n11014) );
  NAND2X0 U12382 ( .IN1(test_so43), .IN2(n8563), .QN(n11908) );
  NAND3X0 U12383 ( .IN1(n11913), .IN2(n11914), .IN3(n11915), .QN(g30431) );
  NAND2X0 U12384 ( .IN1(n11916), .IN2(n3765), .QN(n11915) );
  OR3X1 U12385 ( .IN1(n11916), .IN2(n8050), .IN3(n8541), .Q(n11914) );
  NOR2X0 U12386 ( .IN1(n3983), .IN2(n5645), .QN(n11916) );
  NAND2X0 U12387 ( .IN1(n8593), .IN2(g3598), .QN(n11913) );
  NAND3X0 U12388 ( .IN1(n11917), .IN2(n11918), .IN3(n11919), .QN(g30430) );
  NAND2X0 U12389 ( .IN1(n3984), .IN2(n11920), .QN(n11919) );
  NAND2X0 U12390 ( .IN1(n8593), .IN2(g3594), .QN(n11918) );
  NAND3X0 U12391 ( .IN1(n11921), .IN2(g3610), .IN3(n8487), .QN(n11917) );
  NAND2X0 U12392 ( .IN1(n11024), .IN2(n11920), .QN(n11921) );
  NAND3X0 U12393 ( .IN1(n11922), .IN2(n11923), .IN3(n11924), .QN(g30429) );
  NAND2X0 U12394 ( .IN1(n3984), .IN2(n11016), .QN(n11924) );
  NAND2X0 U12395 ( .IN1(n8592), .IN2(g3590), .QN(n11923) );
  NAND3X0 U12396 ( .IN1(n11925), .IN2(g3606), .IN3(n8487), .QN(n11922) );
  NAND2X0 U12397 ( .IN1(n11024), .IN2(n11016), .QN(n11925) );
  NAND3X0 U12398 ( .IN1(n11926), .IN2(n11927), .IN3(n11928), .QN(g30428) );
  NAND2X0 U12399 ( .IN1(n3984), .IN2(n11912), .QN(n11928) );
  NAND2X0 U12400 ( .IN1(n8592), .IN2(g3586), .QN(n11927) );
  NAND3X0 U12401 ( .IN1(test_so43), .IN2(n11929), .IN3(n8487), .QN(n11926) );
  NAND2X0 U12402 ( .IN1(n11024), .IN2(n11912), .QN(n11929) );
  NAND3X0 U12403 ( .IN1(n11930), .IN2(n11931), .IN3(n11932), .QN(g30427) );
  NAND2X0 U12404 ( .IN1(n3984), .IN2(n11933), .QN(n11932) );
  NAND2X0 U12405 ( .IN1(n8592), .IN2(g3582), .QN(n11931) );
  NAND3X0 U12406 ( .IN1(n11934), .IN2(g3598), .IN3(n8502), .QN(n11930) );
  NAND2X0 U12407 ( .IN1(n11024), .IN2(n11933), .QN(n11934) );
  INVX0 U12408 ( .INP(n3489), .ZN(n11024) );
  NAND2X0 U12409 ( .IN1(g3512), .IN2(g3506), .QN(n3489) );
  NAND3X0 U12410 ( .IN1(n11935), .IN2(n11936), .IN3(n11937), .QN(g30426) );
  NAND2X0 U12411 ( .IN1(n3990), .IN2(n11920), .QN(n11937) );
  NAND2X0 U12412 ( .IN1(n8592), .IN2(g3578), .QN(n11936) );
  NAND3X0 U12413 ( .IN1(n11938), .IN2(g3594), .IN3(n8502), .QN(n11935) );
  NAND2X0 U12414 ( .IN1(n11029), .IN2(n11920), .QN(n11938) );
  NAND3X0 U12415 ( .IN1(n11939), .IN2(n11940), .IN3(n11941), .QN(g30425) );
  NAND2X0 U12416 ( .IN1(n3990), .IN2(n11016), .QN(n11941) );
  NAND2X0 U12417 ( .IN1(n8592), .IN2(g3574), .QN(n11940) );
  NAND3X0 U12418 ( .IN1(n11942), .IN2(g3590), .IN3(n8502), .QN(n11939) );
  NAND2X0 U12419 ( .IN1(n11029), .IN2(n11016), .QN(n11942) );
  NAND3X0 U12420 ( .IN1(n11943), .IN2(n11944), .IN3(n11945), .QN(g30424) );
  NAND2X0 U12421 ( .IN1(n3990), .IN2(n11912), .QN(n11945) );
  NAND2X0 U12422 ( .IN1(n8592), .IN2(g3570), .QN(n11944) );
  NAND3X0 U12423 ( .IN1(n11946), .IN2(g3586), .IN3(n8502), .QN(n11943) );
  NAND2X0 U12424 ( .IN1(n11029), .IN2(n11912), .QN(n11946) );
  NAND3X0 U12425 ( .IN1(n11947), .IN2(n11948), .IN3(n11949), .QN(g30423) );
  NAND2X0 U12426 ( .IN1(n3990), .IN2(n11933), .QN(n11949) );
  NAND2X0 U12427 ( .IN1(n8592), .IN2(g3566), .QN(n11948) );
  NAND3X0 U12428 ( .IN1(n11950), .IN2(g3582), .IN3(n8502), .QN(n11947) );
  NAND2X0 U12429 ( .IN1(n11029), .IN2(n11933), .QN(n11950) );
  INVX0 U12430 ( .INP(n3491), .ZN(n11029) );
  NAND2X0 U12431 ( .IN1(n5576), .IN2(g3512), .QN(n3491) );
  NAND3X0 U12432 ( .IN1(n11951), .IN2(n11952), .IN3(n11953), .QN(g30422) );
  NAND2X0 U12433 ( .IN1(n3995), .IN2(n11920), .QN(n11953) );
  NAND2X0 U12434 ( .IN1(n8591), .IN2(g3558), .QN(n11952) );
  NAND3X0 U12435 ( .IN1(n11954), .IN2(g3578), .IN3(n8501), .QN(n11951) );
  NAND2X0 U12436 ( .IN1(n11955), .IN2(n11920), .QN(n11954) );
  NAND3X0 U12437 ( .IN1(n11956), .IN2(n11957), .IN3(n11958), .QN(g30421) );
  NAND2X0 U12438 ( .IN1(n3995), .IN2(n11016), .QN(n11958) );
  NAND2X0 U12439 ( .IN1(n8591), .IN2(g3550), .QN(n11957) );
  NAND3X0 U12440 ( .IN1(n11959), .IN2(g3574), .IN3(n8502), .QN(n11956) );
  NAND2X0 U12441 ( .IN1(n11955), .IN2(n11016), .QN(n11959) );
  INVX0 U12442 ( .INP(n3978), .ZN(n11016) );
  NAND2X0 U12443 ( .IN1(n5383), .IN2(g3530), .QN(n3978) );
  NAND3X0 U12444 ( .IN1(n11960), .IN2(n11961), .IN3(n11962), .QN(g30420) );
  NAND2X0 U12445 ( .IN1(n3995), .IN2(n11912), .QN(n11962) );
  NAND2X0 U12446 ( .IN1(n8591), .IN2(g3542), .QN(n11961) );
  NAND3X0 U12447 ( .IN1(n11963), .IN2(g3570), .IN3(n8501), .QN(n11960) );
  NAND2X0 U12448 ( .IN1(n11955), .IN2(n11912), .QN(n11963) );
  INVX0 U12449 ( .INP(n3980), .ZN(n11912) );
  NAND2X0 U12450 ( .IN1(n5569), .IN2(g3522), .QN(n3980) );
  NAND3X0 U12451 ( .IN1(n11964), .IN2(n11965), .IN3(n11966), .QN(g30419) );
  NAND2X0 U12452 ( .IN1(n3995), .IN2(n11933), .QN(n11966) );
  NAND2X0 U12453 ( .IN1(n8591), .IN2(g3538), .QN(n11965) );
  NAND3X0 U12454 ( .IN1(n11967), .IN2(g3566), .IN3(n8501), .QN(n11964) );
  NAND2X0 U12455 ( .IN1(n11955), .IN2(n11933), .QN(n11967) );
  INVX0 U12456 ( .INP(n3983), .ZN(n11933) );
  NAND2X0 U12457 ( .IN1(n5569), .IN2(n5383), .QN(n3983) );
  INVX0 U12458 ( .INP(n3492), .ZN(n11955) );
  NAND2X0 U12459 ( .IN1(n8146), .IN2(g3506), .QN(n3492) );
  NAND3X0 U12460 ( .IN1(n11968), .IN2(n11969), .IN3(n11970), .QN(g30418) );
  NAND2X0 U12461 ( .IN1(n8591), .IN2(g3562), .QN(n11970) );
  OR3X1 U12462 ( .IN1(n8534), .IN2(n8025), .IN3(n4000), .Q(n11969) );
  NAND2X0 U12463 ( .IN1(n4000), .IN2(n3765), .QN(n11968) );
  NAND3X0 U12464 ( .IN1(n11971), .IN2(n11972), .IN3(n11973), .QN(g30417) );
  NAND2X0 U12465 ( .IN1(n8591), .IN2(g3554), .QN(n11973) );
  OR3X1 U12466 ( .IN1(n8529), .IN2(n8117), .IN3(n4003), .Q(n11972) );
  NAND2X0 U12467 ( .IN1(n4003), .IN2(n3765), .QN(n11971) );
  NAND3X0 U12468 ( .IN1(n11974), .IN2(n11975), .IN3(n11976), .QN(g30416) );
  NAND2X0 U12469 ( .IN1(n8591), .IN2(g3546), .QN(n11976) );
  OR3X1 U12470 ( .IN1(n8535), .IN2(n7891), .IN3(n4005), .Q(n11975) );
  NAND2X0 U12471 ( .IN1(n4005), .IN2(n3765), .QN(n11974) );
  NAND3X0 U12472 ( .IN1(n11977), .IN2(n11978), .IN3(n11979), .QN(g30415) );
  NAND2X0 U12473 ( .IN1(n8590), .IN2(g3530), .QN(n11979) );
  OR3X1 U12474 ( .IN1(n8533), .IN2(n8051), .IN3(n4007), .Q(n11978) );
  NAND2X0 U12475 ( .IN1(n4007), .IN2(n3765), .QN(n11977) );
  NOR2X0 U12476 ( .IN1(g3506), .IN2(n11021), .QN(g30414) );
  NAND3X0 U12477 ( .IN1(n11012), .IN2(n8481), .IN3(n5645), .QN(n11021) );
  NAND3X0 U12478 ( .IN1(n5480), .IN2(g4093), .IN3(n3799), .QN(n11012) );
  NAND3X0 U12479 ( .IN1(n11980), .IN2(n11981), .IN3(n11982), .QN(g30413) );
  NAND2X0 U12480 ( .IN1(test_so84), .IN2(n8660), .QN(n11982) );
  NAND2X0 U12481 ( .IN1(n11983), .IN2(g3263), .QN(n11981) );
  NAND2X0 U12482 ( .IN1(n3765), .IN2(n10349), .QN(n11980) );
  NAND3X0 U12483 ( .IN1(n11984), .IN2(n11985), .IN3(n11986), .QN(g30412) );
  NAND2X0 U12484 ( .IN1(n11987), .IN2(n3765), .QN(n11986) );
  OR3X1 U12485 ( .IN1(n11987), .IN2(n8095), .IN3(n8542), .Q(n11985) );
  NOR2X0 U12486 ( .IN1(n3495), .IN2(n5652), .QN(n11987) );
  NAND2X0 U12487 ( .IN1(n8590), .IN2(g3255), .QN(n11984) );
  NAND3X0 U12488 ( .IN1(n11988), .IN2(n11989), .IN3(n11990), .QN(g30411) );
  NAND2X0 U12489 ( .IN1(n11991), .IN2(n3765), .QN(n11990) );
  INVX0 U12490 ( .INP(n11036), .ZN(n11991) );
  NAND3X0 U12491 ( .IN1(n11036), .IN2(g3203), .IN3(n8501), .QN(n11989) );
  NAND2X0 U12492 ( .IN1(n11992), .IN2(g3167), .QN(n11036) );
  NAND2X0 U12493 ( .IN1(n8590), .IN2(g3251), .QN(n11988) );
  NAND3X0 U12494 ( .IN1(n11993), .IN2(n11994), .IN3(n11995), .QN(g30410) );
  NAND2X0 U12495 ( .IN1(n11996), .IN2(n3765), .QN(n11995) );
  INVX0 U12496 ( .INP(n11997), .ZN(n11996) );
  NAND3X0 U12497 ( .IN1(test_so88), .IN2(n11997), .IN3(n8501), .QN(n11994) );
  NAND2X0 U12498 ( .IN1(n11998), .IN2(g3167), .QN(n11997) );
  NAND2X0 U12499 ( .IN1(n8590), .IN2(g3247), .QN(n11993) );
  NAND3X0 U12500 ( .IN1(n11999), .IN2(n12000), .IN3(n12001), .QN(g30409) );
  NAND2X0 U12501 ( .IN1(n4015), .IN2(n12002), .QN(n12001) );
  NAND2X0 U12502 ( .IN1(n8590), .IN2(g3243), .QN(n12000) );
  NAND3X0 U12503 ( .IN1(test_so84), .IN2(n12003), .IN3(n8500), .QN(n11999) );
  NAND2X0 U12504 ( .IN1(n11043), .IN2(n12002), .QN(n12003) );
  NAND3X0 U12505 ( .IN1(n12004), .IN2(n12005), .IN3(n12006), .QN(g30408) );
  NAND2X0 U12506 ( .IN1(n4015), .IN2(n12007), .QN(n12006) );
  NAND2X0 U12507 ( .IN1(n8590), .IN2(g3239), .QN(n12005) );
  NAND3X0 U12508 ( .IN1(n12008), .IN2(g3255), .IN3(n8501), .QN(n12004) );
  NAND2X0 U12509 ( .IN1(n12007), .IN2(n11043), .QN(n12008) );
  NAND3X0 U12510 ( .IN1(n12009), .IN2(n12010), .IN3(n12011), .QN(g30407) );
  NAND2X0 U12511 ( .IN1(n4015), .IN2(n11992), .QN(n12011) );
  NAND2X0 U12512 ( .IN1(n8590), .IN2(g3235), .QN(n12010) );
  NAND3X0 U12513 ( .IN1(n12012), .IN2(g3251), .IN3(n8501), .QN(n12009) );
  NAND2X0 U12514 ( .IN1(n11043), .IN2(n11992), .QN(n12012) );
  NAND3X0 U12515 ( .IN1(n12013), .IN2(n12014), .IN3(n12015), .QN(g30406) );
  NAND2X0 U12516 ( .IN1(n4015), .IN2(n11998), .QN(n12015) );
  NAND2X0 U12517 ( .IN1(n8589), .IN2(g3231), .QN(n12014) );
  NAND3X0 U12518 ( .IN1(n12016), .IN2(g3247), .IN3(n8501), .QN(n12013) );
  NAND2X0 U12519 ( .IN1(n11043), .IN2(n11998), .QN(n12016) );
  INVX0 U12520 ( .INP(n3500), .ZN(n11043) );
  NAND2X0 U12521 ( .IN1(g3161), .IN2(g3155), .QN(n3500) );
  NAND3X0 U12522 ( .IN1(n12017), .IN2(n12018), .IN3(n12019), .QN(g30405) );
  NAND2X0 U12523 ( .IN1(n4022), .IN2(n12002), .QN(n12019) );
  NAND2X0 U12524 ( .IN1(n8589), .IN2(g3227), .QN(n12018) );
  NAND3X0 U12525 ( .IN1(n12020), .IN2(g3243), .IN3(n8501), .QN(n12017) );
  NAND2X0 U12526 ( .IN1(n11048), .IN2(n12002), .QN(n12020) );
  NAND3X0 U12527 ( .IN1(n12021), .IN2(n12022), .IN3(n12023), .QN(g30404) );
  NAND2X0 U12528 ( .IN1(n4022), .IN2(n12007), .QN(n12023) );
  NAND2X0 U12529 ( .IN1(n8589), .IN2(g3223), .QN(n12022) );
  NAND3X0 U12530 ( .IN1(n12024), .IN2(g3239), .IN3(n8501), .QN(n12021) );
  NAND2X0 U12531 ( .IN1(n12007), .IN2(n11048), .QN(n12024) );
  NAND3X0 U12532 ( .IN1(n12025), .IN2(n12026), .IN3(n12027), .QN(g30403) );
  NAND2X0 U12533 ( .IN1(n4022), .IN2(n11992), .QN(n12027) );
  NAND2X0 U12534 ( .IN1(n8589), .IN2(g3219), .QN(n12026) );
  NAND3X0 U12535 ( .IN1(n12028), .IN2(g3235), .IN3(n8500), .QN(n12025) );
  NAND2X0 U12536 ( .IN1(n11048), .IN2(n11992), .QN(n12028) );
  NAND3X0 U12537 ( .IN1(n12029), .IN2(n12030), .IN3(n12031), .QN(g30402) );
  NAND2X0 U12538 ( .IN1(n4022), .IN2(n11998), .QN(n12031) );
  NAND2X0 U12539 ( .IN1(n8589), .IN2(g3215), .QN(n12030) );
  NAND3X0 U12540 ( .IN1(n12032), .IN2(g3231), .IN3(n8500), .QN(n12029) );
  NAND2X0 U12541 ( .IN1(n11048), .IN2(n11998), .QN(n12032) );
  INVX0 U12542 ( .INP(n3502), .ZN(n11048) );
  NAND2X0 U12543 ( .IN1(n5366), .IN2(g3161), .QN(n3502) );
  NAND3X0 U12544 ( .IN1(n12033), .IN2(n12034), .IN3(n12035), .QN(g30401) );
  NAND2X0 U12545 ( .IN1(n4027), .IN2(n12002), .QN(n12035) );
  NAND2X0 U12546 ( .IN1(n8589), .IN2(g3207), .QN(n12034) );
  NAND3X0 U12547 ( .IN1(n12036), .IN2(g3227), .IN3(n8499), .QN(n12033) );
  NAND2X0 U12548 ( .IN1(n12037), .IN2(n12002), .QN(n12036) );
  INVX0 U12549 ( .INP(n4017), .ZN(n12002) );
  NAND3X0 U12550 ( .IN1(n12038), .IN2(n12039), .IN3(n12040), .QN(g30400) );
  NAND2X0 U12551 ( .IN1(n4027), .IN2(n12007), .QN(n12040) );
  NAND2X0 U12552 ( .IN1(n8589), .IN2(g3199), .QN(n12039) );
  NAND3X0 U12553 ( .IN1(n12041), .IN2(g3223), .IN3(n8499), .QN(n12038) );
  NAND2X0 U12554 ( .IN1(n12007), .IN2(n12037), .QN(n12041) );
  INVX0 U12555 ( .INP(n3495), .ZN(n12007) );
  NAND2X0 U12556 ( .IN1(n5603), .IN2(g3179), .QN(n3495) );
  NAND3X0 U12557 ( .IN1(n12042), .IN2(n12043), .IN3(n12044), .QN(g30399) );
  NAND2X0 U12558 ( .IN1(n4027), .IN2(n11992), .QN(n12044) );
  NAND2X0 U12559 ( .IN1(n8588), .IN2(g3191), .QN(n12043) );
  NAND3X0 U12560 ( .IN1(n12045), .IN2(g3219), .IN3(n8499), .QN(n12042) );
  NAND2X0 U12561 ( .IN1(n12037), .IN2(n11992), .QN(n12045) );
  INVX0 U12562 ( .INP(n4020), .ZN(n11992) );
  NAND2X0 U12563 ( .IN1(n5390), .IN2(g3171), .QN(n4020) );
  NAND3X0 U12564 ( .IN1(n12046), .IN2(n12047), .IN3(n12048), .QN(g30398) );
  NAND2X0 U12565 ( .IN1(n4027), .IN2(n11998), .QN(n12048) );
  NAND2X0 U12566 ( .IN1(n8588), .IN2(g3187), .QN(n12047) );
  NAND3X0 U12567 ( .IN1(n12049), .IN2(g3215), .IN3(n8498), .QN(n12046) );
  NAND2X0 U12568 ( .IN1(n12037), .IN2(n11998), .QN(n12049) );
  INVX0 U12569 ( .INP(n4014), .ZN(n11998) );
  NAND2X0 U12570 ( .IN1(n5603), .IN2(n5390), .QN(n4014) );
  INVX0 U12571 ( .INP(n3501), .ZN(n12037) );
  NAND2X0 U12572 ( .IN1(n8150), .IN2(g3155), .QN(n3501) );
  NAND3X0 U12573 ( .IN1(n12050), .IN2(n12051), .IN3(n12052), .QN(g30397) );
  NAND2X0 U12574 ( .IN1(n8588), .IN2(g3211), .QN(n12052) );
  OR3X1 U12575 ( .IN1(n8536), .IN2(n8007), .IN3(n4032), .Q(n12051) );
  NAND2X0 U12576 ( .IN1(n4032), .IN2(n3765), .QN(n12050) );
  NAND3X0 U12577 ( .IN1(n12053), .IN2(n12054), .IN3(n12055), .QN(g30396) );
  NAND2X0 U12578 ( .IN1(n8588), .IN2(g3203), .QN(n12055) );
  OR3X1 U12579 ( .IN1(n8535), .IN2(n8097), .IN3(n4035), .Q(n12054) );
  NAND2X0 U12580 ( .IN1(n4035), .IN2(n3765), .QN(n12053) );
  NAND3X0 U12581 ( .IN1(n12056), .IN2(n12057), .IN3(n12058), .QN(g30395) );
  NAND2X0 U12582 ( .IN1(test_so88), .IN2(n8661), .QN(n12058) );
  OR3X1 U12583 ( .IN1(n8533), .IN2(n7880), .IN3(n4037), .Q(n12057) );
  NAND2X0 U12584 ( .IN1(n4037), .IN2(n3765), .QN(n12056) );
  NAND3X0 U12585 ( .IN1(n12059), .IN2(n12060), .IN3(n12061), .QN(g30394) );
  NAND2X0 U12586 ( .IN1(n8588), .IN2(g3179), .QN(n12061) );
  OR3X1 U12587 ( .IN1(n8536), .IN2(n8038), .IN3(n4039), .Q(n12060) );
  NAND2X0 U12588 ( .IN1(n4039), .IN2(n3765), .QN(n12059) );
  AND3X1 U12589 ( .IN1(n5366), .IN2(n8528), .IN3(n11033), .Q(g30393) );
  AND2X1 U12590 ( .IN1(n5652), .IN2(n11035), .Q(n11033) );
  NAND2X0 U12591 ( .IN1(n3799), .IN2(n10340), .QN(n11035) );
  NAND2X0 U12592 ( .IN1(n12062), .IN2(n12063), .QN(g30392) );
  NAND2X0 U12593 ( .IN1(n8588), .IN2(g2803), .QN(n12063) );
  NAND2X0 U12594 ( .IN1(n12064), .IN2(n12065), .QN(g30391) );
  NAND2X0 U12595 ( .IN1(n8588), .IN2(g2771), .QN(n12065) );
  NAND2X0 U12596 ( .IN1(n12062), .IN2(n12066), .QN(g30390) );
  NAND2X0 U12597 ( .IN1(g2834), .IN2(n8660), .QN(n12066) );
  NAND2X0 U12598 ( .IN1(n12067), .IN2(n8527), .QN(n12062) );
  NAND2X0 U12599 ( .IN1(n12068), .IN2(n12069), .QN(n12067) );
  NAND4X0 U12600 ( .IN1(n12070), .IN2(n12071), .IN3(n12072), .IN4(n12073), 
        .QN(n12069) );
  NOR2X0 U12601 ( .IN1(n12074), .IN2(n12075), .QN(n12072) );
  NOR2X0 U12602 ( .IN1(n4411), .IN2(g2370), .QN(n12075) );
  NOR2X0 U12603 ( .IN1(n12076), .IN2(g2504), .QN(n12074) );
  NAND2X0 U12604 ( .IN1(n7908), .IN2(n12077), .QN(n12071) );
  NAND2X0 U12605 ( .IN1(n7918), .IN2(n12078), .QN(n12070) );
  NAND4X0 U12606 ( .IN1(n12079), .IN2(n12080), .IN3(n12081), .IN4(n12082), 
        .QN(n12068) );
  NOR2X0 U12607 ( .IN1(n12083), .IN2(n12084), .QN(n12081) );
  NOR2X0 U12608 ( .IN1(n5609), .IN2(n12085), .QN(n12084) );
  NOR2X0 U12609 ( .IN1(n5545), .IN2(n12086), .QN(n12083) );
  NAND2X0 U12610 ( .IN1(n12087), .IN2(g2815), .QN(n12080) );
  NAND2X0 U12611 ( .IN1(n12088), .IN2(g2807), .QN(n12079) );
  NAND2X0 U12612 ( .IN1(n12064), .IN2(n12089), .QN(g30389) );
  NAND2X0 U12613 ( .IN1(g2831), .IN2(n8661), .QN(n12089) );
  NAND2X0 U12614 ( .IN1(n12090), .IN2(n8527), .QN(n12064) );
  NAND2X0 U12615 ( .IN1(n12091), .IN2(n12092), .QN(n12090) );
  NAND4X0 U12616 ( .IN1(n12093), .IN2(n12094), .IN3(n12095), .IN4(n12073), 
        .QN(n12092) );
  NOR2X0 U12617 ( .IN1(n12096), .IN2(n12097), .QN(n12095) );
  NOR2X0 U12618 ( .IN1(n4411), .IN2(g1811), .QN(n12097) );
  NOR2X0 U12619 ( .IN1(test_so53), .IN2(n12076), .QN(n12096) );
  NAND2X0 U12620 ( .IN1(n7914), .IN2(n12077), .QN(n12094) );
  NAND2X0 U12621 ( .IN1(n7915), .IN2(n12078), .QN(n12093) );
  NAND4X0 U12622 ( .IN1(n12098), .IN2(n12099), .IN3(n12100), .IN4(n12082), 
        .QN(n12091) );
  INVX0 U12623 ( .INP(n12073), .ZN(n12082) );
  NAND3X0 U12624 ( .IN1(n3653), .IN2(n9579), .IN3(n5600), .QN(n12073) );
  NOR2X0 U12625 ( .IN1(g2741), .IN2(n8896), .QN(n3653) );
  NOR2X0 U12626 ( .IN1(n12101), .IN2(n12102), .QN(n12100) );
  NOR2X0 U12627 ( .IN1(n5610), .IN2(n12085), .QN(n12102) );
  NOR2X0 U12628 ( .IN1(n5544), .IN2(n12086), .QN(n12101) );
  NAND2X0 U12629 ( .IN1(n12087), .IN2(g2783), .QN(n12099) );
  NAND2X0 U12630 ( .IN1(n12088), .IN2(g2775), .QN(n12098) );
  NAND2X0 U12631 ( .IN1(n12103), .IN2(n12104), .QN(g30388) );
  NAND2X0 U12632 ( .IN1(n12105), .IN2(n3730), .QN(n12104) );
  XOR2X1 U12633 ( .IN1(g2741), .IN2(n8897), .Q(n12105) );
  NOR2X0 U12634 ( .IN1(n12106), .IN2(n5600), .QN(n8897) );
  NAND2X0 U12635 ( .IN1(n8587), .IN2(g2735), .QN(n12103) );
  NAND3X0 U12636 ( .IN1(n12107), .IN2(n12108), .IN3(n12109), .QN(g30387) );
  OR2X1 U12637 ( .IN1(n12110), .IN2(n14517), .Q(n12109) );
  NAND2X0 U12638 ( .IN1(n12111), .IN2(g2681), .QN(n12108) );
  NAND2X0 U12639 ( .IN1(n12112), .IN2(n8527), .QN(n12111) );
  OR2X1 U12640 ( .IN1(n12113), .IN2(n5457), .Q(n12112) );
  NAND3X0 U12641 ( .IN1(n12114), .IN2(n5457), .IN3(n5777), .QN(n12107) );
  NAND2X0 U12642 ( .IN1(n12115), .IN2(n12116), .QN(g30386) );
  NAND2X0 U12643 ( .IN1(n12117), .IN2(g2681), .QN(n12116) );
  NAND2X0 U12644 ( .IN1(n12110), .IN2(g2675), .QN(n12115) );
  NAND3X0 U12645 ( .IN1(n12118), .IN2(n12119), .IN3(n12120), .QN(g30385) );
  NAND2X0 U12646 ( .IN1(n8587), .IN2(g2657), .QN(n12120) );
  NAND2X0 U12647 ( .IN1(n12117), .IN2(g2661), .QN(n12119) );
  INVX0 U12648 ( .INP(n12110), .ZN(n12117) );
  NAND2X0 U12649 ( .IN1(n12113), .IN2(n8527), .QN(n12110) );
  NAND2X0 U12650 ( .IN1(n12114), .IN2(n5418), .QN(n12118) );
  NAND3X0 U12651 ( .IN1(n12121), .IN2(n12122), .IN3(n12123), .QN(g30384) );
  NAND2X0 U12652 ( .IN1(n8587), .IN2(g2652), .QN(n12123) );
  NAND3X0 U12653 ( .IN1(n3517), .IN2(n12124), .IN3(n326), .QN(n12122) );
  XOR2X1 U12654 ( .IN1(n7919), .IN2(n7753), .Q(n12124) );
  NAND2X0 U12655 ( .IN1(n12125), .IN2(g2657), .QN(n12121) );
  NAND2X0 U12656 ( .IN1(n11060), .IN2(n12126), .QN(n12125) );
  NAND2X0 U12657 ( .IN1(n11072), .IN2(n8527), .QN(n12126) );
  NAND2X0 U12658 ( .IN1(n12127), .IN2(n12128), .QN(g30383) );
  NAND2X0 U12659 ( .IN1(test_so66), .IN2(n8565), .QN(n12128) );
  NAND2X0 U12660 ( .IN1(n12129), .IN2(n8527), .QN(n12127) );
  NAND2X0 U12661 ( .IN1(n12130), .IN2(n12131), .QN(n12129) );
  NAND2X0 U12662 ( .IN1(test_so34), .IN2(n12132), .QN(n12131) );
  NAND2X0 U12663 ( .IN1(n12133), .IN2(n12134), .QN(n12130) );
  NAND2X0 U12664 ( .IN1(n5351), .IN2(g2599), .QN(n12134) );
  INVX0 U12665 ( .INP(n12132), .ZN(n12133) );
  NAND3X0 U12666 ( .IN1(n12135), .IN2(g2610), .IN3(n5508), .QN(n12132) );
  NAND3X0 U12667 ( .IN1(n12136), .IN2(n12137), .IN3(n12138), .QN(g30382) );
  NAND2X0 U12668 ( .IN1(n12139), .IN2(n9295), .QN(n12138) );
  NAND2X0 U12669 ( .IN1(n12140), .IN2(g2547), .QN(n12137) );
  NAND2X0 U12670 ( .IN1(n12141), .IN2(n8527), .QN(n12140) );
  OR2X1 U12671 ( .IN1(n12142), .IN2(n5461), .Q(n12141) );
  NAND3X0 U12672 ( .IN1(n12143), .IN2(n5461), .IN3(n5782), .QN(n12136) );
  NAND2X0 U12673 ( .IN1(n12144), .IN2(n12145), .QN(g30381) );
  NAND2X0 U12674 ( .IN1(n12139), .IN2(g2547), .QN(n12145) );
  NAND2X0 U12675 ( .IN1(n12146), .IN2(g2541), .QN(n12144) );
  NAND3X0 U12676 ( .IN1(n12147), .IN2(n12148), .IN3(n12149), .QN(g30380) );
  NAND2X0 U12677 ( .IN1(n8587), .IN2(g2523), .QN(n12149) );
  NAND2X0 U12678 ( .IN1(n12139), .IN2(g2527), .QN(n12148) );
  INVX0 U12679 ( .INP(n12146), .ZN(n12139) );
  NAND2X0 U12680 ( .IN1(n12142), .IN2(n8527), .QN(n12146) );
  NAND2X0 U12681 ( .IN1(n12143), .IN2(n5420), .QN(n12147) );
  NAND3X0 U12682 ( .IN1(n12150), .IN2(n12151), .IN3(n12152), .QN(g30379) );
  NAND2X0 U12683 ( .IN1(n8586), .IN2(g2518), .QN(n12152) );
  NAND3X0 U12684 ( .IN1(n3536), .IN2(n12153), .IN3(n911), .QN(n12151) );
  XOR2X1 U12685 ( .IN1(n7917), .IN2(n7750), .Q(n12153) );
  NAND2X0 U12686 ( .IN1(n12154), .IN2(g2523), .QN(n12150) );
  NAND2X0 U12687 ( .IN1(n11081), .IN2(n12155), .QN(n12154) );
  NAND2X0 U12688 ( .IN1(n11093), .IN2(n8527), .QN(n12155) );
  NAND2X0 U12689 ( .IN1(n12156), .IN2(n12157), .QN(g30378) );
  NAND2X0 U12690 ( .IN1(n8586), .IN2(g2441), .QN(n12157) );
  NAND2X0 U12691 ( .IN1(n12158), .IN2(n8527), .QN(n12156) );
  NAND2X0 U12692 ( .IN1(n12159), .IN2(n12160), .QN(n12158) );
  NAND2X0 U12693 ( .IN1(n12161), .IN2(g2461), .QN(n12160) );
  NAND2X0 U12694 ( .IN1(n12162), .IN2(n12163), .QN(n12159) );
  NAND2X0 U12695 ( .IN1(g2465), .IN2(n8204), .QN(n12163) );
  INVX0 U12696 ( .INP(n12161), .ZN(n12162) );
  NAND3X0 U12697 ( .IN1(n12164), .IN2(g2476), .IN3(n5509), .QN(n12161) );
  NAND3X0 U12698 ( .IN1(n12165), .IN2(n12166), .IN3(n12167), .QN(g30377) );
  NAND2X0 U12699 ( .IN1(n12168), .IN2(n9324), .QN(n12167) );
  NAND2X0 U12700 ( .IN1(test_so89), .IN2(n12169), .QN(n12166) );
  NAND2X0 U12701 ( .IN1(n12170), .IN2(n8526), .QN(n12169) );
  OR2X1 U12702 ( .IN1(n12171), .IN2(n5459), .Q(n12170) );
  NAND3X0 U12703 ( .IN1(n12172), .IN2(n5459), .IN3(n8234), .QN(n12165) );
  NAND2X0 U12704 ( .IN1(n12173), .IN2(n12174), .QN(g30376) );
  NAND2X0 U12705 ( .IN1(test_so89), .IN2(n12168), .QN(n12174) );
  NAND2X0 U12706 ( .IN1(n12175), .IN2(g2407), .QN(n12173) );
  NAND3X0 U12707 ( .IN1(n12176), .IN2(n12177), .IN3(n12178), .QN(g30375) );
  NAND2X0 U12708 ( .IN1(n8586), .IN2(g2389), .QN(n12178) );
  NAND2X0 U12709 ( .IN1(n12168), .IN2(g2393), .QN(n12177) );
  INVX0 U12710 ( .INP(n12175), .ZN(n12168) );
  NAND2X0 U12711 ( .IN1(n12171), .IN2(n8527), .QN(n12175) );
  NAND2X0 U12712 ( .IN1(n12172), .IN2(n5421), .QN(n12176) );
  NAND3X0 U12713 ( .IN1(n12179), .IN2(n12180), .IN3(n12181), .QN(g30374) );
  NAND2X0 U12714 ( .IN1(n8640), .IN2(g2384), .QN(n12181) );
  NAND3X0 U12715 ( .IN1(n3555), .IN2(n12182), .IN3(n456), .QN(n12180) );
  XOR2X1 U12716 ( .IN1(n7911), .IN2(n7749), .Q(n12182) );
  NAND2X0 U12717 ( .IN1(n12183), .IN2(g2389), .QN(n12179) );
  NAND2X0 U12718 ( .IN1(n11102), .IN2(n12184), .QN(n12183) );
  NAND2X0 U12719 ( .IN1(n11114), .IN2(n8527), .QN(n12184) );
  NAND2X0 U12720 ( .IN1(n12185), .IN2(n12186), .QN(g30373) );
  NAND2X0 U12721 ( .IN1(n8636), .IN2(g2307), .QN(n12186) );
  NAND2X0 U12722 ( .IN1(n12187), .IN2(n8527), .QN(n12185) );
  NAND2X0 U12723 ( .IN1(n12188), .IN2(n12189), .QN(n12187) );
  NAND2X0 U12724 ( .IN1(n12190), .IN2(g2327), .QN(n12189) );
  NAND2X0 U12725 ( .IN1(n12191), .IN2(n12192), .QN(n12188) );
  NAND2X0 U12726 ( .IN1(n5353), .IN2(g2331), .QN(n12192) );
  INVX0 U12727 ( .INP(n12190), .ZN(n12191) );
  NAND3X0 U12728 ( .IN1(n12193), .IN2(test_so21), .IN3(n5511), .QN(n12190) );
  NAND3X0 U12729 ( .IN1(n12194), .IN2(n12195), .IN3(n12196), .QN(g30372) );
  OR2X1 U12730 ( .IN1(n12197), .IN2(n14522), .Q(n12196) );
  NAND2X0 U12731 ( .IN1(n12198), .IN2(g2279), .QN(n12195) );
  NAND2X0 U12732 ( .IN1(n12199), .IN2(n8527), .QN(n12198) );
  OR2X1 U12733 ( .IN1(n12200), .IN2(n5458), .Q(n12199) );
  NAND3X0 U12734 ( .IN1(n12201), .IN2(n5458), .IN3(n5778), .QN(n12194) );
  NAND2X0 U12735 ( .IN1(n12202), .IN2(n12203), .QN(g30371) );
  NAND2X0 U12736 ( .IN1(n12204), .IN2(g2279), .QN(n12203) );
  NAND2X0 U12737 ( .IN1(n12197), .IN2(g2273), .QN(n12202) );
  NAND3X0 U12738 ( .IN1(n12205), .IN2(n12206), .IN3(n12207), .QN(g30370) );
  NAND2X0 U12739 ( .IN1(n8642), .IN2(g2255), .QN(n12207) );
  NAND2X0 U12740 ( .IN1(n12204), .IN2(g2259), .QN(n12206) );
  INVX0 U12741 ( .INP(n12197), .ZN(n12204) );
  NAND2X0 U12742 ( .IN1(n12200), .IN2(n8526), .QN(n12197) );
  NAND2X0 U12743 ( .IN1(n12201), .IN2(n5419), .QN(n12205) );
  NAND3X0 U12744 ( .IN1(n12208), .IN2(n12209), .IN3(n12210), .QN(g30369) );
  NAND2X0 U12745 ( .IN1(n8586), .IN2(g2250), .QN(n12210) );
  NAND3X0 U12746 ( .IN1(n3574), .IN2(n12211), .IN3(n982), .QN(n12209) );
  XOR2X1 U12747 ( .IN1(n7907), .IN2(n7752), .Q(n12211) );
  NAND2X0 U12748 ( .IN1(n12212), .IN2(g2255), .QN(n12208) );
  NAND2X0 U12749 ( .IN1(n11123), .IN2(n12213), .QN(n12212) );
  NAND2X0 U12750 ( .IN1(n11135), .IN2(n8526), .QN(n12213) );
  NAND2X0 U12751 ( .IN1(n12214), .IN2(n12215), .QN(g30368) );
  NAND2X0 U12752 ( .IN1(n8637), .IN2(g2173), .QN(n12215) );
  NAND2X0 U12753 ( .IN1(n12216), .IN2(n8527), .QN(n12214) );
  NAND2X0 U12754 ( .IN1(n12217), .IN2(n12218), .QN(n12216) );
  NAND2X0 U12755 ( .IN1(n12219), .IN2(g2193), .QN(n12218) );
  NAND2X0 U12756 ( .IN1(n12220), .IN2(n12221), .QN(n12217) );
  NAND2X0 U12757 ( .IN1(n5356), .IN2(g2197), .QN(n12221) );
  INVX0 U12758 ( .INP(n12219), .ZN(n12220) );
  NAND3X0 U12759 ( .IN1(n12222), .IN2(g2208), .IN3(n5512), .QN(n12219) );
  NAND3X0 U12760 ( .IN1(n12223), .IN2(n12224), .IN3(n12225), .QN(g30367) );
  NAND2X0 U12761 ( .IN1(n12226), .IN2(g2126), .QN(n12225) );
  NAND2X0 U12762 ( .IN1(n12227), .IN2(g2122), .QN(n12224) );
  NAND2X0 U12763 ( .IN1(n12228), .IN2(n8526), .QN(n12227) );
  OR2X1 U12764 ( .IN1(n12229), .IN2(n5463), .Q(n12228) );
  NAND3X0 U12765 ( .IN1(n12230), .IN2(n5463), .IN3(n5784), .QN(n12223) );
  NAND2X0 U12766 ( .IN1(n12231), .IN2(n12232), .QN(g30366) );
  NAND2X0 U12767 ( .IN1(n12226), .IN2(g2122), .QN(n12232) );
  NAND2X0 U12768 ( .IN1(n12233), .IN2(g2116), .QN(n12231) );
  NAND3X0 U12769 ( .IN1(n12234), .IN2(n12235), .IN3(n12236), .QN(g30365) );
  NAND2X0 U12770 ( .IN1(n8586), .IN2(g2098), .QN(n12236) );
  NAND2X0 U12771 ( .IN1(n12226), .IN2(g2102), .QN(n12235) );
  INVX0 U12772 ( .INP(n12233), .ZN(n12226) );
  NAND2X0 U12773 ( .IN1(n12229), .IN2(n8527), .QN(n12233) );
  NAND2X0 U12774 ( .IN1(n12230), .IN2(n5666), .QN(n12234) );
  NAND3X0 U12775 ( .IN1(n12237), .IN2(n12238), .IN3(n12239), .QN(g30364) );
  NAND2X0 U12776 ( .IN1(test_so78), .IN2(n8564), .QN(n12239) );
  NAND3X0 U12777 ( .IN1(n1136), .IN2(n3593), .IN3(n12240), .QN(n12238) );
  XOR2X1 U12778 ( .IN1(g2089), .IN2(test_so78), .Q(n12240) );
  NAND2X0 U12779 ( .IN1(n12241), .IN2(g2098), .QN(n12237) );
  NAND2X0 U12780 ( .IN1(n11144), .IN2(n12242), .QN(n12241) );
  NAND2X0 U12781 ( .IN1(n11156), .IN2(n8526), .QN(n12242) );
  NAND2X0 U12782 ( .IN1(n12243), .IN2(n12244), .QN(g30363) );
  NAND2X0 U12783 ( .IN1(n8586), .IN2(g2016), .QN(n12244) );
  NAND2X0 U12784 ( .IN1(n12245), .IN2(n8526), .QN(n12243) );
  NAND2X0 U12785 ( .IN1(n12246), .IN2(n12247), .QN(n12245) );
  NAND2X0 U12786 ( .IN1(test_so59), .IN2(n12248), .QN(n12247) );
  NAND2X0 U12787 ( .IN1(n12249), .IN2(n12250), .QN(n12246) );
  NAND2X0 U12788 ( .IN1(n5355), .IN2(g2040), .QN(n12250) );
  INVX0 U12789 ( .INP(n12248), .ZN(n12249) );
  NAND3X0 U12790 ( .IN1(n12251), .IN2(g2051), .IN3(n5507), .QN(n12248) );
  NAND3X0 U12791 ( .IN1(n12252), .IN2(n12253), .IN3(n12254), .QN(g30362) );
  NAND2X0 U12792 ( .IN1(n12255), .IN2(g1992), .QN(n12254) );
  NAND2X0 U12793 ( .IN1(n12256), .IN2(g1988), .QN(n12253) );
  NAND2X0 U12794 ( .IN1(n12257), .IN2(n8526), .QN(n12256) );
  OR2X1 U12795 ( .IN1(n12258), .IN2(n5462), .Q(n12257) );
  NAND3X0 U12796 ( .IN1(n12259), .IN2(n5462), .IN3(n5783), .QN(n12252) );
  NAND2X0 U12797 ( .IN1(n12260), .IN2(n12261), .QN(g30361) );
  NAND2X0 U12798 ( .IN1(n12255), .IN2(g1988), .QN(n12261) );
  NAND2X0 U12799 ( .IN1(n12262), .IN2(g1982), .QN(n12260) );
  NAND3X0 U12800 ( .IN1(n12263), .IN2(n12264), .IN3(n12265), .QN(g30360) );
  NAND2X0 U12801 ( .IN1(n8649), .IN2(g1964), .QN(n12265) );
  NAND2X0 U12802 ( .IN1(n12255), .IN2(g1968), .QN(n12264) );
  INVX0 U12803 ( .INP(n12262), .ZN(n12255) );
  NAND2X0 U12804 ( .IN1(n12258), .IN2(n8526), .QN(n12262) );
  NAND2X0 U12805 ( .IN1(n12259), .IN2(n5664), .QN(n12263) );
  NAND3X0 U12806 ( .IN1(n12266), .IN2(n12267), .IN3(n12268), .QN(g30359) );
  NAND2X0 U12807 ( .IN1(n8650), .IN2(g1959), .QN(n12268) );
  NAND3X0 U12808 ( .IN1(n3611), .IN2(n12269), .IN3(n314), .QN(n12267) );
  XOR2X1 U12809 ( .IN1(n7916), .IN2(n7746), .Q(n12269) );
  NAND2X0 U12810 ( .IN1(n12270), .IN2(g1964), .QN(n12266) );
  NAND2X0 U12811 ( .IN1(n11165), .IN2(n12271), .QN(n12270) );
  NAND2X0 U12812 ( .IN1(n11177), .IN2(n8526), .QN(n12271) );
  NAND2X0 U12813 ( .IN1(n12272), .IN2(n12273), .QN(g30358) );
  NAND2X0 U12814 ( .IN1(n8644), .IN2(g1882), .QN(n12273) );
  NAND2X0 U12815 ( .IN1(n12274), .IN2(n8526), .QN(n12272) );
  NAND2X0 U12816 ( .IN1(n12275), .IN2(n12276), .QN(n12274) );
  NAND2X0 U12817 ( .IN1(n12277), .IN2(g1902), .QN(n12276) );
  NAND2X0 U12818 ( .IN1(n12278), .IN2(n12279), .QN(n12275) );
  NAND2X0 U12819 ( .IN1(g1906), .IN2(n8205), .QN(n12279) );
  INVX0 U12820 ( .INP(n12277), .ZN(n12278) );
  NAND3X0 U12821 ( .IN1(n12280), .IN2(g1917), .IN3(n5510), .QN(n12277) );
  NAND3X0 U12822 ( .IN1(n12281), .IN2(n12282), .IN3(n12283), .QN(g30357) );
  OR2X1 U12823 ( .IN1(n12284), .IN2(n5892), .Q(n12283) );
  NAND2X0 U12824 ( .IN1(n12285), .IN2(g1854), .QN(n12282) );
  NAND2X0 U12825 ( .IN1(n12286), .IN2(n8526), .QN(n12285) );
  OR2X1 U12826 ( .IN1(n12287), .IN2(n5464), .Q(n12286) );
  NAND3X0 U12827 ( .IN1(n12288), .IN2(n5464), .IN3(n5785), .QN(n12281) );
  NAND2X0 U12828 ( .IN1(n12289), .IN2(n12290), .QN(g30356) );
  NAND2X0 U12829 ( .IN1(n12291), .IN2(g1854), .QN(n12290) );
  NAND2X0 U12830 ( .IN1(n12284), .IN2(g1848), .QN(n12289) );
  NAND3X0 U12831 ( .IN1(n12292), .IN2(n12293), .IN3(n12294), .QN(g30355) );
  NAND2X0 U12832 ( .IN1(n8639), .IN2(g1830), .QN(n12294) );
  NAND2X0 U12833 ( .IN1(n12291), .IN2(g1834), .QN(n12293) );
  INVX0 U12834 ( .INP(n12284), .ZN(n12291) );
  NAND2X0 U12835 ( .IN1(n12287), .IN2(n8526), .QN(n12284) );
  NAND2X0 U12836 ( .IN1(n12288), .IN2(n5665), .QN(n12292) );
  NAND3X0 U12837 ( .IN1(n12295), .IN2(n12296), .IN3(n12297), .QN(g30354) );
  NAND2X0 U12838 ( .IN1(n8635), .IN2(g1825), .QN(n12297) );
  NAND3X0 U12839 ( .IN1(n3628), .IN2(n12298), .IN3(n709), .QN(n12296) );
  XOR2X1 U12840 ( .IN1(n7909), .IN2(n7747), .Q(n12298) );
  NAND2X0 U12841 ( .IN1(n12299), .IN2(g1830), .QN(n12295) );
  NAND2X0 U12842 ( .IN1(n11186), .IN2(n12300), .QN(n12299) );
  NAND2X0 U12843 ( .IN1(n11198), .IN2(n8526), .QN(n12300) );
  NAND2X0 U12844 ( .IN1(n12301), .IN2(n12302), .QN(g30353) );
  NAND2X0 U12845 ( .IN1(n8585), .IN2(g1748), .QN(n12302) );
  NAND2X0 U12846 ( .IN1(n12303), .IN2(n8526), .QN(n12301) );
  NAND2X0 U12847 ( .IN1(n12304), .IN2(n12305), .QN(n12303) );
  NAND2X0 U12848 ( .IN1(n12306), .IN2(g1768), .QN(n12305) );
  NAND2X0 U12849 ( .IN1(n12307), .IN2(n12308), .QN(n12304) );
  NAND2X0 U12850 ( .IN1(n5352), .IN2(g1772), .QN(n12308) );
  INVX0 U12851 ( .INP(n12306), .ZN(n12307) );
  NAND3X0 U12852 ( .IN1(n12309), .IN2(g1783), .IN3(n5359), .QN(n12306) );
  NAND3X0 U12853 ( .IN1(n12310), .IN2(n12311), .IN3(n12312), .QN(g30352) );
  OR2X1 U12854 ( .IN1(n12313), .IN2(n14521), .Q(n12312) );
  NAND2X0 U12855 ( .IN1(n12314), .IN2(g1720), .QN(n12311) );
  NAND2X0 U12856 ( .IN1(n12315), .IN2(n8526), .QN(n12314) );
  NAND2X0 U12857 ( .IN1(n12316), .IN2(g1714), .QN(n12315) );
  NAND4X0 U12858 ( .IN1(n5460), .IN2(n8505), .IN3(n12316), .IN4(n5780), .QN(
        n12310) );
  NAND2X0 U12859 ( .IN1(n12317), .IN2(n12318), .QN(g30351) );
  NAND2X0 U12860 ( .IN1(n12319), .IN2(g1720), .QN(n12318) );
  NAND2X0 U12861 ( .IN1(n12313), .IN2(g1714), .QN(n12317) );
  INVX0 U12862 ( .INP(n12319), .ZN(n12313) );
  NAND3X0 U12863 ( .IN1(n12320), .IN2(n12321), .IN3(n12322), .QN(g30350) );
  NAND2X0 U12864 ( .IN1(n12319), .IN2(g1700), .QN(n12322) );
  NOR2X0 U12865 ( .IN1(n12316), .IN2(n8557), .QN(n12319) );
  NAND3X0 U12866 ( .IN1(n12316), .IN2(n5417), .IN3(n8496), .QN(n12321) );
  NAND2X0 U12867 ( .IN1(n8587), .IN2(g1696), .QN(n12320) );
  NAND3X0 U12868 ( .IN1(n12323), .IN2(n12324), .IN3(n12325), .QN(g30349) );
  NAND2X0 U12869 ( .IN1(n8584), .IN2(g1691), .QN(n12325) );
  NAND3X0 U12870 ( .IN1(n3646), .IN2(n12326), .IN3(n1123), .QN(n12324) );
  XOR2X1 U12871 ( .IN1(n7913), .IN2(n7751), .Q(n12326) );
  NAND2X0 U12872 ( .IN1(n12327), .IN2(g1696), .QN(n12323) );
  NAND2X0 U12873 ( .IN1(n11207), .IN2(n12328), .QN(n12327) );
  NAND2X0 U12874 ( .IN1(n11221), .IN2(n8526), .QN(n12328) );
  NAND3X0 U12875 ( .IN1(n12329), .IN2(n12330), .IN3(n12331), .QN(g30348) );
  NAND2X0 U12876 ( .IN1(n8583), .IN2(g1612), .QN(n12331) );
  NAND3X0 U12877 ( .IN1(g31863), .IN2(n10793), .IN3(n3646), .QN(n12330) );
  NAND2X0 U12878 ( .IN1(n5362), .IN2(g1636), .QN(n10793) );
  NAND2X0 U12879 ( .IN1(n12332), .IN2(g1632), .QN(n12329) );
  NAND2X0 U12880 ( .IN1(n11207), .IN2(n12333), .QN(n12332) );
  OR2X1 U12881 ( .IN1(g31863), .IN2(n8545), .Q(n12333) );
  NAND2X0 U12882 ( .IN1(n12334), .IN2(n12335), .QN(g30347) );
  NAND3X0 U12883 ( .IN1(n12336), .IN2(n12337), .IN3(n12338), .QN(n12335) );
  NAND2X0 U12884 ( .IN1(n12339), .IN2(n12340), .QN(n12336) );
  INVX0 U12885 ( .INP(n12341), .ZN(n12340) );
  NAND2X0 U12886 ( .IN1(n8511), .IN2(g1413), .QN(n12339) );
  OR2X1 U12887 ( .IN1(n8477), .IN2(n7862), .Q(n12334) );
  NAND2X0 U12888 ( .IN1(n12342), .IN2(n12343), .QN(g30346) );
  NAND2X0 U12889 ( .IN1(n8582), .IN2(g1536), .QN(n12343) );
  NAND3X0 U12890 ( .IN1(n12338), .IN2(n12344), .IN3(n8496), .QN(n12342) );
  XOR2X1 U12891 ( .IN1(n12345), .IN2(n7862), .Q(n12344) );
  INVX0 U12892 ( .INP(n12346), .ZN(n12338) );
  NAND2X0 U12893 ( .IN1(n12347), .IN2(n12348), .QN(g30345) );
  NAND2X0 U12894 ( .IN1(n12349), .IN2(n8526), .QN(n12348) );
  OR2X1 U12895 ( .IN1(n12346), .IN2(n10598), .Q(n12349) );
  NAND2X0 U12896 ( .IN1(n12350), .IN2(g1514), .QN(n12347) );
  NAND2X0 U12897 ( .IN1(n12351), .IN2(n8526), .QN(n12350) );
  XOR2X1 U12898 ( .IN1(test_so49), .IN2(n5302), .Q(n12351) );
  NOR2X0 U12899 ( .IN1(n8576), .IN2(n12352), .QN(g30344) );
  NOR2X0 U12900 ( .IN1(n12346), .IN2(n12353), .QN(n12352) );
  XOR2X1 U12901 ( .IN1(n5364), .IN2(n5302), .Q(n12353) );
  NAND2X0 U12902 ( .IN1(n12354), .IN2(n12355), .QN(n12346) );
  NAND2X0 U12903 ( .IN1(n4172), .IN2(n10598), .QN(n12355) );
  AND4X1 U12904 ( .IN1(n7995), .IN2(n4895), .IN3(n12356), .IN4(g1521), .Q(
        n4172) );
  NAND3X0 U12905 ( .IN1(n12357), .IN2(n12358), .IN3(n12359), .QN(g30343) );
  NAND2X0 U12906 ( .IN1(n4175), .IN2(n11225), .QN(n12359) );
  NAND2X0 U12907 ( .IN1(n8581), .IN2(g1345), .QN(n12358) );
  NAND3X0 U12908 ( .IN1(n11343), .IN2(g1361), .IN3(n8496), .QN(n12357) );
  NAND2X0 U12909 ( .IN1(n12360), .IN2(n12361), .QN(n11343) );
  NAND2X0 U12910 ( .IN1(n7836), .IN2(n10801), .QN(n12361) );
  NAND3X0 U12911 ( .IN1(n12362), .IN2(n12363), .IN3(n12364), .QN(g30342) );
  OR2X1 U12912 ( .IN1(n8477), .IN2(n5558), .Q(n12364) );
  OR3X1 U12913 ( .IN1(n10807), .IN2(n3736), .IN3(n5553), .Q(n12363) );
  NAND2X0 U12914 ( .IN1(n3736), .IN2(n5553), .QN(n12362) );
  NAND2X0 U12915 ( .IN1(n12365), .IN2(n12366), .QN(g30341) );
  NAND3X0 U12916 ( .IN1(n12367), .IN2(n12368), .IN3(n12369), .QN(n12366) );
  NAND2X0 U12917 ( .IN1(n12370), .IN2(n12371), .QN(n12367) );
  INVX0 U12918 ( .INP(n12372), .ZN(n12371) );
  NAND2X0 U12919 ( .IN1(n8511), .IN2(g1070), .QN(n12370) );
  OR2X1 U12920 ( .IN1(n8477), .IN2(n7863), .Q(n12365) );
  NAND2X0 U12921 ( .IN1(n12373), .IN2(n12374), .QN(g30340) );
  NAND2X0 U12922 ( .IN1(n8641), .IN2(g1193), .QN(n12374) );
  NAND3X0 U12923 ( .IN1(n12369), .IN2(n12375), .IN3(n8496), .QN(n12373) );
  XOR2X1 U12924 ( .IN1(n12376), .IN2(n7863), .Q(n12375) );
  INVX0 U12925 ( .INP(n12377), .ZN(n12369) );
  NAND2X0 U12926 ( .IN1(n12378), .IN2(n12379), .QN(g30339) );
  NAND2X0 U12927 ( .IN1(n12380), .IN2(n8526), .QN(n12379) );
  OR2X1 U12928 ( .IN1(n12377), .IN2(n10756), .Q(n12380) );
  NAND2X0 U12929 ( .IN1(n12381), .IN2(g1171), .QN(n12378) );
  NAND2X0 U12930 ( .IN1(n12382), .IN2(n8526), .QN(n12381) );
  XOR2X1 U12931 ( .IN1(g1183), .IN2(n5304), .Q(n12382) );
  NOR2X0 U12932 ( .IN1(n8576), .IN2(n12383), .QN(g30338) );
  NOR2X0 U12933 ( .IN1(n12377), .IN2(n12384), .QN(n12383) );
  XOR2X1 U12934 ( .IN1(n5363), .IN2(n5304), .Q(n12384) );
  NAND2X0 U12935 ( .IN1(n12385), .IN2(n12386), .QN(n12377) );
  NAND2X0 U12936 ( .IN1(n4190), .IN2(n10756), .QN(n12386) );
  AND4X1 U12937 ( .IN1(n5642), .IN2(n4920), .IN3(n12387), .IN4(g1178), .Q(
        n4190) );
  NAND3X0 U12938 ( .IN1(n12388), .IN2(n12389), .IN3(n12390), .QN(g30337) );
  NAND2X0 U12939 ( .IN1(n4193), .IN2(n11239), .QN(n12390) );
  NAND2X0 U12940 ( .IN1(n8580), .IN2(g1002), .QN(n12389) );
  NAND3X0 U12941 ( .IN1(n11351), .IN2(g1018), .IN3(n8496), .QN(n12388) );
  NAND2X0 U12942 ( .IN1(n12391), .IN2(n12392), .QN(n11351) );
  NAND2X0 U12943 ( .IN1(n7837), .IN2(n10814), .QN(n12392) );
  NAND3X0 U12944 ( .IN1(n12393), .IN2(n12394), .IN3(n12395), .QN(g30336) );
  OR2X1 U12945 ( .IN1(n8478), .IN2(n5559), .Q(n12395) );
  OR3X1 U12946 ( .IN1(n10820), .IN2(n3741), .IN3(n5560), .Q(n12394) );
  NAND2X0 U12947 ( .IN1(n3741), .IN2(n5560), .QN(n12393) );
  NAND3X0 U12948 ( .IN1(n12396), .IN2(n12397), .IN3(n12398), .QN(g30335) );
  NAND2X0 U12949 ( .IN1(test_so60), .IN2(n8567), .QN(n12398) );
  NAND3X0 U12950 ( .IN1(n2404), .IN2(n12399), .IN3(g744), .QN(n12397) );
  NAND2X0 U12951 ( .IN1(n43), .IN2(n5470), .QN(n12396) );
  INVX0 U12952 ( .INP(n12399), .ZN(n43) );
  NAND3X0 U12953 ( .IN1(test_so60), .IN2(n4198), .IN3(n12400), .QN(n12399) );
  OR2X1 U12954 ( .IN1(g736), .IN2(n5482), .Q(n4198) );
  NAND3X0 U12955 ( .IN1(n12401), .IN2(n12402), .IN3(n12403), .QN(g30334) );
  NAND2X0 U12956 ( .IN1(n8579), .IN2(g586), .QN(n12403) );
  NAND3X0 U12957 ( .IN1(n2421), .IN2(n12404), .IN3(g577), .QN(n12402) );
  INVX0 U12958 ( .INP(n3745), .ZN(n12404) );
  NAND2X0 U12959 ( .IN1(n3745), .IN2(n5294), .QN(n12401) );
  NAND2X0 U12960 ( .IN1(n12405), .IN2(n12406), .QN(g30333) );
  NAND2X0 U12961 ( .IN1(n11370), .IN2(n12407), .QN(n12406) );
  XOR2X1 U12962 ( .IN1(test_so73), .IN2(n11373), .Q(n12407) );
  INVX0 U12963 ( .INP(n9761), .ZN(n11370) );
  NAND2X0 U12964 ( .IN1(n11372), .IN2(n8525), .QN(n9761) );
  AND3X1 U12965 ( .IN1(n12408), .IN2(g691), .IN3(n12409), .Q(n11372) );
  NAND2X0 U12966 ( .IN1(n11373), .IN2(n12410), .QN(n12409) );
  OR3X1 U12967 ( .IN1(g174), .IN2(test_so72), .IN3(g168), .Q(n12410) );
  NAND2X0 U12968 ( .IN1(n8646), .IN2(g142), .QN(n12405) );
  NAND3X0 U12969 ( .IN1(n12411), .IN2(n12412), .IN3(n12413), .QN(g29309) );
  NAND2X0 U12970 ( .IN1(n3765), .IN2(n12414), .QN(n12413) );
  OR2X1 U12971 ( .IN1(n5739), .IN2(n10354), .Q(n12414) );
  NAND3X0 U12972 ( .IN1(n12415), .IN2(g6541), .IN3(n11401), .QN(n12411) );
  NAND3X0 U12973 ( .IN1(n12416), .IN2(n12417), .IN3(n12418), .QN(g29308) );
  NAND2X0 U12974 ( .IN1(n8638), .IN2(g6523), .QN(n12418) );
  NAND2X0 U12975 ( .IN1(n12419), .IN2(g6527), .QN(n12417) );
  NAND2X0 U12976 ( .IN1(n5659), .IN2(n12420), .QN(n12416) );
  NAND3X0 U12977 ( .IN1(n12421), .IN2(n12422), .IN3(n12423), .QN(g29307) );
  NAND2X0 U12978 ( .IN1(n12419), .IN2(g6523), .QN(n12423) );
  NAND2X0 U12979 ( .IN1(n12424), .IN2(g6519), .QN(n12422) );
  NAND2X0 U12980 ( .IN1(n12425), .IN2(n8525), .QN(n12424) );
  NAND2X0 U12981 ( .IN1(n12426), .IN2(g6513), .QN(n12425) );
  NAND3X0 U12982 ( .IN1(n5426), .IN2(n12420), .IN3(n5806), .QN(n12421) );
  NAND2X0 U12983 ( .IN1(n12427), .IN2(n12428), .QN(g29306) );
  NAND2X0 U12984 ( .IN1(n12419), .IN2(g6519), .QN(n12428) );
  OR2X1 U12985 ( .IN1(n12419), .IN2(n5426), .Q(n12427) );
  NAND3X0 U12986 ( .IN1(n12429), .IN2(n12430), .IN3(n12431), .QN(g29305) );
  NAND2X0 U12987 ( .IN1(n12419), .IN2(g6509), .QN(n12431) );
  NOR2X0 U12988 ( .IN1(n12426), .IN2(n8557), .QN(n12419) );
  NAND2X0 U12989 ( .IN1(n12432), .IN2(g6500), .QN(n12430) );
  NAND2X0 U12990 ( .IN1(n12433), .IN2(n8525), .QN(n12432) );
  NAND2X0 U12991 ( .IN1(n7792), .IN2(n12426), .QN(n12433) );
  NAND3X0 U12992 ( .IN1(n12420), .IN2(g6505), .IN3(n5748), .QN(n12429) );
  AND2X1 U12993 ( .IN1(n12426), .IN2(n8508), .Q(n12420) );
  NOR2X0 U12994 ( .IN1(n12434), .IN2(n8198), .QN(n12426) );
  NAND3X0 U12995 ( .IN1(n12435), .IN2(n12436), .IN3(n12437), .QN(g29304) );
  NAND2X0 U12996 ( .IN1(n10372), .IN2(g6500), .QN(n12437) );
  NAND2X0 U12997 ( .IN1(n8578), .IN2(g6505), .QN(n12436) );
  NAND3X0 U12998 ( .IN1(n10365), .IN2(n12438), .IN3(n8496), .QN(n12435) );
  XNOR2X1 U12999 ( .IN1(n12439), .IN2(n12440), .Q(n12438) );
  NAND2X0 U13000 ( .IN1(g6500), .IN2(n12434), .QN(n12439) );
  NAND3X0 U13001 ( .IN1(g6727), .IN2(g17722), .IN3(n8821), .QN(n12434) );
  NAND3X0 U13002 ( .IN1(n12441), .IN2(n12412), .IN3(n12442), .QN(g29303) );
  NAND2X0 U13003 ( .IN1(n3765), .IN2(n12443), .QN(n12442) );
  NAND2X0 U13004 ( .IN1(g6195), .IN2(n10344), .QN(n12443) );
  NAND3X0 U13005 ( .IN1(n12415), .IN2(g6195), .IN3(n11482), .QN(n12441) );
  NAND3X0 U13006 ( .IN1(n12444), .IN2(n12445), .IN3(n12446), .QN(g29302) );
  NAND2X0 U13007 ( .IN1(n8645), .IN2(g6177), .QN(n12446) );
  NAND2X0 U13008 ( .IN1(n12447), .IN2(g6181), .QN(n12445) );
  NAND2X0 U13009 ( .IN1(n5667), .IN2(n12448), .QN(n12444) );
  NAND3X0 U13010 ( .IN1(n12449), .IN2(n12450), .IN3(n12451), .QN(g29301) );
  NAND2X0 U13011 ( .IN1(n12447), .IN2(g6177), .QN(n12451) );
  NAND2X0 U13012 ( .IN1(n12452), .IN2(g6173), .QN(n12450) );
  NAND2X0 U13013 ( .IN1(n12453), .IN2(n8525), .QN(n12452) );
  NAND2X0 U13014 ( .IN1(n12454), .IN2(g6167), .QN(n12453) );
  NAND3X0 U13015 ( .IN1(n5430), .IN2(n12448), .IN3(n5810), .QN(n12449) );
  NAND2X0 U13016 ( .IN1(n12455), .IN2(n12456), .QN(g29300) );
  NAND2X0 U13017 ( .IN1(n12447), .IN2(g6173), .QN(n12456) );
  OR2X1 U13018 ( .IN1(n12447), .IN2(n5430), .Q(n12455) );
  NAND3X0 U13019 ( .IN1(n12457), .IN2(n12458), .IN3(n12459), .QN(g29299) );
  NAND2X0 U13020 ( .IN1(n12447), .IN2(g6163), .QN(n12459) );
  NOR2X0 U13021 ( .IN1(n12454), .IN2(n8558), .QN(n12447) );
  NAND2X0 U13022 ( .IN1(n12460), .IN2(g6154), .QN(n12458) );
  NAND2X0 U13023 ( .IN1(n12461), .IN2(n8525), .QN(n12460) );
  NAND2X0 U13024 ( .IN1(n7791), .IN2(n12454), .QN(n12461) );
  INVX0 U13025 ( .INP(n12462), .ZN(n12454) );
  NAND3X0 U13026 ( .IN1(n12448), .IN2(g6159), .IN3(n5747), .QN(n12457) );
  NOR2X0 U13027 ( .IN1(n12462), .IN2(n8562), .QN(n12448) );
  NAND2X0 U13028 ( .IN1(n12463), .IN2(n10377), .QN(n12462) );
  NAND3X0 U13029 ( .IN1(n12464), .IN2(n12465), .IN3(n12466), .QN(g29298) );
  NAND2X0 U13030 ( .IN1(n10387), .IN2(g6154), .QN(n12466) );
  NAND2X0 U13031 ( .IN1(n8587), .IN2(g6159), .QN(n12465) );
  NAND3X0 U13032 ( .IN1(n10377), .IN2(n12467), .IN3(n8495), .QN(n12464) );
  XOR2X1 U13033 ( .IN1(n12468), .IN2(n12469), .Q(n12467) );
  NOR2X0 U13034 ( .IN1(n12463), .IN2(n5747), .QN(n12469) );
  AND3X1 U13035 ( .IN1(n9612), .IN2(g17685), .IN3(test_so69), .Q(n12463) );
  NAND3X0 U13036 ( .IN1(n12470), .IN2(n12412), .IN3(n12471), .QN(g29297) );
  NAND2X0 U13037 ( .IN1(n3765), .IN2(n12472), .QN(n12471) );
  NAND2X0 U13038 ( .IN1(g5849), .IN2(n10343), .QN(n12472) );
  NAND3X0 U13039 ( .IN1(n12415), .IN2(g5849), .IN3(n11563), .QN(n12470) );
  NAND3X0 U13040 ( .IN1(n12473), .IN2(n12474), .IN3(n12475), .QN(g29296) );
  NAND2X0 U13041 ( .IN1(n8586), .IN2(g5831), .QN(n12475) );
  NAND2X0 U13042 ( .IN1(n12476), .IN2(g5835), .QN(n12474) );
  NAND2X0 U13043 ( .IN1(n5663), .IN2(n12477), .QN(n12473) );
  NAND3X0 U13044 ( .IN1(n12478), .IN2(n12479), .IN3(n12480), .QN(g29295) );
  NAND2X0 U13045 ( .IN1(n12476), .IN2(g5831), .QN(n12480) );
  NAND2X0 U13046 ( .IN1(n12481), .IN2(g5827), .QN(n12479) );
  NAND2X0 U13047 ( .IN1(n12482), .IN2(n8525), .QN(n12481) );
  NAND2X0 U13048 ( .IN1(n12483), .IN2(g5821), .QN(n12482) );
  NAND3X0 U13049 ( .IN1(n5429), .IN2(n12477), .IN3(n5809), .QN(n12478) );
  NAND2X0 U13050 ( .IN1(n12484), .IN2(n12485), .QN(g29294) );
  NAND2X0 U13051 ( .IN1(n12476), .IN2(g5827), .QN(n12485) );
  OR2X1 U13052 ( .IN1(n12476), .IN2(n5429), .Q(n12484) );
  NAND3X0 U13053 ( .IN1(n12486), .IN2(n12487), .IN3(n12488), .QN(g29293) );
  NAND2X0 U13054 ( .IN1(n12476), .IN2(g5817), .QN(n12488) );
  NOR2X0 U13055 ( .IN1(n12483), .IN2(n8564), .QN(n12476) );
  NAND2X0 U13056 ( .IN1(n12489), .IN2(g5808), .QN(n12487) );
  NAND2X0 U13057 ( .IN1(n12490), .IN2(n8525), .QN(n12489) );
  NAND2X0 U13058 ( .IN1(n7793), .IN2(n12483), .QN(n12490) );
  INVX0 U13059 ( .INP(n12491), .ZN(n12483) );
  NAND3X0 U13060 ( .IN1(n12477), .IN2(g5813), .IN3(n5749), .QN(n12486) );
  NOR2X0 U13061 ( .IN1(n12491), .IN2(n8560), .QN(n12477) );
  NAND2X0 U13062 ( .IN1(n12492), .IN2(n10392), .QN(n12491) );
  NAND3X0 U13063 ( .IN1(n12493), .IN2(n12494), .IN3(n12495), .QN(g29292) );
  NAND2X0 U13064 ( .IN1(n10402), .IN2(g5808), .QN(n12495) );
  NAND2X0 U13065 ( .IN1(n8571), .IN2(g5813), .QN(n12494) );
  NAND3X0 U13066 ( .IN1(n10392), .IN2(n12496), .IN3(n8495), .QN(n12493) );
  XOR2X1 U13067 ( .IN1(n12497), .IN2(n12498), .Q(n12496) );
  NOR2X0 U13068 ( .IN1(n12492), .IN2(n5749), .QN(n12498) );
  AND3X1 U13069 ( .IN1(g6035), .IN2(g17646), .IN3(n9617), .Q(n12492) );
  NAND3X0 U13070 ( .IN1(n12499), .IN2(n12412), .IN3(n12500), .QN(g29291) );
  NAND2X0 U13071 ( .IN1(n3765), .IN2(n12501), .QN(n12500) );
  OR2X1 U13072 ( .IN1(n5737), .IN2(n10339), .Q(n12501) );
  NAND3X0 U13073 ( .IN1(n12415), .IN2(g5503), .IN3(n11644), .QN(n12499) );
  NAND3X0 U13074 ( .IN1(n12502), .IN2(n12503), .IN3(n12504), .QN(g29290) );
  NAND2X0 U13075 ( .IN1(n8570), .IN2(g5485), .QN(n12504) );
  NAND2X0 U13076 ( .IN1(n12505), .IN2(g5489), .QN(n12503) );
  NAND2X0 U13077 ( .IN1(n5660), .IN2(n12506), .QN(n12502) );
  NAND3X0 U13078 ( .IN1(n12507), .IN2(n12508), .IN3(n12509), .QN(g29289) );
  NAND2X0 U13079 ( .IN1(n12505), .IN2(g5485), .QN(n12509) );
  NAND2X0 U13080 ( .IN1(n12510), .IN2(g5481), .QN(n12508) );
  NAND2X0 U13081 ( .IN1(n12511), .IN2(n8525), .QN(n12510) );
  NAND2X0 U13082 ( .IN1(n12512), .IN2(g5475), .QN(n12511) );
  NAND3X0 U13083 ( .IN1(n5425), .IN2(n12506), .IN3(n5805), .QN(n12507) );
  NAND2X0 U13084 ( .IN1(n12513), .IN2(n12514), .QN(g29288) );
  NAND2X0 U13085 ( .IN1(n12505), .IN2(g5481), .QN(n12514) );
  OR2X1 U13086 ( .IN1(n12505), .IN2(n5425), .Q(n12513) );
  NAND3X0 U13087 ( .IN1(n12515), .IN2(n12516), .IN3(n12517), .QN(g29287) );
  NAND2X0 U13088 ( .IN1(n12505), .IN2(g5471), .QN(n12517) );
  NOR2X0 U13089 ( .IN1(n12512), .IN2(n8564), .QN(n12505) );
  NAND2X0 U13090 ( .IN1(n12518), .IN2(g5462), .QN(n12516) );
  NAND2X0 U13091 ( .IN1(n12519), .IN2(n8525), .QN(n12518) );
  NAND2X0 U13092 ( .IN1(n7775), .IN2(n12512), .QN(n12519) );
  INVX0 U13093 ( .INP(n12520), .ZN(n12512) );
  NAND3X0 U13094 ( .IN1(n12506), .IN2(g5467), .IN3(n5744), .QN(n12515) );
  NOR2X0 U13095 ( .IN1(n12520), .IN2(n8563), .QN(n12506) );
  NAND2X0 U13096 ( .IN1(n12521), .IN2(n10407), .QN(n12520) );
  NAND3X0 U13097 ( .IN1(n12522), .IN2(n12523), .IN3(n12524), .QN(g29286) );
  NAND2X0 U13098 ( .IN1(n10417), .IN2(g5462), .QN(n12524) );
  NAND2X0 U13099 ( .IN1(n8569), .IN2(g5467), .QN(n12523) );
  NAND3X0 U13100 ( .IN1(n10407), .IN2(n12525), .IN3(n8495), .QN(n12522) );
  XOR2X1 U13101 ( .IN1(n12526), .IN2(n12527), .Q(n12525) );
  NOR2X0 U13102 ( .IN1(n12521), .IN2(n5744), .QN(n12527) );
  AND3X1 U13103 ( .IN1(g5689), .IN2(g17604), .IN3(n9625), .Q(n12521) );
  NAND3X0 U13104 ( .IN1(n12528), .IN2(n12412), .IN3(n12529), .QN(g29285) );
  NAND2X0 U13105 ( .IN1(n3765), .IN2(n12530), .QN(n12529) );
  OR2X1 U13106 ( .IN1(n5734), .IN2(g26801), .Q(n12530) );
  NAND3X0 U13107 ( .IN1(n12415), .IN2(g5156), .IN3(n11724), .QN(n12528) );
  NAND3X0 U13108 ( .IN1(n12531), .IN2(n12532), .IN3(n12533), .QN(g29284) );
  NAND2X0 U13109 ( .IN1(n8587), .IN2(g5138), .QN(n12533) );
  NAND2X0 U13110 ( .IN1(n12534), .IN2(g5142), .QN(n12532) );
  NAND2X0 U13111 ( .IN1(n5658), .IN2(n12535), .QN(n12531) );
  NAND3X0 U13112 ( .IN1(n12536), .IN2(n12537), .IN3(n12538), .QN(g29283) );
  NAND2X0 U13113 ( .IN1(n12534), .IN2(g5138), .QN(n12538) );
  NAND2X0 U13114 ( .IN1(n12539), .IN2(g5134), .QN(n12537) );
  NAND2X0 U13115 ( .IN1(n12540), .IN2(n8525), .QN(n12539) );
  NAND2X0 U13116 ( .IN1(test_so96), .IN2(n12541), .QN(n12540) );
  NAND3X0 U13117 ( .IN1(n12535), .IN2(n8211), .IN3(n5807), .QN(n12536) );
  NAND2X0 U13118 ( .IN1(n12542), .IN2(n12543), .QN(g29282) );
  NAND2X0 U13119 ( .IN1(n12534), .IN2(g5134), .QN(n12543) );
  OR2X1 U13120 ( .IN1(n8211), .IN2(n12534), .Q(n12542) );
  NOR2X0 U13121 ( .IN1(n12541), .IN2(n8562), .QN(n12534) );
  NAND3X0 U13122 ( .IN1(n12544), .IN2(n12545), .IN3(n12546), .QN(g29281) );
  NAND2X0 U13123 ( .IN1(n11396), .IN2(n12547), .QN(n12546) );
  NOR2X0 U13124 ( .IN1(n8570), .IN2(n7709), .QN(n11396) );
  NAND2X0 U13125 ( .IN1(n12548), .IN2(g5115), .QN(n12545) );
  NAND2X0 U13126 ( .IN1(n12549), .IN2(n8525), .QN(n12548) );
  NAND2X0 U13127 ( .IN1(n7774), .IN2(n12541), .QN(n12549) );
  INVX0 U13128 ( .INP(n12547), .ZN(n12541) );
  NAND3X0 U13129 ( .IN1(n12535), .IN2(g5120), .IN3(n5743), .QN(n12544) );
  NOR2X0 U13130 ( .IN1(n12547), .IN2(n8563), .QN(n12535) );
  NAND2X0 U13131 ( .IN1(n12550), .IN2(g33959), .QN(n12547) );
  NAND3X0 U13132 ( .IN1(n12551), .IN2(n12552), .IN3(n12553), .QN(g29280) );
  NAND2X0 U13133 ( .IN1(n10429), .IN2(g5115), .QN(n12553) );
  NAND2X0 U13134 ( .IN1(n8658), .IN2(g5120), .QN(n12552) );
  NAND3X0 U13135 ( .IN1(g33959), .IN2(n12554), .IN3(n8495), .QN(n12551) );
  XOR2X1 U13136 ( .IN1(n12555), .IN2(n12556), .Q(n12554) );
  NOR2X0 U13137 ( .IN1(n12550), .IN2(n5743), .QN(n12556) );
  AND3X1 U13138 ( .IN1(g31860), .IN2(g17577), .IN3(test_so10), .Q(n12550) );
  OR2X1 U13139 ( .IN1(n12557), .IN2(g29279), .Q(g29278) );
  NOR2X0 U13140 ( .IN1(n7770), .IN2(n8505), .QN(n12557) );
  OR2X1 U13141 ( .IN1(n12558), .IN2(g29277), .Q(g29276) );
  AND2X1 U13142 ( .IN1(n8568), .IN2(test_so100), .Q(n12558) );
  NAND2X0 U13143 ( .IN1(n12559), .IN2(n12560), .QN(g29275) );
  NAND2X0 U13144 ( .IN1(n12561), .IN2(n11816), .QN(n12560) );
  XOR2X1 U13145 ( .IN1(n11334), .IN2(g4087), .Q(n12561) );
  NOR2X0 U13146 ( .IN1(n8220), .IN2(n12562), .QN(n11334) );
  NAND2X0 U13147 ( .IN1(test_so11), .IN2(n8661), .QN(n12559) );
  NAND3X0 U13148 ( .IN1(n12563), .IN2(n12412), .IN3(n12564), .QN(g29274) );
  NAND2X0 U13149 ( .IN1(n3765), .IN2(n12565), .QN(n12564) );
  NAND2X0 U13150 ( .IN1(g3849), .IN2(n10353), .QN(n12565) );
  NAND3X0 U13151 ( .IN1(n12415), .IN2(g3849), .IN3(n11820), .QN(n12563) );
  NAND3X0 U13152 ( .IN1(n12566), .IN2(n12567), .IN3(n12568), .QN(g29273) );
  NAND2X0 U13153 ( .IN1(n8613), .IN2(g3831), .QN(n12568) );
  NAND2X0 U13154 ( .IN1(n12569), .IN2(g3835), .QN(n12567) );
  NAND2X0 U13155 ( .IN1(n5662), .IN2(n12570), .QN(n12566) );
  NAND3X0 U13156 ( .IN1(n12571), .IN2(n12572), .IN3(n12573), .QN(g29272) );
  NAND2X0 U13157 ( .IN1(n12569), .IN2(g3831), .QN(n12573) );
  NAND2X0 U13158 ( .IN1(n12574), .IN2(g3827), .QN(n12572) );
  NAND2X0 U13159 ( .IN1(n12575), .IN2(n8525), .QN(n12574) );
  NAND2X0 U13160 ( .IN1(n12576), .IN2(g3821), .QN(n12575) );
  NAND3X0 U13161 ( .IN1(n5428), .IN2(n12570), .IN3(n5808), .QN(n12571) );
  NAND2X0 U13162 ( .IN1(n12577), .IN2(n12578), .QN(g29271) );
  NAND2X0 U13163 ( .IN1(n12569), .IN2(g3827), .QN(n12578) );
  OR2X1 U13164 ( .IN1(n12569), .IN2(n5428), .Q(n12577) );
  NOR2X0 U13165 ( .IN1(n12576), .IN2(n8561), .QN(n12569) );
  NAND3X0 U13166 ( .IN1(n12579), .IN2(n12580), .IN3(n12581), .QN(g29270) );
  NAND2X0 U13167 ( .IN1(n11378), .IN2(n12582), .QN(n12581) );
  NOR2X0 U13168 ( .IN1(n8571), .IN2(n7710), .QN(n11378) );
  NAND2X0 U13169 ( .IN1(n12583), .IN2(g3808), .QN(n12580) );
  NAND2X0 U13170 ( .IN1(n12584), .IN2(n8525), .QN(n12583) );
  NAND2X0 U13171 ( .IN1(n7776), .IN2(n12576), .QN(n12584) );
  INVX0 U13172 ( .INP(n12582), .ZN(n12576) );
  NAND3X0 U13173 ( .IN1(n12570), .IN2(g3813), .IN3(n5745), .QN(n12579) );
  NOR2X0 U13174 ( .IN1(n12582), .IN2(n8560), .QN(n12570) );
  NAND2X0 U13175 ( .IN1(n12585), .IN2(n10444), .QN(n12582) );
  NAND3X0 U13176 ( .IN1(n12586), .IN2(n12587), .IN3(n12588), .QN(g29269) );
  NAND2X0 U13177 ( .IN1(n10454), .IN2(g3808), .QN(n12588) );
  NAND2X0 U13178 ( .IN1(n8610), .IN2(g3813), .QN(n12587) );
  NAND3X0 U13179 ( .IN1(n10444), .IN2(n12589), .IN3(n8495), .QN(n12586) );
  XOR2X1 U13180 ( .IN1(n12590), .IN2(n12591), .Q(n12589) );
  NOR2X0 U13181 ( .IN1(n12585), .IN2(n5745), .QN(n12591) );
  AND3X1 U13182 ( .IN1(g4040), .IN2(g16693), .IN3(n9613), .Q(n12585) );
  NAND3X0 U13183 ( .IN1(n12592), .IN2(n12412), .IN3(n12593), .QN(g29268) );
  NAND2X0 U13184 ( .IN1(n3765), .IN2(n12594), .QN(n12593) );
  NAND2X0 U13185 ( .IN1(g3498), .IN2(n10352), .QN(n12594) );
  NAND3X0 U13186 ( .IN1(n12415), .IN2(g3498), .IN3(n11902), .QN(n12592) );
  NAND3X0 U13187 ( .IN1(n12595), .IN2(n12596), .IN3(n12597), .QN(g29267) );
  NAND2X0 U13188 ( .IN1(n8611), .IN2(g3480), .QN(n12597) );
  NAND2X0 U13189 ( .IN1(n12598), .IN2(g3484), .QN(n12596) );
  NAND2X0 U13190 ( .IN1(n5668), .IN2(n12599), .QN(n12595) );
  NAND3X0 U13191 ( .IN1(n12600), .IN2(n12601), .IN3(n12602), .QN(g29266) );
  NAND2X0 U13192 ( .IN1(n12598), .IN2(g3480), .QN(n12602) );
  NAND2X0 U13193 ( .IN1(n12603), .IN2(g3476), .QN(n12601) );
  NAND2X0 U13194 ( .IN1(n12604), .IN2(n8525), .QN(n12603) );
  NAND2X0 U13195 ( .IN1(n12605), .IN2(g3470), .QN(n12604) );
  NAND3X0 U13196 ( .IN1(n5424), .IN2(n12599), .IN3(n5786), .QN(n12600) );
  NAND2X0 U13197 ( .IN1(n12606), .IN2(n12607), .QN(g29265) );
  NAND2X0 U13198 ( .IN1(n12598), .IN2(g3476), .QN(n12607) );
  OR2X1 U13199 ( .IN1(n12598), .IN2(n5424), .Q(n12606) );
  NAND3X0 U13200 ( .IN1(n12608), .IN2(n12609), .IN3(n12610), .QN(g29264) );
  NAND2X0 U13201 ( .IN1(n12598), .IN2(g3466), .QN(n12610) );
  NOR2X0 U13202 ( .IN1(n12605), .IN2(n8561), .QN(n12598) );
  NAND2X0 U13203 ( .IN1(test_so4), .IN2(n12611), .QN(n12609) );
  NAND2X0 U13204 ( .IN1(n12612), .IN2(n8525), .QN(n12611) );
  NAND2X0 U13205 ( .IN1(n7777), .IN2(n12605), .QN(n12612) );
  INVX0 U13206 ( .INP(n12613), .ZN(n12605) );
  NAND3X0 U13207 ( .IN1(n12599), .IN2(g3462), .IN3(n8224), .QN(n12608) );
  NOR2X0 U13208 ( .IN1(n12613), .IN2(n8562), .QN(n12599) );
  NAND2X0 U13209 ( .IN1(n12614), .IN2(n10458), .QN(n12613) );
  NAND3X0 U13210 ( .IN1(n12615), .IN2(n12616), .IN3(n12617), .QN(g29263) );
  NAND2X0 U13211 ( .IN1(test_so4), .IN2(n10468), .QN(n12617) );
  NAND2X0 U13212 ( .IN1(n8608), .IN2(g3462), .QN(n12616) );
  NAND3X0 U13213 ( .IN1(n10458), .IN2(n12618), .IN3(n8495), .QN(n12615) );
  XOR2X1 U13214 ( .IN1(n12619), .IN2(n12620), .Q(n12618) );
  NOR2X0 U13215 ( .IN1(n12614), .IN2(n8224), .QN(n12620) );
  AND3X1 U13216 ( .IN1(g3689), .IN2(g16656), .IN3(n9618), .Q(n12614) );
  NAND3X0 U13217 ( .IN1(n12621), .IN2(n12412), .IN3(n12622), .QN(g29262) );
  NAND2X0 U13218 ( .IN1(n3765), .IN2(n12623), .QN(n12622) );
  OR2X1 U13219 ( .IN1(n5738), .IN2(n10349), .Q(n12623) );
  NAND2X0 U13220 ( .IN1(n3765), .IN2(n12415), .QN(n12412) );
  NAND3X0 U13221 ( .IN1(n12415), .IN2(g3147), .IN3(n11983), .QN(n12621) );
  INVX0 U13222 ( .INP(n4210), .ZN(n12415) );
  NAND2X0 U13223 ( .IN1(n7812), .IN2(g4180), .QN(n4210) );
  NAND3X0 U13224 ( .IN1(n12624), .IN2(n12625), .IN3(n12626), .QN(g29261) );
  NAND2X0 U13225 ( .IN1(n8609), .IN2(g3129), .QN(n12626) );
  NAND2X0 U13226 ( .IN1(n12627), .IN2(g3133), .QN(n12625) );
  NAND2X0 U13227 ( .IN1(n5661), .IN2(n12628), .QN(n12624) );
  NAND3X0 U13228 ( .IN1(n12629), .IN2(n12630), .IN3(n12631), .QN(g29260) );
  NAND2X0 U13229 ( .IN1(n12627), .IN2(g3129), .QN(n12631) );
  NAND2X0 U13230 ( .IN1(n12632), .IN2(g3125), .QN(n12630) );
  NAND2X0 U13231 ( .IN1(n12633), .IN2(n8525), .QN(n12632) );
  NAND2X0 U13232 ( .IN1(n12634), .IN2(g3119), .QN(n12633) );
  NAND3X0 U13233 ( .IN1(n5423), .IN2(n12628), .IN3(n5781), .QN(n12629) );
  NAND2X0 U13234 ( .IN1(n12635), .IN2(n12636), .QN(g29259) );
  NAND2X0 U13235 ( .IN1(n12627), .IN2(g3125), .QN(n12636) );
  OR2X1 U13236 ( .IN1(n12627), .IN2(n5423), .Q(n12635) );
  NAND3X0 U13237 ( .IN1(n12637), .IN2(n12638), .IN3(n12639), .QN(g29258) );
  NAND2X0 U13238 ( .IN1(n12627), .IN2(g3115), .QN(n12639) );
  NOR2X0 U13239 ( .IN1(n12634), .IN2(n8563), .QN(n12627) );
  NAND2X0 U13240 ( .IN1(n12640), .IN2(g3106), .QN(n12638) );
  NAND2X0 U13241 ( .IN1(n12641), .IN2(n8525), .QN(n12640) );
  NAND2X0 U13242 ( .IN1(n7773), .IN2(n12634), .QN(n12641) );
  INVX0 U13243 ( .INP(n12642), .ZN(n12634) );
  NAND3X0 U13244 ( .IN1(n12628), .IN2(g3111), .IN3(n5742), .QN(n12637) );
  NOR2X0 U13245 ( .IN1(n12642), .IN2(n8563), .QN(n12628) );
  NAND2X0 U13246 ( .IN1(n12643), .IN2(n10477), .QN(n12642) );
  NAND3X0 U13247 ( .IN1(n12644), .IN2(n12645), .IN3(n12646), .QN(g29257) );
  NAND2X0 U13248 ( .IN1(n10483), .IN2(g3106), .QN(n12646) );
  NAND2X0 U13249 ( .IN1(n8600), .IN2(g3111), .QN(n12645) );
  NAND3X0 U13250 ( .IN1(n10477), .IN2(n12647), .IN3(n8495), .QN(n12644) );
  XOR2X1 U13251 ( .IN1(n12648), .IN2(n12649), .Q(n12647) );
  NOR2X0 U13252 ( .IN1(n12643), .IN2(n5742), .QN(n12649) );
  AND3X1 U13253 ( .IN1(g3338), .IN2(g16624), .IN3(n9626), .Q(n12643) );
  NAND4X0 U13254 ( .IN1(n12650), .IN2(n8807), .IN3(n12651), .IN4(n12652), .QN(
        g29256) );
  NAND3X0 U13255 ( .IN1(n12106), .IN2(g2735), .IN3(n8495), .QN(n12652) );
  NAND2X0 U13256 ( .IN1(n8601), .IN2(g2729), .QN(n12651) );
  OR2X1 U13257 ( .IN1(g2735), .IN2(n12106), .Q(n12650) );
  NAND2X0 U13258 ( .IN1(n9565), .IN2(n12078), .QN(n12106) );
  NOR2X0 U13259 ( .IN1(n7867), .IN2(n5301), .QN(n9565) );
  NAND2X0 U13260 ( .IN1(n12653), .IN2(n12654), .QN(g29255) );
  NAND2X0 U13261 ( .IN1(n12655), .IN2(g2638), .QN(n12654) );
  NAND2X0 U13262 ( .IN1(n12656), .IN2(n8525), .QN(n12655) );
  OR2X1 U13263 ( .IN1(n11057), .IN2(n8831), .Q(n12656) );
  NOR2X0 U13264 ( .IN1(n7919), .IN2(n326), .QN(n8831) );
  NAND2X0 U13265 ( .IN1(n12657), .IN2(g2652), .QN(n12653) );
  NAND2X0 U13266 ( .IN1(n11060), .IN2(n12658), .QN(n12657) );
  NAND2X0 U13267 ( .IN1(n4379), .IN2(n8525), .QN(n12658) );
  NAND4X0 U13268 ( .IN1(n12659), .IN2(n12660), .IN3(n12661), .IN4(n12662), 
        .QN(g29254) );
  NAND2X0 U13269 ( .IN1(n12114), .IN2(g2567), .QN(n12662) );
  NOR2X0 U13270 ( .IN1(n12113), .IN2(n8562), .QN(n12114) );
  NAND3X0 U13271 ( .IN1(g2587), .IN2(g2619), .IN3(n12135), .QN(n12113) );
  INVX0 U13272 ( .INP(n11057), .ZN(n12135) );
  NAND2X0 U13273 ( .IN1(n3517), .IN2(n12663), .QN(n12661) );
  NAND3X0 U13274 ( .IN1(n12664), .IN2(n12665), .IN3(n12666), .QN(n12663) );
  NAND2X0 U13275 ( .IN1(n326), .IN2(g2563), .QN(n12666) );
  INVX0 U13276 ( .INP(n11072), .ZN(n326) );
  NAND2X0 U13277 ( .IN1(n5372), .IN2(g2610), .QN(n11072) );
  NAND2X0 U13278 ( .IN1(n5508), .IN2(n12667), .QN(n12665) );
  NAND2X0 U13279 ( .IN1(n12668), .IN2(n12669), .QN(n12667) );
  NAND2X0 U13280 ( .IN1(test_so66), .IN2(n5372), .QN(n12669) );
  NAND2X0 U13281 ( .IN1(g2583), .IN2(g2610), .QN(n12668) );
  NAND2X0 U13282 ( .IN1(n8130), .IN2(n12670), .QN(n12664) );
  NAND2X0 U13283 ( .IN1(n12671), .IN2(n12672), .QN(n12670) );
  NAND2X0 U13284 ( .IN1(test_so61), .IN2(g2587), .QN(n12672) );
  NAND2X0 U13285 ( .IN1(g2619), .IN2(g2571), .QN(n12671) );
  NOR2X0 U13286 ( .IN1(n11057), .IN2(n8561), .QN(n3517) );
  NAND2X0 U13287 ( .IN1(n11066), .IN2(g2638), .QN(n12660) );
  INVX0 U13288 ( .INP(n11060), .ZN(n11066) );
  NAND2X0 U13289 ( .IN1(n11057), .IN2(n8525), .QN(n11060) );
  NAND3X0 U13290 ( .IN1(n12673), .IN2(n12674), .IN3(n12078), .QN(n11057) );
  NAND2X0 U13291 ( .IN1(n9579), .IN2(g2819), .QN(n12673) );
  NAND2X0 U13292 ( .IN1(n8595), .IN2(g2619), .QN(n12659) );
  NAND2X0 U13293 ( .IN1(n12675), .IN2(n12676), .QN(g29253) );
  NAND2X0 U13294 ( .IN1(n12677), .IN2(g2518), .QN(n12676) );
  NAND2X0 U13295 ( .IN1(n11081), .IN2(n12678), .QN(n12677) );
  NAND2X0 U13296 ( .IN1(n4391), .IN2(n8525), .QN(n12678) );
  NAND2X0 U13297 ( .IN1(n12679), .IN2(g2504), .QN(n12675) );
  NAND2X0 U13298 ( .IN1(n12680), .IN2(n8524), .QN(n12679) );
  OR2X1 U13299 ( .IN1(n11078), .IN2(n8830), .Q(n12680) );
  NOR2X0 U13300 ( .IN1(n7917), .IN2(n911), .QN(n8830) );
  NAND4X0 U13301 ( .IN1(n12681), .IN2(n12682), .IN3(n12683), .IN4(n12684), 
        .QN(g29252) );
  NAND2X0 U13302 ( .IN1(n12143), .IN2(g2433), .QN(n12684) );
  NOR2X0 U13303 ( .IN1(n12142), .IN2(n8560), .QN(n12143) );
  NAND3X0 U13304 ( .IN1(g2453), .IN2(g2485), .IN3(n12164), .QN(n12142) );
  INVX0 U13305 ( .INP(n11078), .ZN(n12164) );
  NAND2X0 U13306 ( .IN1(n3536), .IN2(n12685), .QN(n12683) );
  NAND3X0 U13307 ( .IN1(n12686), .IN2(n12687), .IN3(n12688), .QN(n12685) );
  NAND2X0 U13308 ( .IN1(n911), .IN2(g2429), .QN(n12688) );
  INVX0 U13309 ( .INP(n11093), .ZN(n911) );
  NAND2X0 U13310 ( .IN1(n5373), .IN2(g2476), .QN(n11093) );
  NAND2X0 U13311 ( .IN1(n5509), .IN2(n12689), .QN(n12687) );
  NAND2X0 U13312 ( .IN1(n12690), .IN2(n12691), .QN(n12689) );
  NAND2X0 U13313 ( .IN1(n5373), .IN2(g2441), .QN(n12691) );
  NAND2X0 U13314 ( .IN1(g2449), .IN2(g2476), .QN(n12690) );
  NAND2X0 U13315 ( .IN1(n8131), .IN2(n12692), .QN(n12686) );
  NAND2X0 U13316 ( .IN1(n12693), .IN2(n12694), .QN(n12692) );
  NAND2X0 U13317 ( .IN1(g2453), .IN2(n9274), .QN(n12694) );
  NAND2X0 U13318 ( .IN1(g2485), .IN2(g2437), .QN(n12693) );
  NOR2X0 U13319 ( .IN1(n11078), .IN2(n8558), .QN(n3536) );
  NAND2X0 U13320 ( .IN1(n11087), .IN2(g2504), .QN(n12682) );
  INVX0 U13321 ( .INP(n11081), .ZN(n11087) );
  NAND2X0 U13322 ( .IN1(n11078), .IN2(n8524), .QN(n11081) );
  NAND3X0 U13323 ( .IN1(n12695), .IN2(n12674), .IN3(n12087), .QN(n11078) );
  NAND2X0 U13324 ( .IN1(n9579), .IN2(g2815), .QN(n12695) );
  NAND2X0 U13325 ( .IN1(n8603), .IN2(g2485), .QN(n12681) );
  NAND2X0 U13326 ( .IN1(n12696), .IN2(n12697), .QN(g29251) );
  NAND2X0 U13327 ( .IN1(n12698), .IN2(g2384), .QN(n12697) );
  NAND2X0 U13328 ( .IN1(n11102), .IN2(n12699), .QN(n12698) );
  NAND2X0 U13329 ( .IN1(n4402), .IN2(n8524), .QN(n12699) );
  NAND2X0 U13330 ( .IN1(n12700), .IN2(g2370), .QN(n12696) );
  NAND2X0 U13331 ( .IN1(n12701), .IN2(n8524), .QN(n12700) );
  OR2X1 U13332 ( .IN1(n11099), .IN2(n8829), .Q(n12701) );
  NOR2X0 U13333 ( .IN1(n7911), .IN2(n456), .QN(n8829) );
  NAND4X0 U13334 ( .IN1(n12702), .IN2(n12703), .IN3(n12704), .IN4(n12705), 
        .QN(g29250) );
  NAND2X0 U13335 ( .IN1(n12172), .IN2(g2299), .QN(n12705) );
  NOR2X0 U13336 ( .IN1(n12171), .IN2(n8561), .QN(n12172) );
  NAND3X0 U13337 ( .IN1(g2319), .IN2(g2351), .IN3(n12193), .QN(n12171) );
  INVX0 U13338 ( .INP(n11099), .ZN(n12193) );
  NAND2X0 U13339 ( .IN1(n3555), .IN2(n12706), .QN(n12704) );
  NAND3X0 U13340 ( .IN1(n12707), .IN2(n12708), .IN3(n12709), .QN(n12706) );
  NAND2X0 U13341 ( .IN1(n456), .IN2(g2295), .QN(n12709) );
  INVX0 U13342 ( .INP(n11114), .ZN(n456) );
  NAND2X0 U13343 ( .IN1(test_so21), .IN2(n5375), .QN(n11114) );
  NAND2X0 U13344 ( .IN1(n5511), .IN2(n12710), .QN(n12708) );
  NAND2X0 U13345 ( .IN1(n12711), .IN2(n12712), .QN(n12710) );
  NAND2X0 U13346 ( .IN1(n5375), .IN2(g2307), .QN(n12712) );
  NAND2X0 U13347 ( .IN1(test_so21), .IN2(g2315), .QN(n12711) );
  NAND2X0 U13348 ( .IN1(n12713), .IN2(n8213), .QN(n12707) );
  NAND2X0 U13349 ( .IN1(n12714), .IN2(n12715), .QN(n12713) );
  NAND2X0 U13350 ( .IN1(g2319), .IN2(n9314), .QN(n12715) );
  NAND2X0 U13351 ( .IN1(g2351), .IN2(g2303), .QN(n12714) );
  NOR2X0 U13352 ( .IN1(n11099), .IN2(n8559), .QN(n3555) );
  NAND2X0 U13353 ( .IN1(n11108), .IN2(g2370), .QN(n12703) );
  INVX0 U13354 ( .INP(n11102), .ZN(n11108) );
  NAND2X0 U13355 ( .IN1(n11099), .IN2(n8524), .QN(n11102) );
  NAND3X0 U13356 ( .IN1(n12674), .IN2(n12088), .IN3(n12716), .QN(n11099) );
  NAND2X0 U13357 ( .IN1(n9579), .IN2(g2807), .QN(n12716) );
  NAND2X0 U13358 ( .IN1(n8586), .IN2(g2351), .QN(n12702) );
  NAND2X0 U13359 ( .IN1(n12717), .IN2(n12718), .QN(g29249) );
  NAND2X0 U13360 ( .IN1(n12719), .IN2(g2250), .QN(n12718) );
  NAND2X0 U13361 ( .IN1(n11123), .IN2(n12720), .QN(n12719) );
  NAND2X0 U13362 ( .IN1(n4414), .IN2(n8524), .QN(n12720) );
  NAND2X0 U13363 ( .IN1(n12721), .IN2(g2236), .QN(n12717) );
  NAND2X0 U13364 ( .IN1(n12722), .IN2(n8524), .QN(n12721) );
  OR2X1 U13365 ( .IN1(n11120), .IN2(n8828), .Q(n12722) );
  NOR2X0 U13366 ( .IN1(n7907), .IN2(n982), .QN(n8828) );
  NAND4X0 U13367 ( .IN1(n12723), .IN2(n12724), .IN3(n12725), .IN4(n12726), 
        .QN(g29248) );
  NAND2X0 U13368 ( .IN1(n12201), .IN2(g2165), .QN(n12726) );
  NOR2X0 U13369 ( .IN1(n12200), .IN2(n8559), .QN(n12201) );
  NAND3X0 U13370 ( .IN1(g2185), .IN2(g2217), .IN3(n12222), .QN(n12200) );
  INVX0 U13371 ( .INP(n11120), .ZN(n12222) );
  NAND2X0 U13372 ( .IN1(n3574), .IN2(n12727), .QN(n12725) );
  NAND3X0 U13373 ( .IN1(n12728), .IN2(n12729), .IN3(n12730), .QN(n12727) );
  NAND2X0 U13374 ( .IN1(n982), .IN2(g2161), .QN(n12730) );
  INVX0 U13375 ( .INP(n11135), .ZN(n982) );
  NAND2X0 U13376 ( .IN1(n5376), .IN2(g2208), .QN(n11135) );
  NAND2X0 U13377 ( .IN1(n5512), .IN2(n12731), .QN(n12729) );
  NAND2X0 U13378 ( .IN1(n12732), .IN2(n12733), .QN(n12731) );
  NAND2X0 U13379 ( .IN1(n5376), .IN2(g2173), .QN(n12733) );
  NAND2X0 U13380 ( .IN1(g2181), .IN2(g2208), .QN(n12732) );
  NAND2X0 U13381 ( .IN1(n8133), .IN2(n12734), .QN(n12728) );
  NAND2X0 U13382 ( .IN1(n12735), .IN2(n12736), .QN(n12734) );
  NAND2X0 U13383 ( .IN1(g2185), .IN2(n9352), .QN(n12736) );
  NAND2X0 U13384 ( .IN1(g2217), .IN2(g2169), .QN(n12735) );
  NOR2X0 U13385 ( .IN1(n11120), .IN2(n8558), .QN(n3574) );
  NAND2X0 U13386 ( .IN1(n11129), .IN2(g2236), .QN(n12724) );
  INVX0 U13387 ( .INP(n11123), .ZN(n11129) );
  NAND2X0 U13388 ( .IN1(n11120), .IN2(n8524), .QN(n11123) );
  NAND3X0 U13389 ( .IN1(n12737), .IN2(n12674), .IN3(n12077), .QN(n11120) );
  NAND2X0 U13390 ( .IN1(n9579), .IN2(g2803), .QN(n12737) );
  NAND2X0 U13391 ( .IN1(n8588), .IN2(g2217), .QN(n12723) );
  NAND2X0 U13392 ( .IN1(n12738), .IN2(n12739), .QN(g29247) );
  NAND2X0 U13393 ( .IN1(n12740), .IN2(g2079), .QN(n12739) );
  NAND2X0 U13394 ( .IN1(n12741), .IN2(n8524), .QN(n12740) );
  NAND2X0 U13395 ( .IN1(n12251), .IN2(n8827), .QN(n12741) );
  NAND2X0 U13396 ( .IN1(test_so78), .IN2(n11156), .QN(n8827) );
  NAND2X0 U13397 ( .IN1(test_so78), .IN2(n12742), .QN(n12738) );
  NAND2X0 U13398 ( .IN1(n11144), .IN2(n12743), .QN(n12742) );
  NAND2X0 U13399 ( .IN1(n4425), .IN2(n8524), .QN(n12743) );
  NAND4X0 U13400 ( .IN1(n12744), .IN2(n12745), .IN3(n12746), .IN4(n12747), 
        .QN(g29246) );
  NAND2X0 U13401 ( .IN1(n12230), .IN2(g2008), .QN(n12747) );
  NOR2X0 U13402 ( .IN1(n12229), .IN2(n8557), .QN(n12230) );
  NAND3X0 U13403 ( .IN1(g2028), .IN2(g2060), .IN3(n12251), .QN(n12229) );
  INVX0 U13404 ( .INP(n11141), .ZN(n12251) );
  NAND2X0 U13405 ( .IN1(n3593), .IN2(n12748), .QN(n12746) );
  NAND3X0 U13406 ( .IN1(n12749), .IN2(n12750), .IN3(n12751), .QN(n12748) );
  NAND2X0 U13407 ( .IN1(n1136), .IN2(g2004), .QN(n12751) );
  INVX0 U13408 ( .INP(n11156), .ZN(n1136) );
  NAND2X0 U13409 ( .IN1(n5371), .IN2(g2051), .QN(n11156) );
  NAND2X0 U13410 ( .IN1(n5507), .IN2(n12752), .QN(n12750) );
  NAND2X0 U13411 ( .IN1(n12753), .IN2(n12754), .QN(n12752) );
  NAND2X0 U13412 ( .IN1(n5371), .IN2(g2016), .QN(n12754) );
  NAND2X0 U13413 ( .IN1(g2024), .IN2(g2051), .QN(n12753) );
  NAND2X0 U13414 ( .IN1(n8129), .IN2(n12755), .QN(n12749) );
  NAND2X0 U13415 ( .IN1(n12756), .IN2(n12757), .QN(n12755) );
  NAND2X0 U13416 ( .IN1(g2028), .IN2(n9312), .QN(n12757) );
  NAND2X0 U13417 ( .IN1(g2060), .IN2(g2012), .QN(n12756) );
  NOR2X0 U13418 ( .IN1(n11141), .IN2(n8549), .QN(n3593) );
  NAND2X0 U13419 ( .IN1(n11150), .IN2(g2079), .QN(n12745) );
  INVX0 U13420 ( .INP(n11144), .ZN(n11150) );
  NAND2X0 U13421 ( .IN1(n11141), .IN2(n8524), .QN(n11144) );
  NAND3X0 U13422 ( .IN1(n12758), .IN2(n12674), .IN3(n12078), .QN(n11141) );
  NAND2X0 U13423 ( .IN1(n9579), .IN2(g2787), .QN(n12758) );
  NAND2X0 U13424 ( .IN1(n8613), .IN2(g2060), .QN(n12744) );
  NAND2X0 U13425 ( .IN1(n12759), .IN2(n12760), .QN(g29245) );
  NAND2X0 U13426 ( .IN1(n12761), .IN2(g1959), .QN(n12760) );
  NAND2X0 U13427 ( .IN1(n11165), .IN2(n12762), .QN(n12761) );
  NAND2X0 U13428 ( .IN1(n4436), .IN2(n8524), .QN(n12762) );
  NAND2X0 U13429 ( .IN1(test_so53), .IN2(n12763), .QN(n12759) );
  NAND2X0 U13430 ( .IN1(n12764), .IN2(n8524), .QN(n12763) );
  OR2X1 U13431 ( .IN1(n11162), .IN2(n8826), .Q(n12764) );
  NOR2X0 U13432 ( .IN1(n7916), .IN2(n314), .QN(n8826) );
  NAND4X0 U13433 ( .IN1(n12765), .IN2(n12766), .IN3(n12767), .IN4(n12768), 
        .QN(g29244) );
  NAND2X0 U13434 ( .IN1(n12259), .IN2(g1874), .QN(n12768) );
  NOR2X0 U13435 ( .IN1(n12258), .IN2(n8556), .QN(n12259) );
  NAND3X0 U13436 ( .IN1(g1894), .IN2(g1926), .IN3(n12280), .QN(n12258) );
  INVX0 U13437 ( .INP(n11162), .ZN(n12280) );
  NAND2X0 U13438 ( .IN1(n3611), .IN2(n12769), .QN(n12767) );
  NAND3X0 U13439 ( .IN1(n12770), .IN2(n12771), .IN3(n12772), .QN(n12769) );
  NAND2X0 U13440 ( .IN1(n314), .IN2(g1870), .QN(n12772) );
  INVX0 U13441 ( .INP(n11177), .ZN(n314) );
  NAND2X0 U13442 ( .IN1(n5374), .IN2(g1917), .QN(n11177) );
  NAND2X0 U13443 ( .IN1(n5510), .IN2(n12773), .QN(n12771) );
  NAND2X0 U13444 ( .IN1(n12774), .IN2(n12775), .QN(n12773) );
  NAND2X0 U13445 ( .IN1(n5374), .IN2(g1882), .QN(n12775) );
  NAND2X0 U13446 ( .IN1(g1890), .IN2(g1917), .QN(n12774) );
  NAND2X0 U13447 ( .IN1(n8132), .IN2(n12776), .QN(n12770) );
  NAND2X0 U13448 ( .IN1(n12777), .IN2(n12778), .QN(n12776) );
  NAND2X0 U13449 ( .IN1(g1894), .IN2(n9280), .QN(n12778) );
  NAND2X0 U13450 ( .IN1(g1926), .IN2(g1878), .QN(n12777) );
  NOR2X0 U13451 ( .IN1(n11162), .IN2(n8556), .QN(n3611) );
  NAND2X0 U13452 ( .IN1(n11171), .IN2(test_so53), .QN(n12766) );
  INVX0 U13453 ( .INP(n11165), .ZN(n11171) );
  NAND2X0 U13454 ( .IN1(n11162), .IN2(n8524), .QN(n11165) );
  NAND3X0 U13455 ( .IN1(n12779), .IN2(n12674), .IN3(n12087), .QN(n11162) );
  INVX0 U13456 ( .INP(n12076), .ZN(n12087) );
  NAND2X0 U13457 ( .IN1(n9579), .IN2(g2783), .QN(n12779) );
  NAND2X0 U13458 ( .IN1(n8613), .IN2(g1926), .QN(n12765) );
  NAND2X0 U13459 ( .IN1(n12780), .IN2(n12781), .QN(g29243) );
  NAND2X0 U13460 ( .IN1(n12782), .IN2(g1825), .QN(n12781) );
  NAND2X0 U13461 ( .IN1(n11186), .IN2(n12783), .QN(n12782) );
  NAND2X0 U13462 ( .IN1(n4447), .IN2(n8524), .QN(n12783) );
  NAND2X0 U13463 ( .IN1(n12784), .IN2(g1811), .QN(n12780) );
  NAND2X0 U13464 ( .IN1(n12785), .IN2(n8524), .QN(n12784) );
  OR2X1 U13465 ( .IN1(n11183), .IN2(n8825), .Q(n12785) );
  NOR2X0 U13466 ( .IN1(n7909), .IN2(n709), .QN(n8825) );
  NAND4X0 U13467 ( .IN1(n12786), .IN2(n12787), .IN3(n12788), .IN4(n12789), 
        .QN(g29242) );
  NAND2X0 U13468 ( .IN1(n12288), .IN2(g1740), .QN(n12789) );
  NOR2X0 U13469 ( .IN1(n12287), .IN2(n8555), .QN(n12288) );
  NAND3X0 U13470 ( .IN1(g1792), .IN2(g1760), .IN3(n12309), .QN(n12287) );
  INVX0 U13471 ( .INP(n11183), .ZN(n12309) );
  NAND2X0 U13472 ( .IN1(n3628), .IN2(n12790), .QN(n12788) );
  NAND3X0 U13473 ( .IN1(n12791), .IN2(n12792), .IN3(n12793), .QN(n12790) );
  NAND2X0 U13474 ( .IN1(n709), .IN2(g1736), .QN(n12793) );
  INVX0 U13475 ( .INP(n11198), .ZN(n709) );
  NAND2X0 U13476 ( .IN1(n5602), .IN2(g1783), .QN(n11198) );
  NAND2X0 U13477 ( .IN1(n5359), .IN2(n12794), .QN(n12792) );
  NAND2X0 U13478 ( .IN1(n12795), .IN2(n12796), .QN(n12794) );
  NAND2X0 U13479 ( .IN1(g1783), .IN2(g1756), .QN(n12796) );
  NAND2X0 U13480 ( .IN1(n5602), .IN2(g1748), .QN(n12795) );
  NAND2X0 U13481 ( .IN1(n5596), .IN2(n12797), .QN(n12791) );
  NAND2X0 U13482 ( .IN1(n12798), .IN2(n12799), .QN(n12797) );
  NAND2X0 U13483 ( .IN1(g1792), .IN2(g1744), .QN(n12799) );
  NAND2X0 U13484 ( .IN1(g1760), .IN2(g1752), .QN(n12798) );
  NOR2X0 U13485 ( .IN1(n11183), .IN2(n8555), .QN(n3628) );
  NAND2X0 U13486 ( .IN1(n11192), .IN2(g1811), .QN(n12787) );
  INVX0 U13487 ( .INP(n11186), .ZN(n11192) );
  NAND2X0 U13488 ( .IN1(n11183), .IN2(n8524), .QN(n11186) );
  NAND3X0 U13489 ( .IN1(n12674), .IN2(n12088), .IN3(n12800), .QN(n11183) );
  NAND2X0 U13490 ( .IN1(n9579), .IN2(g2775), .QN(n12800) );
  INVX0 U13491 ( .INP(n4411), .ZN(n12088) );
  NAND2X0 U13492 ( .IN1(n5465), .IN2(g2715), .QN(n4411) );
  NAND2X0 U13493 ( .IN1(n8612), .IN2(g1792), .QN(n12786) );
  NAND2X0 U13494 ( .IN1(n12801), .IN2(n12802), .QN(g29241) );
  NAND2X0 U13495 ( .IN1(n12803), .IN2(g1691), .QN(n12802) );
  NAND2X0 U13496 ( .IN1(n11207), .IN2(n12804), .QN(n12803) );
  NAND2X0 U13497 ( .IN1(n4458), .IN2(n8524), .QN(n12804) );
  NAND2X0 U13498 ( .IN1(n12805), .IN2(g1677), .QN(n12801) );
  NAND2X0 U13499 ( .IN1(n12806), .IN2(n8524), .QN(n12805) );
  OR2X1 U13500 ( .IN1(n11204), .IN2(n8824), .Q(n12806) );
  NOR2X0 U13501 ( .IN1(n7913), .IN2(n1123), .QN(n8824) );
  NAND4X0 U13502 ( .IN1(n12807), .IN2(n12808), .IN3(n12809), .IN4(n12810), 
        .QN(g29240) );
  NAND2X0 U13503 ( .IN1(n3646), .IN2(n12811), .QN(n12810) );
  NAND4X0 U13504 ( .IN1(n12812), .IN2(n12813), .IN3(n12814), .IN4(n12815), 
        .QN(n12811) );
  NAND3X0 U13505 ( .IN1(n5370), .IN2(g1612), .IN3(n5525), .QN(n12815) );
  NAND2X0 U13506 ( .IN1(n12816), .IN2(n8210), .QN(n12814) );
  NAND2X0 U13507 ( .IN1(n12817), .IN2(n12818), .QN(n12816) );
  NAND2X0 U13508 ( .IN1(g1624), .IN2(n9303), .QN(n12818) );
  NAND2X0 U13509 ( .IN1(g1657), .IN2(g1608), .QN(n12817) );
  NAND2X0 U13510 ( .IN1(n1123), .IN2(g1600), .QN(n12813) );
  INVX0 U13511 ( .INP(n11221), .ZN(n1123) );
  NAND2X0 U13512 ( .IN1(test_so94), .IN2(n5370), .QN(n11221) );
  NAND2X0 U13513 ( .IN1(g31863), .IN2(g1620), .QN(n12812) );
  NOR2X0 U13514 ( .IN1(g1657), .IN2(n8210), .QN(g31863) );
  NOR2X0 U13515 ( .IN1(n11204), .IN2(n8555), .QN(n3646) );
  NAND2X0 U13516 ( .IN1(n12316), .IN2(g1604), .QN(n12809) );
  NOR3X0 U13517 ( .IN1(n5370), .IN2(n5525), .IN3(n11204), .QN(n12316) );
  NAND2X0 U13518 ( .IN1(n11215), .IN2(g1677), .QN(n12808) );
  INVX0 U13519 ( .INP(n11207), .ZN(n11215) );
  NAND2X0 U13520 ( .IN1(n11204), .IN2(n8524), .QN(n11207) );
  NAND3X0 U13521 ( .IN1(n12819), .IN2(n12674), .IN3(n12077), .QN(n11204) );
  INVX0 U13522 ( .INP(n12086), .ZN(n12077) );
  NAND2X0 U13523 ( .IN1(n5299), .IN2(n5465), .QN(n12086) );
  NAND2X0 U13524 ( .IN1(n12820), .IN2(n9579), .QN(n12674) );
  INVX0 U13525 ( .INP(n4388), .ZN(n12820) );
  NAND2X0 U13526 ( .IN1(n9579), .IN2(g2771), .QN(n12819) );
  NOR2X0 U13527 ( .IN1(g2729), .IN2(g2724), .QN(n9579) );
  NAND2X0 U13528 ( .IN1(n8612), .IN2(g1657), .QN(n12807) );
  NAND3X0 U13529 ( .IN1(n12821), .IN2(n12822), .IN3(n12823), .QN(g29239) );
  NAND3X0 U13530 ( .IN1(n12824), .IN2(n10598), .IN3(n12825), .QN(n12823) );
  NAND2X0 U13531 ( .IN1(n8612), .IN2(g1478), .QN(n12822) );
  NAND3X0 U13532 ( .IN1(n12826), .IN2(g1454), .IN3(n8494), .QN(n12821) );
  NAND2X0 U13533 ( .IN1(n12827), .IN2(n12828), .QN(n12826) );
  INVX0 U13534 ( .INP(n12824), .ZN(n12828) );
  XOR2X1 U13535 ( .IN1(g1448), .IN2(n12829), .Q(n12824) );
  NAND3X0 U13536 ( .IN1(n12830), .IN2(n12831), .IN3(n12832), .QN(g29238) );
  NAND2X0 U13537 ( .IN1(n12833), .IN2(g1484), .QN(n12832) );
  NAND2X0 U13538 ( .IN1(n8612), .IN2(g1472), .QN(n12831) );
  NAND3X0 U13539 ( .IN1(n12834), .IN2(n12835), .IN3(n8494), .QN(n12830) );
  NAND2X0 U13540 ( .IN1(n5865), .IN2(n12836), .QN(n12835) );
  NAND3X0 U13541 ( .IN1(n8137), .IN2(n5850), .IN3(n12837), .QN(n12836) );
  XOR2X1 U13542 ( .IN1(g1300), .IN2(n12829), .Q(n12834) );
  NAND3X0 U13543 ( .IN1(n12838), .IN2(n12839), .IN3(n12840), .QN(g29237) );
  NAND3X0 U13544 ( .IN1(n12825), .IN2(n10561), .IN3(n12841), .QN(n12840) );
  NAND2X0 U13545 ( .IN1(n8612), .IN2(g1448), .QN(n12839) );
  NAND3X0 U13546 ( .IN1(n12842), .IN2(g1467), .IN3(n8494), .QN(n12838) );
  NAND3X0 U13547 ( .IN1(n12843), .IN2(g13272), .IN3(n10561), .QN(n12842) );
  INVX0 U13548 ( .INP(n12841), .ZN(n12843) );
  XOR2X1 U13549 ( .IN1(g1472), .IN2(n12829), .Q(n12841) );
  NAND3X0 U13550 ( .IN1(n12844), .IN2(n12845), .IN3(n12846), .QN(g29236) );
  NAND3X0 U13551 ( .IN1(n12825), .IN2(n10636), .IN3(n12847), .QN(n12846) );
  NOR4X0 U13552 ( .IN1(g1442), .IN2(g1489), .IN3(n8545), .IN4(n7832), .QN(
        n12825) );
  NAND2X0 U13553 ( .IN1(n8611), .IN2(g1442), .QN(n12845) );
  NAND3X0 U13554 ( .IN1(n12848), .IN2(g1437), .IN3(n8494), .QN(n12844) );
  NAND3X0 U13555 ( .IN1(n12849), .IN2(g13272), .IN3(n10636), .QN(n12848) );
  INVX0 U13556 ( .INP(n12847), .ZN(n12849) );
  XOR2X1 U13557 ( .IN1(g1478), .IN2(n12829), .Q(n12847) );
  AND2X1 U13558 ( .IN1(n9225), .IN2(DFF_1092_n1), .Q(n12829) );
  INVX0 U13559 ( .INP(n9311), .ZN(n9225) );
  NAND3X0 U13560 ( .IN1(n12850), .IN2(n12851), .IN3(n12852), .QN(g29235) );
  OR2X1 U13561 ( .IN1(n8480), .IN2(n5554), .Q(n12852) );
  OR3X1 U13562 ( .IN1(n10807), .IN2(n4178), .IN3(n5558), .Q(n12851) );
  NAND2X0 U13563 ( .IN1(n4178), .IN2(n5558), .QN(n12850) );
  NAND3X0 U13564 ( .IN1(n12853), .IN2(n12854), .IN3(n12855), .QN(g29234) );
  NAND3X0 U13565 ( .IN1(n12856), .IN2(n10756), .IN3(n12857), .QN(n12855) );
  NAND2X0 U13566 ( .IN1(n8611), .IN2(g1135), .QN(n12854) );
  NAND3X0 U13567 ( .IN1(test_so90), .IN2(n12858), .IN3(n8494), .QN(n12853) );
  NAND2X0 U13568 ( .IN1(n12859), .IN2(n12860), .QN(n12858) );
  INVX0 U13569 ( .INP(n12856), .ZN(n12860) );
  XOR2X1 U13570 ( .IN1(n12861), .IN2(n5478), .Q(n12856) );
  NAND3X0 U13571 ( .IN1(n12862), .IN2(n12863), .IN3(n12864), .QN(g29233) );
  NAND2X0 U13572 ( .IN1(n12865), .IN2(g1141), .QN(n12864) );
  NAND2X0 U13573 ( .IN1(n8611), .IN2(g1129), .QN(n12863) );
  NAND3X0 U13574 ( .IN1(n12866), .IN2(n12867), .IN3(n8494), .QN(n12862) );
  NAND2X0 U13575 ( .IN1(n5691), .IN2(n12868), .QN(n12867) );
  NAND3X0 U13576 ( .IN1(n5851), .IN2(n8207), .IN3(n12869), .QN(n12868) );
  XOR2X1 U13577 ( .IN1(n12861), .IN2(n5341), .Q(n12866) );
  NAND3X0 U13578 ( .IN1(n12870), .IN2(n12871), .IN3(n12872), .QN(g29232) );
  NAND3X0 U13579 ( .IN1(n12857), .IN2(n10718), .IN3(n12873), .QN(n12872) );
  NAND2X0 U13580 ( .IN1(n8611), .IN2(g1105), .QN(n12871) );
  NAND3X0 U13581 ( .IN1(n12874), .IN2(g1124), .IN3(n8493), .QN(n12870) );
  NAND3X0 U13582 ( .IN1(n12875), .IN2(g13259), .IN3(n10718), .QN(n12874) );
  INVX0 U13583 ( .INP(n12873), .ZN(n12875) );
  XOR2X1 U13584 ( .IN1(n12861), .IN2(n5329), .Q(n12873) );
  NAND3X0 U13585 ( .IN1(n12876), .IN2(n12877), .IN3(n12878), .QN(g29231) );
  NAND3X0 U13586 ( .IN1(n12857), .IN2(n10841), .IN3(n12879), .QN(n12878) );
  NOR4X0 U13587 ( .IN1(g1146), .IN2(n8544), .IN3(n7831), .IN4(test_so7), .QN(
        n12857) );
  NAND2X0 U13588 ( .IN1(test_so7), .IN2(n8549), .QN(n12877) );
  NAND3X0 U13589 ( .IN1(n12880), .IN2(g1094), .IN3(n8493), .QN(n12876) );
  NAND3X0 U13590 ( .IN1(n12881), .IN2(g13259), .IN3(n10841), .QN(n12880) );
  INVX0 U13591 ( .INP(n12879), .ZN(n12881) );
  XOR2X1 U13592 ( .IN1(n12861), .IN2(n5328), .Q(n12879) );
  NAND2X0 U13593 ( .IN1(n9224), .IN2(DFF_24_n1), .QN(n12861) );
  INVX0 U13594 ( .INP(n11245), .ZN(n9224) );
  NAND3X0 U13595 ( .IN1(n12882), .IN2(n12883), .IN3(n12884), .QN(g29230) );
  OR2X1 U13596 ( .IN1(n8480), .IN2(n5555), .Q(n12884) );
  OR3X1 U13597 ( .IN1(n10820), .IN2(n4196), .IN3(n5559), .Q(n12883) );
  NAND2X0 U13598 ( .IN1(n4196), .IN2(n5559), .QN(n12882) );
  NAND3X0 U13599 ( .IN1(n12885), .IN2(n12886), .IN3(n12887), .QN(g29229) );
  NAND2X0 U13600 ( .IN1(n8610), .IN2(g827), .QN(n12887) );
  NAND2X0 U13601 ( .IN1(n4517), .IN2(g723), .QN(n12886) );
  NAND3X0 U13602 ( .IN1(n4516), .IN2(n12888), .IN3(n5826), .QN(n12885) );
  NAND2X0 U13603 ( .IN1(n12889), .IN2(n12890), .QN(g29228) );
  NAND2X0 U13604 ( .IN1(n2404), .IN2(n12891), .QN(n12890) );
  XOR2X1 U13605 ( .IN1(test_so60), .IN2(n12400), .Q(n12891) );
  NOR2X0 U13606 ( .IN1(n12408), .IN2(n12892), .QN(n12400) );
  AND2X1 U13607 ( .IN1(n5482), .IN2(g12184), .Q(n12892) );
  NAND2X0 U13608 ( .IN1(n8610), .IN2(g736), .QN(n12889) );
  NAND3X0 U13609 ( .IN1(n12893), .IN2(n12894), .IN3(n12895), .QN(g29227) );
  NAND2X0 U13610 ( .IN1(n8610), .IN2(g676), .QN(n12895) );
  NAND3X0 U13611 ( .IN1(n4523), .IN2(n12896), .IN3(n8225), .QN(n12894) );
  NAND2X0 U13612 ( .IN1(n4524), .IN2(test_so70), .QN(n12893) );
  NAND3X0 U13613 ( .IN1(n12897), .IN2(n12898), .IN3(n12899), .QN(g29226) );
  OR2X1 U13614 ( .IN1(n8480), .IN2(n7718), .Q(n12899) );
  NAND3X0 U13615 ( .IN1(n4525), .IN2(n12900), .IN3(g676), .QN(n12898) );
  INVX0 U13616 ( .INP(n4526), .ZN(n12900) );
  NAND3X0 U13617 ( .IN1(n4526), .IN2(n12896), .IN3(n5751), .QN(n12897) );
  NAND2X0 U13618 ( .IN1(n12901), .IN2(n12902), .QN(g29225) );
  NAND2X0 U13619 ( .IN1(n12903), .IN2(n4525), .QN(n12902) );
  AND2X1 U13620 ( .IN1(n12896), .IN2(n8508), .Q(n4525) );
  AND2X1 U13621 ( .IN1(n12904), .IN2(g703), .Q(n12896) );
  NAND4X0 U13622 ( .IN1(n12905), .IN2(n12906), .IN3(n12907), .IN4(g681), .QN(
        n12904) );
  INVX0 U13623 ( .INP(n4535), .ZN(n12905) );
  XNOR2X1 U13624 ( .IN1(g718), .IN2(n7906), .Q(n4535) );
  XOR2X1 U13625 ( .IN1(n8195), .IN2(n7718), .Q(n12903) );
  NAND2X0 U13626 ( .IN1(n8610), .IN2(g667), .QN(n12901) );
  NAND3X0 U13627 ( .IN1(n12908), .IN2(n12909), .IN3(n12910), .QN(g29224) );
  NAND2X0 U13628 ( .IN1(n8610), .IN2(g572), .QN(n12910) );
  NAND3X0 U13629 ( .IN1(n2421), .IN2(n12911), .IN3(g586), .QN(n12909) );
  INVX0 U13630 ( .INP(n4201), .ZN(n12911) );
  NAND2X0 U13631 ( .IN1(n4201), .IN2(n5336), .QN(n12908) );
  NAND3X0 U13632 ( .IN1(n12912), .IN2(n12913), .IN3(n12914), .QN(g29223) );
  NAND2X0 U13633 ( .IN1(n12915), .IN2(n5708), .QN(n12914) );
  NAND2X0 U13634 ( .IN1(n8609), .IN2(g482), .QN(n12913) );
  NAND2X0 U13635 ( .IN1(n12916), .IN2(n8524), .QN(n12912) );
  NAND2X0 U13636 ( .IN1(n12917), .IN2(n12918), .QN(n12916) );
  OR2X1 U13637 ( .IN1(n12915), .IN2(n5708), .Q(n12918) );
  NOR2X0 U13638 ( .IN1(n12919), .IN2(n5820), .QN(n12915) );
  NAND3X0 U13639 ( .IN1(n12920), .IN2(n12921), .IN3(n12922), .QN(g29222) );
  NAND2X0 U13640 ( .IN1(n12923), .IN2(g411), .QN(n12922) );
  NAND2X0 U13641 ( .IN1(n12924), .IN2(g417), .QN(n12921) );
  NAND2X0 U13642 ( .IN1(n12925), .IN2(n8523), .QN(n12924) );
  OR2X1 U13643 ( .IN1(n12926), .IN2(n3676), .Q(n12925) );
  NAND3X0 U13644 ( .IN1(n12927), .IN2(n3676), .IN3(n5358), .QN(n12920) );
  XOR2X1 U13645 ( .IN1(g417), .IN2(n12928), .Q(n3676) );
  NOR2X0 U13646 ( .IN1(n12929), .IN2(n12930), .QN(n12928) );
  NOR2X0 U13647 ( .IN1(g392), .IN2(n12931), .QN(n12930) );
  NOR2X0 U13648 ( .IN1(n12932), .IN2(n12933), .QN(n12931) );
  NOR2X0 U13649 ( .IN1(n7833), .IN2(g405), .QN(n12933) );
  NOR2X0 U13650 ( .IN1(n7835), .IN2(n7834), .QN(n12932) );
  NOR2X0 U13651 ( .IN1(n7865), .IN2(n12934), .QN(n12929) );
  NOR2X0 U13652 ( .IN1(n12935), .IN2(n12936), .QN(n12934) );
  NOR2X0 U13653 ( .IN1(n7835), .IN2(n7813), .QN(n12936) );
  NOR2X0 U13654 ( .IN1(n7834), .IN2(g405), .QN(n12935) );
  NAND3X0 U13655 ( .IN1(n12937), .IN2(n12938), .IN3(n12939), .QN(g28105) );
  NAND2X0 U13656 ( .IN1(n10372), .IN2(g5011), .QN(n12939) );
  NAND2X0 U13657 ( .IN1(n8609), .IN2(g6657), .QN(n12938) );
  NAND3X0 U13658 ( .IN1(n12440), .IN2(n10365), .IN3(n8493), .QN(n12937) );
  NAND2X0 U13659 ( .IN1(n12940), .IN2(n12941), .QN(n12440) );
  NAND2X0 U13660 ( .IN1(n5531), .IN2(n12942), .QN(n12941) );
  NAND4X0 U13661 ( .IN1(n12943), .IN2(n12944), .IN3(n12945), .IN4(n12946), 
        .QN(n12942) );
  AND3X1 U13662 ( .IN1(n12947), .IN2(n12948), .IN3(n12949), .Q(n12946) );
  NAND2X0 U13663 ( .IN1(n8819), .IN2(n12950), .QN(n12949) );
  NAND2X0 U13664 ( .IN1(n12951), .IN2(n12952), .QN(n12950) );
  NAND2X0 U13665 ( .IN1(g6723), .IN2(g6605), .QN(n12952) );
  NAND2X0 U13666 ( .IN1(g13099), .IN2(g6593), .QN(n12951) );
  NAND3X0 U13667 ( .IN1(g14749), .IN2(g6633), .IN3(n8820), .QN(n12948) );
  NAND3X0 U13668 ( .IN1(g17871), .IN2(g6617), .IN3(n8821), .QN(n12947) );
  NAND2X0 U13669 ( .IN1(n8822), .IN2(n12953), .QN(n12945) );
  NAND2X0 U13670 ( .IN1(n12954), .IN2(n12955), .QN(n12953) );
  NAND2X0 U13671 ( .IN1(g17764), .IN2(g6649), .QN(n12955) );
  NAND2X0 U13672 ( .IN1(g17722), .IN2(g6597), .QN(n12954) );
  NAND2X0 U13673 ( .IN1(n12956), .IN2(n8231), .QN(n12944) );
  NAND2X0 U13674 ( .IN1(test_so80), .IN2(n12957), .QN(n12943) );
  NAND2X0 U13675 ( .IN1(n12958), .IN2(n12959), .QN(n12957) );
  NAND2X0 U13676 ( .IN1(n8821), .IN2(g6601), .QN(n12959) );
  INVX0 U13677 ( .INP(n12960), .ZN(n12958) );
  NAND2X0 U13678 ( .IN1(n12961), .IN2(g6727), .QN(n12940) );
  NAND4X0 U13679 ( .IN1(n12962), .IN2(n12963), .IN3(n12964), .IN4(n12965), 
        .QN(n12961) );
  AND3X1 U13680 ( .IN1(n12966), .IN2(n12967), .IN3(n12968), .Q(n12965) );
  NAND2X0 U13681 ( .IN1(n8820), .IN2(n12969), .QN(n12968) );
  NAND2X0 U13682 ( .IN1(n12970), .IN2(n12971), .QN(n12969) );
  NAND2X0 U13683 ( .IN1(g6589), .IN2(g6723), .QN(n12971) );
  NAND2X0 U13684 ( .IN1(g6581), .IN2(g13099), .QN(n12970) );
  NAND3X0 U13685 ( .IN1(g14749), .IN2(g6625), .IN3(n8819), .QN(n12967) );
  NAND3X0 U13686 ( .IN1(g6609), .IN2(g17871), .IN3(n8822), .QN(n12966) );
  NAND2X0 U13687 ( .IN1(n8821), .IN2(n12972), .QN(n12964) );
  NAND2X0 U13688 ( .IN1(n12973), .IN2(n12974), .QN(n12972) );
  NAND2X0 U13689 ( .IN1(g6657), .IN2(g17722), .QN(n12974) );
  NAND2X0 U13690 ( .IN1(g6641), .IN2(g17764), .QN(n12973) );
  NAND2X0 U13691 ( .IN1(n12960), .IN2(n8231), .QN(n12963) );
  NAND3X0 U13692 ( .IN1(n12975), .IN2(n12976), .IN3(n12977), .QN(n12960) );
  NAND3X0 U13693 ( .IN1(g6637), .IN2(g17778), .IN3(n8822), .QN(n12977) );
  NAND3X0 U13694 ( .IN1(g14828), .IN2(g6621), .IN3(n8820), .QN(n12976) );
  NAND3X0 U13695 ( .IN1(g6653), .IN2(g17688), .IN3(n8819), .QN(n12975) );
  NAND2X0 U13696 ( .IN1(test_so80), .IN2(n12978), .QN(n12962) );
  NAND2X0 U13697 ( .IN1(n12979), .IN2(n12980), .QN(n12978) );
  NAND2X0 U13698 ( .IN1(test_so71), .IN2(n8822), .QN(n12980) );
  NOR2X0 U13699 ( .IN1(g6682), .IN2(n5398), .QN(n8822) );
  INVX0 U13700 ( .INP(n12956), .ZN(n12979) );
  NAND3X0 U13701 ( .IN1(n12981), .IN2(n12982), .IN3(n12983), .QN(n12956) );
  NAND3X0 U13702 ( .IN1(g14828), .IN2(g6613), .IN3(n8819), .QN(n12983) );
  NOR2X0 U13703 ( .IN1(g6741), .IN2(n5590), .QN(n8819) );
  NAND3X0 U13704 ( .IN1(g17688), .IN2(g6645), .IN3(n8820), .QN(n12982) );
  NOR2X0 U13705 ( .IN1(g6682), .IN2(g6741), .QN(n8820) );
  NAND3X0 U13706 ( .IN1(g17778), .IN2(g6629), .IN3(n8821), .QN(n12981) );
  NOR2X0 U13707 ( .IN1(n5398), .IN2(n5590), .QN(n8821) );
  NAND3X0 U13708 ( .IN1(n12984), .IN2(n12985), .IN3(n12986), .QN(g28102) );
  NAND2X0 U13709 ( .IN1(n10387), .IN2(g4826), .QN(n12986) );
  NAND2X0 U13710 ( .IN1(n8609), .IN2(g6311), .QN(n12985) );
  NAND3X0 U13711 ( .IN1(n10377), .IN2(n12468), .IN3(n8493), .QN(n12984) );
  NAND2X0 U13712 ( .IN1(n12987), .IN2(n12988), .QN(n12468) );
  NAND2X0 U13713 ( .IN1(test_so69), .IN2(n12989), .QN(n12988) );
  NAND4X0 U13714 ( .IN1(n12990), .IN2(n12991), .IN3(n12992), .IN4(n12993), 
        .QN(n12989) );
  AND3X1 U13715 ( .IN1(n12994), .IN2(n12995), .IN3(n12996), .Q(n12993) );
  NAND2X0 U13716 ( .IN1(n12997), .IN2(n12998), .QN(n12996) );
  NAND2X0 U13717 ( .IN1(n12999), .IN2(n13000), .QN(n12998) );
  NAND2X0 U13718 ( .IN1(g6243), .IN2(g6377), .QN(n13000) );
  NAND2X0 U13719 ( .IN1(g6235), .IN2(g13085), .QN(n12999) );
  NAND3X0 U13720 ( .IN1(g6263), .IN2(g17845), .IN3(n10379), .QN(n12995) );
  NAND3X0 U13721 ( .IN1(g14705), .IN2(g6279), .IN3(n10383), .QN(n12994) );
  NAND2X0 U13722 ( .IN1(n9612), .IN2(n13001), .QN(n12992) );
  NAND2X0 U13723 ( .IN1(n13002), .IN2(n13003), .QN(n13001) );
  NAND2X0 U13724 ( .IN1(g6311), .IN2(g17685), .QN(n13003) );
  NAND2X0 U13725 ( .IN1(g6295), .IN2(g17743), .QN(n13002) );
  NAND2X0 U13726 ( .IN1(n5437), .IN2(n13004), .QN(n12991) );
  NAND2X0 U13727 ( .IN1(n13005), .IN2(g12422), .QN(n12990) );
  NAND2X0 U13728 ( .IN1(n13006), .IN2(n13007), .QN(n13005) );
  NAND2X0 U13729 ( .IN1(n10379), .IN2(g6239), .QN(n13007) );
  INVX0 U13730 ( .INP(n13008), .ZN(n13006) );
  NAND2X0 U13731 ( .IN1(n13009), .IN2(n8237), .QN(n12987) );
  NAND4X0 U13732 ( .IN1(n13010), .IN2(n13011), .IN3(n13012), .IN4(n13013), 
        .QN(n13009) );
  AND3X1 U13733 ( .IN1(n13014), .IN2(n13015), .IN3(n13016), .Q(n13013) );
  NAND2X0 U13734 ( .IN1(n10379), .IN2(n13017), .QN(n13016) );
  NAND2X0 U13735 ( .IN1(n13018), .IN2(n13019), .QN(n13017) );
  NAND2X0 U13736 ( .IN1(g17743), .IN2(g6303), .QN(n13019) );
  NAND2X0 U13737 ( .IN1(g17685), .IN2(g6251), .QN(n13018) );
  NAND3X0 U13738 ( .IN1(g14705), .IN2(g6287), .IN3(n12997), .QN(n13015) );
  NAND3X0 U13739 ( .IN1(g17845), .IN2(g6271), .IN3(n9612), .QN(n13014) );
  NAND2X0 U13740 ( .IN1(n10383), .IN2(n13020), .QN(n13012) );
  NAND2X0 U13741 ( .IN1(n13021), .IN2(n13022), .QN(n13020) );
  NAND2X0 U13742 ( .IN1(g6377), .IN2(g6259), .QN(n13022) );
  NAND2X0 U13743 ( .IN1(g13085), .IN2(g6247), .QN(n13021) );
  NAND2X0 U13744 ( .IN1(n5437), .IN2(n13008), .QN(n13011) );
  NAND3X0 U13745 ( .IN1(n13023), .IN2(n13024), .IN3(n13025), .QN(n13008) );
  NAND3X0 U13746 ( .IN1(g17760), .IN2(g6283), .IN3(n9612), .QN(n13025) );
  NAND3X0 U13747 ( .IN1(g17649), .IN2(g6299), .IN3(n12997), .QN(n13024) );
  NAND3X0 U13748 ( .IN1(g14779), .IN2(g6267), .IN3(n10383), .QN(n13023) );
  NAND2X0 U13749 ( .IN1(n13026), .IN2(g12422), .QN(n13010) );
  NAND2X0 U13750 ( .IN1(n13027), .IN2(n13028), .QN(n13026) );
  NAND2X0 U13751 ( .IN1(n9612), .IN2(g6255), .QN(n13028) );
  INVX0 U13752 ( .INP(n13004), .ZN(n13027) );
  NAND3X0 U13753 ( .IN1(n13029), .IN2(n13030), .IN3(n13031), .QN(n13004) );
  NAND3X0 U13754 ( .IN1(g6307), .IN2(g17649), .IN3(n10383), .QN(n13031) );
  NAND3X0 U13755 ( .IN1(g6291), .IN2(g17760), .IN3(n10379), .QN(n13030) );
  NAND3X0 U13756 ( .IN1(g14779), .IN2(g6275), .IN3(n12997), .QN(n13029) );
  NAND3X0 U13757 ( .IN1(n13032), .IN2(n13033), .IN3(n13034), .QN(g28099) );
  NAND2X0 U13758 ( .IN1(n10402), .IN2(g4831), .QN(n13034) );
  NAND2X0 U13759 ( .IN1(test_so13), .IN2(n8558), .QN(n13033) );
  NAND3X0 U13760 ( .IN1(n10392), .IN2(n12497), .IN3(n8493), .QN(n13032) );
  NAND2X0 U13761 ( .IN1(n13035), .IN2(n13036), .QN(n12497) );
  NAND2X0 U13762 ( .IN1(n5528), .IN2(n13037), .QN(n13036) );
  NAND4X0 U13763 ( .IN1(n13038), .IN2(n13039), .IN3(n13040), .IN4(n13041), 
        .QN(n13037) );
  AND3X1 U13764 ( .IN1(n13042), .IN2(n13043), .IN3(n13044), .Q(n13041) );
  NAND2X0 U13765 ( .IN1(n10394), .IN2(n13045), .QN(n13044) );
  NAND2X0 U13766 ( .IN1(n13046), .IN2(n13047), .QN(n13045) );
  NAND2X0 U13767 ( .IN1(g17715), .IN2(g5957), .QN(n13047) );
  NAND2X0 U13768 ( .IN1(g17646), .IN2(g5905), .QN(n13046) );
  NAND3X0 U13769 ( .IN1(g14673), .IN2(g5941), .IN3(n13048), .QN(n13043) );
  NAND3X0 U13770 ( .IN1(g17819), .IN2(g5925), .IN3(n9617), .QN(n13042) );
  NAND2X0 U13771 ( .IN1(n10398), .IN2(n13049), .QN(n13040) );
  NAND2X0 U13772 ( .IN1(n13050), .IN2(n13051), .QN(n13049) );
  NAND2X0 U13773 ( .IN1(g6031), .IN2(g5913), .QN(n13051) );
  NAND2X0 U13774 ( .IN1(g13068), .IN2(g5901), .QN(n13050) );
  NAND2X0 U13775 ( .IN1(n5432), .IN2(n13052), .QN(n13039) );
  NAND2X0 U13776 ( .IN1(n13053), .IN2(g12350), .QN(n13038) );
  NAND2X0 U13777 ( .IN1(n13054), .IN2(n13055), .QN(n13053) );
  NAND2X0 U13778 ( .IN1(n9617), .IN2(g5909), .QN(n13055) );
  INVX0 U13779 ( .INP(n13056), .ZN(n13054) );
  NAND2X0 U13780 ( .IN1(n13057), .IN2(g6035), .QN(n13035) );
  NAND4X0 U13781 ( .IN1(n13058), .IN2(n13059), .IN3(n13060), .IN4(n13061), 
        .QN(n13057) );
  AND3X1 U13782 ( .IN1(n13062), .IN2(n13063), .IN3(n13064), .Q(n13061) );
  NAND2X0 U13783 ( .IN1(n13048), .IN2(n13065), .QN(n13064) );
  NAND2X0 U13784 ( .IN1(n13066), .IN2(n13067), .QN(n13065) );
  NAND2X0 U13785 ( .IN1(g5897), .IN2(g6031), .QN(n13067) );
  NAND2X0 U13786 ( .IN1(g5889), .IN2(g13068), .QN(n13066) );
  NAND3X0 U13787 ( .IN1(n10394), .IN2(g17819), .IN3(test_so28), .QN(n13063) );
  NAND3X0 U13788 ( .IN1(g14673), .IN2(g5933), .IN3(n10398), .QN(n13062) );
  NAND2X0 U13789 ( .IN1(n9617), .IN2(n13068), .QN(n13060) );
  NAND2X0 U13790 ( .IN1(n13069), .IN2(n13070), .QN(n13068) );
  NAND2X0 U13791 ( .IN1(g5949), .IN2(g17715), .QN(n13070) );
  NAND2X0 U13792 ( .IN1(test_so13), .IN2(g17646), .QN(n13069) );
  NAND2X0 U13793 ( .IN1(n5432), .IN2(n13056), .QN(n13059) );
  NAND3X0 U13794 ( .IN1(n13071), .IN2(n13072), .IN3(n13073), .QN(n13056) );
  NAND3X0 U13795 ( .IN1(g5961), .IN2(g17607), .IN3(n10398), .QN(n13073) );
  NAND3X0 U13796 ( .IN1(g5945), .IN2(g17739), .IN3(n10394), .QN(n13072) );
  NAND3X0 U13797 ( .IN1(g14738), .IN2(g5929), .IN3(n13048), .QN(n13071) );
  NAND2X0 U13798 ( .IN1(n13074), .IN2(g12350), .QN(n13058) );
  NAND2X0 U13799 ( .IN1(n13075), .IN2(n13076), .QN(n13074) );
  NAND2X0 U13800 ( .IN1(n10394), .IN2(g5893), .QN(n13076) );
  INVX0 U13801 ( .INP(n13052), .ZN(n13075) );
  NAND3X0 U13802 ( .IN1(n13077), .IN2(n13078), .IN3(n13079), .QN(n13052) );
  NAND3X0 U13803 ( .IN1(g17739), .IN2(g5937), .IN3(n9617), .QN(n13079) );
  NAND3X0 U13804 ( .IN1(g17607), .IN2(g5953), .IN3(n13048), .QN(n13078) );
  NAND3X0 U13805 ( .IN1(g14738), .IN2(g5921), .IN3(n10398), .QN(n13077) );
  NAND3X0 U13806 ( .IN1(n13080), .IN2(n13081), .IN3(n13082), .QN(g28096) );
  NAND2X0 U13807 ( .IN1(n10417), .IN2(g4821), .QN(n13082) );
  NAND2X0 U13808 ( .IN1(n8609), .IN2(g5619), .QN(n13081) );
  NAND3X0 U13809 ( .IN1(n10407), .IN2(n12526), .IN3(n8493), .QN(n13080) );
  NAND2X0 U13810 ( .IN1(n13083), .IN2(n13084), .QN(n12526) );
  NAND2X0 U13811 ( .IN1(n5529), .IN2(n13085), .QN(n13084) );
  NAND4X0 U13812 ( .IN1(n13086), .IN2(n13087), .IN3(n13088), .IN4(n13089), 
        .QN(n13085) );
  AND3X1 U13813 ( .IN1(n13090), .IN2(n13091), .IN3(n13092), .Q(n13089) );
  NAND2X0 U13814 ( .IN1(n10409), .IN2(n13093), .QN(n13092) );
  NAND2X0 U13815 ( .IN1(n13094), .IN2(n13095), .QN(n13093) );
  NAND2X0 U13816 ( .IN1(g17678), .IN2(g5611), .QN(n13095) );
  NAND2X0 U13817 ( .IN1(test_so6), .IN2(g17604), .QN(n13094) );
  NAND3X0 U13818 ( .IN1(g14635), .IN2(g5595), .IN3(n13096), .QN(n13091) );
  NAND3X0 U13819 ( .IN1(g17813), .IN2(g5579), .IN3(n9625), .QN(n13090) );
  NAND2X0 U13820 ( .IN1(n10413), .IN2(n13097), .QN(n13088) );
  NAND2X0 U13821 ( .IN1(n13098), .IN2(n13099), .QN(n13097) );
  NAND2X0 U13822 ( .IN1(g5685), .IN2(g5567), .QN(n13099) );
  NAND2X0 U13823 ( .IN1(g13049), .IN2(g5555), .QN(n13098) );
  NAND2X0 U13824 ( .IN1(n5439), .IN2(n13100), .QN(n13087) );
  NAND2X0 U13825 ( .IN1(n13101), .IN2(g12300), .QN(n13086) );
  NAND2X0 U13826 ( .IN1(n13102), .IN2(n13103), .QN(n13101) );
  NAND2X0 U13827 ( .IN1(n9625), .IN2(g5563), .QN(n13103) );
  INVX0 U13828 ( .INP(n13104), .ZN(n13102) );
  NAND2X0 U13829 ( .IN1(n13105), .IN2(g5689), .QN(n13083) );
  NAND4X0 U13830 ( .IN1(n13106), .IN2(n13107), .IN3(n13108), .IN4(n13109), 
        .QN(n13105) );
  AND3X1 U13831 ( .IN1(n13110), .IN2(n13111), .IN3(n13112), .Q(n13109) );
  NAND2X0 U13832 ( .IN1(n13096), .IN2(n13113), .QN(n13112) );
  NAND2X0 U13833 ( .IN1(n13114), .IN2(n13115), .QN(n13113) );
  NAND2X0 U13834 ( .IN1(g5551), .IN2(g5685), .QN(n13115) );
  NAND2X0 U13835 ( .IN1(g5543), .IN2(g13049), .QN(n13114) );
  NAND3X0 U13836 ( .IN1(g5571), .IN2(g17813), .IN3(n10409), .QN(n13111) );
  NAND3X0 U13837 ( .IN1(g14635), .IN2(g5587), .IN3(n10413), .QN(n13110) );
  NAND2X0 U13838 ( .IN1(n9625), .IN2(n13116), .QN(n13108) );
  NAND2X0 U13839 ( .IN1(n13117), .IN2(n13118), .QN(n13116) );
  NAND2X0 U13840 ( .IN1(g5619), .IN2(g17604), .QN(n13118) );
  NAND2X0 U13841 ( .IN1(g5603), .IN2(g17678), .QN(n13117) );
  NAND2X0 U13842 ( .IN1(n5439), .IN2(n13104), .QN(n13107) );
  NAND3X0 U13843 ( .IN1(n13119), .IN2(n13120), .IN3(n13121), .QN(n13104) );
  NAND3X0 U13844 ( .IN1(g5615), .IN2(g17580), .IN3(n10413), .QN(n13121) );
  NAND3X0 U13845 ( .IN1(g5599), .IN2(g17711), .IN3(n10409), .QN(n13120) );
  NAND3X0 U13846 ( .IN1(g14694), .IN2(g5583), .IN3(n13096), .QN(n13119) );
  NAND2X0 U13847 ( .IN1(n13122), .IN2(g12300), .QN(n13106) );
  NAND2X0 U13848 ( .IN1(n13123), .IN2(n13124), .QN(n13122) );
  NAND2X0 U13849 ( .IN1(n10409), .IN2(g5547), .QN(n13124) );
  INVX0 U13850 ( .INP(n13100), .ZN(n13123) );
  NAND3X0 U13851 ( .IN1(n13125), .IN2(n13126), .IN3(n13127), .QN(n13100) );
  NAND3X0 U13852 ( .IN1(n9625), .IN2(g17711), .IN3(test_so5), .QN(n13127) );
  NAND3X0 U13853 ( .IN1(g17580), .IN2(g5607), .IN3(n13096), .QN(n13126) );
  NAND3X0 U13854 ( .IN1(g14694), .IN2(g5575), .IN3(n10413), .QN(n13125) );
  NAND3X0 U13855 ( .IN1(n13128), .IN2(n13129), .IN3(n13130), .QN(g28093) );
  NAND2X0 U13856 ( .IN1(n10429), .IN2(g29220), .QN(n13130) );
  NAND2X0 U13857 ( .IN1(n8609), .IN2(g5272), .QN(n13129) );
  NAND3X0 U13858 ( .IN1(n12555), .IN2(g33959), .IN3(n8493), .QN(n13128) );
  NAND2X0 U13859 ( .IN1(n13131), .IN2(n13132), .QN(n12555) );
  NAND2X0 U13860 ( .IN1(test_so10), .IN2(n13133), .QN(n13132) );
  NAND4X0 U13861 ( .IN1(n13134), .IN2(n13135), .IN3(n13136), .IN4(n13137), 
        .QN(n13133) );
  AND3X1 U13862 ( .IN1(n13138), .IN2(n13139), .IN3(n13140), .Q(n13137) );
  NAND2X0 U13863 ( .IN1(n8813), .IN2(n13141), .QN(n13140) );
  NAND2X0 U13864 ( .IN1(n13142), .IN2(n13143), .QN(n13141) );
  NAND2X0 U13865 ( .IN1(g5339), .IN2(g5204), .QN(n13143) );
  NAND2X0 U13866 ( .IN1(g13039), .IN2(g5196), .QN(n13142) );
  NAND3X0 U13867 ( .IN1(g14597), .IN2(g5240), .IN3(n8812), .QN(n13139) );
  NAND3X0 U13868 ( .IN1(g5224), .IN2(g17787), .IN3(n8814), .QN(n13138) );
  NAND2X0 U13869 ( .IN1(g31860), .IN2(n13144), .QN(n13136) );
  NAND2X0 U13870 ( .IN1(n13145), .IN2(n13146), .QN(n13144) );
  NAND2X0 U13871 ( .IN1(g5272), .IN2(g17577), .QN(n13146) );
  NAND2X0 U13872 ( .IN1(g5256), .IN2(g17639), .QN(n13145) );
  NAND2X0 U13873 ( .IN1(n5438), .IN2(n13147), .QN(n13135) );
  NAND2X0 U13874 ( .IN1(n13148), .IN2(g12238), .QN(n13134) );
  NAND2X0 U13875 ( .IN1(n13149), .IN2(n13150), .QN(n13148) );
  NAND2X0 U13876 ( .IN1(n8814), .IN2(g5200), .QN(n13150) );
  INVX0 U13877 ( .INP(n13151), .ZN(n13149) );
  NAND2X0 U13878 ( .IN1(n13152), .IN2(n8236), .QN(n13131) );
  NAND4X0 U13879 ( .IN1(n13153), .IN2(n13154), .IN3(n13155), .IN4(n13156), 
        .QN(n13152) );
  AND3X1 U13880 ( .IN1(n13157), .IN2(n13158), .IN3(n13159), .Q(n13156) );
  NAND2X0 U13881 ( .IN1(n8812), .IN2(n13160), .QN(n13159) );
  NAND2X0 U13882 ( .IN1(n13161), .IN2(n13162), .QN(n13160) );
  NAND2X0 U13883 ( .IN1(g5220), .IN2(g5339), .QN(n13162) );
  NAND2X0 U13884 ( .IN1(g5208), .IN2(g13039), .QN(n13161) );
  NAND3X0 U13885 ( .IN1(g14597), .IN2(g5248), .IN3(n8813), .QN(n13158) );
  NAND3X0 U13886 ( .IN1(g17787), .IN2(g5232), .IN3(g31860), .QN(n13157) );
  NAND2X0 U13887 ( .IN1(n8814), .IN2(n13163), .QN(n13155) );
  NAND2X0 U13888 ( .IN1(n13164), .IN2(n13165), .QN(n13163) );
  NAND2X0 U13889 ( .IN1(g17639), .IN2(g5264), .QN(n13165) );
  NAND2X0 U13890 ( .IN1(g17577), .IN2(g5212), .QN(n13164) );
  NAND2X0 U13891 ( .IN1(n5438), .IN2(n13151), .QN(n13154) );
  NAND3X0 U13892 ( .IN1(n13166), .IN2(n13167), .IN3(n13168), .QN(n13151) );
  NAND3X0 U13893 ( .IN1(g17674), .IN2(g5244), .IN3(g31860), .QN(n13168) );
  NAND3X0 U13894 ( .IN1(n8812), .IN2(g14662), .IN3(test_so82), .QN(n13167) );
  NAND3X0 U13895 ( .IN1(g17519), .IN2(g5260), .IN3(n8813), .QN(n13166) );
  NAND2X0 U13896 ( .IN1(n13169), .IN2(g12238), .QN(n13153) );
  NAND2X0 U13897 ( .IN1(n13170), .IN2(n13171), .QN(n13169) );
  NAND2X0 U13898 ( .IN1(g31860), .IN2(g5216), .QN(n13171) );
  NOR2X0 U13899 ( .IN1(n5393), .IN2(n5588), .QN(g31860) );
  INVX0 U13900 ( .INP(n13147), .ZN(n13170) );
  NAND3X0 U13901 ( .IN1(n13172), .IN2(n13173), .IN3(n13174), .QN(n13147) );
  NAND3X0 U13902 ( .IN1(g5252), .IN2(g17674), .IN3(n8814), .QN(n13174) );
  NOR2X0 U13903 ( .IN1(g5297), .IN2(n5393), .QN(n8814) );
  NAND3X0 U13904 ( .IN1(g5268), .IN2(g17519), .IN3(n8812), .QN(n13173) );
  NOR2X0 U13905 ( .IN1(g5357), .IN2(n5588), .QN(n8812) );
  NAND3X0 U13906 ( .IN1(g14662), .IN2(g5236), .IN3(n8813), .QN(n13172) );
  NOR2X0 U13907 ( .IN1(g5297), .IN2(g5357), .QN(n8813) );
  NAND2X0 U13908 ( .IN1(n13175), .IN2(n13176), .QN(g28092) );
  NAND2X0 U13909 ( .IN1(n8608), .IN2(g5057), .QN(n13176) );
  NAND2X0 U13910 ( .IN1(n11322), .IN2(n8523), .QN(n13175) );
  NAND2X0 U13911 ( .IN1(n13177), .IN2(n13178), .QN(n11322) );
  INVX0 U13912 ( .INP(n13179), .ZN(n13178) );
  NOR3X0 U13913 ( .IN1(n5615), .IN2(n7871), .IN3(g5046), .QN(n13177) );
  NAND2X0 U13914 ( .IN1(n13180), .IN2(n13181), .QN(g28091) );
  NAND2X0 U13915 ( .IN1(n8608), .IN2(g5069), .QN(n13181) );
  NAND2X0 U13916 ( .IN1(n11321), .IN2(n8523), .QN(n13180) );
  NAND2X0 U13917 ( .IN1(n13182), .IN2(n13179), .QN(n11321) );
  NAND2X0 U13918 ( .IN1(n13183), .IN2(n13184), .QN(n13179) );
  NAND2X0 U13919 ( .IN1(g84), .IN2(g5041), .QN(n13184) );
  OR2X1 U13920 ( .IN1(g84), .IN2(n5607), .Q(n13183) );
  NOR3X0 U13921 ( .IN1(n5578), .IN2(n7842), .IN3(g5057), .QN(n13182) );
  NAND2X0 U13922 ( .IN1(n13185), .IN2(n13186), .QN(g28090) );
  NAND3X0 U13923 ( .IN1(n13187), .IN2(n8482), .IN3(n9668), .QN(n13186) );
  INVX0 U13924 ( .INP(n9666), .ZN(n9668) );
  NAND2X0 U13925 ( .IN1(n13188), .IN2(n8882), .QN(n9666) );
  NAND2X0 U13926 ( .IN1(n5770), .IN2(n13189), .QN(n13187) );
  NAND2X0 U13927 ( .IN1(n10444), .IN2(n13190), .QN(n13189) );
  NAND4X0 U13928 ( .IN1(n13191), .IN2(n13192), .IN3(n13193), .IN4(n13194), 
        .QN(n13190) );
  NAND2X0 U13929 ( .IN1(n10450), .IN2(g4045), .QN(n13194) );
  NAND2X0 U13930 ( .IN1(n7994), .IN2(n13195), .QN(n13193) );
  NAND2X0 U13931 ( .IN1(n9613), .IN2(g4049), .QN(n13192) );
  NAND2X0 U13932 ( .IN1(n7993), .IN2(n10446), .QN(n13191) );
  NAND2X0 U13933 ( .IN1(n10454), .IN2(g4961), .QN(n13185) );
  NAND2X0 U13934 ( .IN1(n13196), .IN2(n13197), .QN(g28089) );
  NAND3X0 U13935 ( .IN1(n13198), .IN2(n8482), .IN3(n9674), .QN(n13197) );
  INVX0 U13936 ( .INP(n9673), .ZN(n9674) );
  NAND2X0 U13937 ( .IN1(n13188), .IN2(n8883), .QN(n9673) );
  NAND2X0 U13938 ( .IN1(n5772), .IN2(n13199), .QN(n13198) );
  NAND2X0 U13939 ( .IN1(n10458), .IN2(n13200), .QN(n13199) );
  NAND4X0 U13940 ( .IN1(n13201), .IN2(n13202), .IN3(n13203), .IN4(n13204), 
        .QN(n13200) );
  NAND2X0 U13941 ( .IN1(n10464), .IN2(g3694), .QN(n13204) );
  NAND2X0 U13942 ( .IN1(n7990), .IN2(n13205), .QN(n13203) );
  NAND2X0 U13943 ( .IN1(n9618), .IN2(g3698), .QN(n13202) );
  NAND2X0 U13944 ( .IN1(n7989), .IN2(n10460), .QN(n13201) );
  NAND2X0 U13945 ( .IN1(n10468), .IN2(g4950), .QN(n13196) );
  NAND2X0 U13946 ( .IN1(n13206), .IN2(n13207), .QN(g28088) );
  NAND3X0 U13947 ( .IN1(n13208), .IN2(n8482), .IN3(n9682), .QN(n13207) );
  INVX0 U13948 ( .INP(n9679), .ZN(n9682) );
  NAND2X0 U13949 ( .IN1(n13188), .IN2(n8880), .QN(n9679) );
  NAND2X0 U13950 ( .IN1(n5776), .IN2(n13209), .QN(n13208) );
  NAND2X0 U13951 ( .IN1(n10477), .IN2(n13210), .QN(n13209) );
  NAND4X0 U13952 ( .IN1(n13211), .IN2(n13212), .IN3(n13213), .IN4(n13214), 
        .QN(n13210) );
  NAND2X0 U13953 ( .IN1(n10478), .IN2(g3343), .QN(n13214) );
  NAND2X0 U13954 ( .IN1(n7985), .IN2(n13215), .QN(n13213) );
  NAND2X0 U13955 ( .IN1(n9626), .IN2(g3347), .QN(n13212) );
  NAND2X0 U13956 ( .IN1(n7984), .IN2(n10479), .QN(n13211) );
  NAND2X0 U13957 ( .IN1(n10483), .IN2(g4939), .QN(n13206) );
  NAND2X0 U13958 ( .IN1(n13216), .IN2(n13217), .QN(g28087) );
  NAND3X0 U13959 ( .IN1(n13218), .IN2(n8482), .IN3(n9288), .QN(n13217) );
  INVX0 U13960 ( .INP(n9689), .ZN(n9288) );
  NAND2X0 U13961 ( .IN1(n13188), .IN2(n8881), .QN(n9689) );
  INVX0 U13962 ( .INP(n8869), .ZN(n13188) );
  NAND3X0 U13963 ( .IN1(g4966), .IN2(n8214), .IN3(g4983), .QN(n8869) );
  OR2X1 U13964 ( .IN1(n4689), .IN2(g4894), .Q(n13218) );
  NAND2X0 U13965 ( .IN1(n10372), .IN2(g4894), .QN(n13216) );
  NOR2X0 U13966 ( .IN1(n10365), .IN2(n8552), .QN(n10372) );
  INVX0 U13967 ( .INP(n8198), .ZN(n10365) );
  NAND2X0 U13968 ( .IN1(g4836), .IN2(n13219), .QN(n8198) );
  NAND3X0 U13969 ( .IN1(n8880), .IN2(g4888), .IN3(n13220), .QN(n13219) );
  NOR2X0 U13970 ( .IN1(g4899), .IN2(g4975), .QN(n8880) );
  NAND2X0 U13971 ( .IN1(n13221), .IN2(n13222), .QN(g28086) );
  NAND3X0 U13972 ( .IN1(n13223), .IN2(n8482), .IN3(n9699), .QN(n13222) );
  INVX0 U13973 ( .INP(n9697), .ZN(n9699) );
  NAND2X0 U13974 ( .IN1(n13224), .IN2(n8852), .QN(n9697) );
  NAND2X0 U13975 ( .IN1(n5769), .IN2(n13225), .QN(n13223) );
  NAND2X0 U13976 ( .IN1(n10377), .IN2(n13226), .QN(n13225) );
  NAND4X0 U13977 ( .IN1(n13227), .IN2(n13228), .IN3(n13229), .IN4(n13230), 
        .QN(n13226) );
  NAND2X0 U13978 ( .IN1(n9612), .IN2(g6390), .QN(n13230) );
  NOR2X0 U13979 ( .IN1(n5396), .IN2(n5592), .QN(n9612) );
  NAND2X0 U13980 ( .IN1(n7986), .IN2(n10379), .QN(n13229) );
  AND2X1 U13981 ( .IN1(n5592), .IN2(g6395), .Q(n10379) );
  NAND2X0 U13982 ( .IN1(n10383), .IN2(g6386), .QN(n13228) );
  NOR2X0 U13983 ( .IN1(g6395), .IN2(n5592), .QN(n10383) );
  NAND2X0 U13984 ( .IN1(n7987), .IN2(n12997), .QN(n13227) );
  AND2X1 U13985 ( .IN1(n5396), .IN2(n5592), .Q(n12997) );
  NAND2X0 U13986 ( .IN1(n10387), .IN2(g4771), .QN(n13221) );
  NOR2X0 U13987 ( .IN1(n10377), .IN2(n8552), .QN(n10387) );
  AND2X1 U13988 ( .IN1(g4688), .IN2(n13231), .Q(n10377) );
  NAND3X0 U13989 ( .IN1(n13232), .IN2(g4765), .IN3(n8854), .QN(n13231) );
  NAND2X0 U13990 ( .IN1(n13233), .IN2(n13234), .QN(g28085) );
  NAND3X0 U13991 ( .IN1(n13235), .IN2(n8482), .IN3(n9705), .QN(n13234) );
  INVX0 U13992 ( .INP(n9704), .ZN(n9705) );
  NAND2X0 U13993 ( .IN1(n13224), .IN2(n8853), .QN(n9704) );
  NAND2X0 U13994 ( .IN1(n5775), .IN2(n13236), .QN(n13235) );
  NAND2X0 U13995 ( .IN1(n10392), .IN2(n13237), .QN(n13236) );
  NAND4X0 U13996 ( .IN1(n13238), .IN2(n13239), .IN3(n13240), .IN4(n13241), 
        .QN(n13237) );
  NAND2X0 U13997 ( .IN1(n10394), .IN2(n8230), .QN(n13241) );
  AND2X1 U13998 ( .IN1(n5589), .IN2(test_so57), .Q(n10394) );
  NAND2X0 U13999 ( .IN1(test_so50), .IN2(n9617), .QN(n13240) );
  NOR2X0 U14000 ( .IN1(n8216), .IN2(n5589), .QN(n9617) );
  NAND2X0 U14001 ( .IN1(n10398), .IN2(g6040), .QN(n13239) );
  NOR2X0 U14002 ( .IN1(test_so57), .IN2(n5589), .QN(n10398) );
  NAND2X0 U14003 ( .IN1(n7988), .IN2(n13048), .QN(n13238) );
  AND2X1 U14004 ( .IN1(n5589), .IN2(n8216), .Q(n13048) );
  NAND2X0 U14005 ( .IN1(n10402), .IN2(g4760), .QN(n13233) );
  NOR2X0 U14006 ( .IN1(n10392), .IN2(n8551), .QN(n10402) );
  AND2X1 U14007 ( .IN1(g4681), .IN2(n13242), .Q(n10392) );
  NAND3X0 U14008 ( .IN1(n13232), .IN2(g4754), .IN3(n8852), .QN(n13242) );
  NOR2X0 U14009 ( .IN1(g4785), .IN2(n5518), .QN(n8852) );
  NAND2X0 U14010 ( .IN1(n13243), .IN2(n13244), .QN(g28084) );
  NAND3X0 U14011 ( .IN1(n13245), .IN2(n8483), .IN3(n9713), .QN(n13244) );
  INVX0 U14012 ( .INP(n9710), .ZN(n9713) );
  NAND2X0 U14013 ( .IN1(n13224), .IN2(n8855), .QN(n9710) );
  NAND2X0 U14014 ( .IN1(n8242), .IN2(n13246), .QN(n13245) );
  NAND2X0 U14015 ( .IN1(n10407), .IN2(n13247), .QN(n13246) );
  NAND4X0 U14016 ( .IN1(n13248), .IN2(n13249), .IN3(n13250), .IN4(n13251), 
        .QN(n13247) );
  NAND2X0 U14017 ( .IN1(n9625), .IN2(g5698), .QN(n13251) );
  NOR2X0 U14018 ( .IN1(n5397), .IN2(n5593), .QN(n9625) );
  NAND2X0 U14019 ( .IN1(n7991), .IN2(n10409), .QN(n13250) );
  AND2X1 U14020 ( .IN1(n5593), .IN2(g5703), .Q(n10409) );
  NAND2X0 U14021 ( .IN1(n10413), .IN2(g5694), .QN(n13249) );
  NOR2X0 U14022 ( .IN1(g5703), .IN2(n5593), .QN(n10413) );
  NAND2X0 U14023 ( .IN1(n7992), .IN2(n13096), .QN(n13248) );
  AND2X1 U14024 ( .IN1(n5397), .IN2(n5593), .Q(n13096) );
  NAND2X0 U14025 ( .IN1(n10417), .IN2(test_so18), .QN(n13243) );
  NOR2X0 U14026 ( .IN1(n10407), .IN2(n8551), .QN(n10417) );
  AND2X1 U14027 ( .IN1(g4674), .IN2(n13252), .Q(n10407) );
  NAND3X0 U14028 ( .IN1(n13232), .IN2(g4743), .IN3(n8853), .QN(n13252) );
  NOR2X0 U14029 ( .IN1(g4709), .IN2(n5361), .QN(n8853) );
  NAND2X0 U14030 ( .IN1(n13253), .IN2(n13254), .QN(g28083) );
  NAND3X0 U14031 ( .IN1(n13255), .IN2(n8483), .IN3(n9291), .QN(n13254) );
  INVX0 U14032 ( .INP(n9720), .ZN(n9291) );
  NAND2X0 U14033 ( .IN1(n13224), .IN2(n8854), .QN(n9720) );
  NOR2X0 U14034 ( .IN1(n5361), .IN2(n5518), .QN(n8854) );
  INVX0 U14035 ( .INP(n8841), .ZN(n13224) );
  NAND3X0 U14036 ( .IN1(g4776), .IN2(n8215), .IN3(g4793), .QN(n8841) );
  OR2X1 U14037 ( .IN1(n4708), .IN2(g4704), .Q(n13255) );
  NAND2X0 U14038 ( .IN1(n10429), .IN2(g4704), .QN(n13253) );
  NOR2X0 U14039 ( .IN1(g33959), .IN2(n8550), .QN(n10429) );
  INVX0 U14040 ( .INP(n8196), .ZN(g33959) );
  NAND2X0 U14041 ( .IN1(g4646), .IN2(n13256), .QN(n8196) );
  NAND3X0 U14042 ( .IN1(n8855), .IN2(g4698), .IN3(n13232), .QN(n13256) );
  AND4X1 U14043 ( .IN1(n5368), .IN2(g4776), .IN3(test_so19), .IN4(n13257), .Q(
        n13232) );
  NOR3X0 U14044 ( .IN1(n7691), .IN2(test_so29), .IN3(n8152), .QN(n13257) );
  NOR2X0 U14045 ( .IN1(g4709), .IN2(g4785), .QN(n8855) );
  NAND2X0 U14046 ( .IN1(n13258), .IN2(n13259), .QN(g28082) );
  NAND2X0 U14047 ( .IN1(n13260), .IN2(g4521), .QN(n13259) );
  NAND2X0 U14048 ( .IN1(n13261), .IN2(n8523), .QN(n13260) );
  XOR2X1 U14049 ( .IN1(g4527), .IN2(n13262), .Q(n13261) );
  NAND3X0 U14050 ( .IN1(n9165), .IN2(n8483), .IN3(n5752), .QN(n13258) );
  NAND3X0 U14051 ( .IN1(n13263), .IN2(n13264), .IN3(n13265), .QN(g28074) );
  NAND2X0 U14052 ( .IN1(n8607), .IN2(g4119), .QN(n13265) );
  OR3X1 U14053 ( .IN1(n8530), .IN2(n7696), .IN3(n4714), .Q(n13264) );
  NAND2X0 U14054 ( .IN1(n4714), .IN2(n4721), .QN(n13263) );
  NAND3X0 U14055 ( .IN1(n13266), .IN2(n13267), .IN3(n13268), .QN(g28073) );
  NAND2X0 U14056 ( .IN1(n13269), .IN2(n4721), .QN(n13268) );
  INVX0 U14057 ( .INP(n13270), .ZN(n13269) );
  NAND3X0 U14058 ( .IN1(n13270), .IN2(g4119), .IN3(n8493), .QN(n13267) );
  NAND2X0 U14059 ( .IN1(n13271), .IN2(g4057), .QN(n13270) );
  NAND2X0 U14060 ( .IN1(n8606), .IN2(g4116), .QN(n13266) );
  NAND3X0 U14061 ( .IN1(n13272), .IN2(n13273), .IN3(n13274), .QN(g28072) );
  NAND2X0 U14062 ( .IN1(n13275), .IN2(n4721), .QN(n13274) );
  INVX0 U14063 ( .INP(n13276), .ZN(n13275) );
  NAND3X0 U14064 ( .IN1(n13276), .IN2(g4116), .IN3(n8493), .QN(n13273) );
  NAND3X0 U14065 ( .IN1(n5711), .IN2(g4064), .IN3(n4722), .QN(n13276) );
  NAND2X0 U14066 ( .IN1(n8606), .IN2(g4112), .QN(n13272) );
  NAND2X0 U14067 ( .IN1(n13277), .IN2(n13278), .QN(g28071) );
  NAND2X0 U14068 ( .IN1(n13279), .IN2(g4112), .QN(n13278) );
  OR2X1 U14069 ( .IN1(n13279), .IN2(n8160), .Q(n13277) );
  AND2X1 U14070 ( .IN1(n13280), .IN2(n8508), .Q(n13279) );
  NAND2X0 U14071 ( .IN1(n13271), .IN2(n5711), .QN(n13280) );
  AND2X1 U14072 ( .IN1(n4722), .IN2(n5416), .Q(n13271) );
  AND4X1 U14073 ( .IN1(n7826), .IN2(n5612), .IN3(n13281), .IN4(n5350), .Q(
        n4722) );
  AND2X1 U14074 ( .IN1(n8220), .IN2(n9602), .Q(n13281) );
  NOR2X0 U14075 ( .IN1(g4093), .IN2(g4087), .QN(n9602) );
  NAND4X0 U14076 ( .IN1(n13282), .IN2(n10984), .IN3(n13283), .IN4(n13284), 
        .QN(g28070) );
  NAND3X0 U14077 ( .IN1(test_so11), .IN2(n12562), .IN3(n8493), .QN(n13284) );
  NAND2X0 U14078 ( .IN1(n8606), .IN2(g4082), .QN(n13283) );
  OR2X1 U14079 ( .IN1(n12562), .IN2(test_so11), .Q(n13282) );
  NAND2X0 U14080 ( .IN1(n13285), .IN2(g4082), .QN(n12562) );
  NAND3X0 U14081 ( .IN1(n13286), .IN2(n13287), .IN3(n13288), .QN(g28069) );
  NAND2X0 U14082 ( .IN1(n10454), .IN2(g4035), .QN(n13288) );
  NOR2X0 U14083 ( .IN1(n10444), .IN2(n8549), .QN(n10454) );
  NAND2X0 U14084 ( .IN1(n8605), .IN2(g3965), .QN(n13287) );
  NAND3X0 U14085 ( .IN1(n10444), .IN2(n12590), .IN3(n8493), .QN(n13286) );
  NAND2X0 U14086 ( .IN1(n13289), .IN2(n13290), .QN(n12590) );
  NAND2X0 U14087 ( .IN1(n5530), .IN2(n13291), .QN(n13290) );
  NAND4X0 U14088 ( .IN1(n13292), .IN2(n13293), .IN3(n13294), .IN4(n13295), 
        .QN(n13291) );
  AND3X1 U14089 ( .IN1(n13296), .IN2(n13297), .IN3(n13298), .Q(n13295) );
  NAND2X0 U14090 ( .IN1(n10450), .IN2(n13299), .QN(n13298) );
  NAND2X0 U14091 ( .IN1(n13300), .IN2(n13301), .QN(n13299) );
  NAND2X0 U14092 ( .IN1(g4031), .IN2(g3913), .QN(n13301) );
  NAND2X0 U14093 ( .IN1(g14518), .IN2(g3901), .QN(n13300) );
  NAND3X0 U14094 ( .IN1(g13906), .IN2(g3941), .IN3(n13195), .QN(n13297) );
  NAND3X0 U14095 ( .IN1(g16955), .IN2(g3925), .IN3(n9613), .QN(n13296) );
  NAND2X0 U14096 ( .IN1(n10446), .IN2(n13302), .QN(n13294) );
  NAND2X0 U14097 ( .IN1(n13303), .IN2(n13304), .QN(n13302) );
  NAND2X0 U14098 ( .IN1(g16748), .IN2(g3957), .QN(n13304) );
  NAND2X0 U14099 ( .IN1(g16693), .IN2(g3905), .QN(n13303) );
  NAND2X0 U14100 ( .IN1(n5435), .IN2(n13305), .QN(n13293) );
  NAND2X0 U14101 ( .IN1(n13306), .IN2(g11418), .QN(n13292) );
  NAND2X0 U14102 ( .IN1(n13307), .IN2(n13308), .QN(n13306) );
  NAND2X0 U14103 ( .IN1(n9613), .IN2(g3909), .QN(n13308) );
  INVX0 U14104 ( .INP(n13309), .ZN(n13307) );
  NAND2X0 U14105 ( .IN1(n13310), .IN2(g4040), .QN(n13289) );
  NAND4X0 U14106 ( .IN1(n13311), .IN2(n13312), .IN3(n13313), .IN4(n13314), 
        .QN(n13310) );
  AND3X1 U14107 ( .IN1(n13315), .IN2(n13316), .IN3(n13317), .Q(n13314) );
  NAND2X0 U14108 ( .IN1(n13195), .IN2(n13318), .QN(n13317) );
  NAND2X0 U14109 ( .IN1(n13319), .IN2(n13320), .QN(n13318) );
  NAND2X0 U14110 ( .IN1(g3897), .IN2(g4031), .QN(n13320) );
  NAND2X0 U14111 ( .IN1(test_so24), .IN2(g14518), .QN(n13319) );
  NAND3X0 U14112 ( .IN1(g13906), .IN2(g3933), .IN3(n10450), .QN(n13316) );
  NAND3X0 U14113 ( .IN1(g3917), .IN2(g16955), .IN3(n10446), .QN(n13315) );
  NAND2X0 U14114 ( .IN1(n9613), .IN2(n13321), .QN(n13313) );
  NAND2X0 U14115 ( .IN1(n13322), .IN2(n13323), .QN(n13321) );
  NAND2X0 U14116 ( .IN1(g3965), .IN2(g16693), .QN(n13323) );
  NAND2X0 U14117 ( .IN1(test_so65), .IN2(g16748), .QN(n13322) );
  NAND2X0 U14118 ( .IN1(n5435), .IN2(n13309), .QN(n13312) );
  NAND3X0 U14119 ( .IN1(n13324), .IN2(n13325), .IN3(n13326), .QN(n13309) );
  NAND3X0 U14120 ( .IN1(g3945), .IN2(g16775), .IN3(n10446), .QN(n13326) );
  NAND3X0 U14121 ( .IN1(g13966), .IN2(g3929), .IN3(n13195), .QN(n13325) );
  NAND3X0 U14122 ( .IN1(g3961), .IN2(g16659), .IN3(n10450), .QN(n13324) );
  NAND2X0 U14123 ( .IN1(n13327), .IN2(g11418), .QN(n13311) );
  NAND2X0 U14124 ( .IN1(n13328), .IN2(n13329), .QN(n13327) );
  NAND2X0 U14125 ( .IN1(n10446), .IN2(g3893), .QN(n13329) );
  AND2X1 U14126 ( .IN1(n5594), .IN2(g4054), .Q(n10446) );
  INVX0 U14127 ( .INP(n13305), .ZN(n13328) );
  NAND3X0 U14128 ( .IN1(n13330), .IN2(n13331), .IN3(n13332), .QN(n13305) );
  NAND3X0 U14129 ( .IN1(g13966), .IN2(g3921), .IN3(n10450), .QN(n13332) );
  NOR2X0 U14130 ( .IN1(g4054), .IN2(n5594), .QN(n10450) );
  NAND3X0 U14131 ( .IN1(g16659), .IN2(g3953), .IN3(n13195), .QN(n13331) );
  AND2X1 U14132 ( .IN1(n5395), .IN2(n5594), .Q(n13195) );
  NAND3X0 U14133 ( .IN1(g16775), .IN2(g3937), .IN3(n9613), .QN(n13330) );
  NOR2X0 U14134 ( .IN1(n5395), .IN2(n5594), .QN(n9613) );
  AND2X1 U14135 ( .IN1(g4878), .IN2(n13333), .Q(n10444) );
  NAND3X0 U14136 ( .IN1(n13220), .IN2(g4955), .IN3(n8881), .QN(n13333) );
  NOR2X0 U14137 ( .IN1(n5360), .IN2(n5517), .QN(n8881) );
  NAND3X0 U14138 ( .IN1(n13334), .IN2(n13335), .IN3(n13336), .QN(g28066) );
  NAND2X0 U14139 ( .IN1(n10468), .IN2(g3684), .QN(n13336) );
  NOR2X0 U14140 ( .IN1(n10458), .IN2(n8551), .QN(n10468) );
  NAND2X0 U14141 ( .IN1(n8605), .IN2(g3614), .QN(n13335) );
  NAND3X0 U14142 ( .IN1(n10458), .IN2(n12619), .IN3(n8492), .QN(n13334) );
  NAND2X0 U14143 ( .IN1(n13337), .IN2(n13338), .QN(n12619) );
  NAND2X0 U14144 ( .IN1(n5532), .IN2(n13339), .QN(n13338) );
  NAND4X0 U14145 ( .IN1(n13340), .IN2(n13341), .IN3(n13342), .IN4(n13343), 
        .QN(n13339) );
  AND3X1 U14146 ( .IN1(n13344), .IN2(n13345), .IN3(n13346), .Q(n13343) );
  NAND2X0 U14147 ( .IN1(n10464), .IN2(n13347), .QN(n13346) );
  NAND2X0 U14148 ( .IN1(n13348), .IN2(n13349), .QN(n13347) );
  NAND2X0 U14149 ( .IN1(g3680), .IN2(g3562), .QN(n13349) );
  NAND2X0 U14150 ( .IN1(g14451), .IN2(g3550), .QN(n13348) );
  NAND3X0 U14151 ( .IN1(test_so26), .IN2(g3590), .IN3(n13205), .QN(n13345) );
  NAND3X0 U14152 ( .IN1(g16924), .IN2(g3574), .IN3(n9618), .QN(n13344) );
  NAND2X0 U14153 ( .IN1(n10460), .IN2(n13350), .QN(n13342) );
  NAND2X0 U14154 ( .IN1(n13351), .IN2(n13352), .QN(n13350) );
  NAND2X0 U14155 ( .IN1(g16722), .IN2(g3606), .QN(n13352) );
  NAND2X0 U14156 ( .IN1(g16656), .IN2(g3554), .QN(n13351) );
  NAND2X0 U14157 ( .IN1(n5433), .IN2(n13353), .QN(n13341) );
  NAND2X0 U14158 ( .IN1(n13354), .IN2(g11388), .QN(n13340) );
  NAND2X0 U14159 ( .IN1(n13355), .IN2(n13356), .QN(n13354) );
  NAND2X0 U14160 ( .IN1(n9618), .IN2(g3558), .QN(n13356) );
  INVX0 U14161 ( .INP(n13357), .ZN(n13355) );
  NAND2X0 U14162 ( .IN1(n13358), .IN2(g3689), .QN(n13337) );
  NAND4X0 U14163 ( .IN1(n13359), .IN2(n13360), .IN3(n13361), .IN4(n13362), 
        .QN(n13358) );
  AND3X1 U14164 ( .IN1(n13363), .IN2(n13364), .IN3(n13365), .Q(n13362) );
  NAND2X0 U14165 ( .IN1(n13205), .IN2(n13366), .QN(n13365) );
  NAND2X0 U14166 ( .IN1(n13367), .IN2(n13368), .QN(n13366) );
  NAND2X0 U14167 ( .IN1(g3546), .IN2(g3680), .QN(n13368) );
  NAND2X0 U14168 ( .IN1(g3538), .IN2(g14451), .QN(n13367) );
  NAND3X0 U14169 ( .IN1(n10464), .IN2(g3582), .IN3(test_so26), .QN(n13364) );
  NAND3X0 U14170 ( .IN1(g3566), .IN2(g16924), .IN3(n10460), .QN(n13363) );
  NAND2X0 U14171 ( .IN1(n9618), .IN2(n13369), .QN(n13361) );
  NAND2X0 U14172 ( .IN1(n13370), .IN2(n13371), .QN(n13369) );
  NAND2X0 U14173 ( .IN1(g3614), .IN2(g16656), .QN(n13371) );
  NAND2X0 U14174 ( .IN1(g3598), .IN2(g16722), .QN(n13370) );
  NAND2X0 U14175 ( .IN1(n5433), .IN2(n13357), .QN(n13360) );
  NAND3X0 U14176 ( .IN1(n13372), .IN2(n13373), .IN3(n13374), .QN(n13357) );
  NAND3X0 U14177 ( .IN1(g3594), .IN2(g16744), .IN3(n10460), .QN(n13374) );
  NAND3X0 U14178 ( .IN1(g13926), .IN2(g3578), .IN3(n13205), .QN(n13373) );
  NAND3X0 U14179 ( .IN1(g3610), .IN2(g16627), .IN3(n10464), .QN(n13372) );
  NAND2X0 U14180 ( .IN1(n13375), .IN2(g11388), .QN(n13359) );
  NAND2X0 U14181 ( .IN1(n13376), .IN2(n13377), .QN(n13375) );
  NAND2X0 U14182 ( .IN1(n10460), .IN2(g3542), .QN(n13377) );
  AND2X1 U14183 ( .IN1(n5591), .IN2(g3703), .Q(n10460) );
  INVX0 U14184 ( .INP(n13353), .ZN(n13376) );
  NAND3X0 U14185 ( .IN1(n13378), .IN2(n13379), .IN3(n13380), .QN(n13353) );
  NAND3X0 U14186 ( .IN1(g13926), .IN2(g3570), .IN3(n10464), .QN(n13380) );
  NOR2X0 U14187 ( .IN1(g3703), .IN2(n5591), .QN(n10464) );
  NAND3X0 U14188 ( .IN1(test_so43), .IN2(g16627), .IN3(n13205), .QN(n13379) );
  AND2X1 U14189 ( .IN1(n5399), .IN2(n5591), .Q(n13205) );
  NAND3X0 U14190 ( .IN1(g16744), .IN2(g3586), .IN3(n9618), .QN(n13378) );
  NOR2X0 U14191 ( .IN1(n5399), .IN2(n5591), .QN(n9618) );
  AND2X1 U14192 ( .IN1(g4871), .IN2(n13381), .Q(n10458) );
  NAND3X0 U14193 ( .IN1(n13220), .IN2(g4944), .IN3(n8882), .QN(n13381) );
  NOR2X0 U14194 ( .IN1(g4975), .IN2(n5517), .QN(n8882) );
  NAND3X0 U14195 ( .IN1(n13382), .IN2(n13383), .IN3(n13384), .QN(g28063) );
  NAND2X0 U14196 ( .IN1(n10483), .IN2(g3333), .QN(n13384) );
  NOR2X0 U14197 ( .IN1(n10477), .IN2(n8551), .QN(n10483) );
  NAND2X0 U14198 ( .IN1(n8605), .IN2(g3263), .QN(n13383) );
  NAND3X0 U14199 ( .IN1(n10477), .IN2(n12648), .IN3(n8492), .QN(n13382) );
  NAND2X0 U14200 ( .IN1(n13385), .IN2(n13386), .QN(n12648) );
  NAND2X0 U14201 ( .IN1(n5527), .IN2(n13387), .QN(n13386) );
  NAND4X0 U14202 ( .IN1(n13388), .IN2(n13389), .IN3(n13390), .IN4(n13391), 
        .QN(n13387) );
  AND3X1 U14203 ( .IN1(n13392), .IN2(n13393), .IN3(n13394), .Q(n13391) );
  NAND2X0 U14204 ( .IN1(n10478), .IN2(n13395), .QN(n13394) );
  NAND2X0 U14205 ( .IN1(n13396), .IN2(n13397), .QN(n13395) );
  NAND2X0 U14206 ( .IN1(test_so91), .IN2(g3211), .QN(n13397) );
  NAND2X0 U14207 ( .IN1(g14421), .IN2(g3199), .QN(n13396) );
  NAND3X0 U14208 ( .IN1(g13865), .IN2(g3239), .IN3(n13215), .QN(n13393) );
  NAND3X0 U14209 ( .IN1(g16874), .IN2(g3223), .IN3(n9626), .QN(n13392) );
  NAND2X0 U14210 ( .IN1(n10479), .IN2(n13398), .QN(n13390) );
  NAND2X0 U14211 ( .IN1(n13399), .IN2(n13400), .QN(n13398) );
  NAND2X0 U14212 ( .IN1(g16686), .IN2(g3255), .QN(n13400) );
  NAND2X0 U14213 ( .IN1(g16624), .IN2(g3203), .QN(n13399) );
  NAND2X0 U14214 ( .IN1(n5436), .IN2(n13401), .QN(n13389) );
  NAND2X0 U14215 ( .IN1(n13402), .IN2(g11349), .QN(n13388) );
  NAND2X0 U14216 ( .IN1(n13403), .IN2(n13404), .QN(n13402) );
  NAND2X0 U14217 ( .IN1(n9626), .IN2(g3207), .QN(n13404) );
  INVX0 U14218 ( .INP(n13405), .ZN(n13403) );
  NAND2X0 U14219 ( .IN1(n13406), .IN2(g3338), .QN(n13385) );
  NAND4X0 U14220 ( .IN1(n13407), .IN2(n13408), .IN3(n13409), .IN4(n13410), 
        .QN(n13406) );
  AND3X1 U14221 ( .IN1(n13411), .IN2(n13412), .IN3(n13413), .Q(n13410) );
  NAND2X0 U14222 ( .IN1(n13215), .IN2(n13414), .QN(n13413) );
  NAND2X0 U14223 ( .IN1(n13415), .IN2(n13416), .QN(n13414) );
  NAND2X0 U14224 ( .IN1(g3187), .IN2(g14421), .QN(n13416) );
  NAND2X0 U14225 ( .IN1(test_so91), .IN2(test_so88), .QN(n13415) );
  NAND3X0 U14226 ( .IN1(g13865), .IN2(g3231), .IN3(n10478), .QN(n13412) );
  NAND3X0 U14227 ( .IN1(g3215), .IN2(g16874), .IN3(n10479), .QN(n13411) );
  NAND2X0 U14228 ( .IN1(n9626), .IN2(n13417), .QN(n13409) );
  NAND2X0 U14229 ( .IN1(n13418), .IN2(n13419), .QN(n13417) );
  NAND2X0 U14230 ( .IN1(g3263), .IN2(g16624), .QN(n13419) );
  NAND2X0 U14231 ( .IN1(g3247), .IN2(g16686), .QN(n13418) );
  NAND2X0 U14232 ( .IN1(n5436), .IN2(n13405), .QN(n13408) );
  NAND3X0 U14233 ( .IN1(n13420), .IN2(n13421), .IN3(n13422), .QN(n13405) );
  NAND3X0 U14234 ( .IN1(g3243), .IN2(g16718), .IN3(n10479), .QN(n13422) );
  NAND3X0 U14235 ( .IN1(g13895), .IN2(g3227), .IN3(n13215), .QN(n13421) );
  NAND3X0 U14236 ( .IN1(test_so84), .IN2(g16603), .IN3(n10478), .QN(n13420) );
  NAND2X0 U14237 ( .IN1(n13423), .IN2(g11349), .QN(n13407) );
  NAND2X0 U14238 ( .IN1(n13424), .IN2(n13425), .QN(n13423) );
  NAND2X0 U14239 ( .IN1(n10479), .IN2(g3191), .QN(n13425) );
  NOR2X0 U14240 ( .IN1(g3288), .IN2(n5604), .QN(n10479) );
  INVX0 U14241 ( .INP(n13401), .ZN(n13424) );
  NAND3X0 U14242 ( .IN1(n13426), .IN2(n13427), .IN3(n13428), .QN(n13401) );
  NAND3X0 U14243 ( .IN1(g13895), .IN2(g3219), .IN3(n10478), .QN(n13428) );
  NOR2X0 U14244 ( .IN1(g3352), .IN2(n5400), .QN(n10478) );
  NAND3X0 U14245 ( .IN1(g16603), .IN2(g3251), .IN3(n13215), .QN(n13427) );
  NOR2X0 U14246 ( .IN1(g3352), .IN2(g3288), .QN(n13215) );
  NAND3X0 U14247 ( .IN1(g16718), .IN2(g3235), .IN3(n9626), .QN(n13426) );
  NOR2X0 U14248 ( .IN1(n5400), .IN2(n5604), .QN(n9626) );
  INVX0 U14249 ( .INP(n10474), .ZN(n10477) );
  NAND2X0 U14250 ( .IN1(g4864), .IN2(n13429), .QN(n10474) );
  NAND3X0 U14251 ( .IN1(n13220), .IN2(g4933), .IN3(n8883), .QN(n13429) );
  NOR2X0 U14252 ( .IN1(g4899), .IN2(n5360), .QN(n8883) );
  AND4X1 U14253 ( .IN1(g4966), .IN2(g4859), .IN3(n5367), .IN4(n13430), .Q(
        n13220) );
  NOR3X0 U14254 ( .IN1(n7796), .IN2(test_so58), .IN3(n8151), .QN(n13430) );
  NAND4X0 U14255 ( .IN1(n13431), .IN2(n8807), .IN3(n13432), .IN4(n13433), .QN(
        g28060) );
  OR3X1 U14256 ( .IN1(n13434), .IN2(n7867), .IN3(n8532), .Q(n13433) );
  NAND2X0 U14257 ( .IN1(n8604), .IN2(g2724), .QN(n13432) );
  NAND2X0 U14258 ( .IN1(n13434), .IN2(n7867), .QN(n13431) );
  NOR2X0 U14259 ( .IN1(n12085), .IN2(n5301), .QN(n13434) );
  NAND3X0 U14260 ( .IN1(n13435), .IN2(n13436), .IN3(n13437), .QN(g28059) );
  NAND2X0 U14261 ( .IN1(n8604), .IN2(g1351), .QN(n13437) );
  NAND3X0 U14262 ( .IN1(n11225), .IN2(n7836), .IN3(n12360), .QN(n13436) );
  AND2X1 U14263 ( .IN1(n10801), .IN2(n8508), .Q(n11225) );
  AND4X1 U14264 ( .IN1(n5466), .IN2(n13438), .IN3(n13439), .IN4(n13440), .Q(
        n10801) );
  OR2X1 U14265 ( .IN1(n13441), .IN2(g1351), .Q(n13440) );
  NAND3X0 U14266 ( .IN1(n13442), .IN2(g1351), .IN3(n13441), .QN(n13439) );
  INVX0 U14267 ( .INP(n13443), .ZN(n13442) );
  NAND2X0 U14268 ( .IN1(n4798), .IN2(n13444), .QN(n13435) );
  NAND3X0 U14269 ( .IN1(n13445), .IN2(n13446), .IN3(n13447), .QN(g28058) );
  NAND2X0 U14270 ( .IN1(test_so77), .IN2(n8577), .QN(n13447) );
  OR3X1 U14271 ( .IN1(n10807), .IN2(n4490), .IN3(n5554), .Q(n13446) );
  NAND2X0 U14272 ( .IN1(n4490), .IN2(n5554), .QN(n13445) );
  NAND3X0 U14273 ( .IN1(n13448), .IN2(n13449), .IN3(n13450), .QN(g28057) );
  NAND2X0 U14274 ( .IN1(n8604), .IN2(g1008), .QN(n13450) );
  NAND3X0 U14275 ( .IN1(n11239), .IN2(n7837), .IN3(n12391), .QN(n13449) );
  AND2X1 U14276 ( .IN1(n10814), .IN2(n8508), .Q(n11239) );
  AND4X1 U14277 ( .IN1(n13451), .IN2(n8223), .IN3(n13452), .IN4(n13453), .Q(
        n10814) );
  NAND3X0 U14278 ( .IN1(n13454), .IN2(n13455), .IN3(g1008), .QN(n13453) );
  NAND2X0 U14279 ( .IN1(n5321), .IN2(n13456), .QN(n13452) );
  NAND2X0 U14280 ( .IN1(n4805), .IN2(n13457), .QN(n13448) );
  INVX0 U14281 ( .INP(n12391), .ZN(n13457) );
  NAND3X0 U14282 ( .IN1(n13458), .IN2(n13459), .IN3(n13460), .QN(g28056) );
  NAND2X0 U14283 ( .IN1(n8604), .IN2(g936), .QN(n13460) );
  OR3X1 U14284 ( .IN1(n10820), .IN2(n4514), .IN3(n5555), .Q(n13459) );
  NAND2X0 U14285 ( .IN1(n4514), .IN2(n5555), .QN(n13458) );
  NAND3X0 U14286 ( .IN1(n13461), .IN2(n13462), .IN3(n13463), .QN(g28055) );
  OR2X1 U14287 ( .IN1(n8481), .IN2(n5422), .Q(n13463) );
  NAND3X0 U14288 ( .IN1(n4518), .IN2(n13464), .IN3(g827), .QN(n13462) );
  INVX0 U14289 ( .INP(n4519), .ZN(n13464) );
  NAND3X0 U14290 ( .IN1(n4519), .IN2(n12888), .IN3(n5728), .QN(n13461) );
  NAND2X0 U14291 ( .IN1(n13465), .IN2(n13466), .QN(g28054) );
  OR2X1 U14292 ( .IN1(n13467), .IN2(n7876), .Q(n13466) );
  NAND2X0 U14293 ( .IN1(n13467), .IN2(g661), .QN(n13465) );
  NAND3X0 U14294 ( .IN1(n13468), .IN2(n13469), .IN3(n13470), .QN(g28053) );
  NAND2X0 U14295 ( .IN1(n8603), .IN2(g681), .QN(n13470) );
  INVX0 U14296 ( .INP(n13471), .ZN(n13469) );
  NAND2X0 U14297 ( .IN1(n12923), .IN2(test_so87), .QN(n13468) );
  NAND2X0 U14298 ( .IN1(n13472), .IN2(n13473), .QN(g28052) );
  NAND2X0 U14299 ( .IN1(n13474), .IN2(g661), .QN(n13473) );
  NAND2X0 U14300 ( .IN1(n13467), .IN2(g718), .QN(n13472) );
  NAND2X0 U14301 ( .IN1(n13475), .IN2(n13476), .QN(g28051) );
  NAND2X0 U14302 ( .IN1(n13474), .IN2(g718), .QN(n13476) );
  NAND2X0 U14303 ( .IN1(n13467), .IN2(g655), .QN(n13475) );
  NAND2X0 U14304 ( .IN1(n13477), .IN2(n13478), .QN(g28050) );
  NAND2X0 U14305 ( .IN1(n13474), .IN2(g655), .QN(n13478) );
  NAND2X0 U14306 ( .IN1(n13467), .IN2(g650), .QN(n13477) );
  NAND3X0 U14307 ( .IN1(n13479), .IN2(n13480), .IN3(n13481), .QN(g28049) );
  NAND2X0 U14308 ( .IN1(test_so87), .IN2(n8566), .QN(n13481) );
  NAND2X0 U14309 ( .IN1(n13471), .IN2(g681), .QN(n13480) );
  NAND2X0 U14310 ( .IN1(n13474), .IN2(g650), .QN(n13479) );
  NAND3X0 U14311 ( .IN1(n13482), .IN2(n13483), .IN3(n13484), .QN(g28048) );
  NAND2X0 U14312 ( .IN1(n8603), .IN2(g29212), .QN(n13484) );
  NAND2X0 U14313 ( .IN1(n13485), .IN2(g691), .QN(n13483) );
  NAND2X0 U14314 ( .IN1(n13486), .IN2(n13487), .QN(n13485) );
  NAND3X0 U14315 ( .IN1(g703), .IN2(n8225), .IN3(n8492), .QN(n13487) );
  NAND2X0 U14316 ( .IN1(n13488), .IN2(n13489), .QN(n13482) );
  INVX0 U14317 ( .INP(n4819), .ZN(n13489) );
  NAND4X0 U14318 ( .IN1(n5520), .IN2(n5112), .IN3(n12906), .IN4(g703), .QN(
        n4819) );
  AND4X1 U14319 ( .IN1(n13490), .IN2(test_so87), .IN3(n7861), .IN4(n7860), .Q(
        n12906) );
  XOR2X1 U14320 ( .IN1(g661), .IN2(n7876), .Q(n13490) );
  NAND2X0 U14321 ( .IN1(n13491), .IN2(n13492), .QN(g28047) );
  NAND2X0 U14322 ( .IN1(n13474), .IN2(g681), .QN(n13492) );
  NAND2X0 U14323 ( .IN1(n13467), .IN2(g645), .QN(n13491) );
  NAND2X0 U14324 ( .IN1(n13493), .IN2(n13494), .QN(g28046) );
  NAND2X0 U14325 ( .IN1(n13471), .IN2(g446), .QN(n13494) );
  NOR2X0 U14326 ( .IN1(n13495), .IN2(n8547), .QN(n13471) );
  NAND2X0 U14327 ( .IN1(n13474), .IN2(g645), .QN(n13493) );
  INVX0 U14328 ( .INP(n13467), .ZN(n13474) );
  NAND2X0 U14329 ( .IN1(n13495), .IN2(n8523), .QN(n13467) );
  NAND3X0 U14330 ( .IN1(n13496), .IN2(n13497), .IN3(n13498), .QN(n13495) );
  NAND2X0 U14331 ( .IN1(n5520), .IN2(n13499), .QN(n13497) );
  NAND3X0 U14332 ( .IN1(n5629), .IN2(g417), .IN3(n7833), .QN(n13499) );
  NAND2X0 U14333 ( .IN1(n13500), .IN2(g691), .QN(n13496) );
  NAND2X0 U14334 ( .IN1(n5287), .IN2(n8221), .QN(n13500) );
  NAND3X0 U14335 ( .IN1(n13501), .IN2(n13502), .IN3(n13503), .QN(g28045) );
  NAND2X0 U14336 ( .IN1(n8603), .IN2(g568), .QN(n13503) );
  NAND3X0 U14337 ( .IN1(n2421), .IN2(n13504), .IN3(g572), .QN(n13502) );
  INVX0 U14338 ( .INP(n4537), .ZN(n13504) );
  NAND2X0 U14339 ( .IN1(n4537), .IN2(n5337), .QN(n13501) );
  NAND2X0 U14340 ( .IN1(n13505), .IN2(n13506), .QN(g28044) );
  NAND2X0 U14341 ( .IN1(n8603), .IN2(g528), .QN(n13506) );
  NAND2X0 U14342 ( .IN1(n13507), .IN2(n8523), .QN(n13505) );
  NAND2X0 U14343 ( .IN1(n13508), .IN2(n12917), .QN(n13507) );
  XOR2X1 U14344 ( .IN1(g482), .IN2(n12919), .Q(n13508) );
  NAND2X0 U14345 ( .IN1(n13509), .IN2(n13510), .QN(n12919) );
  NAND2X0 U14346 ( .IN1(n5327), .IN2(n13511), .QN(n13510) );
  NAND2X0 U14347 ( .IN1(n13512), .IN2(n13513), .QN(g28043) );
  NAND2X0 U14348 ( .IN1(n8194), .IN2(n8228), .QN(n13513) );
  AND2X1 U14349 ( .IN1(n11266), .IN2(n8508), .Q(n8194) );
  AND4X1 U14350 ( .IN1(n13514), .IN2(n12408), .IN3(n13515), .IN4(g691), .Q(
        n11266) );
  NAND4X0 U14351 ( .IN1(n13516), .IN2(n13517), .IN3(n13518), .IN4(n13519), 
        .QN(n12408) );
  NAND3X0 U14352 ( .IN1(g753), .IN2(g718), .IN3(g655), .QN(n13519) );
  NAND3X0 U14353 ( .IN1(n7905), .IN2(n7771), .IN3(n7906), .QN(n13518) );
  NAND2X0 U14354 ( .IN1(g807), .IN2(g554), .QN(n13517) );
  NAND2X0 U14355 ( .IN1(g278), .IN2(n13520), .QN(n13514) );
  NAND2X0 U14356 ( .IN1(n8603), .IN2(g278), .QN(n13512) );
  NAND3X0 U14357 ( .IN1(n5796), .IN2(n8483), .IN3(n5630), .QN(g28042) );
  NAND3X0 U14358 ( .IN1(n11245), .IN2(n8483), .IN3(n9311), .QN(g28041) );
  NAND2X0 U14359 ( .IN1(g1536), .IN2(n4836), .QN(n9311) );
  NAND2X0 U14360 ( .IN1(g1193), .IN2(n4837), .QN(n11245) );
  NAND2X0 U14361 ( .IN1(n13521), .IN2(n13522), .QN(g28030) );
  NAND3X0 U14362 ( .IN1(n5861), .IN2(n13523), .IN3(n5882), .QN(n13522) );
  NAND2X0 U14363 ( .IN1(n13524), .IN2(n13525), .QN(n13523) );
  NAND2X0 U14364 ( .IN1(n13526), .IN2(n9254), .QN(n13525) );
  NAND2X0 U14365 ( .IN1(n13527), .IN2(n13528), .QN(n13526) );
  NAND3X0 U14366 ( .IN1(n5872), .IN2(n13529), .IN3(n5886), .QN(n13528) );
  NAND2X0 U14367 ( .IN1(n13530), .IN2(n13531), .QN(n13529) );
  NAND2X0 U14368 ( .IN1(n13532), .IN2(n13533), .QN(n13531) );
  NAND2X0 U14369 ( .IN1(n13534), .IN2(n13535), .QN(n13532) );
  NAND4X0 U14370 ( .IN1(n5885), .IN2(n5869), .IN3(n13536), .IN4(n13537), .QN(
        n13535) );
  NAND2X0 U14371 ( .IN1(n13538), .IN2(n13539), .QN(n13537) );
  NAND2X0 U14372 ( .IN1(n5873), .IN2(n8233), .QN(n13539) );
  NAND2X0 U14373 ( .IN1(n5888), .IN2(n5874), .QN(n13538) );
  OR2X1 U14374 ( .IN1(n13540), .IN2(n13541), .Q(n13536) );
  NAND2X0 U14375 ( .IN1(n13541), .IN2(n13540), .QN(n13534) );
  NAND2X0 U14376 ( .IN1(n13542), .IN2(n13533), .QN(n13527) );
  NAND2X0 U14377 ( .IN1(n9253), .IN2(n9254), .QN(n13521) );
  NAND2X0 U14378 ( .IN1(n13543), .IN2(n8523), .QN(n9254) );
  NAND2X0 U14379 ( .IN1(n5889), .IN2(n5868), .QN(n13543) );
  INVX0 U14380 ( .INP(n13524), .ZN(n9253) );
  NAND3X0 U14381 ( .IN1(n13544), .IN2(n13533), .IN3(n13542), .QN(n13524) );
  INVX0 U14382 ( .INP(n13530), .ZN(n13542) );
  NAND3X0 U14383 ( .IN1(n13541), .IN2(n13540), .IN3(n13545), .QN(n13530) );
  NAND2X0 U14384 ( .IN1(n13546), .IN2(n8523), .QN(n13545) );
  NAND2X0 U14385 ( .IN1(n5885), .IN2(n5869), .QN(n13546) );
  NAND2X0 U14386 ( .IN1(n13547), .IN2(n8523), .QN(n13540) );
  NAND2X0 U14387 ( .IN1(n5884), .IN2(n5870), .QN(n13547) );
  NAND2X0 U14388 ( .IN1(n13548), .IN2(n8523), .QN(n13541) );
  NAND4X0 U14389 ( .IN1(n5888), .IN2(n5874), .IN3(n5873), .IN4(n8233), .QN(
        n13548) );
  NAND2X0 U14390 ( .IN1(n13549), .IN2(n8523), .QN(n13533) );
  NAND2X0 U14391 ( .IN1(n5883), .IN2(n5871), .QN(n13549) );
  NAND2X0 U14392 ( .IN1(n13550), .IN2(n8523), .QN(n13544) );
  NAND2X0 U14393 ( .IN1(n5886), .IN2(n5872), .QN(n13550) );
  NAND3X0 U14394 ( .IN1(n13551), .IN2(n13552), .IN3(n11329), .QN(g26971) );
  NAND2X0 U14395 ( .IN1(n5670), .IN2(n8523), .QN(n11329) );
  NAND2X0 U14396 ( .IN1(n14516), .IN2(n8523), .QN(n13552) );
  NAND2X0 U14397 ( .IN1(n8603), .IN2(g4512), .QN(n13551) );
  NAND2X0 U14398 ( .IN1(n13553), .IN2(n13554), .QN(g26970) );
  NAND2X0 U14399 ( .IN1(n8511), .IN2(g4473), .QN(n13554) );
  NAND2X0 U14400 ( .IN1(n8602), .IN2(g4459), .QN(n13553) );
  NAND2X0 U14401 ( .IN1(n13555), .IN2(n13556), .QN(g26969) );
  NAND2X0 U14402 ( .IN1(n8602), .IN2(g4462), .QN(n13556) );
  NAND3X0 U14403 ( .IN1(n7794), .IN2(n8222), .IN3(n8492), .QN(n13555) );
  NAND2X0 U14404 ( .IN1(n13557), .IN2(n13558), .QN(g26968) );
  NAND2X0 U14405 ( .IN1(n8602), .IN2(g4558), .QN(n13557) );
  NAND2X0 U14406 ( .IN1(n13559), .IN2(n13560), .QN(g26967) );
  NAND2X0 U14407 ( .IN1(n8602), .IN2(g4561), .QN(n13559) );
  NAND2X0 U14408 ( .IN1(n13561), .IN2(n13562), .QN(g26966) );
  NAND2X0 U14409 ( .IN1(n8602), .IN2(g4555), .QN(n13561) );
  XOR2X1 U14410 ( .IN1(DFF_228_n1), .IN2(n13563), .Q(g26965) );
  NAND2X0 U14411 ( .IN1(n8511), .IN2(g10306), .QN(n13563) );
  NAND2X0 U14412 ( .IN1(n13564), .IN2(n13565), .QN(g26964) );
  NAND3X0 U14413 ( .IN1(n13566), .IN2(n13567), .IN3(n8492), .QN(n13565) );
  NAND2X0 U14414 ( .IN1(n8134), .IN2(g4521), .QN(n13567) );
  NAND2X0 U14415 ( .IN1(n5752), .IN2(n13568), .QN(n13566) );
  NAND2X0 U14416 ( .IN1(n8159), .IN2(n9843), .QN(n13568) );
  INVX0 U14417 ( .INP(n13262), .ZN(n9843) );
  NAND2X0 U14418 ( .IN1(n13569), .IN2(g4527), .QN(n13564) );
  NAND2X0 U14419 ( .IN1(n13570), .IN2(n8523), .QN(n13569) );
  NAND2X0 U14420 ( .IN1(n5752), .IN2(n13262), .QN(n13570) );
  NAND4X0 U14421 ( .IN1(test_so27), .IN2(g4483), .IN3(g4489), .IN4(g4492), 
        .QN(n13262) );
  NAND2X0 U14422 ( .IN1(n13571), .IN2(n13560), .QN(g26963) );
  NAND2X0 U14423 ( .IN1(g6750), .IN2(n8523), .QN(n13560) );
  NAND2X0 U14424 ( .IN1(n8602), .IN2(g4489), .QN(n13571) );
  NAND2X0 U14425 ( .IN1(n13558), .IN2(n13572), .QN(g26962) );
  NAND2X0 U14426 ( .IN1(test_so27), .IN2(n8660), .QN(n13572) );
  NAND2X0 U14427 ( .IN1(g6749), .IN2(n8523), .QN(n13558) );
  NAND2X0 U14428 ( .IN1(n13573), .IN2(n13562), .QN(g26961) );
  NAND2X0 U14429 ( .IN1(g6748), .IN2(n8526), .QN(n13562) );
  NAND2X0 U14430 ( .IN1(n8602), .IN2(g4483), .QN(n13573) );
  NAND2X0 U14431 ( .IN1(n13574), .IN2(n13575), .QN(g26958) );
  NAND2X0 U14432 ( .IN1(n8601), .IN2(g4455), .QN(n13575) );
  NAND2X0 U14433 ( .IN1(n13576), .IN2(n13577), .QN(g26957) );
  NAND2X0 U14434 ( .IN1(n13578), .IN2(g4434), .QN(n13577) );
  NAND2X0 U14435 ( .IN1(n13579), .IN2(n8517), .QN(n13578) );
  NAND2X0 U14436 ( .IN1(n13580), .IN2(g4392), .QN(n13579) );
  NAND2X0 U14437 ( .IN1(test_so47), .IN2(n8513), .QN(n13576) );
  NAND2X0 U14438 ( .IN1(n14518), .IN2(n13581), .QN(g26956) );
  NAND3X0 U14439 ( .IN1(n13580), .IN2(g4430), .IN3(n13582), .QN(n13581) );
  NAND2X0 U14440 ( .IN1(n13583), .IN2(n13584), .QN(g26955) );
  NAND3X0 U14441 ( .IN1(n8502), .IN2(g4392), .IN3(n13580), .QN(n13584) );
  NAND2X0 U14442 ( .IN1(n13585), .IN2(g4438), .QN(n13583) );
  NAND3X0 U14443 ( .IN1(n13586), .IN2(n13587), .IN3(n13588), .QN(g26954) );
  NAND2X0 U14444 ( .IN1(test_so47), .IN2(n8661), .QN(n13588) );
  NAND2X0 U14445 ( .IN1(n13582), .IN2(n13580), .QN(n13587) );
  AND4X1 U14446 ( .IN1(n14518), .IN2(n8139), .IN3(n13589), .IN4(DFF_1225_n1), 
        .Q(n13580) );
  NOR2X0 U14447 ( .IN1(test_so47), .IN2(g7260), .QN(n13589) );
  NAND2X0 U14448 ( .IN1(n13590), .IN2(g4438), .QN(n13586) );
  NAND2X0 U14449 ( .IN1(n13591), .IN2(n13592), .QN(g26952) );
  NAND2X0 U14450 ( .IN1(n13593), .IN2(g4430), .QN(n13592) );
  NAND2X0 U14451 ( .IN1(n8511), .IN2(g4388), .QN(n13593) );
  NAND2X0 U14452 ( .IN1(n13594), .IN2(n8513), .QN(n13591) );
  NAND2X0 U14453 ( .IN1(n13595), .IN2(n13596), .QN(n13594) );
  NAND2X0 U14454 ( .IN1(n7772), .IN2(g4388), .QN(n13596) );
  XOR2X1 U14455 ( .IN1(g4401), .IN2(n7768), .Q(n13595) );
  OR2X1 U14456 ( .IN1(n13597), .IN2(g26953), .Q(g26951) );
  NOR2X0 U14457 ( .IN1(n7856), .IN2(n8504), .QN(n13597) );
  NAND2X0 U14458 ( .IN1(n13574), .IN2(n13598), .QN(g26950) );
  OR2X1 U14459 ( .IN1(n8480), .IN2(n7675), .Q(n13598) );
  NAND2X0 U14460 ( .IN1(n13599), .IN2(n8513), .QN(n13574) );
  NAND2X0 U14461 ( .IN1(n13600), .IN2(n13601), .QN(n13599) );
  NAND2X0 U14462 ( .IN1(n13602), .IN2(g4392), .QN(n13601) );
  NAND2X0 U14463 ( .IN1(n13603), .IN2(n13604), .QN(g26949) );
  NAND2X0 U14464 ( .IN1(n13605), .IN2(g4401), .QN(n13604) );
  NAND2X0 U14465 ( .IN1(n13606), .IN2(n8513), .QN(n13605) );
  NAND2X0 U14466 ( .IN1(n13607), .IN2(g4392), .QN(n13606) );
  NAND2X0 U14467 ( .IN1(n8511), .IN2(g4411), .QN(n13603) );
  NAND2X0 U14468 ( .IN1(n7671), .IN2(n13608), .QN(g26948) );
  NAND3X0 U14469 ( .IN1(n13607), .IN2(g4388), .IN3(n13582), .QN(n13608) );
  NAND2X0 U14470 ( .IN1(n13609), .IN2(n13610), .QN(g26947) );
  NAND2X0 U14471 ( .IN1(n8601), .IN2(g4388), .QN(n13610) );
  NAND2X0 U14472 ( .IN1(n13611), .IN2(n8513), .QN(n13609) );
  NAND2X0 U14473 ( .IN1(n13600), .IN2(n13612), .QN(n13611) );
  NAND2X0 U14474 ( .IN1(n13613), .IN2(n13602), .QN(n13612) );
  XOR2X1 U14475 ( .IN1(n7680), .IN2(n5714), .Q(n13613) );
  NAND3X0 U14476 ( .IN1(n5710), .IN2(n13607), .IN3(n7675), .QN(n13600) );
  NAND2X0 U14477 ( .IN1(n13614), .IN2(n13615), .QN(g26946) );
  NAND3X0 U14478 ( .IN1(n8503), .IN2(g4392), .IN3(n13607), .QN(n13615) );
  NAND2X0 U14479 ( .IN1(n13585), .IN2(g4375), .QN(n13614) );
  NAND3X0 U14480 ( .IN1(n13616), .IN2(n13617), .IN3(n13618), .QN(g26945) );
  NAND2X0 U14481 ( .IN1(n8601), .IN2(g4411), .QN(n13618) );
  NAND2X0 U14482 ( .IN1(n13582), .IN2(n13607), .QN(n13617) );
  INVX0 U14483 ( .INP(n13602), .ZN(n13607) );
  NAND4X0 U14484 ( .IN1(n7680), .IN2(n7671), .IN3(n7681), .IN4(n13619), .QN(
        n13602) );
  NOR2X0 U14485 ( .IN1(g7257), .IN2(g7243), .QN(n13619) );
  NOR2X0 U14486 ( .IN1(g4392), .IN2(n8547), .QN(n13582) );
  NAND2X0 U14487 ( .IN1(n13590), .IN2(g4375), .QN(n13616) );
  INVX0 U14488 ( .INP(n13585), .ZN(n13590) );
  NAND2X0 U14489 ( .IN1(n5714), .IN2(n8513), .QN(n13585) );
  NOR2X0 U14490 ( .IN1(n8574), .IN2(n13620), .QN(g26944) );
  NOR4X0 U14491 ( .IN1(n13621), .IN2(n13622), .IN3(n8208), .IN4(n9724), .QN(
        n13620) );
  INVX0 U14492 ( .INP(n9165), .ZN(n13622) );
  NOR2X0 U14493 ( .IN1(g135), .IN2(n13623), .QN(n9165) );
  AND3X1 U14494 ( .IN1(n13624), .IN2(n13625), .IN3(n13626), .Q(n13623) );
  NAND3X0 U14495 ( .IN1(n13627), .IN2(n5608), .IN3(n13628), .QN(n13626) );
  XOR2X1 U14496 ( .IN1(g4608), .IN2(n5539), .Q(n13628) );
  XOR2X1 U14497 ( .IN1(g4593), .IN2(n5365), .Q(n13627) );
  NAND4X0 U14498 ( .IN1(n5365), .IN2(g4593), .IN3(n5274), .IN4(g4584), .QN(
        n13625) );
  NAND3X0 U14499 ( .IN1(n5303), .IN2(g4608), .IN3(n5539), .QN(n13624) );
  NAND3X0 U14500 ( .IN1(g4340), .IN2(g4633), .IN3(g4358), .QN(n13621) );
  NAND2X0 U14501 ( .IN1(n13629), .IN2(n13630), .QN(g26940) );
  NAND2X0 U14502 ( .IN1(n8601), .IN2(g4153), .QN(n13630) );
  NAND2X0 U14503 ( .IN1(n11812), .IN2(n8514), .QN(n13629) );
  NAND2X0 U14504 ( .IN1(n13631), .IN2(n13632), .QN(n11812) );
  NAND2X0 U14505 ( .IN1(g116), .IN2(g4157), .QN(n13632) );
  NAND2X0 U14506 ( .IN1(g114), .IN2(n5983), .QN(n13631) );
  NAND2X0 U14507 ( .IN1(n13633), .IN2(n13634), .QN(g26939) );
  NAND2X0 U14508 ( .IN1(n8601), .IN2(g4104), .QN(n13634) );
  NAND2X0 U14509 ( .IN1(n11810), .IN2(n8514), .QN(n13633) );
  NAND2X0 U14510 ( .IN1(n13635), .IN2(n13636), .QN(n11810) );
  NAND2X0 U14511 ( .IN1(g124), .IN2(g4146), .QN(n13636) );
  NAND2X0 U14512 ( .IN1(g120), .IN2(n5981), .QN(n13635) );
  NAND3X0 U14513 ( .IN1(n13637), .IN2(n13638), .IN3(n10984), .QN(g26938) );
  OR2X1 U14514 ( .IN1(n8481), .IN2(n5612), .Q(n13638) );
  NAND2X0 U14515 ( .IN1(n13639), .IN2(n8514), .QN(n13637) );
  XOR2X1 U14516 ( .IN1(n13285), .IN2(g4082), .Q(n13639) );
  NOR2X0 U14517 ( .IN1(n4723), .IN2(n5612), .QN(n13285) );
  NAND3X0 U14518 ( .IN1(n13640), .IN2(n13641), .IN3(n13642), .QN(g26934) );
  NAND2X0 U14519 ( .IN1(n4888), .IN2(g2827), .QN(n13642) );
  NAND2X0 U14520 ( .IN1(n13643), .IN2(n8243), .QN(n13641) );
  NAND2X0 U14521 ( .IN1(test_so37), .IN2(n8661), .QN(n13640) );
  NAND3X0 U14522 ( .IN1(n13644), .IN2(n13645), .IN3(n13646), .QN(g26933) );
  NAND2X0 U14523 ( .IN1(n4888), .IN2(test_so37), .QN(n13646) );
  NAND2X0 U14524 ( .IN1(n5840), .IN2(n13643), .QN(n13645) );
  NAND2X0 U14525 ( .IN1(n8600), .IN2(g2811), .QN(n13644) );
  NAND3X0 U14526 ( .IN1(n13647), .IN2(n13648), .IN3(n13649), .QN(g26932) );
  NAND2X0 U14527 ( .IN1(n4888), .IN2(g2811), .QN(n13649) );
  NAND2X0 U14528 ( .IN1(n5841), .IN2(n13643), .QN(n13648) );
  NAND2X0 U14529 ( .IN1(n8600), .IN2(g2799), .QN(n13647) );
  NAND3X0 U14530 ( .IN1(n13650), .IN2(n13651), .IN3(n13652), .QN(g26931) );
  NAND2X0 U14531 ( .IN1(n4888), .IN2(g2799), .QN(n13652) );
  NAND2X0 U14532 ( .IN1(n5839), .IN2(n13643), .QN(n13651) );
  NAND2X0 U14533 ( .IN1(n8600), .IN2(g29219), .QN(n13650) );
  NAND3X0 U14534 ( .IN1(n13653), .IN2(n13654), .IN3(n13655), .QN(g26930) );
  NAND2X0 U14535 ( .IN1(n4888), .IN2(g2795), .QN(n13655) );
  NAND2X0 U14536 ( .IN1(n13643), .IN2(n8244), .QN(n13654) );
  NAND2X0 U14537 ( .IN1(n8600), .IN2(g2791), .QN(n13653) );
  NAND3X0 U14538 ( .IN1(n13656), .IN2(n13657), .IN3(n13658), .QN(g26929) );
  NAND2X0 U14539 ( .IN1(n4888), .IN2(g2791), .QN(n13658) );
  NAND2X0 U14540 ( .IN1(n5837), .IN2(n13643), .QN(n13657) );
  NAND2X0 U14541 ( .IN1(n8600), .IN2(g2779), .QN(n13656) );
  NAND3X0 U14542 ( .IN1(n13659), .IN2(n13660), .IN3(n13661), .QN(g26928) );
  NAND2X0 U14543 ( .IN1(n4888), .IN2(g2779), .QN(n13661) );
  NAND2X0 U14544 ( .IN1(n5834), .IN2(n13643), .QN(n13660) );
  NAND2X0 U14545 ( .IN1(n8600), .IN2(g2767), .QN(n13659) );
  NAND3X0 U14546 ( .IN1(n13662), .IN2(n13663), .IN3(n13664), .QN(g26927) );
  NAND2X0 U14547 ( .IN1(n4888), .IN2(g2767), .QN(n13664) );
  NAND2X0 U14548 ( .IN1(n5836), .IN2(n13643), .QN(n13663) );
  AND3X1 U14549 ( .IN1(n9580), .IN2(n8896), .IN3(n4888), .Q(n13643) );
  NAND2X0 U14550 ( .IN1(n5516), .IN2(n5300), .QN(n8896) );
  NAND3X0 U14551 ( .IN1(n3505), .IN2(g2735), .IN3(test_so30), .QN(n9580) );
  NOR2X0 U14552 ( .IN1(n5349), .IN2(n5516), .QN(n3505) );
  OR2X1 U14553 ( .IN1(n8480), .IN2(n7689), .Q(n13662) );
  NAND2X0 U14554 ( .IN1(n13665), .IN2(n13666), .QN(g26926) );
  NAND2X0 U14555 ( .IN1(n13667), .IN2(n3730), .QN(n13666) );
  XOR2X1 U14556 ( .IN1(g2724), .IN2(n12078), .Q(n13667) );
  INVX0 U14557 ( .INP(n12085), .ZN(n12078) );
  NAND2X0 U14558 ( .IN1(g2719), .IN2(g2715), .QN(n12085) );
  NAND2X0 U14559 ( .IN1(n8599), .IN2(g2719), .QN(n13665) );
  NAND2X0 U14560 ( .IN1(n13668), .IN2(n13669), .QN(g26925) );
  NAND2X0 U14561 ( .IN1(n8599), .IN2(g1532), .QN(n13669) );
  NAND2X0 U14562 ( .IN1(n13670), .IN2(n8514), .QN(n13668) );
  NAND2X0 U14563 ( .IN1(n12354), .IN2(n13671), .QN(n13670) );
  NAND2X0 U14564 ( .IN1(n12337), .IN2(g1536), .QN(n13671) );
  NAND2X0 U14565 ( .IN1(n12341), .IN2(g1413), .QN(n12337) );
  NOR2X0 U14566 ( .IN1(n12345), .IN2(n7862), .QN(n12341) );
  NAND3X0 U14567 ( .IN1(n13672), .IN2(g7946), .IN3(n10598), .QN(n12345) );
  NAND3X0 U14568 ( .IN1(g1339), .IN2(g1521), .IN3(n7995), .QN(n13672) );
  INVX0 U14569 ( .INP(n4173), .ZN(n12354) );
  NAND3X0 U14570 ( .IN1(n13673), .IN2(n13674), .IN3(n13675), .QN(g26924) );
  OR2X1 U14571 ( .IN1(n13676), .IN2(g1478), .Q(n13675) );
  NAND3X0 U14572 ( .IN1(n13676), .IN2(g1478), .IN3(n8494), .QN(n13674) );
  NAND4X0 U14573 ( .IN1(n13677), .IN2(n10636), .IN3(g1437), .IN4(g13272), .QN(
        n13676) );
  NOR2X0 U14574 ( .IN1(test_so49), .IN2(n5364), .QN(n10636) );
  NAND2X0 U14575 ( .IN1(n8599), .IN2(g1437), .QN(n13673) );
  NAND3X0 U14576 ( .IN1(n13678), .IN2(n13679), .IN3(n13680), .QN(g26923) );
  OR2X1 U14577 ( .IN1(n13681), .IN2(g1472), .Q(n13680) );
  NAND3X0 U14578 ( .IN1(n13681), .IN2(g1472), .IN3(n8494), .QN(n13679) );
  NAND4X0 U14579 ( .IN1(n13677), .IN2(n10561), .IN3(g1467), .IN4(g13272), .QN(
        n13681) );
  NAND2X0 U14580 ( .IN1(n8599), .IN2(g1467), .QN(n13678) );
  NAND3X0 U14581 ( .IN1(n13682), .IN2(n13683), .IN3(n13684), .QN(g26922) );
  OR2X1 U14582 ( .IN1(n13685), .IN2(g1448), .Q(n13684) );
  NAND3X0 U14583 ( .IN1(n13685), .IN2(g1448), .IN3(n8494), .QN(n13683) );
  NAND3X0 U14584 ( .IN1(n12827), .IN2(g1454), .IN3(n13677), .QN(n13685) );
  AND2X1 U14585 ( .IN1(n10598), .IN2(g13272), .Q(n12827) );
  NOR2X0 U14586 ( .IN1(n8206), .IN2(g1514), .QN(n10598) );
  NAND2X0 U14587 ( .IN1(n8599), .IN2(g1454), .QN(n13682) );
  NAND2X0 U14588 ( .IN1(n13686), .IN2(n13687), .QN(g26921) );
  NAND2X0 U14589 ( .IN1(n8599), .IN2(g1395), .QN(n13687) );
  NAND3X0 U14590 ( .IN1(n13688), .IN2(n8203), .IN3(n8494), .QN(n13686) );
  XNOR2X1 U14591 ( .IN1(n13689), .IN2(n7839), .Q(n13688) );
  NAND3X0 U14592 ( .IN1(n13690), .IN2(n13691), .IN3(n13692), .QN(g26920) );
  NAND2X0 U14593 ( .IN1(n4913), .IN2(n13693), .QN(n13692) );
  NAND2X0 U14594 ( .IN1(n8598), .IN2(g1384), .QN(n13691) );
  OR3X1 U14595 ( .IN1(n4915), .IN2(n7845), .IN3(n8538), .Q(n13690) );
  AND2X1 U14596 ( .IN1(n13694), .IN2(n13695), .Q(n4915) );
  NAND2X0 U14597 ( .IN1(n7693), .IN2(g1351), .QN(n13695) );
  NAND3X0 U14598 ( .IN1(n13696), .IN2(n13697), .IN3(n13698), .QN(g26919) );
  NAND2X0 U14599 ( .IN1(n8598), .IN2(g1266), .QN(n13698) );
  NAND3X0 U14600 ( .IN1(test_so77), .IN2(n11235), .IN3(n8802), .QN(n13697) );
  OR2X1 U14601 ( .IN1(n8802), .IN2(test_so77), .Q(n13696) );
  NAND3X0 U14602 ( .IN1(g1249), .IN2(g1266), .IN3(g12923), .QN(n8802) );
  NAND2X0 U14603 ( .IN1(n13699), .IN2(n13700), .QN(g26918) );
  NAND2X0 U14604 ( .IN1(n8598), .IN2(g1189), .QN(n13700) );
  NAND2X0 U14605 ( .IN1(n13701), .IN2(n8515), .QN(n13699) );
  NAND2X0 U14606 ( .IN1(n12385), .IN2(n13702), .QN(n13701) );
  NAND2X0 U14607 ( .IN1(n12368), .IN2(g1193), .QN(n13702) );
  NAND2X0 U14608 ( .IN1(n12372), .IN2(g1070), .QN(n12368) );
  NOR2X0 U14609 ( .IN1(n12376), .IN2(n7863), .QN(n12372) );
  NAND3X0 U14610 ( .IN1(n13703), .IN2(g7916), .IN3(n10756), .QN(n12376) );
  NAND3X0 U14611 ( .IN1(g1178), .IN2(g996), .IN3(n5642), .QN(n13703) );
  INVX0 U14612 ( .INP(n4191), .ZN(n12385) );
  NAND3X0 U14613 ( .IN1(n13704), .IN2(n13705), .IN3(n13706), .QN(g26917) );
  OR2X1 U14614 ( .IN1(n13707), .IN2(g1135), .Q(n13706) );
  NAND3X0 U14615 ( .IN1(n13707), .IN2(g1135), .IN3(n8494), .QN(n13705) );
  NAND4X0 U14616 ( .IN1(n13708), .IN2(n10841), .IN3(g1094), .IN4(g13259), .QN(
        n13707) );
  NOR2X0 U14617 ( .IN1(g1183), .IN2(n5363), .QN(n10841) );
  NAND2X0 U14618 ( .IN1(n8598), .IN2(g1094), .QN(n13704) );
  NAND3X0 U14619 ( .IN1(n13709), .IN2(n13710), .IN3(n13711), .QN(g26916) );
  OR2X1 U14620 ( .IN1(n13712), .IN2(g1129), .Q(n13711) );
  NAND3X0 U14621 ( .IN1(n13712), .IN2(g1129), .IN3(n8494), .QN(n13710) );
  NAND4X0 U14622 ( .IN1(n13708), .IN2(n10718), .IN3(g1124), .IN4(g13259), .QN(
        n13712) );
  NAND2X0 U14623 ( .IN1(n8598), .IN2(g1124), .QN(n13709) );
  NAND3X0 U14624 ( .IN1(n13713), .IN2(n13714), .IN3(n13715), .QN(g26915) );
  OR2X1 U14625 ( .IN1(n13716), .IN2(g1105), .Q(n13715) );
  NAND3X0 U14626 ( .IN1(n13716), .IN2(g1105), .IN3(n8494), .QN(n13714) );
  NAND3X0 U14627 ( .IN1(test_so90), .IN2(n12859), .IN3(n13708), .QN(n13716) );
  AND2X1 U14628 ( .IN1(n10756), .IN2(g13259), .Q(n12859) );
  NOR2X0 U14629 ( .IN1(g1171), .IN2(n5599), .QN(n10756) );
  NAND2X0 U14630 ( .IN1(test_so90), .IN2(n8542), .QN(n13713) );
  NAND2X0 U14631 ( .IN1(n13717), .IN2(n13718), .QN(g26914) );
  NAND2X0 U14632 ( .IN1(n8597), .IN2(g1052), .QN(n13718) );
  NAND3X0 U14633 ( .IN1(n5320), .IN2(n13719), .IN3(n8495), .QN(n13717) );
  XNOR2X1 U14634 ( .IN1(n13720), .IN2(n7840), .Q(n13719) );
  NAND3X0 U14635 ( .IN1(n13721), .IN2(n13722), .IN3(n13723), .QN(g26913) );
  NAND2X0 U14636 ( .IN1(n4938), .IN2(n13724), .QN(n13723) );
  NAND2X0 U14637 ( .IN1(n8597), .IN2(g1041), .QN(n13722) );
  NAND3X0 U14638 ( .IN1(n8823), .IN2(g1046), .IN3(n8497), .QN(n13721) );
  NAND2X0 U14639 ( .IN1(n13725), .IN2(n13726), .QN(n8823) );
  NAND2X0 U14640 ( .IN1(n7692), .IN2(g1008), .QN(n13726) );
  NAND3X0 U14641 ( .IN1(n13727), .IN2(n13728), .IN3(n13729), .QN(g26912) );
  NAND2X0 U14642 ( .IN1(n8597), .IN2(g921), .QN(n13729) );
  NAND3X0 U14643 ( .IN1(n11250), .IN2(n13730), .IN3(g936), .QN(n13728) );
  NAND2X0 U14644 ( .IN1(n220), .IN2(n5557), .QN(n13727) );
  INVX0 U14645 ( .INP(n13730), .ZN(n220) );
  NAND3X0 U14646 ( .IN1(g921), .IN2(g904), .IN3(g12919), .QN(n13730) );
  XOR2X1 U14647 ( .IN1(n13731), .IN2(n5682), .Q(g26910) );
  NAND2X0 U14648 ( .IN1(n5305), .IN2(n8515), .QN(n13731) );
  NAND2X0 U14649 ( .IN1(n13732), .IN2(n13733), .QN(g26909) );
  NAND2X0 U14650 ( .IN1(n8597), .IN2(g890), .QN(n13733) );
  NAND2X0 U14651 ( .IN1(n13734), .IN2(n8517), .QN(n13732) );
  NAND2X0 U14652 ( .IN1(n13735), .IN2(n13736), .QN(n13734) );
  NAND2X0 U14653 ( .IN1(n5431), .IN2(g862), .QN(n13736) );
  NAND2X0 U14654 ( .IN1(n5305), .IN2(g896), .QN(n13735) );
  NAND3X0 U14655 ( .IN1(n13737), .IN2(n13738), .IN3(n13739), .QN(g26908) );
  NAND2X0 U14656 ( .IN1(n4945), .IN2(g446), .QN(n13739) );
  NAND2X0 U14657 ( .IN1(n13740), .IN2(g872), .QN(n13738) );
  NAND2X0 U14658 ( .IN1(n8597), .IN2(g246), .QN(n13737) );
  NAND3X0 U14659 ( .IN1(n13741), .IN2(n13742), .IN3(n13743), .QN(g26907) );
  NAND2X0 U14660 ( .IN1(n4945), .IN2(g246), .QN(n13743) );
  NAND2X0 U14661 ( .IN1(n13740), .IN2(g14167), .QN(n13742) );
  NAND2X0 U14662 ( .IN1(n8596), .IN2(g269), .QN(n13741) );
  NAND3X0 U14663 ( .IN1(n13744), .IN2(n13745), .IN3(n13746), .QN(g26906) );
  NAND2X0 U14664 ( .IN1(n4945), .IN2(g269), .QN(n13746) );
  NAND2X0 U14665 ( .IN1(n13740), .IN2(g14147), .QN(n13745) );
  NAND2X0 U14666 ( .IN1(n8596), .IN2(g239), .QN(n13744) );
  NAND3X0 U14667 ( .IN1(n13747), .IN2(n13748), .IN3(n13749), .QN(g26905) );
  NAND2X0 U14668 ( .IN1(n4945), .IN2(g239), .QN(n13749) );
  NAND2X0 U14669 ( .IN1(n13740), .IN2(g14125), .QN(n13748) );
  NAND2X0 U14670 ( .IN1(n8596), .IN2(g262), .QN(n13747) );
  NAND3X0 U14671 ( .IN1(n13750), .IN2(n13751), .IN3(n13752), .QN(g26904) );
  NAND2X0 U14672 ( .IN1(n4945), .IN2(g262), .QN(n13752) );
  NAND2X0 U14673 ( .IN1(n13740), .IN2(g14096), .QN(n13751) );
  NAND2X0 U14674 ( .IN1(n8607), .IN2(g232), .QN(n13750) );
  NAND3X0 U14675 ( .IN1(n13753), .IN2(n13754), .IN3(n13755), .QN(g26903) );
  NAND2X0 U14676 ( .IN1(n4945), .IN2(g232), .QN(n13755) );
  NAND2X0 U14677 ( .IN1(n13740), .IN2(g14217), .QN(n13754) );
  NAND2X0 U14678 ( .IN1(n8544), .IN2(g255), .QN(n13753) );
  NAND3X0 U14679 ( .IN1(n13756), .IN2(n13757), .IN3(n13758), .QN(g26902) );
  NAND2X0 U14680 ( .IN1(n4945), .IN2(g255), .QN(n13758) );
  NAND2X0 U14681 ( .IN1(n13740), .IN2(g14201), .QN(n13757) );
  NAND2X0 U14682 ( .IN1(n8596), .IN2(g225), .QN(n13756) );
  NAND3X0 U14683 ( .IN1(n13759), .IN2(n13760), .IN3(n13761), .QN(g26901) );
  NAND2X0 U14684 ( .IN1(n4945), .IN2(g225), .QN(n13761) );
  NAND2X0 U14685 ( .IN1(n13740), .IN2(g14189), .QN(n13760) );
  NOR2X0 U14686 ( .IN1(n8576), .IN2(n4946), .QN(n13740) );
  NAND3X0 U14687 ( .IN1(n5431), .IN2(g890), .IN3(n5682), .QN(n4946) );
  NAND2X0 U14688 ( .IN1(n8597), .IN2(g872), .QN(n13759) );
  NAND2X0 U14689 ( .IN1(n13762), .IN2(n13763), .QN(g26899) );
  NAND2X0 U14690 ( .IN1(n13764), .IN2(n4518), .QN(n13763) );
  XNOR2X1 U14691 ( .IN1(n4814), .IN2(n5422), .Q(n13764) );
  AND3X1 U14692 ( .IN1(g817), .IN2(g832), .IN3(n4948), .Q(n4814) );
  NAND2X0 U14693 ( .IN1(n8597), .IN2(g832), .QN(n13762) );
  NAND2X0 U14694 ( .IN1(n13765), .IN2(n13766), .QN(g26898) );
  NAND2X0 U14695 ( .IN1(n13767), .IN2(n13768), .QN(n13766) );
  NAND2X0 U14696 ( .IN1(n13769), .IN2(n13770), .QN(n13768) );
  NAND2X0 U14697 ( .IN1(n7804), .IN2(n8515), .QN(n13770) );
  NAND2X0 U14698 ( .IN1(n13771), .IN2(g843), .QN(n13765) );
  NAND2X0 U14699 ( .IN1(n13772), .IN2(n8515), .QN(n13771) );
  NAND3X0 U14700 ( .IN1(n5733), .IN2(g837), .IN3(n13773), .QN(n13772) );
  NAND2X0 U14701 ( .IN1(n13774), .IN2(n13775), .QN(g26897) );
  NAND2X0 U14702 ( .IN1(n13776), .IN2(g753), .QN(n13775) );
  OR2X1 U14703 ( .IN1(n13776), .IN2(n5732), .Q(n13774) );
  NOR2X0 U14704 ( .IN1(n13516), .IN2(n8549), .QN(n13776) );
  NAND3X0 U14705 ( .IN1(n13777), .IN2(n13778), .IN3(n13779), .QN(g26896) );
  NAND2X0 U14706 ( .IN1(n4956), .IN2(n12907), .QN(n13779) );
  NAND2X0 U14707 ( .IN1(n13780), .IN2(g29212), .QN(n13778) );
  OR2X1 U14708 ( .IN1(n13780), .IN2(n7876), .Q(n13777) );
  NOR2X0 U14709 ( .IN1(n12907), .IN2(n8547), .QN(n13780) );
  INVX0 U14710 ( .INP(n8195), .ZN(n12907) );
  NAND4X0 U14711 ( .IN1(n4948), .IN2(n13781), .IN3(n5327), .IN4(n13782), .QN(
        n8195) );
  NOR2X0 U14712 ( .IN1(g504), .IN2(n8221), .QN(n13782) );
  INVX0 U14713 ( .INP(n13511), .ZN(n13781) );
  NAND3X0 U14714 ( .IN1(n13783), .IN2(n13784), .IN3(n13785), .QN(g26895) );
  NAND2X0 U14715 ( .IN1(n8598), .IN2(g562), .QN(n13785) );
  NAND3X0 U14716 ( .IN1(n2421), .IN2(n13786), .IN3(g568), .QN(n13784) );
  NAND2X0 U14717 ( .IN1(n5), .IN2(n5335), .QN(n13783) );
  INVX0 U14718 ( .INP(n13786), .ZN(n5) );
  NAND3X0 U14719 ( .IN1(n13787), .IN2(g562), .IN3(n4959), .QN(n13786) );
  NAND2X0 U14720 ( .IN1(n13788), .IN2(n13789), .QN(g26894) );
  NAND2X0 U14721 ( .IN1(n8598), .IN2(g518), .QN(n13789) );
  NAND4X0 U14722 ( .IN1(n13790), .IN2(n13791), .IN3(n12917), .IN4(n8506), .QN(
        n13788) );
  NAND2X0 U14723 ( .IN1(n13509), .IN2(g528), .QN(n13791) );
  NAND2X0 U14724 ( .IN1(n5327), .IN2(n13792), .QN(n13790) );
  NAND2X0 U14725 ( .IN1(n13509), .IN2(n13511), .QN(n13792) );
  NAND2X0 U14726 ( .IN1(g482), .IN2(g490), .QN(n13511) );
  NOR3X0 U14727 ( .IN1(g513), .IN2(n5287), .IN3(n13793), .QN(n13509) );
  NAND2X0 U14728 ( .IN1(n13794), .IN2(n13795), .QN(g26893) );
  OR2X1 U14729 ( .IN1(n8479), .IN2(n8136), .Q(n13795) );
  NAND2X0 U14730 ( .IN1(n13796), .IN2(n8515), .QN(n13794) );
  NAND2X0 U14731 ( .IN1(n13797), .IN2(n13798), .QN(n13796) );
  NAND2X0 U14732 ( .IN1(g29211), .IN2(n8229), .QN(n13798) );
  NAND2X0 U14733 ( .IN1(test_so17), .IN2(n13799), .QN(n13797) );
  NAND2X0 U14734 ( .IN1(n13800), .IN2(n13801), .QN(g26892) );
  NAND3X0 U14735 ( .IN1(n8503), .IN2(n13799), .IN3(n8229), .QN(n13801) );
  NAND2X0 U14736 ( .IN1(n8136), .IN2(n8135), .QN(n13799) );
  NAND2X0 U14737 ( .IN1(test_so17), .IN2(n8576), .QN(n13800) );
  NAND2X0 U14738 ( .IN1(n13802), .IN2(n13803), .QN(g26891) );
  OR2X1 U14739 ( .IN1(n8478), .IN2(n5860), .Q(n13803) );
  NAND3X0 U14740 ( .IN1(n8502), .IN2(g7540), .IN3(n5860), .QN(n13802) );
  NAND2X0 U14741 ( .IN1(n13804), .IN2(n13805), .QN(g26890) );
  NAND2X0 U14742 ( .IN1(n5860), .IN2(n8516), .QN(n13805) );
  OR2X1 U14743 ( .IN1(n8478), .IN2(n8135), .Q(n13804) );
  NAND2X0 U14744 ( .IN1(n13806), .IN2(n13807), .QN(g26889) );
  NAND2X0 U14745 ( .IN1(n8599), .IN2(g29211), .QN(n13807) );
  NAND4X0 U14746 ( .IN1(g329), .IN2(DFF_709_n1), .IN3(n13808), .IN4(n8507), 
        .QN(n13806) );
  NAND2X0 U14747 ( .IN1(n13809), .IN2(n13810), .QN(g26888) );
  NAND2X0 U14748 ( .IN1(n8510), .IN2(g316), .QN(n13810) );
  NAND2X0 U14749 ( .IN1(n8600), .IN2(g29216), .QN(n13809) );
  NAND3X0 U14750 ( .IN1(n13811), .IN2(n13812), .IN3(n13813), .QN(g26887) );
  NAND2X0 U14751 ( .IN1(n8601), .IN2(g336), .QN(n13812) );
  NAND3X0 U14752 ( .IN1(n5317), .IN2(g324), .IN3(n8495), .QN(n13811) );
  NAND3X0 U14753 ( .IN1(n13814), .IN2(n13815), .IN3(n13816), .QN(g26886) );
  OR2X1 U14754 ( .IN1(n13813), .IN2(n13808), .Q(n13816) );
  NAND3X0 U14755 ( .IN1(n13808), .IN2(g336), .IN3(n8495), .QN(n13815) );
  NAND2X0 U14756 ( .IN1(n8601), .IN2(g311), .QN(n13814) );
  NAND2X0 U14757 ( .IN1(n13817), .IN2(n13818), .QN(g26884) );
  NAND2X0 U14758 ( .IN1(n8603), .IN2(g329), .QN(n13818) );
  NAND2X0 U14759 ( .IN1(n13819), .IN2(n8516), .QN(n13817) );
  NAND2X0 U14760 ( .IN1(n13820), .IN2(n13821), .QN(n13819) );
  NAND4X0 U14761 ( .IN1(n5766), .IN2(n5456), .IN3(n5282), .IN4(n5317), .QN(
        n13821) );
  NAND2X0 U14762 ( .IN1(n13822), .IN2(n13823), .QN(n13820) );
  NAND3X0 U14763 ( .IN1(n13824), .IN2(n13825), .IN3(n5456), .QN(n13823) );
  NAND2X0 U14764 ( .IN1(n5824), .IN2(g311), .QN(n13825) );
  NAND2X0 U14765 ( .IN1(g305), .IN2(g336), .QN(n13824) );
  NAND2X0 U14766 ( .IN1(n13826), .IN2(n13827), .QN(g26883) );
  NAND2X0 U14767 ( .IN1(n8604), .IN2(g324), .QN(n13827) );
  NAND2X0 U14768 ( .IN1(n13822), .IN2(n8516), .QN(n13826) );
  INVX0 U14769 ( .INP(n13808), .ZN(n13822) );
  NAND2X0 U14770 ( .IN1(n13828), .IN2(n13829), .QN(n13808) );
  NAND2X0 U14771 ( .IN1(n5282), .IN2(g324), .QN(n13829) );
  NAND2X0 U14772 ( .IN1(n5827), .IN2(n5317), .QN(n13828) );
  NAND3X0 U14773 ( .IN1(n13830), .IN2(n13831), .IN3(n13813), .QN(g26882) );
  NAND2X0 U14774 ( .IN1(n8510), .IN2(g305), .QN(n13813) );
  NAND2X0 U14775 ( .IN1(n8510), .IN2(g311), .QN(n13831) );
  NAND2X0 U14776 ( .IN1(n8604), .IN2(g316), .QN(n13830) );
  NAND2X0 U14777 ( .IN1(n13832), .IN2(n13833), .QN(g26881) );
  NAND2X0 U14778 ( .IN1(g6744), .IN2(n8516), .QN(n13833) );
  NAND2X0 U14779 ( .IN1(n8604), .IN2(g305), .QN(n13832) );
  NAND3X0 U14780 ( .IN1(n9248), .IN2(n8481), .IN3(n9249), .QN(g26877) );
  NAND4X0 U14781 ( .IN1(n5620), .IN2(n5619), .IN3(n13834), .IN4(n13835), .QN(
        n9249) );
  NOR4X0 U14782 ( .IN1(test_so40), .IN2(g2357), .IN3(g2338), .IN4(g2606), .QN(
        n13835) );
  NOR2X0 U14783 ( .IN1(g2491), .IN2(g2223), .QN(n13834) );
  NAND4X0 U14784 ( .IN1(n5833), .IN2(n5832), .IN3(n13836), .IN4(n13837), .QN(
        n9248) );
  NOR4X0 U14785 ( .IN1(test_so75), .IN2(g1664), .IN3(g1913), .IN4(g1932), .QN(
        n13837) );
  NOR2X0 U14786 ( .IN1(g1779), .IN2(g2047), .QN(n13836) );
  NAND2X0 U14787 ( .IN1(n9266), .IN2(n9207), .QN(g26876) );
  NAND4X0 U14788 ( .IN1(n14521), .IN2(n5892), .IN3(n13838), .IN4(n13839), .QN(
        n9207) );
  NOR4X0 U14789 ( .IN1(g1710), .IN2(g1978), .IN3(g1844), .IN4(g2112), .QN(
        n13839) );
  NOR2X0 U14790 ( .IN1(g1992), .IN2(g2126), .QN(n13838) );
  INVX0 U14791 ( .INP(n9203), .ZN(n9266) );
  NAND2X0 U14792 ( .IN1(n13840), .IN2(n8516), .QN(n9203) );
  NAND4X0 U14793 ( .IN1(n14517), .IN2(n14522), .IN3(n13841), .IN4(n13842), 
        .QN(n13840) );
  NOR4X0 U14794 ( .IN1(test_so31), .IN2(g2671), .IN3(g2269), .IN4(g2537), .QN(
        n13842) );
  NOR2X0 U14795 ( .IN1(n9324), .IN2(n9295), .QN(n13841) );
  NAND2X0 U14796 ( .IN1(n9271), .IN2(n9208), .QN(g26875) );
  NAND4X0 U14797 ( .IN1(n5628), .IN2(n5413), .IN3(n5315), .IN4(n5280), .QN(
        n9208) );
  INVX0 U14798 ( .INP(n9204), .ZN(n9271) );
  NAND2X0 U14799 ( .IN1(n13843), .IN2(n8516), .QN(n9204) );
  NAND4X0 U14800 ( .IN1(n5631), .IN2(n5414), .IN3(n5316), .IN4(n5281), .QN(
        n13843) );
  NAND2X0 U14801 ( .IN1(n13844), .IN2(n13845), .QN(g25764) );
  NAND2X0 U14802 ( .IN1(n11401), .IN2(g6505), .QN(n13845) );
  NAND2X0 U14803 ( .IN1(n13846), .IN2(g6541), .QN(n13844) );
  NAND3X0 U14804 ( .IN1(n13847), .IN2(n13848), .IN3(n13849), .QN(g25763) );
  OR2X1 U14805 ( .IN1(n13846), .IN2(n5884), .Q(n13849) );
  NAND2X0 U14806 ( .IN1(n13850), .IN2(g6533), .QN(n13848) );
  NAND2X0 U14807 ( .IN1(n13851), .IN2(n8516), .QN(n13850) );
  NAND2X0 U14808 ( .IN1(n10354), .IN2(g6527), .QN(n13851) );
  NAND4X0 U14809 ( .IN1(n10354), .IN2(n8505), .IN3(n5659), .IN4(n5445), .QN(
        n13847) );
  NAND2X0 U14810 ( .IN1(n13852), .IN2(n13853), .QN(g25762) );
  NAND2X0 U14811 ( .IN1(n11401), .IN2(g6533), .QN(n13853) );
  NAND2X0 U14812 ( .IN1(n13846), .IN2(g6527), .QN(n13852) );
  INVX0 U14813 ( .INP(n11401), .ZN(n13846) );
  NAND3X0 U14814 ( .IN1(n13854), .IN2(n13855), .IN3(n13856), .QN(g25761) );
  NAND2X0 U14815 ( .IN1(n11401), .IN2(g6513), .QN(n13856) );
  NOR2X0 U14816 ( .IN1(n10354), .IN2(n8553), .QN(n11401) );
  NAND3X0 U14817 ( .IN1(n5426), .IN2(n10354), .IN3(n8492), .QN(n13855) );
  NOR2X0 U14818 ( .IN1(n3776), .IN2(n5646), .QN(n10354) );
  NAND2X0 U14819 ( .IN1(g6573), .IN2(g6565), .QN(n3776) );
  NAND2X0 U14820 ( .IN1(n8605), .IN2(g6509), .QN(n13854) );
  NAND2X0 U14821 ( .IN1(n13857), .IN2(n13858), .QN(g25758) );
  OR2X1 U14822 ( .IN1(n8478), .IN2(n7729), .Q(n13858) );
  NAND3X0 U14823 ( .IN1(n7728), .IN2(n13859), .IN3(n8496), .QN(n13857) );
  NAND2X0 U14824 ( .IN1(n5990), .IN2(n13860), .QN(n13859) );
  NAND2X0 U14825 ( .IN1(n7729), .IN2(g9743), .QN(n13860) );
  NAND2X0 U14826 ( .IN1(n13861), .IN2(n13862), .QN(g25757) );
  NAND2X0 U14827 ( .IN1(n8510), .IN2(g6727), .QN(n13862) );
  OR2X1 U14828 ( .IN1(n8478), .IN2(n5990), .Q(n13861) );
  NOR2X0 U14829 ( .IN1(n8572), .IN2(n5563), .QN(g25756) );
  NAND2X0 U14830 ( .IN1(n13863), .IN2(n13864), .QN(g25750) );
  NAND2X0 U14831 ( .IN1(n11482), .IN2(g6159), .QN(n13864) );
  NAND2X0 U14832 ( .IN1(n13865), .IN2(g6195), .QN(n13863) );
  NAND3X0 U14833 ( .IN1(n13866), .IN2(n13867), .IN3(n13868), .QN(g25749) );
  OR2X1 U14834 ( .IN1(n13865), .IN2(n5888), .Q(n13868) );
  NAND2X0 U14835 ( .IN1(n13869), .IN2(g6187), .QN(n13867) );
  NAND2X0 U14836 ( .IN1(n13870), .IN2(n8517), .QN(n13869) );
  NAND2X0 U14837 ( .IN1(n11483), .IN2(g6181), .QN(n13870) );
  NAND4X0 U14838 ( .IN1(n11483), .IN2(n8505), .IN3(n5667), .IN4(n5453), .QN(
        n13866) );
  NAND2X0 U14839 ( .IN1(n13871), .IN2(n13872), .QN(g25748) );
  NAND2X0 U14840 ( .IN1(n11482), .IN2(g6187), .QN(n13872) );
  NAND2X0 U14841 ( .IN1(n13865), .IN2(g6181), .QN(n13871) );
  NAND3X0 U14842 ( .IN1(n13873), .IN2(n13874), .IN3(n13875), .QN(g25747) );
  NAND2X0 U14843 ( .IN1(n11482), .IN2(g6167), .QN(n13875) );
  INVX0 U14844 ( .INP(n13865), .ZN(n11482) );
  NAND2X0 U14845 ( .IN1(n10344), .IN2(n8512), .QN(n13865) );
  NAND3X0 U14846 ( .IN1(n5430), .IN2(n11483), .IN3(n8496), .QN(n13874) );
  INVX0 U14847 ( .INP(n10344), .ZN(n11483) );
  NAND2X0 U14848 ( .IN1(n11500), .IN2(g6215), .QN(n10344) );
  INVX0 U14849 ( .INP(n3810), .ZN(n11500) );
  NAND2X0 U14850 ( .IN1(g6227), .IN2(g6219), .QN(n3810) );
  NAND2X0 U14851 ( .IN1(n8605), .IN2(g6163), .QN(n13873) );
  NAND2X0 U14852 ( .IN1(n13876), .IN2(n13877), .QN(g25744) );
  OR2X1 U14853 ( .IN1(n8477), .IN2(n7724), .Q(n13877) );
  NAND3X0 U14854 ( .IN1(n7723), .IN2(n13878), .IN3(n8496), .QN(n13876) );
  NAND2X0 U14855 ( .IN1(n5988), .IN2(n13879), .QN(n13878) );
  NAND2X0 U14856 ( .IN1(test_so92), .IN2(n7724), .QN(n13879) );
  NAND2X0 U14857 ( .IN1(n13880), .IN2(n13881), .QN(g25743) );
  NAND2X0 U14858 ( .IN1(test_so69), .IN2(n8517), .QN(n13881) );
  OR2X1 U14859 ( .IN1(n8477), .IN2(n5988), .Q(n13880) );
  NOR2X0 U14860 ( .IN1(n8571), .IN2(n5568), .QN(g25742) );
  NAND2X0 U14861 ( .IN1(n13882), .IN2(n13883), .QN(g25736) );
  NAND2X0 U14862 ( .IN1(n11563), .IN2(g5813), .QN(n13883) );
  NAND2X0 U14863 ( .IN1(n13884), .IN2(g5849), .QN(n13882) );
  NAND3X0 U14864 ( .IN1(n13885), .IN2(n13886), .IN3(n13887), .QN(g25735) );
  NAND2X0 U14865 ( .IN1(test_so83), .IN2(n11563), .QN(n13887) );
  NAND2X0 U14866 ( .IN1(n13888), .IN2(g5841), .QN(n13886) );
  NAND2X0 U14867 ( .IN1(n13889), .IN2(n8517), .QN(n13888) );
  NAND2X0 U14868 ( .IN1(n11564), .IN2(g5835), .QN(n13889) );
  NAND4X0 U14869 ( .IN1(n11564), .IN2(n8505), .IN3(n5663), .IN4(n5449), .QN(
        n13885) );
  NAND2X0 U14870 ( .IN1(n13890), .IN2(n13891), .QN(g25734) );
  NAND2X0 U14871 ( .IN1(n11563), .IN2(g5841), .QN(n13891) );
  NAND2X0 U14872 ( .IN1(n13884), .IN2(g5835), .QN(n13890) );
  NAND3X0 U14873 ( .IN1(n13892), .IN2(n13893), .IN3(n13894), .QN(g25733) );
  NAND2X0 U14874 ( .IN1(n11563), .IN2(g5821), .QN(n13894) );
  INVX0 U14875 ( .INP(n13884), .ZN(n11563) );
  NAND2X0 U14876 ( .IN1(n10343), .IN2(n8517), .QN(n13884) );
  NAND3X0 U14877 ( .IN1(n5429), .IN2(n11564), .IN3(n8496), .QN(n13893) );
  INVX0 U14878 ( .INP(n10343), .ZN(n11564) );
  NAND2X0 U14879 ( .IN1(n11581), .IN2(g5869), .QN(n10343) );
  INVX0 U14880 ( .INP(n3844), .ZN(n11581) );
  NAND2X0 U14881 ( .IN1(test_so36), .IN2(g5873), .QN(n3844) );
  NAND2X0 U14882 ( .IN1(n8605), .IN2(g5817), .QN(n13892) );
  NAND2X0 U14883 ( .IN1(n13895), .IN2(n13896), .QN(g25730) );
  OR2X1 U14884 ( .IN1(n8477), .IN2(n7740), .Q(n13896) );
  NAND3X0 U14885 ( .IN1(n7739), .IN2(n13897), .IN3(n8497), .QN(n13895) );
  NAND2X0 U14886 ( .IN1(n5996), .IN2(n13898), .QN(n13897) );
  NAND2X0 U14887 ( .IN1(n7740), .IN2(g9617), .QN(n13898) );
  NAND2X0 U14888 ( .IN1(n13899), .IN2(n13900), .QN(g25729) );
  NAND2X0 U14889 ( .IN1(n8511), .IN2(g6035), .QN(n13900) );
  OR2X1 U14890 ( .IN1(n8476), .IN2(n5996), .Q(n13899) );
  NOR2X0 U14891 ( .IN1(n8217), .IN2(n8557), .QN(g25728) );
  NAND2X0 U14892 ( .IN1(n13901), .IN2(n13902), .QN(g25722) );
  NAND2X0 U14893 ( .IN1(n11644), .IN2(g5467), .QN(n13902) );
  NAND2X0 U14894 ( .IN1(n13903), .IN2(g5503), .QN(n13901) );
  NAND3X0 U14895 ( .IN1(n13904), .IN2(n13905), .IN3(n13906), .QN(g25721) );
  OR2X1 U14896 ( .IN1(n13903), .IN2(n5885), .Q(n13906) );
  NAND2X0 U14897 ( .IN1(n13907), .IN2(g5495), .QN(n13905) );
  NAND2X0 U14898 ( .IN1(n13908), .IN2(n8517), .QN(n13907) );
  NAND2X0 U14899 ( .IN1(n10339), .IN2(g5489), .QN(n13908) );
  NAND4X0 U14900 ( .IN1(n10339), .IN2(n8505), .IN3(n5660), .IN4(n5446), .QN(
        n13904) );
  NAND2X0 U14901 ( .IN1(n13909), .IN2(n13910), .QN(g25720) );
  NAND2X0 U14902 ( .IN1(n11644), .IN2(g5495), .QN(n13910) );
  NAND2X0 U14903 ( .IN1(n13903), .IN2(g5489), .QN(n13909) );
  INVX0 U14904 ( .INP(n11644), .ZN(n13903) );
  NAND3X0 U14905 ( .IN1(n13911), .IN2(n13912), .IN3(n13913), .QN(g25719) );
  NAND2X0 U14906 ( .IN1(n11644), .IN2(g5475), .QN(n13913) );
  NOR2X0 U14907 ( .IN1(n10339), .IN2(n8548), .QN(n11644) );
  NAND3X0 U14908 ( .IN1(n5425), .IN2(n10339), .IN3(n8497), .QN(n13912) );
  NOR2X0 U14909 ( .IN1(n3877), .IN2(n5647), .QN(n10339) );
  NAND2X0 U14910 ( .IN1(g5535), .IN2(g5527), .QN(n3877) );
  NAND2X0 U14911 ( .IN1(n8605), .IN2(g5471), .QN(n13911) );
  NAND2X0 U14912 ( .IN1(n13914), .IN2(n13915), .QN(g25716) );
  OR2X1 U14913 ( .IN1(n8476), .IN2(n7733), .Q(n13915) );
  NAND3X0 U14914 ( .IN1(n13916), .IN2(n7732), .IN3(n8497), .QN(n13914) );
  NAND2X0 U14915 ( .IN1(n5992), .IN2(n13917), .QN(n13916) );
  NAND2X0 U14916 ( .IN1(n7733), .IN2(g9555), .QN(n13917) );
  NAND2X0 U14917 ( .IN1(n13918), .IN2(n13919), .QN(g25715) );
  NAND2X0 U14918 ( .IN1(n8511), .IN2(g5689), .QN(n13919) );
  OR2X1 U14919 ( .IN1(n8476), .IN2(n5992), .Q(n13918) );
  NOR2X0 U14920 ( .IN1(n8570), .IN2(n5566), .QN(g25714) );
  NAND2X0 U14921 ( .IN1(n13920), .IN2(n13921), .QN(g25708) );
  NAND2X0 U14922 ( .IN1(n11724), .IN2(g5120), .QN(n13921) );
  NAND2X0 U14923 ( .IN1(n13922), .IN2(g5156), .QN(n13920) );
  NAND3X0 U14924 ( .IN1(n13923), .IN2(n13924), .IN3(n13925), .QN(g25707) );
  OR2X1 U14925 ( .IN1(n13922), .IN2(n5883), .Q(n13925) );
  NAND2X0 U14926 ( .IN1(test_so98), .IN2(n13926), .QN(n13924) );
  NAND2X0 U14927 ( .IN1(n13927), .IN2(n8517), .QN(n13926) );
  NAND2X0 U14928 ( .IN1(g26801), .IN2(g5142), .QN(n13927) );
  NAND4X0 U14929 ( .IN1(g26801), .IN2(n8505), .IN3(n5658), .IN4(n8238), .QN(
        n13923) );
  NAND2X0 U14930 ( .IN1(n13928), .IN2(n13929), .QN(g25706) );
  NAND2X0 U14931 ( .IN1(test_so98), .IN2(n11724), .QN(n13929) );
  NAND2X0 U14932 ( .IN1(n13922), .IN2(g5142), .QN(n13928) );
  INVX0 U14933 ( .INP(n11724), .ZN(n13922) );
  NAND3X0 U14934 ( .IN1(n13930), .IN2(n13931), .IN3(n13932), .QN(g25705) );
  NAND2X0 U14935 ( .IN1(test_so96), .IN2(n11724), .QN(n13932) );
  NOR2X0 U14936 ( .IN1(g26801), .IN2(n8548), .QN(n11724) );
  NAND3X0 U14937 ( .IN1(g26801), .IN2(n8211), .IN3(n8497), .QN(n13931) );
  NOR2X0 U14938 ( .IN1(n3910), .IN2(n5650), .QN(g26801) );
  NAND2X0 U14939 ( .IN1(g5188), .IN2(g5180), .QN(n3910) );
  OR2X1 U14940 ( .IN1(n8476), .IN2(n7709), .Q(n13930) );
  NOR2X0 U14941 ( .IN1(n7781), .IN2(n13933), .QN(g25704) );
  NOR2X0 U14942 ( .IN1(n8570), .IN2(g5069), .QN(n13933) );
  NAND2X0 U14943 ( .IN1(n13934), .IN2(n13935), .QN(g25703) );
  NAND2X0 U14944 ( .IN1(n8606), .IN2(g5112), .QN(n13935) );
  NAND3X0 U14945 ( .IN1(n5689), .IN2(n13936), .IN3(n8497), .QN(n13934) );
  NAND2X0 U14946 ( .IN1(n7871), .IN2(n13937), .QN(n13936) );
  OR2X1 U14947 ( .IN1(g5112), .IN2(n5690), .Q(n13937) );
  NAND2X0 U14948 ( .IN1(n13938), .IN2(n13939), .QN(g25702) );
  NAND2X0 U14949 ( .IN1(test_so32), .IN2(n8535), .QN(n13939) );
  NAND3X0 U14950 ( .IN1(n5690), .IN2(n13940), .IN3(n8497), .QN(n13938) );
  NAND2X0 U14951 ( .IN1(n7842), .IN2(n13941), .QN(n13940) );
  OR2X1 U14952 ( .IN1(n5689), .IN2(test_so32), .Q(n13941) );
  NAND2X0 U14953 ( .IN1(n13942), .IN2(n13943), .QN(g25701) );
  NAND2X0 U14954 ( .IN1(test_so10), .IN2(n8516), .QN(n13943) );
  NAND2X0 U14955 ( .IN1(n8606), .IN2(g5062), .QN(n13942) );
  NOR2X0 U14956 ( .IN1(n8569), .IN2(n5567), .QN(g25700) );
  NAND3X0 U14957 ( .IN1(n13944), .IN2(n13945), .IN3(n13946), .QN(g25699) );
  OR2X1 U14958 ( .IN1(n8476), .IN2(n5753), .Q(n13946) );
  OR3X1 U14959 ( .IN1(n8531), .IN2(n5014), .IN3(n5669), .Q(n13945) );
  NAND2X0 U14960 ( .IN1(n5014), .IN2(n5669), .QN(n13944) );
  NAND3X0 U14961 ( .IN1(n13947), .IN2(n13948), .IN3(n13949), .QN(g25698) );
  NAND2X0 U14962 ( .IN1(n8606), .IN2(g5092), .QN(n13949) );
  OR3X1 U14963 ( .IN1(n8530), .IN2(n5016), .IN3(n5753), .Q(n13948) );
  NAND2X0 U14964 ( .IN1(n5016), .IN2(n5753), .QN(n13947) );
  XOR2X1 U14965 ( .IN1(n13950), .IN2(n5681), .Q(g25697) );
  NAND2X0 U14966 ( .IN1(n8512), .IN2(g5092), .QN(n13950) );
  NAND3X0 U14967 ( .IN1(n13951), .IN2(n13952), .IN3(n13953), .QN(g25696) );
  NAND3X0 U14968 ( .IN1(n8502), .IN2(g5077), .IN3(n7781), .QN(n13953) );
  OR2X1 U14969 ( .IN1(n13954), .IN2(n5893), .Q(n13952) );
  NAND3X0 U14970 ( .IN1(n13954), .IN2(n13955), .IN3(n5893), .QN(n13951) );
  NAND2X0 U14971 ( .IN1(n7780), .IN2(g5077), .QN(n13955) );
  NOR2X0 U14972 ( .IN1(g5084), .IN2(n8552), .QN(n13954) );
  NOR2X0 U14973 ( .IN1(n5455), .IN2(n13956), .QN(g25695) );
  AND3X1 U14974 ( .IN1(n13957), .IN2(n13958), .IN3(n8528), .Q(n13956) );
  NAND2X0 U14975 ( .IN1(n7780), .IN2(g5084), .QN(n13958) );
  NAND2X0 U14976 ( .IN1(n7781), .IN2(n5681), .QN(n13957) );
  NAND2X0 U14977 ( .IN1(n13959), .IN2(n13960), .QN(g25691) );
  NAND2X0 U14978 ( .IN1(n616), .IN2(n13961), .QN(n13960) );
  NAND4X0 U14979 ( .IN1(n5416), .IN2(test_so11), .IN3(n5711), .IN4(n13962), 
        .QN(n13961) );
  AND4X1 U14980 ( .IN1(g4098), .IN2(n10340), .IN3(n5612), .IN4(n7826), .Q(
        n13962) );
  NOR2X0 U14981 ( .IN1(g4093), .IN2(n5480), .QN(n10340) );
  INVX0 U14982 ( .INP(n10984), .ZN(n616) );
  NAND2X0 U14983 ( .IN1(n8606), .IN2(g4125), .QN(n13959) );
  NAND2X0 U14984 ( .IN1(n13963), .IN2(n13964), .QN(g25690) );
  NAND2X0 U14985 ( .IN1(n8607), .IN2(g4169), .QN(n13964) );
  NAND3X0 U14986 ( .IN1(n8122), .IN2(g25689), .IN3(n8498), .QN(n13963) );
  NAND3X0 U14987 ( .IN1(n13965), .IN2(n13966), .IN3(n13967), .QN(g25687) );
  NAND2X0 U14988 ( .IN1(n8596), .IN2(g4057), .QN(n13967) );
  NAND3X0 U14989 ( .IN1(n13968), .IN2(g4169), .IN3(n5612), .QN(n13966) );
  INVX0 U14990 ( .INP(n4723), .ZN(n13968) );
  NAND2X0 U14991 ( .IN1(g4057), .IN2(g4064), .QN(n4723) );
  NAND2X0 U14992 ( .IN1(n5026), .IN2(n11816), .QN(n13965) );
  NAND2X0 U14993 ( .IN1(n13969), .IN2(n13970), .QN(g25686) );
  NAND2X0 U14994 ( .IN1(n13971), .IN2(g4064), .QN(n13970) );
  NAND2X0 U14995 ( .IN1(n13972), .IN2(n8516), .QN(n13971) );
  NAND2X0 U14996 ( .IN1(n5711), .IN2(g4169), .QN(n13972) );
  NAND3X0 U14997 ( .IN1(n11816), .IN2(g4057), .IN3(n5416), .QN(n13969) );
  NOR2X0 U14998 ( .IN1(n8569), .IN2(n5729), .QN(n11816) );
  NAND3X0 U14999 ( .IN1(n13973), .IN2(n13974), .IN3(n10984), .QN(g25685) );
  NAND2X0 U15000 ( .IN1(n5729), .IN2(n8516), .QN(n10984) );
  NAND2X0 U15001 ( .IN1(n5416), .IN2(n8516), .QN(n13974) );
  OR2X1 U15002 ( .IN1(n8478), .IN2(n8181), .Q(n13973) );
  NAND2X0 U15003 ( .IN1(n13975), .IN2(n13976), .QN(g25684) );
  NAND2X0 U15004 ( .IN1(n11820), .IN2(g3813), .QN(n13976) );
  NAND2X0 U15005 ( .IN1(n13977), .IN2(g3849), .QN(n13975) );
  NAND3X0 U15006 ( .IN1(n13978), .IN2(n13979), .IN3(n13980), .QN(g25683) );
  OR2X1 U15007 ( .IN1(n13977), .IN2(n5886), .Q(n13980) );
  NAND2X0 U15008 ( .IN1(test_so97), .IN2(n13981), .QN(n13979) );
  NAND2X0 U15009 ( .IN1(n13982), .IN2(n8514), .QN(n13981) );
  NAND2X0 U15010 ( .IN1(n11821), .IN2(g3835), .QN(n13982) );
  OR4X1 U15011 ( .IN1(n10353), .IN2(n8544), .IN3(g3835), .IN4(test_so97), .Q(
        n13978) );
  NAND2X0 U15012 ( .IN1(n13983), .IN2(n13984), .QN(g25682) );
  NAND2X0 U15013 ( .IN1(test_so97), .IN2(n11820), .QN(n13984) );
  NAND2X0 U15014 ( .IN1(n13977), .IN2(g3835), .QN(n13983) );
  NAND3X0 U15015 ( .IN1(n13985), .IN2(n13986), .IN3(n13987), .QN(g25681) );
  NAND2X0 U15016 ( .IN1(n11820), .IN2(g3821), .QN(n13987) );
  INVX0 U15017 ( .INP(n13977), .ZN(n11820) );
  NAND2X0 U15018 ( .IN1(n10353), .IN2(n8513), .QN(n13977) );
  NAND3X0 U15019 ( .IN1(n5428), .IN2(n11821), .IN3(n8490), .QN(n13986) );
  INVX0 U15020 ( .INP(n10353), .ZN(n11821) );
  NAND2X0 U15021 ( .IN1(test_so33), .IN2(n11838), .QN(n10353) );
  INVX0 U15022 ( .INP(n3953), .ZN(n11838) );
  NAND2X0 U15023 ( .IN1(g3881), .IN2(g3873), .QN(n3953) );
  OR2X1 U15024 ( .IN1(n8479), .IN2(n7710), .Q(n13985) );
  NAND2X0 U15025 ( .IN1(n13988), .IN2(n13989), .QN(g25678) );
  OR2X1 U15026 ( .IN1(n8479), .IN2(n7735), .Q(n13989) );
  NAND3X0 U15027 ( .IN1(n7734), .IN2(n13990), .IN3(n8490), .QN(n13988) );
  NAND2X0 U15028 ( .IN1(n5994), .IN2(n13991), .QN(n13990) );
  NAND2X0 U15029 ( .IN1(n7735), .IN2(g8344), .QN(n13991) );
  NAND2X0 U15030 ( .IN1(n13992), .IN2(n13993), .QN(g25677) );
  NAND2X0 U15031 ( .IN1(n8511), .IN2(g4040), .QN(n13993) );
  OR2X1 U15032 ( .IN1(n8478), .IN2(n5994), .Q(n13992) );
  NOR2X0 U15033 ( .IN1(n8570), .IN2(n5564), .QN(g25676) );
  NAND2X0 U15034 ( .IN1(n13994), .IN2(n13995), .QN(g25670) );
  NAND2X0 U15035 ( .IN1(n11902), .IN2(g3462), .QN(n13995) );
  NAND2X0 U15036 ( .IN1(n13996), .IN2(g3498), .QN(n13994) );
  NAND3X0 U15037 ( .IN1(n13997), .IN2(n13998), .IN3(n13999), .QN(g25669) );
  OR2X1 U15038 ( .IN1(n13996), .IN2(n5889), .Q(n13999) );
  NAND2X0 U15039 ( .IN1(n14000), .IN2(g3490), .QN(n13998) );
  NAND2X0 U15040 ( .IN1(n14001), .IN2(n8513), .QN(n14000) );
  NAND2X0 U15041 ( .IN1(n11903), .IN2(g3484), .QN(n14001) );
  NAND4X0 U15042 ( .IN1(n11903), .IN2(n8505), .IN3(n5668), .IN4(n5454), .QN(
        n13997) );
  NAND2X0 U15043 ( .IN1(n14002), .IN2(n14003), .QN(g25668) );
  NAND2X0 U15044 ( .IN1(n11902), .IN2(g3490), .QN(n14003) );
  NAND2X0 U15045 ( .IN1(n13996), .IN2(g3484), .QN(n14002) );
  NAND3X0 U15046 ( .IN1(n14004), .IN2(n14005), .IN3(n14006), .QN(g25667) );
  NAND2X0 U15047 ( .IN1(n11902), .IN2(g3470), .QN(n14006) );
  INVX0 U15048 ( .INP(n13996), .ZN(n11902) );
  NAND2X0 U15049 ( .IN1(n10352), .IN2(n8513), .QN(n13996) );
  NAND3X0 U15050 ( .IN1(n5424), .IN2(n11903), .IN3(n8489), .QN(n14005) );
  INVX0 U15051 ( .INP(n10352), .ZN(n11903) );
  NAND2X0 U15052 ( .IN1(n11920), .IN2(g3518), .QN(n10352) );
  INVX0 U15053 ( .INP(n3986), .ZN(n11920) );
  NAND2X0 U15054 ( .IN1(g3530), .IN2(g3522), .QN(n3986) );
  NAND2X0 U15055 ( .IN1(n8607), .IN2(g3466), .QN(n14004) );
  NAND2X0 U15056 ( .IN1(n14007), .IN2(n14008), .QN(g25664) );
  OR2X1 U15057 ( .IN1(n8477), .IN2(n7713), .Q(n14008) );
  NAND3X0 U15058 ( .IN1(n7712), .IN2(n14009), .IN3(n8489), .QN(n14007) );
  NAND2X0 U15059 ( .IN1(n5986), .IN2(n14010), .QN(n14009) );
  NAND2X0 U15060 ( .IN1(n7713), .IN2(g8279), .QN(n14010) );
  NAND2X0 U15061 ( .IN1(n14011), .IN2(n14012), .QN(g25663) );
  NAND2X0 U15062 ( .IN1(n8512), .IN2(g3689), .QN(n14012) );
  OR2X1 U15063 ( .IN1(n8477), .IN2(n5986), .Q(n14011) );
  NOR2X0 U15064 ( .IN1(n8570), .IN2(n5569), .QN(g25662) );
  NAND2X0 U15065 ( .IN1(n14013), .IN2(n14014), .QN(g25656) );
  NAND2X0 U15066 ( .IN1(n11983), .IN2(g3111), .QN(n14014) );
  NAND2X0 U15067 ( .IN1(n14015), .IN2(g3147), .QN(n14013) );
  NAND3X0 U15068 ( .IN1(n14016), .IN2(n14017), .IN3(n14018), .QN(g25655) );
  OR2X1 U15069 ( .IN1(n14015), .IN2(n5882), .Q(n14018) );
  NAND2X0 U15070 ( .IN1(n14019), .IN2(g3139), .QN(n14017) );
  NAND2X0 U15071 ( .IN1(n14020), .IN2(n8513), .QN(n14019) );
  NAND2X0 U15072 ( .IN1(n10349), .IN2(g3133), .QN(n14020) );
  NAND4X0 U15073 ( .IN1(n10349), .IN2(n8505), .IN3(n5661), .IN4(n5447), .QN(
        n14016) );
  NAND2X0 U15074 ( .IN1(n14021), .IN2(n14022), .QN(g25654) );
  NAND2X0 U15075 ( .IN1(n11983), .IN2(g3139), .QN(n14022) );
  NAND2X0 U15076 ( .IN1(n14015), .IN2(g3133), .QN(n14021) );
  INVX0 U15077 ( .INP(n11983), .ZN(n14015) );
  NAND3X0 U15078 ( .IN1(n14023), .IN2(n14024), .IN3(n14025), .QN(g25653) );
  NAND2X0 U15079 ( .IN1(n11983), .IN2(g3119), .QN(n14025) );
  NOR2X0 U15080 ( .IN1(n10349), .IN2(n8550), .QN(n11983) );
  NAND3X0 U15081 ( .IN1(n5423), .IN2(n10349), .IN3(n8489), .QN(n14024) );
  NOR2X0 U15082 ( .IN1(n4017), .IN2(n5652), .QN(n10349) );
  NAND2X0 U15083 ( .IN1(g3171), .IN2(g3179), .QN(n4017) );
  NAND2X0 U15084 ( .IN1(n8607), .IN2(g3115), .QN(n14023) );
  NAND2X0 U15085 ( .IN1(n14026), .IN2(n14027), .QN(g25650) );
  OR2X1 U15086 ( .IN1(n8476), .IN2(n7743), .Q(n14027) );
  NAND3X0 U15087 ( .IN1(n7742), .IN2(n14028), .IN3(n8488), .QN(n14026) );
  NAND2X0 U15088 ( .IN1(n5998), .IN2(n14029), .QN(n14028) );
  NAND2X0 U15089 ( .IN1(n7743), .IN2(g8215), .QN(n14029) );
  NAND2X0 U15090 ( .IN1(n14030), .IN2(n14031), .QN(g25649) );
  NAND2X0 U15091 ( .IN1(n8512), .IN2(g3338), .QN(n14031) );
  OR2X1 U15092 ( .IN1(n8476), .IN2(n5998), .Q(n14030) );
  NOR2X0 U15093 ( .IN1(n8571), .IN2(n5390), .QN(g25648) );
  OR3X1 U15094 ( .IN1(n14032), .IN2(n14033), .IN3(n5045), .Q(g25639) );
  NOR2X0 U15095 ( .IN1(n8571), .IN2(n12076), .QN(n14033) );
  NAND2X0 U15096 ( .IN1(n5299), .IN2(g2719), .QN(n12076) );
  NOR2X0 U15097 ( .IN1(n5299), .IN2(n8504), .QN(n14032) );
  NAND2X0 U15098 ( .IN1(n14034), .IN2(n14035), .QN(g25638) );
  NAND2X0 U15099 ( .IN1(n8607), .IN2(g1564), .QN(n14035) );
  NAND2X0 U15100 ( .IN1(n14036), .IN2(n8514), .QN(n14034) );
  NAND2X0 U15101 ( .IN1(n14037), .IN2(n14038), .QN(n14036) );
  NAND2X0 U15102 ( .IN1(n14039), .IN2(g1559), .QN(n14038) );
  NAND3X0 U15103 ( .IN1(n14040), .IN2(n5768), .IN3(n5441), .QN(n14037) );
  NAND2X0 U15104 ( .IN1(n14041), .IN2(n14042), .QN(g25637) );
  NAND3X0 U15105 ( .IN1(n8504), .IN2(g1554), .IN3(n14039), .QN(n14042) );
  NAND2X0 U15106 ( .IN1(n14043), .IN2(g1559), .QN(n14041) );
  NAND2X0 U15107 ( .IN1(n14044), .IN2(n8514), .QN(n14043) );
  NAND2X0 U15108 ( .IN1(n14040), .IN2(n5768), .QN(n14044) );
  NAND2X0 U15109 ( .IN1(n14045), .IN2(n14046), .QN(g25636) );
  NAND2X0 U15110 ( .IN1(n8607), .IN2(g1521), .QN(n14046) );
  NAND2X0 U15111 ( .IN1(n14047), .IN2(n8514), .QN(n14045) );
  NAND2X0 U15112 ( .IN1(n14048), .IN2(n14049), .QN(n14047) );
  NAND2X0 U15113 ( .IN1(n10561), .IN2(n12356), .QN(n14049) );
  INVX0 U15114 ( .INP(n14050), .ZN(n12356) );
  NAND2X0 U15115 ( .IN1(n14051), .IN2(g1306), .QN(n14048) );
  NAND2X0 U15116 ( .IN1(n10561), .IN2(g7946), .QN(n14051) );
  NOR2X0 U15117 ( .IN1(n8206), .IN2(n5364), .QN(n10561) );
  NAND2X0 U15118 ( .IN1(n14052), .IN2(n14053), .QN(g25635) );
  NAND2X0 U15119 ( .IN1(n14054), .IN2(g1484), .QN(n14053) );
  NAND2X0 U15120 ( .IN1(n14055), .IN2(n8514), .QN(n14054) );
  NAND3X0 U15121 ( .IN1(n5483), .IN2(n12837), .IN3(n13677), .QN(n14055) );
  NAND2X0 U15122 ( .IN1(n14056), .IN2(g1300), .QN(n14052) );
  NAND2X0 U15123 ( .IN1(n14057), .IN2(n14058), .QN(n14056) );
  NAND2X0 U15124 ( .IN1(n14059), .IN2(n8514), .QN(n14058) );
  NAND2X0 U15125 ( .IN1(n13677), .IN2(g1484), .QN(n14059) );
  NOR2X0 U15126 ( .IN1(n8137), .IN2(test_so12), .QN(n13677) );
  NOR3X0 U15127 ( .IN1(n14060), .IN2(test_so68), .IN3(n13689), .QN(g25634) );
  NOR3X0 U15128 ( .IN1(n5655), .IN2(n8054), .IN3(n14061), .QN(n13689) );
  NOR2X0 U15129 ( .IN1(n14062), .IN2(n14063), .QN(n14060) );
  NOR2X0 U15130 ( .IN1(n8054), .IN2(n8556), .QN(n14063) );
  NOR2X0 U15131 ( .IN1(n14061), .IN2(n10807), .QN(n14062) );
  NAND3X0 U15132 ( .IN1(n14064), .IN2(n14065), .IN3(n14066), .QN(g25633) );
  NAND3X0 U15133 ( .IN1(n13694), .IN2(n7693), .IN3(n13693), .QN(n14066) );
  NAND3X0 U15134 ( .IN1(n14067), .IN2(g1384), .IN3(n8486), .QN(n14065) );
  NAND2X0 U15135 ( .IN1(n8608), .IN2(g1379), .QN(n14064) );
  NAND2X0 U15136 ( .IN1(n14068), .IN2(n14069), .QN(g25632) );
  NAND2X0 U15137 ( .IN1(n13693), .IN2(n14070), .QN(n14069) );
  NAND2X0 U15138 ( .IN1(n12360), .IN2(n14071), .QN(n14070) );
  NAND2X0 U15139 ( .IN1(n13443), .IN2(n13438), .QN(n14071) );
  INVX0 U15140 ( .INP(n14072), .ZN(n13438) );
  NOR2X0 U15141 ( .IN1(n8571), .IN2(n5322), .QN(n13693) );
  NAND2X0 U15142 ( .IN1(n14073), .IN2(g1312), .QN(n14068) );
  NAND2X0 U15143 ( .IN1(n14067), .IN2(n8514), .QN(n14073) );
  INVX0 U15144 ( .INP(n13694), .ZN(n14067) );
  NOR2X0 U15145 ( .IN1(n8572), .IN2(n14074), .QN(g25631) );
  NOR2X0 U15146 ( .IN1(n14075), .IN2(n14076), .QN(n14074) );
  NOR2X0 U15147 ( .IN1(n5466), .IN2(n13694), .QN(n14076) );
  NOR3X0 U15148 ( .IN1(n13444), .IN2(n14077), .IN3(n14078), .QN(n14075) );
  NOR2X0 U15149 ( .IN1(n5322), .IN2(n14079), .QN(n14078) );
  NOR2X0 U15150 ( .IN1(n14072), .IN2(n13443), .QN(n14079) );
  NAND2X0 U15151 ( .IN1(g1373), .IN2(g1361), .QN(n13443) );
  NOR2X0 U15152 ( .IN1(n13441), .IN2(n7845), .QN(n14072) );
  AND2X1 U15153 ( .IN1(n4896), .IN2(n5322), .Q(n14077) );
  NAND4X0 U15154 ( .IN1(n13441), .IN2(g1379), .IN3(g1367), .IN4(g1345), .QN(
        n4896) );
  NAND2X0 U15155 ( .IN1(n14080), .IN2(n14081), .QN(g25630) );
  NAND2X0 U15156 ( .IN1(n14082), .IN2(g1249), .QN(n14081) );
  NAND2X0 U15157 ( .IN1(n14083), .IN2(n8514), .QN(n14082) );
  NAND2X0 U15158 ( .IN1(n7830), .IN2(g12923), .QN(n14083) );
  NAND2X0 U15159 ( .IN1(g24247), .IN2(g1266), .QN(n14080) );
  NAND2X0 U15160 ( .IN1(n14084), .IN2(n14085), .QN(g25629) );
  NAND2X0 U15161 ( .IN1(n8608), .IN2(g1221), .QN(n14085) );
  NAND2X0 U15162 ( .IN1(n14086), .IN2(n8514), .QN(n14084) );
  NAND2X0 U15163 ( .IN1(n14087), .IN2(n14088), .QN(n14086) );
  NAND2X0 U15164 ( .IN1(n14089), .IN2(g1216), .QN(n14088) );
  NAND3X0 U15165 ( .IN1(n14090), .IN2(n8212), .IN3(n5442), .QN(n14087) );
  NAND2X0 U15166 ( .IN1(n14091), .IN2(n14092), .QN(g25628) );
  NAND3X0 U15167 ( .IN1(n14089), .IN2(n8482), .IN3(test_so76), .QN(n14092) );
  NAND2X0 U15168 ( .IN1(n14093), .IN2(g1216), .QN(n14091) );
  NAND2X0 U15169 ( .IN1(n14094), .IN2(n8514), .QN(n14093) );
  NAND2X0 U15170 ( .IN1(n14090), .IN2(n8212), .QN(n14094) );
  INVX0 U15171 ( .INP(n14089), .ZN(n14090) );
  NAND2X0 U15172 ( .IN1(n14095), .IN2(n14096), .QN(g25627) );
  NAND2X0 U15173 ( .IN1(n8608), .IN2(g1178), .QN(n14096) );
  NAND2X0 U15174 ( .IN1(n14097), .IN2(n8514), .QN(n14095) );
  NAND2X0 U15175 ( .IN1(n14098), .IN2(n14099), .QN(n14097) );
  NAND2X0 U15176 ( .IN1(n10718), .IN2(n12387), .QN(n14099) );
  INVX0 U15177 ( .INP(n14100), .ZN(n12387) );
  NAND2X0 U15178 ( .IN1(n14101), .IN2(g962), .QN(n14098) );
  NAND2X0 U15179 ( .IN1(n10718), .IN2(g7916), .QN(n14101) );
  NOR2X0 U15180 ( .IN1(n5599), .IN2(n5363), .QN(n10718) );
  NAND2X0 U15181 ( .IN1(n14102), .IN2(n14103), .QN(g25626) );
  NAND2X0 U15182 ( .IN1(n14104), .IN2(g1141), .QN(n14103) );
  NAND2X0 U15183 ( .IN1(n14105), .IN2(n8514), .QN(n14104) );
  NAND3X0 U15184 ( .IN1(n5341), .IN2(n12869), .IN3(n13708), .QN(n14105) );
  NAND2X0 U15185 ( .IN1(n14106), .IN2(g956), .QN(n14102) );
  NAND2X0 U15186 ( .IN1(n14107), .IN2(n14108), .QN(n14106) );
  NAND2X0 U15187 ( .IN1(n14109), .IN2(n8515), .QN(n14108) );
  NAND2X0 U15188 ( .IN1(n13708), .IN2(g1141), .QN(n14109) );
  NOR2X0 U15189 ( .IN1(g1152), .IN2(n8207), .QN(n13708) );
  NOR3X0 U15190 ( .IN1(g979), .IN2(n13720), .IN3(n14110), .QN(g25625) );
  NOR2X0 U15191 ( .IN1(n14111), .IN2(n14112), .QN(n14110) );
  NOR2X0 U15192 ( .IN1(n8055), .IN2(n8554), .QN(n14112) );
  NOR2X0 U15193 ( .IN1(n14113), .IN2(n10820), .QN(n14111) );
  NOR3X0 U15194 ( .IN1(n5654), .IN2(n8055), .IN3(n14113), .QN(n13720) );
  NAND3X0 U15195 ( .IN1(n14114), .IN2(n14115), .IN3(n14116), .QN(g25624) );
  NAND3X0 U15196 ( .IN1(n13725), .IN2(n7692), .IN3(n13724), .QN(n14116) );
  NAND3X0 U15197 ( .IN1(n14117), .IN2(g1041), .IN3(n8485), .QN(n14115) );
  NAND2X0 U15198 ( .IN1(n8608), .IN2(g1036), .QN(n14114) );
  NAND2X0 U15199 ( .IN1(n14118), .IN2(n14119), .QN(g25623) );
  NAND2X0 U15200 ( .IN1(n13724), .IN2(n14120), .QN(n14119) );
  NAND2X0 U15201 ( .IN1(n12391), .IN2(n14121), .QN(n14120) );
  NAND2X0 U15202 ( .IN1(n14122), .IN2(n13451), .QN(n14121) );
  NOR2X0 U15203 ( .IN1(n8572), .IN2(n5321), .QN(n13724) );
  NAND2X0 U15204 ( .IN1(test_so20), .IN2(n14123), .QN(n14118) );
  NAND2X0 U15205 ( .IN1(n14117), .IN2(n8515), .QN(n14123) );
  NOR2X0 U15206 ( .IN1(n8573), .IN2(n14124), .QN(g25622) );
  NOR2X0 U15207 ( .IN1(n14125), .IN2(n14126), .QN(n14124) );
  NOR2X0 U15208 ( .IN1(n13725), .IN2(n8223), .QN(n14126) );
  AND3X1 U15209 ( .IN1(n14127), .IN2(n14128), .IN3(n12391), .Q(n14125) );
  NAND2X0 U15210 ( .IN1(n5321), .IN2(n4921), .QN(n14128) );
  NAND4X0 U15211 ( .IN1(n13455), .IN2(g1036), .IN3(g1024), .IN4(g1002), .QN(
        n4921) );
  INVX0 U15212 ( .INP(n13456), .ZN(n13455) );
  NAND2X0 U15213 ( .IN1(n14129), .IN2(g1008), .QN(n14127) );
  NAND2X0 U15214 ( .IN1(n13454), .IN2(n13451), .QN(n14129) );
  NAND2X0 U15215 ( .IN1(n13456), .IN2(g1046), .QN(n13451) );
  INVX0 U15216 ( .INP(n14122), .ZN(n13454) );
  NAND2X0 U15217 ( .IN1(g1030), .IN2(g1018), .QN(n14122) );
  NAND2X0 U15218 ( .IN1(n14130), .IN2(n14131), .QN(g25621) );
  NAND2X0 U15219 ( .IN1(n14132), .IN2(g904), .QN(n14131) );
  NAND2X0 U15220 ( .IN1(n14133), .IN2(n8515), .QN(n14132) );
  NAND2X0 U15221 ( .IN1(n7827), .IN2(g12919), .QN(n14133) );
  NAND2X0 U15222 ( .IN1(g24231), .IN2(g921), .QN(n14130) );
  NOR2X0 U15223 ( .IN1(n5562), .IN2(n14134), .QN(g25619) );
  NOR2X0 U15224 ( .IN1(n8573), .IN2(n14135), .QN(n14134) );
  XOR2X1 U15225 ( .IN1(n13773), .IN2(g843), .Q(n14135) );
  NAND2X0 U15226 ( .IN1(n14136), .IN2(n14137), .QN(g25618) );
  NAND2X0 U15227 ( .IN1(n14138), .IN2(g817), .QN(n14137) );
  NAND2X0 U15228 ( .IN1(n14139), .IN2(n8515), .QN(n14138) );
  NAND3X0 U15229 ( .IN1(n4948), .IN2(n12888), .IN3(n8153), .QN(n14139) );
  NAND2X0 U15230 ( .IN1(n14140), .IN2(g832), .QN(n14136) );
  NAND2X0 U15231 ( .IN1(n14141), .IN2(n14142), .QN(n14140) );
  NAND2X0 U15232 ( .IN1(n12923), .IN2(n12888), .QN(n14142) );
  NAND2X0 U15233 ( .IN1(n5822), .IN2(n4518), .QN(n14141) );
  AND2X1 U15234 ( .IN1(n12888), .IN2(n8508), .Q(n4518) );
  NAND2X0 U15235 ( .IN1(n14143), .IN2(n14144), .QN(g25617) );
  NAND3X0 U15236 ( .IN1(n14145), .IN2(n14146), .IN3(n12888), .QN(n14144) );
  NAND2X0 U15237 ( .IN1(g847), .IN2(n14147), .QN(n12888) );
  NAND2X0 U15238 ( .IN1(n5733), .IN2(g837), .QN(n14147) );
  NAND2X0 U15239 ( .IN1(n5822), .IN2(n14148), .QN(n14146) );
  NAND2X0 U15240 ( .IN1(n14149), .IN2(g817), .QN(n14145) );
  NAND2X0 U15241 ( .IN1(n8608), .IN2(g812), .QN(n14143) );
  NOR2X0 U15242 ( .IN1(n8572), .IN2(n14150), .QN(g25616) );
  XOR3X1 U15243 ( .IN1(n14151), .IN2(n14152), .IN3(n14153), .Q(n14150) );
  XOR2X1 U15244 ( .IN1(n14154), .IN2(n5597), .Q(n14153) );
  OR2X1 U15245 ( .IN1(n5732), .IN2(n13516), .Q(n14154) );
  AND4X1 U15246 ( .IN1(n5327), .IN2(n8221), .IN3(n13498), .IN4(n14155), .Q(
        n13516) );
  AND3X1 U15247 ( .IN1(n5708), .IN2(n5287), .IN3(n5820), .Q(n14155) );
  XOR2X1 U15248 ( .IN1(g255), .IN2(n6008), .Q(n14152) );
  XOR3X1 U15249 ( .IN1(n7870), .IN2(n7869), .IN3(n14156), .Q(n14151) );
  XOR2X1 U15250 ( .IN1(n7997), .IN2(n7996), .Q(n14156) );
  NAND2X0 U15251 ( .IN1(n14157), .IN2(n14158), .QN(g25615) );
  NAND2X0 U15252 ( .IN1(n14159), .IN2(g667), .QN(n14158) );
  NAND2X0 U15253 ( .IN1(n13486), .IN2(g686), .QN(n14157) );
  NAND3X0 U15254 ( .IN1(n14160), .IN2(n14161), .IN3(n14162), .QN(g25614) );
  NAND2X0 U15255 ( .IN1(n8609), .IN2(g691), .QN(n14162) );
  NAND2X0 U15256 ( .IN1(n14159), .IN2(g686), .QN(n14161) );
  NAND2X0 U15257 ( .IN1(n5111), .IN2(n14163), .QN(n14160) );
  NAND2X0 U15258 ( .IN1(n14164), .IN2(n14165), .QN(g25613) );
  NAND2X0 U15259 ( .IN1(n8609), .IN2(g559), .QN(n14165) );
  NAND3X0 U15260 ( .IN1(n2421), .IN2(n14166), .IN3(n14167), .QN(n14164) );
  XOR2X1 U15261 ( .IN1(n13787), .IN2(g562), .Q(n14167) );
  AND2X1 U15262 ( .IN1(n14168), .IN2(g29211), .Q(n13787) );
  NAND2X0 U15263 ( .IN1(n7672), .IN2(g12368), .QN(n14168) );
  NAND2X0 U15264 ( .IN1(g626), .IN2(n9340), .QN(n14166) );
  NAND2X0 U15265 ( .IN1(n14169), .IN2(n14170), .QN(g25612) );
  NAND2X0 U15266 ( .IN1(n14171), .IN2(g513), .QN(n14170) );
  NAND2X0 U15267 ( .IN1(n14159), .IN2(g518), .QN(n14169) );
  NAND2X0 U15268 ( .IN1(n14172), .IN2(n14173), .QN(g25611) );
  NAND2X0 U15269 ( .IN1(n14171), .IN2(g504), .QN(n14173) );
  NAND2X0 U15270 ( .IN1(n14174), .IN2(n8515), .QN(n14171) );
  NAND2X0 U15271 ( .IN1(n14163), .IN2(n12917), .QN(n14174) );
  INVX0 U15272 ( .INP(n4962), .ZN(n12917) );
  INVX0 U15273 ( .INP(n13793), .ZN(n14163) );
  NAND2X0 U15274 ( .IN1(n14159), .IN2(g513), .QN(n14172) );
  NAND3X0 U15275 ( .IN1(n14175), .IN2(n14176), .IN3(n14177), .QN(g25610) );
  NAND2X0 U15276 ( .IN1(n14159), .IN2(g504), .QN(n14176) );
  INVX0 U15277 ( .INP(n13486), .ZN(n14159) );
  NAND2X0 U15278 ( .IN1(test_so54), .IN2(n13486), .QN(n14175) );
  NAND3X0 U15279 ( .IN1(n14178), .IN2(n14177), .IN3(n14179), .QN(g25609) );
  NAND2X0 U15280 ( .IN1(n13488), .IN2(n5287), .QN(n14179) );
  NAND2X0 U15281 ( .IN1(n4962), .IN2(n13488), .QN(n14177) );
  NOR2X0 U15282 ( .IN1(n13793), .IN2(n8553), .QN(n13488) );
  NAND2X0 U15283 ( .IN1(test_so54), .IN2(n14180), .QN(n14178) );
  NAND2X0 U15284 ( .IN1(n13486), .IN2(n14181), .QN(n14180) );
  NAND2X0 U15285 ( .IN1(n5548), .IN2(n8515), .QN(n14181) );
  NAND2X0 U15286 ( .IN1(n13793), .IN2(n8515), .QN(n13486) );
  NAND3X0 U15287 ( .IN1(g385), .IN2(g358), .IN3(n5633), .QN(n13793) );
  NAND3X0 U15288 ( .IN1(n14182), .IN2(n14183), .IN3(n14184), .QN(g25605) );
  NAND2X0 U15289 ( .IN1(n14185), .IN2(g460), .QN(n14184) );
  NAND2X0 U15290 ( .IN1(n8610), .IN2(g168), .QN(n14183) );
  NAND3X0 U15291 ( .IN1(n13498), .IN2(g246), .IN3(n8502), .QN(n14182) );
  NAND2X0 U15292 ( .IN1(n14186), .IN2(n14187), .QN(g25604) );
  OR2X1 U15293 ( .IN1(n14188), .IN2(n8002), .Q(n14187) );
  NAND2X0 U15294 ( .IN1(n14188), .IN2(g460), .QN(n14186) );
  NAND3X0 U15295 ( .IN1(n14189), .IN2(n14190), .IN3(n14191), .QN(g25602) );
  NAND2X0 U15296 ( .IN1(n14185), .IN2(test_so72), .QN(n14191) );
  NAND2X0 U15297 ( .IN1(n8610), .IN2(g405), .QN(n14190) );
  NAND3X0 U15298 ( .IN1(n13498), .IN2(g446), .IN3(n8502), .QN(n14189) );
  NAND2X0 U15299 ( .IN1(n14192), .IN2(n14193), .QN(g25601) );
  NAND2X0 U15300 ( .IN1(n14185), .IN2(g174), .QN(n14193) );
  NAND2X0 U15301 ( .IN1(test_so72), .IN2(n14188), .QN(n14192) );
  NAND2X0 U15302 ( .IN1(n14194), .IN2(n14195), .QN(g25600) );
  NAND2X0 U15303 ( .IN1(n14185), .IN2(g168), .QN(n14195) );
  NAND2X0 U15304 ( .IN1(n14188), .IN2(g174), .QN(n14194) );
  INVX0 U15305 ( .INP(n14185), .ZN(n14188) );
  NOR2X0 U15306 ( .IN1(n13498), .IN2(n8554), .QN(n14185) );
  NOR2X0 U15307 ( .IN1(g370), .IN2(n917), .QN(n13498) );
  NAND2X0 U15308 ( .IN1(n9590), .IN2(n14196), .QN(g25599) );
  NAND2X0 U15309 ( .IN1(n8611), .IN2(g385), .QN(n14196) );
  NAND2X0 U15310 ( .IN1(n14197), .IN2(n14198), .QN(g25598) );
  NAND3X0 U15311 ( .IN1(n8504), .IN2(g385), .IN3(n917), .QN(n14198) );
  NAND2X0 U15312 ( .IN1(n14199), .IN2(g376), .QN(n14197) );
  NAND2X0 U15313 ( .IN1(n14200), .IN2(n8515), .QN(n14199) );
  NAND2X0 U15314 ( .IN1(n917), .IN2(g358), .QN(n14200) );
  NAND3X0 U15315 ( .IN1(g376), .IN2(g358), .IN3(g385), .QN(n917) );
  NAND2X0 U15316 ( .IN1(n14201), .IN2(n14202), .QN(g25597) );
  NAND2X0 U15317 ( .IN1(n8611), .IN2(g358), .QN(n14202) );
  NAND2X0 U15318 ( .IN1(n14203), .IN2(n8515), .QN(n14201) );
  XOR2X1 U15319 ( .IN1(n7874), .IN2(n9590), .Q(n14203) );
  NAND3X0 U15320 ( .IN1(g376), .IN2(g8719), .IN3(g385), .QN(n9590) );
  NAND2X0 U15321 ( .IN1(n14204), .IN2(n14205), .QN(g25596) );
  NAND2X0 U15322 ( .IN1(n8611), .IN2(g370), .QN(n14205) );
  NAND2X0 U15323 ( .IN1(n14206), .IN2(n8515), .QN(n14204) );
  XOR2X1 U15324 ( .IN1(n7872), .IN2(n5633), .Q(n14206) );
  AND3X1 U15325 ( .IN1(n7872), .IN2(n8528), .IN3(n7873), .Q(g25595) );
  AND3X1 U15326 ( .IN1(n13515), .IN2(n8528), .IN3(n13520), .Q(g25594) );
  NAND4X0 U15327 ( .IN1(n7869), .IN2(n7868), .IN3(n7870), .IN4(n14207), .QN(
        n13520) );
  NOR4X0 U15328 ( .IN1(n7997), .IN2(n7996), .IN3(n6008), .IN4(n5597), .QN(
        n14207) );
  NAND2X0 U15329 ( .IN1(n5627), .IN2(n14208), .QN(n13515) );
  NAND4X0 U15330 ( .IN1(n7996), .IN2(n6008), .IN3(n7997), .IN4(n14209), .QN(
        n14208) );
  NOR4X0 U15331 ( .IN1(n7870), .IN2(n7869), .IN3(n7868), .IN4(g225), .QN(
        n14209) );
  NAND2X0 U15332 ( .IN1(n14210), .IN2(n14211), .QN(g25593) );
  OR2X1 U15333 ( .IN1(n8480), .IN2(n7847), .Q(n14211) );
  NAND2X0 U15334 ( .IN1(n14212), .IN2(n8515), .QN(n14210) );
  NAND2X0 U15335 ( .IN1(n14213), .IN2(n14214), .QN(n14212) );
  NAND2X0 U15336 ( .IN1(n14215), .IN2(g209), .QN(n14214) );
  NAND2X0 U15337 ( .IN1(n14216), .IN2(n14217), .QN(n14213) );
  INVX0 U15338 ( .INP(n14215), .ZN(n14217) );
  NAND2X0 U15339 ( .IN1(n14218), .IN2(n14219), .QN(g25592) );
  OR2X1 U15340 ( .IN1(n8479), .IN2(n8187), .Q(n14219) );
  NAND2X0 U15341 ( .IN1(n14220), .IN2(n8515), .QN(n14218) );
  XNOR2X1 U15342 ( .IN1(n7846), .IN2(n14221), .Q(n14220) );
  NOR2X0 U15343 ( .IN1(n14215), .IN2(n14216), .QN(n14221) );
  XOR2X1 U15344 ( .IN1(n7846), .IN2(n7847), .Q(n14216) );
  NAND2X0 U15345 ( .IN1(test_so42), .IN2(g218), .QN(n14215) );
  NAND2X0 U15346 ( .IN1(n14222), .IN2(n14223), .QN(g25591) );
  NAND2X0 U15347 ( .IN1(n8138), .IN2(n8515), .QN(n14223) );
  NAND2X0 U15348 ( .IN1(n8612), .IN2(g209), .QN(n14222) );
  NOR2X0 U15349 ( .IN1(n8125), .IN2(n14224), .QN(g24355) );
  NOR2X0 U15350 ( .IN1(n8574), .IN2(n14225), .QN(n14224) );
  NAND2X0 U15351 ( .IN1(n14226), .IN2(n14227), .QN(g24354) );
  NAND2X0 U15352 ( .IN1(n8612), .IN2(g6727), .QN(n14227) );
  NAND3X0 U15353 ( .IN1(n8124), .IN2(n14225), .IN3(n8500), .QN(n14226) );
  OR2X1 U15354 ( .IN1(n14228), .IN2(n5531), .Q(n14225) );
  NAND2X0 U15355 ( .IN1(n14229), .IN2(n14230), .QN(g24353) );
  NAND2X0 U15356 ( .IN1(n8613), .IN2(g6723), .QN(n14230) );
  NAND2X0 U15357 ( .IN1(n14231), .IN2(n8515), .QN(n14229) );
  XOR2X1 U15358 ( .IN1(n14228), .IN2(n5531), .Q(n14231) );
  NAND4X0 U15359 ( .IN1(test_so80), .IN2(g14828), .IN3(g17688), .IN4(g17778), 
        .QN(n14228) );
  NOR4X0 U15360 ( .IN1(n14232), .IN2(g13099), .IN3(n14233), .IN4(n14234), .QN(
        g24352) );
  NOR2X0 U15361 ( .IN1(test_so80), .IN2(n5700), .QN(n14234) );
  NOR2X0 U15362 ( .IN1(n7978), .IN2(g14828), .QN(n14233) );
  NAND3X0 U15363 ( .IN1(n7964), .IN2(n8482), .IN3(n8083), .QN(n14232) );
  NOR2X0 U15364 ( .IN1(n7987), .IN2(n14235), .QN(g24351) );
  NOR2X0 U15365 ( .IN1(n8575), .IN2(n14236), .QN(n14235) );
  NAND2X0 U15366 ( .IN1(n14237), .IN2(n14238), .QN(g24350) );
  NAND2X0 U15367 ( .IN1(test_so69), .IN2(n8659), .QN(n14238) );
  NAND3X0 U15368 ( .IN1(n7986), .IN2(n14236), .IN3(n8500), .QN(n14237) );
  NAND2X0 U15369 ( .IN1(n14239), .IN2(test_so69), .QN(n14236) );
  NAND2X0 U15370 ( .IN1(n14240), .IN2(n14241), .QN(g24349) );
  NAND2X0 U15371 ( .IN1(n8613), .IN2(g6377), .QN(n14241) );
  NAND2X0 U15372 ( .IN1(n14242), .IN2(n8515), .QN(n14240) );
  XOR2X1 U15373 ( .IN1(test_so69), .IN2(n14239), .Q(n14242) );
  NOR4X0 U15374 ( .IN1(n5437), .IN2(n5703), .IN3(n7967), .IN4(n7982), .QN(
        n14239) );
  NOR4X0 U15375 ( .IN1(n14243), .IN2(g13085), .IN3(n14244), .IN4(n14245), .QN(
        g24348) );
  NOR2X0 U15376 ( .IN1(n5703), .IN2(g12422), .QN(n14245) );
  NOR2X0 U15377 ( .IN1(n7982), .IN2(g14779), .QN(n14244) );
  NAND3X0 U15378 ( .IN1(n7967), .IN2(n8483), .IN3(n8093), .QN(n14243) );
  NOR2X0 U15379 ( .IN1(n7988), .IN2(n14246), .QN(g24347) );
  NOR2X0 U15380 ( .IN1(n8573), .IN2(n14247), .QN(n14246) );
  NAND2X0 U15381 ( .IN1(n14248), .IN2(n14249), .QN(g24346) );
  NAND2X0 U15382 ( .IN1(n8613), .IN2(g6035), .QN(n14249) );
  NAND3X0 U15383 ( .IN1(n14247), .IN2(n8230), .IN3(n8500), .QN(n14248) );
  OR2X1 U15384 ( .IN1(n14250), .IN2(n5528), .Q(n14247) );
  NAND2X0 U15385 ( .IN1(n14251), .IN2(n14252), .QN(g24345) );
  NAND2X0 U15386 ( .IN1(n8613), .IN2(g6031), .QN(n14252) );
  NAND2X0 U15387 ( .IN1(n14253), .IN2(n8515), .QN(n14251) );
  XOR2X1 U15388 ( .IN1(n14250), .IN2(n5528), .Q(n14253) );
  NAND4X0 U15389 ( .IN1(g12350), .IN2(g14738), .IN3(g17607), .IN4(g17739), 
        .QN(n14250) );
  NOR4X0 U15390 ( .IN1(n14254), .IN2(g13068), .IN3(n14255), .IN4(n14256), .QN(
        g24344) );
  NOR2X0 U15391 ( .IN1(n5698), .IN2(g12350), .QN(n14256) );
  NOR2X0 U15392 ( .IN1(n7973), .IN2(g14738), .QN(n14255) );
  NAND3X0 U15393 ( .IN1(n7958), .IN2(n8484), .IN3(n8069), .QN(n14254) );
  NOR2X0 U15394 ( .IN1(n7992), .IN2(n14257), .QN(g24343) );
  NOR2X0 U15395 ( .IN1(n8575), .IN2(n14258), .QN(n14257) );
  NAND2X0 U15396 ( .IN1(n14259), .IN2(n14260), .QN(g24342) );
  NAND2X0 U15397 ( .IN1(n8613), .IN2(g5689), .QN(n14260) );
  NAND3X0 U15398 ( .IN1(n7991), .IN2(n14258), .IN3(n8499), .QN(n14259) );
  OR2X1 U15399 ( .IN1(n14261), .IN2(n5529), .Q(n14258) );
  NAND2X0 U15400 ( .IN1(n14262), .IN2(n14263), .QN(g24341) );
  NAND2X0 U15401 ( .IN1(n8589), .IN2(g5685), .QN(n14263) );
  NAND2X0 U15402 ( .IN1(n14264), .IN2(n8516), .QN(n14262) );
  XOR2X1 U15403 ( .IN1(n14261), .IN2(n5529), .Q(n14264) );
  NAND4X0 U15404 ( .IN1(g12300), .IN2(g14694), .IN3(g17580), .IN4(g17711), 
        .QN(n14261) );
  NOR4X0 U15405 ( .IN1(n14265), .IN2(g13049), .IN3(n14266), .IN4(n14267), .QN(
        g24340) );
  NOR2X0 U15406 ( .IN1(n5705), .IN2(g12300), .QN(n14267) );
  NOR2X0 U15407 ( .IN1(n7975), .IN2(g14694), .QN(n14266) );
  NAND3X0 U15408 ( .IN1(n7960), .IN2(n8484), .IN3(n8074), .QN(n14265) );
  NOR2X0 U15409 ( .IN1(n8127), .IN2(n14268), .QN(g24339) );
  NOR2X0 U15410 ( .IN1(n8575), .IN2(n14269), .QN(n14268) );
  NAND2X0 U15411 ( .IN1(n14270), .IN2(n14271), .QN(g24338) );
  NAND2X0 U15412 ( .IN1(test_so10), .IN2(n8659), .QN(n14271) );
  NAND3X0 U15413 ( .IN1(n8126), .IN2(n14269), .IN3(n8499), .QN(n14270) );
  NAND2X0 U15414 ( .IN1(n14272), .IN2(test_so10), .QN(n14269) );
  NAND2X0 U15415 ( .IN1(n14273), .IN2(n14274), .QN(g24337) );
  NAND2X0 U15416 ( .IN1(n8591), .IN2(g5339), .QN(n14274) );
  NAND2X0 U15417 ( .IN1(n14275), .IN2(n8516), .QN(n14273) );
  XOR2X1 U15418 ( .IN1(test_so10), .IN2(n14272), .Q(n14275) );
  NOR4X0 U15419 ( .IN1(n5438), .IN2(n5704), .IN3(n7956), .IN4(n7971), .QN(
        n14272) );
  NOR4X0 U15420 ( .IN1(n14276), .IN2(g17577), .IN3(n14277), .IN4(n14278), .QN(
        g24336) );
  NOR2X0 U15421 ( .IN1(n5704), .IN2(g12238), .QN(n14278) );
  NOR2X0 U15422 ( .IN1(n7971), .IN2(g14662), .QN(n14277) );
  NAND3X0 U15423 ( .IN1(n7956), .IN2(n8483), .IN3(n8041), .QN(n14276) );
  NAND2X0 U15424 ( .IN1(n14279), .IN2(n14280), .QN(g24335) );
  OR3X1 U15425 ( .IN1(g4340), .IN2(n5382), .IN3(n14281), .Q(n14280) );
  OR2X1 U15426 ( .IN1(n8476), .IN2(n5541), .Q(n14279) );
  NAND2X0 U15427 ( .IN1(n14282), .IN2(n14283), .QN(g24334) );
  NAND4X0 U15428 ( .IN1(n5303), .IN2(n5365), .IN3(n14284), .IN4(n14285), .QN(
        n14283) );
  NOR4X0 U15429 ( .IN1(g4584), .IN2(g4608), .IN3(g4616), .IN4(n14281), .QN(
        n14285) );
  NAND4X0 U15430 ( .IN1(n8508), .IN2(n8208), .IN3(n5506), .IN4(n14286), .QN(
        n14281) );
  AND3X1 U15431 ( .IN1(n5323), .IN2(n5540), .IN3(n5348), .Q(n14286) );
  NOR3X0 U15432 ( .IN1(n9724), .IN2(n5844), .IN3(n5653), .QN(n14284) );
  NAND2X0 U15433 ( .IN1(test_so3), .IN2(n5727), .QN(n9724) );
  NAND2X0 U15434 ( .IN1(n8590), .IN2(g4358), .QN(n14282) );
  NOR2X0 U15435 ( .IN1(n5710), .IN2(n8505), .QN(g24298) );
  NAND2X0 U15436 ( .IN1(n14287), .IN2(n14288), .QN(g24282) );
  NAND2X0 U15437 ( .IN1(n14289), .IN2(g4308), .QN(n14288) );
  NAND2X0 U15438 ( .IN1(n8512), .IN2(g9251), .QN(n14289) );
  NAND2X0 U15439 ( .IN1(g24281), .IN2(g9251), .QN(n14287) );
  NOR2X0 U15440 ( .IN1(g4308), .IN2(n8558), .QN(g24281) );
  NAND2X0 U15441 ( .IN1(n14290), .IN2(n14291), .QN(g24280) );
  NAND2X0 U15442 ( .IN1(n14292), .IN2(g4269), .QN(n14291) );
  NAND2X0 U15443 ( .IN1(n14293), .IN2(n8516), .QN(n14292) );
  NAND3X0 U15444 ( .IN1(g4264), .IN2(g4258), .IN3(n5764), .QN(n14293) );
  NAND2X0 U15445 ( .IN1(n14294), .IN2(g4273), .QN(n14290) );
  NAND2X0 U15446 ( .IN1(n14295), .IN2(n14296), .QN(n14294) );
  NAND2X0 U15447 ( .IN1(n5763), .IN2(n8516), .QN(n14296) );
  NAND3X0 U15448 ( .IN1(n14297), .IN2(n14298), .IN3(n14299), .QN(g24279) );
  NAND2X0 U15449 ( .IN1(n14300), .IN2(n14301), .QN(n14299) );
  OR2X1 U15450 ( .IN1(n8476), .IN2(n7920), .Q(n14298) );
  NAND2X0 U15451 ( .IN1(n14302), .IN2(n8517), .QN(n14297) );
  NAND2X0 U15452 ( .IN1(n14303), .IN2(n14304), .QN(n14302) );
  NAND3X0 U15453 ( .IN1(n14305), .IN2(n14306), .IN3(n14307), .QN(n14304) );
  INVX0 U15454 ( .INP(n14300), .ZN(n14306) );
  NOR2X0 U15455 ( .IN1(n7920), .IN2(n5726), .QN(n14300) );
  OR2X1 U15456 ( .IN1(n14307), .IN2(n14305), .Q(n14303) );
  INVX0 U15457 ( .INP(n14301), .ZN(n14305) );
  NAND3X0 U15458 ( .IN1(n5726), .IN2(n14308), .IN3(n7920), .QN(n14307) );
  NAND4X0 U15459 ( .IN1(n14524), .IN2(n14525), .IN3(n14523), .IN4(n14309), 
        .QN(n14308) );
  NOR4X0 U15460 ( .IN1(g8915), .IN2(g8916), .IN3(g11770), .IN4(g8920), .QN(
        n14309) );
  NOR2X0 U15461 ( .IN1(n7994), .IN2(n14310), .QN(g24278) );
  NOR2X0 U15462 ( .IN1(n8575), .IN2(n14311), .QN(n14310) );
  NAND2X0 U15463 ( .IN1(n14312), .IN2(n14313), .QN(g24277) );
  NAND2X0 U15464 ( .IN1(n8587), .IN2(g4040), .QN(n14313) );
  NAND3X0 U15465 ( .IN1(n7993), .IN2(n14311), .IN3(n8497), .QN(n14312) );
  OR2X1 U15466 ( .IN1(n14314), .IN2(n5530), .Q(n14311) );
  NAND2X0 U15467 ( .IN1(n14315), .IN2(n14316), .QN(g24276) );
  NAND2X0 U15468 ( .IN1(n8592), .IN2(g4031), .QN(n14316) );
  NAND2X0 U15469 ( .IN1(n14317), .IN2(n8517), .QN(n14315) );
  XOR2X1 U15470 ( .IN1(n14314), .IN2(n5530), .Q(n14317) );
  NAND4X0 U15471 ( .IN1(g11418), .IN2(g13966), .IN3(g16659), .IN4(g16775), 
        .QN(n14314) );
  NOR4X0 U15472 ( .IN1(n14318), .IN2(g14518), .IN3(n14319), .IN4(n14320), .QN(
        g24275) );
  NOR2X0 U15473 ( .IN1(n5701), .IN2(g11418), .QN(n14320) );
  NOR2X0 U15474 ( .IN1(n7976), .IN2(g13966), .QN(n14319) );
  NAND3X0 U15475 ( .IN1(n7962), .IN2(n8482), .IN3(n8078), .QN(n14318) );
  NOR2X0 U15476 ( .IN1(n7990), .IN2(n14321), .QN(g24274) );
  NOR2X0 U15477 ( .IN1(n8574), .IN2(n14322), .QN(n14321) );
  NAND2X0 U15478 ( .IN1(n14323), .IN2(n14324), .QN(g24273) );
  NAND2X0 U15479 ( .IN1(n8593), .IN2(g3689), .QN(n14324) );
  NAND3X0 U15480 ( .IN1(n7989), .IN2(n14322), .IN3(n8497), .QN(n14323) );
  OR2X1 U15481 ( .IN1(n14325), .IN2(n5532), .Q(n14322) );
  NAND2X0 U15482 ( .IN1(n14326), .IN2(n14327), .QN(g24272) );
  NAND2X0 U15483 ( .IN1(n8602), .IN2(g3680), .QN(n14327) );
  NAND2X0 U15484 ( .IN1(n14328), .IN2(n8517), .QN(n14326) );
  XOR2X1 U15485 ( .IN1(n14325), .IN2(n5532), .Q(n14328) );
  NAND4X0 U15486 ( .IN1(g11388), .IN2(g13926), .IN3(g16627), .IN4(g16744), 
        .QN(n14325) );
  NOR4X0 U15487 ( .IN1(n14329), .IN2(g14451), .IN3(n14330), .IN4(n14331), .QN(
        g24271) );
  NOR2X0 U15488 ( .IN1(n5699), .IN2(g11388), .QN(n14331) );
  NOR2X0 U15489 ( .IN1(n7980), .IN2(g13926), .QN(n14330) );
  NAND3X0 U15490 ( .IN1(n7966), .IN2(n8483), .IN3(n8088), .QN(n14329) );
  NOR2X0 U15491 ( .IN1(n7985), .IN2(n14332), .QN(g24270) );
  NOR2X0 U15492 ( .IN1(n8574), .IN2(n14333), .QN(n14332) );
  NAND2X0 U15493 ( .IN1(n14334), .IN2(n14335), .QN(g24269) );
  NAND2X0 U15494 ( .IN1(n8594), .IN2(g3338), .QN(n14335) );
  NAND3X0 U15495 ( .IN1(n7984), .IN2(n14333), .IN3(n8497), .QN(n14334) );
  OR2X1 U15496 ( .IN1(n14336), .IN2(n5527), .Q(n14333) );
  NAND2X0 U15497 ( .IN1(n14337), .IN2(n14338), .QN(g24268) );
  NAND2X0 U15498 ( .IN1(test_so91), .IN2(n8559), .QN(n14338) );
  NAND2X0 U15499 ( .IN1(n14339), .IN2(n8517), .QN(n14337) );
  XOR2X1 U15500 ( .IN1(n14336), .IN2(n5527), .Q(n14339) );
  NAND4X0 U15501 ( .IN1(g11349), .IN2(g13895), .IN3(g16603), .IN4(g16718), 
        .QN(n14336) );
  NOR4X0 U15502 ( .IN1(n14340), .IN2(g14421), .IN3(n14341), .IN4(n14342), .QN(
        g24267) );
  NOR2X0 U15503 ( .IN1(n5702), .IN2(g11349), .QN(n14342) );
  NOR2X0 U15504 ( .IN1(n7969), .IN2(g13895), .QN(n14341) );
  NAND3X0 U15505 ( .IN1(n7954), .IN2(n8483), .IN3(n8059), .QN(n14340) );
  NAND2X0 U15506 ( .IN1(n14343), .IN2(n14344), .QN(g24266) );
  OR2X1 U15507 ( .IN1(n8477), .IN2(n5963), .Q(n14344) );
  NAND3X0 U15508 ( .IN1(test_so9), .IN2(n7722), .IN3(n8496), .QN(n14343) );
  NAND3X0 U15509 ( .IN1(n14345), .IN2(n14346), .IN3(n8807), .QN(g24263) );
  NAND2X0 U15510 ( .IN1(n5963), .IN2(n8517), .QN(n8807) );
  NAND2X0 U15511 ( .IN1(n5299), .IN2(n8517), .QN(n14346) );
  OR2X1 U15512 ( .IN1(n8477), .IN2(n7722), .Q(n14345) );
  NAND3X0 U15513 ( .IN1(n14347), .IN2(n14348), .IN3(n14349), .QN(g24262) );
  NAND2X0 U15514 ( .IN1(n14350), .IN2(n8154), .QN(n14349) );
  NAND3X0 U15515 ( .IN1(n14351), .IN2(g1564), .IN3(n8496), .QN(n14348) );
  NAND2X0 U15516 ( .IN1(n8598), .IN2(g1548), .QN(n14347) );
  NAND2X0 U15517 ( .IN1(n10807), .IN2(n14352), .QN(g24261) );
  NAND2X0 U15518 ( .IN1(n8599), .IN2(g1585), .QN(n14352) );
  XOR2X1 U15519 ( .IN1(n14353), .IN2(n8155), .Q(g24260) );
  NAND2X0 U15520 ( .IN1(n8511), .IN2(g1548), .QN(n14353) );
  NAND2X0 U15521 ( .IN1(n10807), .IN2(n14354), .QN(g24259) );
  OR2X1 U15522 ( .IN1(n8478), .IN2(n7809), .Q(n14354) );
  NAND2X0 U15523 ( .IN1(n14355), .IN2(n14356), .QN(g24258) );
  NAND2X0 U15524 ( .IN1(n8510), .IN2(g496), .QN(n14356) );
  NAND2X0 U15525 ( .IN1(n8596), .IN2(g1554), .QN(n14355) );
  XOR2X1 U15526 ( .IN1(n14357), .IN2(n5616), .Q(g24257) );
  OR2X1 U15527 ( .IN1(n14358), .IN2(n8546), .Q(n14357) );
  NAND2X0 U15528 ( .IN1(n14359), .IN2(n14360), .QN(g24256) );
  NAND2X0 U15529 ( .IN1(n8597), .IN2(g1339), .QN(n14360) );
  NAND2X0 U15530 ( .IN1(n14361), .IN2(n8516), .QN(n14359) );
  XOR2X1 U15531 ( .IN1(n14358), .IN2(n14362), .Q(n14361) );
  NAND3X0 U15532 ( .IN1(n7744), .IN2(n14061), .IN3(n7832), .QN(n14362) );
  AND3X1 U15533 ( .IN1(n5302), .IN2(n5616), .IN3(n5401), .Q(n14061) );
  NAND3X0 U15534 ( .IN1(n13694), .IN2(n14363), .IN3(n14364), .QN(n14358) );
  XOR2X1 U15535 ( .IN1(n7809), .IN2(n8203), .Q(n14364) );
  NAND3X0 U15536 ( .IN1(n14365), .IN2(n14366), .IN3(n14367), .QN(g24255) );
  NAND2X0 U15537 ( .IN1(n11235), .IN2(g17423), .QN(n14367) );
  NAND3X0 U15538 ( .IN1(n7822), .IN2(g10527), .IN3(n8495), .QN(n14366) );
  NAND2X0 U15539 ( .IN1(n8604), .IN2(g1589), .QN(n14365) );
  NOR4X0 U15540 ( .IN1(g17423), .IN2(n14368), .IN3(g17404), .IN4(g17320), .QN(
        g24254) );
  NAND2X0 U15541 ( .IN1(n14369), .IN2(n8516), .QN(n14368) );
  NAND3X0 U15542 ( .IN1(n14370), .IN2(g1554), .IN3(n14040), .QN(n14369) );
  INVX0 U15543 ( .INP(n14039), .ZN(n14040) );
  NAND2X0 U15544 ( .IN1(n14350), .IN2(g1564), .QN(n14039) );
  INVX0 U15545 ( .INP(n14351), .ZN(n14350) );
  NAND2X0 U15546 ( .IN1(g1430), .IN2(g1548), .QN(n14351) );
  NAND2X0 U15547 ( .IN1(n13694), .IN2(n14363), .QN(n14370) );
  INVX0 U15548 ( .INP(n4836), .ZN(n14363) );
  NAND2X0 U15549 ( .IN1(n5466), .IN2(n5322), .QN(n4836) );
  NOR2X0 U15550 ( .IN1(n13441), .IN2(n13444), .QN(n13694) );
  INVX0 U15551 ( .INP(n12360), .ZN(n13444) );
  NAND2X0 U15552 ( .IN1(n5616), .IN2(n8203), .QN(n12360) );
  XOR2X1 U15553 ( .IN1(g1339), .IN2(n8203), .Q(n13441) );
  NAND2X0 U15554 ( .IN1(n14371), .IN2(n14372), .QN(g24253) );
  NAND2X0 U15555 ( .IN1(n8605), .IN2(g1306), .QN(n14372) );
  NAND2X0 U15556 ( .IN1(n14373), .IN2(n8516), .QN(n14371) );
  NAND2X0 U15557 ( .IN1(n14374), .IN2(n14375), .QN(n14373) );
  NAND2X0 U15558 ( .IN1(n5302), .IN2(g1532), .QN(n14375) );
  NAND2X0 U15559 ( .IN1(g7946), .IN2(g1521), .QN(n14374) );
  NAND2X0 U15560 ( .IN1(n14376), .IN2(n14377), .QN(g24252) );
  NAND2X0 U15561 ( .IN1(test_so49), .IN2(n8560), .QN(n14377) );
  NAND2X0 U15562 ( .IN1(n14378), .IN2(n8516), .QN(n14376) );
  NAND2X0 U15563 ( .IN1(n14050), .IN2(n14379), .QN(n14378) );
  NAND2X0 U15564 ( .IN1(n5302), .IN2(g1521), .QN(n14379) );
  NAND2X0 U15565 ( .IN1(g7946), .IN2(g1339), .QN(n14050) );
  NAND2X0 U15566 ( .IN1(n14380), .IN2(n14381), .QN(g24251) );
  NAND2X0 U15567 ( .IN1(n12833), .IN2(g1442), .QN(n14381) );
  NAND2X0 U15568 ( .IN1(test_so12), .IN2(n14057), .QN(n14380) );
  NAND2X0 U15569 ( .IN1(n14382), .IN2(n14383), .QN(g24250) );
  NAND2X0 U15570 ( .IN1(test_so12), .IN2(n12833), .QN(n14383) );
  NAND2X0 U15571 ( .IN1(n14057), .IN2(g1489), .QN(n14382) );
  NAND2X0 U15572 ( .IN1(n14384), .IN2(n14385), .QN(g24249) );
  NAND3X0 U15573 ( .IN1(n8137), .IN2(n8482), .IN3(n12837), .QN(n14385) );
  NAND2X0 U15574 ( .IN1(n14386), .IN2(g1489), .QN(n14384) );
  NAND2X0 U15575 ( .IN1(n14057), .IN2(n14387), .QN(n14386) );
  OR2X1 U15576 ( .IN1(n8547), .IN2(test_so12), .Q(n14387) );
  INVX0 U15577 ( .INP(n12833), .ZN(n14057) );
  NOR2X0 U15578 ( .IN1(n12837), .IN2(n8563), .QN(n12833) );
  AND3X1 U15579 ( .IN1(g13272), .IN2(n8206), .IN3(n5364), .Q(n12837) );
  NAND3X0 U15580 ( .IN1(n14388), .IN2(n14389), .IN3(n14390), .QN(g24248) );
  XNOR2X1 U15581 ( .IN1(n7839), .IN2(n14391), .Q(n14390) );
  NAND2X0 U15582 ( .IN1(n5655), .IN2(n8516), .QN(n14391) );
  NAND2X0 U15583 ( .IN1(n11235), .IN2(g1395), .QN(n14389) );
  INVX0 U15584 ( .INP(n10807), .ZN(n11235) );
  NAND2X0 U15585 ( .IN1(n5401), .IN2(n8516), .QN(n14388) );
  NOR2X0 U15586 ( .IN1(g1249), .IN2(n10807), .QN(g24247) );
  NAND2X0 U15587 ( .IN1(n8510), .IN2(g12923), .QN(n10807) );
  NAND3X0 U15588 ( .IN1(n14392), .IN2(n14393), .IN3(n14394), .QN(g24246) );
  NAND2X0 U15589 ( .IN1(n14395), .IN2(n8156), .QN(n14394) );
  NAND3X0 U15590 ( .IN1(n14396), .IN2(g1221), .IN3(n8495), .QN(n14393) );
  NAND2X0 U15591 ( .IN1(n8606), .IN2(g1205), .QN(n14392) );
  NAND2X0 U15592 ( .IN1(n10820), .IN2(n14397), .QN(g24245) );
  NAND2X0 U15593 ( .IN1(n8607), .IN2(g30332), .QN(n14397) );
  XOR2X1 U15594 ( .IN1(n14398), .IN2(n8157), .Q(g24244) );
  NAND2X0 U15595 ( .IN1(n8509), .IN2(g1205), .QN(n14398) );
  NAND2X0 U15596 ( .IN1(n10820), .IN2(n14399), .QN(g24243) );
  OR2X1 U15597 ( .IN1(n8479), .IN2(n7808), .Q(n14399) );
  NAND2X0 U15598 ( .IN1(n14400), .IN2(n14401), .QN(g24242) );
  NAND2X0 U15599 ( .IN1(n8509), .IN2(g29215), .QN(n14401) );
  NAND2X0 U15600 ( .IN1(test_so76), .IN2(n8553), .QN(n14400) );
  XOR2X1 U15601 ( .IN1(n14402), .IN2(n5622), .Q(g24241) );
  OR2X1 U15602 ( .IN1(n14403), .IN2(n8546), .Q(n14402) );
  NAND2X0 U15603 ( .IN1(n14404), .IN2(n14405), .QN(g24240) );
  NAND2X0 U15604 ( .IN1(n8612), .IN2(g996), .QN(n14405) );
  NAND2X0 U15605 ( .IN1(n14406), .IN2(n8514), .QN(n14404) );
  XOR2X1 U15606 ( .IN1(n14403), .IN2(n14407), .Q(n14406) );
  NAND3X0 U15607 ( .IN1(n7730), .IN2(n14113), .IN3(n7831), .QN(n14407) );
  AND3X1 U15608 ( .IN1(n5304), .IN2(n5622), .IN3(n5392), .Q(n14113) );
  NAND3X0 U15609 ( .IN1(n14408), .IN2(n14409), .IN3(n13725), .QN(n14403) );
  INVX0 U15610 ( .INP(n14117), .ZN(n13725) );
  INVX0 U15611 ( .INP(n4837), .ZN(n14409) );
  XOR2X1 U15612 ( .IN1(n7808), .IN2(n5320), .Q(n14408) );
  NAND3X0 U15613 ( .IN1(n14410), .IN2(n14411), .IN3(n14412), .QN(g24239) );
  NAND2X0 U15614 ( .IN1(n11250), .IN2(g17400), .QN(n14412) );
  NAND3X0 U15615 ( .IN1(n7811), .IN2(g10500), .IN3(n8493), .QN(n14411) );
  NAND2X0 U15616 ( .IN1(n8655), .IN2(g1246), .QN(n14410) );
  NOR4X0 U15617 ( .IN1(n14413), .IN2(n14414), .IN3(g17400), .IN4(g17291), .QN(
        g24238) );
  OR2X1 U15618 ( .IN1(n8547), .IN2(test_so44), .Q(n14414) );
  NOR3X0 U15619 ( .IN1(n8212), .IN2(n14415), .IN3(n14089), .QN(n14413) );
  NAND2X0 U15620 ( .IN1(n14395), .IN2(g1221), .QN(n14089) );
  INVX0 U15621 ( .INP(n14396), .ZN(n14395) );
  NAND2X0 U15622 ( .IN1(g1087), .IN2(g1205), .QN(n14396) );
  NOR2X0 U15623 ( .IN1(n4837), .IN2(n14117), .QN(n14415) );
  NAND2X0 U15624 ( .IN1(n13456), .IN2(n12391), .QN(n14117) );
  NAND2X0 U15625 ( .IN1(n5622), .IN2(n5320), .QN(n12391) );
  XNOR2X1 U15626 ( .IN1(g996), .IN2(n5320), .Q(n13456) );
  NAND2X0 U15627 ( .IN1(n5321), .IN2(n8223), .QN(n4837) );
  NAND2X0 U15628 ( .IN1(n14416), .IN2(n14417), .QN(g24237) );
  NAND2X0 U15629 ( .IN1(n8656), .IN2(g962), .QN(n14417) );
  NAND2X0 U15630 ( .IN1(n14418), .IN2(n8514), .QN(n14416) );
  NAND2X0 U15631 ( .IN1(n14419), .IN2(n14420), .QN(n14418) );
  NAND2X0 U15632 ( .IN1(n5304), .IN2(g1189), .QN(n14420) );
  NAND2X0 U15633 ( .IN1(g7916), .IN2(g1178), .QN(n14419) );
  NAND2X0 U15634 ( .IN1(n14421), .IN2(n14422), .QN(g24236) );
  NAND2X0 U15635 ( .IN1(n8538), .IN2(g1183), .QN(n14422) );
  NAND2X0 U15636 ( .IN1(n14423), .IN2(n8514), .QN(n14421) );
  NAND2X0 U15637 ( .IN1(n14100), .IN2(n14424), .QN(n14423) );
  NAND2X0 U15638 ( .IN1(n5304), .IN2(g1178), .QN(n14424) );
  NAND2X0 U15639 ( .IN1(g7916), .IN2(g996), .QN(n14100) );
  NAND2X0 U15640 ( .IN1(n14425), .IN2(n14426), .QN(g24235) );
  NAND2X0 U15641 ( .IN1(test_so7), .IN2(n12865), .QN(n14426) );
  NAND2X0 U15642 ( .IN1(n14107), .IN2(g1152), .QN(n14425) );
  NAND2X0 U15643 ( .IN1(n14427), .IN2(n14428), .QN(g24234) );
  NAND2X0 U15644 ( .IN1(n12865), .IN2(g1152), .QN(n14428) );
  NAND2X0 U15645 ( .IN1(n14107), .IN2(g1146), .QN(n14427) );
  NAND2X0 U15646 ( .IN1(n14429), .IN2(n14430), .QN(g24233) );
  NAND3X0 U15647 ( .IN1(n8504), .IN2(n8207), .IN3(n12869), .QN(n14430) );
  NAND2X0 U15648 ( .IN1(n14431), .IN2(g1146), .QN(n14429) );
  NAND2X0 U15649 ( .IN1(n14107), .IN2(n14432), .QN(n14431) );
  NAND2X0 U15650 ( .IN1(n5618), .IN2(n8514), .QN(n14432) );
  INVX0 U15651 ( .INP(n12865), .ZN(n14107) );
  NOR2X0 U15652 ( .IN1(n12869), .IN2(n8562), .QN(n12865) );
  AND3X1 U15653 ( .IN1(n5363), .IN2(g13259), .IN3(n5599), .Q(n12869) );
  NAND3X0 U15654 ( .IN1(n14433), .IN2(n14434), .IN3(n14435), .QN(g24232) );
  XNOR2X1 U15655 ( .IN1(n7840), .IN2(n14436), .Q(n14435) );
  NAND2X0 U15656 ( .IN1(n5654), .IN2(n8514), .QN(n14436) );
  NAND2X0 U15657 ( .IN1(n11250), .IN2(g1052), .QN(n14434) );
  INVX0 U15658 ( .INP(n10820), .ZN(n11250) );
  NAND2X0 U15659 ( .IN1(n5392), .IN2(n8513), .QN(n14433) );
  NOR2X0 U15660 ( .IN1(g904), .IN2(n10820), .QN(g24231) );
  NAND2X0 U15661 ( .IN1(n8510), .IN2(g12919), .QN(n10820) );
  NAND2X0 U15662 ( .IN1(n14437), .IN2(n14438), .QN(g24216) );
  NAND2X0 U15663 ( .IN1(n12923), .IN2(g847), .QN(n14438) );
  NAND2X0 U15664 ( .IN1(n14149), .IN2(g854), .QN(n14437) );
  NAND2X0 U15665 ( .IN1(n14439), .IN2(n14440), .QN(g24215) );
  NAND2X0 U15666 ( .IN1(n14441), .IN2(g837), .QN(n14440) );
  NAND2X0 U15667 ( .IN1(n14149), .IN2(n14442), .QN(n14441) );
  NAND3X0 U15668 ( .IN1(n14443), .IN2(n8483), .IN3(n14444), .QN(n14442) );
  NAND2X0 U15669 ( .IN1(g827), .IN2(g832), .QN(n14444) );
  NAND2X0 U15670 ( .IN1(g847), .IN2(g812), .QN(n14443) );
  NAND2X0 U15671 ( .IN1(n14445), .IN2(g703), .QN(n14439) );
  NAND2X0 U15672 ( .IN1(n14446), .IN2(n8513), .QN(n14445) );
  NAND2X0 U15673 ( .IN1(n5562), .IN2(n13773), .QN(n14446) );
  NOR2X0 U15674 ( .IN1(n12926), .IN2(n5709), .QN(n13773) );
  NAND3X0 U15675 ( .IN1(n14447), .IN2(n14448), .IN3(n14449), .QN(g24214) );
  NAND2X0 U15676 ( .IN1(n14450), .IN2(g703), .QN(n14449) );
  NAND2X0 U15677 ( .IN1(n13769), .IN2(n14451), .QN(n14450) );
  OR2X1 U15678 ( .IN1(n13767), .IN2(n8546), .Q(n14451) );
  NOR2X0 U15679 ( .IN1(n5733), .IN2(n5562), .QN(n13767) );
  AND2X1 U15680 ( .IN1(n14149), .IN2(n14452), .Q(n13769) );
  NAND2X0 U15681 ( .IN1(n5709), .IN2(n8513), .QN(n14452) );
  NAND2X0 U15682 ( .IN1(n8585), .IN2(g847), .QN(n14448) );
  NAND4X0 U15683 ( .IN1(g817), .IN2(g723), .IN3(n14453), .IN4(n5709), .QN(
        n14447) );
  NOR2X0 U15684 ( .IN1(n5422), .IN2(n14148), .QN(n14453) );
  OR2X1 U15685 ( .IN1(n14454), .IN2(g24212), .Q(g24213) );
  NOR2X0 U15686 ( .IN1(n7771), .IN2(n8504), .QN(n14454) );
  NAND2X0 U15687 ( .IN1(n14455), .IN2(n14456), .QN(g24211) );
  NAND2X0 U15688 ( .IN1(n2404), .IN2(n14457), .QN(n14456) );
  NAND2X0 U15689 ( .IN1(n8232), .IN2(g691), .QN(n14457) );
  NAND2X0 U15690 ( .IN1(n8585), .IN2(g546), .QN(n14455) );
  AND3X1 U15691 ( .IN1(n14458), .IN2(n8528), .IN3(n11373), .Q(g24210) );
  AND3X1 U15692 ( .IN1(g518), .IN2(g203), .IN3(n5548), .Q(n11373) );
  NAND2X0 U15693 ( .IN1(n14459), .IN2(n14460), .QN(n14458) );
  NAND2X0 U15694 ( .IN1(test_so72), .IN2(n14461), .QN(n14460) );
  NAND2X0 U15695 ( .IN1(n5606), .IN2(n5402), .QN(n14461) );
  NAND2X0 U15696 ( .IN1(g174), .IN2(g168), .QN(n14459) );
  NAND2X0 U15697 ( .IN1(n14462), .IN2(n14463), .QN(g24209) );
  NAND2X0 U15698 ( .IN1(n12927), .IN2(g446), .QN(n14463) );
  NAND2X0 U15699 ( .IN1(n12923), .IN2(g417), .QN(n14462) );
  NAND3X0 U15700 ( .IN1(n14464), .IN2(n14465), .IN3(n14466), .QN(g24208) );
  NAND2X0 U15701 ( .IN1(n8572), .IN2(g424), .QN(n14466) );
  NAND2X0 U15702 ( .IN1(n12927), .IN2(g246), .QN(n14465) );
  NAND2X0 U15703 ( .IN1(n12923), .IN2(g475), .QN(n14464) );
  NAND2X0 U15704 ( .IN1(n14467), .IN2(n14468), .QN(g24207) );
  NAND2X0 U15705 ( .IN1(n12923), .IN2(g441), .QN(n14468) );
  NAND2X0 U15706 ( .IN1(n14149), .IN2(g475), .QN(n14467) );
  NAND2X0 U15707 ( .IN1(n14469), .IN2(n14470), .QN(g24206) );
  NAND2X0 U15708 ( .IN1(n12923), .IN2(g437), .QN(n14470) );
  NAND2X0 U15709 ( .IN1(n14149), .IN2(g441), .QN(n14469) );
  NAND3X0 U15710 ( .IN1(n14471), .IN2(n14472), .IN3(n14473), .QN(g24205) );
  NAND2X0 U15711 ( .IN1(n8643), .IN2(g437), .QN(n14473) );
  NAND2X0 U15712 ( .IN1(n12927), .IN2(g269), .QN(n14472) );
  NAND2X0 U15713 ( .IN1(test_so23), .IN2(n12923), .QN(n14471) );
  NAND2X0 U15714 ( .IN1(n14474), .IN2(n14475), .QN(g24204) );
  NAND2X0 U15715 ( .IN1(n12923), .IN2(g429), .QN(n14475) );
  NAND2X0 U15716 ( .IN1(test_so23), .IN2(n14149), .QN(n14474) );
  NAND2X0 U15717 ( .IN1(n14476), .IN2(n14477), .QN(g24203) );
  NAND2X0 U15718 ( .IN1(n12923), .IN2(g401), .QN(n14477) );
  NAND2X0 U15719 ( .IN1(n14149), .IN2(g429), .QN(n14476) );
  NAND2X0 U15720 ( .IN1(n14478), .IN2(n14479), .QN(g24202) );
  NAND2X0 U15721 ( .IN1(n12923), .IN2(g424), .QN(n14479) );
  NAND2X0 U15722 ( .IN1(n14149), .IN2(g411), .QN(n14478) );
  NAND2X0 U15723 ( .IN1(n14480), .IN2(n14481), .QN(g24201) );
  NAND2X0 U15724 ( .IN1(n12923), .IN2(g405), .QN(n14481) );
  NAND2X0 U15725 ( .IN1(n14149), .IN2(g392), .QN(n14480) );
  NAND3X0 U15726 ( .IN1(n14482), .IN2(n14483), .IN3(n14484), .QN(g24200) );
  NAND2X0 U15727 ( .IN1(n8573), .IN2(g401), .QN(n14484) );
  NAND3X0 U15728 ( .IN1(n5821), .IN2(g854), .IN3(n12927), .QN(n14483) );
  INVX0 U15729 ( .INP(n14148), .ZN(n12927) );
  NAND2X0 U15730 ( .IN1(n4948), .IN2(n8513), .QN(n14148) );
  NAND2X0 U15731 ( .IN1(n12923), .IN2(g392), .QN(n14482) );
  INVX0 U15732 ( .INP(n14149), .ZN(n12923) );
  NAND2X0 U15733 ( .IN1(n8510), .IN2(n12926), .QN(n14149) );
  INVX0 U15734 ( .INP(n4948), .ZN(n12926) );
  NOR2X0 U15735 ( .IN1(g22), .IN2(g25), .QN(g23190) );
  NAND2X0 U15736 ( .IN1(n14485), .IN2(n14486), .QN(g21901) );
  NAND2X0 U15737 ( .IN1(n8574), .IN2(g2946), .QN(n14486) );
  NAND2X0 U15738 ( .IN1(n14487), .IN2(n8513), .QN(n14485) );
  NAND2X0 U15739 ( .IN1(n14488), .IN2(n14489), .QN(n14487) );
  NAND2X0 U15740 ( .IN1(n5694), .IN2(g4180), .QN(n14489) );
  NAND2X0 U15741 ( .IN1(n5380), .IN2(n14490), .QN(n14488) );
  NAND2X0 U15742 ( .IN1(n5694), .IN2(n14491), .QN(n14490) );
  NAND4X0 U15743 ( .IN1(n14527), .IN2(n7854), .IN3(n14526), .IN4(n14492), .QN(
        n14491) );
  NOR4X0 U15744 ( .IN1(test_so86), .IN2(test_so39), .IN3(g8787), .IN4(g8788), 
        .QN(n14492) );
  NAND2X0 U15745 ( .IN1(n14493), .IN2(n14494), .QN(g21900) );
  OR2X1 U15746 ( .IN1(n8481), .IN2(n7797), .Q(n14494) );
  NAND3X0 U15747 ( .IN1(n7727), .IN2(n7726), .IN3(n8493), .QN(n14493) );
  XOR2X1 U15748 ( .IN1(n14495), .IN2(n8189), .Q(g21899) );
  NAND2X0 U15749 ( .IN1(n8511), .IN2(g9019), .QN(n14495) );
  NAND2X0 U15750 ( .IN1(n14496), .IN2(n14497), .QN(g21898) );
  NAND2X0 U15751 ( .IN1(n8189), .IN2(n8513), .QN(n14497) );
  OR2X1 U15752 ( .IN1(n8481), .IN2(n7812), .Q(n14496) );
  XOR2X1 U15753 ( .IN1(n14498), .IN2(n8190), .Q(g21897) );
  NAND2X0 U15754 ( .IN1(n8511), .IN2(g8839), .QN(n14498) );
  NAND2X0 U15755 ( .IN1(n14499), .IN2(n14500), .QN(g21896) );
  NAND2X0 U15756 ( .IN1(n8190), .IN2(n8513), .QN(n14500) );
  NAND2X0 U15757 ( .IN1(n8575), .IN2(g4245), .QN(n14499) );
  NAND2X0 U15758 ( .IN1(n14501), .IN2(n14502), .QN(g21895) );
  NAND2X0 U15759 ( .IN1(n14503), .IN2(g4264), .QN(n14502) );
  NAND2X0 U15760 ( .IN1(n14504), .IN2(n8513), .QN(n14503) );
  NAND2X0 U15761 ( .IN1(n5763), .IN2(g4258), .QN(n14504) );
  OR2X1 U15762 ( .IN1(n14295), .IN2(n5763), .Q(n14501) );
  NOR2X0 U15763 ( .IN1(g21893), .IN2(n14505), .QN(n14295) );
  NOR2X0 U15764 ( .IN1(g4264), .IN2(n8561), .QN(n14505) );
  NAND2X0 U15765 ( .IN1(n14506), .IN2(n14507), .QN(g21894) );
  NAND2X0 U15766 ( .IN1(n14508), .IN2(g4258), .QN(n14507) );
  NAND2X0 U15767 ( .IN1(n8511), .IN2(g4264), .QN(n14508) );
  NAND2X0 U15768 ( .IN1(g21893), .IN2(g4264), .QN(n14506) );
  NOR2X0 U15769 ( .IN1(g4258), .IN2(n8564), .QN(g21893) );
  NAND2X0 U15770 ( .IN1(n14509), .IN2(n14510), .QN(g21892) );
  NAND2X0 U15771 ( .IN1(n7797), .IN2(n8513), .QN(n14510) );
  NAND2X0 U15772 ( .IN1(n8577), .IN2(g4273), .QN(n14509) );
  NAND2X0 U15773 ( .IN1(n14511), .IN2(n14512), .QN(g21891) );
  NAND2X0 U15774 ( .IN1(n8539), .IN2(g4180), .QN(n14512) );
  NAND2X0 U15775 ( .IN1(n14301), .IN2(n8513), .QN(n14511) );
  NAND2X0 U15776 ( .IN1(n14513), .IN2(n14514), .QN(n14301) );
  NAND2X0 U15777 ( .IN1(n8161), .IN2(g4253), .QN(n14514) );
  NAND2X0 U15778 ( .IN1(n8160), .IN2(n5484), .QN(n14513) );
  NOR2X0 U15779 ( .IN1(n8506), .IN2(DFF_1381_n1), .QN(g21727) );
  NOR2X0 U15780 ( .IN1(n5750), .IN2(n8504), .QN(g18597) );
  INVX0 U15781 ( .INP(g5), .ZN(g12833) );
  OR2X1 U5116_U1 ( .IN1(g34783), .IN2(n2730), .Q(g34221) );
  OR2X1 U5126_U1 ( .IN1(n4836), .IN2(n4896), .Q(n4895) );
  OR2X1 U5127_U1 ( .IN1(n4837), .IN2(n4921), .Q(n4920) );
  OR2X1 U5128_U1 ( .IN1(n628), .IN2(n4411), .Q(n5045) );
  OR2X1 U5129_U1 ( .IN1(g559), .IN2(g9048), .Q(n4959) );
  INVX0 U5353_U2 ( .INP(n5960), .ZN(U5353_n1) );
  NOR2X0 U5353_U1 ( .IN1(n8198), .IN2(U5353_n1), .QN(n4689) );
  INVX0 U5355_U2 ( .INP(n5961), .ZN(U5355_n1) );
  NOR2X0 U5355_U1 ( .IN1(n8196), .IN2(U5355_n1), .QN(n4708) );
  INVX0 U5961_U2 ( .INP(n3593), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n3589), .IN2(U5961_n1), .QN(n3595) );
  INVX0 U5962_U2 ( .INP(n3574), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n3570), .IN2(U5962_n1), .QN(n3576) );
  INVX0 U5963_U2 ( .INP(n3517), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n3513), .IN2(U5963_n1), .QN(n3519) );
  INVX0 U5964_U2 ( .INP(n3628), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n3624), .IN2(U5964_n1), .QN(n3630) );
  INVX0 U5965_U2 ( .INP(n3555), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n3551), .IN2(U5965_n1), .QN(n3557) );
  INVX0 U5966_U2 ( .INP(n3646), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n3642), .IN2(U5966_n1), .QN(n3648) );
  INVX0 U5967_U2 ( .INP(n3536), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n3532), .IN2(U5967_n1), .QN(n3538) );
  INVX0 U5968_U2 ( .INP(n3611), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n3607), .IN2(U5968_n1), .QN(n3613) );
  INVX0 U6100_U2 ( .INP(n3635), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n8564), .IN2(U6100_n1), .QN(n4888) );
  INVX0 U6211_U2 ( .INP(n3623), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n1413), .IN2(U6211_n1), .QN(n3622) );
  INVX0 U6212_U2 ( .INP(n3587), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n3588), .IN2(U6212_n1), .QN(n3586) );
  INVX0 U6213_U2 ( .INP(n3605), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n3606), .IN2(U6213_n1), .QN(n3604) );
  INVX0 U6214_U2 ( .INP(n3568), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n3569), .IN2(U6214_n1), .QN(n3567) );
  INVX0 U6215_U2 ( .INP(n3549), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n3550), .IN2(U6215_n1), .QN(n3548) );
  INVX0 U6216_U2 ( .INP(n3512), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n3006), .IN2(U6216_n1), .QN(n3511) );
  INVX0 U6217_U2 ( .INP(n3531), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n3007), .IN2(U6217_n1), .QN(n3530) );
  INVX0 U6218_U2 ( .INP(n3641), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n3003), .IN2(U6218_n1), .QN(n3640) );
  INVX0 U6279_U2 ( .INP(n4537), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n5337), .IN2(U6279_n1), .QN(n4201) );
  INVX0 U6280_U2 ( .INP(n4201), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n5336), .IN2(U6280_n1), .QN(n3745) );
  INVX0 U6281_U2 ( .INP(n3745), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n5294), .IN2(U6281_n1), .QN(n3684) );
  INVX0 U6282_U2 ( .INP(n3684), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n5552), .IN2(U6282_n1), .QN(n3274) );
  INVX0 U6283_U2 ( .INP(n3274), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n5472), .IN2(U6283_n1), .QN(n2982) );
  INVX0 U6284_U2 ( .INP(n2982), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n5476), .IN2(U6284_n1), .QN(n2706) );
  INVX0 U6285_U2 ( .INP(n2706), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n5550), .IN2(U6285_n1), .QN(n2649) );
  INVX0 U6286_U2 ( .INP(n2649), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n5473), .IN2(U6286_n1), .QN(n2556) );
  INVX0 U6287_U2 ( .INP(n2556), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n5475), .IN2(U6287_n1), .QN(n2509) );
  INVX0 U6288_U2 ( .INP(n2509), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n5474), .IN2(U6288_n1), .QN(n2487) );
  INVX0 U6289_U2 ( .INP(n2487), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n5339), .IN2(U6289_n1), .QN(n2427) );
  INVX0 U6290_U2 ( .INP(n2427), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n5672), .IN2(U6290_n1), .QN(n2423) );
  INVX0 U6291_U2 ( .INP(n5), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n5335), .IN2(U6291_n1), .QN(n4537) );
  INVX0 U6292_U2 ( .INP(n4959), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n8565), .IN2(U6292_n1), .QN(n2421) );
  INVX0 U6338_U2 ( .INP(n4210), .ZN(U6338_n1) );
  NOR2X1 U6338_U1 ( .IN1(n8565), .IN2(U6338_n1), .QN(n3765) );
  INVX0 U6341_U2 ( .INP(n3765), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n3479), .IN2(U6341_n1), .QN(n3951) );
  INVX0 U6342_U2 ( .INP(n3765), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n3404), .IN2(U6342_n1), .QN(n3774) );
  INVX0 U6343_U2 ( .INP(n3765), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n3424), .IN2(U6343_n1), .QN(n3842) );
  INVX0 U6344_U2 ( .INP(n3765), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n3414), .IN2(U6344_n1), .QN(n3808) );
  INVX0 U6345_U2 ( .INP(n3765), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n3444), .IN2(U6345_n1), .QN(n3908) );
  INVX0 U6346_U2 ( .INP(n3765), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n3489), .IN2(U6346_n1), .QN(n3984) );
  INVX0 U6347_U2 ( .INP(n3765), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n3434), .IN2(U6347_n1), .QN(n3875) );
  INVX0 U6348_U2 ( .INP(n3765), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n3500), .IN2(U6348_n1), .QN(n4015) );
  INVX0 U6349_U2 ( .INP(n3765), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n3446), .IN2(U6349_n1), .QN(n3914) );
  INVX0 U6350_U2 ( .INP(n3765), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n3406), .IN2(U6350_n1), .QN(n3780) );
  INVX0 U6351_U2 ( .INP(n3765), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n3481), .IN2(U6351_n1), .QN(n3957) );
  INVX0 U6352_U2 ( .INP(n3765), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n3426), .IN2(U6352_n1), .QN(n3848) );
  INVX0 U6353_U2 ( .INP(n3765), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n3491), .IN2(U6353_n1), .QN(n3990) );
  INVX0 U6354_U2 ( .INP(n3765), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n3416), .IN2(U6354_n1), .QN(n3814) );
  INVX0 U6355_U2 ( .INP(n3765), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n3436), .IN2(U6355_n1), .QN(n3881) );
  INVX0 U6356_U2 ( .INP(n3765), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n3502), .IN2(U6356_n1), .QN(n4022) );
  INVX0 U6357_U2 ( .INP(n3765), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n3501), .IN2(U6357_n1), .QN(n4027) );
  INVX0 U6358_U2 ( .INP(n3765), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n3407), .IN2(U6358_n1), .QN(n3785) );
  INVX0 U6359_U2 ( .INP(n3765), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n3482), .IN2(U6359_n1), .QN(n3962) );
  INVX0 U6360_U2 ( .INP(n3765), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n3427), .IN2(U6360_n1), .QN(n3853) );
  INVX0 U6361_U2 ( .INP(n3765), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n3437), .IN2(U6361_n1), .QN(n3886) );
  INVX0 U6362_U2 ( .INP(n3765), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n3417), .IN2(U6362_n1), .QN(n3819) );
  INVX0 U6363_U2 ( .INP(n3765), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n3492), .IN2(U6363_n1), .QN(n3995) );
  INVX0 U6364_U2 ( .INP(n3765), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n3447), .IN2(U6364_n1), .QN(n3919) );
  INVX0 U6365_U2 ( .INP(n3682), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n5471), .IN2(U6365_n1), .QN(n3272) );
  INVX0 U6366_U2 ( .INP(n3272), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n5331), .IN2(U6366_n1), .QN(n2980) );
  INVX0 U6367_U2 ( .INP(n2980), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n5332), .IN2(U6367_n1), .QN(n2704) );
  INVX0 U6368_U2 ( .INP(n2704), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n5333), .IN2(U6368_n1), .QN(n2647) );
  INVX0 U6369_U2 ( .INP(n2647), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n5334), .IN2(U6369_n1), .QN(n2554) );
  INVX0 U6370_U2 ( .INP(n2554), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n5330), .IN2(U6370_n1), .QN(n2507) );
  INVX0 U6371_U2 ( .INP(n2507), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n5551), .IN2(U6371_n1), .QN(n2485) );
  INVX0 U6372_U2 ( .INP(n2485), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n5293), .IN2(U6372_n1), .QN(n2425) );
  INVX0 U6373_U2 ( .INP(n2425), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n5292), .IN2(U6373_n1), .QN(n2419) );
  INVX0 U6374_U2 ( .INP(n43), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n5470), .IN2(U6374_n1), .QN(n3682) );
  INVX0 U6375_U2 ( .INP(n2419), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n5291), .IN2(U6375_n1), .QN(n2405) );
  INVX0 U6417_U2 ( .INP(n4198), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n8567), .IN2(U6417_n1), .QN(n2404) );
  INVX0 U6446_U2 ( .INP(g110), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n1430), .IN2(U6446_n1), .QN(n3524) );
  INVX0 U6465_U2 ( .INP(n3653), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n5600), .IN2(U6465_n1), .QN(n4388) );
  INVX0 U6497_U2 ( .INP(n3581), .ZN(U6497_n1) );
  NOR2X0 U6497_U1 ( .IN1(n3635), .IN2(U6497_n1), .QN(n3005) );
  INVX0 U6523_U2 ( .INP(n4946), .ZN(U6523_n1) );
  NOR2X0 U6523_U1 ( .IN1(n8564), .IN2(U6523_n1), .QN(n4945) );
  INVX0 U6542_U2 ( .INP(n3581), .ZN(U6542_n1) );
  NOR2X0 U6542_U1 ( .IN1(n5300), .IN2(U6542_n1), .QN(n3525) );
  INVX0 U6552_U2 ( .INP(n3281), .ZN(U6552_n1) );
  NOR2X0 U6552_U1 ( .IN1(n5676), .IN2(U6552_n1), .QN(n3277) );
  INVX0 U6553_U2 ( .INP(n3276), .ZN(U6553_n1) );
  NOR2X0 U6553_U1 ( .IN1(n5680), .IN2(U6553_n1), .QN(n2989) );
  INVX0 U6554_U2 ( .INP(n3277), .ZN(U6554_n1) );
  NOR2X0 U6554_U1 ( .IN1(n5677), .IN2(U6554_n1), .QN(n2991) );
  INVX0 U6555_U2 ( .INP(n45), .ZN(U6555_n1) );
  NOR2X0 U6555_U1 ( .IN1(n5561), .IN2(U6555_n1), .QN(n3281) );
  INVX0 U6556_U2 ( .INP(n42), .ZN(U6556_n1) );
  NOR2X0 U6556_U1 ( .IN1(n5679), .IN2(U6556_n1), .QN(n3276) );
  INVX0 U6559_U2 ( .INP(n2991), .ZN(U6559_n1) );
  NOR2X0 U6559_U1 ( .IN1(n5678), .IN2(U6559_n1), .QN(n2710) );
  INVX0 U6560_U2 ( .INP(n2989), .ZN(U6560_n1) );
  NOR2X0 U6560_U1 ( .IN1(n5675), .IN2(U6560_n1), .QN(n2707) );
  INVX0 U6561_U2 ( .INP(n3174), .ZN(U6561_n1) );
  NOR2X0 U6561_U1 ( .IN1(n5327), .IN2(U6561_n1), .QN(n3116) );
  INVX0 U6570_U2 ( .INP(n3362), .ZN(U6570_n1) );
  NOR2X0 U6570_U1 ( .IN1(n5477), .IN2(U6570_n1), .QN(n2527) );
  INVX0 U6911_U2 ( .INP(n3115), .ZN(U6911_n1) );
  NOR2X0 U6911_U1 ( .IN1(n2726), .IN2(U6911_n1), .QN(n3111) );
  INVX0 U6912_U2 ( .INP(n3115), .ZN(U6912_n1) );
  NOR2X0 U6912_U1 ( .IN1(n2727), .IN2(U6912_n1), .QN(n3131) );
  INVX0 U6917_U2 ( .INP(n3933), .ZN(U6917_n1) );
  NOR2X0 U6917_U1 ( .IN1(n5350), .IN2(U6917_n1), .QN(n3799) );
  INVX0 U6926_U2 ( .INP(n3664), .ZN(U6926_n1) );
  NOR2X0 U6926_U1 ( .IN1(n5674), .IN2(U6926_n1), .QN(n3662) );
  INVX0 U6927_U2 ( .INP(n3673), .ZN(U6927_n1) );
  NOR2X0 U6927_U1 ( .IN1(n5673), .IN2(U6927_n1), .QN(n3671) );
  INVX0 U6929_U2 ( .INP(n3505), .ZN(U6929_n1) );
  NOR2X0 U6929_U1 ( .IN1(n3506), .IN2(U6929_n1), .QN(n2790) );
  INVX0 U6931_U2 ( .INP(n4490), .ZN(U6931_n1) );
  NOR2X0 U6931_U1 ( .IN1(n5554), .IN2(U6931_n1), .QN(n4178) );
  INVX0 U6932_U2 ( .INP(n4514), .ZN(U6932_n1) );
  NOR2X0 U6932_U1 ( .IN1(n5555), .IN2(U6932_n1), .QN(n4196) );
  INVX0 U6933_U2 ( .INP(n4178), .ZN(U6933_n1) );
  NOR2X0 U6933_U1 ( .IN1(n5558), .IN2(U6933_n1), .QN(n3736) );
  INVX0 U6934_U2 ( .INP(n4196), .ZN(U6934_n1) );
  NOR2X0 U6934_U1 ( .IN1(n5559), .IN2(U6934_n1), .QN(n3741) );
  INVX0 U6935_U2 ( .INP(n3736), .ZN(U6935_n1) );
  NOR2X0 U6935_U1 ( .IN1(n5553), .IN2(U6935_n1), .QN(n3664) );
  INVX0 U6936_U2 ( .INP(n3741), .ZN(U6936_n1) );
  NOR2X0 U6936_U1 ( .IN1(n5560), .IN2(U6936_n1), .QN(n3673) );
  INVX0 U6937_U2 ( .INP(n2601), .ZN(U6937_n1) );
  NOR2X0 U6937_U1 ( .IN1(n5303), .IN2(U6937_n1), .QN(n2598) );
  INVX0 U6938_U2 ( .INP(n965), .ZN(U6938_n1) );
  NOR2X0 U6938_U1 ( .IN1(n5556), .IN2(U6938_n1), .QN(n4490) );
  INVX0 U6939_U2 ( .INP(n220), .ZN(U6939_n1) );
  NOR2X0 U6939_U1 ( .IN1(n5557), .IN2(U6939_n1), .QN(n4514) );
  INVX0 U6940_U2 ( .INP(n4814), .ZN(U6940_n1) );
  NOR2X0 U6940_U1 ( .IN1(n5422), .IN2(U6940_n1), .QN(n4519) );
  INVX0 U6941_U2 ( .INP(n2607), .ZN(U6941_n1) );
  NOR2X0 U6941_U1 ( .IN1(n5323), .IN2(U6941_n1), .QN(n2594) );
  INVX0 U6944_U2 ( .INP(n3084), .ZN(U6944_n1) );
  NOR2X0 U6944_U1 ( .IN1(n5348), .IN2(U6944_n1), .QN(n3033) );
  INVX0 U6950_U2 ( .INP(n2598), .ZN(U6950_n1) );
  NOR2X0 U6950_U1 ( .IN1(n5365), .IN2(U6950_n1), .QN(n2590) );
  INVX0 U6954_U2 ( .INP(n3122), .ZN(U6954_n1) );
  NOR2X0 U6954_U1 ( .IN1(n2727), .IN2(U6954_n1), .QN(n3125) );
  INVX0 U6955_U2 ( .INP(n3102), .ZN(U6955_n1) );
  NOR2X0 U6955_U1 ( .IN1(n2726), .IN2(U6955_n1), .QN(n3105) );
  INVX0 U6956_U2 ( .INP(n3141), .ZN(U6956_n1) );
  NOR2X0 U6956_U1 ( .IN1(n3146), .IN2(U6956_n1), .QN(n3145) );
  INVX0 U6957_U2 ( .INP(n3160), .ZN(U6957_n1) );
  NOR2X0 U6957_U1 ( .IN1(n3165), .IN2(U6957_n1), .QN(n3164) );
  INVX0 U7174_U2 ( .INP(n2423), .ZN(U7174_n1) );
  NOR2X0 U7174_U1 ( .IN1(n5288), .IN2(U7174_n1), .QN(n2422) );
  INVX0 U7248_U2 ( .INP(n4172), .ZN(U7248_n1) );
  NOR2X0 U7248_U1 ( .IN1(g1536), .IN2(U7248_n1), .QN(n4173) );
  INVX0 U7249_U2 ( .INP(n4190), .ZN(U7249_n1) );
  NOR2X0 U7249_U1 ( .IN1(g1193), .IN2(U7249_n1), .QN(n4191) );
  INVX0 U7402_U2 ( .INP(n4034), .ZN(U7402_n1) );
  NOR2X0 U7402_U1 ( .IN1(n4020), .IN2(U7402_n1), .QN(n4037) );
  INVX0 U7405_U2 ( .INP(n4034), .ZN(U7405_n1) );
  NOR2X0 U7405_U1 ( .IN1(n4014), .IN2(U7405_n1), .QN(n4039) );
  INVX0 U7413_U2 ( .INP(n3969), .ZN(U7413_n1) );
  NOR2X0 U7413_U1 ( .IN1(n3947), .IN2(U7413_n1), .QN(n3972) );
  INVX0 U7416_U2 ( .INP(n3926), .ZN(U7416_n1) );
  NOR2X0 U7416_U1 ( .IN1(n3904), .IN2(U7416_n1), .QN(n3929) );
  INVX0 U7427_U2 ( .INP(n3860), .ZN(U7427_n1) );
  NOR2X0 U7427_U1 ( .IN1(n3838), .IN2(U7427_n1), .QN(n3863) );
  INVX0 U7438_U2 ( .INP(n4002), .ZN(U7438_n1) );
  NOR2X0 U7438_U1 ( .IN1(n3978), .IN2(U7438_n1), .QN(n4003) );
  INVX0 U7449_U2 ( .INP(n4034), .ZN(U7449_n1) );
  NOR2X0 U7449_U1 ( .IN1(n4017), .IN2(U7449_n1), .QN(n4032) );
  INVX0 U7455_U2 ( .INP(n4034), .ZN(U7455_n1) );
  NOR2X0 U7455_U1 ( .IN1(n3495), .IN2(U7455_n1), .QN(n4035) );
  INVX0 U7464_U2 ( .INP(n3792), .ZN(U7464_n1) );
  NOR2X0 U7464_U1 ( .IN1(n3773), .IN2(U7464_n1), .QN(n3797) );
  INVX0 U7467_U2 ( .INP(n3792), .ZN(U7467_n1) );
  NOR2X0 U7467_U1 ( .IN1(n3776), .IN2(U7467_n1), .QN(n3790) );
  INVX0 U7482_U2 ( .INP(n3792), .ZN(U7482_n1) );
  NOR2X0 U7482_U1 ( .IN1(n3770), .IN2(U7482_n1), .QN(n3795) );
  INVX0 U7492_U2 ( .INP(n3893), .ZN(U7492_n1) );
  NOR2X0 U7492_U1 ( .IN1(n3877), .IN2(U7492_n1), .QN(n3891) );
  INVX0 U7513_U2 ( .INP(n3826), .ZN(U7513_n1) );
  NOR2X0 U7513_U1 ( .IN1(n3802), .IN2(U7513_n1), .QN(n3827) );
  INVX0 U7516_U2 ( .INP(n3893), .ZN(U7516_n1) );
  NOR2X0 U7516_U1 ( .IN1(n3871), .IN2(U7516_n1), .QN(n3896) );
  INVX0 U7549_U2 ( .INP(n4002), .ZN(U7549_n1) );
  NOR2X0 U7549_U1 ( .IN1(n3983), .IN2(U7549_n1), .QN(n4007) );
  INVX0 U7561_U2 ( .INP(n3926), .ZN(U7561_n1) );
  NOR2X0 U7561_U1 ( .IN1(n3907), .IN2(U7561_n1), .QN(n3931) );
  INVX0 U7574_U2 ( .INP(n3792), .ZN(U7574_n1) );
  NOR2X0 U7574_U1 ( .IN1(n3768), .IN2(U7574_n1), .QN(n3793) );
  INVX0 U7577_U2 ( .INP(n3926), .ZN(U7577_n1) );
  NOR2X0 U7577_U1 ( .IN1(n3910), .IN2(U7577_n1), .QN(n3924) );
  INVX0 U7585_U2 ( .INP(n3826), .ZN(U7585_n1) );
  NOR2X0 U7585_U1 ( .IN1(n3807), .IN2(U7585_n1), .QN(n3831) );
  INVX0 U7595_U2 ( .INP(n3826), .ZN(U7595_n1) );
  NOR2X0 U7595_U1 ( .IN1(n3804), .IN2(U7595_n1), .QN(n3829) );
  INVX0 U7614_U2 ( .INP(n3926), .ZN(U7614_n1) );
  NOR2X0 U7614_U1 ( .IN1(n3902), .IN2(U7614_n1), .QN(n3927) );
  INVX0 U7621_U2 ( .INP(n3969), .ZN(U7621_n1) );
  NOR2X0 U7621_U1 ( .IN1(n3950), .IN2(U7621_n1), .QN(n3974) );
  INVX0 U7629_U2 ( .INP(n3893), .ZN(U7629_n1) );
  NOR2X0 U7629_U1 ( .IN1(n3874), .IN2(U7629_n1), .QN(n3898) );
  INVX0 U7636_U2 ( .INP(n3969), .ZN(U7636_n1) );
  NOR2X0 U7636_U1 ( .IN1(n3945), .IN2(U7636_n1), .QN(n3970) );
  INVX0 U7639_U2 ( .INP(n4002), .ZN(U7639_n1) );
  NOR2X0 U7639_U1 ( .IN1(n3986), .IN2(U7639_n1), .QN(n4000) );
  INVX0 U7649_U2 ( .INP(n3860), .ZN(U7649_n1) );
  NOR2X0 U7649_U1 ( .IN1(n3841), .IN2(U7649_n1), .QN(n3865) );
  INVX0 U7652_U2 ( .INP(n3860), .ZN(U7652_n1) );
  NOR2X0 U7652_U1 ( .IN1(n3836), .IN2(U7652_n1), .QN(n3861) );
  INVX0 U7668_U2 ( .INP(n3826), .ZN(U7668_n1) );
  NOR2X0 U7668_U1 ( .IN1(n3810), .IN2(U7668_n1), .QN(n3824) );
  INVX0 U7673_U2 ( .INP(n3893), .ZN(U7673_n1) );
  NOR2X0 U7673_U1 ( .IN1(n3869), .IN2(U7673_n1), .QN(n3894) );
  INVX0 U7690_U2 ( .INP(n3969), .ZN(U7690_n1) );
  NOR2X0 U7690_U1 ( .IN1(n3953), .IN2(U7690_n1), .QN(n3967) );
  INVX0 U7707_U2 ( .INP(n3860), .ZN(U7707_n1) );
  NOR2X0 U7707_U1 ( .IN1(n3844), .IN2(U7707_n1), .QN(n3858) );
  INVX0 U7712_U2 ( .INP(n4002), .ZN(U7712_n1) );
  NOR2X0 U7712_U1 ( .IN1(n3980), .IN2(U7712_n1), .QN(n4005) );
  INVX0 U7792_U2 ( .INP(g952), .ZN(U7792_n1) );
  NOR2X0 U7792_U1 ( .IN1(n8565), .IN2(U7792_n1), .QN(n2505) );
  INVX0 U7794_U2 ( .INP(g1296), .ZN(U7794_n1) );
  NOR2X0 U7794_U1 ( .IN1(n8566), .IN2(U7794_n1), .QN(n2499) );
  INVX0 U7895_U2 ( .INP(n2668), .ZN(U7895_n1) );
  NOR2X0 U7895_U1 ( .IN1(g113), .IN2(U7895_n1), .QN(n2760) );
  INVX0 U7897_U2 ( .INP(g6), .ZN(U7897_n1) );
  NOR2X0 U7897_U1 ( .IN1(g31), .IN2(U7897_n1), .QN(n3395) );
  INVX0 U7977_U2 ( .INP(g661), .ZN(U7977_n1) );
  NOR2X0 U7977_U1 ( .IN1(n8567), .IN2(U7977_n1), .QN(n4956) );
  INVX0 U8034_U2 ( .INP(n4723), .ZN(U8034_n1) );
  NOR2X0 U8034_U1 ( .IN1(n5612), .IN2(U8034_n1), .QN(n5026) );
  INVX0 U8036_U2 ( .INP(n3729), .ZN(U8036_n1) );
  NOR2X0 U8036_U1 ( .IN1(n5340), .IN2(U8036_n1), .QN(n3941) );
  INVX0 U8050_U2 ( .INP(n155), .ZN(U8050_n1) );
  NOR2X0 U8050_U1 ( .IN1(g1367), .IN2(U8050_n1), .QN(n3733) );
  INVX0 U8055_U2 ( .INP(g1345), .ZN(U8055_n1) );
  NOR2X0 U8055_U1 ( .IN1(n8566), .IN2(U8055_n1), .QN(n4798) );
  INVX0 U8060_U2 ( .INP(g1002), .ZN(U8060_n1) );
  NOR2X0 U8060_U1 ( .IN1(n8565), .IN2(U8060_n1), .QN(n4805) );
  INVX0 U8070_U2 ( .INP(n156), .ZN(U8070_n1) );
  NOR2X0 U8070_U1 ( .IN1(g1361), .IN2(U8070_n1), .QN(n4175) );
  INVX0 U8074_U2 ( .INP(n436), .ZN(U8074_n1) );
  NOR2X0 U8074_U1 ( .IN1(g1018), .IN2(U8074_n1), .QN(n4193) );
  INVX0 U8088_U2 ( .INP(n435), .ZN(U8088_n1) );
  NOR2X0 U8088_U1 ( .IN1(g1024), .IN2(U8088_n1), .QN(n3738) );
  INVX0 U8112_U2 ( .INP(n4525), .ZN(U8112_n1) );
  NOR2X0 U8112_U1 ( .IN1(n4523), .IN2(U8112_n1), .QN(n4524) );
  INVX0 U8113_U2 ( .INP(n4526), .ZN(U8113_n1) );
  NOR2X0 U8113_U1 ( .IN1(n5751), .IN2(U8113_n1), .QN(n4523) );
  INVX0 U8147_U2 ( .INP(g4659), .ZN(U8147_n1) );
  NOR2X0 U8147_U1 ( .IN1(n2573), .IN2(U8147_n1), .QN(n2577) );
  INVX0 U8165_U2 ( .INP(g4849), .ZN(U8165_n1) );
  NOR2X0 U8165_U1 ( .IN1(n2563), .IN2(U8165_n1), .QN(n2567) );
  INVX0 U8185_U2 ( .INP(n4940), .ZN(U8185_n1) );
  NOR2X0 U8185_U1 ( .IN1(g1046), .IN2(U8185_n1), .QN(n4938) );
  INVX0 U8192_U2 ( .INP(n4915), .ZN(U8192_n1) );
  NOR2X0 U8192_U1 ( .IN1(g1389), .IN2(U8192_n1), .QN(n4913) );
  INVX0 U8210_U2 ( .INP(n4722), .ZN(U8210_n1) );
  NOR2X0 U8210_U1 ( .IN1(n4723), .IN2(U8210_n1), .QN(n4714) );
  INVX0 U8223_U2 ( .INP(n4518), .ZN(U8223_n1) );
  NOR2X0 U8223_U1 ( .IN1(n4516), .IN2(U8223_n1), .QN(n4517) );
  INVX0 U8224_U2 ( .INP(n4519), .ZN(U8224_n1) );
  NOR2X0 U8224_U1 ( .IN1(n5728), .IN2(U8224_n1), .QN(n4516) );
  INVX0 U8281_U2 ( .INP(n4819), .ZN(U8281_n1) );
  NOR2X0 U8281_U1 ( .IN1(n8566), .IN2(U8281_n1), .QN(n5111) );
  INVX0 U8307_U2 ( .INP(g29216), .ZN(U8307_n1) );
  NOR2X0 U8307_U1 ( .IN1(n8568), .IN2(U8307_n1), .QN(g26900) );
  INVX0 U8974_U2 ( .INP(n3362), .ZN(U8974_n1) );
  NOR2X0 U8974_U1 ( .IN1(test_so25), .IN2(U8974_n1), .QN(n2552) );
  INVX0 U8975_U2 ( .INP(n3174), .ZN(U8975_n1) );
  NOR2X0 U8975_U1 ( .IN1(g528), .IN2(U8975_n1), .QN(n3195) );
  INVX0 U9065_U2 ( .INP(g4145), .ZN(U9065_n1) );
  NOR2X0 U9065_U1 ( .IN1(n8567), .IN2(U9065_n1), .QN(n4721) );
  INVX0 U9070_U2 ( .INP(g2841), .ZN(U9070_n1) );
  NOR2X0 U9070_U1 ( .IN1(n8566), .IN2(U9070_n1), .QN(n3730) );
  INVX0 U9075_U2 ( .INP(g19), .ZN(U9075_n1) );
  NOR2X0 U9075_U1 ( .IN1(g9), .IN2(U9075_n1), .QN(n3362) );
  INVX0 U9076_U2 ( .INP(g113), .ZN(U9076_n1) );
  NOR2X0 U9076_U1 ( .IN1(n8568), .IN2(U9076_n1), .QN(g25694) );
  INVX0 U9080_U2 ( .INP(n4305), .ZN(U9080_n1) );
  NOR2X0 U9080_U1 ( .IN1(n8565), .IN2(U9080_n1), .QN(g29277) );
  INVX0 U9084_U2 ( .INP(g4423), .ZN(U9084_n1) );
  NOR2X0 U9084_U1 ( .IN1(n8567), .IN2(U9084_n1), .QN(g26953) );
  INVX0 U9085_U2 ( .INP(g64), .ZN(U9085_n1) );
  NOR2X0 U9085_U1 ( .IN1(n8568), .IN2(U9085_n1), .QN(g24212) );
  INVX0 U9086_U2 ( .INP(n4283), .ZN(U9086_n1) );
  NOR2X0 U9086_U1 ( .IN1(n8566), .IN2(U9086_n1), .QN(g29279) );
  INVX0 U9090_U2 ( .INP(g125), .ZN(U9090_n1) );
  NOR2X0 U9090_U1 ( .IN1(n8568), .IN2(U9090_n1), .QN(g25688) );
  INVX0 U9098_U2 ( .INP(g4681), .ZN(U9098_n1) );
  NOR2X0 U9098_U1 ( .IN1(n2774), .IN2(U9098_n1), .QN(g34028) );
  INVX0 U9099_U2 ( .INP(n2595), .ZN(U9099_n1) );
  NOR2X0 U9099_U1 ( .IN1(n2608), .IN2(U9099_n1), .QN(g34449) );
  INVX0 U9101_U2 ( .INP(g6745), .ZN(U9101_n1) );
  NOR2X0 U9101_U1 ( .IN1(n8567), .IN2(U9101_n1), .QN(g26880) );
  INVX0 U9107_U2 ( .INP(n4448), .ZN(U9107_n1) );
  NOR2X0 U9107_U1 ( .IN1(n709), .IN2(U9107_n1), .QN(n4447) );
  INVX0 U9111_U2 ( .INP(n4403), .ZN(U9111_n1) );
  NOR2X0 U9111_U1 ( .IN1(n456), .IN2(U9111_n1), .QN(n4402) );
  INVX0 U9116_U2 ( .INP(n4426), .ZN(U9116_n1) );
  NOR2X0 U9116_U1 ( .IN1(n1136), .IN2(U9116_n1), .QN(n4425) );
  INVX0 U9120_U2 ( .INP(n4437), .ZN(U9120_n1) );
  NOR2X0 U9120_U1 ( .IN1(n314), .IN2(U9120_n1), .QN(n4436) );
  INVX0 U9124_U2 ( .INP(n4392), .ZN(U9124_n1) );
  NOR2X0 U9124_U1 ( .IN1(n911), .IN2(U9124_n1), .QN(n4391) );
  INVX0 U9128_U2 ( .INP(n4380), .ZN(U9128_n1) );
  NOR2X0 U9128_U1 ( .IN1(n326), .IN2(U9128_n1), .QN(n4379) );
  INVX0 U9132_U2 ( .INP(n4415), .ZN(U9132_n1) );
  NOR2X0 U9132_U1 ( .IN1(n982), .IN2(U9132_n1), .QN(n4414) );
  INVX0 U9136_U2 ( .INP(n4459), .ZN(U9136_n1) );
  NOR2X0 U9136_U1 ( .IN1(n1123), .IN2(U9136_n1), .QN(n4458) );
  INVX0 U9315_U2 ( .INP(n5016), .ZN(U9315_n1) );
  NOR2X0 U9315_U1 ( .IN1(n5753), .IN2(U9315_n1), .QN(n5014) );
  INVX0 U9453_U2 ( .INP(n3065), .ZN(U9453_n1) );
  NOR2X0 U9453_U1 ( .IN1(n616), .IN2(U9453_n1), .QN(n3064) );
  INVX0 U9825_U2 ( .INP(g112), .ZN(U9825_n1) );
  NOR2X0 U9825_U1 ( .IN1(n1430), .IN2(U9825_n1), .QN(n3115) );
  INVX0 U9886_U2 ( .INP(g370), .ZN(U9886_n1) );
  NOR2X0 U9886_U1 ( .IN1(n917), .IN2(U9886_n1), .QN(n4948) );
  INVX0 U9927_U2 ( .INP(n3933), .ZN(U9927_n1) );
  NOR2X0 U9927_U1 ( .IN1(g4098), .IN2(U9927_n1), .QN(n3833) );
  INVX0 U9953_U2 ( .INP(g671), .ZN(U9953_n1) );
  NOR2X0 U9953_U1 ( .IN1(n8195), .IN2(U9953_n1), .QN(n4526) );
  INVX0 U9957_U2 ( .INP(g4843), .ZN(U9957_n1) );
  NOR2X0 U9957_U1 ( .IN1(n5283), .IN2(U9957_n1), .QN(n2563) );
  INVX0 U9958_U2 ( .INP(test_so19), .ZN(U9958_n1) );
  NOR2X0 U9958_U1 ( .IN1(n5656), .IN2(U9958_n1), .QN(n2573) );
  INVX0 U9968_U2 ( .INP(n3084), .ZN(U9968_n1) );
  NOR2X0 U9968_U1 ( .IN1(g4358), .IN2(U9968_n1), .QN(n3023) );
  INVX0 U9972_U2 ( .INP(g681), .ZN(U9972_n1) );
  NOR2X0 U9972_U1 ( .IN1(n4535), .IN2(U9972_n1), .QN(n5112) );
  INVX0 U9992_U2 ( .INP(n3675), .ZN(U9992_n1) );
  NOR2X0 U9992_U1 ( .IN1(n3676), .IN2(U9992_n1), .QN(n2644) );
  INVX0 U10314_U2 ( .INP(g667), .ZN(U10314_n1) );
  NOR2X0 U10314_U1 ( .IN1(g686), .IN2(U10314_n1), .QN(n4962) );
  INVX0 U10318_U2 ( .INP(g5092), .ZN(U10318_n1) );
  NOR2X0 U10318_U1 ( .IN1(n5681), .IN2(U10318_n1), .QN(n5016) );
endmodule

