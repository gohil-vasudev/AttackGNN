module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n350_, new_n352_, new_n353_, new_n355_, new_n356_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n377_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n388_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n402_, new_n404_, new_n406_, new_n407_, new_n409_, new_n410_, new_n412_, new_n414_, new_n416_, new_n417_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n441_, new_n442_, new_n444_, new_n445_, new_n447_, new_n448_, new_n450_, new_n451_, new_n453_, new_n454_, new_n455_, new_n457_, new_n459_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n483_, new_n485_, new_n486_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n500_, new_n501_, new_n503_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_;
  XNOR2_X1 g000 ( .A(G155GAT), .B(KEYINPUT3), .ZN(new_n138_) );
  XNOR2_X1 g001 ( .A(G141GAT), .B(KEYINPUT2), .ZN(new_n139_) );
  XNOR2_X1 g002 ( .A(new_n138_), .B(new_n139_), .ZN(new_n140_) );
  XNOR2_X1 g003 ( .A(G57GAT), .B(KEYINPUT1), .ZN(new_n141_) );
  NAND2_X1 g004 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n142_) );
  XNOR2_X1 g005 ( .A(new_n141_), .B(new_n142_), .ZN(new_n143_) );
  XNOR2_X1 g006 ( .A(new_n140_), .B(new_n143_), .ZN(new_n144_) );
  XNOR2_X1 g007 ( .A(G120GAT), .B(G127GAT), .ZN(new_n145_) );
  XNOR2_X1 g008 ( .A(G113GAT), .B(KEYINPUT0), .ZN(new_n146_) );
  XNOR2_X1 g009 ( .A(new_n145_), .B(new_n146_), .ZN(new_n147_) );
  XNOR2_X1 g010 ( .A(new_n147_), .B(G1GAT), .ZN(new_n148_) );
  XNOR2_X1 g011 ( .A(new_n144_), .B(new_n148_), .ZN(new_n149_) );
  XNOR2_X1 g012 ( .A(G29GAT), .B(G134GAT), .ZN(new_n150_) );
  XNOR2_X1 g013 ( .A(new_n149_), .B(new_n150_), .ZN(new_n151_) );
  XOR2_X1 g014 ( .A(G85GAT), .B(G162GAT), .Z(new_n152_) );
  XNOR2_X1 g015 ( .A(new_n151_), .B(new_n152_), .ZN(new_n153_) );
  XOR2_X1 g016 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(new_n154_) );
  XNOR2_X1 g017 ( .A(G148GAT), .B(KEYINPUT6), .ZN(new_n155_) );
  XNOR2_X1 g018 ( .A(new_n154_), .B(new_n155_), .ZN(new_n156_) );
  XNOR2_X1 g019 ( .A(new_n153_), .B(new_n156_), .ZN(new_n157_) );
  INV_X1 g020 ( .A(new_n157_), .ZN(new_n158_) );
  INV_X1 g021 ( .A(KEYINPUT26), .ZN(new_n159_) );
  XOR2_X1 g022 ( .A(G211GAT), .B(G218GAT), .Z(new_n160_) );
  XNOR2_X1 g023 ( .A(G204GAT), .B(KEYINPUT21), .ZN(new_n161_) );
  XNOR2_X1 g024 ( .A(new_n160_), .B(new_n161_), .ZN(new_n162_) );
  XNOR2_X1 g025 ( .A(new_n162_), .B(G197GAT), .ZN(new_n163_) );
  XNOR2_X1 g026 ( .A(new_n163_), .B(new_n140_), .ZN(new_n164_) );
  XNOR2_X1 g027 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(new_n165_) );
  XNOR2_X1 g028 ( .A(G22GAT), .B(KEYINPUT22), .ZN(new_n166_) );
  XOR2_X1 g029 ( .A(new_n165_), .B(new_n166_), .Z(new_n167_) );
  INV_X1 g030 ( .A(G78GAT), .ZN(new_n168_) );
  NAND2_X1 g031 ( .A1(new_n168_), .A2(G106GAT), .ZN(new_n169_) );
  INV_X1 g032 ( .A(G106GAT), .ZN(new_n170_) );
  NAND2_X1 g033 ( .A1(new_n170_), .A2(G78GAT), .ZN(new_n171_) );
  NAND3_X1 g034 ( .A1(new_n169_), .A2(new_n171_), .A3(G148GAT), .ZN(new_n172_) );
  INV_X1 g035 ( .A(G148GAT), .ZN(new_n173_) );
  NAND2_X1 g036 ( .A1(new_n169_), .A2(new_n171_), .ZN(new_n174_) );
  NAND2_X1 g037 ( .A1(new_n174_), .A2(new_n173_), .ZN(new_n175_) );
  NAND2_X1 g038 ( .A1(new_n175_), .A2(new_n172_), .ZN(new_n176_) );
  XNOR2_X1 g039 ( .A(new_n167_), .B(new_n176_), .ZN(new_n177_) );
  NAND2_X1 g040 ( .A1(new_n164_), .A2(new_n177_), .ZN(new_n178_) );
  OR2_X1 g041 ( .A1(new_n164_), .A2(new_n177_), .ZN(new_n179_) );
  NAND2_X1 g042 ( .A1(new_n179_), .A2(new_n178_), .ZN(new_n180_) );
  XNOR2_X1 g043 ( .A(G50GAT), .B(G162GAT), .ZN(new_n181_) );
  NAND2_X1 g044 ( .A1(new_n180_), .A2(new_n181_), .ZN(new_n182_) );
  INV_X1 g045 ( .A(new_n181_), .ZN(new_n183_) );
  NAND3_X1 g046 ( .A1(new_n179_), .A2(new_n178_), .A3(new_n183_), .ZN(new_n184_) );
  NAND2_X1 g047 ( .A1(new_n182_), .A2(new_n184_), .ZN(new_n185_) );
  NAND2_X1 g048 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n186_) );
  INV_X1 g049 ( .A(new_n186_), .ZN(new_n187_) );
  NAND2_X1 g050 ( .A1(new_n185_), .A2(new_n187_), .ZN(new_n188_) );
  NAND3_X1 g051 ( .A1(new_n182_), .A2(new_n184_), .A3(new_n186_), .ZN(new_n189_) );
  XNOR2_X1 g052 ( .A(new_n147_), .B(G15GAT), .ZN(new_n190_) );
  NAND2_X1 g053 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n191_) );
  XNOR2_X1 g054 ( .A(new_n190_), .B(new_n191_), .ZN(new_n192_) );
  XOR2_X1 g055 ( .A(G176GAT), .B(G183GAT), .Z(new_n193_) );
  XNOR2_X1 g056 ( .A(G71GAT), .B(KEYINPUT20), .ZN(new_n194_) );
  XNOR2_X1 g057 ( .A(new_n193_), .B(new_n194_), .ZN(new_n195_) );
  XNOR2_X1 g058 ( .A(new_n192_), .B(new_n195_), .ZN(new_n196_) );
  XOR2_X1 g059 ( .A(G134GAT), .B(G190GAT), .Z(new_n197_) );
  XNOR2_X1 g060 ( .A(G43GAT), .B(G99GAT), .ZN(new_n198_) );
  XNOR2_X1 g061 ( .A(new_n197_), .B(new_n198_), .ZN(new_n199_) );
  XNOR2_X1 g062 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(new_n200_) );
  XNOR2_X1 g063 ( .A(G169GAT), .B(KEYINPUT19), .ZN(new_n201_) );
  XNOR2_X1 g064 ( .A(new_n200_), .B(new_n201_), .ZN(new_n202_) );
  XNOR2_X1 g065 ( .A(new_n199_), .B(new_n202_), .ZN(new_n203_) );
  XNOR2_X1 g066 ( .A(new_n196_), .B(new_n203_), .ZN(new_n204_) );
  NAND3_X1 g067 ( .A1(new_n188_), .A2(new_n189_), .A3(new_n204_), .ZN(new_n205_) );
  NAND2_X1 g068 ( .A1(new_n205_), .A2(new_n159_), .ZN(new_n206_) );
  NAND4_X1 g069 ( .A1(new_n188_), .A2(KEYINPUT26), .A3(new_n189_), .A4(new_n204_), .ZN(new_n207_) );
  NAND2_X1 g070 ( .A1(new_n206_), .A2(new_n207_), .ZN(new_n208_) );
  XOR2_X1 g071 ( .A(G36GAT), .B(G190GAT), .Z(new_n209_) );
  XNOR2_X1 g072 ( .A(new_n163_), .B(new_n209_), .ZN(new_n210_) );
  INV_X1 g073 ( .A(G92GAT), .ZN(new_n211_) );
  XNOR2_X1 g074 ( .A(G64GAT), .B(G176GAT), .ZN(new_n212_) );
  XNOR2_X1 g075 ( .A(new_n212_), .B(new_n211_), .ZN(new_n213_) );
  NAND2_X1 g076 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n214_) );
  XNOR2_X1 g077 ( .A(new_n213_), .B(new_n214_), .ZN(new_n215_) );
  XOR2_X1 g078 ( .A(G8GAT), .B(G183GAT), .Z(new_n216_) );
  XNOR2_X1 g079 ( .A(new_n215_), .B(new_n216_), .ZN(new_n217_) );
  XNOR2_X1 g080 ( .A(new_n210_), .B(new_n217_), .ZN(new_n218_) );
  XNOR2_X1 g081 ( .A(new_n218_), .B(new_n202_), .ZN(new_n219_) );
  XNOR2_X1 g082 ( .A(new_n219_), .B(KEYINPUT27), .ZN(new_n220_) );
  NAND2_X1 g083 ( .A1(new_n208_), .A2(new_n220_), .ZN(new_n221_) );
  INV_X1 g084 ( .A(KEYINPUT25), .ZN(new_n222_) );
  NAND2_X1 g085 ( .A1(new_n188_), .A2(new_n189_), .ZN(new_n223_) );
  INV_X1 g086 ( .A(new_n204_), .ZN(new_n224_) );
  NAND2_X1 g087 ( .A1(new_n224_), .A2(new_n219_), .ZN(new_n225_) );
  NAND2_X1 g088 ( .A1(new_n223_), .A2(new_n225_), .ZN(new_n226_) );
  NAND2_X1 g089 ( .A1(new_n226_), .A2(new_n222_), .ZN(new_n227_) );
  NAND3_X1 g090 ( .A1(new_n223_), .A2(new_n225_), .A3(KEYINPUT25), .ZN(new_n228_) );
  NAND2_X1 g091 ( .A1(new_n227_), .A2(new_n228_), .ZN(new_n229_) );
  NAND2_X1 g092 ( .A1(new_n221_), .A2(new_n229_), .ZN(new_n230_) );
  NAND2_X1 g093 ( .A1(new_n230_), .A2(new_n158_), .ZN(new_n231_) );
  XNOR2_X1 g094 ( .A(new_n223_), .B(KEYINPUT28), .ZN(new_n232_) );
  AND2_X1 g095 ( .A1(new_n220_), .A2(new_n157_), .ZN(new_n233_) );
  NAND3_X1 g096 ( .A1(new_n232_), .A2(new_n233_), .A3(new_n204_), .ZN(new_n234_) );
  NAND2_X1 g097 ( .A1(new_n231_), .A2(new_n234_), .ZN(new_n235_) );
  INV_X1 g098 ( .A(new_n209_), .ZN(new_n236_) );
  XNOR2_X1 g099 ( .A(G106GAT), .B(G218GAT), .ZN(new_n237_) );
  XNOR2_X1 g100 ( .A(new_n150_), .B(new_n237_), .ZN(new_n238_) );
  XOR2_X1 g101 ( .A(new_n238_), .B(KEYINPUT9), .Z(new_n239_) );
  XNOR2_X1 g102 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(new_n240_) );
  NAND2_X1 g103 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n241_) );
  XNOR2_X1 g104 ( .A(new_n240_), .B(new_n241_), .ZN(new_n242_) );
  XNOR2_X1 g105 ( .A(G85GAT), .B(G99GAT), .ZN(new_n243_) );
  NAND2_X1 g106 ( .A1(new_n243_), .A2(G92GAT), .ZN(new_n244_) );
  NAND2_X1 g107 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n245_) );
  OR2_X1 g108 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n246_) );
  NAND3_X1 g109 ( .A1(new_n246_), .A2(new_n211_), .A3(new_n245_), .ZN(new_n247_) );
  NAND2_X1 g110 ( .A1(new_n244_), .A2(new_n247_), .ZN(new_n248_) );
  XNOR2_X1 g111 ( .A(G43GAT), .B(KEYINPUT8), .ZN(new_n249_) );
  NAND2_X1 g112 ( .A1(new_n249_), .A2(KEYINPUT7), .ZN(new_n250_) );
  INV_X1 g113 ( .A(KEYINPUT7), .ZN(new_n251_) );
  NAND2_X1 g114 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n252_) );
  OR2_X1 g115 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n253_) );
  NAND3_X1 g116 ( .A1(new_n253_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n254_) );
  NAND2_X1 g117 ( .A1(new_n250_), .A2(new_n254_), .ZN(new_n255_) );
  XNOR2_X1 g118 ( .A(new_n248_), .B(new_n255_), .ZN(new_n256_) );
  XNOR2_X1 g119 ( .A(new_n256_), .B(new_n242_), .ZN(new_n257_) );
  NAND2_X1 g120 ( .A1(new_n257_), .A2(new_n239_), .ZN(new_n258_) );
  INV_X1 g121 ( .A(new_n239_), .ZN(new_n259_) );
  OR2_X1 g122 ( .A1(new_n256_), .A2(new_n242_), .ZN(new_n260_) );
  NAND2_X1 g123 ( .A1(new_n256_), .A2(new_n242_), .ZN(new_n261_) );
  NAND3_X1 g124 ( .A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_) );
  NAND2_X1 g125 ( .A1(new_n258_), .A2(new_n262_), .ZN(new_n263_) );
  NAND2_X1 g126 ( .A1(new_n263_), .A2(new_n183_), .ZN(new_n264_) );
  NAND3_X1 g127 ( .A1(new_n258_), .A2(new_n181_), .A3(new_n262_), .ZN(new_n265_) );
  NAND2_X1 g128 ( .A1(new_n264_), .A2(new_n265_), .ZN(new_n266_) );
  NAND2_X1 g129 ( .A1(new_n266_), .A2(new_n236_), .ZN(new_n267_) );
  NAND3_X1 g130 ( .A1(new_n264_), .A2(new_n209_), .A3(new_n265_), .ZN(new_n268_) );
  XOR2_X1 g131 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(new_n269_) );
  XNOR2_X1 g132 ( .A(G64GAT), .B(KEYINPUT15), .ZN(new_n270_) );
  XNOR2_X1 g133 ( .A(new_n269_), .B(new_n270_), .ZN(new_n271_) );
  XNOR2_X1 g134 ( .A(G78GAT), .B(G155GAT), .ZN(new_n272_) );
  XNOR2_X1 g135 ( .A(G127GAT), .B(G211GAT), .ZN(new_n273_) );
  XNOR2_X1 g136 ( .A(new_n272_), .B(new_n273_), .ZN(new_n274_) );
  XNOR2_X1 g137 ( .A(new_n271_), .B(new_n274_), .ZN(new_n275_) );
  XNOR2_X1 g138 ( .A(G57GAT), .B(G71GAT), .ZN(new_n276_) );
  XOR2_X1 g139 ( .A(new_n276_), .B(KEYINPUT13), .Z(new_n277_) );
  INV_X1 g140 ( .A(G1GAT), .ZN(new_n278_) );
  XNOR2_X1 g141 ( .A(G15GAT), .B(G22GAT), .ZN(new_n279_) );
  XNOR2_X1 g142 ( .A(new_n279_), .B(new_n278_), .ZN(new_n280_) );
  XNOR2_X1 g143 ( .A(new_n277_), .B(new_n280_), .ZN(new_n281_) );
  XNOR2_X1 g144 ( .A(new_n281_), .B(new_n275_), .ZN(new_n282_) );
  XNOR2_X1 g145 ( .A(new_n282_), .B(new_n216_), .ZN(new_n283_) );
  NAND2_X1 g146 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n284_) );
  XOR2_X1 g147 ( .A(new_n283_), .B(new_n284_), .Z(new_n285_) );
  NAND3_X1 g148 ( .A1(new_n285_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n286_) );
  XOR2_X1 g149 ( .A(new_n286_), .B(KEYINPUT16), .Z(new_n287_) );
  AND2_X1 g150 ( .A1(new_n235_), .A2(new_n287_), .ZN(new_n288_) );
  XOR2_X1 g151 ( .A(new_n280_), .B(new_n255_), .Z(new_n289_) );
  XNOR2_X1 g152 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(new_n290_) );
  XNOR2_X1 g153 ( .A(G8GAT), .B(G169GAT), .ZN(new_n291_) );
  XNOR2_X1 g154 ( .A(new_n290_), .B(new_n291_), .ZN(new_n292_) );
  XNOR2_X1 g155 ( .A(G113GAT), .B(G197GAT), .ZN(new_n293_) );
  XNOR2_X1 g156 ( .A(G29GAT), .B(G141GAT), .ZN(new_n294_) );
  XNOR2_X1 g157 ( .A(new_n293_), .B(new_n294_), .ZN(new_n295_) );
  XNOR2_X1 g158 ( .A(new_n292_), .B(new_n295_), .ZN(new_n296_) );
  XNOR2_X1 g159 ( .A(new_n289_), .B(new_n296_), .ZN(new_n297_) );
  XOR2_X1 g160 ( .A(G36GAT), .B(G50GAT), .Z(new_n298_) );
  NAND2_X1 g161 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n299_) );
  XNOR2_X1 g162 ( .A(new_n298_), .B(new_n299_), .ZN(new_n300_) );
  XNOR2_X1 g163 ( .A(new_n297_), .B(new_n300_), .ZN(new_n301_) );
  INV_X1 g164 ( .A(new_n301_), .ZN(new_n302_) );
  XOR2_X1 g165 ( .A(G120GAT), .B(G204GAT), .Z(new_n303_) );
  INV_X1 g166 ( .A(new_n303_), .ZN(new_n304_) );
  NAND2_X1 g167 ( .A1(new_n176_), .A2(new_n248_), .ZN(new_n305_) );
  NAND4_X1 g168 ( .A1(new_n175_), .A2(new_n244_), .A3(new_n172_), .A4(new_n247_), .ZN(new_n306_) );
  NAND2_X1 g169 ( .A1(new_n305_), .A2(new_n306_), .ZN(new_n307_) );
  INV_X1 g170 ( .A(KEYINPUT32), .ZN(new_n308_) );
  NAND2_X1 g171 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n309_) );
  INV_X1 g172 ( .A(KEYINPUT31), .ZN(new_n310_) );
  NAND2_X1 g173 ( .A1(new_n310_), .A2(KEYINPUT33), .ZN(new_n311_) );
  INV_X1 g174 ( .A(KEYINPUT33), .ZN(new_n312_) );
  NAND2_X1 g175 ( .A1(new_n312_), .A2(KEYINPUT31), .ZN(new_n313_) );
  NAND2_X1 g176 ( .A1(new_n311_), .A2(new_n313_), .ZN(new_n314_) );
  NAND2_X1 g177 ( .A1(new_n314_), .A2(new_n309_), .ZN(new_n315_) );
  NAND4_X1 g178 ( .A1(new_n311_), .A2(new_n313_), .A3(G230GAT), .A4(G233GAT), .ZN(new_n316_) );
  NAND3_X1 g179 ( .A1(new_n315_), .A2(new_n308_), .A3(new_n316_), .ZN(new_n317_) );
  NAND2_X1 g180 ( .A1(new_n315_), .A2(new_n316_), .ZN(new_n318_) );
  NAND2_X1 g181 ( .A1(new_n318_), .A2(KEYINPUT32), .ZN(new_n319_) );
  NAND2_X1 g182 ( .A1(new_n319_), .A2(new_n317_), .ZN(new_n320_) );
  NAND2_X1 g183 ( .A1(new_n307_), .A2(new_n320_), .ZN(new_n321_) );
  NAND4_X1 g184 ( .A1(new_n311_), .A2(new_n313_), .A3(G230GAT), .A4(G233GAT), .ZN(new_n322_) );
  NAND3_X1 g185 ( .A1(new_n315_), .A2(new_n308_), .A3(new_n322_), .ZN(new_n323_) );
  NAND4_X1 g186 ( .A1(new_n305_), .A2(new_n319_), .A3(new_n306_), .A4(new_n323_), .ZN(new_n324_) );
  NAND2_X1 g187 ( .A1(new_n321_), .A2(new_n324_), .ZN(new_n325_) );
  NAND2_X1 g188 ( .A1(new_n325_), .A2(new_n212_), .ZN(new_n326_) );
  INV_X1 g189 ( .A(new_n212_), .ZN(new_n327_) );
  NAND3_X1 g190 ( .A1(new_n321_), .A2(new_n327_), .A3(new_n324_), .ZN(new_n328_) );
  NAND2_X1 g191 ( .A1(new_n326_), .A2(new_n328_), .ZN(new_n329_) );
  NAND2_X1 g192 ( .A1(new_n329_), .A2(new_n304_), .ZN(new_n330_) );
  NAND4_X1 g193 ( .A1(new_n305_), .A2(new_n319_), .A3(new_n306_), .A4(new_n317_), .ZN(new_n331_) );
  NAND2_X1 g194 ( .A1(new_n319_), .A2(new_n323_), .ZN(new_n332_) );
  NAND2_X1 g195 ( .A1(new_n307_), .A2(new_n332_), .ZN(new_n333_) );
  NAND2_X1 g196 ( .A1(new_n333_), .A2(new_n331_), .ZN(new_n334_) );
  NAND2_X1 g197 ( .A1(new_n334_), .A2(new_n212_), .ZN(new_n335_) );
  NAND3_X1 g198 ( .A1(new_n335_), .A2(new_n303_), .A3(new_n328_), .ZN(new_n336_) );
  NAND3_X1 g199 ( .A1(new_n330_), .A2(new_n277_), .A3(new_n336_), .ZN(new_n337_) );
  INV_X1 g200 ( .A(new_n277_), .ZN(new_n338_) );
  NAND2_X1 g201 ( .A1(new_n335_), .A2(new_n328_), .ZN(new_n339_) );
  NAND2_X1 g202 ( .A1(new_n339_), .A2(new_n304_), .ZN(new_n340_) );
  NAND2_X1 g203 ( .A1(new_n340_), .A2(new_n336_), .ZN(new_n341_) );
  NAND2_X1 g204 ( .A1(new_n341_), .A2(new_n338_), .ZN(new_n342_) );
  NAND2_X1 g205 ( .A1(new_n342_), .A2(new_n337_), .ZN(new_n343_) );
  INV_X1 g206 ( .A(new_n343_), .ZN(new_n344_) );
  NOR2_X1 g207 ( .A1(new_n344_), .A2(new_n302_), .ZN(new_n345_) );
  AND2_X1 g208 ( .A1(new_n288_), .A2(new_n345_), .ZN(new_n346_) );
  NAND2_X1 g209 ( .A1(new_n346_), .A2(new_n157_), .ZN(new_n347_) );
  XNOR2_X1 g210 ( .A(new_n347_), .B(KEYINPUT34), .ZN(new_n348_) );
  XNOR2_X1 g211 ( .A(new_n348_), .B(G1GAT), .ZN(G1324GAT) );
  NAND2_X1 g212 ( .A1(new_n346_), .A2(new_n219_), .ZN(new_n350_) );
  XNOR2_X1 g213 ( .A(new_n350_), .B(G8GAT), .ZN(G1325GAT) );
  NAND2_X1 g214 ( .A1(new_n346_), .A2(new_n224_), .ZN(new_n352_) );
  XOR2_X1 g215 ( .A(G15GAT), .B(KEYINPUT35), .Z(new_n353_) );
  XNOR2_X1 g216 ( .A(new_n352_), .B(new_n353_), .ZN(G1326GAT) );
  INV_X1 g217 ( .A(new_n232_), .ZN(new_n355_) );
  NAND2_X1 g218 ( .A1(new_n346_), .A2(new_n355_), .ZN(new_n356_) );
  XNOR2_X1 g219 ( .A(new_n356_), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 g220 ( .A(KEYINPUT38), .ZN(new_n358_) );
  INV_X1 g221 ( .A(KEYINPUT36), .ZN(new_n359_) );
  NAND2_X1 g222 ( .A1(new_n267_), .A2(new_n268_), .ZN(new_n360_) );
  NAND2_X1 g223 ( .A1(new_n360_), .A2(new_n359_), .ZN(new_n361_) );
  NAND3_X1 g224 ( .A1(new_n267_), .A2(KEYINPUT36), .A3(new_n268_), .ZN(new_n362_) );
  NAND2_X1 g225 ( .A1(new_n361_), .A2(new_n362_), .ZN(new_n363_) );
  NOR2_X1 g226 ( .A1(new_n363_), .A2(new_n285_), .ZN(new_n364_) );
  NAND2_X1 g227 ( .A1(new_n235_), .A2(new_n364_), .ZN(new_n365_) );
  NAND2_X1 g228 ( .A1(new_n365_), .A2(KEYINPUT37), .ZN(new_n366_) );
  INV_X1 g229 ( .A(KEYINPUT37), .ZN(new_n367_) );
  NAND3_X1 g230 ( .A1(new_n235_), .A2(new_n367_), .A3(new_n364_), .ZN(new_n368_) );
  NAND2_X1 g231 ( .A1(new_n366_), .A2(new_n368_), .ZN(new_n369_) );
  NAND2_X1 g232 ( .A1(new_n369_), .A2(new_n345_), .ZN(new_n370_) );
  NAND2_X1 g233 ( .A1(new_n370_), .A2(new_n358_), .ZN(new_n371_) );
  NAND3_X1 g234 ( .A1(new_n369_), .A2(KEYINPUT38), .A3(new_n345_), .ZN(new_n372_) );
  NAND2_X1 g235 ( .A1(new_n371_), .A2(new_n372_), .ZN(new_n373_) );
  NAND2_X1 g236 ( .A1(new_n373_), .A2(new_n157_), .ZN(new_n374_) );
  XOR2_X1 g237 ( .A(G29GAT), .B(KEYINPUT39), .Z(new_n375_) );
  XNOR2_X1 g238 ( .A(new_n374_), .B(new_n375_), .ZN(G1328GAT) );
  NAND2_X1 g239 ( .A1(new_n373_), .A2(new_n219_), .ZN(new_n377_) );
  XNOR2_X1 g240 ( .A(new_n377_), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 g241 ( .A1(new_n373_), .A2(new_n224_), .ZN(new_n379_) );
  NAND2_X1 g242 ( .A1(new_n379_), .A2(KEYINPUT40), .ZN(new_n380_) );
  INV_X1 g243 ( .A(KEYINPUT40), .ZN(new_n381_) );
  NAND3_X1 g244 ( .A1(new_n373_), .A2(new_n381_), .A3(new_n224_), .ZN(new_n382_) );
  NAND2_X1 g245 ( .A1(new_n380_), .A2(new_n382_), .ZN(new_n383_) );
  NAND2_X1 g246 ( .A1(new_n383_), .A2(G43GAT), .ZN(new_n384_) );
  INV_X1 g247 ( .A(G43GAT), .ZN(new_n385_) );
  NAND3_X1 g248 ( .A1(new_n380_), .A2(new_n385_), .A3(new_n382_), .ZN(new_n386_) );
  NAND2_X1 g249 ( .A1(new_n384_), .A2(new_n386_), .ZN(G1330GAT) );
  NAND2_X1 g250 ( .A1(new_n373_), .A2(new_n355_), .ZN(new_n388_) );
  XNOR2_X1 g251 ( .A(new_n388_), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 g252 ( .A1(new_n330_), .A2(new_n336_), .ZN(new_n390_) );
  NAND2_X1 g253 ( .A1(new_n390_), .A2(new_n338_), .ZN(new_n391_) );
  NAND2_X1 g254 ( .A1(new_n391_), .A2(new_n337_), .ZN(new_n392_) );
  NAND2_X1 g255 ( .A1(new_n392_), .A2(KEYINPUT41), .ZN(new_n393_) );
  INV_X1 g256 ( .A(KEYINPUT41), .ZN(new_n394_) );
  NAND3_X1 g257 ( .A1(new_n342_), .A2(new_n394_), .A3(new_n337_), .ZN(new_n395_) );
  NAND2_X1 g258 ( .A1(new_n393_), .A2(new_n395_), .ZN(new_n396_) );
  AND2_X1 g259 ( .A1(new_n396_), .A2(new_n302_), .ZN(new_n397_) );
  AND2_X1 g260 ( .A1(new_n288_), .A2(new_n397_), .ZN(new_n398_) );
  NAND2_X1 g261 ( .A1(new_n398_), .A2(new_n157_), .ZN(new_n399_) );
  XNOR2_X1 g262 ( .A(G57GAT), .B(KEYINPUT42), .ZN(new_n400_) );
  XNOR2_X1 g263 ( .A(new_n399_), .B(new_n400_), .ZN(G1332GAT) );
  NAND2_X1 g264 ( .A1(new_n398_), .A2(new_n219_), .ZN(new_n402_) );
  XNOR2_X1 g265 ( .A(new_n402_), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 g266 ( .A1(new_n398_), .A2(new_n224_), .ZN(new_n404_) );
  XNOR2_X1 g267 ( .A(new_n404_), .B(G71GAT), .ZN(G1334GAT) );
  NAND2_X1 g268 ( .A1(new_n398_), .A2(new_n355_), .ZN(new_n406_) );
  XOR2_X1 g269 ( .A(G78GAT), .B(KEYINPUT43), .Z(new_n407_) );
  XNOR2_X1 g270 ( .A(new_n406_), .B(new_n407_), .ZN(G1335GAT) );
  AND2_X1 g271 ( .A1(new_n369_), .A2(new_n397_), .ZN(new_n409_) );
  NAND2_X1 g272 ( .A1(new_n409_), .A2(new_n157_), .ZN(new_n410_) );
  XNOR2_X1 g273 ( .A(new_n410_), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 g274 ( .A1(new_n409_), .A2(new_n219_), .ZN(new_n412_) );
  XNOR2_X1 g275 ( .A(new_n412_), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 g276 ( .A1(new_n409_), .A2(new_n224_), .ZN(new_n414_) );
  XNOR2_X1 g277 ( .A(new_n414_), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 g278 ( .A1(new_n409_), .A2(new_n355_), .ZN(new_n416_) );
  XNOR2_X1 g279 ( .A(new_n416_), .B(KEYINPUT44), .ZN(new_n417_) );
  XNOR2_X1 g280 ( .A(new_n417_), .B(G106GAT), .ZN(G1339GAT) );
  INV_X1 g281 ( .A(KEYINPUT47), .ZN(new_n419_) );
  NAND3_X1 g282 ( .A1(new_n396_), .A2(KEYINPUT46), .A3(new_n301_), .ZN(new_n420_) );
  INV_X1 g283 ( .A(KEYINPUT46), .ZN(new_n421_) );
  NAND2_X1 g284 ( .A1(new_n396_), .A2(new_n301_), .ZN(new_n422_) );
  NAND2_X1 g285 ( .A1(new_n422_), .A2(new_n421_), .ZN(new_n423_) );
  NOR2_X1 g286 ( .A1(new_n285_), .A2(new_n360_), .ZN(new_n424_) );
  NAND4_X1 g287 ( .A1(new_n423_), .A2(new_n419_), .A3(new_n420_), .A4(new_n424_), .ZN(new_n425_) );
  NAND3_X1 g288 ( .A1(new_n423_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n426_) );
  NAND2_X1 g289 ( .A1(new_n426_), .A2(KEYINPUT47), .ZN(new_n427_) );
  NAND3_X1 g290 ( .A1(new_n361_), .A2(new_n285_), .A3(new_n362_), .ZN(new_n428_) );
  NAND2_X1 g291 ( .A1(new_n428_), .A2(KEYINPUT45), .ZN(new_n429_) );
  INV_X1 g292 ( .A(KEYINPUT45), .ZN(new_n430_) );
  NAND4_X1 g293 ( .A1(new_n361_), .A2(new_n285_), .A3(new_n430_), .A4(new_n362_), .ZN(new_n431_) );
  NAND4_X1 g294 ( .A1(new_n429_), .A2(new_n302_), .A3(new_n343_), .A4(new_n431_), .ZN(new_n432_) );
  NAND4_X1 g295 ( .A1(new_n427_), .A2(new_n432_), .A3(KEYINPUT48), .A4(new_n425_), .ZN(new_n433_) );
  INV_X1 g296 ( .A(KEYINPUT48), .ZN(new_n434_) );
  NAND3_X1 g297 ( .A1(new_n427_), .A2(new_n425_), .A3(new_n432_), .ZN(new_n435_) );
  NAND2_X1 g298 ( .A1(new_n435_), .A2(new_n434_), .ZN(new_n436_) );
  AND3_X1 g299 ( .A1(new_n436_), .A2(new_n233_), .A3(new_n433_), .ZN(new_n437_) );
  AND3_X1 g300 ( .A1(new_n437_), .A2(new_n224_), .A3(new_n232_), .ZN(new_n438_) );
  NAND2_X1 g301 ( .A1(new_n438_), .A2(new_n301_), .ZN(new_n439_) );
  XNOR2_X1 g302 ( .A(new_n439_), .B(G113GAT), .ZN(G1340GAT) );
  NAND2_X1 g303 ( .A1(new_n438_), .A2(new_n396_), .ZN(new_n441_) );
  XOR2_X1 g304 ( .A(G120GAT), .B(KEYINPUT49), .Z(new_n442_) );
  XNOR2_X1 g305 ( .A(new_n441_), .B(new_n442_), .ZN(G1341GAT) );
  NAND2_X1 g306 ( .A1(new_n438_), .A2(new_n285_), .ZN(new_n444_) );
  XNOR2_X1 g307 ( .A(new_n444_), .B(KEYINPUT50), .ZN(new_n445_) );
  XNOR2_X1 g308 ( .A(new_n445_), .B(G127GAT), .ZN(G1342GAT) );
  NAND2_X1 g309 ( .A1(new_n438_), .A2(new_n360_), .ZN(new_n447_) );
  XOR2_X1 g310 ( .A(G134GAT), .B(KEYINPUT51), .Z(new_n448_) );
  XNOR2_X1 g311 ( .A(new_n447_), .B(new_n448_), .ZN(G1343GAT) );
  AND2_X1 g312 ( .A1(new_n437_), .A2(new_n208_), .ZN(new_n450_) );
  NAND2_X1 g313 ( .A1(new_n450_), .A2(new_n301_), .ZN(new_n451_) );
  XNOR2_X1 g314 ( .A(new_n451_), .B(G141GAT), .ZN(G1344GAT) );
  NAND2_X1 g315 ( .A1(new_n450_), .A2(new_n396_), .ZN(new_n453_) );
  XOR2_X1 g316 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(new_n454_) );
  XNOR2_X1 g317 ( .A(new_n453_), .B(new_n454_), .ZN(new_n455_) );
  XNOR2_X1 g318 ( .A(new_n455_), .B(G148GAT), .ZN(G1345GAT) );
  NAND2_X1 g319 ( .A1(new_n450_), .A2(new_n285_), .ZN(new_n457_) );
  XNOR2_X1 g320 ( .A(new_n457_), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 g321 ( .A1(new_n450_), .A2(new_n360_), .ZN(new_n459_) );
  XNOR2_X1 g322 ( .A(new_n459_), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 g323 ( .A(KEYINPUT55), .ZN(new_n461_) );
  INV_X1 g324 ( .A(KEYINPUT54), .ZN(new_n462_) );
  NAND4_X1 g325 ( .A1(new_n436_), .A2(new_n462_), .A3(new_n219_), .A4(new_n433_), .ZN(new_n463_) );
  NAND3_X1 g326 ( .A1(new_n436_), .A2(new_n219_), .A3(new_n433_), .ZN(new_n464_) );
  NAND2_X1 g327 ( .A1(new_n464_), .A2(KEYINPUT54), .ZN(new_n465_) );
  AND2_X1 g328 ( .A1(new_n465_), .A2(new_n158_), .ZN(new_n466_) );
  NAND4_X1 g329 ( .A1(new_n466_), .A2(new_n461_), .A3(new_n223_), .A4(new_n463_), .ZN(new_n467_) );
  NAND4_X1 g330 ( .A1(new_n465_), .A2(new_n158_), .A3(new_n223_), .A4(new_n463_), .ZN(new_n468_) );
  NAND2_X1 g331 ( .A1(new_n468_), .A2(KEYINPUT55), .ZN(new_n469_) );
  NAND2_X1 g332 ( .A1(new_n467_), .A2(new_n469_), .ZN(new_n470_) );
  NAND3_X1 g333 ( .A1(new_n470_), .A2(new_n224_), .A3(new_n301_), .ZN(new_n471_) );
  XNOR2_X1 g334 ( .A(new_n471_), .B(G169GAT), .ZN(G1348GAT) );
  INV_X1 g335 ( .A(G176GAT), .ZN(new_n473_) );
  NAND3_X1 g336 ( .A1(new_n470_), .A2(new_n224_), .A3(new_n396_), .ZN(new_n474_) );
  XOR2_X1 g337 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(new_n475_) );
  INV_X1 g338 ( .A(new_n475_), .ZN(new_n476_) );
  NAND2_X1 g339 ( .A1(new_n474_), .A2(new_n476_), .ZN(new_n477_) );
  NAND4_X1 g340 ( .A1(new_n470_), .A2(new_n224_), .A3(new_n396_), .A4(new_n475_), .ZN(new_n478_) );
  NAND2_X1 g341 ( .A1(new_n477_), .A2(new_n478_), .ZN(new_n479_) );
  NAND2_X1 g342 ( .A1(new_n479_), .A2(new_n473_), .ZN(new_n480_) );
  NAND3_X1 g343 ( .A1(new_n477_), .A2(G176GAT), .A3(new_n478_), .ZN(new_n481_) );
  NAND2_X1 g344 ( .A1(new_n480_), .A2(new_n481_), .ZN(G1349GAT) );
  NAND3_X1 g345 ( .A1(new_n470_), .A2(new_n224_), .A3(new_n285_), .ZN(new_n483_) );
  XNOR2_X1 g346 ( .A(new_n483_), .B(G183GAT), .ZN(G1350GAT) );
  NAND3_X1 g347 ( .A1(new_n470_), .A2(new_n224_), .A3(new_n360_), .ZN(new_n485_) );
  XNOR2_X1 g348 ( .A(G190GAT), .B(KEYINPUT58), .ZN(new_n486_) );
  XNOR2_X1 g349 ( .A(new_n485_), .B(new_n486_), .ZN(G1351GAT) );
  AND2_X1 g350 ( .A1(new_n466_), .A2(new_n463_), .ZN(new_n488_) );
  NAND3_X1 g351 ( .A1(new_n488_), .A2(new_n208_), .A3(new_n301_), .ZN(new_n489_) );
  XNOR2_X1 g352 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(new_n490_) );
  INV_X1 g353 ( .A(new_n490_), .ZN(new_n491_) );
  NAND2_X1 g354 ( .A1(new_n489_), .A2(new_n491_), .ZN(new_n492_) );
  AND2_X1 g355 ( .A1(new_n488_), .A2(new_n208_), .ZN(new_n493_) );
  NAND3_X1 g356 ( .A1(new_n493_), .A2(new_n301_), .A3(new_n490_), .ZN(new_n494_) );
  NAND2_X1 g357 ( .A1(new_n494_), .A2(new_n492_), .ZN(new_n495_) );
  NAND2_X1 g358 ( .A1(new_n495_), .A2(G197GAT), .ZN(new_n496_) );
  INV_X1 g359 ( .A(G197GAT), .ZN(new_n497_) );
  NAND3_X1 g360 ( .A1(new_n494_), .A2(new_n497_), .A3(new_n492_), .ZN(new_n498_) );
  NAND2_X1 g361 ( .A1(new_n496_), .A2(new_n498_), .ZN(G1352GAT) );
  NAND2_X1 g362 ( .A1(new_n493_), .A2(new_n344_), .ZN(new_n500_) );
  XOR2_X1 g363 ( .A(G204GAT), .B(KEYINPUT61), .Z(new_n501_) );
  XNOR2_X1 g364 ( .A(new_n500_), .B(new_n501_), .ZN(G1353GAT) );
  NAND2_X1 g365 ( .A1(new_n493_), .A2(new_n285_), .ZN(new_n503_) );
  XNOR2_X1 g366 ( .A(new_n503_), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 g367 ( .A(new_n363_), .ZN(new_n505_) );
  NAND3_X1 g368 ( .A1(new_n488_), .A2(new_n208_), .A3(new_n505_), .ZN(new_n506_) );
  OR2_X1 g369 ( .A1(new_n506_), .A2(KEYINPUT62), .ZN(new_n507_) );
  NAND2_X1 g370 ( .A1(new_n506_), .A2(KEYINPUT62), .ZN(new_n508_) );
  NAND2_X1 g371 ( .A1(new_n507_), .A2(new_n508_), .ZN(new_n509_) );
  NAND2_X1 g372 ( .A1(new_n509_), .A2(G218GAT), .ZN(new_n510_) );
  INV_X1 g373 ( .A(G218GAT), .ZN(new_n511_) );
  NAND3_X1 g374 ( .A1(new_n507_), .A2(new_n511_), .A3(new_n508_), .ZN(new_n512_) );
  NAND2_X1 g375 ( .A1(new_n510_), .A2(new_n512_), .ZN(G1355GAT) );
endmodule


