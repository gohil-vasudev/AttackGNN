module add_mul_comp_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, Result_0_, Result_1_, Result_2_, 
        Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, 
        Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, 
        Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, 
        Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, 
        Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, Result_32_, 
        Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, Result_38_, 
        Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, Result_44_, 
        Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, Result_50_, 
        Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, Result_56_, 
        Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, Result_62_, 
        Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088;

  INV_X2 U7618 ( .A(n7584), .ZN(n7554) );
  INV_X2 U7619 ( .A(b_9_), .ZN(n8049) );
  INV_X2 U7620 ( .A(b_29_), .ZN(n7611) );
  INV_X2 U7621 ( .A(b_21_), .ZN(n8103) );
  INV_X2 U7622 ( .A(b_17_), .ZN(n8085) );
  INV_X2 U7623 ( .A(b_13_), .ZN(n8067) );
  INV_X2 U7624 ( .A(b_19_), .ZN(n8094) );
  INV_X2 U7625 ( .A(b_15_), .ZN(n8076) );
  INV_X2 U7626 ( .A(b_5_), .ZN(n8031) );
  INV_X2 U7627 ( .A(b_11_), .ZN(n8058) );
  INV_X2 U7628 ( .A(b_7_), .ZN(n8040) );
  INV_X2 U7629 ( .A(b_3_), .ZN(n8022) );
  AND2_X1 U7630 ( .A1(n7554), .A2(n7555), .ZN(Result_9_) );
  XOR2_X1 U7631 ( .A(n7556), .B(n7557), .Z(n7555) );
  AND2_X1 U7632 ( .A1(n7558), .A2(n7559), .ZN(n7557) );
  OR2_X1 U7633 ( .A1(n7560), .A2(n7561), .ZN(n7559) );
  AND2_X1 U7634 ( .A1(n7562), .A2(n7563), .ZN(n7561) );
  INV_X1 U7635 ( .A(n7564), .ZN(n7558) );
  AND2_X1 U7636 ( .A1(n7565), .A2(n7554), .ZN(Result_8_) );
  XOR2_X1 U7637 ( .A(n7566), .B(n7567), .Z(n7565) );
  AND2_X1 U7638 ( .A1(n7554), .A2(n7568), .ZN(Result_7_) );
  XOR2_X1 U7639 ( .A(n7569), .B(n7570), .Z(n7568) );
  AND2_X1 U7640 ( .A1(n7571), .A2(n7572), .ZN(n7570) );
  OR2_X1 U7641 ( .A1(n7573), .A2(n7574), .ZN(n7572) );
  AND2_X1 U7642 ( .A1(n7575), .A2(n7576), .ZN(n7574) );
  INV_X1 U7643 ( .A(n7577), .ZN(n7571) );
  AND2_X1 U7644 ( .A1(n7578), .A2(n7554), .ZN(Result_6_) );
  XOR2_X1 U7645 ( .A(n7579), .B(n7580), .Z(n7578) );
  OR2_X1 U7646 ( .A1(n7581), .A2(n7582), .ZN(Result_63_) );
  AND2_X1 U7647 ( .A1(n7583), .A2(n7584), .ZN(n7582) );
  OR2_X1 U7648 ( .A1(n7585), .A2(n7586), .ZN(n7583) );
  AND2_X1 U7649 ( .A1(b_31_), .A2(n7587), .ZN(n7585) );
  AND2_X1 U7650 ( .A1(n7588), .A2(n7554), .ZN(n7581) );
  OR2_X1 U7651 ( .A1(n7589), .A2(n7590), .ZN(Result_62_) );
  AND2_X1 U7652 ( .A1(n7591), .A2(n7584), .ZN(n7590) );
  XOR2_X1 U7653 ( .A(n7588), .B(n7592), .Z(n7591) );
  XOR2_X1 U7654 ( .A(b_30_), .B(a_30_), .Z(n7592) );
  AND2_X1 U7655 ( .A1(n7554), .A2(n7593), .ZN(n7589) );
  OR2_X1 U7656 ( .A1(n7594), .A2(n7595), .ZN(n7593) );
  AND2_X1 U7657 ( .A1(b_31_), .A2(n7596), .ZN(n7595) );
  OR2_X1 U7658 ( .A1(n7597), .A2(n7598), .ZN(n7596) );
  AND2_X1 U7659 ( .A1(a_30_), .A2(n7599), .ZN(n7597) );
  AND2_X1 U7660 ( .A1(b_30_), .A2(n7600), .ZN(n7594) );
  OR2_X1 U7661 ( .A1(n7586), .A2(n7601), .ZN(n7600) );
  OR2_X1 U7662 ( .A1(n7602), .A2(n7603), .ZN(Result_61_) );
  AND2_X1 U7663 ( .A1(n7604), .A2(n7584), .ZN(n7603) );
  OR2_X1 U7664 ( .A1(n7605), .A2(n7606), .ZN(n7604) );
  AND2_X1 U7665 ( .A1(n7607), .A2(n7608), .ZN(n7606) );
  OR2_X1 U7666 ( .A1(n7609), .A2(n7610), .ZN(n7608) );
  AND2_X1 U7667 ( .A1(a_29_), .A2(n7611), .ZN(n7609) );
  AND2_X1 U7668 ( .A1(n7612), .A2(n7613), .ZN(n7605) );
  OR2_X1 U7669 ( .A1(n7614), .A2(n7615), .ZN(n7612) );
  INV_X1 U7670 ( .A(n7616), .ZN(n7615) );
  AND2_X1 U7671 ( .A1(n7617), .A2(n7554), .ZN(n7602) );
  XOR2_X1 U7672 ( .A(n7618), .B(n7619), .Z(n7617) );
  XOR2_X1 U7673 ( .A(n7620), .B(n7621), .Z(n7619) );
  OR2_X1 U7674 ( .A1(n7622), .A2(n7623), .ZN(Result_60_) );
  AND2_X1 U7675 ( .A1(n7624), .A2(n7554), .ZN(n7623) );
  XNOR2_X1 U7676 ( .A(n7625), .B(n7626), .ZN(n7624) );
  XOR2_X1 U7677 ( .A(n7627), .B(n7628), .Z(n7626) );
  AND2_X1 U7678 ( .A1(n7629), .A2(n7584), .ZN(n7622) );
  XOR2_X1 U7679 ( .A(n7630), .B(n7631), .Z(n7629) );
  OR2_X1 U7680 ( .A1(n7632), .A2(n7633), .ZN(n7631) );
  INV_X1 U7681 ( .A(n7634), .ZN(n7632) );
  AND2_X1 U7682 ( .A1(n7554), .A2(n7635), .ZN(Result_5_) );
  XOR2_X1 U7683 ( .A(n7636), .B(n7637), .Z(n7635) );
  AND2_X1 U7684 ( .A1(n7638), .A2(n7639), .ZN(n7637) );
  OR2_X1 U7685 ( .A1(n7640), .A2(n7641), .ZN(n7639) );
  AND2_X1 U7686 ( .A1(n7642), .A2(n7643), .ZN(n7641) );
  INV_X1 U7687 ( .A(n7644), .ZN(n7638) );
  OR2_X1 U7688 ( .A1(n7645), .A2(n7646), .ZN(Result_59_) );
  AND2_X1 U7689 ( .A1(n7647), .A2(n7584), .ZN(n7646) );
  OR2_X1 U7690 ( .A1(n7648), .A2(n7649), .ZN(n7647) );
  AND2_X1 U7691 ( .A1(n7650), .A2(n7651), .ZN(n7649) );
  XOR2_X1 U7692 ( .A(b_27_), .B(a_27_), .Z(n7650) );
  AND2_X1 U7693 ( .A1(n7652), .A2(n7653), .ZN(n7648) );
  OR2_X1 U7694 ( .A1(n7654), .A2(n7655), .ZN(n7653) );
  INV_X1 U7695 ( .A(n7656), .ZN(n7655) );
  INV_X1 U7696 ( .A(n7651), .ZN(n7652) );
  AND2_X1 U7697 ( .A1(n7657), .A2(n7554), .ZN(n7645) );
  XNOR2_X1 U7698 ( .A(n7658), .B(n7659), .ZN(n7657) );
  XOR2_X1 U7699 ( .A(n7660), .B(n7661), .Z(n7659) );
  OR2_X1 U7700 ( .A1(n7662), .A2(n7663), .ZN(Result_58_) );
  AND2_X1 U7701 ( .A1(n7664), .A2(n7554), .ZN(n7663) );
  XNOR2_X1 U7702 ( .A(n7665), .B(n7666), .ZN(n7664) );
  XOR2_X1 U7703 ( .A(n7667), .B(n7668), .Z(n7666) );
  AND2_X1 U7704 ( .A1(n7669), .A2(n7584), .ZN(n7662) );
  XOR2_X1 U7705 ( .A(n7670), .B(n7671), .Z(n7669) );
  OR2_X1 U7706 ( .A1(n7672), .A2(n7673), .ZN(n7671) );
  INV_X1 U7707 ( .A(n7674), .ZN(n7672) );
  OR2_X1 U7708 ( .A1(n7675), .A2(n7676), .ZN(Result_57_) );
  AND2_X1 U7709 ( .A1(n7677), .A2(n7584), .ZN(n7676) );
  OR2_X1 U7710 ( .A1(n7678), .A2(n7679), .ZN(n7677) );
  AND2_X1 U7711 ( .A1(n7680), .A2(n7681), .ZN(n7679) );
  XOR2_X1 U7712 ( .A(b_25_), .B(a_25_), .Z(n7680) );
  AND2_X1 U7713 ( .A1(n7682), .A2(n7683), .ZN(n7678) );
  OR2_X1 U7714 ( .A1(n7684), .A2(n7685), .ZN(n7683) );
  INV_X1 U7715 ( .A(n7686), .ZN(n7685) );
  INV_X1 U7716 ( .A(n7681), .ZN(n7682) );
  AND2_X1 U7717 ( .A1(n7687), .A2(n7554), .ZN(n7675) );
  XNOR2_X1 U7718 ( .A(n7688), .B(n7689), .ZN(n7687) );
  XOR2_X1 U7719 ( .A(n7690), .B(n7691), .Z(n7689) );
  OR2_X1 U7720 ( .A1(n7692), .A2(n7693), .ZN(Result_56_) );
  AND2_X1 U7721 ( .A1(n7694), .A2(n7554), .ZN(n7693) );
  XNOR2_X1 U7722 ( .A(n7695), .B(n7696), .ZN(n7694) );
  XOR2_X1 U7723 ( .A(n7697), .B(n7698), .Z(n7696) );
  AND2_X1 U7724 ( .A1(n7699), .A2(n7584), .ZN(n7692) );
  XOR2_X1 U7725 ( .A(n7700), .B(n7701), .Z(n7699) );
  OR2_X1 U7726 ( .A1(n7702), .A2(n7703), .ZN(n7701) );
  INV_X1 U7727 ( .A(n7704), .ZN(n7702) );
  OR2_X1 U7728 ( .A1(n7705), .A2(n7706), .ZN(Result_55_) );
  AND2_X1 U7729 ( .A1(n7707), .A2(n7584), .ZN(n7706) );
  OR2_X1 U7730 ( .A1(n7708), .A2(n7709), .ZN(n7707) );
  AND2_X1 U7731 ( .A1(n7710), .A2(n7711), .ZN(n7709) );
  XOR2_X1 U7732 ( .A(b_23_), .B(a_23_), .Z(n7710) );
  AND2_X1 U7733 ( .A1(n7712), .A2(n7713), .ZN(n7708) );
  OR2_X1 U7734 ( .A1(n7714), .A2(n7715), .ZN(n7713) );
  INV_X1 U7735 ( .A(n7716), .ZN(n7715) );
  INV_X1 U7736 ( .A(n7711), .ZN(n7712) );
  AND2_X1 U7737 ( .A1(n7717), .A2(n7554), .ZN(n7705) );
  XNOR2_X1 U7738 ( .A(n7718), .B(n7719), .ZN(n7717) );
  XOR2_X1 U7739 ( .A(n7720), .B(n7721), .Z(n7719) );
  OR2_X1 U7740 ( .A1(n7722), .A2(n7723), .ZN(Result_54_) );
  AND2_X1 U7741 ( .A1(n7724), .A2(n7554), .ZN(n7723) );
  XNOR2_X1 U7742 ( .A(n7725), .B(n7726), .ZN(n7724) );
  XOR2_X1 U7743 ( .A(n7727), .B(n7728), .Z(n7726) );
  AND2_X1 U7744 ( .A1(n7729), .A2(n7584), .ZN(n7722) );
  XOR2_X1 U7745 ( .A(n7730), .B(n7731), .Z(n7729) );
  OR2_X1 U7746 ( .A1(n7732), .A2(n7733), .ZN(n7731) );
  INV_X1 U7747 ( .A(n7734), .ZN(n7732) );
  OR2_X1 U7748 ( .A1(n7735), .A2(n7736), .ZN(Result_53_) );
  AND2_X1 U7749 ( .A1(n7737), .A2(n7554), .ZN(n7736) );
  XNOR2_X1 U7750 ( .A(n7738), .B(n7739), .ZN(n7737) );
  XOR2_X1 U7751 ( .A(n7740), .B(n7741), .Z(n7739) );
  AND2_X1 U7752 ( .A1(n7742), .A2(n7584), .ZN(n7735) );
  XOR2_X1 U7753 ( .A(n7743), .B(n7744), .Z(n7742) );
  AND2_X1 U7754 ( .A1(n7745), .A2(n7746), .ZN(n7744) );
  OR2_X1 U7755 ( .A1(n7747), .A2(n7748), .ZN(Result_52_) );
  AND2_X1 U7756 ( .A1(n7749), .A2(n7554), .ZN(n7748) );
  XNOR2_X1 U7757 ( .A(n7750), .B(n7751), .ZN(n7749) );
  XOR2_X1 U7758 ( .A(n7752), .B(n7753), .Z(n7751) );
  AND2_X1 U7759 ( .A1(n7754), .A2(n7584), .ZN(n7747) );
  XOR2_X1 U7760 ( .A(n7755), .B(n7756), .Z(n7754) );
  OR2_X1 U7761 ( .A1(n7757), .A2(n7758), .ZN(n7756) );
  OR2_X1 U7762 ( .A1(n7759), .A2(n7760), .ZN(Result_51_) );
  AND2_X1 U7763 ( .A1(n7761), .A2(n7554), .ZN(n7760) );
  XNOR2_X1 U7764 ( .A(n7762), .B(n7763), .ZN(n7761) );
  XOR2_X1 U7765 ( .A(n7764), .B(n7765), .Z(n7763) );
  AND2_X1 U7766 ( .A1(n7766), .A2(n7584), .ZN(n7759) );
  XOR2_X1 U7767 ( .A(n7767), .B(n7768), .Z(n7766) );
  AND2_X1 U7768 ( .A1(n7769), .A2(n7770), .ZN(n7768) );
  OR2_X1 U7769 ( .A1(n7771), .A2(n7772), .ZN(Result_50_) );
  AND2_X1 U7770 ( .A1(n7773), .A2(n7554), .ZN(n7772) );
  XNOR2_X1 U7771 ( .A(n7774), .B(n7775), .ZN(n7773) );
  XOR2_X1 U7772 ( .A(n7776), .B(n7777), .Z(n7775) );
  AND2_X1 U7773 ( .A1(n7778), .A2(n7584), .ZN(n7771) );
  XOR2_X1 U7774 ( .A(n7779), .B(n7780), .Z(n7778) );
  OR2_X1 U7775 ( .A1(n7781), .A2(n7782), .ZN(n7780) );
  AND2_X1 U7776 ( .A1(n7783), .A2(n7554), .ZN(Result_4_) );
  XOR2_X1 U7777 ( .A(n7784), .B(n7785), .Z(n7783) );
  OR2_X1 U7778 ( .A1(n7786), .A2(n7787), .ZN(Result_49_) );
  AND2_X1 U7779 ( .A1(n7788), .A2(n7554), .ZN(n7787) );
  XNOR2_X1 U7780 ( .A(n7789), .B(n7790), .ZN(n7788) );
  XOR2_X1 U7781 ( .A(n7791), .B(n7792), .Z(n7790) );
  AND2_X1 U7782 ( .A1(n7793), .A2(n7584), .ZN(n7786) );
  XOR2_X1 U7783 ( .A(n7794), .B(n7795), .Z(n7793) );
  AND2_X1 U7784 ( .A1(n7796), .A2(n7797), .ZN(n7795) );
  OR2_X1 U7785 ( .A1(n7798), .A2(n7799), .ZN(Result_48_) );
  AND2_X1 U7786 ( .A1(n7800), .A2(n7554), .ZN(n7799) );
  XNOR2_X1 U7787 ( .A(n7801), .B(n7802), .ZN(n7800) );
  XOR2_X1 U7788 ( .A(n7803), .B(n7804), .Z(n7802) );
  AND2_X1 U7789 ( .A1(n7805), .A2(n7584), .ZN(n7798) );
  XOR2_X1 U7790 ( .A(n7806), .B(n7807), .Z(n7805) );
  OR2_X1 U7791 ( .A1(n7808), .A2(n7809), .ZN(n7807) );
  OR2_X1 U7792 ( .A1(n7810), .A2(n7811), .ZN(Result_47_) );
  AND2_X1 U7793 ( .A1(n7812), .A2(n7554), .ZN(n7811) );
  XNOR2_X1 U7794 ( .A(n7813), .B(n7814), .ZN(n7812) );
  XOR2_X1 U7795 ( .A(n7815), .B(n7816), .Z(n7814) );
  AND2_X1 U7796 ( .A1(n7817), .A2(n7584), .ZN(n7810) );
  XOR2_X1 U7797 ( .A(n7818), .B(n7819), .Z(n7817) );
  AND2_X1 U7798 ( .A1(n7820), .A2(n7821), .ZN(n7819) );
  OR2_X1 U7799 ( .A1(n7822), .A2(n7823), .ZN(Result_46_) );
  AND2_X1 U7800 ( .A1(n7824), .A2(n7554), .ZN(n7823) );
  XNOR2_X1 U7801 ( .A(n7825), .B(n7826), .ZN(n7824) );
  XOR2_X1 U7802 ( .A(n7827), .B(n7828), .Z(n7826) );
  AND2_X1 U7803 ( .A1(n7829), .A2(n7584), .ZN(n7822) );
  XOR2_X1 U7804 ( .A(n7830), .B(n7831), .Z(n7829) );
  OR2_X1 U7805 ( .A1(n7832), .A2(n7833), .ZN(n7831) );
  OR2_X1 U7806 ( .A1(n7834), .A2(n7835), .ZN(Result_45_) );
  AND2_X1 U7807 ( .A1(n7836), .A2(n7554), .ZN(n7835) );
  XNOR2_X1 U7808 ( .A(n7837), .B(n7838), .ZN(n7836) );
  XOR2_X1 U7809 ( .A(n7839), .B(n7840), .Z(n7838) );
  AND2_X1 U7810 ( .A1(n7841), .A2(n7584), .ZN(n7834) );
  XOR2_X1 U7811 ( .A(n7842), .B(n7843), .Z(n7841) );
  AND2_X1 U7812 ( .A1(n7844), .A2(n7845), .ZN(n7843) );
  OR2_X1 U7813 ( .A1(n7846), .A2(n7847), .ZN(Result_44_) );
  AND2_X1 U7814 ( .A1(n7848), .A2(n7554), .ZN(n7847) );
  XNOR2_X1 U7815 ( .A(n7849), .B(n7850), .ZN(n7848) );
  XOR2_X1 U7816 ( .A(n7851), .B(n7852), .Z(n7850) );
  AND2_X1 U7817 ( .A1(n7853), .A2(n7584), .ZN(n7846) );
  XOR2_X1 U7818 ( .A(n7854), .B(n7855), .Z(n7853) );
  OR2_X1 U7819 ( .A1(n7856), .A2(n7857), .ZN(n7855) );
  OR2_X1 U7820 ( .A1(n7858), .A2(n7859), .ZN(Result_43_) );
  AND2_X1 U7821 ( .A1(n7860), .A2(n7554), .ZN(n7859) );
  XNOR2_X1 U7822 ( .A(n7861), .B(n7862), .ZN(n7860) );
  XOR2_X1 U7823 ( .A(n7863), .B(n7864), .Z(n7862) );
  AND2_X1 U7824 ( .A1(n7865), .A2(n7584), .ZN(n7858) );
  XOR2_X1 U7825 ( .A(n7866), .B(n7867), .Z(n7865) );
  AND2_X1 U7826 ( .A1(n7868), .A2(n7869), .ZN(n7867) );
  OR2_X1 U7827 ( .A1(n7870), .A2(n7871), .ZN(Result_42_) );
  AND2_X1 U7828 ( .A1(n7872), .A2(n7554), .ZN(n7871) );
  XNOR2_X1 U7829 ( .A(n7873), .B(n7874), .ZN(n7872) );
  XOR2_X1 U7830 ( .A(n7875), .B(n7876), .Z(n7874) );
  AND2_X1 U7831 ( .A1(n7877), .A2(n7584), .ZN(n7870) );
  XOR2_X1 U7832 ( .A(n7878), .B(n7879), .Z(n7877) );
  OR2_X1 U7833 ( .A1(n7880), .A2(n7881), .ZN(n7879) );
  OR2_X1 U7834 ( .A1(n7882), .A2(n7883), .ZN(Result_41_) );
  AND2_X1 U7835 ( .A1(n7884), .A2(n7554), .ZN(n7883) );
  XNOR2_X1 U7836 ( .A(n7885), .B(n7886), .ZN(n7884) );
  XOR2_X1 U7837 ( .A(n7887), .B(n7888), .Z(n7886) );
  AND2_X1 U7838 ( .A1(n7889), .A2(n7584), .ZN(n7882) );
  XOR2_X1 U7839 ( .A(n7890), .B(n7891), .Z(n7889) );
  AND2_X1 U7840 ( .A1(n7892), .A2(n7893), .ZN(n7891) );
  OR2_X1 U7841 ( .A1(n7894), .A2(n7895), .ZN(Result_40_) );
  AND2_X1 U7842 ( .A1(n7896), .A2(n7554), .ZN(n7895) );
  XNOR2_X1 U7843 ( .A(n7897), .B(n7898), .ZN(n7896) );
  XOR2_X1 U7844 ( .A(n7899), .B(n7900), .Z(n7898) );
  AND2_X1 U7845 ( .A1(n7901), .A2(n7584), .ZN(n7894) );
  XOR2_X1 U7846 ( .A(n7902), .B(n7903), .Z(n7901) );
  OR2_X1 U7847 ( .A1(n7904), .A2(n7905), .ZN(n7903) );
  AND2_X1 U7848 ( .A1(n7554), .A2(n7906), .ZN(Result_3_) );
  XOR2_X1 U7849 ( .A(n7907), .B(n7908), .Z(n7906) );
  AND2_X1 U7850 ( .A1(n7909), .A2(n7910), .ZN(n7908) );
  OR2_X1 U7851 ( .A1(n7911), .A2(n7912), .ZN(n7910) );
  AND2_X1 U7852 ( .A1(n7913), .A2(n7914), .ZN(n7912) );
  INV_X1 U7853 ( .A(n7915), .ZN(n7909) );
  OR2_X1 U7854 ( .A1(n7916), .A2(n7917), .ZN(Result_39_) );
  AND2_X1 U7855 ( .A1(n7918), .A2(n7554), .ZN(n7917) );
  XNOR2_X1 U7856 ( .A(n7919), .B(n7920), .ZN(n7918) );
  XOR2_X1 U7857 ( .A(n7921), .B(n7922), .Z(n7920) );
  AND2_X1 U7858 ( .A1(n7923), .A2(n7584), .ZN(n7916) );
  XOR2_X1 U7859 ( .A(n7924), .B(n7925), .Z(n7923) );
  AND2_X1 U7860 ( .A1(n7926), .A2(n7927), .ZN(n7925) );
  OR2_X1 U7861 ( .A1(n7928), .A2(n7929), .ZN(Result_38_) );
  AND2_X1 U7862 ( .A1(n7930), .A2(n7554), .ZN(n7929) );
  XNOR2_X1 U7863 ( .A(n7931), .B(n7932), .ZN(n7930) );
  XOR2_X1 U7864 ( .A(n7933), .B(n7934), .Z(n7932) );
  AND2_X1 U7865 ( .A1(n7935), .A2(n7584), .ZN(n7928) );
  XOR2_X1 U7866 ( .A(n7936), .B(n7937), .Z(n7935) );
  OR2_X1 U7867 ( .A1(n7938), .A2(n7939), .ZN(n7937) );
  OR2_X1 U7868 ( .A1(n7940), .A2(n7941), .ZN(Result_37_) );
  AND2_X1 U7869 ( .A1(n7942), .A2(n7554), .ZN(n7941) );
  XNOR2_X1 U7870 ( .A(n7943), .B(n7944), .ZN(n7942) );
  XOR2_X1 U7871 ( .A(n7945), .B(n7946), .Z(n7944) );
  AND2_X1 U7872 ( .A1(n7947), .A2(n7584), .ZN(n7940) );
  XOR2_X1 U7873 ( .A(n7948), .B(n7949), .Z(n7947) );
  AND2_X1 U7874 ( .A1(n7950), .A2(n7951), .ZN(n7949) );
  OR2_X1 U7875 ( .A1(n7952), .A2(n7953), .ZN(Result_36_) );
  AND2_X1 U7876 ( .A1(n7954), .A2(n7554), .ZN(n7953) );
  XNOR2_X1 U7877 ( .A(n7955), .B(n7956), .ZN(n7954) );
  XOR2_X1 U7878 ( .A(n7957), .B(n7958), .Z(n7956) );
  AND2_X1 U7879 ( .A1(n7959), .A2(n7584), .ZN(n7952) );
  XOR2_X1 U7880 ( .A(n7960), .B(n7961), .Z(n7959) );
  OR2_X1 U7881 ( .A1(n7962), .A2(n7963), .ZN(n7961) );
  OR2_X1 U7882 ( .A1(n7964), .A2(n7965), .ZN(Result_35_) );
  AND2_X1 U7883 ( .A1(n7966), .A2(n7554), .ZN(n7965) );
  XNOR2_X1 U7884 ( .A(n7967), .B(n7968), .ZN(n7966) );
  XOR2_X1 U7885 ( .A(n7969), .B(n7970), .Z(n7968) );
  AND2_X1 U7886 ( .A1(n7971), .A2(n7584), .ZN(n7964) );
  XOR2_X1 U7887 ( .A(n7972), .B(n7973), .Z(n7971) );
  AND2_X1 U7888 ( .A1(n7974), .A2(n7975), .ZN(n7973) );
  OR2_X1 U7889 ( .A1(n7976), .A2(n7977), .ZN(Result_34_) );
  AND2_X1 U7890 ( .A1(n7978), .A2(n7554), .ZN(n7977) );
  XNOR2_X1 U7891 ( .A(n7979), .B(n7980), .ZN(n7978) );
  XOR2_X1 U7892 ( .A(n7981), .B(n7982), .Z(n7980) );
  AND2_X1 U7893 ( .A1(n7983), .A2(n7584), .ZN(n7976) );
  XOR2_X1 U7894 ( .A(n7984), .B(n7985), .Z(n7983) );
  OR2_X1 U7895 ( .A1(n7986), .A2(n7987), .ZN(n7985) );
  OR2_X1 U7896 ( .A1(n7988), .A2(n7989), .ZN(Result_33_) );
  AND2_X1 U7897 ( .A1(n7990), .A2(n7554), .ZN(n7989) );
  XNOR2_X1 U7898 ( .A(n7991), .B(n7992), .ZN(n7990) );
  XOR2_X1 U7899 ( .A(n7993), .B(n7994), .Z(n7992) );
  AND2_X1 U7900 ( .A1(n7995), .A2(n7584), .ZN(n7988) );
  XOR2_X1 U7901 ( .A(n7996), .B(n7997), .Z(n7995) );
  AND2_X1 U7902 ( .A1(n7998), .A2(n7999), .ZN(n7997) );
  OR2_X1 U7903 ( .A1(n8000), .A2(n8001), .ZN(Result_32_) );
  AND2_X1 U7904 ( .A1(n8002), .A2(n7554), .ZN(n8001) );
  XNOR2_X1 U7905 ( .A(n8003), .B(n8004), .ZN(n8002) );
  XOR2_X1 U7906 ( .A(n8005), .B(n8006), .Z(n8004) );
  AND2_X1 U7907 ( .A1(n8007), .A2(n7584), .ZN(n8000) );
  XNOR2_X1 U7908 ( .A(n8008), .B(n8009), .ZN(n8007) );
  OR2_X1 U7909 ( .A1(n8010), .A2(n8011), .ZN(n8009) );
  AND2_X1 U7910 ( .A1(n8012), .A2(n8013), .ZN(n8011) );
  AND2_X1 U7911 ( .A1(n7996), .A2(n8014), .ZN(n8010) );
  OR2_X1 U7912 ( .A1(n8015), .A2(n7986), .ZN(n7996) );
  AND2_X1 U7913 ( .A1(n8016), .A2(n8017), .ZN(n7986) );
  AND2_X1 U7914 ( .A1(n7984), .A2(n8018), .ZN(n8015) );
  OR2_X1 U7915 ( .A1(n8019), .A2(n8020), .ZN(n7984) );
  AND2_X1 U7916 ( .A1(n8021), .A2(n8022), .ZN(n8020) );
  AND2_X1 U7917 ( .A1(n7972), .A2(n8023), .ZN(n8019) );
  OR2_X1 U7918 ( .A1(n8024), .A2(n7962), .ZN(n7972) );
  AND2_X1 U7919 ( .A1(n8025), .A2(n8026), .ZN(n7962) );
  AND2_X1 U7920 ( .A1(n7960), .A2(n8027), .ZN(n8024) );
  OR2_X1 U7921 ( .A1(n8028), .A2(n8029), .ZN(n7960) );
  AND2_X1 U7922 ( .A1(n8030), .A2(n8031), .ZN(n8029) );
  AND2_X1 U7923 ( .A1(n7948), .A2(n8032), .ZN(n8028) );
  OR2_X1 U7924 ( .A1(n8033), .A2(n7938), .ZN(n7948) );
  AND2_X1 U7925 ( .A1(n8034), .A2(n8035), .ZN(n7938) );
  AND2_X1 U7926 ( .A1(n7936), .A2(n8036), .ZN(n8033) );
  OR2_X1 U7927 ( .A1(n8037), .A2(n8038), .ZN(n7936) );
  AND2_X1 U7928 ( .A1(n8039), .A2(n8040), .ZN(n8038) );
  AND2_X1 U7929 ( .A1(n7924), .A2(n8041), .ZN(n8037) );
  OR2_X1 U7930 ( .A1(n8042), .A2(n7904), .ZN(n7924) );
  AND2_X1 U7931 ( .A1(n8043), .A2(n8044), .ZN(n7904) );
  AND2_X1 U7932 ( .A1(n7902), .A2(n8045), .ZN(n8042) );
  OR2_X1 U7933 ( .A1(n8046), .A2(n8047), .ZN(n7902) );
  AND2_X1 U7934 ( .A1(n8048), .A2(n8049), .ZN(n8047) );
  AND2_X1 U7935 ( .A1(n7890), .A2(n8050), .ZN(n8046) );
  OR2_X1 U7936 ( .A1(n8051), .A2(n7880), .ZN(n7890) );
  AND2_X1 U7937 ( .A1(n8052), .A2(n8053), .ZN(n7880) );
  AND2_X1 U7938 ( .A1(n7878), .A2(n8054), .ZN(n8051) );
  OR2_X1 U7939 ( .A1(n8055), .A2(n8056), .ZN(n7878) );
  AND2_X1 U7940 ( .A1(n8057), .A2(n8058), .ZN(n8056) );
  AND2_X1 U7941 ( .A1(n7866), .A2(n8059), .ZN(n8055) );
  OR2_X1 U7942 ( .A1(n8060), .A2(n7856), .ZN(n7866) );
  AND2_X1 U7943 ( .A1(n8061), .A2(n8062), .ZN(n7856) );
  AND2_X1 U7944 ( .A1(n7854), .A2(n8063), .ZN(n8060) );
  OR2_X1 U7945 ( .A1(n8064), .A2(n8065), .ZN(n7854) );
  AND2_X1 U7946 ( .A1(n8066), .A2(n8067), .ZN(n8065) );
  AND2_X1 U7947 ( .A1(n7842), .A2(n8068), .ZN(n8064) );
  OR2_X1 U7948 ( .A1(n8069), .A2(n7832), .ZN(n7842) );
  AND2_X1 U7949 ( .A1(n8070), .A2(n8071), .ZN(n7832) );
  AND2_X1 U7950 ( .A1(n7830), .A2(n8072), .ZN(n8069) );
  OR2_X1 U7951 ( .A1(n8073), .A2(n8074), .ZN(n7830) );
  AND2_X1 U7952 ( .A1(n8075), .A2(n8076), .ZN(n8074) );
  AND2_X1 U7953 ( .A1(n7818), .A2(n8077), .ZN(n8073) );
  OR2_X1 U7954 ( .A1(n8078), .A2(n7808), .ZN(n7818) );
  AND2_X1 U7955 ( .A1(n8079), .A2(n8080), .ZN(n7808) );
  AND2_X1 U7956 ( .A1(n7806), .A2(n8081), .ZN(n8078) );
  OR2_X1 U7957 ( .A1(n8082), .A2(n8083), .ZN(n7806) );
  AND2_X1 U7958 ( .A1(n8084), .A2(n8085), .ZN(n8083) );
  AND2_X1 U7959 ( .A1(n7794), .A2(n8086), .ZN(n8082) );
  OR2_X1 U7960 ( .A1(n8087), .A2(n7781), .ZN(n7794) );
  AND2_X1 U7961 ( .A1(n8088), .A2(n8089), .ZN(n7781) );
  AND2_X1 U7962 ( .A1(n7779), .A2(n8090), .ZN(n8087) );
  OR2_X1 U7963 ( .A1(n8091), .A2(n8092), .ZN(n7779) );
  AND2_X1 U7964 ( .A1(n8093), .A2(n8094), .ZN(n8092) );
  AND2_X1 U7965 ( .A1(n7767), .A2(n8095), .ZN(n8091) );
  OR2_X1 U7966 ( .A1(n8096), .A2(n7757), .ZN(n7767) );
  AND2_X1 U7967 ( .A1(n8097), .A2(n8098), .ZN(n7757) );
  AND2_X1 U7968 ( .A1(n7755), .A2(n8099), .ZN(n8096) );
  OR2_X1 U7969 ( .A1(n8100), .A2(n8101), .ZN(n7755) );
  AND2_X1 U7970 ( .A1(n8102), .A2(n8103), .ZN(n8101) );
  AND2_X1 U7971 ( .A1(n7743), .A2(n8104), .ZN(n8100) );
  OR2_X1 U7972 ( .A1(n8105), .A2(n7733), .ZN(n7743) );
  AND2_X1 U7973 ( .A1(n8106), .A2(n8107), .ZN(n7733) );
  AND2_X1 U7974 ( .A1(n7730), .A2(n7734), .ZN(n8105) );
  OR2_X1 U7975 ( .A1(n8108), .A2(n7714), .ZN(n7730) );
  AND2_X1 U7976 ( .A1(n8109), .A2(n8110), .ZN(n7714) );
  AND2_X1 U7977 ( .A1(n7711), .A2(n7716), .ZN(n8108) );
  OR2_X1 U7978 ( .A1(n8111), .A2(n7703), .ZN(n7711) );
  AND2_X1 U7979 ( .A1(n8112), .A2(n8113), .ZN(n7703) );
  AND2_X1 U7980 ( .A1(n7700), .A2(n7704), .ZN(n8111) );
  OR2_X1 U7981 ( .A1(n8114), .A2(n7684), .ZN(n7700) );
  AND2_X1 U7982 ( .A1(n8115), .A2(n8116), .ZN(n7684) );
  AND2_X1 U7983 ( .A1(n7681), .A2(n7686), .ZN(n8114) );
  OR2_X1 U7984 ( .A1(n8117), .A2(n7673), .ZN(n7681) );
  AND2_X1 U7985 ( .A1(n8118), .A2(n8119), .ZN(n7673) );
  AND2_X1 U7986 ( .A1(n7670), .A2(n7674), .ZN(n8117) );
  OR2_X1 U7987 ( .A1(n8120), .A2(n7654), .ZN(n7670) );
  AND2_X1 U7988 ( .A1(n8121), .A2(n8122), .ZN(n7654) );
  AND2_X1 U7989 ( .A1(n7651), .A2(n7656), .ZN(n8120) );
  OR2_X1 U7990 ( .A1(n8123), .A2(n7633), .ZN(n7651) );
  AND2_X1 U7991 ( .A1(n8124), .A2(n8125), .ZN(n7633) );
  AND2_X1 U7992 ( .A1(n7630), .A2(n7634), .ZN(n8123) );
  OR2_X1 U7993 ( .A1(n8126), .A2(n7614), .ZN(n7630) );
  AND2_X1 U7994 ( .A1(n8127), .A2(n7611), .ZN(n7614) );
  AND2_X1 U7995 ( .A1(n7607), .A2(n7616), .ZN(n8126) );
  INV_X1 U7996 ( .A(n7613), .ZN(n7607) );
  OR2_X1 U7997 ( .A1(n8128), .A2(n8129), .ZN(n7613) );
  AND2_X1 U7998 ( .A1(b_31_), .A2(n8130), .ZN(n8129) );
  AND2_X1 U7999 ( .A1(b_30_), .A2(n8131), .ZN(n8128) );
  OR2_X1 U8000 ( .A1(n7588), .A2(a_30_), .ZN(n8131) );
  AND2_X1 U8001 ( .A1(a_31_), .A2(b_31_), .ZN(n7588) );
  AND2_X1 U8002 ( .A1(n7554), .A2(n8132), .ZN(Result_31_) );
  XOR2_X1 U8003 ( .A(n8133), .B(n8134), .Z(n8132) );
  AND3_X1 U8004 ( .A1(n8135), .A2(n8136), .A3(n7554), .ZN(Result_30_) );
  INV_X1 U8005 ( .A(n8137), .ZN(n8136) );
  OR2_X1 U8006 ( .A1(n8138), .A2(n8139), .ZN(n8135) );
  AND2_X1 U8007 ( .A1(n8133), .A2(n8134), .ZN(n8138) );
  AND2_X1 U8008 ( .A1(n8140), .A2(n7554), .ZN(Result_2_) );
  XOR2_X1 U8009 ( .A(n8141), .B(n8142), .Z(n8140) );
  AND2_X1 U8010 ( .A1(n7554), .A2(n8143), .ZN(Result_29_) );
  XOR2_X1 U8011 ( .A(n8137), .B(n8144), .Z(n8143) );
  AND2_X1 U8012 ( .A1(n8145), .A2(n8146), .ZN(n8144) );
  AND2_X1 U8013 ( .A1(n8147), .A2(n7554), .ZN(Result_28_) );
  XOR2_X1 U8014 ( .A(n8148), .B(n8149), .Z(n8147) );
  AND2_X1 U8015 ( .A1(n8150), .A2(n8151), .ZN(n8149) );
  INV_X1 U8016 ( .A(n8152), .ZN(n8151) );
  AND2_X1 U8017 ( .A1(n8153), .A2(n7554), .ZN(Result_27_) );
  XOR2_X1 U8018 ( .A(n8154), .B(n8155), .Z(n8153) );
  AND2_X1 U8019 ( .A1(n8156), .A2(n8157), .ZN(n8155) );
  INV_X1 U8020 ( .A(n8158), .ZN(n8157) );
  AND2_X1 U8021 ( .A1(n8159), .A2(n7554), .ZN(Result_26_) );
  XOR2_X1 U8022 ( .A(n8160), .B(n8161), .Z(n8159) );
  AND2_X1 U8023 ( .A1(n8162), .A2(n8163), .ZN(n8161) );
  INV_X1 U8024 ( .A(n8164), .ZN(n8163) );
  AND2_X1 U8025 ( .A1(n8165), .A2(n7554), .ZN(Result_25_) );
  XOR2_X1 U8026 ( .A(n8166), .B(n8167), .Z(n8165) );
  AND2_X1 U8027 ( .A1(n8168), .A2(n8169), .ZN(n8167) );
  INV_X1 U8028 ( .A(n8170), .ZN(n8168) );
  AND2_X1 U8029 ( .A1(n8171), .A2(n7554), .ZN(Result_24_) );
  XOR2_X1 U8030 ( .A(n8172), .B(n8173), .Z(n8171) );
  AND2_X1 U8031 ( .A1(n8174), .A2(n8175), .ZN(n8173) );
  AND2_X1 U8032 ( .A1(n8176), .A2(n7554), .ZN(Result_23_) );
  XOR2_X1 U8033 ( .A(n8177), .B(n8178), .Z(n8176) );
  AND2_X1 U8034 ( .A1(n8179), .A2(n8180), .ZN(n8178) );
  AND2_X1 U8035 ( .A1(n8181), .A2(n7554), .ZN(Result_22_) );
  XOR2_X1 U8036 ( .A(n8182), .B(n8183), .Z(n8181) );
  AND2_X1 U8037 ( .A1(n8184), .A2(n8185), .ZN(n8183) );
  AND2_X1 U8038 ( .A1(n8186), .A2(n7554), .ZN(Result_21_) );
  XOR2_X1 U8039 ( .A(n8187), .B(n8188), .Z(n8186) );
  AND2_X1 U8040 ( .A1(n8189), .A2(n8190), .ZN(n8188) );
  INV_X1 U8041 ( .A(n8191), .ZN(n8189) );
  AND2_X1 U8042 ( .A1(n8192), .A2(n7554), .ZN(Result_20_) );
  XOR2_X1 U8043 ( .A(n8193), .B(n8194), .Z(n8192) );
  AND2_X1 U8044 ( .A1(n8195), .A2(n8196), .ZN(n8194) );
  AND2_X1 U8045 ( .A1(n7554), .A2(n8197), .ZN(Result_1_) );
  XOR2_X1 U8046 ( .A(n8198), .B(n8199), .Z(n8197) );
  AND2_X1 U8047 ( .A1(n8200), .A2(n8201), .ZN(n8199) );
  OR2_X1 U8048 ( .A1(n8202), .A2(n8203), .ZN(n8201) );
  AND2_X1 U8049 ( .A1(n8204), .A2(n8205), .ZN(n8203) );
  INV_X1 U8050 ( .A(n8206), .ZN(n8200) );
  AND2_X1 U8051 ( .A1(n8207), .A2(n7554), .ZN(Result_19_) );
  XOR2_X1 U8052 ( .A(n8208), .B(n8209), .Z(n8207) );
  AND2_X1 U8053 ( .A1(n8210), .A2(n8211), .ZN(n8209) );
  AND2_X1 U8054 ( .A1(n8212), .A2(n7554), .ZN(Result_18_) );
  XOR2_X1 U8055 ( .A(n8213), .B(n8214), .Z(n8212) );
  AND2_X1 U8056 ( .A1(n8215), .A2(n8216), .ZN(n8214) );
  AND2_X1 U8057 ( .A1(n8217), .A2(n7554), .ZN(Result_17_) );
  XOR2_X1 U8058 ( .A(n8218), .B(n8219), .Z(n8217) );
  AND2_X1 U8059 ( .A1(n8220), .A2(n8221), .ZN(n8219) );
  AND2_X1 U8060 ( .A1(n8222), .A2(n7554), .ZN(Result_16_) );
  XOR2_X1 U8061 ( .A(n8223), .B(n8224), .Z(n8222) );
  AND2_X1 U8062 ( .A1(n8225), .A2(n8226), .ZN(n8224) );
  AND2_X1 U8063 ( .A1(n8227), .A2(n7554), .ZN(Result_15_) );
  XOR2_X1 U8064 ( .A(n8228), .B(n8229), .Z(n8227) );
  AND2_X1 U8065 ( .A1(n8230), .A2(n8231), .ZN(n8229) );
  AND2_X1 U8066 ( .A1(n8232), .A2(n7554), .ZN(Result_14_) );
  XOR2_X1 U8067 ( .A(n8233), .B(n8234), .Z(n8232) );
  AND2_X1 U8068 ( .A1(n8235), .A2(n8236), .ZN(n8234) );
  INV_X1 U8069 ( .A(n8237), .ZN(n8236) );
  OR2_X1 U8070 ( .A1(n8238), .A2(n8239), .ZN(n8235) );
  AND2_X1 U8071 ( .A1(n8240), .A2(n8241), .ZN(n8238) );
  AND2_X1 U8072 ( .A1(n8242), .A2(n7554), .ZN(Result_13_) );
  XOR2_X1 U8073 ( .A(n8243), .B(n8244), .Z(n8242) );
  AND2_X1 U8074 ( .A1(n8245), .A2(n8246), .ZN(n8244) );
  INV_X1 U8075 ( .A(n8247), .ZN(n8246) );
  OR2_X1 U8076 ( .A1(n8248), .A2(n8249), .ZN(n8245) );
  AND2_X1 U8077 ( .A1(n8250), .A2(n8251), .ZN(n8248) );
  AND2_X1 U8078 ( .A1(n8252), .A2(n7554), .ZN(Result_12_) );
  XOR2_X1 U8079 ( .A(n8253), .B(n8254), .Z(n8252) );
  AND2_X1 U8080 ( .A1(n7554), .A2(n8255), .ZN(Result_11_) );
  XOR2_X1 U8081 ( .A(n8256), .B(n8257), .Z(n8255) );
  AND2_X1 U8082 ( .A1(n8258), .A2(n8259), .ZN(n8257) );
  INV_X1 U8083 ( .A(n8260), .ZN(n8259) );
  OR2_X1 U8084 ( .A1(n8261), .A2(n8262), .ZN(n8258) );
  AND2_X1 U8085 ( .A1(n8263), .A2(n8264), .ZN(n8261) );
  AND2_X1 U8086 ( .A1(n8265), .A2(n7554), .ZN(Result_10_) );
  XOR2_X1 U8087 ( .A(n8266), .B(n8267), .Z(n8265) );
  AND2_X1 U8088 ( .A1(n7554), .A2(n8268), .ZN(Result_0_) );
  OR3_X1 U8089 ( .A1(n8206), .A2(n8269), .A3(n8270), .ZN(n8268) );
  AND2_X1 U8090 ( .A1(n8198), .A2(n8202), .ZN(n8270) );
  AND2_X1 U8091 ( .A1(n8141), .A2(n8142), .ZN(n8198) );
  XOR2_X1 U8092 ( .A(n8205), .B(n8204), .Z(n8142) );
  OR2_X1 U8093 ( .A1(n8271), .A2(n8272), .ZN(n8141) );
  INV_X1 U8094 ( .A(n8273), .ZN(n8272) );
  OR2_X1 U8095 ( .A1(n8274), .A2(n7915), .ZN(n8271) );
  AND3_X1 U8096 ( .A1(n7914), .A2(n7913), .A3(n7911), .ZN(n7915) );
  AND2_X1 U8097 ( .A1(n7907), .A2(n7911), .ZN(n8274) );
  AND2_X1 U8098 ( .A1(n8275), .A2(n8273), .ZN(n7911) );
  OR2_X1 U8099 ( .A1(n8276), .A2(n8277), .ZN(n8273) );
  INV_X1 U8100 ( .A(n8278), .ZN(n8275) );
  AND2_X1 U8101 ( .A1(n8276), .A2(n8277), .ZN(n8278) );
  OR2_X1 U8102 ( .A1(n8279), .A2(n8280), .ZN(n8277) );
  AND2_X1 U8103 ( .A1(n8281), .A2(n8282), .ZN(n8280) );
  AND2_X1 U8104 ( .A1(n8283), .A2(n8284), .ZN(n8279) );
  OR2_X1 U8105 ( .A1(n8282), .A2(n8281), .ZN(n8284) );
  XNOR2_X1 U8106 ( .A(n8285), .B(n8286), .ZN(n8276) );
  XNOR2_X1 U8107 ( .A(n8287), .B(n8288), .ZN(n8286) );
  AND2_X1 U8108 ( .A1(n7784), .A2(n7785), .ZN(n7907) );
  XOR2_X1 U8109 ( .A(n7914), .B(n7913), .Z(n7785) );
  INV_X1 U8110 ( .A(n8289), .ZN(n7913) );
  OR2_X1 U8111 ( .A1(n8290), .A2(n8291), .ZN(n8289) );
  AND2_X1 U8112 ( .A1(n8292), .A2(n8293), .ZN(n8291) );
  AND2_X1 U8113 ( .A1(n8294), .A2(n8295), .ZN(n8290) );
  OR2_X1 U8114 ( .A1(n8293), .A2(n8292), .ZN(n8295) );
  XNOR2_X1 U8115 ( .A(n8283), .B(n8296), .ZN(n7914) );
  XOR2_X1 U8116 ( .A(n8282), .B(n8281), .Z(n8296) );
  OR2_X1 U8117 ( .A1(n8022), .A2(n8297), .ZN(n8281) );
  OR2_X1 U8118 ( .A1(n8298), .A2(n8299), .ZN(n8282) );
  AND2_X1 U8119 ( .A1(n8300), .A2(n8301), .ZN(n8299) );
  AND2_X1 U8120 ( .A1(n8302), .A2(n8303), .ZN(n8298) );
  OR2_X1 U8121 ( .A1(n8301), .A2(n8300), .ZN(n8303) );
  XOR2_X1 U8122 ( .A(n8304), .B(n8305), .Z(n8283) );
  XOR2_X1 U8123 ( .A(n8306), .B(n8307), .Z(n8305) );
  OR2_X1 U8124 ( .A1(n8308), .A2(n8309), .ZN(n7784) );
  INV_X1 U8125 ( .A(n8310), .ZN(n8309) );
  OR2_X1 U8126 ( .A1(n8311), .A2(n7644), .ZN(n8308) );
  AND3_X1 U8127 ( .A1(n7643), .A2(n7642), .A3(n7640), .ZN(n7644) );
  AND2_X1 U8128 ( .A1(n7636), .A2(n7640), .ZN(n8311) );
  AND2_X1 U8129 ( .A1(n8312), .A2(n8310), .ZN(n7640) );
  OR2_X1 U8130 ( .A1(n8313), .A2(n8314), .ZN(n8310) );
  INV_X1 U8131 ( .A(n8315), .ZN(n8312) );
  AND2_X1 U8132 ( .A1(n8313), .A2(n8314), .ZN(n8315) );
  OR2_X1 U8133 ( .A1(n8316), .A2(n8317), .ZN(n8314) );
  AND2_X1 U8134 ( .A1(n8318), .A2(n8319), .ZN(n8317) );
  AND2_X1 U8135 ( .A1(n8320), .A2(n8321), .ZN(n8316) );
  OR2_X1 U8136 ( .A1(n8319), .A2(n8318), .ZN(n8321) );
  XOR2_X1 U8137 ( .A(n8294), .B(n8322), .Z(n8313) );
  XOR2_X1 U8138 ( .A(n8293), .B(n8292), .Z(n8322) );
  OR2_X1 U8139 ( .A1(n8026), .A2(n8297), .ZN(n8292) );
  OR2_X1 U8140 ( .A1(n8323), .A2(n8324), .ZN(n8293) );
  AND2_X1 U8141 ( .A1(n8325), .A2(n8326), .ZN(n8324) );
  AND2_X1 U8142 ( .A1(n8327), .A2(n8328), .ZN(n8323) );
  OR2_X1 U8143 ( .A1(n8326), .A2(n8325), .ZN(n8328) );
  XOR2_X1 U8144 ( .A(n8302), .B(n8329), .Z(n8294) );
  XOR2_X1 U8145 ( .A(n8301), .B(n8300), .Z(n8329) );
  OR2_X1 U8146 ( .A1(n8022), .A2(n8012), .ZN(n8300) );
  OR2_X1 U8147 ( .A1(n8330), .A2(n8331), .ZN(n8301) );
  AND2_X1 U8148 ( .A1(n8332), .A2(n8333), .ZN(n8331) );
  AND2_X1 U8149 ( .A1(n8334), .A2(n8335), .ZN(n8330) );
  OR2_X1 U8150 ( .A1(n8333), .A2(n8332), .ZN(n8335) );
  XNOR2_X1 U8151 ( .A(n8336), .B(n8337), .ZN(n8302) );
  XOR2_X1 U8152 ( .A(n7987), .B(n8338), .Z(n8336) );
  INV_X1 U8153 ( .A(n8018), .ZN(n7987) );
  AND2_X1 U8154 ( .A1(n7579), .A2(n7580), .ZN(n7636) );
  XOR2_X1 U8155 ( .A(n7643), .B(n7642), .Z(n7580) );
  INV_X1 U8156 ( .A(n8339), .ZN(n7642) );
  OR2_X1 U8157 ( .A1(n8340), .A2(n8341), .ZN(n8339) );
  AND2_X1 U8158 ( .A1(n8342), .A2(n8343), .ZN(n8341) );
  AND2_X1 U8159 ( .A1(n8344), .A2(n8345), .ZN(n8340) );
  OR2_X1 U8160 ( .A1(n8343), .A2(n8342), .ZN(n8345) );
  XNOR2_X1 U8161 ( .A(n8320), .B(n8346), .ZN(n7643) );
  XOR2_X1 U8162 ( .A(n8319), .B(n8318), .Z(n8346) );
  OR2_X1 U8163 ( .A1(n8031), .A2(n8297), .ZN(n8318) );
  OR2_X1 U8164 ( .A1(n8347), .A2(n8348), .ZN(n8319) );
  AND2_X1 U8165 ( .A1(n8349), .A2(n8350), .ZN(n8348) );
  AND2_X1 U8166 ( .A1(n8351), .A2(n8352), .ZN(n8347) );
  OR2_X1 U8167 ( .A1(n8350), .A2(n8349), .ZN(n8352) );
  XOR2_X1 U8168 ( .A(n8327), .B(n8353), .Z(n8320) );
  XOR2_X1 U8169 ( .A(n8326), .B(n8325), .Z(n8353) );
  OR2_X1 U8170 ( .A1(n8026), .A2(n8012), .ZN(n8325) );
  OR2_X1 U8171 ( .A1(n8354), .A2(n8355), .ZN(n8326) );
  AND2_X1 U8172 ( .A1(n8356), .A2(n8357), .ZN(n8355) );
  AND2_X1 U8173 ( .A1(n8358), .A2(n8359), .ZN(n8354) );
  OR2_X1 U8174 ( .A1(n8357), .A2(n8356), .ZN(n8359) );
  XOR2_X1 U8175 ( .A(n8334), .B(n8360), .Z(n8327) );
  XOR2_X1 U8176 ( .A(n8333), .B(n8332), .Z(n8360) );
  OR2_X1 U8177 ( .A1(n8022), .A2(n8016), .ZN(n8332) );
  OR2_X1 U8178 ( .A1(n8361), .A2(n8362), .ZN(n8333) );
  AND2_X1 U8179 ( .A1(n8023), .A2(n8363), .ZN(n8362) );
  AND2_X1 U8180 ( .A1(n8364), .A2(n8365), .ZN(n8361) );
  OR2_X1 U8181 ( .A1(n8363), .A2(n8023), .ZN(n8365) );
  XOR2_X1 U8182 ( .A(n8366), .B(n8367), .Z(n8334) );
  XOR2_X1 U8183 ( .A(n8368), .B(n8369), .Z(n8367) );
  OR2_X1 U8184 ( .A1(n8370), .A2(n8371), .ZN(n7579) );
  INV_X1 U8185 ( .A(n8372), .ZN(n8371) );
  OR2_X1 U8186 ( .A1(n8373), .A2(n7577), .ZN(n8370) );
  AND3_X1 U8187 ( .A1(n7576), .A2(n7575), .A3(n7573), .ZN(n7577) );
  AND2_X1 U8188 ( .A1(n7569), .A2(n7573), .ZN(n8373) );
  AND2_X1 U8189 ( .A1(n8374), .A2(n8372), .ZN(n7573) );
  OR2_X1 U8190 ( .A1(n8375), .A2(n8376), .ZN(n8372) );
  INV_X1 U8191 ( .A(n8377), .ZN(n8374) );
  AND2_X1 U8192 ( .A1(n8375), .A2(n8376), .ZN(n8377) );
  OR2_X1 U8193 ( .A1(n8378), .A2(n8379), .ZN(n8376) );
  AND2_X1 U8194 ( .A1(n8380), .A2(n8381), .ZN(n8379) );
  AND2_X1 U8195 ( .A1(n8382), .A2(n8383), .ZN(n8378) );
  OR2_X1 U8196 ( .A1(n8381), .A2(n8380), .ZN(n8383) );
  XOR2_X1 U8197 ( .A(n8344), .B(n8384), .Z(n8375) );
  XOR2_X1 U8198 ( .A(n8343), .B(n8342), .Z(n8384) );
  OR2_X1 U8199 ( .A1(n8035), .A2(n8297), .ZN(n8342) );
  OR2_X1 U8200 ( .A1(n8385), .A2(n8386), .ZN(n8343) );
  AND2_X1 U8201 ( .A1(n8387), .A2(n8388), .ZN(n8386) );
  AND2_X1 U8202 ( .A1(n8389), .A2(n8390), .ZN(n8385) );
  OR2_X1 U8203 ( .A1(n8388), .A2(n8387), .ZN(n8390) );
  XOR2_X1 U8204 ( .A(n8351), .B(n8391), .Z(n8344) );
  XOR2_X1 U8205 ( .A(n8350), .B(n8349), .Z(n8391) );
  OR2_X1 U8206 ( .A1(n8031), .A2(n8012), .ZN(n8349) );
  OR2_X1 U8207 ( .A1(n8392), .A2(n8393), .ZN(n8350) );
  AND2_X1 U8208 ( .A1(n8394), .A2(n8395), .ZN(n8393) );
  AND2_X1 U8209 ( .A1(n8396), .A2(n8397), .ZN(n8392) );
  OR2_X1 U8210 ( .A1(n8395), .A2(n8394), .ZN(n8397) );
  XOR2_X1 U8211 ( .A(n8358), .B(n8398), .Z(n8351) );
  XOR2_X1 U8212 ( .A(n8357), .B(n8356), .Z(n8398) );
  OR2_X1 U8213 ( .A1(n8026), .A2(n8016), .ZN(n8356) );
  OR2_X1 U8214 ( .A1(n8399), .A2(n8400), .ZN(n8357) );
  AND2_X1 U8215 ( .A1(n8401), .A2(n8402), .ZN(n8400) );
  AND2_X1 U8216 ( .A1(n8403), .A2(n8404), .ZN(n8399) );
  OR2_X1 U8217 ( .A1(n8402), .A2(n8401), .ZN(n8404) );
  XOR2_X1 U8218 ( .A(n8364), .B(n8405), .Z(n8358) );
  XOR2_X1 U8219 ( .A(n8363), .B(n8023), .Z(n8405) );
  OR2_X1 U8220 ( .A1(n8021), .A2(n8022), .ZN(n8023) );
  OR2_X1 U8221 ( .A1(n8406), .A2(n8407), .ZN(n8363) );
  AND2_X1 U8222 ( .A1(n8408), .A2(n8409), .ZN(n8407) );
  AND2_X1 U8223 ( .A1(n8410), .A2(n8411), .ZN(n8406) );
  OR2_X1 U8224 ( .A1(n8409), .A2(n8408), .ZN(n8411) );
  XOR2_X1 U8225 ( .A(n8412), .B(n8413), .Z(n8364) );
  XOR2_X1 U8226 ( .A(n8414), .B(n8415), .Z(n8413) );
  AND2_X1 U8227 ( .A1(n7566), .A2(n7567), .ZN(n7569) );
  XOR2_X1 U8228 ( .A(n7576), .B(n7575), .Z(n7567) );
  INV_X1 U8229 ( .A(n8416), .ZN(n7575) );
  OR2_X1 U8230 ( .A1(n8417), .A2(n8418), .ZN(n8416) );
  AND2_X1 U8231 ( .A1(n8419), .A2(n8420), .ZN(n8418) );
  AND2_X1 U8232 ( .A1(n8421), .A2(n8422), .ZN(n8417) );
  OR2_X1 U8233 ( .A1(n8420), .A2(n8419), .ZN(n8422) );
  XNOR2_X1 U8234 ( .A(n8382), .B(n8423), .ZN(n7576) );
  XOR2_X1 U8235 ( .A(n8381), .B(n8380), .Z(n8423) );
  OR2_X1 U8236 ( .A1(n8040), .A2(n8297), .ZN(n8380) );
  OR2_X1 U8237 ( .A1(n8424), .A2(n8425), .ZN(n8381) );
  AND2_X1 U8238 ( .A1(n8426), .A2(n8427), .ZN(n8425) );
  AND2_X1 U8239 ( .A1(n8428), .A2(n8429), .ZN(n8424) );
  OR2_X1 U8240 ( .A1(n8427), .A2(n8426), .ZN(n8429) );
  XOR2_X1 U8241 ( .A(n8389), .B(n8430), .Z(n8382) );
  XOR2_X1 U8242 ( .A(n8388), .B(n8387), .Z(n8430) );
  OR2_X1 U8243 ( .A1(n8035), .A2(n8012), .ZN(n8387) );
  OR2_X1 U8244 ( .A1(n8431), .A2(n8432), .ZN(n8388) );
  AND2_X1 U8245 ( .A1(n8433), .A2(n8434), .ZN(n8432) );
  AND2_X1 U8246 ( .A1(n8435), .A2(n8436), .ZN(n8431) );
  OR2_X1 U8247 ( .A1(n8434), .A2(n8433), .ZN(n8436) );
  XOR2_X1 U8248 ( .A(n8396), .B(n8437), .Z(n8389) );
  XOR2_X1 U8249 ( .A(n8395), .B(n8394), .Z(n8437) );
  OR2_X1 U8250 ( .A1(n8031), .A2(n8016), .ZN(n8394) );
  OR2_X1 U8251 ( .A1(n8438), .A2(n8439), .ZN(n8395) );
  AND2_X1 U8252 ( .A1(n8440), .A2(n8441), .ZN(n8439) );
  AND2_X1 U8253 ( .A1(n8442), .A2(n8443), .ZN(n8438) );
  OR2_X1 U8254 ( .A1(n8441), .A2(n8440), .ZN(n8443) );
  XOR2_X1 U8255 ( .A(n8403), .B(n8444), .Z(n8396) );
  XOR2_X1 U8256 ( .A(n8402), .B(n8401), .Z(n8444) );
  OR2_X1 U8257 ( .A1(n8021), .A2(n8026), .ZN(n8401) );
  OR2_X1 U8258 ( .A1(n8445), .A2(n8446), .ZN(n8402) );
  AND2_X1 U8259 ( .A1(n8447), .A2(n8027), .ZN(n8446) );
  AND2_X1 U8260 ( .A1(n8448), .A2(n8449), .ZN(n8445) );
  OR2_X1 U8261 ( .A1(n8027), .A2(n8447), .ZN(n8449) );
  XOR2_X1 U8262 ( .A(n8410), .B(n8450), .Z(n8403) );
  XOR2_X1 U8263 ( .A(n8409), .B(n8408), .Z(n8450) );
  OR2_X1 U8264 ( .A1(n8022), .A2(n8025), .ZN(n8408) );
  OR2_X1 U8265 ( .A1(n8451), .A2(n8452), .ZN(n8409) );
  AND2_X1 U8266 ( .A1(n8453), .A2(n8454), .ZN(n8452) );
  AND2_X1 U8267 ( .A1(n8455), .A2(n8456), .ZN(n8451) );
  OR2_X1 U8268 ( .A1(n8454), .A2(n8453), .ZN(n8456) );
  XOR2_X1 U8269 ( .A(n8457), .B(n8458), .Z(n8410) );
  XOR2_X1 U8270 ( .A(n8459), .B(n8460), .Z(n8458) );
  OR2_X1 U8271 ( .A1(n8461), .A2(n8462), .ZN(n7566) );
  INV_X1 U8272 ( .A(n8463), .ZN(n8462) );
  OR2_X1 U8273 ( .A1(n8464), .A2(n7564), .ZN(n8461) );
  AND3_X1 U8274 ( .A1(n7563), .A2(n7562), .A3(n7560), .ZN(n7564) );
  AND2_X1 U8275 ( .A1(n7556), .A2(n7560), .ZN(n8464) );
  AND2_X1 U8276 ( .A1(n8465), .A2(n8463), .ZN(n7560) );
  OR2_X1 U8277 ( .A1(n8466), .A2(n8467), .ZN(n8463) );
  INV_X1 U8278 ( .A(n8468), .ZN(n8465) );
  AND2_X1 U8279 ( .A1(n8466), .A2(n8467), .ZN(n8468) );
  OR2_X1 U8280 ( .A1(n8469), .A2(n8470), .ZN(n8467) );
  AND2_X1 U8281 ( .A1(n8471), .A2(n8472), .ZN(n8470) );
  AND2_X1 U8282 ( .A1(n8473), .A2(n8474), .ZN(n8469) );
  OR2_X1 U8283 ( .A1(n8472), .A2(n8471), .ZN(n8474) );
  XOR2_X1 U8284 ( .A(n8421), .B(n8475), .Z(n8466) );
  XOR2_X1 U8285 ( .A(n8420), .B(n8419), .Z(n8475) );
  OR2_X1 U8286 ( .A1(n8044), .A2(n8297), .ZN(n8419) );
  OR2_X1 U8287 ( .A1(n8476), .A2(n8477), .ZN(n8420) );
  AND2_X1 U8288 ( .A1(n8478), .A2(n8479), .ZN(n8477) );
  AND2_X1 U8289 ( .A1(n8480), .A2(n8481), .ZN(n8476) );
  OR2_X1 U8290 ( .A1(n8479), .A2(n8478), .ZN(n8481) );
  XOR2_X1 U8291 ( .A(n8428), .B(n8482), .Z(n8421) );
  XOR2_X1 U8292 ( .A(n8427), .B(n8426), .Z(n8482) );
  OR2_X1 U8293 ( .A1(n8040), .A2(n8012), .ZN(n8426) );
  OR2_X1 U8294 ( .A1(n8483), .A2(n8484), .ZN(n8427) );
  AND2_X1 U8295 ( .A1(n8485), .A2(n8486), .ZN(n8484) );
  AND2_X1 U8296 ( .A1(n8487), .A2(n8488), .ZN(n8483) );
  OR2_X1 U8297 ( .A1(n8486), .A2(n8485), .ZN(n8488) );
  XOR2_X1 U8298 ( .A(n8435), .B(n8489), .Z(n8428) );
  XOR2_X1 U8299 ( .A(n8434), .B(n8433), .Z(n8489) );
  OR2_X1 U8300 ( .A1(n8035), .A2(n8016), .ZN(n8433) );
  OR2_X1 U8301 ( .A1(n8490), .A2(n8491), .ZN(n8434) );
  AND2_X1 U8302 ( .A1(n8492), .A2(n8493), .ZN(n8491) );
  AND2_X1 U8303 ( .A1(n8494), .A2(n8495), .ZN(n8490) );
  OR2_X1 U8304 ( .A1(n8493), .A2(n8492), .ZN(n8495) );
  XOR2_X1 U8305 ( .A(n8442), .B(n8496), .Z(n8435) );
  XOR2_X1 U8306 ( .A(n8441), .B(n8440), .Z(n8496) );
  OR2_X1 U8307 ( .A1(n8021), .A2(n8031), .ZN(n8440) );
  OR2_X1 U8308 ( .A1(n8497), .A2(n8498), .ZN(n8441) );
  AND2_X1 U8309 ( .A1(n8499), .A2(n8500), .ZN(n8498) );
  AND2_X1 U8310 ( .A1(n8501), .A2(n8502), .ZN(n8497) );
  OR2_X1 U8311 ( .A1(n8500), .A2(n8499), .ZN(n8502) );
  XNOR2_X1 U8312 ( .A(n8503), .B(n8448), .ZN(n8442) );
  XOR2_X1 U8313 ( .A(n8455), .B(n8504), .Z(n8448) );
  XOR2_X1 U8314 ( .A(n8454), .B(n8453), .Z(n8504) );
  OR2_X1 U8315 ( .A1(n8022), .A2(n8030), .ZN(n8453) );
  OR2_X1 U8316 ( .A1(n8505), .A2(n8506), .ZN(n8454) );
  AND2_X1 U8317 ( .A1(n8507), .A2(n8508), .ZN(n8506) );
  AND2_X1 U8318 ( .A1(n8509), .A2(n8510), .ZN(n8505) );
  OR2_X1 U8319 ( .A1(n8508), .A2(n8507), .ZN(n8510) );
  XOR2_X1 U8320 ( .A(n8511), .B(n8512), .Z(n8455) );
  XOR2_X1 U8321 ( .A(n8513), .B(n8514), .Z(n8512) );
  XOR2_X1 U8322 ( .A(n7963), .B(n8447), .Z(n8503) );
  OR2_X1 U8323 ( .A1(n8515), .A2(n8516), .ZN(n8447) );
  AND2_X1 U8324 ( .A1(n8517), .A2(n8518), .ZN(n8516) );
  AND2_X1 U8325 ( .A1(n8519), .A2(n8520), .ZN(n8515) );
  OR2_X1 U8326 ( .A1(n8518), .A2(n8517), .ZN(n8520) );
  INV_X1 U8327 ( .A(n8027), .ZN(n7963) );
  OR2_X1 U8328 ( .A1(n8026), .A2(n8025), .ZN(n8027) );
  AND2_X1 U8329 ( .A1(n8266), .A2(n8267), .ZN(n7556) );
  XOR2_X1 U8330 ( .A(n7563), .B(n7562), .Z(n8267) );
  INV_X1 U8331 ( .A(n8521), .ZN(n7562) );
  OR2_X1 U8332 ( .A1(n8522), .A2(n8523), .ZN(n8521) );
  AND2_X1 U8333 ( .A1(n8524), .A2(n8525), .ZN(n8523) );
  AND2_X1 U8334 ( .A1(n8526), .A2(n8527), .ZN(n8522) );
  OR2_X1 U8335 ( .A1(n8525), .A2(n8524), .ZN(n8527) );
  XNOR2_X1 U8336 ( .A(n8473), .B(n8528), .ZN(n7563) );
  XOR2_X1 U8337 ( .A(n8472), .B(n8471), .Z(n8528) );
  OR2_X1 U8338 ( .A1(n8049), .A2(n8297), .ZN(n8471) );
  OR2_X1 U8339 ( .A1(n8529), .A2(n8530), .ZN(n8472) );
  AND2_X1 U8340 ( .A1(n8531), .A2(n8532), .ZN(n8530) );
  AND2_X1 U8341 ( .A1(n8533), .A2(n8534), .ZN(n8529) );
  OR2_X1 U8342 ( .A1(n8532), .A2(n8531), .ZN(n8534) );
  XOR2_X1 U8343 ( .A(n8480), .B(n8535), .Z(n8473) );
  XOR2_X1 U8344 ( .A(n8479), .B(n8478), .Z(n8535) );
  OR2_X1 U8345 ( .A1(n8044), .A2(n8012), .ZN(n8478) );
  OR2_X1 U8346 ( .A1(n8536), .A2(n8537), .ZN(n8479) );
  AND2_X1 U8347 ( .A1(n8538), .A2(n8539), .ZN(n8537) );
  AND2_X1 U8348 ( .A1(n8540), .A2(n8541), .ZN(n8536) );
  OR2_X1 U8349 ( .A1(n8539), .A2(n8538), .ZN(n8541) );
  XOR2_X1 U8350 ( .A(n8487), .B(n8542), .Z(n8480) );
  XOR2_X1 U8351 ( .A(n8486), .B(n8485), .Z(n8542) );
  OR2_X1 U8352 ( .A1(n8040), .A2(n8016), .ZN(n8485) );
  OR2_X1 U8353 ( .A1(n8543), .A2(n8544), .ZN(n8486) );
  AND2_X1 U8354 ( .A1(n8545), .A2(n8546), .ZN(n8544) );
  AND2_X1 U8355 ( .A1(n8547), .A2(n8548), .ZN(n8543) );
  OR2_X1 U8356 ( .A1(n8546), .A2(n8545), .ZN(n8548) );
  XOR2_X1 U8357 ( .A(n8494), .B(n8549), .Z(n8487) );
  XOR2_X1 U8358 ( .A(n8493), .B(n8492), .Z(n8549) );
  OR2_X1 U8359 ( .A1(n8021), .A2(n8035), .ZN(n8492) );
  OR2_X1 U8360 ( .A1(n8550), .A2(n8551), .ZN(n8493) );
  AND2_X1 U8361 ( .A1(n8552), .A2(n8553), .ZN(n8551) );
  AND2_X1 U8362 ( .A1(n8554), .A2(n8555), .ZN(n8550) );
  OR2_X1 U8363 ( .A1(n8553), .A2(n8552), .ZN(n8555) );
  XOR2_X1 U8364 ( .A(n8501), .B(n8556), .Z(n8494) );
  XOR2_X1 U8365 ( .A(n8500), .B(n8499), .Z(n8556) );
  OR2_X1 U8366 ( .A1(n8031), .A2(n8025), .ZN(n8499) );
  OR2_X1 U8367 ( .A1(n8557), .A2(n8558), .ZN(n8500) );
  AND2_X1 U8368 ( .A1(n8032), .A2(n8559), .ZN(n8558) );
  AND2_X1 U8369 ( .A1(n8560), .A2(n8561), .ZN(n8557) );
  OR2_X1 U8370 ( .A1(n8559), .A2(n8032), .ZN(n8561) );
  XOR2_X1 U8371 ( .A(n8519), .B(n8562), .Z(n8501) );
  XOR2_X1 U8372 ( .A(n8518), .B(n8517), .Z(n8562) );
  OR2_X1 U8373 ( .A1(n8026), .A2(n8030), .ZN(n8517) );
  OR2_X1 U8374 ( .A1(n8563), .A2(n8564), .ZN(n8518) );
  AND2_X1 U8375 ( .A1(n8565), .A2(n8566), .ZN(n8564) );
  AND2_X1 U8376 ( .A1(n8567), .A2(n8568), .ZN(n8563) );
  OR2_X1 U8377 ( .A1(n8566), .A2(n8565), .ZN(n8568) );
  XOR2_X1 U8378 ( .A(n8509), .B(n8569), .Z(n8519) );
  XOR2_X1 U8379 ( .A(n8508), .B(n8507), .Z(n8569) );
  OR2_X1 U8380 ( .A1(n8022), .A2(n8034), .ZN(n8507) );
  OR2_X1 U8381 ( .A1(n8570), .A2(n8571), .ZN(n8508) );
  AND2_X1 U8382 ( .A1(n8572), .A2(n8573), .ZN(n8571) );
  AND2_X1 U8383 ( .A1(n8574), .A2(n8575), .ZN(n8570) );
  OR2_X1 U8384 ( .A1(n8573), .A2(n8572), .ZN(n8575) );
  XOR2_X1 U8385 ( .A(n8576), .B(n8577), .Z(n8509) );
  XOR2_X1 U8386 ( .A(n8578), .B(n8579), .Z(n8577) );
  OR2_X1 U8387 ( .A1(n8580), .A2(n8581), .ZN(n8266) );
  OR2_X1 U8388 ( .A1(n8582), .A2(n8260), .ZN(n8581) );
  AND3_X1 U8389 ( .A1(n8264), .A2(n8263), .A3(n8262), .ZN(n8260) );
  AND2_X1 U8390 ( .A1(n8256), .A2(n8262), .ZN(n8582) );
  AND2_X1 U8391 ( .A1(n8583), .A2(n8584), .ZN(n8262) );
  INV_X1 U8392 ( .A(n8585), .ZN(n8583) );
  AND2_X1 U8393 ( .A1(n8586), .A2(n8587), .ZN(n8585) );
  AND2_X1 U8394 ( .A1(n8253), .A2(n8254), .ZN(n8256) );
  XOR2_X1 U8395 ( .A(n8264), .B(n8263), .Z(n8254) );
  INV_X1 U8396 ( .A(n8588), .ZN(n8263) );
  OR2_X1 U8397 ( .A1(n8589), .A2(n8590), .ZN(n8588) );
  AND2_X1 U8398 ( .A1(n8591), .A2(n8592), .ZN(n8590) );
  AND2_X1 U8399 ( .A1(n8593), .A2(n8594), .ZN(n8589) );
  OR2_X1 U8400 ( .A1(n8592), .A2(n8591), .ZN(n8594) );
  XNOR2_X1 U8401 ( .A(n8595), .B(n8596), .ZN(n8264) );
  XOR2_X1 U8402 ( .A(n8597), .B(n8598), .Z(n8596) );
  OR2_X1 U8403 ( .A1(n8599), .A2(n8600), .ZN(n8253) );
  OR2_X1 U8404 ( .A1(n8601), .A2(n8247), .ZN(n8600) );
  AND3_X1 U8405 ( .A1(n8251), .A2(n8250), .A3(n8249), .ZN(n8247) );
  AND2_X1 U8406 ( .A1(n8249), .A2(n8243), .ZN(n8601) );
  OR2_X1 U8407 ( .A1(n8602), .A2(n8237), .ZN(n8243) );
  AND3_X1 U8408 ( .A1(n8241), .A2(n8239), .A3(n8240), .ZN(n8237) );
  INV_X1 U8409 ( .A(n8603), .ZN(n8240) );
  AND2_X1 U8410 ( .A1(n8239), .A2(n8233), .ZN(n8602) );
  OR2_X1 U8411 ( .A1(n8604), .A2(n8605), .ZN(n8233) );
  INV_X1 U8412 ( .A(n8231), .ZN(n8605) );
  OR3_X1 U8413 ( .A1(n8606), .A2(n8607), .A3(n8608), .ZN(n8231) );
  AND2_X1 U8414 ( .A1(n8228), .A2(n8230), .ZN(n8604) );
  INV_X1 U8415 ( .A(n8609), .ZN(n8230) );
  AND2_X1 U8416 ( .A1(n8610), .A2(n8607), .ZN(n8609) );
  XOR2_X1 U8417 ( .A(n8241), .B(n8603), .Z(n8607) );
  OR2_X1 U8418 ( .A1(n8611), .A2(n8612), .ZN(n8603) );
  AND2_X1 U8419 ( .A1(n8613), .A2(n8614), .ZN(n8612) );
  AND2_X1 U8420 ( .A1(n8615), .A2(n8616), .ZN(n8611) );
  OR2_X1 U8421 ( .A1(n8614), .A2(n8613), .ZN(n8616) );
  XNOR2_X1 U8422 ( .A(n8617), .B(n8618), .ZN(n8241) );
  XOR2_X1 U8423 ( .A(n8619), .B(n8620), .Z(n8618) );
  OR2_X1 U8424 ( .A1(n8608), .A2(n8606), .ZN(n8610) );
  OR2_X1 U8425 ( .A1(n8621), .A2(n8622), .ZN(n8228) );
  INV_X1 U8426 ( .A(n8225), .ZN(n8622) );
  OR3_X1 U8427 ( .A1(n8623), .A2(n8624), .A3(n8625), .ZN(n8225) );
  AND2_X1 U8428 ( .A1(n8223), .A2(n8226), .ZN(n8621) );
  INV_X1 U8429 ( .A(n8626), .ZN(n8226) );
  AND2_X1 U8430 ( .A1(n8627), .A2(n8624), .ZN(n8626) );
  XNOR2_X1 U8431 ( .A(n8606), .B(n8608), .ZN(n8624) );
  OR2_X1 U8432 ( .A1(n8628), .A2(n8629), .ZN(n8608) );
  AND2_X1 U8433 ( .A1(n8630), .A2(n8631), .ZN(n8629) );
  AND2_X1 U8434 ( .A1(n8632), .A2(n8633), .ZN(n8628) );
  OR2_X1 U8435 ( .A1(n8630), .A2(n8631), .ZN(n8633) );
  XOR2_X1 U8436 ( .A(n8615), .B(n8634), .Z(n8606) );
  XOR2_X1 U8437 ( .A(n8614), .B(n8613), .Z(n8634) );
  OR2_X1 U8438 ( .A1(n8076), .A2(n8297), .ZN(n8613) );
  OR2_X1 U8439 ( .A1(n8635), .A2(n8636), .ZN(n8614) );
  AND2_X1 U8440 ( .A1(n8637), .A2(n8638), .ZN(n8636) );
  AND2_X1 U8441 ( .A1(n8639), .A2(n8640), .ZN(n8635) );
  OR2_X1 U8442 ( .A1(n8638), .A2(n8637), .ZN(n8640) );
  XOR2_X1 U8443 ( .A(n8641), .B(n8642), .Z(n8615) );
  XOR2_X1 U8444 ( .A(n8643), .B(n8644), .Z(n8642) );
  OR2_X1 U8445 ( .A1(n8625), .A2(n8623), .ZN(n8627) );
  OR2_X1 U8446 ( .A1(n8645), .A2(n8646), .ZN(n8223) );
  INV_X1 U8447 ( .A(n8220), .ZN(n8646) );
  OR3_X1 U8448 ( .A1(n8647), .A2(n8648), .A3(n8649), .ZN(n8220) );
  AND2_X1 U8449 ( .A1(n8218), .A2(n8221), .ZN(n8645) );
  INV_X1 U8450 ( .A(n8650), .ZN(n8221) );
  AND2_X1 U8451 ( .A1(n8651), .A2(n8648), .ZN(n8650) );
  XNOR2_X1 U8452 ( .A(n8623), .B(n8625), .ZN(n8648) );
  OR2_X1 U8453 ( .A1(n8652), .A2(n8653), .ZN(n8625) );
  AND2_X1 U8454 ( .A1(n8654), .A2(n8655), .ZN(n8653) );
  AND2_X1 U8455 ( .A1(n8656), .A2(n8657), .ZN(n8652) );
  OR2_X1 U8456 ( .A1(n8654), .A2(n8655), .ZN(n8657) );
  XOR2_X1 U8457 ( .A(n8632), .B(n8658), .Z(n8623) );
  XOR2_X1 U8458 ( .A(n8631), .B(n8630), .Z(n8658) );
  OR2_X1 U8459 ( .A1(n8080), .A2(n8297), .ZN(n8630) );
  OR2_X1 U8460 ( .A1(n8659), .A2(n8660), .ZN(n8631) );
  AND2_X1 U8461 ( .A1(n8661), .A2(n8662), .ZN(n8660) );
  AND2_X1 U8462 ( .A1(n8663), .A2(n8664), .ZN(n8659) );
  OR2_X1 U8463 ( .A1(n8661), .A2(n8662), .ZN(n8664) );
  XOR2_X1 U8464 ( .A(n8639), .B(n8665), .Z(n8632) );
  XOR2_X1 U8465 ( .A(n8638), .B(n8637), .Z(n8665) );
  OR2_X1 U8466 ( .A1(n8076), .A2(n8012), .ZN(n8637) );
  OR2_X1 U8467 ( .A1(n8666), .A2(n8667), .ZN(n8638) );
  AND2_X1 U8468 ( .A1(n8668), .A2(n8669), .ZN(n8667) );
  AND2_X1 U8469 ( .A1(n8670), .A2(n8671), .ZN(n8666) );
  OR2_X1 U8470 ( .A1(n8669), .A2(n8668), .ZN(n8671) );
  XOR2_X1 U8471 ( .A(n8672), .B(n8673), .Z(n8639) );
  XOR2_X1 U8472 ( .A(n8674), .B(n8675), .Z(n8673) );
  OR2_X1 U8473 ( .A1(n8649), .A2(n8647), .ZN(n8651) );
  OR2_X1 U8474 ( .A1(n8676), .A2(n8677), .ZN(n8218) );
  INV_X1 U8475 ( .A(n8216), .ZN(n8677) );
  OR3_X1 U8476 ( .A1(n8678), .A2(n8679), .A3(n8680), .ZN(n8216) );
  AND2_X1 U8477 ( .A1(n8213), .A2(n8215), .ZN(n8676) );
  INV_X1 U8478 ( .A(n8681), .ZN(n8215) );
  AND2_X1 U8479 ( .A1(n8682), .A2(n8679), .ZN(n8681) );
  XNOR2_X1 U8480 ( .A(n8647), .B(n8649), .ZN(n8679) );
  OR2_X1 U8481 ( .A1(n8683), .A2(n8684), .ZN(n8649) );
  AND2_X1 U8482 ( .A1(n8685), .A2(n8686), .ZN(n8684) );
  AND2_X1 U8483 ( .A1(n8687), .A2(n8688), .ZN(n8683) );
  OR2_X1 U8484 ( .A1(n8685), .A2(n8686), .ZN(n8688) );
  XOR2_X1 U8485 ( .A(n8656), .B(n8689), .Z(n8647) );
  XOR2_X1 U8486 ( .A(n8655), .B(n8654), .Z(n8689) );
  OR2_X1 U8487 ( .A1(n8085), .A2(n8297), .ZN(n8654) );
  OR2_X1 U8488 ( .A1(n8690), .A2(n8691), .ZN(n8655) );
  AND2_X1 U8489 ( .A1(n8692), .A2(n8693), .ZN(n8691) );
  AND2_X1 U8490 ( .A1(n8694), .A2(n8695), .ZN(n8690) );
  OR2_X1 U8491 ( .A1(n8692), .A2(n8693), .ZN(n8695) );
  XOR2_X1 U8492 ( .A(n8663), .B(n8696), .Z(n8656) );
  XOR2_X1 U8493 ( .A(n8662), .B(n8661), .Z(n8696) );
  OR2_X1 U8494 ( .A1(n8080), .A2(n8012), .ZN(n8661) );
  OR2_X1 U8495 ( .A1(n8697), .A2(n8698), .ZN(n8662) );
  AND2_X1 U8496 ( .A1(n8699), .A2(n8700), .ZN(n8698) );
  AND2_X1 U8497 ( .A1(n8701), .A2(n8702), .ZN(n8697) );
  OR2_X1 U8498 ( .A1(n8699), .A2(n8700), .ZN(n8702) );
  XOR2_X1 U8499 ( .A(n8670), .B(n8703), .Z(n8663) );
  XOR2_X1 U8500 ( .A(n8669), .B(n8668), .Z(n8703) );
  OR2_X1 U8501 ( .A1(n8076), .A2(n8016), .ZN(n8668) );
  OR2_X1 U8502 ( .A1(n8704), .A2(n8705), .ZN(n8669) );
  AND2_X1 U8503 ( .A1(n8706), .A2(n8707), .ZN(n8705) );
  AND2_X1 U8504 ( .A1(n8708), .A2(n8709), .ZN(n8704) );
  OR2_X1 U8505 ( .A1(n8707), .A2(n8706), .ZN(n8709) );
  XOR2_X1 U8506 ( .A(n8710), .B(n8711), .Z(n8670) );
  XOR2_X1 U8507 ( .A(n8712), .B(n8713), .Z(n8711) );
  OR2_X1 U8508 ( .A1(n8680), .A2(n8678), .ZN(n8682) );
  OR2_X1 U8509 ( .A1(n8714), .A2(n8715), .ZN(n8213) );
  INV_X1 U8510 ( .A(n8210), .ZN(n8715) );
  OR3_X1 U8511 ( .A1(n8716), .A2(n8717), .A3(n8718), .ZN(n8210) );
  AND2_X1 U8512 ( .A1(n8208), .A2(n8211), .ZN(n8714) );
  INV_X1 U8513 ( .A(n8719), .ZN(n8211) );
  AND2_X1 U8514 ( .A1(n8720), .A2(n8717), .ZN(n8719) );
  XNOR2_X1 U8515 ( .A(n8678), .B(n8680), .ZN(n8717) );
  OR2_X1 U8516 ( .A1(n8721), .A2(n8722), .ZN(n8680) );
  AND2_X1 U8517 ( .A1(n8723), .A2(n8724), .ZN(n8722) );
  AND2_X1 U8518 ( .A1(n8725), .A2(n8726), .ZN(n8721) );
  OR2_X1 U8519 ( .A1(n8723), .A2(n8724), .ZN(n8726) );
  XOR2_X1 U8520 ( .A(n8687), .B(n8727), .Z(n8678) );
  XOR2_X1 U8521 ( .A(n8686), .B(n8685), .Z(n8727) );
  OR2_X1 U8522 ( .A1(n8089), .A2(n8297), .ZN(n8685) );
  OR2_X1 U8523 ( .A1(n8728), .A2(n8729), .ZN(n8686) );
  AND2_X1 U8524 ( .A1(n8730), .A2(n8731), .ZN(n8729) );
  AND2_X1 U8525 ( .A1(n8732), .A2(n8733), .ZN(n8728) );
  OR2_X1 U8526 ( .A1(n8730), .A2(n8731), .ZN(n8733) );
  XOR2_X1 U8527 ( .A(n8694), .B(n8734), .Z(n8687) );
  XOR2_X1 U8528 ( .A(n8693), .B(n8692), .Z(n8734) );
  OR2_X1 U8529 ( .A1(n8085), .A2(n8012), .ZN(n8692) );
  OR2_X1 U8530 ( .A1(n8735), .A2(n8736), .ZN(n8693) );
  AND2_X1 U8531 ( .A1(n8737), .A2(n8738), .ZN(n8736) );
  AND2_X1 U8532 ( .A1(n8739), .A2(n8740), .ZN(n8735) );
  OR2_X1 U8533 ( .A1(n8737), .A2(n8738), .ZN(n8740) );
  XOR2_X1 U8534 ( .A(n8701), .B(n8741), .Z(n8694) );
  XOR2_X1 U8535 ( .A(n8700), .B(n8699), .Z(n8741) );
  OR2_X1 U8536 ( .A1(n8080), .A2(n8016), .ZN(n8699) );
  OR2_X1 U8537 ( .A1(n8742), .A2(n8743), .ZN(n8700) );
  AND2_X1 U8538 ( .A1(n8744), .A2(n8745), .ZN(n8743) );
  AND2_X1 U8539 ( .A1(n8746), .A2(n8747), .ZN(n8742) );
  OR2_X1 U8540 ( .A1(n8744), .A2(n8745), .ZN(n8747) );
  XOR2_X1 U8541 ( .A(n8708), .B(n8748), .Z(n8701) );
  XOR2_X1 U8542 ( .A(n8707), .B(n8706), .Z(n8748) );
  OR2_X1 U8543 ( .A1(n8021), .A2(n8076), .ZN(n8706) );
  OR2_X1 U8544 ( .A1(n8749), .A2(n8750), .ZN(n8707) );
  AND2_X1 U8545 ( .A1(n8751), .A2(n8752), .ZN(n8750) );
  AND2_X1 U8546 ( .A1(n8753), .A2(n8754), .ZN(n8749) );
  OR2_X1 U8547 ( .A1(n8752), .A2(n8751), .ZN(n8754) );
  XOR2_X1 U8548 ( .A(n8755), .B(n8756), .Z(n8708) );
  XOR2_X1 U8549 ( .A(n8757), .B(n8758), .Z(n8756) );
  OR2_X1 U8550 ( .A1(n8718), .A2(n8716), .ZN(n8720) );
  OR2_X1 U8551 ( .A1(n8759), .A2(n8760), .ZN(n8208) );
  INV_X1 U8552 ( .A(n8195), .ZN(n8760) );
  OR3_X1 U8553 ( .A1(n8761), .A2(n8762), .A3(n8763), .ZN(n8195) );
  AND2_X1 U8554 ( .A1(n8193), .A2(n8196), .ZN(n8759) );
  INV_X1 U8555 ( .A(n8764), .ZN(n8196) );
  AND2_X1 U8556 ( .A1(n8765), .A2(n8762), .ZN(n8764) );
  XNOR2_X1 U8557 ( .A(n8716), .B(n8718), .ZN(n8762) );
  OR2_X1 U8558 ( .A1(n8766), .A2(n8767), .ZN(n8718) );
  AND2_X1 U8559 ( .A1(n8768), .A2(n8769), .ZN(n8767) );
  AND2_X1 U8560 ( .A1(n8770), .A2(n8771), .ZN(n8766) );
  OR2_X1 U8561 ( .A1(n8768), .A2(n8769), .ZN(n8771) );
  XOR2_X1 U8562 ( .A(n8725), .B(n8772), .Z(n8716) );
  XOR2_X1 U8563 ( .A(n8724), .B(n8723), .Z(n8772) );
  OR2_X1 U8564 ( .A1(n8094), .A2(n8297), .ZN(n8723) );
  OR2_X1 U8565 ( .A1(n8773), .A2(n8774), .ZN(n8724) );
  AND2_X1 U8566 ( .A1(n8775), .A2(n8776), .ZN(n8774) );
  AND2_X1 U8567 ( .A1(n8777), .A2(n8778), .ZN(n8773) );
  OR2_X1 U8568 ( .A1(n8775), .A2(n8776), .ZN(n8778) );
  XOR2_X1 U8569 ( .A(n8732), .B(n8779), .Z(n8725) );
  XOR2_X1 U8570 ( .A(n8731), .B(n8730), .Z(n8779) );
  OR2_X1 U8571 ( .A1(n8089), .A2(n8012), .ZN(n8730) );
  OR2_X1 U8572 ( .A1(n8780), .A2(n8781), .ZN(n8731) );
  AND2_X1 U8573 ( .A1(n8782), .A2(n8783), .ZN(n8781) );
  AND2_X1 U8574 ( .A1(n8784), .A2(n8785), .ZN(n8780) );
  OR2_X1 U8575 ( .A1(n8782), .A2(n8783), .ZN(n8785) );
  XOR2_X1 U8576 ( .A(n8739), .B(n8786), .Z(n8732) );
  XOR2_X1 U8577 ( .A(n8738), .B(n8737), .Z(n8786) );
  OR2_X1 U8578 ( .A1(n8085), .A2(n8016), .ZN(n8737) );
  OR2_X1 U8579 ( .A1(n8787), .A2(n8788), .ZN(n8738) );
  AND2_X1 U8580 ( .A1(n8789), .A2(n8790), .ZN(n8788) );
  AND2_X1 U8581 ( .A1(n8791), .A2(n8792), .ZN(n8787) );
  OR2_X1 U8582 ( .A1(n8789), .A2(n8790), .ZN(n8792) );
  XOR2_X1 U8583 ( .A(n8746), .B(n8793), .Z(n8739) );
  XOR2_X1 U8584 ( .A(n8745), .B(n8744), .Z(n8793) );
  OR2_X1 U8585 ( .A1(n8021), .A2(n8080), .ZN(n8744) );
  OR2_X1 U8586 ( .A1(n8794), .A2(n8795), .ZN(n8745) );
  AND2_X1 U8587 ( .A1(n8796), .A2(n8797), .ZN(n8795) );
  AND2_X1 U8588 ( .A1(n8798), .A2(n8799), .ZN(n8794) );
  OR2_X1 U8589 ( .A1(n8796), .A2(n8797), .ZN(n8799) );
  XOR2_X1 U8590 ( .A(n8753), .B(n8800), .Z(n8746) );
  XOR2_X1 U8591 ( .A(n8752), .B(n8751), .Z(n8800) );
  OR2_X1 U8592 ( .A1(n8076), .A2(n8025), .ZN(n8751) );
  OR2_X1 U8593 ( .A1(n8801), .A2(n8802), .ZN(n8752) );
  AND2_X1 U8594 ( .A1(n8803), .A2(n8804), .ZN(n8802) );
  AND2_X1 U8595 ( .A1(n8805), .A2(n8806), .ZN(n8801) );
  OR2_X1 U8596 ( .A1(n8804), .A2(n8803), .ZN(n8806) );
  XOR2_X1 U8597 ( .A(n8807), .B(n8808), .Z(n8753) );
  XOR2_X1 U8598 ( .A(n8809), .B(n8810), .Z(n8808) );
  OR2_X1 U8599 ( .A1(n8763), .A2(n8761), .ZN(n8765) );
  OR2_X1 U8600 ( .A1(n8811), .A2(n8191), .ZN(n8193) );
  AND3_X1 U8601 ( .A1(n8812), .A2(n8813), .A3(n8814), .ZN(n8191) );
  AND2_X1 U8602 ( .A1(n8190), .A2(n8187), .ZN(n8811) );
  OR2_X1 U8603 ( .A1(n8815), .A2(n8816), .ZN(n8187) );
  INV_X1 U8604 ( .A(n8185), .ZN(n8816) );
  OR3_X1 U8605 ( .A1(n8817), .A2(n8818), .A3(n8819), .ZN(n8185) );
  AND2_X1 U8606 ( .A1(n8182), .A2(n8184), .ZN(n8815) );
  INV_X1 U8607 ( .A(n8820), .ZN(n8184) );
  AND2_X1 U8608 ( .A1(n8821), .A2(n8818), .ZN(n8820) );
  XOR2_X1 U8609 ( .A(n8812), .B(n8822), .Z(n8818) );
  OR2_X1 U8610 ( .A1(n8819), .A2(n8817), .ZN(n8821) );
  OR2_X1 U8611 ( .A1(n8823), .A2(n8824), .ZN(n8182) );
  INV_X1 U8612 ( .A(n8179), .ZN(n8824) );
  OR3_X1 U8613 ( .A1(n8825), .A2(n8826), .A3(n8827), .ZN(n8179) );
  AND2_X1 U8614 ( .A1(n8177), .A2(n8180), .ZN(n8823) );
  INV_X1 U8615 ( .A(n8828), .ZN(n8180) );
  AND2_X1 U8616 ( .A1(n8829), .A2(n8826), .ZN(n8828) );
  XNOR2_X1 U8617 ( .A(n8817), .B(n8819), .ZN(n8826) );
  OR2_X1 U8618 ( .A1(n8830), .A2(n8831), .ZN(n8819) );
  AND2_X1 U8619 ( .A1(n8832), .A2(n8833), .ZN(n8831) );
  AND2_X1 U8620 ( .A1(n8834), .A2(n8835), .ZN(n8830) );
  OR2_X1 U8621 ( .A1(n8832), .A2(n8833), .ZN(n8835) );
  XOR2_X1 U8622 ( .A(n8836), .B(n8837), .Z(n8817) );
  XOR2_X1 U8623 ( .A(n8838), .B(n8839), .Z(n8837) );
  OR2_X1 U8624 ( .A1(n8827), .A2(n8825), .ZN(n8829) );
  OR2_X1 U8625 ( .A1(n8840), .A2(n8841), .ZN(n8177) );
  INV_X1 U8626 ( .A(n8174), .ZN(n8841) );
  OR3_X1 U8627 ( .A1(n8842), .A2(n8843), .A3(n8844), .ZN(n8174) );
  AND2_X1 U8628 ( .A1(n8172), .A2(n8175), .ZN(n8840) );
  INV_X1 U8629 ( .A(n8845), .ZN(n8175) );
  AND2_X1 U8630 ( .A1(n8846), .A2(n8843), .ZN(n8845) );
  XNOR2_X1 U8631 ( .A(n8825), .B(n8827), .ZN(n8843) );
  OR2_X1 U8632 ( .A1(n8847), .A2(n8848), .ZN(n8827) );
  AND2_X1 U8633 ( .A1(n8849), .A2(n8850), .ZN(n8848) );
  AND2_X1 U8634 ( .A1(n8851), .A2(n8852), .ZN(n8847) );
  OR2_X1 U8635 ( .A1(n8849), .A2(n8850), .ZN(n8852) );
  XOR2_X1 U8636 ( .A(n8834), .B(n8853), .Z(n8825) );
  XOR2_X1 U8637 ( .A(n8833), .B(n8832), .Z(n8853) );
  OR2_X1 U8638 ( .A1(n8297), .A2(n8110), .ZN(n8832) );
  OR2_X1 U8639 ( .A1(n8854), .A2(n8855), .ZN(n8833) );
  AND2_X1 U8640 ( .A1(n8856), .A2(n8857), .ZN(n8855) );
  AND2_X1 U8641 ( .A1(n8858), .A2(n8859), .ZN(n8854) );
  OR2_X1 U8642 ( .A1(n8856), .A2(n8857), .ZN(n8859) );
  XOR2_X1 U8643 ( .A(n8860), .B(n8861), .Z(n8834) );
  XOR2_X1 U8644 ( .A(n8862), .B(n8863), .Z(n8861) );
  OR2_X1 U8645 ( .A1(n8844), .A2(n8842), .ZN(n8846) );
  OR2_X1 U8646 ( .A1(n8864), .A2(n8170), .ZN(n8172) );
  AND3_X1 U8647 ( .A1(n8865), .A2(n8866), .A3(n8867), .ZN(n8170) );
  AND2_X1 U8648 ( .A1(n8169), .A2(n8166), .ZN(n8864) );
  OR2_X1 U8649 ( .A1(n8868), .A2(n8164), .ZN(n8166) );
  AND2_X1 U8650 ( .A1(n8869), .A2(n8870), .ZN(n8164) );
  AND2_X1 U8651 ( .A1(n8162), .A2(n8160), .ZN(n8868) );
  OR2_X1 U8652 ( .A1(n8871), .A2(n8158), .ZN(n8160) );
  AND3_X1 U8653 ( .A1(n8872), .A2(n8873), .A3(n8874), .ZN(n8158) );
  AND2_X1 U8654 ( .A1(n8156), .A2(n8154), .ZN(n8871) );
  OR2_X1 U8655 ( .A1(n8875), .A2(n8152), .ZN(n8154) );
  AND3_X1 U8656 ( .A1(n8876), .A2(n8877), .A3(n8878), .ZN(n8152) );
  AND2_X1 U8657 ( .A1(n8150), .A2(n8148), .ZN(n8875) );
  OR2_X1 U8658 ( .A1(n8879), .A2(n8880), .ZN(n8148) );
  INV_X1 U8659 ( .A(n8146), .ZN(n8880) );
  OR3_X1 U8660 ( .A1(n8881), .A2(n8882), .A3(n8883), .ZN(n8146) );
  XOR2_X1 U8661 ( .A(n8876), .B(n8884), .Z(n8881) );
  AND2_X1 U8662 ( .A1(n8137), .A2(n8145), .ZN(n8879) );
  OR2_X1 U8663 ( .A1(n8885), .A2(n8886), .ZN(n8145) );
  XOR2_X1 U8664 ( .A(n8878), .B(n8876), .Z(n8886) );
  INV_X1 U8665 ( .A(n8887), .ZN(n8885) );
  OR2_X1 U8666 ( .A1(n8883), .A2(n8882), .ZN(n8887) );
  AND3_X1 U8667 ( .A1(n8134), .A2(n8139), .A3(n8133), .ZN(n8137) );
  INV_X1 U8668 ( .A(n8888), .ZN(n8133) );
  OR2_X1 U8669 ( .A1(n8889), .A2(n8890), .ZN(n8888) );
  AND2_X1 U8670 ( .A1(n8006), .A2(n8005), .ZN(n8890) );
  AND2_X1 U8671 ( .A1(n8003), .A2(n8891), .ZN(n8889) );
  OR2_X1 U8672 ( .A1(n8006), .A2(n8005), .ZN(n8891) );
  OR2_X1 U8673 ( .A1(n8892), .A2(n8893), .ZN(n8005) );
  AND2_X1 U8674 ( .A1(n7994), .A2(n7993), .ZN(n8893) );
  AND2_X1 U8675 ( .A1(n7991), .A2(n8894), .ZN(n8892) );
  OR2_X1 U8676 ( .A1(n7994), .A2(n7993), .ZN(n8894) );
  OR2_X1 U8677 ( .A1(n8895), .A2(n8896), .ZN(n7993) );
  AND2_X1 U8678 ( .A1(n7982), .A2(n7981), .ZN(n8896) );
  AND2_X1 U8679 ( .A1(n7979), .A2(n8897), .ZN(n8895) );
  OR2_X1 U8680 ( .A1(n7982), .A2(n7981), .ZN(n8897) );
  OR2_X1 U8681 ( .A1(n8898), .A2(n8899), .ZN(n7981) );
  AND2_X1 U8682 ( .A1(n7970), .A2(n7969), .ZN(n8899) );
  AND2_X1 U8683 ( .A1(n7967), .A2(n8900), .ZN(n8898) );
  OR2_X1 U8684 ( .A1(n7970), .A2(n7969), .ZN(n8900) );
  OR2_X1 U8685 ( .A1(n8901), .A2(n8902), .ZN(n7969) );
  AND2_X1 U8686 ( .A1(n7958), .A2(n7957), .ZN(n8902) );
  AND2_X1 U8687 ( .A1(n7955), .A2(n8903), .ZN(n8901) );
  OR2_X1 U8688 ( .A1(n7958), .A2(n7957), .ZN(n8903) );
  OR2_X1 U8689 ( .A1(n8904), .A2(n8905), .ZN(n7957) );
  AND2_X1 U8690 ( .A1(n7946), .A2(n7945), .ZN(n8905) );
  AND2_X1 U8691 ( .A1(n7943), .A2(n8906), .ZN(n8904) );
  OR2_X1 U8692 ( .A1(n7946), .A2(n7945), .ZN(n8906) );
  OR2_X1 U8693 ( .A1(n8907), .A2(n8908), .ZN(n7945) );
  AND2_X1 U8694 ( .A1(n7934), .A2(n7933), .ZN(n8908) );
  AND2_X1 U8695 ( .A1(n7931), .A2(n8909), .ZN(n8907) );
  OR2_X1 U8696 ( .A1(n7934), .A2(n7933), .ZN(n8909) );
  OR2_X1 U8697 ( .A1(n8910), .A2(n8911), .ZN(n7933) );
  AND2_X1 U8698 ( .A1(n7922), .A2(n7921), .ZN(n8911) );
  AND2_X1 U8699 ( .A1(n7919), .A2(n8912), .ZN(n8910) );
  OR2_X1 U8700 ( .A1(n7922), .A2(n7921), .ZN(n8912) );
  OR2_X1 U8701 ( .A1(n8913), .A2(n8914), .ZN(n7921) );
  AND2_X1 U8702 ( .A1(n7900), .A2(n7899), .ZN(n8914) );
  AND2_X1 U8703 ( .A1(n7897), .A2(n8915), .ZN(n8913) );
  OR2_X1 U8704 ( .A1(n7900), .A2(n7899), .ZN(n8915) );
  OR2_X1 U8705 ( .A1(n8916), .A2(n8917), .ZN(n7899) );
  AND2_X1 U8706 ( .A1(n7888), .A2(n7887), .ZN(n8917) );
  AND2_X1 U8707 ( .A1(n7885), .A2(n8918), .ZN(n8916) );
  OR2_X1 U8708 ( .A1(n7888), .A2(n7887), .ZN(n8918) );
  OR2_X1 U8709 ( .A1(n8919), .A2(n8920), .ZN(n7887) );
  AND2_X1 U8710 ( .A1(n7876), .A2(n7875), .ZN(n8920) );
  AND2_X1 U8711 ( .A1(n7873), .A2(n8921), .ZN(n8919) );
  OR2_X1 U8712 ( .A1(n7876), .A2(n7875), .ZN(n8921) );
  OR2_X1 U8713 ( .A1(n8922), .A2(n8923), .ZN(n7875) );
  AND2_X1 U8714 ( .A1(n7864), .A2(n7863), .ZN(n8923) );
  AND2_X1 U8715 ( .A1(n7861), .A2(n8924), .ZN(n8922) );
  OR2_X1 U8716 ( .A1(n7864), .A2(n7863), .ZN(n8924) );
  OR2_X1 U8717 ( .A1(n8925), .A2(n8926), .ZN(n7863) );
  AND2_X1 U8718 ( .A1(n7852), .A2(n7851), .ZN(n8926) );
  AND2_X1 U8719 ( .A1(n7849), .A2(n8927), .ZN(n8925) );
  OR2_X1 U8720 ( .A1(n7852), .A2(n7851), .ZN(n8927) );
  OR2_X1 U8721 ( .A1(n8928), .A2(n8929), .ZN(n7851) );
  AND2_X1 U8722 ( .A1(n7840), .A2(n7839), .ZN(n8929) );
  AND2_X1 U8723 ( .A1(n7837), .A2(n8930), .ZN(n8928) );
  OR2_X1 U8724 ( .A1(n7840), .A2(n7839), .ZN(n8930) );
  OR2_X1 U8725 ( .A1(n8931), .A2(n8932), .ZN(n7839) );
  AND2_X1 U8726 ( .A1(n7828), .A2(n7827), .ZN(n8932) );
  AND2_X1 U8727 ( .A1(n7825), .A2(n8933), .ZN(n8931) );
  OR2_X1 U8728 ( .A1(n7828), .A2(n7827), .ZN(n8933) );
  OR2_X1 U8729 ( .A1(n8934), .A2(n8935), .ZN(n7827) );
  AND2_X1 U8730 ( .A1(n7816), .A2(n7815), .ZN(n8935) );
  AND2_X1 U8731 ( .A1(n7813), .A2(n8936), .ZN(n8934) );
  OR2_X1 U8732 ( .A1(n7816), .A2(n7815), .ZN(n8936) );
  OR2_X1 U8733 ( .A1(n8937), .A2(n8938), .ZN(n7815) );
  AND2_X1 U8734 ( .A1(n7804), .A2(n7803), .ZN(n8938) );
  AND2_X1 U8735 ( .A1(n7801), .A2(n8939), .ZN(n8937) );
  OR2_X1 U8736 ( .A1(n7804), .A2(n7803), .ZN(n8939) );
  OR2_X1 U8737 ( .A1(n8940), .A2(n8941), .ZN(n7803) );
  AND2_X1 U8738 ( .A1(n7792), .A2(n7791), .ZN(n8941) );
  AND2_X1 U8739 ( .A1(n7789), .A2(n8942), .ZN(n8940) );
  OR2_X1 U8740 ( .A1(n7792), .A2(n7791), .ZN(n8942) );
  OR2_X1 U8741 ( .A1(n8943), .A2(n8944), .ZN(n7791) );
  AND2_X1 U8742 ( .A1(n7777), .A2(n7776), .ZN(n8944) );
  AND2_X1 U8743 ( .A1(n7774), .A2(n8945), .ZN(n8943) );
  OR2_X1 U8744 ( .A1(n7777), .A2(n7776), .ZN(n8945) );
  OR2_X1 U8745 ( .A1(n8946), .A2(n8947), .ZN(n7776) );
  AND2_X1 U8746 ( .A1(n7765), .A2(n7764), .ZN(n8947) );
  AND2_X1 U8747 ( .A1(n7762), .A2(n8948), .ZN(n8946) );
  OR2_X1 U8748 ( .A1(n7765), .A2(n7764), .ZN(n8948) );
  OR2_X1 U8749 ( .A1(n8949), .A2(n8950), .ZN(n7764) );
  AND2_X1 U8750 ( .A1(n7753), .A2(n7752), .ZN(n8950) );
  AND2_X1 U8751 ( .A1(n7750), .A2(n8951), .ZN(n8949) );
  OR2_X1 U8752 ( .A1(n7753), .A2(n7752), .ZN(n8951) );
  OR2_X1 U8753 ( .A1(n8952), .A2(n8953), .ZN(n7752) );
  AND2_X1 U8754 ( .A1(n7741), .A2(n7740), .ZN(n8953) );
  AND2_X1 U8755 ( .A1(n7738), .A2(n8954), .ZN(n8952) );
  OR2_X1 U8756 ( .A1(n7741), .A2(n7740), .ZN(n8954) );
  OR2_X1 U8757 ( .A1(n8955), .A2(n8956), .ZN(n7740) );
  AND2_X1 U8758 ( .A1(n7728), .A2(n7727), .ZN(n8956) );
  AND2_X1 U8759 ( .A1(n7725), .A2(n8957), .ZN(n8955) );
  OR2_X1 U8760 ( .A1(n7728), .A2(n7727), .ZN(n8957) );
  OR2_X1 U8761 ( .A1(n8958), .A2(n8959), .ZN(n7727) );
  AND2_X1 U8762 ( .A1(n7721), .A2(n7720), .ZN(n8959) );
  AND2_X1 U8763 ( .A1(n7718), .A2(n8960), .ZN(n8958) );
  OR2_X1 U8764 ( .A1(n7721), .A2(n7720), .ZN(n8960) );
  OR2_X1 U8765 ( .A1(n8961), .A2(n8962), .ZN(n7720) );
  AND2_X1 U8766 ( .A1(n7698), .A2(n7697), .ZN(n8962) );
  AND2_X1 U8767 ( .A1(n7695), .A2(n8963), .ZN(n8961) );
  OR2_X1 U8768 ( .A1(n7698), .A2(n7697), .ZN(n8963) );
  OR2_X1 U8769 ( .A1(n8964), .A2(n8965), .ZN(n7697) );
  AND2_X1 U8770 ( .A1(n7691), .A2(n7690), .ZN(n8965) );
  AND2_X1 U8771 ( .A1(n7688), .A2(n8966), .ZN(n8964) );
  OR2_X1 U8772 ( .A1(n7691), .A2(n7690), .ZN(n8966) );
  OR2_X1 U8773 ( .A1(n8967), .A2(n8968), .ZN(n7690) );
  AND2_X1 U8774 ( .A1(n7668), .A2(n7667), .ZN(n8968) );
  AND2_X1 U8775 ( .A1(n7665), .A2(n8969), .ZN(n8967) );
  OR2_X1 U8776 ( .A1(n7668), .A2(n7667), .ZN(n8969) );
  OR2_X1 U8777 ( .A1(n8970), .A2(n8971), .ZN(n7667) );
  AND2_X1 U8778 ( .A1(n7661), .A2(n7660), .ZN(n8971) );
  AND2_X1 U8779 ( .A1(n7658), .A2(n8972), .ZN(n8970) );
  OR2_X1 U8780 ( .A1(n7661), .A2(n7660), .ZN(n8972) );
  OR2_X1 U8781 ( .A1(n8973), .A2(n8974), .ZN(n7660) );
  AND2_X1 U8782 ( .A1(n7628), .A2(n7627), .ZN(n8974) );
  AND2_X1 U8783 ( .A1(n7625), .A2(n8975), .ZN(n8973) );
  OR2_X1 U8784 ( .A1(n7628), .A2(n7627), .ZN(n8975) );
  OR2_X1 U8785 ( .A1(n8976), .A2(n8977), .ZN(n7627) );
  AND2_X1 U8786 ( .A1(n7618), .A2(n7621), .ZN(n8977) );
  AND2_X1 U8787 ( .A1(n8978), .A2(n8979), .ZN(n8976) );
  OR2_X1 U8788 ( .A1(n7618), .A2(n7621), .ZN(n8979) );
  OR2_X1 U8789 ( .A1(n8127), .A2(n8980), .ZN(n7621) );
  OR3_X1 U8790 ( .A1(n8981), .A2(n7599), .A3(n8980), .ZN(n7618) );
  INV_X1 U8791 ( .A(n7620), .ZN(n8978) );
  OR2_X1 U8792 ( .A1(n8982), .A2(n8983), .ZN(n7620) );
  AND2_X1 U8793 ( .A1(b_30_), .A2(n8984), .ZN(n8983) );
  OR2_X1 U8794 ( .A1(n8985), .A2(n7598), .ZN(n8984) );
  AND2_X1 U8795 ( .A1(a_30_), .A2(n7611), .ZN(n8985) );
  AND2_X1 U8796 ( .A1(b_29_), .A2(n8986), .ZN(n8982) );
  OR2_X1 U8797 ( .A1(n8987), .A2(n7601), .ZN(n8986) );
  AND2_X1 U8798 ( .A1(a_31_), .A2(n7599), .ZN(n8987) );
  OR2_X1 U8799 ( .A1(n8124), .A2(n8980), .ZN(n7628) );
  XNOR2_X1 U8800 ( .A(n8988), .B(n8989), .ZN(n7625) );
  XOR2_X1 U8801 ( .A(n8990), .B(n8991), .Z(n8989) );
  OR2_X1 U8802 ( .A1(n8121), .A2(n8980), .ZN(n7661) );
  XOR2_X1 U8803 ( .A(n8992), .B(n8993), .Z(n7658) );
  XOR2_X1 U8804 ( .A(n8994), .B(n8995), .Z(n8993) );
  OR2_X1 U8805 ( .A1(n8118), .A2(n8980), .ZN(n7668) );
  XOR2_X1 U8806 ( .A(n8996), .B(n8997), .Z(n7665) );
  XOR2_X1 U8807 ( .A(n8998), .B(n8999), .Z(n8997) );
  OR2_X1 U8808 ( .A1(n8115), .A2(n8980), .ZN(n7691) );
  XOR2_X1 U8809 ( .A(n9000), .B(n9001), .Z(n7688) );
  XOR2_X1 U8810 ( .A(n9002), .B(n9003), .Z(n9001) );
  OR2_X1 U8811 ( .A1(n8112), .A2(n8980), .ZN(n7698) );
  XOR2_X1 U8812 ( .A(n9004), .B(n9005), .Z(n7695) );
  XOR2_X1 U8813 ( .A(n9006), .B(n9007), .Z(n9005) );
  OR2_X1 U8814 ( .A1(n8109), .A2(n8980), .ZN(n7721) );
  XOR2_X1 U8815 ( .A(n9008), .B(n9009), .Z(n7718) );
  XOR2_X1 U8816 ( .A(n9010), .B(n9011), .Z(n9009) );
  OR2_X1 U8817 ( .A1(n8106), .A2(n8980), .ZN(n7728) );
  XOR2_X1 U8818 ( .A(n9012), .B(n9013), .Z(n7725) );
  XOR2_X1 U8819 ( .A(n9014), .B(n9015), .Z(n9013) );
  OR2_X1 U8820 ( .A1(n8102), .A2(n8980), .ZN(n7741) );
  XOR2_X1 U8821 ( .A(n9016), .B(n9017), .Z(n7738) );
  XOR2_X1 U8822 ( .A(n9018), .B(n9019), .Z(n9017) );
  OR2_X1 U8823 ( .A1(n8097), .A2(n8980), .ZN(n7753) );
  XOR2_X1 U8824 ( .A(n9020), .B(n9021), .Z(n7750) );
  XOR2_X1 U8825 ( .A(n9022), .B(n9023), .Z(n9021) );
  OR2_X1 U8826 ( .A1(n8093), .A2(n8980), .ZN(n7765) );
  XOR2_X1 U8827 ( .A(n9024), .B(n9025), .Z(n7762) );
  XOR2_X1 U8828 ( .A(n9026), .B(n9027), .Z(n9025) );
  OR2_X1 U8829 ( .A1(n8088), .A2(n8980), .ZN(n7777) );
  XOR2_X1 U8830 ( .A(n9028), .B(n9029), .Z(n7774) );
  XOR2_X1 U8831 ( .A(n9030), .B(n9031), .Z(n9029) );
  OR2_X1 U8832 ( .A1(n8084), .A2(n8980), .ZN(n7792) );
  XOR2_X1 U8833 ( .A(n9032), .B(n9033), .Z(n7789) );
  XOR2_X1 U8834 ( .A(n9034), .B(n9035), .Z(n9033) );
  OR2_X1 U8835 ( .A1(n8079), .A2(n8980), .ZN(n7804) );
  XOR2_X1 U8836 ( .A(n9036), .B(n9037), .Z(n7801) );
  XOR2_X1 U8837 ( .A(n9038), .B(n9039), .Z(n9037) );
  OR2_X1 U8838 ( .A1(n8075), .A2(n8980), .ZN(n7816) );
  XOR2_X1 U8839 ( .A(n9040), .B(n9041), .Z(n7813) );
  XOR2_X1 U8840 ( .A(n9042), .B(n9043), .Z(n9041) );
  OR2_X1 U8841 ( .A1(n8070), .A2(n8980), .ZN(n7828) );
  XOR2_X1 U8842 ( .A(n9044), .B(n9045), .Z(n7825) );
  XOR2_X1 U8843 ( .A(n9046), .B(n9047), .Z(n9045) );
  OR2_X1 U8844 ( .A1(n8066), .A2(n8980), .ZN(n7840) );
  XOR2_X1 U8845 ( .A(n9048), .B(n9049), .Z(n7837) );
  XOR2_X1 U8846 ( .A(n9050), .B(n9051), .Z(n9049) );
  OR2_X1 U8847 ( .A1(n8061), .A2(n8980), .ZN(n7852) );
  XOR2_X1 U8848 ( .A(n9052), .B(n9053), .Z(n7849) );
  XOR2_X1 U8849 ( .A(n9054), .B(n9055), .Z(n9053) );
  OR2_X1 U8850 ( .A1(n8057), .A2(n8980), .ZN(n7864) );
  XOR2_X1 U8851 ( .A(n9056), .B(n9057), .Z(n7861) );
  XOR2_X1 U8852 ( .A(n9058), .B(n9059), .Z(n9057) );
  OR2_X1 U8853 ( .A1(n8052), .A2(n8980), .ZN(n7876) );
  XOR2_X1 U8854 ( .A(n9060), .B(n9061), .Z(n7873) );
  XOR2_X1 U8855 ( .A(n9062), .B(n9063), .Z(n9061) );
  OR2_X1 U8856 ( .A1(n8048), .A2(n8980), .ZN(n7888) );
  XOR2_X1 U8857 ( .A(n9064), .B(n9065), .Z(n7885) );
  XOR2_X1 U8858 ( .A(n9066), .B(n9067), .Z(n9065) );
  OR2_X1 U8859 ( .A1(n8043), .A2(n8980), .ZN(n7900) );
  XOR2_X1 U8860 ( .A(n9068), .B(n9069), .Z(n7897) );
  XOR2_X1 U8861 ( .A(n9070), .B(n9071), .Z(n9069) );
  OR2_X1 U8862 ( .A1(n8039), .A2(n8980), .ZN(n7922) );
  XOR2_X1 U8863 ( .A(n9072), .B(n9073), .Z(n7919) );
  XOR2_X1 U8864 ( .A(n9074), .B(n9075), .Z(n9073) );
  OR2_X1 U8865 ( .A1(n8034), .A2(n8980), .ZN(n7934) );
  XOR2_X1 U8866 ( .A(n9076), .B(n9077), .Z(n7931) );
  XOR2_X1 U8867 ( .A(n9078), .B(n9079), .Z(n9077) );
  OR2_X1 U8868 ( .A1(n8030), .A2(n8980), .ZN(n7946) );
  XOR2_X1 U8869 ( .A(n9080), .B(n9081), .Z(n7943) );
  XOR2_X1 U8870 ( .A(n9082), .B(n9083), .Z(n9081) );
  OR2_X1 U8871 ( .A1(n8025), .A2(n8980), .ZN(n7958) );
  XOR2_X1 U8872 ( .A(n9084), .B(n9085), .Z(n7955) );
  XOR2_X1 U8873 ( .A(n9086), .B(n9087), .Z(n9085) );
  OR2_X1 U8874 ( .A1(n8021), .A2(n8980), .ZN(n7970) );
  XOR2_X1 U8875 ( .A(n9088), .B(n9089), .Z(n7967) );
  XOR2_X1 U8876 ( .A(n9090), .B(n9091), .Z(n9089) );
  OR2_X1 U8877 ( .A1(n8016), .A2(n8980), .ZN(n7982) );
  XOR2_X1 U8878 ( .A(n9092), .B(n9093), .Z(n7979) );
  XOR2_X1 U8879 ( .A(n9094), .B(n9095), .Z(n9093) );
  OR2_X1 U8880 ( .A1(n8012), .A2(n8980), .ZN(n7994) );
  XOR2_X1 U8881 ( .A(n9096), .B(n9097), .Z(n7991) );
  XOR2_X1 U8882 ( .A(n9098), .B(n9099), .Z(n9097) );
  OR2_X1 U8883 ( .A1(n8297), .A2(n8980), .ZN(n8006) );
  XOR2_X1 U8884 ( .A(n9100), .B(n9101), .Z(n8003) );
  XOR2_X1 U8885 ( .A(n9102), .B(n9103), .Z(n9101) );
  XOR2_X1 U8886 ( .A(n8882), .B(n8883), .Z(n8139) );
  OR2_X1 U8887 ( .A1(n9104), .A2(n9105), .ZN(n8883) );
  AND2_X1 U8888 ( .A1(n9106), .A2(n9107), .ZN(n9105) );
  AND2_X1 U8889 ( .A1(n9108), .A2(n9109), .ZN(n9104) );
  OR2_X1 U8890 ( .A1(n9106), .A2(n9107), .ZN(n9109) );
  XOR2_X1 U8891 ( .A(n9110), .B(n9111), .Z(n8882) );
  XOR2_X1 U8892 ( .A(n9112), .B(n9113), .Z(n9111) );
  XNOR2_X1 U8893 ( .A(n9108), .B(n9114), .ZN(n8134) );
  XOR2_X1 U8894 ( .A(n9107), .B(n9106), .Z(n9114) );
  OR2_X1 U8895 ( .A1(n7599), .A2(n8297), .ZN(n9106) );
  OR2_X1 U8896 ( .A1(n9115), .A2(n9116), .ZN(n9107) );
  AND2_X1 U8897 ( .A1(n9100), .A2(n9103), .ZN(n9116) );
  AND2_X1 U8898 ( .A1(n9117), .A2(n9102), .ZN(n9115) );
  OR2_X1 U8899 ( .A1(n9118), .A2(n9119), .ZN(n9102) );
  AND2_X1 U8900 ( .A1(n9096), .A2(n9099), .ZN(n9119) );
  AND2_X1 U8901 ( .A1(n9120), .A2(n9098), .ZN(n9118) );
  OR2_X1 U8902 ( .A1(n9121), .A2(n9122), .ZN(n9098) );
  AND2_X1 U8903 ( .A1(n9092), .A2(n9095), .ZN(n9122) );
  AND2_X1 U8904 ( .A1(n9123), .A2(n9094), .ZN(n9121) );
  OR2_X1 U8905 ( .A1(n9124), .A2(n9125), .ZN(n9094) );
  AND2_X1 U8906 ( .A1(n9088), .A2(n9091), .ZN(n9125) );
  AND2_X1 U8907 ( .A1(n9126), .A2(n9090), .ZN(n9124) );
  OR2_X1 U8908 ( .A1(n9127), .A2(n9128), .ZN(n9090) );
  AND2_X1 U8909 ( .A1(n9084), .A2(n9087), .ZN(n9128) );
  AND2_X1 U8910 ( .A1(n9129), .A2(n9086), .ZN(n9127) );
  OR2_X1 U8911 ( .A1(n9130), .A2(n9131), .ZN(n9086) );
  AND2_X1 U8912 ( .A1(n9080), .A2(n9083), .ZN(n9131) );
  AND2_X1 U8913 ( .A1(n9132), .A2(n9082), .ZN(n9130) );
  OR2_X1 U8914 ( .A1(n9133), .A2(n9134), .ZN(n9082) );
  AND2_X1 U8915 ( .A1(n9076), .A2(n9079), .ZN(n9134) );
  AND2_X1 U8916 ( .A1(n9135), .A2(n9078), .ZN(n9133) );
  OR2_X1 U8917 ( .A1(n9136), .A2(n9137), .ZN(n9078) );
  AND2_X1 U8918 ( .A1(n9072), .A2(n9075), .ZN(n9137) );
  AND2_X1 U8919 ( .A1(n9138), .A2(n9074), .ZN(n9136) );
  OR2_X1 U8920 ( .A1(n9139), .A2(n9140), .ZN(n9074) );
  AND2_X1 U8921 ( .A1(n9068), .A2(n9071), .ZN(n9140) );
  AND2_X1 U8922 ( .A1(n9141), .A2(n9070), .ZN(n9139) );
  OR2_X1 U8923 ( .A1(n9142), .A2(n9143), .ZN(n9070) );
  AND2_X1 U8924 ( .A1(n9064), .A2(n9067), .ZN(n9143) );
  AND2_X1 U8925 ( .A1(n9144), .A2(n9066), .ZN(n9142) );
  OR2_X1 U8926 ( .A1(n9145), .A2(n9146), .ZN(n9066) );
  AND2_X1 U8927 ( .A1(n9060), .A2(n9063), .ZN(n9146) );
  AND2_X1 U8928 ( .A1(n9147), .A2(n9062), .ZN(n9145) );
  OR2_X1 U8929 ( .A1(n9148), .A2(n9149), .ZN(n9062) );
  AND2_X1 U8930 ( .A1(n9056), .A2(n9059), .ZN(n9149) );
  AND2_X1 U8931 ( .A1(n9150), .A2(n9058), .ZN(n9148) );
  OR2_X1 U8932 ( .A1(n9151), .A2(n9152), .ZN(n9058) );
  AND2_X1 U8933 ( .A1(n9052), .A2(n9055), .ZN(n9152) );
  AND2_X1 U8934 ( .A1(n9153), .A2(n9054), .ZN(n9151) );
  OR2_X1 U8935 ( .A1(n9154), .A2(n9155), .ZN(n9054) );
  AND2_X1 U8936 ( .A1(n9048), .A2(n9051), .ZN(n9155) );
  AND2_X1 U8937 ( .A1(n9156), .A2(n9050), .ZN(n9154) );
  OR2_X1 U8938 ( .A1(n9157), .A2(n9158), .ZN(n9050) );
  AND2_X1 U8939 ( .A1(n9044), .A2(n9047), .ZN(n9158) );
  AND2_X1 U8940 ( .A1(n9159), .A2(n9046), .ZN(n9157) );
  OR2_X1 U8941 ( .A1(n9160), .A2(n9161), .ZN(n9046) );
  AND2_X1 U8942 ( .A1(n9040), .A2(n9043), .ZN(n9161) );
  AND2_X1 U8943 ( .A1(n9162), .A2(n9042), .ZN(n9160) );
  OR2_X1 U8944 ( .A1(n9163), .A2(n9164), .ZN(n9042) );
  AND2_X1 U8945 ( .A1(n9036), .A2(n9039), .ZN(n9164) );
  AND2_X1 U8946 ( .A1(n9165), .A2(n9038), .ZN(n9163) );
  OR2_X1 U8947 ( .A1(n9166), .A2(n9167), .ZN(n9038) );
  AND2_X1 U8948 ( .A1(n9032), .A2(n9035), .ZN(n9167) );
  AND2_X1 U8949 ( .A1(n9168), .A2(n9034), .ZN(n9166) );
  OR2_X1 U8950 ( .A1(n9169), .A2(n9170), .ZN(n9034) );
  AND2_X1 U8951 ( .A1(n9028), .A2(n9031), .ZN(n9170) );
  AND2_X1 U8952 ( .A1(n9171), .A2(n9030), .ZN(n9169) );
  OR2_X1 U8953 ( .A1(n9172), .A2(n9173), .ZN(n9030) );
  AND2_X1 U8954 ( .A1(n9024), .A2(n9027), .ZN(n9173) );
  AND2_X1 U8955 ( .A1(n9174), .A2(n9026), .ZN(n9172) );
  OR2_X1 U8956 ( .A1(n9175), .A2(n9176), .ZN(n9026) );
  AND2_X1 U8957 ( .A1(n9020), .A2(n9023), .ZN(n9176) );
  AND2_X1 U8958 ( .A1(n9177), .A2(n9022), .ZN(n9175) );
  OR2_X1 U8959 ( .A1(n9178), .A2(n9179), .ZN(n9022) );
  AND2_X1 U8960 ( .A1(n9016), .A2(n9019), .ZN(n9179) );
  AND2_X1 U8961 ( .A1(n9180), .A2(n9018), .ZN(n9178) );
  OR2_X1 U8962 ( .A1(n9181), .A2(n9182), .ZN(n9018) );
  AND2_X1 U8963 ( .A1(n9012), .A2(n9015), .ZN(n9182) );
  AND2_X1 U8964 ( .A1(n9183), .A2(n9014), .ZN(n9181) );
  OR2_X1 U8965 ( .A1(n9184), .A2(n9185), .ZN(n9014) );
  AND2_X1 U8966 ( .A1(n9008), .A2(n9011), .ZN(n9185) );
  AND2_X1 U8967 ( .A1(n9186), .A2(n9010), .ZN(n9184) );
  OR2_X1 U8968 ( .A1(n9187), .A2(n9188), .ZN(n9010) );
  AND2_X1 U8969 ( .A1(n9004), .A2(n9007), .ZN(n9188) );
  AND2_X1 U8970 ( .A1(n9189), .A2(n9006), .ZN(n9187) );
  OR2_X1 U8971 ( .A1(n9190), .A2(n9191), .ZN(n9006) );
  AND2_X1 U8972 ( .A1(n9000), .A2(n9003), .ZN(n9191) );
  AND2_X1 U8973 ( .A1(n9192), .A2(n9002), .ZN(n9190) );
  OR2_X1 U8974 ( .A1(n9193), .A2(n9194), .ZN(n9002) );
  AND2_X1 U8975 ( .A1(n8996), .A2(n8999), .ZN(n9194) );
  AND2_X1 U8976 ( .A1(n9195), .A2(n8998), .ZN(n9193) );
  OR2_X1 U8977 ( .A1(n9196), .A2(n9197), .ZN(n8998) );
  AND2_X1 U8978 ( .A1(n8992), .A2(n8995), .ZN(n9197) );
  AND2_X1 U8979 ( .A1(n9198), .A2(n8994), .ZN(n9196) );
  OR2_X1 U8980 ( .A1(n9199), .A2(n9200), .ZN(n8994) );
  AND2_X1 U8981 ( .A1(n8988), .A2(n8991), .ZN(n9200) );
  AND2_X1 U8982 ( .A1(n9201), .A2(n9202), .ZN(n9199) );
  OR2_X1 U8983 ( .A1(n8991), .A2(n8988), .ZN(n9202) );
  OR2_X1 U8984 ( .A1(n7599), .A2(n8127), .ZN(n8988) );
  OR3_X1 U8985 ( .A1(n8981), .A2(n7599), .A3(n7611), .ZN(n8991) );
  INV_X1 U8986 ( .A(n8990), .ZN(n9201) );
  OR2_X1 U8987 ( .A1(n9203), .A2(n9204), .ZN(n8990) );
  AND2_X1 U8988 ( .A1(b_29_), .A2(n9205), .ZN(n9204) );
  OR2_X1 U8989 ( .A1(n9206), .A2(n7598), .ZN(n9205) );
  AND2_X1 U8990 ( .A1(a_30_), .A2(n8125), .ZN(n9206) );
  AND2_X1 U8991 ( .A1(b_28_), .A2(n9207), .ZN(n9203) );
  OR2_X1 U8992 ( .A1(n9208), .A2(n7601), .ZN(n9207) );
  AND2_X1 U8993 ( .A1(a_31_), .A2(n7611), .ZN(n9208) );
  OR2_X1 U8994 ( .A1(n8995), .A2(n8992), .ZN(n9198) );
  XNOR2_X1 U8995 ( .A(n7616), .B(n9209), .ZN(n8992) );
  XOR2_X1 U8996 ( .A(n9210), .B(n9211), .Z(n9209) );
  OR2_X1 U8997 ( .A1(n7599), .A2(n8124), .ZN(n8995) );
  OR2_X1 U8998 ( .A1(n8999), .A2(n8996), .ZN(n9195) );
  XOR2_X1 U8999 ( .A(n9212), .B(n9213), .Z(n8996) );
  XOR2_X1 U9000 ( .A(n9214), .B(n9215), .Z(n9213) );
  OR2_X1 U9001 ( .A1(n7599), .A2(n8121), .ZN(n8999) );
  OR2_X1 U9002 ( .A1(n9003), .A2(n9000), .ZN(n9192) );
  XOR2_X1 U9003 ( .A(n9216), .B(n9217), .Z(n9000) );
  XOR2_X1 U9004 ( .A(n9218), .B(n9219), .Z(n9217) );
  OR2_X1 U9005 ( .A1(n7599), .A2(n8118), .ZN(n9003) );
  OR2_X1 U9006 ( .A1(n9007), .A2(n9004), .ZN(n9189) );
  XOR2_X1 U9007 ( .A(n9220), .B(n9221), .Z(n9004) );
  XOR2_X1 U9008 ( .A(n9222), .B(n9223), .Z(n9221) );
  OR2_X1 U9009 ( .A1(n7599), .A2(n8115), .ZN(n9007) );
  OR2_X1 U9010 ( .A1(n9011), .A2(n9008), .ZN(n9186) );
  XOR2_X1 U9011 ( .A(n9224), .B(n9225), .Z(n9008) );
  XOR2_X1 U9012 ( .A(n9226), .B(n9227), .Z(n9225) );
  OR2_X1 U9013 ( .A1(n7599), .A2(n8112), .ZN(n9011) );
  OR2_X1 U9014 ( .A1(n9015), .A2(n9012), .ZN(n9183) );
  XOR2_X1 U9015 ( .A(n9228), .B(n9229), .Z(n9012) );
  XOR2_X1 U9016 ( .A(n9230), .B(n9231), .Z(n9229) );
  OR2_X1 U9017 ( .A1(n7599), .A2(n8109), .ZN(n9015) );
  OR2_X1 U9018 ( .A1(n9019), .A2(n9016), .ZN(n9180) );
  XOR2_X1 U9019 ( .A(n9232), .B(n9233), .Z(n9016) );
  XOR2_X1 U9020 ( .A(n9234), .B(n9235), .Z(n9233) );
  OR2_X1 U9021 ( .A1(n7599), .A2(n8106), .ZN(n9019) );
  OR2_X1 U9022 ( .A1(n9023), .A2(n9020), .ZN(n9177) );
  XOR2_X1 U9023 ( .A(n9236), .B(n9237), .Z(n9020) );
  XOR2_X1 U9024 ( .A(n9238), .B(n9239), .Z(n9237) );
  OR2_X1 U9025 ( .A1(n8102), .A2(n7599), .ZN(n9023) );
  OR2_X1 U9026 ( .A1(n9027), .A2(n9024), .ZN(n9174) );
  XOR2_X1 U9027 ( .A(n9240), .B(n9241), .Z(n9024) );
  XOR2_X1 U9028 ( .A(n9242), .B(n9243), .Z(n9241) );
  OR2_X1 U9029 ( .A1(n7599), .A2(n8097), .ZN(n9027) );
  OR2_X1 U9030 ( .A1(n9031), .A2(n9028), .ZN(n9171) );
  XOR2_X1 U9031 ( .A(n9244), .B(n9245), .Z(n9028) );
  XOR2_X1 U9032 ( .A(n9246), .B(n9247), .Z(n9245) );
  OR2_X1 U9033 ( .A1(n8093), .A2(n7599), .ZN(n9031) );
  OR2_X1 U9034 ( .A1(n9035), .A2(n9032), .ZN(n9168) );
  XOR2_X1 U9035 ( .A(n9248), .B(n9249), .Z(n9032) );
  XOR2_X1 U9036 ( .A(n9250), .B(n9251), .Z(n9249) );
  OR2_X1 U9037 ( .A1(n7599), .A2(n8088), .ZN(n9035) );
  OR2_X1 U9038 ( .A1(n9039), .A2(n9036), .ZN(n9165) );
  XOR2_X1 U9039 ( .A(n9252), .B(n9253), .Z(n9036) );
  XOR2_X1 U9040 ( .A(n9254), .B(n9255), .Z(n9253) );
  OR2_X1 U9041 ( .A1(n8084), .A2(n7599), .ZN(n9039) );
  OR2_X1 U9042 ( .A1(n9043), .A2(n9040), .ZN(n9162) );
  XOR2_X1 U9043 ( .A(n9256), .B(n9257), .Z(n9040) );
  XOR2_X1 U9044 ( .A(n9258), .B(n9259), .Z(n9257) );
  OR2_X1 U9045 ( .A1(n7599), .A2(n8079), .ZN(n9043) );
  OR2_X1 U9046 ( .A1(n9047), .A2(n9044), .ZN(n9159) );
  XOR2_X1 U9047 ( .A(n9260), .B(n9261), .Z(n9044) );
  XOR2_X1 U9048 ( .A(n9262), .B(n9263), .Z(n9261) );
  OR2_X1 U9049 ( .A1(n8075), .A2(n7599), .ZN(n9047) );
  OR2_X1 U9050 ( .A1(n9051), .A2(n9048), .ZN(n9156) );
  XOR2_X1 U9051 ( .A(n9264), .B(n9265), .Z(n9048) );
  XOR2_X1 U9052 ( .A(n9266), .B(n9267), .Z(n9265) );
  OR2_X1 U9053 ( .A1(n7599), .A2(n8070), .ZN(n9051) );
  OR2_X1 U9054 ( .A1(n9055), .A2(n9052), .ZN(n9153) );
  XOR2_X1 U9055 ( .A(n9268), .B(n9269), .Z(n9052) );
  XOR2_X1 U9056 ( .A(n9270), .B(n9271), .Z(n9269) );
  OR2_X1 U9057 ( .A1(n8066), .A2(n7599), .ZN(n9055) );
  OR2_X1 U9058 ( .A1(n9059), .A2(n9056), .ZN(n9150) );
  XOR2_X1 U9059 ( .A(n9272), .B(n9273), .Z(n9056) );
  XOR2_X1 U9060 ( .A(n9274), .B(n9275), .Z(n9273) );
  OR2_X1 U9061 ( .A1(n7599), .A2(n8061), .ZN(n9059) );
  OR2_X1 U9062 ( .A1(n9063), .A2(n9060), .ZN(n9147) );
  XOR2_X1 U9063 ( .A(n9276), .B(n9277), .Z(n9060) );
  XOR2_X1 U9064 ( .A(n9278), .B(n9279), .Z(n9277) );
  OR2_X1 U9065 ( .A1(n8057), .A2(n7599), .ZN(n9063) );
  OR2_X1 U9066 ( .A1(n9067), .A2(n9064), .ZN(n9144) );
  XOR2_X1 U9067 ( .A(n9280), .B(n9281), .Z(n9064) );
  XOR2_X1 U9068 ( .A(n9282), .B(n9283), .Z(n9281) );
  OR2_X1 U9069 ( .A1(n7599), .A2(n8052), .ZN(n9067) );
  OR2_X1 U9070 ( .A1(n9071), .A2(n9068), .ZN(n9141) );
  XOR2_X1 U9071 ( .A(n9284), .B(n9285), .Z(n9068) );
  XOR2_X1 U9072 ( .A(n9286), .B(n9287), .Z(n9285) );
  OR2_X1 U9073 ( .A1(n8048), .A2(n7599), .ZN(n9071) );
  OR2_X1 U9074 ( .A1(n9075), .A2(n9072), .ZN(n9138) );
  XOR2_X1 U9075 ( .A(n9288), .B(n9289), .Z(n9072) );
  XOR2_X1 U9076 ( .A(n9290), .B(n9291), .Z(n9289) );
  OR2_X1 U9077 ( .A1(n7599), .A2(n8043), .ZN(n9075) );
  OR2_X1 U9078 ( .A1(n9079), .A2(n9076), .ZN(n9135) );
  XOR2_X1 U9079 ( .A(n9292), .B(n9293), .Z(n9076) );
  XOR2_X1 U9080 ( .A(n9294), .B(n9295), .Z(n9293) );
  OR2_X1 U9081 ( .A1(n8039), .A2(n7599), .ZN(n9079) );
  OR2_X1 U9082 ( .A1(n9083), .A2(n9080), .ZN(n9132) );
  XOR2_X1 U9083 ( .A(n9296), .B(n9297), .Z(n9080) );
  XOR2_X1 U9084 ( .A(n9298), .B(n9299), .Z(n9297) );
  OR2_X1 U9085 ( .A1(n7599), .A2(n8034), .ZN(n9083) );
  OR2_X1 U9086 ( .A1(n9087), .A2(n9084), .ZN(n9129) );
  XOR2_X1 U9087 ( .A(n9300), .B(n9301), .Z(n9084) );
  XOR2_X1 U9088 ( .A(n9302), .B(n9303), .Z(n9301) );
  OR2_X1 U9089 ( .A1(n8030), .A2(n7599), .ZN(n9087) );
  OR2_X1 U9090 ( .A1(n9091), .A2(n9088), .ZN(n9126) );
  XOR2_X1 U9091 ( .A(n9304), .B(n9305), .Z(n9088) );
  XOR2_X1 U9092 ( .A(n9306), .B(n9307), .Z(n9305) );
  OR2_X1 U9093 ( .A1(n7599), .A2(n8025), .ZN(n9091) );
  OR2_X1 U9094 ( .A1(n9095), .A2(n9092), .ZN(n9123) );
  XOR2_X1 U9095 ( .A(n9308), .B(n9309), .Z(n9092) );
  XOR2_X1 U9096 ( .A(n9310), .B(n9311), .Z(n9309) );
  OR2_X1 U9097 ( .A1(n8021), .A2(n7599), .ZN(n9095) );
  OR2_X1 U9098 ( .A1(n9099), .A2(n9096), .ZN(n9120) );
  XOR2_X1 U9099 ( .A(n9312), .B(n9313), .Z(n9096) );
  XOR2_X1 U9100 ( .A(n9314), .B(n9315), .Z(n9313) );
  OR2_X1 U9101 ( .A1(n7599), .A2(n8016), .ZN(n9099) );
  OR2_X1 U9102 ( .A1(n9103), .A2(n9100), .ZN(n9117) );
  XNOR2_X1 U9103 ( .A(n9316), .B(n9317), .ZN(n9100) );
  XNOR2_X1 U9104 ( .A(n9318), .B(n9319), .ZN(n9316) );
  OR2_X1 U9105 ( .A1(n7599), .A2(n8012), .ZN(n9103) );
  INV_X1 U9106 ( .A(b_30_), .ZN(n7599) );
  XOR2_X1 U9107 ( .A(n9320), .B(n9321), .Z(n9108) );
  XOR2_X1 U9108 ( .A(n9322), .B(n9323), .Z(n9321) );
  OR2_X1 U9109 ( .A1(n9324), .A2(n8877), .ZN(n8150) );
  XOR2_X1 U9110 ( .A(n8872), .B(n8873), .Z(n8877) );
  AND2_X1 U9111 ( .A1(n8878), .A2(n8876), .ZN(n9324) );
  XNOR2_X1 U9112 ( .A(n9325), .B(n9326), .ZN(n8876) );
  XOR2_X1 U9113 ( .A(n9327), .B(n9328), .Z(n9326) );
  INV_X1 U9114 ( .A(n8884), .ZN(n8878) );
  OR2_X1 U9115 ( .A1(n9329), .A2(n9330), .ZN(n8884) );
  AND2_X1 U9116 ( .A1(n9113), .A2(n9112), .ZN(n9330) );
  AND2_X1 U9117 ( .A1(n9110), .A2(n9331), .ZN(n9329) );
  OR2_X1 U9118 ( .A1(n9112), .A2(n9113), .ZN(n9331) );
  OR2_X1 U9119 ( .A1(n7611), .A2(n8297), .ZN(n9113) );
  OR2_X1 U9120 ( .A1(n9332), .A2(n9333), .ZN(n9112) );
  AND2_X1 U9121 ( .A1(n9323), .A2(n9322), .ZN(n9333) );
  AND2_X1 U9122 ( .A1(n9320), .A2(n9334), .ZN(n9332) );
  OR2_X1 U9123 ( .A1(n9322), .A2(n9323), .ZN(n9334) );
  OR2_X1 U9124 ( .A1(n7611), .A2(n8012), .ZN(n9323) );
  OR2_X1 U9125 ( .A1(n9335), .A2(n9336), .ZN(n9322) );
  AND2_X1 U9126 ( .A1(n9319), .A2(n9318), .ZN(n9336) );
  AND2_X1 U9127 ( .A1(n9317), .A2(n9337), .ZN(n9335) );
  OR2_X1 U9128 ( .A1(n9318), .A2(n9319), .ZN(n9337) );
  OR2_X1 U9129 ( .A1(n9338), .A2(n9339), .ZN(n9319) );
  AND2_X1 U9130 ( .A1(n9315), .A2(n9314), .ZN(n9339) );
  AND2_X1 U9131 ( .A1(n9312), .A2(n9340), .ZN(n9338) );
  OR2_X1 U9132 ( .A1(n9314), .A2(n9315), .ZN(n9340) );
  OR2_X1 U9133 ( .A1(n8021), .A2(n7611), .ZN(n9315) );
  OR2_X1 U9134 ( .A1(n9341), .A2(n9342), .ZN(n9314) );
  AND2_X1 U9135 ( .A1(n9311), .A2(n9310), .ZN(n9342) );
  AND2_X1 U9136 ( .A1(n9308), .A2(n9343), .ZN(n9341) );
  OR2_X1 U9137 ( .A1(n9310), .A2(n9311), .ZN(n9343) );
  OR2_X1 U9138 ( .A1(n7611), .A2(n8025), .ZN(n9311) );
  OR2_X1 U9139 ( .A1(n9344), .A2(n9345), .ZN(n9310) );
  AND2_X1 U9140 ( .A1(n9307), .A2(n9306), .ZN(n9345) );
  AND2_X1 U9141 ( .A1(n9304), .A2(n9346), .ZN(n9344) );
  OR2_X1 U9142 ( .A1(n9306), .A2(n9307), .ZN(n9346) );
  OR2_X1 U9143 ( .A1(n8030), .A2(n7611), .ZN(n9307) );
  OR2_X1 U9144 ( .A1(n9347), .A2(n9348), .ZN(n9306) );
  AND2_X1 U9145 ( .A1(n9303), .A2(n9302), .ZN(n9348) );
  AND2_X1 U9146 ( .A1(n9300), .A2(n9349), .ZN(n9347) );
  OR2_X1 U9147 ( .A1(n9302), .A2(n9303), .ZN(n9349) );
  OR2_X1 U9148 ( .A1(n7611), .A2(n8034), .ZN(n9303) );
  OR2_X1 U9149 ( .A1(n9350), .A2(n9351), .ZN(n9302) );
  AND2_X1 U9150 ( .A1(n9299), .A2(n9298), .ZN(n9351) );
  AND2_X1 U9151 ( .A1(n9296), .A2(n9352), .ZN(n9350) );
  OR2_X1 U9152 ( .A1(n9298), .A2(n9299), .ZN(n9352) );
  OR2_X1 U9153 ( .A1(n8039), .A2(n7611), .ZN(n9299) );
  OR2_X1 U9154 ( .A1(n9353), .A2(n9354), .ZN(n9298) );
  AND2_X1 U9155 ( .A1(n9295), .A2(n9294), .ZN(n9354) );
  AND2_X1 U9156 ( .A1(n9292), .A2(n9355), .ZN(n9353) );
  OR2_X1 U9157 ( .A1(n9294), .A2(n9295), .ZN(n9355) );
  OR2_X1 U9158 ( .A1(n7611), .A2(n8043), .ZN(n9295) );
  OR2_X1 U9159 ( .A1(n9356), .A2(n9357), .ZN(n9294) );
  AND2_X1 U9160 ( .A1(n9291), .A2(n9290), .ZN(n9357) );
  AND2_X1 U9161 ( .A1(n9288), .A2(n9358), .ZN(n9356) );
  OR2_X1 U9162 ( .A1(n9290), .A2(n9291), .ZN(n9358) );
  OR2_X1 U9163 ( .A1(n8048), .A2(n7611), .ZN(n9291) );
  OR2_X1 U9164 ( .A1(n9359), .A2(n9360), .ZN(n9290) );
  AND2_X1 U9165 ( .A1(n9287), .A2(n9286), .ZN(n9360) );
  AND2_X1 U9166 ( .A1(n9284), .A2(n9361), .ZN(n9359) );
  OR2_X1 U9167 ( .A1(n9286), .A2(n9287), .ZN(n9361) );
  OR2_X1 U9168 ( .A1(n7611), .A2(n8052), .ZN(n9287) );
  OR2_X1 U9169 ( .A1(n9362), .A2(n9363), .ZN(n9286) );
  AND2_X1 U9170 ( .A1(n9283), .A2(n9282), .ZN(n9363) );
  AND2_X1 U9171 ( .A1(n9280), .A2(n9364), .ZN(n9362) );
  OR2_X1 U9172 ( .A1(n9282), .A2(n9283), .ZN(n9364) );
  OR2_X1 U9173 ( .A1(n8057), .A2(n7611), .ZN(n9283) );
  OR2_X1 U9174 ( .A1(n9365), .A2(n9366), .ZN(n9282) );
  AND2_X1 U9175 ( .A1(n9279), .A2(n9278), .ZN(n9366) );
  AND2_X1 U9176 ( .A1(n9276), .A2(n9367), .ZN(n9365) );
  OR2_X1 U9177 ( .A1(n9278), .A2(n9279), .ZN(n9367) );
  OR2_X1 U9178 ( .A1(n7611), .A2(n8061), .ZN(n9279) );
  OR2_X1 U9179 ( .A1(n9368), .A2(n9369), .ZN(n9278) );
  AND2_X1 U9180 ( .A1(n9275), .A2(n9274), .ZN(n9369) );
  AND2_X1 U9181 ( .A1(n9272), .A2(n9370), .ZN(n9368) );
  OR2_X1 U9182 ( .A1(n9274), .A2(n9275), .ZN(n9370) );
  OR2_X1 U9183 ( .A1(n8066), .A2(n7611), .ZN(n9275) );
  OR2_X1 U9184 ( .A1(n9371), .A2(n9372), .ZN(n9274) );
  AND2_X1 U9185 ( .A1(n9271), .A2(n9270), .ZN(n9372) );
  AND2_X1 U9186 ( .A1(n9268), .A2(n9373), .ZN(n9371) );
  OR2_X1 U9187 ( .A1(n9270), .A2(n9271), .ZN(n9373) );
  OR2_X1 U9188 ( .A1(n7611), .A2(n8070), .ZN(n9271) );
  OR2_X1 U9189 ( .A1(n9374), .A2(n9375), .ZN(n9270) );
  AND2_X1 U9190 ( .A1(n9267), .A2(n9266), .ZN(n9375) );
  AND2_X1 U9191 ( .A1(n9264), .A2(n9376), .ZN(n9374) );
  OR2_X1 U9192 ( .A1(n9266), .A2(n9267), .ZN(n9376) );
  OR2_X1 U9193 ( .A1(n8075), .A2(n7611), .ZN(n9267) );
  OR2_X1 U9194 ( .A1(n9377), .A2(n9378), .ZN(n9266) );
  AND2_X1 U9195 ( .A1(n9263), .A2(n9262), .ZN(n9378) );
  AND2_X1 U9196 ( .A1(n9260), .A2(n9379), .ZN(n9377) );
  OR2_X1 U9197 ( .A1(n9262), .A2(n9263), .ZN(n9379) );
  OR2_X1 U9198 ( .A1(n7611), .A2(n8079), .ZN(n9263) );
  OR2_X1 U9199 ( .A1(n9380), .A2(n9381), .ZN(n9262) );
  AND2_X1 U9200 ( .A1(n9259), .A2(n9258), .ZN(n9381) );
  AND2_X1 U9201 ( .A1(n9256), .A2(n9382), .ZN(n9380) );
  OR2_X1 U9202 ( .A1(n9258), .A2(n9259), .ZN(n9382) );
  OR2_X1 U9203 ( .A1(n8084), .A2(n7611), .ZN(n9259) );
  OR2_X1 U9204 ( .A1(n9383), .A2(n9384), .ZN(n9258) );
  AND2_X1 U9205 ( .A1(n9255), .A2(n9254), .ZN(n9384) );
  AND2_X1 U9206 ( .A1(n9252), .A2(n9385), .ZN(n9383) );
  OR2_X1 U9207 ( .A1(n9254), .A2(n9255), .ZN(n9385) );
  OR2_X1 U9208 ( .A1(n7611), .A2(n8088), .ZN(n9255) );
  OR2_X1 U9209 ( .A1(n9386), .A2(n9387), .ZN(n9254) );
  AND2_X1 U9210 ( .A1(n9251), .A2(n9250), .ZN(n9387) );
  AND2_X1 U9211 ( .A1(n9248), .A2(n9388), .ZN(n9386) );
  OR2_X1 U9212 ( .A1(n9250), .A2(n9251), .ZN(n9388) );
  OR2_X1 U9213 ( .A1(n8093), .A2(n7611), .ZN(n9251) );
  OR2_X1 U9214 ( .A1(n9389), .A2(n9390), .ZN(n9250) );
  AND2_X1 U9215 ( .A1(n9247), .A2(n9246), .ZN(n9390) );
  AND2_X1 U9216 ( .A1(n9244), .A2(n9391), .ZN(n9389) );
  OR2_X1 U9217 ( .A1(n9246), .A2(n9247), .ZN(n9391) );
  OR2_X1 U9218 ( .A1(n7611), .A2(n8097), .ZN(n9247) );
  OR2_X1 U9219 ( .A1(n9392), .A2(n9393), .ZN(n9246) );
  AND2_X1 U9220 ( .A1(n9243), .A2(n9242), .ZN(n9393) );
  AND2_X1 U9221 ( .A1(n9240), .A2(n9394), .ZN(n9392) );
  OR2_X1 U9222 ( .A1(n9242), .A2(n9243), .ZN(n9394) );
  OR2_X1 U9223 ( .A1(n8102), .A2(n7611), .ZN(n9243) );
  OR2_X1 U9224 ( .A1(n9395), .A2(n9396), .ZN(n9242) );
  AND2_X1 U9225 ( .A1(n9239), .A2(n9238), .ZN(n9396) );
  AND2_X1 U9226 ( .A1(n9236), .A2(n9397), .ZN(n9395) );
  OR2_X1 U9227 ( .A1(n9238), .A2(n9239), .ZN(n9397) );
  OR2_X1 U9228 ( .A1(n7611), .A2(n8106), .ZN(n9239) );
  OR2_X1 U9229 ( .A1(n9398), .A2(n9399), .ZN(n9238) );
  AND2_X1 U9230 ( .A1(n9235), .A2(n9234), .ZN(n9399) );
  AND2_X1 U9231 ( .A1(n9232), .A2(n9400), .ZN(n9398) );
  OR2_X1 U9232 ( .A1(n9234), .A2(n9235), .ZN(n9400) );
  OR2_X1 U9233 ( .A1(n7611), .A2(n8109), .ZN(n9235) );
  OR2_X1 U9234 ( .A1(n9401), .A2(n9402), .ZN(n9234) );
  AND2_X1 U9235 ( .A1(n9231), .A2(n9230), .ZN(n9402) );
  AND2_X1 U9236 ( .A1(n9228), .A2(n9403), .ZN(n9401) );
  OR2_X1 U9237 ( .A1(n9230), .A2(n9231), .ZN(n9403) );
  OR2_X1 U9238 ( .A1(n7611), .A2(n8112), .ZN(n9231) );
  OR2_X1 U9239 ( .A1(n9404), .A2(n9405), .ZN(n9230) );
  AND2_X1 U9240 ( .A1(n9227), .A2(n9226), .ZN(n9405) );
  AND2_X1 U9241 ( .A1(n9224), .A2(n9406), .ZN(n9404) );
  OR2_X1 U9242 ( .A1(n9226), .A2(n9227), .ZN(n9406) );
  OR2_X1 U9243 ( .A1(n7611), .A2(n8115), .ZN(n9227) );
  OR2_X1 U9244 ( .A1(n9407), .A2(n9408), .ZN(n9226) );
  AND2_X1 U9245 ( .A1(n9223), .A2(n9222), .ZN(n9408) );
  AND2_X1 U9246 ( .A1(n9220), .A2(n9409), .ZN(n9407) );
  OR2_X1 U9247 ( .A1(n9222), .A2(n9223), .ZN(n9409) );
  OR2_X1 U9248 ( .A1(n7611), .A2(n8118), .ZN(n9223) );
  OR2_X1 U9249 ( .A1(n9410), .A2(n9411), .ZN(n9222) );
  AND2_X1 U9250 ( .A1(n9219), .A2(n9218), .ZN(n9411) );
  AND2_X1 U9251 ( .A1(n9216), .A2(n9412), .ZN(n9410) );
  OR2_X1 U9252 ( .A1(n9218), .A2(n9219), .ZN(n9412) );
  OR2_X1 U9253 ( .A1(n7611), .A2(n8121), .ZN(n9219) );
  OR2_X1 U9254 ( .A1(n9413), .A2(n9414), .ZN(n9218) );
  AND2_X1 U9255 ( .A1(n9215), .A2(n9214), .ZN(n9414) );
  AND2_X1 U9256 ( .A1(n9212), .A2(n9415), .ZN(n9413) );
  OR2_X1 U9257 ( .A1(n9214), .A2(n9215), .ZN(n9415) );
  OR2_X1 U9258 ( .A1(n7611), .A2(n8124), .ZN(n9215) );
  OR2_X1 U9259 ( .A1(n9416), .A2(n9417), .ZN(n9214) );
  AND2_X1 U9260 ( .A1(n7616), .A2(n9211), .ZN(n9417) );
  AND2_X1 U9261 ( .A1(n9418), .A2(n9419), .ZN(n9416) );
  OR2_X1 U9262 ( .A1(n9211), .A2(n7616), .ZN(n9419) );
  OR2_X1 U9263 ( .A1(n7611), .A2(n8127), .ZN(n7616) );
  OR3_X1 U9264 ( .A1(n8981), .A2(n7611), .A3(n8125), .ZN(n9211) );
  INV_X1 U9265 ( .A(n9210), .ZN(n9418) );
  OR2_X1 U9266 ( .A1(n9420), .A2(n9421), .ZN(n9210) );
  AND2_X1 U9267 ( .A1(b_28_), .A2(n9422), .ZN(n9421) );
  OR2_X1 U9268 ( .A1(n9423), .A2(n7598), .ZN(n9422) );
  AND2_X1 U9269 ( .A1(a_30_), .A2(n8122), .ZN(n9423) );
  AND2_X1 U9270 ( .A1(b_27_), .A2(n9424), .ZN(n9420) );
  OR2_X1 U9271 ( .A1(n9425), .A2(n7601), .ZN(n9424) );
  AND2_X1 U9272 ( .A1(a_31_), .A2(n8125), .ZN(n9425) );
  XNOR2_X1 U9273 ( .A(n9426), .B(n9427), .ZN(n9212) );
  XOR2_X1 U9274 ( .A(n9428), .B(n9429), .Z(n9427) );
  XOR2_X1 U9275 ( .A(n9430), .B(n9431), .Z(n9216) );
  XOR2_X1 U9276 ( .A(n9432), .B(n7634), .Z(n9431) );
  XOR2_X1 U9277 ( .A(n9433), .B(n9434), .Z(n9220) );
  XOR2_X1 U9278 ( .A(n9435), .B(n9436), .Z(n9434) );
  XOR2_X1 U9279 ( .A(n9437), .B(n9438), .Z(n9224) );
  XOR2_X1 U9280 ( .A(n9439), .B(n9440), .Z(n9438) );
  XOR2_X1 U9281 ( .A(n9441), .B(n9442), .Z(n9228) );
  XOR2_X1 U9282 ( .A(n9443), .B(n9444), .Z(n9442) );
  XOR2_X1 U9283 ( .A(n9445), .B(n9446), .Z(n9232) );
  XOR2_X1 U9284 ( .A(n9447), .B(n9448), .Z(n9446) );
  XOR2_X1 U9285 ( .A(n9449), .B(n9450), .Z(n9236) );
  XOR2_X1 U9286 ( .A(n9451), .B(n9452), .Z(n9450) );
  XOR2_X1 U9287 ( .A(n9453), .B(n9454), .Z(n9240) );
  XOR2_X1 U9288 ( .A(n9455), .B(n9456), .Z(n9454) );
  XOR2_X1 U9289 ( .A(n9457), .B(n9458), .Z(n9244) );
  XOR2_X1 U9290 ( .A(n9459), .B(n9460), .Z(n9458) );
  XOR2_X1 U9291 ( .A(n9461), .B(n9462), .Z(n9248) );
  XOR2_X1 U9292 ( .A(n9463), .B(n9464), .Z(n9462) );
  XOR2_X1 U9293 ( .A(n9465), .B(n9466), .Z(n9252) );
  XOR2_X1 U9294 ( .A(n9467), .B(n9468), .Z(n9466) );
  XOR2_X1 U9295 ( .A(n9469), .B(n9470), .Z(n9256) );
  XOR2_X1 U9296 ( .A(n9471), .B(n9472), .Z(n9470) );
  XOR2_X1 U9297 ( .A(n9473), .B(n9474), .Z(n9260) );
  XOR2_X1 U9298 ( .A(n9475), .B(n9476), .Z(n9474) );
  XOR2_X1 U9299 ( .A(n9477), .B(n9478), .Z(n9264) );
  XOR2_X1 U9300 ( .A(n9479), .B(n9480), .Z(n9478) );
  XOR2_X1 U9301 ( .A(n9481), .B(n9482), .Z(n9268) );
  XOR2_X1 U9302 ( .A(n9483), .B(n9484), .Z(n9482) );
  XOR2_X1 U9303 ( .A(n9485), .B(n9486), .Z(n9272) );
  XOR2_X1 U9304 ( .A(n9487), .B(n9488), .Z(n9486) );
  XOR2_X1 U9305 ( .A(n9489), .B(n9490), .Z(n9276) );
  XOR2_X1 U9306 ( .A(n9491), .B(n9492), .Z(n9490) );
  XOR2_X1 U9307 ( .A(n9493), .B(n9494), .Z(n9280) );
  XOR2_X1 U9308 ( .A(n9495), .B(n9496), .Z(n9494) );
  XOR2_X1 U9309 ( .A(n9497), .B(n9498), .Z(n9284) );
  XOR2_X1 U9310 ( .A(n9499), .B(n9500), .Z(n9498) );
  XOR2_X1 U9311 ( .A(n9501), .B(n9502), .Z(n9288) );
  XOR2_X1 U9312 ( .A(n9503), .B(n9504), .Z(n9502) );
  XOR2_X1 U9313 ( .A(n9505), .B(n9506), .Z(n9292) );
  XOR2_X1 U9314 ( .A(n9507), .B(n9508), .Z(n9506) );
  XOR2_X1 U9315 ( .A(n9509), .B(n9510), .Z(n9296) );
  XOR2_X1 U9316 ( .A(n9511), .B(n9512), .Z(n9510) );
  XOR2_X1 U9317 ( .A(n9513), .B(n9514), .Z(n9300) );
  XOR2_X1 U9318 ( .A(n9515), .B(n9516), .Z(n9514) );
  XOR2_X1 U9319 ( .A(n9517), .B(n9518), .Z(n9304) );
  XOR2_X1 U9320 ( .A(n9519), .B(n9520), .Z(n9518) );
  XOR2_X1 U9321 ( .A(n9521), .B(n9522), .Z(n9308) );
  XOR2_X1 U9322 ( .A(n9523), .B(n9524), .Z(n9522) );
  XOR2_X1 U9323 ( .A(n9525), .B(n9526), .Z(n9312) );
  XOR2_X1 U9324 ( .A(n9527), .B(n9528), .Z(n9526) );
  OR2_X1 U9325 ( .A1(n7611), .A2(n8016), .ZN(n9318) );
  XOR2_X1 U9326 ( .A(n9529), .B(n9530), .Z(n9317) );
  XOR2_X1 U9327 ( .A(n9531), .B(n9532), .Z(n9530) );
  XNOR2_X1 U9328 ( .A(n9533), .B(n9534), .ZN(n9320) );
  XNOR2_X1 U9329 ( .A(n9535), .B(n9536), .ZN(n9533) );
  XOR2_X1 U9330 ( .A(n9537), .B(n9538), .Z(n9110) );
  XOR2_X1 U9331 ( .A(n9539), .B(n9540), .Z(n9538) );
  OR2_X1 U9332 ( .A1(n9541), .A2(n8874), .ZN(n8156) );
  AND2_X1 U9333 ( .A1(n9542), .A2(n9543), .ZN(n8874) );
  INV_X1 U9334 ( .A(n9544), .ZN(n9542) );
  AND2_X1 U9335 ( .A1(n9545), .A2(n9546), .ZN(n9544) );
  AND2_X1 U9336 ( .A1(n8873), .A2(n8872), .ZN(n9541) );
  XNOR2_X1 U9337 ( .A(n9547), .B(n9548), .ZN(n8872) );
  XOR2_X1 U9338 ( .A(n9549), .B(n9550), .Z(n9548) );
  INV_X1 U9339 ( .A(n9551), .ZN(n8873) );
  OR2_X1 U9340 ( .A1(n9552), .A2(n9553), .ZN(n9551) );
  AND2_X1 U9341 ( .A1(n9328), .A2(n9327), .ZN(n9553) );
  AND2_X1 U9342 ( .A1(n9325), .A2(n9554), .ZN(n9552) );
  OR2_X1 U9343 ( .A1(n9327), .A2(n9328), .ZN(n9554) );
  OR2_X1 U9344 ( .A1(n8125), .A2(n8297), .ZN(n9328) );
  OR2_X1 U9345 ( .A1(n9555), .A2(n9556), .ZN(n9327) );
  AND2_X1 U9346 ( .A1(n9540), .A2(n9539), .ZN(n9556) );
  AND2_X1 U9347 ( .A1(n9537), .A2(n9557), .ZN(n9555) );
  OR2_X1 U9348 ( .A1(n9539), .A2(n9540), .ZN(n9557) );
  OR2_X1 U9349 ( .A1(n8125), .A2(n8012), .ZN(n9540) );
  OR2_X1 U9350 ( .A1(n9558), .A2(n9559), .ZN(n9539) );
  AND2_X1 U9351 ( .A1(n9536), .A2(n9535), .ZN(n9559) );
  AND2_X1 U9352 ( .A1(n9534), .A2(n9560), .ZN(n9558) );
  OR2_X1 U9353 ( .A1(n9535), .A2(n9536), .ZN(n9560) );
  OR2_X1 U9354 ( .A1(n9561), .A2(n9562), .ZN(n9536) );
  AND2_X1 U9355 ( .A1(n9532), .A2(n9531), .ZN(n9562) );
  AND2_X1 U9356 ( .A1(n9529), .A2(n9563), .ZN(n9561) );
  OR2_X1 U9357 ( .A1(n9531), .A2(n9532), .ZN(n9563) );
  OR2_X1 U9358 ( .A1(n8021), .A2(n8125), .ZN(n9532) );
  OR2_X1 U9359 ( .A1(n9564), .A2(n9565), .ZN(n9531) );
  AND2_X1 U9360 ( .A1(n9528), .A2(n9527), .ZN(n9565) );
  AND2_X1 U9361 ( .A1(n9525), .A2(n9566), .ZN(n9564) );
  OR2_X1 U9362 ( .A1(n9527), .A2(n9528), .ZN(n9566) );
  OR2_X1 U9363 ( .A1(n8125), .A2(n8025), .ZN(n9528) );
  OR2_X1 U9364 ( .A1(n9567), .A2(n9568), .ZN(n9527) );
  AND2_X1 U9365 ( .A1(n9524), .A2(n9523), .ZN(n9568) );
  AND2_X1 U9366 ( .A1(n9521), .A2(n9569), .ZN(n9567) );
  OR2_X1 U9367 ( .A1(n9523), .A2(n9524), .ZN(n9569) );
  OR2_X1 U9368 ( .A1(n8030), .A2(n8125), .ZN(n9524) );
  OR2_X1 U9369 ( .A1(n9570), .A2(n9571), .ZN(n9523) );
  AND2_X1 U9370 ( .A1(n9520), .A2(n9519), .ZN(n9571) );
  AND2_X1 U9371 ( .A1(n9517), .A2(n9572), .ZN(n9570) );
  OR2_X1 U9372 ( .A1(n9519), .A2(n9520), .ZN(n9572) );
  OR2_X1 U9373 ( .A1(n8125), .A2(n8034), .ZN(n9520) );
  OR2_X1 U9374 ( .A1(n9573), .A2(n9574), .ZN(n9519) );
  AND2_X1 U9375 ( .A1(n9516), .A2(n9515), .ZN(n9574) );
  AND2_X1 U9376 ( .A1(n9513), .A2(n9575), .ZN(n9573) );
  OR2_X1 U9377 ( .A1(n9515), .A2(n9516), .ZN(n9575) );
  OR2_X1 U9378 ( .A1(n8039), .A2(n8125), .ZN(n9516) );
  OR2_X1 U9379 ( .A1(n9576), .A2(n9577), .ZN(n9515) );
  AND2_X1 U9380 ( .A1(n9512), .A2(n9511), .ZN(n9577) );
  AND2_X1 U9381 ( .A1(n9509), .A2(n9578), .ZN(n9576) );
  OR2_X1 U9382 ( .A1(n9511), .A2(n9512), .ZN(n9578) );
  OR2_X1 U9383 ( .A1(n8125), .A2(n8043), .ZN(n9512) );
  OR2_X1 U9384 ( .A1(n9579), .A2(n9580), .ZN(n9511) );
  AND2_X1 U9385 ( .A1(n9508), .A2(n9507), .ZN(n9580) );
  AND2_X1 U9386 ( .A1(n9505), .A2(n9581), .ZN(n9579) );
  OR2_X1 U9387 ( .A1(n9507), .A2(n9508), .ZN(n9581) );
  OR2_X1 U9388 ( .A1(n8048), .A2(n8125), .ZN(n9508) );
  OR2_X1 U9389 ( .A1(n9582), .A2(n9583), .ZN(n9507) );
  AND2_X1 U9390 ( .A1(n9504), .A2(n9503), .ZN(n9583) );
  AND2_X1 U9391 ( .A1(n9501), .A2(n9584), .ZN(n9582) );
  OR2_X1 U9392 ( .A1(n9503), .A2(n9504), .ZN(n9584) );
  OR2_X1 U9393 ( .A1(n8125), .A2(n8052), .ZN(n9504) );
  OR2_X1 U9394 ( .A1(n9585), .A2(n9586), .ZN(n9503) );
  AND2_X1 U9395 ( .A1(n9500), .A2(n9499), .ZN(n9586) );
  AND2_X1 U9396 ( .A1(n9497), .A2(n9587), .ZN(n9585) );
  OR2_X1 U9397 ( .A1(n9499), .A2(n9500), .ZN(n9587) );
  OR2_X1 U9398 ( .A1(n8057), .A2(n8125), .ZN(n9500) );
  OR2_X1 U9399 ( .A1(n9588), .A2(n9589), .ZN(n9499) );
  AND2_X1 U9400 ( .A1(n9496), .A2(n9495), .ZN(n9589) );
  AND2_X1 U9401 ( .A1(n9493), .A2(n9590), .ZN(n9588) );
  OR2_X1 U9402 ( .A1(n9495), .A2(n9496), .ZN(n9590) );
  OR2_X1 U9403 ( .A1(n8125), .A2(n8061), .ZN(n9496) );
  OR2_X1 U9404 ( .A1(n9591), .A2(n9592), .ZN(n9495) );
  AND2_X1 U9405 ( .A1(n9492), .A2(n9491), .ZN(n9592) );
  AND2_X1 U9406 ( .A1(n9489), .A2(n9593), .ZN(n9591) );
  OR2_X1 U9407 ( .A1(n9491), .A2(n9492), .ZN(n9593) );
  OR2_X1 U9408 ( .A1(n8066), .A2(n8125), .ZN(n9492) );
  OR2_X1 U9409 ( .A1(n9594), .A2(n9595), .ZN(n9491) );
  AND2_X1 U9410 ( .A1(n9488), .A2(n9487), .ZN(n9595) );
  AND2_X1 U9411 ( .A1(n9485), .A2(n9596), .ZN(n9594) );
  OR2_X1 U9412 ( .A1(n9487), .A2(n9488), .ZN(n9596) );
  OR2_X1 U9413 ( .A1(n8125), .A2(n8070), .ZN(n9488) );
  OR2_X1 U9414 ( .A1(n9597), .A2(n9598), .ZN(n9487) );
  AND2_X1 U9415 ( .A1(n9484), .A2(n9483), .ZN(n9598) );
  AND2_X1 U9416 ( .A1(n9481), .A2(n9599), .ZN(n9597) );
  OR2_X1 U9417 ( .A1(n9483), .A2(n9484), .ZN(n9599) );
  OR2_X1 U9418 ( .A1(n8075), .A2(n8125), .ZN(n9484) );
  OR2_X1 U9419 ( .A1(n9600), .A2(n9601), .ZN(n9483) );
  AND2_X1 U9420 ( .A1(n9480), .A2(n9479), .ZN(n9601) );
  AND2_X1 U9421 ( .A1(n9477), .A2(n9602), .ZN(n9600) );
  OR2_X1 U9422 ( .A1(n9479), .A2(n9480), .ZN(n9602) );
  OR2_X1 U9423 ( .A1(n8125), .A2(n8079), .ZN(n9480) );
  OR2_X1 U9424 ( .A1(n9603), .A2(n9604), .ZN(n9479) );
  AND2_X1 U9425 ( .A1(n9476), .A2(n9475), .ZN(n9604) );
  AND2_X1 U9426 ( .A1(n9473), .A2(n9605), .ZN(n9603) );
  OR2_X1 U9427 ( .A1(n9475), .A2(n9476), .ZN(n9605) );
  OR2_X1 U9428 ( .A1(n8084), .A2(n8125), .ZN(n9476) );
  OR2_X1 U9429 ( .A1(n9606), .A2(n9607), .ZN(n9475) );
  AND2_X1 U9430 ( .A1(n9472), .A2(n9471), .ZN(n9607) );
  AND2_X1 U9431 ( .A1(n9469), .A2(n9608), .ZN(n9606) );
  OR2_X1 U9432 ( .A1(n9471), .A2(n9472), .ZN(n9608) );
  OR2_X1 U9433 ( .A1(n8125), .A2(n8088), .ZN(n9472) );
  OR2_X1 U9434 ( .A1(n9609), .A2(n9610), .ZN(n9471) );
  AND2_X1 U9435 ( .A1(n9468), .A2(n9467), .ZN(n9610) );
  AND2_X1 U9436 ( .A1(n9465), .A2(n9611), .ZN(n9609) );
  OR2_X1 U9437 ( .A1(n9467), .A2(n9468), .ZN(n9611) );
  OR2_X1 U9438 ( .A1(n8093), .A2(n8125), .ZN(n9468) );
  OR2_X1 U9439 ( .A1(n9612), .A2(n9613), .ZN(n9467) );
  AND2_X1 U9440 ( .A1(n9464), .A2(n9463), .ZN(n9613) );
  AND2_X1 U9441 ( .A1(n9461), .A2(n9614), .ZN(n9612) );
  OR2_X1 U9442 ( .A1(n9463), .A2(n9464), .ZN(n9614) );
  OR2_X1 U9443 ( .A1(n8125), .A2(n8097), .ZN(n9464) );
  OR2_X1 U9444 ( .A1(n9615), .A2(n9616), .ZN(n9463) );
  AND2_X1 U9445 ( .A1(n9460), .A2(n9459), .ZN(n9616) );
  AND2_X1 U9446 ( .A1(n9457), .A2(n9617), .ZN(n9615) );
  OR2_X1 U9447 ( .A1(n9459), .A2(n9460), .ZN(n9617) );
  OR2_X1 U9448 ( .A1(n8102), .A2(n8125), .ZN(n9460) );
  OR2_X1 U9449 ( .A1(n9618), .A2(n9619), .ZN(n9459) );
  AND2_X1 U9450 ( .A1(n9456), .A2(n9455), .ZN(n9619) );
  AND2_X1 U9451 ( .A1(n9453), .A2(n9620), .ZN(n9618) );
  OR2_X1 U9452 ( .A1(n9455), .A2(n9456), .ZN(n9620) );
  OR2_X1 U9453 ( .A1(n8125), .A2(n8106), .ZN(n9456) );
  OR2_X1 U9454 ( .A1(n9621), .A2(n9622), .ZN(n9455) );
  AND2_X1 U9455 ( .A1(n9452), .A2(n9451), .ZN(n9622) );
  AND2_X1 U9456 ( .A1(n9449), .A2(n9623), .ZN(n9621) );
  OR2_X1 U9457 ( .A1(n9451), .A2(n9452), .ZN(n9623) );
  OR2_X1 U9458 ( .A1(n8125), .A2(n8109), .ZN(n9452) );
  OR2_X1 U9459 ( .A1(n9624), .A2(n9625), .ZN(n9451) );
  AND2_X1 U9460 ( .A1(n9448), .A2(n9447), .ZN(n9625) );
  AND2_X1 U9461 ( .A1(n9445), .A2(n9626), .ZN(n9624) );
  OR2_X1 U9462 ( .A1(n9447), .A2(n9448), .ZN(n9626) );
  OR2_X1 U9463 ( .A1(n8125), .A2(n8112), .ZN(n9448) );
  OR2_X1 U9464 ( .A1(n9627), .A2(n9628), .ZN(n9447) );
  AND2_X1 U9465 ( .A1(n9444), .A2(n9443), .ZN(n9628) );
  AND2_X1 U9466 ( .A1(n9441), .A2(n9629), .ZN(n9627) );
  OR2_X1 U9467 ( .A1(n9443), .A2(n9444), .ZN(n9629) );
  OR2_X1 U9468 ( .A1(n8125), .A2(n8115), .ZN(n9444) );
  OR2_X1 U9469 ( .A1(n9630), .A2(n9631), .ZN(n9443) );
  AND2_X1 U9470 ( .A1(n9440), .A2(n9439), .ZN(n9631) );
  AND2_X1 U9471 ( .A1(n9437), .A2(n9632), .ZN(n9630) );
  OR2_X1 U9472 ( .A1(n9439), .A2(n9440), .ZN(n9632) );
  OR2_X1 U9473 ( .A1(n8125), .A2(n8118), .ZN(n9440) );
  OR2_X1 U9474 ( .A1(n9633), .A2(n9634), .ZN(n9439) );
  AND2_X1 U9475 ( .A1(n9436), .A2(n9435), .ZN(n9634) );
  AND2_X1 U9476 ( .A1(n9433), .A2(n9635), .ZN(n9633) );
  OR2_X1 U9477 ( .A1(n9435), .A2(n9436), .ZN(n9635) );
  OR2_X1 U9478 ( .A1(n8125), .A2(n8121), .ZN(n9436) );
  OR2_X1 U9479 ( .A1(n9636), .A2(n9637), .ZN(n9435) );
  AND2_X1 U9480 ( .A1(n7634), .A2(n9432), .ZN(n9637) );
  AND2_X1 U9481 ( .A1(n9430), .A2(n9638), .ZN(n9636) );
  OR2_X1 U9482 ( .A1(n9432), .A2(n7634), .ZN(n9638) );
  OR2_X1 U9483 ( .A1(n8124), .A2(n8125), .ZN(n7634) );
  OR2_X1 U9484 ( .A1(n9639), .A2(n9640), .ZN(n9432) );
  AND2_X1 U9485 ( .A1(n9426), .A2(n9429), .ZN(n9640) );
  AND2_X1 U9486 ( .A1(n9641), .A2(n9642), .ZN(n9639) );
  OR2_X1 U9487 ( .A1(n9429), .A2(n9426), .ZN(n9642) );
  OR2_X1 U9488 ( .A1(n8127), .A2(n8125), .ZN(n9426) );
  OR3_X1 U9489 ( .A1(n8981), .A2(n8125), .A3(n8122), .ZN(n9429) );
  INV_X1 U9490 ( .A(n9428), .ZN(n9641) );
  OR2_X1 U9491 ( .A1(n9643), .A2(n9644), .ZN(n9428) );
  AND2_X1 U9492 ( .A1(b_27_), .A2(n9645), .ZN(n9644) );
  OR2_X1 U9493 ( .A1(n9646), .A2(n7598), .ZN(n9645) );
  AND2_X1 U9494 ( .A1(a_30_), .A2(n8119), .ZN(n9646) );
  AND2_X1 U9495 ( .A1(b_26_), .A2(n9647), .ZN(n9643) );
  OR2_X1 U9496 ( .A1(n9648), .A2(n7601), .ZN(n9647) );
  AND2_X1 U9497 ( .A1(a_31_), .A2(n8122), .ZN(n9648) );
  XNOR2_X1 U9498 ( .A(n9649), .B(n9650), .ZN(n9430) );
  XOR2_X1 U9499 ( .A(n9651), .B(n9652), .Z(n9650) );
  XOR2_X1 U9500 ( .A(n9653), .B(n9654), .Z(n9433) );
  XOR2_X1 U9501 ( .A(n9655), .B(n9656), .Z(n9654) );
  XOR2_X1 U9502 ( .A(n9657), .B(n9658), .Z(n9437) );
  XOR2_X1 U9503 ( .A(n9659), .B(n7656), .Z(n9658) );
  XOR2_X1 U9504 ( .A(n9660), .B(n9661), .Z(n9441) );
  XOR2_X1 U9505 ( .A(n9662), .B(n9663), .Z(n9661) );
  XOR2_X1 U9506 ( .A(n9664), .B(n9665), .Z(n9445) );
  XOR2_X1 U9507 ( .A(n9666), .B(n9667), .Z(n9665) );
  XOR2_X1 U9508 ( .A(n9668), .B(n9669), .Z(n9449) );
  XOR2_X1 U9509 ( .A(n9670), .B(n9671), .Z(n9669) );
  XOR2_X1 U9510 ( .A(n9672), .B(n9673), .Z(n9453) );
  XOR2_X1 U9511 ( .A(n9674), .B(n9675), .Z(n9673) );
  XOR2_X1 U9512 ( .A(n9676), .B(n9677), .Z(n9457) );
  XOR2_X1 U9513 ( .A(n9678), .B(n9679), .Z(n9677) );
  XOR2_X1 U9514 ( .A(n9680), .B(n9681), .Z(n9461) );
  XOR2_X1 U9515 ( .A(n9682), .B(n9683), .Z(n9681) );
  XOR2_X1 U9516 ( .A(n9684), .B(n9685), .Z(n9465) );
  XOR2_X1 U9517 ( .A(n9686), .B(n9687), .Z(n9685) );
  XOR2_X1 U9518 ( .A(n9688), .B(n9689), .Z(n9469) );
  XOR2_X1 U9519 ( .A(n9690), .B(n9691), .Z(n9689) );
  XOR2_X1 U9520 ( .A(n9692), .B(n9693), .Z(n9473) );
  XOR2_X1 U9521 ( .A(n9694), .B(n9695), .Z(n9693) );
  XOR2_X1 U9522 ( .A(n9696), .B(n9697), .Z(n9477) );
  XOR2_X1 U9523 ( .A(n9698), .B(n9699), .Z(n9697) );
  XOR2_X1 U9524 ( .A(n9700), .B(n9701), .Z(n9481) );
  XOR2_X1 U9525 ( .A(n9702), .B(n9703), .Z(n9701) );
  XOR2_X1 U9526 ( .A(n9704), .B(n9705), .Z(n9485) );
  XOR2_X1 U9527 ( .A(n9706), .B(n9707), .Z(n9705) );
  XOR2_X1 U9528 ( .A(n9708), .B(n9709), .Z(n9489) );
  XOR2_X1 U9529 ( .A(n9710), .B(n9711), .Z(n9709) );
  XOR2_X1 U9530 ( .A(n9712), .B(n9713), .Z(n9493) );
  XOR2_X1 U9531 ( .A(n9714), .B(n9715), .Z(n9713) );
  XOR2_X1 U9532 ( .A(n9716), .B(n9717), .Z(n9497) );
  XOR2_X1 U9533 ( .A(n9718), .B(n9719), .Z(n9717) );
  XOR2_X1 U9534 ( .A(n9720), .B(n9721), .Z(n9501) );
  XOR2_X1 U9535 ( .A(n9722), .B(n9723), .Z(n9721) );
  XOR2_X1 U9536 ( .A(n9724), .B(n9725), .Z(n9505) );
  XOR2_X1 U9537 ( .A(n9726), .B(n9727), .Z(n9725) );
  XOR2_X1 U9538 ( .A(n9728), .B(n9729), .Z(n9509) );
  XOR2_X1 U9539 ( .A(n9730), .B(n9731), .Z(n9729) );
  XOR2_X1 U9540 ( .A(n9732), .B(n9733), .Z(n9513) );
  XOR2_X1 U9541 ( .A(n9734), .B(n9735), .Z(n9733) );
  XOR2_X1 U9542 ( .A(n9736), .B(n9737), .Z(n9517) );
  XOR2_X1 U9543 ( .A(n9738), .B(n9739), .Z(n9737) );
  XNOR2_X1 U9544 ( .A(n9740), .B(n9741), .ZN(n9521) );
  XNOR2_X1 U9545 ( .A(n9742), .B(n9743), .ZN(n9740) );
  XOR2_X1 U9546 ( .A(n9744), .B(n9745), .Z(n9525) );
  XOR2_X1 U9547 ( .A(n9746), .B(n9747), .Z(n9745) );
  XOR2_X1 U9548 ( .A(n9748), .B(n9749), .Z(n9529) );
  XOR2_X1 U9549 ( .A(n9750), .B(n9751), .Z(n9749) );
  OR2_X1 U9550 ( .A1(n8125), .A2(n8016), .ZN(n9535) );
  INV_X1 U9551 ( .A(b_28_), .ZN(n8125) );
  XOR2_X1 U9552 ( .A(n9752), .B(n9753), .Z(n9534) );
  XOR2_X1 U9553 ( .A(n9754), .B(n9755), .Z(n9753) );
  XNOR2_X1 U9554 ( .A(n9756), .B(n9757), .ZN(n9537) );
  XNOR2_X1 U9555 ( .A(n9758), .B(n9759), .ZN(n9756) );
  XOR2_X1 U9556 ( .A(n9760), .B(n9761), .Z(n9325) );
  XOR2_X1 U9557 ( .A(n9762), .B(n9763), .Z(n9761) );
  OR2_X1 U9558 ( .A1(n8870), .A2(n8869), .ZN(n8162) );
  XOR2_X1 U9559 ( .A(n8865), .B(n8867), .Z(n8869) );
  INV_X1 U9560 ( .A(n9543), .ZN(n8870) );
  OR2_X1 U9561 ( .A1(n9545), .A2(n9546), .ZN(n9543) );
  OR2_X1 U9562 ( .A1(n9764), .A2(n9765), .ZN(n9546) );
  AND2_X1 U9563 ( .A1(n9547), .A2(n9550), .ZN(n9765) );
  AND2_X1 U9564 ( .A1(n9766), .A2(n9549), .ZN(n9764) );
  OR2_X1 U9565 ( .A1(n9767), .A2(n9768), .ZN(n9549) );
  AND2_X1 U9566 ( .A1(n9760), .A2(n9763), .ZN(n9768) );
  AND2_X1 U9567 ( .A1(n9769), .A2(n9762), .ZN(n9767) );
  OR2_X1 U9568 ( .A1(n9770), .A2(n9771), .ZN(n9762) );
  AND2_X1 U9569 ( .A1(n9759), .A2(n9758), .ZN(n9771) );
  AND2_X1 U9570 ( .A1(n9757), .A2(n9772), .ZN(n9770) );
  OR2_X1 U9571 ( .A1(n9758), .A2(n9759), .ZN(n9772) );
  OR2_X1 U9572 ( .A1(n9773), .A2(n9774), .ZN(n9759) );
  AND2_X1 U9573 ( .A1(n9755), .A2(n9754), .ZN(n9774) );
  AND2_X1 U9574 ( .A1(n9752), .A2(n9775), .ZN(n9773) );
  OR2_X1 U9575 ( .A1(n9754), .A2(n9755), .ZN(n9775) );
  OR2_X1 U9576 ( .A1(n8021), .A2(n8122), .ZN(n9755) );
  OR2_X1 U9577 ( .A1(n9776), .A2(n9777), .ZN(n9754) );
  AND2_X1 U9578 ( .A1(n9751), .A2(n9750), .ZN(n9777) );
  AND2_X1 U9579 ( .A1(n9748), .A2(n9778), .ZN(n9776) );
  OR2_X1 U9580 ( .A1(n9750), .A2(n9751), .ZN(n9778) );
  OR2_X1 U9581 ( .A1(n8025), .A2(n8122), .ZN(n9751) );
  OR2_X1 U9582 ( .A1(n9779), .A2(n9780), .ZN(n9750) );
  AND2_X1 U9583 ( .A1(n9747), .A2(n9746), .ZN(n9780) );
  AND2_X1 U9584 ( .A1(n9744), .A2(n9781), .ZN(n9779) );
  OR2_X1 U9585 ( .A1(n9746), .A2(n9747), .ZN(n9781) );
  OR2_X1 U9586 ( .A1(n8030), .A2(n8122), .ZN(n9747) );
  OR2_X1 U9587 ( .A1(n9782), .A2(n9783), .ZN(n9746) );
  AND2_X1 U9588 ( .A1(n9743), .A2(n9742), .ZN(n9783) );
  AND2_X1 U9589 ( .A1(n9741), .A2(n9784), .ZN(n9782) );
  OR2_X1 U9590 ( .A1(n9742), .A2(n9743), .ZN(n9784) );
  OR2_X1 U9591 ( .A1(n9785), .A2(n9786), .ZN(n9743) );
  AND2_X1 U9592 ( .A1(n9739), .A2(n9738), .ZN(n9786) );
  AND2_X1 U9593 ( .A1(n9736), .A2(n9787), .ZN(n9785) );
  OR2_X1 U9594 ( .A1(n9738), .A2(n9739), .ZN(n9787) );
  OR2_X1 U9595 ( .A1(n8039), .A2(n8122), .ZN(n9739) );
  OR2_X1 U9596 ( .A1(n9788), .A2(n9789), .ZN(n9738) );
  AND2_X1 U9597 ( .A1(n9735), .A2(n9734), .ZN(n9789) );
  AND2_X1 U9598 ( .A1(n9732), .A2(n9790), .ZN(n9788) );
  OR2_X1 U9599 ( .A1(n9734), .A2(n9735), .ZN(n9790) );
  OR2_X1 U9600 ( .A1(n8043), .A2(n8122), .ZN(n9735) );
  OR2_X1 U9601 ( .A1(n9791), .A2(n9792), .ZN(n9734) );
  AND2_X1 U9602 ( .A1(n9731), .A2(n9730), .ZN(n9792) );
  AND2_X1 U9603 ( .A1(n9728), .A2(n9793), .ZN(n9791) );
  OR2_X1 U9604 ( .A1(n9730), .A2(n9731), .ZN(n9793) );
  OR2_X1 U9605 ( .A1(n8048), .A2(n8122), .ZN(n9731) );
  OR2_X1 U9606 ( .A1(n9794), .A2(n9795), .ZN(n9730) );
  AND2_X1 U9607 ( .A1(n9727), .A2(n9726), .ZN(n9795) );
  AND2_X1 U9608 ( .A1(n9724), .A2(n9796), .ZN(n9794) );
  OR2_X1 U9609 ( .A1(n9726), .A2(n9727), .ZN(n9796) );
  OR2_X1 U9610 ( .A1(n8052), .A2(n8122), .ZN(n9727) );
  OR2_X1 U9611 ( .A1(n9797), .A2(n9798), .ZN(n9726) );
  AND2_X1 U9612 ( .A1(n9723), .A2(n9722), .ZN(n9798) );
  AND2_X1 U9613 ( .A1(n9720), .A2(n9799), .ZN(n9797) );
  OR2_X1 U9614 ( .A1(n9722), .A2(n9723), .ZN(n9799) );
  OR2_X1 U9615 ( .A1(n8057), .A2(n8122), .ZN(n9723) );
  OR2_X1 U9616 ( .A1(n9800), .A2(n9801), .ZN(n9722) );
  AND2_X1 U9617 ( .A1(n9719), .A2(n9718), .ZN(n9801) );
  AND2_X1 U9618 ( .A1(n9716), .A2(n9802), .ZN(n9800) );
  OR2_X1 U9619 ( .A1(n9718), .A2(n9719), .ZN(n9802) );
  OR2_X1 U9620 ( .A1(n8061), .A2(n8122), .ZN(n9719) );
  OR2_X1 U9621 ( .A1(n9803), .A2(n9804), .ZN(n9718) );
  AND2_X1 U9622 ( .A1(n9715), .A2(n9714), .ZN(n9804) );
  AND2_X1 U9623 ( .A1(n9712), .A2(n9805), .ZN(n9803) );
  OR2_X1 U9624 ( .A1(n9714), .A2(n9715), .ZN(n9805) );
  OR2_X1 U9625 ( .A1(n8066), .A2(n8122), .ZN(n9715) );
  OR2_X1 U9626 ( .A1(n9806), .A2(n9807), .ZN(n9714) );
  AND2_X1 U9627 ( .A1(n9711), .A2(n9710), .ZN(n9807) );
  AND2_X1 U9628 ( .A1(n9708), .A2(n9808), .ZN(n9806) );
  OR2_X1 U9629 ( .A1(n9710), .A2(n9711), .ZN(n9808) );
  OR2_X1 U9630 ( .A1(n8070), .A2(n8122), .ZN(n9711) );
  OR2_X1 U9631 ( .A1(n9809), .A2(n9810), .ZN(n9710) );
  AND2_X1 U9632 ( .A1(n9707), .A2(n9706), .ZN(n9810) );
  AND2_X1 U9633 ( .A1(n9704), .A2(n9811), .ZN(n9809) );
  OR2_X1 U9634 ( .A1(n9706), .A2(n9707), .ZN(n9811) );
  OR2_X1 U9635 ( .A1(n8075), .A2(n8122), .ZN(n9707) );
  OR2_X1 U9636 ( .A1(n9812), .A2(n9813), .ZN(n9706) );
  AND2_X1 U9637 ( .A1(n9703), .A2(n9702), .ZN(n9813) );
  AND2_X1 U9638 ( .A1(n9700), .A2(n9814), .ZN(n9812) );
  OR2_X1 U9639 ( .A1(n9702), .A2(n9703), .ZN(n9814) );
  OR2_X1 U9640 ( .A1(n8079), .A2(n8122), .ZN(n9703) );
  OR2_X1 U9641 ( .A1(n9815), .A2(n9816), .ZN(n9702) );
  AND2_X1 U9642 ( .A1(n9699), .A2(n9698), .ZN(n9816) );
  AND2_X1 U9643 ( .A1(n9696), .A2(n9817), .ZN(n9815) );
  OR2_X1 U9644 ( .A1(n9698), .A2(n9699), .ZN(n9817) );
  OR2_X1 U9645 ( .A1(n8084), .A2(n8122), .ZN(n9699) );
  OR2_X1 U9646 ( .A1(n9818), .A2(n9819), .ZN(n9698) );
  AND2_X1 U9647 ( .A1(n9695), .A2(n9694), .ZN(n9819) );
  AND2_X1 U9648 ( .A1(n9692), .A2(n9820), .ZN(n9818) );
  OR2_X1 U9649 ( .A1(n9694), .A2(n9695), .ZN(n9820) );
  OR2_X1 U9650 ( .A1(n8088), .A2(n8122), .ZN(n9695) );
  OR2_X1 U9651 ( .A1(n9821), .A2(n9822), .ZN(n9694) );
  AND2_X1 U9652 ( .A1(n9691), .A2(n9690), .ZN(n9822) );
  AND2_X1 U9653 ( .A1(n9688), .A2(n9823), .ZN(n9821) );
  OR2_X1 U9654 ( .A1(n9690), .A2(n9691), .ZN(n9823) );
  OR2_X1 U9655 ( .A1(n8093), .A2(n8122), .ZN(n9691) );
  OR2_X1 U9656 ( .A1(n9824), .A2(n9825), .ZN(n9690) );
  AND2_X1 U9657 ( .A1(n9687), .A2(n9686), .ZN(n9825) );
  AND2_X1 U9658 ( .A1(n9684), .A2(n9826), .ZN(n9824) );
  OR2_X1 U9659 ( .A1(n9686), .A2(n9687), .ZN(n9826) );
  OR2_X1 U9660 ( .A1(n8097), .A2(n8122), .ZN(n9687) );
  OR2_X1 U9661 ( .A1(n9827), .A2(n9828), .ZN(n9686) );
  AND2_X1 U9662 ( .A1(n9683), .A2(n9682), .ZN(n9828) );
  AND2_X1 U9663 ( .A1(n9680), .A2(n9829), .ZN(n9827) );
  OR2_X1 U9664 ( .A1(n9682), .A2(n9683), .ZN(n9829) );
  OR2_X1 U9665 ( .A1(n8102), .A2(n8122), .ZN(n9683) );
  OR2_X1 U9666 ( .A1(n9830), .A2(n9831), .ZN(n9682) );
  AND2_X1 U9667 ( .A1(n9679), .A2(n9678), .ZN(n9831) );
  AND2_X1 U9668 ( .A1(n9676), .A2(n9832), .ZN(n9830) );
  OR2_X1 U9669 ( .A1(n9678), .A2(n9679), .ZN(n9832) );
  OR2_X1 U9670 ( .A1(n8106), .A2(n8122), .ZN(n9679) );
  OR2_X1 U9671 ( .A1(n9833), .A2(n9834), .ZN(n9678) );
  AND2_X1 U9672 ( .A1(n9675), .A2(n9674), .ZN(n9834) );
  AND2_X1 U9673 ( .A1(n9672), .A2(n9835), .ZN(n9833) );
  OR2_X1 U9674 ( .A1(n9674), .A2(n9675), .ZN(n9835) );
  OR2_X1 U9675 ( .A1(n8109), .A2(n8122), .ZN(n9675) );
  OR2_X1 U9676 ( .A1(n9836), .A2(n9837), .ZN(n9674) );
  AND2_X1 U9677 ( .A1(n9671), .A2(n9670), .ZN(n9837) );
  AND2_X1 U9678 ( .A1(n9668), .A2(n9838), .ZN(n9836) );
  OR2_X1 U9679 ( .A1(n9670), .A2(n9671), .ZN(n9838) );
  OR2_X1 U9680 ( .A1(n8112), .A2(n8122), .ZN(n9671) );
  OR2_X1 U9681 ( .A1(n9839), .A2(n9840), .ZN(n9670) );
  AND2_X1 U9682 ( .A1(n9667), .A2(n9666), .ZN(n9840) );
  AND2_X1 U9683 ( .A1(n9664), .A2(n9841), .ZN(n9839) );
  OR2_X1 U9684 ( .A1(n9666), .A2(n9667), .ZN(n9841) );
  OR2_X1 U9685 ( .A1(n8115), .A2(n8122), .ZN(n9667) );
  OR2_X1 U9686 ( .A1(n9842), .A2(n9843), .ZN(n9666) );
  AND2_X1 U9687 ( .A1(n9663), .A2(n9662), .ZN(n9843) );
  AND2_X1 U9688 ( .A1(n9660), .A2(n9844), .ZN(n9842) );
  OR2_X1 U9689 ( .A1(n9662), .A2(n9663), .ZN(n9844) );
  OR2_X1 U9690 ( .A1(n8118), .A2(n8122), .ZN(n9663) );
  OR2_X1 U9691 ( .A1(n9845), .A2(n9846), .ZN(n9662) );
  AND2_X1 U9692 ( .A1(n7656), .A2(n9659), .ZN(n9846) );
  AND2_X1 U9693 ( .A1(n9657), .A2(n9847), .ZN(n9845) );
  OR2_X1 U9694 ( .A1(n9659), .A2(n7656), .ZN(n9847) );
  OR2_X1 U9695 ( .A1(n8121), .A2(n8122), .ZN(n7656) );
  OR2_X1 U9696 ( .A1(n9848), .A2(n9849), .ZN(n9659) );
  AND2_X1 U9697 ( .A1(n9656), .A2(n9655), .ZN(n9849) );
  AND2_X1 U9698 ( .A1(n9653), .A2(n9850), .ZN(n9848) );
  OR2_X1 U9699 ( .A1(n9655), .A2(n9656), .ZN(n9850) );
  OR2_X1 U9700 ( .A1(n8124), .A2(n8122), .ZN(n9656) );
  OR2_X1 U9701 ( .A1(n9851), .A2(n9852), .ZN(n9655) );
  AND2_X1 U9702 ( .A1(n9649), .A2(n9652), .ZN(n9852) );
  AND2_X1 U9703 ( .A1(n9853), .A2(n9854), .ZN(n9851) );
  OR2_X1 U9704 ( .A1(n9652), .A2(n9649), .ZN(n9854) );
  OR2_X1 U9705 ( .A1(n8127), .A2(n8122), .ZN(n9649) );
  OR3_X1 U9706 ( .A1(n8981), .A2(n8119), .A3(n8122), .ZN(n9652) );
  INV_X1 U9707 ( .A(n9651), .ZN(n9853) );
  OR2_X1 U9708 ( .A1(n9855), .A2(n9856), .ZN(n9651) );
  AND2_X1 U9709 ( .A1(b_26_), .A2(n9857), .ZN(n9856) );
  OR2_X1 U9710 ( .A1(n9858), .A2(n7598), .ZN(n9857) );
  AND2_X1 U9711 ( .A1(a_30_), .A2(n8116), .ZN(n9858) );
  AND2_X1 U9712 ( .A1(b_25_), .A2(n9859), .ZN(n9855) );
  OR2_X1 U9713 ( .A1(n9860), .A2(n7601), .ZN(n9859) );
  AND2_X1 U9714 ( .A1(a_31_), .A2(n8119), .ZN(n9860) );
  XNOR2_X1 U9715 ( .A(n9861), .B(n9862), .ZN(n9653) );
  XOR2_X1 U9716 ( .A(n9863), .B(n9864), .Z(n9862) );
  XOR2_X1 U9717 ( .A(n9865), .B(n9866), .Z(n9657) );
  XOR2_X1 U9718 ( .A(n9867), .B(n9868), .Z(n9866) );
  XOR2_X1 U9719 ( .A(n9869), .B(n9870), .Z(n9660) );
  XOR2_X1 U9720 ( .A(n9871), .B(n9872), .Z(n9870) );
  XOR2_X1 U9721 ( .A(n9873), .B(n9874), .Z(n9664) );
  XOR2_X1 U9722 ( .A(n9875), .B(n7674), .Z(n9874) );
  XOR2_X1 U9723 ( .A(n9876), .B(n9877), .Z(n9668) );
  XOR2_X1 U9724 ( .A(n9878), .B(n9879), .Z(n9877) );
  XOR2_X1 U9725 ( .A(n9880), .B(n9881), .Z(n9672) );
  XOR2_X1 U9726 ( .A(n9882), .B(n9883), .Z(n9881) );
  XOR2_X1 U9727 ( .A(n9884), .B(n9885), .Z(n9676) );
  XOR2_X1 U9728 ( .A(n9886), .B(n9887), .Z(n9885) );
  XOR2_X1 U9729 ( .A(n9888), .B(n9889), .Z(n9680) );
  XOR2_X1 U9730 ( .A(n9890), .B(n9891), .Z(n9889) );
  XOR2_X1 U9731 ( .A(n9892), .B(n9893), .Z(n9684) );
  XOR2_X1 U9732 ( .A(n9894), .B(n9895), .Z(n9893) );
  XOR2_X1 U9733 ( .A(n9896), .B(n9897), .Z(n9688) );
  XOR2_X1 U9734 ( .A(n9898), .B(n9899), .Z(n9897) );
  XOR2_X1 U9735 ( .A(n9900), .B(n9901), .Z(n9692) );
  XOR2_X1 U9736 ( .A(n9902), .B(n9903), .Z(n9901) );
  XOR2_X1 U9737 ( .A(n9904), .B(n9905), .Z(n9696) );
  XOR2_X1 U9738 ( .A(n9906), .B(n9907), .Z(n9905) );
  XOR2_X1 U9739 ( .A(n9908), .B(n9909), .Z(n9700) );
  XOR2_X1 U9740 ( .A(n9910), .B(n9911), .Z(n9909) );
  XOR2_X1 U9741 ( .A(n9912), .B(n9913), .Z(n9704) );
  XOR2_X1 U9742 ( .A(n9914), .B(n9915), .Z(n9913) );
  XOR2_X1 U9743 ( .A(n9916), .B(n9917), .Z(n9708) );
  XOR2_X1 U9744 ( .A(n9918), .B(n9919), .Z(n9917) );
  XOR2_X1 U9745 ( .A(n9920), .B(n9921), .Z(n9712) );
  XOR2_X1 U9746 ( .A(n9922), .B(n9923), .Z(n9921) );
  XOR2_X1 U9747 ( .A(n9924), .B(n9925), .Z(n9716) );
  XOR2_X1 U9748 ( .A(n9926), .B(n9927), .Z(n9925) );
  XOR2_X1 U9749 ( .A(n9928), .B(n9929), .Z(n9720) );
  XOR2_X1 U9750 ( .A(n9930), .B(n9931), .Z(n9929) );
  XOR2_X1 U9751 ( .A(n9932), .B(n9933), .Z(n9724) );
  XOR2_X1 U9752 ( .A(n9934), .B(n9935), .Z(n9933) );
  XOR2_X1 U9753 ( .A(n9936), .B(n9937), .Z(n9728) );
  XOR2_X1 U9754 ( .A(n9938), .B(n9939), .Z(n9937) );
  XOR2_X1 U9755 ( .A(n9940), .B(n9941), .Z(n9732) );
  XOR2_X1 U9756 ( .A(n9942), .B(n9943), .Z(n9941) );
  XOR2_X1 U9757 ( .A(n9944), .B(n9945), .Z(n9736) );
  XOR2_X1 U9758 ( .A(n9946), .B(n9947), .Z(n9945) );
  OR2_X1 U9759 ( .A1(n8034), .A2(n8122), .ZN(n9742) );
  XOR2_X1 U9760 ( .A(n9948), .B(n9949), .Z(n9741) );
  XOR2_X1 U9761 ( .A(n9950), .B(n9951), .Z(n9949) );
  XNOR2_X1 U9762 ( .A(n9952), .B(n9953), .ZN(n9744) );
  XNOR2_X1 U9763 ( .A(n9954), .B(n9955), .ZN(n9952) );
  XOR2_X1 U9764 ( .A(n9956), .B(n9957), .Z(n9748) );
  XOR2_X1 U9765 ( .A(n9958), .B(n9959), .Z(n9957) );
  XOR2_X1 U9766 ( .A(n9960), .B(n9961), .Z(n9752) );
  XOR2_X1 U9767 ( .A(n9962), .B(n9963), .Z(n9961) );
  OR2_X1 U9768 ( .A1(n8016), .A2(n8122), .ZN(n9758) );
  XOR2_X1 U9769 ( .A(n9964), .B(n9965), .Z(n9757) );
  XOR2_X1 U9770 ( .A(n9966), .B(n9967), .Z(n9965) );
  OR2_X1 U9771 ( .A1(n9760), .A2(n9763), .ZN(n9769) );
  OR2_X1 U9772 ( .A1(n8012), .A2(n8122), .ZN(n9763) );
  XOR2_X1 U9773 ( .A(n9968), .B(n9969), .Z(n9760) );
  XOR2_X1 U9774 ( .A(n9970), .B(n9971), .Z(n9969) );
  OR2_X1 U9775 ( .A1(n9547), .A2(n9550), .ZN(n9766) );
  OR2_X1 U9776 ( .A1(n8297), .A2(n8122), .ZN(n9550) );
  INV_X1 U9777 ( .A(b_27_), .ZN(n8122) );
  XOR2_X1 U9778 ( .A(n9972), .B(n9973), .Z(n9547) );
  XOR2_X1 U9779 ( .A(n9974), .B(n9975), .Z(n9973) );
  XOR2_X1 U9780 ( .A(n9976), .B(n9977), .Z(n9545) );
  XOR2_X1 U9781 ( .A(n9978), .B(n9979), .Z(n9977) );
  OR2_X1 U9782 ( .A1(n9980), .A2(n8866), .ZN(n8169) );
  XOR2_X1 U9783 ( .A(n8842), .B(n8844), .Z(n8866) );
  OR2_X1 U9784 ( .A1(n9981), .A2(n9982), .ZN(n8844) );
  AND2_X1 U9785 ( .A1(n9983), .A2(n9984), .ZN(n9982) );
  AND2_X1 U9786 ( .A1(n9985), .A2(n9986), .ZN(n9981) );
  OR2_X1 U9787 ( .A1(n9983), .A2(n9984), .ZN(n9986) );
  XOR2_X1 U9788 ( .A(n8851), .B(n9987), .Z(n8842) );
  XOR2_X1 U9789 ( .A(n8850), .B(n8849), .Z(n9987) );
  OR2_X1 U9790 ( .A1(n8113), .A2(n8297), .ZN(n8849) );
  OR2_X1 U9791 ( .A1(n9988), .A2(n9989), .ZN(n8850) );
  AND2_X1 U9792 ( .A1(n9990), .A2(n9991), .ZN(n9989) );
  AND2_X1 U9793 ( .A1(n9992), .A2(n9993), .ZN(n9988) );
  OR2_X1 U9794 ( .A1(n9990), .A2(n9991), .ZN(n9993) );
  XOR2_X1 U9795 ( .A(n8858), .B(n9994), .Z(n8851) );
  XOR2_X1 U9796 ( .A(n8857), .B(n8856), .Z(n9994) );
  OR2_X1 U9797 ( .A1(n8012), .A2(n8110), .ZN(n8856) );
  OR2_X1 U9798 ( .A1(n9995), .A2(n9996), .ZN(n8857) );
  AND2_X1 U9799 ( .A1(n9997), .A2(n9998), .ZN(n9996) );
  AND2_X1 U9800 ( .A1(n9999), .A2(n10000), .ZN(n9995) );
  OR2_X1 U9801 ( .A1(n9997), .A2(n9998), .ZN(n10000) );
  XOR2_X1 U9802 ( .A(n10001), .B(n10002), .Z(n8858) );
  XOR2_X1 U9803 ( .A(n10003), .B(n10004), .Z(n10002) );
  AND2_X1 U9804 ( .A1(n8867), .A2(n8865), .ZN(n9980) );
  XNOR2_X1 U9805 ( .A(n9985), .B(n10005), .ZN(n8865) );
  XOR2_X1 U9806 ( .A(n9984), .B(n9983), .Z(n10005) );
  OR2_X1 U9807 ( .A1(n8297), .A2(n8116), .ZN(n9983) );
  OR2_X1 U9808 ( .A1(n10006), .A2(n10007), .ZN(n9984) );
  AND2_X1 U9809 ( .A1(n10008), .A2(n10009), .ZN(n10007) );
  AND2_X1 U9810 ( .A1(n10010), .A2(n10011), .ZN(n10006) );
  OR2_X1 U9811 ( .A1(n10008), .A2(n10009), .ZN(n10011) );
  XNOR2_X1 U9812 ( .A(n10012), .B(n9992), .ZN(n9985) );
  XOR2_X1 U9813 ( .A(n9999), .B(n10013), .Z(n9992) );
  XOR2_X1 U9814 ( .A(n9998), .B(n9997), .Z(n10013) );
  OR2_X1 U9815 ( .A1(n8016), .A2(n8110), .ZN(n9997) );
  OR2_X1 U9816 ( .A1(n10014), .A2(n10015), .ZN(n9998) );
  AND2_X1 U9817 ( .A1(n10016), .A2(n10017), .ZN(n10015) );
  AND2_X1 U9818 ( .A1(n10018), .A2(n10019), .ZN(n10014) );
  OR2_X1 U9819 ( .A1(n10016), .A2(n10017), .ZN(n10019) );
  XOR2_X1 U9820 ( .A(n10020), .B(n10021), .Z(n9999) );
  XOR2_X1 U9821 ( .A(n10022), .B(n10023), .Z(n10021) );
  XNOR2_X1 U9822 ( .A(n9991), .B(n9990), .ZN(n10012) );
  OR2_X1 U9823 ( .A1(n10024), .A2(n10025), .ZN(n9990) );
  AND2_X1 U9824 ( .A1(n10026), .A2(n10027), .ZN(n10025) );
  AND2_X1 U9825 ( .A1(n10028), .A2(n10029), .ZN(n10024) );
  OR2_X1 U9826 ( .A1(n10026), .A2(n10027), .ZN(n10029) );
  OR2_X1 U9827 ( .A1(n8113), .A2(n8012), .ZN(n9991) );
  INV_X1 U9828 ( .A(n10030), .ZN(n8867) );
  OR2_X1 U9829 ( .A1(n10031), .A2(n10032), .ZN(n10030) );
  AND2_X1 U9830 ( .A1(n9979), .A2(n9978), .ZN(n10032) );
  AND2_X1 U9831 ( .A1(n9976), .A2(n10033), .ZN(n10031) );
  OR2_X1 U9832 ( .A1(n9978), .A2(n9979), .ZN(n10033) );
  OR2_X1 U9833 ( .A1(n8119), .A2(n8297), .ZN(n9979) );
  OR2_X1 U9834 ( .A1(n10034), .A2(n10035), .ZN(n9978) );
  AND2_X1 U9835 ( .A1(n9975), .A2(n9974), .ZN(n10035) );
  AND2_X1 U9836 ( .A1(n9972), .A2(n10036), .ZN(n10034) );
  OR2_X1 U9837 ( .A1(n9974), .A2(n9975), .ZN(n10036) );
  OR2_X1 U9838 ( .A1(n8119), .A2(n8012), .ZN(n9975) );
  OR2_X1 U9839 ( .A1(n10037), .A2(n10038), .ZN(n9974) );
  AND2_X1 U9840 ( .A1(n9971), .A2(n9970), .ZN(n10038) );
  AND2_X1 U9841 ( .A1(n9968), .A2(n10039), .ZN(n10037) );
  OR2_X1 U9842 ( .A1(n9970), .A2(n9971), .ZN(n10039) );
  OR2_X1 U9843 ( .A1(n8119), .A2(n8016), .ZN(n9971) );
  OR2_X1 U9844 ( .A1(n10040), .A2(n10041), .ZN(n9970) );
  AND2_X1 U9845 ( .A1(n9967), .A2(n9966), .ZN(n10041) );
  AND2_X1 U9846 ( .A1(n9964), .A2(n10042), .ZN(n10040) );
  OR2_X1 U9847 ( .A1(n9966), .A2(n9967), .ZN(n10042) );
  OR2_X1 U9848 ( .A1(n8021), .A2(n8119), .ZN(n9967) );
  OR2_X1 U9849 ( .A1(n10043), .A2(n10044), .ZN(n9966) );
  AND2_X1 U9850 ( .A1(n9963), .A2(n9962), .ZN(n10044) );
  AND2_X1 U9851 ( .A1(n9960), .A2(n10045), .ZN(n10043) );
  OR2_X1 U9852 ( .A1(n9962), .A2(n9963), .ZN(n10045) );
  OR2_X1 U9853 ( .A1(n8119), .A2(n8025), .ZN(n9963) );
  OR2_X1 U9854 ( .A1(n10046), .A2(n10047), .ZN(n9962) );
  AND2_X1 U9855 ( .A1(n9959), .A2(n9958), .ZN(n10047) );
  AND2_X1 U9856 ( .A1(n9956), .A2(n10048), .ZN(n10046) );
  OR2_X1 U9857 ( .A1(n9958), .A2(n9959), .ZN(n10048) );
  OR2_X1 U9858 ( .A1(n8030), .A2(n8119), .ZN(n9959) );
  OR2_X1 U9859 ( .A1(n10049), .A2(n10050), .ZN(n9958) );
  AND2_X1 U9860 ( .A1(n9955), .A2(n9954), .ZN(n10050) );
  AND2_X1 U9861 ( .A1(n9953), .A2(n10051), .ZN(n10049) );
  OR2_X1 U9862 ( .A1(n9954), .A2(n9955), .ZN(n10051) );
  OR2_X1 U9863 ( .A1(n10052), .A2(n10053), .ZN(n9955) );
  AND2_X1 U9864 ( .A1(n9951), .A2(n9950), .ZN(n10053) );
  AND2_X1 U9865 ( .A1(n9948), .A2(n10054), .ZN(n10052) );
  OR2_X1 U9866 ( .A1(n9950), .A2(n9951), .ZN(n10054) );
  OR2_X1 U9867 ( .A1(n8039), .A2(n8119), .ZN(n9951) );
  OR2_X1 U9868 ( .A1(n10055), .A2(n10056), .ZN(n9950) );
  AND2_X1 U9869 ( .A1(n9947), .A2(n9946), .ZN(n10056) );
  AND2_X1 U9870 ( .A1(n9944), .A2(n10057), .ZN(n10055) );
  OR2_X1 U9871 ( .A1(n9946), .A2(n9947), .ZN(n10057) );
  OR2_X1 U9872 ( .A1(n8119), .A2(n8043), .ZN(n9947) );
  OR2_X1 U9873 ( .A1(n10058), .A2(n10059), .ZN(n9946) );
  AND2_X1 U9874 ( .A1(n9943), .A2(n9942), .ZN(n10059) );
  AND2_X1 U9875 ( .A1(n9940), .A2(n10060), .ZN(n10058) );
  OR2_X1 U9876 ( .A1(n9942), .A2(n9943), .ZN(n10060) );
  OR2_X1 U9877 ( .A1(n8048), .A2(n8119), .ZN(n9943) );
  OR2_X1 U9878 ( .A1(n10061), .A2(n10062), .ZN(n9942) );
  AND2_X1 U9879 ( .A1(n9939), .A2(n9938), .ZN(n10062) );
  AND2_X1 U9880 ( .A1(n9936), .A2(n10063), .ZN(n10061) );
  OR2_X1 U9881 ( .A1(n9938), .A2(n9939), .ZN(n10063) );
  OR2_X1 U9882 ( .A1(n8119), .A2(n8052), .ZN(n9939) );
  OR2_X1 U9883 ( .A1(n10064), .A2(n10065), .ZN(n9938) );
  AND2_X1 U9884 ( .A1(n9935), .A2(n9934), .ZN(n10065) );
  AND2_X1 U9885 ( .A1(n9932), .A2(n10066), .ZN(n10064) );
  OR2_X1 U9886 ( .A1(n9934), .A2(n9935), .ZN(n10066) );
  OR2_X1 U9887 ( .A1(n8057), .A2(n8119), .ZN(n9935) );
  OR2_X1 U9888 ( .A1(n10067), .A2(n10068), .ZN(n9934) );
  AND2_X1 U9889 ( .A1(n9931), .A2(n9930), .ZN(n10068) );
  AND2_X1 U9890 ( .A1(n9928), .A2(n10069), .ZN(n10067) );
  OR2_X1 U9891 ( .A1(n9930), .A2(n9931), .ZN(n10069) );
  OR2_X1 U9892 ( .A1(n8119), .A2(n8061), .ZN(n9931) );
  OR2_X1 U9893 ( .A1(n10070), .A2(n10071), .ZN(n9930) );
  AND2_X1 U9894 ( .A1(n9927), .A2(n9926), .ZN(n10071) );
  AND2_X1 U9895 ( .A1(n9924), .A2(n10072), .ZN(n10070) );
  OR2_X1 U9896 ( .A1(n9926), .A2(n9927), .ZN(n10072) );
  OR2_X1 U9897 ( .A1(n8066), .A2(n8119), .ZN(n9927) );
  OR2_X1 U9898 ( .A1(n10073), .A2(n10074), .ZN(n9926) );
  AND2_X1 U9899 ( .A1(n9923), .A2(n9922), .ZN(n10074) );
  AND2_X1 U9900 ( .A1(n9920), .A2(n10075), .ZN(n10073) );
  OR2_X1 U9901 ( .A1(n9922), .A2(n9923), .ZN(n10075) );
  OR2_X1 U9902 ( .A1(n8119), .A2(n8070), .ZN(n9923) );
  OR2_X1 U9903 ( .A1(n10076), .A2(n10077), .ZN(n9922) );
  AND2_X1 U9904 ( .A1(n9919), .A2(n9918), .ZN(n10077) );
  AND2_X1 U9905 ( .A1(n9916), .A2(n10078), .ZN(n10076) );
  OR2_X1 U9906 ( .A1(n9918), .A2(n9919), .ZN(n10078) );
  OR2_X1 U9907 ( .A1(n8075), .A2(n8119), .ZN(n9919) );
  OR2_X1 U9908 ( .A1(n10079), .A2(n10080), .ZN(n9918) );
  AND2_X1 U9909 ( .A1(n9915), .A2(n9914), .ZN(n10080) );
  AND2_X1 U9910 ( .A1(n9912), .A2(n10081), .ZN(n10079) );
  OR2_X1 U9911 ( .A1(n9914), .A2(n9915), .ZN(n10081) );
  OR2_X1 U9912 ( .A1(n8119), .A2(n8079), .ZN(n9915) );
  OR2_X1 U9913 ( .A1(n10082), .A2(n10083), .ZN(n9914) );
  AND2_X1 U9914 ( .A1(n9911), .A2(n9910), .ZN(n10083) );
  AND2_X1 U9915 ( .A1(n9908), .A2(n10084), .ZN(n10082) );
  OR2_X1 U9916 ( .A1(n9910), .A2(n9911), .ZN(n10084) );
  OR2_X1 U9917 ( .A1(n8084), .A2(n8119), .ZN(n9911) );
  OR2_X1 U9918 ( .A1(n10085), .A2(n10086), .ZN(n9910) );
  AND2_X1 U9919 ( .A1(n9907), .A2(n9906), .ZN(n10086) );
  AND2_X1 U9920 ( .A1(n9904), .A2(n10087), .ZN(n10085) );
  OR2_X1 U9921 ( .A1(n9906), .A2(n9907), .ZN(n10087) );
  OR2_X1 U9922 ( .A1(n8119), .A2(n8088), .ZN(n9907) );
  OR2_X1 U9923 ( .A1(n10088), .A2(n10089), .ZN(n9906) );
  AND2_X1 U9924 ( .A1(n9903), .A2(n9902), .ZN(n10089) );
  AND2_X1 U9925 ( .A1(n9900), .A2(n10090), .ZN(n10088) );
  OR2_X1 U9926 ( .A1(n9902), .A2(n9903), .ZN(n10090) );
  OR2_X1 U9927 ( .A1(n8093), .A2(n8119), .ZN(n9903) );
  OR2_X1 U9928 ( .A1(n10091), .A2(n10092), .ZN(n9902) );
  AND2_X1 U9929 ( .A1(n9899), .A2(n9898), .ZN(n10092) );
  AND2_X1 U9930 ( .A1(n9896), .A2(n10093), .ZN(n10091) );
  OR2_X1 U9931 ( .A1(n9898), .A2(n9899), .ZN(n10093) );
  OR2_X1 U9932 ( .A1(n8119), .A2(n8097), .ZN(n9899) );
  OR2_X1 U9933 ( .A1(n10094), .A2(n10095), .ZN(n9898) );
  AND2_X1 U9934 ( .A1(n9895), .A2(n9894), .ZN(n10095) );
  AND2_X1 U9935 ( .A1(n9892), .A2(n10096), .ZN(n10094) );
  OR2_X1 U9936 ( .A1(n9894), .A2(n9895), .ZN(n10096) );
  OR2_X1 U9937 ( .A1(n8102), .A2(n8119), .ZN(n9895) );
  OR2_X1 U9938 ( .A1(n10097), .A2(n10098), .ZN(n9894) );
  AND2_X1 U9939 ( .A1(n9891), .A2(n9890), .ZN(n10098) );
  AND2_X1 U9940 ( .A1(n9888), .A2(n10099), .ZN(n10097) );
  OR2_X1 U9941 ( .A1(n9890), .A2(n9891), .ZN(n10099) );
  OR2_X1 U9942 ( .A1(n8119), .A2(n8106), .ZN(n9891) );
  OR2_X1 U9943 ( .A1(n10100), .A2(n10101), .ZN(n9890) );
  AND2_X1 U9944 ( .A1(n9887), .A2(n9886), .ZN(n10101) );
  AND2_X1 U9945 ( .A1(n9884), .A2(n10102), .ZN(n10100) );
  OR2_X1 U9946 ( .A1(n9886), .A2(n9887), .ZN(n10102) );
  OR2_X1 U9947 ( .A1(n8119), .A2(n8109), .ZN(n9887) );
  OR2_X1 U9948 ( .A1(n10103), .A2(n10104), .ZN(n9886) );
  AND2_X1 U9949 ( .A1(n9883), .A2(n9882), .ZN(n10104) );
  AND2_X1 U9950 ( .A1(n9880), .A2(n10105), .ZN(n10103) );
  OR2_X1 U9951 ( .A1(n9882), .A2(n9883), .ZN(n10105) );
  OR2_X1 U9952 ( .A1(n8119), .A2(n8112), .ZN(n9883) );
  OR2_X1 U9953 ( .A1(n10106), .A2(n10107), .ZN(n9882) );
  AND2_X1 U9954 ( .A1(n9879), .A2(n9878), .ZN(n10107) );
  AND2_X1 U9955 ( .A1(n9876), .A2(n10108), .ZN(n10106) );
  OR2_X1 U9956 ( .A1(n9878), .A2(n9879), .ZN(n10108) );
  OR2_X1 U9957 ( .A1(n8119), .A2(n8115), .ZN(n9879) );
  OR2_X1 U9958 ( .A1(n10109), .A2(n10110), .ZN(n9878) );
  AND2_X1 U9959 ( .A1(n7674), .A2(n9875), .ZN(n10110) );
  AND2_X1 U9960 ( .A1(n9873), .A2(n10111), .ZN(n10109) );
  OR2_X1 U9961 ( .A1(n9875), .A2(n7674), .ZN(n10111) );
  OR2_X1 U9962 ( .A1(n8118), .A2(n8119), .ZN(n7674) );
  OR2_X1 U9963 ( .A1(n10112), .A2(n10113), .ZN(n9875) );
  AND2_X1 U9964 ( .A1(n9872), .A2(n9871), .ZN(n10113) );
  AND2_X1 U9965 ( .A1(n9869), .A2(n10114), .ZN(n10112) );
  OR2_X1 U9966 ( .A1(n9871), .A2(n9872), .ZN(n10114) );
  OR2_X1 U9967 ( .A1(n8121), .A2(n8119), .ZN(n9872) );
  OR2_X1 U9968 ( .A1(n10115), .A2(n10116), .ZN(n9871) );
  AND2_X1 U9969 ( .A1(n9868), .A2(n9867), .ZN(n10116) );
  AND2_X1 U9970 ( .A1(n9865), .A2(n10117), .ZN(n10115) );
  OR2_X1 U9971 ( .A1(n9867), .A2(n9868), .ZN(n10117) );
  OR2_X1 U9972 ( .A1(n8124), .A2(n8119), .ZN(n9868) );
  OR2_X1 U9973 ( .A1(n10118), .A2(n10119), .ZN(n9867) );
  AND2_X1 U9974 ( .A1(n9861), .A2(n9864), .ZN(n10119) );
  AND2_X1 U9975 ( .A1(n10120), .A2(n10121), .ZN(n10118) );
  OR2_X1 U9976 ( .A1(n9864), .A2(n9861), .ZN(n10121) );
  OR2_X1 U9977 ( .A1(n8127), .A2(n8119), .ZN(n9861) );
  OR3_X1 U9978 ( .A1(n8981), .A2(n8119), .A3(n8116), .ZN(n9864) );
  INV_X1 U9979 ( .A(n9863), .ZN(n10120) );
  OR2_X1 U9980 ( .A1(n10122), .A2(n10123), .ZN(n9863) );
  AND2_X1 U9981 ( .A1(b_25_), .A2(n10124), .ZN(n10123) );
  OR2_X1 U9982 ( .A1(n10125), .A2(n7598), .ZN(n10124) );
  AND2_X1 U9983 ( .A1(a_30_), .A2(n8113), .ZN(n10125) );
  AND2_X1 U9984 ( .A1(b_24_), .A2(n10126), .ZN(n10122) );
  OR2_X1 U9985 ( .A1(n10127), .A2(n7601), .ZN(n10126) );
  AND2_X1 U9986 ( .A1(a_31_), .A2(n8116), .ZN(n10127) );
  XNOR2_X1 U9987 ( .A(n10128), .B(n10129), .ZN(n9865) );
  XOR2_X1 U9988 ( .A(n10130), .B(n10131), .Z(n10129) );
  XOR2_X1 U9989 ( .A(n10132), .B(n10133), .Z(n9869) );
  XOR2_X1 U9990 ( .A(n10134), .B(n10135), .Z(n10133) );
  XOR2_X1 U9991 ( .A(n10136), .B(n10137), .Z(n9873) );
  XOR2_X1 U9992 ( .A(n10138), .B(n10139), .Z(n10137) );
  XOR2_X1 U9993 ( .A(n10140), .B(n10141), .Z(n9876) );
  XOR2_X1 U9994 ( .A(n10142), .B(n10143), .Z(n10141) );
  XOR2_X1 U9995 ( .A(n10144), .B(n10145), .Z(n9880) );
  XOR2_X1 U9996 ( .A(n10146), .B(n7686), .Z(n10145) );
  XOR2_X1 U9997 ( .A(n10147), .B(n10148), .Z(n9884) );
  XOR2_X1 U9998 ( .A(n10149), .B(n10150), .Z(n10148) );
  XOR2_X1 U9999 ( .A(n10151), .B(n10152), .Z(n9888) );
  XOR2_X1 U10000 ( .A(n10153), .B(n10154), .Z(n10152) );
  XOR2_X1 U10001 ( .A(n10155), .B(n10156), .Z(n9892) );
  XOR2_X1 U10002 ( .A(n10157), .B(n10158), .Z(n10156) );
  XOR2_X1 U10003 ( .A(n10159), .B(n10160), .Z(n9896) );
  XOR2_X1 U10004 ( .A(n10161), .B(n10162), .Z(n10160) );
  XOR2_X1 U10005 ( .A(n10163), .B(n10164), .Z(n9900) );
  XOR2_X1 U10006 ( .A(n10165), .B(n10166), .Z(n10164) );
  XOR2_X1 U10007 ( .A(n10167), .B(n10168), .Z(n9904) );
  XOR2_X1 U10008 ( .A(n10169), .B(n10170), .Z(n10168) );
  XOR2_X1 U10009 ( .A(n10171), .B(n10172), .Z(n9908) );
  XOR2_X1 U10010 ( .A(n10173), .B(n10174), .Z(n10172) );
  XOR2_X1 U10011 ( .A(n10175), .B(n10176), .Z(n9912) );
  XOR2_X1 U10012 ( .A(n10177), .B(n10178), .Z(n10176) );
  XOR2_X1 U10013 ( .A(n10179), .B(n10180), .Z(n9916) );
  XOR2_X1 U10014 ( .A(n10181), .B(n10182), .Z(n10180) );
  XOR2_X1 U10015 ( .A(n10183), .B(n10184), .Z(n9920) );
  XOR2_X1 U10016 ( .A(n10185), .B(n10186), .Z(n10184) );
  XOR2_X1 U10017 ( .A(n10187), .B(n10188), .Z(n9924) );
  XOR2_X1 U10018 ( .A(n10189), .B(n10190), .Z(n10188) );
  XOR2_X1 U10019 ( .A(n10191), .B(n10192), .Z(n9928) );
  XOR2_X1 U10020 ( .A(n10193), .B(n10194), .Z(n10192) );
  XOR2_X1 U10021 ( .A(n10195), .B(n10196), .Z(n9932) );
  XOR2_X1 U10022 ( .A(n10197), .B(n10198), .Z(n10196) );
  XOR2_X1 U10023 ( .A(n10199), .B(n10200), .Z(n9936) );
  XOR2_X1 U10024 ( .A(n10201), .B(n10202), .Z(n10200) );
  XNOR2_X1 U10025 ( .A(n10203), .B(n10204), .ZN(n9940) );
  XNOR2_X1 U10026 ( .A(n10205), .B(n10206), .ZN(n10203) );
  XOR2_X1 U10027 ( .A(n10207), .B(n10208), .Z(n9944) );
  XOR2_X1 U10028 ( .A(n10209), .B(n10210), .Z(n10208) );
  XOR2_X1 U10029 ( .A(n10211), .B(n10212), .Z(n9948) );
  XOR2_X1 U10030 ( .A(n10213), .B(n10214), .Z(n10212) );
  OR2_X1 U10031 ( .A1(n8119), .A2(n8034), .ZN(n9954) );
  INV_X1 U10032 ( .A(b_26_), .ZN(n8119) );
  XOR2_X1 U10033 ( .A(n10215), .B(n10216), .Z(n9953) );
  XOR2_X1 U10034 ( .A(n10217), .B(n10218), .Z(n10216) );
  XNOR2_X1 U10035 ( .A(n10219), .B(n10220), .ZN(n9956) );
  XNOR2_X1 U10036 ( .A(n10221), .B(n10222), .ZN(n10219) );
  XOR2_X1 U10037 ( .A(n10223), .B(n10224), .Z(n9960) );
  XOR2_X1 U10038 ( .A(n10225), .B(n10226), .Z(n10224) );
  XOR2_X1 U10039 ( .A(n10227), .B(n10228), .Z(n9964) );
  XOR2_X1 U10040 ( .A(n10229), .B(n10230), .Z(n10228) );
  XOR2_X1 U10041 ( .A(n10231), .B(n10232), .Z(n9968) );
  XOR2_X1 U10042 ( .A(n10233), .B(n10234), .Z(n10232) );
  XOR2_X1 U10043 ( .A(n10235), .B(n10236), .Z(n9972) );
  XOR2_X1 U10044 ( .A(n10237), .B(n10238), .Z(n10236) );
  XOR2_X1 U10045 ( .A(n10010), .B(n10239), .Z(n9976) );
  XOR2_X1 U10046 ( .A(n10009), .B(n10008), .Z(n10239) );
  OR2_X1 U10047 ( .A1(n8012), .A2(n8116), .ZN(n10008) );
  OR2_X1 U10048 ( .A1(n10240), .A2(n10241), .ZN(n10009) );
  AND2_X1 U10049 ( .A1(n10238), .A2(n10237), .ZN(n10241) );
  AND2_X1 U10050 ( .A1(n10235), .A2(n10242), .ZN(n10240) );
  OR2_X1 U10051 ( .A1(n10238), .A2(n10237), .ZN(n10242) );
  OR2_X1 U10052 ( .A1(n10243), .A2(n10244), .ZN(n10237) );
  AND2_X1 U10053 ( .A1(n10234), .A2(n10233), .ZN(n10244) );
  AND2_X1 U10054 ( .A1(n10231), .A2(n10245), .ZN(n10243) );
  OR2_X1 U10055 ( .A1(n10234), .A2(n10233), .ZN(n10245) );
  OR2_X1 U10056 ( .A1(n10246), .A2(n10247), .ZN(n10233) );
  AND2_X1 U10057 ( .A1(n10230), .A2(n10229), .ZN(n10247) );
  AND2_X1 U10058 ( .A1(n10227), .A2(n10248), .ZN(n10246) );
  OR2_X1 U10059 ( .A1(n10230), .A2(n10229), .ZN(n10248) );
  OR2_X1 U10060 ( .A1(n10249), .A2(n10250), .ZN(n10229) );
  AND2_X1 U10061 ( .A1(n10226), .A2(n10225), .ZN(n10250) );
  AND2_X1 U10062 ( .A1(n10223), .A2(n10251), .ZN(n10249) );
  OR2_X1 U10063 ( .A1(n10226), .A2(n10225), .ZN(n10251) );
  OR2_X1 U10064 ( .A1(n10252), .A2(n10253), .ZN(n10225) );
  AND2_X1 U10065 ( .A1(n10222), .A2(n10221), .ZN(n10253) );
  AND2_X1 U10066 ( .A1(n10220), .A2(n10254), .ZN(n10252) );
  OR2_X1 U10067 ( .A1(n10222), .A2(n10221), .ZN(n10254) );
  OR2_X1 U10068 ( .A1(n8034), .A2(n8116), .ZN(n10221) );
  OR2_X1 U10069 ( .A1(n10255), .A2(n10256), .ZN(n10222) );
  AND2_X1 U10070 ( .A1(n10218), .A2(n10217), .ZN(n10256) );
  AND2_X1 U10071 ( .A1(n10215), .A2(n10257), .ZN(n10255) );
  OR2_X1 U10072 ( .A1(n10218), .A2(n10217), .ZN(n10257) );
  OR2_X1 U10073 ( .A1(n10258), .A2(n10259), .ZN(n10217) );
  AND2_X1 U10074 ( .A1(n10214), .A2(n10213), .ZN(n10259) );
  AND2_X1 U10075 ( .A1(n10211), .A2(n10260), .ZN(n10258) );
  OR2_X1 U10076 ( .A1(n10214), .A2(n10213), .ZN(n10260) );
  OR2_X1 U10077 ( .A1(n10261), .A2(n10262), .ZN(n10213) );
  AND2_X1 U10078 ( .A1(n10210), .A2(n10209), .ZN(n10262) );
  AND2_X1 U10079 ( .A1(n10207), .A2(n10263), .ZN(n10261) );
  OR2_X1 U10080 ( .A1(n10210), .A2(n10209), .ZN(n10263) );
  OR2_X1 U10081 ( .A1(n10264), .A2(n10265), .ZN(n10209) );
  AND2_X1 U10082 ( .A1(n10206), .A2(n10205), .ZN(n10265) );
  AND2_X1 U10083 ( .A1(n10204), .A2(n10266), .ZN(n10264) );
  OR2_X1 U10084 ( .A1(n10206), .A2(n10205), .ZN(n10266) );
  OR2_X1 U10085 ( .A1(n8052), .A2(n8116), .ZN(n10205) );
  OR2_X1 U10086 ( .A1(n10267), .A2(n10268), .ZN(n10206) );
  AND2_X1 U10087 ( .A1(n10202), .A2(n10201), .ZN(n10268) );
  AND2_X1 U10088 ( .A1(n10199), .A2(n10269), .ZN(n10267) );
  OR2_X1 U10089 ( .A1(n10202), .A2(n10201), .ZN(n10269) );
  OR2_X1 U10090 ( .A1(n10270), .A2(n10271), .ZN(n10201) );
  AND2_X1 U10091 ( .A1(n10198), .A2(n10197), .ZN(n10271) );
  AND2_X1 U10092 ( .A1(n10195), .A2(n10272), .ZN(n10270) );
  OR2_X1 U10093 ( .A1(n10198), .A2(n10197), .ZN(n10272) );
  OR2_X1 U10094 ( .A1(n10273), .A2(n10274), .ZN(n10197) );
  AND2_X1 U10095 ( .A1(n10194), .A2(n10193), .ZN(n10274) );
  AND2_X1 U10096 ( .A1(n10191), .A2(n10275), .ZN(n10273) );
  OR2_X1 U10097 ( .A1(n10194), .A2(n10193), .ZN(n10275) );
  OR2_X1 U10098 ( .A1(n10276), .A2(n10277), .ZN(n10193) );
  AND2_X1 U10099 ( .A1(n10190), .A2(n10189), .ZN(n10277) );
  AND2_X1 U10100 ( .A1(n10187), .A2(n10278), .ZN(n10276) );
  OR2_X1 U10101 ( .A1(n10190), .A2(n10189), .ZN(n10278) );
  OR2_X1 U10102 ( .A1(n10279), .A2(n10280), .ZN(n10189) );
  AND2_X1 U10103 ( .A1(n10186), .A2(n10185), .ZN(n10280) );
  AND2_X1 U10104 ( .A1(n10183), .A2(n10281), .ZN(n10279) );
  OR2_X1 U10105 ( .A1(n10186), .A2(n10185), .ZN(n10281) );
  OR2_X1 U10106 ( .A1(n10282), .A2(n10283), .ZN(n10185) );
  AND2_X1 U10107 ( .A1(n10182), .A2(n10181), .ZN(n10283) );
  AND2_X1 U10108 ( .A1(n10179), .A2(n10284), .ZN(n10282) );
  OR2_X1 U10109 ( .A1(n10182), .A2(n10181), .ZN(n10284) );
  OR2_X1 U10110 ( .A1(n10285), .A2(n10286), .ZN(n10181) );
  AND2_X1 U10111 ( .A1(n10178), .A2(n10177), .ZN(n10286) );
  AND2_X1 U10112 ( .A1(n10175), .A2(n10287), .ZN(n10285) );
  OR2_X1 U10113 ( .A1(n10178), .A2(n10177), .ZN(n10287) );
  OR2_X1 U10114 ( .A1(n10288), .A2(n10289), .ZN(n10177) );
  AND2_X1 U10115 ( .A1(n10174), .A2(n10173), .ZN(n10289) );
  AND2_X1 U10116 ( .A1(n10171), .A2(n10290), .ZN(n10288) );
  OR2_X1 U10117 ( .A1(n10174), .A2(n10173), .ZN(n10290) );
  OR2_X1 U10118 ( .A1(n10291), .A2(n10292), .ZN(n10173) );
  AND2_X1 U10119 ( .A1(n10170), .A2(n10169), .ZN(n10292) );
  AND2_X1 U10120 ( .A1(n10167), .A2(n10293), .ZN(n10291) );
  OR2_X1 U10121 ( .A1(n10170), .A2(n10169), .ZN(n10293) );
  OR2_X1 U10122 ( .A1(n10294), .A2(n10295), .ZN(n10169) );
  AND2_X1 U10123 ( .A1(n10166), .A2(n10165), .ZN(n10295) );
  AND2_X1 U10124 ( .A1(n10163), .A2(n10296), .ZN(n10294) );
  OR2_X1 U10125 ( .A1(n10166), .A2(n10165), .ZN(n10296) );
  OR2_X1 U10126 ( .A1(n10297), .A2(n10298), .ZN(n10165) );
  AND2_X1 U10127 ( .A1(n10162), .A2(n10161), .ZN(n10298) );
  AND2_X1 U10128 ( .A1(n10159), .A2(n10299), .ZN(n10297) );
  OR2_X1 U10129 ( .A1(n10162), .A2(n10161), .ZN(n10299) );
  OR2_X1 U10130 ( .A1(n10300), .A2(n10301), .ZN(n10161) );
  AND2_X1 U10131 ( .A1(n10158), .A2(n10157), .ZN(n10301) );
  AND2_X1 U10132 ( .A1(n10155), .A2(n10302), .ZN(n10300) );
  OR2_X1 U10133 ( .A1(n10158), .A2(n10157), .ZN(n10302) );
  OR2_X1 U10134 ( .A1(n10303), .A2(n10304), .ZN(n10157) );
  AND2_X1 U10135 ( .A1(n10154), .A2(n10153), .ZN(n10304) );
  AND2_X1 U10136 ( .A1(n10151), .A2(n10305), .ZN(n10303) );
  OR2_X1 U10137 ( .A1(n10154), .A2(n10153), .ZN(n10305) );
  OR2_X1 U10138 ( .A1(n10306), .A2(n10307), .ZN(n10153) );
  AND2_X1 U10139 ( .A1(n10150), .A2(n10149), .ZN(n10307) );
  AND2_X1 U10140 ( .A1(n10147), .A2(n10308), .ZN(n10306) );
  OR2_X1 U10141 ( .A1(n10150), .A2(n10149), .ZN(n10308) );
  OR2_X1 U10142 ( .A1(n10309), .A2(n10310), .ZN(n10149) );
  AND2_X1 U10143 ( .A1(n7686), .A2(n10146), .ZN(n10310) );
  AND2_X1 U10144 ( .A1(n10144), .A2(n10311), .ZN(n10309) );
  OR2_X1 U10145 ( .A1(n7686), .A2(n10146), .ZN(n10311) );
  OR2_X1 U10146 ( .A1(n10312), .A2(n10313), .ZN(n10146) );
  AND2_X1 U10147 ( .A1(n10143), .A2(n10142), .ZN(n10313) );
  AND2_X1 U10148 ( .A1(n10140), .A2(n10314), .ZN(n10312) );
  OR2_X1 U10149 ( .A1(n10143), .A2(n10142), .ZN(n10314) );
  OR2_X1 U10150 ( .A1(n10315), .A2(n10316), .ZN(n10142) );
  AND2_X1 U10151 ( .A1(n10139), .A2(n10138), .ZN(n10316) );
  AND2_X1 U10152 ( .A1(n10136), .A2(n10317), .ZN(n10315) );
  OR2_X1 U10153 ( .A1(n10139), .A2(n10138), .ZN(n10317) );
  OR2_X1 U10154 ( .A1(n10318), .A2(n10319), .ZN(n10138) );
  AND2_X1 U10155 ( .A1(n10135), .A2(n10134), .ZN(n10319) );
  AND2_X1 U10156 ( .A1(n10132), .A2(n10320), .ZN(n10318) );
  OR2_X1 U10157 ( .A1(n10135), .A2(n10134), .ZN(n10320) );
  OR2_X1 U10158 ( .A1(n10321), .A2(n10322), .ZN(n10134) );
  AND2_X1 U10159 ( .A1(n10128), .A2(n10131), .ZN(n10322) );
  AND2_X1 U10160 ( .A1(n10323), .A2(n10324), .ZN(n10321) );
  OR2_X1 U10161 ( .A1(n10128), .A2(n10131), .ZN(n10324) );
  OR3_X1 U10162 ( .A1(n8981), .A2(n8113), .A3(n8116), .ZN(n10131) );
  OR2_X1 U10163 ( .A1(n8127), .A2(n8116), .ZN(n10128) );
  INV_X1 U10164 ( .A(n10130), .ZN(n10323) );
  OR2_X1 U10165 ( .A1(n10325), .A2(n10326), .ZN(n10130) );
  AND2_X1 U10166 ( .A1(b_24_), .A2(n10327), .ZN(n10326) );
  OR2_X1 U10167 ( .A1(n10328), .A2(n7598), .ZN(n10327) );
  AND2_X1 U10168 ( .A1(a_30_), .A2(n8110), .ZN(n10328) );
  AND2_X1 U10169 ( .A1(b_23_), .A2(n10329), .ZN(n10325) );
  OR2_X1 U10170 ( .A1(n10330), .A2(n7601), .ZN(n10329) );
  AND2_X1 U10171 ( .A1(a_31_), .A2(n8113), .ZN(n10330) );
  OR2_X1 U10172 ( .A1(n8124), .A2(n8116), .ZN(n10135) );
  XNOR2_X1 U10173 ( .A(n10331), .B(n10332), .ZN(n10132) );
  XOR2_X1 U10174 ( .A(n10333), .B(n10334), .Z(n10332) );
  OR2_X1 U10175 ( .A1(n8121), .A2(n8116), .ZN(n10139) );
  XOR2_X1 U10176 ( .A(n10335), .B(n10336), .Z(n10136) );
  XOR2_X1 U10177 ( .A(n10337), .B(n10338), .Z(n10336) );
  OR2_X1 U10178 ( .A1(n8118), .A2(n8116), .ZN(n10143) );
  XOR2_X1 U10179 ( .A(n10339), .B(n10340), .Z(n10140) );
  XOR2_X1 U10180 ( .A(n10341), .B(n10342), .Z(n10340) );
  OR2_X1 U10181 ( .A1(n8115), .A2(n8116), .ZN(n7686) );
  XOR2_X1 U10182 ( .A(n10343), .B(n10344), .Z(n10144) );
  XOR2_X1 U10183 ( .A(n10345), .B(n10346), .Z(n10344) );
  OR2_X1 U10184 ( .A1(n8112), .A2(n8116), .ZN(n10150) );
  XOR2_X1 U10185 ( .A(n10347), .B(n10348), .Z(n10147) );
  XOR2_X1 U10186 ( .A(n10349), .B(n10350), .Z(n10348) );
  OR2_X1 U10187 ( .A1(n8109), .A2(n8116), .ZN(n10154) );
  XOR2_X1 U10188 ( .A(n10351), .B(n10352), .Z(n10151) );
  XOR2_X1 U10189 ( .A(n10353), .B(n7704), .Z(n10352) );
  OR2_X1 U10190 ( .A1(n8106), .A2(n8116), .ZN(n10158) );
  XOR2_X1 U10191 ( .A(n10354), .B(n10355), .Z(n10155) );
  XOR2_X1 U10192 ( .A(n10356), .B(n10357), .Z(n10355) );
  OR2_X1 U10193 ( .A1(n8102), .A2(n8116), .ZN(n10162) );
  XOR2_X1 U10194 ( .A(n10358), .B(n10359), .Z(n10159) );
  XOR2_X1 U10195 ( .A(n10360), .B(n10361), .Z(n10359) );
  OR2_X1 U10196 ( .A1(n8097), .A2(n8116), .ZN(n10166) );
  XOR2_X1 U10197 ( .A(n10362), .B(n10363), .Z(n10163) );
  XOR2_X1 U10198 ( .A(n10364), .B(n10365), .Z(n10363) );
  OR2_X1 U10199 ( .A1(n8093), .A2(n8116), .ZN(n10170) );
  XOR2_X1 U10200 ( .A(n10366), .B(n10367), .Z(n10167) );
  XOR2_X1 U10201 ( .A(n10368), .B(n10369), .Z(n10367) );
  OR2_X1 U10202 ( .A1(n8088), .A2(n8116), .ZN(n10174) );
  XOR2_X1 U10203 ( .A(n10370), .B(n10371), .Z(n10171) );
  XOR2_X1 U10204 ( .A(n10372), .B(n10373), .Z(n10371) );
  OR2_X1 U10205 ( .A1(n8084), .A2(n8116), .ZN(n10178) );
  XOR2_X1 U10206 ( .A(n10374), .B(n10375), .Z(n10175) );
  XOR2_X1 U10207 ( .A(n10376), .B(n10377), .Z(n10375) );
  OR2_X1 U10208 ( .A1(n8079), .A2(n8116), .ZN(n10182) );
  XOR2_X1 U10209 ( .A(n10378), .B(n10379), .Z(n10179) );
  XOR2_X1 U10210 ( .A(n10380), .B(n10381), .Z(n10379) );
  OR2_X1 U10211 ( .A1(n8075), .A2(n8116), .ZN(n10186) );
  XOR2_X1 U10212 ( .A(n10382), .B(n10383), .Z(n10183) );
  XOR2_X1 U10213 ( .A(n10384), .B(n10385), .Z(n10383) );
  OR2_X1 U10214 ( .A1(n8070), .A2(n8116), .ZN(n10190) );
  XOR2_X1 U10215 ( .A(n10386), .B(n10387), .Z(n10187) );
  XOR2_X1 U10216 ( .A(n10388), .B(n10389), .Z(n10387) );
  OR2_X1 U10217 ( .A1(n8066), .A2(n8116), .ZN(n10194) );
  XOR2_X1 U10218 ( .A(n10390), .B(n10391), .Z(n10191) );
  XOR2_X1 U10219 ( .A(n10392), .B(n10393), .Z(n10391) );
  OR2_X1 U10220 ( .A1(n8061), .A2(n8116), .ZN(n10198) );
  XOR2_X1 U10221 ( .A(n10394), .B(n10395), .Z(n10195) );
  XOR2_X1 U10222 ( .A(n10396), .B(n10397), .Z(n10395) );
  OR2_X1 U10223 ( .A1(n8057), .A2(n8116), .ZN(n10202) );
  XOR2_X1 U10224 ( .A(n10398), .B(n10399), .Z(n10199) );
  XOR2_X1 U10225 ( .A(n10400), .B(n10401), .Z(n10399) );
  XOR2_X1 U10226 ( .A(n10402), .B(n10403), .Z(n10204) );
  XOR2_X1 U10227 ( .A(n10404), .B(n10405), .Z(n10403) );
  OR2_X1 U10228 ( .A1(n8048), .A2(n8116), .ZN(n10210) );
  XNOR2_X1 U10229 ( .A(n10406), .B(n10407), .ZN(n10207) );
  XNOR2_X1 U10230 ( .A(n10408), .B(n10409), .ZN(n10406) );
  OR2_X1 U10231 ( .A1(n8043), .A2(n8116), .ZN(n10214) );
  XOR2_X1 U10232 ( .A(n10410), .B(n10411), .Z(n10211) );
  XOR2_X1 U10233 ( .A(n10412), .B(n10413), .Z(n10411) );
  OR2_X1 U10234 ( .A1(n8039), .A2(n8116), .ZN(n10218) );
  XOR2_X1 U10235 ( .A(n10414), .B(n10415), .Z(n10215) );
  XOR2_X1 U10236 ( .A(n10416), .B(n10417), .Z(n10415) );
  XOR2_X1 U10237 ( .A(n10418), .B(n10419), .Z(n10220) );
  XOR2_X1 U10238 ( .A(n10420), .B(n10421), .Z(n10419) );
  OR2_X1 U10239 ( .A1(n8030), .A2(n8116), .ZN(n10226) );
  XNOR2_X1 U10240 ( .A(n10422), .B(n10423), .ZN(n10223) );
  XNOR2_X1 U10241 ( .A(n10424), .B(n10425), .ZN(n10422) );
  OR2_X1 U10242 ( .A1(n8025), .A2(n8116), .ZN(n10230) );
  XOR2_X1 U10243 ( .A(n10426), .B(n10427), .Z(n10227) );
  XOR2_X1 U10244 ( .A(n10428), .B(n10429), .Z(n10427) );
  OR2_X1 U10245 ( .A1(n8021), .A2(n8116), .ZN(n10234) );
  XOR2_X1 U10246 ( .A(n10430), .B(n10431), .Z(n10231) );
  XOR2_X1 U10247 ( .A(n10432), .B(n10433), .Z(n10431) );
  OR2_X1 U10248 ( .A1(n8016), .A2(n8116), .ZN(n10238) );
  INV_X1 U10249 ( .A(b_25_), .ZN(n8116) );
  XNOR2_X1 U10250 ( .A(n10434), .B(n10435), .ZN(n10235) );
  XNOR2_X1 U10251 ( .A(n10436), .B(n10437), .ZN(n10434) );
  XOR2_X1 U10252 ( .A(n10028), .B(n10438), .Z(n10010) );
  XOR2_X1 U10253 ( .A(n10027), .B(n10026), .Z(n10438) );
  OR2_X1 U10254 ( .A1(n8113), .A2(n8016), .ZN(n10026) );
  OR2_X1 U10255 ( .A1(n10439), .A2(n10440), .ZN(n10027) );
  AND2_X1 U10256 ( .A1(n10437), .A2(n10436), .ZN(n10440) );
  AND2_X1 U10257 ( .A1(n10435), .A2(n10441), .ZN(n10439) );
  OR2_X1 U10258 ( .A1(n10437), .A2(n10436), .ZN(n10441) );
  OR2_X1 U10259 ( .A1(n8021), .A2(n8113), .ZN(n10436) );
  OR2_X1 U10260 ( .A1(n10442), .A2(n10443), .ZN(n10437) );
  AND2_X1 U10261 ( .A1(n10433), .A2(n10432), .ZN(n10443) );
  AND2_X1 U10262 ( .A1(n10430), .A2(n10444), .ZN(n10442) );
  OR2_X1 U10263 ( .A1(n10433), .A2(n10432), .ZN(n10444) );
  OR2_X1 U10264 ( .A1(n10445), .A2(n10446), .ZN(n10432) );
  AND2_X1 U10265 ( .A1(n10429), .A2(n10428), .ZN(n10446) );
  AND2_X1 U10266 ( .A1(n10426), .A2(n10447), .ZN(n10445) );
  OR2_X1 U10267 ( .A1(n10429), .A2(n10428), .ZN(n10447) );
  OR2_X1 U10268 ( .A1(n10448), .A2(n10449), .ZN(n10428) );
  AND2_X1 U10269 ( .A1(n10425), .A2(n10424), .ZN(n10449) );
  AND2_X1 U10270 ( .A1(n10423), .A2(n10450), .ZN(n10448) );
  OR2_X1 U10271 ( .A1(n10425), .A2(n10424), .ZN(n10450) );
  OR2_X1 U10272 ( .A1(n8113), .A2(n8034), .ZN(n10424) );
  OR2_X1 U10273 ( .A1(n10451), .A2(n10452), .ZN(n10425) );
  AND2_X1 U10274 ( .A1(n10421), .A2(n10420), .ZN(n10452) );
  AND2_X1 U10275 ( .A1(n10418), .A2(n10453), .ZN(n10451) );
  OR2_X1 U10276 ( .A1(n10421), .A2(n10420), .ZN(n10453) );
  OR2_X1 U10277 ( .A1(n10454), .A2(n10455), .ZN(n10420) );
  AND2_X1 U10278 ( .A1(n10417), .A2(n10416), .ZN(n10455) );
  AND2_X1 U10279 ( .A1(n10414), .A2(n10456), .ZN(n10454) );
  OR2_X1 U10280 ( .A1(n10417), .A2(n10416), .ZN(n10456) );
  OR2_X1 U10281 ( .A1(n10457), .A2(n10458), .ZN(n10416) );
  AND2_X1 U10282 ( .A1(n10413), .A2(n10412), .ZN(n10458) );
  AND2_X1 U10283 ( .A1(n10410), .A2(n10459), .ZN(n10457) );
  OR2_X1 U10284 ( .A1(n10413), .A2(n10412), .ZN(n10459) );
  OR2_X1 U10285 ( .A1(n10460), .A2(n10461), .ZN(n10412) );
  AND2_X1 U10286 ( .A1(n10409), .A2(n10408), .ZN(n10461) );
  AND2_X1 U10287 ( .A1(n10407), .A2(n10462), .ZN(n10460) );
  OR2_X1 U10288 ( .A1(n10409), .A2(n10408), .ZN(n10462) );
  OR2_X1 U10289 ( .A1(n8113), .A2(n8052), .ZN(n10408) );
  OR2_X1 U10290 ( .A1(n10463), .A2(n10464), .ZN(n10409) );
  AND2_X1 U10291 ( .A1(n10405), .A2(n10404), .ZN(n10464) );
  AND2_X1 U10292 ( .A1(n10402), .A2(n10465), .ZN(n10463) );
  OR2_X1 U10293 ( .A1(n10405), .A2(n10404), .ZN(n10465) );
  OR2_X1 U10294 ( .A1(n10466), .A2(n10467), .ZN(n10404) );
  AND2_X1 U10295 ( .A1(n10401), .A2(n10400), .ZN(n10467) );
  AND2_X1 U10296 ( .A1(n10398), .A2(n10468), .ZN(n10466) );
  OR2_X1 U10297 ( .A1(n10401), .A2(n10400), .ZN(n10468) );
  OR2_X1 U10298 ( .A1(n10469), .A2(n10470), .ZN(n10400) );
  AND2_X1 U10299 ( .A1(n10397), .A2(n10396), .ZN(n10470) );
  AND2_X1 U10300 ( .A1(n10394), .A2(n10471), .ZN(n10469) );
  OR2_X1 U10301 ( .A1(n10397), .A2(n10396), .ZN(n10471) );
  OR2_X1 U10302 ( .A1(n10472), .A2(n10473), .ZN(n10396) );
  AND2_X1 U10303 ( .A1(n10393), .A2(n10392), .ZN(n10473) );
  AND2_X1 U10304 ( .A1(n10390), .A2(n10474), .ZN(n10472) );
  OR2_X1 U10305 ( .A1(n10393), .A2(n10392), .ZN(n10474) );
  OR2_X1 U10306 ( .A1(n10475), .A2(n10476), .ZN(n10392) );
  AND2_X1 U10307 ( .A1(n10389), .A2(n10388), .ZN(n10476) );
  AND2_X1 U10308 ( .A1(n10386), .A2(n10477), .ZN(n10475) );
  OR2_X1 U10309 ( .A1(n10389), .A2(n10388), .ZN(n10477) );
  OR2_X1 U10310 ( .A1(n10478), .A2(n10479), .ZN(n10388) );
  AND2_X1 U10311 ( .A1(n10385), .A2(n10384), .ZN(n10479) );
  AND2_X1 U10312 ( .A1(n10382), .A2(n10480), .ZN(n10478) );
  OR2_X1 U10313 ( .A1(n10385), .A2(n10384), .ZN(n10480) );
  OR2_X1 U10314 ( .A1(n10481), .A2(n10482), .ZN(n10384) );
  AND2_X1 U10315 ( .A1(n10381), .A2(n10380), .ZN(n10482) );
  AND2_X1 U10316 ( .A1(n10378), .A2(n10483), .ZN(n10481) );
  OR2_X1 U10317 ( .A1(n10381), .A2(n10380), .ZN(n10483) );
  OR2_X1 U10318 ( .A1(n10484), .A2(n10485), .ZN(n10380) );
  AND2_X1 U10319 ( .A1(n10377), .A2(n10376), .ZN(n10485) );
  AND2_X1 U10320 ( .A1(n10374), .A2(n10486), .ZN(n10484) );
  OR2_X1 U10321 ( .A1(n10377), .A2(n10376), .ZN(n10486) );
  OR2_X1 U10322 ( .A1(n10487), .A2(n10488), .ZN(n10376) );
  AND2_X1 U10323 ( .A1(n10373), .A2(n10372), .ZN(n10488) );
  AND2_X1 U10324 ( .A1(n10370), .A2(n10489), .ZN(n10487) );
  OR2_X1 U10325 ( .A1(n10373), .A2(n10372), .ZN(n10489) );
  OR2_X1 U10326 ( .A1(n10490), .A2(n10491), .ZN(n10372) );
  AND2_X1 U10327 ( .A1(n10369), .A2(n10368), .ZN(n10491) );
  AND2_X1 U10328 ( .A1(n10366), .A2(n10492), .ZN(n10490) );
  OR2_X1 U10329 ( .A1(n10369), .A2(n10368), .ZN(n10492) );
  OR2_X1 U10330 ( .A1(n10493), .A2(n10494), .ZN(n10368) );
  AND2_X1 U10331 ( .A1(n10365), .A2(n10364), .ZN(n10494) );
  AND2_X1 U10332 ( .A1(n10362), .A2(n10495), .ZN(n10493) );
  OR2_X1 U10333 ( .A1(n10365), .A2(n10364), .ZN(n10495) );
  OR2_X1 U10334 ( .A1(n10496), .A2(n10497), .ZN(n10364) );
  AND2_X1 U10335 ( .A1(n10361), .A2(n10360), .ZN(n10497) );
  AND2_X1 U10336 ( .A1(n10358), .A2(n10498), .ZN(n10496) );
  OR2_X1 U10337 ( .A1(n10361), .A2(n10360), .ZN(n10498) );
  OR2_X1 U10338 ( .A1(n10499), .A2(n10500), .ZN(n10360) );
  AND2_X1 U10339 ( .A1(n10357), .A2(n10356), .ZN(n10500) );
  AND2_X1 U10340 ( .A1(n10354), .A2(n10501), .ZN(n10499) );
  OR2_X1 U10341 ( .A1(n10357), .A2(n10356), .ZN(n10501) );
  OR2_X1 U10342 ( .A1(n10502), .A2(n10503), .ZN(n10356) );
  AND2_X1 U10343 ( .A1(n7704), .A2(n10353), .ZN(n10503) );
  AND2_X1 U10344 ( .A1(n10351), .A2(n10504), .ZN(n10502) );
  OR2_X1 U10345 ( .A1(n7704), .A2(n10353), .ZN(n10504) );
  OR2_X1 U10346 ( .A1(n10505), .A2(n10506), .ZN(n10353) );
  AND2_X1 U10347 ( .A1(n10350), .A2(n10349), .ZN(n10506) );
  AND2_X1 U10348 ( .A1(n10347), .A2(n10507), .ZN(n10505) );
  OR2_X1 U10349 ( .A1(n10350), .A2(n10349), .ZN(n10507) );
  OR2_X1 U10350 ( .A1(n10508), .A2(n10509), .ZN(n10349) );
  AND2_X1 U10351 ( .A1(n10346), .A2(n10345), .ZN(n10509) );
  AND2_X1 U10352 ( .A1(n10343), .A2(n10510), .ZN(n10508) );
  OR2_X1 U10353 ( .A1(n10346), .A2(n10345), .ZN(n10510) );
  OR2_X1 U10354 ( .A1(n10511), .A2(n10512), .ZN(n10345) );
  AND2_X1 U10355 ( .A1(n10342), .A2(n10341), .ZN(n10512) );
  AND2_X1 U10356 ( .A1(n10339), .A2(n10513), .ZN(n10511) );
  OR2_X1 U10357 ( .A1(n10342), .A2(n10341), .ZN(n10513) );
  OR2_X1 U10358 ( .A1(n10514), .A2(n10515), .ZN(n10341) );
  AND2_X1 U10359 ( .A1(n10338), .A2(n10337), .ZN(n10515) );
  AND2_X1 U10360 ( .A1(n10335), .A2(n10516), .ZN(n10514) );
  OR2_X1 U10361 ( .A1(n10338), .A2(n10337), .ZN(n10516) );
  OR2_X1 U10362 ( .A1(n10517), .A2(n10518), .ZN(n10337) );
  AND2_X1 U10363 ( .A1(n10331), .A2(n10334), .ZN(n10518) );
  AND2_X1 U10364 ( .A1(n10519), .A2(n10520), .ZN(n10517) );
  OR2_X1 U10365 ( .A1(n10331), .A2(n10334), .ZN(n10520) );
  OR3_X1 U10366 ( .A1(n8981), .A2(n8113), .A3(n8110), .ZN(n10334) );
  OR2_X1 U10367 ( .A1(n8127), .A2(n8113), .ZN(n10331) );
  INV_X1 U10368 ( .A(n10333), .ZN(n10519) );
  OR2_X1 U10369 ( .A1(n10521), .A2(n10522), .ZN(n10333) );
  AND2_X1 U10370 ( .A1(b_23_), .A2(n10523), .ZN(n10522) );
  OR2_X1 U10371 ( .A1(n10524), .A2(n7598), .ZN(n10523) );
  AND2_X1 U10372 ( .A1(a_30_), .A2(n8107), .ZN(n10524) );
  AND2_X1 U10373 ( .A1(b_22_), .A2(n10525), .ZN(n10521) );
  OR2_X1 U10374 ( .A1(n10526), .A2(n7601), .ZN(n10525) );
  AND2_X1 U10375 ( .A1(a_31_), .A2(n8110), .ZN(n10526) );
  OR2_X1 U10376 ( .A1(n8124), .A2(n8113), .ZN(n10338) );
  XNOR2_X1 U10377 ( .A(n10527), .B(n10528), .ZN(n10335) );
  XOR2_X1 U10378 ( .A(n10529), .B(n10530), .Z(n10528) );
  OR2_X1 U10379 ( .A1(n8121), .A2(n8113), .ZN(n10342) );
  XOR2_X1 U10380 ( .A(n10531), .B(n10532), .Z(n10339) );
  XOR2_X1 U10381 ( .A(n10533), .B(n10534), .Z(n10532) );
  OR2_X1 U10382 ( .A1(n8118), .A2(n8113), .ZN(n10346) );
  XOR2_X1 U10383 ( .A(n10535), .B(n10536), .Z(n10343) );
  XOR2_X1 U10384 ( .A(n10537), .B(n10538), .Z(n10536) );
  OR2_X1 U10385 ( .A1(n8115), .A2(n8113), .ZN(n10350) );
  XOR2_X1 U10386 ( .A(n10539), .B(n10540), .Z(n10347) );
  XOR2_X1 U10387 ( .A(n10541), .B(n10542), .Z(n10540) );
  OR2_X1 U10388 ( .A1(n8112), .A2(n8113), .ZN(n7704) );
  XOR2_X1 U10389 ( .A(n10543), .B(n10544), .Z(n10351) );
  XOR2_X1 U10390 ( .A(n10545), .B(n10546), .Z(n10544) );
  OR2_X1 U10391 ( .A1(n8113), .A2(n8109), .ZN(n10357) );
  XOR2_X1 U10392 ( .A(n10547), .B(n10548), .Z(n10354) );
  XOR2_X1 U10393 ( .A(n10549), .B(n10550), .Z(n10548) );
  OR2_X1 U10394 ( .A1(n8113), .A2(n8106), .ZN(n10361) );
  XOR2_X1 U10395 ( .A(n10551), .B(n10552), .Z(n10358) );
  XOR2_X1 U10396 ( .A(n10553), .B(n7716), .Z(n10552) );
  OR2_X1 U10397 ( .A1(n8102), .A2(n8113), .ZN(n10365) );
  XOR2_X1 U10398 ( .A(n10554), .B(n10555), .Z(n10362) );
  XOR2_X1 U10399 ( .A(n10556), .B(n10557), .Z(n10555) );
  OR2_X1 U10400 ( .A1(n8113), .A2(n8097), .ZN(n10369) );
  XOR2_X1 U10401 ( .A(n10558), .B(n10559), .Z(n10366) );
  XOR2_X1 U10402 ( .A(n10560), .B(n10561), .Z(n10559) );
  OR2_X1 U10403 ( .A1(n8093), .A2(n8113), .ZN(n10373) );
  XOR2_X1 U10404 ( .A(n10562), .B(n10563), .Z(n10370) );
  XOR2_X1 U10405 ( .A(n10564), .B(n10565), .Z(n10563) );
  OR2_X1 U10406 ( .A1(n8113), .A2(n8088), .ZN(n10377) );
  XOR2_X1 U10407 ( .A(n10566), .B(n10567), .Z(n10374) );
  XOR2_X1 U10408 ( .A(n10568), .B(n10569), .Z(n10567) );
  OR2_X1 U10409 ( .A1(n8084), .A2(n8113), .ZN(n10381) );
  XOR2_X1 U10410 ( .A(n10570), .B(n10571), .Z(n10378) );
  XOR2_X1 U10411 ( .A(n10572), .B(n10573), .Z(n10571) );
  OR2_X1 U10412 ( .A1(n8113), .A2(n8079), .ZN(n10385) );
  XOR2_X1 U10413 ( .A(n10574), .B(n10575), .Z(n10382) );
  XOR2_X1 U10414 ( .A(n10576), .B(n10577), .Z(n10575) );
  OR2_X1 U10415 ( .A1(n8075), .A2(n8113), .ZN(n10389) );
  XOR2_X1 U10416 ( .A(n10578), .B(n10579), .Z(n10386) );
  XOR2_X1 U10417 ( .A(n10580), .B(n10581), .Z(n10579) );
  OR2_X1 U10418 ( .A1(n8113), .A2(n8070), .ZN(n10393) );
  XOR2_X1 U10419 ( .A(n10582), .B(n10583), .Z(n10390) );
  XOR2_X1 U10420 ( .A(n10584), .B(n10585), .Z(n10583) );
  OR2_X1 U10421 ( .A1(n8066), .A2(n8113), .ZN(n10397) );
  XNOR2_X1 U10422 ( .A(n10586), .B(n10587), .ZN(n10394) );
  XNOR2_X1 U10423 ( .A(n10588), .B(n10589), .ZN(n10586) );
  OR2_X1 U10424 ( .A1(n8113), .A2(n8061), .ZN(n10401) );
  XOR2_X1 U10425 ( .A(n10590), .B(n10591), .Z(n10398) );
  XOR2_X1 U10426 ( .A(n10592), .B(n10593), .Z(n10591) );
  OR2_X1 U10427 ( .A1(n8057), .A2(n8113), .ZN(n10405) );
  XOR2_X1 U10428 ( .A(n10594), .B(n10595), .Z(n10402) );
  XOR2_X1 U10429 ( .A(n10596), .B(n10597), .Z(n10595) );
  XOR2_X1 U10430 ( .A(n10598), .B(n10599), .Z(n10407) );
  XOR2_X1 U10431 ( .A(n10600), .B(n10601), .Z(n10599) );
  OR2_X1 U10432 ( .A1(n8048), .A2(n8113), .ZN(n10413) );
  XNOR2_X1 U10433 ( .A(n10602), .B(n10603), .ZN(n10410) );
  XNOR2_X1 U10434 ( .A(n10604), .B(n10605), .ZN(n10602) );
  OR2_X1 U10435 ( .A1(n8113), .A2(n8043), .ZN(n10417) );
  XOR2_X1 U10436 ( .A(n10606), .B(n10607), .Z(n10414) );
  XOR2_X1 U10437 ( .A(n10608), .B(n10609), .Z(n10607) );
  OR2_X1 U10438 ( .A1(n8039), .A2(n8113), .ZN(n10421) );
  XOR2_X1 U10439 ( .A(n10610), .B(n10611), .Z(n10418) );
  XOR2_X1 U10440 ( .A(n10612), .B(n10613), .Z(n10611) );
  XOR2_X1 U10441 ( .A(n10614), .B(n10615), .Z(n10423) );
  XOR2_X1 U10442 ( .A(n10616), .B(n10617), .Z(n10615) );
  OR2_X1 U10443 ( .A1(n8030), .A2(n8113), .ZN(n10429) );
  XNOR2_X1 U10444 ( .A(n10618), .B(n10619), .ZN(n10426) );
  XNOR2_X1 U10445 ( .A(n10620), .B(n10621), .ZN(n10618) );
  OR2_X1 U10446 ( .A1(n8113), .A2(n8025), .ZN(n10433) );
  INV_X1 U10447 ( .A(b_24_), .ZN(n8113) );
  XOR2_X1 U10448 ( .A(n10622), .B(n10623), .Z(n10430) );
  XOR2_X1 U10449 ( .A(n10624), .B(n10625), .Z(n10623) );
  XOR2_X1 U10450 ( .A(n10626), .B(n10627), .Z(n10435) );
  XOR2_X1 U10451 ( .A(n10628), .B(n10629), .Z(n10627) );
  XOR2_X1 U10452 ( .A(n10018), .B(n10630), .Z(n10028) );
  XOR2_X1 U10453 ( .A(n10017), .B(n10016), .Z(n10630) );
  OR2_X1 U10454 ( .A1(n8021), .A2(n8110), .ZN(n10016) );
  OR2_X1 U10455 ( .A1(n10631), .A2(n10632), .ZN(n10017) );
  AND2_X1 U10456 ( .A1(n10629), .A2(n10628), .ZN(n10632) );
  AND2_X1 U10457 ( .A1(n10626), .A2(n10633), .ZN(n10631) );
  OR2_X1 U10458 ( .A1(n10629), .A2(n10628), .ZN(n10633) );
  OR2_X1 U10459 ( .A1(n10634), .A2(n10635), .ZN(n10628) );
  AND2_X1 U10460 ( .A1(n10625), .A2(n10624), .ZN(n10635) );
  AND2_X1 U10461 ( .A1(n10622), .A2(n10636), .ZN(n10634) );
  OR2_X1 U10462 ( .A1(n10625), .A2(n10624), .ZN(n10636) );
  OR2_X1 U10463 ( .A1(n10637), .A2(n10638), .ZN(n10624) );
  AND2_X1 U10464 ( .A1(n10621), .A2(n10620), .ZN(n10638) );
  AND2_X1 U10465 ( .A1(n10619), .A2(n10639), .ZN(n10637) );
  OR2_X1 U10466 ( .A1(n10621), .A2(n10620), .ZN(n10639) );
  OR2_X1 U10467 ( .A1(n8034), .A2(n8110), .ZN(n10620) );
  OR2_X1 U10468 ( .A1(n10640), .A2(n10641), .ZN(n10621) );
  AND2_X1 U10469 ( .A1(n10617), .A2(n10616), .ZN(n10641) );
  AND2_X1 U10470 ( .A1(n10614), .A2(n10642), .ZN(n10640) );
  OR2_X1 U10471 ( .A1(n10617), .A2(n10616), .ZN(n10642) );
  OR2_X1 U10472 ( .A1(n10643), .A2(n10644), .ZN(n10616) );
  AND2_X1 U10473 ( .A1(n10613), .A2(n10612), .ZN(n10644) );
  AND2_X1 U10474 ( .A1(n10610), .A2(n10645), .ZN(n10643) );
  OR2_X1 U10475 ( .A1(n10613), .A2(n10612), .ZN(n10645) );
  OR2_X1 U10476 ( .A1(n10646), .A2(n10647), .ZN(n10612) );
  AND2_X1 U10477 ( .A1(n10609), .A2(n10608), .ZN(n10647) );
  AND2_X1 U10478 ( .A1(n10606), .A2(n10648), .ZN(n10646) );
  OR2_X1 U10479 ( .A1(n10609), .A2(n10608), .ZN(n10648) );
  OR2_X1 U10480 ( .A1(n10649), .A2(n10650), .ZN(n10608) );
  AND2_X1 U10481 ( .A1(n10605), .A2(n10604), .ZN(n10650) );
  AND2_X1 U10482 ( .A1(n10603), .A2(n10651), .ZN(n10649) );
  OR2_X1 U10483 ( .A1(n10605), .A2(n10604), .ZN(n10651) );
  OR2_X1 U10484 ( .A1(n8052), .A2(n8110), .ZN(n10604) );
  OR2_X1 U10485 ( .A1(n10652), .A2(n10653), .ZN(n10605) );
  AND2_X1 U10486 ( .A1(n10601), .A2(n10600), .ZN(n10653) );
  AND2_X1 U10487 ( .A1(n10598), .A2(n10654), .ZN(n10652) );
  OR2_X1 U10488 ( .A1(n10601), .A2(n10600), .ZN(n10654) );
  OR2_X1 U10489 ( .A1(n10655), .A2(n10656), .ZN(n10600) );
  AND2_X1 U10490 ( .A1(n10597), .A2(n10596), .ZN(n10656) );
  AND2_X1 U10491 ( .A1(n10594), .A2(n10657), .ZN(n10655) );
  OR2_X1 U10492 ( .A1(n10597), .A2(n10596), .ZN(n10657) );
  OR2_X1 U10493 ( .A1(n10658), .A2(n10659), .ZN(n10596) );
  AND2_X1 U10494 ( .A1(n10593), .A2(n10592), .ZN(n10659) );
  AND2_X1 U10495 ( .A1(n10590), .A2(n10660), .ZN(n10658) );
  OR2_X1 U10496 ( .A1(n10593), .A2(n10592), .ZN(n10660) );
  OR2_X1 U10497 ( .A1(n10661), .A2(n10662), .ZN(n10592) );
  AND2_X1 U10498 ( .A1(n10589), .A2(n10588), .ZN(n10662) );
  AND2_X1 U10499 ( .A1(n10587), .A2(n10663), .ZN(n10661) );
  OR2_X1 U10500 ( .A1(n10589), .A2(n10588), .ZN(n10663) );
  OR2_X1 U10501 ( .A1(n8070), .A2(n8110), .ZN(n10588) );
  OR2_X1 U10502 ( .A1(n10664), .A2(n10665), .ZN(n10589) );
  AND2_X1 U10503 ( .A1(n10585), .A2(n10584), .ZN(n10665) );
  AND2_X1 U10504 ( .A1(n10582), .A2(n10666), .ZN(n10664) );
  OR2_X1 U10505 ( .A1(n10585), .A2(n10584), .ZN(n10666) );
  OR2_X1 U10506 ( .A1(n10667), .A2(n10668), .ZN(n10584) );
  AND2_X1 U10507 ( .A1(n10581), .A2(n10580), .ZN(n10668) );
  AND2_X1 U10508 ( .A1(n10578), .A2(n10669), .ZN(n10667) );
  OR2_X1 U10509 ( .A1(n10581), .A2(n10580), .ZN(n10669) );
  OR2_X1 U10510 ( .A1(n10670), .A2(n10671), .ZN(n10580) );
  AND2_X1 U10511 ( .A1(n10577), .A2(n10576), .ZN(n10671) );
  AND2_X1 U10512 ( .A1(n10574), .A2(n10672), .ZN(n10670) );
  OR2_X1 U10513 ( .A1(n10577), .A2(n10576), .ZN(n10672) );
  OR2_X1 U10514 ( .A1(n10673), .A2(n10674), .ZN(n10576) );
  AND2_X1 U10515 ( .A1(n10573), .A2(n10572), .ZN(n10674) );
  AND2_X1 U10516 ( .A1(n10570), .A2(n10675), .ZN(n10673) );
  OR2_X1 U10517 ( .A1(n10573), .A2(n10572), .ZN(n10675) );
  OR2_X1 U10518 ( .A1(n10676), .A2(n10677), .ZN(n10572) );
  AND2_X1 U10519 ( .A1(n10569), .A2(n10568), .ZN(n10677) );
  AND2_X1 U10520 ( .A1(n10566), .A2(n10678), .ZN(n10676) );
  OR2_X1 U10521 ( .A1(n10569), .A2(n10568), .ZN(n10678) );
  OR2_X1 U10522 ( .A1(n10679), .A2(n10680), .ZN(n10568) );
  AND2_X1 U10523 ( .A1(n10565), .A2(n10564), .ZN(n10680) );
  AND2_X1 U10524 ( .A1(n10562), .A2(n10681), .ZN(n10679) );
  OR2_X1 U10525 ( .A1(n10565), .A2(n10564), .ZN(n10681) );
  OR2_X1 U10526 ( .A1(n10682), .A2(n10683), .ZN(n10564) );
  AND2_X1 U10527 ( .A1(n10561), .A2(n10560), .ZN(n10683) );
  AND2_X1 U10528 ( .A1(n10558), .A2(n10684), .ZN(n10682) );
  OR2_X1 U10529 ( .A1(n10561), .A2(n10560), .ZN(n10684) );
  OR2_X1 U10530 ( .A1(n10685), .A2(n10686), .ZN(n10560) );
  AND2_X1 U10531 ( .A1(n10557), .A2(n10556), .ZN(n10686) );
  AND2_X1 U10532 ( .A1(n10554), .A2(n10687), .ZN(n10685) );
  OR2_X1 U10533 ( .A1(n10557), .A2(n10556), .ZN(n10687) );
  OR2_X1 U10534 ( .A1(n10688), .A2(n10689), .ZN(n10556) );
  AND2_X1 U10535 ( .A1(n7716), .A2(n10553), .ZN(n10689) );
  AND2_X1 U10536 ( .A1(n10551), .A2(n10690), .ZN(n10688) );
  OR2_X1 U10537 ( .A1(n7716), .A2(n10553), .ZN(n10690) );
  OR2_X1 U10538 ( .A1(n10691), .A2(n10692), .ZN(n10553) );
  AND2_X1 U10539 ( .A1(n10550), .A2(n10549), .ZN(n10692) );
  AND2_X1 U10540 ( .A1(n10547), .A2(n10693), .ZN(n10691) );
  OR2_X1 U10541 ( .A1(n10550), .A2(n10549), .ZN(n10693) );
  OR2_X1 U10542 ( .A1(n10694), .A2(n10695), .ZN(n10549) );
  AND2_X1 U10543 ( .A1(n10546), .A2(n10545), .ZN(n10695) );
  AND2_X1 U10544 ( .A1(n10543), .A2(n10696), .ZN(n10694) );
  OR2_X1 U10545 ( .A1(n10546), .A2(n10545), .ZN(n10696) );
  OR2_X1 U10546 ( .A1(n10697), .A2(n10698), .ZN(n10545) );
  AND2_X1 U10547 ( .A1(n10542), .A2(n10541), .ZN(n10698) );
  AND2_X1 U10548 ( .A1(n10539), .A2(n10699), .ZN(n10697) );
  OR2_X1 U10549 ( .A1(n10542), .A2(n10541), .ZN(n10699) );
  OR2_X1 U10550 ( .A1(n10700), .A2(n10701), .ZN(n10541) );
  AND2_X1 U10551 ( .A1(n10538), .A2(n10537), .ZN(n10701) );
  AND2_X1 U10552 ( .A1(n10535), .A2(n10702), .ZN(n10700) );
  OR2_X1 U10553 ( .A1(n10538), .A2(n10537), .ZN(n10702) );
  OR2_X1 U10554 ( .A1(n10703), .A2(n10704), .ZN(n10537) );
  AND2_X1 U10555 ( .A1(n10534), .A2(n10533), .ZN(n10704) );
  AND2_X1 U10556 ( .A1(n10531), .A2(n10705), .ZN(n10703) );
  OR2_X1 U10557 ( .A1(n10534), .A2(n10533), .ZN(n10705) );
  OR2_X1 U10558 ( .A1(n10706), .A2(n10707), .ZN(n10533) );
  AND2_X1 U10559 ( .A1(n10527), .A2(n10530), .ZN(n10707) );
  AND2_X1 U10560 ( .A1(n10708), .A2(n10709), .ZN(n10706) );
  OR2_X1 U10561 ( .A1(n10527), .A2(n10530), .ZN(n10709) );
  OR3_X1 U10562 ( .A1(n8981), .A2(n8107), .A3(n8110), .ZN(n10530) );
  OR2_X1 U10563 ( .A1(n8127), .A2(n8110), .ZN(n10527) );
  INV_X1 U10564 ( .A(n10529), .ZN(n10708) );
  OR2_X1 U10565 ( .A1(n10710), .A2(n10711), .ZN(n10529) );
  AND2_X1 U10566 ( .A1(b_22_), .A2(n10712), .ZN(n10711) );
  OR2_X1 U10567 ( .A1(n10713), .A2(n7598), .ZN(n10712) );
  AND2_X1 U10568 ( .A1(a_30_), .A2(n8103), .ZN(n10713) );
  AND2_X1 U10569 ( .A1(b_21_), .A2(n10714), .ZN(n10710) );
  OR2_X1 U10570 ( .A1(n10715), .A2(n7601), .ZN(n10714) );
  AND2_X1 U10571 ( .A1(a_31_), .A2(n8107), .ZN(n10715) );
  OR2_X1 U10572 ( .A1(n8124), .A2(n8110), .ZN(n10534) );
  XNOR2_X1 U10573 ( .A(n10716), .B(n10717), .ZN(n10531) );
  XOR2_X1 U10574 ( .A(n10718), .B(n10719), .Z(n10717) );
  OR2_X1 U10575 ( .A1(n8121), .A2(n8110), .ZN(n10538) );
  XOR2_X1 U10576 ( .A(n10720), .B(n10721), .Z(n10535) );
  XOR2_X1 U10577 ( .A(n10722), .B(n10723), .Z(n10721) );
  OR2_X1 U10578 ( .A1(n8118), .A2(n8110), .ZN(n10542) );
  XOR2_X1 U10579 ( .A(n10724), .B(n10725), .Z(n10539) );
  XOR2_X1 U10580 ( .A(n10726), .B(n10727), .Z(n10725) );
  OR2_X1 U10581 ( .A1(n8115), .A2(n8110), .ZN(n10546) );
  XOR2_X1 U10582 ( .A(n10728), .B(n10729), .Z(n10543) );
  XOR2_X1 U10583 ( .A(n10730), .B(n10731), .Z(n10729) );
  OR2_X1 U10584 ( .A1(n8112), .A2(n8110), .ZN(n10550) );
  XOR2_X1 U10585 ( .A(n10732), .B(n10733), .Z(n10547) );
  XOR2_X1 U10586 ( .A(n10734), .B(n10735), .Z(n10733) );
  OR2_X1 U10587 ( .A1(n8109), .A2(n8110), .ZN(n7716) );
  XOR2_X1 U10588 ( .A(n10736), .B(n10737), .Z(n10551) );
  XOR2_X1 U10589 ( .A(n10738), .B(n10739), .Z(n10737) );
  OR2_X1 U10590 ( .A1(n8106), .A2(n8110), .ZN(n10557) );
  XOR2_X1 U10591 ( .A(n10740), .B(n10741), .Z(n10554) );
  XOR2_X1 U10592 ( .A(n10742), .B(n10743), .Z(n10741) );
  OR2_X1 U10593 ( .A1(n8102), .A2(n8110), .ZN(n10561) );
  XOR2_X1 U10594 ( .A(n10744), .B(n10745), .Z(n10558) );
  XOR2_X1 U10595 ( .A(n10746), .B(n7734), .Z(n10745) );
  OR2_X1 U10596 ( .A1(n8097), .A2(n8110), .ZN(n10565) );
  XOR2_X1 U10597 ( .A(n10747), .B(n10748), .Z(n10562) );
  XOR2_X1 U10598 ( .A(n10749), .B(n10750), .Z(n10748) );
  OR2_X1 U10599 ( .A1(n8093), .A2(n8110), .ZN(n10569) );
  XOR2_X1 U10600 ( .A(n10751), .B(n10752), .Z(n10566) );
  XOR2_X1 U10601 ( .A(n10753), .B(n10754), .Z(n10752) );
  OR2_X1 U10602 ( .A1(n8088), .A2(n8110), .ZN(n10573) );
  XOR2_X1 U10603 ( .A(n10755), .B(n10756), .Z(n10570) );
  XOR2_X1 U10604 ( .A(n10757), .B(n10758), .Z(n10756) );
  OR2_X1 U10605 ( .A1(n8084), .A2(n8110), .ZN(n10577) );
  XOR2_X1 U10606 ( .A(n10759), .B(n10760), .Z(n10574) );
  XOR2_X1 U10607 ( .A(n10761), .B(n10762), .Z(n10760) );
  OR2_X1 U10608 ( .A1(n8079), .A2(n8110), .ZN(n10581) );
  XOR2_X1 U10609 ( .A(n10763), .B(n10764), .Z(n10578) );
  XOR2_X1 U10610 ( .A(n10765), .B(n10766), .Z(n10764) );
  OR2_X1 U10611 ( .A1(n8075), .A2(n8110), .ZN(n10585) );
  XOR2_X1 U10612 ( .A(n10767), .B(n10768), .Z(n10582) );
  XOR2_X1 U10613 ( .A(n10769), .B(n10770), .Z(n10768) );
  XOR2_X1 U10614 ( .A(n10771), .B(n10772), .Z(n10587) );
  XOR2_X1 U10615 ( .A(n10773), .B(n10774), .Z(n10772) );
  OR2_X1 U10616 ( .A1(n8066), .A2(n8110), .ZN(n10593) );
  XOR2_X1 U10617 ( .A(n10775), .B(n10776), .Z(n10590) );
  XOR2_X1 U10618 ( .A(n10777), .B(n10778), .Z(n10776) );
  OR2_X1 U10619 ( .A1(n8061), .A2(n8110), .ZN(n10597) );
  XOR2_X1 U10620 ( .A(n10779), .B(n10780), .Z(n10594) );
  XOR2_X1 U10621 ( .A(n10781), .B(n10782), .Z(n10780) );
  OR2_X1 U10622 ( .A1(n8057), .A2(n8110), .ZN(n10601) );
  XOR2_X1 U10623 ( .A(n10783), .B(n10784), .Z(n10598) );
  XOR2_X1 U10624 ( .A(n10785), .B(n10786), .Z(n10784) );
  XOR2_X1 U10625 ( .A(n10787), .B(n10788), .Z(n10603) );
  XOR2_X1 U10626 ( .A(n10789), .B(n10790), .Z(n10788) );
  OR2_X1 U10627 ( .A1(n8048), .A2(n8110), .ZN(n10609) );
  XOR2_X1 U10628 ( .A(n10791), .B(n10792), .Z(n10606) );
  XOR2_X1 U10629 ( .A(n10793), .B(n10794), .Z(n10792) );
  OR2_X1 U10630 ( .A1(n8043), .A2(n8110), .ZN(n10613) );
  XOR2_X1 U10631 ( .A(n10795), .B(n10796), .Z(n10610) );
  XOR2_X1 U10632 ( .A(n10797), .B(n10798), .Z(n10796) );
  OR2_X1 U10633 ( .A1(n8039), .A2(n8110), .ZN(n10617) );
  XOR2_X1 U10634 ( .A(n10799), .B(n10800), .Z(n10614) );
  XOR2_X1 U10635 ( .A(n10801), .B(n10802), .Z(n10800) );
  XOR2_X1 U10636 ( .A(n10803), .B(n10804), .Z(n10619) );
  XOR2_X1 U10637 ( .A(n10805), .B(n10806), .Z(n10804) );
  OR2_X1 U10638 ( .A1(n8030), .A2(n8110), .ZN(n10625) );
  XOR2_X1 U10639 ( .A(n10807), .B(n10808), .Z(n10622) );
  XOR2_X1 U10640 ( .A(n10809), .B(n10810), .Z(n10808) );
  OR2_X1 U10641 ( .A1(n8025), .A2(n8110), .ZN(n10629) );
  INV_X1 U10642 ( .A(b_23_), .ZN(n8110) );
  XOR2_X1 U10643 ( .A(n10811), .B(n10812), .Z(n10626) );
  XOR2_X1 U10644 ( .A(n10813), .B(n10814), .Z(n10812) );
  XOR2_X1 U10645 ( .A(n10815), .B(n10816), .Z(n10018) );
  XOR2_X1 U10646 ( .A(n10817), .B(n10818), .Z(n10816) );
  OR2_X1 U10647 ( .A1(n10819), .A2(n8813), .ZN(n8190) );
  XOR2_X1 U10648 ( .A(n8761), .B(n8763), .Z(n8813) );
  OR2_X1 U10649 ( .A1(n10820), .A2(n10821), .ZN(n8763) );
  AND2_X1 U10650 ( .A1(n10822), .A2(n10823), .ZN(n10821) );
  AND2_X1 U10651 ( .A1(n10824), .A2(n10825), .ZN(n10820) );
  OR2_X1 U10652 ( .A1(n10822), .A2(n10823), .ZN(n10825) );
  XOR2_X1 U10653 ( .A(n8770), .B(n10826), .Z(n8761) );
  XOR2_X1 U10654 ( .A(n8769), .B(n8768), .Z(n10826) );
  OR2_X1 U10655 ( .A1(n8098), .A2(n8297), .ZN(n8768) );
  OR2_X1 U10656 ( .A1(n10827), .A2(n10828), .ZN(n8769) );
  AND2_X1 U10657 ( .A1(n10829), .A2(n10830), .ZN(n10828) );
  AND2_X1 U10658 ( .A1(n10831), .A2(n10832), .ZN(n10827) );
  OR2_X1 U10659 ( .A1(n10829), .A2(n10830), .ZN(n10832) );
  XOR2_X1 U10660 ( .A(n8777), .B(n10833), .Z(n8770) );
  XOR2_X1 U10661 ( .A(n8776), .B(n8775), .Z(n10833) );
  OR2_X1 U10662 ( .A1(n8094), .A2(n8012), .ZN(n8775) );
  OR2_X1 U10663 ( .A1(n10834), .A2(n10835), .ZN(n8776) );
  AND2_X1 U10664 ( .A1(n10836), .A2(n10837), .ZN(n10835) );
  AND2_X1 U10665 ( .A1(n10838), .A2(n10839), .ZN(n10834) );
  OR2_X1 U10666 ( .A1(n10836), .A2(n10837), .ZN(n10839) );
  XOR2_X1 U10667 ( .A(n8784), .B(n10840), .Z(n8777) );
  XOR2_X1 U10668 ( .A(n8783), .B(n8782), .Z(n10840) );
  OR2_X1 U10669 ( .A1(n8089), .A2(n8016), .ZN(n8782) );
  OR2_X1 U10670 ( .A1(n10841), .A2(n10842), .ZN(n8783) );
  AND2_X1 U10671 ( .A1(n10843), .A2(n10844), .ZN(n10842) );
  AND2_X1 U10672 ( .A1(n10845), .A2(n10846), .ZN(n10841) );
  OR2_X1 U10673 ( .A1(n10843), .A2(n10844), .ZN(n10846) );
  XOR2_X1 U10674 ( .A(n8791), .B(n10847), .Z(n8784) );
  XOR2_X1 U10675 ( .A(n8790), .B(n8789), .Z(n10847) );
  OR2_X1 U10676 ( .A1(n8021), .A2(n8085), .ZN(n8789) );
  OR2_X1 U10677 ( .A1(n10848), .A2(n10849), .ZN(n8790) );
  AND2_X1 U10678 ( .A1(n10850), .A2(n10851), .ZN(n10849) );
  AND2_X1 U10679 ( .A1(n10852), .A2(n10853), .ZN(n10848) );
  OR2_X1 U10680 ( .A1(n10850), .A2(n10851), .ZN(n10853) );
  XOR2_X1 U10681 ( .A(n8798), .B(n10854), .Z(n8791) );
  XOR2_X1 U10682 ( .A(n8797), .B(n8796), .Z(n10854) );
  OR2_X1 U10683 ( .A1(n8080), .A2(n8025), .ZN(n8796) );
  OR2_X1 U10684 ( .A1(n10855), .A2(n10856), .ZN(n8797) );
  AND2_X1 U10685 ( .A1(n10857), .A2(n10858), .ZN(n10856) );
  AND2_X1 U10686 ( .A1(n10859), .A2(n10860), .ZN(n10855) );
  OR2_X1 U10687 ( .A1(n10857), .A2(n10858), .ZN(n10860) );
  XOR2_X1 U10688 ( .A(n8805), .B(n10861), .Z(n8798) );
  XOR2_X1 U10689 ( .A(n8804), .B(n8803), .Z(n10861) );
  OR2_X1 U10690 ( .A1(n8030), .A2(n8076), .ZN(n8803) );
  OR2_X1 U10691 ( .A1(n10862), .A2(n10863), .ZN(n8804) );
  AND2_X1 U10692 ( .A1(n10864), .A2(n10865), .ZN(n10863) );
  AND2_X1 U10693 ( .A1(n10866), .A2(n10867), .ZN(n10862) );
  OR2_X1 U10694 ( .A1(n10865), .A2(n10864), .ZN(n10867) );
  XOR2_X1 U10695 ( .A(n10868), .B(n10869), .Z(n8805) );
  XOR2_X1 U10696 ( .A(n10870), .B(n10871), .Z(n10869) );
  AND2_X1 U10697 ( .A1(n8814), .A2(n8812), .ZN(n10819) );
  XNOR2_X1 U10698 ( .A(n10824), .B(n10872), .ZN(n8812) );
  XOR2_X1 U10699 ( .A(n10823), .B(n10822), .Z(n10872) );
  OR2_X1 U10700 ( .A1(n8103), .A2(n8297), .ZN(n10822) );
  OR2_X1 U10701 ( .A1(n10873), .A2(n10874), .ZN(n10823) );
  AND2_X1 U10702 ( .A1(n10875), .A2(n10876), .ZN(n10874) );
  AND2_X1 U10703 ( .A1(n10877), .A2(n10878), .ZN(n10873) );
  OR2_X1 U10704 ( .A1(n10875), .A2(n10876), .ZN(n10878) );
  XOR2_X1 U10705 ( .A(n10831), .B(n10879), .Z(n10824) );
  XOR2_X1 U10706 ( .A(n10830), .B(n10829), .Z(n10879) );
  OR2_X1 U10707 ( .A1(n8098), .A2(n8012), .ZN(n10829) );
  OR2_X1 U10708 ( .A1(n10880), .A2(n10881), .ZN(n10830) );
  AND2_X1 U10709 ( .A1(n10882), .A2(n10883), .ZN(n10881) );
  AND2_X1 U10710 ( .A1(n10884), .A2(n10885), .ZN(n10880) );
  OR2_X1 U10711 ( .A1(n10882), .A2(n10883), .ZN(n10885) );
  XOR2_X1 U10712 ( .A(n10838), .B(n10886), .Z(n10831) );
  XOR2_X1 U10713 ( .A(n10837), .B(n10836), .Z(n10886) );
  OR2_X1 U10714 ( .A1(n8094), .A2(n8016), .ZN(n10836) );
  OR2_X1 U10715 ( .A1(n10887), .A2(n10888), .ZN(n10837) );
  AND2_X1 U10716 ( .A1(n10889), .A2(n10890), .ZN(n10888) );
  AND2_X1 U10717 ( .A1(n10891), .A2(n10892), .ZN(n10887) );
  OR2_X1 U10718 ( .A1(n10889), .A2(n10890), .ZN(n10892) );
  XOR2_X1 U10719 ( .A(n10845), .B(n10893), .Z(n10838) );
  XOR2_X1 U10720 ( .A(n10844), .B(n10843), .Z(n10893) );
  OR2_X1 U10721 ( .A1(n8021), .A2(n8089), .ZN(n10843) );
  OR2_X1 U10722 ( .A1(n10894), .A2(n10895), .ZN(n10844) );
  AND2_X1 U10723 ( .A1(n10896), .A2(n10897), .ZN(n10895) );
  AND2_X1 U10724 ( .A1(n10898), .A2(n10899), .ZN(n10894) );
  OR2_X1 U10725 ( .A1(n10896), .A2(n10897), .ZN(n10899) );
  XOR2_X1 U10726 ( .A(n10852), .B(n10900), .Z(n10845) );
  XOR2_X1 U10727 ( .A(n10851), .B(n10850), .Z(n10900) );
  OR2_X1 U10728 ( .A1(n8085), .A2(n8025), .ZN(n10850) );
  OR2_X1 U10729 ( .A1(n10901), .A2(n10902), .ZN(n10851) );
  AND2_X1 U10730 ( .A1(n10903), .A2(n10904), .ZN(n10902) );
  AND2_X1 U10731 ( .A1(n10905), .A2(n10906), .ZN(n10901) );
  OR2_X1 U10732 ( .A1(n10903), .A2(n10904), .ZN(n10906) );
  XOR2_X1 U10733 ( .A(n10859), .B(n10907), .Z(n10852) );
  XOR2_X1 U10734 ( .A(n10858), .B(n10857), .Z(n10907) );
  OR2_X1 U10735 ( .A1(n8030), .A2(n8080), .ZN(n10857) );
  OR2_X1 U10736 ( .A1(n10908), .A2(n10909), .ZN(n10858) );
  AND2_X1 U10737 ( .A1(n10910), .A2(n10911), .ZN(n10909) );
  AND2_X1 U10738 ( .A1(n10912), .A2(n10913), .ZN(n10908) );
  OR2_X1 U10739 ( .A1(n10910), .A2(n10911), .ZN(n10913) );
  XOR2_X1 U10740 ( .A(n10866), .B(n10914), .Z(n10859) );
  XOR2_X1 U10741 ( .A(n10865), .B(n10864), .Z(n10914) );
  OR2_X1 U10742 ( .A1(n8076), .A2(n8034), .ZN(n10864) );
  OR2_X1 U10743 ( .A1(n10915), .A2(n10916), .ZN(n10865) );
  AND2_X1 U10744 ( .A1(n10917), .A2(n10918), .ZN(n10916) );
  AND2_X1 U10745 ( .A1(n10919), .A2(n10920), .ZN(n10915) );
  OR2_X1 U10746 ( .A1(n10918), .A2(n10917), .ZN(n10920) );
  XOR2_X1 U10747 ( .A(n10921), .B(n10922), .Z(n10866) );
  XOR2_X1 U10748 ( .A(n10923), .B(n10924), .Z(n10922) );
  INV_X1 U10749 ( .A(n8822), .ZN(n8814) );
  OR2_X1 U10750 ( .A1(n10925), .A2(n10926), .ZN(n8822) );
  AND2_X1 U10751 ( .A1(n8839), .A2(n8838), .ZN(n10926) );
  AND2_X1 U10752 ( .A1(n8836), .A2(n10927), .ZN(n10925) );
  OR2_X1 U10753 ( .A1(n8838), .A2(n8839), .ZN(n10927) );
  OR2_X1 U10754 ( .A1(n8107), .A2(n8297), .ZN(n8839) );
  OR2_X1 U10755 ( .A1(n10928), .A2(n10929), .ZN(n8838) );
  AND2_X1 U10756 ( .A1(n8863), .A2(n8862), .ZN(n10929) );
  AND2_X1 U10757 ( .A1(n8860), .A2(n10930), .ZN(n10928) );
  OR2_X1 U10758 ( .A1(n8862), .A2(n8863), .ZN(n10930) );
  OR2_X1 U10759 ( .A1(n8107), .A2(n8012), .ZN(n8863) );
  OR2_X1 U10760 ( .A1(n10931), .A2(n10932), .ZN(n8862) );
  AND2_X1 U10761 ( .A1(n10004), .A2(n10003), .ZN(n10932) );
  AND2_X1 U10762 ( .A1(n10001), .A2(n10933), .ZN(n10931) );
  OR2_X1 U10763 ( .A1(n10003), .A2(n10004), .ZN(n10933) );
  OR2_X1 U10764 ( .A1(n8107), .A2(n8016), .ZN(n10004) );
  OR2_X1 U10765 ( .A1(n10934), .A2(n10935), .ZN(n10003) );
  AND2_X1 U10766 ( .A1(n10023), .A2(n10022), .ZN(n10935) );
  AND2_X1 U10767 ( .A1(n10020), .A2(n10936), .ZN(n10934) );
  OR2_X1 U10768 ( .A1(n10022), .A2(n10023), .ZN(n10936) );
  OR2_X1 U10769 ( .A1(n8021), .A2(n8107), .ZN(n10023) );
  OR2_X1 U10770 ( .A1(n10937), .A2(n10938), .ZN(n10022) );
  AND2_X1 U10771 ( .A1(n10818), .A2(n10817), .ZN(n10938) );
  AND2_X1 U10772 ( .A1(n10815), .A2(n10939), .ZN(n10937) );
  OR2_X1 U10773 ( .A1(n10817), .A2(n10818), .ZN(n10939) );
  OR2_X1 U10774 ( .A1(n8107), .A2(n8025), .ZN(n10818) );
  OR2_X1 U10775 ( .A1(n10940), .A2(n10941), .ZN(n10817) );
  AND2_X1 U10776 ( .A1(n10814), .A2(n10813), .ZN(n10941) );
  AND2_X1 U10777 ( .A1(n10811), .A2(n10942), .ZN(n10940) );
  OR2_X1 U10778 ( .A1(n10813), .A2(n10814), .ZN(n10942) );
  OR2_X1 U10779 ( .A1(n8030), .A2(n8107), .ZN(n10814) );
  OR2_X1 U10780 ( .A1(n10943), .A2(n10944), .ZN(n10813) );
  AND2_X1 U10781 ( .A1(n10810), .A2(n10809), .ZN(n10944) );
  AND2_X1 U10782 ( .A1(n10807), .A2(n10945), .ZN(n10943) );
  OR2_X1 U10783 ( .A1(n10809), .A2(n10810), .ZN(n10945) );
  OR2_X1 U10784 ( .A1(n8107), .A2(n8034), .ZN(n10810) );
  OR2_X1 U10785 ( .A1(n10946), .A2(n10947), .ZN(n10809) );
  AND2_X1 U10786 ( .A1(n10806), .A2(n10805), .ZN(n10947) );
  AND2_X1 U10787 ( .A1(n10803), .A2(n10948), .ZN(n10946) );
  OR2_X1 U10788 ( .A1(n10805), .A2(n10806), .ZN(n10948) );
  OR2_X1 U10789 ( .A1(n8039), .A2(n8107), .ZN(n10806) );
  OR2_X1 U10790 ( .A1(n10949), .A2(n10950), .ZN(n10805) );
  AND2_X1 U10791 ( .A1(n10802), .A2(n10801), .ZN(n10950) );
  AND2_X1 U10792 ( .A1(n10799), .A2(n10951), .ZN(n10949) );
  OR2_X1 U10793 ( .A1(n10801), .A2(n10802), .ZN(n10951) );
  OR2_X1 U10794 ( .A1(n8107), .A2(n8043), .ZN(n10802) );
  OR2_X1 U10795 ( .A1(n10952), .A2(n10953), .ZN(n10801) );
  AND2_X1 U10796 ( .A1(n10798), .A2(n10797), .ZN(n10953) );
  AND2_X1 U10797 ( .A1(n10795), .A2(n10954), .ZN(n10952) );
  OR2_X1 U10798 ( .A1(n10797), .A2(n10798), .ZN(n10954) );
  OR2_X1 U10799 ( .A1(n8048), .A2(n8107), .ZN(n10798) );
  OR2_X1 U10800 ( .A1(n10955), .A2(n10956), .ZN(n10797) );
  AND2_X1 U10801 ( .A1(n10794), .A2(n10793), .ZN(n10956) );
  AND2_X1 U10802 ( .A1(n10791), .A2(n10957), .ZN(n10955) );
  OR2_X1 U10803 ( .A1(n10793), .A2(n10794), .ZN(n10957) );
  OR2_X1 U10804 ( .A1(n8107), .A2(n8052), .ZN(n10794) );
  OR2_X1 U10805 ( .A1(n10958), .A2(n10959), .ZN(n10793) );
  AND2_X1 U10806 ( .A1(n10790), .A2(n10789), .ZN(n10959) );
  AND2_X1 U10807 ( .A1(n10787), .A2(n10960), .ZN(n10958) );
  OR2_X1 U10808 ( .A1(n10789), .A2(n10790), .ZN(n10960) );
  OR2_X1 U10809 ( .A1(n8057), .A2(n8107), .ZN(n10790) );
  OR2_X1 U10810 ( .A1(n10961), .A2(n10962), .ZN(n10789) );
  AND2_X1 U10811 ( .A1(n10786), .A2(n10785), .ZN(n10962) );
  AND2_X1 U10812 ( .A1(n10783), .A2(n10963), .ZN(n10961) );
  OR2_X1 U10813 ( .A1(n10785), .A2(n10786), .ZN(n10963) );
  OR2_X1 U10814 ( .A1(n8107), .A2(n8061), .ZN(n10786) );
  OR2_X1 U10815 ( .A1(n10964), .A2(n10965), .ZN(n10785) );
  AND2_X1 U10816 ( .A1(n10782), .A2(n10781), .ZN(n10965) );
  AND2_X1 U10817 ( .A1(n10779), .A2(n10966), .ZN(n10964) );
  OR2_X1 U10818 ( .A1(n10781), .A2(n10782), .ZN(n10966) );
  OR2_X1 U10819 ( .A1(n8066), .A2(n8107), .ZN(n10782) );
  OR2_X1 U10820 ( .A1(n10967), .A2(n10968), .ZN(n10781) );
  AND2_X1 U10821 ( .A1(n10778), .A2(n10777), .ZN(n10968) );
  AND2_X1 U10822 ( .A1(n10775), .A2(n10969), .ZN(n10967) );
  OR2_X1 U10823 ( .A1(n10777), .A2(n10778), .ZN(n10969) );
  OR2_X1 U10824 ( .A1(n8107), .A2(n8070), .ZN(n10778) );
  OR2_X1 U10825 ( .A1(n10970), .A2(n10971), .ZN(n10777) );
  AND2_X1 U10826 ( .A1(n10774), .A2(n10773), .ZN(n10971) );
  AND2_X1 U10827 ( .A1(n10771), .A2(n10972), .ZN(n10970) );
  OR2_X1 U10828 ( .A1(n10773), .A2(n10774), .ZN(n10972) );
  OR2_X1 U10829 ( .A1(n8075), .A2(n8107), .ZN(n10774) );
  OR2_X1 U10830 ( .A1(n10973), .A2(n10974), .ZN(n10773) );
  AND2_X1 U10831 ( .A1(n10770), .A2(n10769), .ZN(n10974) );
  AND2_X1 U10832 ( .A1(n10767), .A2(n10975), .ZN(n10973) );
  OR2_X1 U10833 ( .A1(n10769), .A2(n10770), .ZN(n10975) );
  OR2_X1 U10834 ( .A1(n8107), .A2(n8079), .ZN(n10770) );
  OR2_X1 U10835 ( .A1(n10976), .A2(n10977), .ZN(n10769) );
  AND2_X1 U10836 ( .A1(n10766), .A2(n10765), .ZN(n10977) );
  AND2_X1 U10837 ( .A1(n10763), .A2(n10978), .ZN(n10976) );
  OR2_X1 U10838 ( .A1(n10765), .A2(n10766), .ZN(n10978) );
  OR2_X1 U10839 ( .A1(n8084), .A2(n8107), .ZN(n10766) );
  OR2_X1 U10840 ( .A1(n10979), .A2(n10980), .ZN(n10765) );
  AND2_X1 U10841 ( .A1(n10762), .A2(n10761), .ZN(n10980) );
  AND2_X1 U10842 ( .A1(n10759), .A2(n10981), .ZN(n10979) );
  OR2_X1 U10843 ( .A1(n10761), .A2(n10762), .ZN(n10981) );
  OR2_X1 U10844 ( .A1(n8107), .A2(n8088), .ZN(n10762) );
  OR2_X1 U10845 ( .A1(n10982), .A2(n10983), .ZN(n10761) );
  AND2_X1 U10846 ( .A1(n10758), .A2(n10757), .ZN(n10983) );
  AND2_X1 U10847 ( .A1(n10755), .A2(n10984), .ZN(n10982) );
  OR2_X1 U10848 ( .A1(n10757), .A2(n10758), .ZN(n10984) );
  OR2_X1 U10849 ( .A1(n8093), .A2(n8107), .ZN(n10758) );
  OR2_X1 U10850 ( .A1(n10985), .A2(n10986), .ZN(n10757) );
  AND2_X1 U10851 ( .A1(n10754), .A2(n10753), .ZN(n10986) );
  AND2_X1 U10852 ( .A1(n10751), .A2(n10987), .ZN(n10985) );
  OR2_X1 U10853 ( .A1(n10753), .A2(n10754), .ZN(n10987) );
  OR2_X1 U10854 ( .A1(n8107), .A2(n8097), .ZN(n10754) );
  OR2_X1 U10855 ( .A1(n10988), .A2(n10989), .ZN(n10753) );
  AND2_X1 U10856 ( .A1(n10750), .A2(n10749), .ZN(n10989) );
  AND2_X1 U10857 ( .A1(n10747), .A2(n10990), .ZN(n10988) );
  OR2_X1 U10858 ( .A1(n10749), .A2(n10750), .ZN(n10990) );
  OR2_X1 U10859 ( .A1(n8102), .A2(n8107), .ZN(n10750) );
  OR2_X1 U10860 ( .A1(n10991), .A2(n10992), .ZN(n10749) );
  AND2_X1 U10861 ( .A1(n7734), .A2(n10746), .ZN(n10992) );
  AND2_X1 U10862 ( .A1(n10744), .A2(n10993), .ZN(n10991) );
  OR2_X1 U10863 ( .A1(n10746), .A2(n7734), .ZN(n10993) );
  OR2_X1 U10864 ( .A1(n8106), .A2(n8107), .ZN(n7734) );
  OR2_X1 U10865 ( .A1(n10994), .A2(n10995), .ZN(n10746) );
  AND2_X1 U10866 ( .A1(n10743), .A2(n10742), .ZN(n10995) );
  AND2_X1 U10867 ( .A1(n10740), .A2(n10996), .ZN(n10994) );
  OR2_X1 U10868 ( .A1(n10742), .A2(n10743), .ZN(n10996) );
  OR2_X1 U10869 ( .A1(n8109), .A2(n8107), .ZN(n10743) );
  OR2_X1 U10870 ( .A1(n10997), .A2(n10998), .ZN(n10742) );
  AND2_X1 U10871 ( .A1(n10739), .A2(n10738), .ZN(n10998) );
  AND2_X1 U10872 ( .A1(n10736), .A2(n10999), .ZN(n10997) );
  OR2_X1 U10873 ( .A1(n10738), .A2(n10739), .ZN(n10999) );
  OR2_X1 U10874 ( .A1(n8112), .A2(n8107), .ZN(n10739) );
  OR2_X1 U10875 ( .A1(n11000), .A2(n11001), .ZN(n10738) );
  AND2_X1 U10876 ( .A1(n10735), .A2(n10734), .ZN(n11001) );
  AND2_X1 U10877 ( .A1(n10732), .A2(n11002), .ZN(n11000) );
  OR2_X1 U10878 ( .A1(n10734), .A2(n10735), .ZN(n11002) );
  OR2_X1 U10879 ( .A1(n8115), .A2(n8107), .ZN(n10735) );
  OR2_X1 U10880 ( .A1(n11003), .A2(n11004), .ZN(n10734) );
  AND2_X1 U10881 ( .A1(n10731), .A2(n10730), .ZN(n11004) );
  AND2_X1 U10882 ( .A1(n10728), .A2(n11005), .ZN(n11003) );
  OR2_X1 U10883 ( .A1(n10730), .A2(n10731), .ZN(n11005) );
  OR2_X1 U10884 ( .A1(n8118), .A2(n8107), .ZN(n10731) );
  OR2_X1 U10885 ( .A1(n11006), .A2(n11007), .ZN(n10730) );
  AND2_X1 U10886 ( .A1(n10727), .A2(n10726), .ZN(n11007) );
  AND2_X1 U10887 ( .A1(n10724), .A2(n11008), .ZN(n11006) );
  OR2_X1 U10888 ( .A1(n10726), .A2(n10727), .ZN(n11008) );
  OR2_X1 U10889 ( .A1(n8121), .A2(n8107), .ZN(n10727) );
  OR2_X1 U10890 ( .A1(n11009), .A2(n11010), .ZN(n10726) );
  AND2_X1 U10891 ( .A1(n10723), .A2(n10722), .ZN(n11010) );
  AND2_X1 U10892 ( .A1(n10720), .A2(n11011), .ZN(n11009) );
  OR2_X1 U10893 ( .A1(n10722), .A2(n10723), .ZN(n11011) );
  OR2_X1 U10894 ( .A1(n8124), .A2(n8107), .ZN(n10723) );
  OR2_X1 U10895 ( .A1(n11012), .A2(n11013), .ZN(n10722) );
  AND2_X1 U10896 ( .A1(n10716), .A2(n10719), .ZN(n11013) );
  AND2_X1 U10897 ( .A1(n11014), .A2(n11015), .ZN(n11012) );
  OR2_X1 U10898 ( .A1(n10719), .A2(n10716), .ZN(n11015) );
  OR2_X1 U10899 ( .A1(n8127), .A2(n8107), .ZN(n10716) );
  OR3_X1 U10900 ( .A1(n8103), .A2(n8981), .A3(n8107), .ZN(n10719) );
  INV_X1 U10901 ( .A(b_22_), .ZN(n8107) );
  INV_X1 U10902 ( .A(n10718), .ZN(n11014) );
  OR2_X1 U10903 ( .A1(n11016), .A2(n11017), .ZN(n10718) );
  AND2_X1 U10904 ( .A1(b_21_), .A2(n11018), .ZN(n11017) );
  OR2_X1 U10905 ( .A1(n11019), .A2(n7598), .ZN(n11018) );
  AND2_X1 U10906 ( .A1(a_30_), .A2(n8098), .ZN(n11019) );
  AND2_X1 U10907 ( .A1(b_20_), .A2(n11020), .ZN(n11016) );
  OR2_X1 U10908 ( .A1(n11021), .A2(n7601), .ZN(n11020) );
  AND2_X1 U10909 ( .A1(a_31_), .A2(n8103), .ZN(n11021) );
  XNOR2_X1 U10910 ( .A(n11022), .B(n11023), .ZN(n10720) );
  XOR2_X1 U10911 ( .A(n11024), .B(n11025), .Z(n11023) );
  XOR2_X1 U10912 ( .A(n11026), .B(n11027), .Z(n10724) );
  XOR2_X1 U10913 ( .A(n11028), .B(n11029), .Z(n11027) );
  XOR2_X1 U10914 ( .A(n11030), .B(n11031), .Z(n10728) );
  XOR2_X1 U10915 ( .A(n11032), .B(n11033), .Z(n11031) );
  XOR2_X1 U10916 ( .A(n11034), .B(n11035), .Z(n10732) );
  XOR2_X1 U10917 ( .A(n11036), .B(n11037), .Z(n11035) );
  XOR2_X1 U10918 ( .A(n11038), .B(n11039), .Z(n10736) );
  XOR2_X1 U10919 ( .A(n11040), .B(n11041), .Z(n11039) );
  XOR2_X1 U10920 ( .A(n11042), .B(n11043), .Z(n10740) );
  XOR2_X1 U10921 ( .A(n11044), .B(n11045), .Z(n11043) );
  XOR2_X1 U10922 ( .A(n11046), .B(n11047), .Z(n10744) );
  XOR2_X1 U10923 ( .A(n11048), .B(n11049), .Z(n11047) );
  XOR2_X1 U10924 ( .A(n11050), .B(n11051), .Z(n10747) );
  XOR2_X1 U10925 ( .A(n11052), .B(n11053), .Z(n11051) );
  XOR2_X1 U10926 ( .A(n11054), .B(n11055), .Z(n10751) );
  XOR2_X1 U10927 ( .A(n11056), .B(n8104), .Z(n11055) );
  XOR2_X1 U10928 ( .A(n11057), .B(n11058), .Z(n10755) );
  XOR2_X1 U10929 ( .A(n11059), .B(n11060), .Z(n11058) );
  XOR2_X1 U10930 ( .A(n11061), .B(n11062), .Z(n10759) );
  XOR2_X1 U10931 ( .A(n11063), .B(n11064), .Z(n11062) );
  XOR2_X1 U10932 ( .A(n11065), .B(n11066), .Z(n10763) );
  XOR2_X1 U10933 ( .A(n11067), .B(n11068), .Z(n11066) );
  XOR2_X1 U10934 ( .A(n11069), .B(n11070), .Z(n10767) );
  XOR2_X1 U10935 ( .A(n11071), .B(n11072), .Z(n11070) );
  XOR2_X1 U10936 ( .A(n11073), .B(n11074), .Z(n10771) );
  XOR2_X1 U10937 ( .A(n11075), .B(n11076), .Z(n11074) );
  XOR2_X1 U10938 ( .A(n11077), .B(n11078), .Z(n10775) );
  XOR2_X1 U10939 ( .A(n11079), .B(n11080), .Z(n11078) );
  XOR2_X1 U10940 ( .A(n11081), .B(n11082), .Z(n10779) );
  XOR2_X1 U10941 ( .A(n11083), .B(n11084), .Z(n11082) );
  XOR2_X1 U10942 ( .A(n11085), .B(n11086), .Z(n10783) );
  XOR2_X1 U10943 ( .A(n11087), .B(n11088), .Z(n11086) );
  XOR2_X1 U10944 ( .A(n11089), .B(n11090), .Z(n10787) );
  XOR2_X1 U10945 ( .A(n11091), .B(n11092), .Z(n11090) );
  XOR2_X1 U10946 ( .A(n11093), .B(n11094), .Z(n10791) );
  XOR2_X1 U10947 ( .A(n11095), .B(n11096), .Z(n11094) );
  XOR2_X1 U10948 ( .A(n11097), .B(n11098), .Z(n10795) );
  XOR2_X1 U10949 ( .A(n11099), .B(n11100), .Z(n11098) );
  XOR2_X1 U10950 ( .A(n11101), .B(n11102), .Z(n10799) );
  XOR2_X1 U10951 ( .A(n11103), .B(n11104), .Z(n11102) );
  XOR2_X1 U10952 ( .A(n11105), .B(n11106), .Z(n10803) );
  XOR2_X1 U10953 ( .A(n11107), .B(n11108), .Z(n11106) );
  XOR2_X1 U10954 ( .A(n11109), .B(n11110), .Z(n10807) );
  XOR2_X1 U10955 ( .A(n11111), .B(n11112), .Z(n11110) );
  XOR2_X1 U10956 ( .A(n11113), .B(n11114), .Z(n10811) );
  XOR2_X1 U10957 ( .A(n11115), .B(n11116), .Z(n11114) );
  XOR2_X1 U10958 ( .A(n11117), .B(n11118), .Z(n10815) );
  XOR2_X1 U10959 ( .A(n11119), .B(n11120), .Z(n11118) );
  XOR2_X1 U10960 ( .A(n11121), .B(n11122), .Z(n10020) );
  XOR2_X1 U10961 ( .A(n11123), .B(n11124), .Z(n11122) );
  XOR2_X1 U10962 ( .A(n11125), .B(n11126), .Z(n10001) );
  XOR2_X1 U10963 ( .A(n11127), .B(n11128), .Z(n11126) );
  XOR2_X1 U10964 ( .A(n11129), .B(n11130), .Z(n8860) );
  XOR2_X1 U10965 ( .A(n11131), .B(n11132), .Z(n11130) );
  XOR2_X1 U10966 ( .A(n10877), .B(n11133), .Z(n8836) );
  XOR2_X1 U10967 ( .A(n10876), .B(n10875), .Z(n11133) );
  OR2_X1 U10968 ( .A1(n8103), .A2(n8012), .ZN(n10875) );
  OR2_X1 U10969 ( .A1(n11134), .A2(n11135), .ZN(n10876) );
  AND2_X1 U10970 ( .A1(n11132), .A2(n11131), .ZN(n11135) );
  AND2_X1 U10971 ( .A1(n11129), .A2(n11136), .ZN(n11134) );
  OR2_X1 U10972 ( .A1(n11132), .A2(n11131), .ZN(n11136) );
  OR2_X1 U10973 ( .A1(n11137), .A2(n11138), .ZN(n11131) );
  AND2_X1 U10974 ( .A1(n11128), .A2(n11127), .ZN(n11138) );
  AND2_X1 U10975 ( .A1(n11125), .A2(n11139), .ZN(n11137) );
  OR2_X1 U10976 ( .A1(n11128), .A2(n11127), .ZN(n11139) );
  OR2_X1 U10977 ( .A1(n11140), .A2(n11141), .ZN(n11127) );
  AND2_X1 U10978 ( .A1(n11124), .A2(n11123), .ZN(n11141) );
  AND2_X1 U10979 ( .A1(n11121), .A2(n11142), .ZN(n11140) );
  OR2_X1 U10980 ( .A1(n11124), .A2(n11123), .ZN(n11142) );
  OR2_X1 U10981 ( .A1(n11143), .A2(n11144), .ZN(n11123) );
  AND2_X1 U10982 ( .A1(n11120), .A2(n11119), .ZN(n11144) );
  AND2_X1 U10983 ( .A1(n11117), .A2(n11145), .ZN(n11143) );
  OR2_X1 U10984 ( .A1(n11120), .A2(n11119), .ZN(n11145) );
  OR2_X1 U10985 ( .A1(n11146), .A2(n11147), .ZN(n11119) );
  AND2_X1 U10986 ( .A1(n11116), .A2(n11115), .ZN(n11147) );
  AND2_X1 U10987 ( .A1(n11113), .A2(n11148), .ZN(n11146) );
  OR2_X1 U10988 ( .A1(n11116), .A2(n11115), .ZN(n11148) );
  OR2_X1 U10989 ( .A1(n11149), .A2(n11150), .ZN(n11115) );
  AND2_X1 U10990 ( .A1(n11112), .A2(n11111), .ZN(n11150) );
  AND2_X1 U10991 ( .A1(n11109), .A2(n11151), .ZN(n11149) );
  OR2_X1 U10992 ( .A1(n11112), .A2(n11111), .ZN(n11151) );
  OR2_X1 U10993 ( .A1(n11152), .A2(n11153), .ZN(n11111) );
  AND2_X1 U10994 ( .A1(n11108), .A2(n11107), .ZN(n11153) );
  AND2_X1 U10995 ( .A1(n11105), .A2(n11154), .ZN(n11152) );
  OR2_X1 U10996 ( .A1(n11108), .A2(n11107), .ZN(n11154) );
  OR2_X1 U10997 ( .A1(n11155), .A2(n11156), .ZN(n11107) );
  AND2_X1 U10998 ( .A1(n11104), .A2(n11103), .ZN(n11156) );
  AND2_X1 U10999 ( .A1(n11101), .A2(n11157), .ZN(n11155) );
  OR2_X1 U11000 ( .A1(n11104), .A2(n11103), .ZN(n11157) );
  OR2_X1 U11001 ( .A1(n11158), .A2(n11159), .ZN(n11103) );
  AND2_X1 U11002 ( .A1(n11100), .A2(n11099), .ZN(n11159) );
  AND2_X1 U11003 ( .A1(n11097), .A2(n11160), .ZN(n11158) );
  OR2_X1 U11004 ( .A1(n11100), .A2(n11099), .ZN(n11160) );
  OR2_X1 U11005 ( .A1(n11161), .A2(n11162), .ZN(n11099) );
  AND2_X1 U11006 ( .A1(n11096), .A2(n11095), .ZN(n11162) );
  AND2_X1 U11007 ( .A1(n11093), .A2(n11163), .ZN(n11161) );
  OR2_X1 U11008 ( .A1(n11096), .A2(n11095), .ZN(n11163) );
  OR2_X1 U11009 ( .A1(n11164), .A2(n11165), .ZN(n11095) );
  AND2_X1 U11010 ( .A1(n11092), .A2(n11091), .ZN(n11165) );
  AND2_X1 U11011 ( .A1(n11089), .A2(n11166), .ZN(n11164) );
  OR2_X1 U11012 ( .A1(n11092), .A2(n11091), .ZN(n11166) );
  OR2_X1 U11013 ( .A1(n11167), .A2(n11168), .ZN(n11091) );
  AND2_X1 U11014 ( .A1(n11088), .A2(n11087), .ZN(n11168) );
  AND2_X1 U11015 ( .A1(n11085), .A2(n11169), .ZN(n11167) );
  OR2_X1 U11016 ( .A1(n11088), .A2(n11087), .ZN(n11169) );
  OR2_X1 U11017 ( .A1(n11170), .A2(n11171), .ZN(n11087) );
  AND2_X1 U11018 ( .A1(n11084), .A2(n11083), .ZN(n11171) );
  AND2_X1 U11019 ( .A1(n11081), .A2(n11172), .ZN(n11170) );
  OR2_X1 U11020 ( .A1(n11084), .A2(n11083), .ZN(n11172) );
  OR2_X1 U11021 ( .A1(n11173), .A2(n11174), .ZN(n11083) );
  AND2_X1 U11022 ( .A1(n11080), .A2(n11079), .ZN(n11174) );
  AND2_X1 U11023 ( .A1(n11077), .A2(n11175), .ZN(n11173) );
  OR2_X1 U11024 ( .A1(n11080), .A2(n11079), .ZN(n11175) );
  OR2_X1 U11025 ( .A1(n11176), .A2(n11177), .ZN(n11079) );
  AND2_X1 U11026 ( .A1(n11076), .A2(n11075), .ZN(n11177) );
  AND2_X1 U11027 ( .A1(n11073), .A2(n11178), .ZN(n11176) );
  OR2_X1 U11028 ( .A1(n11076), .A2(n11075), .ZN(n11178) );
  OR2_X1 U11029 ( .A1(n11179), .A2(n11180), .ZN(n11075) );
  AND2_X1 U11030 ( .A1(n11072), .A2(n11071), .ZN(n11180) );
  AND2_X1 U11031 ( .A1(n11069), .A2(n11181), .ZN(n11179) );
  OR2_X1 U11032 ( .A1(n11072), .A2(n11071), .ZN(n11181) );
  OR2_X1 U11033 ( .A1(n11182), .A2(n11183), .ZN(n11071) );
  AND2_X1 U11034 ( .A1(n11068), .A2(n11067), .ZN(n11183) );
  AND2_X1 U11035 ( .A1(n11065), .A2(n11184), .ZN(n11182) );
  OR2_X1 U11036 ( .A1(n11068), .A2(n11067), .ZN(n11184) );
  OR2_X1 U11037 ( .A1(n11185), .A2(n11186), .ZN(n11067) );
  AND2_X1 U11038 ( .A1(n11064), .A2(n11063), .ZN(n11186) );
  AND2_X1 U11039 ( .A1(n11061), .A2(n11187), .ZN(n11185) );
  OR2_X1 U11040 ( .A1(n11064), .A2(n11063), .ZN(n11187) );
  OR2_X1 U11041 ( .A1(n11188), .A2(n11189), .ZN(n11063) );
  AND2_X1 U11042 ( .A1(n11060), .A2(n11059), .ZN(n11189) );
  AND2_X1 U11043 ( .A1(n11057), .A2(n11190), .ZN(n11188) );
  OR2_X1 U11044 ( .A1(n11060), .A2(n11059), .ZN(n11190) );
  OR2_X1 U11045 ( .A1(n11191), .A2(n11192), .ZN(n11059) );
  AND2_X1 U11046 ( .A1(n8104), .A2(n11056), .ZN(n11192) );
  AND2_X1 U11047 ( .A1(n11054), .A2(n11193), .ZN(n11191) );
  OR2_X1 U11048 ( .A1(n8104), .A2(n11056), .ZN(n11193) );
  OR2_X1 U11049 ( .A1(n11194), .A2(n11195), .ZN(n11056) );
  AND2_X1 U11050 ( .A1(n11053), .A2(n11052), .ZN(n11195) );
  AND2_X1 U11051 ( .A1(n11050), .A2(n11196), .ZN(n11194) );
  OR2_X1 U11052 ( .A1(n11053), .A2(n11052), .ZN(n11196) );
  OR2_X1 U11053 ( .A1(n11197), .A2(n11198), .ZN(n11052) );
  AND2_X1 U11054 ( .A1(n11049), .A2(n11048), .ZN(n11198) );
  AND2_X1 U11055 ( .A1(n11046), .A2(n11199), .ZN(n11197) );
  OR2_X1 U11056 ( .A1(n11049), .A2(n11048), .ZN(n11199) );
  OR2_X1 U11057 ( .A1(n11200), .A2(n11201), .ZN(n11048) );
  AND2_X1 U11058 ( .A1(n11045), .A2(n11044), .ZN(n11201) );
  AND2_X1 U11059 ( .A1(n11042), .A2(n11202), .ZN(n11200) );
  OR2_X1 U11060 ( .A1(n11045), .A2(n11044), .ZN(n11202) );
  OR2_X1 U11061 ( .A1(n11203), .A2(n11204), .ZN(n11044) );
  AND2_X1 U11062 ( .A1(n11041), .A2(n11040), .ZN(n11204) );
  AND2_X1 U11063 ( .A1(n11038), .A2(n11205), .ZN(n11203) );
  OR2_X1 U11064 ( .A1(n11041), .A2(n11040), .ZN(n11205) );
  OR2_X1 U11065 ( .A1(n11206), .A2(n11207), .ZN(n11040) );
  AND2_X1 U11066 ( .A1(n11037), .A2(n11036), .ZN(n11207) );
  AND2_X1 U11067 ( .A1(n11034), .A2(n11208), .ZN(n11206) );
  OR2_X1 U11068 ( .A1(n11037), .A2(n11036), .ZN(n11208) );
  OR2_X1 U11069 ( .A1(n11209), .A2(n11210), .ZN(n11036) );
  AND2_X1 U11070 ( .A1(n11033), .A2(n11032), .ZN(n11210) );
  AND2_X1 U11071 ( .A1(n11030), .A2(n11211), .ZN(n11209) );
  OR2_X1 U11072 ( .A1(n11033), .A2(n11032), .ZN(n11211) );
  OR2_X1 U11073 ( .A1(n11212), .A2(n11213), .ZN(n11032) );
  AND2_X1 U11074 ( .A1(n11029), .A2(n11028), .ZN(n11213) );
  AND2_X1 U11075 ( .A1(n11026), .A2(n11214), .ZN(n11212) );
  OR2_X1 U11076 ( .A1(n11029), .A2(n11028), .ZN(n11214) );
  OR2_X1 U11077 ( .A1(n11215), .A2(n11216), .ZN(n11028) );
  AND2_X1 U11078 ( .A1(n11022), .A2(n11025), .ZN(n11216) );
  AND2_X1 U11079 ( .A1(n11217), .A2(n11218), .ZN(n11215) );
  OR2_X1 U11080 ( .A1(n11022), .A2(n11025), .ZN(n11218) );
  OR3_X1 U11081 ( .A1(n8098), .A2(n8103), .A3(n8981), .ZN(n11025) );
  OR2_X1 U11082 ( .A1(n8103), .A2(n8127), .ZN(n11022) );
  INV_X1 U11083 ( .A(n11024), .ZN(n11217) );
  OR2_X1 U11084 ( .A1(n11219), .A2(n11220), .ZN(n11024) );
  AND2_X1 U11085 ( .A1(b_20_), .A2(n11221), .ZN(n11220) );
  OR2_X1 U11086 ( .A1(n11222), .A2(n7598), .ZN(n11221) );
  AND2_X1 U11087 ( .A1(a_30_), .A2(n8094), .ZN(n11222) );
  AND2_X1 U11088 ( .A1(b_19_), .A2(n11223), .ZN(n11219) );
  OR2_X1 U11089 ( .A1(n11224), .A2(n7601), .ZN(n11223) );
  AND2_X1 U11090 ( .A1(a_31_), .A2(n8098), .ZN(n11224) );
  OR2_X1 U11091 ( .A1(n8103), .A2(n8124), .ZN(n11029) );
  XNOR2_X1 U11092 ( .A(n11225), .B(n11226), .ZN(n11026) );
  XOR2_X1 U11093 ( .A(n11227), .B(n11228), .Z(n11226) );
  OR2_X1 U11094 ( .A1(n8103), .A2(n8121), .ZN(n11033) );
  XOR2_X1 U11095 ( .A(n11229), .B(n11230), .Z(n11030) );
  XOR2_X1 U11096 ( .A(n11231), .B(n11232), .Z(n11230) );
  OR2_X1 U11097 ( .A1(n8103), .A2(n8118), .ZN(n11037) );
  XOR2_X1 U11098 ( .A(n11233), .B(n11234), .Z(n11034) );
  XOR2_X1 U11099 ( .A(n11235), .B(n11236), .Z(n11234) );
  OR2_X1 U11100 ( .A1(n8103), .A2(n8115), .ZN(n11041) );
  XOR2_X1 U11101 ( .A(n11237), .B(n11238), .Z(n11038) );
  XOR2_X1 U11102 ( .A(n11239), .B(n11240), .Z(n11238) );
  OR2_X1 U11103 ( .A1(n8103), .A2(n8112), .ZN(n11045) );
  XOR2_X1 U11104 ( .A(n11241), .B(n11242), .Z(n11042) );
  XOR2_X1 U11105 ( .A(n11243), .B(n11244), .Z(n11242) );
  OR2_X1 U11106 ( .A1(n8103), .A2(n8109), .ZN(n11049) );
  XOR2_X1 U11107 ( .A(n11245), .B(n11246), .Z(n11046) );
  XOR2_X1 U11108 ( .A(n11247), .B(n11248), .Z(n11246) );
  OR2_X1 U11109 ( .A1(n8103), .A2(n8106), .ZN(n11053) );
  XOR2_X1 U11110 ( .A(n11249), .B(n11250), .Z(n11050) );
  XOR2_X1 U11111 ( .A(n11251), .B(n11252), .Z(n11250) );
  OR2_X1 U11112 ( .A1(n8102), .A2(n8103), .ZN(n8104) );
  XOR2_X1 U11113 ( .A(n11253), .B(n11254), .Z(n11054) );
  XOR2_X1 U11114 ( .A(n11255), .B(n11256), .Z(n11254) );
  OR2_X1 U11115 ( .A1(n8103), .A2(n8097), .ZN(n11060) );
  XOR2_X1 U11116 ( .A(n11257), .B(n11258), .Z(n11057) );
  XOR2_X1 U11117 ( .A(n11259), .B(n11260), .Z(n11258) );
  OR2_X1 U11118 ( .A1(n8093), .A2(n8103), .ZN(n11064) );
  XNOR2_X1 U11119 ( .A(n11261), .B(n11262), .ZN(n11061) );
  XOR2_X1 U11120 ( .A(n7758), .B(n11263), .Z(n11261) );
  INV_X1 U11121 ( .A(n8099), .ZN(n7758) );
  OR2_X1 U11122 ( .A1(n8103), .A2(n8088), .ZN(n11068) );
  XOR2_X1 U11123 ( .A(n11264), .B(n11265), .Z(n11065) );
  XOR2_X1 U11124 ( .A(n11266), .B(n11267), .Z(n11265) );
  OR2_X1 U11125 ( .A1(n8084), .A2(n8103), .ZN(n11072) );
  XOR2_X1 U11126 ( .A(n11268), .B(n11269), .Z(n11069) );
  XOR2_X1 U11127 ( .A(n11270), .B(n11271), .Z(n11269) );
  OR2_X1 U11128 ( .A1(n8103), .A2(n8079), .ZN(n11076) );
  XOR2_X1 U11129 ( .A(n11272), .B(n11273), .Z(n11073) );
  XOR2_X1 U11130 ( .A(n11274), .B(n11275), .Z(n11273) );
  OR2_X1 U11131 ( .A1(n8075), .A2(n8103), .ZN(n11080) );
  XOR2_X1 U11132 ( .A(n11276), .B(n11277), .Z(n11077) );
  XOR2_X1 U11133 ( .A(n11278), .B(n11279), .Z(n11277) );
  OR2_X1 U11134 ( .A1(n8103), .A2(n8070), .ZN(n11084) );
  XOR2_X1 U11135 ( .A(n11280), .B(n11281), .Z(n11081) );
  XOR2_X1 U11136 ( .A(n11282), .B(n11283), .Z(n11281) );
  OR2_X1 U11137 ( .A1(n8066), .A2(n8103), .ZN(n11088) );
  XOR2_X1 U11138 ( .A(n11284), .B(n11285), .Z(n11085) );
  XOR2_X1 U11139 ( .A(n11286), .B(n11287), .Z(n11285) );
  OR2_X1 U11140 ( .A1(n8103), .A2(n8061), .ZN(n11092) );
  XOR2_X1 U11141 ( .A(n11288), .B(n11289), .Z(n11089) );
  XOR2_X1 U11142 ( .A(n11290), .B(n11291), .Z(n11289) );
  OR2_X1 U11143 ( .A1(n8057), .A2(n8103), .ZN(n11096) );
  XOR2_X1 U11144 ( .A(n11292), .B(n11293), .Z(n11093) );
  XOR2_X1 U11145 ( .A(n11294), .B(n11295), .Z(n11293) );
  OR2_X1 U11146 ( .A1(n8103), .A2(n8052), .ZN(n11100) );
  XOR2_X1 U11147 ( .A(n11296), .B(n11297), .Z(n11097) );
  XOR2_X1 U11148 ( .A(n11298), .B(n11299), .Z(n11297) );
  OR2_X1 U11149 ( .A1(n8048), .A2(n8103), .ZN(n11104) );
  XOR2_X1 U11150 ( .A(n11300), .B(n11301), .Z(n11101) );
  XOR2_X1 U11151 ( .A(n11302), .B(n11303), .Z(n11301) );
  OR2_X1 U11152 ( .A1(n8103), .A2(n8043), .ZN(n11108) );
  XOR2_X1 U11153 ( .A(n11304), .B(n11305), .Z(n11105) );
  XOR2_X1 U11154 ( .A(n11306), .B(n11307), .Z(n11305) );
  OR2_X1 U11155 ( .A1(n8039), .A2(n8103), .ZN(n11112) );
  XOR2_X1 U11156 ( .A(n11308), .B(n11309), .Z(n11109) );
  XOR2_X1 U11157 ( .A(n11310), .B(n11311), .Z(n11309) );
  OR2_X1 U11158 ( .A1(n8103), .A2(n8034), .ZN(n11116) );
  XOR2_X1 U11159 ( .A(n11312), .B(n11313), .Z(n11113) );
  XOR2_X1 U11160 ( .A(n11314), .B(n11315), .Z(n11313) );
  OR2_X1 U11161 ( .A1(n8030), .A2(n8103), .ZN(n11120) );
  XOR2_X1 U11162 ( .A(n11316), .B(n11317), .Z(n11117) );
  XOR2_X1 U11163 ( .A(n11318), .B(n11319), .Z(n11317) );
  OR2_X1 U11164 ( .A1(n8103), .A2(n8025), .ZN(n11124) );
  XOR2_X1 U11165 ( .A(n11320), .B(n11321), .Z(n11121) );
  XOR2_X1 U11166 ( .A(n11322), .B(n11323), .Z(n11321) );
  OR2_X1 U11167 ( .A1(n8021), .A2(n8103), .ZN(n11128) );
  XOR2_X1 U11168 ( .A(n11324), .B(n11325), .Z(n11125) );
  XOR2_X1 U11169 ( .A(n11326), .B(n11327), .Z(n11325) );
  OR2_X1 U11170 ( .A1(n8103), .A2(n8016), .ZN(n11132) );
  XOR2_X1 U11171 ( .A(n11328), .B(n11329), .Z(n11129) );
  XOR2_X1 U11172 ( .A(n11330), .B(n11331), .Z(n11329) );
  XOR2_X1 U11173 ( .A(n10884), .B(n11332), .Z(n10877) );
  XOR2_X1 U11174 ( .A(n10883), .B(n10882), .Z(n11332) );
  OR2_X1 U11175 ( .A1(n8098), .A2(n8016), .ZN(n10882) );
  OR2_X1 U11176 ( .A1(n11333), .A2(n11334), .ZN(n10883) );
  AND2_X1 U11177 ( .A1(n11331), .A2(n11330), .ZN(n11334) );
  AND2_X1 U11178 ( .A1(n11328), .A2(n11335), .ZN(n11333) );
  OR2_X1 U11179 ( .A1(n11331), .A2(n11330), .ZN(n11335) );
  OR2_X1 U11180 ( .A1(n11336), .A2(n11337), .ZN(n11330) );
  AND2_X1 U11181 ( .A1(n11327), .A2(n11326), .ZN(n11337) );
  AND2_X1 U11182 ( .A1(n11324), .A2(n11338), .ZN(n11336) );
  OR2_X1 U11183 ( .A1(n11327), .A2(n11326), .ZN(n11338) );
  OR2_X1 U11184 ( .A1(n11339), .A2(n11340), .ZN(n11326) );
  AND2_X1 U11185 ( .A1(n11323), .A2(n11322), .ZN(n11340) );
  AND2_X1 U11186 ( .A1(n11320), .A2(n11341), .ZN(n11339) );
  OR2_X1 U11187 ( .A1(n11323), .A2(n11322), .ZN(n11341) );
  OR2_X1 U11188 ( .A1(n11342), .A2(n11343), .ZN(n11322) );
  AND2_X1 U11189 ( .A1(n11319), .A2(n11318), .ZN(n11343) );
  AND2_X1 U11190 ( .A1(n11316), .A2(n11344), .ZN(n11342) );
  OR2_X1 U11191 ( .A1(n11319), .A2(n11318), .ZN(n11344) );
  OR2_X1 U11192 ( .A1(n11345), .A2(n11346), .ZN(n11318) );
  AND2_X1 U11193 ( .A1(n11315), .A2(n11314), .ZN(n11346) );
  AND2_X1 U11194 ( .A1(n11312), .A2(n11347), .ZN(n11345) );
  OR2_X1 U11195 ( .A1(n11315), .A2(n11314), .ZN(n11347) );
  OR2_X1 U11196 ( .A1(n11348), .A2(n11349), .ZN(n11314) );
  AND2_X1 U11197 ( .A1(n11311), .A2(n11310), .ZN(n11349) );
  AND2_X1 U11198 ( .A1(n11308), .A2(n11350), .ZN(n11348) );
  OR2_X1 U11199 ( .A1(n11311), .A2(n11310), .ZN(n11350) );
  OR2_X1 U11200 ( .A1(n11351), .A2(n11352), .ZN(n11310) );
  AND2_X1 U11201 ( .A1(n11307), .A2(n11306), .ZN(n11352) );
  AND2_X1 U11202 ( .A1(n11304), .A2(n11353), .ZN(n11351) );
  OR2_X1 U11203 ( .A1(n11307), .A2(n11306), .ZN(n11353) );
  OR2_X1 U11204 ( .A1(n11354), .A2(n11355), .ZN(n11306) );
  AND2_X1 U11205 ( .A1(n11303), .A2(n11302), .ZN(n11355) );
  AND2_X1 U11206 ( .A1(n11300), .A2(n11356), .ZN(n11354) );
  OR2_X1 U11207 ( .A1(n11303), .A2(n11302), .ZN(n11356) );
  OR2_X1 U11208 ( .A1(n11357), .A2(n11358), .ZN(n11302) );
  AND2_X1 U11209 ( .A1(n11299), .A2(n11298), .ZN(n11358) );
  AND2_X1 U11210 ( .A1(n11296), .A2(n11359), .ZN(n11357) );
  OR2_X1 U11211 ( .A1(n11299), .A2(n11298), .ZN(n11359) );
  OR2_X1 U11212 ( .A1(n11360), .A2(n11361), .ZN(n11298) );
  AND2_X1 U11213 ( .A1(n11295), .A2(n11294), .ZN(n11361) );
  AND2_X1 U11214 ( .A1(n11292), .A2(n11362), .ZN(n11360) );
  OR2_X1 U11215 ( .A1(n11295), .A2(n11294), .ZN(n11362) );
  OR2_X1 U11216 ( .A1(n11363), .A2(n11364), .ZN(n11294) );
  AND2_X1 U11217 ( .A1(n11291), .A2(n11290), .ZN(n11364) );
  AND2_X1 U11218 ( .A1(n11288), .A2(n11365), .ZN(n11363) );
  OR2_X1 U11219 ( .A1(n11291), .A2(n11290), .ZN(n11365) );
  OR2_X1 U11220 ( .A1(n11366), .A2(n11367), .ZN(n11290) );
  AND2_X1 U11221 ( .A1(n11287), .A2(n11286), .ZN(n11367) );
  AND2_X1 U11222 ( .A1(n11284), .A2(n11368), .ZN(n11366) );
  OR2_X1 U11223 ( .A1(n11287), .A2(n11286), .ZN(n11368) );
  OR2_X1 U11224 ( .A1(n11369), .A2(n11370), .ZN(n11286) );
  AND2_X1 U11225 ( .A1(n11283), .A2(n11282), .ZN(n11370) );
  AND2_X1 U11226 ( .A1(n11280), .A2(n11371), .ZN(n11369) );
  OR2_X1 U11227 ( .A1(n11283), .A2(n11282), .ZN(n11371) );
  OR2_X1 U11228 ( .A1(n11372), .A2(n11373), .ZN(n11282) );
  AND2_X1 U11229 ( .A1(n11279), .A2(n11278), .ZN(n11373) );
  AND2_X1 U11230 ( .A1(n11276), .A2(n11374), .ZN(n11372) );
  OR2_X1 U11231 ( .A1(n11279), .A2(n11278), .ZN(n11374) );
  OR2_X1 U11232 ( .A1(n11375), .A2(n11376), .ZN(n11278) );
  AND2_X1 U11233 ( .A1(n11275), .A2(n11274), .ZN(n11376) );
  AND2_X1 U11234 ( .A1(n11272), .A2(n11377), .ZN(n11375) );
  OR2_X1 U11235 ( .A1(n11275), .A2(n11274), .ZN(n11377) );
  OR2_X1 U11236 ( .A1(n11378), .A2(n11379), .ZN(n11274) );
  AND2_X1 U11237 ( .A1(n11271), .A2(n11270), .ZN(n11379) );
  AND2_X1 U11238 ( .A1(n11268), .A2(n11380), .ZN(n11378) );
  OR2_X1 U11239 ( .A1(n11271), .A2(n11270), .ZN(n11380) );
  OR2_X1 U11240 ( .A1(n11381), .A2(n11382), .ZN(n11270) );
  AND2_X1 U11241 ( .A1(n11267), .A2(n11266), .ZN(n11382) );
  AND2_X1 U11242 ( .A1(n11264), .A2(n11383), .ZN(n11381) );
  OR2_X1 U11243 ( .A1(n11267), .A2(n11266), .ZN(n11383) );
  OR2_X1 U11244 ( .A1(n11384), .A2(n11385), .ZN(n11266) );
  AND2_X1 U11245 ( .A1(n11263), .A2(n8099), .ZN(n11385) );
  AND2_X1 U11246 ( .A1(n11262), .A2(n11386), .ZN(n11384) );
  OR2_X1 U11247 ( .A1(n11263), .A2(n8099), .ZN(n11386) );
  OR2_X1 U11248 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  OR2_X1 U11249 ( .A1(n11387), .A2(n11388), .ZN(n11263) );
  AND2_X1 U11250 ( .A1(n11260), .A2(n11259), .ZN(n11388) );
  AND2_X1 U11251 ( .A1(n11257), .A2(n11389), .ZN(n11387) );
  OR2_X1 U11252 ( .A1(n11260), .A2(n11259), .ZN(n11389) );
  OR2_X1 U11253 ( .A1(n11390), .A2(n11391), .ZN(n11259) );
  AND2_X1 U11254 ( .A1(n11256), .A2(n11255), .ZN(n11391) );
  AND2_X1 U11255 ( .A1(n11253), .A2(n11392), .ZN(n11390) );
  OR2_X1 U11256 ( .A1(n11256), .A2(n11255), .ZN(n11392) );
  OR2_X1 U11257 ( .A1(n11393), .A2(n11394), .ZN(n11255) );
  AND2_X1 U11258 ( .A1(n11252), .A2(n11251), .ZN(n11394) );
  AND2_X1 U11259 ( .A1(n11249), .A2(n11395), .ZN(n11393) );
  OR2_X1 U11260 ( .A1(n11252), .A2(n11251), .ZN(n11395) );
  OR2_X1 U11261 ( .A1(n11396), .A2(n11397), .ZN(n11251) );
  AND2_X1 U11262 ( .A1(n11248), .A2(n11247), .ZN(n11397) );
  AND2_X1 U11263 ( .A1(n11245), .A2(n11398), .ZN(n11396) );
  OR2_X1 U11264 ( .A1(n11248), .A2(n11247), .ZN(n11398) );
  OR2_X1 U11265 ( .A1(n11399), .A2(n11400), .ZN(n11247) );
  AND2_X1 U11266 ( .A1(n11244), .A2(n11243), .ZN(n11400) );
  AND2_X1 U11267 ( .A1(n11241), .A2(n11401), .ZN(n11399) );
  OR2_X1 U11268 ( .A1(n11244), .A2(n11243), .ZN(n11401) );
  OR2_X1 U11269 ( .A1(n11402), .A2(n11403), .ZN(n11243) );
  AND2_X1 U11270 ( .A1(n11240), .A2(n11239), .ZN(n11403) );
  AND2_X1 U11271 ( .A1(n11237), .A2(n11404), .ZN(n11402) );
  OR2_X1 U11272 ( .A1(n11240), .A2(n11239), .ZN(n11404) );
  OR2_X1 U11273 ( .A1(n11405), .A2(n11406), .ZN(n11239) );
  AND2_X1 U11274 ( .A1(n11236), .A2(n11235), .ZN(n11406) );
  AND2_X1 U11275 ( .A1(n11233), .A2(n11407), .ZN(n11405) );
  OR2_X1 U11276 ( .A1(n11236), .A2(n11235), .ZN(n11407) );
  OR2_X1 U11277 ( .A1(n11408), .A2(n11409), .ZN(n11235) );
  AND2_X1 U11278 ( .A1(n11232), .A2(n11231), .ZN(n11409) );
  AND2_X1 U11279 ( .A1(n11229), .A2(n11410), .ZN(n11408) );
  OR2_X1 U11280 ( .A1(n11232), .A2(n11231), .ZN(n11410) );
  OR2_X1 U11281 ( .A1(n11411), .A2(n11412), .ZN(n11231) );
  AND2_X1 U11282 ( .A1(n11225), .A2(n11228), .ZN(n11412) );
  AND2_X1 U11283 ( .A1(n11413), .A2(n11414), .ZN(n11411) );
  OR2_X1 U11284 ( .A1(n11225), .A2(n11228), .ZN(n11414) );
  OR3_X1 U11285 ( .A1(n8094), .A2(n8098), .A3(n8981), .ZN(n11228) );
  OR2_X1 U11286 ( .A1(n8098), .A2(n8127), .ZN(n11225) );
  INV_X1 U11287 ( .A(n11227), .ZN(n11413) );
  OR2_X1 U11288 ( .A1(n11415), .A2(n11416), .ZN(n11227) );
  AND2_X1 U11289 ( .A1(b_19_), .A2(n11417), .ZN(n11416) );
  OR2_X1 U11290 ( .A1(n11418), .A2(n7598), .ZN(n11417) );
  AND2_X1 U11291 ( .A1(a_30_), .A2(n8089), .ZN(n11418) );
  AND2_X1 U11292 ( .A1(b_18_), .A2(n11419), .ZN(n11415) );
  OR2_X1 U11293 ( .A1(n11420), .A2(n7601), .ZN(n11419) );
  AND2_X1 U11294 ( .A1(a_31_), .A2(n8094), .ZN(n11420) );
  OR2_X1 U11295 ( .A1(n8098), .A2(n8124), .ZN(n11232) );
  XNOR2_X1 U11296 ( .A(n11421), .B(n11422), .ZN(n11229) );
  XOR2_X1 U11297 ( .A(n11423), .B(n11424), .Z(n11422) );
  OR2_X1 U11298 ( .A1(n8098), .A2(n8121), .ZN(n11236) );
  XOR2_X1 U11299 ( .A(n11425), .B(n11426), .Z(n11233) );
  XOR2_X1 U11300 ( .A(n11427), .B(n11428), .Z(n11426) );
  OR2_X1 U11301 ( .A1(n8098), .A2(n8118), .ZN(n11240) );
  XOR2_X1 U11302 ( .A(n11429), .B(n11430), .Z(n11237) );
  XOR2_X1 U11303 ( .A(n11431), .B(n11432), .Z(n11430) );
  OR2_X1 U11304 ( .A1(n8098), .A2(n8115), .ZN(n11244) );
  XOR2_X1 U11305 ( .A(n11433), .B(n11434), .Z(n11241) );
  XOR2_X1 U11306 ( .A(n11435), .B(n11436), .Z(n11434) );
  OR2_X1 U11307 ( .A1(n8098), .A2(n8112), .ZN(n11248) );
  XOR2_X1 U11308 ( .A(n11437), .B(n11438), .Z(n11245) );
  XOR2_X1 U11309 ( .A(n11439), .B(n11440), .Z(n11438) );
  OR2_X1 U11310 ( .A1(n8098), .A2(n8109), .ZN(n11252) );
  XOR2_X1 U11311 ( .A(n11441), .B(n11442), .Z(n11249) );
  XOR2_X1 U11312 ( .A(n11443), .B(n11444), .Z(n11442) );
  OR2_X1 U11313 ( .A1(n8098), .A2(n8106), .ZN(n11256) );
  XOR2_X1 U11314 ( .A(n11445), .B(n11446), .Z(n11253) );
  XOR2_X1 U11315 ( .A(n11447), .B(n11448), .Z(n11446) );
  OR2_X1 U11316 ( .A1(n8098), .A2(n8102), .ZN(n11260) );
  XOR2_X1 U11317 ( .A(n11449), .B(n11450), .Z(n11257) );
  XOR2_X1 U11318 ( .A(n11451), .B(n11452), .Z(n11450) );
  XOR2_X1 U11319 ( .A(n11453), .B(n11454), .Z(n11262) );
  XOR2_X1 U11320 ( .A(n11455), .B(n11456), .Z(n11454) );
  OR2_X1 U11321 ( .A1(n8093), .A2(n8098), .ZN(n11267) );
  XOR2_X1 U11322 ( .A(n11457), .B(n11458), .Z(n11264) );
  XOR2_X1 U11323 ( .A(n11459), .B(n11460), .Z(n11458) );
  OR2_X1 U11324 ( .A1(n8098), .A2(n8088), .ZN(n11271) );
  XOR2_X1 U11325 ( .A(n11461), .B(n11462), .Z(n11268) );
  XOR2_X1 U11326 ( .A(n11463), .B(n8095), .Z(n11462) );
  OR2_X1 U11327 ( .A1(n8084), .A2(n8098), .ZN(n11275) );
  XOR2_X1 U11328 ( .A(n11464), .B(n11465), .Z(n11272) );
  XOR2_X1 U11329 ( .A(n11466), .B(n11467), .Z(n11465) );
  OR2_X1 U11330 ( .A1(n8098), .A2(n8079), .ZN(n11279) );
  XOR2_X1 U11331 ( .A(n11468), .B(n11469), .Z(n11276) );
  XOR2_X1 U11332 ( .A(n11470), .B(n11471), .Z(n11469) );
  OR2_X1 U11333 ( .A1(n8075), .A2(n8098), .ZN(n11283) );
  XOR2_X1 U11334 ( .A(n11472), .B(n11473), .Z(n11280) );
  XOR2_X1 U11335 ( .A(n11474), .B(n11475), .Z(n11473) );
  OR2_X1 U11336 ( .A1(n8098), .A2(n8070), .ZN(n11287) );
  XOR2_X1 U11337 ( .A(n11476), .B(n11477), .Z(n11284) );
  XOR2_X1 U11338 ( .A(n11478), .B(n11479), .Z(n11477) );
  OR2_X1 U11339 ( .A1(n8066), .A2(n8098), .ZN(n11291) );
  XOR2_X1 U11340 ( .A(n11480), .B(n11481), .Z(n11288) );
  XOR2_X1 U11341 ( .A(n11482), .B(n11483), .Z(n11481) );
  OR2_X1 U11342 ( .A1(n8098), .A2(n8061), .ZN(n11295) );
  XOR2_X1 U11343 ( .A(n11484), .B(n11485), .Z(n11292) );
  XOR2_X1 U11344 ( .A(n11486), .B(n11487), .Z(n11485) );
  OR2_X1 U11345 ( .A1(n8057), .A2(n8098), .ZN(n11299) );
  XOR2_X1 U11346 ( .A(n11488), .B(n11489), .Z(n11296) );
  XOR2_X1 U11347 ( .A(n11490), .B(n11491), .Z(n11489) );
  OR2_X1 U11348 ( .A1(n8098), .A2(n8052), .ZN(n11303) );
  XOR2_X1 U11349 ( .A(n11492), .B(n11493), .Z(n11300) );
  XOR2_X1 U11350 ( .A(n11494), .B(n11495), .Z(n11493) );
  OR2_X1 U11351 ( .A1(n8048), .A2(n8098), .ZN(n11307) );
  XOR2_X1 U11352 ( .A(n11496), .B(n11497), .Z(n11304) );
  XOR2_X1 U11353 ( .A(n11498), .B(n11499), .Z(n11497) );
  OR2_X1 U11354 ( .A1(n8098), .A2(n8043), .ZN(n11311) );
  XOR2_X1 U11355 ( .A(n11500), .B(n11501), .Z(n11308) );
  XOR2_X1 U11356 ( .A(n11502), .B(n11503), .Z(n11501) );
  OR2_X1 U11357 ( .A1(n8039), .A2(n8098), .ZN(n11315) );
  XOR2_X1 U11358 ( .A(n11504), .B(n11505), .Z(n11312) );
  XOR2_X1 U11359 ( .A(n11506), .B(n11507), .Z(n11505) );
  OR2_X1 U11360 ( .A1(n8098), .A2(n8034), .ZN(n11319) );
  XOR2_X1 U11361 ( .A(n11508), .B(n11509), .Z(n11316) );
  XOR2_X1 U11362 ( .A(n11510), .B(n11511), .Z(n11509) );
  OR2_X1 U11363 ( .A1(n8030), .A2(n8098), .ZN(n11323) );
  XOR2_X1 U11364 ( .A(n11512), .B(n11513), .Z(n11320) );
  XOR2_X1 U11365 ( .A(n11514), .B(n11515), .Z(n11513) );
  OR2_X1 U11366 ( .A1(n8098), .A2(n8025), .ZN(n11327) );
  XOR2_X1 U11367 ( .A(n11516), .B(n11517), .Z(n11324) );
  XOR2_X1 U11368 ( .A(n11518), .B(n11519), .Z(n11517) );
  OR2_X1 U11369 ( .A1(n8021), .A2(n8098), .ZN(n11331) );
  INV_X1 U11370 ( .A(b_20_), .ZN(n8098) );
  XOR2_X1 U11371 ( .A(n11520), .B(n11521), .Z(n11328) );
  XOR2_X1 U11372 ( .A(n11522), .B(n11523), .Z(n11521) );
  XOR2_X1 U11373 ( .A(n10891), .B(n11524), .Z(n10884) );
  XOR2_X1 U11374 ( .A(n10890), .B(n10889), .Z(n11524) );
  OR2_X1 U11375 ( .A1(n8021), .A2(n8094), .ZN(n10889) );
  OR2_X1 U11376 ( .A1(n11525), .A2(n11526), .ZN(n10890) );
  AND2_X1 U11377 ( .A1(n11523), .A2(n11522), .ZN(n11526) );
  AND2_X1 U11378 ( .A1(n11520), .A2(n11527), .ZN(n11525) );
  OR2_X1 U11379 ( .A1(n11523), .A2(n11522), .ZN(n11527) );
  OR2_X1 U11380 ( .A1(n11528), .A2(n11529), .ZN(n11522) );
  AND2_X1 U11381 ( .A1(n11519), .A2(n11518), .ZN(n11529) );
  AND2_X1 U11382 ( .A1(n11516), .A2(n11530), .ZN(n11528) );
  OR2_X1 U11383 ( .A1(n11519), .A2(n11518), .ZN(n11530) );
  OR2_X1 U11384 ( .A1(n11531), .A2(n11532), .ZN(n11518) );
  AND2_X1 U11385 ( .A1(n11515), .A2(n11514), .ZN(n11532) );
  AND2_X1 U11386 ( .A1(n11512), .A2(n11533), .ZN(n11531) );
  OR2_X1 U11387 ( .A1(n11515), .A2(n11514), .ZN(n11533) );
  OR2_X1 U11388 ( .A1(n11534), .A2(n11535), .ZN(n11514) );
  AND2_X1 U11389 ( .A1(n11511), .A2(n11510), .ZN(n11535) );
  AND2_X1 U11390 ( .A1(n11508), .A2(n11536), .ZN(n11534) );
  OR2_X1 U11391 ( .A1(n11511), .A2(n11510), .ZN(n11536) );
  OR2_X1 U11392 ( .A1(n11537), .A2(n11538), .ZN(n11510) );
  AND2_X1 U11393 ( .A1(n11507), .A2(n11506), .ZN(n11538) );
  AND2_X1 U11394 ( .A1(n11504), .A2(n11539), .ZN(n11537) );
  OR2_X1 U11395 ( .A1(n11507), .A2(n11506), .ZN(n11539) );
  OR2_X1 U11396 ( .A1(n11540), .A2(n11541), .ZN(n11506) );
  AND2_X1 U11397 ( .A1(n11503), .A2(n11502), .ZN(n11541) );
  AND2_X1 U11398 ( .A1(n11500), .A2(n11542), .ZN(n11540) );
  OR2_X1 U11399 ( .A1(n11503), .A2(n11502), .ZN(n11542) );
  OR2_X1 U11400 ( .A1(n11543), .A2(n11544), .ZN(n11502) );
  AND2_X1 U11401 ( .A1(n11499), .A2(n11498), .ZN(n11544) );
  AND2_X1 U11402 ( .A1(n11496), .A2(n11545), .ZN(n11543) );
  OR2_X1 U11403 ( .A1(n11499), .A2(n11498), .ZN(n11545) );
  OR2_X1 U11404 ( .A1(n11546), .A2(n11547), .ZN(n11498) );
  AND2_X1 U11405 ( .A1(n11495), .A2(n11494), .ZN(n11547) );
  AND2_X1 U11406 ( .A1(n11492), .A2(n11548), .ZN(n11546) );
  OR2_X1 U11407 ( .A1(n11495), .A2(n11494), .ZN(n11548) );
  OR2_X1 U11408 ( .A1(n11549), .A2(n11550), .ZN(n11494) );
  AND2_X1 U11409 ( .A1(n11491), .A2(n11490), .ZN(n11550) );
  AND2_X1 U11410 ( .A1(n11488), .A2(n11551), .ZN(n11549) );
  OR2_X1 U11411 ( .A1(n11491), .A2(n11490), .ZN(n11551) );
  OR2_X1 U11412 ( .A1(n11552), .A2(n11553), .ZN(n11490) );
  AND2_X1 U11413 ( .A1(n11487), .A2(n11486), .ZN(n11553) );
  AND2_X1 U11414 ( .A1(n11484), .A2(n11554), .ZN(n11552) );
  OR2_X1 U11415 ( .A1(n11487), .A2(n11486), .ZN(n11554) );
  OR2_X1 U11416 ( .A1(n11555), .A2(n11556), .ZN(n11486) );
  AND2_X1 U11417 ( .A1(n11483), .A2(n11482), .ZN(n11556) );
  AND2_X1 U11418 ( .A1(n11480), .A2(n11557), .ZN(n11555) );
  OR2_X1 U11419 ( .A1(n11483), .A2(n11482), .ZN(n11557) );
  OR2_X1 U11420 ( .A1(n11558), .A2(n11559), .ZN(n11482) );
  AND2_X1 U11421 ( .A1(n11479), .A2(n11478), .ZN(n11559) );
  AND2_X1 U11422 ( .A1(n11476), .A2(n11560), .ZN(n11558) );
  OR2_X1 U11423 ( .A1(n11479), .A2(n11478), .ZN(n11560) );
  OR2_X1 U11424 ( .A1(n11561), .A2(n11562), .ZN(n11478) );
  AND2_X1 U11425 ( .A1(n11475), .A2(n11474), .ZN(n11562) );
  AND2_X1 U11426 ( .A1(n11472), .A2(n11563), .ZN(n11561) );
  OR2_X1 U11427 ( .A1(n11475), .A2(n11474), .ZN(n11563) );
  OR2_X1 U11428 ( .A1(n11564), .A2(n11565), .ZN(n11474) );
  AND2_X1 U11429 ( .A1(n11471), .A2(n11470), .ZN(n11565) );
  AND2_X1 U11430 ( .A1(n11468), .A2(n11566), .ZN(n11564) );
  OR2_X1 U11431 ( .A1(n11471), .A2(n11470), .ZN(n11566) );
  OR2_X1 U11432 ( .A1(n11567), .A2(n11568), .ZN(n11470) );
  AND2_X1 U11433 ( .A1(n11467), .A2(n11466), .ZN(n11568) );
  AND2_X1 U11434 ( .A1(n11464), .A2(n11569), .ZN(n11567) );
  OR2_X1 U11435 ( .A1(n11467), .A2(n11466), .ZN(n11569) );
  OR2_X1 U11436 ( .A1(n11570), .A2(n11571), .ZN(n11466) );
  AND2_X1 U11437 ( .A1(n8095), .A2(n11463), .ZN(n11571) );
  AND2_X1 U11438 ( .A1(n11461), .A2(n11572), .ZN(n11570) );
  OR2_X1 U11439 ( .A1(n8095), .A2(n11463), .ZN(n11572) );
  OR2_X1 U11440 ( .A1(n11573), .A2(n11574), .ZN(n11463) );
  AND2_X1 U11441 ( .A1(n11460), .A2(n11459), .ZN(n11574) );
  AND2_X1 U11442 ( .A1(n11457), .A2(n11575), .ZN(n11573) );
  OR2_X1 U11443 ( .A1(n11460), .A2(n11459), .ZN(n11575) );
  OR2_X1 U11444 ( .A1(n11576), .A2(n11577), .ZN(n11459) );
  AND2_X1 U11445 ( .A1(n11456), .A2(n11455), .ZN(n11577) );
  AND2_X1 U11446 ( .A1(n11453), .A2(n11578), .ZN(n11576) );
  OR2_X1 U11447 ( .A1(n11456), .A2(n11455), .ZN(n11578) );
  OR2_X1 U11448 ( .A1(n11579), .A2(n11580), .ZN(n11455) );
  AND2_X1 U11449 ( .A1(n11452), .A2(n11451), .ZN(n11580) );
  AND2_X1 U11450 ( .A1(n11449), .A2(n11581), .ZN(n11579) );
  OR2_X1 U11451 ( .A1(n11452), .A2(n11451), .ZN(n11581) );
  OR2_X1 U11452 ( .A1(n11582), .A2(n11583), .ZN(n11451) );
  AND2_X1 U11453 ( .A1(n11448), .A2(n11447), .ZN(n11583) );
  AND2_X1 U11454 ( .A1(n11445), .A2(n11584), .ZN(n11582) );
  OR2_X1 U11455 ( .A1(n11448), .A2(n11447), .ZN(n11584) );
  OR2_X1 U11456 ( .A1(n11585), .A2(n11586), .ZN(n11447) );
  AND2_X1 U11457 ( .A1(n11444), .A2(n11443), .ZN(n11586) );
  AND2_X1 U11458 ( .A1(n11441), .A2(n11587), .ZN(n11585) );
  OR2_X1 U11459 ( .A1(n11444), .A2(n11443), .ZN(n11587) );
  OR2_X1 U11460 ( .A1(n11588), .A2(n11589), .ZN(n11443) );
  AND2_X1 U11461 ( .A1(n11440), .A2(n11439), .ZN(n11589) );
  AND2_X1 U11462 ( .A1(n11437), .A2(n11590), .ZN(n11588) );
  OR2_X1 U11463 ( .A1(n11440), .A2(n11439), .ZN(n11590) );
  OR2_X1 U11464 ( .A1(n11591), .A2(n11592), .ZN(n11439) );
  AND2_X1 U11465 ( .A1(n11436), .A2(n11435), .ZN(n11592) );
  AND2_X1 U11466 ( .A1(n11433), .A2(n11593), .ZN(n11591) );
  OR2_X1 U11467 ( .A1(n11436), .A2(n11435), .ZN(n11593) );
  OR2_X1 U11468 ( .A1(n11594), .A2(n11595), .ZN(n11435) );
  AND2_X1 U11469 ( .A1(n11432), .A2(n11431), .ZN(n11595) );
  AND2_X1 U11470 ( .A1(n11429), .A2(n11596), .ZN(n11594) );
  OR2_X1 U11471 ( .A1(n11432), .A2(n11431), .ZN(n11596) );
  OR2_X1 U11472 ( .A1(n11597), .A2(n11598), .ZN(n11431) );
  AND2_X1 U11473 ( .A1(n11428), .A2(n11427), .ZN(n11598) );
  AND2_X1 U11474 ( .A1(n11425), .A2(n11599), .ZN(n11597) );
  OR2_X1 U11475 ( .A1(n11428), .A2(n11427), .ZN(n11599) );
  OR2_X1 U11476 ( .A1(n11600), .A2(n11601), .ZN(n11427) );
  AND2_X1 U11477 ( .A1(n11421), .A2(n11424), .ZN(n11601) );
  AND2_X1 U11478 ( .A1(n11602), .A2(n11603), .ZN(n11600) );
  OR2_X1 U11479 ( .A1(n11421), .A2(n11424), .ZN(n11603) );
  OR3_X1 U11480 ( .A1(n8094), .A2(n8981), .A3(n8089), .ZN(n11424) );
  OR2_X1 U11481 ( .A1(n8094), .A2(n8127), .ZN(n11421) );
  INV_X1 U11482 ( .A(n11423), .ZN(n11602) );
  OR2_X1 U11483 ( .A1(n11604), .A2(n11605), .ZN(n11423) );
  AND2_X1 U11484 ( .A1(b_18_), .A2(n11606), .ZN(n11605) );
  OR2_X1 U11485 ( .A1(n11607), .A2(n7598), .ZN(n11606) );
  AND2_X1 U11486 ( .A1(a_30_), .A2(n8085), .ZN(n11607) );
  AND2_X1 U11487 ( .A1(b_17_), .A2(n11608), .ZN(n11604) );
  OR2_X1 U11488 ( .A1(n11609), .A2(n7601), .ZN(n11608) );
  AND2_X1 U11489 ( .A1(a_31_), .A2(n8089), .ZN(n11609) );
  OR2_X1 U11490 ( .A1(n8094), .A2(n8124), .ZN(n11428) );
  XNOR2_X1 U11491 ( .A(n11610), .B(n11611), .ZN(n11425) );
  XOR2_X1 U11492 ( .A(n11612), .B(n11613), .Z(n11611) );
  OR2_X1 U11493 ( .A1(n8094), .A2(n8121), .ZN(n11432) );
  XOR2_X1 U11494 ( .A(n11614), .B(n11615), .Z(n11429) );
  XOR2_X1 U11495 ( .A(n11616), .B(n11617), .Z(n11615) );
  OR2_X1 U11496 ( .A1(n8094), .A2(n8118), .ZN(n11436) );
  XOR2_X1 U11497 ( .A(n11618), .B(n11619), .Z(n11433) );
  XOR2_X1 U11498 ( .A(n11620), .B(n11621), .Z(n11619) );
  OR2_X1 U11499 ( .A1(n8094), .A2(n8115), .ZN(n11440) );
  XOR2_X1 U11500 ( .A(n11622), .B(n11623), .Z(n11437) );
  XOR2_X1 U11501 ( .A(n11624), .B(n11625), .Z(n11623) );
  OR2_X1 U11502 ( .A1(n8094), .A2(n8112), .ZN(n11444) );
  XOR2_X1 U11503 ( .A(n11626), .B(n11627), .Z(n11441) );
  XOR2_X1 U11504 ( .A(n11628), .B(n11629), .Z(n11627) );
  OR2_X1 U11505 ( .A1(n8094), .A2(n8109), .ZN(n11448) );
  XOR2_X1 U11506 ( .A(n11630), .B(n11631), .Z(n11445) );
  XOR2_X1 U11507 ( .A(n11632), .B(n11633), .Z(n11631) );
  OR2_X1 U11508 ( .A1(n8094), .A2(n8106), .ZN(n11452) );
  XOR2_X1 U11509 ( .A(n11634), .B(n11635), .Z(n11449) );
  XOR2_X1 U11510 ( .A(n11636), .B(n11637), .Z(n11635) );
  OR2_X1 U11511 ( .A1(n8094), .A2(n8102), .ZN(n11456) );
  XOR2_X1 U11512 ( .A(n11638), .B(n11639), .Z(n11453) );
  XOR2_X1 U11513 ( .A(n11640), .B(n11641), .Z(n11639) );
  OR2_X1 U11514 ( .A1(n8094), .A2(n8097), .ZN(n11460) );
  XOR2_X1 U11515 ( .A(n11642), .B(n11643), .Z(n11457) );
  XOR2_X1 U11516 ( .A(n11644), .B(n11645), .Z(n11643) );
  OR2_X1 U11517 ( .A1(n8093), .A2(n8094), .ZN(n8095) );
  XOR2_X1 U11518 ( .A(n11646), .B(n11647), .Z(n11461) );
  XOR2_X1 U11519 ( .A(n11648), .B(n11649), .Z(n11647) );
  OR2_X1 U11520 ( .A1(n8094), .A2(n8088), .ZN(n11467) );
  XOR2_X1 U11521 ( .A(n11650), .B(n11651), .Z(n11464) );
  XOR2_X1 U11522 ( .A(n11652), .B(n11653), .Z(n11651) );
  OR2_X1 U11523 ( .A1(n8084), .A2(n8094), .ZN(n11471) );
  XNOR2_X1 U11524 ( .A(n11654), .B(n11655), .ZN(n11468) );
  XOR2_X1 U11525 ( .A(n7782), .B(n11656), .Z(n11654) );
  INV_X1 U11526 ( .A(n8090), .ZN(n7782) );
  OR2_X1 U11527 ( .A1(n8094), .A2(n8079), .ZN(n11475) );
  XOR2_X1 U11528 ( .A(n11657), .B(n11658), .Z(n11472) );
  XOR2_X1 U11529 ( .A(n11659), .B(n11660), .Z(n11658) );
  OR2_X1 U11530 ( .A1(n8075), .A2(n8094), .ZN(n11479) );
  XOR2_X1 U11531 ( .A(n11661), .B(n11662), .Z(n11476) );
  XOR2_X1 U11532 ( .A(n11663), .B(n11664), .Z(n11662) );
  OR2_X1 U11533 ( .A1(n8094), .A2(n8070), .ZN(n11483) );
  XOR2_X1 U11534 ( .A(n11665), .B(n11666), .Z(n11480) );
  XOR2_X1 U11535 ( .A(n11667), .B(n11668), .Z(n11666) );
  OR2_X1 U11536 ( .A1(n8066), .A2(n8094), .ZN(n11487) );
  XOR2_X1 U11537 ( .A(n11669), .B(n11670), .Z(n11484) );
  XOR2_X1 U11538 ( .A(n11671), .B(n11672), .Z(n11670) );
  OR2_X1 U11539 ( .A1(n8094), .A2(n8061), .ZN(n11491) );
  XOR2_X1 U11540 ( .A(n11673), .B(n11674), .Z(n11488) );
  XOR2_X1 U11541 ( .A(n11675), .B(n11676), .Z(n11674) );
  OR2_X1 U11542 ( .A1(n8057), .A2(n8094), .ZN(n11495) );
  XOR2_X1 U11543 ( .A(n11677), .B(n11678), .Z(n11492) );
  XOR2_X1 U11544 ( .A(n11679), .B(n11680), .Z(n11678) );
  OR2_X1 U11545 ( .A1(n8094), .A2(n8052), .ZN(n11499) );
  XOR2_X1 U11546 ( .A(n11681), .B(n11682), .Z(n11496) );
  XOR2_X1 U11547 ( .A(n11683), .B(n11684), .Z(n11682) );
  OR2_X1 U11548 ( .A1(n8048), .A2(n8094), .ZN(n11503) );
  XOR2_X1 U11549 ( .A(n11685), .B(n11686), .Z(n11500) );
  XOR2_X1 U11550 ( .A(n11687), .B(n11688), .Z(n11686) );
  OR2_X1 U11551 ( .A1(n8094), .A2(n8043), .ZN(n11507) );
  XOR2_X1 U11552 ( .A(n11689), .B(n11690), .Z(n11504) );
  XOR2_X1 U11553 ( .A(n11691), .B(n11692), .Z(n11690) );
  OR2_X1 U11554 ( .A1(n8039), .A2(n8094), .ZN(n11511) );
  XOR2_X1 U11555 ( .A(n11693), .B(n11694), .Z(n11508) );
  XOR2_X1 U11556 ( .A(n11695), .B(n11696), .Z(n11694) );
  OR2_X1 U11557 ( .A1(n8094), .A2(n8034), .ZN(n11515) );
  XOR2_X1 U11558 ( .A(n11697), .B(n11698), .Z(n11512) );
  XOR2_X1 U11559 ( .A(n11699), .B(n11700), .Z(n11698) );
  OR2_X1 U11560 ( .A1(n8030), .A2(n8094), .ZN(n11519) );
  XOR2_X1 U11561 ( .A(n11701), .B(n11702), .Z(n11516) );
  XOR2_X1 U11562 ( .A(n11703), .B(n11704), .Z(n11702) );
  OR2_X1 U11563 ( .A1(n8094), .A2(n8025), .ZN(n11523) );
  XOR2_X1 U11564 ( .A(n11705), .B(n11706), .Z(n11520) );
  XOR2_X1 U11565 ( .A(n11707), .B(n11708), .Z(n11706) );
  XOR2_X1 U11566 ( .A(n10898), .B(n11709), .Z(n10891) );
  XOR2_X1 U11567 ( .A(n10897), .B(n10896), .Z(n11709) );
  OR2_X1 U11568 ( .A1(n8089), .A2(n8025), .ZN(n10896) );
  OR2_X1 U11569 ( .A1(n11710), .A2(n11711), .ZN(n10897) );
  AND2_X1 U11570 ( .A1(n11708), .A2(n11707), .ZN(n11711) );
  AND2_X1 U11571 ( .A1(n11705), .A2(n11712), .ZN(n11710) );
  OR2_X1 U11572 ( .A1(n11708), .A2(n11707), .ZN(n11712) );
  OR2_X1 U11573 ( .A1(n11713), .A2(n11714), .ZN(n11707) );
  AND2_X1 U11574 ( .A1(n11704), .A2(n11703), .ZN(n11714) );
  AND2_X1 U11575 ( .A1(n11701), .A2(n11715), .ZN(n11713) );
  OR2_X1 U11576 ( .A1(n11704), .A2(n11703), .ZN(n11715) );
  OR2_X1 U11577 ( .A1(n11716), .A2(n11717), .ZN(n11703) );
  AND2_X1 U11578 ( .A1(n11700), .A2(n11699), .ZN(n11717) );
  AND2_X1 U11579 ( .A1(n11697), .A2(n11718), .ZN(n11716) );
  OR2_X1 U11580 ( .A1(n11700), .A2(n11699), .ZN(n11718) );
  OR2_X1 U11581 ( .A1(n11719), .A2(n11720), .ZN(n11699) );
  AND2_X1 U11582 ( .A1(n11696), .A2(n11695), .ZN(n11720) );
  AND2_X1 U11583 ( .A1(n11693), .A2(n11721), .ZN(n11719) );
  OR2_X1 U11584 ( .A1(n11696), .A2(n11695), .ZN(n11721) );
  OR2_X1 U11585 ( .A1(n11722), .A2(n11723), .ZN(n11695) );
  AND2_X1 U11586 ( .A1(n11692), .A2(n11691), .ZN(n11723) );
  AND2_X1 U11587 ( .A1(n11689), .A2(n11724), .ZN(n11722) );
  OR2_X1 U11588 ( .A1(n11692), .A2(n11691), .ZN(n11724) );
  OR2_X1 U11589 ( .A1(n11725), .A2(n11726), .ZN(n11691) );
  AND2_X1 U11590 ( .A1(n11688), .A2(n11687), .ZN(n11726) );
  AND2_X1 U11591 ( .A1(n11685), .A2(n11727), .ZN(n11725) );
  OR2_X1 U11592 ( .A1(n11688), .A2(n11687), .ZN(n11727) );
  OR2_X1 U11593 ( .A1(n11728), .A2(n11729), .ZN(n11687) );
  AND2_X1 U11594 ( .A1(n11684), .A2(n11683), .ZN(n11729) );
  AND2_X1 U11595 ( .A1(n11681), .A2(n11730), .ZN(n11728) );
  OR2_X1 U11596 ( .A1(n11684), .A2(n11683), .ZN(n11730) );
  OR2_X1 U11597 ( .A1(n11731), .A2(n11732), .ZN(n11683) );
  AND2_X1 U11598 ( .A1(n11680), .A2(n11679), .ZN(n11732) );
  AND2_X1 U11599 ( .A1(n11677), .A2(n11733), .ZN(n11731) );
  OR2_X1 U11600 ( .A1(n11680), .A2(n11679), .ZN(n11733) );
  OR2_X1 U11601 ( .A1(n11734), .A2(n11735), .ZN(n11679) );
  AND2_X1 U11602 ( .A1(n11676), .A2(n11675), .ZN(n11735) );
  AND2_X1 U11603 ( .A1(n11673), .A2(n11736), .ZN(n11734) );
  OR2_X1 U11604 ( .A1(n11676), .A2(n11675), .ZN(n11736) );
  OR2_X1 U11605 ( .A1(n11737), .A2(n11738), .ZN(n11675) );
  AND2_X1 U11606 ( .A1(n11672), .A2(n11671), .ZN(n11738) );
  AND2_X1 U11607 ( .A1(n11669), .A2(n11739), .ZN(n11737) );
  OR2_X1 U11608 ( .A1(n11672), .A2(n11671), .ZN(n11739) );
  OR2_X1 U11609 ( .A1(n11740), .A2(n11741), .ZN(n11671) );
  AND2_X1 U11610 ( .A1(n11668), .A2(n11667), .ZN(n11741) );
  AND2_X1 U11611 ( .A1(n11665), .A2(n11742), .ZN(n11740) );
  OR2_X1 U11612 ( .A1(n11668), .A2(n11667), .ZN(n11742) );
  OR2_X1 U11613 ( .A1(n11743), .A2(n11744), .ZN(n11667) );
  AND2_X1 U11614 ( .A1(n11664), .A2(n11663), .ZN(n11744) );
  AND2_X1 U11615 ( .A1(n11661), .A2(n11745), .ZN(n11743) );
  OR2_X1 U11616 ( .A1(n11664), .A2(n11663), .ZN(n11745) );
  OR2_X1 U11617 ( .A1(n11746), .A2(n11747), .ZN(n11663) );
  AND2_X1 U11618 ( .A1(n11660), .A2(n11659), .ZN(n11747) );
  AND2_X1 U11619 ( .A1(n11657), .A2(n11748), .ZN(n11746) );
  OR2_X1 U11620 ( .A1(n11660), .A2(n11659), .ZN(n11748) );
  OR2_X1 U11621 ( .A1(n11749), .A2(n11750), .ZN(n11659) );
  AND2_X1 U11622 ( .A1(n11656), .A2(n8090), .ZN(n11750) );
  AND2_X1 U11623 ( .A1(n11655), .A2(n11751), .ZN(n11749) );
  OR2_X1 U11624 ( .A1(n11656), .A2(n8090), .ZN(n11751) );
  OR2_X1 U11625 ( .A1(n8088), .A2(n8089), .ZN(n8090) );
  OR2_X1 U11626 ( .A1(n11752), .A2(n11753), .ZN(n11656) );
  AND2_X1 U11627 ( .A1(n11653), .A2(n11652), .ZN(n11753) );
  AND2_X1 U11628 ( .A1(n11650), .A2(n11754), .ZN(n11752) );
  OR2_X1 U11629 ( .A1(n11653), .A2(n11652), .ZN(n11754) );
  OR2_X1 U11630 ( .A1(n11755), .A2(n11756), .ZN(n11652) );
  AND2_X1 U11631 ( .A1(n11649), .A2(n11648), .ZN(n11756) );
  AND2_X1 U11632 ( .A1(n11646), .A2(n11757), .ZN(n11755) );
  OR2_X1 U11633 ( .A1(n11649), .A2(n11648), .ZN(n11757) );
  OR2_X1 U11634 ( .A1(n11758), .A2(n11759), .ZN(n11648) );
  AND2_X1 U11635 ( .A1(n11645), .A2(n11644), .ZN(n11759) );
  AND2_X1 U11636 ( .A1(n11642), .A2(n11760), .ZN(n11758) );
  OR2_X1 U11637 ( .A1(n11645), .A2(n11644), .ZN(n11760) );
  OR2_X1 U11638 ( .A1(n11761), .A2(n11762), .ZN(n11644) );
  AND2_X1 U11639 ( .A1(n11641), .A2(n11640), .ZN(n11762) );
  AND2_X1 U11640 ( .A1(n11638), .A2(n11763), .ZN(n11761) );
  OR2_X1 U11641 ( .A1(n11641), .A2(n11640), .ZN(n11763) );
  OR2_X1 U11642 ( .A1(n11764), .A2(n11765), .ZN(n11640) );
  AND2_X1 U11643 ( .A1(n11637), .A2(n11636), .ZN(n11765) );
  AND2_X1 U11644 ( .A1(n11634), .A2(n11766), .ZN(n11764) );
  OR2_X1 U11645 ( .A1(n11637), .A2(n11636), .ZN(n11766) );
  OR2_X1 U11646 ( .A1(n11767), .A2(n11768), .ZN(n11636) );
  AND2_X1 U11647 ( .A1(n11633), .A2(n11632), .ZN(n11768) );
  AND2_X1 U11648 ( .A1(n11630), .A2(n11769), .ZN(n11767) );
  OR2_X1 U11649 ( .A1(n11633), .A2(n11632), .ZN(n11769) );
  OR2_X1 U11650 ( .A1(n11770), .A2(n11771), .ZN(n11632) );
  AND2_X1 U11651 ( .A1(n11629), .A2(n11628), .ZN(n11771) );
  AND2_X1 U11652 ( .A1(n11626), .A2(n11772), .ZN(n11770) );
  OR2_X1 U11653 ( .A1(n11629), .A2(n11628), .ZN(n11772) );
  OR2_X1 U11654 ( .A1(n11773), .A2(n11774), .ZN(n11628) );
  AND2_X1 U11655 ( .A1(n11625), .A2(n11624), .ZN(n11774) );
  AND2_X1 U11656 ( .A1(n11622), .A2(n11775), .ZN(n11773) );
  OR2_X1 U11657 ( .A1(n11625), .A2(n11624), .ZN(n11775) );
  OR2_X1 U11658 ( .A1(n11776), .A2(n11777), .ZN(n11624) );
  AND2_X1 U11659 ( .A1(n11621), .A2(n11620), .ZN(n11777) );
  AND2_X1 U11660 ( .A1(n11618), .A2(n11778), .ZN(n11776) );
  OR2_X1 U11661 ( .A1(n11621), .A2(n11620), .ZN(n11778) );
  OR2_X1 U11662 ( .A1(n11779), .A2(n11780), .ZN(n11620) );
  AND2_X1 U11663 ( .A1(n11617), .A2(n11616), .ZN(n11780) );
  AND2_X1 U11664 ( .A1(n11614), .A2(n11781), .ZN(n11779) );
  OR2_X1 U11665 ( .A1(n11617), .A2(n11616), .ZN(n11781) );
  OR2_X1 U11666 ( .A1(n11782), .A2(n11783), .ZN(n11616) );
  AND2_X1 U11667 ( .A1(n11610), .A2(n11613), .ZN(n11783) );
  AND2_X1 U11668 ( .A1(n11784), .A2(n11785), .ZN(n11782) );
  OR2_X1 U11669 ( .A1(n11610), .A2(n11613), .ZN(n11785) );
  OR3_X1 U11670 ( .A1(n8085), .A2(n8981), .A3(n8089), .ZN(n11613) );
  OR2_X1 U11671 ( .A1(n8127), .A2(n8089), .ZN(n11610) );
  INV_X1 U11672 ( .A(n11612), .ZN(n11784) );
  OR2_X1 U11673 ( .A1(n11786), .A2(n11787), .ZN(n11612) );
  AND2_X1 U11674 ( .A1(b_17_), .A2(n11788), .ZN(n11787) );
  OR2_X1 U11675 ( .A1(n11789), .A2(n7598), .ZN(n11788) );
  AND2_X1 U11676 ( .A1(a_30_), .A2(n8080), .ZN(n11789) );
  AND2_X1 U11677 ( .A1(b_16_), .A2(n11790), .ZN(n11786) );
  OR2_X1 U11678 ( .A1(n11791), .A2(n7601), .ZN(n11790) );
  AND2_X1 U11679 ( .A1(a_31_), .A2(n8085), .ZN(n11791) );
  OR2_X1 U11680 ( .A1(n8124), .A2(n8089), .ZN(n11617) );
  XNOR2_X1 U11681 ( .A(n11792), .B(n11793), .ZN(n11614) );
  XOR2_X1 U11682 ( .A(n11794), .B(n11795), .Z(n11793) );
  OR2_X1 U11683 ( .A1(n8121), .A2(n8089), .ZN(n11621) );
  XOR2_X1 U11684 ( .A(n11796), .B(n11797), .Z(n11618) );
  XOR2_X1 U11685 ( .A(n11798), .B(n11799), .Z(n11797) );
  OR2_X1 U11686 ( .A1(n8118), .A2(n8089), .ZN(n11625) );
  XOR2_X1 U11687 ( .A(n11800), .B(n11801), .Z(n11622) );
  XOR2_X1 U11688 ( .A(n11802), .B(n11803), .Z(n11801) );
  OR2_X1 U11689 ( .A1(n8115), .A2(n8089), .ZN(n11629) );
  XOR2_X1 U11690 ( .A(n11804), .B(n11805), .Z(n11626) );
  XOR2_X1 U11691 ( .A(n11806), .B(n11807), .Z(n11805) );
  OR2_X1 U11692 ( .A1(n8112), .A2(n8089), .ZN(n11633) );
  XOR2_X1 U11693 ( .A(n11808), .B(n11809), .Z(n11630) );
  XOR2_X1 U11694 ( .A(n11810), .B(n11811), .Z(n11809) );
  OR2_X1 U11695 ( .A1(n8109), .A2(n8089), .ZN(n11637) );
  XOR2_X1 U11696 ( .A(n11812), .B(n11813), .Z(n11634) );
  XOR2_X1 U11697 ( .A(n11814), .B(n11815), .Z(n11813) );
  OR2_X1 U11698 ( .A1(n8106), .A2(n8089), .ZN(n11641) );
  XOR2_X1 U11699 ( .A(n11816), .B(n11817), .Z(n11638) );
  XOR2_X1 U11700 ( .A(n11818), .B(n11819), .Z(n11817) );
  OR2_X1 U11701 ( .A1(n8102), .A2(n8089), .ZN(n11645) );
  XOR2_X1 U11702 ( .A(n11820), .B(n11821), .Z(n11642) );
  XOR2_X1 U11703 ( .A(n11822), .B(n11823), .Z(n11821) );
  OR2_X1 U11704 ( .A1(n8097), .A2(n8089), .ZN(n11649) );
  XOR2_X1 U11705 ( .A(n11824), .B(n11825), .Z(n11646) );
  XOR2_X1 U11706 ( .A(n11826), .B(n11827), .Z(n11825) );
  OR2_X1 U11707 ( .A1(n8093), .A2(n8089), .ZN(n11653) );
  XOR2_X1 U11708 ( .A(n11828), .B(n11829), .Z(n11650) );
  XOR2_X1 U11709 ( .A(n11830), .B(n11831), .Z(n11829) );
  XOR2_X1 U11710 ( .A(n11832), .B(n11833), .Z(n11655) );
  XOR2_X1 U11711 ( .A(n11834), .B(n11835), .Z(n11833) );
  OR2_X1 U11712 ( .A1(n8084), .A2(n8089), .ZN(n11660) );
  XOR2_X1 U11713 ( .A(n11836), .B(n11837), .Z(n11657) );
  XOR2_X1 U11714 ( .A(n11838), .B(n11839), .Z(n11837) );
  OR2_X1 U11715 ( .A1(n8089), .A2(n8079), .ZN(n11664) );
  XOR2_X1 U11716 ( .A(n11840), .B(n11841), .Z(n11661) );
  XOR2_X1 U11717 ( .A(n11842), .B(n8086), .Z(n11841) );
  OR2_X1 U11718 ( .A1(n8075), .A2(n8089), .ZN(n11668) );
  XOR2_X1 U11719 ( .A(n11843), .B(n11844), .Z(n11665) );
  XOR2_X1 U11720 ( .A(n11845), .B(n11846), .Z(n11844) );
  OR2_X1 U11721 ( .A1(n8089), .A2(n8070), .ZN(n11672) );
  XOR2_X1 U11722 ( .A(n11847), .B(n11848), .Z(n11669) );
  XOR2_X1 U11723 ( .A(n11849), .B(n11850), .Z(n11848) );
  OR2_X1 U11724 ( .A1(n8066), .A2(n8089), .ZN(n11676) );
  XOR2_X1 U11725 ( .A(n11851), .B(n11852), .Z(n11673) );
  XOR2_X1 U11726 ( .A(n11853), .B(n11854), .Z(n11852) );
  OR2_X1 U11727 ( .A1(n8089), .A2(n8061), .ZN(n11680) );
  XOR2_X1 U11728 ( .A(n11855), .B(n11856), .Z(n11677) );
  XOR2_X1 U11729 ( .A(n11857), .B(n11858), .Z(n11856) );
  OR2_X1 U11730 ( .A1(n8057), .A2(n8089), .ZN(n11684) );
  XOR2_X1 U11731 ( .A(n11859), .B(n11860), .Z(n11681) );
  XOR2_X1 U11732 ( .A(n11861), .B(n11862), .Z(n11860) );
  OR2_X1 U11733 ( .A1(n8089), .A2(n8052), .ZN(n11688) );
  XOR2_X1 U11734 ( .A(n11863), .B(n11864), .Z(n11685) );
  XOR2_X1 U11735 ( .A(n11865), .B(n11866), .Z(n11864) );
  OR2_X1 U11736 ( .A1(n8048), .A2(n8089), .ZN(n11692) );
  XOR2_X1 U11737 ( .A(n11867), .B(n11868), .Z(n11689) );
  XOR2_X1 U11738 ( .A(n11869), .B(n11870), .Z(n11868) );
  OR2_X1 U11739 ( .A1(n8089), .A2(n8043), .ZN(n11696) );
  XOR2_X1 U11740 ( .A(n11871), .B(n11872), .Z(n11693) );
  XOR2_X1 U11741 ( .A(n11873), .B(n11874), .Z(n11872) );
  OR2_X1 U11742 ( .A1(n8039), .A2(n8089), .ZN(n11700) );
  XOR2_X1 U11743 ( .A(n11875), .B(n11876), .Z(n11697) );
  XOR2_X1 U11744 ( .A(n11877), .B(n11878), .Z(n11876) );
  OR2_X1 U11745 ( .A1(n8089), .A2(n8034), .ZN(n11704) );
  XOR2_X1 U11746 ( .A(n11879), .B(n11880), .Z(n11701) );
  XOR2_X1 U11747 ( .A(n11881), .B(n11882), .Z(n11880) );
  OR2_X1 U11748 ( .A1(n8030), .A2(n8089), .ZN(n11708) );
  INV_X1 U11749 ( .A(b_18_), .ZN(n8089) );
  XOR2_X1 U11750 ( .A(n11883), .B(n11884), .Z(n11705) );
  XOR2_X1 U11751 ( .A(n11885), .B(n11886), .Z(n11884) );
  XOR2_X1 U11752 ( .A(n10905), .B(n11887), .Z(n10898) );
  XOR2_X1 U11753 ( .A(n10904), .B(n10903), .Z(n11887) );
  OR2_X1 U11754 ( .A1(n8030), .A2(n8085), .ZN(n10903) );
  OR2_X1 U11755 ( .A1(n11888), .A2(n11889), .ZN(n10904) );
  AND2_X1 U11756 ( .A1(n11886), .A2(n11885), .ZN(n11889) );
  AND2_X1 U11757 ( .A1(n11883), .A2(n11890), .ZN(n11888) );
  OR2_X1 U11758 ( .A1(n11886), .A2(n11885), .ZN(n11890) );
  OR2_X1 U11759 ( .A1(n11891), .A2(n11892), .ZN(n11885) );
  AND2_X1 U11760 ( .A1(n11882), .A2(n11881), .ZN(n11892) );
  AND2_X1 U11761 ( .A1(n11879), .A2(n11893), .ZN(n11891) );
  OR2_X1 U11762 ( .A1(n11882), .A2(n11881), .ZN(n11893) );
  OR2_X1 U11763 ( .A1(n11894), .A2(n11895), .ZN(n11881) );
  AND2_X1 U11764 ( .A1(n11878), .A2(n11877), .ZN(n11895) );
  AND2_X1 U11765 ( .A1(n11875), .A2(n11896), .ZN(n11894) );
  OR2_X1 U11766 ( .A1(n11878), .A2(n11877), .ZN(n11896) );
  OR2_X1 U11767 ( .A1(n11897), .A2(n11898), .ZN(n11877) );
  AND2_X1 U11768 ( .A1(n11874), .A2(n11873), .ZN(n11898) );
  AND2_X1 U11769 ( .A1(n11871), .A2(n11899), .ZN(n11897) );
  OR2_X1 U11770 ( .A1(n11874), .A2(n11873), .ZN(n11899) );
  OR2_X1 U11771 ( .A1(n11900), .A2(n11901), .ZN(n11873) );
  AND2_X1 U11772 ( .A1(n11870), .A2(n11869), .ZN(n11901) );
  AND2_X1 U11773 ( .A1(n11867), .A2(n11902), .ZN(n11900) );
  OR2_X1 U11774 ( .A1(n11870), .A2(n11869), .ZN(n11902) );
  OR2_X1 U11775 ( .A1(n11903), .A2(n11904), .ZN(n11869) );
  AND2_X1 U11776 ( .A1(n11866), .A2(n11865), .ZN(n11904) );
  AND2_X1 U11777 ( .A1(n11863), .A2(n11905), .ZN(n11903) );
  OR2_X1 U11778 ( .A1(n11866), .A2(n11865), .ZN(n11905) );
  OR2_X1 U11779 ( .A1(n11906), .A2(n11907), .ZN(n11865) );
  AND2_X1 U11780 ( .A1(n11862), .A2(n11861), .ZN(n11907) );
  AND2_X1 U11781 ( .A1(n11859), .A2(n11908), .ZN(n11906) );
  OR2_X1 U11782 ( .A1(n11862), .A2(n11861), .ZN(n11908) );
  OR2_X1 U11783 ( .A1(n11909), .A2(n11910), .ZN(n11861) );
  AND2_X1 U11784 ( .A1(n11858), .A2(n11857), .ZN(n11910) );
  AND2_X1 U11785 ( .A1(n11855), .A2(n11911), .ZN(n11909) );
  OR2_X1 U11786 ( .A1(n11858), .A2(n11857), .ZN(n11911) );
  OR2_X1 U11787 ( .A1(n11912), .A2(n11913), .ZN(n11857) );
  AND2_X1 U11788 ( .A1(n11854), .A2(n11853), .ZN(n11913) );
  AND2_X1 U11789 ( .A1(n11851), .A2(n11914), .ZN(n11912) );
  OR2_X1 U11790 ( .A1(n11854), .A2(n11853), .ZN(n11914) );
  OR2_X1 U11791 ( .A1(n11915), .A2(n11916), .ZN(n11853) );
  AND2_X1 U11792 ( .A1(n11850), .A2(n11849), .ZN(n11916) );
  AND2_X1 U11793 ( .A1(n11847), .A2(n11917), .ZN(n11915) );
  OR2_X1 U11794 ( .A1(n11850), .A2(n11849), .ZN(n11917) );
  OR2_X1 U11795 ( .A1(n11918), .A2(n11919), .ZN(n11849) );
  AND2_X1 U11796 ( .A1(n11846), .A2(n11845), .ZN(n11919) );
  AND2_X1 U11797 ( .A1(n11843), .A2(n11920), .ZN(n11918) );
  OR2_X1 U11798 ( .A1(n11846), .A2(n11845), .ZN(n11920) );
  OR2_X1 U11799 ( .A1(n11921), .A2(n11922), .ZN(n11845) );
  AND2_X1 U11800 ( .A1(n8086), .A2(n11842), .ZN(n11922) );
  AND2_X1 U11801 ( .A1(n11840), .A2(n11923), .ZN(n11921) );
  OR2_X1 U11802 ( .A1(n8086), .A2(n11842), .ZN(n11923) );
  OR2_X1 U11803 ( .A1(n11924), .A2(n11925), .ZN(n11842) );
  AND2_X1 U11804 ( .A1(n11839), .A2(n11838), .ZN(n11925) );
  AND2_X1 U11805 ( .A1(n11836), .A2(n11926), .ZN(n11924) );
  OR2_X1 U11806 ( .A1(n11839), .A2(n11838), .ZN(n11926) );
  OR2_X1 U11807 ( .A1(n11927), .A2(n11928), .ZN(n11838) );
  AND2_X1 U11808 ( .A1(n11835), .A2(n11834), .ZN(n11928) );
  AND2_X1 U11809 ( .A1(n11832), .A2(n11929), .ZN(n11927) );
  OR2_X1 U11810 ( .A1(n11835), .A2(n11834), .ZN(n11929) );
  OR2_X1 U11811 ( .A1(n11930), .A2(n11931), .ZN(n11834) );
  AND2_X1 U11812 ( .A1(n11831), .A2(n11830), .ZN(n11931) );
  AND2_X1 U11813 ( .A1(n11828), .A2(n11932), .ZN(n11930) );
  OR2_X1 U11814 ( .A1(n11831), .A2(n11830), .ZN(n11932) );
  OR2_X1 U11815 ( .A1(n11933), .A2(n11934), .ZN(n11830) );
  AND2_X1 U11816 ( .A1(n11827), .A2(n11826), .ZN(n11934) );
  AND2_X1 U11817 ( .A1(n11824), .A2(n11935), .ZN(n11933) );
  OR2_X1 U11818 ( .A1(n11827), .A2(n11826), .ZN(n11935) );
  OR2_X1 U11819 ( .A1(n11936), .A2(n11937), .ZN(n11826) );
  AND2_X1 U11820 ( .A1(n11823), .A2(n11822), .ZN(n11937) );
  AND2_X1 U11821 ( .A1(n11820), .A2(n11938), .ZN(n11936) );
  OR2_X1 U11822 ( .A1(n11823), .A2(n11822), .ZN(n11938) );
  OR2_X1 U11823 ( .A1(n11939), .A2(n11940), .ZN(n11822) );
  AND2_X1 U11824 ( .A1(n11819), .A2(n11818), .ZN(n11940) );
  AND2_X1 U11825 ( .A1(n11816), .A2(n11941), .ZN(n11939) );
  OR2_X1 U11826 ( .A1(n11819), .A2(n11818), .ZN(n11941) );
  OR2_X1 U11827 ( .A1(n11942), .A2(n11943), .ZN(n11818) );
  AND2_X1 U11828 ( .A1(n11815), .A2(n11814), .ZN(n11943) );
  AND2_X1 U11829 ( .A1(n11812), .A2(n11944), .ZN(n11942) );
  OR2_X1 U11830 ( .A1(n11815), .A2(n11814), .ZN(n11944) );
  OR2_X1 U11831 ( .A1(n11945), .A2(n11946), .ZN(n11814) );
  AND2_X1 U11832 ( .A1(n11811), .A2(n11810), .ZN(n11946) );
  AND2_X1 U11833 ( .A1(n11808), .A2(n11947), .ZN(n11945) );
  OR2_X1 U11834 ( .A1(n11811), .A2(n11810), .ZN(n11947) );
  OR2_X1 U11835 ( .A1(n11948), .A2(n11949), .ZN(n11810) );
  AND2_X1 U11836 ( .A1(n11807), .A2(n11806), .ZN(n11949) );
  AND2_X1 U11837 ( .A1(n11804), .A2(n11950), .ZN(n11948) );
  OR2_X1 U11838 ( .A1(n11807), .A2(n11806), .ZN(n11950) );
  OR2_X1 U11839 ( .A1(n11951), .A2(n11952), .ZN(n11806) );
  AND2_X1 U11840 ( .A1(n11803), .A2(n11802), .ZN(n11952) );
  AND2_X1 U11841 ( .A1(n11800), .A2(n11953), .ZN(n11951) );
  OR2_X1 U11842 ( .A1(n11803), .A2(n11802), .ZN(n11953) );
  OR2_X1 U11843 ( .A1(n11954), .A2(n11955), .ZN(n11802) );
  AND2_X1 U11844 ( .A1(n11799), .A2(n11798), .ZN(n11955) );
  AND2_X1 U11845 ( .A1(n11796), .A2(n11956), .ZN(n11954) );
  OR2_X1 U11846 ( .A1(n11799), .A2(n11798), .ZN(n11956) );
  OR2_X1 U11847 ( .A1(n11957), .A2(n11958), .ZN(n11798) );
  AND2_X1 U11848 ( .A1(n11792), .A2(n11795), .ZN(n11958) );
  AND2_X1 U11849 ( .A1(n11959), .A2(n11960), .ZN(n11957) );
  OR2_X1 U11850 ( .A1(n11792), .A2(n11795), .ZN(n11960) );
  OR3_X1 U11851 ( .A1(n8080), .A2(n8085), .A3(n8981), .ZN(n11795) );
  OR2_X1 U11852 ( .A1(n8085), .A2(n8127), .ZN(n11792) );
  INV_X1 U11853 ( .A(n11794), .ZN(n11959) );
  OR2_X1 U11854 ( .A1(n11961), .A2(n11962), .ZN(n11794) );
  AND2_X1 U11855 ( .A1(b_16_), .A2(n11963), .ZN(n11962) );
  OR2_X1 U11856 ( .A1(n11964), .A2(n7598), .ZN(n11963) );
  AND2_X1 U11857 ( .A1(a_30_), .A2(n8076), .ZN(n11964) );
  AND2_X1 U11858 ( .A1(b_15_), .A2(n11965), .ZN(n11961) );
  OR2_X1 U11859 ( .A1(n11966), .A2(n7601), .ZN(n11965) );
  AND2_X1 U11860 ( .A1(a_31_), .A2(n8080), .ZN(n11966) );
  OR2_X1 U11861 ( .A1(n8085), .A2(n8124), .ZN(n11799) );
  XNOR2_X1 U11862 ( .A(n11967), .B(n11968), .ZN(n11796) );
  XOR2_X1 U11863 ( .A(n11969), .B(n11970), .Z(n11968) );
  OR2_X1 U11864 ( .A1(n8085), .A2(n8121), .ZN(n11803) );
  XOR2_X1 U11865 ( .A(n11971), .B(n11972), .Z(n11800) );
  XOR2_X1 U11866 ( .A(n11973), .B(n11974), .Z(n11972) );
  OR2_X1 U11867 ( .A1(n8085), .A2(n8118), .ZN(n11807) );
  XOR2_X1 U11868 ( .A(n11975), .B(n11976), .Z(n11804) );
  XOR2_X1 U11869 ( .A(n11977), .B(n11978), .Z(n11976) );
  OR2_X1 U11870 ( .A1(n8085), .A2(n8115), .ZN(n11811) );
  XOR2_X1 U11871 ( .A(n11979), .B(n11980), .Z(n11808) );
  XOR2_X1 U11872 ( .A(n11981), .B(n11982), .Z(n11980) );
  OR2_X1 U11873 ( .A1(n8085), .A2(n8112), .ZN(n11815) );
  XOR2_X1 U11874 ( .A(n11983), .B(n11984), .Z(n11812) );
  XOR2_X1 U11875 ( .A(n11985), .B(n11986), .Z(n11984) );
  OR2_X1 U11876 ( .A1(n8085), .A2(n8109), .ZN(n11819) );
  XOR2_X1 U11877 ( .A(n11987), .B(n11988), .Z(n11816) );
  XOR2_X1 U11878 ( .A(n11989), .B(n11990), .Z(n11988) );
  OR2_X1 U11879 ( .A1(n8085), .A2(n8106), .ZN(n11823) );
  XOR2_X1 U11880 ( .A(n11991), .B(n11992), .Z(n11820) );
  XOR2_X1 U11881 ( .A(n11993), .B(n11994), .Z(n11992) );
  OR2_X1 U11882 ( .A1(n8085), .A2(n8102), .ZN(n11827) );
  XOR2_X1 U11883 ( .A(n11995), .B(n11996), .Z(n11824) );
  XOR2_X1 U11884 ( .A(n11997), .B(n11998), .Z(n11996) );
  OR2_X1 U11885 ( .A1(n8085), .A2(n8097), .ZN(n11831) );
  XOR2_X1 U11886 ( .A(n11999), .B(n12000), .Z(n11828) );
  XOR2_X1 U11887 ( .A(n12001), .B(n12002), .Z(n12000) );
  OR2_X1 U11888 ( .A1(n8085), .A2(n8093), .ZN(n11835) );
  XOR2_X1 U11889 ( .A(n12003), .B(n12004), .Z(n11832) );
  XOR2_X1 U11890 ( .A(n12005), .B(n12006), .Z(n12004) );
  OR2_X1 U11891 ( .A1(n8085), .A2(n8088), .ZN(n11839) );
  XOR2_X1 U11892 ( .A(n12007), .B(n12008), .Z(n11836) );
  XOR2_X1 U11893 ( .A(n12009), .B(n12010), .Z(n12008) );
  OR2_X1 U11894 ( .A1(n8084), .A2(n8085), .ZN(n8086) );
  XOR2_X1 U11895 ( .A(n12011), .B(n12012), .Z(n11840) );
  XOR2_X1 U11896 ( .A(n12013), .B(n12014), .Z(n12012) );
  OR2_X1 U11897 ( .A1(n8085), .A2(n8079), .ZN(n11846) );
  XOR2_X1 U11898 ( .A(n12015), .B(n12016), .Z(n11843) );
  XOR2_X1 U11899 ( .A(n12017), .B(n12018), .Z(n12016) );
  OR2_X1 U11900 ( .A1(n8075), .A2(n8085), .ZN(n11850) );
  XNOR2_X1 U11901 ( .A(n12019), .B(n12020), .ZN(n11847) );
  XOR2_X1 U11902 ( .A(n7809), .B(n12021), .Z(n12019) );
  INV_X1 U11903 ( .A(n8081), .ZN(n7809) );
  OR2_X1 U11904 ( .A1(n8085), .A2(n8070), .ZN(n11854) );
  XOR2_X1 U11905 ( .A(n12022), .B(n12023), .Z(n11851) );
  XOR2_X1 U11906 ( .A(n12024), .B(n12025), .Z(n12023) );
  OR2_X1 U11907 ( .A1(n8066), .A2(n8085), .ZN(n11858) );
  XOR2_X1 U11908 ( .A(n12026), .B(n12027), .Z(n11855) );
  XOR2_X1 U11909 ( .A(n12028), .B(n12029), .Z(n12027) );
  OR2_X1 U11910 ( .A1(n8085), .A2(n8061), .ZN(n11862) );
  XOR2_X1 U11911 ( .A(n12030), .B(n12031), .Z(n11859) );
  XOR2_X1 U11912 ( .A(n12032), .B(n12033), .Z(n12031) );
  OR2_X1 U11913 ( .A1(n8057), .A2(n8085), .ZN(n11866) );
  XOR2_X1 U11914 ( .A(n12034), .B(n12035), .Z(n11863) );
  XOR2_X1 U11915 ( .A(n12036), .B(n12037), .Z(n12035) );
  OR2_X1 U11916 ( .A1(n8085), .A2(n8052), .ZN(n11870) );
  XOR2_X1 U11917 ( .A(n12038), .B(n12039), .Z(n11867) );
  XOR2_X1 U11918 ( .A(n12040), .B(n12041), .Z(n12039) );
  OR2_X1 U11919 ( .A1(n8048), .A2(n8085), .ZN(n11874) );
  XOR2_X1 U11920 ( .A(n12042), .B(n12043), .Z(n11871) );
  XOR2_X1 U11921 ( .A(n12044), .B(n12045), .Z(n12043) );
  OR2_X1 U11922 ( .A1(n8085), .A2(n8043), .ZN(n11878) );
  XOR2_X1 U11923 ( .A(n12046), .B(n12047), .Z(n11875) );
  XOR2_X1 U11924 ( .A(n12048), .B(n12049), .Z(n12047) );
  OR2_X1 U11925 ( .A1(n8039), .A2(n8085), .ZN(n11882) );
  XOR2_X1 U11926 ( .A(n12050), .B(n12051), .Z(n11879) );
  XOR2_X1 U11927 ( .A(n12052), .B(n12053), .Z(n12051) );
  OR2_X1 U11928 ( .A1(n8085), .A2(n8034), .ZN(n11886) );
  XOR2_X1 U11929 ( .A(n12054), .B(n12055), .Z(n11883) );
  XOR2_X1 U11930 ( .A(n12056), .B(n12057), .Z(n12055) );
  XOR2_X1 U11931 ( .A(n10912), .B(n12058), .Z(n10905) );
  XOR2_X1 U11932 ( .A(n10911), .B(n10910), .Z(n12058) );
  OR2_X1 U11933 ( .A1(n8080), .A2(n8034), .ZN(n10910) );
  OR2_X1 U11934 ( .A1(n12059), .A2(n12060), .ZN(n10911) );
  AND2_X1 U11935 ( .A1(n12057), .A2(n12056), .ZN(n12060) );
  AND2_X1 U11936 ( .A1(n12054), .A2(n12061), .ZN(n12059) );
  OR2_X1 U11937 ( .A1(n12057), .A2(n12056), .ZN(n12061) );
  OR2_X1 U11938 ( .A1(n12062), .A2(n12063), .ZN(n12056) );
  AND2_X1 U11939 ( .A1(n12053), .A2(n12052), .ZN(n12063) );
  AND2_X1 U11940 ( .A1(n12050), .A2(n12064), .ZN(n12062) );
  OR2_X1 U11941 ( .A1(n12053), .A2(n12052), .ZN(n12064) );
  OR2_X1 U11942 ( .A1(n12065), .A2(n12066), .ZN(n12052) );
  AND2_X1 U11943 ( .A1(n12049), .A2(n12048), .ZN(n12066) );
  AND2_X1 U11944 ( .A1(n12046), .A2(n12067), .ZN(n12065) );
  OR2_X1 U11945 ( .A1(n12049), .A2(n12048), .ZN(n12067) );
  OR2_X1 U11946 ( .A1(n12068), .A2(n12069), .ZN(n12048) );
  AND2_X1 U11947 ( .A1(n12045), .A2(n12044), .ZN(n12069) );
  AND2_X1 U11948 ( .A1(n12042), .A2(n12070), .ZN(n12068) );
  OR2_X1 U11949 ( .A1(n12045), .A2(n12044), .ZN(n12070) );
  OR2_X1 U11950 ( .A1(n12071), .A2(n12072), .ZN(n12044) );
  AND2_X1 U11951 ( .A1(n12041), .A2(n12040), .ZN(n12072) );
  AND2_X1 U11952 ( .A1(n12038), .A2(n12073), .ZN(n12071) );
  OR2_X1 U11953 ( .A1(n12041), .A2(n12040), .ZN(n12073) );
  OR2_X1 U11954 ( .A1(n12074), .A2(n12075), .ZN(n12040) );
  AND2_X1 U11955 ( .A1(n12037), .A2(n12036), .ZN(n12075) );
  AND2_X1 U11956 ( .A1(n12034), .A2(n12076), .ZN(n12074) );
  OR2_X1 U11957 ( .A1(n12037), .A2(n12036), .ZN(n12076) );
  OR2_X1 U11958 ( .A1(n12077), .A2(n12078), .ZN(n12036) );
  AND2_X1 U11959 ( .A1(n12030), .A2(n12033), .ZN(n12078) );
  AND2_X1 U11960 ( .A1(n12079), .A2(n12032), .ZN(n12077) );
  OR2_X1 U11961 ( .A1(n12080), .A2(n12081), .ZN(n12032) );
  AND2_X1 U11962 ( .A1(n12029), .A2(n12028), .ZN(n12081) );
  AND2_X1 U11963 ( .A1(n12026), .A2(n12082), .ZN(n12080) );
  OR2_X1 U11964 ( .A1(n12029), .A2(n12028), .ZN(n12082) );
  OR2_X1 U11965 ( .A1(n12083), .A2(n12084), .ZN(n12028) );
  AND2_X1 U11966 ( .A1(n12022), .A2(n12025), .ZN(n12084) );
  AND2_X1 U11967 ( .A1(n12085), .A2(n12024), .ZN(n12083) );
  OR2_X1 U11968 ( .A1(n12086), .A2(n12087), .ZN(n12024) );
  AND2_X1 U11969 ( .A1(n12020), .A2(n8081), .ZN(n12087) );
  AND2_X1 U11970 ( .A1(n12088), .A2(n12021), .ZN(n12086) );
  OR2_X1 U11971 ( .A1(n12089), .A2(n12090), .ZN(n12021) );
  AND2_X1 U11972 ( .A1(n12015), .A2(n12018), .ZN(n12090) );
  AND2_X1 U11973 ( .A1(n12091), .A2(n12017), .ZN(n12089) );
  OR2_X1 U11974 ( .A1(n12092), .A2(n12093), .ZN(n12017) );
  AND2_X1 U11975 ( .A1(n12011), .A2(n12014), .ZN(n12093) );
  AND2_X1 U11976 ( .A1(n12094), .A2(n12013), .ZN(n12092) );
  OR2_X1 U11977 ( .A1(n12095), .A2(n12096), .ZN(n12013) );
  AND2_X1 U11978 ( .A1(n12007), .A2(n12010), .ZN(n12096) );
  AND2_X1 U11979 ( .A1(n12097), .A2(n12009), .ZN(n12095) );
  OR2_X1 U11980 ( .A1(n12098), .A2(n12099), .ZN(n12009) );
  AND2_X1 U11981 ( .A1(n12003), .A2(n12006), .ZN(n12099) );
  AND2_X1 U11982 ( .A1(n12100), .A2(n12005), .ZN(n12098) );
  OR2_X1 U11983 ( .A1(n12101), .A2(n12102), .ZN(n12005) );
  AND2_X1 U11984 ( .A1(n11999), .A2(n12002), .ZN(n12102) );
  AND2_X1 U11985 ( .A1(n12103), .A2(n12001), .ZN(n12101) );
  OR2_X1 U11986 ( .A1(n12104), .A2(n12105), .ZN(n12001) );
  AND2_X1 U11987 ( .A1(n11995), .A2(n11998), .ZN(n12105) );
  AND2_X1 U11988 ( .A1(n12106), .A2(n11997), .ZN(n12104) );
  OR2_X1 U11989 ( .A1(n12107), .A2(n12108), .ZN(n11997) );
  AND2_X1 U11990 ( .A1(n11991), .A2(n11994), .ZN(n12108) );
  AND2_X1 U11991 ( .A1(n12109), .A2(n11993), .ZN(n12107) );
  OR2_X1 U11992 ( .A1(n12110), .A2(n12111), .ZN(n11993) );
  AND2_X1 U11993 ( .A1(n11987), .A2(n11990), .ZN(n12111) );
  AND2_X1 U11994 ( .A1(n12112), .A2(n11989), .ZN(n12110) );
  OR2_X1 U11995 ( .A1(n12113), .A2(n12114), .ZN(n11989) );
  AND2_X1 U11996 ( .A1(n11983), .A2(n11986), .ZN(n12114) );
  AND2_X1 U11997 ( .A1(n12115), .A2(n11985), .ZN(n12113) );
  OR2_X1 U11998 ( .A1(n12116), .A2(n12117), .ZN(n11985) );
  AND2_X1 U11999 ( .A1(n11979), .A2(n11982), .ZN(n12117) );
  AND2_X1 U12000 ( .A1(n12118), .A2(n11981), .ZN(n12116) );
  OR2_X1 U12001 ( .A1(n12119), .A2(n12120), .ZN(n11981) );
  AND2_X1 U12002 ( .A1(n11975), .A2(n11978), .ZN(n12120) );
  AND2_X1 U12003 ( .A1(n12121), .A2(n11977), .ZN(n12119) );
  OR2_X1 U12004 ( .A1(n12122), .A2(n12123), .ZN(n11977) );
  AND2_X1 U12005 ( .A1(n11971), .A2(n11974), .ZN(n12123) );
  AND2_X1 U12006 ( .A1(n12124), .A2(n11973), .ZN(n12122) );
  OR2_X1 U12007 ( .A1(n12125), .A2(n12126), .ZN(n11973) );
  AND2_X1 U12008 ( .A1(n11967), .A2(n11970), .ZN(n12126) );
  AND2_X1 U12009 ( .A1(n12127), .A2(n12128), .ZN(n12125) );
  OR2_X1 U12010 ( .A1(n11967), .A2(n11970), .ZN(n12128) );
  OR3_X1 U12011 ( .A1(n8076), .A2(n8080), .A3(n8981), .ZN(n11970) );
  OR2_X1 U12012 ( .A1(n8080), .A2(n8127), .ZN(n11967) );
  INV_X1 U12013 ( .A(n11969), .ZN(n12127) );
  OR2_X1 U12014 ( .A1(n12129), .A2(n12130), .ZN(n11969) );
  AND2_X1 U12015 ( .A1(b_15_), .A2(n12131), .ZN(n12130) );
  OR2_X1 U12016 ( .A1(n12132), .A2(n7598), .ZN(n12131) );
  AND2_X1 U12017 ( .A1(a_30_), .A2(n8071), .ZN(n12132) );
  AND2_X1 U12018 ( .A1(b_14_), .A2(n12133), .ZN(n12129) );
  OR2_X1 U12019 ( .A1(n12134), .A2(n7601), .ZN(n12133) );
  AND2_X1 U12020 ( .A1(a_31_), .A2(n8076), .ZN(n12134) );
  OR2_X1 U12021 ( .A1(n11971), .A2(n11974), .ZN(n12124) );
  OR2_X1 U12022 ( .A1(n8080), .A2(n8124), .ZN(n11974) );
  XNOR2_X1 U12023 ( .A(n12135), .B(n12136), .ZN(n11971) );
  XOR2_X1 U12024 ( .A(n12137), .B(n12138), .Z(n12136) );
  OR2_X1 U12025 ( .A1(n11975), .A2(n11978), .ZN(n12121) );
  OR2_X1 U12026 ( .A1(n8080), .A2(n8121), .ZN(n11978) );
  XOR2_X1 U12027 ( .A(n12139), .B(n12140), .Z(n11975) );
  XOR2_X1 U12028 ( .A(n12141), .B(n12142), .Z(n12140) );
  OR2_X1 U12029 ( .A1(n11979), .A2(n11982), .ZN(n12118) );
  OR2_X1 U12030 ( .A1(n8080), .A2(n8118), .ZN(n11982) );
  XOR2_X1 U12031 ( .A(n12143), .B(n12144), .Z(n11979) );
  XOR2_X1 U12032 ( .A(n12145), .B(n12146), .Z(n12144) );
  OR2_X1 U12033 ( .A1(n11983), .A2(n11986), .ZN(n12115) );
  OR2_X1 U12034 ( .A1(n8080), .A2(n8115), .ZN(n11986) );
  XOR2_X1 U12035 ( .A(n12147), .B(n12148), .Z(n11983) );
  XOR2_X1 U12036 ( .A(n12149), .B(n12150), .Z(n12148) );
  OR2_X1 U12037 ( .A1(n11987), .A2(n11990), .ZN(n12112) );
  OR2_X1 U12038 ( .A1(n8080), .A2(n8112), .ZN(n11990) );
  XOR2_X1 U12039 ( .A(n12151), .B(n12152), .Z(n11987) );
  XOR2_X1 U12040 ( .A(n12153), .B(n12154), .Z(n12152) );
  OR2_X1 U12041 ( .A1(n11991), .A2(n11994), .ZN(n12109) );
  OR2_X1 U12042 ( .A1(n8080), .A2(n8109), .ZN(n11994) );
  XOR2_X1 U12043 ( .A(n12155), .B(n12156), .Z(n11991) );
  XOR2_X1 U12044 ( .A(n12157), .B(n12158), .Z(n12156) );
  OR2_X1 U12045 ( .A1(n11995), .A2(n11998), .ZN(n12106) );
  OR2_X1 U12046 ( .A1(n8080), .A2(n8106), .ZN(n11998) );
  XOR2_X1 U12047 ( .A(n12159), .B(n12160), .Z(n11995) );
  XOR2_X1 U12048 ( .A(n12161), .B(n12162), .Z(n12160) );
  OR2_X1 U12049 ( .A1(n11999), .A2(n12002), .ZN(n12103) );
  OR2_X1 U12050 ( .A1(n8080), .A2(n8102), .ZN(n12002) );
  XOR2_X1 U12051 ( .A(n12163), .B(n12164), .Z(n11999) );
  XOR2_X1 U12052 ( .A(n12165), .B(n12166), .Z(n12164) );
  OR2_X1 U12053 ( .A1(n12003), .A2(n12006), .ZN(n12100) );
  OR2_X1 U12054 ( .A1(n8080), .A2(n8097), .ZN(n12006) );
  XOR2_X1 U12055 ( .A(n12167), .B(n12168), .Z(n12003) );
  XOR2_X1 U12056 ( .A(n12169), .B(n12170), .Z(n12168) );
  OR2_X1 U12057 ( .A1(n12007), .A2(n12010), .ZN(n12097) );
  OR2_X1 U12058 ( .A1(n8080), .A2(n8093), .ZN(n12010) );
  XOR2_X1 U12059 ( .A(n12171), .B(n12172), .Z(n12007) );
  XOR2_X1 U12060 ( .A(n12173), .B(n12174), .Z(n12172) );
  OR2_X1 U12061 ( .A1(n12011), .A2(n12014), .ZN(n12094) );
  OR2_X1 U12062 ( .A1(n8080), .A2(n8088), .ZN(n12014) );
  XOR2_X1 U12063 ( .A(n12175), .B(n12176), .Z(n12011) );
  XOR2_X1 U12064 ( .A(n12177), .B(n12178), .Z(n12176) );
  OR2_X1 U12065 ( .A1(n12015), .A2(n12018), .ZN(n12091) );
  OR2_X1 U12066 ( .A1(n8080), .A2(n8084), .ZN(n12018) );
  XOR2_X1 U12067 ( .A(n12179), .B(n12180), .Z(n12015) );
  XOR2_X1 U12068 ( .A(n12181), .B(n12182), .Z(n12180) );
  OR2_X1 U12069 ( .A1(n12020), .A2(n8081), .ZN(n12088) );
  OR2_X1 U12070 ( .A1(n8080), .A2(n8079), .ZN(n8081) );
  XOR2_X1 U12071 ( .A(n12183), .B(n12184), .Z(n12020) );
  XOR2_X1 U12072 ( .A(n12185), .B(n12186), .Z(n12184) );
  OR2_X1 U12073 ( .A1(n12022), .A2(n12025), .ZN(n12085) );
  OR2_X1 U12074 ( .A1(n8075), .A2(n8080), .ZN(n12025) );
  XOR2_X1 U12075 ( .A(n12187), .B(n12188), .Z(n12022) );
  XOR2_X1 U12076 ( .A(n12189), .B(n12190), .Z(n12188) );
  OR2_X1 U12077 ( .A1(n8080), .A2(n8070), .ZN(n12029) );
  XOR2_X1 U12078 ( .A(n12191), .B(n12192), .Z(n12026) );
  XOR2_X1 U12079 ( .A(n12193), .B(n8077), .Z(n12192) );
  OR2_X1 U12080 ( .A1(n12030), .A2(n12033), .ZN(n12079) );
  OR2_X1 U12081 ( .A1(n8066), .A2(n8080), .ZN(n12033) );
  XOR2_X1 U12082 ( .A(n12194), .B(n12195), .Z(n12030) );
  XOR2_X1 U12083 ( .A(n12196), .B(n12197), .Z(n12195) );
  OR2_X1 U12084 ( .A1(n8080), .A2(n8061), .ZN(n12037) );
  XOR2_X1 U12085 ( .A(n12198), .B(n12199), .Z(n12034) );
  XOR2_X1 U12086 ( .A(n12200), .B(n12201), .Z(n12199) );
  OR2_X1 U12087 ( .A1(n8057), .A2(n8080), .ZN(n12041) );
  XOR2_X1 U12088 ( .A(n12202), .B(n12203), .Z(n12038) );
  XOR2_X1 U12089 ( .A(n12204), .B(n12205), .Z(n12203) );
  OR2_X1 U12090 ( .A1(n8080), .A2(n8052), .ZN(n12045) );
  XOR2_X1 U12091 ( .A(n12206), .B(n12207), .Z(n12042) );
  XOR2_X1 U12092 ( .A(n12208), .B(n12209), .Z(n12207) );
  OR2_X1 U12093 ( .A1(n8048), .A2(n8080), .ZN(n12049) );
  XOR2_X1 U12094 ( .A(n12210), .B(n12211), .Z(n12046) );
  XOR2_X1 U12095 ( .A(n12212), .B(n12213), .Z(n12211) );
  OR2_X1 U12096 ( .A1(n8080), .A2(n8043), .ZN(n12053) );
  XOR2_X1 U12097 ( .A(n12214), .B(n12215), .Z(n12050) );
  XOR2_X1 U12098 ( .A(n12216), .B(n12217), .Z(n12215) );
  OR2_X1 U12099 ( .A1(n8039), .A2(n8080), .ZN(n12057) );
  INV_X1 U12100 ( .A(b_16_), .ZN(n8080) );
  XOR2_X1 U12101 ( .A(n12218), .B(n12219), .Z(n12054) );
  XOR2_X1 U12102 ( .A(n12220), .B(n12221), .Z(n12219) );
  XOR2_X1 U12103 ( .A(n10919), .B(n12222), .Z(n10912) );
  XOR2_X1 U12104 ( .A(n10918), .B(n10917), .Z(n12222) );
  OR2_X1 U12105 ( .A1(n8039), .A2(n8076), .ZN(n10917) );
  OR2_X1 U12106 ( .A1(n12223), .A2(n12224), .ZN(n10918) );
  AND2_X1 U12107 ( .A1(n12221), .A2(n12220), .ZN(n12224) );
  AND2_X1 U12108 ( .A1(n12218), .A2(n12225), .ZN(n12223) );
  OR2_X1 U12109 ( .A1(n12220), .A2(n12221), .ZN(n12225) );
  OR2_X1 U12110 ( .A1(n8076), .A2(n8043), .ZN(n12221) );
  OR2_X1 U12111 ( .A1(n12226), .A2(n12227), .ZN(n12220) );
  AND2_X1 U12112 ( .A1(n12217), .A2(n12216), .ZN(n12227) );
  AND2_X1 U12113 ( .A1(n12214), .A2(n12228), .ZN(n12226) );
  OR2_X1 U12114 ( .A1(n12216), .A2(n12217), .ZN(n12228) );
  OR2_X1 U12115 ( .A1(n8048), .A2(n8076), .ZN(n12217) );
  OR2_X1 U12116 ( .A1(n12229), .A2(n12230), .ZN(n12216) );
  AND2_X1 U12117 ( .A1(n12213), .A2(n12212), .ZN(n12230) );
  AND2_X1 U12118 ( .A1(n12210), .A2(n12231), .ZN(n12229) );
  OR2_X1 U12119 ( .A1(n12212), .A2(n12213), .ZN(n12231) );
  OR2_X1 U12120 ( .A1(n8076), .A2(n8052), .ZN(n12213) );
  OR2_X1 U12121 ( .A1(n12232), .A2(n12233), .ZN(n12212) );
  AND2_X1 U12122 ( .A1(n12209), .A2(n12208), .ZN(n12233) );
  AND2_X1 U12123 ( .A1(n12206), .A2(n12234), .ZN(n12232) );
  OR2_X1 U12124 ( .A1(n12208), .A2(n12209), .ZN(n12234) );
  OR2_X1 U12125 ( .A1(n8057), .A2(n8076), .ZN(n12209) );
  OR2_X1 U12126 ( .A1(n12235), .A2(n12236), .ZN(n12208) );
  AND2_X1 U12127 ( .A1(n12205), .A2(n12204), .ZN(n12236) );
  AND2_X1 U12128 ( .A1(n12202), .A2(n12237), .ZN(n12235) );
  OR2_X1 U12129 ( .A1(n12204), .A2(n12205), .ZN(n12237) );
  OR2_X1 U12130 ( .A1(n8076), .A2(n8061), .ZN(n12205) );
  OR2_X1 U12131 ( .A1(n12238), .A2(n12239), .ZN(n12204) );
  AND2_X1 U12132 ( .A1(n12201), .A2(n12200), .ZN(n12239) );
  AND2_X1 U12133 ( .A1(n12198), .A2(n12240), .ZN(n12238) );
  OR2_X1 U12134 ( .A1(n12200), .A2(n12201), .ZN(n12240) );
  OR2_X1 U12135 ( .A1(n8066), .A2(n8076), .ZN(n12201) );
  OR2_X1 U12136 ( .A1(n12241), .A2(n12242), .ZN(n12200) );
  AND2_X1 U12137 ( .A1(n12197), .A2(n12196), .ZN(n12242) );
  AND2_X1 U12138 ( .A1(n12194), .A2(n12243), .ZN(n12241) );
  OR2_X1 U12139 ( .A1(n12196), .A2(n12197), .ZN(n12243) );
  OR2_X1 U12140 ( .A1(n8076), .A2(n8070), .ZN(n12197) );
  OR2_X1 U12141 ( .A1(n12244), .A2(n12245), .ZN(n12196) );
  AND2_X1 U12142 ( .A1(n8077), .A2(n12193), .ZN(n12245) );
  AND2_X1 U12143 ( .A1(n12191), .A2(n12246), .ZN(n12244) );
  OR2_X1 U12144 ( .A1(n12193), .A2(n8077), .ZN(n12246) );
  OR2_X1 U12145 ( .A1(n8075), .A2(n8076), .ZN(n8077) );
  OR2_X1 U12146 ( .A1(n12247), .A2(n12248), .ZN(n12193) );
  AND2_X1 U12147 ( .A1(n12190), .A2(n12189), .ZN(n12248) );
  AND2_X1 U12148 ( .A1(n12187), .A2(n12249), .ZN(n12247) );
  OR2_X1 U12149 ( .A1(n12189), .A2(n12190), .ZN(n12249) );
  OR2_X1 U12150 ( .A1(n8076), .A2(n8079), .ZN(n12190) );
  OR2_X1 U12151 ( .A1(n12250), .A2(n12251), .ZN(n12189) );
  AND2_X1 U12152 ( .A1(n12186), .A2(n12185), .ZN(n12251) );
  AND2_X1 U12153 ( .A1(n12183), .A2(n12252), .ZN(n12250) );
  OR2_X1 U12154 ( .A1(n12185), .A2(n12186), .ZN(n12252) );
  OR2_X1 U12155 ( .A1(n8076), .A2(n8084), .ZN(n12186) );
  OR2_X1 U12156 ( .A1(n12253), .A2(n12254), .ZN(n12185) );
  AND2_X1 U12157 ( .A1(n12182), .A2(n12181), .ZN(n12254) );
  AND2_X1 U12158 ( .A1(n12179), .A2(n12255), .ZN(n12253) );
  OR2_X1 U12159 ( .A1(n12181), .A2(n12182), .ZN(n12255) );
  OR2_X1 U12160 ( .A1(n8076), .A2(n8088), .ZN(n12182) );
  OR2_X1 U12161 ( .A1(n12256), .A2(n12257), .ZN(n12181) );
  AND2_X1 U12162 ( .A1(n12178), .A2(n12177), .ZN(n12257) );
  AND2_X1 U12163 ( .A1(n12175), .A2(n12258), .ZN(n12256) );
  OR2_X1 U12164 ( .A1(n12177), .A2(n12178), .ZN(n12258) );
  OR2_X1 U12165 ( .A1(n8076), .A2(n8093), .ZN(n12178) );
  OR2_X1 U12166 ( .A1(n12259), .A2(n12260), .ZN(n12177) );
  AND2_X1 U12167 ( .A1(n12174), .A2(n12173), .ZN(n12260) );
  AND2_X1 U12168 ( .A1(n12171), .A2(n12261), .ZN(n12259) );
  OR2_X1 U12169 ( .A1(n12173), .A2(n12174), .ZN(n12261) );
  OR2_X1 U12170 ( .A1(n8076), .A2(n8097), .ZN(n12174) );
  OR2_X1 U12171 ( .A1(n12262), .A2(n12263), .ZN(n12173) );
  AND2_X1 U12172 ( .A1(n12170), .A2(n12169), .ZN(n12263) );
  AND2_X1 U12173 ( .A1(n12167), .A2(n12264), .ZN(n12262) );
  OR2_X1 U12174 ( .A1(n12169), .A2(n12170), .ZN(n12264) );
  OR2_X1 U12175 ( .A1(n8076), .A2(n8102), .ZN(n12170) );
  OR2_X1 U12176 ( .A1(n12265), .A2(n12266), .ZN(n12169) );
  AND2_X1 U12177 ( .A1(n12166), .A2(n12165), .ZN(n12266) );
  AND2_X1 U12178 ( .A1(n12163), .A2(n12267), .ZN(n12265) );
  OR2_X1 U12179 ( .A1(n12165), .A2(n12166), .ZN(n12267) );
  OR2_X1 U12180 ( .A1(n8076), .A2(n8106), .ZN(n12166) );
  OR2_X1 U12181 ( .A1(n12268), .A2(n12269), .ZN(n12165) );
  AND2_X1 U12182 ( .A1(n12162), .A2(n12161), .ZN(n12269) );
  AND2_X1 U12183 ( .A1(n12159), .A2(n12270), .ZN(n12268) );
  OR2_X1 U12184 ( .A1(n12161), .A2(n12162), .ZN(n12270) );
  OR2_X1 U12185 ( .A1(n8076), .A2(n8109), .ZN(n12162) );
  OR2_X1 U12186 ( .A1(n12271), .A2(n12272), .ZN(n12161) );
  AND2_X1 U12187 ( .A1(n12158), .A2(n12157), .ZN(n12272) );
  AND2_X1 U12188 ( .A1(n12155), .A2(n12273), .ZN(n12271) );
  OR2_X1 U12189 ( .A1(n12157), .A2(n12158), .ZN(n12273) );
  OR2_X1 U12190 ( .A1(n8076), .A2(n8112), .ZN(n12158) );
  OR2_X1 U12191 ( .A1(n12274), .A2(n12275), .ZN(n12157) );
  AND2_X1 U12192 ( .A1(n12154), .A2(n12153), .ZN(n12275) );
  AND2_X1 U12193 ( .A1(n12151), .A2(n12276), .ZN(n12274) );
  OR2_X1 U12194 ( .A1(n12153), .A2(n12154), .ZN(n12276) );
  OR2_X1 U12195 ( .A1(n8076), .A2(n8115), .ZN(n12154) );
  OR2_X1 U12196 ( .A1(n12277), .A2(n12278), .ZN(n12153) );
  AND2_X1 U12197 ( .A1(n12150), .A2(n12149), .ZN(n12278) );
  AND2_X1 U12198 ( .A1(n12147), .A2(n12279), .ZN(n12277) );
  OR2_X1 U12199 ( .A1(n12149), .A2(n12150), .ZN(n12279) );
  OR2_X1 U12200 ( .A1(n8076), .A2(n8118), .ZN(n12150) );
  OR2_X1 U12201 ( .A1(n12280), .A2(n12281), .ZN(n12149) );
  AND2_X1 U12202 ( .A1(n12146), .A2(n12145), .ZN(n12281) );
  AND2_X1 U12203 ( .A1(n12143), .A2(n12282), .ZN(n12280) );
  OR2_X1 U12204 ( .A1(n12145), .A2(n12146), .ZN(n12282) );
  OR2_X1 U12205 ( .A1(n8076), .A2(n8121), .ZN(n12146) );
  OR2_X1 U12206 ( .A1(n12283), .A2(n12284), .ZN(n12145) );
  AND2_X1 U12207 ( .A1(n12142), .A2(n12141), .ZN(n12284) );
  AND2_X1 U12208 ( .A1(n12139), .A2(n12285), .ZN(n12283) );
  OR2_X1 U12209 ( .A1(n12141), .A2(n12142), .ZN(n12285) );
  OR2_X1 U12210 ( .A1(n8076), .A2(n8124), .ZN(n12142) );
  OR2_X1 U12211 ( .A1(n12286), .A2(n12287), .ZN(n12141) );
  AND2_X1 U12212 ( .A1(n12135), .A2(n12138), .ZN(n12287) );
  AND2_X1 U12213 ( .A1(n12288), .A2(n12289), .ZN(n12286) );
  OR2_X1 U12214 ( .A1(n12138), .A2(n12135), .ZN(n12289) );
  OR2_X1 U12215 ( .A1(n8076), .A2(n8127), .ZN(n12135) );
  OR3_X1 U12216 ( .A1(n8076), .A2(n8981), .A3(n8071), .ZN(n12138) );
  INV_X1 U12217 ( .A(n12137), .ZN(n12288) );
  OR2_X1 U12218 ( .A1(n12290), .A2(n12291), .ZN(n12137) );
  AND2_X1 U12219 ( .A1(b_14_), .A2(n12292), .ZN(n12291) );
  OR2_X1 U12220 ( .A1(n12293), .A2(n7598), .ZN(n12292) );
  AND2_X1 U12221 ( .A1(a_30_), .A2(n8067), .ZN(n12293) );
  AND2_X1 U12222 ( .A1(b_13_), .A2(n12294), .ZN(n12290) );
  OR2_X1 U12223 ( .A1(n12295), .A2(n7601), .ZN(n12294) );
  AND2_X1 U12224 ( .A1(a_31_), .A2(n8071), .ZN(n12295) );
  XNOR2_X1 U12225 ( .A(n12296), .B(n12297), .ZN(n12139) );
  XOR2_X1 U12226 ( .A(n12298), .B(n12299), .Z(n12297) );
  XOR2_X1 U12227 ( .A(n12300), .B(n12301), .Z(n12143) );
  XOR2_X1 U12228 ( .A(n12302), .B(n12303), .Z(n12301) );
  XOR2_X1 U12229 ( .A(n12304), .B(n12305), .Z(n12147) );
  XOR2_X1 U12230 ( .A(n12306), .B(n12307), .Z(n12305) );
  XOR2_X1 U12231 ( .A(n12308), .B(n12309), .Z(n12151) );
  XOR2_X1 U12232 ( .A(n12310), .B(n12311), .Z(n12309) );
  XOR2_X1 U12233 ( .A(n12312), .B(n12313), .Z(n12155) );
  XOR2_X1 U12234 ( .A(n12314), .B(n12315), .Z(n12313) );
  XOR2_X1 U12235 ( .A(n12316), .B(n12317), .Z(n12159) );
  XOR2_X1 U12236 ( .A(n12318), .B(n12319), .Z(n12317) );
  XOR2_X1 U12237 ( .A(n12320), .B(n12321), .Z(n12163) );
  XOR2_X1 U12238 ( .A(n12322), .B(n12323), .Z(n12321) );
  XOR2_X1 U12239 ( .A(n12324), .B(n12325), .Z(n12167) );
  XOR2_X1 U12240 ( .A(n12326), .B(n12327), .Z(n12325) );
  XOR2_X1 U12241 ( .A(n12328), .B(n12329), .Z(n12171) );
  XOR2_X1 U12242 ( .A(n12330), .B(n12331), .Z(n12329) );
  XOR2_X1 U12243 ( .A(n12332), .B(n12333), .Z(n12175) );
  XOR2_X1 U12244 ( .A(n12334), .B(n12335), .Z(n12333) );
  XOR2_X1 U12245 ( .A(n12336), .B(n12337), .Z(n12179) );
  XOR2_X1 U12246 ( .A(n12338), .B(n12339), .Z(n12337) );
  XOR2_X1 U12247 ( .A(n12340), .B(n12341), .Z(n12183) );
  XOR2_X1 U12248 ( .A(n12342), .B(n12343), .Z(n12341) );
  XOR2_X1 U12249 ( .A(n12344), .B(n12345), .Z(n12187) );
  XOR2_X1 U12250 ( .A(n12346), .B(n12347), .Z(n12345) );
  XOR2_X1 U12251 ( .A(n12348), .B(n12349), .Z(n12191) );
  XOR2_X1 U12252 ( .A(n12350), .B(n12351), .Z(n12349) );
  XOR2_X1 U12253 ( .A(n12352), .B(n12353), .Z(n12194) );
  XOR2_X1 U12254 ( .A(n12354), .B(n12355), .Z(n12353) );
  XNOR2_X1 U12255 ( .A(n12356), .B(n12357), .ZN(n12198) );
  XOR2_X1 U12256 ( .A(n7833), .B(n12358), .Z(n12356) );
  INV_X1 U12257 ( .A(n8072), .ZN(n7833) );
  XOR2_X1 U12258 ( .A(n12359), .B(n12360), .Z(n12202) );
  XOR2_X1 U12259 ( .A(n12361), .B(n12362), .Z(n12360) );
  XOR2_X1 U12260 ( .A(n12363), .B(n12364), .Z(n12206) );
  XOR2_X1 U12261 ( .A(n12365), .B(n12366), .Z(n12364) );
  XOR2_X1 U12262 ( .A(n12367), .B(n12368), .Z(n12210) );
  XOR2_X1 U12263 ( .A(n12369), .B(n12370), .Z(n12368) );
  XOR2_X1 U12264 ( .A(n12371), .B(n12372), .Z(n12214) );
  XOR2_X1 U12265 ( .A(n12373), .B(n12374), .Z(n12372) );
  XOR2_X1 U12266 ( .A(n12375), .B(n12376), .Z(n12218) );
  XOR2_X1 U12267 ( .A(n12377), .B(n12378), .Z(n12376) );
  XOR2_X1 U12268 ( .A(n12379), .B(n12380), .Z(n10919) );
  XOR2_X1 U12269 ( .A(n12381), .B(n12382), .Z(n12380) );
  XOR2_X1 U12270 ( .A(n8251), .B(n8250), .Z(n8239) );
  INV_X1 U12271 ( .A(n12383), .ZN(n8250) );
  OR2_X1 U12272 ( .A1(n12384), .A2(n12385), .ZN(n12383) );
  AND2_X1 U12273 ( .A1(n8620), .A2(n8619), .ZN(n12385) );
  AND2_X1 U12274 ( .A1(n8617), .A2(n12386), .ZN(n12384) );
  OR2_X1 U12275 ( .A1(n8619), .A2(n8620), .ZN(n12386) );
  OR2_X1 U12276 ( .A1(n8071), .A2(n8297), .ZN(n8620) );
  OR2_X1 U12277 ( .A1(n12387), .A2(n12388), .ZN(n8619) );
  AND2_X1 U12278 ( .A1(n8644), .A2(n8643), .ZN(n12388) );
  AND2_X1 U12279 ( .A1(n8641), .A2(n12389), .ZN(n12387) );
  OR2_X1 U12280 ( .A1(n8643), .A2(n8644), .ZN(n12389) );
  OR2_X1 U12281 ( .A1(n8071), .A2(n8012), .ZN(n8644) );
  OR2_X1 U12282 ( .A1(n12390), .A2(n12391), .ZN(n8643) );
  AND2_X1 U12283 ( .A1(n8675), .A2(n8674), .ZN(n12391) );
  AND2_X1 U12284 ( .A1(n8672), .A2(n12392), .ZN(n12390) );
  OR2_X1 U12285 ( .A1(n8674), .A2(n8675), .ZN(n12392) );
  OR2_X1 U12286 ( .A1(n8071), .A2(n8016), .ZN(n8675) );
  OR2_X1 U12287 ( .A1(n12393), .A2(n12394), .ZN(n8674) );
  AND2_X1 U12288 ( .A1(n8713), .A2(n8712), .ZN(n12394) );
  AND2_X1 U12289 ( .A1(n8710), .A2(n12395), .ZN(n12393) );
  OR2_X1 U12290 ( .A1(n8712), .A2(n8713), .ZN(n12395) );
  OR2_X1 U12291 ( .A1(n8021), .A2(n8071), .ZN(n8713) );
  OR2_X1 U12292 ( .A1(n12396), .A2(n12397), .ZN(n8712) );
  AND2_X1 U12293 ( .A1(n8758), .A2(n8757), .ZN(n12397) );
  AND2_X1 U12294 ( .A1(n8755), .A2(n12398), .ZN(n12396) );
  OR2_X1 U12295 ( .A1(n8757), .A2(n8758), .ZN(n12398) );
  OR2_X1 U12296 ( .A1(n8071), .A2(n8025), .ZN(n8758) );
  OR2_X1 U12297 ( .A1(n12399), .A2(n12400), .ZN(n8757) );
  AND2_X1 U12298 ( .A1(n8810), .A2(n8809), .ZN(n12400) );
  AND2_X1 U12299 ( .A1(n8807), .A2(n12401), .ZN(n12399) );
  OR2_X1 U12300 ( .A1(n8809), .A2(n8810), .ZN(n12401) );
  OR2_X1 U12301 ( .A1(n8030), .A2(n8071), .ZN(n8810) );
  OR2_X1 U12302 ( .A1(n12402), .A2(n12403), .ZN(n8809) );
  AND2_X1 U12303 ( .A1(n10871), .A2(n10870), .ZN(n12403) );
  AND2_X1 U12304 ( .A1(n10868), .A2(n12404), .ZN(n12402) );
  OR2_X1 U12305 ( .A1(n10870), .A2(n10871), .ZN(n12404) );
  OR2_X1 U12306 ( .A1(n8071), .A2(n8034), .ZN(n10871) );
  OR2_X1 U12307 ( .A1(n12405), .A2(n12406), .ZN(n10870) );
  AND2_X1 U12308 ( .A1(n10924), .A2(n10923), .ZN(n12406) );
  AND2_X1 U12309 ( .A1(n10921), .A2(n12407), .ZN(n12405) );
  OR2_X1 U12310 ( .A1(n10923), .A2(n10924), .ZN(n12407) );
  OR2_X1 U12311 ( .A1(n8039), .A2(n8071), .ZN(n10924) );
  OR2_X1 U12312 ( .A1(n12408), .A2(n12409), .ZN(n10923) );
  AND2_X1 U12313 ( .A1(n12382), .A2(n12381), .ZN(n12409) );
  AND2_X1 U12314 ( .A1(n12379), .A2(n12410), .ZN(n12408) );
  OR2_X1 U12315 ( .A1(n12381), .A2(n12382), .ZN(n12410) );
  OR2_X1 U12316 ( .A1(n8071), .A2(n8043), .ZN(n12382) );
  OR2_X1 U12317 ( .A1(n12411), .A2(n12412), .ZN(n12381) );
  AND2_X1 U12318 ( .A1(n12378), .A2(n12377), .ZN(n12412) );
  AND2_X1 U12319 ( .A1(n12375), .A2(n12413), .ZN(n12411) );
  OR2_X1 U12320 ( .A1(n12377), .A2(n12378), .ZN(n12413) );
  OR2_X1 U12321 ( .A1(n8048), .A2(n8071), .ZN(n12378) );
  OR2_X1 U12322 ( .A1(n12414), .A2(n12415), .ZN(n12377) );
  AND2_X1 U12323 ( .A1(n12374), .A2(n12373), .ZN(n12415) );
  AND2_X1 U12324 ( .A1(n12371), .A2(n12416), .ZN(n12414) );
  OR2_X1 U12325 ( .A1(n12373), .A2(n12374), .ZN(n12416) );
  OR2_X1 U12326 ( .A1(n8071), .A2(n8052), .ZN(n12374) );
  OR2_X1 U12327 ( .A1(n12417), .A2(n12418), .ZN(n12373) );
  AND2_X1 U12328 ( .A1(n12370), .A2(n12369), .ZN(n12418) );
  AND2_X1 U12329 ( .A1(n12367), .A2(n12419), .ZN(n12417) );
  OR2_X1 U12330 ( .A1(n12369), .A2(n12370), .ZN(n12419) );
  OR2_X1 U12331 ( .A1(n8057), .A2(n8071), .ZN(n12370) );
  OR2_X1 U12332 ( .A1(n12420), .A2(n12421), .ZN(n12369) );
  AND2_X1 U12333 ( .A1(n12366), .A2(n12365), .ZN(n12421) );
  AND2_X1 U12334 ( .A1(n12363), .A2(n12422), .ZN(n12420) );
  OR2_X1 U12335 ( .A1(n12365), .A2(n12366), .ZN(n12422) );
  OR2_X1 U12336 ( .A1(n8071), .A2(n8061), .ZN(n12366) );
  OR2_X1 U12337 ( .A1(n12423), .A2(n12424), .ZN(n12365) );
  AND2_X1 U12338 ( .A1(n12362), .A2(n12361), .ZN(n12424) );
  AND2_X1 U12339 ( .A1(n12359), .A2(n12425), .ZN(n12423) );
  OR2_X1 U12340 ( .A1(n12361), .A2(n12362), .ZN(n12425) );
  OR2_X1 U12341 ( .A1(n8066), .A2(n8071), .ZN(n12362) );
  OR2_X1 U12342 ( .A1(n12426), .A2(n12427), .ZN(n12361) );
  AND2_X1 U12343 ( .A1(n12358), .A2(n8072), .ZN(n12427) );
  AND2_X1 U12344 ( .A1(n12357), .A2(n12428), .ZN(n12426) );
  OR2_X1 U12345 ( .A1(n8072), .A2(n12358), .ZN(n12428) );
  OR2_X1 U12346 ( .A1(n12429), .A2(n12430), .ZN(n12358) );
  AND2_X1 U12347 ( .A1(n12355), .A2(n12354), .ZN(n12430) );
  AND2_X1 U12348 ( .A1(n12352), .A2(n12431), .ZN(n12429) );
  OR2_X1 U12349 ( .A1(n12354), .A2(n12355), .ZN(n12431) );
  OR2_X1 U12350 ( .A1(n8075), .A2(n8071), .ZN(n12355) );
  OR2_X1 U12351 ( .A1(n12432), .A2(n12433), .ZN(n12354) );
  AND2_X1 U12352 ( .A1(n12351), .A2(n12350), .ZN(n12433) );
  AND2_X1 U12353 ( .A1(n12348), .A2(n12434), .ZN(n12432) );
  OR2_X1 U12354 ( .A1(n12350), .A2(n12351), .ZN(n12434) );
  OR2_X1 U12355 ( .A1(n8079), .A2(n8071), .ZN(n12351) );
  OR2_X1 U12356 ( .A1(n12435), .A2(n12436), .ZN(n12350) );
  AND2_X1 U12357 ( .A1(n12347), .A2(n12346), .ZN(n12436) );
  AND2_X1 U12358 ( .A1(n12344), .A2(n12437), .ZN(n12435) );
  OR2_X1 U12359 ( .A1(n12346), .A2(n12347), .ZN(n12437) );
  OR2_X1 U12360 ( .A1(n8084), .A2(n8071), .ZN(n12347) );
  OR2_X1 U12361 ( .A1(n12438), .A2(n12439), .ZN(n12346) );
  AND2_X1 U12362 ( .A1(n12343), .A2(n12342), .ZN(n12439) );
  AND2_X1 U12363 ( .A1(n12340), .A2(n12440), .ZN(n12438) );
  OR2_X1 U12364 ( .A1(n12342), .A2(n12343), .ZN(n12440) );
  OR2_X1 U12365 ( .A1(n8088), .A2(n8071), .ZN(n12343) );
  OR2_X1 U12366 ( .A1(n12441), .A2(n12442), .ZN(n12342) );
  AND2_X1 U12367 ( .A1(n12339), .A2(n12338), .ZN(n12442) );
  AND2_X1 U12368 ( .A1(n12336), .A2(n12443), .ZN(n12441) );
  OR2_X1 U12369 ( .A1(n12338), .A2(n12339), .ZN(n12443) );
  OR2_X1 U12370 ( .A1(n8093), .A2(n8071), .ZN(n12339) );
  OR2_X1 U12371 ( .A1(n12444), .A2(n12445), .ZN(n12338) );
  AND2_X1 U12372 ( .A1(n12335), .A2(n12334), .ZN(n12445) );
  AND2_X1 U12373 ( .A1(n12332), .A2(n12446), .ZN(n12444) );
  OR2_X1 U12374 ( .A1(n12334), .A2(n12335), .ZN(n12446) );
  OR2_X1 U12375 ( .A1(n8097), .A2(n8071), .ZN(n12335) );
  OR2_X1 U12376 ( .A1(n12447), .A2(n12448), .ZN(n12334) );
  AND2_X1 U12377 ( .A1(n12331), .A2(n12330), .ZN(n12448) );
  AND2_X1 U12378 ( .A1(n12328), .A2(n12449), .ZN(n12447) );
  OR2_X1 U12379 ( .A1(n12330), .A2(n12331), .ZN(n12449) );
  OR2_X1 U12380 ( .A1(n8102), .A2(n8071), .ZN(n12331) );
  OR2_X1 U12381 ( .A1(n12450), .A2(n12451), .ZN(n12330) );
  AND2_X1 U12382 ( .A1(n12327), .A2(n12326), .ZN(n12451) );
  AND2_X1 U12383 ( .A1(n12324), .A2(n12452), .ZN(n12450) );
  OR2_X1 U12384 ( .A1(n12326), .A2(n12327), .ZN(n12452) );
  OR2_X1 U12385 ( .A1(n8106), .A2(n8071), .ZN(n12327) );
  OR2_X1 U12386 ( .A1(n12453), .A2(n12454), .ZN(n12326) );
  AND2_X1 U12387 ( .A1(n12323), .A2(n12322), .ZN(n12454) );
  AND2_X1 U12388 ( .A1(n12320), .A2(n12455), .ZN(n12453) );
  OR2_X1 U12389 ( .A1(n12322), .A2(n12323), .ZN(n12455) );
  OR2_X1 U12390 ( .A1(n8109), .A2(n8071), .ZN(n12323) );
  OR2_X1 U12391 ( .A1(n12456), .A2(n12457), .ZN(n12322) );
  AND2_X1 U12392 ( .A1(n12319), .A2(n12318), .ZN(n12457) );
  AND2_X1 U12393 ( .A1(n12316), .A2(n12458), .ZN(n12456) );
  OR2_X1 U12394 ( .A1(n12318), .A2(n12319), .ZN(n12458) );
  OR2_X1 U12395 ( .A1(n8112), .A2(n8071), .ZN(n12319) );
  OR2_X1 U12396 ( .A1(n12459), .A2(n12460), .ZN(n12318) );
  AND2_X1 U12397 ( .A1(n12315), .A2(n12314), .ZN(n12460) );
  AND2_X1 U12398 ( .A1(n12312), .A2(n12461), .ZN(n12459) );
  OR2_X1 U12399 ( .A1(n12314), .A2(n12315), .ZN(n12461) );
  OR2_X1 U12400 ( .A1(n8115), .A2(n8071), .ZN(n12315) );
  OR2_X1 U12401 ( .A1(n12462), .A2(n12463), .ZN(n12314) );
  AND2_X1 U12402 ( .A1(n12311), .A2(n12310), .ZN(n12463) );
  AND2_X1 U12403 ( .A1(n12308), .A2(n12464), .ZN(n12462) );
  OR2_X1 U12404 ( .A1(n12310), .A2(n12311), .ZN(n12464) );
  OR2_X1 U12405 ( .A1(n8118), .A2(n8071), .ZN(n12311) );
  OR2_X1 U12406 ( .A1(n12465), .A2(n12466), .ZN(n12310) );
  AND2_X1 U12407 ( .A1(n12307), .A2(n12306), .ZN(n12466) );
  AND2_X1 U12408 ( .A1(n12304), .A2(n12467), .ZN(n12465) );
  OR2_X1 U12409 ( .A1(n12306), .A2(n12307), .ZN(n12467) );
  OR2_X1 U12410 ( .A1(n8121), .A2(n8071), .ZN(n12307) );
  OR2_X1 U12411 ( .A1(n12468), .A2(n12469), .ZN(n12306) );
  AND2_X1 U12412 ( .A1(n12303), .A2(n12302), .ZN(n12469) );
  AND2_X1 U12413 ( .A1(n12300), .A2(n12470), .ZN(n12468) );
  OR2_X1 U12414 ( .A1(n12302), .A2(n12303), .ZN(n12470) );
  OR2_X1 U12415 ( .A1(n8124), .A2(n8071), .ZN(n12303) );
  OR2_X1 U12416 ( .A1(n12471), .A2(n12472), .ZN(n12302) );
  AND2_X1 U12417 ( .A1(n12296), .A2(n12299), .ZN(n12472) );
  AND2_X1 U12418 ( .A1(n12473), .A2(n12474), .ZN(n12471) );
  OR2_X1 U12419 ( .A1(n12299), .A2(n12296), .ZN(n12474) );
  OR2_X1 U12420 ( .A1(n8127), .A2(n8071), .ZN(n12296) );
  OR3_X1 U12421 ( .A1(n8067), .A2(n8981), .A3(n8071), .ZN(n12299) );
  INV_X1 U12422 ( .A(n12298), .ZN(n12473) );
  OR2_X1 U12423 ( .A1(n12475), .A2(n12476), .ZN(n12298) );
  AND2_X1 U12424 ( .A1(b_13_), .A2(n12477), .ZN(n12476) );
  OR2_X1 U12425 ( .A1(n12478), .A2(n7598), .ZN(n12477) );
  AND2_X1 U12426 ( .A1(a_30_), .A2(n8062), .ZN(n12478) );
  AND2_X1 U12427 ( .A1(b_12_), .A2(n12479), .ZN(n12475) );
  OR2_X1 U12428 ( .A1(n12480), .A2(n7601), .ZN(n12479) );
  AND2_X1 U12429 ( .A1(a_31_), .A2(n8067), .ZN(n12480) );
  XNOR2_X1 U12430 ( .A(n12481), .B(n12482), .ZN(n12300) );
  XOR2_X1 U12431 ( .A(n12483), .B(n12484), .Z(n12482) );
  XOR2_X1 U12432 ( .A(n12485), .B(n12486), .Z(n12304) );
  XOR2_X1 U12433 ( .A(n12487), .B(n12488), .Z(n12486) );
  XOR2_X1 U12434 ( .A(n12489), .B(n12490), .Z(n12308) );
  XOR2_X1 U12435 ( .A(n12491), .B(n12492), .Z(n12490) );
  XOR2_X1 U12436 ( .A(n12493), .B(n12494), .Z(n12312) );
  XOR2_X1 U12437 ( .A(n12495), .B(n12496), .Z(n12494) );
  XOR2_X1 U12438 ( .A(n12497), .B(n12498), .Z(n12316) );
  XOR2_X1 U12439 ( .A(n12499), .B(n12500), .Z(n12498) );
  XOR2_X1 U12440 ( .A(n12501), .B(n12502), .Z(n12320) );
  XOR2_X1 U12441 ( .A(n12503), .B(n12504), .Z(n12502) );
  XOR2_X1 U12442 ( .A(n12505), .B(n12506), .Z(n12324) );
  XOR2_X1 U12443 ( .A(n12507), .B(n12508), .Z(n12506) );
  XOR2_X1 U12444 ( .A(n12509), .B(n12510), .Z(n12328) );
  XOR2_X1 U12445 ( .A(n12511), .B(n12512), .Z(n12510) );
  XOR2_X1 U12446 ( .A(n12513), .B(n12514), .Z(n12332) );
  XOR2_X1 U12447 ( .A(n12515), .B(n12516), .Z(n12514) );
  XOR2_X1 U12448 ( .A(n12517), .B(n12518), .Z(n12336) );
  XOR2_X1 U12449 ( .A(n12519), .B(n12520), .Z(n12518) );
  XOR2_X1 U12450 ( .A(n12521), .B(n12522), .Z(n12340) );
  XOR2_X1 U12451 ( .A(n12523), .B(n12524), .Z(n12522) );
  XOR2_X1 U12452 ( .A(n12525), .B(n12526), .Z(n12344) );
  XOR2_X1 U12453 ( .A(n12527), .B(n12528), .Z(n12526) );
  XOR2_X1 U12454 ( .A(n12529), .B(n12530), .Z(n12348) );
  XOR2_X1 U12455 ( .A(n12531), .B(n12532), .Z(n12530) );
  XOR2_X1 U12456 ( .A(n12533), .B(n12534), .Z(n12352) );
  XOR2_X1 U12457 ( .A(n12535), .B(n12536), .Z(n12534) );
  OR2_X1 U12458 ( .A1(n8070), .A2(n8071), .ZN(n8072) );
  INV_X1 U12459 ( .A(b_14_), .ZN(n8071) );
  XOR2_X1 U12460 ( .A(n12537), .B(n12538), .Z(n12357) );
  XOR2_X1 U12461 ( .A(n12539), .B(n12540), .Z(n12538) );
  XOR2_X1 U12462 ( .A(n12541), .B(n12542), .Z(n12359) );
  XOR2_X1 U12463 ( .A(n12543), .B(n12544), .Z(n12542) );
  XOR2_X1 U12464 ( .A(n12545), .B(n12546), .Z(n12363) );
  XOR2_X1 U12465 ( .A(n12547), .B(n8068), .Z(n12546) );
  XOR2_X1 U12466 ( .A(n12548), .B(n12549), .Z(n12367) );
  XOR2_X1 U12467 ( .A(n12550), .B(n12551), .Z(n12549) );
  XOR2_X1 U12468 ( .A(n12552), .B(n12553), .Z(n12371) );
  XOR2_X1 U12469 ( .A(n12554), .B(n12555), .Z(n12553) );
  XOR2_X1 U12470 ( .A(n12556), .B(n12557), .Z(n12375) );
  XOR2_X1 U12471 ( .A(n12558), .B(n12559), .Z(n12557) );
  XOR2_X1 U12472 ( .A(n12560), .B(n12561), .Z(n12379) );
  XOR2_X1 U12473 ( .A(n12562), .B(n12563), .Z(n12561) );
  XOR2_X1 U12474 ( .A(n12564), .B(n12565), .Z(n10921) );
  XOR2_X1 U12475 ( .A(n12566), .B(n12567), .Z(n12565) );
  XOR2_X1 U12476 ( .A(n12568), .B(n12569), .Z(n10868) );
  XOR2_X1 U12477 ( .A(n12570), .B(n12571), .Z(n12569) );
  XOR2_X1 U12478 ( .A(n12572), .B(n12573), .Z(n8807) );
  XOR2_X1 U12479 ( .A(n12574), .B(n12575), .Z(n12573) );
  XOR2_X1 U12480 ( .A(n12576), .B(n12577), .Z(n8755) );
  XOR2_X1 U12481 ( .A(n12578), .B(n12579), .Z(n12577) );
  XOR2_X1 U12482 ( .A(n12580), .B(n12581), .Z(n8710) );
  XOR2_X1 U12483 ( .A(n12582), .B(n12583), .Z(n12581) );
  XOR2_X1 U12484 ( .A(n12584), .B(n12585), .Z(n8672) );
  XOR2_X1 U12485 ( .A(n12586), .B(n12587), .Z(n12585) );
  XOR2_X1 U12486 ( .A(n12588), .B(n12589), .Z(n8641) );
  XOR2_X1 U12487 ( .A(n12590), .B(n12591), .Z(n12589) );
  XOR2_X1 U12488 ( .A(n12592), .B(n12593), .Z(n8617) );
  XOR2_X1 U12489 ( .A(n12594), .B(n12595), .Z(n12593) );
  XNOR2_X1 U12490 ( .A(n12596), .B(n12597), .ZN(n8251) );
  XOR2_X1 U12491 ( .A(n12598), .B(n12599), .Z(n12597) );
  AND2_X1 U12492 ( .A1(n12600), .A2(n12601), .ZN(n8249) );
  INV_X1 U12493 ( .A(n12602), .ZN(n12600) );
  AND2_X1 U12494 ( .A1(n12603), .A2(n12604), .ZN(n12602) );
  INV_X1 U12495 ( .A(n12601), .ZN(n8599) );
  OR2_X1 U12496 ( .A1(n12603), .A2(n12604), .ZN(n12601) );
  OR2_X1 U12497 ( .A1(n12605), .A2(n12606), .ZN(n12604) );
  AND2_X1 U12498 ( .A1(n12599), .A2(n12598), .ZN(n12606) );
  AND2_X1 U12499 ( .A1(n12596), .A2(n12607), .ZN(n12605) );
  OR2_X1 U12500 ( .A1(n12599), .A2(n12598), .ZN(n12607) );
  OR2_X1 U12501 ( .A1(n12608), .A2(n12609), .ZN(n12598) );
  AND2_X1 U12502 ( .A1(n12595), .A2(n12594), .ZN(n12609) );
  AND2_X1 U12503 ( .A1(n12592), .A2(n12610), .ZN(n12608) );
  OR2_X1 U12504 ( .A1(n12595), .A2(n12594), .ZN(n12610) );
  OR2_X1 U12505 ( .A1(n12611), .A2(n12612), .ZN(n12594) );
  AND2_X1 U12506 ( .A1(n12591), .A2(n12590), .ZN(n12612) );
  AND2_X1 U12507 ( .A1(n12588), .A2(n12613), .ZN(n12611) );
  OR2_X1 U12508 ( .A1(n12591), .A2(n12590), .ZN(n12613) );
  OR2_X1 U12509 ( .A1(n12614), .A2(n12615), .ZN(n12590) );
  AND2_X1 U12510 ( .A1(n12587), .A2(n12586), .ZN(n12615) );
  AND2_X1 U12511 ( .A1(n12584), .A2(n12616), .ZN(n12614) );
  OR2_X1 U12512 ( .A1(n12587), .A2(n12586), .ZN(n12616) );
  OR2_X1 U12513 ( .A1(n12617), .A2(n12618), .ZN(n12586) );
  AND2_X1 U12514 ( .A1(n12583), .A2(n12582), .ZN(n12618) );
  AND2_X1 U12515 ( .A1(n12580), .A2(n12619), .ZN(n12617) );
  OR2_X1 U12516 ( .A1(n12583), .A2(n12582), .ZN(n12619) );
  OR2_X1 U12517 ( .A1(n12620), .A2(n12621), .ZN(n12582) );
  AND2_X1 U12518 ( .A1(n12579), .A2(n12578), .ZN(n12621) );
  AND2_X1 U12519 ( .A1(n12576), .A2(n12622), .ZN(n12620) );
  OR2_X1 U12520 ( .A1(n12579), .A2(n12578), .ZN(n12622) );
  OR2_X1 U12521 ( .A1(n12623), .A2(n12624), .ZN(n12578) );
  AND2_X1 U12522 ( .A1(n12575), .A2(n12574), .ZN(n12624) );
  AND2_X1 U12523 ( .A1(n12572), .A2(n12625), .ZN(n12623) );
  OR2_X1 U12524 ( .A1(n12575), .A2(n12574), .ZN(n12625) );
  OR2_X1 U12525 ( .A1(n12626), .A2(n12627), .ZN(n12574) );
  AND2_X1 U12526 ( .A1(n12571), .A2(n12570), .ZN(n12627) );
  AND2_X1 U12527 ( .A1(n12568), .A2(n12628), .ZN(n12626) );
  OR2_X1 U12528 ( .A1(n12571), .A2(n12570), .ZN(n12628) );
  OR2_X1 U12529 ( .A1(n12629), .A2(n12630), .ZN(n12570) );
  AND2_X1 U12530 ( .A1(n12567), .A2(n12566), .ZN(n12630) );
  AND2_X1 U12531 ( .A1(n12564), .A2(n12631), .ZN(n12629) );
  OR2_X1 U12532 ( .A1(n12567), .A2(n12566), .ZN(n12631) );
  OR2_X1 U12533 ( .A1(n12632), .A2(n12633), .ZN(n12566) );
  AND2_X1 U12534 ( .A1(n12563), .A2(n12562), .ZN(n12633) );
  AND2_X1 U12535 ( .A1(n12560), .A2(n12634), .ZN(n12632) );
  OR2_X1 U12536 ( .A1(n12563), .A2(n12562), .ZN(n12634) );
  OR2_X1 U12537 ( .A1(n12635), .A2(n12636), .ZN(n12562) );
  AND2_X1 U12538 ( .A1(n12559), .A2(n12558), .ZN(n12636) );
  AND2_X1 U12539 ( .A1(n12556), .A2(n12637), .ZN(n12635) );
  OR2_X1 U12540 ( .A1(n12559), .A2(n12558), .ZN(n12637) );
  OR2_X1 U12541 ( .A1(n12638), .A2(n12639), .ZN(n12558) );
  AND2_X1 U12542 ( .A1(n12555), .A2(n12554), .ZN(n12639) );
  AND2_X1 U12543 ( .A1(n12552), .A2(n12640), .ZN(n12638) );
  OR2_X1 U12544 ( .A1(n12555), .A2(n12554), .ZN(n12640) );
  OR2_X1 U12545 ( .A1(n12641), .A2(n12642), .ZN(n12554) );
  AND2_X1 U12546 ( .A1(n12551), .A2(n12550), .ZN(n12642) );
  AND2_X1 U12547 ( .A1(n12548), .A2(n12643), .ZN(n12641) );
  OR2_X1 U12548 ( .A1(n12551), .A2(n12550), .ZN(n12643) );
  OR2_X1 U12549 ( .A1(n12644), .A2(n12645), .ZN(n12550) );
  AND2_X1 U12550 ( .A1(n8068), .A2(n12547), .ZN(n12645) );
  AND2_X1 U12551 ( .A1(n12545), .A2(n12646), .ZN(n12644) );
  OR2_X1 U12552 ( .A1(n8068), .A2(n12547), .ZN(n12646) );
  OR2_X1 U12553 ( .A1(n12647), .A2(n12648), .ZN(n12547) );
  AND2_X1 U12554 ( .A1(n12544), .A2(n12543), .ZN(n12648) );
  AND2_X1 U12555 ( .A1(n12541), .A2(n12649), .ZN(n12647) );
  OR2_X1 U12556 ( .A1(n12544), .A2(n12543), .ZN(n12649) );
  OR2_X1 U12557 ( .A1(n12650), .A2(n12651), .ZN(n12543) );
  AND2_X1 U12558 ( .A1(n12540), .A2(n12539), .ZN(n12651) );
  AND2_X1 U12559 ( .A1(n12537), .A2(n12652), .ZN(n12650) );
  OR2_X1 U12560 ( .A1(n12540), .A2(n12539), .ZN(n12652) );
  OR2_X1 U12561 ( .A1(n12653), .A2(n12654), .ZN(n12539) );
  AND2_X1 U12562 ( .A1(n12536), .A2(n12535), .ZN(n12654) );
  AND2_X1 U12563 ( .A1(n12533), .A2(n12655), .ZN(n12653) );
  OR2_X1 U12564 ( .A1(n12536), .A2(n12535), .ZN(n12655) );
  OR2_X1 U12565 ( .A1(n12656), .A2(n12657), .ZN(n12535) );
  AND2_X1 U12566 ( .A1(n12532), .A2(n12531), .ZN(n12657) );
  AND2_X1 U12567 ( .A1(n12529), .A2(n12658), .ZN(n12656) );
  OR2_X1 U12568 ( .A1(n12532), .A2(n12531), .ZN(n12658) );
  OR2_X1 U12569 ( .A1(n12659), .A2(n12660), .ZN(n12531) );
  AND2_X1 U12570 ( .A1(n12528), .A2(n12527), .ZN(n12660) );
  AND2_X1 U12571 ( .A1(n12525), .A2(n12661), .ZN(n12659) );
  OR2_X1 U12572 ( .A1(n12528), .A2(n12527), .ZN(n12661) );
  OR2_X1 U12573 ( .A1(n12662), .A2(n12663), .ZN(n12527) );
  AND2_X1 U12574 ( .A1(n12524), .A2(n12523), .ZN(n12663) );
  AND2_X1 U12575 ( .A1(n12521), .A2(n12664), .ZN(n12662) );
  OR2_X1 U12576 ( .A1(n12524), .A2(n12523), .ZN(n12664) );
  OR2_X1 U12577 ( .A1(n12665), .A2(n12666), .ZN(n12523) );
  AND2_X1 U12578 ( .A1(n12520), .A2(n12519), .ZN(n12666) );
  AND2_X1 U12579 ( .A1(n12517), .A2(n12667), .ZN(n12665) );
  OR2_X1 U12580 ( .A1(n12520), .A2(n12519), .ZN(n12667) );
  OR2_X1 U12581 ( .A1(n12668), .A2(n12669), .ZN(n12519) );
  AND2_X1 U12582 ( .A1(n12516), .A2(n12515), .ZN(n12669) );
  AND2_X1 U12583 ( .A1(n12513), .A2(n12670), .ZN(n12668) );
  OR2_X1 U12584 ( .A1(n12516), .A2(n12515), .ZN(n12670) );
  OR2_X1 U12585 ( .A1(n12671), .A2(n12672), .ZN(n12515) );
  AND2_X1 U12586 ( .A1(n12512), .A2(n12511), .ZN(n12672) );
  AND2_X1 U12587 ( .A1(n12509), .A2(n12673), .ZN(n12671) );
  OR2_X1 U12588 ( .A1(n12512), .A2(n12511), .ZN(n12673) );
  OR2_X1 U12589 ( .A1(n12674), .A2(n12675), .ZN(n12511) );
  AND2_X1 U12590 ( .A1(n12508), .A2(n12507), .ZN(n12675) );
  AND2_X1 U12591 ( .A1(n12505), .A2(n12676), .ZN(n12674) );
  OR2_X1 U12592 ( .A1(n12508), .A2(n12507), .ZN(n12676) );
  OR2_X1 U12593 ( .A1(n12677), .A2(n12678), .ZN(n12507) );
  AND2_X1 U12594 ( .A1(n12504), .A2(n12503), .ZN(n12678) );
  AND2_X1 U12595 ( .A1(n12501), .A2(n12679), .ZN(n12677) );
  OR2_X1 U12596 ( .A1(n12504), .A2(n12503), .ZN(n12679) );
  OR2_X1 U12597 ( .A1(n12680), .A2(n12681), .ZN(n12503) );
  AND2_X1 U12598 ( .A1(n12500), .A2(n12499), .ZN(n12681) );
  AND2_X1 U12599 ( .A1(n12497), .A2(n12682), .ZN(n12680) );
  OR2_X1 U12600 ( .A1(n12500), .A2(n12499), .ZN(n12682) );
  OR2_X1 U12601 ( .A1(n12683), .A2(n12684), .ZN(n12499) );
  AND2_X1 U12602 ( .A1(n12496), .A2(n12495), .ZN(n12684) );
  AND2_X1 U12603 ( .A1(n12493), .A2(n12685), .ZN(n12683) );
  OR2_X1 U12604 ( .A1(n12496), .A2(n12495), .ZN(n12685) );
  OR2_X1 U12605 ( .A1(n12686), .A2(n12687), .ZN(n12495) );
  AND2_X1 U12606 ( .A1(n12492), .A2(n12491), .ZN(n12687) );
  AND2_X1 U12607 ( .A1(n12489), .A2(n12688), .ZN(n12686) );
  OR2_X1 U12608 ( .A1(n12492), .A2(n12491), .ZN(n12688) );
  OR2_X1 U12609 ( .A1(n12689), .A2(n12690), .ZN(n12491) );
  AND2_X1 U12610 ( .A1(n12488), .A2(n12487), .ZN(n12690) );
  AND2_X1 U12611 ( .A1(n12485), .A2(n12691), .ZN(n12689) );
  OR2_X1 U12612 ( .A1(n12488), .A2(n12487), .ZN(n12691) );
  OR2_X1 U12613 ( .A1(n12692), .A2(n12693), .ZN(n12487) );
  AND2_X1 U12614 ( .A1(n12481), .A2(n12484), .ZN(n12693) );
  AND2_X1 U12615 ( .A1(n12694), .A2(n12695), .ZN(n12692) );
  OR2_X1 U12616 ( .A1(n12481), .A2(n12484), .ZN(n12695) );
  OR3_X1 U12617 ( .A1(n8062), .A2(n8067), .A3(n8981), .ZN(n12484) );
  OR2_X1 U12618 ( .A1(n8067), .A2(n8127), .ZN(n12481) );
  INV_X1 U12619 ( .A(n12483), .ZN(n12694) );
  OR2_X1 U12620 ( .A1(n12696), .A2(n12697), .ZN(n12483) );
  AND2_X1 U12621 ( .A1(b_12_), .A2(n12698), .ZN(n12697) );
  OR2_X1 U12622 ( .A1(n12699), .A2(n7598), .ZN(n12698) );
  AND2_X1 U12623 ( .A1(a_30_), .A2(n8058), .ZN(n12699) );
  AND2_X1 U12624 ( .A1(b_11_), .A2(n12700), .ZN(n12696) );
  OR2_X1 U12625 ( .A1(n12701), .A2(n7601), .ZN(n12700) );
  AND2_X1 U12626 ( .A1(a_31_), .A2(n8062), .ZN(n12701) );
  OR2_X1 U12627 ( .A1(n8067), .A2(n8124), .ZN(n12488) );
  XNOR2_X1 U12628 ( .A(n12702), .B(n12703), .ZN(n12485) );
  XOR2_X1 U12629 ( .A(n12704), .B(n12705), .Z(n12703) );
  OR2_X1 U12630 ( .A1(n8067), .A2(n8121), .ZN(n12492) );
  XOR2_X1 U12631 ( .A(n12706), .B(n12707), .Z(n12489) );
  XOR2_X1 U12632 ( .A(n12708), .B(n12709), .Z(n12707) );
  OR2_X1 U12633 ( .A1(n8067), .A2(n8118), .ZN(n12496) );
  XOR2_X1 U12634 ( .A(n12710), .B(n12711), .Z(n12493) );
  XOR2_X1 U12635 ( .A(n12712), .B(n12713), .Z(n12711) );
  OR2_X1 U12636 ( .A1(n8067), .A2(n8115), .ZN(n12500) );
  XOR2_X1 U12637 ( .A(n12714), .B(n12715), .Z(n12497) );
  XOR2_X1 U12638 ( .A(n12716), .B(n12717), .Z(n12715) );
  OR2_X1 U12639 ( .A1(n8067), .A2(n8112), .ZN(n12504) );
  XOR2_X1 U12640 ( .A(n12718), .B(n12719), .Z(n12501) );
  XOR2_X1 U12641 ( .A(n12720), .B(n12721), .Z(n12719) );
  OR2_X1 U12642 ( .A1(n8067), .A2(n8109), .ZN(n12508) );
  XOR2_X1 U12643 ( .A(n12722), .B(n12723), .Z(n12505) );
  XOR2_X1 U12644 ( .A(n12724), .B(n12725), .Z(n12723) );
  OR2_X1 U12645 ( .A1(n8067), .A2(n8106), .ZN(n12512) );
  XOR2_X1 U12646 ( .A(n12726), .B(n12727), .Z(n12509) );
  XOR2_X1 U12647 ( .A(n12728), .B(n12729), .Z(n12727) );
  OR2_X1 U12648 ( .A1(n8067), .A2(n8102), .ZN(n12516) );
  XOR2_X1 U12649 ( .A(n12730), .B(n12731), .Z(n12513) );
  XOR2_X1 U12650 ( .A(n12732), .B(n12733), .Z(n12731) );
  OR2_X1 U12651 ( .A1(n8067), .A2(n8097), .ZN(n12520) );
  XOR2_X1 U12652 ( .A(n12734), .B(n12735), .Z(n12517) );
  XOR2_X1 U12653 ( .A(n12736), .B(n12737), .Z(n12735) );
  OR2_X1 U12654 ( .A1(n8067), .A2(n8093), .ZN(n12524) );
  XOR2_X1 U12655 ( .A(n12738), .B(n12739), .Z(n12521) );
  XOR2_X1 U12656 ( .A(n12740), .B(n12741), .Z(n12739) );
  OR2_X1 U12657 ( .A1(n8067), .A2(n8088), .ZN(n12528) );
  XOR2_X1 U12658 ( .A(n12742), .B(n12743), .Z(n12525) );
  XOR2_X1 U12659 ( .A(n12744), .B(n12745), .Z(n12743) );
  OR2_X1 U12660 ( .A1(n8067), .A2(n8084), .ZN(n12532) );
  XOR2_X1 U12661 ( .A(n12746), .B(n12747), .Z(n12529) );
  XOR2_X1 U12662 ( .A(n12748), .B(n12749), .Z(n12747) );
  OR2_X1 U12663 ( .A1(n8067), .A2(n8079), .ZN(n12536) );
  XOR2_X1 U12664 ( .A(n12750), .B(n12751), .Z(n12533) );
  XOR2_X1 U12665 ( .A(n12752), .B(n12753), .Z(n12751) );
  OR2_X1 U12666 ( .A1(n8067), .A2(n8075), .ZN(n12540) );
  XOR2_X1 U12667 ( .A(n12754), .B(n12755), .Z(n12537) );
  XOR2_X1 U12668 ( .A(n12756), .B(n12757), .Z(n12755) );
  OR2_X1 U12669 ( .A1(n8067), .A2(n8070), .ZN(n12544) );
  XOR2_X1 U12670 ( .A(n12758), .B(n12759), .Z(n12541) );
  XOR2_X1 U12671 ( .A(n12760), .B(n12761), .Z(n12759) );
  OR2_X1 U12672 ( .A1(n8066), .A2(n8067), .ZN(n8068) );
  XOR2_X1 U12673 ( .A(n12762), .B(n12763), .Z(n12545) );
  XOR2_X1 U12674 ( .A(n12764), .B(n12765), .Z(n12763) );
  OR2_X1 U12675 ( .A1(n8067), .A2(n8061), .ZN(n12551) );
  XOR2_X1 U12676 ( .A(n12766), .B(n12767), .Z(n12548) );
  XOR2_X1 U12677 ( .A(n12768), .B(n12769), .Z(n12767) );
  OR2_X1 U12678 ( .A1(n8057), .A2(n8067), .ZN(n12555) );
  XNOR2_X1 U12679 ( .A(n12770), .B(n12771), .ZN(n12552) );
  XOR2_X1 U12680 ( .A(n7857), .B(n12772), .Z(n12770) );
  INV_X1 U12681 ( .A(n8063), .ZN(n7857) );
  OR2_X1 U12682 ( .A1(n8067), .A2(n8052), .ZN(n12559) );
  XOR2_X1 U12683 ( .A(n12773), .B(n12774), .Z(n12556) );
  XOR2_X1 U12684 ( .A(n12775), .B(n12776), .Z(n12774) );
  OR2_X1 U12685 ( .A1(n8048), .A2(n8067), .ZN(n12563) );
  XOR2_X1 U12686 ( .A(n12777), .B(n12778), .Z(n12560) );
  XOR2_X1 U12687 ( .A(n12779), .B(n12780), .Z(n12778) );
  OR2_X1 U12688 ( .A1(n8067), .A2(n8043), .ZN(n12567) );
  XOR2_X1 U12689 ( .A(n12781), .B(n12782), .Z(n12564) );
  XOR2_X1 U12690 ( .A(n12783), .B(n12784), .Z(n12782) );
  OR2_X1 U12691 ( .A1(n8039), .A2(n8067), .ZN(n12571) );
  XOR2_X1 U12692 ( .A(n12785), .B(n12786), .Z(n12568) );
  XOR2_X1 U12693 ( .A(n12787), .B(n12788), .Z(n12786) );
  OR2_X1 U12694 ( .A1(n8067), .A2(n8034), .ZN(n12575) );
  XOR2_X1 U12695 ( .A(n12789), .B(n12790), .Z(n12572) );
  XOR2_X1 U12696 ( .A(n12791), .B(n12792), .Z(n12790) );
  OR2_X1 U12697 ( .A1(n8030), .A2(n8067), .ZN(n12579) );
  XOR2_X1 U12698 ( .A(n12793), .B(n12794), .Z(n12576) );
  XOR2_X1 U12699 ( .A(n12795), .B(n12796), .Z(n12794) );
  OR2_X1 U12700 ( .A1(n8067), .A2(n8025), .ZN(n12583) );
  XOR2_X1 U12701 ( .A(n12797), .B(n12798), .Z(n12580) );
  XOR2_X1 U12702 ( .A(n12799), .B(n12800), .Z(n12798) );
  OR2_X1 U12703 ( .A1(n8021), .A2(n8067), .ZN(n12587) );
  XOR2_X1 U12704 ( .A(n12801), .B(n12802), .Z(n12584) );
  XOR2_X1 U12705 ( .A(n12803), .B(n12804), .Z(n12802) );
  OR2_X1 U12706 ( .A1(n8067), .A2(n8016), .ZN(n12591) );
  XOR2_X1 U12707 ( .A(n12805), .B(n12806), .Z(n12588) );
  XOR2_X1 U12708 ( .A(n12807), .B(n12808), .Z(n12806) );
  OR2_X1 U12709 ( .A1(n8067), .A2(n8012), .ZN(n12595) );
  XOR2_X1 U12710 ( .A(n12809), .B(n12810), .Z(n12592) );
  XOR2_X1 U12711 ( .A(n12811), .B(n12812), .Z(n12810) );
  OR2_X1 U12712 ( .A1(n8067), .A2(n8297), .ZN(n12599) );
  XOR2_X1 U12713 ( .A(n12813), .B(n12814), .Z(n12596) );
  XOR2_X1 U12714 ( .A(n12815), .B(n12816), .Z(n12814) );
  XOR2_X1 U12715 ( .A(n8593), .B(n12817), .Z(n12603) );
  XOR2_X1 U12716 ( .A(n8592), .B(n8591), .Z(n12817) );
  OR2_X1 U12717 ( .A1(n8062), .A2(n8297), .ZN(n8591) );
  OR2_X1 U12718 ( .A1(n12818), .A2(n12819), .ZN(n8592) );
  AND2_X1 U12719 ( .A1(n12816), .A2(n12815), .ZN(n12819) );
  AND2_X1 U12720 ( .A1(n12813), .A2(n12820), .ZN(n12818) );
  OR2_X1 U12721 ( .A1(n12815), .A2(n12816), .ZN(n12820) );
  OR2_X1 U12722 ( .A1(n8062), .A2(n8012), .ZN(n12816) );
  OR2_X1 U12723 ( .A1(n12821), .A2(n12822), .ZN(n12815) );
  AND2_X1 U12724 ( .A1(n12812), .A2(n12811), .ZN(n12822) );
  AND2_X1 U12725 ( .A1(n12809), .A2(n12823), .ZN(n12821) );
  OR2_X1 U12726 ( .A1(n12811), .A2(n12812), .ZN(n12823) );
  OR2_X1 U12727 ( .A1(n8062), .A2(n8016), .ZN(n12812) );
  OR2_X1 U12728 ( .A1(n12824), .A2(n12825), .ZN(n12811) );
  AND2_X1 U12729 ( .A1(n12808), .A2(n12807), .ZN(n12825) );
  AND2_X1 U12730 ( .A1(n12805), .A2(n12826), .ZN(n12824) );
  OR2_X1 U12731 ( .A1(n12807), .A2(n12808), .ZN(n12826) );
  OR2_X1 U12732 ( .A1(n8021), .A2(n8062), .ZN(n12808) );
  OR2_X1 U12733 ( .A1(n12827), .A2(n12828), .ZN(n12807) );
  AND2_X1 U12734 ( .A1(n12804), .A2(n12803), .ZN(n12828) );
  AND2_X1 U12735 ( .A1(n12801), .A2(n12829), .ZN(n12827) );
  OR2_X1 U12736 ( .A1(n12803), .A2(n12804), .ZN(n12829) );
  OR2_X1 U12737 ( .A1(n8062), .A2(n8025), .ZN(n12804) );
  OR2_X1 U12738 ( .A1(n12830), .A2(n12831), .ZN(n12803) );
  AND2_X1 U12739 ( .A1(n12800), .A2(n12799), .ZN(n12831) );
  AND2_X1 U12740 ( .A1(n12797), .A2(n12832), .ZN(n12830) );
  OR2_X1 U12741 ( .A1(n12799), .A2(n12800), .ZN(n12832) );
  OR2_X1 U12742 ( .A1(n8030), .A2(n8062), .ZN(n12800) );
  OR2_X1 U12743 ( .A1(n12833), .A2(n12834), .ZN(n12799) );
  AND2_X1 U12744 ( .A1(n12796), .A2(n12795), .ZN(n12834) );
  AND2_X1 U12745 ( .A1(n12793), .A2(n12835), .ZN(n12833) );
  OR2_X1 U12746 ( .A1(n12795), .A2(n12796), .ZN(n12835) );
  OR2_X1 U12747 ( .A1(n8062), .A2(n8034), .ZN(n12796) );
  OR2_X1 U12748 ( .A1(n12836), .A2(n12837), .ZN(n12795) );
  AND2_X1 U12749 ( .A1(n12792), .A2(n12791), .ZN(n12837) );
  AND2_X1 U12750 ( .A1(n12789), .A2(n12838), .ZN(n12836) );
  OR2_X1 U12751 ( .A1(n12791), .A2(n12792), .ZN(n12838) );
  OR2_X1 U12752 ( .A1(n8039), .A2(n8062), .ZN(n12792) );
  OR2_X1 U12753 ( .A1(n12839), .A2(n12840), .ZN(n12791) );
  AND2_X1 U12754 ( .A1(n12788), .A2(n12787), .ZN(n12840) );
  AND2_X1 U12755 ( .A1(n12785), .A2(n12841), .ZN(n12839) );
  OR2_X1 U12756 ( .A1(n12787), .A2(n12788), .ZN(n12841) );
  OR2_X1 U12757 ( .A1(n8062), .A2(n8043), .ZN(n12788) );
  OR2_X1 U12758 ( .A1(n12842), .A2(n12843), .ZN(n12787) );
  AND2_X1 U12759 ( .A1(n12784), .A2(n12783), .ZN(n12843) );
  AND2_X1 U12760 ( .A1(n12781), .A2(n12844), .ZN(n12842) );
  OR2_X1 U12761 ( .A1(n12783), .A2(n12784), .ZN(n12844) );
  OR2_X1 U12762 ( .A1(n8048), .A2(n8062), .ZN(n12784) );
  OR2_X1 U12763 ( .A1(n12845), .A2(n12846), .ZN(n12783) );
  AND2_X1 U12764 ( .A1(n12780), .A2(n12779), .ZN(n12846) );
  AND2_X1 U12765 ( .A1(n12777), .A2(n12847), .ZN(n12845) );
  OR2_X1 U12766 ( .A1(n12779), .A2(n12780), .ZN(n12847) );
  OR2_X1 U12767 ( .A1(n8062), .A2(n8052), .ZN(n12780) );
  OR2_X1 U12768 ( .A1(n12848), .A2(n12849), .ZN(n12779) );
  AND2_X1 U12769 ( .A1(n12776), .A2(n12775), .ZN(n12849) );
  AND2_X1 U12770 ( .A1(n12773), .A2(n12850), .ZN(n12848) );
  OR2_X1 U12771 ( .A1(n12775), .A2(n12776), .ZN(n12850) );
  OR2_X1 U12772 ( .A1(n8057), .A2(n8062), .ZN(n12776) );
  OR2_X1 U12773 ( .A1(n12851), .A2(n12852), .ZN(n12775) );
  AND2_X1 U12774 ( .A1(n12772), .A2(n8063), .ZN(n12852) );
  AND2_X1 U12775 ( .A1(n12771), .A2(n12853), .ZN(n12851) );
  OR2_X1 U12776 ( .A1(n8063), .A2(n12772), .ZN(n12853) );
  OR2_X1 U12777 ( .A1(n12854), .A2(n12855), .ZN(n12772) );
  AND2_X1 U12778 ( .A1(n12769), .A2(n12768), .ZN(n12855) );
  AND2_X1 U12779 ( .A1(n12766), .A2(n12856), .ZN(n12854) );
  OR2_X1 U12780 ( .A1(n12768), .A2(n12769), .ZN(n12856) );
  OR2_X1 U12781 ( .A1(n8062), .A2(n8066), .ZN(n12769) );
  OR2_X1 U12782 ( .A1(n12857), .A2(n12858), .ZN(n12768) );
  AND2_X1 U12783 ( .A1(n12765), .A2(n12764), .ZN(n12858) );
  AND2_X1 U12784 ( .A1(n12762), .A2(n12859), .ZN(n12857) );
  OR2_X1 U12785 ( .A1(n12764), .A2(n12765), .ZN(n12859) );
  OR2_X1 U12786 ( .A1(n8062), .A2(n8070), .ZN(n12765) );
  OR2_X1 U12787 ( .A1(n12860), .A2(n12861), .ZN(n12764) );
  AND2_X1 U12788 ( .A1(n12761), .A2(n12760), .ZN(n12861) );
  AND2_X1 U12789 ( .A1(n12758), .A2(n12862), .ZN(n12860) );
  OR2_X1 U12790 ( .A1(n12760), .A2(n12761), .ZN(n12862) );
  OR2_X1 U12791 ( .A1(n8062), .A2(n8075), .ZN(n12761) );
  OR2_X1 U12792 ( .A1(n12863), .A2(n12864), .ZN(n12760) );
  AND2_X1 U12793 ( .A1(n12757), .A2(n12756), .ZN(n12864) );
  AND2_X1 U12794 ( .A1(n12754), .A2(n12865), .ZN(n12863) );
  OR2_X1 U12795 ( .A1(n12756), .A2(n12757), .ZN(n12865) );
  OR2_X1 U12796 ( .A1(n8062), .A2(n8079), .ZN(n12757) );
  OR2_X1 U12797 ( .A1(n12866), .A2(n12867), .ZN(n12756) );
  AND2_X1 U12798 ( .A1(n12753), .A2(n12752), .ZN(n12867) );
  AND2_X1 U12799 ( .A1(n12750), .A2(n12868), .ZN(n12866) );
  OR2_X1 U12800 ( .A1(n12752), .A2(n12753), .ZN(n12868) );
  OR2_X1 U12801 ( .A1(n8062), .A2(n8084), .ZN(n12753) );
  OR2_X1 U12802 ( .A1(n12869), .A2(n12870), .ZN(n12752) );
  AND2_X1 U12803 ( .A1(n12749), .A2(n12748), .ZN(n12870) );
  AND2_X1 U12804 ( .A1(n12746), .A2(n12871), .ZN(n12869) );
  OR2_X1 U12805 ( .A1(n12748), .A2(n12749), .ZN(n12871) );
  OR2_X1 U12806 ( .A1(n8062), .A2(n8088), .ZN(n12749) );
  OR2_X1 U12807 ( .A1(n12872), .A2(n12873), .ZN(n12748) );
  AND2_X1 U12808 ( .A1(n12745), .A2(n12744), .ZN(n12873) );
  AND2_X1 U12809 ( .A1(n12742), .A2(n12874), .ZN(n12872) );
  OR2_X1 U12810 ( .A1(n12744), .A2(n12745), .ZN(n12874) );
  OR2_X1 U12811 ( .A1(n8062), .A2(n8093), .ZN(n12745) );
  OR2_X1 U12812 ( .A1(n12875), .A2(n12876), .ZN(n12744) );
  AND2_X1 U12813 ( .A1(n12741), .A2(n12740), .ZN(n12876) );
  AND2_X1 U12814 ( .A1(n12738), .A2(n12877), .ZN(n12875) );
  OR2_X1 U12815 ( .A1(n12740), .A2(n12741), .ZN(n12877) );
  OR2_X1 U12816 ( .A1(n8062), .A2(n8097), .ZN(n12741) );
  OR2_X1 U12817 ( .A1(n12878), .A2(n12879), .ZN(n12740) );
  AND2_X1 U12818 ( .A1(n12737), .A2(n12736), .ZN(n12879) );
  AND2_X1 U12819 ( .A1(n12734), .A2(n12880), .ZN(n12878) );
  OR2_X1 U12820 ( .A1(n12736), .A2(n12737), .ZN(n12880) );
  OR2_X1 U12821 ( .A1(n8062), .A2(n8102), .ZN(n12737) );
  OR2_X1 U12822 ( .A1(n12881), .A2(n12882), .ZN(n12736) );
  AND2_X1 U12823 ( .A1(n12733), .A2(n12732), .ZN(n12882) );
  AND2_X1 U12824 ( .A1(n12730), .A2(n12883), .ZN(n12881) );
  OR2_X1 U12825 ( .A1(n12732), .A2(n12733), .ZN(n12883) );
  OR2_X1 U12826 ( .A1(n8062), .A2(n8106), .ZN(n12733) );
  OR2_X1 U12827 ( .A1(n12884), .A2(n12885), .ZN(n12732) );
  AND2_X1 U12828 ( .A1(n12729), .A2(n12728), .ZN(n12885) );
  AND2_X1 U12829 ( .A1(n12726), .A2(n12886), .ZN(n12884) );
  OR2_X1 U12830 ( .A1(n12728), .A2(n12729), .ZN(n12886) );
  OR2_X1 U12831 ( .A1(n8062), .A2(n8109), .ZN(n12729) );
  OR2_X1 U12832 ( .A1(n12887), .A2(n12888), .ZN(n12728) );
  AND2_X1 U12833 ( .A1(n12725), .A2(n12724), .ZN(n12888) );
  AND2_X1 U12834 ( .A1(n12722), .A2(n12889), .ZN(n12887) );
  OR2_X1 U12835 ( .A1(n12724), .A2(n12725), .ZN(n12889) );
  OR2_X1 U12836 ( .A1(n8062), .A2(n8112), .ZN(n12725) );
  OR2_X1 U12837 ( .A1(n12890), .A2(n12891), .ZN(n12724) );
  AND2_X1 U12838 ( .A1(n12721), .A2(n12720), .ZN(n12891) );
  AND2_X1 U12839 ( .A1(n12718), .A2(n12892), .ZN(n12890) );
  OR2_X1 U12840 ( .A1(n12720), .A2(n12721), .ZN(n12892) );
  OR2_X1 U12841 ( .A1(n8062), .A2(n8115), .ZN(n12721) );
  OR2_X1 U12842 ( .A1(n12893), .A2(n12894), .ZN(n12720) );
  AND2_X1 U12843 ( .A1(n12717), .A2(n12716), .ZN(n12894) );
  AND2_X1 U12844 ( .A1(n12714), .A2(n12895), .ZN(n12893) );
  OR2_X1 U12845 ( .A1(n12716), .A2(n12717), .ZN(n12895) );
  OR2_X1 U12846 ( .A1(n8062), .A2(n8118), .ZN(n12717) );
  OR2_X1 U12847 ( .A1(n12896), .A2(n12897), .ZN(n12716) );
  AND2_X1 U12848 ( .A1(n12713), .A2(n12712), .ZN(n12897) );
  AND2_X1 U12849 ( .A1(n12710), .A2(n12898), .ZN(n12896) );
  OR2_X1 U12850 ( .A1(n12712), .A2(n12713), .ZN(n12898) );
  OR2_X1 U12851 ( .A1(n8062), .A2(n8121), .ZN(n12713) );
  OR2_X1 U12852 ( .A1(n12899), .A2(n12900), .ZN(n12712) );
  AND2_X1 U12853 ( .A1(n12709), .A2(n12708), .ZN(n12900) );
  AND2_X1 U12854 ( .A1(n12706), .A2(n12901), .ZN(n12899) );
  OR2_X1 U12855 ( .A1(n12708), .A2(n12709), .ZN(n12901) );
  OR2_X1 U12856 ( .A1(n8062), .A2(n8124), .ZN(n12709) );
  OR2_X1 U12857 ( .A1(n12902), .A2(n12903), .ZN(n12708) );
  AND2_X1 U12858 ( .A1(n12702), .A2(n12705), .ZN(n12903) );
  AND2_X1 U12859 ( .A1(n12904), .A2(n12905), .ZN(n12902) );
  OR2_X1 U12860 ( .A1(n12705), .A2(n12702), .ZN(n12905) );
  OR2_X1 U12861 ( .A1(n8062), .A2(n8127), .ZN(n12702) );
  OR3_X1 U12862 ( .A1(n8058), .A2(n8062), .A3(n8981), .ZN(n12705) );
  INV_X1 U12863 ( .A(n12704), .ZN(n12904) );
  OR2_X1 U12864 ( .A1(n12906), .A2(n12907), .ZN(n12704) );
  AND2_X1 U12865 ( .A1(b_11_), .A2(n12908), .ZN(n12907) );
  OR2_X1 U12866 ( .A1(n12909), .A2(n7598), .ZN(n12908) );
  AND2_X1 U12867 ( .A1(a_30_), .A2(n8053), .ZN(n12909) );
  AND2_X1 U12868 ( .A1(b_10_), .A2(n12910), .ZN(n12906) );
  OR2_X1 U12869 ( .A1(n12911), .A2(n7601), .ZN(n12910) );
  AND2_X1 U12870 ( .A1(a_31_), .A2(n8058), .ZN(n12911) );
  XNOR2_X1 U12871 ( .A(n12912), .B(n12913), .ZN(n12706) );
  XOR2_X1 U12872 ( .A(n12914), .B(n12915), .Z(n12913) );
  XOR2_X1 U12873 ( .A(n12916), .B(n12917), .Z(n12710) );
  XOR2_X1 U12874 ( .A(n12918), .B(n12919), .Z(n12917) );
  XOR2_X1 U12875 ( .A(n12920), .B(n12921), .Z(n12714) );
  XOR2_X1 U12876 ( .A(n12922), .B(n12923), .Z(n12921) );
  XOR2_X1 U12877 ( .A(n12924), .B(n12925), .Z(n12718) );
  XOR2_X1 U12878 ( .A(n12926), .B(n12927), .Z(n12925) );
  XOR2_X1 U12879 ( .A(n12928), .B(n12929), .Z(n12722) );
  XOR2_X1 U12880 ( .A(n12930), .B(n12931), .Z(n12929) );
  XOR2_X1 U12881 ( .A(n12932), .B(n12933), .Z(n12726) );
  XOR2_X1 U12882 ( .A(n12934), .B(n12935), .Z(n12933) );
  XOR2_X1 U12883 ( .A(n12936), .B(n12937), .Z(n12730) );
  XOR2_X1 U12884 ( .A(n12938), .B(n12939), .Z(n12937) );
  XOR2_X1 U12885 ( .A(n12940), .B(n12941), .Z(n12734) );
  XOR2_X1 U12886 ( .A(n12942), .B(n12943), .Z(n12941) );
  XOR2_X1 U12887 ( .A(n12944), .B(n12945), .Z(n12738) );
  XOR2_X1 U12888 ( .A(n12946), .B(n12947), .Z(n12945) );
  XOR2_X1 U12889 ( .A(n12948), .B(n12949), .Z(n12742) );
  XOR2_X1 U12890 ( .A(n12950), .B(n12951), .Z(n12949) );
  XOR2_X1 U12891 ( .A(n12952), .B(n12953), .Z(n12746) );
  XOR2_X1 U12892 ( .A(n12954), .B(n12955), .Z(n12953) );
  XOR2_X1 U12893 ( .A(n12956), .B(n12957), .Z(n12750) );
  XOR2_X1 U12894 ( .A(n12958), .B(n12959), .Z(n12957) );
  XOR2_X1 U12895 ( .A(n12960), .B(n12961), .Z(n12754) );
  XOR2_X1 U12896 ( .A(n12962), .B(n12963), .Z(n12961) );
  XOR2_X1 U12897 ( .A(n12964), .B(n12965), .Z(n12758) );
  XOR2_X1 U12898 ( .A(n12966), .B(n12967), .Z(n12965) );
  XOR2_X1 U12899 ( .A(n12968), .B(n12969), .Z(n12762) );
  XOR2_X1 U12900 ( .A(n12970), .B(n12971), .Z(n12969) );
  XOR2_X1 U12901 ( .A(n12972), .B(n12973), .Z(n12766) );
  XOR2_X1 U12902 ( .A(n12974), .B(n12975), .Z(n12973) );
  OR2_X1 U12903 ( .A1(n8062), .A2(n8061), .ZN(n8063) );
  INV_X1 U12904 ( .A(b_12_), .ZN(n8062) );
  XOR2_X1 U12905 ( .A(n12976), .B(n12977), .Z(n12771) );
  XOR2_X1 U12906 ( .A(n12978), .B(n12979), .Z(n12977) );
  XOR2_X1 U12907 ( .A(n12980), .B(n12981), .Z(n12773) );
  XOR2_X1 U12908 ( .A(n12982), .B(n12983), .Z(n12981) );
  XOR2_X1 U12909 ( .A(n12984), .B(n12985), .Z(n12777) );
  XOR2_X1 U12910 ( .A(n12986), .B(n8059), .Z(n12985) );
  XOR2_X1 U12911 ( .A(n12987), .B(n12988), .Z(n12781) );
  XOR2_X1 U12912 ( .A(n12989), .B(n12990), .Z(n12988) );
  XOR2_X1 U12913 ( .A(n12991), .B(n12992), .Z(n12785) );
  XOR2_X1 U12914 ( .A(n12993), .B(n12994), .Z(n12992) );
  XOR2_X1 U12915 ( .A(n12995), .B(n12996), .Z(n12789) );
  XOR2_X1 U12916 ( .A(n12997), .B(n12998), .Z(n12996) );
  XOR2_X1 U12917 ( .A(n12999), .B(n13000), .Z(n12793) );
  XOR2_X1 U12918 ( .A(n13001), .B(n13002), .Z(n13000) );
  XOR2_X1 U12919 ( .A(n13003), .B(n13004), .Z(n12797) );
  XOR2_X1 U12920 ( .A(n13005), .B(n13006), .Z(n13004) );
  XOR2_X1 U12921 ( .A(n13007), .B(n13008), .Z(n12801) );
  XOR2_X1 U12922 ( .A(n13009), .B(n13010), .Z(n13008) );
  XOR2_X1 U12923 ( .A(n13011), .B(n13012), .Z(n12805) );
  XOR2_X1 U12924 ( .A(n13013), .B(n13014), .Z(n13012) );
  XOR2_X1 U12925 ( .A(n13015), .B(n13016), .Z(n12809) );
  XOR2_X1 U12926 ( .A(n13017), .B(n13018), .Z(n13016) );
  XOR2_X1 U12927 ( .A(n13019), .B(n13020), .Z(n12813) );
  XOR2_X1 U12928 ( .A(n13021), .B(n13022), .Z(n13020) );
  XOR2_X1 U12929 ( .A(n13023), .B(n13024), .Z(n8593) );
  XOR2_X1 U12930 ( .A(n13025), .B(n13026), .Z(n13024) );
  INV_X1 U12931 ( .A(n8584), .ZN(n8580) );
  OR2_X1 U12932 ( .A1(n8586), .A2(n8587), .ZN(n8584) );
  OR2_X1 U12933 ( .A1(n13027), .A2(n13028), .ZN(n8587) );
  AND2_X1 U12934 ( .A1(n8598), .A2(n8597), .ZN(n13028) );
  AND2_X1 U12935 ( .A1(n8595), .A2(n13029), .ZN(n13027) );
  OR2_X1 U12936 ( .A1(n8598), .A2(n8597), .ZN(n13029) );
  OR2_X1 U12937 ( .A1(n13030), .A2(n13031), .ZN(n8597) );
  AND2_X1 U12938 ( .A1(n13026), .A2(n13025), .ZN(n13031) );
  AND2_X1 U12939 ( .A1(n13023), .A2(n13032), .ZN(n13030) );
  OR2_X1 U12940 ( .A1(n13026), .A2(n13025), .ZN(n13032) );
  OR2_X1 U12941 ( .A1(n13033), .A2(n13034), .ZN(n13025) );
  AND2_X1 U12942 ( .A1(n13022), .A2(n13021), .ZN(n13034) );
  AND2_X1 U12943 ( .A1(n13019), .A2(n13035), .ZN(n13033) );
  OR2_X1 U12944 ( .A1(n13022), .A2(n13021), .ZN(n13035) );
  OR2_X1 U12945 ( .A1(n13036), .A2(n13037), .ZN(n13021) );
  AND2_X1 U12946 ( .A1(n13018), .A2(n13017), .ZN(n13037) );
  AND2_X1 U12947 ( .A1(n13015), .A2(n13038), .ZN(n13036) );
  OR2_X1 U12948 ( .A1(n13018), .A2(n13017), .ZN(n13038) );
  OR2_X1 U12949 ( .A1(n13039), .A2(n13040), .ZN(n13017) );
  AND2_X1 U12950 ( .A1(n13014), .A2(n13013), .ZN(n13040) );
  AND2_X1 U12951 ( .A1(n13011), .A2(n13041), .ZN(n13039) );
  OR2_X1 U12952 ( .A1(n13014), .A2(n13013), .ZN(n13041) );
  OR2_X1 U12953 ( .A1(n13042), .A2(n13043), .ZN(n13013) );
  AND2_X1 U12954 ( .A1(n13010), .A2(n13009), .ZN(n13043) );
  AND2_X1 U12955 ( .A1(n13007), .A2(n13044), .ZN(n13042) );
  OR2_X1 U12956 ( .A1(n13010), .A2(n13009), .ZN(n13044) );
  OR2_X1 U12957 ( .A1(n13045), .A2(n13046), .ZN(n13009) );
  AND2_X1 U12958 ( .A1(n13006), .A2(n13005), .ZN(n13046) );
  AND2_X1 U12959 ( .A1(n13003), .A2(n13047), .ZN(n13045) );
  OR2_X1 U12960 ( .A1(n13006), .A2(n13005), .ZN(n13047) );
  OR2_X1 U12961 ( .A1(n13048), .A2(n13049), .ZN(n13005) );
  AND2_X1 U12962 ( .A1(n13002), .A2(n13001), .ZN(n13049) );
  AND2_X1 U12963 ( .A1(n12999), .A2(n13050), .ZN(n13048) );
  OR2_X1 U12964 ( .A1(n13002), .A2(n13001), .ZN(n13050) );
  OR2_X1 U12965 ( .A1(n13051), .A2(n13052), .ZN(n13001) );
  AND2_X1 U12966 ( .A1(n12998), .A2(n12997), .ZN(n13052) );
  AND2_X1 U12967 ( .A1(n12995), .A2(n13053), .ZN(n13051) );
  OR2_X1 U12968 ( .A1(n12998), .A2(n12997), .ZN(n13053) );
  OR2_X1 U12969 ( .A1(n13054), .A2(n13055), .ZN(n12997) );
  AND2_X1 U12970 ( .A1(n12994), .A2(n12993), .ZN(n13055) );
  AND2_X1 U12971 ( .A1(n12991), .A2(n13056), .ZN(n13054) );
  OR2_X1 U12972 ( .A1(n12994), .A2(n12993), .ZN(n13056) );
  OR2_X1 U12973 ( .A1(n13057), .A2(n13058), .ZN(n12993) );
  AND2_X1 U12974 ( .A1(n12990), .A2(n12989), .ZN(n13058) );
  AND2_X1 U12975 ( .A1(n12987), .A2(n13059), .ZN(n13057) );
  OR2_X1 U12976 ( .A1(n12990), .A2(n12989), .ZN(n13059) );
  OR2_X1 U12977 ( .A1(n13060), .A2(n13061), .ZN(n12989) );
  AND2_X1 U12978 ( .A1(n8059), .A2(n12986), .ZN(n13061) );
  AND2_X1 U12979 ( .A1(n12984), .A2(n13062), .ZN(n13060) );
  OR2_X1 U12980 ( .A1(n8059), .A2(n12986), .ZN(n13062) );
  OR2_X1 U12981 ( .A1(n13063), .A2(n13064), .ZN(n12986) );
  AND2_X1 U12982 ( .A1(n12983), .A2(n12982), .ZN(n13064) );
  AND2_X1 U12983 ( .A1(n12980), .A2(n13065), .ZN(n13063) );
  OR2_X1 U12984 ( .A1(n12983), .A2(n12982), .ZN(n13065) );
  OR2_X1 U12985 ( .A1(n13066), .A2(n13067), .ZN(n12982) );
  AND2_X1 U12986 ( .A1(n12979), .A2(n12978), .ZN(n13067) );
  AND2_X1 U12987 ( .A1(n12976), .A2(n13068), .ZN(n13066) );
  OR2_X1 U12988 ( .A1(n12979), .A2(n12978), .ZN(n13068) );
  OR2_X1 U12989 ( .A1(n13069), .A2(n13070), .ZN(n12978) );
  AND2_X1 U12990 ( .A1(n12975), .A2(n12974), .ZN(n13070) );
  AND2_X1 U12991 ( .A1(n12972), .A2(n13071), .ZN(n13069) );
  OR2_X1 U12992 ( .A1(n12975), .A2(n12974), .ZN(n13071) );
  OR2_X1 U12993 ( .A1(n13072), .A2(n13073), .ZN(n12974) );
  AND2_X1 U12994 ( .A1(n12971), .A2(n12970), .ZN(n13073) );
  AND2_X1 U12995 ( .A1(n12968), .A2(n13074), .ZN(n13072) );
  OR2_X1 U12996 ( .A1(n12971), .A2(n12970), .ZN(n13074) );
  OR2_X1 U12997 ( .A1(n13075), .A2(n13076), .ZN(n12970) );
  AND2_X1 U12998 ( .A1(n12967), .A2(n12966), .ZN(n13076) );
  AND2_X1 U12999 ( .A1(n12964), .A2(n13077), .ZN(n13075) );
  OR2_X1 U13000 ( .A1(n12967), .A2(n12966), .ZN(n13077) );
  OR2_X1 U13001 ( .A1(n13078), .A2(n13079), .ZN(n12966) );
  AND2_X1 U13002 ( .A1(n12963), .A2(n12962), .ZN(n13079) );
  AND2_X1 U13003 ( .A1(n12960), .A2(n13080), .ZN(n13078) );
  OR2_X1 U13004 ( .A1(n12963), .A2(n12962), .ZN(n13080) );
  OR2_X1 U13005 ( .A1(n13081), .A2(n13082), .ZN(n12962) );
  AND2_X1 U13006 ( .A1(n12959), .A2(n12958), .ZN(n13082) );
  AND2_X1 U13007 ( .A1(n12956), .A2(n13083), .ZN(n13081) );
  OR2_X1 U13008 ( .A1(n12959), .A2(n12958), .ZN(n13083) );
  OR2_X1 U13009 ( .A1(n13084), .A2(n13085), .ZN(n12958) );
  AND2_X1 U13010 ( .A1(n12955), .A2(n12954), .ZN(n13085) );
  AND2_X1 U13011 ( .A1(n12952), .A2(n13086), .ZN(n13084) );
  OR2_X1 U13012 ( .A1(n12955), .A2(n12954), .ZN(n13086) );
  OR2_X1 U13013 ( .A1(n13087), .A2(n13088), .ZN(n12954) );
  AND2_X1 U13014 ( .A1(n12951), .A2(n12950), .ZN(n13088) );
  AND2_X1 U13015 ( .A1(n12948), .A2(n13089), .ZN(n13087) );
  OR2_X1 U13016 ( .A1(n12951), .A2(n12950), .ZN(n13089) );
  OR2_X1 U13017 ( .A1(n13090), .A2(n13091), .ZN(n12950) );
  AND2_X1 U13018 ( .A1(n12947), .A2(n12946), .ZN(n13091) );
  AND2_X1 U13019 ( .A1(n12944), .A2(n13092), .ZN(n13090) );
  OR2_X1 U13020 ( .A1(n12947), .A2(n12946), .ZN(n13092) );
  OR2_X1 U13021 ( .A1(n13093), .A2(n13094), .ZN(n12946) );
  AND2_X1 U13022 ( .A1(n12943), .A2(n12942), .ZN(n13094) );
  AND2_X1 U13023 ( .A1(n12940), .A2(n13095), .ZN(n13093) );
  OR2_X1 U13024 ( .A1(n12943), .A2(n12942), .ZN(n13095) );
  OR2_X1 U13025 ( .A1(n13096), .A2(n13097), .ZN(n12942) );
  AND2_X1 U13026 ( .A1(n12939), .A2(n12938), .ZN(n13097) );
  AND2_X1 U13027 ( .A1(n12936), .A2(n13098), .ZN(n13096) );
  OR2_X1 U13028 ( .A1(n12939), .A2(n12938), .ZN(n13098) );
  OR2_X1 U13029 ( .A1(n13099), .A2(n13100), .ZN(n12938) );
  AND2_X1 U13030 ( .A1(n12935), .A2(n12934), .ZN(n13100) );
  AND2_X1 U13031 ( .A1(n12932), .A2(n13101), .ZN(n13099) );
  OR2_X1 U13032 ( .A1(n12935), .A2(n12934), .ZN(n13101) );
  OR2_X1 U13033 ( .A1(n13102), .A2(n13103), .ZN(n12934) );
  AND2_X1 U13034 ( .A1(n12931), .A2(n12930), .ZN(n13103) );
  AND2_X1 U13035 ( .A1(n12928), .A2(n13104), .ZN(n13102) );
  OR2_X1 U13036 ( .A1(n12931), .A2(n12930), .ZN(n13104) );
  OR2_X1 U13037 ( .A1(n13105), .A2(n13106), .ZN(n12930) );
  AND2_X1 U13038 ( .A1(n12927), .A2(n12926), .ZN(n13106) );
  AND2_X1 U13039 ( .A1(n12924), .A2(n13107), .ZN(n13105) );
  OR2_X1 U13040 ( .A1(n12927), .A2(n12926), .ZN(n13107) );
  OR2_X1 U13041 ( .A1(n13108), .A2(n13109), .ZN(n12926) );
  AND2_X1 U13042 ( .A1(n12923), .A2(n12922), .ZN(n13109) );
  AND2_X1 U13043 ( .A1(n12920), .A2(n13110), .ZN(n13108) );
  OR2_X1 U13044 ( .A1(n12923), .A2(n12922), .ZN(n13110) );
  OR2_X1 U13045 ( .A1(n13111), .A2(n13112), .ZN(n12922) );
  AND2_X1 U13046 ( .A1(n12919), .A2(n12918), .ZN(n13112) );
  AND2_X1 U13047 ( .A1(n12916), .A2(n13113), .ZN(n13111) );
  OR2_X1 U13048 ( .A1(n12919), .A2(n12918), .ZN(n13113) );
  OR2_X1 U13049 ( .A1(n13114), .A2(n13115), .ZN(n12918) );
  AND2_X1 U13050 ( .A1(n12912), .A2(n12915), .ZN(n13115) );
  AND2_X1 U13051 ( .A1(n13116), .A2(n13117), .ZN(n13114) );
  OR2_X1 U13052 ( .A1(n12912), .A2(n12915), .ZN(n13117) );
  OR3_X1 U13053 ( .A1(n8058), .A2(n8981), .A3(n8053), .ZN(n12915) );
  OR2_X1 U13054 ( .A1(n8058), .A2(n8127), .ZN(n12912) );
  INV_X1 U13055 ( .A(n12914), .ZN(n13116) );
  OR2_X1 U13056 ( .A1(n13118), .A2(n13119), .ZN(n12914) );
  AND2_X1 U13057 ( .A1(b_9_), .A2(n13120), .ZN(n13119) );
  OR2_X1 U13058 ( .A1(n13121), .A2(n7601), .ZN(n13120) );
  AND2_X1 U13059 ( .A1(a_31_), .A2(n8053), .ZN(n13121) );
  AND2_X1 U13060 ( .A1(b_10_), .A2(n13122), .ZN(n13118) );
  OR2_X1 U13061 ( .A1(n13123), .A2(n7598), .ZN(n13122) );
  AND2_X1 U13062 ( .A1(a_30_), .A2(n8049), .ZN(n13123) );
  OR2_X1 U13063 ( .A1(n8058), .A2(n8124), .ZN(n12919) );
  XNOR2_X1 U13064 ( .A(n13124), .B(n13125), .ZN(n12916) );
  XOR2_X1 U13065 ( .A(n13126), .B(n13127), .Z(n13125) );
  OR2_X1 U13066 ( .A1(n8058), .A2(n8121), .ZN(n12923) );
  XOR2_X1 U13067 ( .A(n13128), .B(n13129), .Z(n12920) );
  XOR2_X1 U13068 ( .A(n13130), .B(n13131), .Z(n13129) );
  OR2_X1 U13069 ( .A1(n8058), .A2(n8118), .ZN(n12927) );
  XOR2_X1 U13070 ( .A(n13132), .B(n13133), .Z(n12924) );
  XOR2_X1 U13071 ( .A(n13134), .B(n13135), .Z(n13133) );
  OR2_X1 U13072 ( .A1(n8058), .A2(n8115), .ZN(n12931) );
  XOR2_X1 U13073 ( .A(n13136), .B(n13137), .Z(n12928) );
  XOR2_X1 U13074 ( .A(n13138), .B(n13139), .Z(n13137) );
  OR2_X1 U13075 ( .A1(n8058), .A2(n8112), .ZN(n12935) );
  XOR2_X1 U13076 ( .A(n13140), .B(n13141), .Z(n12932) );
  XOR2_X1 U13077 ( .A(n13142), .B(n13143), .Z(n13141) );
  OR2_X1 U13078 ( .A1(n8058), .A2(n8109), .ZN(n12939) );
  XOR2_X1 U13079 ( .A(n13144), .B(n13145), .Z(n12936) );
  XOR2_X1 U13080 ( .A(n13146), .B(n13147), .Z(n13145) );
  OR2_X1 U13081 ( .A1(n8058), .A2(n8106), .ZN(n12943) );
  XOR2_X1 U13082 ( .A(n13148), .B(n13149), .Z(n12940) );
  XOR2_X1 U13083 ( .A(n13150), .B(n13151), .Z(n13149) );
  OR2_X1 U13084 ( .A1(n8058), .A2(n8102), .ZN(n12947) );
  XOR2_X1 U13085 ( .A(n13152), .B(n13153), .Z(n12944) );
  XOR2_X1 U13086 ( .A(n13154), .B(n13155), .Z(n13153) );
  OR2_X1 U13087 ( .A1(n8058), .A2(n8097), .ZN(n12951) );
  XOR2_X1 U13088 ( .A(n13156), .B(n13157), .Z(n12948) );
  XOR2_X1 U13089 ( .A(n13158), .B(n13159), .Z(n13157) );
  OR2_X1 U13090 ( .A1(n8058), .A2(n8093), .ZN(n12955) );
  XOR2_X1 U13091 ( .A(n13160), .B(n13161), .Z(n12952) );
  XOR2_X1 U13092 ( .A(n13162), .B(n13163), .Z(n13161) );
  OR2_X1 U13093 ( .A1(n8058), .A2(n8088), .ZN(n12959) );
  XOR2_X1 U13094 ( .A(n13164), .B(n13165), .Z(n12956) );
  XOR2_X1 U13095 ( .A(n13166), .B(n13167), .Z(n13165) );
  OR2_X1 U13096 ( .A1(n8058), .A2(n8084), .ZN(n12963) );
  XOR2_X1 U13097 ( .A(n13168), .B(n13169), .Z(n12960) );
  XOR2_X1 U13098 ( .A(n13170), .B(n13171), .Z(n13169) );
  OR2_X1 U13099 ( .A1(n8058), .A2(n8079), .ZN(n12967) );
  XOR2_X1 U13100 ( .A(n13172), .B(n13173), .Z(n12964) );
  XOR2_X1 U13101 ( .A(n13174), .B(n13175), .Z(n13173) );
  OR2_X1 U13102 ( .A1(n8058), .A2(n8075), .ZN(n12971) );
  XOR2_X1 U13103 ( .A(n13176), .B(n13177), .Z(n12968) );
  XOR2_X1 U13104 ( .A(n13178), .B(n13179), .Z(n13177) );
  OR2_X1 U13105 ( .A1(n8058), .A2(n8070), .ZN(n12975) );
  XOR2_X1 U13106 ( .A(n13180), .B(n13181), .Z(n12972) );
  XOR2_X1 U13107 ( .A(n13182), .B(n13183), .Z(n13181) );
  OR2_X1 U13108 ( .A1(n8058), .A2(n8066), .ZN(n12979) );
  XOR2_X1 U13109 ( .A(n13184), .B(n13185), .Z(n12976) );
  XOR2_X1 U13110 ( .A(n13186), .B(n13187), .Z(n13185) );
  OR2_X1 U13111 ( .A1(n8058), .A2(n8061), .ZN(n12983) );
  XOR2_X1 U13112 ( .A(n13188), .B(n13189), .Z(n12980) );
  XOR2_X1 U13113 ( .A(n13190), .B(n13191), .Z(n13189) );
  OR2_X1 U13114 ( .A1(n8057), .A2(n8058), .ZN(n8059) );
  XOR2_X1 U13115 ( .A(n13192), .B(n13193), .Z(n12984) );
  XOR2_X1 U13116 ( .A(n13194), .B(n13195), .Z(n13193) );
  OR2_X1 U13117 ( .A1(n8058), .A2(n8052), .ZN(n12990) );
  XOR2_X1 U13118 ( .A(n13196), .B(n13197), .Z(n12987) );
  XOR2_X1 U13119 ( .A(n13198), .B(n13199), .Z(n13197) );
  OR2_X1 U13120 ( .A1(n8048), .A2(n8058), .ZN(n12994) );
  XNOR2_X1 U13121 ( .A(n13200), .B(n13201), .ZN(n12991) );
  XOR2_X1 U13122 ( .A(n7881), .B(n13202), .Z(n13200) );
  INV_X1 U13123 ( .A(n8054), .ZN(n7881) );
  OR2_X1 U13124 ( .A1(n8058), .A2(n8043), .ZN(n12998) );
  XOR2_X1 U13125 ( .A(n13203), .B(n13204), .Z(n12995) );
  XOR2_X1 U13126 ( .A(n13205), .B(n13206), .Z(n13204) );
  OR2_X1 U13127 ( .A1(n8039), .A2(n8058), .ZN(n13002) );
  XOR2_X1 U13128 ( .A(n13207), .B(n13208), .Z(n12999) );
  XOR2_X1 U13129 ( .A(n13209), .B(n13210), .Z(n13208) );
  OR2_X1 U13130 ( .A1(n8058), .A2(n8034), .ZN(n13006) );
  XOR2_X1 U13131 ( .A(n13211), .B(n13212), .Z(n13003) );
  XOR2_X1 U13132 ( .A(n13213), .B(n13214), .Z(n13212) );
  OR2_X1 U13133 ( .A1(n8030), .A2(n8058), .ZN(n13010) );
  XOR2_X1 U13134 ( .A(n13215), .B(n13216), .Z(n13007) );
  XOR2_X1 U13135 ( .A(n13217), .B(n13218), .Z(n13216) );
  OR2_X1 U13136 ( .A1(n8058), .A2(n8025), .ZN(n13014) );
  XOR2_X1 U13137 ( .A(n13219), .B(n13220), .Z(n13011) );
  XOR2_X1 U13138 ( .A(n13221), .B(n13222), .Z(n13220) );
  OR2_X1 U13139 ( .A1(n8021), .A2(n8058), .ZN(n13018) );
  XOR2_X1 U13140 ( .A(n13223), .B(n13224), .Z(n13015) );
  XOR2_X1 U13141 ( .A(n13225), .B(n13226), .Z(n13224) );
  OR2_X1 U13142 ( .A1(n8058), .A2(n8016), .ZN(n13022) );
  XOR2_X1 U13143 ( .A(n13227), .B(n13228), .Z(n13019) );
  XOR2_X1 U13144 ( .A(n13229), .B(n13230), .Z(n13228) );
  OR2_X1 U13145 ( .A1(n8058), .A2(n8012), .ZN(n13026) );
  XOR2_X1 U13146 ( .A(n13231), .B(n13232), .Z(n13023) );
  XOR2_X1 U13147 ( .A(n13233), .B(n13234), .Z(n13232) );
  OR2_X1 U13148 ( .A1(n8058), .A2(n8297), .ZN(n8598) );
  XOR2_X1 U13149 ( .A(n13235), .B(n13236), .Z(n8595) );
  XOR2_X1 U13150 ( .A(n13237), .B(n13238), .Z(n13236) );
  XOR2_X1 U13151 ( .A(n8526), .B(n13239), .Z(n8586) );
  XOR2_X1 U13152 ( .A(n8525), .B(n8524), .Z(n13239) );
  OR2_X1 U13153 ( .A1(n8053), .A2(n8297), .ZN(n8524) );
  OR2_X1 U13154 ( .A1(n13240), .A2(n13241), .ZN(n8525) );
  AND2_X1 U13155 ( .A1(n13238), .A2(n13237), .ZN(n13241) );
  AND2_X1 U13156 ( .A1(n13235), .A2(n13242), .ZN(n13240) );
  OR2_X1 U13157 ( .A1(n13237), .A2(n13238), .ZN(n13242) );
  OR2_X1 U13158 ( .A1(n8053), .A2(n8012), .ZN(n13238) );
  OR2_X1 U13159 ( .A1(n13243), .A2(n13244), .ZN(n13237) );
  AND2_X1 U13160 ( .A1(n13234), .A2(n13233), .ZN(n13244) );
  AND2_X1 U13161 ( .A1(n13231), .A2(n13245), .ZN(n13243) );
  OR2_X1 U13162 ( .A1(n13233), .A2(n13234), .ZN(n13245) );
  OR2_X1 U13163 ( .A1(n8053), .A2(n8016), .ZN(n13234) );
  OR2_X1 U13164 ( .A1(n13246), .A2(n13247), .ZN(n13233) );
  AND2_X1 U13165 ( .A1(n13230), .A2(n13229), .ZN(n13247) );
  AND2_X1 U13166 ( .A1(n13227), .A2(n13248), .ZN(n13246) );
  OR2_X1 U13167 ( .A1(n13229), .A2(n13230), .ZN(n13248) );
  OR2_X1 U13168 ( .A1(n8021), .A2(n8053), .ZN(n13230) );
  OR2_X1 U13169 ( .A1(n13249), .A2(n13250), .ZN(n13229) );
  AND2_X1 U13170 ( .A1(n13226), .A2(n13225), .ZN(n13250) );
  AND2_X1 U13171 ( .A1(n13223), .A2(n13251), .ZN(n13249) );
  OR2_X1 U13172 ( .A1(n13225), .A2(n13226), .ZN(n13251) );
  OR2_X1 U13173 ( .A1(n8053), .A2(n8025), .ZN(n13226) );
  OR2_X1 U13174 ( .A1(n13252), .A2(n13253), .ZN(n13225) );
  AND2_X1 U13175 ( .A1(n13222), .A2(n13221), .ZN(n13253) );
  AND2_X1 U13176 ( .A1(n13219), .A2(n13254), .ZN(n13252) );
  OR2_X1 U13177 ( .A1(n13221), .A2(n13222), .ZN(n13254) );
  OR2_X1 U13178 ( .A1(n8030), .A2(n8053), .ZN(n13222) );
  OR2_X1 U13179 ( .A1(n13255), .A2(n13256), .ZN(n13221) );
  AND2_X1 U13180 ( .A1(n13218), .A2(n13217), .ZN(n13256) );
  AND2_X1 U13181 ( .A1(n13215), .A2(n13257), .ZN(n13255) );
  OR2_X1 U13182 ( .A1(n13217), .A2(n13218), .ZN(n13257) );
  OR2_X1 U13183 ( .A1(n8053), .A2(n8034), .ZN(n13218) );
  OR2_X1 U13184 ( .A1(n13258), .A2(n13259), .ZN(n13217) );
  AND2_X1 U13185 ( .A1(n13214), .A2(n13213), .ZN(n13259) );
  AND2_X1 U13186 ( .A1(n13211), .A2(n13260), .ZN(n13258) );
  OR2_X1 U13187 ( .A1(n13213), .A2(n13214), .ZN(n13260) );
  OR2_X1 U13188 ( .A1(n8039), .A2(n8053), .ZN(n13214) );
  OR2_X1 U13189 ( .A1(n13261), .A2(n13262), .ZN(n13213) );
  AND2_X1 U13190 ( .A1(n13210), .A2(n13209), .ZN(n13262) );
  AND2_X1 U13191 ( .A1(n13207), .A2(n13263), .ZN(n13261) );
  OR2_X1 U13192 ( .A1(n13209), .A2(n13210), .ZN(n13263) );
  OR2_X1 U13193 ( .A1(n8053), .A2(n8043), .ZN(n13210) );
  OR2_X1 U13194 ( .A1(n13264), .A2(n13265), .ZN(n13209) );
  AND2_X1 U13195 ( .A1(n13206), .A2(n13205), .ZN(n13265) );
  AND2_X1 U13196 ( .A1(n13203), .A2(n13266), .ZN(n13264) );
  OR2_X1 U13197 ( .A1(n13205), .A2(n13206), .ZN(n13266) );
  OR2_X1 U13198 ( .A1(n8048), .A2(n8053), .ZN(n13206) );
  OR2_X1 U13199 ( .A1(n13267), .A2(n13268), .ZN(n13205) );
  AND2_X1 U13200 ( .A1(n13202), .A2(n8054), .ZN(n13268) );
  AND2_X1 U13201 ( .A1(n13201), .A2(n13269), .ZN(n13267) );
  OR2_X1 U13202 ( .A1(n8054), .A2(n13202), .ZN(n13269) );
  OR2_X1 U13203 ( .A1(n13270), .A2(n13271), .ZN(n13202) );
  AND2_X1 U13204 ( .A1(n13199), .A2(n13198), .ZN(n13271) );
  AND2_X1 U13205 ( .A1(n13196), .A2(n13272), .ZN(n13270) );
  OR2_X1 U13206 ( .A1(n13198), .A2(n13199), .ZN(n13272) );
  OR2_X1 U13207 ( .A1(n8057), .A2(n8053), .ZN(n13199) );
  OR2_X1 U13208 ( .A1(n13273), .A2(n13274), .ZN(n13198) );
  AND2_X1 U13209 ( .A1(n13195), .A2(n13194), .ZN(n13274) );
  AND2_X1 U13210 ( .A1(n13192), .A2(n13275), .ZN(n13273) );
  OR2_X1 U13211 ( .A1(n13194), .A2(n13195), .ZN(n13275) );
  OR2_X1 U13212 ( .A1(n8061), .A2(n8053), .ZN(n13195) );
  OR2_X1 U13213 ( .A1(n13276), .A2(n13277), .ZN(n13194) );
  AND2_X1 U13214 ( .A1(n13191), .A2(n13190), .ZN(n13277) );
  AND2_X1 U13215 ( .A1(n13188), .A2(n13278), .ZN(n13276) );
  OR2_X1 U13216 ( .A1(n13190), .A2(n13191), .ZN(n13278) );
  OR2_X1 U13217 ( .A1(n8066), .A2(n8053), .ZN(n13191) );
  OR2_X1 U13218 ( .A1(n13279), .A2(n13280), .ZN(n13190) );
  AND2_X1 U13219 ( .A1(n13187), .A2(n13186), .ZN(n13280) );
  AND2_X1 U13220 ( .A1(n13184), .A2(n13281), .ZN(n13279) );
  OR2_X1 U13221 ( .A1(n13186), .A2(n13187), .ZN(n13281) );
  OR2_X1 U13222 ( .A1(n8070), .A2(n8053), .ZN(n13187) );
  OR2_X1 U13223 ( .A1(n13282), .A2(n13283), .ZN(n13186) );
  AND2_X1 U13224 ( .A1(n13183), .A2(n13182), .ZN(n13283) );
  AND2_X1 U13225 ( .A1(n13180), .A2(n13284), .ZN(n13282) );
  OR2_X1 U13226 ( .A1(n13182), .A2(n13183), .ZN(n13284) );
  OR2_X1 U13227 ( .A1(n8075), .A2(n8053), .ZN(n13183) );
  OR2_X1 U13228 ( .A1(n13285), .A2(n13286), .ZN(n13182) );
  AND2_X1 U13229 ( .A1(n13179), .A2(n13178), .ZN(n13286) );
  AND2_X1 U13230 ( .A1(n13176), .A2(n13287), .ZN(n13285) );
  OR2_X1 U13231 ( .A1(n13178), .A2(n13179), .ZN(n13287) );
  OR2_X1 U13232 ( .A1(n8079), .A2(n8053), .ZN(n13179) );
  OR2_X1 U13233 ( .A1(n13288), .A2(n13289), .ZN(n13178) );
  AND2_X1 U13234 ( .A1(n13175), .A2(n13174), .ZN(n13289) );
  AND2_X1 U13235 ( .A1(n13172), .A2(n13290), .ZN(n13288) );
  OR2_X1 U13236 ( .A1(n13174), .A2(n13175), .ZN(n13290) );
  OR2_X1 U13237 ( .A1(n8084), .A2(n8053), .ZN(n13175) );
  OR2_X1 U13238 ( .A1(n13291), .A2(n13292), .ZN(n13174) );
  AND2_X1 U13239 ( .A1(n13171), .A2(n13170), .ZN(n13292) );
  AND2_X1 U13240 ( .A1(n13168), .A2(n13293), .ZN(n13291) );
  OR2_X1 U13241 ( .A1(n13170), .A2(n13171), .ZN(n13293) );
  OR2_X1 U13242 ( .A1(n8088), .A2(n8053), .ZN(n13171) );
  OR2_X1 U13243 ( .A1(n13294), .A2(n13295), .ZN(n13170) );
  AND2_X1 U13244 ( .A1(n13164), .A2(n13167), .ZN(n13295) );
  AND2_X1 U13245 ( .A1(n13296), .A2(n13166), .ZN(n13294) );
  OR2_X1 U13246 ( .A1(n13297), .A2(n13298), .ZN(n13166) );
  AND2_X1 U13247 ( .A1(n13163), .A2(n13162), .ZN(n13298) );
  AND2_X1 U13248 ( .A1(n13160), .A2(n13299), .ZN(n13297) );
  OR2_X1 U13249 ( .A1(n13162), .A2(n13163), .ZN(n13299) );
  OR2_X1 U13250 ( .A1(n8097), .A2(n8053), .ZN(n13163) );
  OR2_X1 U13251 ( .A1(n13300), .A2(n13301), .ZN(n13162) );
  AND2_X1 U13252 ( .A1(n13156), .A2(n13159), .ZN(n13301) );
  AND2_X1 U13253 ( .A1(n13302), .A2(n13158), .ZN(n13300) );
  OR2_X1 U13254 ( .A1(n13303), .A2(n13304), .ZN(n13158) );
  AND2_X1 U13255 ( .A1(n13152), .A2(n13155), .ZN(n13304) );
  AND2_X1 U13256 ( .A1(n13305), .A2(n13154), .ZN(n13303) );
  OR2_X1 U13257 ( .A1(n13306), .A2(n13307), .ZN(n13154) );
  AND2_X1 U13258 ( .A1(n13148), .A2(n13151), .ZN(n13307) );
  AND2_X1 U13259 ( .A1(n13308), .A2(n13150), .ZN(n13306) );
  OR2_X1 U13260 ( .A1(n13309), .A2(n13310), .ZN(n13150) );
  AND2_X1 U13261 ( .A1(n13144), .A2(n13147), .ZN(n13310) );
  AND2_X1 U13262 ( .A1(n13311), .A2(n13146), .ZN(n13309) );
  OR2_X1 U13263 ( .A1(n13312), .A2(n13313), .ZN(n13146) );
  AND2_X1 U13264 ( .A1(n13140), .A2(n13143), .ZN(n13313) );
  AND2_X1 U13265 ( .A1(n13314), .A2(n13142), .ZN(n13312) );
  OR2_X1 U13266 ( .A1(n13315), .A2(n13316), .ZN(n13142) );
  AND2_X1 U13267 ( .A1(n13136), .A2(n13139), .ZN(n13316) );
  AND2_X1 U13268 ( .A1(n13317), .A2(n13138), .ZN(n13315) );
  OR2_X1 U13269 ( .A1(n13318), .A2(n13319), .ZN(n13138) );
  AND2_X1 U13270 ( .A1(n13132), .A2(n13135), .ZN(n13319) );
  AND2_X1 U13271 ( .A1(n13320), .A2(n13134), .ZN(n13318) );
  OR2_X1 U13272 ( .A1(n13321), .A2(n13322), .ZN(n13134) );
  AND2_X1 U13273 ( .A1(n13128), .A2(n13131), .ZN(n13322) );
  AND2_X1 U13274 ( .A1(n13323), .A2(n13130), .ZN(n13321) );
  OR2_X1 U13275 ( .A1(n13324), .A2(n13325), .ZN(n13130) );
  AND2_X1 U13276 ( .A1(n13124), .A2(n13127), .ZN(n13325) );
  AND2_X1 U13277 ( .A1(n13326), .A2(n13327), .ZN(n13324) );
  OR2_X1 U13278 ( .A1(n13127), .A2(n13124), .ZN(n13327) );
  OR2_X1 U13279 ( .A1(n8127), .A2(n8053), .ZN(n13124) );
  OR3_X1 U13280 ( .A1(n8981), .A2(n8049), .A3(n8053), .ZN(n13127) );
  INV_X1 U13281 ( .A(n13126), .ZN(n13326) );
  OR2_X1 U13282 ( .A1(n13328), .A2(n13329), .ZN(n13126) );
  AND2_X1 U13283 ( .A1(b_9_), .A2(n13330), .ZN(n13329) );
  OR2_X1 U13284 ( .A1(n13331), .A2(n7598), .ZN(n13330) );
  AND2_X1 U13285 ( .A1(a_30_), .A2(n8044), .ZN(n13331) );
  AND2_X1 U13286 ( .A1(b_8_), .A2(n13332), .ZN(n13328) );
  OR2_X1 U13287 ( .A1(n13333), .A2(n7601), .ZN(n13332) );
  AND2_X1 U13288 ( .A1(a_31_), .A2(n8049), .ZN(n13333) );
  OR2_X1 U13289 ( .A1(n13131), .A2(n13128), .ZN(n13323) );
  XNOR2_X1 U13290 ( .A(n13334), .B(n13335), .ZN(n13128) );
  XOR2_X1 U13291 ( .A(n13336), .B(n13337), .Z(n13335) );
  OR2_X1 U13292 ( .A1(n8124), .A2(n8053), .ZN(n13131) );
  OR2_X1 U13293 ( .A1(n13135), .A2(n13132), .ZN(n13320) );
  XOR2_X1 U13294 ( .A(n13338), .B(n13339), .Z(n13132) );
  XOR2_X1 U13295 ( .A(n13340), .B(n13341), .Z(n13339) );
  OR2_X1 U13296 ( .A1(n8121), .A2(n8053), .ZN(n13135) );
  OR2_X1 U13297 ( .A1(n13139), .A2(n13136), .ZN(n13317) );
  XOR2_X1 U13298 ( .A(n13342), .B(n13343), .Z(n13136) );
  XOR2_X1 U13299 ( .A(n13344), .B(n13345), .Z(n13343) );
  OR2_X1 U13300 ( .A1(n8118), .A2(n8053), .ZN(n13139) );
  OR2_X1 U13301 ( .A1(n13143), .A2(n13140), .ZN(n13314) );
  XOR2_X1 U13302 ( .A(n13346), .B(n13347), .Z(n13140) );
  XOR2_X1 U13303 ( .A(n13348), .B(n13349), .Z(n13347) );
  OR2_X1 U13304 ( .A1(n8115), .A2(n8053), .ZN(n13143) );
  OR2_X1 U13305 ( .A1(n13147), .A2(n13144), .ZN(n13311) );
  XOR2_X1 U13306 ( .A(n13350), .B(n13351), .Z(n13144) );
  XOR2_X1 U13307 ( .A(n13352), .B(n13353), .Z(n13351) );
  OR2_X1 U13308 ( .A1(n8112), .A2(n8053), .ZN(n13147) );
  OR2_X1 U13309 ( .A1(n13151), .A2(n13148), .ZN(n13308) );
  XOR2_X1 U13310 ( .A(n13354), .B(n13355), .Z(n13148) );
  XOR2_X1 U13311 ( .A(n13356), .B(n13357), .Z(n13355) );
  OR2_X1 U13312 ( .A1(n8109), .A2(n8053), .ZN(n13151) );
  OR2_X1 U13313 ( .A1(n13155), .A2(n13152), .ZN(n13305) );
  XOR2_X1 U13314 ( .A(n13358), .B(n13359), .Z(n13152) );
  XOR2_X1 U13315 ( .A(n13360), .B(n13361), .Z(n13359) );
  OR2_X1 U13316 ( .A1(n8106), .A2(n8053), .ZN(n13155) );
  OR2_X1 U13317 ( .A1(n13159), .A2(n13156), .ZN(n13302) );
  XOR2_X1 U13318 ( .A(n13362), .B(n13363), .Z(n13156) );
  XOR2_X1 U13319 ( .A(n13364), .B(n13365), .Z(n13363) );
  OR2_X1 U13320 ( .A1(n8102), .A2(n8053), .ZN(n13159) );
  XOR2_X1 U13321 ( .A(n13366), .B(n13367), .Z(n13160) );
  XOR2_X1 U13322 ( .A(n13368), .B(n13369), .Z(n13367) );
  OR2_X1 U13323 ( .A1(n13167), .A2(n13164), .ZN(n13296) );
  XOR2_X1 U13324 ( .A(n13370), .B(n13371), .Z(n13164) );
  XOR2_X1 U13325 ( .A(n13372), .B(n13373), .Z(n13371) );
  OR2_X1 U13326 ( .A1(n8093), .A2(n8053), .ZN(n13167) );
  XOR2_X1 U13327 ( .A(n13374), .B(n13375), .Z(n13168) );
  XOR2_X1 U13328 ( .A(n13376), .B(n13377), .Z(n13375) );
  XOR2_X1 U13329 ( .A(n13378), .B(n13379), .Z(n13172) );
  XOR2_X1 U13330 ( .A(n13380), .B(n13381), .Z(n13379) );
  XOR2_X1 U13331 ( .A(n13382), .B(n13383), .Z(n13176) );
  XOR2_X1 U13332 ( .A(n13384), .B(n13385), .Z(n13383) );
  XOR2_X1 U13333 ( .A(n13386), .B(n13387), .Z(n13180) );
  XOR2_X1 U13334 ( .A(n13388), .B(n13389), .Z(n13387) );
  XOR2_X1 U13335 ( .A(n13390), .B(n13391), .Z(n13184) );
  XOR2_X1 U13336 ( .A(n13392), .B(n13393), .Z(n13391) );
  XOR2_X1 U13337 ( .A(n13394), .B(n13395), .Z(n13188) );
  XOR2_X1 U13338 ( .A(n13396), .B(n13397), .Z(n13395) );
  XOR2_X1 U13339 ( .A(n13398), .B(n13399), .Z(n13192) );
  XOR2_X1 U13340 ( .A(n13400), .B(n13401), .Z(n13399) );
  XOR2_X1 U13341 ( .A(n13402), .B(n13403), .Z(n13196) );
  XOR2_X1 U13342 ( .A(n13404), .B(n13405), .Z(n13403) );
  OR2_X1 U13343 ( .A1(n8052), .A2(n8053), .ZN(n8054) );
  INV_X1 U13344 ( .A(b_10_), .ZN(n8053) );
  XOR2_X1 U13345 ( .A(n13406), .B(n13407), .Z(n13201) );
  XOR2_X1 U13346 ( .A(n13408), .B(n13409), .Z(n13407) );
  XOR2_X1 U13347 ( .A(n13410), .B(n13411), .Z(n13203) );
  XOR2_X1 U13348 ( .A(n13412), .B(n13413), .Z(n13411) );
  XOR2_X1 U13349 ( .A(n13414), .B(n13415), .Z(n13207) );
  XOR2_X1 U13350 ( .A(n13416), .B(n8050), .Z(n13415) );
  XOR2_X1 U13351 ( .A(n13417), .B(n13418), .Z(n13211) );
  XOR2_X1 U13352 ( .A(n13419), .B(n13420), .Z(n13418) );
  XOR2_X1 U13353 ( .A(n13421), .B(n13422), .Z(n13215) );
  XOR2_X1 U13354 ( .A(n13423), .B(n13424), .Z(n13422) );
  XOR2_X1 U13355 ( .A(n13425), .B(n13426), .Z(n13219) );
  XOR2_X1 U13356 ( .A(n13427), .B(n13428), .Z(n13426) );
  XOR2_X1 U13357 ( .A(n13429), .B(n13430), .Z(n13223) );
  XOR2_X1 U13358 ( .A(n13431), .B(n13432), .Z(n13430) );
  XOR2_X1 U13359 ( .A(n13433), .B(n13434), .Z(n13227) );
  XOR2_X1 U13360 ( .A(n13435), .B(n13436), .Z(n13434) );
  XOR2_X1 U13361 ( .A(n13437), .B(n13438), .Z(n13231) );
  XOR2_X1 U13362 ( .A(n13439), .B(n13440), .Z(n13438) );
  XOR2_X1 U13363 ( .A(n13441), .B(n13442), .Z(n13235) );
  XOR2_X1 U13364 ( .A(n13443), .B(n13444), .Z(n13442) );
  XOR2_X1 U13365 ( .A(n8533), .B(n13445), .Z(n8526) );
  XOR2_X1 U13366 ( .A(n8532), .B(n8531), .Z(n13445) );
  OR2_X1 U13367 ( .A1(n8049), .A2(n8012), .ZN(n8531) );
  OR2_X1 U13368 ( .A1(n13446), .A2(n13447), .ZN(n8532) );
  AND2_X1 U13369 ( .A1(n13444), .A2(n13443), .ZN(n13447) );
  AND2_X1 U13370 ( .A1(n13441), .A2(n13448), .ZN(n13446) );
  OR2_X1 U13371 ( .A1(n13443), .A2(n13444), .ZN(n13448) );
  OR2_X1 U13372 ( .A1(n8049), .A2(n8016), .ZN(n13444) );
  OR2_X1 U13373 ( .A1(n13449), .A2(n13450), .ZN(n13443) );
  AND2_X1 U13374 ( .A1(n13440), .A2(n13439), .ZN(n13450) );
  AND2_X1 U13375 ( .A1(n13437), .A2(n13451), .ZN(n13449) );
  OR2_X1 U13376 ( .A1(n13439), .A2(n13440), .ZN(n13451) );
  OR2_X1 U13377 ( .A1(n8021), .A2(n8049), .ZN(n13440) );
  OR2_X1 U13378 ( .A1(n13452), .A2(n13453), .ZN(n13439) );
  AND2_X1 U13379 ( .A1(n13436), .A2(n13435), .ZN(n13453) );
  AND2_X1 U13380 ( .A1(n13433), .A2(n13454), .ZN(n13452) );
  OR2_X1 U13381 ( .A1(n13435), .A2(n13436), .ZN(n13454) );
  OR2_X1 U13382 ( .A1(n8049), .A2(n8025), .ZN(n13436) );
  OR2_X1 U13383 ( .A1(n13455), .A2(n13456), .ZN(n13435) );
  AND2_X1 U13384 ( .A1(n13432), .A2(n13431), .ZN(n13456) );
  AND2_X1 U13385 ( .A1(n13429), .A2(n13457), .ZN(n13455) );
  OR2_X1 U13386 ( .A1(n13431), .A2(n13432), .ZN(n13457) );
  OR2_X1 U13387 ( .A1(n8030), .A2(n8049), .ZN(n13432) );
  OR2_X1 U13388 ( .A1(n13458), .A2(n13459), .ZN(n13431) );
  AND2_X1 U13389 ( .A1(n13428), .A2(n13427), .ZN(n13459) );
  AND2_X1 U13390 ( .A1(n13425), .A2(n13460), .ZN(n13458) );
  OR2_X1 U13391 ( .A1(n13427), .A2(n13428), .ZN(n13460) );
  OR2_X1 U13392 ( .A1(n8049), .A2(n8034), .ZN(n13428) );
  OR2_X1 U13393 ( .A1(n13461), .A2(n13462), .ZN(n13427) );
  AND2_X1 U13394 ( .A1(n13424), .A2(n13423), .ZN(n13462) );
  AND2_X1 U13395 ( .A1(n13421), .A2(n13463), .ZN(n13461) );
  OR2_X1 U13396 ( .A1(n13423), .A2(n13424), .ZN(n13463) );
  OR2_X1 U13397 ( .A1(n8039), .A2(n8049), .ZN(n13424) );
  OR2_X1 U13398 ( .A1(n13464), .A2(n13465), .ZN(n13423) );
  AND2_X1 U13399 ( .A1(n13420), .A2(n13419), .ZN(n13465) );
  AND2_X1 U13400 ( .A1(n13417), .A2(n13466), .ZN(n13464) );
  OR2_X1 U13401 ( .A1(n13419), .A2(n13420), .ZN(n13466) );
  OR2_X1 U13402 ( .A1(n8049), .A2(n8043), .ZN(n13420) );
  OR2_X1 U13403 ( .A1(n13467), .A2(n13468), .ZN(n13419) );
  AND2_X1 U13404 ( .A1(n8050), .A2(n13416), .ZN(n13468) );
  AND2_X1 U13405 ( .A1(n13414), .A2(n13469), .ZN(n13467) );
  OR2_X1 U13406 ( .A1(n13416), .A2(n8050), .ZN(n13469) );
  OR2_X1 U13407 ( .A1(n8048), .A2(n8049), .ZN(n8050) );
  OR2_X1 U13408 ( .A1(n13470), .A2(n13471), .ZN(n13416) );
  AND2_X1 U13409 ( .A1(n13413), .A2(n13412), .ZN(n13471) );
  AND2_X1 U13410 ( .A1(n13410), .A2(n13472), .ZN(n13470) );
  OR2_X1 U13411 ( .A1(n13412), .A2(n13413), .ZN(n13472) );
  OR2_X1 U13412 ( .A1(n8052), .A2(n8049), .ZN(n13413) );
  OR2_X1 U13413 ( .A1(n13473), .A2(n13474), .ZN(n13412) );
  AND2_X1 U13414 ( .A1(n13409), .A2(n13408), .ZN(n13474) );
  AND2_X1 U13415 ( .A1(n13406), .A2(n13475), .ZN(n13473) );
  OR2_X1 U13416 ( .A1(n13408), .A2(n13409), .ZN(n13475) );
  OR2_X1 U13417 ( .A1(n8057), .A2(n8049), .ZN(n13409) );
  OR2_X1 U13418 ( .A1(n13476), .A2(n13477), .ZN(n13408) );
  AND2_X1 U13419 ( .A1(n13405), .A2(n13404), .ZN(n13477) );
  AND2_X1 U13420 ( .A1(n13402), .A2(n13478), .ZN(n13476) );
  OR2_X1 U13421 ( .A1(n13404), .A2(n13405), .ZN(n13478) );
  OR2_X1 U13422 ( .A1(n8061), .A2(n8049), .ZN(n13405) );
  OR2_X1 U13423 ( .A1(n13479), .A2(n13480), .ZN(n13404) );
  AND2_X1 U13424 ( .A1(n13401), .A2(n13400), .ZN(n13480) );
  AND2_X1 U13425 ( .A1(n13398), .A2(n13481), .ZN(n13479) );
  OR2_X1 U13426 ( .A1(n13400), .A2(n13401), .ZN(n13481) );
  OR2_X1 U13427 ( .A1(n8066), .A2(n8049), .ZN(n13401) );
  OR2_X1 U13428 ( .A1(n13482), .A2(n13483), .ZN(n13400) );
  AND2_X1 U13429 ( .A1(n13397), .A2(n13396), .ZN(n13483) );
  AND2_X1 U13430 ( .A1(n13394), .A2(n13484), .ZN(n13482) );
  OR2_X1 U13431 ( .A1(n13396), .A2(n13397), .ZN(n13484) );
  OR2_X1 U13432 ( .A1(n8070), .A2(n8049), .ZN(n13397) );
  OR2_X1 U13433 ( .A1(n13485), .A2(n13486), .ZN(n13396) );
  AND2_X1 U13434 ( .A1(n13393), .A2(n13392), .ZN(n13486) );
  AND2_X1 U13435 ( .A1(n13390), .A2(n13487), .ZN(n13485) );
  OR2_X1 U13436 ( .A1(n13392), .A2(n13393), .ZN(n13487) );
  OR2_X1 U13437 ( .A1(n8075), .A2(n8049), .ZN(n13393) );
  OR2_X1 U13438 ( .A1(n13488), .A2(n13489), .ZN(n13392) );
  AND2_X1 U13439 ( .A1(n13389), .A2(n13388), .ZN(n13489) );
  AND2_X1 U13440 ( .A1(n13386), .A2(n13490), .ZN(n13488) );
  OR2_X1 U13441 ( .A1(n13388), .A2(n13389), .ZN(n13490) );
  OR2_X1 U13442 ( .A1(n8079), .A2(n8049), .ZN(n13389) );
  OR2_X1 U13443 ( .A1(n13491), .A2(n13492), .ZN(n13388) );
  AND2_X1 U13444 ( .A1(n13385), .A2(n13384), .ZN(n13492) );
  AND2_X1 U13445 ( .A1(n13382), .A2(n13493), .ZN(n13491) );
  OR2_X1 U13446 ( .A1(n13384), .A2(n13385), .ZN(n13493) );
  OR2_X1 U13447 ( .A1(n8084), .A2(n8049), .ZN(n13385) );
  OR2_X1 U13448 ( .A1(n13494), .A2(n13495), .ZN(n13384) );
  AND2_X1 U13449 ( .A1(n13381), .A2(n13380), .ZN(n13495) );
  AND2_X1 U13450 ( .A1(n13378), .A2(n13496), .ZN(n13494) );
  OR2_X1 U13451 ( .A1(n13380), .A2(n13381), .ZN(n13496) );
  OR2_X1 U13452 ( .A1(n8088), .A2(n8049), .ZN(n13381) );
  OR2_X1 U13453 ( .A1(n13497), .A2(n13498), .ZN(n13380) );
  AND2_X1 U13454 ( .A1(n13377), .A2(n13376), .ZN(n13498) );
  AND2_X1 U13455 ( .A1(n13374), .A2(n13499), .ZN(n13497) );
  OR2_X1 U13456 ( .A1(n13376), .A2(n13377), .ZN(n13499) );
  OR2_X1 U13457 ( .A1(n8093), .A2(n8049), .ZN(n13377) );
  OR2_X1 U13458 ( .A1(n13500), .A2(n13501), .ZN(n13376) );
  AND2_X1 U13459 ( .A1(n13370), .A2(n13373), .ZN(n13501) );
  AND2_X1 U13460 ( .A1(n13502), .A2(n13372), .ZN(n13500) );
  OR2_X1 U13461 ( .A1(n13503), .A2(n13504), .ZN(n13372) );
  AND2_X1 U13462 ( .A1(n13369), .A2(n13368), .ZN(n13504) );
  AND2_X1 U13463 ( .A1(n13366), .A2(n13505), .ZN(n13503) );
  OR2_X1 U13464 ( .A1(n13368), .A2(n13369), .ZN(n13505) );
  OR2_X1 U13465 ( .A1(n8102), .A2(n8049), .ZN(n13369) );
  OR2_X1 U13466 ( .A1(n13506), .A2(n13507), .ZN(n13368) );
  AND2_X1 U13467 ( .A1(n13362), .A2(n13365), .ZN(n13507) );
  AND2_X1 U13468 ( .A1(n13508), .A2(n13364), .ZN(n13506) );
  OR2_X1 U13469 ( .A1(n13509), .A2(n13510), .ZN(n13364) );
  AND2_X1 U13470 ( .A1(n13358), .A2(n13361), .ZN(n13510) );
  AND2_X1 U13471 ( .A1(n13511), .A2(n13360), .ZN(n13509) );
  OR2_X1 U13472 ( .A1(n13512), .A2(n13513), .ZN(n13360) );
  AND2_X1 U13473 ( .A1(n13354), .A2(n13357), .ZN(n13513) );
  AND2_X1 U13474 ( .A1(n13514), .A2(n13356), .ZN(n13512) );
  OR2_X1 U13475 ( .A1(n13515), .A2(n13516), .ZN(n13356) );
  AND2_X1 U13476 ( .A1(n13350), .A2(n13353), .ZN(n13516) );
  AND2_X1 U13477 ( .A1(n13517), .A2(n13352), .ZN(n13515) );
  OR2_X1 U13478 ( .A1(n13518), .A2(n13519), .ZN(n13352) );
  AND2_X1 U13479 ( .A1(n13346), .A2(n13349), .ZN(n13519) );
  AND2_X1 U13480 ( .A1(n13520), .A2(n13348), .ZN(n13518) );
  OR2_X1 U13481 ( .A1(n13521), .A2(n13522), .ZN(n13348) );
  AND2_X1 U13482 ( .A1(n13342), .A2(n13345), .ZN(n13522) );
  AND2_X1 U13483 ( .A1(n13523), .A2(n13344), .ZN(n13521) );
  OR2_X1 U13484 ( .A1(n13524), .A2(n13525), .ZN(n13344) );
  AND2_X1 U13485 ( .A1(n13338), .A2(n13341), .ZN(n13525) );
  AND2_X1 U13486 ( .A1(n13526), .A2(n13340), .ZN(n13524) );
  OR2_X1 U13487 ( .A1(n13527), .A2(n13528), .ZN(n13340) );
  AND2_X1 U13488 ( .A1(n13334), .A2(n13337), .ZN(n13528) );
  AND2_X1 U13489 ( .A1(n13529), .A2(n13530), .ZN(n13527) );
  OR2_X1 U13490 ( .A1(n13337), .A2(n13334), .ZN(n13530) );
  OR2_X1 U13491 ( .A1(n8127), .A2(n8049), .ZN(n13334) );
  OR3_X1 U13492 ( .A1(n8044), .A2(n8981), .A3(n8049), .ZN(n13337) );
  INV_X1 U13493 ( .A(n13336), .ZN(n13529) );
  OR2_X1 U13494 ( .A1(n13531), .A2(n13532), .ZN(n13336) );
  AND2_X1 U13495 ( .A1(b_8_), .A2(n13533), .ZN(n13532) );
  OR2_X1 U13496 ( .A1(n13534), .A2(n7598), .ZN(n13533) );
  AND2_X1 U13497 ( .A1(a_30_), .A2(n8040), .ZN(n13534) );
  AND2_X1 U13498 ( .A1(b_7_), .A2(n13535), .ZN(n13531) );
  OR2_X1 U13499 ( .A1(n13536), .A2(n7601), .ZN(n13535) );
  AND2_X1 U13500 ( .A1(a_31_), .A2(n8044), .ZN(n13536) );
  OR2_X1 U13501 ( .A1(n13341), .A2(n13338), .ZN(n13526) );
  XNOR2_X1 U13502 ( .A(n13537), .B(n13538), .ZN(n13338) );
  XOR2_X1 U13503 ( .A(n13539), .B(n13540), .Z(n13538) );
  OR2_X1 U13504 ( .A1(n8124), .A2(n8049), .ZN(n13341) );
  OR2_X1 U13505 ( .A1(n13345), .A2(n13342), .ZN(n13523) );
  XOR2_X1 U13506 ( .A(n13541), .B(n13542), .Z(n13342) );
  XOR2_X1 U13507 ( .A(n13543), .B(n13544), .Z(n13542) );
  OR2_X1 U13508 ( .A1(n8121), .A2(n8049), .ZN(n13345) );
  OR2_X1 U13509 ( .A1(n13349), .A2(n13346), .ZN(n13520) );
  XOR2_X1 U13510 ( .A(n13545), .B(n13546), .Z(n13346) );
  XOR2_X1 U13511 ( .A(n13547), .B(n13548), .Z(n13546) );
  OR2_X1 U13512 ( .A1(n8118), .A2(n8049), .ZN(n13349) );
  OR2_X1 U13513 ( .A1(n13353), .A2(n13350), .ZN(n13517) );
  XOR2_X1 U13514 ( .A(n13549), .B(n13550), .Z(n13350) );
  XOR2_X1 U13515 ( .A(n13551), .B(n13552), .Z(n13550) );
  OR2_X1 U13516 ( .A1(n8115), .A2(n8049), .ZN(n13353) );
  OR2_X1 U13517 ( .A1(n13357), .A2(n13354), .ZN(n13514) );
  XOR2_X1 U13518 ( .A(n13553), .B(n13554), .Z(n13354) );
  XOR2_X1 U13519 ( .A(n13555), .B(n13556), .Z(n13554) );
  OR2_X1 U13520 ( .A1(n8112), .A2(n8049), .ZN(n13357) );
  OR2_X1 U13521 ( .A1(n13361), .A2(n13358), .ZN(n13511) );
  XOR2_X1 U13522 ( .A(n13557), .B(n13558), .Z(n13358) );
  XOR2_X1 U13523 ( .A(n13559), .B(n13560), .Z(n13558) );
  OR2_X1 U13524 ( .A1(n8109), .A2(n8049), .ZN(n13361) );
  OR2_X1 U13525 ( .A1(n13365), .A2(n13362), .ZN(n13508) );
  XOR2_X1 U13526 ( .A(n13561), .B(n13562), .Z(n13362) );
  XOR2_X1 U13527 ( .A(n13563), .B(n13564), .Z(n13562) );
  OR2_X1 U13528 ( .A1(n8106), .A2(n8049), .ZN(n13365) );
  XOR2_X1 U13529 ( .A(n13565), .B(n13566), .Z(n13366) );
  XOR2_X1 U13530 ( .A(n13567), .B(n13568), .Z(n13566) );
  OR2_X1 U13531 ( .A1(n13373), .A2(n13370), .ZN(n13502) );
  XOR2_X1 U13532 ( .A(n13569), .B(n13570), .Z(n13370) );
  XOR2_X1 U13533 ( .A(n13571), .B(n13572), .Z(n13570) );
  OR2_X1 U13534 ( .A1(n8097), .A2(n8049), .ZN(n13373) );
  XOR2_X1 U13535 ( .A(n13573), .B(n13574), .Z(n13374) );
  XOR2_X1 U13536 ( .A(n13575), .B(n13576), .Z(n13574) );
  XOR2_X1 U13537 ( .A(n13577), .B(n13578), .Z(n13378) );
  XOR2_X1 U13538 ( .A(n13579), .B(n13580), .Z(n13578) );
  XOR2_X1 U13539 ( .A(n13581), .B(n13582), .Z(n13382) );
  XOR2_X1 U13540 ( .A(n13583), .B(n13584), .Z(n13582) );
  XOR2_X1 U13541 ( .A(n13585), .B(n13586), .Z(n13386) );
  XOR2_X1 U13542 ( .A(n13587), .B(n13588), .Z(n13586) );
  XOR2_X1 U13543 ( .A(n13589), .B(n13590), .Z(n13390) );
  XOR2_X1 U13544 ( .A(n13591), .B(n13592), .Z(n13590) );
  XOR2_X1 U13545 ( .A(n13593), .B(n13594), .Z(n13394) );
  XOR2_X1 U13546 ( .A(n13595), .B(n13596), .Z(n13594) );
  XOR2_X1 U13547 ( .A(n13597), .B(n13598), .Z(n13398) );
  XOR2_X1 U13548 ( .A(n13599), .B(n13600), .Z(n13598) );
  XOR2_X1 U13549 ( .A(n13601), .B(n13602), .Z(n13402) );
  XOR2_X1 U13550 ( .A(n13603), .B(n13604), .Z(n13602) );
  XOR2_X1 U13551 ( .A(n13605), .B(n13606), .Z(n13406) );
  XOR2_X1 U13552 ( .A(n13607), .B(n13608), .Z(n13606) );
  XOR2_X1 U13553 ( .A(n13609), .B(n13610), .Z(n13410) );
  XOR2_X1 U13554 ( .A(n13611), .B(n13612), .Z(n13610) );
  XOR2_X1 U13555 ( .A(n13613), .B(n13614), .Z(n13414) );
  XOR2_X1 U13556 ( .A(n13615), .B(n13616), .Z(n13614) );
  XOR2_X1 U13557 ( .A(n13617), .B(n13618), .Z(n13417) );
  XOR2_X1 U13558 ( .A(n13619), .B(n13620), .Z(n13618) );
  XNOR2_X1 U13559 ( .A(n13621), .B(n13622), .ZN(n13421) );
  XOR2_X1 U13560 ( .A(n7905), .B(n13623), .Z(n13621) );
  INV_X1 U13561 ( .A(n8045), .ZN(n7905) );
  XOR2_X1 U13562 ( .A(n13624), .B(n13625), .Z(n13425) );
  XOR2_X1 U13563 ( .A(n13626), .B(n13627), .Z(n13625) );
  XOR2_X1 U13564 ( .A(n13628), .B(n13629), .Z(n13429) );
  XOR2_X1 U13565 ( .A(n13630), .B(n13631), .Z(n13629) );
  XOR2_X1 U13566 ( .A(n13632), .B(n13633), .Z(n13433) );
  XOR2_X1 U13567 ( .A(n13634), .B(n13635), .Z(n13633) );
  XOR2_X1 U13568 ( .A(n13636), .B(n13637), .Z(n13437) );
  XOR2_X1 U13569 ( .A(n13638), .B(n13639), .Z(n13637) );
  XOR2_X1 U13570 ( .A(n13640), .B(n13641), .Z(n13441) );
  XOR2_X1 U13571 ( .A(n13642), .B(n13643), .Z(n13641) );
  XOR2_X1 U13572 ( .A(n8540), .B(n13644), .Z(n8533) );
  XOR2_X1 U13573 ( .A(n8539), .B(n8538), .Z(n13644) );
  OR2_X1 U13574 ( .A1(n8044), .A2(n8016), .ZN(n8538) );
  OR2_X1 U13575 ( .A1(n13645), .A2(n13646), .ZN(n8539) );
  AND2_X1 U13576 ( .A1(n13643), .A2(n13642), .ZN(n13646) );
  AND2_X1 U13577 ( .A1(n13640), .A2(n13647), .ZN(n13645) );
  OR2_X1 U13578 ( .A1(n13642), .A2(n13643), .ZN(n13647) );
  OR2_X1 U13579 ( .A1(n8021), .A2(n8044), .ZN(n13643) );
  OR2_X1 U13580 ( .A1(n13648), .A2(n13649), .ZN(n13642) );
  AND2_X1 U13581 ( .A1(n13639), .A2(n13638), .ZN(n13649) );
  AND2_X1 U13582 ( .A1(n13636), .A2(n13650), .ZN(n13648) );
  OR2_X1 U13583 ( .A1(n13638), .A2(n13639), .ZN(n13650) );
  OR2_X1 U13584 ( .A1(n8044), .A2(n8025), .ZN(n13639) );
  OR2_X1 U13585 ( .A1(n13651), .A2(n13652), .ZN(n13638) );
  AND2_X1 U13586 ( .A1(n13635), .A2(n13634), .ZN(n13652) );
  AND2_X1 U13587 ( .A1(n13632), .A2(n13653), .ZN(n13651) );
  OR2_X1 U13588 ( .A1(n13634), .A2(n13635), .ZN(n13653) );
  OR2_X1 U13589 ( .A1(n8030), .A2(n8044), .ZN(n13635) );
  OR2_X1 U13590 ( .A1(n13654), .A2(n13655), .ZN(n13634) );
  AND2_X1 U13591 ( .A1(n13631), .A2(n13630), .ZN(n13655) );
  AND2_X1 U13592 ( .A1(n13628), .A2(n13656), .ZN(n13654) );
  OR2_X1 U13593 ( .A1(n13630), .A2(n13631), .ZN(n13656) );
  OR2_X1 U13594 ( .A1(n8044), .A2(n8034), .ZN(n13631) );
  OR2_X1 U13595 ( .A1(n13657), .A2(n13658), .ZN(n13630) );
  AND2_X1 U13596 ( .A1(n13627), .A2(n13626), .ZN(n13658) );
  AND2_X1 U13597 ( .A1(n13624), .A2(n13659), .ZN(n13657) );
  OR2_X1 U13598 ( .A1(n13626), .A2(n13627), .ZN(n13659) );
  OR2_X1 U13599 ( .A1(n8039), .A2(n8044), .ZN(n13627) );
  OR2_X1 U13600 ( .A1(n13660), .A2(n13661), .ZN(n13626) );
  AND2_X1 U13601 ( .A1(n13623), .A2(n8045), .ZN(n13661) );
  AND2_X1 U13602 ( .A1(n13622), .A2(n13662), .ZN(n13660) );
  OR2_X1 U13603 ( .A1(n8045), .A2(n13623), .ZN(n13662) );
  OR2_X1 U13604 ( .A1(n13663), .A2(n13664), .ZN(n13623) );
  AND2_X1 U13605 ( .A1(n13620), .A2(n13619), .ZN(n13664) );
  AND2_X1 U13606 ( .A1(n13617), .A2(n13665), .ZN(n13663) );
  OR2_X1 U13607 ( .A1(n13619), .A2(n13620), .ZN(n13665) );
  OR2_X1 U13608 ( .A1(n8044), .A2(n8048), .ZN(n13620) );
  OR2_X1 U13609 ( .A1(n13666), .A2(n13667), .ZN(n13619) );
  AND2_X1 U13610 ( .A1(n13616), .A2(n13615), .ZN(n13667) );
  AND2_X1 U13611 ( .A1(n13613), .A2(n13668), .ZN(n13666) );
  OR2_X1 U13612 ( .A1(n13615), .A2(n13616), .ZN(n13668) );
  OR2_X1 U13613 ( .A1(n8044), .A2(n8052), .ZN(n13616) );
  OR2_X1 U13614 ( .A1(n13669), .A2(n13670), .ZN(n13615) );
  AND2_X1 U13615 ( .A1(n13612), .A2(n13611), .ZN(n13670) );
  AND2_X1 U13616 ( .A1(n13609), .A2(n13671), .ZN(n13669) );
  OR2_X1 U13617 ( .A1(n13611), .A2(n13612), .ZN(n13671) );
  OR2_X1 U13618 ( .A1(n8044), .A2(n8057), .ZN(n13612) );
  OR2_X1 U13619 ( .A1(n13672), .A2(n13673), .ZN(n13611) );
  AND2_X1 U13620 ( .A1(n13608), .A2(n13607), .ZN(n13673) );
  AND2_X1 U13621 ( .A1(n13605), .A2(n13674), .ZN(n13672) );
  OR2_X1 U13622 ( .A1(n13607), .A2(n13608), .ZN(n13674) );
  OR2_X1 U13623 ( .A1(n8044), .A2(n8061), .ZN(n13608) );
  OR2_X1 U13624 ( .A1(n13675), .A2(n13676), .ZN(n13607) );
  AND2_X1 U13625 ( .A1(n13604), .A2(n13603), .ZN(n13676) );
  AND2_X1 U13626 ( .A1(n13601), .A2(n13677), .ZN(n13675) );
  OR2_X1 U13627 ( .A1(n13603), .A2(n13604), .ZN(n13677) );
  OR2_X1 U13628 ( .A1(n8044), .A2(n8066), .ZN(n13604) );
  OR2_X1 U13629 ( .A1(n13678), .A2(n13679), .ZN(n13603) );
  AND2_X1 U13630 ( .A1(n13600), .A2(n13599), .ZN(n13679) );
  AND2_X1 U13631 ( .A1(n13597), .A2(n13680), .ZN(n13678) );
  OR2_X1 U13632 ( .A1(n13599), .A2(n13600), .ZN(n13680) );
  OR2_X1 U13633 ( .A1(n8044), .A2(n8070), .ZN(n13600) );
  OR2_X1 U13634 ( .A1(n13681), .A2(n13682), .ZN(n13599) );
  AND2_X1 U13635 ( .A1(n13596), .A2(n13595), .ZN(n13682) );
  AND2_X1 U13636 ( .A1(n13593), .A2(n13683), .ZN(n13681) );
  OR2_X1 U13637 ( .A1(n13595), .A2(n13596), .ZN(n13683) );
  OR2_X1 U13638 ( .A1(n8044), .A2(n8075), .ZN(n13596) );
  OR2_X1 U13639 ( .A1(n13684), .A2(n13685), .ZN(n13595) );
  AND2_X1 U13640 ( .A1(n13592), .A2(n13591), .ZN(n13685) );
  AND2_X1 U13641 ( .A1(n13589), .A2(n13686), .ZN(n13684) );
  OR2_X1 U13642 ( .A1(n13591), .A2(n13592), .ZN(n13686) );
  OR2_X1 U13643 ( .A1(n8044), .A2(n8079), .ZN(n13592) );
  OR2_X1 U13644 ( .A1(n13687), .A2(n13688), .ZN(n13591) );
  AND2_X1 U13645 ( .A1(n13588), .A2(n13587), .ZN(n13688) );
  AND2_X1 U13646 ( .A1(n13585), .A2(n13689), .ZN(n13687) );
  OR2_X1 U13647 ( .A1(n13587), .A2(n13588), .ZN(n13689) );
  OR2_X1 U13648 ( .A1(n8044), .A2(n8084), .ZN(n13588) );
  OR2_X1 U13649 ( .A1(n13690), .A2(n13691), .ZN(n13587) );
  AND2_X1 U13650 ( .A1(n13584), .A2(n13583), .ZN(n13691) );
  AND2_X1 U13651 ( .A1(n13581), .A2(n13692), .ZN(n13690) );
  OR2_X1 U13652 ( .A1(n13583), .A2(n13584), .ZN(n13692) );
  OR2_X1 U13653 ( .A1(n8044), .A2(n8088), .ZN(n13584) );
  OR2_X1 U13654 ( .A1(n13693), .A2(n13694), .ZN(n13583) );
  AND2_X1 U13655 ( .A1(n13580), .A2(n13579), .ZN(n13694) );
  AND2_X1 U13656 ( .A1(n13577), .A2(n13695), .ZN(n13693) );
  OR2_X1 U13657 ( .A1(n13579), .A2(n13580), .ZN(n13695) );
  OR2_X1 U13658 ( .A1(n8044), .A2(n8093), .ZN(n13580) );
  OR2_X1 U13659 ( .A1(n13696), .A2(n13697), .ZN(n13579) );
  AND2_X1 U13660 ( .A1(n13576), .A2(n13575), .ZN(n13697) );
  AND2_X1 U13661 ( .A1(n13573), .A2(n13698), .ZN(n13696) );
  OR2_X1 U13662 ( .A1(n13575), .A2(n13576), .ZN(n13698) );
  OR2_X1 U13663 ( .A1(n8044), .A2(n8097), .ZN(n13576) );
  OR2_X1 U13664 ( .A1(n13699), .A2(n13700), .ZN(n13575) );
  AND2_X1 U13665 ( .A1(n13569), .A2(n13572), .ZN(n13700) );
  AND2_X1 U13666 ( .A1(n13701), .A2(n13571), .ZN(n13699) );
  OR2_X1 U13667 ( .A1(n13702), .A2(n13703), .ZN(n13571) );
  AND2_X1 U13668 ( .A1(n13568), .A2(n13567), .ZN(n13703) );
  AND2_X1 U13669 ( .A1(n13565), .A2(n13704), .ZN(n13702) );
  OR2_X1 U13670 ( .A1(n13567), .A2(n13568), .ZN(n13704) );
  OR2_X1 U13671 ( .A1(n8044), .A2(n8106), .ZN(n13568) );
  OR2_X1 U13672 ( .A1(n13705), .A2(n13706), .ZN(n13567) );
  AND2_X1 U13673 ( .A1(n13561), .A2(n13564), .ZN(n13706) );
  AND2_X1 U13674 ( .A1(n13707), .A2(n13563), .ZN(n13705) );
  OR2_X1 U13675 ( .A1(n13708), .A2(n13709), .ZN(n13563) );
  AND2_X1 U13676 ( .A1(n13557), .A2(n13560), .ZN(n13709) );
  AND2_X1 U13677 ( .A1(n13710), .A2(n13559), .ZN(n13708) );
  OR2_X1 U13678 ( .A1(n13711), .A2(n13712), .ZN(n13559) );
  AND2_X1 U13679 ( .A1(n13553), .A2(n13556), .ZN(n13712) );
  AND2_X1 U13680 ( .A1(n13713), .A2(n13555), .ZN(n13711) );
  OR2_X1 U13681 ( .A1(n13714), .A2(n13715), .ZN(n13555) );
  AND2_X1 U13682 ( .A1(n13549), .A2(n13552), .ZN(n13715) );
  AND2_X1 U13683 ( .A1(n13716), .A2(n13551), .ZN(n13714) );
  OR2_X1 U13684 ( .A1(n13717), .A2(n13718), .ZN(n13551) );
  AND2_X1 U13685 ( .A1(n13545), .A2(n13548), .ZN(n13718) );
  AND2_X1 U13686 ( .A1(n13719), .A2(n13547), .ZN(n13717) );
  OR2_X1 U13687 ( .A1(n13720), .A2(n13721), .ZN(n13547) );
  AND2_X1 U13688 ( .A1(n13541), .A2(n13544), .ZN(n13721) );
  AND2_X1 U13689 ( .A1(n13722), .A2(n13543), .ZN(n13720) );
  OR2_X1 U13690 ( .A1(n13723), .A2(n13724), .ZN(n13543) );
  AND2_X1 U13691 ( .A1(n13537), .A2(n13540), .ZN(n13724) );
  AND2_X1 U13692 ( .A1(n13725), .A2(n13726), .ZN(n13723) );
  OR2_X1 U13693 ( .A1(n13540), .A2(n13537), .ZN(n13726) );
  OR2_X1 U13694 ( .A1(n8044), .A2(n8127), .ZN(n13537) );
  OR3_X1 U13695 ( .A1(n8040), .A2(n8044), .A3(n8981), .ZN(n13540) );
  INV_X1 U13696 ( .A(n13539), .ZN(n13725) );
  OR2_X1 U13697 ( .A1(n13727), .A2(n13728), .ZN(n13539) );
  AND2_X1 U13698 ( .A1(b_7_), .A2(n13729), .ZN(n13728) );
  OR2_X1 U13699 ( .A1(n13730), .A2(n7598), .ZN(n13729) );
  AND2_X1 U13700 ( .A1(a_30_), .A2(n8035), .ZN(n13730) );
  AND2_X1 U13701 ( .A1(b_6_), .A2(n13731), .ZN(n13727) );
  OR2_X1 U13702 ( .A1(n13732), .A2(n7601), .ZN(n13731) );
  AND2_X1 U13703 ( .A1(a_31_), .A2(n8040), .ZN(n13732) );
  OR2_X1 U13704 ( .A1(n13544), .A2(n13541), .ZN(n13722) );
  XNOR2_X1 U13705 ( .A(n13733), .B(n13734), .ZN(n13541) );
  XOR2_X1 U13706 ( .A(n13735), .B(n13736), .Z(n13734) );
  OR2_X1 U13707 ( .A1(n8044), .A2(n8124), .ZN(n13544) );
  OR2_X1 U13708 ( .A1(n13548), .A2(n13545), .ZN(n13719) );
  XOR2_X1 U13709 ( .A(n13737), .B(n13738), .Z(n13545) );
  XOR2_X1 U13710 ( .A(n13739), .B(n13740), .Z(n13738) );
  OR2_X1 U13711 ( .A1(n8044), .A2(n8121), .ZN(n13548) );
  OR2_X1 U13712 ( .A1(n13552), .A2(n13549), .ZN(n13716) );
  XOR2_X1 U13713 ( .A(n13741), .B(n13742), .Z(n13549) );
  XOR2_X1 U13714 ( .A(n13743), .B(n13744), .Z(n13742) );
  OR2_X1 U13715 ( .A1(n8044), .A2(n8118), .ZN(n13552) );
  OR2_X1 U13716 ( .A1(n13556), .A2(n13553), .ZN(n13713) );
  XOR2_X1 U13717 ( .A(n13745), .B(n13746), .Z(n13553) );
  XOR2_X1 U13718 ( .A(n13747), .B(n13748), .Z(n13746) );
  OR2_X1 U13719 ( .A1(n8044), .A2(n8115), .ZN(n13556) );
  OR2_X1 U13720 ( .A1(n13560), .A2(n13557), .ZN(n13710) );
  XOR2_X1 U13721 ( .A(n13749), .B(n13750), .Z(n13557) );
  XOR2_X1 U13722 ( .A(n13751), .B(n13752), .Z(n13750) );
  OR2_X1 U13723 ( .A1(n8044), .A2(n8112), .ZN(n13560) );
  OR2_X1 U13724 ( .A1(n13564), .A2(n13561), .ZN(n13707) );
  XOR2_X1 U13725 ( .A(n13753), .B(n13754), .Z(n13561) );
  XOR2_X1 U13726 ( .A(n13755), .B(n13756), .Z(n13754) );
  OR2_X1 U13727 ( .A1(n8044), .A2(n8109), .ZN(n13564) );
  XOR2_X1 U13728 ( .A(n13757), .B(n13758), .Z(n13565) );
  XOR2_X1 U13729 ( .A(n13759), .B(n13760), .Z(n13758) );
  OR2_X1 U13730 ( .A1(n13572), .A2(n13569), .ZN(n13701) );
  XOR2_X1 U13731 ( .A(n13761), .B(n13762), .Z(n13569) );
  XOR2_X1 U13732 ( .A(n13763), .B(n13764), .Z(n13762) );
  OR2_X1 U13733 ( .A1(n8044), .A2(n8102), .ZN(n13572) );
  XOR2_X1 U13734 ( .A(n13765), .B(n13766), .Z(n13573) );
  XOR2_X1 U13735 ( .A(n13767), .B(n13768), .Z(n13766) );
  XOR2_X1 U13736 ( .A(n13769), .B(n13770), .Z(n13577) );
  XOR2_X1 U13737 ( .A(n13771), .B(n13772), .Z(n13770) );
  XOR2_X1 U13738 ( .A(n13773), .B(n13774), .Z(n13581) );
  XOR2_X1 U13739 ( .A(n13775), .B(n13776), .Z(n13774) );
  XOR2_X1 U13740 ( .A(n13777), .B(n13778), .Z(n13585) );
  XOR2_X1 U13741 ( .A(n13779), .B(n13780), .Z(n13778) );
  XOR2_X1 U13742 ( .A(n13781), .B(n13782), .Z(n13589) );
  XOR2_X1 U13743 ( .A(n13783), .B(n13784), .Z(n13782) );
  XOR2_X1 U13744 ( .A(n13785), .B(n13786), .Z(n13593) );
  XOR2_X1 U13745 ( .A(n13787), .B(n13788), .Z(n13786) );
  XOR2_X1 U13746 ( .A(n13789), .B(n13790), .Z(n13597) );
  XOR2_X1 U13747 ( .A(n13791), .B(n13792), .Z(n13790) );
  XOR2_X1 U13748 ( .A(n13793), .B(n13794), .Z(n13601) );
  XOR2_X1 U13749 ( .A(n13795), .B(n13796), .Z(n13794) );
  XOR2_X1 U13750 ( .A(n13797), .B(n13798), .Z(n13605) );
  XOR2_X1 U13751 ( .A(n13799), .B(n13800), .Z(n13798) );
  XOR2_X1 U13752 ( .A(n13801), .B(n13802), .Z(n13609) );
  XOR2_X1 U13753 ( .A(n13803), .B(n13804), .Z(n13802) );
  XOR2_X1 U13754 ( .A(n13805), .B(n13806), .Z(n13613) );
  XOR2_X1 U13755 ( .A(n13807), .B(n13808), .Z(n13806) );
  XOR2_X1 U13756 ( .A(n13809), .B(n13810), .Z(n13617) );
  XOR2_X1 U13757 ( .A(n13811), .B(n13812), .Z(n13810) );
  OR2_X1 U13758 ( .A1(n8044), .A2(n8043), .ZN(n8045) );
  INV_X1 U13759 ( .A(b_8_), .ZN(n8044) );
  XOR2_X1 U13760 ( .A(n13813), .B(n13814), .Z(n13622) );
  XOR2_X1 U13761 ( .A(n13815), .B(n13816), .Z(n13814) );
  XOR2_X1 U13762 ( .A(n13817), .B(n13818), .Z(n13624) );
  XOR2_X1 U13763 ( .A(n13819), .B(n13820), .Z(n13818) );
  XOR2_X1 U13764 ( .A(n13821), .B(n13822), .Z(n13628) );
  XOR2_X1 U13765 ( .A(n13823), .B(n8041), .Z(n13822) );
  XOR2_X1 U13766 ( .A(n13824), .B(n13825), .Z(n13632) );
  XOR2_X1 U13767 ( .A(n13826), .B(n13827), .Z(n13825) );
  XOR2_X1 U13768 ( .A(n13828), .B(n13829), .Z(n13636) );
  XOR2_X1 U13769 ( .A(n13830), .B(n13831), .Z(n13829) );
  XOR2_X1 U13770 ( .A(n13832), .B(n13833), .Z(n13640) );
  XOR2_X1 U13771 ( .A(n13834), .B(n13835), .Z(n13833) );
  XOR2_X1 U13772 ( .A(n8547), .B(n13836), .Z(n8540) );
  XOR2_X1 U13773 ( .A(n8546), .B(n8545), .Z(n13836) );
  OR2_X1 U13774 ( .A1(n8021), .A2(n8040), .ZN(n8545) );
  OR2_X1 U13775 ( .A1(n13837), .A2(n13838), .ZN(n8546) );
  AND2_X1 U13776 ( .A1(n13835), .A2(n13834), .ZN(n13838) );
  AND2_X1 U13777 ( .A1(n13832), .A2(n13839), .ZN(n13837) );
  OR2_X1 U13778 ( .A1(n13834), .A2(n13835), .ZN(n13839) );
  OR2_X1 U13779 ( .A1(n8040), .A2(n8025), .ZN(n13835) );
  OR2_X1 U13780 ( .A1(n13840), .A2(n13841), .ZN(n13834) );
  AND2_X1 U13781 ( .A1(n13831), .A2(n13830), .ZN(n13841) );
  AND2_X1 U13782 ( .A1(n13828), .A2(n13842), .ZN(n13840) );
  OR2_X1 U13783 ( .A1(n13830), .A2(n13831), .ZN(n13842) );
  OR2_X1 U13784 ( .A1(n8030), .A2(n8040), .ZN(n13831) );
  OR2_X1 U13785 ( .A1(n13843), .A2(n13844), .ZN(n13830) );
  AND2_X1 U13786 ( .A1(n13827), .A2(n13826), .ZN(n13844) );
  AND2_X1 U13787 ( .A1(n13824), .A2(n13845), .ZN(n13843) );
  OR2_X1 U13788 ( .A1(n13826), .A2(n13827), .ZN(n13845) );
  OR2_X1 U13789 ( .A1(n8040), .A2(n8034), .ZN(n13827) );
  OR2_X1 U13790 ( .A1(n13846), .A2(n13847), .ZN(n13826) );
  AND2_X1 U13791 ( .A1(n8041), .A2(n13823), .ZN(n13847) );
  AND2_X1 U13792 ( .A1(n13821), .A2(n13848), .ZN(n13846) );
  OR2_X1 U13793 ( .A1(n13823), .A2(n8041), .ZN(n13848) );
  OR2_X1 U13794 ( .A1(n8039), .A2(n8040), .ZN(n8041) );
  OR2_X1 U13795 ( .A1(n13849), .A2(n13850), .ZN(n13823) );
  AND2_X1 U13796 ( .A1(n13820), .A2(n13819), .ZN(n13850) );
  AND2_X1 U13797 ( .A1(n13817), .A2(n13851), .ZN(n13849) );
  OR2_X1 U13798 ( .A1(n13819), .A2(n13820), .ZN(n13851) );
  OR2_X1 U13799 ( .A1(n8040), .A2(n8043), .ZN(n13820) );
  OR2_X1 U13800 ( .A1(n13852), .A2(n13853), .ZN(n13819) );
  AND2_X1 U13801 ( .A1(n13816), .A2(n13815), .ZN(n13853) );
  AND2_X1 U13802 ( .A1(n13813), .A2(n13854), .ZN(n13852) );
  OR2_X1 U13803 ( .A1(n13815), .A2(n13816), .ZN(n13854) );
  OR2_X1 U13804 ( .A1(n8040), .A2(n8048), .ZN(n13816) );
  OR2_X1 U13805 ( .A1(n13855), .A2(n13856), .ZN(n13815) );
  AND2_X1 U13806 ( .A1(n13812), .A2(n13811), .ZN(n13856) );
  AND2_X1 U13807 ( .A1(n13809), .A2(n13857), .ZN(n13855) );
  OR2_X1 U13808 ( .A1(n13811), .A2(n13812), .ZN(n13857) );
  OR2_X1 U13809 ( .A1(n8040), .A2(n8052), .ZN(n13812) );
  OR2_X1 U13810 ( .A1(n13858), .A2(n13859), .ZN(n13811) );
  AND2_X1 U13811 ( .A1(n13808), .A2(n13807), .ZN(n13859) );
  AND2_X1 U13812 ( .A1(n13805), .A2(n13860), .ZN(n13858) );
  OR2_X1 U13813 ( .A1(n13807), .A2(n13808), .ZN(n13860) );
  OR2_X1 U13814 ( .A1(n8040), .A2(n8057), .ZN(n13808) );
  OR2_X1 U13815 ( .A1(n13861), .A2(n13862), .ZN(n13807) );
  AND2_X1 U13816 ( .A1(n13804), .A2(n13803), .ZN(n13862) );
  AND2_X1 U13817 ( .A1(n13801), .A2(n13863), .ZN(n13861) );
  OR2_X1 U13818 ( .A1(n13803), .A2(n13804), .ZN(n13863) );
  OR2_X1 U13819 ( .A1(n8040), .A2(n8061), .ZN(n13804) );
  OR2_X1 U13820 ( .A1(n13864), .A2(n13865), .ZN(n13803) );
  AND2_X1 U13821 ( .A1(n13800), .A2(n13799), .ZN(n13865) );
  AND2_X1 U13822 ( .A1(n13797), .A2(n13866), .ZN(n13864) );
  OR2_X1 U13823 ( .A1(n13799), .A2(n13800), .ZN(n13866) );
  OR2_X1 U13824 ( .A1(n8040), .A2(n8066), .ZN(n13800) );
  OR2_X1 U13825 ( .A1(n13867), .A2(n13868), .ZN(n13799) );
  AND2_X1 U13826 ( .A1(n13796), .A2(n13795), .ZN(n13868) );
  AND2_X1 U13827 ( .A1(n13793), .A2(n13869), .ZN(n13867) );
  OR2_X1 U13828 ( .A1(n13795), .A2(n13796), .ZN(n13869) );
  OR2_X1 U13829 ( .A1(n8040), .A2(n8070), .ZN(n13796) );
  OR2_X1 U13830 ( .A1(n13870), .A2(n13871), .ZN(n13795) );
  AND2_X1 U13831 ( .A1(n13792), .A2(n13791), .ZN(n13871) );
  AND2_X1 U13832 ( .A1(n13789), .A2(n13872), .ZN(n13870) );
  OR2_X1 U13833 ( .A1(n13791), .A2(n13792), .ZN(n13872) );
  OR2_X1 U13834 ( .A1(n8040), .A2(n8075), .ZN(n13792) );
  OR2_X1 U13835 ( .A1(n13873), .A2(n13874), .ZN(n13791) );
  AND2_X1 U13836 ( .A1(n13788), .A2(n13787), .ZN(n13874) );
  AND2_X1 U13837 ( .A1(n13785), .A2(n13875), .ZN(n13873) );
  OR2_X1 U13838 ( .A1(n13787), .A2(n13788), .ZN(n13875) );
  OR2_X1 U13839 ( .A1(n8040), .A2(n8079), .ZN(n13788) );
  OR2_X1 U13840 ( .A1(n13876), .A2(n13877), .ZN(n13787) );
  AND2_X1 U13841 ( .A1(n13784), .A2(n13783), .ZN(n13877) );
  AND2_X1 U13842 ( .A1(n13781), .A2(n13878), .ZN(n13876) );
  OR2_X1 U13843 ( .A1(n13783), .A2(n13784), .ZN(n13878) );
  OR2_X1 U13844 ( .A1(n8040), .A2(n8084), .ZN(n13784) );
  OR2_X1 U13845 ( .A1(n13879), .A2(n13880), .ZN(n13783) );
  AND2_X1 U13846 ( .A1(n13780), .A2(n13779), .ZN(n13880) );
  AND2_X1 U13847 ( .A1(n13777), .A2(n13881), .ZN(n13879) );
  OR2_X1 U13848 ( .A1(n13779), .A2(n13780), .ZN(n13881) );
  OR2_X1 U13849 ( .A1(n8040), .A2(n8088), .ZN(n13780) );
  OR2_X1 U13850 ( .A1(n13882), .A2(n13883), .ZN(n13779) );
  AND2_X1 U13851 ( .A1(n13776), .A2(n13775), .ZN(n13883) );
  AND2_X1 U13852 ( .A1(n13773), .A2(n13884), .ZN(n13882) );
  OR2_X1 U13853 ( .A1(n13775), .A2(n13776), .ZN(n13884) );
  OR2_X1 U13854 ( .A1(n8040), .A2(n8093), .ZN(n13776) );
  OR2_X1 U13855 ( .A1(n13885), .A2(n13886), .ZN(n13775) );
  AND2_X1 U13856 ( .A1(n13772), .A2(n13771), .ZN(n13886) );
  AND2_X1 U13857 ( .A1(n13769), .A2(n13887), .ZN(n13885) );
  OR2_X1 U13858 ( .A1(n13771), .A2(n13772), .ZN(n13887) );
  OR2_X1 U13859 ( .A1(n8040), .A2(n8097), .ZN(n13772) );
  OR2_X1 U13860 ( .A1(n13888), .A2(n13889), .ZN(n13771) );
  AND2_X1 U13861 ( .A1(n13768), .A2(n13767), .ZN(n13889) );
  AND2_X1 U13862 ( .A1(n13765), .A2(n13890), .ZN(n13888) );
  OR2_X1 U13863 ( .A1(n13767), .A2(n13768), .ZN(n13890) );
  OR2_X1 U13864 ( .A1(n8040), .A2(n8102), .ZN(n13768) );
  OR2_X1 U13865 ( .A1(n13891), .A2(n13892), .ZN(n13767) );
  AND2_X1 U13866 ( .A1(n13761), .A2(n13764), .ZN(n13892) );
  AND2_X1 U13867 ( .A1(n13893), .A2(n13763), .ZN(n13891) );
  OR2_X1 U13868 ( .A1(n13894), .A2(n13895), .ZN(n13763) );
  AND2_X1 U13869 ( .A1(n13760), .A2(n13759), .ZN(n13895) );
  AND2_X1 U13870 ( .A1(n13757), .A2(n13896), .ZN(n13894) );
  OR2_X1 U13871 ( .A1(n13759), .A2(n13760), .ZN(n13896) );
  OR2_X1 U13872 ( .A1(n8040), .A2(n8109), .ZN(n13760) );
  OR2_X1 U13873 ( .A1(n13897), .A2(n13898), .ZN(n13759) );
  AND2_X1 U13874 ( .A1(n13753), .A2(n13756), .ZN(n13898) );
  AND2_X1 U13875 ( .A1(n13899), .A2(n13755), .ZN(n13897) );
  OR2_X1 U13876 ( .A1(n13900), .A2(n13901), .ZN(n13755) );
  AND2_X1 U13877 ( .A1(n13749), .A2(n13752), .ZN(n13901) );
  AND2_X1 U13878 ( .A1(n13902), .A2(n13751), .ZN(n13900) );
  OR2_X1 U13879 ( .A1(n13903), .A2(n13904), .ZN(n13751) );
  AND2_X1 U13880 ( .A1(n13745), .A2(n13748), .ZN(n13904) );
  AND2_X1 U13881 ( .A1(n13905), .A2(n13747), .ZN(n13903) );
  OR2_X1 U13882 ( .A1(n13906), .A2(n13907), .ZN(n13747) );
  AND2_X1 U13883 ( .A1(n13741), .A2(n13744), .ZN(n13907) );
  AND2_X1 U13884 ( .A1(n13908), .A2(n13743), .ZN(n13906) );
  OR2_X1 U13885 ( .A1(n13909), .A2(n13910), .ZN(n13743) );
  AND2_X1 U13886 ( .A1(n13737), .A2(n13740), .ZN(n13910) );
  AND2_X1 U13887 ( .A1(n13911), .A2(n13739), .ZN(n13909) );
  OR2_X1 U13888 ( .A1(n13912), .A2(n13913), .ZN(n13739) );
  AND2_X1 U13889 ( .A1(n13733), .A2(n13736), .ZN(n13913) );
  AND2_X1 U13890 ( .A1(n13914), .A2(n13915), .ZN(n13912) );
  OR2_X1 U13891 ( .A1(n13736), .A2(n13733), .ZN(n13915) );
  OR2_X1 U13892 ( .A1(n8040), .A2(n8127), .ZN(n13733) );
  OR3_X1 U13893 ( .A1(n8040), .A2(n8981), .A3(n8035), .ZN(n13736) );
  INV_X1 U13894 ( .A(n13735), .ZN(n13914) );
  OR2_X1 U13895 ( .A1(n13916), .A2(n13917), .ZN(n13735) );
  AND2_X1 U13896 ( .A1(b_6_), .A2(n13918), .ZN(n13917) );
  OR2_X1 U13897 ( .A1(n13919), .A2(n7598), .ZN(n13918) );
  AND2_X1 U13898 ( .A1(a_30_), .A2(n8031), .ZN(n13919) );
  AND2_X1 U13899 ( .A1(b_5_), .A2(n13920), .ZN(n13916) );
  OR2_X1 U13900 ( .A1(n13921), .A2(n7601), .ZN(n13920) );
  AND2_X1 U13901 ( .A1(a_31_), .A2(n8035), .ZN(n13921) );
  OR2_X1 U13902 ( .A1(n13740), .A2(n13737), .ZN(n13911) );
  XNOR2_X1 U13903 ( .A(n13922), .B(n13923), .ZN(n13737) );
  XOR2_X1 U13904 ( .A(n13924), .B(n13925), .Z(n13923) );
  OR2_X1 U13905 ( .A1(n8040), .A2(n8124), .ZN(n13740) );
  OR2_X1 U13906 ( .A1(n13744), .A2(n13741), .ZN(n13908) );
  XOR2_X1 U13907 ( .A(n13926), .B(n13927), .Z(n13741) );
  XOR2_X1 U13908 ( .A(n13928), .B(n13929), .Z(n13927) );
  OR2_X1 U13909 ( .A1(n8040), .A2(n8121), .ZN(n13744) );
  OR2_X1 U13910 ( .A1(n13748), .A2(n13745), .ZN(n13905) );
  XOR2_X1 U13911 ( .A(n13930), .B(n13931), .Z(n13745) );
  XOR2_X1 U13912 ( .A(n13932), .B(n13933), .Z(n13931) );
  OR2_X1 U13913 ( .A1(n8040), .A2(n8118), .ZN(n13748) );
  OR2_X1 U13914 ( .A1(n13752), .A2(n13749), .ZN(n13902) );
  XOR2_X1 U13915 ( .A(n13934), .B(n13935), .Z(n13749) );
  XOR2_X1 U13916 ( .A(n13936), .B(n13937), .Z(n13935) );
  OR2_X1 U13917 ( .A1(n8040), .A2(n8115), .ZN(n13752) );
  OR2_X1 U13918 ( .A1(n13756), .A2(n13753), .ZN(n13899) );
  XOR2_X1 U13919 ( .A(n13938), .B(n13939), .Z(n13753) );
  XOR2_X1 U13920 ( .A(n13940), .B(n13941), .Z(n13939) );
  OR2_X1 U13921 ( .A1(n8040), .A2(n8112), .ZN(n13756) );
  XOR2_X1 U13922 ( .A(n13942), .B(n13943), .Z(n13757) );
  XOR2_X1 U13923 ( .A(n13944), .B(n13945), .Z(n13943) );
  OR2_X1 U13924 ( .A1(n13764), .A2(n13761), .ZN(n13893) );
  XOR2_X1 U13925 ( .A(n13946), .B(n13947), .Z(n13761) );
  XOR2_X1 U13926 ( .A(n13948), .B(n13949), .Z(n13947) );
  OR2_X1 U13927 ( .A1(n8040), .A2(n8106), .ZN(n13764) );
  XOR2_X1 U13928 ( .A(n13950), .B(n13951), .Z(n13765) );
  XOR2_X1 U13929 ( .A(n13952), .B(n13953), .Z(n13951) );
  XOR2_X1 U13930 ( .A(n13954), .B(n13955), .Z(n13769) );
  XOR2_X1 U13931 ( .A(n13956), .B(n13957), .Z(n13955) );
  XOR2_X1 U13932 ( .A(n13958), .B(n13959), .Z(n13773) );
  XOR2_X1 U13933 ( .A(n13960), .B(n13961), .Z(n13959) );
  XOR2_X1 U13934 ( .A(n13962), .B(n13963), .Z(n13777) );
  XOR2_X1 U13935 ( .A(n13964), .B(n13965), .Z(n13963) );
  XOR2_X1 U13936 ( .A(n13966), .B(n13967), .Z(n13781) );
  XOR2_X1 U13937 ( .A(n13968), .B(n13969), .Z(n13967) );
  XOR2_X1 U13938 ( .A(n13970), .B(n13971), .Z(n13785) );
  XOR2_X1 U13939 ( .A(n13972), .B(n13973), .Z(n13971) );
  XOR2_X1 U13940 ( .A(n13974), .B(n13975), .Z(n13789) );
  XOR2_X1 U13941 ( .A(n13976), .B(n13977), .Z(n13975) );
  XOR2_X1 U13942 ( .A(n13978), .B(n13979), .Z(n13793) );
  XOR2_X1 U13943 ( .A(n13980), .B(n13981), .Z(n13979) );
  XOR2_X1 U13944 ( .A(n13982), .B(n13983), .Z(n13797) );
  XOR2_X1 U13945 ( .A(n13984), .B(n13985), .Z(n13983) );
  XOR2_X1 U13946 ( .A(n13986), .B(n13987), .Z(n13801) );
  XOR2_X1 U13947 ( .A(n13988), .B(n13989), .Z(n13987) );
  XOR2_X1 U13948 ( .A(n13990), .B(n13991), .Z(n13805) );
  XOR2_X1 U13949 ( .A(n13992), .B(n13993), .Z(n13991) );
  XOR2_X1 U13950 ( .A(n13994), .B(n13995), .Z(n13809) );
  XOR2_X1 U13951 ( .A(n13996), .B(n13997), .Z(n13995) );
  XOR2_X1 U13952 ( .A(n13998), .B(n13999), .Z(n13813) );
  XOR2_X1 U13953 ( .A(n14000), .B(n14001), .Z(n13999) );
  XOR2_X1 U13954 ( .A(n14002), .B(n14003), .Z(n13817) );
  XOR2_X1 U13955 ( .A(n14004), .B(n14005), .Z(n14003) );
  XOR2_X1 U13956 ( .A(n14006), .B(n14007), .Z(n13821) );
  XOR2_X1 U13957 ( .A(n14008), .B(n14009), .Z(n14007) );
  XOR2_X1 U13958 ( .A(n14010), .B(n14011), .Z(n13824) );
  XOR2_X1 U13959 ( .A(n14012), .B(n14013), .Z(n14011) );
  XNOR2_X1 U13960 ( .A(n14014), .B(n14015), .ZN(n13828) );
  XOR2_X1 U13961 ( .A(n7939), .B(n14016), .Z(n14014) );
  INV_X1 U13962 ( .A(n8036), .ZN(n7939) );
  XOR2_X1 U13963 ( .A(n14017), .B(n14018), .Z(n13832) );
  XOR2_X1 U13964 ( .A(n14019), .B(n14020), .Z(n14018) );
  XOR2_X1 U13965 ( .A(n8554), .B(n14021), .Z(n8547) );
  XOR2_X1 U13966 ( .A(n8553), .B(n8552), .Z(n14021) );
  OR2_X1 U13967 ( .A1(n8035), .A2(n8025), .ZN(n8552) );
  OR2_X1 U13968 ( .A1(n14022), .A2(n14023), .ZN(n8553) );
  AND2_X1 U13969 ( .A1(n14020), .A2(n14019), .ZN(n14023) );
  AND2_X1 U13970 ( .A1(n14017), .A2(n14024), .ZN(n14022) );
  OR2_X1 U13971 ( .A1(n14019), .A2(n14020), .ZN(n14024) );
  OR2_X1 U13972 ( .A1(n8030), .A2(n8035), .ZN(n14020) );
  OR2_X1 U13973 ( .A1(n14025), .A2(n14026), .ZN(n14019) );
  AND2_X1 U13974 ( .A1(n14016), .A2(n8036), .ZN(n14026) );
  AND2_X1 U13975 ( .A1(n14015), .A2(n14027), .ZN(n14025) );
  OR2_X1 U13976 ( .A1(n8036), .A2(n14016), .ZN(n14027) );
  OR2_X1 U13977 ( .A1(n14028), .A2(n14029), .ZN(n14016) );
  AND2_X1 U13978 ( .A1(n14013), .A2(n14012), .ZN(n14029) );
  AND2_X1 U13979 ( .A1(n14010), .A2(n14030), .ZN(n14028) );
  OR2_X1 U13980 ( .A1(n14012), .A2(n14013), .ZN(n14030) );
  OR2_X1 U13981 ( .A1(n8039), .A2(n8035), .ZN(n14013) );
  OR2_X1 U13982 ( .A1(n14031), .A2(n14032), .ZN(n14012) );
  AND2_X1 U13983 ( .A1(n14009), .A2(n14008), .ZN(n14032) );
  AND2_X1 U13984 ( .A1(n14006), .A2(n14033), .ZN(n14031) );
  OR2_X1 U13985 ( .A1(n14008), .A2(n14009), .ZN(n14033) );
  OR2_X1 U13986 ( .A1(n8043), .A2(n8035), .ZN(n14009) );
  OR2_X1 U13987 ( .A1(n14034), .A2(n14035), .ZN(n14008) );
  AND2_X1 U13988 ( .A1(n14005), .A2(n14004), .ZN(n14035) );
  AND2_X1 U13989 ( .A1(n14002), .A2(n14036), .ZN(n14034) );
  OR2_X1 U13990 ( .A1(n14004), .A2(n14005), .ZN(n14036) );
  OR2_X1 U13991 ( .A1(n8048), .A2(n8035), .ZN(n14005) );
  OR2_X1 U13992 ( .A1(n14037), .A2(n14038), .ZN(n14004) );
  AND2_X1 U13993 ( .A1(n14001), .A2(n14000), .ZN(n14038) );
  AND2_X1 U13994 ( .A1(n13998), .A2(n14039), .ZN(n14037) );
  OR2_X1 U13995 ( .A1(n14000), .A2(n14001), .ZN(n14039) );
  OR2_X1 U13996 ( .A1(n8052), .A2(n8035), .ZN(n14001) );
  OR2_X1 U13997 ( .A1(n14040), .A2(n14041), .ZN(n14000) );
  AND2_X1 U13998 ( .A1(n13997), .A2(n13996), .ZN(n14041) );
  AND2_X1 U13999 ( .A1(n13994), .A2(n14042), .ZN(n14040) );
  OR2_X1 U14000 ( .A1(n13996), .A2(n13997), .ZN(n14042) );
  OR2_X1 U14001 ( .A1(n8057), .A2(n8035), .ZN(n13997) );
  OR2_X1 U14002 ( .A1(n14043), .A2(n14044), .ZN(n13996) );
  AND2_X1 U14003 ( .A1(n13993), .A2(n13992), .ZN(n14044) );
  AND2_X1 U14004 ( .A1(n13990), .A2(n14045), .ZN(n14043) );
  OR2_X1 U14005 ( .A1(n13992), .A2(n13993), .ZN(n14045) );
  OR2_X1 U14006 ( .A1(n8061), .A2(n8035), .ZN(n13993) );
  OR2_X1 U14007 ( .A1(n14046), .A2(n14047), .ZN(n13992) );
  AND2_X1 U14008 ( .A1(n13989), .A2(n13988), .ZN(n14047) );
  AND2_X1 U14009 ( .A1(n13986), .A2(n14048), .ZN(n14046) );
  OR2_X1 U14010 ( .A1(n13988), .A2(n13989), .ZN(n14048) );
  OR2_X1 U14011 ( .A1(n8066), .A2(n8035), .ZN(n13989) );
  OR2_X1 U14012 ( .A1(n14049), .A2(n14050), .ZN(n13988) );
  AND2_X1 U14013 ( .A1(n13985), .A2(n13984), .ZN(n14050) );
  AND2_X1 U14014 ( .A1(n13982), .A2(n14051), .ZN(n14049) );
  OR2_X1 U14015 ( .A1(n13984), .A2(n13985), .ZN(n14051) );
  OR2_X1 U14016 ( .A1(n8070), .A2(n8035), .ZN(n13985) );
  OR2_X1 U14017 ( .A1(n14052), .A2(n14053), .ZN(n13984) );
  AND2_X1 U14018 ( .A1(n13981), .A2(n13980), .ZN(n14053) );
  AND2_X1 U14019 ( .A1(n13978), .A2(n14054), .ZN(n14052) );
  OR2_X1 U14020 ( .A1(n13980), .A2(n13981), .ZN(n14054) );
  OR2_X1 U14021 ( .A1(n8075), .A2(n8035), .ZN(n13981) );
  OR2_X1 U14022 ( .A1(n14055), .A2(n14056), .ZN(n13980) );
  AND2_X1 U14023 ( .A1(n13977), .A2(n13976), .ZN(n14056) );
  AND2_X1 U14024 ( .A1(n13974), .A2(n14057), .ZN(n14055) );
  OR2_X1 U14025 ( .A1(n13976), .A2(n13977), .ZN(n14057) );
  OR2_X1 U14026 ( .A1(n8079), .A2(n8035), .ZN(n13977) );
  OR2_X1 U14027 ( .A1(n14058), .A2(n14059), .ZN(n13976) );
  AND2_X1 U14028 ( .A1(n13973), .A2(n13972), .ZN(n14059) );
  AND2_X1 U14029 ( .A1(n13970), .A2(n14060), .ZN(n14058) );
  OR2_X1 U14030 ( .A1(n13972), .A2(n13973), .ZN(n14060) );
  OR2_X1 U14031 ( .A1(n8084), .A2(n8035), .ZN(n13973) );
  OR2_X1 U14032 ( .A1(n14061), .A2(n14062), .ZN(n13972) );
  AND2_X1 U14033 ( .A1(n13969), .A2(n13968), .ZN(n14062) );
  AND2_X1 U14034 ( .A1(n13966), .A2(n14063), .ZN(n14061) );
  OR2_X1 U14035 ( .A1(n13968), .A2(n13969), .ZN(n14063) );
  OR2_X1 U14036 ( .A1(n8088), .A2(n8035), .ZN(n13969) );
  OR2_X1 U14037 ( .A1(n14064), .A2(n14065), .ZN(n13968) );
  AND2_X1 U14038 ( .A1(n13965), .A2(n13964), .ZN(n14065) );
  AND2_X1 U14039 ( .A1(n13962), .A2(n14066), .ZN(n14064) );
  OR2_X1 U14040 ( .A1(n13964), .A2(n13965), .ZN(n14066) );
  OR2_X1 U14041 ( .A1(n8093), .A2(n8035), .ZN(n13965) );
  OR2_X1 U14042 ( .A1(n14067), .A2(n14068), .ZN(n13964) );
  AND2_X1 U14043 ( .A1(n13961), .A2(n13960), .ZN(n14068) );
  AND2_X1 U14044 ( .A1(n13958), .A2(n14069), .ZN(n14067) );
  OR2_X1 U14045 ( .A1(n13960), .A2(n13961), .ZN(n14069) );
  OR2_X1 U14046 ( .A1(n8097), .A2(n8035), .ZN(n13961) );
  OR2_X1 U14047 ( .A1(n14070), .A2(n14071), .ZN(n13960) );
  AND2_X1 U14048 ( .A1(n13957), .A2(n13956), .ZN(n14071) );
  AND2_X1 U14049 ( .A1(n13954), .A2(n14072), .ZN(n14070) );
  OR2_X1 U14050 ( .A1(n13956), .A2(n13957), .ZN(n14072) );
  OR2_X1 U14051 ( .A1(n8102), .A2(n8035), .ZN(n13957) );
  OR2_X1 U14052 ( .A1(n14073), .A2(n14074), .ZN(n13956) );
  AND2_X1 U14053 ( .A1(n13953), .A2(n13952), .ZN(n14074) );
  AND2_X1 U14054 ( .A1(n13950), .A2(n14075), .ZN(n14073) );
  OR2_X1 U14055 ( .A1(n13952), .A2(n13953), .ZN(n14075) );
  OR2_X1 U14056 ( .A1(n8106), .A2(n8035), .ZN(n13953) );
  OR2_X1 U14057 ( .A1(n14076), .A2(n14077), .ZN(n13952) );
  AND2_X1 U14058 ( .A1(n13946), .A2(n13949), .ZN(n14077) );
  AND2_X1 U14059 ( .A1(n14078), .A2(n13948), .ZN(n14076) );
  OR2_X1 U14060 ( .A1(n14079), .A2(n14080), .ZN(n13948) );
  AND2_X1 U14061 ( .A1(n13945), .A2(n13944), .ZN(n14080) );
  AND2_X1 U14062 ( .A1(n13942), .A2(n14081), .ZN(n14079) );
  OR2_X1 U14063 ( .A1(n13944), .A2(n13945), .ZN(n14081) );
  OR2_X1 U14064 ( .A1(n8112), .A2(n8035), .ZN(n13945) );
  OR2_X1 U14065 ( .A1(n14082), .A2(n14083), .ZN(n13944) );
  AND2_X1 U14066 ( .A1(n13938), .A2(n13941), .ZN(n14083) );
  AND2_X1 U14067 ( .A1(n14084), .A2(n13940), .ZN(n14082) );
  OR2_X1 U14068 ( .A1(n14085), .A2(n14086), .ZN(n13940) );
  AND2_X1 U14069 ( .A1(n13934), .A2(n13937), .ZN(n14086) );
  AND2_X1 U14070 ( .A1(n14087), .A2(n13936), .ZN(n14085) );
  OR2_X1 U14071 ( .A1(n14088), .A2(n14089), .ZN(n13936) );
  AND2_X1 U14072 ( .A1(n13930), .A2(n13933), .ZN(n14089) );
  AND2_X1 U14073 ( .A1(n14090), .A2(n13932), .ZN(n14088) );
  OR2_X1 U14074 ( .A1(n14091), .A2(n14092), .ZN(n13932) );
  AND2_X1 U14075 ( .A1(n13926), .A2(n13929), .ZN(n14092) );
  AND2_X1 U14076 ( .A1(n14093), .A2(n13928), .ZN(n14091) );
  OR2_X1 U14077 ( .A1(n14094), .A2(n14095), .ZN(n13928) );
  AND2_X1 U14078 ( .A1(n13922), .A2(n13925), .ZN(n14095) );
  AND2_X1 U14079 ( .A1(n14096), .A2(n14097), .ZN(n14094) );
  OR2_X1 U14080 ( .A1(n13925), .A2(n13922), .ZN(n14097) );
  OR2_X1 U14081 ( .A1(n8127), .A2(n8035), .ZN(n13922) );
  OR3_X1 U14082 ( .A1(n8031), .A2(n8981), .A3(n8035), .ZN(n13925) );
  INV_X1 U14083 ( .A(n13924), .ZN(n14096) );
  OR2_X1 U14084 ( .A1(n14098), .A2(n14099), .ZN(n13924) );
  AND2_X1 U14085 ( .A1(b_5_), .A2(n14100), .ZN(n14099) );
  OR2_X1 U14086 ( .A1(n14101), .A2(n7598), .ZN(n14100) );
  AND2_X1 U14087 ( .A1(a_30_), .A2(n8026), .ZN(n14101) );
  AND2_X1 U14088 ( .A1(b_4_), .A2(n14102), .ZN(n14098) );
  OR2_X1 U14089 ( .A1(n14103), .A2(n7601), .ZN(n14102) );
  AND2_X1 U14090 ( .A1(a_31_), .A2(n8031), .ZN(n14103) );
  OR2_X1 U14091 ( .A1(n13929), .A2(n13926), .ZN(n14093) );
  XNOR2_X1 U14092 ( .A(n14104), .B(n14105), .ZN(n13926) );
  XOR2_X1 U14093 ( .A(n14106), .B(n14107), .Z(n14105) );
  OR2_X1 U14094 ( .A1(n8124), .A2(n8035), .ZN(n13929) );
  OR2_X1 U14095 ( .A1(n13933), .A2(n13930), .ZN(n14090) );
  XOR2_X1 U14096 ( .A(n14108), .B(n14109), .Z(n13930) );
  XOR2_X1 U14097 ( .A(n14110), .B(n14111), .Z(n14109) );
  OR2_X1 U14098 ( .A1(n8121), .A2(n8035), .ZN(n13933) );
  OR2_X1 U14099 ( .A1(n13937), .A2(n13934), .ZN(n14087) );
  XOR2_X1 U14100 ( .A(n14112), .B(n14113), .Z(n13934) );
  XOR2_X1 U14101 ( .A(n14114), .B(n14115), .Z(n14113) );
  OR2_X1 U14102 ( .A1(n8118), .A2(n8035), .ZN(n13937) );
  OR2_X1 U14103 ( .A1(n13941), .A2(n13938), .ZN(n14084) );
  XOR2_X1 U14104 ( .A(n14116), .B(n14117), .Z(n13938) );
  XOR2_X1 U14105 ( .A(n14118), .B(n14119), .Z(n14117) );
  OR2_X1 U14106 ( .A1(n8115), .A2(n8035), .ZN(n13941) );
  XOR2_X1 U14107 ( .A(n14120), .B(n14121), .Z(n13942) );
  XOR2_X1 U14108 ( .A(n14122), .B(n14123), .Z(n14121) );
  OR2_X1 U14109 ( .A1(n13949), .A2(n13946), .ZN(n14078) );
  XOR2_X1 U14110 ( .A(n14124), .B(n14125), .Z(n13946) );
  XOR2_X1 U14111 ( .A(n14126), .B(n14127), .Z(n14125) );
  OR2_X1 U14112 ( .A1(n8109), .A2(n8035), .ZN(n13949) );
  XOR2_X1 U14113 ( .A(n14128), .B(n14129), .Z(n13950) );
  XOR2_X1 U14114 ( .A(n14130), .B(n14131), .Z(n14129) );
  XOR2_X1 U14115 ( .A(n14132), .B(n14133), .Z(n13954) );
  XOR2_X1 U14116 ( .A(n14134), .B(n14135), .Z(n14133) );
  XOR2_X1 U14117 ( .A(n14136), .B(n14137), .Z(n13958) );
  XOR2_X1 U14118 ( .A(n14138), .B(n14139), .Z(n14137) );
  XOR2_X1 U14119 ( .A(n14140), .B(n14141), .Z(n13962) );
  XOR2_X1 U14120 ( .A(n14142), .B(n14143), .Z(n14141) );
  XOR2_X1 U14121 ( .A(n14144), .B(n14145), .Z(n13966) );
  XOR2_X1 U14122 ( .A(n14146), .B(n14147), .Z(n14145) );
  XOR2_X1 U14123 ( .A(n14148), .B(n14149), .Z(n13970) );
  XOR2_X1 U14124 ( .A(n14150), .B(n14151), .Z(n14149) );
  XOR2_X1 U14125 ( .A(n14152), .B(n14153), .Z(n13974) );
  XOR2_X1 U14126 ( .A(n14154), .B(n14155), .Z(n14153) );
  XOR2_X1 U14127 ( .A(n14156), .B(n14157), .Z(n13978) );
  XOR2_X1 U14128 ( .A(n14158), .B(n14159), .Z(n14157) );
  XOR2_X1 U14129 ( .A(n14160), .B(n14161), .Z(n13982) );
  XOR2_X1 U14130 ( .A(n14162), .B(n14163), .Z(n14161) );
  XOR2_X1 U14131 ( .A(n14164), .B(n14165), .Z(n13986) );
  XOR2_X1 U14132 ( .A(n14166), .B(n14167), .Z(n14165) );
  XOR2_X1 U14133 ( .A(n14168), .B(n14169), .Z(n13990) );
  XOR2_X1 U14134 ( .A(n14170), .B(n14171), .Z(n14169) );
  XOR2_X1 U14135 ( .A(n14172), .B(n14173), .Z(n13994) );
  XOR2_X1 U14136 ( .A(n14174), .B(n14175), .Z(n14173) );
  XOR2_X1 U14137 ( .A(n14176), .B(n14177), .Z(n13998) );
  XOR2_X1 U14138 ( .A(n14178), .B(n14179), .Z(n14177) );
  XOR2_X1 U14139 ( .A(n14180), .B(n14181), .Z(n14002) );
  XOR2_X1 U14140 ( .A(n14182), .B(n14183), .Z(n14181) );
  XOR2_X1 U14141 ( .A(n14184), .B(n14185), .Z(n14006) );
  XOR2_X1 U14142 ( .A(n14186), .B(n14187), .Z(n14185) );
  XOR2_X1 U14143 ( .A(n14188), .B(n14189), .Z(n14010) );
  XOR2_X1 U14144 ( .A(n14190), .B(n14191), .Z(n14189) );
  OR2_X1 U14145 ( .A1(n8034), .A2(n8035), .ZN(n8036) );
  INV_X1 U14146 ( .A(b_6_), .ZN(n8035) );
  XOR2_X1 U14147 ( .A(n14192), .B(n14193), .Z(n14015) );
  XOR2_X1 U14148 ( .A(n14194), .B(n14195), .Z(n14193) );
  XOR2_X1 U14149 ( .A(n14196), .B(n14197), .Z(n14017) );
  XOR2_X1 U14150 ( .A(n14198), .B(n14199), .Z(n14197) );
  XOR2_X1 U14151 ( .A(n8560), .B(n14200), .Z(n8554) );
  XOR2_X1 U14152 ( .A(n8559), .B(n8032), .Z(n14200) );
  OR2_X1 U14153 ( .A1(n8030), .A2(n8031), .ZN(n8032) );
  OR2_X1 U14154 ( .A1(n14201), .A2(n14202), .ZN(n8559) );
  AND2_X1 U14155 ( .A1(n14199), .A2(n14198), .ZN(n14202) );
  AND2_X1 U14156 ( .A1(n14196), .A2(n14203), .ZN(n14201) );
  OR2_X1 U14157 ( .A1(n14198), .A2(n14199), .ZN(n14203) );
  OR2_X1 U14158 ( .A1(n8031), .A2(n8034), .ZN(n14199) );
  OR2_X1 U14159 ( .A1(n14204), .A2(n14205), .ZN(n14198) );
  AND2_X1 U14160 ( .A1(n14195), .A2(n14194), .ZN(n14205) );
  AND2_X1 U14161 ( .A1(n14192), .A2(n14206), .ZN(n14204) );
  OR2_X1 U14162 ( .A1(n14194), .A2(n14195), .ZN(n14206) );
  OR2_X1 U14163 ( .A1(n8031), .A2(n8039), .ZN(n14195) );
  OR2_X1 U14164 ( .A1(n14207), .A2(n14208), .ZN(n14194) );
  AND2_X1 U14165 ( .A1(n14191), .A2(n14190), .ZN(n14208) );
  AND2_X1 U14166 ( .A1(n14188), .A2(n14209), .ZN(n14207) );
  OR2_X1 U14167 ( .A1(n14190), .A2(n14191), .ZN(n14209) );
  OR2_X1 U14168 ( .A1(n8031), .A2(n8043), .ZN(n14191) );
  OR2_X1 U14169 ( .A1(n14210), .A2(n14211), .ZN(n14190) );
  AND2_X1 U14170 ( .A1(n14187), .A2(n14186), .ZN(n14211) );
  AND2_X1 U14171 ( .A1(n14184), .A2(n14212), .ZN(n14210) );
  OR2_X1 U14172 ( .A1(n14186), .A2(n14187), .ZN(n14212) );
  OR2_X1 U14173 ( .A1(n8031), .A2(n8048), .ZN(n14187) );
  OR2_X1 U14174 ( .A1(n14213), .A2(n14214), .ZN(n14186) );
  AND2_X1 U14175 ( .A1(n14183), .A2(n14182), .ZN(n14214) );
  AND2_X1 U14176 ( .A1(n14180), .A2(n14215), .ZN(n14213) );
  OR2_X1 U14177 ( .A1(n14182), .A2(n14183), .ZN(n14215) );
  OR2_X1 U14178 ( .A1(n8031), .A2(n8052), .ZN(n14183) );
  OR2_X1 U14179 ( .A1(n14216), .A2(n14217), .ZN(n14182) );
  AND2_X1 U14180 ( .A1(n14179), .A2(n14178), .ZN(n14217) );
  AND2_X1 U14181 ( .A1(n14176), .A2(n14218), .ZN(n14216) );
  OR2_X1 U14182 ( .A1(n14178), .A2(n14179), .ZN(n14218) );
  OR2_X1 U14183 ( .A1(n8031), .A2(n8057), .ZN(n14179) );
  OR2_X1 U14184 ( .A1(n14219), .A2(n14220), .ZN(n14178) );
  AND2_X1 U14185 ( .A1(n14175), .A2(n14174), .ZN(n14220) );
  AND2_X1 U14186 ( .A1(n14172), .A2(n14221), .ZN(n14219) );
  OR2_X1 U14187 ( .A1(n14174), .A2(n14175), .ZN(n14221) );
  OR2_X1 U14188 ( .A1(n8031), .A2(n8061), .ZN(n14175) );
  OR2_X1 U14189 ( .A1(n14222), .A2(n14223), .ZN(n14174) );
  AND2_X1 U14190 ( .A1(n14171), .A2(n14170), .ZN(n14223) );
  AND2_X1 U14191 ( .A1(n14168), .A2(n14224), .ZN(n14222) );
  OR2_X1 U14192 ( .A1(n14170), .A2(n14171), .ZN(n14224) );
  OR2_X1 U14193 ( .A1(n8031), .A2(n8066), .ZN(n14171) );
  OR2_X1 U14194 ( .A1(n14225), .A2(n14226), .ZN(n14170) );
  AND2_X1 U14195 ( .A1(n14167), .A2(n14166), .ZN(n14226) );
  AND2_X1 U14196 ( .A1(n14164), .A2(n14227), .ZN(n14225) );
  OR2_X1 U14197 ( .A1(n14166), .A2(n14167), .ZN(n14227) );
  OR2_X1 U14198 ( .A1(n8031), .A2(n8070), .ZN(n14167) );
  OR2_X1 U14199 ( .A1(n14228), .A2(n14229), .ZN(n14166) );
  AND2_X1 U14200 ( .A1(n14163), .A2(n14162), .ZN(n14229) );
  AND2_X1 U14201 ( .A1(n14160), .A2(n14230), .ZN(n14228) );
  OR2_X1 U14202 ( .A1(n14162), .A2(n14163), .ZN(n14230) );
  OR2_X1 U14203 ( .A1(n8031), .A2(n8075), .ZN(n14163) );
  OR2_X1 U14204 ( .A1(n14231), .A2(n14232), .ZN(n14162) );
  AND2_X1 U14205 ( .A1(n14159), .A2(n14158), .ZN(n14232) );
  AND2_X1 U14206 ( .A1(n14156), .A2(n14233), .ZN(n14231) );
  OR2_X1 U14207 ( .A1(n14158), .A2(n14159), .ZN(n14233) );
  OR2_X1 U14208 ( .A1(n8031), .A2(n8079), .ZN(n14159) );
  OR2_X1 U14209 ( .A1(n14234), .A2(n14235), .ZN(n14158) );
  AND2_X1 U14210 ( .A1(n14155), .A2(n14154), .ZN(n14235) );
  AND2_X1 U14211 ( .A1(n14152), .A2(n14236), .ZN(n14234) );
  OR2_X1 U14212 ( .A1(n14154), .A2(n14155), .ZN(n14236) );
  OR2_X1 U14213 ( .A1(n8031), .A2(n8084), .ZN(n14155) );
  OR2_X1 U14214 ( .A1(n14237), .A2(n14238), .ZN(n14154) );
  AND2_X1 U14215 ( .A1(n14151), .A2(n14150), .ZN(n14238) );
  AND2_X1 U14216 ( .A1(n14148), .A2(n14239), .ZN(n14237) );
  OR2_X1 U14217 ( .A1(n14150), .A2(n14151), .ZN(n14239) );
  OR2_X1 U14218 ( .A1(n8031), .A2(n8088), .ZN(n14151) );
  OR2_X1 U14219 ( .A1(n14240), .A2(n14241), .ZN(n14150) );
  AND2_X1 U14220 ( .A1(n14147), .A2(n14146), .ZN(n14241) );
  AND2_X1 U14221 ( .A1(n14144), .A2(n14242), .ZN(n14240) );
  OR2_X1 U14222 ( .A1(n14146), .A2(n14147), .ZN(n14242) );
  OR2_X1 U14223 ( .A1(n8031), .A2(n8093), .ZN(n14147) );
  OR2_X1 U14224 ( .A1(n14243), .A2(n14244), .ZN(n14146) );
  AND2_X1 U14225 ( .A1(n14143), .A2(n14142), .ZN(n14244) );
  AND2_X1 U14226 ( .A1(n14140), .A2(n14245), .ZN(n14243) );
  OR2_X1 U14227 ( .A1(n14142), .A2(n14143), .ZN(n14245) );
  OR2_X1 U14228 ( .A1(n8031), .A2(n8097), .ZN(n14143) );
  OR2_X1 U14229 ( .A1(n14246), .A2(n14247), .ZN(n14142) );
  AND2_X1 U14230 ( .A1(n14139), .A2(n14138), .ZN(n14247) );
  AND2_X1 U14231 ( .A1(n14136), .A2(n14248), .ZN(n14246) );
  OR2_X1 U14232 ( .A1(n14138), .A2(n14139), .ZN(n14248) );
  OR2_X1 U14233 ( .A1(n8031), .A2(n8102), .ZN(n14139) );
  OR2_X1 U14234 ( .A1(n14249), .A2(n14250), .ZN(n14138) );
  AND2_X1 U14235 ( .A1(n14135), .A2(n14134), .ZN(n14250) );
  AND2_X1 U14236 ( .A1(n14132), .A2(n14251), .ZN(n14249) );
  OR2_X1 U14237 ( .A1(n14134), .A2(n14135), .ZN(n14251) );
  OR2_X1 U14238 ( .A1(n8031), .A2(n8106), .ZN(n14135) );
  OR2_X1 U14239 ( .A1(n14252), .A2(n14253), .ZN(n14134) );
  AND2_X1 U14240 ( .A1(n14131), .A2(n14130), .ZN(n14253) );
  AND2_X1 U14241 ( .A1(n14128), .A2(n14254), .ZN(n14252) );
  OR2_X1 U14242 ( .A1(n14130), .A2(n14131), .ZN(n14254) );
  OR2_X1 U14243 ( .A1(n8031), .A2(n8109), .ZN(n14131) );
  OR2_X1 U14244 ( .A1(n14255), .A2(n14256), .ZN(n14130) );
  AND2_X1 U14245 ( .A1(n14124), .A2(n14127), .ZN(n14256) );
  AND2_X1 U14246 ( .A1(n14257), .A2(n14126), .ZN(n14255) );
  OR2_X1 U14247 ( .A1(n14258), .A2(n14259), .ZN(n14126) );
  AND2_X1 U14248 ( .A1(n14123), .A2(n14122), .ZN(n14259) );
  AND2_X1 U14249 ( .A1(n14120), .A2(n14260), .ZN(n14258) );
  OR2_X1 U14250 ( .A1(n14122), .A2(n14123), .ZN(n14260) );
  OR2_X1 U14251 ( .A1(n8031), .A2(n8115), .ZN(n14123) );
  OR2_X1 U14252 ( .A1(n14261), .A2(n14262), .ZN(n14122) );
  AND2_X1 U14253 ( .A1(n14116), .A2(n14119), .ZN(n14262) );
  AND2_X1 U14254 ( .A1(n14263), .A2(n14118), .ZN(n14261) );
  OR2_X1 U14255 ( .A1(n14264), .A2(n14265), .ZN(n14118) );
  AND2_X1 U14256 ( .A1(n14112), .A2(n14115), .ZN(n14265) );
  AND2_X1 U14257 ( .A1(n14266), .A2(n14114), .ZN(n14264) );
  OR2_X1 U14258 ( .A1(n14267), .A2(n14268), .ZN(n14114) );
  AND2_X1 U14259 ( .A1(n14108), .A2(n14111), .ZN(n14268) );
  AND2_X1 U14260 ( .A1(n14269), .A2(n14110), .ZN(n14267) );
  OR2_X1 U14261 ( .A1(n14270), .A2(n14271), .ZN(n14110) );
  AND2_X1 U14262 ( .A1(n14104), .A2(n14107), .ZN(n14271) );
  AND2_X1 U14263 ( .A1(n14272), .A2(n14273), .ZN(n14270) );
  OR2_X1 U14264 ( .A1(n14107), .A2(n14104), .ZN(n14273) );
  OR2_X1 U14265 ( .A1(n8031), .A2(n8127), .ZN(n14104) );
  OR3_X1 U14266 ( .A1(n8026), .A2(n8031), .A3(n8981), .ZN(n14107) );
  INV_X1 U14267 ( .A(n14106), .ZN(n14272) );
  OR2_X1 U14268 ( .A1(n14274), .A2(n14275), .ZN(n14106) );
  AND2_X1 U14269 ( .A1(b_4_), .A2(n14276), .ZN(n14275) );
  OR2_X1 U14270 ( .A1(n14277), .A2(n7598), .ZN(n14276) );
  AND2_X1 U14271 ( .A1(a_30_), .A2(n8022), .ZN(n14277) );
  AND2_X1 U14272 ( .A1(b_3_), .A2(n14278), .ZN(n14274) );
  OR2_X1 U14273 ( .A1(n14279), .A2(n7601), .ZN(n14278) );
  AND2_X1 U14274 ( .A1(a_31_), .A2(n8026), .ZN(n14279) );
  OR2_X1 U14275 ( .A1(n14111), .A2(n14108), .ZN(n14269) );
  XNOR2_X1 U14276 ( .A(n14280), .B(n14281), .ZN(n14108) );
  XOR2_X1 U14277 ( .A(n14282), .B(n14283), .Z(n14281) );
  OR2_X1 U14278 ( .A1(n8031), .A2(n8124), .ZN(n14111) );
  OR2_X1 U14279 ( .A1(n14115), .A2(n14112), .ZN(n14266) );
  XOR2_X1 U14280 ( .A(n14284), .B(n14285), .Z(n14112) );
  XOR2_X1 U14281 ( .A(n14286), .B(n14287), .Z(n14285) );
  OR2_X1 U14282 ( .A1(n8031), .A2(n8121), .ZN(n14115) );
  OR2_X1 U14283 ( .A1(n14119), .A2(n14116), .ZN(n14263) );
  XOR2_X1 U14284 ( .A(n14288), .B(n14289), .Z(n14116) );
  XOR2_X1 U14285 ( .A(n14290), .B(n14291), .Z(n14289) );
  OR2_X1 U14286 ( .A1(n8031), .A2(n8118), .ZN(n14119) );
  XOR2_X1 U14287 ( .A(n14292), .B(n14293), .Z(n14120) );
  XOR2_X1 U14288 ( .A(n14294), .B(n14295), .Z(n14293) );
  OR2_X1 U14289 ( .A1(n14127), .A2(n14124), .ZN(n14257) );
  XOR2_X1 U14290 ( .A(n14296), .B(n14297), .Z(n14124) );
  XOR2_X1 U14291 ( .A(n14298), .B(n14299), .Z(n14297) );
  OR2_X1 U14292 ( .A1(n8031), .A2(n8112), .ZN(n14127) );
  XOR2_X1 U14293 ( .A(n14300), .B(n14301), .Z(n14128) );
  XOR2_X1 U14294 ( .A(n14302), .B(n14303), .Z(n14301) );
  XOR2_X1 U14295 ( .A(n14304), .B(n14305), .Z(n14132) );
  XOR2_X1 U14296 ( .A(n14306), .B(n14307), .Z(n14305) );
  XOR2_X1 U14297 ( .A(n14308), .B(n14309), .Z(n14136) );
  XOR2_X1 U14298 ( .A(n14310), .B(n14311), .Z(n14309) );
  XOR2_X1 U14299 ( .A(n14312), .B(n14313), .Z(n14140) );
  XOR2_X1 U14300 ( .A(n14314), .B(n14315), .Z(n14313) );
  XOR2_X1 U14301 ( .A(n14316), .B(n14317), .Z(n14144) );
  XOR2_X1 U14302 ( .A(n14318), .B(n14319), .Z(n14317) );
  XOR2_X1 U14303 ( .A(n14320), .B(n14321), .Z(n14148) );
  XOR2_X1 U14304 ( .A(n14322), .B(n14323), .Z(n14321) );
  XOR2_X1 U14305 ( .A(n14324), .B(n14325), .Z(n14152) );
  XOR2_X1 U14306 ( .A(n14326), .B(n14327), .Z(n14325) );
  XOR2_X1 U14307 ( .A(n14328), .B(n14329), .Z(n14156) );
  XOR2_X1 U14308 ( .A(n14330), .B(n14331), .Z(n14329) );
  XOR2_X1 U14309 ( .A(n14332), .B(n14333), .Z(n14160) );
  XOR2_X1 U14310 ( .A(n14334), .B(n14335), .Z(n14333) );
  XOR2_X1 U14311 ( .A(n14336), .B(n14337), .Z(n14164) );
  XOR2_X1 U14312 ( .A(n14338), .B(n14339), .Z(n14337) );
  XOR2_X1 U14313 ( .A(n14340), .B(n14341), .Z(n14168) );
  XOR2_X1 U14314 ( .A(n14342), .B(n14343), .Z(n14341) );
  XOR2_X1 U14315 ( .A(n14344), .B(n14345), .Z(n14172) );
  XOR2_X1 U14316 ( .A(n14346), .B(n14347), .Z(n14345) );
  XOR2_X1 U14317 ( .A(n14348), .B(n14349), .Z(n14176) );
  XOR2_X1 U14318 ( .A(n14350), .B(n14351), .Z(n14349) );
  XOR2_X1 U14319 ( .A(n14352), .B(n14353), .Z(n14180) );
  XOR2_X1 U14320 ( .A(n14354), .B(n14355), .Z(n14353) );
  XOR2_X1 U14321 ( .A(n14356), .B(n14357), .Z(n14184) );
  XOR2_X1 U14322 ( .A(n14358), .B(n14359), .Z(n14357) );
  XOR2_X1 U14323 ( .A(n14360), .B(n14361), .Z(n14188) );
  XOR2_X1 U14324 ( .A(n14362), .B(n14363), .Z(n14361) );
  XOR2_X1 U14325 ( .A(n14364), .B(n14365), .Z(n14192) );
  XOR2_X1 U14326 ( .A(n14366), .B(n14367), .Z(n14365) );
  XOR2_X1 U14327 ( .A(n14368), .B(n14369), .Z(n14196) );
  XOR2_X1 U14328 ( .A(n14370), .B(n14371), .Z(n14369) );
  XOR2_X1 U14329 ( .A(n8567), .B(n14372), .Z(n8560) );
  XOR2_X1 U14330 ( .A(n8566), .B(n8565), .Z(n14372) );
  OR2_X1 U14331 ( .A1(n8026), .A2(n8034), .ZN(n8565) );
  OR2_X1 U14332 ( .A1(n14373), .A2(n14374), .ZN(n8566) );
  AND2_X1 U14333 ( .A1(n14371), .A2(n14370), .ZN(n14374) );
  AND2_X1 U14334 ( .A1(n14368), .A2(n14375), .ZN(n14373) );
  OR2_X1 U14335 ( .A1(n14370), .A2(n14371), .ZN(n14375) );
  OR2_X1 U14336 ( .A1(n8026), .A2(n8039), .ZN(n14371) );
  OR2_X1 U14337 ( .A1(n14376), .A2(n14377), .ZN(n14370) );
  AND2_X1 U14338 ( .A1(n14367), .A2(n14366), .ZN(n14377) );
  AND2_X1 U14339 ( .A1(n14364), .A2(n14378), .ZN(n14376) );
  OR2_X1 U14340 ( .A1(n14366), .A2(n14367), .ZN(n14378) );
  OR2_X1 U14341 ( .A1(n8026), .A2(n8043), .ZN(n14367) );
  OR2_X1 U14342 ( .A1(n14379), .A2(n14380), .ZN(n14366) );
  AND2_X1 U14343 ( .A1(n14363), .A2(n14362), .ZN(n14380) );
  AND2_X1 U14344 ( .A1(n14360), .A2(n14381), .ZN(n14379) );
  OR2_X1 U14345 ( .A1(n14362), .A2(n14363), .ZN(n14381) );
  OR2_X1 U14346 ( .A1(n8026), .A2(n8048), .ZN(n14363) );
  OR2_X1 U14347 ( .A1(n14382), .A2(n14383), .ZN(n14362) );
  AND2_X1 U14348 ( .A1(n14359), .A2(n14358), .ZN(n14383) );
  AND2_X1 U14349 ( .A1(n14356), .A2(n14384), .ZN(n14382) );
  OR2_X1 U14350 ( .A1(n14358), .A2(n14359), .ZN(n14384) );
  OR2_X1 U14351 ( .A1(n8026), .A2(n8052), .ZN(n14359) );
  OR2_X1 U14352 ( .A1(n14385), .A2(n14386), .ZN(n14358) );
  AND2_X1 U14353 ( .A1(n14355), .A2(n14354), .ZN(n14386) );
  AND2_X1 U14354 ( .A1(n14352), .A2(n14387), .ZN(n14385) );
  OR2_X1 U14355 ( .A1(n14354), .A2(n14355), .ZN(n14387) );
  OR2_X1 U14356 ( .A1(n8026), .A2(n8057), .ZN(n14355) );
  OR2_X1 U14357 ( .A1(n14388), .A2(n14389), .ZN(n14354) );
  AND2_X1 U14358 ( .A1(n14351), .A2(n14350), .ZN(n14389) );
  AND2_X1 U14359 ( .A1(n14348), .A2(n14390), .ZN(n14388) );
  OR2_X1 U14360 ( .A1(n14350), .A2(n14351), .ZN(n14390) );
  OR2_X1 U14361 ( .A1(n8026), .A2(n8061), .ZN(n14351) );
  OR2_X1 U14362 ( .A1(n14391), .A2(n14392), .ZN(n14350) );
  AND2_X1 U14363 ( .A1(n14347), .A2(n14346), .ZN(n14392) );
  AND2_X1 U14364 ( .A1(n14344), .A2(n14393), .ZN(n14391) );
  OR2_X1 U14365 ( .A1(n14346), .A2(n14347), .ZN(n14393) );
  OR2_X1 U14366 ( .A1(n8026), .A2(n8066), .ZN(n14347) );
  OR2_X1 U14367 ( .A1(n14394), .A2(n14395), .ZN(n14346) );
  AND2_X1 U14368 ( .A1(n14343), .A2(n14342), .ZN(n14395) );
  AND2_X1 U14369 ( .A1(n14340), .A2(n14396), .ZN(n14394) );
  OR2_X1 U14370 ( .A1(n14342), .A2(n14343), .ZN(n14396) );
  OR2_X1 U14371 ( .A1(n8026), .A2(n8070), .ZN(n14343) );
  OR2_X1 U14372 ( .A1(n14397), .A2(n14398), .ZN(n14342) );
  AND2_X1 U14373 ( .A1(n14339), .A2(n14338), .ZN(n14398) );
  AND2_X1 U14374 ( .A1(n14336), .A2(n14399), .ZN(n14397) );
  OR2_X1 U14375 ( .A1(n14338), .A2(n14339), .ZN(n14399) );
  OR2_X1 U14376 ( .A1(n8026), .A2(n8075), .ZN(n14339) );
  OR2_X1 U14377 ( .A1(n14400), .A2(n14401), .ZN(n14338) );
  AND2_X1 U14378 ( .A1(n14335), .A2(n14334), .ZN(n14401) );
  AND2_X1 U14379 ( .A1(n14332), .A2(n14402), .ZN(n14400) );
  OR2_X1 U14380 ( .A1(n14334), .A2(n14335), .ZN(n14402) );
  OR2_X1 U14381 ( .A1(n8026), .A2(n8079), .ZN(n14335) );
  OR2_X1 U14382 ( .A1(n14403), .A2(n14404), .ZN(n14334) );
  AND2_X1 U14383 ( .A1(n14331), .A2(n14330), .ZN(n14404) );
  AND2_X1 U14384 ( .A1(n14328), .A2(n14405), .ZN(n14403) );
  OR2_X1 U14385 ( .A1(n14330), .A2(n14331), .ZN(n14405) );
  OR2_X1 U14386 ( .A1(n8026), .A2(n8084), .ZN(n14331) );
  OR2_X1 U14387 ( .A1(n14406), .A2(n14407), .ZN(n14330) );
  AND2_X1 U14388 ( .A1(n14327), .A2(n14326), .ZN(n14407) );
  AND2_X1 U14389 ( .A1(n14324), .A2(n14408), .ZN(n14406) );
  OR2_X1 U14390 ( .A1(n14326), .A2(n14327), .ZN(n14408) );
  OR2_X1 U14391 ( .A1(n8026), .A2(n8088), .ZN(n14327) );
  OR2_X1 U14392 ( .A1(n14409), .A2(n14410), .ZN(n14326) );
  AND2_X1 U14393 ( .A1(n14323), .A2(n14322), .ZN(n14410) );
  AND2_X1 U14394 ( .A1(n14320), .A2(n14411), .ZN(n14409) );
  OR2_X1 U14395 ( .A1(n14322), .A2(n14323), .ZN(n14411) );
  OR2_X1 U14396 ( .A1(n8026), .A2(n8093), .ZN(n14323) );
  OR2_X1 U14397 ( .A1(n14412), .A2(n14413), .ZN(n14322) );
  AND2_X1 U14398 ( .A1(n14319), .A2(n14318), .ZN(n14413) );
  AND2_X1 U14399 ( .A1(n14316), .A2(n14414), .ZN(n14412) );
  OR2_X1 U14400 ( .A1(n14318), .A2(n14319), .ZN(n14414) );
  OR2_X1 U14401 ( .A1(n8026), .A2(n8097), .ZN(n14319) );
  OR2_X1 U14402 ( .A1(n14415), .A2(n14416), .ZN(n14318) );
  AND2_X1 U14403 ( .A1(n14315), .A2(n14314), .ZN(n14416) );
  AND2_X1 U14404 ( .A1(n14312), .A2(n14417), .ZN(n14415) );
  OR2_X1 U14405 ( .A1(n14314), .A2(n14315), .ZN(n14417) );
  OR2_X1 U14406 ( .A1(n8026), .A2(n8102), .ZN(n14315) );
  OR2_X1 U14407 ( .A1(n14418), .A2(n14419), .ZN(n14314) );
  AND2_X1 U14408 ( .A1(n14311), .A2(n14310), .ZN(n14419) );
  AND2_X1 U14409 ( .A1(n14308), .A2(n14420), .ZN(n14418) );
  OR2_X1 U14410 ( .A1(n14310), .A2(n14311), .ZN(n14420) );
  OR2_X1 U14411 ( .A1(n8026), .A2(n8106), .ZN(n14311) );
  OR2_X1 U14412 ( .A1(n14421), .A2(n14422), .ZN(n14310) );
  AND2_X1 U14413 ( .A1(n14307), .A2(n14306), .ZN(n14422) );
  AND2_X1 U14414 ( .A1(n14304), .A2(n14423), .ZN(n14421) );
  OR2_X1 U14415 ( .A1(n14306), .A2(n14307), .ZN(n14423) );
  OR2_X1 U14416 ( .A1(n8026), .A2(n8109), .ZN(n14307) );
  OR2_X1 U14417 ( .A1(n14424), .A2(n14425), .ZN(n14306) );
  AND2_X1 U14418 ( .A1(n14303), .A2(n14302), .ZN(n14425) );
  AND2_X1 U14419 ( .A1(n14300), .A2(n14426), .ZN(n14424) );
  OR2_X1 U14420 ( .A1(n14302), .A2(n14303), .ZN(n14426) );
  OR2_X1 U14421 ( .A1(n8026), .A2(n8112), .ZN(n14303) );
  OR2_X1 U14422 ( .A1(n14427), .A2(n14428), .ZN(n14302) );
  AND2_X1 U14423 ( .A1(n14296), .A2(n14299), .ZN(n14428) );
  AND2_X1 U14424 ( .A1(n14429), .A2(n14298), .ZN(n14427) );
  OR2_X1 U14425 ( .A1(n14430), .A2(n14431), .ZN(n14298) );
  AND2_X1 U14426 ( .A1(n14295), .A2(n14294), .ZN(n14431) );
  AND2_X1 U14427 ( .A1(n14292), .A2(n14432), .ZN(n14430) );
  OR2_X1 U14428 ( .A1(n14294), .A2(n14295), .ZN(n14432) );
  OR2_X1 U14429 ( .A1(n8026), .A2(n8118), .ZN(n14295) );
  OR2_X1 U14430 ( .A1(n14433), .A2(n14434), .ZN(n14294) );
  AND2_X1 U14431 ( .A1(n14288), .A2(n14291), .ZN(n14434) );
  AND2_X1 U14432 ( .A1(n14435), .A2(n14290), .ZN(n14433) );
  OR2_X1 U14433 ( .A1(n14436), .A2(n14437), .ZN(n14290) );
  AND2_X1 U14434 ( .A1(n14284), .A2(n14287), .ZN(n14437) );
  AND2_X1 U14435 ( .A1(n14438), .A2(n14286), .ZN(n14436) );
  OR2_X1 U14436 ( .A1(n14439), .A2(n14440), .ZN(n14286) );
  AND2_X1 U14437 ( .A1(n14280), .A2(n14283), .ZN(n14440) );
  AND2_X1 U14438 ( .A1(n14441), .A2(n14442), .ZN(n14439) );
  OR2_X1 U14439 ( .A1(n14283), .A2(n14280), .ZN(n14442) );
  OR2_X1 U14440 ( .A1(n8026), .A2(n8127), .ZN(n14280) );
  OR3_X1 U14441 ( .A1(n8022), .A2(n8026), .A3(n8981), .ZN(n14283) );
  INV_X1 U14442 ( .A(n14282), .ZN(n14441) );
  OR2_X1 U14443 ( .A1(n14443), .A2(n14444), .ZN(n14282) );
  AND2_X1 U14444 ( .A1(b_3_), .A2(n14445), .ZN(n14444) );
  OR2_X1 U14445 ( .A1(n14446), .A2(n7598), .ZN(n14445) );
  AND2_X1 U14446 ( .A1(a_30_), .A2(n8017), .ZN(n14446) );
  AND2_X1 U14447 ( .A1(b_2_), .A2(n14447), .ZN(n14443) );
  OR2_X1 U14448 ( .A1(n14448), .A2(n7601), .ZN(n14447) );
  AND2_X1 U14449 ( .A1(a_31_), .A2(n8022), .ZN(n14448) );
  OR2_X1 U14450 ( .A1(n14287), .A2(n14284), .ZN(n14438) );
  XNOR2_X1 U14451 ( .A(n14449), .B(n14450), .ZN(n14284) );
  XOR2_X1 U14452 ( .A(n14451), .B(n14452), .Z(n14450) );
  OR2_X1 U14453 ( .A1(n8026), .A2(n8124), .ZN(n14287) );
  OR2_X1 U14454 ( .A1(n14291), .A2(n14288), .ZN(n14435) );
  XOR2_X1 U14455 ( .A(n14453), .B(n14454), .Z(n14288) );
  XOR2_X1 U14456 ( .A(n14455), .B(n14456), .Z(n14454) );
  OR2_X1 U14457 ( .A1(n8026), .A2(n8121), .ZN(n14291) );
  XOR2_X1 U14458 ( .A(n14457), .B(n14458), .Z(n14292) );
  XOR2_X1 U14459 ( .A(n14459), .B(n14460), .Z(n14458) );
  OR2_X1 U14460 ( .A1(n14299), .A2(n14296), .ZN(n14429) );
  XOR2_X1 U14461 ( .A(n14461), .B(n14462), .Z(n14296) );
  XOR2_X1 U14462 ( .A(n14463), .B(n14464), .Z(n14462) );
  OR2_X1 U14463 ( .A1(n8026), .A2(n8115), .ZN(n14299) );
  INV_X1 U14464 ( .A(b_4_), .ZN(n8026) );
  XOR2_X1 U14465 ( .A(n14465), .B(n14466), .Z(n14300) );
  XOR2_X1 U14466 ( .A(n14467), .B(n14468), .Z(n14466) );
  XOR2_X1 U14467 ( .A(n14469), .B(n14470), .Z(n14304) );
  XOR2_X1 U14468 ( .A(n14471), .B(n14472), .Z(n14470) );
  XOR2_X1 U14469 ( .A(n14473), .B(n14474), .Z(n14308) );
  XOR2_X1 U14470 ( .A(n14475), .B(n14476), .Z(n14474) );
  XOR2_X1 U14471 ( .A(n14477), .B(n14478), .Z(n14312) );
  XOR2_X1 U14472 ( .A(n14479), .B(n14480), .Z(n14478) );
  XOR2_X1 U14473 ( .A(n14481), .B(n14482), .Z(n14316) );
  XOR2_X1 U14474 ( .A(n14483), .B(n14484), .Z(n14482) );
  XOR2_X1 U14475 ( .A(n14485), .B(n14486), .Z(n14320) );
  XOR2_X1 U14476 ( .A(n14487), .B(n14488), .Z(n14486) );
  XOR2_X1 U14477 ( .A(n14489), .B(n14490), .Z(n14324) );
  XOR2_X1 U14478 ( .A(n14491), .B(n14492), .Z(n14490) );
  XOR2_X1 U14479 ( .A(n14493), .B(n14494), .Z(n14328) );
  XOR2_X1 U14480 ( .A(n14495), .B(n14496), .Z(n14494) );
  XOR2_X1 U14481 ( .A(n14497), .B(n14498), .Z(n14332) );
  XOR2_X1 U14482 ( .A(n14499), .B(n14500), .Z(n14498) );
  XOR2_X1 U14483 ( .A(n14501), .B(n14502), .Z(n14336) );
  XOR2_X1 U14484 ( .A(n14503), .B(n14504), .Z(n14502) );
  XOR2_X1 U14485 ( .A(n14505), .B(n14506), .Z(n14340) );
  XOR2_X1 U14486 ( .A(n14507), .B(n14508), .Z(n14506) );
  XOR2_X1 U14487 ( .A(n14509), .B(n14510), .Z(n14344) );
  XOR2_X1 U14488 ( .A(n14511), .B(n14512), .Z(n14510) );
  XOR2_X1 U14489 ( .A(n14513), .B(n14514), .Z(n14348) );
  XOR2_X1 U14490 ( .A(n14515), .B(n14516), .Z(n14514) );
  XOR2_X1 U14491 ( .A(n14517), .B(n14518), .Z(n14352) );
  XOR2_X1 U14492 ( .A(n14519), .B(n14520), .Z(n14518) );
  XOR2_X1 U14493 ( .A(n14521), .B(n14522), .Z(n14356) );
  XOR2_X1 U14494 ( .A(n14523), .B(n14524), .Z(n14522) );
  XOR2_X1 U14495 ( .A(n14525), .B(n14526), .Z(n14360) );
  XOR2_X1 U14496 ( .A(n14527), .B(n14528), .Z(n14526) );
  XOR2_X1 U14497 ( .A(n14529), .B(n14530), .Z(n14364) );
  XOR2_X1 U14498 ( .A(n14531), .B(n14532), .Z(n14530) );
  XOR2_X1 U14499 ( .A(n14533), .B(n14534), .Z(n14368) );
  XOR2_X1 U14500 ( .A(n14535), .B(n14536), .Z(n14534) );
  XOR2_X1 U14501 ( .A(n8574), .B(n14537), .Z(n8567) );
  XOR2_X1 U14502 ( .A(n8573), .B(n8572), .Z(n14537) );
  OR2_X1 U14503 ( .A1(n8022), .A2(n8039), .ZN(n8572) );
  OR2_X1 U14504 ( .A1(n14538), .A2(n14539), .ZN(n8573) );
  AND2_X1 U14505 ( .A1(n14536), .A2(n14535), .ZN(n14539) );
  AND2_X1 U14506 ( .A1(n14533), .A2(n14540), .ZN(n14538) );
  OR2_X1 U14507 ( .A1(n14535), .A2(n14536), .ZN(n14540) );
  OR2_X1 U14508 ( .A1(n8022), .A2(n8043), .ZN(n14536) );
  OR2_X1 U14509 ( .A1(n14541), .A2(n14542), .ZN(n14535) );
  AND2_X1 U14510 ( .A1(n14532), .A2(n14531), .ZN(n14542) );
  AND2_X1 U14511 ( .A1(n14529), .A2(n14543), .ZN(n14541) );
  OR2_X1 U14512 ( .A1(n14531), .A2(n14532), .ZN(n14543) );
  OR2_X1 U14513 ( .A1(n8022), .A2(n8048), .ZN(n14532) );
  OR2_X1 U14514 ( .A1(n14544), .A2(n14545), .ZN(n14531) );
  AND2_X1 U14515 ( .A1(n14528), .A2(n14527), .ZN(n14545) );
  AND2_X1 U14516 ( .A1(n14525), .A2(n14546), .ZN(n14544) );
  OR2_X1 U14517 ( .A1(n14527), .A2(n14528), .ZN(n14546) );
  OR2_X1 U14518 ( .A1(n8022), .A2(n8052), .ZN(n14528) );
  OR2_X1 U14519 ( .A1(n14547), .A2(n14548), .ZN(n14527) );
  AND2_X1 U14520 ( .A1(n14524), .A2(n14523), .ZN(n14548) );
  AND2_X1 U14521 ( .A1(n14521), .A2(n14549), .ZN(n14547) );
  OR2_X1 U14522 ( .A1(n14523), .A2(n14524), .ZN(n14549) );
  OR2_X1 U14523 ( .A1(n8022), .A2(n8057), .ZN(n14524) );
  OR2_X1 U14524 ( .A1(n14550), .A2(n14551), .ZN(n14523) );
  AND2_X1 U14525 ( .A1(n14520), .A2(n14519), .ZN(n14551) );
  AND2_X1 U14526 ( .A1(n14517), .A2(n14552), .ZN(n14550) );
  OR2_X1 U14527 ( .A1(n14519), .A2(n14520), .ZN(n14552) );
  OR2_X1 U14528 ( .A1(n8022), .A2(n8061), .ZN(n14520) );
  OR2_X1 U14529 ( .A1(n14553), .A2(n14554), .ZN(n14519) );
  AND2_X1 U14530 ( .A1(n14516), .A2(n14515), .ZN(n14554) );
  AND2_X1 U14531 ( .A1(n14513), .A2(n14555), .ZN(n14553) );
  OR2_X1 U14532 ( .A1(n14515), .A2(n14516), .ZN(n14555) );
  OR2_X1 U14533 ( .A1(n8022), .A2(n8066), .ZN(n14516) );
  OR2_X1 U14534 ( .A1(n14556), .A2(n14557), .ZN(n14515) );
  AND2_X1 U14535 ( .A1(n14512), .A2(n14511), .ZN(n14557) );
  AND2_X1 U14536 ( .A1(n14509), .A2(n14558), .ZN(n14556) );
  OR2_X1 U14537 ( .A1(n14511), .A2(n14512), .ZN(n14558) );
  OR2_X1 U14538 ( .A1(n8022), .A2(n8070), .ZN(n14512) );
  OR2_X1 U14539 ( .A1(n14559), .A2(n14560), .ZN(n14511) );
  AND2_X1 U14540 ( .A1(n14508), .A2(n14507), .ZN(n14560) );
  AND2_X1 U14541 ( .A1(n14505), .A2(n14561), .ZN(n14559) );
  OR2_X1 U14542 ( .A1(n14507), .A2(n14508), .ZN(n14561) );
  OR2_X1 U14543 ( .A1(n8022), .A2(n8075), .ZN(n14508) );
  OR2_X1 U14544 ( .A1(n14562), .A2(n14563), .ZN(n14507) );
  AND2_X1 U14545 ( .A1(n14504), .A2(n14503), .ZN(n14563) );
  AND2_X1 U14546 ( .A1(n14501), .A2(n14564), .ZN(n14562) );
  OR2_X1 U14547 ( .A1(n14503), .A2(n14504), .ZN(n14564) );
  OR2_X1 U14548 ( .A1(n8022), .A2(n8079), .ZN(n14504) );
  OR2_X1 U14549 ( .A1(n14565), .A2(n14566), .ZN(n14503) );
  AND2_X1 U14550 ( .A1(n14500), .A2(n14499), .ZN(n14566) );
  AND2_X1 U14551 ( .A1(n14497), .A2(n14567), .ZN(n14565) );
  OR2_X1 U14552 ( .A1(n14499), .A2(n14500), .ZN(n14567) );
  OR2_X1 U14553 ( .A1(n8022), .A2(n8084), .ZN(n14500) );
  OR2_X1 U14554 ( .A1(n14568), .A2(n14569), .ZN(n14499) );
  AND2_X1 U14555 ( .A1(n14496), .A2(n14495), .ZN(n14569) );
  AND2_X1 U14556 ( .A1(n14493), .A2(n14570), .ZN(n14568) );
  OR2_X1 U14557 ( .A1(n14495), .A2(n14496), .ZN(n14570) );
  OR2_X1 U14558 ( .A1(n8022), .A2(n8088), .ZN(n14496) );
  OR2_X1 U14559 ( .A1(n14571), .A2(n14572), .ZN(n14495) );
  AND2_X1 U14560 ( .A1(n14492), .A2(n14491), .ZN(n14572) );
  AND2_X1 U14561 ( .A1(n14489), .A2(n14573), .ZN(n14571) );
  OR2_X1 U14562 ( .A1(n14491), .A2(n14492), .ZN(n14573) );
  OR2_X1 U14563 ( .A1(n8022), .A2(n8093), .ZN(n14492) );
  OR2_X1 U14564 ( .A1(n14574), .A2(n14575), .ZN(n14491) );
  AND2_X1 U14565 ( .A1(n14488), .A2(n14487), .ZN(n14575) );
  AND2_X1 U14566 ( .A1(n14485), .A2(n14576), .ZN(n14574) );
  OR2_X1 U14567 ( .A1(n14487), .A2(n14488), .ZN(n14576) );
  OR2_X1 U14568 ( .A1(n8022), .A2(n8097), .ZN(n14488) );
  OR2_X1 U14569 ( .A1(n14577), .A2(n14578), .ZN(n14487) );
  AND2_X1 U14570 ( .A1(n14484), .A2(n14483), .ZN(n14578) );
  AND2_X1 U14571 ( .A1(n14481), .A2(n14579), .ZN(n14577) );
  OR2_X1 U14572 ( .A1(n14483), .A2(n14484), .ZN(n14579) );
  OR2_X1 U14573 ( .A1(n8022), .A2(n8102), .ZN(n14484) );
  OR2_X1 U14574 ( .A1(n14580), .A2(n14581), .ZN(n14483) );
  AND2_X1 U14575 ( .A1(n14480), .A2(n14479), .ZN(n14581) );
  AND2_X1 U14576 ( .A1(n14477), .A2(n14582), .ZN(n14580) );
  OR2_X1 U14577 ( .A1(n14479), .A2(n14480), .ZN(n14582) );
  OR2_X1 U14578 ( .A1(n8022), .A2(n8106), .ZN(n14480) );
  OR2_X1 U14579 ( .A1(n14583), .A2(n14584), .ZN(n14479) );
  AND2_X1 U14580 ( .A1(n14476), .A2(n14475), .ZN(n14584) );
  AND2_X1 U14581 ( .A1(n14473), .A2(n14585), .ZN(n14583) );
  OR2_X1 U14582 ( .A1(n14475), .A2(n14476), .ZN(n14585) );
  OR2_X1 U14583 ( .A1(n8022), .A2(n8109), .ZN(n14476) );
  OR2_X1 U14584 ( .A1(n14586), .A2(n14587), .ZN(n14475) );
  AND2_X1 U14585 ( .A1(n14472), .A2(n14471), .ZN(n14587) );
  AND2_X1 U14586 ( .A1(n14469), .A2(n14588), .ZN(n14586) );
  OR2_X1 U14587 ( .A1(n14471), .A2(n14472), .ZN(n14588) );
  OR2_X1 U14588 ( .A1(n8022), .A2(n8112), .ZN(n14472) );
  OR2_X1 U14589 ( .A1(n14589), .A2(n14590), .ZN(n14471) );
  AND2_X1 U14590 ( .A1(n14468), .A2(n14467), .ZN(n14590) );
  AND2_X1 U14591 ( .A1(n14465), .A2(n14591), .ZN(n14589) );
  OR2_X1 U14592 ( .A1(n14467), .A2(n14468), .ZN(n14591) );
  OR2_X1 U14593 ( .A1(n8022), .A2(n8115), .ZN(n14468) );
  OR2_X1 U14594 ( .A1(n14592), .A2(n14593), .ZN(n14467) );
  AND2_X1 U14595 ( .A1(n14461), .A2(n14464), .ZN(n14593) );
  AND2_X1 U14596 ( .A1(n14594), .A2(n14463), .ZN(n14592) );
  OR2_X1 U14597 ( .A1(n14595), .A2(n14596), .ZN(n14463) );
  AND2_X1 U14598 ( .A1(n14460), .A2(n14459), .ZN(n14596) );
  AND2_X1 U14599 ( .A1(n14457), .A2(n14597), .ZN(n14595) );
  OR2_X1 U14600 ( .A1(n14459), .A2(n14460), .ZN(n14597) );
  OR2_X1 U14601 ( .A1(n8022), .A2(n8121), .ZN(n14460) );
  OR2_X1 U14602 ( .A1(n14598), .A2(n14599), .ZN(n14459) );
  AND2_X1 U14603 ( .A1(n14453), .A2(n14456), .ZN(n14599) );
  AND2_X1 U14604 ( .A1(n14600), .A2(n14455), .ZN(n14598) );
  OR2_X1 U14605 ( .A1(n14601), .A2(n14602), .ZN(n14455) );
  AND2_X1 U14606 ( .A1(n14449), .A2(n14452), .ZN(n14602) );
  AND2_X1 U14607 ( .A1(n14603), .A2(n14604), .ZN(n14601) );
  OR2_X1 U14608 ( .A1(n14452), .A2(n14449), .ZN(n14604) );
  OR2_X1 U14609 ( .A1(n8022), .A2(n8127), .ZN(n14449) );
  OR3_X1 U14610 ( .A1(n8022), .A2(n8981), .A3(n8017), .ZN(n14452) );
  INV_X1 U14611 ( .A(n14451), .ZN(n14603) );
  OR2_X1 U14612 ( .A1(n14605), .A2(n14606), .ZN(n14451) );
  AND2_X1 U14613 ( .A1(b_2_), .A2(n14607), .ZN(n14606) );
  OR2_X1 U14614 ( .A1(n14608), .A2(n7598), .ZN(n14607) );
  AND2_X1 U14615 ( .A1(a_30_), .A2(n8013), .ZN(n14608) );
  AND2_X1 U14616 ( .A1(b_1_), .A2(n14609), .ZN(n14605) );
  OR2_X1 U14617 ( .A1(n14610), .A2(n7601), .ZN(n14609) );
  AND2_X1 U14618 ( .A1(a_31_), .A2(n8017), .ZN(n14610) );
  OR2_X1 U14619 ( .A1(n14456), .A2(n14453), .ZN(n14600) );
  XNOR2_X1 U14620 ( .A(n14611), .B(n14612), .ZN(n14453) );
  XOR2_X1 U14621 ( .A(n14613), .B(n14614), .Z(n14612) );
  OR2_X1 U14622 ( .A1(n8022), .A2(n8124), .ZN(n14456) );
  XOR2_X1 U14623 ( .A(n14615), .B(n14616), .Z(n14457) );
  XOR2_X1 U14624 ( .A(n14617), .B(n14618), .Z(n14616) );
  OR2_X1 U14625 ( .A1(n14464), .A2(n14461), .ZN(n14594) );
  XOR2_X1 U14626 ( .A(n14619), .B(n14620), .Z(n14461) );
  XOR2_X1 U14627 ( .A(n14621), .B(n14622), .Z(n14620) );
  OR2_X1 U14628 ( .A1(n8022), .A2(n8118), .ZN(n14464) );
  XOR2_X1 U14629 ( .A(n14623), .B(n14624), .Z(n14465) );
  XOR2_X1 U14630 ( .A(n14625), .B(n14626), .Z(n14624) );
  XOR2_X1 U14631 ( .A(n14627), .B(n14628), .Z(n14469) );
  XOR2_X1 U14632 ( .A(n14629), .B(n14630), .Z(n14628) );
  XOR2_X1 U14633 ( .A(n14631), .B(n14632), .Z(n14473) );
  XOR2_X1 U14634 ( .A(n14633), .B(n14634), .Z(n14632) );
  XOR2_X1 U14635 ( .A(n14635), .B(n14636), .Z(n14477) );
  XOR2_X1 U14636 ( .A(n14637), .B(n14638), .Z(n14636) );
  XOR2_X1 U14637 ( .A(n14639), .B(n14640), .Z(n14481) );
  XOR2_X1 U14638 ( .A(n14641), .B(n14642), .Z(n14640) );
  XOR2_X1 U14639 ( .A(n14643), .B(n14644), .Z(n14485) );
  XOR2_X1 U14640 ( .A(n14645), .B(n14646), .Z(n14644) );
  XOR2_X1 U14641 ( .A(n14647), .B(n14648), .Z(n14489) );
  XOR2_X1 U14642 ( .A(n14649), .B(n14650), .Z(n14648) );
  XOR2_X1 U14643 ( .A(n14651), .B(n14652), .Z(n14493) );
  XOR2_X1 U14644 ( .A(n14653), .B(n14654), .Z(n14652) );
  XOR2_X1 U14645 ( .A(n14655), .B(n14656), .Z(n14497) );
  XOR2_X1 U14646 ( .A(n14657), .B(n14658), .Z(n14656) );
  XOR2_X1 U14647 ( .A(n14659), .B(n14660), .Z(n14501) );
  XOR2_X1 U14648 ( .A(n14661), .B(n14662), .Z(n14660) );
  XOR2_X1 U14649 ( .A(n14663), .B(n14664), .Z(n14505) );
  XOR2_X1 U14650 ( .A(n14665), .B(n14666), .Z(n14664) );
  XOR2_X1 U14651 ( .A(n14667), .B(n14668), .Z(n14509) );
  XOR2_X1 U14652 ( .A(n14669), .B(n14670), .Z(n14668) );
  XOR2_X1 U14653 ( .A(n14671), .B(n14672), .Z(n14513) );
  XOR2_X1 U14654 ( .A(n14673), .B(n14674), .Z(n14672) );
  XOR2_X1 U14655 ( .A(n14675), .B(n14676), .Z(n14517) );
  XOR2_X1 U14656 ( .A(n14677), .B(n14678), .Z(n14676) );
  XOR2_X1 U14657 ( .A(n14679), .B(n14680), .Z(n14521) );
  XOR2_X1 U14658 ( .A(n14681), .B(n14682), .Z(n14680) );
  XOR2_X1 U14659 ( .A(n14683), .B(n14684), .Z(n14525) );
  XOR2_X1 U14660 ( .A(n14685), .B(n14686), .Z(n14684) );
  XOR2_X1 U14661 ( .A(n14687), .B(n14688), .Z(n14529) );
  XOR2_X1 U14662 ( .A(n14689), .B(n14690), .Z(n14688) );
  XOR2_X1 U14663 ( .A(n14691), .B(n14692), .Z(n14533) );
  XOR2_X1 U14664 ( .A(n14693), .B(n14694), .Z(n14692) );
  XOR2_X1 U14665 ( .A(n14695), .B(n14696), .Z(n8574) );
  XOR2_X1 U14666 ( .A(n14697), .B(n14698), .Z(n14696) );
  AND2_X1 U14667 ( .A1(n14699), .A2(b_0_), .ZN(n8269) );
  INV_X1 U14668 ( .A(n14700), .ZN(n14699) );
  AND3_X1 U14669 ( .A1(n8205), .A2(n8204), .A3(n8202), .ZN(n8206) );
  AND2_X1 U14670 ( .A1(n14700), .A2(b_0_), .ZN(n8202) );
  OR3_X1 U14671 ( .A1(n14701), .A2(n14702), .A3(n14703), .ZN(n8204) );
  XNOR2_X1 U14672 ( .A(n14700), .B(n14704), .ZN(n14703) );
  AND2_X1 U14673 ( .A1(b_0_), .A2(a_1_), .ZN(n14704) );
  OR2_X1 U14674 ( .A1(n8013), .A2(n8297), .ZN(n14700) );
  OR2_X1 U14675 ( .A1(n14705), .A2(n14706), .ZN(n8205) );
  AND2_X1 U14676 ( .A1(n8288), .A2(n8285), .ZN(n14706) );
  XNOR2_X1 U14677 ( .A(n14707), .B(n14702), .ZN(n8285) );
  INV_X1 U14678 ( .A(n14708), .ZN(n14702) );
  OR2_X1 U14679 ( .A1(n14709), .A2(n14710), .ZN(n14708) );
  AND2_X1 U14680 ( .A1(n14711), .A2(n14712), .ZN(n14710) );
  AND2_X1 U14681 ( .A1(n14713), .A2(n14714), .ZN(n14709) );
  OR2_X1 U14682 ( .A1(n14712), .A2(n14711), .ZN(n14713) );
  OR2_X1 U14683 ( .A1(n14715), .A2(n14701), .ZN(n14707) );
  AND3_X1 U14684 ( .A1(a_2_), .A2(b_0_), .A3(n14716), .ZN(n14701) );
  INV_X1 U14685 ( .A(n8014), .ZN(n14716) );
  AND2_X1 U14686 ( .A1(n14717), .A2(n8014), .ZN(n14715) );
  OR2_X1 U14687 ( .A1(n8013), .A2(n8012), .ZN(n8014) );
  OR2_X1 U14688 ( .A1(n8016), .A2(n14718), .ZN(n14717) );
  AND2_X1 U14689 ( .A1(b_2_), .A2(a_0_), .ZN(n8288) );
  INV_X1 U14690 ( .A(n8287), .ZN(n14705) );
  OR2_X1 U14691 ( .A1(n14719), .A2(n14720), .ZN(n8287) );
  AND2_X1 U14692 ( .A1(n8307), .A2(n8306), .ZN(n14720) );
  AND2_X1 U14693 ( .A1(n8304), .A2(n14721), .ZN(n14719) );
  OR2_X1 U14694 ( .A1(n8306), .A2(n8307), .ZN(n14721) );
  OR2_X1 U14695 ( .A1(n8017), .A2(n8012), .ZN(n8307) );
  OR2_X1 U14696 ( .A1(n14722), .A2(n14723), .ZN(n8306) );
  AND2_X1 U14697 ( .A1(n8338), .A2(n8018), .ZN(n14723) );
  AND2_X1 U14698 ( .A1(n8337), .A2(n14724), .ZN(n14722) );
  OR2_X1 U14699 ( .A1(n8018), .A2(n8338), .ZN(n14724) );
  OR2_X1 U14700 ( .A1(n14725), .A2(n14726), .ZN(n8338) );
  AND2_X1 U14701 ( .A1(n8369), .A2(n8368), .ZN(n14726) );
  AND2_X1 U14702 ( .A1(n8366), .A2(n14727), .ZN(n14725) );
  OR2_X1 U14703 ( .A1(n8368), .A2(n8369), .ZN(n14727) );
  OR2_X1 U14704 ( .A1(n8021), .A2(n8017), .ZN(n8369) );
  OR2_X1 U14705 ( .A1(n14728), .A2(n14729), .ZN(n8368) );
  AND2_X1 U14706 ( .A1(n8415), .A2(n8414), .ZN(n14729) );
  AND2_X1 U14707 ( .A1(n8412), .A2(n14730), .ZN(n14728) );
  OR2_X1 U14708 ( .A1(n8414), .A2(n8415), .ZN(n14730) );
  OR2_X1 U14709 ( .A1(n8025), .A2(n8017), .ZN(n8415) );
  OR2_X1 U14710 ( .A1(n14731), .A2(n14732), .ZN(n8414) );
  AND2_X1 U14711 ( .A1(n8460), .A2(n8459), .ZN(n14732) );
  AND2_X1 U14712 ( .A1(n8457), .A2(n14733), .ZN(n14731) );
  OR2_X1 U14713 ( .A1(n8459), .A2(n8460), .ZN(n14733) );
  OR2_X1 U14714 ( .A1(n8030), .A2(n8017), .ZN(n8460) );
  OR2_X1 U14715 ( .A1(n14734), .A2(n14735), .ZN(n8459) );
  AND2_X1 U14716 ( .A1(n8514), .A2(n8513), .ZN(n14735) );
  AND2_X1 U14717 ( .A1(n8511), .A2(n14736), .ZN(n14734) );
  OR2_X1 U14718 ( .A1(n8513), .A2(n8514), .ZN(n14736) );
  OR2_X1 U14719 ( .A1(n8034), .A2(n8017), .ZN(n8514) );
  OR2_X1 U14720 ( .A1(n14737), .A2(n14738), .ZN(n8513) );
  AND2_X1 U14721 ( .A1(n8579), .A2(n8578), .ZN(n14738) );
  AND2_X1 U14722 ( .A1(n8576), .A2(n14739), .ZN(n14737) );
  OR2_X1 U14723 ( .A1(n8578), .A2(n8579), .ZN(n14739) );
  OR2_X1 U14724 ( .A1(n8039), .A2(n8017), .ZN(n8579) );
  OR2_X1 U14725 ( .A1(n14740), .A2(n14741), .ZN(n8578) );
  AND2_X1 U14726 ( .A1(n14698), .A2(n14697), .ZN(n14741) );
  AND2_X1 U14727 ( .A1(n14695), .A2(n14742), .ZN(n14740) );
  OR2_X1 U14728 ( .A1(n14697), .A2(n14698), .ZN(n14742) );
  OR2_X1 U14729 ( .A1(n8043), .A2(n8017), .ZN(n14698) );
  OR2_X1 U14730 ( .A1(n14743), .A2(n14744), .ZN(n14697) );
  AND2_X1 U14731 ( .A1(n14694), .A2(n14693), .ZN(n14744) );
  AND2_X1 U14732 ( .A1(n14691), .A2(n14745), .ZN(n14743) );
  OR2_X1 U14733 ( .A1(n14693), .A2(n14694), .ZN(n14745) );
  OR2_X1 U14734 ( .A1(n8048), .A2(n8017), .ZN(n14694) );
  OR2_X1 U14735 ( .A1(n14746), .A2(n14747), .ZN(n14693) );
  AND2_X1 U14736 ( .A1(n14690), .A2(n14689), .ZN(n14747) );
  AND2_X1 U14737 ( .A1(n14687), .A2(n14748), .ZN(n14746) );
  OR2_X1 U14738 ( .A1(n14689), .A2(n14690), .ZN(n14748) );
  OR2_X1 U14739 ( .A1(n8052), .A2(n8017), .ZN(n14690) );
  OR2_X1 U14740 ( .A1(n14749), .A2(n14750), .ZN(n14689) );
  AND2_X1 U14741 ( .A1(n14686), .A2(n14685), .ZN(n14750) );
  AND2_X1 U14742 ( .A1(n14683), .A2(n14751), .ZN(n14749) );
  OR2_X1 U14743 ( .A1(n14685), .A2(n14686), .ZN(n14751) );
  OR2_X1 U14744 ( .A1(n8057), .A2(n8017), .ZN(n14686) );
  OR2_X1 U14745 ( .A1(n14752), .A2(n14753), .ZN(n14685) );
  AND2_X1 U14746 ( .A1(n14682), .A2(n14681), .ZN(n14753) );
  AND2_X1 U14747 ( .A1(n14679), .A2(n14754), .ZN(n14752) );
  OR2_X1 U14748 ( .A1(n14681), .A2(n14682), .ZN(n14754) );
  OR2_X1 U14749 ( .A1(n8061), .A2(n8017), .ZN(n14682) );
  OR2_X1 U14750 ( .A1(n14755), .A2(n14756), .ZN(n14681) );
  AND2_X1 U14751 ( .A1(n14678), .A2(n14677), .ZN(n14756) );
  AND2_X1 U14752 ( .A1(n14675), .A2(n14757), .ZN(n14755) );
  OR2_X1 U14753 ( .A1(n14677), .A2(n14678), .ZN(n14757) );
  OR2_X1 U14754 ( .A1(n8066), .A2(n8017), .ZN(n14678) );
  OR2_X1 U14755 ( .A1(n14758), .A2(n14759), .ZN(n14677) );
  AND2_X1 U14756 ( .A1(n14674), .A2(n14673), .ZN(n14759) );
  AND2_X1 U14757 ( .A1(n14671), .A2(n14760), .ZN(n14758) );
  OR2_X1 U14758 ( .A1(n14673), .A2(n14674), .ZN(n14760) );
  OR2_X1 U14759 ( .A1(n8070), .A2(n8017), .ZN(n14674) );
  OR2_X1 U14760 ( .A1(n14761), .A2(n14762), .ZN(n14673) );
  AND2_X1 U14761 ( .A1(n14670), .A2(n14669), .ZN(n14762) );
  AND2_X1 U14762 ( .A1(n14667), .A2(n14763), .ZN(n14761) );
  OR2_X1 U14763 ( .A1(n14669), .A2(n14670), .ZN(n14763) );
  OR2_X1 U14764 ( .A1(n8075), .A2(n8017), .ZN(n14670) );
  OR2_X1 U14765 ( .A1(n14764), .A2(n14765), .ZN(n14669) );
  AND2_X1 U14766 ( .A1(n14666), .A2(n14665), .ZN(n14765) );
  AND2_X1 U14767 ( .A1(n14663), .A2(n14766), .ZN(n14764) );
  OR2_X1 U14768 ( .A1(n14665), .A2(n14666), .ZN(n14766) );
  OR2_X1 U14769 ( .A1(n8079), .A2(n8017), .ZN(n14666) );
  OR2_X1 U14770 ( .A1(n14767), .A2(n14768), .ZN(n14665) );
  AND2_X1 U14771 ( .A1(n14662), .A2(n14661), .ZN(n14768) );
  AND2_X1 U14772 ( .A1(n14659), .A2(n14769), .ZN(n14767) );
  OR2_X1 U14773 ( .A1(n14661), .A2(n14662), .ZN(n14769) );
  OR2_X1 U14774 ( .A1(n8084), .A2(n8017), .ZN(n14662) );
  OR2_X1 U14775 ( .A1(n14770), .A2(n14771), .ZN(n14661) );
  AND2_X1 U14776 ( .A1(n14658), .A2(n14657), .ZN(n14771) );
  AND2_X1 U14777 ( .A1(n14655), .A2(n14772), .ZN(n14770) );
  OR2_X1 U14778 ( .A1(n14657), .A2(n14658), .ZN(n14772) );
  OR2_X1 U14779 ( .A1(n8088), .A2(n8017), .ZN(n14658) );
  OR2_X1 U14780 ( .A1(n14773), .A2(n14774), .ZN(n14657) );
  AND2_X1 U14781 ( .A1(n14654), .A2(n14653), .ZN(n14774) );
  AND2_X1 U14782 ( .A1(n14651), .A2(n14775), .ZN(n14773) );
  OR2_X1 U14783 ( .A1(n14653), .A2(n14654), .ZN(n14775) );
  OR2_X1 U14784 ( .A1(n8093), .A2(n8017), .ZN(n14654) );
  OR2_X1 U14785 ( .A1(n14776), .A2(n14777), .ZN(n14653) );
  AND2_X1 U14786 ( .A1(n14650), .A2(n14649), .ZN(n14777) );
  AND2_X1 U14787 ( .A1(n14647), .A2(n14778), .ZN(n14776) );
  OR2_X1 U14788 ( .A1(n14649), .A2(n14650), .ZN(n14778) );
  OR2_X1 U14789 ( .A1(n8097), .A2(n8017), .ZN(n14650) );
  OR2_X1 U14790 ( .A1(n14779), .A2(n14780), .ZN(n14649) );
  AND2_X1 U14791 ( .A1(n14646), .A2(n14645), .ZN(n14780) );
  AND2_X1 U14792 ( .A1(n14643), .A2(n14781), .ZN(n14779) );
  OR2_X1 U14793 ( .A1(n14645), .A2(n14646), .ZN(n14781) );
  OR2_X1 U14794 ( .A1(n8102), .A2(n8017), .ZN(n14646) );
  OR2_X1 U14795 ( .A1(n14782), .A2(n14783), .ZN(n14645) );
  AND2_X1 U14796 ( .A1(n14642), .A2(n14641), .ZN(n14783) );
  AND2_X1 U14797 ( .A1(n14639), .A2(n14784), .ZN(n14782) );
  OR2_X1 U14798 ( .A1(n14641), .A2(n14642), .ZN(n14784) );
  OR2_X1 U14799 ( .A1(n8106), .A2(n8017), .ZN(n14642) );
  OR2_X1 U14800 ( .A1(n14785), .A2(n14786), .ZN(n14641) );
  AND2_X1 U14801 ( .A1(n14638), .A2(n14637), .ZN(n14786) );
  AND2_X1 U14802 ( .A1(n14635), .A2(n14787), .ZN(n14785) );
  OR2_X1 U14803 ( .A1(n14637), .A2(n14638), .ZN(n14787) );
  OR2_X1 U14804 ( .A1(n8109), .A2(n8017), .ZN(n14638) );
  OR2_X1 U14805 ( .A1(n14788), .A2(n14789), .ZN(n14637) );
  AND2_X1 U14806 ( .A1(n14634), .A2(n14633), .ZN(n14789) );
  AND2_X1 U14807 ( .A1(n14631), .A2(n14790), .ZN(n14788) );
  OR2_X1 U14808 ( .A1(n14633), .A2(n14634), .ZN(n14790) );
  OR2_X1 U14809 ( .A1(n8112), .A2(n8017), .ZN(n14634) );
  OR2_X1 U14810 ( .A1(n14791), .A2(n14792), .ZN(n14633) );
  AND2_X1 U14811 ( .A1(n14630), .A2(n14629), .ZN(n14792) );
  AND2_X1 U14812 ( .A1(n14627), .A2(n14793), .ZN(n14791) );
  OR2_X1 U14813 ( .A1(n14629), .A2(n14630), .ZN(n14793) );
  OR2_X1 U14814 ( .A1(n8115), .A2(n8017), .ZN(n14630) );
  OR2_X1 U14815 ( .A1(n14794), .A2(n14795), .ZN(n14629) );
  AND2_X1 U14816 ( .A1(n14626), .A2(n14625), .ZN(n14795) );
  AND2_X1 U14817 ( .A1(n14623), .A2(n14796), .ZN(n14794) );
  OR2_X1 U14818 ( .A1(n14625), .A2(n14626), .ZN(n14796) );
  OR2_X1 U14819 ( .A1(n8118), .A2(n8017), .ZN(n14626) );
  OR2_X1 U14820 ( .A1(n14797), .A2(n14798), .ZN(n14625) );
  AND2_X1 U14821 ( .A1(n14619), .A2(n14622), .ZN(n14798) );
  AND2_X1 U14822 ( .A1(n14799), .A2(n14621), .ZN(n14797) );
  OR2_X1 U14823 ( .A1(n14800), .A2(n14801), .ZN(n14621) );
  AND2_X1 U14824 ( .A1(n14618), .A2(n14617), .ZN(n14801) );
  AND2_X1 U14825 ( .A1(n14615), .A2(n14802), .ZN(n14800) );
  OR2_X1 U14826 ( .A1(n14617), .A2(n14618), .ZN(n14802) );
  OR2_X1 U14827 ( .A1(n8124), .A2(n8017), .ZN(n14618) );
  OR2_X1 U14828 ( .A1(n14803), .A2(n14804), .ZN(n14617) );
  AND2_X1 U14829 ( .A1(n14611), .A2(n14614), .ZN(n14804) );
  AND2_X1 U14830 ( .A1(n14805), .A2(n14806), .ZN(n14803) );
  OR2_X1 U14831 ( .A1(n14614), .A2(n14611), .ZN(n14806) );
  OR2_X1 U14832 ( .A1(n8127), .A2(n8017), .ZN(n14611) );
  OR3_X1 U14833 ( .A1(n8013), .A2(n8981), .A3(n8017), .ZN(n14614) );
  INV_X1 U14834 ( .A(n14613), .ZN(n14805) );
  OR2_X1 U14835 ( .A1(n14807), .A2(n14808), .ZN(n14613) );
  AND2_X1 U14836 ( .A1(b_1_), .A2(n14809), .ZN(n14808) );
  OR2_X1 U14837 ( .A1(n14810), .A2(n7598), .ZN(n14809) );
  AND2_X1 U14838 ( .A1(n7587), .A2(a_30_), .ZN(n7598) );
  AND2_X1 U14839 ( .A1(a_30_), .A2(n14718), .ZN(n14810) );
  AND2_X1 U14840 ( .A1(b_0_), .A2(n14811), .ZN(n14807) );
  OR2_X1 U14841 ( .A1(n14812), .A2(n7601), .ZN(n14811) );
  AND2_X1 U14842 ( .A1(n14813), .A2(a_31_), .ZN(n7601) );
  AND2_X1 U14843 ( .A1(a_31_), .A2(n8013), .ZN(n14812) );
  XOR2_X1 U14844 ( .A(n14814), .B(n14815), .Z(n14615) );
  OR2_X1 U14845 ( .A1(n14816), .A2(n14817), .ZN(n14814) );
  AND2_X1 U14846 ( .A1(n14818), .A2(n14819), .ZN(n14816) );
  OR2_X1 U14847 ( .A1(n14813), .A2(n14718), .ZN(n14818) );
  OR2_X1 U14848 ( .A1(n14622), .A2(n14619), .ZN(n14799) );
  XNOR2_X1 U14849 ( .A(n14820), .B(n14821), .ZN(n14619) );
  XOR2_X1 U14850 ( .A(n14822), .B(n14823), .Z(n14821) );
  OR2_X1 U14851 ( .A1(n8121), .A2(n8017), .ZN(n14622) );
  XNOR2_X1 U14852 ( .A(n14824), .B(n14825), .ZN(n14623) );
  XNOR2_X1 U14853 ( .A(n14826), .B(n14827), .ZN(n14824) );
  XNOR2_X1 U14854 ( .A(n14828), .B(n14829), .ZN(n14627) );
  XNOR2_X1 U14855 ( .A(n14830), .B(n14831), .ZN(n14828) );
  XNOR2_X1 U14856 ( .A(n14832), .B(n14833), .ZN(n14631) );
  XNOR2_X1 U14857 ( .A(n14834), .B(n14835), .ZN(n14832) );
  XNOR2_X1 U14858 ( .A(n14836), .B(n14837), .ZN(n14635) );
  XNOR2_X1 U14859 ( .A(n14838), .B(n14839), .ZN(n14836) );
  XNOR2_X1 U14860 ( .A(n14840), .B(n14841), .ZN(n14639) );
  XNOR2_X1 U14861 ( .A(n14842), .B(n14843), .ZN(n14840) );
  XNOR2_X1 U14862 ( .A(n14844), .B(n14845), .ZN(n14643) );
  XNOR2_X1 U14863 ( .A(n14846), .B(n14847), .ZN(n14844) );
  XNOR2_X1 U14864 ( .A(n14848), .B(n14849), .ZN(n14647) );
  XNOR2_X1 U14865 ( .A(n14850), .B(n14851), .ZN(n14848) );
  XNOR2_X1 U14866 ( .A(n14852), .B(n14853), .ZN(n14651) );
  XNOR2_X1 U14867 ( .A(n14854), .B(n14855), .ZN(n14852) );
  XNOR2_X1 U14868 ( .A(n14856), .B(n14857), .ZN(n14655) );
  XNOR2_X1 U14869 ( .A(n14858), .B(n14859), .ZN(n14856) );
  XNOR2_X1 U14870 ( .A(n14860), .B(n14861), .ZN(n14659) );
  XNOR2_X1 U14871 ( .A(n14862), .B(n14863), .ZN(n14860) );
  XNOR2_X1 U14872 ( .A(n14864), .B(n14865), .ZN(n14663) );
  XNOR2_X1 U14873 ( .A(n14866), .B(n14867), .ZN(n14864) );
  XNOR2_X1 U14874 ( .A(n14868), .B(n14869), .ZN(n14667) );
  XNOR2_X1 U14875 ( .A(n14870), .B(n14871), .ZN(n14868) );
  XNOR2_X1 U14876 ( .A(n14872), .B(n14873), .ZN(n14671) );
  XNOR2_X1 U14877 ( .A(n14874), .B(n14875), .ZN(n14872) );
  XNOR2_X1 U14878 ( .A(n14876), .B(n14877), .ZN(n14675) );
  XNOR2_X1 U14879 ( .A(n14878), .B(n14879), .ZN(n14876) );
  XNOR2_X1 U14880 ( .A(n14880), .B(n14881), .ZN(n14679) );
  XNOR2_X1 U14881 ( .A(n14882), .B(n14883), .ZN(n14880) );
  XNOR2_X1 U14882 ( .A(n14884), .B(n14885), .ZN(n14683) );
  XNOR2_X1 U14883 ( .A(n14886), .B(n14887), .ZN(n14884) );
  XNOR2_X1 U14884 ( .A(n14888), .B(n14889), .ZN(n14687) );
  XNOR2_X1 U14885 ( .A(n14890), .B(n14891), .ZN(n14888) );
  XNOR2_X1 U14886 ( .A(n14892), .B(n14893), .ZN(n14691) );
  XNOR2_X1 U14887 ( .A(n14894), .B(n14895), .ZN(n14892) );
  XNOR2_X1 U14888 ( .A(n14896), .B(n14897), .ZN(n14695) );
  XNOR2_X1 U14889 ( .A(n14898), .B(n14899), .ZN(n14896) );
  XOR2_X1 U14890 ( .A(n14900), .B(n14901), .Z(n8576) );
  XOR2_X1 U14891 ( .A(n14902), .B(n14903), .Z(n14901) );
  XOR2_X1 U14892 ( .A(n14904), .B(n14905), .Z(n8511) );
  XOR2_X1 U14893 ( .A(n14906), .B(n14907), .Z(n14905) );
  XOR2_X1 U14894 ( .A(n14908), .B(n14909), .Z(n8457) );
  XOR2_X1 U14895 ( .A(n14910), .B(n14911), .Z(n14909) );
  XOR2_X1 U14896 ( .A(n14912), .B(n14913), .Z(n8412) );
  XOR2_X1 U14897 ( .A(n14914), .B(n14915), .Z(n14913) );
  XOR2_X1 U14898 ( .A(n14916), .B(n14917), .Z(n8366) );
  XOR2_X1 U14899 ( .A(n14918), .B(n14919), .Z(n14917) );
  OR2_X1 U14900 ( .A1(n8016), .A2(n8017), .ZN(n8018) );
  INV_X1 U14901 ( .A(b_2_), .ZN(n8017) );
  XOR2_X1 U14902 ( .A(n14920), .B(n14921), .Z(n8337) );
  XOR2_X1 U14903 ( .A(n14922), .B(n14923), .Z(n14921) );
  XOR2_X1 U14904 ( .A(n14711), .B(n14924), .Z(n8304) );
  XOR2_X1 U14905 ( .A(n14712), .B(n14714), .Z(n14924) );
  OR2_X1 U14906 ( .A1(n8021), .A2(n14718), .ZN(n14714) );
  OR2_X1 U14907 ( .A1(n14925), .A2(n14926), .ZN(n14712) );
  AND2_X1 U14908 ( .A1(n14920), .A2(n14922), .ZN(n14926) );
  AND2_X1 U14909 ( .A1(n14927), .A2(n14923), .ZN(n14925) );
  OR2_X1 U14910 ( .A1(n8025), .A2(n14718), .ZN(n14923) );
  OR2_X1 U14911 ( .A1(n14922), .A2(n14920), .ZN(n14927) );
  OR2_X1 U14912 ( .A1(n8013), .A2(n8021), .ZN(n14920) );
  OR2_X1 U14913 ( .A1(n14928), .A2(n14929), .ZN(n14922) );
  AND2_X1 U14914 ( .A1(n14916), .A2(n14918), .ZN(n14929) );
  AND2_X1 U14915 ( .A1(n14930), .A2(n14919), .ZN(n14928) );
  OR2_X1 U14916 ( .A1(n8030), .A2(n14718), .ZN(n14919) );
  OR2_X1 U14917 ( .A1(n14918), .A2(n14916), .ZN(n14930) );
  OR2_X1 U14918 ( .A1(n8013), .A2(n8025), .ZN(n14916) );
  OR2_X1 U14919 ( .A1(n14931), .A2(n14932), .ZN(n14918) );
  AND2_X1 U14920 ( .A1(n14912), .A2(n14914), .ZN(n14932) );
  AND2_X1 U14921 ( .A1(n14933), .A2(n14915), .ZN(n14931) );
  OR2_X1 U14922 ( .A1(n8034), .A2(n14718), .ZN(n14915) );
  OR2_X1 U14923 ( .A1(n14914), .A2(n14912), .ZN(n14933) );
  OR2_X1 U14924 ( .A1(n8013), .A2(n8030), .ZN(n14912) );
  OR2_X1 U14925 ( .A1(n14934), .A2(n14935), .ZN(n14914) );
  AND2_X1 U14926 ( .A1(n14908), .A2(n14910), .ZN(n14935) );
  AND2_X1 U14927 ( .A1(n14936), .A2(n14911), .ZN(n14934) );
  OR2_X1 U14928 ( .A1(n8039), .A2(n14718), .ZN(n14911) );
  OR2_X1 U14929 ( .A1(n14910), .A2(n14908), .ZN(n14936) );
  OR2_X1 U14930 ( .A1(n8013), .A2(n8034), .ZN(n14908) );
  OR2_X1 U14931 ( .A1(n14937), .A2(n14938), .ZN(n14910) );
  AND2_X1 U14932 ( .A1(n14904), .A2(n14906), .ZN(n14938) );
  AND2_X1 U14933 ( .A1(n14939), .A2(n14907), .ZN(n14937) );
  OR2_X1 U14934 ( .A1(n8043), .A2(n14718), .ZN(n14907) );
  OR2_X1 U14935 ( .A1(n14906), .A2(n14904), .ZN(n14939) );
  OR2_X1 U14936 ( .A1(n8013), .A2(n8039), .ZN(n14904) );
  OR2_X1 U14937 ( .A1(n14940), .A2(n14941), .ZN(n14906) );
  AND2_X1 U14938 ( .A1(n14900), .A2(n14902), .ZN(n14941) );
  AND2_X1 U14939 ( .A1(n14942), .A2(n14903), .ZN(n14940) );
  OR2_X1 U14940 ( .A1(n8048), .A2(n14718), .ZN(n14903) );
  OR2_X1 U14941 ( .A1(n14902), .A2(n14900), .ZN(n14942) );
  OR2_X1 U14942 ( .A1(n8013), .A2(n8043), .ZN(n14900) );
  OR2_X1 U14943 ( .A1(n14943), .A2(n14944), .ZN(n14902) );
  AND2_X1 U14944 ( .A1(n14897), .A2(n14899), .ZN(n14944) );
  AND2_X1 U14945 ( .A1(n14945), .A2(n14898), .ZN(n14943) );
  OR2_X1 U14946 ( .A1(n8052), .A2(n14718), .ZN(n14898) );
  OR2_X1 U14947 ( .A1(n14899), .A2(n14897), .ZN(n14945) );
  OR2_X1 U14948 ( .A1(n8013), .A2(n8048), .ZN(n14897) );
  OR2_X1 U14949 ( .A1(n14946), .A2(n14947), .ZN(n14899) );
  AND2_X1 U14950 ( .A1(n14893), .A2(n14895), .ZN(n14947) );
  AND2_X1 U14951 ( .A1(n14948), .A2(n14894), .ZN(n14946) );
  OR2_X1 U14952 ( .A1(n8057), .A2(n14718), .ZN(n14894) );
  OR2_X1 U14953 ( .A1(n14895), .A2(n14893), .ZN(n14948) );
  OR2_X1 U14954 ( .A1(n8013), .A2(n8052), .ZN(n14893) );
  OR2_X1 U14955 ( .A1(n14949), .A2(n14950), .ZN(n14895) );
  AND2_X1 U14956 ( .A1(n14889), .A2(n14891), .ZN(n14950) );
  AND2_X1 U14957 ( .A1(n14951), .A2(n14890), .ZN(n14949) );
  OR2_X1 U14958 ( .A1(n8061), .A2(n14718), .ZN(n14890) );
  OR2_X1 U14959 ( .A1(n14891), .A2(n14889), .ZN(n14951) );
  OR2_X1 U14960 ( .A1(n8013), .A2(n8057), .ZN(n14889) );
  OR2_X1 U14961 ( .A1(n14952), .A2(n14953), .ZN(n14891) );
  AND2_X1 U14962 ( .A1(n14885), .A2(n14887), .ZN(n14953) );
  AND2_X1 U14963 ( .A1(n14954), .A2(n14886), .ZN(n14952) );
  OR2_X1 U14964 ( .A1(n8066), .A2(n14718), .ZN(n14886) );
  OR2_X1 U14965 ( .A1(n14887), .A2(n14885), .ZN(n14954) );
  OR2_X1 U14966 ( .A1(n8013), .A2(n8061), .ZN(n14885) );
  OR2_X1 U14967 ( .A1(n14955), .A2(n14956), .ZN(n14887) );
  AND2_X1 U14968 ( .A1(n14881), .A2(n14883), .ZN(n14956) );
  AND2_X1 U14969 ( .A1(n14957), .A2(n14882), .ZN(n14955) );
  OR2_X1 U14970 ( .A1(n8070), .A2(n14718), .ZN(n14882) );
  OR2_X1 U14971 ( .A1(n14883), .A2(n14881), .ZN(n14957) );
  OR2_X1 U14972 ( .A1(n8013), .A2(n8066), .ZN(n14881) );
  OR2_X1 U14973 ( .A1(n14958), .A2(n14959), .ZN(n14883) );
  AND2_X1 U14974 ( .A1(n14877), .A2(n14879), .ZN(n14959) );
  AND2_X1 U14975 ( .A1(n14960), .A2(n14878), .ZN(n14958) );
  OR2_X1 U14976 ( .A1(n8075), .A2(n14718), .ZN(n14878) );
  OR2_X1 U14977 ( .A1(n14879), .A2(n14877), .ZN(n14960) );
  OR2_X1 U14978 ( .A1(n8013), .A2(n8070), .ZN(n14877) );
  OR2_X1 U14979 ( .A1(n14961), .A2(n14962), .ZN(n14879) );
  AND2_X1 U14980 ( .A1(n14873), .A2(n14875), .ZN(n14962) );
  AND2_X1 U14981 ( .A1(n14963), .A2(n14874), .ZN(n14961) );
  OR2_X1 U14982 ( .A1(n8079), .A2(n14718), .ZN(n14874) );
  OR2_X1 U14983 ( .A1(n14875), .A2(n14873), .ZN(n14963) );
  OR2_X1 U14984 ( .A1(n8013), .A2(n8075), .ZN(n14873) );
  OR2_X1 U14985 ( .A1(n14964), .A2(n14965), .ZN(n14875) );
  AND2_X1 U14986 ( .A1(n14869), .A2(n14871), .ZN(n14965) );
  AND2_X1 U14987 ( .A1(n14966), .A2(n14870), .ZN(n14964) );
  OR2_X1 U14988 ( .A1(n8084), .A2(n14718), .ZN(n14870) );
  OR2_X1 U14989 ( .A1(n14871), .A2(n14869), .ZN(n14966) );
  OR2_X1 U14990 ( .A1(n8013), .A2(n8079), .ZN(n14869) );
  OR2_X1 U14991 ( .A1(n14967), .A2(n14968), .ZN(n14871) );
  AND2_X1 U14992 ( .A1(n14865), .A2(n14867), .ZN(n14968) );
  AND2_X1 U14993 ( .A1(n14969), .A2(n14866), .ZN(n14967) );
  OR2_X1 U14994 ( .A1(n8088), .A2(n14718), .ZN(n14866) );
  OR2_X1 U14995 ( .A1(n14867), .A2(n14865), .ZN(n14969) );
  OR2_X1 U14996 ( .A1(n8013), .A2(n8084), .ZN(n14865) );
  OR2_X1 U14997 ( .A1(n14970), .A2(n14971), .ZN(n14867) );
  AND2_X1 U14998 ( .A1(n14861), .A2(n14863), .ZN(n14971) );
  AND2_X1 U14999 ( .A1(n14972), .A2(n14862), .ZN(n14970) );
  OR2_X1 U15000 ( .A1(n8093), .A2(n14718), .ZN(n14862) );
  OR2_X1 U15001 ( .A1(n14863), .A2(n14861), .ZN(n14972) );
  OR2_X1 U15002 ( .A1(n8013), .A2(n8088), .ZN(n14861) );
  OR2_X1 U15003 ( .A1(n14973), .A2(n14974), .ZN(n14863) );
  AND2_X1 U15004 ( .A1(n14857), .A2(n14859), .ZN(n14974) );
  AND2_X1 U15005 ( .A1(n14975), .A2(n14858), .ZN(n14973) );
  OR2_X1 U15006 ( .A1(n8097), .A2(n14718), .ZN(n14858) );
  OR2_X1 U15007 ( .A1(n14859), .A2(n14857), .ZN(n14975) );
  OR2_X1 U15008 ( .A1(n8013), .A2(n8093), .ZN(n14857) );
  OR2_X1 U15009 ( .A1(n14976), .A2(n14977), .ZN(n14859) );
  AND2_X1 U15010 ( .A1(n14853), .A2(n14855), .ZN(n14977) );
  AND2_X1 U15011 ( .A1(n14978), .A2(n14854), .ZN(n14976) );
  OR2_X1 U15012 ( .A1(n8102), .A2(n14718), .ZN(n14854) );
  OR2_X1 U15013 ( .A1(n14855), .A2(n14853), .ZN(n14978) );
  OR2_X1 U15014 ( .A1(n8013), .A2(n8097), .ZN(n14853) );
  OR2_X1 U15015 ( .A1(n14979), .A2(n14980), .ZN(n14855) );
  AND2_X1 U15016 ( .A1(n14849), .A2(n14851), .ZN(n14980) );
  AND2_X1 U15017 ( .A1(n14981), .A2(n14850), .ZN(n14979) );
  OR2_X1 U15018 ( .A1(n8106), .A2(n14718), .ZN(n14850) );
  OR2_X1 U15019 ( .A1(n14851), .A2(n14849), .ZN(n14981) );
  OR2_X1 U15020 ( .A1(n8013), .A2(n8102), .ZN(n14849) );
  OR2_X1 U15021 ( .A1(n14982), .A2(n14983), .ZN(n14851) );
  AND2_X1 U15022 ( .A1(n14845), .A2(n14847), .ZN(n14983) );
  AND2_X1 U15023 ( .A1(n14984), .A2(n14846), .ZN(n14982) );
  OR2_X1 U15024 ( .A1(n8109), .A2(n14718), .ZN(n14846) );
  OR2_X1 U15025 ( .A1(n14847), .A2(n14845), .ZN(n14984) );
  OR2_X1 U15026 ( .A1(n8013), .A2(n8106), .ZN(n14845) );
  OR2_X1 U15027 ( .A1(n14985), .A2(n14986), .ZN(n14847) );
  AND2_X1 U15028 ( .A1(n14841), .A2(n14843), .ZN(n14986) );
  AND2_X1 U15029 ( .A1(n14987), .A2(n14842), .ZN(n14985) );
  OR2_X1 U15030 ( .A1(n8112), .A2(n14718), .ZN(n14842) );
  OR2_X1 U15031 ( .A1(n14843), .A2(n14841), .ZN(n14987) );
  OR2_X1 U15032 ( .A1(n8013), .A2(n8109), .ZN(n14841) );
  OR2_X1 U15033 ( .A1(n14988), .A2(n14989), .ZN(n14843) );
  AND2_X1 U15034 ( .A1(n14837), .A2(n14839), .ZN(n14989) );
  AND2_X1 U15035 ( .A1(n14990), .A2(n14838), .ZN(n14988) );
  OR2_X1 U15036 ( .A1(n8115), .A2(n14718), .ZN(n14838) );
  OR2_X1 U15037 ( .A1(n14839), .A2(n14837), .ZN(n14990) );
  OR2_X1 U15038 ( .A1(n8013), .A2(n8112), .ZN(n14837) );
  OR2_X1 U15039 ( .A1(n14991), .A2(n14992), .ZN(n14839) );
  AND2_X1 U15040 ( .A1(n14833), .A2(n14835), .ZN(n14992) );
  AND2_X1 U15041 ( .A1(n14993), .A2(n14834), .ZN(n14991) );
  OR2_X1 U15042 ( .A1(n8118), .A2(n14718), .ZN(n14834) );
  OR2_X1 U15043 ( .A1(n14835), .A2(n14833), .ZN(n14993) );
  OR2_X1 U15044 ( .A1(n8013), .A2(n8115), .ZN(n14833) );
  OR2_X1 U15045 ( .A1(n14994), .A2(n14995), .ZN(n14835) );
  AND2_X1 U15046 ( .A1(n14829), .A2(n14831), .ZN(n14995) );
  AND2_X1 U15047 ( .A1(n14996), .A2(n14830), .ZN(n14994) );
  OR2_X1 U15048 ( .A1(n8121), .A2(n14718), .ZN(n14830) );
  OR2_X1 U15049 ( .A1(n14831), .A2(n14829), .ZN(n14996) );
  OR2_X1 U15050 ( .A1(n8013), .A2(n8118), .ZN(n14829) );
  OR2_X1 U15051 ( .A1(n14997), .A2(n14998), .ZN(n14831) );
  AND2_X1 U15052 ( .A1(n14825), .A2(n14827), .ZN(n14998) );
  AND2_X1 U15053 ( .A1(n14999), .A2(n14826), .ZN(n14997) );
  OR2_X1 U15054 ( .A1(n8124), .A2(n14718), .ZN(n14826) );
  OR2_X1 U15055 ( .A1(n14827), .A2(n14825), .ZN(n14999) );
  OR2_X1 U15056 ( .A1(n8013), .A2(n8121), .ZN(n14825) );
  OR2_X1 U15057 ( .A1(n15000), .A2(n15001), .ZN(n14827) );
  AND2_X1 U15058 ( .A1(n14820), .A2(n14823), .ZN(n15001) );
  AND2_X1 U15059 ( .A1(n15002), .A2(n15003), .ZN(n15000) );
  OR2_X1 U15060 ( .A1(n14823), .A2(n14820), .ZN(n15003) );
  OR2_X1 U15061 ( .A1(n8013), .A2(n8124), .ZN(n14820) );
  OR2_X1 U15062 ( .A1(n8127), .A2(n14718), .ZN(n14823) );
  INV_X1 U15063 ( .A(b_0_), .ZN(n14718) );
  INV_X1 U15064 ( .A(n14822), .ZN(n15002) );
  OR2_X1 U15065 ( .A1(n14817), .A2(n14815), .ZN(n14822) );
  AND3_X1 U15066 ( .A1(b_1_), .A2(n8130), .A3(b_0_), .ZN(n14815) );
  INV_X1 U15067 ( .A(n8981), .ZN(n8130) );
  AND3_X1 U15068 ( .A1(a_30_), .A2(b_0_), .A3(n15004), .ZN(n14817) );
  INV_X1 U15069 ( .A(n14819), .ZN(n15004) );
  OR2_X1 U15070 ( .A1(n8013), .A2(n8127), .ZN(n14819) );
  OR2_X1 U15071 ( .A1(n8013), .A2(n8016), .ZN(n14711) );
  OR2_X1 U15072 ( .A1(n15005), .A2(n8008), .ZN(n7584) );
  AND2_X1 U15073 ( .A1(n8297), .A2(b_0_), .ZN(n8008) );
  AND3_X1 U15074 ( .A1(n7999), .A2(n15006), .A3(n15007), .ZN(n15005) );
  OR2_X1 U15075 ( .A1(b_0_), .A2(n8297), .ZN(n15007) );
  INV_X1 U15076 ( .A(a_0_), .ZN(n8297) );
  OR3_X1 U15077 ( .A1(n15008), .A2(n15009), .A3(n15010), .ZN(n15006) );
  AND2_X1 U15078 ( .A1(b_2_), .A2(n8016), .ZN(n15010) );
  AND3_X1 U15079 ( .A1(n15011), .A2(n7975), .A3(n15012), .ZN(n15009) );
  OR2_X1 U15080 ( .A1(b_2_), .A2(n8016), .ZN(n15012) );
  INV_X1 U15081 ( .A(a_2_), .ZN(n8016) );
  OR2_X1 U15082 ( .A1(b_3_), .A2(n8021), .ZN(n7975) );
  INV_X1 U15083 ( .A(a_3_), .ZN(n8021) );
  OR3_X1 U15084 ( .A1(n15013), .A2(n15014), .A3(n15015), .ZN(n15011) );
  AND3_X1 U15085 ( .A1(n15016), .A2(n7951), .A3(n15017), .ZN(n15015) );
  OR2_X1 U15086 ( .A1(b_4_), .A2(n8025), .ZN(n15017) );
  OR2_X1 U15087 ( .A1(b_5_), .A2(n8030), .ZN(n7951) );
  INV_X1 U15088 ( .A(a_5_), .ZN(n8030) );
  OR3_X1 U15089 ( .A1(n15018), .A2(n15019), .A3(n15020), .ZN(n15016) );
  AND2_X1 U15090 ( .A1(b_6_), .A2(n8034), .ZN(n15020) );
  AND3_X1 U15091 ( .A1(n15021), .A2(n7927), .A3(n15022), .ZN(n15019) );
  OR2_X1 U15092 ( .A1(b_6_), .A2(n8034), .ZN(n15022) );
  INV_X1 U15093 ( .A(a_6_), .ZN(n8034) );
  OR2_X1 U15094 ( .A1(b_7_), .A2(n8039), .ZN(n7927) );
  INV_X1 U15095 ( .A(a_7_), .ZN(n8039) );
  OR3_X1 U15096 ( .A1(n15023), .A2(n15024), .A3(n15025), .ZN(n15021) );
  AND3_X1 U15097 ( .A1(n15026), .A2(n7893), .A3(n15027), .ZN(n15025) );
  OR2_X1 U15098 ( .A1(b_8_), .A2(n8043), .ZN(n15027) );
  OR2_X1 U15099 ( .A1(b_9_), .A2(n8048), .ZN(n7893) );
  INV_X1 U15100 ( .A(a_9_), .ZN(n8048) );
  OR3_X1 U15101 ( .A1(n15028), .A2(n15029), .A3(n15030), .ZN(n15026) );
  AND2_X1 U15102 ( .A1(b_10_), .A2(n8052), .ZN(n15030) );
  INV_X1 U15103 ( .A(n7892), .ZN(n15029) );
  OR2_X1 U15104 ( .A1(a_9_), .A2(n8049), .ZN(n7892) );
  AND3_X1 U15105 ( .A1(n15031), .A2(n7869), .A3(n15032), .ZN(n15028) );
  OR2_X1 U15106 ( .A1(b_10_), .A2(n8052), .ZN(n15032) );
  INV_X1 U15107 ( .A(a_10_), .ZN(n8052) );
  OR2_X1 U15108 ( .A1(b_11_), .A2(n8057), .ZN(n7869) );
  INV_X1 U15109 ( .A(a_11_), .ZN(n8057) );
  OR3_X1 U15110 ( .A1(n15033), .A2(n15034), .A3(n15035), .ZN(n15031) );
  AND3_X1 U15111 ( .A1(n15036), .A2(n7845), .A3(n15037), .ZN(n15035) );
  OR2_X1 U15112 ( .A1(b_12_), .A2(n8061), .ZN(n15037) );
  OR2_X1 U15113 ( .A1(b_13_), .A2(n8066), .ZN(n7845) );
  INV_X1 U15114 ( .A(a_13_), .ZN(n8066) );
  OR3_X1 U15115 ( .A1(n15038), .A2(n15039), .A3(n15040), .ZN(n15036) );
  AND2_X1 U15116 ( .A1(b_14_), .A2(n8070), .ZN(n15040) );
  AND3_X1 U15117 ( .A1(n15041), .A2(n7821), .A3(n15042), .ZN(n15039) );
  OR2_X1 U15118 ( .A1(b_14_), .A2(n8070), .ZN(n15042) );
  INV_X1 U15119 ( .A(a_14_), .ZN(n8070) );
  OR2_X1 U15120 ( .A1(b_15_), .A2(n8075), .ZN(n7821) );
  INV_X1 U15121 ( .A(a_15_), .ZN(n8075) );
  OR3_X1 U15122 ( .A1(n15043), .A2(n15044), .A3(n15045), .ZN(n15041) );
  AND3_X1 U15123 ( .A1(n15046), .A2(n7797), .A3(n15047), .ZN(n15045) );
  OR2_X1 U15124 ( .A1(b_16_), .A2(n8079), .ZN(n15047) );
  OR2_X1 U15125 ( .A1(b_17_), .A2(n8084), .ZN(n7797) );
  INV_X1 U15126 ( .A(a_17_), .ZN(n8084) );
  OR3_X1 U15127 ( .A1(n15048), .A2(n15049), .A3(n15050), .ZN(n15046) );
  AND2_X1 U15128 ( .A1(b_18_), .A2(n8088), .ZN(n15050) );
  AND3_X1 U15129 ( .A1(n15051), .A2(n7770), .A3(n15052), .ZN(n15049) );
  OR2_X1 U15130 ( .A1(b_18_), .A2(n8088), .ZN(n15052) );
  INV_X1 U15131 ( .A(a_18_), .ZN(n8088) );
  OR2_X1 U15132 ( .A1(b_19_), .A2(n8093), .ZN(n7770) );
  INV_X1 U15133 ( .A(a_19_), .ZN(n8093) );
  OR3_X1 U15134 ( .A1(n15053), .A2(n15054), .A3(n15055), .ZN(n15051) );
  AND3_X1 U15135 ( .A1(n15056), .A2(n7746), .A3(n15057), .ZN(n15055) );
  OR2_X1 U15136 ( .A1(b_20_), .A2(n8097), .ZN(n15057) );
  OR2_X1 U15137 ( .A1(b_21_), .A2(n8102), .ZN(n7746) );
  INV_X1 U15138 ( .A(a_21_), .ZN(n8102) );
  OR3_X1 U15139 ( .A1(n15058), .A2(n15059), .A3(n15060), .ZN(n15056) );
  AND2_X1 U15140 ( .A1(b_22_), .A2(n8106), .ZN(n15060) );
  AND3_X1 U15141 ( .A1(n15061), .A2(n15062), .A3(n15063), .ZN(n15059) );
  OR2_X1 U15142 ( .A1(b_22_), .A2(n8106), .ZN(n15063) );
  INV_X1 U15143 ( .A(a_22_), .ZN(n8106) );
  OR2_X1 U15144 ( .A1(b_23_), .A2(n15064), .ZN(n15062) );
  AND2_X1 U15145 ( .A1(n8109), .A2(n15065), .ZN(n15064) );
  OR2_X1 U15146 ( .A1(n15065), .A2(n8109), .ZN(n15061) );
  INV_X1 U15147 ( .A(a_23_), .ZN(n8109) );
  OR2_X1 U15148 ( .A1(n15066), .A2(n15067), .ZN(n15065) );
  AND2_X1 U15149 ( .A1(b_24_), .A2(n8112), .ZN(n15067) );
  AND3_X1 U15150 ( .A1(n15068), .A2(n15069), .A3(n15070), .ZN(n15066) );
  OR2_X1 U15151 ( .A1(b_24_), .A2(n8112), .ZN(n15070) );
  INV_X1 U15152 ( .A(a_24_), .ZN(n8112) );
  OR2_X1 U15153 ( .A1(b_25_), .A2(n15071), .ZN(n15069) );
  AND2_X1 U15154 ( .A1(n8115), .A2(n15072), .ZN(n15071) );
  OR2_X1 U15155 ( .A1(n15072), .A2(n8115), .ZN(n15068) );
  INV_X1 U15156 ( .A(a_25_), .ZN(n8115) );
  OR2_X1 U15157 ( .A1(n15073), .A2(n15074), .ZN(n15072) );
  AND2_X1 U15158 ( .A1(b_26_), .A2(n8118), .ZN(n15074) );
  AND3_X1 U15159 ( .A1(n15075), .A2(n15076), .A3(n15077), .ZN(n15073) );
  OR2_X1 U15160 ( .A1(b_26_), .A2(n8118), .ZN(n15077) );
  INV_X1 U15161 ( .A(a_26_), .ZN(n8118) );
  OR2_X1 U15162 ( .A1(b_27_), .A2(n15078), .ZN(n15076) );
  AND2_X1 U15163 ( .A1(n8121), .A2(n15079), .ZN(n15078) );
  OR2_X1 U15164 ( .A1(n15079), .A2(n8121), .ZN(n15075) );
  INV_X1 U15165 ( .A(a_27_), .ZN(n8121) );
  OR2_X1 U15166 ( .A1(n15080), .A2(n15081), .ZN(n15079) );
  AND2_X1 U15167 ( .A1(b_28_), .A2(n8124), .ZN(n15081) );
  AND3_X1 U15168 ( .A1(n15082), .A2(n15083), .A3(n15084), .ZN(n15080) );
  OR2_X1 U15169 ( .A1(b_29_), .A2(n8127), .ZN(n15084) );
  OR3_X1 U15170 ( .A1(n15085), .A2(n7610), .A3(n15086), .ZN(n15083) );
  INV_X1 U15171 ( .A(n15087), .ZN(n15086) );
  OR2_X1 U15172 ( .A1(a_30_), .A2(n7586), .ZN(n15087) );
  AND2_X1 U15173 ( .A1(n8980), .A2(a_31_), .ZN(n7586) );
  INV_X1 U15174 ( .A(b_31_), .ZN(n8980) );
  AND2_X1 U15175 ( .A1(n8127), .A2(b_29_), .ZN(n7610) );
  INV_X1 U15176 ( .A(a_29_), .ZN(n8127) );
  AND2_X1 U15177 ( .A1(b_30_), .A2(n15088), .ZN(n15085) );
  OR2_X1 U15178 ( .A1(b_31_), .A2(n8981), .ZN(n15088) );
  OR2_X1 U15179 ( .A1(n14813), .A2(n7587), .ZN(n8981) );
  INV_X1 U15180 ( .A(a_31_), .ZN(n7587) );
  INV_X1 U15181 ( .A(a_30_), .ZN(n14813) );
  OR2_X1 U15182 ( .A1(b_28_), .A2(n8124), .ZN(n15082) );
  INV_X1 U15183 ( .A(a_28_), .ZN(n8124) );
  INV_X1 U15184 ( .A(n7745), .ZN(n15058) );
  OR2_X1 U15185 ( .A1(a_21_), .A2(n8103), .ZN(n7745) );
  AND2_X1 U15186 ( .A1(b_20_), .A2(n8097), .ZN(n15054) );
  INV_X1 U15187 ( .A(a_20_), .ZN(n8097) );
  INV_X1 U15188 ( .A(n7769), .ZN(n15053) );
  OR2_X1 U15189 ( .A1(a_19_), .A2(n8094), .ZN(n7769) );
  INV_X1 U15190 ( .A(n7796), .ZN(n15048) );
  OR2_X1 U15191 ( .A1(a_17_), .A2(n8085), .ZN(n7796) );
  AND2_X1 U15192 ( .A1(b_16_), .A2(n8079), .ZN(n15044) );
  INV_X1 U15193 ( .A(a_16_), .ZN(n8079) );
  INV_X1 U15194 ( .A(n7820), .ZN(n15043) );
  OR2_X1 U15195 ( .A1(a_15_), .A2(n8076), .ZN(n7820) );
  INV_X1 U15196 ( .A(n7844), .ZN(n15038) );
  OR2_X1 U15197 ( .A1(a_13_), .A2(n8067), .ZN(n7844) );
  AND2_X1 U15198 ( .A1(b_12_), .A2(n8061), .ZN(n15034) );
  INV_X1 U15199 ( .A(a_12_), .ZN(n8061) );
  INV_X1 U15200 ( .A(n7868), .ZN(n15033) );
  OR2_X1 U15201 ( .A1(a_11_), .A2(n8058), .ZN(n7868) );
  AND2_X1 U15202 ( .A1(b_8_), .A2(n8043), .ZN(n15024) );
  INV_X1 U15203 ( .A(a_8_), .ZN(n8043) );
  INV_X1 U15204 ( .A(n7926), .ZN(n15023) );
  OR2_X1 U15205 ( .A1(a_7_), .A2(n8040), .ZN(n7926) );
  INV_X1 U15206 ( .A(n7950), .ZN(n15018) );
  OR2_X1 U15207 ( .A1(a_5_), .A2(n8031), .ZN(n7950) );
  AND2_X1 U15208 ( .A1(b_4_), .A2(n8025), .ZN(n15014) );
  INV_X1 U15209 ( .A(a_4_), .ZN(n8025) );
  INV_X1 U15210 ( .A(n7974), .ZN(n15013) );
  OR2_X1 U15211 ( .A1(a_3_), .A2(n8022), .ZN(n7974) );
  INV_X1 U15212 ( .A(n7998), .ZN(n15008) );
  OR2_X1 U15213 ( .A1(a_1_), .A2(n8013), .ZN(n7998) );
  INV_X1 U15214 ( .A(b_1_), .ZN(n8013) );
  OR2_X1 U15215 ( .A1(b_1_), .A2(n8012), .ZN(n7999) );
  INV_X1 U15216 ( .A(a_1_), .ZN(n8012) );
endmodule

