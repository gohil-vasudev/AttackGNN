module add_mul_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, operation_0_, operation_1_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, Result_17_, 
        Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, Result_23_, 
        Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, Result_29_, 
        Result_30_, Result_31_, Result_32_, Result_33_, Result_34_, Result_35_, 
        Result_36_, Result_37_, Result_38_, Result_39_, Result_40_, Result_41_, 
        Result_42_, Result_43_, Result_44_, Result_45_, Result_46_, Result_47_, 
        Result_48_, Result_49_, Result_50_, Result_51_, Result_52_, Result_53_, 
        Result_54_, Result_55_, Result_56_, Result_57_, Result_58_, Result_59_, 
        Result_60_, Result_61_, Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
         n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
         n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
         n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
         n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
         n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403,
         n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
         n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
         n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
         n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
         n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
         n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
         n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
         n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
         n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
         n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
         n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
         n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
         n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571,
         n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
         n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595,
         n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
         n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
         n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619,
         n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
         n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
         n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643,
         n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
         n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
         n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
         n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
         n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
         n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691,
         n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699,
         n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
         n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715,
         n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723,
         n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
         n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739,
         n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
         n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
         n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763,
         n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771,
         n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
         n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787,
         n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795,
         n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
         n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811,
         n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
         n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
         n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835,
         n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843,
         n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
         n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859,
         n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867,
         n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
         n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
         n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
         n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899,
         n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907,
         n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
         n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
         n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931,
         n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939,
         n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
         n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955,
         n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
         n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971,
         n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979,
         n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
         n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
         n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003,
         n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011,
         n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
         n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027,
         n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
         n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043,
         n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
         n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
         n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
         n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075,
         n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083,
         n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
         n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
         n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
         n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
         n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147,
         n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
         n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
         n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171,
         n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
         n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
         n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195,
         n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
         n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211,
         n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219,
         n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227,
         n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
         n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
         n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
         n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259,
         n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
         n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
         n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283,
         n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
         n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299,
         n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
         n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315,
         n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
         n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
         n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
         n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
         n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
         n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
         n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
         n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
         n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
         n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
         n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
         n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427,
         n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435,
         n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443,
         n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
         n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459,
         n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
         n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475,
         n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483,
         n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
         n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499,
         n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507,
         n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
         n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
         n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
         n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
         n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
         n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
         n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
         n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
         n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
         n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
         n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627,
         n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
         n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
         n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651,
         n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659,
         n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
         n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675,
         n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
         n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
         n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699,
         n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
         n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723,
         n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731,
         n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
         n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747,
         n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
         n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
         n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771,
         n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779,
         n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
         n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795,
         n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803,
         n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
         n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
         n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
         n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
         n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843,
         n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
         n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
         n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867,
         n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875,
         n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
         n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891,
         n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
         n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
         n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
         n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
         n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
         n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
         n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947,
         n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
         n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
         n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
         n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
         n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987,
         n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011,
         n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
         n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
         n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
         n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
         n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
         n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
         n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
         n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163,
         n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
         n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227,
         n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
         n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
         n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
         n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371,
         n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
         n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
         n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
         n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491,
         n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
         n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
         n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
         n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
         n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659,
         n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
         n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
         n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
         n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
         n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
         n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707,
         n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
         n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
         n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
         n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739,
         n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
         n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
         n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
         n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
         n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883,
         n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
         n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
         n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
         n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
         n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923,
         n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931,
         n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
         n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947,
         n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955,
         n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
         n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
         n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
         n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987,
         n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995,
         n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003,
         n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
         n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019,
         n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027,
         n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
         n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
         n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
         n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059,
         n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067,
         n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
         n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
         n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
         n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131,
         n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139,
         n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
         n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
         n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163,
         n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171,
         n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
         n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
         n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
         n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
         n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
         n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
         n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
         n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235,
         n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243,
         n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
         n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
         n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
         n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
         n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283,
         n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
         n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299,
         n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307,
         n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315,
         n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
         n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331,
         n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
         n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347,
         n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355,
         n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
         n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419,
         n29420, n29421, n29422, n29423, n29424;

  AND2_X2 U14804 ( .A1(n15862), .A2(n15863), .ZN(n14793) );
  AND2_X2 U14805 ( .A1(n15862), .A2(operation_0_), .ZN(n14792) );
  AND2_X2 U14806 ( .A1(n15863), .A2(operation_1_), .ZN(n14791) );
  AND2_X2 U14807 ( .A1(operation_0_), .A2(operation_1_), .ZN(n14744) );
  INV_X2 U14808 ( .A(a_28_), .ZN(n14891) );
  INV_X2 U14809 ( .A(a_2_), .ZN(n15808) );
  OR2_X1 U14810 ( .A1(n14740), .A2(n14741), .ZN(Result_9_) );
  AND3_X1 U14811 ( .A1(n14742), .A2(n14743), .A3(n14744), .ZN(n14740) );
  OR3_X1 U14812 ( .A1(n14745), .A2(n14746), .A3(n14747), .ZN(n14743) );
  INV_X1 U14813 ( .A(n14748), .ZN(n14747) );
  AND2_X1 U14814 ( .A1(n14749), .A2(n14750), .ZN(n14746) );
  AND2_X1 U14815 ( .A1(n14751), .A2(n14752), .ZN(n14745) );
  INV_X1 U14816 ( .A(n14750), .ZN(n14751) );
  OR2_X1 U14817 ( .A1(n14750), .A2(n14748), .ZN(n14742) );
  OR2_X1 U14818 ( .A1(n14753), .A2(n14741), .ZN(Result_8_) );
  AND3_X1 U14819 ( .A1(n14754), .A2(n14755), .A3(n14744), .ZN(n14753) );
  OR3_X1 U14820 ( .A1(n14756), .A2(n14757), .A3(n14758), .ZN(n14755) );
  INV_X1 U14821 ( .A(n14759), .ZN(n14758) );
  AND2_X1 U14822 ( .A1(n14760), .A2(n14761), .ZN(n14757) );
  INV_X1 U14823 ( .A(n14762), .ZN(n14760) );
  AND2_X1 U14824 ( .A1(n14763), .A2(n14762), .ZN(n14756) );
  OR2_X1 U14825 ( .A1(n14762), .A2(n14759), .ZN(n14754) );
  OR2_X1 U14826 ( .A1(n14764), .A2(n14741), .ZN(Result_7_) );
  AND3_X1 U14827 ( .A1(n14765), .A2(n14766), .A3(n14744), .ZN(n14764) );
  OR3_X1 U14828 ( .A1(n14767), .A2(n14768), .A3(n14769), .ZN(n14766) );
  INV_X1 U14829 ( .A(n14770), .ZN(n14769) );
  AND2_X1 U14830 ( .A1(n14771), .A2(n14772), .ZN(n14768) );
  INV_X1 U14831 ( .A(n14773), .ZN(n14771) );
  AND2_X1 U14832 ( .A1(n14774), .A2(n14773), .ZN(n14767) );
  OR2_X1 U14833 ( .A1(n14773), .A2(n14770), .ZN(n14765) );
  OR2_X1 U14834 ( .A1(n14775), .A2(n14741), .ZN(Result_6_) );
  AND3_X1 U14835 ( .A1(n14776), .A2(n14777), .A3(n14744), .ZN(n14775) );
  OR3_X1 U14836 ( .A1(n14778), .A2(n14779), .A3(n14780), .ZN(n14777) );
  INV_X1 U14837 ( .A(n14781), .ZN(n14780) );
  AND2_X1 U14838 ( .A1(n14782), .A2(n14783), .ZN(n14779) );
  INV_X1 U14839 ( .A(n14784), .ZN(n14782) );
  AND2_X1 U14840 ( .A1(n14785), .A2(n14784), .ZN(n14778) );
  OR2_X1 U14841 ( .A1(n14784), .A2(n14781), .ZN(n14776) );
  OR2_X1 U14842 ( .A1(n14786), .A2(n14787), .ZN(Result_63_) );
  AND2_X1 U14843 ( .A1(n14788), .A2(n14744), .ZN(n14787) );
  AND2_X1 U14844 ( .A1(n14789), .A2(n14790), .ZN(n14786) );
  OR3_X1 U14845 ( .A1(n14791), .A2(n14792), .A3(n14793), .ZN(n14790) );
  OR2_X1 U14846 ( .A1(n14794), .A2(n14795), .ZN(n14789) );
  OR4_X1 U14847 ( .A1(n14796), .A2(n14797), .A3(n14798), .A4(n14799), .ZN(
        Result_62_) );
  AND2_X1 U14848 ( .A1(n14800), .A2(n14801), .ZN(n14799) );
  OR2_X1 U14849 ( .A1(n14802), .A2(n14803), .ZN(n14800) );
  AND2_X1 U14850 ( .A1(a_30_), .A2(n14804), .ZN(n14803) );
  AND2_X1 U14851 ( .A1(n14805), .A2(n14806), .ZN(n14802) );
  AND2_X1 U14852 ( .A1(b_30_), .A2(n14807), .ZN(n14798) );
  OR2_X1 U14853 ( .A1(n14808), .A2(n14809), .ZN(n14807) );
  AND2_X1 U14854 ( .A1(n14804), .A2(n14806), .ZN(n14809) );
  OR3_X1 U14855 ( .A1(n14810), .A2(n14811), .A3(n14812), .ZN(n14804) );
  AND2_X1 U14856 ( .A1(n14791), .A2(n14813), .ZN(n14812) );
  AND2_X1 U14857 ( .A1(n14792), .A2(n14814), .ZN(n14811) );
  AND2_X1 U14858 ( .A1(n14793), .A2(n14815), .ZN(n14810) );
  AND2_X1 U14859 ( .A1(n14744), .A2(n14816), .ZN(n14808) );
  OR2_X1 U14860 ( .A1(n14794), .A2(n14817), .ZN(n14816) );
  AND2_X1 U14861 ( .A1(n14818), .A2(n14805), .ZN(n14797) );
  OR3_X1 U14862 ( .A1(n14819), .A2(n14820), .A3(n14821), .ZN(n14805) );
  AND2_X1 U14863 ( .A1(n14791), .A2(n14795), .ZN(n14821) );
  AND2_X1 U14864 ( .A1(n14792), .A2(n14794), .ZN(n14820) );
  AND2_X1 U14865 ( .A1(n14793), .A2(n14788), .ZN(n14819) );
  AND3_X1 U14866 ( .A1(a_30_), .A2(n14822), .A3(n14744), .ZN(n14796) );
  OR2_X1 U14867 ( .A1(n14823), .A2(n14795), .ZN(n14822) );
  AND2_X1 U14868 ( .A1(b_31_), .A2(n14801), .ZN(n14823) );
  OR3_X1 U14869 ( .A1(n14824), .A2(n14825), .A3(n14826), .ZN(Result_61_) );
  AND3_X1 U14870 ( .A1(n14827), .A2(n14828), .A3(n14744), .ZN(n14826) );
  OR2_X1 U14871 ( .A1(n14829), .A2(n14830), .ZN(n14828) );
  AND2_X1 U14872 ( .A1(n14831), .A2(n14832), .ZN(n14830) );
  INV_X1 U14873 ( .A(n14833), .ZN(n14827) );
  AND3_X1 U14874 ( .A1(n14832), .A2(n14831), .A3(n14829), .ZN(n14833) );
  OR2_X1 U14875 ( .A1(n14834), .A2(n14835), .ZN(n14831) );
  OR2_X1 U14876 ( .A1(n14836), .A2(n14837), .ZN(n14832) );
  AND2_X1 U14877 ( .A1(n14838), .A2(n14839), .ZN(n14825) );
  OR3_X1 U14878 ( .A1(n14840), .A2(n14841), .A3(n14842), .ZN(n14839) );
  AND2_X1 U14879 ( .A1(n14791), .A2(n14843), .ZN(n14842) );
  AND2_X1 U14880 ( .A1(n14792), .A2(n14844), .ZN(n14841) );
  AND2_X1 U14881 ( .A1(n14793), .A2(n14845), .ZN(n14840) );
  INV_X1 U14882 ( .A(n14846), .ZN(n14838) );
  AND2_X1 U14883 ( .A1(n14846), .A2(n14847), .ZN(n14824) );
  OR3_X1 U14884 ( .A1(n14848), .A2(n14849), .A3(n14850), .ZN(n14847) );
  AND2_X1 U14885 ( .A1(n14791), .A2(n14851), .ZN(n14850) );
  INV_X1 U14886 ( .A(n14843), .ZN(n14851) );
  AND2_X1 U14887 ( .A1(n14792), .A2(n14852), .ZN(n14849) );
  INV_X1 U14888 ( .A(n14844), .ZN(n14852) );
  AND2_X1 U14889 ( .A1(n14853), .A2(n14793), .ZN(n14848) );
  OR2_X1 U14890 ( .A1(n14854), .A2(n14855), .ZN(n14846) );
  AND2_X1 U14891 ( .A1(a_29_), .A2(n14856), .ZN(n14855) );
  AND2_X1 U14892 ( .A1(b_29_), .A2(n14857), .ZN(n14854) );
  OR3_X1 U14893 ( .A1(n14858), .A2(n14859), .A3(n14860), .ZN(Result_60_) );
  AND3_X1 U14894 ( .A1(n14861), .A2(n14862), .A3(n14744), .ZN(n14860) );
  INV_X1 U14895 ( .A(n14863), .ZN(n14862) );
  AND2_X1 U14896 ( .A1(n14864), .A2(n14865), .ZN(n14863) );
  OR2_X1 U14897 ( .A1(n14865), .A2(n14864), .ZN(n14861) );
  AND2_X1 U14898 ( .A1(n14866), .A2(n14867), .ZN(n14864) );
  OR2_X1 U14899 ( .A1(n14868), .A2(n14869), .ZN(n14867) );
  INV_X1 U14900 ( .A(n14870), .ZN(n14869) );
  OR2_X1 U14901 ( .A1(n14870), .A2(n14871), .ZN(n14866) );
  INV_X1 U14902 ( .A(n14868), .ZN(n14871) );
  AND2_X1 U14903 ( .A1(n14872), .A2(n14873), .ZN(n14859) );
  OR3_X1 U14904 ( .A1(n14874), .A2(n14875), .A3(n14876), .ZN(n14873) );
  AND2_X1 U14905 ( .A1(n14791), .A2(n14877), .ZN(n14876) );
  AND2_X1 U14906 ( .A1(n14792), .A2(n14878), .ZN(n14875) );
  AND2_X1 U14907 ( .A1(n14879), .A2(n14793), .ZN(n14874) );
  INV_X1 U14908 ( .A(n14880), .ZN(n14879) );
  INV_X1 U14909 ( .A(n14881), .ZN(n14872) );
  AND2_X1 U14910 ( .A1(n14881), .A2(n14882), .ZN(n14858) );
  OR3_X1 U14911 ( .A1(n14883), .A2(n14884), .A3(n14885), .ZN(n14882) );
  AND2_X1 U14912 ( .A1(n14791), .A2(n14886), .ZN(n14885) );
  INV_X1 U14913 ( .A(n14877), .ZN(n14886) );
  AND2_X1 U14914 ( .A1(n14792), .A2(n14887), .ZN(n14884) );
  INV_X1 U14915 ( .A(n14878), .ZN(n14887) );
  AND2_X1 U14916 ( .A1(n14793), .A2(n14880), .ZN(n14883) );
  OR2_X1 U14917 ( .A1(n14888), .A2(n14889), .ZN(n14881) );
  AND2_X1 U14918 ( .A1(a_28_), .A2(n14890), .ZN(n14889) );
  AND2_X1 U14919 ( .A1(b_28_), .A2(n14891), .ZN(n14888) );
  OR2_X1 U14920 ( .A1(n14892), .A2(n14741), .ZN(Result_5_) );
  AND3_X1 U14921 ( .A1(n14893), .A2(n14894), .A3(n14744), .ZN(n14892) );
  OR3_X1 U14922 ( .A1(n14895), .A2(n14896), .A3(n14897), .ZN(n14894) );
  INV_X1 U14923 ( .A(n14898), .ZN(n14897) );
  AND2_X1 U14924 ( .A1(n14899), .A2(n14900), .ZN(n14896) );
  INV_X1 U14925 ( .A(n14901), .ZN(n14899) );
  AND2_X1 U14926 ( .A1(n14902), .A2(n14901), .ZN(n14895) );
  OR2_X1 U14927 ( .A1(n14901), .A2(n14898), .ZN(n14893) );
  OR3_X1 U14928 ( .A1(n14903), .A2(n14904), .A3(n14905), .ZN(Result_59_) );
  AND3_X1 U14929 ( .A1(n14906), .A2(n14907), .A3(n14744), .ZN(n14905) );
  INV_X1 U14930 ( .A(n14908), .ZN(n14907) );
  AND2_X1 U14931 ( .A1(n14909), .A2(n14910), .ZN(n14908) );
  OR2_X1 U14932 ( .A1(n14910), .A2(n14909), .ZN(n14906) );
  AND2_X1 U14933 ( .A1(n14911), .A2(n14912), .ZN(n14909) );
  OR2_X1 U14934 ( .A1(n14913), .A2(n14914), .ZN(n14912) );
  INV_X1 U14935 ( .A(n14915), .ZN(n14914) );
  OR2_X1 U14936 ( .A1(n14915), .A2(n14916), .ZN(n14911) );
  INV_X1 U14937 ( .A(n14913), .ZN(n14916) );
  AND2_X1 U14938 ( .A1(n14917), .A2(n14918), .ZN(n14904) );
  OR3_X1 U14939 ( .A1(n14919), .A2(n14920), .A3(n14921), .ZN(n14918) );
  AND2_X1 U14940 ( .A1(n14791), .A2(n14922), .ZN(n14921) );
  AND2_X1 U14941 ( .A1(n14792), .A2(n14923), .ZN(n14920) );
  AND2_X1 U14942 ( .A1(n14924), .A2(n14793), .ZN(n14919) );
  INV_X1 U14943 ( .A(n14925), .ZN(n14924) );
  INV_X1 U14944 ( .A(n14926), .ZN(n14917) );
  AND2_X1 U14945 ( .A1(n14926), .A2(n14927), .ZN(n14903) );
  OR3_X1 U14946 ( .A1(n14928), .A2(n14929), .A3(n14930), .ZN(n14927) );
  AND2_X1 U14947 ( .A1(n14791), .A2(n14931), .ZN(n14930) );
  INV_X1 U14948 ( .A(n14922), .ZN(n14931) );
  AND2_X1 U14949 ( .A1(n14792), .A2(n14932), .ZN(n14929) );
  INV_X1 U14950 ( .A(n14923), .ZN(n14932) );
  AND2_X1 U14951 ( .A1(n14793), .A2(n14925), .ZN(n14928) );
  OR2_X1 U14952 ( .A1(n14933), .A2(n14934), .ZN(n14926) );
  AND2_X1 U14953 ( .A1(a_27_), .A2(n14935), .ZN(n14934) );
  AND2_X1 U14954 ( .A1(b_27_), .A2(n14936), .ZN(n14933) );
  OR3_X1 U14955 ( .A1(n14937), .A2(n14938), .A3(n14939), .ZN(Result_58_) );
  AND3_X1 U14956 ( .A1(n14940), .A2(n14941), .A3(n14744), .ZN(n14939) );
  INV_X1 U14957 ( .A(n14942), .ZN(n14941) );
  AND2_X1 U14958 ( .A1(n14943), .A2(n14944), .ZN(n14942) );
  OR2_X1 U14959 ( .A1(n14944), .A2(n14943), .ZN(n14940) );
  AND2_X1 U14960 ( .A1(n14945), .A2(n14946), .ZN(n14943) );
  OR2_X1 U14961 ( .A1(n14947), .A2(n14948), .ZN(n14946) );
  INV_X1 U14962 ( .A(n14949), .ZN(n14948) );
  OR2_X1 U14963 ( .A1(n14949), .A2(n14950), .ZN(n14945) );
  INV_X1 U14964 ( .A(n14947), .ZN(n14950) );
  AND2_X1 U14965 ( .A1(n14951), .A2(n14952), .ZN(n14938) );
  OR3_X1 U14966 ( .A1(n14953), .A2(n14954), .A3(n14955), .ZN(n14952) );
  AND2_X1 U14967 ( .A1(n14791), .A2(n14956), .ZN(n14955) );
  AND2_X1 U14968 ( .A1(n14792), .A2(n14957), .ZN(n14954) );
  AND2_X1 U14969 ( .A1(n14958), .A2(n14793), .ZN(n14953) );
  INV_X1 U14970 ( .A(n14959), .ZN(n14958) );
  INV_X1 U14971 ( .A(n14960), .ZN(n14951) );
  AND2_X1 U14972 ( .A1(n14960), .A2(n14961), .ZN(n14937) );
  OR3_X1 U14973 ( .A1(n14962), .A2(n14963), .A3(n14964), .ZN(n14961) );
  AND2_X1 U14974 ( .A1(n14791), .A2(n14965), .ZN(n14964) );
  INV_X1 U14975 ( .A(n14956), .ZN(n14965) );
  AND2_X1 U14976 ( .A1(n14792), .A2(n14966), .ZN(n14963) );
  INV_X1 U14977 ( .A(n14957), .ZN(n14966) );
  AND2_X1 U14978 ( .A1(n14793), .A2(n14959), .ZN(n14962) );
  OR2_X1 U14979 ( .A1(n14967), .A2(n14968), .ZN(n14960) );
  AND2_X1 U14980 ( .A1(a_26_), .A2(n14969), .ZN(n14968) );
  AND2_X1 U14981 ( .A1(b_26_), .A2(n14970), .ZN(n14967) );
  OR3_X1 U14982 ( .A1(n14971), .A2(n14972), .A3(n14973), .ZN(Result_57_) );
  AND3_X1 U14983 ( .A1(n14974), .A2(n14975), .A3(n14744), .ZN(n14973) );
  INV_X1 U14984 ( .A(n14976), .ZN(n14975) );
  AND2_X1 U14985 ( .A1(n14977), .A2(n14978), .ZN(n14976) );
  OR2_X1 U14986 ( .A1(n14978), .A2(n14977), .ZN(n14974) );
  AND2_X1 U14987 ( .A1(n14979), .A2(n14980), .ZN(n14977) );
  OR2_X1 U14988 ( .A1(n14981), .A2(n14982), .ZN(n14980) );
  INV_X1 U14989 ( .A(n14983), .ZN(n14982) );
  OR2_X1 U14990 ( .A1(n14983), .A2(n14984), .ZN(n14979) );
  INV_X1 U14991 ( .A(n14981), .ZN(n14984) );
  AND2_X1 U14992 ( .A1(n14985), .A2(n14986), .ZN(n14972) );
  OR3_X1 U14993 ( .A1(n14987), .A2(n14988), .A3(n14989), .ZN(n14986) );
  AND2_X1 U14994 ( .A1(n14791), .A2(n14990), .ZN(n14989) );
  AND2_X1 U14995 ( .A1(n14792), .A2(n14991), .ZN(n14988) );
  AND2_X1 U14996 ( .A1(n14992), .A2(n14793), .ZN(n14987) );
  INV_X1 U14997 ( .A(n14993), .ZN(n14992) );
  INV_X1 U14998 ( .A(n14994), .ZN(n14985) );
  AND2_X1 U14999 ( .A1(n14994), .A2(n14995), .ZN(n14971) );
  OR3_X1 U15000 ( .A1(n14996), .A2(n14997), .A3(n14998), .ZN(n14995) );
  AND2_X1 U15001 ( .A1(n14791), .A2(n14999), .ZN(n14998) );
  INV_X1 U15002 ( .A(n14990), .ZN(n14999) );
  AND2_X1 U15003 ( .A1(n14792), .A2(n15000), .ZN(n14997) );
  INV_X1 U15004 ( .A(n14991), .ZN(n15000) );
  AND2_X1 U15005 ( .A1(n14793), .A2(n14993), .ZN(n14996) );
  OR2_X1 U15006 ( .A1(n15001), .A2(n15002), .ZN(n14994) );
  AND2_X1 U15007 ( .A1(a_25_), .A2(n15003), .ZN(n15002) );
  AND2_X1 U15008 ( .A1(b_25_), .A2(n15004), .ZN(n15001) );
  OR3_X1 U15009 ( .A1(n15005), .A2(n15006), .A3(n15007), .ZN(Result_56_) );
  AND3_X1 U15010 ( .A1(n15008), .A2(n15009), .A3(n14744), .ZN(n15007) );
  INV_X1 U15011 ( .A(n15010), .ZN(n15009) );
  AND2_X1 U15012 ( .A1(n15011), .A2(n15012), .ZN(n15010) );
  OR2_X1 U15013 ( .A1(n15012), .A2(n15011), .ZN(n15008) );
  AND2_X1 U15014 ( .A1(n15013), .A2(n15014), .ZN(n15011) );
  OR2_X1 U15015 ( .A1(n15015), .A2(n15016), .ZN(n15014) );
  INV_X1 U15016 ( .A(n15017), .ZN(n15016) );
  OR2_X1 U15017 ( .A1(n15017), .A2(n15018), .ZN(n15013) );
  INV_X1 U15018 ( .A(n15015), .ZN(n15018) );
  AND2_X1 U15019 ( .A1(n15019), .A2(n15020), .ZN(n15006) );
  OR3_X1 U15020 ( .A1(n15021), .A2(n15022), .A3(n15023), .ZN(n15020) );
  AND2_X1 U15021 ( .A1(n14791), .A2(n15024), .ZN(n15023) );
  AND2_X1 U15022 ( .A1(n14792), .A2(n15025), .ZN(n15022) );
  AND2_X1 U15023 ( .A1(n15026), .A2(n14793), .ZN(n15021) );
  INV_X1 U15024 ( .A(n15027), .ZN(n15026) );
  INV_X1 U15025 ( .A(n15028), .ZN(n15019) );
  AND2_X1 U15026 ( .A1(n15028), .A2(n15029), .ZN(n15005) );
  OR3_X1 U15027 ( .A1(n15030), .A2(n15031), .A3(n15032), .ZN(n15029) );
  AND2_X1 U15028 ( .A1(n14791), .A2(n15033), .ZN(n15032) );
  INV_X1 U15029 ( .A(n15024), .ZN(n15033) );
  AND2_X1 U15030 ( .A1(n14792), .A2(n15034), .ZN(n15031) );
  INV_X1 U15031 ( .A(n15025), .ZN(n15034) );
  AND2_X1 U15032 ( .A1(n14793), .A2(n15027), .ZN(n15030) );
  OR2_X1 U15033 ( .A1(n15035), .A2(n15036), .ZN(n15028) );
  AND2_X1 U15034 ( .A1(a_24_), .A2(n15037), .ZN(n15036) );
  AND2_X1 U15035 ( .A1(b_24_), .A2(n15038), .ZN(n15035) );
  OR3_X1 U15036 ( .A1(n15039), .A2(n15040), .A3(n15041), .ZN(Result_55_) );
  AND3_X1 U15037 ( .A1(n15042), .A2(n15043), .A3(n14744), .ZN(n15041) );
  INV_X1 U15038 ( .A(n15044), .ZN(n15043) );
  AND2_X1 U15039 ( .A1(n15045), .A2(n15046), .ZN(n15044) );
  OR2_X1 U15040 ( .A1(n15046), .A2(n15045), .ZN(n15042) );
  AND2_X1 U15041 ( .A1(n15047), .A2(n15048), .ZN(n15045) );
  OR2_X1 U15042 ( .A1(n15049), .A2(n15050), .ZN(n15048) );
  INV_X1 U15043 ( .A(n15051), .ZN(n15050) );
  OR2_X1 U15044 ( .A1(n15051), .A2(n15052), .ZN(n15047) );
  INV_X1 U15045 ( .A(n15049), .ZN(n15052) );
  AND2_X1 U15046 ( .A1(n15053), .A2(n15054), .ZN(n15040) );
  OR3_X1 U15047 ( .A1(n15055), .A2(n15056), .A3(n15057), .ZN(n15054) );
  AND2_X1 U15048 ( .A1(n14791), .A2(n15058), .ZN(n15057) );
  AND2_X1 U15049 ( .A1(n14792), .A2(n15059), .ZN(n15056) );
  AND2_X1 U15050 ( .A1(n15060), .A2(n14793), .ZN(n15055) );
  INV_X1 U15051 ( .A(n15061), .ZN(n15060) );
  INV_X1 U15052 ( .A(n15062), .ZN(n15053) );
  AND2_X1 U15053 ( .A1(n15062), .A2(n15063), .ZN(n15039) );
  OR3_X1 U15054 ( .A1(n15064), .A2(n15065), .A3(n15066), .ZN(n15063) );
  AND2_X1 U15055 ( .A1(n14791), .A2(n15067), .ZN(n15066) );
  INV_X1 U15056 ( .A(n15058), .ZN(n15067) );
  AND2_X1 U15057 ( .A1(n14792), .A2(n15068), .ZN(n15065) );
  INV_X1 U15058 ( .A(n15059), .ZN(n15068) );
  AND2_X1 U15059 ( .A1(n14793), .A2(n15061), .ZN(n15064) );
  OR2_X1 U15060 ( .A1(n15069), .A2(n15070), .ZN(n15062) );
  AND2_X1 U15061 ( .A1(a_23_), .A2(n15071), .ZN(n15070) );
  AND2_X1 U15062 ( .A1(b_23_), .A2(n15072), .ZN(n15069) );
  OR3_X1 U15063 ( .A1(n15073), .A2(n15074), .A3(n15075), .ZN(Result_54_) );
  AND3_X1 U15064 ( .A1(n15076), .A2(n15077), .A3(n14744), .ZN(n15075) );
  INV_X1 U15065 ( .A(n15078), .ZN(n15077) );
  AND2_X1 U15066 ( .A1(n15079), .A2(n15080), .ZN(n15078) );
  OR2_X1 U15067 ( .A1(n15080), .A2(n15079), .ZN(n15076) );
  AND2_X1 U15068 ( .A1(n15081), .A2(n15082), .ZN(n15079) );
  OR2_X1 U15069 ( .A1(n15083), .A2(n15084), .ZN(n15082) );
  INV_X1 U15070 ( .A(n15085), .ZN(n15084) );
  OR2_X1 U15071 ( .A1(n15085), .A2(n15086), .ZN(n15081) );
  INV_X1 U15072 ( .A(n15083), .ZN(n15086) );
  AND2_X1 U15073 ( .A1(n15087), .A2(n15088), .ZN(n15074) );
  OR3_X1 U15074 ( .A1(n15089), .A2(n15090), .A3(n15091), .ZN(n15088) );
  AND2_X1 U15075 ( .A1(n14791), .A2(n15092), .ZN(n15091) );
  AND2_X1 U15076 ( .A1(n14792), .A2(n15093), .ZN(n15090) );
  AND2_X1 U15077 ( .A1(n15094), .A2(n14793), .ZN(n15089) );
  INV_X1 U15078 ( .A(n15095), .ZN(n15094) );
  INV_X1 U15079 ( .A(n15096), .ZN(n15087) );
  AND2_X1 U15080 ( .A1(n15096), .A2(n15097), .ZN(n15073) );
  OR3_X1 U15081 ( .A1(n15098), .A2(n15099), .A3(n15100), .ZN(n15097) );
  AND2_X1 U15082 ( .A1(n14791), .A2(n15101), .ZN(n15100) );
  INV_X1 U15083 ( .A(n15092), .ZN(n15101) );
  AND2_X1 U15084 ( .A1(n14792), .A2(n15102), .ZN(n15099) );
  INV_X1 U15085 ( .A(n15093), .ZN(n15102) );
  AND2_X1 U15086 ( .A1(n14793), .A2(n15095), .ZN(n15098) );
  OR2_X1 U15087 ( .A1(n15103), .A2(n15104), .ZN(n15096) );
  AND2_X1 U15088 ( .A1(a_22_), .A2(n15105), .ZN(n15104) );
  AND2_X1 U15089 ( .A1(b_22_), .A2(n15106), .ZN(n15103) );
  OR3_X1 U15090 ( .A1(n15107), .A2(n15108), .A3(n15109), .ZN(Result_53_) );
  AND3_X1 U15091 ( .A1(n15110), .A2(n15111), .A3(n14744), .ZN(n15109) );
  INV_X1 U15092 ( .A(n15112), .ZN(n15111) );
  AND2_X1 U15093 ( .A1(n15113), .A2(n15114), .ZN(n15112) );
  OR2_X1 U15094 ( .A1(n15114), .A2(n15113), .ZN(n15110) );
  AND2_X1 U15095 ( .A1(n15115), .A2(n15116), .ZN(n15113) );
  OR2_X1 U15096 ( .A1(n15117), .A2(n15118), .ZN(n15116) );
  INV_X1 U15097 ( .A(n15119), .ZN(n15118) );
  OR2_X1 U15098 ( .A1(n15119), .A2(n15120), .ZN(n15115) );
  INV_X1 U15099 ( .A(n15117), .ZN(n15120) );
  AND2_X1 U15100 ( .A1(n15121), .A2(n15122), .ZN(n15108) );
  OR3_X1 U15101 ( .A1(n15123), .A2(n15124), .A3(n15125), .ZN(n15122) );
  AND2_X1 U15102 ( .A1(n14791), .A2(n15126), .ZN(n15125) );
  AND2_X1 U15103 ( .A1(n14792), .A2(n15127), .ZN(n15124) );
  AND2_X1 U15104 ( .A1(n15128), .A2(n14793), .ZN(n15123) );
  INV_X1 U15105 ( .A(n15129), .ZN(n15128) );
  INV_X1 U15106 ( .A(n15130), .ZN(n15121) );
  AND2_X1 U15107 ( .A1(n15130), .A2(n15131), .ZN(n15107) );
  OR3_X1 U15108 ( .A1(n15132), .A2(n15133), .A3(n15134), .ZN(n15131) );
  AND2_X1 U15109 ( .A1(n14791), .A2(n15135), .ZN(n15134) );
  INV_X1 U15110 ( .A(n15126), .ZN(n15135) );
  AND2_X1 U15111 ( .A1(n14792), .A2(n15136), .ZN(n15133) );
  INV_X1 U15112 ( .A(n15127), .ZN(n15136) );
  AND2_X1 U15113 ( .A1(n14793), .A2(n15129), .ZN(n15132) );
  OR2_X1 U15114 ( .A1(n15137), .A2(n15138), .ZN(n15130) );
  AND2_X1 U15115 ( .A1(a_21_), .A2(n15139), .ZN(n15138) );
  AND2_X1 U15116 ( .A1(b_21_), .A2(n15140), .ZN(n15137) );
  OR3_X1 U15117 ( .A1(n15141), .A2(n15142), .A3(n15143), .ZN(Result_52_) );
  AND3_X1 U15118 ( .A1(n15144), .A2(n15145), .A3(n14744), .ZN(n15143) );
  INV_X1 U15119 ( .A(n15146), .ZN(n15145) );
  AND2_X1 U15120 ( .A1(n15147), .A2(n15148), .ZN(n15146) );
  OR2_X1 U15121 ( .A1(n15148), .A2(n15147), .ZN(n15144) );
  AND2_X1 U15122 ( .A1(n15149), .A2(n15150), .ZN(n15147) );
  OR2_X1 U15123 ( .A1(n15151), .A2(n15152), .ZN(n15150) );
  INV_X1 U15124 ( .A(n15153), .ZN(n15152) );
  OR2_X1 U15125 ( .A1(n15153), .A2(n15154), .ZN(n15149) );
  INV_X1 U15126 ( .A(n15151), .ZN(n15154) );
  AND2_X1 U15127 ( .A1(n15155), .A2(n15156), .ZN(n15142) );
  OR3_X1 U15128 ( .A1(n15157), .A2(n15158), .A3(n15159), .ZN(n15156) );
  AND2_X1 U15129 ( .A1(n14791), .A2(n15160), .ZN(n15159) );
  AND2_X1 U15130 ( .A1(n14792), .A2(n15161), .ZN(n15158) );
  AND2_X1 U15131 ( .A1(n15162), .A2(n14793), .ZN(n15157) );
  INV_X1 U15132 ( .A(n15163), .ZN(n15162) );
  INV_X1 U15133 ( .A(n15164), .ZN(n15155) );
  AND2_X1 U15134 ( .A1(n15164), .A2(n15165), .ZN(n15141) );
  OR3_X1 U15135 ( .A1(n15166), .A2(n15167), .A3(n15168), .ZN(n15165) );
  AND2_X1 U15136 ( .A1(n14791), .A2(n15169), .ZN(n15168) );
  INV_X1 U15137 ( .A(n15160), .ZN(n15169) );
  AND2_X1 U15138 ( .A1(n14792), .A2(n15170), .ZN(n15167) );
  INV_X1 U15139 ( .A(n15161), .ZN(n15170) );
  AND2_X1 U15140 ( .A1(n14793), .A2(n15163), .ZN(n15166) );
  OR2_X1 U15141 ( .A1(n15171), .A2(n15172), .ZN(n15164) );
  AND2_X1 U15142 ( .A1(a_20_), .A2(n15173), .ZN(n15172) );
  AND2_X1 U15143 ( .A1(b_20_), .A2(n15174), .ZN(n15171) );
  OR3_X1 U15144 ( .A1(n15175), .A2(n15176), .A3(n15177), .ZN(Result_51_) );
  AND3_X1 U15145 ( .A1(n15178), .A2(n15179), .A3(n14744), .ZN(n15177) );
  INV_X1 U15146 ( .A(n15180), .ZN(n15179) );
  AND2_X1 U15147 ( .A1(n15181), .A2(n15182), .ZN(n15180) );
  OR2_X1 U15148 ( .A1(n15182), .A2(n15181), .ZN(n15178) );
  AND2_X1 U15149 ( .A1(n15183), .A2(n15184), .ZN(n15181) );
  OR2_X1 U15150 ( .A1(n15185), .A2(n15186), .ZN(n15184) );
  INV_X1 U15151 ( .A(n15187), .ZN(n15186) );
  OR2_X1 U15152 ( .A1(n15187), .A2(n15188), .ZN(n15183) );
  INV_X1 U15153 ( .A(n15185), .ZN(n15188) );
  AND2_X1 U15154 ( .A1(n15189), .A2(n15190), .ZN(n15176) );
  OR3_X1 U15155 ( .A1(n15191), .A2(n15192), .A3(n15193), .ZN(n15190) );
  AND2_X1 U15156 ( .A1(n14791), .A2(n15194), .ZN(n15193) );
  AND2_X1 U15157 ( .A1(n14792), .A2(n15195), .ZN(n15192) );
  AND2_X1 U15158 ( .A1(n15196), .A2(n14793), .ZN(n15191) );
  INV_X1 U15159 ( .A(n15197), .ZN(n15196) );
  INV_X1 U15160 ( .A(n15198), .ZN(n15189) );
  AND2_X1 U15161 ( .A1(n15198), .A2(n15199), .ZN(n15175) );
  OR3_X1 U15162 ( .A1(n15200), .A2(n15201), .A3(n15202), .ZN(n15199) );
  AND2_X1 U15163 ( .A1(n14791), .A2(n15203), .ZN(n15202) );
  INV_X1 U15164 ( .A(n15194), .ZN(n15203) );
  AND2_X1 U15165 ( .A1(n14792), .A2(n15204), .ZN(n15201) );
  INV_X1 U15166 ( .A(n15195), .ZN(n15204) );
  AND2_X1 U15167 ( .A1(n14793), .A2(n15197), .ZN(n15200) );
  OR2_X1 U15168 ( .A1(n15205), .A2(n15206), .ZN(n15198) );
  AND2_X1 U15169 ( .A1(a_19_), .A2(n15207), .ZN(n15206) );
  AND2_X1 U15170 ( .A1(b_19_), .A2(n15208), .ZN(n15205) );
  OR3_X1 U15171 ( .A1(n15209), .A2(n15210), .A3(n15211), .ZN(Result_50_) );
  AND3_X1 U15172 ( .A1(n15212), .A2(n15213), .A3(n14744), .ZN(n15211) );
  INV_X1 U15173 ( .A(n15214), .ZN(n15213) );
  AND2_X1 U15174 ( .A1(n15215), .A2(n15216), .ZN(n15214) );
  OR2_X1 U15175 ( .A1(n15216), .A2(n15215), .ZN(n15212) );
  AND2_X1 U15176 ( .A1(n15217), .A2(n15218), .ZN(n15215) );
  OR2_X1 U15177 ( .A1(n15219), .A2(n15220), .ZN(n15218) );
  INV_X1 U15178 ( .A(n15221), .ZN(n15220) );
  OR2_X1 U15179 ( .A1(n15221), .A2(n15222), .ZN(n15217) );
  INV_X1 U15180 ( .A(n15219), .ZN(n15222) );
  AND2_X1 U15181 ( .A1(n15223), .A2(n15224), .ZN(n15210) );
  OR3_X1 U15182 ( .A1(n15225), .A2(n15226), .A3(n15227), .ZN(n15224) );
  AND2_X1 U15183 ( .A1(n14791), .A2(n15228), .ZN(n15227) );
  AND2_X1 U15184 ( .A1(n14792), .A2(n15229), .ZN(n15226) );
  AND2_X1 U15185 ( .A1(n15230), .A2(n14793), .ZN(n15225) );
  INV_X1 U15186 ( .A(n15231), .ZN(n15230) );
  INV_X1 U15187 ( .A(n15232), .ZN(n15223) );
  AND2_X1 U15188 ( .A1(n15232), .A2(n15233), .ZN(n15209) );
  OR3_X1 U15189 ( .A1(n15234), .A2(n15235), .A3(n15236), .ZN(n15233) );
  AND2_X1 U15190 ( .A1(n14791), .A2(n15237), .ZN(n15236) );
  INV_X1 U15191 ( .A(n15228), .ZN(n15237) );
  AND2_X1 U15192 ( .A1(n14792), .A2(n15238), .ZN(n15235) );
  INV_X1 U15193 ( .A(n15229), .ZN(n15238) );
  AND2_X1 U15194 ( .A1(n14793), .A2(n15231), .ZN(n15234) );
  OR2_X1 U15195 ( .A1(n15239), .A2(n15240), .ZN(n15232) );
  AND2_X1 U15196 ( .A1(a_18_), .A2(n15241), .ZN(n15240) );
  AND2_X1 U15197 ( .A1(b_18_), .A2(n15242), .ZN(n15239) );
  OR2_X1 U15198 ( .A1(n15243), .A2(n14741), .ZN(Result_4_) );
  AND3_X1 U15199 ( .A1(n15244), .A2(n15245), .A3(n14744), .ZN(n15243) );
  OR3_X1 U15200 ( .A1(n15246), .A2(n15247), .A3(n15248), .ZN(n15245) );
  INV_X1 U15201 ( .A(n15249), .ZN(n15248) );
  AND2_X1 U15202 ( .A1(n15250), .A2(n15251), .ZN(n15247) );
  INV_X1 U15203 ( .A(n15252), .ZN(n15250) );
  AND2_X1 U15204 ( .A1(n15253), .A2(n15252), .ZN(n15246) );
  OR2_X1 U15205 ( .A1(n15252), .A2(n15249), .ZN(n15244) );
  OR3_X1 U15206 ( .A1(n15254), .A2(n15255), .A3(n15256), .ZN(Result_49_) );
  AND3_X1 U15207 ( .A1(n15257), .A2(n15258), .A3(n14744), .ZN(n15256) );
  INV_X1 U15208 ( .A(n15259), .ZN(n15258) );
  AND2_X1 U15209 ( .A1(n15260), .A2(n15261), .ZN(n15259) );
  OR2_X1 U15210 ( .A1(n15261), .A2(n15260), .ZN(n15257) );
  AND2_X1 U15211 ( .A1(n15262), .A2(n15263), .ZN(n15260) );
  OR2_X1 U15212 ( .A1(n15264), .A2(n15265), .ZN(n15263) );
  INV_X1 U15213 ( .A(n15266), .ZN(n15265) );
  OR2_X1 U15214 ( .A1(n15266), .A2(n15267), .ZN(n15262) );
  INV_X1 U15215 ( .A(n15264), .ZN(n15267) );
  AND2_X1 U15216 ( .A1(n15268), .A2(n15269), .ZN(n15255) );
  OR3_X1 U15217 ( .A1(n15270), .A2(n15271), .A3(n15272), .ZN(n15269) );
  AND2_X1 U15218 ( .A1(n14791), .A2(n15273), .ZN(n15272) );
  AND2_X1 U15219 ( .A1(n14792), .A2(n15274), .ZN(n15271) );
  AND2_X1 U15220 ( .A1(n15275), .A2(n14793), .ZN(n15270) );
  INV_X1 U15221 ( .A(n15276), .ZN(n15275) );
  INV_X1 U15222 ( .A(n15277), .ZN(n15268) );
  AND2_X1 U15223 ( .A1(n15277), .A2(n15278), .ZN(n15254) );
  OR3_X1 U15224 ( .A1(n15279), .A2(n15280), .A3(n15281), .ZN(n15278) );
  AND2_X1 U15225 ( .A1(n14791), .A2(n15282), .ZN(n15281) );
  INV_X1 U15226 ( .A(n15273), .ZN(n15282) );
  AND2_X1 U15227 ( .A1(n14792), .A2(n15283), .ZN(n15280) );
  INV_X1 U15228 ( .A(n15274), .ZN(n15283) );
  AND2_X1 U15229 ( .A1(n14793), .A2(n15276), .ZN(n15279) );
  OR2_X1 U15230 ( .A1(n15284), .A2(n15285), .ZN(n15277) );
  AND2_X1 U15231 ( .A1(a_17_), .A2(n15286), .ZN(n15285) );
  AND2_X1 U15232 ( .A1(b_17_), .A2(n15287), .ZN(n15284) );
  OR3_X1 U15233 ( .A1(n15288), .A2(n15289), .A3(n15290), .ZN(Result_48_) );
  AND3_X1 U15234 ( .A1(n15291), .A2(n15292), .A3(n14744), .ZN(n15290) );
  INV_X1 U15235 ( .A(n15293), .ZN(n15292) );
  AND2_X1 U15236 ( .A1(n15294), .A2(n15295), .ZN(n15293) );
  OR2_X1 U15237 ( .A1(n15295), .A2(n15294), .ZN(n15291) );
  AND2_X1 U15238 ( .A1(n15296), .A2(n15297), .ZN(n15294) );
  OR2_X1 U15239 ( .A1(n15298), .A2(n15299), .ZN(n15297) );
  INV_X1 U15240 ( .A(n15300), .ZN(n15299) );
  OR2_X1 U15241 ( .A1(n15300), .A2(n15301), .ZN(n15296) );
  INV_X1 U15242 ( .A(n15298), .ZN(n15301) );
  AND2_X1 U15243 ( .A1(n15302), .A2(n15303), .ZN(n15289) );
  OR3_X1 U15244 ( .A1(n15304), .A2(n15305), .A3(n15306), .ZN(n15303) );
  AND2_X1 U15245 ( .A1(n14791), .A2(n15307), .ZN(n15306) );
  AND2_X1 U15246 ( .A1(n14792), .A2(n15308), .ZN(n15305) );
  AND2_X1 U15247 ( .A1(n15309), .A2(n14793), .ZN(n15304) );
  INV_X1 U15248 ( .A(n15310), .ZN(n15309) );
  INV_X1 U15249 ( .A(n15311), .ZN(n15302) );
  AND2_X1 U15250 ( .A1(n15311), .A2(n15312), .ZN(n15288) );
  OR3_X1 U15251 ( .A1(n15313), .A2(n15314), .A3(n15315), .ZN(n15312) );
  AND2_X1 U15252 ( .A1(n14791), .A2(n15316), .ZN(n15315) );
  INV_X1 U15253 ( .A(n15307), .ZN(n15316) );
  AND2_X1 U15254 ( .A1(n14792), .A2(n15317), .ZN(n15314) );
  INV_X1 U15255 ( .A(n15308), .ZN(n15317) );
  AND2_X1 U15256 ( .A1(n14793), .A2(n15310), .ZN(n15313) );
  OR2_X1 U15257 ( .A1(n15318), .A2(n15319), .ZN(n15311) );
  AND2_X1 U15258 ( .A1(a_16_), .A2(n15320), .ZN(n15319) );
  AND2_X1 U15259 ( .A1(b_16_), .A2(n15321), .ZN(n15318) );
  OR3_X1 U15260 ( .A1(n15322), .A2(n15323), .A3(n15324), .ZN(Result_47_) );
  AND3_X1 U15261 ( .A1(n15325), .A2(n15326), .A3(n14744), .ZN(n15324) );
  INV_X1 U15262 ( .A(n15327), .ZN(n15326) );
  AND2_X1 U15263 ( .A1(n15328), .A2(n15329), .ZN(n15327) );
  OR2_X1 U15264 ( .A1(n15329), .A2(n15328), .ZN(n15325) );
  AND2_X1 U15265 ( .A1(n15330), .A2(n15331), .ZN(n15328) );
  OR2_X1 U15266 ( .A1(n15332), .A2(n15333), .ZN(n15331) );
  INV_X1 U15267 ( .A(n15334), .ZN(n15333) );
  OR2_X1 U15268 ( .A1(n15334), .A2(n15335), .ZN(n15330) );
  INV_X1 U15269 ( .A(n15332), .ZN(n15335) );
  AND2_X1 U15270 ( .A1(n15336), .A2(n15337), .ZN(n15323) );
  OR3_X1 U15271 ( .A1(n15338), .A2(n15339), .A3(n15340), .ZN(n15337) );
  AND2_X1 U15272 ( .A1(n14791), .A2(n15341), .ZN(n15340) );
  AND2_X1 U15273 ( .A1(n14792), .A2(n15342), .ZN(n15339) );
  AND2_X1 U15274 ( .A1(n15343), .A2(n14793), .ZN(n15338) );
  INV_X1 U15275 ( .A(n15344), .ZN(n15343) );
  INV_X1 U15276 ( .A(n15345), .ZN(n15336) );
  AND2_X1 U15277 ( .A1(n15345), .A2(n15346), .ZN(n15322) );
  OR3_X1 U15278 ( .A1(n15347), .A2(n15348), .A3(n15349), .ZN(n15346) );
  AND2_X1 U15279 ( .A1(n14791), .A2(n15350), .ZN(n15349) );
  INV_X1 U15280 ( .A(n15341), .ZN(n15350) );
  AND2_X1 U15281 ( .A1(n14792), .A2(n15351), .ZN(n15348) );
  INV_X1 U15282 ( .A(n15342), .ZN(n15351) );
  AND2_X1 U15283 ( .A1(n14793), .A2(n15344), .ZN(n15347) );
  OR2_X1 U15284 ( .A1(n15352), .A2(n15353), .ZN(n15345) );
  AND2_X1 U15285 ( .A1(a_15_), .A2(n15354), .ZN(n15353) );
  AND2_X1 U15286 ( .A1(b_15_), .A2(n15355), .ZN(n15352) );
  OR3_X1 U15287 ( .A1(n15356), .A2(n15357), .A3(n15358), .ZN(Result_46_) );
  AND3_X1 U15288 ( .A1(n15359), .A2(n15360), .A3(n14744), .ZN(n15358) );
  INV_X1 U15289 ( .A(n15361), .ZN(n15360) );
  AND2_X1 U15290 ( .A1(n15362), .A2(n15363), .ZN(n15361) );
  OR2_X1 U15291 ( .A1(n15363), .A2(n15362), .ZN(n15359) );
  AND2_X1 U15292 ( .A1(n15364), .A2(n15365), .ZN(n15362) );
  OR2_X1 U15293 ( .A1(n15366), .A2(n15367), .ZN(n15365) );
  INV_X1 U15294 ( .A(n15368), .ZN(n15367) );
  OR2_X1 U15295 ( .A1(n15368), .A2(n15369), .ZN(n15364) );
  INV_X1 U15296 ( .A(n15366), .ZN(n15369) );
  AND2_X1 U15297 ( .A1(n15370), .A2(n15371), .ZN(n15357) );
  OR3_X1 U15298 ( .A1(n15372), .A2(n15373), .A3(n15374), .ZN(n15371) );
  AND2_X1 U15299 ( .A1(n14791), .A2(n15375), .ZN(n15374) );
  AND2_X1 U15300 ( .A1(n14792), .A2(n15376), .ZN(n15373) );
  AND2_X1 U15301 ( .A1(n15377), .A2(n14793), .ZN(n15372) );
  INV_X1 U15302 ( .A(n15378), .ZN(n15377) );
  INV_X1 U15303 ( .A(n15379), .ZN(n15370) );
  AND2_X1 U15304 ( .A1(n15379), .A2(n15380), .ZN(n15356) );
  OR3_X1 U15305 ( .A1(n15381), .A2(n15382), .A3(n15383), .ZN(n15380) );
  AND2_X1 U15306 ( .A1(n14791), .A2(n15384), .ZN(n15383) );
  INV_X1 U15307 ( .A(n15375), .ZN(n15384) );
  AND2_X1 U15308 ( .A1(n14792), .A2(n15385), .ZN(n15382) );
  INV_X1 U15309 ( .A(n15376), .ZN(n15385) );
  AND2_X1 U15310 ( .A1(n14793), .A2(n15378), .ZN(n15381) );
  OR2_X1 U15311 ( .A1(n15386), .A2(n15387), .ZN(n15379) );
  AND2_X1 U15312 ( .A1(a_14_), .A2(n15388), .ZN(n15387) );
  AND2_X1 U15313 ( .A1(b_14_), .A2(n15389), .ZN(n15386) );
  OR3_X1 U15314 ( .A1(n15390), .A2(n15391), .A3(n15392), .ZN(Result_45_) );
  AND3_X1 U15315 ( .A1(n15393), .A2(n15394), .A3(n14744), .ZN(n15392) );
  INV_X1 U15316 ( .A(n15395), .ZN(n15394) );
  AND2_X1 U15317 ( .A1(n15396), .A2(n15397), .ZN(n15395) );
  OR2_X1 U15318 ( .A1(n15397), .A2(n15396), .ZN(n15393) );
  AND2_X1 U15319 ( .A1(n15398), .A2(n15399), .ZN(n15396) );
  OR2_X1 U15320 ( .A1(n15400), .A2(n15401), .ZN(n15399) );
  INV_X1 U15321 ( .A(n15402), .ZN(n15401) );
  OR2_X1 U15322 ( .A1(n15402), .A2(n15403), .ZN(n15398) );
  INV_X1 U15323 ( .A(n15400), .ZN(n15403) );
  AND2_X1 U15324 ( .A1(n15404), .A2(n15405), .ZN(n15391) );
  OR3_X1 U15325 ( .A1(n15406), .A2(n15407), .A3(n15408), .ZN(n15405) );
  AND2_X1 U15326 ( .A1(n14791), .A2(n15409), .ZN(n15408) );
  AND2_X1 U15327 ( .A1(n14792), .A2(n15410), .ZN(n15407) );
  AND2_X1 U15328 ( .A1(n15411), .A2(n14793), .ZN(n15406) );
  INV_X1 U15329 ( .A(n15412), .ZN(n15411) );
  INV_X1 U15330 ( .A(n15413), .ZN(n15404) );
  AND2_X1 U15331 ( .A1(n15413), .A2(n15414), .ZN(n15390) );
  OR3_X1 U15332 ( .A1(n15415), .A2(n15416), .A3(n15417), .ZN(n15414) );
  AND2_X1 U15333 ( .A1(n14791), .A2(n15418), .ZN(n15417) );
  INV_X1 U15334 ( .A(n15409), .ZN(n15418) );
  AND2_X1 U15335 ( .A1(n14792), .A2(n15419), .ZN(n15416) );
  INV_X1 U15336 ( .A(n15410), .ZN(n15419) );
  AND2_X1 U15337 ( .A1(n14793), .A2(n15412), .ZN(n15415) );
  OR2_X1 U15338 ( .A1(n15420), .A2(n15421), .ZN(n15413) );
  AND2_X1 U15339 ( .A1(a_13_), .A2(n15422), .ZN(n15421) );
  AND2_X1 U15340 ( .A1(b_13_), .A2(n15423), .ZN(n15420) );
  OR3_X1 U15341 ( .A1(n15424), .A2(n15425), .A3(n15426), .ZN(Result_44_) );
  AND3_X1 U15342 ( .A1(n15427), .A2(n15428), .A3(n14744), .ZN(n15426) );
  INV_X1 U15343 ( .A(n15429), .ZN(n15428) );
  AND2_X1 U15344 ( .A1(n15430), .A2(n15431), .ZN(n15429) );
  OR2_X1 U15345 ( .A1(n15431), .A2(n15430), .ZN(n15427) );
  AND2_X1 U15346 ( .A1(n15432), .A2(n15433), .ZN(n15430) );
  OR2_X1 U15347 ( .A1(n15434), .A2(n15435), .ZN(n15433) );
  INV_X1 U15348 ( .A(n15436), .ZN(n15435) );
  OR2_X1 U15349 ( .A1(n15436), .A2(n15437), .ZN(n15432) );
  INV_X1 U15350 ( .A(n15434), .ZN(n15437) );
  AND2_X1 U15351 ( .A1(n15438), .A2(n15439), .ZN(n15425) );
  OR3_X1 U15352 ( .A1(n15440), .A2(n15441), .A3(n15442), .ZN(n15439) );
  AND2_X1 U15353 ( .A1(n14791), .A2(n15443), .ZN(n15442) );
  AND2_X1 U15354 ( .A1(n14792), .A2(n15444), .ZN(n15441) );
  AND2_X1 U15355 ( .A1(n15445), .A2(n14793), .ZN(n15440) );
  INV_X1 U15356 ( .A(n15446), .ZN(n15445) );
  INV_X1 U15357 ( .A(n15447), .ZN(n15438) );
  AND2_X1 U15358 ( .A1(n15447), .A2(n15448), .ZN(n15424) );
  OR3_X1 U15359 ( .A1(n15449), .A2(n15450), .A3(n15451), .ZN(n15448) );
  AND2_X1 U15360 ( .A1(n14791), .A2(n15452), .ZN(n15451) );
  INV_X1 U15361 ( .A(n15443), .ZN(n15452) );
  AND2_X1 U15362 ( .A1(n14792), .A2(n15453), .ZN(n15450) );
  INV_X1 U15363 ( .A(n15444), .ZN(n15453) );
  AND2_X1 U15364 ( .A1(n14793), .A2(n15446), .ZN(n15449) );
  OR2_X1 U15365 ( .A1(n15454), .A2(n15455), .ZN(n15447) );
  AND2_X1 U15366 ( .A1(a_12_), .A2(n15456), .ZN(n15455) );
  AND2_X1 U15367 ( .A1(b_12_), .A2(n15457), .ZN(n15454) );
  OR3_X1 U15368 ( .A1(n15458), .A2(n15459), .A3(n15460), .ZN(Result_43_) );
  AND3_X1 U15369 ( .A1(n15461), .A2(n15462), .A3(n14744), .ZN(n15460) );
  INV_X1 U15370 ( .A(n15463), .ZN(n15462) );
  AND2_X1 U15371 ( .A1(n15464), .A2(n15465), .ZN(n15463) );
  OR2_X1 U15372 ( .A1(n15465), .A2(n15464), .ZN(n15461) );
  AND2_X1 U15373 ( .A1(n15466), .A2(n15467), .ZN(n15464) );
  OR2_X1 U15374 ( .A1(n15468), .A2(n15469), .ZN(n15467) );
  INV_X1 U15375 ( .A(n15470), .ZN(n15469) );
  OR2_X1 U15376 ( .A1(n15470), .A2(n15471), .ZN(n15466) );
  INV_X1 U15377 ( .A(n15468), .ZN(n15471) );
  AND2_X1 U15378 ( .A1(n15472), .A2(n15473), .ZN(n15459) );
  OR3_X1 U15379 ( .A1(n15474), .A2(n15475), .A3(n15476), .ZN(n15473) );
  AND2_X1 U15380 ( .A1(n14791), .A2(n15477), .ZN(n15476) );
  AND2_X1 U15381 ( .A1(n14792), .A2(n15478), .ZN(n15475) );
  AND2_X1 U15382 ( .A1(n15479), .A2(n14793), .ZN(n15474) );
  INV_X1 U15383 ( .A(n15480), .ZN(n15479) );
  INV_X1 U15384 ( .A(n15481), .ZN(n15472) );
  AND2_X1 U15385 ( .A1(n15481), .A2(n15482), .ZN(n15458) );
  OR3_X1 U15386 ( .A1(n15483), .A2(n15484), .A3(n15485), .ZN(n15482) );
  AND2_X1 U15387 ( .A1(n14791), .A2(n15486), .ZN(n15485) );
  INV_X1 U15388 ( .A(n15477), .ZN(n15486) );
  AND2_X1 U15389 ( .A1(n14792), .A2(n15487), .ZN(n15484) );
  INV_X1 U15390 ( .A(n15478), .ZN(n15487) );
  AND2_X1 U15391 ( .A1(n14793), .A2(n15480), .ZN(n15483) );
  OR2_X1 U15392 ( .A1(n15488), .A2(n15489), .ZN(n15481) );
  AND2_X1 U15393 ( .A1(a_11_), .A2(n15490), .ZN(n15489) );
  AND2_X1 U15394 ( .A1(b_11_), .A2(n15491), .ZN(n15488) );
  OR3_X1 U15395 ( .A1(n15492), .A2(n15493), .A3(n15494), .ZN(Result_42_) );
  AND3_X1 U15396 ( .A1(n15495), .A2(n15496), .A3(n14744), .ZN(n15494) );
  INV_X1 U15397 ( .A(n15497), .ZN(n15496) );
  AND2_X1 U15398 ( .A1(n15498), .A2(n15499), .ZN(n15497) );
  OR2_X1 U15399 ( .A1(n15499), .A2(n15498), .ZN(n15495) );
  AND2_X1 U15400 ( .A1(n15500), .A2(n15501), .ZN(n15498) );
  OR2_X1 U15401 ( .A1(n15502), .A2(n15503), .ZN(n15501) );
  INV_X1 U15402 ( .A(n15504), .ZN(n15503) );
  OR2_X1 U15403 ( .A1(n15504), .A2(n15505), .ZN(n15500) );
  INV_X1 U15404 ( .A(n15502), .ZN(n15505) );
  AND2_X1 U15405 ( .A1(n15506), .A2(n15507), .ZN(n15493) );
  OR3_X1 U15406 ( .A1(n15508), .A2(n15509), .A3(n15510), .ZN(n15507) );
  AND2_X1 U15407 ( .A1(n14791), .A2(n15511), .ZN(n15510) );
  AND2_X1 U15408 ( .A1(n14792), .A2(n15512), .ZN(n15509) );
  AND2_X1 U15409 ( .A1(n15513), .A2(n14793), .ZN(n15508) );
  INV_X1 U15410 ( .A(n15514), .ZN(n15513) );
  INV_X1 U15411 ( .A(n15515), .ZN(n15506) );
  AND2_X1 U15412 ( .A1(n15515), .A2(n15516), .ZN(n15492) );
  OR3_X1 U15413 ( .A1(n15517), .A2(n15518), .A3(n15519), .ZN(n15516) );
  AND2_X1 U15414 ( .A1(n14791), .A2(n15520), .ZN(n15519) );
  INV_X1 U15415 ( .A(n15511), .ZN(n15520) );
  AND2_X1 U15416 ( .A1(n14792), .A2(n15521), .ZN(n15518) );
  INV_X1 U15417 ( .A(n15512), .ZN(n15521) );
  AND2_X1 U15418 ( .A1(n14793), .A2(n15514), .ZN(n15517) );
  OR2_X1 U15419 ( .A1(n15522), .A2(n15523), .ZN(n15515) );
  AND2_X1 U15420 ( .A1(a_10_), .A2(n15524), .ZN(n15523) );
  AND2_X1 U15421 ( .A1(b_10_), .A2(n15525), .ZN(n15522) );
  OR3_X1 U15422 ( .A1(n15526), .A2(n15527), .A3(n15528), .ZN(Result_41_) );
  AND3_X1 U15423 ( .A1(n15529), .A2(n15530), .A3(n14744), .ZN(n15528) );
  INV_X1 U15424 ( .A(n15531), .ZN(n15530) );
  AND2_X1 U15425 ( .A1(n15532), .A2(n15533), .ZN(n15531) );
  OR2_X1 U15426 ( .A1(n15533), .A2(n15532), .ZN(n15529) );
  AND2_X1 U15427 ( .A1(n15534), .A2(n15535), .ZN(n15532) );
  OR2_X1 U15428 ( .A1(n15536), .A2(n15537), .ZN(n15535) );
  INV_X1 U15429 ( .A(n15538), .ZN(n15537) );
  OR2_X1 U15430 ( .A1(n15538), .A2(n15539), .ZN(n15534) );
  INV_X1 U15431 ( .A(n15536), .ZN(n15539) );
  AND2_X1 U15432 ( .A1(n15540), .A2(n15541), .ZN(n15527) );
  OR3_X1 U15433 ( .A1(n15542), .A2(n15543), .A3(n15544), .ZN(n15541) );
  AND2_X1 U15434 ( .A1(n14791), .A2(n15545), .ZN(n15544) );
  AND2_X1 U15435 ( .A1(n14792), .A2(n15546), .ZN(n15543) );
  AND2_X1 U15436 ( .A1(n15547), .A2(n14793), .ZN(n15542) );
  INV_X1 U15437 ( .A(n15548), .ZN(n15547) );
  INV_X1 U15438 ( .A(n15549), .ZN(n15540) );
  AND2_X1 U15439 ( .A1(n15549), .A2(n15550), .ZN(n15526) );
  OR3_X1 U15440 ( .A1(n15551), .A2(n15552), .A3(n15553), .ZN(n15550) );
  AND2_X1 U15441 ( .A1(n14791), .A2(n15554), .ZN(n15553) );
  INV_X1 U15442 ( .A(n15545), .ZN(n15554) );
  AND2_X1 U15443 ( .A1(n14792), .A2(n15555), .ZN(n15552) );
  INV_X1 U15444 ( .A(n15546), .ZN(n15555) );
  AND2_X1 U15445 ( .A1(n14793), .A2(n15548), .ZN(n15551) );
  OR2_X1 U15446 ( .A1(n15556), .A2(n15557), .ZN(n15549) );
  AND2_X1 U15447 ( .A1(a_9_), .A2(n15558), .ZN(n15557) );
  AND2_X1 U15448 ( .A1(b_9_), .A2(n15559), .ZN(n15556) );
  OR3_X1 U15449 ( .A1(n15560), .A2(n15561), .A3(n15562), .ZN(Result_40_) );
  AND3_X1 U15450 ( .A1(n15563), .A2(n15564), .A3(n14744), .ZN(n15562) );
  INV_X1 U15451 ( .A(n15565), .ZN(n15564) );
  AND2_X1 U15452 ( .A1(n15566), .A2(n15567), .ZN(n15565) );
  OR2_X1 U15453 ( .A1(n15567), .A2(n15566), .ZN(n15563) );
  AND2_X1 U15454 ( .A1(n15568), .A2(n15569), .ZN(n15566) );
  OR2_X1 U15455 ( .A1(n15570), .A2(n15571), .ZN(n15569) );
  INV_X1 U15456 ( .A(n15572), .ZN(n15571) );
  OR2_X1 U15457 ( .A1(n15572), .A2(n15573), .ZN(n15568) );
  INV_X1 U15458 ( .A(n15570), .ZN(n15573) );
  AND2_X1 U15459 ( .A1(n15574), .A2(n15575), .ZN(n15561) );
  OR3_X1 U15460 ( .A1(n15576), .A2(n15577), .A3(n15578), .ZN(n15575) );
  AND2_X1 U15461 ( .A1(n14791), .A2(n15579), .ZN(n15578) );
  AND2_X1 U15462 ( .A1(n14792), .A2(n15580), .ZN(n15577) );
  AND2_X1 U15463 ( .A1(n15581), .A2(n14793), .ZN(n15576) );
  INV_X1 U15464 ( .A(n15582), .ZN(n15581) );
  INV_X1 U15465 ( .A(n15583), .ZN(n15574) );
  AND2_X1 U15466 ( .A1(n15583), .A2(n15584), .ZN(n15560) );
  OR3_X1 U15467 ( .A1(n15585), .A2(n15586), .A3(n15587), .ZN(n15584) );
  AND2_X1 U15468 ( .A1(n14791), .A2(n15588), .ZN(n15587) );
  INV_X1 U15469 ( .A(n15579), .ZN(n15588) );
  AND2_X1 U15470 ( .A1(n14792), .A2(n15589), .ZN(n15586) );
  INV_X1 U15471 ( .A(n15580), .ZN(n15589) );
  AND2_X1 U15472 ( .A1(n14793), .A2(n15582), .ZN(n15585) );
  OR2_X1 U15473 ( .A1(n15590), .A2(n15591), .ZN(n15583) );
  AND2_X1 U15474 ( .A1(a_8_), .A2(n15592), .ZN(n15591) );
  AND2_X1 U15475 ( .A1(b_8_), .A2(n15593), .ZN(n15590) );
  OR2_X1 U15476 ( .A1(n15594), .A2(n14741), .ZN(Result_3_) );
  AND3_X1 U15477 ( .A1(n15595), .A2(n15596), .A3(n14744), .ZN(n15594) );
  OR3_X1 U15478 ( .A1(n15597), .A2(n15598), .A3(n15599), .ZN(n15596) );
  INV_X1 U15479 ( .A(n15600), .ZN(n15599) );
  AND2_X1 U15480 ( .A1(n15601), .A2(n15602), .ZN(n15598) );
  INV_X1 U15481 ( .A(n15603), .ZN(n15601) );
  AND2_X1 U15482 ( .A1(n15604), .A2(n15603), .ZN(n15597) );
  OR2_X1 U15483 ( .A1(n15603), .A2(n15600), .ZN(n15595) );
  OR3_X1 U15484 ( .A1(n15605), .A2(n15606), .A3(n15607), .ZN(Result_39_) );
  AND3_X1 U15485 ( .A1(n15608), .A2(n15609), .A3(n14744), .ZN(n15607) );
  INV_X1 U15486 ( .A(n15610), .ZN(n15609) );
  AND2_X1 U15487 ( .A1(n15611), .A2(n15612), .ZN(n15610) );
  OR2_X1 U15488 ( .A1(n15612), .A2(n15611), .ZN(n15608) );
  AND2_X1 U15489 ( .A1(n15613), .A2(n15614), .ZN(n15611) );
  OR2_X1 U15490 ( .A1(n15615), .A2(n15616), .ZN(n15614) );
  INV_X1 U15491 ( .A(n15617), .ZN(n15616) );
  OR2_X1 U15492 ( .A1(n15617), .A2(n15618), .ZN(n15613) );
  INV_X1 U15493 ( .A(n15615), .ZN(n15618) );
  AND2_X1 U15494 ( .A1(n15619), .A2(n15620), .ZN(n15606) );
  OR3_X1 U15495 ( .A1(n15621), .A2(n15622), .A3(n15623), .ZN(n15620) );
  AND2_X1 U15496 ( .A1(n14791), .A2(n15624), .ZN(n15623) );
  AND2_X1 U15497 ( .A1(n14792), .A2(n15625), .ZN(n15622) );
  AND2_X1 U15498 ( .A1(n15626), .A2(n14793), .ZN(n15621) );
  INV_X1 U15499 ( .A(n15627), .ZN(n15626) );
  INV_X1 U15500 ( .A(n15628), .ZN(n15619) );
  AND2_X1 U15501 ( .A1(n15628), .A2(n15629), .ZN(n15605) );
  OR3_X1 U15502 ( .A1(n15630), .A2(n15631), .A3(n15632), .ZN(n15629) );
  AND2_X1 U15503 ( .A1(n14791), .A2(n15633), .ZN(n15632) );
  INV_X1 U15504 ( .A(n15624), .ZN(n15633) );
  AND2_X1 U15505 ( .A1(n14792), .A2(n15634), .ZN(n15631) );
  INV_X1 U15506 ( .A(n15625), .ZN(n15634) );
  AND2_X1 U15507 ( .A1(n14793), .A2(n15627), .ZN(n15630) );
  OR2_X1 U15508 ( .A1(n15635), .A2(n15636), .ZN(n15628) );
  AND2_X1 U15509 ( .A1(a_7_), .A2(n15637), .ZN(n15636) );
  AND2_X1 U15510 ( .A1(b_7_), .A2(n15638), .ZN(n15635) );
  OR3_X1 U15511 ( .A1(n15639), .A2(n15640), .A3(n15641), .ZN(Result_38_) );
  AND3_X1 U15512 ( .A1(n15642), .A2(n15643), .A3(n14744), .ZN(n15641) );
  INV_X1 U15513 ( .A(n15644), .ZN(n15643) );
  AND2_X1 U15514 ( .A1(n15645), .A2(n15646), .ZN(n15644) );
  OR2_X1 U15515 ( .A1(n15646), .A2(n15645), .ZN(n15642) );
  AND2_X1 U15516 ( .A1(n15647), .A2(n15648), .ZN(n15645) );
  OR2_X1 U15517 ( .A1(n15649), .A2(n15650), .ZN(n15648) );
  INV_X1 U15518 ( .A(n15651), .ZN(n15650) );
  OR2_X1 U15519 ( .A1(n15651), .A2(n15652), .ZN(n15647) );
  INV_X1 U15520 ( .A(n15649), .ZN(n15652) );
  AND2_X1 U15521 ( .A1(n15653), .A2(n15654), .ZN(n15640) );
  OR3_X1 U15522 ( .A1(n15655), .A2(n15656), .A3(n15657), .ZN(n15654) );
  AND2_X1 U15523 ( .A1(n14791), .A2(n15658), .ZN(n15657) );
  AND2_X1 U15524 ( .A1(n14792), .A2(n15659), .ZN(n15656) );
  AND2_X1 U15525 ( .A1(n15660), .A2(n14793), .ZN(n15655) );
  INV_X1 U15526 ( .A(n15661), .ZN(n15660) );
  INV_X1 U15527 ( .A(n15662), .ZN(n15653) );
  AND2_X1 U15528 ( .A1(n15662), .A2(n15663), .ZN(n15639) );
  OR3_X1 U15529 ( .A1(n15664), .A2(n15665), .A3(n15666), .ZN(n15663) );
  AND2_X1 U15530 ( .A1(n14791), .A2(n15667), .ZN(n15666) );
  INV_X1 U15531 ( .A(n15658), .ZN(n15667) );
  AND2_X1 U15532 ( .A1(n14792), .A2(n15668), .ZN(n15665) );
  INV_X1 U15533 ( .A(n15659), .ZN(n15668) );
  AND2_X1 U15534 ( .A1(n14793), .A2(n15661), .ZN(n15664) );
  OR2_X1 U15535 ( .A1(n15669), .A2(n15670), .ZN(n15662) );
  AND2_X1 U15536 ( .A1(a_6_), .A2(n15671), .ZN(n15670) );
  AND2_X1 U15537 ( .A1(b_6_), .A2(n15672), .ZN(n15669) );
  OR3_X1 U15538 ( .A1(n15673), .A2(n15674), .A3(n15675), .ZN(Result_37_) );
  AND3_X1 U15539 ( .A1(n15676), .A2(n15677), .A3(n14744), .ZN(n15675) );
  INV_X1 U15540 ( .A(n15678), .ZN(n15677) );
  AND2_X1 U15541 ( .A1(n15679), .A2(n15680), .ZN(n15678) );
  OR2_X1 U15542 ( .A1(n15680), .A2(n15679), .ZN(n15676) );
  AND2_X1 U15543 ( .A1(n15681), .A2(n15682), .ZN(n15679) );
  OR2_X1 U15544 ( .A1(n15683), .A2(n15684), .ZN(n15682) );
  INV_X1 U15545 ( .A(n15685), .ZN(n15684) );
  OR2_X1 U15546 ( .A1(n15685), .A2(n15686), .ZN(n15681) );
  INV_X1 U15547 ( .A(n15683), .ZN(n15686) );
  AND2_X1 U15548 ( .A1(n15687), .A2(n15688), .ZN(n15674) );
  OR3_X1 U15549 ( .A1(n15689), .A2(n15690), .A3(n15691), .ZN(n15688) );
  AND2_X1 U15550 ( .A1(n14791), .A2(n15692), .ZN(n15691) );
  AND2_X1 U15551 ( .A1(n14792), .A2(n15693), .ZN(n15690) );
  AND2_X1 U15552 ( .A1(n15694), .A2(n14793), .ZN(n15689) );
  INV_X1 U15553 ( .A(n15695), .ZN(n15694) );
  INV_X1 U15554 ( .A(n15696), .ZN(n15687) );
  AND2_X1 U15555 ( .A1(n15696), .A2(n15697), .ZN(n15673) );
  OR3_X1 U15556 ( .A1(n15698), .A2(n15699), .A3(n15700), .ZN(n15697) );
  AND2_X1 U15557 ( .A1(n14791), .A2(n15701), .ZN(n15700) );
  INV_X1 U15558 ( .A(n15692), .ZN(n15701) );
  AND2_X1 U15559 ( .A1(n14792), .A2(n15702), .ZN(n15699) );
  INV_X1 U15560 ( .A(n15693), .ZN(n15702) );
  AND2_X1 U15561 ( .A1(n14793), .A2(n15695), .ZN(n15698) );
  OR2_X1 U15562 ( .A1(n15703), .A2(n15704), .ZN(n15696) );
  AND2_X1 U15563 ( .A1(a_5_), .A2(n15705), .ZN(n15704) );
  AND2_X1 U15564 ( .A1(b_5_), .A2(n15706), .ZN(n15703) );
  OR3_X1 U15565 ( .A1(n15707), .A2(n15708), .A3(n15709), .ZN(Result_36_) );
  AND3_X1 U15566 ( .A1(n15710), .A2(n15711), .A3(n14744), .ZN(n15709) );
  INV_X1 U15567 ( .A(n15712), .ZN(n15711) );
  AND2_X1 U15568 ( .A1(n15713), .A2(n15714), .ZN(n15712) );
  OR2_X1 U15569 ( .A1(n15714), .A2(n15713), .ZN(n15710) );
  AND2_X1 U15570 ( .A1(n15715), .A2(n15716), .ZN(n15713) );
  OR2_X1 U15571 ( .A1(n15717), .A2(n15718), .ZN(n15716) );
  INV_X1 U15572 ( .A(n15719), .ZN(n15718) );
  OR2_X1 U15573 ( .A1(n15719), .A2(n15720), .ZN(n15715) );
  INV_X1 U15574 ( .A(n15717), .ZN(n15720) );
  AND2_X1 U15575 ( .A1(n15721), .A2(n15722), .ZN(n15708) );
  OR3_X1 U15576 ( .A1(n15723), .A2(n15724), .A3(n15725), .ZN(n15722) );
  AND2_X1 U15577 ( .A1(n14791), .A2(n15726), .ZN(n15725) );
  AND2_X1 U15578 ( .A1(n14792), .A2(n15727), .ZN(n15724) );
  AND2_X1 U15579 ( .A1(n15728), .A2(n14793), .ZN(n15723) );
  INV_X1 U15580 ( .A(n15729), .ZN(n15728) );
  INV_X1 U15581 ( .A(n15730), .ZN(n15721) );
  AND2_X1 U15582 ( .A1(n15730), .A2(n15731), .ZN(n15707) );
  OR3_X1 U15583 ( .A1(n15732), .A2(n15733), .A3(n15734), .ZN(n15731) );
  AND2_X1 U15584 ( .A1(n14791), .A2(n15735), .ZN(n15734) );
  INV_X1 U15585 ( .A(n15726), .ZN(n15735) );
  AND2_X1 U15586 ( .A1(n14792), .A2(n15736), .ZN(n15733) );
  INV_X1 U15587 ( .A(n15727), .ZN(n15736) );
  AND2_X1 U15588 ( .A1(n14793), .A2(n15729), .ZN(n15732) );
  OR2_X1 U15589 ( .A1(n15737), .A2(n15738), .ZN(n15730) );
  AND2_X1 U15590 ( .A1(a_4_), .A2(n15739), .ZN(n15738) );
  AND2_X1 U15591 ( .A1(b_4_), .A2(n15740), .ZN(n15737) );
  OR3_X1 U15592 ( .A1(n15741), .A2(n15742), .A3(n15743), .ZN(Result_35_) );
  AND3_X1 U15593 ( .A1(n15744), .A2(n15745), .A3(n14744), .ZN(n15743) );
  INV_X1 U15594 ( .A(n15746), .ZN(n15745) );
  AND2_X1 U15595 ( .A1(n15747), .A2(n15748), .ZN(n15746) );
  OR2_X1 U15596 ( .A1(n15748), .A2(n15747), .ZN(n15744) );
  AND2_X1 U15597 ( .A1(n15749), .A2(n15750), .ZN(n15747) );
  OR2_X1 U15598 ( .A1(n15751), .A2(n15752), .ZN(n15750) );
  INV_X1 U15599 ( .A(n15753), .ZN(n15752) );
  OR2_X1 U15600 ( .A1(n15753), .A2(n15754), .ZN(n15749) );
  INV_X1 U15601 ( .A(n15751), .ZN(n15754) );
  AND2_X1 U15602 ( .A1(n15755), .A2(n15756), .ZN(n15742) );
  OR3_X1 U15603 ( .A1(n15757), .A2(n15758), .A3(n15759), .ZN(n15756) );
  AND2_X1 U15604 ( .A1(n14791), .A2(n15760), .ZN(n15759) );
  AND2_X1 U15605 ( .A1(n14792), .A2(n15761), .ZN(n15758) );
  AND2_X1 U15606 ( .A1(n15762), .A2(n14793), .ZN(n15757) );
  INV_X1 U15607 ( .A(n15763), .ZN(n15762) );
  INV_X1 U15608 ( .A(n15764), .ZN(n15755) );
  AND2_X1 U15609 ( .A1(n15764), .A2(n15765), .ZN(n15741) );
  OR3_X1 U15610 ( .A1(n15766), .A2(n15767), .A3(n15768), .ZN(n15765) );
  AND2_X1 U15611 ( .A1(n14791), .A2(n15769), .ZN(n15768) );
  INV_X1 U15612 ( .A(n15760), .ZN(n15769) );
  AND2_X1 U15613 ( .A1(n14792), .A2(n15770), .ZN(n15767) );
  INV_X1 U15614 ( .A(n15761), .ZN(n15770) );
  AND2_X1 U15615 ( .A1(n14793), .A2(n15763), .ZN(n15766) );
  OR2_X1 U15616 ( .A1(n15771), .A2(n15772), .ZN(n15764) );
  AND2_X1 U15617 ( .A1(a_3_), .A2(n15773), .ZN(n15772) );
  AND2_X1 U15618 ( .A1(b_3_), .A2(n15774), .ZN(n15771) );
  OR3_X1 U15619 ( .A1(n15775), .A2(n15776), .A3(n15777), .ZN(Result_34_) );
  AND3_X1 U15620 ( .A1(n15778), .A2(n15779), .A3(n14744), .ZN(n15777) );
  INV_X1 U15621 ( .A(n15780), .ZN(n15779) );
  AND2_X1 U15622 ( .A1(n15781), .A2(n15782), .ZN(n15780) );
  OR2_X1 U15623 ( .A1(n15782), .A2(n15781), .ZN(n15778) );
  AND2_X1 U15624 ( .A1(n15783), .A2(n15784), .ZN(n15781) );
  OR2_X1 U15625 ( .A1(n15785), .A2(n15786), .ZN(n15784) );
  INV_X1 U15626 ( .A(n15787), .ZN(n15786) );
  OR2_X1 U15627 ( .A1(n15787), .A2(n15788), .ZN(n15783) );
  INV_X1 U15628 ( .A(n15785), .ZN(n15788) );
  AND2_X1 U15629 ( .A1(n15789), .A2(n15790), .ZN(n15776) );
  OR3_X1 U15630 ( .A1(n15791), .A2(n15792), .A3(n15793), .ZN(n15790) );
  AND2_X1 U15631 ( .A1(n14791), .A2(n15794), .ZN(n15793) );
  AND2_X1 U15632 ( .A1(n14792), .A2(n15795), .ZN(n15792) );
  AND2_X1 U15633 ( .A1(n15796), .A2(n14793), .ZN(n15791) );
  INV_X1 U15634 ( .A(n15797), .ZN(n15796) );
  INV_X1 U15635 ( .A(n15798), .ZN(n15789) );
  AND2_X1 U15636 ( .A1(n15798), .A2(n15799), .ZN(n15775) );
  OR3_X1 U15637 ( .A1(n15800), .A2(n15801), .A3(n15802), .ZN(n15799) );
  AND2_X1 U15638 ( .A1(n14791), .A2(n15803), .ZN(n15802) );
  INV_X1 U15639 ( .A(n15794), .ZN(n15803) );
  AND2_X1 U15640 ( .A1(n14792), .A2(n15804), .ZN(n15801) );
  INV_X1 U15641 ( .A(n15795), .ZN(n15804) );
  AND2_X1 U15642 ( .A1(n14793), .A2(n15797), .ZN(n15800) );
  OR2_X1 U15643 ( .A1(n15805), .A2(n15806), .ZN(n15798) );
  AND2_X1 U15644 ( .A1(a_2_), .A2(n15807), .ZN(n15806) );
  AND2_X1 U15645 ( .A1(b_2_), .A2(n15808), .ZN(n15805) );
  OR3_X1 U15646 ( .A1(n15809), .A2(n15810), .A3(n15811), .ZN(Result_33_) );
  AND3_X1 U15647 ( .A1(n15812), .A2(n15813), .A3(n14744), .ZN(n15811) );
  INV_X1 U15648 ( .A(n15814), .ZN(n15813) );
  AND2_X1 U15649 ( .A1(n15815), .A2(n15816), .ZN(n15814) );
  OR2_X1 U15650 ( .A1(n15816), .A2(n15815), .ZN(n15812) );
  AND2_X1 U15651 ( .A1(n15817), .A2(n15818), .ZN(n15815) );
  OR2_X1 U15652 ( .A1(n15819), .A2(n15820), .ZN(n15818) );
  INV_X1 U15653 ( .A(n15821), .ZN(n15820) );
  OR2_X1 U15654 ( .A1(n15821), .A2(n15822), .ZN(n15817) );
  INV_X1 U15655 ( .A(n15819), .ZN(n15822) );
  AND2_X1 U15656 ( .A1(n15823), .A2(n15824), .ZN(n15810) );
  OR3_X1 U15657 ( .A1(n15825), .A2(n15826), .A3(n15827), .ZN(n15824) );
  AND2_X1 U15658 ( .A1(n14791), .A2(n15828), .ZN(n15827) );
  AND2_X1 U15659 ( .A1(n14792), .A2(n15829), .ZN(n15826) );
  AND2_X1 U15660 ( .A1(n15830), .A2(n14793), .ZN(n15825) );
  INV_X1 U15661 ( .A(n15831), .ZN(n15830) );
  INV_X1 U15662 ( .A(n15832), .ZN(n15823) );
  AND2_X1 U15663 ( .A1(n15832), .A2(n15833), .ZN(n15809) );
  OR3_X1 U15664 ( .A1(n15834), .A2(n15835), .A3(n15836), .ZN(n15833) );
  AND2_X1 U15665 ( .A1(n14791), .A2(n15837), .ZN(n15836) );
  INV_X1 U15666 ( .A(n15828), .ZN(n15837) );
  AND2_X1 U15667 ( .A1(n14792), .A2(n15838), .ZN(n15835) );
  INV_X1 U15668 ( .A(n15829), .ZN(n15838) );
  AND2_X1 U15669 ( .A1(n14793), .A2(n15831), .ZN(n15834) );
  OR2_X1 U15670 ( .A1(n15839), .A2(n15840), .ZN(n15832) );
  AND2_X1 U15671 ( .A1(a_1_), .A2(n15841), .ZN(n15840) );
  AND2_X1 U15672 ( .A1(b_1_), .A2(n15842), .ZN(n15839) );
  OR4_X1 U15673 ( .A1(n15843), .A2(n15844), .A3(n15845), .A4(n15846), .ZN(
        Result_32_) );
  AND2_X1 U15674 ( .A1(n15847), .A2(n15848), .ZN(n15846) );
  OR2_X1 U15675 ( .A1(n15849), .A2(n15850), .ZN(n15847) );
  AND2_X1 U15676 ( .A1(n15851), .A2(n14791), .ZN(n15850) );
  AND2_X1 U15677 ( .A1(n14792), .A2(n15852), .ZN(n15849) );
  INV_X1 U15678 ( .A(n15853), .ZN(n15852) );
  AND2_X1 U15679 ( .A1(n15854), .A2(n15855), .ZN(n15845) );
  OR3_X1 U15680 ( .A1(n15856), .A2(n15857), .A3(n15858), .ZN(n15855) );
  AND2_X1 U15681 ( .A1(n14791), .A2(n15859), .ZN(n15858) );
  AND2_X1 U15682 ( .A1(n14792), .A2(n15853), .ZN(n15857) );
  AND2_X1 U15683 ( .A1(n14793), .A2(n15860), .ZN(n15856) );
  INV_X1 U15684 ( .A(n15848), .ZN(n15854) );
  AND3_X1 U15685 ( .A1(n15861), .A2(n15860), .A3(n14793), .ZN(n15844) );
  OR2_X1 U15686 ( .A1(n15864), .A2(n15848), .ZN(n15860) );
  OR2_X1 U15687 ( .A1(n15865), .A2(n15866), .ZN(n15848) );
  INV_X1 U15688 ( .A(n15867), .ZN(n15865) );
  INV_X1 U15689 ( .A(n15861), .ZN(n15864) );
  OR2_X1 U15690 ( .A1(n15868), .A2(n15869), .ZN(n15861) );
  AND2_X1 U15691 ( .A1(n15842), .A2(n15841), .ZN(n15869) );
  AND2_X1 U15692 ( .A1(n15831), .A2(n15870), .ZN(n15868) );
  OR2_X1 U15693 ( .A1(n15871), .A2(n15872), .ZN(n15831) );
  AND2_X1 U15694 ( .A1(n15808), .A2(n15807), .ZN(n15872) );
  AND2_X1 U15695 ( .A1(n15797), .A2(n15873), .ZN(n15871) );
  OR2_X1 U15696 ( .A1(n15874), .A2(n15875), .ZN(n15797) );
  AND2_X1 U15697 ( .A1(n15774), .A2(n15773), .ZN(n15875) );
  AND2_X1 U15698 ( .A1(n15763), .A2(n15876), .ZN(n15874) );
  OR2_X1 U15699 ( .A1(n15877), .A2(n15878), .ZN(n15763) );
  AND2_X1 U15700 ( .A1(n15740), .A2(n15739), .ZN(n15878) );
  AND2_X1 U15701 ( .A1(n15729), .A2(n15879), .ZN(n15877) );
  OR2_X1 U15702 ( .A1(n15880), .A2(n15881), .ZN(n15729) );
  AND2_X1 U15703 ( .A1(n15706), .A2(n15705), .ZN(n15881) );
  AND2_X1 U15704 ( .A1(n15695), .A2(n15882), .ZN(n15880) );
  OR2_X1 U15705 ( .A1(n15883), .A2(n15884), .ZN(n15695) );
  AND2_X1 U15706 ( .A1(n15672), .A2(n15671), .ZN(n15884) );
  AND2_X1 U15707 ( .A1(n15661), .A2(n15885), .ZN(n15883) );
  OR2_X1 U15708 ( .A1(n15886), .A2(n15887), .ZN(n15661) );
  AND2_X1 U15709 ( .A1(n15638), .A2(n15637), .ZN(n15887) );
  AND2_X1 U15710 ( .A1(n15627), .A2(n15888), .ZN(n15886) );
  OR2_X1 U15711 ( .A1(n15889), .A2(n15890), .ZN(n15627) );
  AND2_X1 U15712 ( .A1(n15593), .A2(n15592), .ZN(n15890) );
  AND2_X1 U15713 ( .A1(n15582), .A2(n15891), .ZN(n15889) );
  OR2_X1 U15714 ( .A1(n15892), .A2(n15893), .ZN(n15582) );
  AND2_X1 U15715 ( .A1(n15559), .A2(n15558), .ZN(n15893) );
  AND2_X1 U15716 ( .A1(n15548), .A2(n15894), .ZN(n15892) );
  OR2_X1 U15717 ( .A1(n15895), .A2(n15896), .ZN(n15548) );
  AND2_X1 U15718 ( .A1(n15525), .A2(n15524), .ZN(n15896) );
  AND2_X1 U15719 ( .A1(n15514), .A2(n15897), .ZN(n15895) );
  OR2_X1 U15720 ( .A1(n15898), .A2(n15899), .ZN(n15514) );
  AND2_X1 U15721 ( .A1(n15491), .A2(n15490), .ZN(n15899) );
  AND2_X1 U15722 ( .A1(n15480), .A2(n15900), .ZN(n15898) );
  OR2_X1 U15723 ( .A1(n15901), .A2(n15902), .ZN(n15480) );
  AND2_X1 U15724 ( .A1(n15457), .A2(n15456), .ZN(n15902) );
  AND2_X1 U15725 ( .A1(n15446), .A2(n15903), .ZN(n15901) );
  OR2_X1 U15726 ( .A1(n15904), .A2(n15905), .ZN(n15446) );
  AND2_X1 U15727 ( .A1(n15423), .A2(n15422), .ZN(n15905) );
  AND2_X1 U15728 ( .A1(n15412), .A2(n15906), .ZN(n15904) );
  OR2_X1 U15729 ( .A1(n15907), .A2(n15908), .ZN(n15412) );
  AND2_X1 U15730 ( .A1(n15389), .A2(n15388), .ZN(n15908) );
  AND2_X1 U15731 ( .A1(n15378), .A2(n15909), .ZN(n15907) );
  OR2_X1 U15732 ( .A1(n15910), .A2(n15911), .ZN(n15378) );
  AND2_X1 U15733 ( .A1(n15355), .A2(n15354), .ZN(n15911) );
  AND2_X1 U15734 ( .A1(n15344), .A2(n15912), .ZN(n15910) );
  OR2_X1 U15735 ( .A1(n15913), .A2(n15914), .ZN(n15344) );
  AND2_X1 U15736 ( .A1(n15321), .A2(n15320), .ZN(n15914) );
  AND2_X1 U15737 ( .A1(n15310), .A2(n15915), .ZN(n15913) );
  OR2_X1 U15738 ( .A1(n15916), .A2(n15917), .ZN(n15310) );
  AND2_X1 U15739 ( .A1(n15287), .A2(n15286), .ZN(n15917) );
  AND2_X1 U15740 ( .A1(n15276), .A2(n15918), .ZN(n15916) );
  OR2_X1 U15741 ( .A1(n15919), .A2(n15920), .ZN(n15276) );
  AND2_X1 U15742 ( .A1(n15242), .A2(n15241), .ZN(n15920) );
  AND2_X1 U15743 ( .A1(n15231), .A2(n15921), .ZN(n15919) );
  OR2_X1 U15744 ( .A1(n15922), .A2(n15923), .ZN(n15231) );
  AND2_X1 U15745 ( .A1(n15208), .A2(n15207), .ZN(n15923) );
  AND2_X1 U15746 ( .A1(n15197), .A2(n15924), .ZN(n15922) );
  OR2_X1 U15747 ( .A1(n15925), .A2(n15926), .ZN(n15197) );
  AND2_X1 U15748 ( .A1(n15174), .A2(n15173), .ZN(n15926) );
  AND2_X1 U15749 ( .A1(n15163), .A2(n15927), .ZN(n15925) );
  OR2_X1 U15750 ( .A1(n15928), .A2(n15929), .ZN(n15163) );
  AND2_X1 U15751 ( .A1(n15140), .A2(n15139), .ZN(n15929) );
  AND2_X1 U15752 ( .A1(n15129), .A2(n15930), .ZN(n15928) );
  OR2_X1 U15753 ( .A1(n15931), .A2(n15932), .ZN(n15129) );
  AND2_X1 U15754 ( .A1(n15106), .A2(n15105), .ZN(n15932) );
  AND2_X1 U15755 ( .A1(n15095), .A2(n15933), .ZN(n15931) );
  OR2_X1 U15756 ( .A1(n15934), .A2(n15935), .ZN(n15095) );
  AND2_X1 U15757 ( .A1(n15072), .A2(n15071), .ZN(n15935) );
  AND2_X1 U15758 ( .A1(n15061), .A2(n15936), .ZN(n15934) );
  OR2_X1 U15759 ( .A1(n15937), .A2(n15938), .ZN(n15061) );
  AND2_X1 U15760 ( .A1(n15038), .A2(n15037), .ZN(n15938) );
  AND2_X1 U15761 ( .A1(n15027), .A2(n15939), .ZN(n15937) );
  OR2_X1 U15762 ( .A1(n15940), .A2(n15941), .ZN(n15027) );
  AND2_X1 U15763 ( .A1(n15004), .A2(n15003), .ZN(n15941) );
  AND2_X1 U15764 ( .A1(n14993), .A2(n15942), .ZN(n15940) );
  OR2_X1 U15765 ( .A1(n15943), .A2(n15944), .ZN(n14993) );
  AND2_X1 U15766 ( .A1(n14970), .A2(n14969), .ZN(n15944) );
  AND2_X1 U15767 ( .A1(n14959), .A2(n15945), .ZN(n15943) );
  OR2_X1 U15768 ( .A1(n15946), .A2(n15947), .ZN(n14959) );
  AND2_X1 U15769 ( .A1(n14936), .A2(n14935), .ZN(n15947) );
  AND2_X1 U15770 ( .A1(n14925), .A2(n15948), .ZN(n15946) );
  OR2_X1 U15771 ( .A1(n15949), .A2(n15950), .ZN(n14925) );
  AND2_X1 U15772 ( .A1(n14891), .A2(n14890), .ZN(n15950) );
  AND2_X1 U15773 ( .A1(n14880), .A2(n15951), .ZN(n15949) );
  OR2_X1 U15774 ( .A1(n15952), .A2(n15953), .ZN(n14880) );
  AND2_X1 U15775 ( .A1(n14857), .A2(n14856), .ZN(n15953) );
  AND2_X1 U15776 ( .A1(n14853), .A2(n15954), .ZN(n15952) );
  INV_X1 U15777 ( .A(n14845), .ZN(n14853) );
  OR3_X1 U15778 ( .A1(n14818), .A2(n15955), .A3(n15956), .ZN(n14845) );
  AND2_X1 U15779 ( .A1(n15957), .A2(b_31_), .ZN(n15956) );
  AND2_X1 U15780 ( .A1(n14788), .A2(b_30_), .ZN(n15955) );
  INV_X1 U15781 ( .A(n14815), .ZN(n14788) );
  OR2_X1 U15782 ( .A1(n15958), .A2(n15959), .ZN(n14815) );
  AND3_X1 U15783 ( .A1(n15960), .A2(n15961), .A3(n14744), .ZN(n15843) );
  INV_X1 U15784 ( .A(n15962), .ZN(n15961) );
  AND2_X1 U15785 ( .A1(n15963), .A2(n15964), .ZN(n15962) );
  OR2_X1 U15786 ( .A1(n15964), .A2(n15963), .ZN(n15960) );
  AND2_X1 U15787 ( .A1(n15965), .A2(n15966), .ZN(n15963) );
  OR2_X1 U15788 ( .A1(n15967), .A2(n15968), .ZN(n15966) );
  INV_X1 U15789 ( .A(n15969), .ZN(n15968) );
  OR2_X1 U15790 ( .A1(n15969), .A2(n15970), .ZN(n15965) );
  INV_X1 U15791 ( .A(n15967), .ZN(n15970) );
  OR2_X1 U15792 ( .A1(n15971), .A2(n14741), .ZN(Result_31_) );
  AND3_X1 U15793 ( .A1(n15972), .A2(n15973), .A3(n14744), .ZN(n15971) );
  OR2_X1 U15794 ( .A1(n15974), .A2(n15975), .ZN(n15973) );
  INV_X1 U15795 ( .A(n15976), .ZN(n15975) );
  OR2_X1 U15796 ( .A1(n15977), .A2(n15976), .ZN(n15972) );
  OR2_X1 U15797 ( .A1(n15978), .A2(n14741), .ZN(Result_30_) );
  AND2_X1 U15798 ( .A1(n15979), .A2(n15980), .ZN(n15978) );
  OR2_X1 U15799 ( .A1(n15981), .A2(n15982), .ZN(n15980) );
  AND2_X1 U15800 ( .A1(n15977), .A2(n15976), .ZN(n15981) );
  OR2_X1 U15801 ( .A1(n15983), .A2(n14741), .ZN(Result_2_) );
  AND3_X1 U15802 ( .A1(n15984), .A2(n15985), .A3(n14744), .ZN(n15983) );
  OR3_X1 U15803 ( .A1(n15986), .A2(n15987), .A3(n15988), .ZN(n15985) );
  INV_X1 U15804 ( .A(n15989), .ZN(n15988) );
  AND2_X1 U15805 ( .A1(n15990), .A2(n15991), .ZN(n15987) );
  INV_X1 U15806 ( .A(n15992), .ZN(n15990) );
  AND2_X1 U15807 ( .A1(n15993), .A2(n15992), .ZN(n15986) );
  OR2_X1 U15808 ( .A1(n15992), .A2(n15989), .ZN(n15984) );
  OR3_X1 U15809 ( .A1(n15994), .A2(n15995), .A3(n14741), .ZN(Result_29_) );
  AND2_X1 U15810 ( .A1(n15996), .A2(n15979), .ZN(n15995) );
  AND2_X1 U15811 ( .A1(n15997), .A2(n14744), .ZN(n15979) );
  INV_X1 U15812 ( .A(n15998), .ZN(n15997) );
  INV_X1 U15813 ( .A(n15999), .ZN(n15996) );
  AND3_X1 U15814 ( .A1(n14744), .A2(n15998), .A3(n15999), .ZN(n15994) );
  OR2_X1 U15815 ( .A1(n16000), .A2(n16001), .ZN(n15999) );
  INV_X1 U15816 ( .A(n16002), .ZN(n16000) );
  OR2_X1 U15817 ( .A1(n16003), .A2(n14741), .ZN(Result_28_) );
  AND3_X1 U15818 ( .A1(n16004), .A2(n16005), .A3(n14744), .ZN(n16003) );
  INV_X1 U15819 ( .A(n16006), .ZN(n16005) );
  OR2_X1 U15820 ( .A1(n16007), .A2(n16008), .ZN(n16004) );
  AND2_X1 U15821 ( .A1(n16009), .A2(n16010), .ZN(n16007) );
  INV_X1 U15822 ( .A(n16011), .ZN(n16010) );
  OR2_X1 U15823 ( .A1(n16012), .A2(n14741), .ZN(Result_27_) );
  AND3_X1 U15824 ( .A1(n16013), .A2(n16014), .A3(n14744), .ZN(n16012) );
  INV_X1 U15825 ( .A(n16015), .ZN(n16014) );
  OR2_X1 U15826 ( .A1(n16016), .A2(n16017), .ZN(n16013) );
  AND2_X1 U15827 ( .A1(n16018), .A2(n16019), .ZN(n16016) );
  INV_X1 U15828 ( .A(n16020), .ZN(n16018) );
  OR2_X1 U15829 ( .A1(n16021), .A2(n14741), .ZN(Result_26_) );
  AND3_X1 U15830 ( .A1(n16022), .A2(n16023), .A3(n14744), .ZN(n16021) );
  OR2_X1 U15831 ( .A1(n16024), .A2(n16025), .ZN(n16023) );
  INV_X1 U15832 ( .A(n16026), .ZN(n16022) );
  AND2_X1 U15833 ( .A1(n16025), .A2(n16024), .ZN(n16026) );
  AND2_X1 U15834 ( .A1(n16027), .A2(n16028), .ZN(n16024) );
  INV_X1 U15835 ( .A(n16029), .ZN(n16027) );
  OR2_X1 U15836 ( .A1(n16030), .A2(n14741), .ZN(Result_25_) );
  AND3_X1 U15837 ( .A1(n16031), .A2(n16032), .A3(n14744), .ZN(n16030) );
  OR2_X1 U15838 ( .A1(n16033), .A2(n16034), .ZN(n16032) );
  AND2_X1 U15839 ( .A1(n16035), .A2(n16036), .ZN(n16033) );
  INV_X1 U15840 ( .A(n16037), .ZN(n16036) );
  INV_X1 U15841 ( .A(n16038), .ZN(n16031) );
  OR2_X1 U15842 ( .A1(n16039), .A2(n14741), .ZN(Result_24_) );
  AND3_X1 U15843 ( .A1(n16040), .A2(n16041), .A3(n14744), .ZN(n16039) );
  OR2_X1 U15844 ( .A1(n16042), .A2(n16043), .ZN(n16041) );
  INV_X1 U15845 ( .A(n16044), .ZN(n16040) );
  AND2_X1 U15846 ( .A1(n16043), .A2(n16042), .ZN(n16044) );
  AND2_X1 U15847 ( .A1(n16045), .A2(n16046), .ZN(n16042) );
  INV_X1 U15848 ( .A(n16047), .ZN(n16046) );
  OR2_X1 U15849 ( .A1(n16048), .A2(n14741), .ZN(Result_23_) );
  AND3_X1 U15850 ( .A1(n16049), .A2(n16050), .A3(n14744), .ZN(n16048) );
  OR2_X1 U15851 ( .A1(n16051), .A2(n16052), .ZN(n16050) );
  INV_X1 U15852 ( .A(n16053), .ZN(n16049) );
  AND2_X1 U15853 ( .A1(n16052), .A2(n16051), .ZN(n16053) );
  AND2_X1 U15854 ( .A1(n16054), .A2(n16055), .ZN(n16051) );
  INV_X1 U15855 ( .A(n16056), .ZN(n16055) );
  OR2_X1 U15856 ( .A1(n16057), .A2(n14741), .ZN(Result_22_) );
  AND3_X1 U15857 ( .A1(n16058), .A2(n16059), .A3(n14744), .ZN(n16057) );
  OR2_X1 U15858 ( .A1(n16060), .A2(n16061), .ZN(n16059) );
  AND2_X1 U15859 ( .A1(n16062), .A2(n16063), .ZN(n16060) );
  INV_X1 U15860 ( .A(n16064), .ZN(n16063) );
  INV_X1 U15861 ( .A(n16065), .ZN(n16058) );
  OR2_X1 U15862 ( .A1(n16066), .A2(n14741), .ZN(Result_21_) );
  AND3_X1 U15863 ( .A1(n16067), .A2(n16068), .A3(n14744), .ZN(n16066) );
  OR2_X1 U15864 ( .A1(n16069), .A2(n16070), .ZN(n16068) );
  AND2_X1 U15865 ( .A1(n16071), .A2(n16072), .ZN(n16069) );
  INV_X1 U15866 ( .A(n16073), .ZN(n16072) );
  INV_X1 U15867 ( .A(n16074), .ZN(n16067) );
  OR2_X1 U15868 ( .A1(n16075), .A2(n14741), .ZN(Result_20_) );
  AND3_X1 U15869 ( .A1(n16076), .A2(n16077), .A3(n14744), .ZN(n16075) );
  OR2_X1 U15870 ( .A1(n16078), .A2(n16079), .ZN(n16077) );
  INV_X1 U15871 ( .A(n16080), .ZN(n16076) );
  AND2_X1 U15872 ( .A1(n16079), .A2(n16078), .ZN(n16080) );
  AND2_X1 U15873 ( .A1(n16081), .A2(n16082), .ZN(n16078) );
  INV_X1 U15874 ( .A(n16083), .ZN(n16082) );
  OR2_X1 U15875 ( .A1(n16084), .A2(n14741), .ZN(Result_1_) );
  AND3_X1 U15876 ( .A1(n16085), .A2(n16086), .A3(n14744), .ZN(n16084) );
  OR3_X1 U15877 ( .A1(n16087), .A2(n16088), .A3(n16089), .ZN(n16086) );
  AND2_X1 U15878 ( .A1(n16090), .A2(n16091), .ZN(n16088) );
  AND2_X1 U15879 ( .A1(n16092), .A2(n16093), .ZN(n16087) );
  OR2_X1 U15880 ( .A1(n16094), .A2(n16092), .ZN(n16085) );
  OR2_X1 U15881 ( .A1(n16095), .A2(n14741), .ZN(Result_19_) );
  AND3_X1 U15882 ( .A1(n16096), .A2(n16097), .A3(n14744), .ZN(n16095) );
  OR2_X1 U15883 ( .A1(n16098), .A2(n16099), .ZN(n16097) );
  INV_X1 U15884 ( .A(n16100), .ZN(n16096) );
  AND2_X1 U15885 ( .A1(n16099), .A2(n16098), .ZN(n16100) );
  AND2_X1 U15886 ( .A1(n16101), .A2(n16102), .ZN(n16098) );
  INV_X1 U15887 ( .A(n16103), .ZN(n16102) );
  OR2_X1 U15888 ( .A1(n16104), .A2(n14741), .ZN(Result_18_) );
  AND3_X1 U15889 ( .A1(n16105), .A2(n16106), .A3(n14744), .ZN(n16104) );
  OR2_X1 U15890 ( .A1(n16107), .A2(n16108), .ZN(n16106) );
  AND2_X1 U15891 ( .A1(n16109), .A2(n16110), .ZN(n16107) );
  OR2_X1 U15892 ( .A1(n16111), .A2(n14741), .ZN(Result_17_) );
  AND3_X1 U15893 ( .A1(n16112), .A2(n16113), .A3(n14744), .ZN(n16111) );
  INV_X1 U15894 ( .A(n16114), .ZN(n16113) );
  AND2_X1 U15895 ( .A1(n16115), .A2(n16116), .ZN(n16114) );
  OR2_X1 U15896 ( .A1(n16116), .A2(n16115), .ZN(n16112) );
  OR2_X1 U15897 ( .A1(n16117), .A2(n16118), .ZN(n16115) );
  OR2_X1 U15898 ( .A1(n16119), .A2(n14741), .ZN(Result_16_) );
  AND3_X1 U15899 ( .A1(n16120), .A2(n16121), .A3(n14744), .ZN(n16119) );
  OR2_X1 U15900 ( .A1(n16122), .A2(n16123), .ZN(n16121) );
  INV_X1 U15901 ( .A(n16124), .ZN(n16120) );
  AND2_X1 U15902 ( .A1(n16123), .A2(n16122), .ZN(n16124) );
  AND2_X1 U15903 ( .A1(n16125), .A2(n16126), .ZN(n16122) );
  INV_X1 U15904 ( .A(n16127), .ZN(n16126) );
  OR2_X1 U15905 ( .A1(n16128), .A2(n16129), .ZN(n16125) );
  OR2_X1 U15906 ( .A1(n16130), .A2(n14741), .ZN(Result_15_) );
  AND3_X1 U15907 ( .A1(n16131), .A2(n16132), .A3(n14744), .ZN(n16130) );
  OR2_X1 U15908 ( .A1(n16133), .A2(n16134), .ZN(n16132) );
  INV_X1 U15909 ( .A(n16135), .ZN(n16131) );
  AND2_X1 U15910 ( .A1(n16134), .A2(n16133), .ZN(n16135) );
  AND2_X1 U15911 ( .A1(n16136), .A2(n16137), .ZN(n16133) );
  INV_X1 U15912 ( .A(n16138), .ZN(n16136) );
  AND2_X1 U15913 ( .A1(n16139), .A2(n16140), .ZN(n16138) );
  OR2_X1 U15914 ( .A1(n16141), .A2(n14741), .ZN(Result_14_) );
  AND3_X1 U15915 ( .A1(n16142), .A2(n16143), .A3(n14744), .ZN(n16141) );
  INV_X1 U15916 ( .A(n16144), .ZN(n16143) );
  AND2_X1 U15917 ( .A1(n16145), .A2(n16146), .ZN(n16144) );
  OR2_X1 U15918 ( .A1(n16146), .A2(n16145), .ZN(n16142) );
  OR2_X1 U15919 ( .A1(n16147), .A2(n16148), .ZN(n16145) );
  AND2_X1 U15920 ( .A1(n16149), .A2(n16150), .ZN(n16148) );
  INV_X1 U15921 ( .A(n16151), .ZN(n16147) );
  OR2_X1 U15922 ( .A1(n16152), .A2(n14741), .ZN(Result_13_) );
  AND3_X1 U15923 ( .A1(n16153), .A2(n16154), .A3(n14744), .ZN(n16152) );
  OR2_X1 U15924 ( .A1(n16155), .A2(n16156), .ZN(n16154) );
  OR3_X1 U15925 ( .A1(n16157), .A2(n16158), .A3(n16159), .ZN(n16153) );
  INV_X1 U15926 ( .A(n16155), .ZN(n16159) );
  AND2_X1 U15927 ( .A1(n16160), .A2(n16156), .ZN(n16158) );
  AND2_X1 U15928 ( .A1(n16161), .A2(n16162), .ZN(n16157) );
  INV_X1 U15929 ( .A(n16156), .ZN(n16161) );
  OR2_X1 U15930 ( .A1(n16163), .A2(n14741), .ZN(Result_12_) );
  AND2_X1 U15931 ( .A1(n14744), .A2(n16164), .ZN(n16163) );
  OR2_X1 U15932 ( .A1(n16165), .A2(n16166), .ZN(n16164) );
  AND2_X1 U15933 ( .A1(n16167), .A2(n16168), .ZN(n16166) );
  INV_X1 U15934 ( .A(n16169), .ZN(n16165) );
  OR2_X1 U15935 ( .A1(n16168), .A2(n16167), .ZN(n16169) );
  AND2_X1 U15936 ( .A1(n16170), .A2(n16171), .ZN(n16167) );
  OR2_X1 U15937 ( .A1(n16172), .A2(n16173), .ZN(n16171) );
  INV_X1 U15938 ( .A(n16174), .ZN(n16172) );
  OR2_X1 U15939 ( .A1(n16175), .A2(n14741), .ZN(Result_11_) );
  AND3_X1 U15940 ( .A1(n16176), .A2(n16177), .A3(n14744), .ZN(n16175) );
  OR2_X1 U15941 ( .A1(n16178), .A2(n16179), .ZN(n16177) );
  OR3_X1 U15942 ( .A1(n16180), .A2(n16181), .A3(n16182), .ZN(n16176) );
  INV_X1 U15943 ( .A(n16178), .ZN(n16182) );
  AND2_X1 U15944 ( .A1(n16183), .A2(n16179), .ZN(n16181) );
  INV_X1 U15945 ( .A(n16184), .ZN(n16183) );
  AND2_X1 U15946 ( .A1(n16185), .A2(n16184), .ZN(n16180) );
  INV_X1 U15947 ( .A(n16179), .ZN(n16185) );
  OR2_X1 U15948 ( .A1(n16186), .A2(n14741), .ZN(Result_10_) );
  AND3_X1 U15949 ( .A1(n16187), .A2(n16188), .A3(n14744), .ZN(n16186) );
  OR3_X1 U15950 ( .A1(n16189), .A2(n16190), .A3(n16191), .ZN(n16188) );
  INV_X1 U15951 ( .A(n16192), .ZN(n16191) );
  AND2_X1 U15952 ( .A1(n16193), .A2(n16194), .ZN(n16190) );
  AND2_X1 U15953 ( .A1(n16195), .A2(n16196), .ZN(n16189) );
  INV_X1 U15954 ( .A(n16194), .ZN(n16195) );
  OR2_X1 U15955 ( .A1(n16194), .A2(n16192), .ZN(n16187) );
  OR2_X1 U15956 ( .A1(n16197), .A2(n14741), .ZN(Result_0_) );
  OR2_X1 U15957 ( .A1(n16198), .A2(n16199), .ZN(n14741) );
  AND2_X1 U15958 ( .A1(n14791), .A2(n16200), .ZN(n16199) );
  INV_X1 U15959 ( .A(n16201), .ZN(n16200) );
  AND2_X1 U15960 ( .A1(n16202), .A2(n15867), .ZN(n16201) );
  OR2_X1 U15961 ( .A1(n15851), .A2(n15866), .ZN(n16202) );
  INV_X1 U15962 ( .A(n15859), .ZN(n15851) );
  OR2_X1 U15963 ( .A1(n16203), .A2(n16204), .ZN(n15859) );
  AND2_X1 U15964 ( .A1(n15828), .A2(n15842), .ZN(n16204) );
  AND2_X1 U15965 ( .A1(b_1_), .A2(n16205), .ZN(n16203) );
  OR2_X1 U15966 ( .A1(n15842), .A2(n15828), .ZN(n16205) );
  OR2_X1 U15967 ( .A1(n16206), .A2(n16207), .ZN(n15828) );
  AND2_X1 U15968 ( .A1(n15794), .A2(n15808), .ZN(n16207) );
  AND2_X1 U15969 ( .A1(b_2_), .A2(n16208), .ZN(n16206) );
  OR2_X1 U15970 ( .A1(n15808), .A2(n15794), .ZN(n16208) );
  OR2_X1 U15971 ( .A1(n16209), .A2(n16210), .ZN(n15794) );
  AND2_X1 U15972 ( .A1(n15760), .A2(n15774), .ZN(n16210) );
  AND2_X1 U15973 ( .A1(b_3_), .A2(n16211), .ZN(n16209) );
  OR2_X1 U15974 ( .A1(n15774), .A2(n15760), .ZN(n16211) );
  OR2_X1 U15975 ( .A1(n16212), .A2(n16213), .ZN(n15760) );
  AND2_X1 U15976 ( .A1(n15726), .A2(n15740), .ZN(n16213) );
  AND2_X1 U15977 ( .A1(b_4_), .A2(n16214), .ZN(n16212) );
  OR2_X1 U15978 ( .A1(n15740), .A2(n15726), .ZN(n16214) );
  OR2_X1 U15979 ( .A1(n16215), .A2(n16216), .ZN(n15726) );
  AND2_X1 U15980 ( .A1(n15692), .A2(n15706), .ZN(n16216) );
  AND2_X1 U15981 ( .A1(b_5_), .A2(n16217), .ZN(n16215) );
  OR2_X1 U15982 ( .A1(n15706), .A2(n15692), .ZN(n16217) );
  OR2_X1 U15983 ( .A1(n16218), .A2(n16219), .ZN(n15692) );
  AND2_X1 U15984 ( .A1(n15658), .A2(n15672), .ZN(n16219) );
  AND2_X1 U15985 ( .A1(b_6_), .A2(n16220), .ZN(n16218) );
  OR2_X1 U15986 ( .A1(n15672), .A2(n15658), .ZN(n16220) );
  OR2_X1 U15987 ( .A1(n16221), .A2(n16222), .ZN(n15658) );
  AND2_X1 U15988 ( .A1(n15624), .A2(n15638), .ZN(n16222) );
  AND2_X1 U15989 ( .A1(b_7_), .A2(n16223), .ZN(n16221) );
  OR2_X1 U15990 ( .A1(n15638), .A2(n15624), .ZN(n16223) );
  OR2_X1 U15991 ( .A1(n16224), .A2(n16225), .ZN(n15624) );
  AND2_X1 U15992 ( .A1(n15579), .A2(n15593), .ZN(n16225) );
  AND2_X1 U15993 ( .A1(b_8_), .A2(n16226), .ZN(n16224) );
  OR2_X1 U15994 ( .A1(n15593), .A2(n15579), .ZN(n16226) );
  OR2_X1 U15995 ( .A1(n16227), .A2(n16228), .ZN(n15579) );
  AND2_X1 U15996 ( .A1(n15545), .A2(n15559), .ZN(n16228) );
  AND2_X1 U15997 ( .A1(b_9_), .A2(n16229), .ZN(n16227) );
  OR2_X1 U15998 ( .A1(n15559), .A2(n15545), .ZN(n16229) );
  OR2_X1 U15999 ( .A1(n16230), .A2(n16231), .ZN(n15545) );
  AND2_X1 U16000 ( .A1(n15511), .A2(n15525), .ZN(n16231) );
  AND2_X1 U16001 ( .A1(b_10_), .A2(n16232), .ZN(n16230) );
  OR2_X1 U16002 ( .A1(n15525), .A2(n15511), .ZN(n16232) );
  OR2_X1 U16003 ( .A1(n16233), .A2(n16234), .ZN(n15511) );
  AND2_X1 U16004 ( .A1(n15477), .A2(n15491), .ZN(n16234) );
  AND2_X1 U16005 ( .A1(b_11_), .A2(n16235), .ZN(n16233) );
  OR2_X1 U16006 ( .A1(n15491), .A2(n15477), .ZN(n16235) );
  OR2_X1 U16007 ( .A1(n16236), .A2(n16237), .ZN(n15477) );
  AND2_X1 U16008 ( .A1(n15443), .A2(n15457), .ZN(n16237) );
  AND2_X1 U16009 ( .A1(b_12_), .A2(n16238), .ZN(n16236) );
  OR2_X1 U16010 ( .A1(n15457), .A2(n15443), .ZN(n16238) );
  OR2_X1 U16011 ( .A1(n16239), .A2(n16240), .ZN(n15443) );
  AND2_X1 U16012 ( .A1(n15409), .A2(n15423), .ZN(n16240) );
  AND2_X1 U16013 ( .A1(b_13_), .A2(n16241), .ZN(n16239) );
  OR2_X1 U16014 ( .A1(n15423), .A2(n15409), .ZN(n16241) );
  OR2_X1 U16015 ( .A1(n16242), .A2(n16243), .ZN(n15409) );
  AND2_X1 U16016 ( .A1(n15375), .A2(n15389), .ZN(n16243) );
  AND2_X1 U16017 ( .A1(b_14_), .A2(n16244), .ZN(n16242) );
  OR2_X1 U16018 ( .A1(n15389), .A2(n15375), .ZN(n16244) );
  OR2_X1 U16019 ( .A1(n16245), .A2(n16246), .ZN(n15375) );
  AND2_X1 U16020 ( .A1(n15341), .A2(n15355), .ZN(n16246) );
  AND2_X1 U16021 ( .A1(b_15_), .A2(n16247), .ZN(n16245) );
  OR2_X1 U16022 ( .A1(n15355), .A2(n15341), .ZN(n16247) );
  OR2_X1 U16023 ( .A1(n16248), .A2(n16249), .ZN(n15341) );
  AND2_X1 U16024 ( .A1(n15307), .A2(n15321), .ZN(n16249) );
  AND2_X1 U16025 ( .A1(b_16_), .A2(n16250), .ZN(n16248) );
  OR2_X1 U16026 ( .A1(n15321), .A2(n15307), .ZN(n16250) );
  OR2_X1 U16027 ( .A1(n16251), .A2(n16252), .ZN(n15307) );
  AND2_X1 U16028 ( .A1(n15273), .A2(n15287), .ZN(n16252) );
  AND2_X1 U16029 ( .A1(b_17_), .A2(n16253), .ZN(n16251) );
  OR2_X1 U16030 ( .A1(n15287), .A2(n15273), .ZN(n16253) );
  OR2_X1 U16031 ( .A1(n16254), .A2(n16255), .ZN(n15273) );
  AND2_X1 U16032 ( .A1(n15228), .A2(n15242), .ZN(n16255) );
  AND2_X1 U16033 ( .A1(b_18_), .A2(n16256), .ZN(n16254) );
  OR2_X1 U16034 ( .A1(n15242), .A2(n15228), .ZN(n16256) );
  OR2_X1 U16035 ( .A1(n16257), .A2(n16258), .ZN(n15228) );
  AND2_X1 U16036 ( .A1(n15194), .A2(n15208), .ZN(n16258) );
  AND2_X1 U16037 ( .A1(b_19_), .A2(n16259), .ZN(n16257) );
  OR2_X1 U16038 ( .A1(n15208), .A2(n15194), .ZN(n16259) );
  OR2_X1 U16039 ( .A1(n16260), .A2(n16261), .ZN(n15194) );
  AND2_X1 U16040 ( .A1(n15160), .A2(n15174), .ZN(n16261) );
  AND2_X1 U16041 ( .A1(b_20_), .A2(n16262), .ZN(n16260) );
  OR2_X1 U16042 ( .A1(n15174), .A2(n15160), .ZN(n16262) );
  OR2_X1 U16043 ( .A1(n16263), .A2(n16264), .ZN(n15160) );
  AND2_X1 U16044 ( .A1(n15126), .A2(n15140), .ZN(n16264) );
  AND2_X1 U16045 ( .A1(b_21_), .A2(n16265), .ZN(n16263) );
  OR2_X1 U16046 ( .A1(n15140), .A2(n15126), .ZN(n16265) );
  OR2_X1 U16047 ( .A1(n16266), .A2(n16267), .ZN(n15126) );
  AND2_X1 U16048 ( .A1(n15092), .A2(n15106), .ZN(n16267) );
  AND2_X1 U16049 ( .A1(b_22_), .A2(n16268), .ZN(n16266) );
  OR2_X1 U16050 ( .A1(n15106), .A2(n15092), .ZN(n16268) );
  OR2_X1 U16051 ( .A1(n16269), .A2(n16270), .ZN(n15092) );
  AND2_X1 U16052 ( .A1(n15058), .A2(n15072), .ZN(n16270) );
  AND2_X1 U16053 ( .A1(b_23_), .A2(n16271), .ZN(n16269) );
  OR2_X1 U16054 ( .A1(n15072), .A2(n15058), .ZN(n16271) );
  OR2_X1 U16055 ( .A1(n16272), .A2(n16273), .ZN(n15058) );
  AND2_X1 U16056 ( .A1(n15024), .A2(n15038), .ZN(n16273) );
  AND2_X1 U16057 ( .A1(b_24_), .A2(n16274), .ZN(n16272) );
  OR2_X1 U16058 ( .A1(n15038), .A2(n15024), .ZN(n16274) );
  OR2_X1 U16059 ( .A1(n16275), .A2(n16276), .ZN(n15024) );
  AND2_X1 U16060 ( .A1(n14990), .A2(n15004), .ZN(n16276) );
  AND2_X1 U16061 ( .A1(b_25_), .A2(n16277), .ZN(n16275) );
  OR2_X1 U16062 ( .A1(n15004), .A2(n14990), .ZN(n16277) );
  OR2_X1 U16063 ( .A1(n16278), .A2(n16279), .ZN(n14990) );
  AND2_X1 U16064 ( .A1(n14956), .A2(n14970), .ZN(n16279) );
  AND2_X1 U16065 ( .A1(b_26_), .A2(n16280), .ZN(n16278) );
  OR2_X1 U16066 ( .A1(n14970), .A2(n14956), .ZN(n16280) );
  OR2_X1 U16067 ( .A1(n16281), .A2(n16282), .ZN(n14956) );
  AND2_X1 U16068 ( .A1(n14922), .A2(n14936), .ZN(n16282) );
  AND2_X1 U16069 ( .A1(b_27_), .A2(n16283), .ZN(n16281) );
  OR2_X1 U16070 ( .A1(n14936), .A2(n14922), .ZN(n16283) );
  OR2_X1 U16071 ( .A1(n16284), .A2(n16285), .ZN(n14922) );
  AND2_X1 U16072 ( .A1(n14877), .A2(n14891), .ZN(n16285) );
  AND2_X1 U16073 ( .A1(b_28_), .A2(n16286), .ZN(n16284) );
  OR2_X1 U16074 ( .A1(n14891), .A2(n14877), .ZN(n16286) );
  OR2_X1 U16075 ( .A1(n16287), .A2(n16288), .ZN(n14877) );
  AND2_X1 U16076 ( .A1(n14843), .A2(n14857), .ZN(n16288) );
  AND2_X1 U16077 ( .A1(b_29_), .A2(n16289), .ZN(n16287) );
  OR2_X1 U16078 ( .A1(n14857), .A2(n14843), .ZN(n16289) );
  OR2_X1 U16079 ( .A1(n16290), .A2(n16291), .ZN(n14843) );
  AND2_X1 U16080 ( .A1(n14795), .A2(n14806), .ZN(n16291) );
  AND2_X1 U16081 ( .A1(b_30_), .A2(n16292), .ZN(n16290) );
  OR2_X1 U16082 ( .A1(n14795), .A2(n14806), .ZN(n16292) );
  INV_X1 U16083 ( .A(n14813), .ZN(n14795) );
  OR2_X1 U16084 ( .A1(a_31_), .A2(n15959), .ZN(n14813) );
  INV_X1 U16085 ( .A(operation_0_), .ZN(n15863) );
  AND3_X1 U16086 ( .A1(n16293), .A2(n15867), .A3(n14792), .ZN(n16198) );
  INV_X1 U16087 ( .A(operation_1_), .ZN(n15862) );
  OR2_X1 U16088 ( .A1(a_0_), .A2(n16294), .ZN(n15867) );
  OR2_X1 U16089 ( .A1(n15866), .A2(n15853), .ZN(n16293) );
  OR2_X1 U16090 ( .A1(n16295), .A2(n16296), .ZN(n15853) );
  AND2_X1 U16091 ( .A1(a_1_), .A2(n15829), .ZN(n16296) );
  AND2_X1 U16092 ( .A1(n16297), .A2(n15841), .ZN(n16295) );
  OR2_X1 U16093 ( .A1(a_1_), .A2(n15829), .ZN(n16297) );
  OR2_X1 U16094 ( .A1(n16298), .A2(n16299), .ZN(n15829) );
  AND2_X1 U16095 ( .A1(a_2_), .A2(n15795), .ZN(n16299) );
  AND2_X1 U16096 ( .A1(n16300), .A2(n15807), .ZN(n16298) );
  OR2_X1 U16097 ( .A1(a_2_), .A2(n15795), .ZN(n16300) );
  OR2_X1 U16098 ( .A1(n16301), .A2(n16302), .ZN(n15795) );
  AND2_X1 U16099 ( .A1(a_3_), .A2(n15761), .ZN(n16302) );
  AND2_X1 U16100 ( .A1(n16303), .A2(n15773), .ZN(n16301) );
  OR2_X1 U16101 ( .A1(a_3_), .A2(n15761), .ZN(n16303) );
  OR2_X1 U16102 ( .A1(n16304), .A2(n16305), .ZN(n15761) );
  AND2_X1 U16103 ( .A1(a_4_), .A2(n15727), .ZN(n16305) );
  AND2_X1 U16104 ( .A1(n16306), .A2(n15739), .ZN(n16304) );
  OR2_X1 U16105 ( .A1(a_4_), .A2(n15727), .ZN(n16306) );
  OR2_X1 U16106 ( .A1(n16307), .A2(n16308), .ZN(n15727) );
  AND2_X1 U16107 ( .A1(a_5_), .A2(n15693), .ZN(n16308) );
  AND2_X1 U16108 ( .A1(n16309), .A2(n15705), .ZN(n16307) );
  OR2_X1 U16109 ( .A1(a_5_), .A2(n15693), .ZN(n16309) );
  OR2_X1 U16110 ( .A1(n16310), .A2(n16311), .ZN(n15693) );
  AND2_X1 U16111 ( .A1(a_6_), .A2(n15659), .ZN(n16311) );
  AND2_X1 U16112 ( .A1(n16312), .A2(n15671), .ZN(n16310) );
  OR2_X1 U16113 ( .A1(a_6_), .A2(n15659), .ZN(n16312) );
  OR2_X1 U16114 ( .A1(n16313), .A2(n16314), .ZN(n15659) );
  AND2_X1 U16115 ( .A1(a_7_), .A2(n15625), .ZN(n16314) );
  AND2_X1 U16116 ( .A1(n16315), .A2(n15637), .ZN(n16313) );
  OR2_X1 U16117 ( .A1(a_7_), .A2(n15625), .ZN(n16315) );
  OR2_X1 U16118 ( .A1(n16316), .A2(n16317), .ZN(n15625) );
  AND2_X1 U16119 ( .A1(a_8_), .A2(n15580), .ZN(n16317) );
  AND2_X1 U16120 ( .A1(n16318), .A2(n15592), .ZN(n16316) );
  OR2_X1 U16121 ( .A1(a_8_), .A2(n15580), .ZN(n16318) );
  OR2_X1 U16122 ( .A1(n16319), .A2(n16320), .ZN(n15580) );
  AND2_X1 U16123 ( .A1(a_9_), .A2(n15546), .ZN(n16320) );
  AND2_X1 U16124 ( .A1(n16321), .A2(n15558), .ZN(n16319) );
  OR2_X1 U16125 ( .A1(a_9_), .A2(n15546), .ZN(n16321) );
  OR2_X1 U16126 ( .A1(n16322), .A2(n16323), .ZN(n15546) );
  AND2_X1 U16127 ( .A1(a_10_), .A2(n15512), .ZN(n16323) );
  AND2_X1 U16128 ( .A1(n16324), .A2(n15524), .ZN(n16322) );
  OR2_X1 U16129 ( .A1(a_10_), .A2(n15512), .ZN(n16324) );
  OR2_X1 U16130 ( .A1(n16325), .A2(n16326), .ZN(n15512) );
  AND2_X1 U16131 ( .A1(a_11_), .A2(n15478), .ZN(n16326) );
  AND2_X1 U16132 ( .A1(n16327), .A2(n15490), .ZN(n16325) );
  OR2_X1 U16133 ( .A1(a_11_), .A2(n15478), .ZN(n16327) );
  OR2_X1 U16134 ( .A1(n16328), .A2(n16329), .ZN(n15478) );
  AND2_X1 U16135 ( .A1(a_12_), .A2(n15444), .ZN(n16329) );
  AND2_X1 U16136 ( .A1(n16330), .A2(n15456), .ZN(n16328) );
  OR2_X1 U16137 ( .A1(a_12_), .A2(n15444), .ZN(n16330) );
  OR2_X1 U16138 ( .A1(n16331), .A2(n16332), .ZN(n15444) );
  AND2_X1 U16139 ( .A1(a_13_), .A2(n15410), .ZN(n16332) );
  AND2_X1 U16140 ( .A1(n16333), .A2(n15422), .ZN(n16331) );
  OR2_X1 U16141 ( .A1(a_13_), .A2(n15410), .ZN(n16333) );
  OR2_X1 U16142 ( .A1(n16334), .A2(n16335), .ZN(n15410) );
  AND2_X1 U16143 ( .A1(a_14_), .A2(n15376), .ZN(n16335) );
  AND2_X1 U16144 ( .A1(n16336), .A2(n15388), .ZN(n16334) );
  OR2_X1 U16145 ( .A1(a_14_), .A2(n15376), .ZN(n16336) );
  OR2_X1 U16146 ( .A1(n16337), .A2(n16338), .ZN(n15376) );
  AND2_X1 U16147 ( .A1(a_15_), .A2(n15342), .ZN(n16338) );
  AND2_X1 U16148 ( .A1(n16339), .A2(n15354), .ZN(n16337) );
  OR2_X1 U16149 ( .A1(a_15_), .A2(n15342), .ZN(n16339) );
  OR2_X1 U16150 ( .A1(n16340), .A2(n16341), .ZN(n15342) );
  AND2_X1 U16151 ( .A1(a_16_), .A2(n15308), .ZN(n16341) );
  AND2_X1 U16152 ( .A1(n16342), .A2(n15320), .ZN(n16340) );
  OR2_X1 U16153 ( .A1(a_16_), .A2(n15308), .ZN(n16342) );
  OR2_X1 U16154 ( .A1(n16343), .A2(n16344), .ZN(n15308) );
  AND2_X1 U16155 ( .A1(a_17_), .A2(n15274), .ZN(n16344) );
  AND2_X1 U16156 ( .A1(n16345), .A2(n15286), .ZN(n16343) );
  OR2_X1 U16157 ( .A1(a_17_), .A2(n15274), .ZN(n16345) );
  OR2_X1 U16158 ( .A1(n16346), .A2(n16347), .ZN(n15274) );
  AND2_X1 U16159 ( .A1(a_18_), .A2(n15229), .ZN(n16347) );
  AND2_X1 U16160 ( .A1(n16348), .A2(n15241), .ZN(n16346) );
  OR2_X1 U16161 ( .A1(a_18_), .A2(n15229), .ZN(n16348) );
  OR2_X1 U16162 ( .A1(n16349), .A2(n16350), .ZN(n15229) );
  AND2_X1 U16163 ( .A1(a_19_), .A2(n15195), .ZN(n16350) );
  AND2_X1 U16164 ( .A1(n16351), .A2(n15207), .ZN(n16349) );
  OR2_X1 U16165 ( .A1(a_19_), .A2(n15195), .ZN(n16351) );
  OR2_X1 U16166 ( .A1(n16352), .A2(n16353), .ZN(n15195) );
  AND2_X1 U16167 ( .A1(a_20_), .A2(n15161), .ZN(n16353) );
  AND2_X1 U16168 ( .A1(n16354), .A2(n15173), .ZN(n16352) );
  OR2_X1 U16169 ( .A1(a_20_), .A2(n15161), .ZN(n16354) );
  OR2_X1 U16170 ( .A1(n16355), .A2(n16356), .ZN(n15161) );
  AND2_X1 U16171 ( .A1(a_21_), .A2(n15127), .ZN(n16356) );
  AND2_X1 U16172 ( .A1(n16357), .A2(n15139), .ZN(n16355) );
  OR2_X1 U16173 ( .A1(a_21_), .A2(n15127), .ZN(n16357) );
  OR2_X1 U16174 ( .A1(n16358), .A2(n16359), .ZN(n15127) );
  AND2_X1 U16175 ( .A1(a_22_), .A2(n15093), .ZN(n16359) );
  AND2_X1 U16176 ( .A1(n16360), .A2(n15105), .ZN(n16358) );
  OR2_X1 U16177 ( .A1(a_22_), .A2(n15093), .ZN(n16360) );
  OR2_X1 U16178 ( .A1(n16361), .A2(n16362), .ZN(n15093) );
  AND2_X1 U16179 ( .A1(a_23_), .A2(n15059), .ZN(n16362) );
  AND2_X1 U16180 ( .A1(n16363), .A2(n15071), .ZN(n16361) );
  OR2_X1 U16181 ( .A1(a_23_), .A2(n15059), .ZN(n16363) );
  OR2_X1 U16182 ( .A1(n16364), .A2(n16365), .ZN(n15059) );
  AND2_X1 U16183 ( .A1(a_24_), .A2(n15025), .ZN(n16365) );
  AND2_X1 U16184 ( .A1(n16366), .A2(n15037), .ZN(n16364) );
  OR2_X1 U16185 ( .A1(a_24_), .A2(n15025), .ZN(n16366) );
  OR2_X1 U16186 ( .A1(n16367), .A2(n16368), .ZN(n15025) );
  AND2_X1 U16187 ( .A1(a_25_), .A2(n14991), .ZN(n16368) );
  AND2_X1 U16188 ( .A1(n16369), .A2(n15003), .ZN(n16367) );
  OR2_X1 U16189 ( .A1(a_25_), .A2(n14991), .ZN(n16369) );
  OR2_X1 U16190 ( .A1(n16370), .A2(n16371), .ZN(n14991) );
  AND2_X1 U16191 ( .A1(a_26_), .A2(n14957), .ZN(n16371) );
  AND2_X1 U16192 ( .A1(n16372), .A2(n14969), .ZN(n16370) );
  OR2_X1 U16193 ( .A1(a_26_), .A2(n14957), .ZN(n16372) );
  OR2_X1 U16194 ( .A1(n16373), .A2(n16374), .ZN(n14957) );
  AND2_X1 U16195 ( .A1(a_27_), .A2(n14923), .ZN(n16374) );
  AND2_X1 U16196 ( .A1(n16375), .A2(n14935), .ZN(n16373) );
  OR2_X1 U16197 ( .A1(a_27_), .A2(n14923), .ZN(n16375) );
  OR2_X1 U16198 ( .A1(n16376), .A2(n16377), .ZN(n14923) );
  AND2_X1 U16199 ( .A1(a_28_), .A2(n14878), .ZN(n16377) );
  AND2_X1 U16200 ( .A1(n16378), .A2(n14890), .ZN(n16376) );
  OR2_X1 U16201 ( .A1(a_28_), .A2(n14878), .ZN(n16378) );
  OR2_X1 U16202 ( .A1(n16379), .A2(n16380), .ZN(n14878) );
  AND2_X1 U16203 ( .A1(a_29_), .A2(n14844), .ZN(n16380) );
  AND2_X1 U16204 ( .A1(n16381), .A2(n14856), .ZN(n16379) );
  OR2_X1 U16205 ( .A1(a_29_), .A2(n14844), .ZN(n16381) );
  OR2_X1 U16206 ( .A1(n16382), .A2(n16383), .ZN(n14844) );
  AND2_X1 U16207 ( .A1(a_30_), .A2(n14794), .ZN(n16383) );
  AND2_X1 U16208 ( .A1(n16384), .A2(n14801), .ZN(n16382) );
  OR2_X1 U16209 ( .A1(n14794), .A2(a_30_), .ZN(n16384) );
  INV_X1 U16210 ( .A(n14814), .ZN(n14794) );
  OR2_X1 U16211 ( .A1(b_31_), .A2(n15958), .ZN(n14814) );
  AND2_X1 U16212 ( .A1(n16294), .A2(a_0_), .ZN(n15866) );
  AND2_X1 U16213 ( .A1(n14744), .A2(n16385), .ZN(n16197) );
  OR3_X1 U16214 ( .A1(n16386), .A2(n16387), .A3(n16388), .ZN(n16385) );
  AND2_X1 U16215 ( .A1(n16389), .A2(a_0_), .ZN(n16388) );
  AND2_X1 U16216 ( .A1(n16089), .A2(n16090), .ZN(n16387) );
  INV_X1 U16217 ( .A(n16094), .ZN(n16089) );
  OR2_X1 U16218 ( .A1(n16390), .A2(n15992), .ZN(n16094) );
  OR2_X1 U16219 ( .A1(n16391), .A2(n16093), .ZN(n15992) );
  AND2_X1 U16220 ( .A1(n16392), .A2(n16393), .ZN(n16391) );
  AND2_X1 U16221 ( .A1(n15991), .A2(n15989), .ZN(n16390) );
  OR2_X1 U16222 ( .A1(n16394), .A2(n15603), .ZN(n15989) );
  OR2_X1 U16223 ( .A1(n16395), .A2(n15993), .ZN(n15603) );
  INV_X1 U16224 ( .A(n15991), .ZN(n15993) );
  AND2_X1 U16225 ( .A1(n16396), .A2(n16397), .ZN(n16395) );
  AND2_X1 U16226 ( .A1(n15600), .A2(n15602), .ZN(n16394) );
  OR2_X1 U16227 ( .A1(n16398), .A2(n15252), .ZN(n15600) );
  OR2_X1 U16228 ( .A1(n16399), .A2(n15604), .ZN(n15252) );
  INV_X1 U16229 ( .A(n15602), .ZN(n15604) );
  OR2_X1 U16230 ( .A1(n16400), .A2(n16401), .ZN(n15602) );
  AND2_X1 U16231 ( .A1(n16400), .A2(n16401), .ZN(n16399) );
  OR2_X1 U16232 ( .A1(n16402), .A2(n16403), .ZN(n16401) );
  AND2_X1 U16233 ( .A1(n16404), .A2(n16405), .ZN(n16403) );
  AND2_X1 U16234 ( .A1(n16406), .A2(n16407), .ZN(n16402) );
  OR2_X1 U16235 ( .A1(n16405), .A2(n16404), .ZN(n16407) );
  AND2_X1 U16236 ( .A1(n16408), .A2(n16409), .ZN(n16400) );
  INV_X1 U16237 ( .A(n16410), .ZN(n16409) );
  AND2_X1 U16238 ( .A1(n16411), .A2(n16412), .ZN(n16410) );
  OR2_X1 U16239 ( .A1(n16412), .A2(n16411), .ZN(n16408) );
  OR2_X1 U16240 ( .A1(n16413), .A2(n16414), .ZN(n16411) );
  AND2_X1 U16241 ( .A1(n16415), .A2(n16416), .ZN(n16414) );
  INV_X1 U16242 ( .A(n16417), .ZN(n16415) );
  AND2_X1 U16243 ( .A1(n16418), .A2(n16417), .ZN(n16413) );
  INV_X1 U16244 ( .A(n16416), .ZN(n16418) );
  AND2_X1 U16245 ( .A1(n15251), .A2(n15249), .ZN(n16398) );
  OR2_X1 U16246 ( .A1(n16419), .A2(n14901), .ZN(n15249) );
  OR2_X1 U16247 ( .A1(n16420), .A2(n15253), .ZN(n14901) );
  INV_X1 U16248 ( .A(n15251), .ZN(n15253) );
  AND2_X1 U16249 ( .A1(n16421), .A2(n16422), .ZN(n16420) );
  AND2_X1 U16250 ( .A1(n14898), .A2(n14900), .ZN(n16419) );
  OR2_X1 U16251 ( .A1(n16423), .A2(n14784), .ZN(n14898) );
  OR2_X1 U16252 ( .A1(n16424), .A2(n14902), .ZN(n14784) );
  INV_X1 U16253 ( .A(n14900), .ZN(n14902) );
  OR2_X1 U16254 ( .A1(n16425), .A2(n16426), .ZN(n14900) );
  AND2_X1 U16255 ( .A1(n16425), .A2(n16426), .ZN(n16424) );
  OR2_X1 U16256 ( .A1(n16427), .A2(n16428), .ZN(n16426) );
  AND2_X1 U16257 ( .A1(n16429), .A2(n16430), .ZN(n16428) );
  AND2_X1 U16258 ( .A1(n16431), .A2(n16432), .ZN(n16427) );
  OR2_X1 U16259 ( .A1(n16430), .A2(n16429), .ZN(n16432) );
  AND2_X1 U16260 ( .A1(n16433), .A2(n16434), .ZN(n16425) );
  INV_X1 U16261 ( .A(n16435), .ZN(n16434) );
  AND2_X1 U16262 ( .A1(n16436), .A2(n16437), .ZN(n16435) );
  OR2_X1 U16263 ( .A1(n16437), .A2(n16436), .ZN(n16433) );
  OR2_X1 U16264 ( .A1(n16438), .A2(n16439), .ZN(n16436) );
  AND2_X1 U16265 ( .A1(n16440), .A2(n16441), .ZN(n16439) );
  INV_X1 U16266 ( .A(n16442), .ZN(n16440) );
  AND2_X1 U16267 ( .A1(n16443), .A2(n16442), .ZN(n16438) );
  INV_X1 U16268 ( .A(n16441), .ZN(n16443) );
  AND2_X1 U16269 ( .A1(n14783), .A2(n14781), .ZN(n16423) );
  OR2_X1 U16270 ( .A1(n16444), .A2(n14773), .ZN(n14781) );
  OR2_X1 U16271 ( .A1(n16445), .A2(n14785), .ZN(n14773) );
  INV_X1 U16272 ( .A(n14783), .ZN(n14785) );
  AND2_X1 U16273 ( .A1(n16446), .A2(n16447), .ZN(n16445) );
  AND2_X1 U16274 ( .A1(n14770), .A2(n14772), .ZN(n16444) );
  OR2_X1 U16275 ( .A1(n16448), .A2(n14762), .ZN(n14770) );
  OR2_X1 U16276 ( .A1(n16449), .A2(n14774), .ZN(n14762) );
  INV_X1 U16277 ( .A(n14772), .ZN(n14774) );
  OR2_X1 U16278 ( .A1(n16450), .A2(n16451), .ZN(n14772) );
  AND2_X1 U16279 ( .A1(n16450), .A2(n16451), .ZN(n16449) );
  OR2_X1 U16280 ( .A1(n16452), .A2(n16453), .ZN(n16451) );
  AND2_X1 U16281 ( .A1(n16454), .A2(n16455), .ZN(n16453) );
  AND2_X1 U16282 ( .A1(n16456), .A2(n16457), .ZN(n16452) );
  OR2_X1 U16283 ( .A1(n16455), .A2(n16454), .ZN(n16457) );
  AND2_X1 U16284 ( .A1(n16458), .A2(n16459), .ZN(n16450) );
  INV_X1 U16285 ( .A(n16460), .ZN(n16459) );
  AND2_X1 U16286 ( .A1(n16461), .A2(n16462), .ZN(n16460) );
  OR2_X1 U16287 ( .A1(n16462), .A2(n16461), .ZN(n16458) );
  OR2_X1 U16288 ( .A1(n16463), .A2(n16464), .ZN(n16461) );
  AND2_X1 U16289 ( .A1(n16465), .A2(n16466), .ZN(n16464) );
  INV_X1 U16290 ( .A(n16467), .ZN(n16465) );
  AND2_X1 U16291 ( .A1(n16468), .A2(n16467), .ZN(n16463) );
  INV_X1 U16292 ( .A(n16466), .ZN(n16468) );
  AND2_X1 U16293 ( .A1(n14761), .A2(n14759), .ZN(n16448) );
  OR2_X1 U16294 ( .A1(n16469), .A2(n14750), .ZN(n14759) );
  OR2_X1 U16295 ( .A1(n16470), .A2(n14763), .ZN(n14750) );
  INV_X1 U16296 ( .A(n14761), .ZN(n14763) );
  AND2_X1 U16297 ( .A1(n16471), .A2(n16472), .ZN(n16470) );
  AND2_X1 U16298 ( .A1(n14748), .A2(n14752), .ZN(n16469) );
  OR2_X1 U16299 ( .A1(n16473), .A2(n16194), .ZN(n14748) );
  OR2_X1 U16300 ( .A1(n16474), .A2(n14749), .ZN(n16194) );
  INV_X1 U16301 ( .A(n14752), .ZN(n14749) );
  OR2_X1 U16302 ( .A1(n16475), .A2(n16476), .ZN(n14752) );
  AND2_X1 U16303 ( .A1(n16475), .A2(n16476), .ZN(n16474) );
  OR2_X1 U16304 ( .A1(n16477), .A2(n16478), .ZN(n16476) );
  AND2_X1 U16305 ( .A1(n16479), .A2(n16480), .ZN(n16478) );
  AND2_X1 U16306 ( .A1(n16481), .A2(n16482), .ZN(n16477) );
  OR2_X1 U16307 ( .A1(n16479), .A2(n16480), .ZN(n16482) );
  AND2_X1 U16308 ( .A1(n16483), .A2(n16484), .ZN(n16475) );
  INV_X1 U16309 ( .A(n16485), .ZN(n16484) );
  AND2_X1 U16310 ( .A1(n16486), .A2(n16487), .ZN(n16485) );
  OR2_X1 U16311 ( .A1(n16487), .A2(n16486), .ZN(n16483) );
  OR2_X1 U16312 ( .A1(n16488), .A2(n16489), .ZN(n16486) );
  AND2_X1 U16313 ( .A1(n16490), .A2(n16491), .ZN(n16489) );
  INV_X1 U16314 ( .A(n16492), .ZN(n16490) );
  AND2_X1 U16315 ( .A1(n16493), .A2(n16492), .ZN(n16488) );
  INV_X1 U16316 ( .A(n16491), .ZN(n16493) );
  AND2_X1 U16317 ( .A1(n16192), .A2(n16196), .ZN(n16473) );
  OR2_X1 U16318 ( .A1(n16494), .A2(n16179), .ZN(n16192) );
  OR2_X1 U16319 ( .A1(n16495), .A2(n16193), .ZN(n16179) );
  INV_X1 U16320 ( .A(n16196), .ZN(n16193) );
  OR2_X1 U16321 ( .A1(n16496), .A2(n16497), .ZN(n16196) );
  AND2_X1 U16322 ( .A1(n16496), .A2(n16497), .ZN(n16495) );
  OR2_X1 U16323 ( .A1(n16498), .A2(n16499), .ZN(n16497) );
  AND2_X1 U16324 ( .A1(n16500), .A2(n16501), .ZN(n16499) );
  AND2_X1 U16325 ( .A1(n16502), .A2(n16503), .ZN(n16498) );
  OR2_X1 U16326 ( .A1(n16500), .A2(n16501), .ZN(n16503) );
  AND2_X1 U16327 ( .A1(n16504), .A2(n16505), .ZN(n16496) );
  INV_X1 U16328 ( .A(n16506), .ZN(n16505) );
  AND2_X1 U16329 ( .A1(n16507), .A2(n16481), .ZN(n16506) );
  OR2_X1 U16330 ( .A1(n16481), .A2(n16507), .ZN(n16504) );
  OR2_X1 U16331 ( .A1(n16508), .A2(n16509), .ZN(n16507) );
  AND2_X1 U16332 ( .A1(n16510), .A2(n16480), .ZN(n16509) );
  INV_X1 U16333 ( .A(n16479), .ZN(n16510) );
  AND2_X1 U16334 ( .A1(n16511), .A2(n16479), .ZN(n16508) );
  OR2_X1 U16335 ( .A1(n16512), .A2(n15524), .ZN(n16479) );
  INV_X1 U16336 ( .A(n16480), .ZN(n16511) );
  OR2_X1 U16337 ( .A1(n16513), .A2(n16514), .ZN(n16480) );
  AND2_X1 U16338 ( .A1(n16515), .A2(n16516), .ZN(n16514) );
  AND2_X1 U16339 ( .A1(n16517), .A2(n16518), .ZN(n16513) );
  OR2_X1 U16340 ( .A1(n16515), .A2(n16516), .ZN(n16518) );
  AND2_X1 U16341 ( .A1(n16519), .A2(n16520), .ZN(n16481) );
  INV_X1 U16342 ( .A(n16521), .ZN(n16520) );
  AND2_X1 U16343 ( .A1(n16522), .A2(n16523), .ZN(n16521) );
  OR2_X1 U16344 ( .A1(n16523), .A2(n16522), .ZN(n16519) );
  OR2_X1 U16345 ( .A1(n16524), .A2(n16525), .ZN(n16522) );
  AND2_X1 U16346 ( .A1(n16526), .A2(n16527), .ZN(n16525) );
  INV_X1 U16347 ( .A(n16528), .ZN(n16526) );
  AND2_X1 U16348 ( .A1(n16529), .A2(n16528), .ZN(n16524) );
  INV_X1 U16349 ( .A(n16527), .ZN(n16529) );
  AND2_X1 U16350 ( .A1(n16178), .A2(n16184), .ZN(n16494) );
  OR2_X1 U16351 ( .A1(n16530), .A2(n16531), .ZN(n16184) );
  INV_X1 U16352 ( .A(n16532), .ZN(n16530) );
  AND2_X1 U16353 ( .A1(n16533), .A2(n16170), .ZN(n16178) );
  OR2_X1 U16354 ( .A1(n16174), .A2(n16534), .ZN(n16170) );
  OR2_X1 U16355 ( .A1(n16168), .A2(n16174), .ZN(n16533) );
  AND2_X1 U16356 ( .A1(n16535), .A2(n16536), .ZN(n16174) );
  INV_X1 U16357 ( .A(n16537), .ZN(n16536) );
  AND2_X1 U16358 ( .A1(n16532), .A2(n16531), .ZN(n16537) );
  OR2_X1 U16359 ( .A1(n16532), .A2(n16531), .ZN(n16535) );
  OR2_X1 U16360 ( .A1(n16538), .A2(n16539), .ZN(n16531) );
  AND2_X1 U16361 ( .A1(n16540), .A2(n16541), .ZN(n16539) );
  AND2_X1 U16362 ( .A1(n16542), .A2(n16543), .ZN(n16538) );
  OR2_X1 U16363 ( .A1(n16541), .A2(n16540), .ZN(n16543) );
  OR2_X1 U16364 ( .A1(n16544), .A2(n16545), .ZN(n16532) );
  AND2_X1 U16365 ( .A1(n16546), .A2(n16502), .ZN(n16545) );
  INV_X1 U16366 ( .A(n16547), .ZN(n16544) );
  OR2_X1 U16367 ( .A1(n16502), .A2(n16546), .ZN(n16547) );
  OR2_X1 U16368 ( .A1(n16548), .A2(n16549), .ZN(n16546) );
  AND2_X1 U16369 ( .A1(n16550), .A2(n16501), .ZN(n16549) );
  INV_X1 U16370 ( .A(n16500), .ZN(n16550) );
  AND2_X1 U16371 ( .A1(n16551), .A2(n16500), .ZN(n16548) );
  OR2_X1 U16372 ( .A1(n16512), .A2(n15490), .ZN(n16500) );
  INV_X1 U16373 ( .A(n16501), .ZN(n16551) );
  OR2_X1 U16374 ( .A1(n16552), .A2(n16553), .ZN(n16501) );
  AND2_X1 U16375 ( .A1(n16554), .A2(n16555), .ZN(n16553) );
  AND2_X1 U16376 ( .A1(n16556), .A2(n16557), .ZN(n16552) );
  OR2_X1 U16377 ( .A1(n16554), .A2(n16555), .ZN(n16557) );
  AND2_X1 U16378 ( .A1(n16558), .A2(n16559), .ZN(n16502) );
  INV_X1 U16379 ( .A(n16560), .ZN(n16559) );
  AND2_X1 U16380 ( .A1(n16561), .A2(n16517), .ZN(n16560) );
  OR2_X1 U16381 ( .A1(n16517), .A2(n16561), .ZN(n16558) );
  OR2_X1 U16382 ( .A1(n16562), .A2(n16563), .ZN(n16561) );
  AND2_X1 U16383 ( .A1(n16564), .A2(n16516), .ZN(n16563) );
  INV_X1 U16384 ( .A(n16515), .ZN(n16564) );
  AND2_X1 U16385 ( .A1(n16565), .A2(n16515), .ZN(n16562) );
  OR2_X1 U16386 ( .A1(n15842), .A2(n15524), .ZN(n16515) );
  INV_X1 U16387 ( .A(n16516), .ZN(n16565) );
  OR2_X1 U16388 ( .A1(n16566), .A2(n16567), .ZN(n16516) );
  AND2_X1 U16389 ( .A1(n16568), .A2(n16569), .ZN(n16567) );
  AND2_X1 U16390 ( .A1(n16570), .A2(n16571), .ZN(n16566) );
  OR2_X1 U16391 ( .A1(n16568), .A2(n16569), .ZN(n16571) );
  AND2_X1 U16392 ( .A1(n16572), .A2(n16573), .ZN(n16517) );
  INV_X1 U16393 ( .A(n16574), .ZN(n16573) );
  AND2_X1 U16394 ( .A1(n16575), .A2(n16576), .ZN(n16574) );
  OR2_X1 U16395 ( .A1(n16576), .A2(n16575), .ZN(n16572) );
  OR2_X1 U16396 ( .A1(n16577), .A2(n16578), .ZN(n16575) );
  AND2_X1 U16397 ( .A1(n16579), .A2(n16580), .ZN(n16578) );
  INV_X1 U16398 ( .A(n16581), .ZN(n16579) );
  AND2_X1 U16399 ( .A1(n16582), .A2(n16581), .ZN(n16577) );
  INV_X1 U16400 ( .A(n16580), .ZN(n16582) );
  OR2_X1 U16401 ( .A1(n16583), .A2(n16156), .ZN(n16168) );
  OR2_X1 U16402 ( .A1(n16584), .A2(n16173), .ZN(n16156) );
  INV_X1 U16403 ( .A(n16534), .ZN(n16173) );
  OR2_X1 U16404 ( .A1(n16585), .A2(n16586), .ZN(n16534) );
  AND2_X1 U16405 ( .A1(n16585), .A2(n16586), .ZN(n16584) );
  OR2_X1 U16406 ( .A1(n16587), .A2(n16588), .ZN(n16586) );
  AND2_X1 U16407 ( .A1(n16589), .A2(n16590), .ZN(n16588) );
  AND2_X1 U16408 ( .A1(n16591), .A2(n16592), .ZN(n16587) );
  OR2_X1 U16409 ( .A1(n16589), .A2(n16590), .ZN(n16592) );
  AND2_X1 U16410 ( .A1(n16593), .A2(n16594), .ZN(n16585) );
  INV_X1 U16411 ( .A(n16595), .ZN(n16594) );
  AND2_X1 U16412 ( .A1(n16596), .A2(n16542), .ZN(n16595) );
  OR2_X1 U16413 ( .A1(n16542), .A2(n16596), .ZN(n16593) );
  OR2_X1 U16414 ( .A1(n16597), .A2(n16598), .ZN(n16596) );
  AND2_X1 U16415 ( .A1(n16599), .A2(n16541), .ZN(n16598) );
  INV_X1 U16416 ( .A(n16540), .ZN(n16599) );
  AND2_X1 U16417 ( .A1(n16600), .A2(n16540), .ZN(n16597) );
  OR2_X1 U16418 ( .A1(n16512), .A2(n15456), .ZN(n16540) );
  INV_X1 U16419 ( .A(n16541), .ZN(n16600) );
  OR2_X1 U16420 ( .A1(n16601), .A2(n16602), .ZN(n16541) );
  AND2_X1 U16421 ( .A1(n16603), .A2(n16604), .ZN(n16602) );
  AND2_X1 U16422 ( .A1(n16605), .A2(n16606), .ZN(n16601) );
  OR2_X1 U16423 ( .A1(n16604), .A2(n16603), .ZN(n16606) );
  AND2_X1 U16424 ( .A1(n16607), .A2(n16608), .ZN(n16542) );
  INV_X1 U16425 ( .A(n16609), .ZN(n16608) );
  AND2_X1 U16426 ( .A1(n16610), .A2(n16556), .ZN(n16609) );
  OR2_X1 U16427 ( .A1(n16556), .A2(n16610), .ZN(n16607) );
  OR2_X1 U16428 ( .A1(n16611), .A2(n16612), .ZN(n16610) );
  AND2_X1 U16429 ( .A1(n16613), .A2(n16555), .ZN(n16612) );
  INV_X1 U16430 ( .A(n16554), .ZN(n16613) );
  AND2_X1 U16431 ( .A1(n16614), .A2(n16554), .ZN(n16611) );
  OR2_X1 U16432 ( .A1(n15842), .A2(n15490), .ZN(n16554) );
  INV_X1 U16433 ( .A(n16555), .ZN(n16614) );
  OR2_X1 U16434 ( .A1(n16615), .A2(n16616), .ZN(n16555) );
  AND2_X1 U16435 ( .A1(n16617), .A2(n16618), .ZN(n16616) );
  AND2_X1 U16436 ( .A1(n16619), .A2(n16620), .ZN(n16615) );
  OR2_X1 U16437 ( .A1(n16617), .A2(n16618), .ZN(n16620) );
  AND2_X1 U16438 ( .A1(n16621), .A2(n16622), .ZN(n16556) );
  INV_X1 U16439 ( .A(n16623), .ZN(n16622) );
  AND2_X1 U16440 ( .A1(n16624), .A2(n16570), .ZN(n16623) );
  OR2_X1 U16441 ( .A1(n16570), .A2(n16624), .ZN(n16621) );
  OR2_X1 U16442 ( .A1(n16625), .A2(n16626), .ZN(n16624) );
  AND2_X1 U16443 ( .A1(n16627), .A2(n16569), .ZN(n16626) );
  INV_X1 U16444 ( .A(n16568), .ZN(n16627) );
  AND2_X1 U16445 ( .A1(n16628), .A2(n16568), .ZN(n16625) );
  OR2_X1 U16446 ( .A1(n15808), .A2(n15524), .ZN(n16568) );
  INV_X1 U16447 ( .A(n16569), .ZN(n16628) );
  OR2_X1 U16448 ( .A1(n16629), .A2(n16630), .ZN(n16569) );
  AND2_X1 U16449 ( .A1(n16631), .A2(n16632), .ZN(n16630) );
  AND2_X1 U16450 ( .A1(n16633), .A2(n16634), .ZN(n16629) );
  OR2_X1 U16451 ( .A1(n16631), .A2(n16632), .ZN(n16634) );
  AND2_X1 U16452 ( .A1(n16635), .A2(n16636), .ZN(n16570) );
  INV_X1 U16453 ( .A(n16637), .ZN(n16636) );
  AND2_X1 U16454 ( .A1(n16638), .A2(n16639), .ZN(n16637) );
  OR2_X1 U16455 ( .A1(n16639), .A2(n16638), .ZN(n16635) );
  OR2_X1 U16456 ( .A1(n16640), .A2(n16641), .ZN(n16638) );
  AND2_X1 U16457 ( .A1(n16642), .A2(n16643), .ZN(n16641) );
  INV_X1 U16458 ( .A(n16644), .ZN(n16642) );
  AND2_X1 U16459 ( .A1(n16645), .A2(n16644), .ZN(n16640) );
  INV_X1 U16460 ( .A(n16643), .ZN(n16645) );
  AND2_X1 U16461 ( .A1(n16155), .A2(n16162), .ZN(n16583) );
  INV_X1 U16462 ( .A(n16160), .ZN(n16162) );
  AND2_X1 U16463 ( .A1(n16646), .A2(n16647), .ZN(n16160) );
  INV_X1 U16464 ( .A(n16648), .ZN(n16647) );
  AND2_X1 U16465 ( .A1(n16649), .A2(n16151), .ZN(n16155) );
  OR2_X1 U16466 ( .A1(n16149), .A2(n16150), .ZN(n16151) );
  OR2_X1 U16467 ( .A1(n16149), .A2(n16146), .ZN(n16649) );
  AND2_X1 U16468 ( .A1(n16137), .A2(n16650), .ZN(n16146) );
  OR2_X1 U16469 ( .A1(n16140), .A2(n16651), .ZN(n16650) );
  INV_X1 U16470 ( .A(n16134), .ZN(n16651) );
  OR2_X1 U16471 ( .A1(n16127), .A2(n16652), .ZN(n16134) );
  AND2_X1 U16472 ( .A1(n16128), .A2(n16123), .ZN(n16652) );
  OR2_X1 U16473 ( .A1(n16653), .A2(n16118), .ZN(n16123) );
  INV_X1 U16474 ( .A(n16654), .ZN(n16118) );
  OR4_X1 U16475 ( .A1(n16655), .A2(n16656), .A3(n16129), .A4(n16657), .ZN(
        n16654) );
  INV_X1 U16476 ( .A(n16658), .ZN(n16653) );
  OR2_X1 U16477 ( .A1(n16116), .A2(n16117), .ZN(n16658) );
  AND2_X1 U16478 ( .A1(n16659), .A2(n16660), .ZN(n16117) );
  OR2_X1 U16479 ( .A1(n16656), .A2(n16655), .ZN(n16660) );
  OR2_X1 U16480 ( .A1(n16657), .A2(n16129), .ZN(n16659) );
  AND2_X1 U16481 ( .A1(n16661), .A2(n16662), .ZN(n16657) );
  AND2_X1 U16482 ( .A1(n16105), .A2(n16110), .ZN(n16116) );
  INV_X1 U16483 ( .A(n16663), .ZN(n16110) );
  AND3_X1 U16484 ( .A1(n16664), .A2(n16665), .A3(n16666), .ZN(n16663) );
  INV_X1 U16485 ( .A(n16667), .ZN(n16105) );
  AND2_X1 U16486 ( .A1(n16109), .A2(n16108), .ZN(n16667) );
  OR2_X1 U16487 ( .A1(n16668), .A2(n16103), .ZN(n16108) );
  AND3_X1 U16488 ( .A1(n16669), .A2(n16670), .A3(n16671), .ZN(n16103) );
  AND2_X1 U16489 ( .A1(n16099), .A2(n16101), .ZN(n16668) );
  OR2_X1 U16490 ( .A1(n16672), .A2(n16670), .ZN(n16101) );
  OR2_X1 U16491 ( .A1(n16673), .A2(n16674), .ZN(n16670) );
  AND2_X1 U16492 ( .A1(n16664), .A2(n16675), .ZN(n16674) );
  AND2_X1 U16493 ( .A1(n16676), .A2(n16666), .ZN(n16673) );
  AND2_X1 U16494 ( .A1(n16671), .A2(n16669), .ZN(n16672) );
  OR2_X1 U16495 ( .A1(n16677), .A2(n16083), .ZN(n16099) );
  AND3_X1 U16496 ( .A1(n16678), .A2(n16679), .A3(n16680), .ZN(n16083) );
  AND2_X1 U16497 ( .A1(n16079), .A2(n16081), .ZN(n16677) );
  OR2_X1 U16498 ( .A1(n16681), .A2(n16679), .ZN(n16081) );
  OR2_X1 U16499 ( .A1(n16682), .A2(n16683), .ZN(n16679) );
  AND2_X1 U16500 ( .A1(n16669), .A2(n16684), .ZN(n16683) );
  INV_X1 U16501 ( .A(n16685), .ZN(n16669) );
  AND2_X1 U16502 ( .A1(n16685), .A2(n16671), .ZN(n16682) );
  INV_X1 U16503 ( .A(n16684), .ZN(n16671) );
  OR2_X1 U16504 ( .A1(n16686), .A2(n16687), .ZN(n16684) );
  AND2_X1 U16505 ( .A1(n16688), .A2(n16689), .ZN(n16687) );
  AND2_X1 U16506 ( .A1(n16690), .A2(n16691), .ZN(n16686) );
  OR2_X1 U16507 ( .A1(n16688), .A2(n16689), .ZN(n16691) );
  AND2_X1 U16508 ( .A1(n16692), .A2(n16693), .ZN(n16685) );
  INV_X1 U16509 ( .A(n16694), .ZN(n16693) );
  AND2_X1 U16510 ( .A1(n16695), .A2(n16696), .ZN(n16694) );
  OR2_X1 U16511 ( .A1(n16696), .A2(n16695), .ZN(n16692) );
  OR2_X1 U16512 ( .A1(n16697), .A2(n16698), .ZN(n16695) );
  AND2_X1 U16513 ( .A1(n16699), .A2(n16700), .ZN(n16698) );
  INV_X1 U16514 ( .A(n16701), .ZN(n16699) );
  AND2_X1 U16515 ( .A1(n16702), .A2(n16701), .ZN(n16697) );
  INV_X1 U16516 ( .A(n16700), .ZN(n16702) );
  AND2_X1 U16517 ( .A1(n16680), .A2(n16678), .ZN(n16681) );
  OR2_X1 U16518 ( .A1(n16074), .A2(n16073), .ZN(n16079) );
  AND3_X1 U16519 ( .A1(n16703), .A2(n16704), .A3(n16705), .ZN(n16073) );
  AND2_X1 U16520 ( .A1(n16070), .A2(n16071), .ZN(n16074) );
  OR2_X1 U16521 ( .A1(n16706), .A2(n16704), .ZN(n16071) );
  OR2_X1 U16522 ( .A1(n16707), .A2(n16708), .ZN(n16704) );
  AND2_X1 U16523 ( .A1(n16678), .A2(n16709), .ZN(n16708) );
  INV_X1 U16524 ( .A(n16710), .ZN(n16678) );
  AND2_X1 U16525 ( .A1(n16710), .A2(n16680), .ZN(n16707) );
  INV_X1 U16526 ( .A(n16709), .ZN(n16680) );
  OR2_X1 U16527 ( .A1(n16711), .A2(n16712), .ZN(n16709) );
  AND2_X1 U16528 ( .A1(n16713), .A2(n16714), .ZN(n16712) );
  AND2_X1 U16529 ( .A1(n16715), .A2(n16716), .ZN(n16711) );
  OR2_X1 U16530 ( .A1(n16713), .A2(n16714), .ZN(n16716) );
  AND2_X1 U16531 ( .A1(n16717), .A2(n16718), .ZN(n16710) );
  INV_X1 U16532 ( .A(n16719), .ZN(n16718) );
  AND2_X1 U16533 ( .A1(n16720), .A2(n16690), .ZN(n16719) );
  OR2_X1 U16534 ( .A1(n16690), .A2(n16720), .ZN(n16717) );
  OR2_X1 U16535 ( .A1(n16721), .A2(n16722), .ZN(n16720) );
  AND2_X1 U16536 ( .A1(n16723), .A2(n16689), .ZN(n16722) );
  INV_X1 U16537 ( .A(n16688), .ZN(n16723) );
  AND2_X1 U16538 ( .A1(n16724), .A2(n16688), .ZN(n16721) );
  OR2_X1 U16539 ( .A1(n16512), .A2(n15173), .ZN(n16688) );
  INV_X1 U16540 ( .A(n16689), .ZN(n16724) );
  OR2_X1 U16541 ( .A1(n16725), .A2(n16726), .ZN(n16689) );
  AND2_X1 U16542 ( .A1(n16727), .A2(n16728), .ZN(n16726) );
  AND2_X1 U16543 ( .A1(n16729), .A2(n16730), .ZN(n16725) );
  OR2_X1 U16544 ( .A1(n16727), .A2(n16728), .ZN(n16730) );
  AND2_X1 U16545 ( .A1(n16731), .A2(n16732), .ZN(n16690) );
  INV_X1 U16546 ( .A(n16733), .ZN(n16732) );
  AND2_X1 U16547 ( .A1(n16734), .A2(n16735), .ZN(n16733) );
  OR2_X1 U16548 ( .A1(n16735), .A2(n16734), .ZN(n16731) );
  OR2_X1 U16549 ( .A1(n16736), .A2(n16737), .ZN(n16734) );
  AND2_X1 U16550 ( .A1(n16738), .A2(n16739), .ZN(n16737) );
  INV_X1 U16551 ( .A(n16740), .ZN(n16738) );
  AND2_X1 U16552 ( .A1(n16741), .A2(n16740), .ZN(n16736) );
  INV_X1 U16553 ( .A(n16739), .ZN(n16741) );
  AND2_X1 U16554 ( .A1(n16705), .A2(n16703), .ZN(n16706) );
  OR2_X1 U16555 ( .A1(n16065), .A2(n16064), .ZN(n16070) );
  AND3_X1 U16556 ( .A1(n16742), .A2(n16743), .A3(n16744), .ZN(n16064) );
  AND2_X1 U16557 ( .A1(n16062), .A2(n16061), .ZN(n16065) );
  OR2_X1 U16558 ( .A1(n16745), .A2(n16056), .ZN(n16061) );
  AND3_X1 U16559 ( .A1(n16746), .A2(n16747), .A3(n16748), .ZN(n16056) );
  AND2_X1 U16560 ( .A1(n16052), .A2(n16054), .ZN(n16745) );
  OR2_X1 U16561 ( .A1(n16749), .A2(n16747), .ZN(n16054) );
  OR2_X1 U16562 ( .A1(n16750), .A2(n16751), .ZN(n16747) );
  AND2_X1 U16563 ( .A1(n16742), .A2(n16752), .ZN(n16751) );
  AND2_X1 U16564 ( .A1(n16753), .A2(n16744), .ZN(n16750) );
  AND2_X1 U16565 ( .A1(n16748), .A2(n16746), .ZN(n16749) );
  OR2_X1 U16566 ( .A1(n16754), .A2(n16047), .ZN(n16052) );
  AND3_X1 U16567 ( .A1(n16755), .A2(n16756), .A3(n16757), .ZN(n16047) );
  AND2_X1 U16568 ( .A1(n16043), .A2(n16045), .ZN(n16754) );
  OR2_X1 U16569 ( .A1(n16758), .A2(n16756), .ZN(n16045) );
  OR2_X1 U16570 ( .A1(n16759), .A2(n16760), .ZN(n16756) );
  AND2_X1 U16571 ( .A1(n16746), .A2(n16761), .ZN(n16760) );
  INV_X1 U16572 ( .A(n16762), .ZN(n16746) );
  AND2_X1 U16573 ( .A1(n16762), .A2(n16748), .ZN(n16759) );
  INV_X1 U16574 ( .A(n16761), .ZN(n16748) );
  OR2_X1 U16575 ( .A1(n16763), .A2(n16764), .ZN(n16761) );
  AND2_X1 U16576 ( .A1(n16765), .A2(n16766), .ZN(n16764) );
  AND2_X1 U16577 ( .A1(n16767), .A2(n16768), .ZN(n16763) );
  OR2_X1 U16578 ( .A1(n16765), .A2(n16766), .ZN(n16768) );
  AND2_X1 U16579 ( .A1(n16769), .A2(n16770), .ZN(n16762) );
  INV_X1 U16580 ( .A(n16771), .ZN(n16770) );
  AND2_X1 U16581 ( .A1(n16772), .A2(n16773), .ZN(n16771) );
  OR2_X1 U16582 ( .A1(n16773), .A2(n16772), .ZN(n16769) );
  OR2_X1 U16583 ( .A1(n16774), .A2(n16775), .ZN(n16772) );
  AND2_X1 U16584 ( .A1(n16776), .A2(n16777), .ZN(n16775) );
  INV_X1 U16585 ( .A(n16778), .ZN(n16776) );
  AND2_X1 U16586 ( .A1(n16779), .A2(n16778), .ZN(n16774) );
  INV_X1 U16587 ( .A(n16777), .ZN(n16779) );
  AND2_X1 U16588 ( .A1(n16757), .A2(n16755), .ZN(n16758) );
  OR2_X1 U16589 ( .A1(n16038), .A2(n16037), .ZN(n16043) );
  AND2_X1 U16590 ( .A1(n16780), .A2(n16781), .ZN(n16037) );
  AND2_X1 U16591 ( .A1(n16034), .A2(n16035), .ZN(n16038) );
  OR2_X1 U16592 ( .A1(n16781), .A2(n16780), .ZN(n16035) );
  OR2_X1 U16593 ( .A1(n16782), .A2(n16783), .ZN(n16780) );
  AND2_X1 U16594 ( .A1(n16755), .A2(n16784), .ZN(n16783) );
  INV_X1 U16595 ( .A(n16785), .ZN(n16755) );
  AND2_X1 U16596 ( .A1(n16785), .A2(n16757), .ZN(n16782) );
  INV_X1 U16597 ( .A(n16784), .ZN(n16757) );
  OR2_X1 U16598 ( .A1(n16786), .A2(n16787), .ZN(n16784) );
  AND2_X1 U16599 ( .A1(n16788), .A2(n16789), .ZN(n16787) );
  AND2_X1 U16600 ( .A1(n16790), .A2(n16791), .ZN(n16786) );
  OR2_X1 U16601 ( .A1(n16788), .A2(n16789), .ZN(n16791) );
  AND2_X1 U16602 ( .A1(n16792), .A2(n16793), .ZN(n16785) );
  INV_X1 U16603 ( .A(n16794), .ZN(n16793) );
  AND2_X1 U16604 ( .A1(n16795), .A2(n16767), .ZN(n16794) );
  OR2_X1 U16605 ( .A1(n16767), .A2(n16795), .ZN(n16792) );
  OR2_X1 U16606 ( .A1(n16796), .A2(n16797), .ZN(n16795) );
  AND2_X1 U16607 ( .A1(n16798), .A2(n16766), .ZN(n16797) );
  INV_X1 U16608 ( .A(n16765), .ZN(n16798) );
  AND2_X1 U16609 ( .A1(n16799), .A2(n16765), .ZN(n16796) );
  OR2_X1 U16610 ( .A1(n16512), .A2(n15037), .ZN(n16765) );
  INV_X1 U16611 ( .A(n16766), .ZN(n16799) );
  OR2_X1 U16612 ( .A1(n16800), .A2(n16801), .ZN(n16766) );
  AND2_X1 U16613 ( .A1(n16802), .A2(n16803), .ZN(n16801) );
  AND2_X1 U16614 ( .A1(n16804), .A2(n16805), .ZN(n16800) );
  OR2_X1 U16615 ( .A1(n16802), .A2(n16803), .ZN(n16805) );
  AND2_X1 U16616 ( .A1(n16806), .A2(n16807), .ZN(n16767) );
  INV_X1 U16617 ( .A(n16808), .ZN(n16807) );
  AND2_X1 U16618 ( .A1(n16809), .A2(n16810), .ZN(n16808) );
  OR2_X1 U16619 ( .A1(n16810), .A2(n16809), .ZN(n16806) );
  OR2_X1 U16620 ( .A1(n16811), .A2(n16812), .ZN(n16809) );
  AND2_X1 U16621 ( .A1(n16813), .A2(n16814), .ZN(n16812) );
  INV_X1 U16622 ( .A(n16815), .ZN(n16813) );
  AND2_X1 U16623 ( .A1(n16816), .A2(n16815), .ZN(n16811) );
  INV_X1 U16624 ( .A(n16814), .ZN(n16816) );
  OR2_X1 U16625 ( .A1(n16817), .A2(n16029), .ZN(n16034) );
  AND3_X1 U16626 ( .A1(n16818), .A2(n16819), .A3(n16820), .ZN(n16029) );
  AND2_X1 U16627 ( .A1(n16025), .A2(n16028), .ZN(n16817) );
  OR2_X1 U16628 ( .A1(n16820), .A2(n16821), .ZN(n16028) );
  AND2_X1 U16629 ( .A1(n16819), .A2(n16818), .ZN(n16821) );
  INV_X1 U16630 ( .A(n16822), .ZN(n16820) );
  OR2_X1 U16631 ( .A1(n16823), .A2(n16781), .ZN(n16822) );
  INV_X1 U16632 ( .A(n16824), .ZN(n16781) );
  OR2_X1 U16633 ( .A1(n16825), .A2(n16826), .ZN(n16824) );
  AND2_X1 U16634 ( .A1(n16825), .A2(n16826), .ZN(n16823) );
  OR2_X1 U16635 ( .A1(n16827), .A2(n16828), .ZN(n16826) );
  AND2_X1 U16636 ( .A1(n16829), .A2(n16830), .ZN(n16828) );
  AND2_X1 U16637 ( .A1(n16831), .A2(n16832), .ZN(n16827) );
  OR2_X1 U16638 ( .A1(n16829), .A2(n16830), .ZN(n16832) );
  AND2_X1 U16639 ( .A1(n16833), .A2(n16834), .ZN(n16825) );
  INV_X1 U16640 ( .A(n16835), .ZN(n16834) );
  AND2_X1 U16641 ( .A1(n16836), .A2(n16790), .ZN(n16835) );
  OR2_X1 U16642 ( .A1(n16790), .A2(n16836), .ZN(n16833) );
  OR2_X1 U16643 ( .A1(n16837), .A2(n16838), .ZN(n16836) );
  AND2_X1 U16644 ( .A1(n16839), .A2(n16789), .ZN(n16838) );
  INV_X1 U16645 ( .A(n16788), .ZN(n16839) );
  AND2_X1 U16646 ( .A1(n16840), .A2(n16788), .ZN(n16837) );
  OR2_X1 U16647 ( .A1(n16512), .A2(n15003), .ZN(n16788) );
  INV_X1 U16648 ( .A(n16789), .ZN(n16840) );
  OR2_X1 U16649 ( .A1(n16841), .A2(n16842), .ZN(n16789) );
  AND2_X1 U16650 ( .A1(n16843), .A2(n16844), .ZN(n16842) );
  AND2_X1 U16651 ( .A1(n16845), .A2(n16846), .ZN(n16841) );
  OR2_X1 U16652 ( .A1(n16843), .A2(n16844), .ZN(n16846) );
  AND2_X1 U16653 ( .A1(n16847), .A2(n16848), .ZN(n16790) );
  INV_X1 U16654 ( .A(n16849), .ZN(n16848) );
  AND2_X1 U16655 ( .A1(n16850), .A2(n16804), .ZN(n16849) );
  OR2_X1 U16656 ( .A1(n16804), .A2(n16850), .ZN(n16847) );
  OR2_X1 U16657 ( .A1(n16851), .A2(n16852), .ZN(n16850) );
  AND2_X1 U16658 ( .A1(n16853), .A2(n16803), .ZN(n16852) );
  INV_X1 U16659 ( .A(n16802), .ZN(n16853) );
  AND2_X1 U16660 ( .A1(n16854), .A2(n16802), .ZN(n16851) );
  OR2_X1 U16661 ( .A1(n15842), .A2(n15037), .ZN(n16802) );
  INV_X1 U16662 ( .A(n16803), .ZN(n16854) );
  OR2_X1 U16663 ( .A1(n16855), .A2(n16856), .ZN(n16803) );
  AND2_X1 U16664 ( .A1(n16857), .A2(n16858), .ZN(n16856) );
  AND2_X1 U16665 ( .A1(n16859), .A2(n16860), .ZN(n16855) );
  OR2_X1 U16666 ( .A1(n16857), .A2(n16858), .ZN(n16860) );
  AND2_X1 U16667 ( .A1(n16861), .A2(n16862), .ZN(n16804) );
  INV_X1 U16668 ( .A(n16863), .ZN(n16862) );
  AND2_X1 U16669 ( .A1(n16864), .A2(n16865), .ZN(n16863) );
  OR2_X1 U16670 ( .A1(n16865), .A2(n16864), .ZN(n16861) );
  OR2_X1 U16671 ( .A1(n16866), .A2(n16867), .ZN(n16864) );
  AND2_X1 U16672 ( .A1(n16868), .A2(n16869), .ZN(n16867) );
  INV_X1 U16673 ( .A(n16870), .ZN(n16868) );
  AND2_X1 U16674 ( .A1(n16871), .A2(n16870), .ZN(n16866) );
  INV_X1 U16675 ( .A(n16869), .ZN(n16871) );
  OR2_X1 U16676 ( .A1(n16020), .A2(n16015), .ZN(n16025) );
  AND2_X1 U16677 ( .A1(n16017), .A2(n16019), .ZN(n16015) );
  OR2_X1 U16678 ( .A1(n16872), .A2(n16873), .ZN(n16019) );
  OR2_X1 U16679 ( .A1(n16011), .A2(n16006), .ZN(n16017) );
  AND2_X1 U16680 ( .A1(n16008), .A2(n16009), .ZN(n16006) );
  OR2_X1 U16681 ( .A1(n16874), .A2(n16875), .ZN(n16009) );
  AND2_X1 U16682 ( .A1(n16876), .A2(n16877), .ZN(n16874) );
  OR2_X1 U16683 ( .A1(n16878), .A2(n16001), .ZN(n16008) );
  AND3_X1 U16684 ( .A1(n16879), .A2(n16880), .A3(n16881), .ZN(n16001) );
  AND2_X1 U16685 ( .A1(n15998), .A2(n16002), .ZN(n16878) );
  OR2_X1 U16686 ( .A1(n16882), .A2(n16879), .ZN(n16002) );
  OR2_X1 U16687 ( .A1(n16883), .A2(n16884), .ZN(n16879) );
  AND2_X1 U16688 ( .A1(n16877), .A2(n16885), .ZN(n16884) );
  AND2_X1 U16689 ( .A1(n16886), .A2(n16876), .ZN(n16883) );
  AND3_X1 U16690 ( .A1(n15976), .A2(n15982), .A3(n15977), .ZN(n15998) );
  INV_X1 U16691 ( .A(n15974), .ZN(n15977) );
  OR2_X1 U16692 ( .A1(n16887), .A2(n16888), .ZN(n15974) );
  AND2_X1 U16693 ( .A1(n15967), .A2(n15969), .ZN(n16888) );
  AND2_X1 U16694 ( .A1(n15964), .A2(n16889), .ZN(n16887) );
  OR2_X1 U16695 ( .A1(n15967), .A2(n15969), .ZN(n16889) );
  OR2_X1 U16696 ( .A1(n16890), .A2(n16891), .ZN(n15969) );
  AND2_X1 U16697 ( .A1(n15819), .A2(n15821), .ZN(n16891) );
  AND2_X1 U16698 ( .A1(n15816), .A2(n16892), .ZN(n16890) );
  OR2_X1 U16699 ( .A1(n15819), .A2(n15821), .ZN(n16892) );
  OR2_X1 U16700 ( .A1(n16893), .A2(n16894), .ZN(n15821) );
  AND2_X1 U16701 ( .A1(n15785), .A2(n15787), .ZN(n16894) );
  AND2_X1 U16702 ( .A1(n15782), .A2(n16895), .ZN(n16893) );
  OR2_X1 U16703 ( .A1(n15785), .A2(n15787), .ZN(n16895) );
  OR2_X1 U16704 ( .A1(n16896), .A2(n16897), .ZN(n15787) );
  AND2_X1 U16705 ( .A1(n15751), .A2(n15753), .ZN(n16897) );
  AND2_X1 U16706 ( .A1(n15748), .A2(n16898), .ZN(n16896) );
  OR2_X1 U16707 ( .A1(n15751), .A2(n15753), .ZN(n16898) );
  OR2_X1 U16708 ( .A1(n16899), .A2(n16900), .ZN(n15753) );
  AND2_X1 U16709 ( .A1(n15717), .A2(n15719), .ZN(n16900) );
  AND2_X1 U16710 ( .A1(n15714), .A2(n16901), .ZN(n16899) );
  OR2_X1 U16711 ( .A1(n15717), .A2(n15719), .ZN(n16901) );
  OR2_X1 U16712 ( .A1(n16902), .A2(n16903), .ZN(n15719) );
  AND2_X1 U16713 ( .A1(n15683), .A2(n15685), .ZN(n16903) );
  AND2_X1 U16714 ( .A1(n15680), .A2(n16904), .ZN(n16902) );
  OR2_X1 U16715 ( .A1(n15683), .A2(n15685), .ZN(n16904) );
  OR2_X1 U16716 ( .A1(n16905), .A2(n16906), .ZN(n15685) );
  AND2_X1 U16717 ( .A1(n15649), .A2(n15651), .ZN(n16906) );
  AND2_X1 U16718 ( .A1(n15646), .A2(n16907), .ZN(n16905) );
  OR2_X1 U16719 ( .A1(n15649), .A2(n15651), .ZN(n16907) );
  OR2_X1 U16720 ( .A1(n16908), .A2(n16909), .ZN(n15651) );
  AND2_X1 U16721 ( .A1(n15615), .A2(n15617), .ZN(n16909) );
  AND2_X1 U16722 ( .A1(n15612), .A2(n16910), .ZN(n16908) );
  OR2_X1 U16723 ( .A1(n15615), .A2(n15617), .ZN(n16910) );
  OR2_X1 U16724 ( .A1(n16911), .A2(n16912), .ZN(n15617) );
  AND2_X1 U16725 ( .A1(n15570), .A2(n15572), .ZN(n16912) );
  AND2_X1 U16726 ( .A1(n15567), .A2(n16913), .ZN(n16911) );
  OR2_X1 U16727 ( .A1(n15570), .A2(n15572), .ZN(n16913) );
  OR2_X1 U16728 ( .A1(n16914), .A2(n16915), .ZN(n15572) );
  AND2_X1 U16729 ( .A1(n15536), .A2(n15538), .ZN(n16915) );
  AND2_X1 U16730 ( .A1(n15533), .A2(n16916), .ZN(n16914) );
  OR2_X1 U16731 ( .A1(n15536), .A2(n15538), .ZN(n16916) );
  OR2_X1 U16732 ( .A1(n16917), .A2(n16918), .ZN(n15538) );
  AND2_X1 U16733 ( .A1(n15502), .A2(n15504), .ZN(n16918) );
  AND2_X1 U16734 ( .A1(n15499), .A2(n16919), .ZN(n16917) );
  OR2_X1 U16735 ( .A1(n15502), .A2(n15504), .ZN(n16919) );
  OR2_X1 U16736 ( .A1(n16920), .A2(n16921), .ZN(n15504) );
  AND2_X1 U16737 ( .A1(n15468), .A2(n15470), .ZN(n16921) );
  AND2_X1 U16738 ( .A1(n15465), .A2(n16922), .ZN(n16920) );
  OR2_X1 U16739 ( .A1(n15468), .A2(n15470), .ZN(n16922) );
  OR2_X1 U16740 ( .A1(n16923), .A2(n16924), .ZN(n15470) );
  AND2_X1 U16741 ( .A1(n15434), .A2(n15436), .ZN(n16924) );
  AND2_X1 U16742 ( .A1(n15431), .A2(n16925), .ZN(n16923) );
  OR2_X1 U16743 ( .A1(n15434), .A2(n15436), .ZN(n16925) );
  OR2_X1 U16744 ( .A1(n16926), .A2(n16927), .ZN(n15436) );
  AND2_X1 U16745 ( .A1(n15400), .A2(n15402), .ZN(n16927) );
  AND2_X1 U16746 ( .A1(n15397), .A2(n16928), .ZN(n16926) );
  OR2_X1 U16747 ( .A1(n15400), .A2(n15402), .ZN(n16928) );
  OR2_X1 U16748 ( .A1(n16929), .A2(n16930), .ZN(n15402) );
  AND2_X1 U16749 ( .A1(n15366), .A2(n15368), .ZN(n16930) );
  AND2_X1 U16750 ( .A1(n15363), .A2(n16931), .ZN(n16929) );
  OR2_X1 U16751 ( .A1(n15366), .A2(n15368), .ZN(n16931) );
  OR2_X1 U16752 ( .A1(n16932), .A2(n16933), .ZN(n15368) );
  AND2_X1 U16753 ( .A1(n15332), .A2(n15334), .ZN(n16933) );
  AND2_X1 U16754 ( .A1(n15329), .A2(n16934), .ZN(n16932) );
  OR2_X1 U16755 ( .A1(n15332), .A2(n15334), .ZN(n16934) );
  OR2_X1 U16756 ( .A1(n16935), .A2(n16936), .ZN(n15334) );
  AND2_X1 U16757 ( .A1(n15298), .A2(n15300), .ZN(n16936) );
  AND2_X1 U16758 ( .A1(n15295), .A2(n16937), .ZN(n16935) );
  OR2_X1 U16759 ( .A1(n15298), .A2(n15300), .ZN(n16937) );
  OR2_X1 U16760 ( .A1(n16938), .A2(n16939), .ZN(n15300) );
  AND2_X1 U16761 ( .A1(n15264), .A2(n15266), .ZN(n16939) );
  AND2_X1 U16762 ( .A1(n15261), .A2(n16940), .ZN(n16938) );
  OR2_X1 U16763 ( .A1(n15264), .A2(n15266), .ZN(n16940) );
  OR2_X1 U16764 ( .A1(n16941), .A2(n16942), .ZN(n15266) );
  AND2_X1 U16765 ( .A1(n15219), .A2(n15221), .ZN(n16942) );
  AND2_X1 U16766 ( .A1(n15216), .A2(n16943), .ZN(n16941) );
  OR2_X1 U16767 ( .A1(n15219), .A2(n15221), .ZN(n16943) );
  OR2_X1 U16768 ( .A1(n16944), .A2(n16945), .ZN(n15221) );
  AND2_X1 U16769 ( .A1(n15185), .A2(n15187), .ZN(n16945) );
  AND2_X1 U16770 ( .A1(n15182), .A2(n16946), .ZN(n16944) );
  OR2_X1 U16771 ( .A1(n15185), .A2(n15187), .ZN(n16946) );
  OR2_X1 U16772 ( .A1(n16947), .A2(n16948), .ZN(n15187) );
  AND2_X1 U16773 ( .A1(n15151), .A2(n15153), .ZN(n16948) );
  AND2_X1 U16774 ( .A1(n15148), .A2(n16949), .ZN(n16947) );
  OR2_X1 U16775 ( .A1(n15151), .A2(n15153), .ZN(n16949) );
  OR2_X1 U16776 ( .A1(n16950), .A2(n16951), .ZN(n15153) );
  AND2_X1 U16777 ( .A1(n15117), .A2(n15119), .ZN(n16951) );
  AND2_X1 U16778 ( .A1(n15114), .A2(n16952), .ZN(n16950) );
  OR2_X1 U16779 ( .A1(n15117), .A2(n15119), .ZN(n16952) );
  OR2_X1 U16780 ( .A1(n16953), .A2(n16954), .ZN(n15119) );
  AND2_X1 U16781 ( .A1(n15083), .A2(n15085), .ZN(n16954) );
  AND2_X1 U16782 ( .A1(n15080), .A2(n16955), .ZN(n16953) );
  OR2_X1 U16783 ( .A1(n15083), .A2(n15085), .ZN(n16955) );
  OR2_X1 U16784 ( .A1(n16956), .A2(n16957), .ZN(n15085) );
  AND2_X1 U16785 ( .A1(n15049), .A2(n15051), .ZN(n16957) );
  AND2_X1 U16786 ( .A1(n15046), .A2(n16958), .ZN(n16956) );
  OR2_X1 U16787 ( .A1(n15049), .A2(n15051), .ZN(n16958) );
  OR2_X1 U16788 ( .A1(n16959), .A2(n16960), .ZN(n15051) );
  AND2_X1 U16789 ( .A1(n15015), .A2(n15017), .ZN(n16960) );
  AND2_X1 U16790 ( .A1(n15012), .A2(n16961), .ZN(n16959) );
  OR2_X1 U16791 ( .A1(n15015), .A2(n15017), .ZN(n16961) );
  OR2_X1 U16792 ( .A1(n16962), .A2(n16963), .ZN(n15017) );
  AND2_X1 U16793 ( .A1(n14981), .A2(n14983), .ZN(n16963) );
  AND2_X1 U16794 ( .A1(n14978), .A2(n16964), .ZN(n16962) );
  OR2_X1 U16795 ( .A1(n14981), .A2(n14983), .ZN(n16964) );
  OR2_X1 U16796 ( .A1(n16965), .A2(n16966), .ZN(n14983) );
  AND2_X1 U16797 ( .A1(n14947), .A2(n14949), .ZN(n16966) );
  AND2_X1 U16798 ( .A1(n14944), .A2(n16967), .ZN(n16965) );
  OR2_X1 U16799 ( .A1(n14947), .A2(n14949), .ZN(n16967) );
  OR2_X1 U16800 ( .A1(n16968), .A2(n16969), .ZN(n14949) );
  AND2_X1 U16801 ( .A1(n14913), .A2(n14915), .ZN(n16969) );
  AND2_X1 U16802 ( .A1(n14910), .A2(n16970), .ZN(n16968) );
  OR2_X1 U16803 ( .A1(n14913), .A2(n14915), .ZN(n16970) );
  OR2_X1 U16804 ( .A1(n16971), .A2(n16972), .ZN(n14915) );
  AND2_X1 U16805 ( .A1(n14868), .A2(n14870), .ZN(n16972) );
  AND2_X1 U16806 ( .A1(n14865), .A2(n16973), .ZN(n16971) );
  OR2_X1 U16807 ( .A1(n14868), .A2(n14870), .ZN(n16973) );
  OR2_X1 U16808 ( .A1(n16974), .A2(n16975), .ZN(n14870) );
  AND2_X1 U16809 ( .A1(n14837), .A2(n14835), .ZN(n16975) );
  AND2_X1 U16810 ( .A1(n14829), .A2(n16976), .ZN(n16974) );
  OR2_X1 U16811 ( .A1(n14837), .A2(n14835), .ZN(n16976) );
  INV_X1 U16812 ( .A(n14836), .ZN(n14835) );
  AND3_X1 U16813 ( .A1(b_31_), .A2(b_30_), .A3(n15957), .ZN(n14836) );
  INV_X1 U16814 ( .A(n14834), .ZN(n14837) );
  AND2_X1 U16815 ( .A1(a_29_), .A2(b_31_), .ZN(n14834) );
  INV_X1 U16816 ( .A(n16977), .ZN(n14829) );
  OR3_X1 U16817 ( .A1(n16978), .A2(n16979), .A3(n16980), .ZN(n16977) );
  AND2_X1 U16818 ( .A1(n16981), .A2(b_30_), .ZN(n16980) );
  AND2_X1 U16819 ( .A1(b_29_), .A2(n16982), .ZN(n16979) );
  OR2_X1 U16820 ( .A1(n16983), .A2(n14817), .ZN(n16982) );
  AND2_X1 U16821 ( .A1(a_31_), .A2(n14801), .ZN(n16983) );
  AND2_X1 U16822 ( .A1(n14818), .A2(n14856), .ZN(n16978) );
  AND2_X1 U16823 ( .A1(a_30_), .A2(b_30_), .ZN(n14818) );
  OR2_X1 U16824 ( .A1(n14891), .A2(n15959), .ZN(n14868) );
  OR2_X1 U16825 ( .A1(n16984), .A2(n16985), .ZN(n14865) );
  AND2_X1 U16826 ( .A1(n16986), .A2(n16987), .ZN(n16985) );
  INV_X1 U16827 ( .A(n16988), .ZN(n16984) );
  OR2_X1 U16828 ( .A1(n16986), .A2(n16987), .ZN(n16988) );
  OR2_X1 U16829 ( .A1(n16989), .A2(n16990), .ZN(n16986) );
  AND2_X1 U16830 ( .A1(n16991), .A2(n16992), .ZN(n16990) );
  AND2_X1 U16831 ( .A1(n16993), .A2(n16994), .ZN(n16989) );
  OR2_X1 U16832 ( .A1(n14936), .A2(n15959), .ZN(n14913) );
  OR2_X1 U16833 ( .A1(n16995), .A2(n16996), .ZN(n14910) );
  INV_X1 U16834 ( .A(n16997), .ZN(n16996) );
  OR2_X1 U16835 ( .A1(n16998), .A2(n16999), .ZN(n16997) );
  AND2_X1 U16836 ( .A1(n16999), .A2(n16998), .ZN(n16995) );
  AND2_X1 U16837 ( .A1(n17000), .A2(n17001), .ZN(n16998) );
  OR2_X1 U16838 ( .A1(n17002), .A2(n17003), .ZN(n17001) );
  INV_X1 U16839 ( .A(n17004), .ZN(n17003) );
  OR2_X1 U16840 ( .A1(n17004), .A2(n17005), .ZN(n17000) );
  INV_X1 U16841 ( .A(n17002), .ZN(n17005) );
  OR2_X1 U16842 ( .A1(n14970), .A2(n15959), .ZN(n14947) );
  OR2_X1 U16843 ( .A1(n17006), .A2(n17007), .ZN(n14944) );
  INV_X1 U16844 ( .A(n17008), .ZN(n17007) );
  OR2_X1 U16845 ( .A1(n17009), .A2(n17010), .ZN(n17008) );
  AND2_X1 U16846 ( .A1(n17010), .A2(n17009), .ZN(n17006) );
  AND2_X1 U16847 ( .A1(n17011), .A2(n17012), .ZN(n17009) );
  OR2_X1 U16848 ( .A1(n17013), .A2(n17014), .ZN(n17012) );
  INV_X1 U16849 ( .A(n17015), .ZN(n17014) );
  OR2_X1 U16850 ( .A1(n17015), .A2(n17016), .ZN(n17011) );
  INV_X1 U16851 ( .A(n17013), .ZN(n17016) );
  OR2_X1 U16852 ( .A1(n15004), .A2(n15959), .ZN(n14981) );
  OR2_X1 U16853 ( .A1(n17017), .A2(n17018), .ZN(n14978) );
  INV_X1 U16854 ( .A(n17019), .ZN(n17018) );
  OR2_X1 U16855 ( .A1(n17020), .A2(n17021), .ZN(n17019) );
  AND2_X1 U16856 ( .A1(n17021), .A2(n17020), .ZN(n17017) );
  AND2_X1 U16857 ( .A1(n17022), .A2(n17023), .ZN(n17020) );
  OR2_X1 U16858 ( .A1(n17024), .A2(n17025), .ZN(n17023) );
  INV_X1 U16859 ( .A(n17026), .ZN(n17025) );
  OR2_X1 U16860 ( .A1(n17026), .A2(n17027), .ZN(n17022) );
  INV_X1 U16861 ( .A(n17024), .ZN(n17027) );
  OR2_X1 U16862 ( .A1(n15038), .A2(n15959), .ZN(n15015) );
  OR2_X1 U16863 ( .A1(n17028), .A2(n17029), .ZN(n15012) );
  INV_X1 U16864 ( .A(n17030), .ZN(n17029) );
  OR2_X1 U16865 ( .A1(n17031), .A2(n17032), .ZN(n17030) );
  AND2_X1 U16866 ( .A1(n17032), .A2(n17031), .ZN(n17028) );
  AND2_X1 U16867 ( .A1(n17033), .A2(n17034), .ZN(n17031) );
  OR2_X1 U16868 ( .A1(n17035), .A2(n17036), .ZN(n17034) );
  INV_X1 U16869 ( .A(n17037), .ZN(n17036) );
  OR2_X1 U16870 ( .A1(n17037), .A2(n17038), .ZN(n17033) );
  INV_X1 U16871 ( .A(n17035), .ZN(n17038) );
  OR2_X1 U16872 ( .A1(n15072), .A2(n15959), .ZN(n15049) );
  OR2_X1 U16873 ( .A1(n17039), .A2(n17040), .ZN(n15046) );
  INV_X1 U16874 ( .A(n17041), .ZN(n17040) );
  OR2_X1 U16875 ( .A1(n17042), .A2(n17043), .ZN(n17041) );
  AND2_X1 U16876 ( .A1(n17043), .A2(n17042), .ZN(n17039) );
  AND2_X1 U16877 ( .A1(n17044), .A2(n17045), .ZN(n17042) );
  OR2_X1 U16878 ( .A1(n17046), .A2(n17047), .ZN(n17045) );
  INV_X1 U16879 ( .A(n17048), .ZN(n17047) );
  OR2_X1 U16880 ( .A1(n17048), .A2(n17049), .ZN(n17044) );
  INV_X1 U16881 ( .A(n17046), .ZN(n17049) );
  OR2_X1 U16882 ( .A1(n15106), .A2(n15959), .ZN(n15083) );
  OR2_X1 U16883 ( .A1(n17050), .A2(n17051), .ZN(n15080) );
  INV_X1 U16884 ( .A(n17052), .ZN(n17051) );
  OR2_X1 U16885 ( .A1(n17053), .A2(n17054), .ZN(n17052) );
  AND2_X1 U16886 ( .A1(n17054), .A2(n17053), .ZN(n17050) );
  AND2_X1 U16887 ( .A1(n17055), .A2(n17056), .ZN(n17053) );
  OR2_X1 U16888 ( .A1(n17057), .A2(n17058), .ZN(n17056) );
  INV_X1 U16889 ( .A(n17059), .ZN(n17058) );
  OR2_X1 U16890 ( .A1(n17059), .A2(n17060), .ZN(n17055) );
  INV_X1 U16891 ( .A(n17057), .ZN(n17060) );
  OR2_X1 U16892 ( .A1(n15140), .A2(n15959), .ZN(n15117) );
  OR2_X1 U16893 ( .A1(n17061), .A2(n17062), .ZN(n15114) );
  INV_X1 U16894 ( .A(n17063), .ZN(n17062) );
  OR2_X1 U16895 ( .A1(n17064), .A2(n17065), .ZN(n17063) );
  AND2_X1 U16896 ( .A1(n17065), .A2(n17064), .ZN(n17061) );
  AND2_X1 U16897 ( .A1(n17066), .A2(n17067), .ZN(n17064) );
  OR2_X1 U16898 ( .A1(n17068), .A2(n17069), .ZN(n17067) );
  INV_X1 U16899 ( .A(n17070), .ZN(n17069) );
  OR2_X1 U16900 ( .A1(n17070), .A2(n17071), .ZN(n17066) );
  INV_X1 U16901 ( .A(n17068), .ZN(n17071) );
  OR2_X1 U16902 ( .A1(n15174), .A2(n15959), .ZN(n15151) );
  OR2_X1 U16903 ( .A1(n17072), .A2(n17073), .ZN(n15148) );
  INV_X1 U16904 ( .A(n17074), .ZN(n17073) );
  OR2_X1 U16905 ( .A1(n17075), .A2(n17076), .ZN(n17074) );
  AND2_X1 U16906 ( .A1(n17076), .A2(n17075), .ZN(n17072) );
  AND2_X1 U16907 ( .A1(n17077), .A2(n17078), .ZN(n17075) );
  OR2_X1 U16908 ( .A1(n17079), .A2(n17080), .ZN(n17078) );
  INV_X1 U16909 ( .A(n17081), .ZN(n17080) );
  OR2_X1 U16910 ( .A1(n17081), .A2(n17082), .ZN(n17077) );
  INV_X1 U16911 ( .A(n17079), .ZN(n17082) );
  OR2_X1 U16912 ( .A1(n15208), .A2(n15959), .ZN(n15185) );
  OR2_X1 U16913 ( .A1(n17083), .A2(n17084), .ZN(n15182) );
  INV_X1 U16914 ( .A(n17085), .ZN(n17084) );
  OR2_X1 U16915 ( .A1(n17086), .A2(n17087), .ZN(n17085) );
  AND2_X1 U16916 ( .A1(n17087), .A2(n17086), .ZN(n17083) );
  AND2_X1 U16917 ( .A1(n17088), .A2(n17089), .ZN(n17086) );
  OR2_X1 U16918 ( .A1(n17090), .A2(n17091), .ZN(n17089) );
  INV_X1 U16919 ( .A(n17092), .ZN(n17091) );
  OR2_X1 U16920 ( .A1(n17092), .A2(n17093), .ZN(n17088) );
  INV_X1 U16921 ( .A(n17090), .ZN(n17093) );
  OR2_X1 U16922 ( .A1(n15242), .A2(n15959), .ZN(n15219) );
  OR2_X1 U16923 ( .A1(n17094), .A2(n17095), .ZN(n15216) );
  INV_X1 U16924 ( .A(n17096), .ZN(n17095) );
  OR2_X1 U16925 ( .A1(n17097), .A2(n17098), .ZN(n17096) );
  AND2_X1 U16926 ( .A1(n17098), .A2(n17097), .ZN(n17094) );
  AND2_X1 U16927 ( .A1(n17099), .A2(n17100), .ZN(n17097) );
  OR2_X1 U16928 ( .A1(n17101), .A2(n17102), .ZN(n17100) );
  INV_X1 U16929 ( .A(n17103), .ZN(n17102) );
  OR2_X1 U16930 ( .A1(n17103), .A2(n17104), .ZN(n17099) );
  INV_X1 U16931 ( .A(n17101), .ZN(n17104) );
  OR2_X1 U16932 ( .A1(n15287), .A2(n15959), .ZN(n15264) );
  OR2_X1 U16933 ( .A1(n17105), .A2(n17106), .ZN(n15261) );
  INV_X1 U16934 ( .A(n17107), .ZN(n17106) );
  OR2_X1 U16935 ( .A1(n17108), .A2(n17109), .ZN(n17107) );
  AND2_X1 U16936 ( .A1(n17109), .A2(n17108), .ZN(n17105) );
  AND2_X1 U16937 ( .A1(n17110), .A2(n17111), .ZN(n17108) );
  OR2_X1 U16938 ( .A1(n17112), .A2(n17113), .ZN(n17111) );
  INV_X1 U16939 ( .A(n17114), .ZN(n17113) );
  OR2_X1 U16940 ( .A1(n17114), .A2(n17115), .ZN(n17110) );
  INV_X1 U16941 ( .A(n17112), .ZN(n17115) );
  OR2_X1 U16942 ( .A1(n15321), .A2(n15959), .ZN(n15298) );
  OR2_X1 U16943 ( .A1(n17116), .A2(n17117), .ZN(n15295) );
  INV_X1 U16944 ( .A(n17118), .ZN(n17117) );
  OR2_X1 U16945 ( .A1(n17119), .A2(n17120), .ZN(n17118) );
  AND2_X1 U16946 ( .A1(n17120), .A2(n17119), .ZN(n17116) );
  AND2_X1 U16947 ( .A1(n17121), .A2(n17122), .ZN(n17119) );
  OR2_X1 U16948 ( .A1(n17123), .A2(n17124), .ZN(n17122) );
  INV_X1 U16949 ( .A(n17125), .ZN(n17124) );
  OR2_X1 U16950 ( .A1(n17125), .A2(n17126), .ZN(n17121) );
  INV_X1 U16951 ( .A(n17123), .ZN(n17126) );
  OR2_X1 U16952 ( .A1(n15355), .A2(n15959), .ZN(n15332) );
  OR2_X1 U16953 ( .A1(n17127), .A2(n17128), .ZN(n15329) );
  INV_X1 U16954 ( .A(n17129), .ZN(n17128) );
  OR2_X1 U16955 ( .A1(n17130), .A2(n17131), .ZN(n17129) );
  AND2_X1 U16956 ( .A1(n17131), .A2(n17130), .ZN(n17127) );
  AND2_X1 U16957 ( .A1(n17132), .A2(n17133), .ZN(n17130) );
  OR2_X1 U16958 ( .A1(n17134), .A2(n17135), .ZN(n17133) );
  INV_X1 U16959 ( .A(n17136), .ZN(n17135) );
  OR2_X1 U16960 ( .A1(n17136), .A2(n17137), .ZN(n17132) );
  INV_X1 U16961 ( .A(n17134), .ZN(n17137) );
  OR2_X1 U16962 ( .A1(n15389), .A2(n15959), .ZN(n15366) );
  OR2_X1 U16963 ( .A1(n17138), .A2(n17139), .ZN(n15363) );
  INV_X1 U16964 ( .A(n17140), .ZN(n17139) );
  OR2_X1 U16965 ( .A1(n17141), .A2(n17142), .ZN(n17140) );
  AND2_X1 U16966 ( .A1(n17142), .A2(n17141), .ZN(n17138) );
  AND2_X1 U16967 ( .A1(n17143), .A2(n17144), .ZN(n17141) );
  OR2_X1 U16968 ( .A1(n17145), .A2(n17146), .ZN(n17144) );
  INV_X1 U16969 ( .A(n17147), .ZN(n17146) );
  OR2_X1 U16970 ( .A1(n17147), .A2(n17148), .ZN(n17143) );
  INV_X1 U16971 ( .A(n17145), .ZN(n17148) );
  OR2_X1 U16972 ( .A1(n15423), .A2(n15959), .ZN(n15400) );
  OR2_X1 U16973 ( .A1(n17149), .A2(n17150), .ZN(n15397) );
  INV_X1 U16974 ( .A(n17151), .ZN(n17150) );
  OR2_X1 U16975 ( .A1(n17152), .A2(n17153), .ZN(n17151) );
  AND2_X1 U16976 ( .A1(n17153), .A2(n17152), .ZN(n17149) );
  AND2_X1 U16977 ( .A1(n17154), .A2(n17155), .ZN(n17152) );
  OR2_X1 U16978 ( .A1(n17156), .A2(n17157), .ZN(n17155) );
  INV_X1 U16979 ( .A(n17158), .ZN(n17157) );
  OR2_X1 U16980 ( .A1(n17158), .A2(n17159), .ZN(n17154) );
  INV_X1 U16981 ( .A(n17156), .ZN(n17159) );
  OR2_X1 U16982 ( .A1(n15457), .A2(n15959), .ZN(n15434) );
  OR2_X1 U16983 ( .A1(n17160), .A2(n17161), .ZN(n15431) );
  INV_X1 U16984 ( .A(n17162), .ZN(n17161) );
  OR2_X1 U16985 ( .A1(n17163), .A2(n17164), .ZN(n17162) );
  AND2_X1 U16986 ( .A1(n17164), .A2(n17163), .ZN(n17160) );
  AND2_X1 U16987 ( .A1(n17165), .A2(n17166), .ZN(n17163) );
  OR2_X1 U16988 ( .A1(n17167), .A2(n17168), .ZN(n17166) );
  INV_X1 U16989 ( .A(n17169), .ZN(n17168) );
  OR2_X1 U16990 ( .A1(n17169), .A2(n17170), .ZN(n17165) );
  INV_X1 U16991 ( .A(n17167), .ZN(n17170) );
  OR2_X1 U16992 ( .A1(n15491), .A2(n15959), .ZN(n15468) );
  OR2_X1 U16993 ( .A1(n17171), .A2(n17172), .ZN(n15465) );
  INV_X1 U16994 ( .A(n17173), .ZN(n17172) );
  OR2_X1 U16995 ( .A1(n17174), .A2(n17175), .ZN(n17173) );
  AND2_X1 U16996 ( .A1(n17175), .A2(n17174), .ZN(n17171) );
  AND2_X1 U16997 ( .A1(n17176), .A2(n17177), .ZN(n17174) );
  OR2_X1 U16998 ( .A1(n17178), .A2(n17179), .ZN(n17177) );
  INV_X1 U16999 ( .A(n17180), .ZN(n17179) );
  OR2_X1 U17000 ( .A1(n17180), .A2(n17181), .ZN(n17176) );
  INV_X1 U17001 ( .A(n17178), .ZN(n17181) );
  OR2_X1 U17002 ( .A1(n15525), .A2(n15959), .ZN(n15502) );
  OR2_X1 U17003 ( .A1(n17182), .A2(n17183), .ZN(n15499) );
  INV_X1 U17004 ( .A(n17184), .ZN(n17183) );
  OR2_X1 U17005 ( .A1(n17185), .A2(n17186), .ZN(n17184) );
  AND2_X1 U17006 ( .A1(n17186), .A2(n17185), .ZN(n17182) );
  AND2_X1 U17007 ( .A1(n17187), .A2(n17188), .ZN(n17185) );
  OR2_X1 U17008 ( .A1(n17189), .A2(n17190), .ZN(n17188) );
  INV_X1 U17009 ( .A(n17191), .ZN(n17190) );
  OR2_X1 U17010 ( .A1(n17191), .A2(n17192), .ZN(n17187) );
  INV_X1 U17011 ( .A(n17189), .ZN(n17192) );
  OR2_X1 U17012 ( .A1(n15559), .A2(n15959), .ZN(n15536) );
  OR2_X1 U17013 ( .A1(n17193), .A2(n17194), .ZN(n15533) );
  INV_X1 U17014 ( .A(n17195), .ZN(n17194) );
  OR2_X1 U17015 ( .A1(n17196), .A2(n17197), .ZN(n17195) );
  AND2_X1 U17016 ( .A1(n17197), .A2(n17196), .ZN(n17193) );
  AND2_X1 U17017 ( .A1(n17198), .A2(n17199), .ZN(n17196) );
  OR2_X1 U17018 ( .A1(n17200), .A2(n17201), .ZN(n17199) );
  INV_X1 U17019 ( .A(n17202), .ZN(n17201) );
  OR2_X1 U17020 ( .A1(n17202), .A2(n17203), .ZN(n17198) );
  INV_X1 U17021 ( .A(n17200), .ZN(n17203) );
  OR2_X1 U17022 ( .A1(n15593), .A2(n15959), .ZN(n15570) );
  OR2_X1 U17023 ( .A1(n17204), .A2(n17205), .ZN(n15567) );
  INV_X1 U17024 ( .A(n17206), .ZN(n17205) );
  OR2_X1 U17025 ( .A1(n17207), .A2(n17208), .ZN(n17206) );
  AND2_X1 U17026 ( .A1(n17208), .A2(n17207), .ZN(n17204) );
  AND2_X1 U17027 ( .A1(n17209), .A2(n17210), .ZN(n17207) );
  OR2_X1 U17028 ( .A1(n17211), .A2(n17212), .ZN(n17210) );
  INV_X1 U17029 ( .A(n17213), .ZN(n17212) );
  OR2_X1 U17030 ( .A1(n17213), .A2(n17214), .ZN(n17209) );
  INV_X1 U17031 ( .A(n17211), .ZN(n17214) );
  OR2_X1 U17032 ( .A1(n15638), .A2(n15959), .ZN(n15615) );
  OR2_X1 U17033 ( .A1(n17215), .A2(n17216), .ZN(n15612) );
  INV_X1 U17034 ( .A(n17217), .ZN(n17216) );
  OR2_X1 U17035 ( .A1(n17218), .A2(n17219), .ZN(n17217) );
  AND2_X1 U17036 ( .A1(n17219), .A2(n17218), .ZN(n17215) );
  AND2_X1 U17037 ( .A1(n17220), .A2(n17221), .ZN(n17218) );
  OR2_X1 U17038 ( .A1(n17222), .A2(n17223), .ZN(n17221) );
  INV_X1 U17039 ( .A(n17224), .ZN(n17223) );
  OR2_X1 U17040 ( .A1(n17224), .A2(n17225), .ZN(n17220) );
  INV_X1 U17041 ( .A(n17222), .ZN(n17225) );
  OR2_X1 U17042 ( .A1(n15672), .A2(n15959), .ZN(n15649) );
  OR2_X1 U17043 ( .A1(n17226), .A2(n17227), .ZN(n15646) );
  INV_X1 U17044 ( .A(n17228), .ZN(n17227) );
  OR2_X1 U17045 ( .A1(n17229), .A2(n17230), .ZN(n17228) );
  AND2_X1 U17046 ( .A1(n17230), .A2(n17229), .ZN(n17226) );
  AND2_X1 U17047 ( .A1(n17231), .A2(n17232), .ZN(n17229) );
  OR2_X1 U17048 ( .A1(n17233), .A2(n17234), .ZN(n17232) );
  INV_X1 U17049 ( .A(n17235), .ZN(n17234) );
  OR2_X1 U17050 ( .A1(n17235), .A2(n17236), .ZN(n17231) );
  INV_X1 U17051 ( .A(n17233), .ZN(n17236) );
  OR2_X1 U17052 ( .A1(n15706), .A2(n15959), .ZN(n15683) );
  OR2_X1 U17053 ( .A1(n17237), .A2(n17238), .ZN(n15680) );
  INV_X1 U17054 ( .A(n17239), .ZN(n17238) );
  OR2_X1 U17055 ( .A1(n17240), .A2(n17241), .ZN(n17239) );
  AND2_X1 U17056 ( .A1(n17241), .A2(n17240), .ZN(n17237) );
  AND2_X1 U17057 ( .A1(n17242), .A2(n17243), .ZN(n17240) );
  OR2_X1 U17058 ( .A1(n17244), .A2(n17245), .ZN(n17243) );
  INV_X1 U17059 ( .A(n17246), .ZN(n17245) );
  OR2_X1 U17060 ( .A1(n17246), .A2(n17247), .ZN(n17242) );
  INV_X1 U17061 ( .A(n17244), .ZN(n17247) );
  OR2_X1 U17062 ( .A1(n15740), .A2(n15959), .ZN(n15717) );
  OR2_X1 U17063 ( .A1(n17248), .A2(n17249), .ZN(n15714) );
  INV_X1 U17064 ( .A(n17250), .ZN(n17249) );
  OR2_X1 U17065 ( .A1(n17251), .A2(n17252), .ZN(n17250) );
  AND2_X1 U17066 ( .A1(n17252), .A2(n17251), .ZN(n17248) );
  AND2_X1 U17067 ( .A1(n17253), .A2(n17254), .ZN(n17251) );
  OR2_X1 U17068 ( .A1(n17255), .A2(n17256), .ZN(n17254) );
  INV_X1 U17069 ( .A(n17257), .ZN(n17256) );
  OR2_X1 U17070 ( .A1(n17257), .A2(n17258), .ZN(n17253) );
  INV_X1 U17071 ( .A(n17255), .ZN(n17258) );
  OR2_X1 U17072 ( .A1(n15774), .A2(n15959), .ZN(n15751) );
  OR2_X1 U17073 ( .A1(n17259), .A2(n17260), .ZN(n15748) );
  INV_X1 U17074 ( .A(n17261), .ZN(n17260) );
  OR2_X1 U17075 ( .A1(n17262), .A2(n17263), .ZN(n17261) );
  AND2_X1 U17076 ( .A1(n17263), .A2(n17262), .ZN(n17259) );
  AND2_X1 U17077 ( .A1(n17264), .A2(n17265), .ZN(n17262) );
  OR2_X1 U17078 ( .A1(n17266), .A2(n17267), .ZN(n17265) );
  INV_X1 U17079 ( .A(n17268), .ZN(n17267) );
  OR2_X1 U17080 ( .A1(n17268), .A2(n17269), .ZN(n17264) );
  INV_X1 U17081 ( .A(n17266), .ZN(n17269) );
  OR2_X1 U17082 ( .A1(n15808), .A2(n15959), .ZN(n15785) );
  OR2_X1 U17083 ( .A1(n17270), .A2(n17271), .ZN(n15782) );
  INV_X1 U17084 ( .A(n17272), .ZN(n17271) );
  OR2_X1 U17085 ( .A1(n17273), .A2(n17274), .ZN(n17272) );
  AND2_X1 U17086 ( .A1(n17274), .A2(n17273), .ZN(n17270) );
  AND2_X1 U17087 ( .A1(n17275), .A2(n17276), .ZN(n17273) );
  OR2_X1 U17088 ( .A1(n17277), .A2(n17278), .ZN(n17276) );
  INV_X1 U17089 ( .A(n17279), .ZN(n17278) );
  OR2_X1 U17090 ( .A1(n17279), .A2(n17280), .ZN(n17275) );
  INV_X1 U17091 ( .A(n17277), .ZN(n17280) );
  OR2_X1 U17092 ( .A1(n15842), .A2(n15959), .ZN(n15819) );
  OR2_X1 U17093 ( .A1(n17281), .A2(n17282), .ZN(n15816) );
  INV_X1 U17094 ( .A(n17283), .ZN(n17282) );
  OR2_X1 U17095 ( .A1(n17284), .A2(n17285), .ZN(n17283) );
  AND2_X1 U17096 ( .A1(n17285), .A2(n17284), .ZN(n17281) );
  AND2_X1 U17097 ( .A1(n17286), .A2(n17287), .ZN(n17284) );
  OR2_X1 U17098 ( .A1(n17288), .A2(n17289), .ZN(n17287) );
  INV_X1 U17099 ( .A(n17290), .ZN(n17289) );
  OR2_X1 U17100 ( .A1(n17290), .A2(n17291), .ZN(n17286) );
  INV_X1 U17101 ( .A(n17288), .ZN(n17291) );
  OR2_X1 U17102 ( .A1(n16512), .A2(n15959), .ZN(n15967) );
  INV_X1 U17103 ( .A(b_31_), .ZN(n15959) );
  OR2_X1 U17104 ( .A1(n17292), .A2(n17293), .ZN(n15964) );
  INV_X1 U17105 ( .A(n17294), .ZN(n17293) );
  OR2_X1 U17106 ( .A1(n17295), .A2(n17296), .ZN(n17294) );
  AND2_X1 U17107 ( .A1(n17296), .A2(n17295), .ZN(n17292) );
  AND2_X1 U17108 ( .A1(n17297), .A2(n17298), .ZN(n17295) );
  OR2_X1 U17109 ( .A1(n17299), .A2(n17300), .ZN(n17298) );
  INV_X1 U17110 ( .A(n17301), .ZN(n17300) );
  OR2_X1 U17111 ( .A1(n17301), .A2(n17302), .ZN(n17297) );
  INV_X1 U17112 ( .A(n17299), .ZN(n17302) );
  INV_X1 U17113 ( .A(n17303), .ZN(n15982) );
  OR2_X1 U17114 ( .A1(n16882), .A2(n17304), .ZN(n17303) );
  AND2_X1 U17115 ( .A1(n17305), .A2(n17306), .ZN(n17304) );
  AND2_X1 U17116 ( .A1(n16881), .A2(n16880), .ZN(n16882) );
  INV_X1 U17117 ( .A(n17305), .ZN(n16880) );
  OR2_X1 U17118 ( .A1(n17307), .A2(n17308), .ZN(n17305) );
  AND3_X1 U17119 ( .A1(n17309), .A2(n17310), .A3(n17311), .ZN(n17308) );
  OR2_X1 U17120 ( .A1(n17312), .A2(n17313), .ZN(n17310) );
  OR2_X1 U17121 ( .A1(n17314), .A2(n17315), .ZN(n17309) );
  AND2_X1 U17122 ( .A1(n17316), .A2(n17317), .ZN(n17307) );
  OR2_X1 U17123 ( .A1(n17318), .A2(n17319), .ZN(n17316) );
  AND2_X1 U17124 ( .A1(n17312), .A2(n17313), .ZN(n17319) );
  INV_X1 U17125 ( .A(n17315), .ZN(n17312) );
  AND2_X1 U17126 ( .A1(n17314), .A2(n17315), .ZN(n17318) );
  INV_X1 U17127 ( .A(n17313), .ZN(n17314) );
  INV_X1 U17128 ( .A(n17306), .ZN(n16881) );
  OR2_X1 U17129 ( .A1(n17320), .A2(n17321), .ZN(n17306) );
  AND2_X1 U17130 ( .A1(n17322), .A2(n17323), .ZN(n17321) );
  AND2_X1 U17131 ( .A1(n17324), .A2(n17325), .ZN(n17320) );
  OR2_X1 U17132 ( .A1(n17322), .A2(n17323), .ZN(n17325) );
  AND2_X1 U17133 ( .A1(n17326), .A2(n17327), .ZN(n15976) );
  OR2_X1 U17134 ( .A1(n17328), .A2(n17324), .ZN(n17327) );
  INV_X1 U17135 ( .A(n17329), .ZN(n17326) );
  AND2_X1 U17136 ( .A1(n17324), .A2(n17328), .ZN(n17329) );
  AND2_X1 U17137 ( .A1(n17330), .A2(n17331), .ZN(n17328) );
  OR2_X1 U17138 ( .A1(n17322), .A2(n17332), .ZN(n17331) );
  INV_X1 U17139 ( .A(n17323), .ZN(n17332) );
  OR2_X1 U17140 ( .A1(n17323), .A2(n17333), .ZN(n17330) );
  INV_X1 U17141 ( .A(n17322), .ZN(n17333) );
  OR2_X1 U17142 ( .A1(n16512), .A2(n14801), .ZN(n17322) );
  OR2_X1 U17143 ( .A1(n17334), .A2(n17335), .ZN(n17323) );
  AND2_X1 U17144 ( .A1(n17296), .A2(n17299), .ZN(n17335) );
  AND2_X1 U17145 ( .A1(n17336), .A2(n17301), .ZN(n17334) );
  OR2_X1 U17146 ( .A1(n17337), .A2(n17338), .ZN(n17301) );
  AND2_X1 U17147 ( .A1(n17285), .A2(n17288), .ZN(n17338) );
  AND2_X1 U17148 ( .A1(n17339), .A2(n17290), .ZN(n17337) );
  OR2_X1 U17149 ( .A1(n17340), .A2(n17341), .ZN(n17290) );
  AND2_X1 U17150 ( .A1(n17274), .A2(n17277), .ZN(n17341) );
  AND2_X1 U17151 ( .A1(n17342), .A2(n17279), .ZN(n17340) );
  OR2_X1 U17152 ( .A1(n17343), .A2(n17344), .ZN(n17279) );
  AND2_X1 U17153 ( .A1(n17263), .A2(n17266), .ZN(n17344) );
  AND2_X1 U17154 ( .A1(n17345), .A2(n17268), .ZN(n17343) );
  OR2_X1 U17155 ( .A1(n17346), .A2(n17347), .ZN(n17268) );
  AND2_X1 U17156 ( .A1(n17252), .A2(n17255), .ZN(n17347) );
  AND2_X1 U17157 ( .A1(n17348), .A2(n17257), .ZN(n17346) );
  OR2_X1 U17158 ( .A1(n17349), .A2(n17350), .ZN(n17257) );
  AND2_X1 U17159 ( .A1(n17241), .A2(n17244), .ZN(n17350) );
  AND2_X1 U17160 ( .A1(n17351), .A2(n17246), .ZN(n17349) );
  OR2_X1 U17161 ( .A1(n17352), .A2(n17353), .ZN(n17246) );
  AND2_X1 U17162 ( .A1(n17230), .A2(n17233), .ZN(n17353) );
  AND2_X1 U17163 ( .A1(n17354), .A2(n17235), .ZN(n17352) );
  OR2_X1 U17164 ( .A1(n17355), .A2(n17356), .ZN(n17235) );
  AND2_X1 U17165 ( .A1(n17219), .A2(n17222), .ZN(n17356) );
  AND2_X1 U17166 ( .A1(n17357), .A2(n17224), .ZN(n17355) );
  OR2_X1 U17167 ( .A1(n17358), .A2(n17359), .ZN(n17224) );
  AND2_X1 U17168 ( .A1(n17208), .A2(n17211), .ZN(n17359) );
  AND2_X1 U17169 ( .A1(n17360), .A2(n17213), .ZN(n17358) );
  OR2_X1 U17170 ( .A1(n17361), .A2(n17362), .ZN(n17213) );
  AND2_X1 U17171 ( .A1(n17197), .A2(n17200), .ZN(n17362) );
  AND2_X1 U17172 ( .A1(n17363), .A2(n17202), .ZN(n17361) );
  OR2_X1 U17173 ( .A1(n17364), .A2(n17365), .ZN(n17202) );
  AND2_X1 U17174 ( .A1(n17186), .A2(n17189), .ZN(n17365) );
  AND2_X1 U17175 ( .A1(n17366), .A2(n17191), .ZN(n17364) );
  OR2_X1 U17176 ( .A1(n17367), .A2(n17368), .ZN(n17191) );
  AND2_X1 U17177 ( .A1(n17175), .A2(n17178), .ZN(n17368) );
  AND2_X1 U17178 ( .A1(n17369), .A2(n17180), .ZN(n17367) );
  OR2_X1 U17179 ( .A1(n17370), .A2(n17371), .ZN(n17180) );
  AND2_X1 U17180 ( .A1(n17164), .A2(n17167), .ZN(n17371) );
  AND2_X1 U17181 ( .A1(n17372), .A2(n17169), .ZN(n17370) );
  OR2_X1 U17182 ( .A1(n17373), .A2(n17374), .ZN(n17169) );
  AND2_X1 U17183 ( .A1(n17153), .A2(n17156), .ZN(n17374) );
  AND2_X1 U17184 ( .A1(n17375), .A2(n17158), .ZN(n17373) );
  OR2_X1 U17185 ( .A1(n17376), .A2(n17377), .ZN(n17158) );
  AND2_X1 U17186 ( .A1(n17142), .A2(n17145), .ZN(n17377) );
  AND2_X1 U17187 ( .A1(n17378), .A2(n17147), .ZN(n17376) );
  OR2_X1 U17188 ( .A1(n17379), .A2(n17380), .ZN(n17147) );
  AND2_X1 U17189 ( .A1(n17131), .A2(n17134), .ZN(n17380) );
  AND2_X1 U17190 ( .A1(n17381), .A2(n17136), .ZN(n17379) );
  OR2_X1 U17191 ( .A1(n17382), .A2(n17383), .ZN(n17136) );
  AND2_X1 U17192 ( .A1(n17120), .A2(n17123), .ZN(n17383) );
  AND2_X1 U17193 ( .A1(n17384), .A2(n17125), .ZN(n17382) );
  OR2_X1 U17194 ( .A1(n17385), .A2(n17386), .ZN(n17125) );
  AND2_X1 U17195 ( .A1(n17109), .A2(n17112), .ZN(n17386) );
  AND2_X1 U17196 ( .A1(n17387), .A2(n17114), .ZN(n17385) );
  OR2_X1 U17197 ( .A1(n17388), .A2(n17389), .ZN(n17114) );
  AND2_X1 U17198 ( .A1(n17098), .A2(n17101), .ZN(n17389) );
  AND2_X1 U17199 ( .A1(n17390), .A2(n17103), .ZN(n17388) );
  OR2_X1 U17200 ( .A1(n17391), .A2(n17392), .ZN(n17103) );
  AND2_X1 U17201 ( .A1(n17087), .A2(n17090), .ZN(n17392) );
  AND2_X1 U17202 ( .A1(n17393), .A2(n17092), .ZN(n17391) );
  OR2_X1 U17203 ( .A1(n17394), .A2(n17395), .ZN(n17092) );
  AND2_X1 U17204 ( .A1(n17076), .A2(n17079), .ZN(n17395) );
  AND2_X1 U17205 ( .A1(n17396), .A2(n17081), .ZN(n17394) );
  OR2_X1 U17206 ( .A1(n17397), .A2(n17398), .ZN(n17081) );
  AND2_X1 U17207 ( .A1(n17065), .A2(n17068), .ZN(n17398) );
  AND2_X1 U17208 ( .A1(n17399), .A2(n17070), .ZN(n17397) );
  OR2_X1 U17209 ( .A1(n17400), .A2(n17401), .ZN(n17070) );
  AND2_X1 U17210 ( .A1(n17054), .A2(n17057), .ZN(n17401) );
  AND2_X1 U17211 ( .A1(n17402), .A2(n17059), .ZN(n17400) );
  OR2_X1 U17212 ( .A1(n17403), .A2(n17404), .ZN(n17059) );
  AND2_X1 U17213 ( .A1(n17043), .A2(n17046), .ZN(n17404) );
  AND2_X1 U17214 ( .A1(n17405), .A2(n17048), .ZN(n17403) );
  OR2_X1 U17215 ( .A1(n17406), .A2(n17407), .ZN(n17048) );
  AND2_X1 U17216 ( .A1(n17032), .A2(n17035), .ZN(n17407) );
  AND2_X1 U17217 ( .A1(n17408), .A2(n17037), .ZN(n17406) );
  OR2_X1 U17218 ( .A1(n17409), .A2(n17410), .ZN(n17037) );
  AND2_X1 U17219 ( .A1(n17021), .A2(n17024), .ZN(n17410) );
  AND2_X1 U17220 ( .A1(n17411), .A2(n17026), .ZN(n17409) );
  OR2_X1 U17221 ( .A1(n17412), .A2(n17413), .ZN(n17026) );
  AND2_X1 U17222 ( .A1(n17010), .A2(n17013), .ZN(n17413) );
  AND2_X1 U17223 ( .A1(n17414), .A2(n17015), .ZN(n17412) );
  OR2_X1 U17224 ( .A1(n17415), .A2(n17416), .ZN(n17015) );
  AND2_X1 U17225 ( .A1(n16999), .A2(n17002), .ZN(n17416) );
  AND2_X1 U17226 ( .A1(n17417), .A2(n17004), .ZN(n17415) );
  OR2_X1 U17227 ( .A1(n17418), .A2(n17419), .ZN(n17004) );
  AND2_X1 U17228 ( .A1(n16987), .A2(n16992), .ZN(n17419) );
  AND2_X1 U17229 ( .A1(n16991), .A2(n17420), .ZN(n17418) );
  OR2_X1 U17230 ( .A1(n16992), .A2(n16987), .ZN(n17420) );
  OR2_X1 U17231 ( .A1(n14857), .A2(n14801), .ZN(n16987) );
  INV_X1 U17232 ( .A(n16993), .ZN(n16992) );
  AND3_X1 U17233 ( .A1(b_30_), .A2(b_29_), .A3(n15957), .ZN(n16993) );
  INV_X1 U17234 ( .A(n16994), .ZN(n16991) );
  OR2_X1 U17235 ( .A1(n17421), .A2(n17422), .ZN(n16994) );
  AND2_X1 U17236 ( .A1(b_29_), .A2(n17423), .ZN(n17422) );
  OR2_X1 U17237 ( .A1(n17424), .A2(n16981), .ZN(n17423) );
  AND2_X1 U17238 ( .A1(a_30_), .A2(n14890), .ZN(n17424) );
  AND2_X1 U17239 ( .A1(b_28_), .A2(n17425), .ZN(n17421) );
  OR2_X1 U17240 ( .A1(n17426), .A2(n14817), .ZN(n17425) );
  AND2_X1 U17241 ( .A1(a_31_), .A2(n14856), .ZN(n17426) );
  OR2_X1 U17242 ( .A1(n17002), .A2(n16999), .ZN(n17417) );
  OR2_X1 U17243 ( .A1(n17427), .A2(n17428), .ZN(n16999) );
  AND2_X1 U17244 ( .A1(n17429), .A2(n15954), .ZN(n17428) );
  INV_X1 U17245 ( .A(n17430), .ZN(n17427) );
  OR2_X1 U17246 ( .A1(n17429), .A2(n15954), .ZN(n17430) );
  OR2_X1 U17247 ( .A1(n17431), .A2(n17432), .ZN(n17429) );
  AND2_X1 U17248 ( .A1(n17433), .A2(n17434), .ZN(n17432) );
  AND2_X1 U17249 ( .A1(n17435), .A2(n17436), .ZN(n17431) );
  OR2_X1 U17250 ( .A1(n14891), .A2(n14801), .ZN(n17002) );
  OR2_X1 U17251 ( .A1(n17013), .A2(n17010), .ZN(n17414) );
  OR2_X1 U17252 ( .A1(n17437), .A2(n17438), .ZN(n17010) );
  INV_X1 U17253 ( .A(n17439), .ZN(n17438) );
  OR2_X1 U17254 ( .A1(n17440), .A2(n17441), .ZN(n17439) );
  AND2_X1 U17255 ( .A1(n17441), .A2(n17440), .ZN(n17437) );
  AND2_X1 U17256 ( .A1(n17442), .A2(n17443), .ZN(n17440) );
  OR2_X1 U17257 ( .A1(n17444), .A2(n17445), .ZN(n17443) );
  INV_X1 U17258 ( .A(n17446), .ZN(n17445) );
  OR2_X1 U17259 ( .A1(n17446), .A2(n17447), .ZN(n17442) );
  INV_X1 U17260 ( .A(n17444), .ZN(n17447) );
  OR2_X1 U17261 ( .A1(n14936), .A2(n14801), .ZN(n17013) );
  OR2_X1 U17262 ( .A1(n17024), .A2(n17021), .ZN(n17411) );
  OR2_X1 U17263 ( .A1(n17448), .A2(n17449), .ZN(n17021) );
  INV_X1 U17264 ( .A(n17450), .ZN(n17449) );
  OR2_X1 U17265 ( .A1(n17451), .A2(n17452), .ZN(n17450) );
  AND2_X1 U17266 ( .A1(n17452), .A2(n17451), .ZN(n17448) );
  AND2_X1 U17267 ( .A1(n17453), .A2(n17454), .ZN(n17451) );
  OR2_X1 U17268 ( .A1(n17455), .A2(n17456), .ZN(n17454) );
  INV_X1 U17269 ( .A(n17457), .ZN(n17456) );
  OR2_X1 U17270 ( .A1(n17457), .A2(n17458), .ZN(n17453) );
  INV_X1 U17271 ( .A(n17455), .ZN(n17458) );
  OR2_X1 U17272 ( .A1(n14970), .A2(n14801), .ZN(n17024) );
  OR2_X1 U17273 ( .A1(n17035), .A2(n17032), .ZN(n17408) );
  OR2_X1 U17274 ( .A1(n17459), .A2(n17460), .ZN(n17032) );
  INV_X1 U17275 ( .A(n17461), .ZN(n17460) );
  OR2_X1 U17276 ( .A1(n17462), .A2(n17463), .ZN(n17461) );
  AND2_X1 U17277 ( .A1(n17463), .A2(n17462), .ZN(n17459) );
  AND2_X1 U17278 ( .A1(n17464), .A2(n17465), .ZN(n17462) );
  OR2_X1 U17279 ( .A1(n17466), .A2(n17467), .ZN(n17465) );
  INV_X1 U17280 ( .A(n17468), .ZN(n17467) );
  OR2_X1 U17281 ( .A1(n17468), .A2(n17469), .ZN(n17464) );
  INV_X1 U17282 ( .A(n17466), .ZN(n17469) );
  OR2_X1 U17283 ( .A1(n15004), .A2(n14801), .ZN(n17035) );
  OR2_X1 U17284 ( .A1(n17046), .A2(n17043), .ZN(n17405) );
  OR2_X1 U17285 ( .A1(n17470), .A2(n17471), .ZN(n17043) );
  INV_X1 U17286 ( .A(n17472), .ZN(n17471) );
  OR2_X1 U17287 ( .A1(n17473), .A2(n17474), .ZN(n17472) );
  AND2_X1 U17288 ( .A1(n17474), .A2(n17473), .ZN(n17470) );
  AND2_X1 U17289 ( .A1(n17475), .A2(n17476), .ZN(n17473) );
  OR2_X1 U17290 ( .A1(n17477), .A2(n17478), .ZN(n17476) );
  INV_X1 U17291 ( .A(n17479), .ZN(n17478) );
  OR2_X1 U17292 ( .A1(n17479), .A2(n17480), .ZN(n17475) );
  INV_X1 U17293 ( .A(n17477), .ZN(n17480) );
  OR2_X1 U17294 ( .A1(n15038), .A2(n14801), .ZN(n17046) );
  OR2_X1 U17295 ( .A1(n17057), .A2(n17054), .ZN(n17402) );
  OR2_X1 U17296 ( .A1(n17481), .A2(n17482), .ZN(n17054) );
  INV_X1 U17297 ( .A(n17483), .ZN(n17482) );
  OR2_X1 U17298 ( .A1(n17484), .A2(n17485), .ZN(n17483) );
  AND2_X1 U17299 ( .A1(n17485), .A2(n17484), .ZN(n17481) );
  AND2_X1 U17300 ( .A1(n17486), .A2(n17487), .ZN(n17484) );
  OR2_X1 U17301 ( .A1(n17488), .A2(n17489), .ZN(n17487) );
  INV_X1 U17302 ( .A(n17490), .ZN(n17489) );
  OR2_X1 U17303 ( .A1(n17490), .A2(n17491), .ZN(n17486) );
  INV_X1 U17304 ( .A(n17488), .ZN(n17491) );
  OR2_X1 U17305 ( .A1(n15072), .A2(n14801), .ZN(n17057) );
  OR2_X1 U17306 ( .A1(n17068), .A2(n17065), .ZN(n17399) );
  OR2_X1 U17307 ( .A1(n17492), .A2(n17493), .ZN(n17065) );
  INV_X1 U17308 ( .A(n17494), .ZN(n17493) );
  OR2_X1 U17309 ( .A1(n17495), .A2(n17496), .ZN(n17494) );
  AND2_X1 U17310 ( .A1(n17496), .A2(n17495), .ZN(n17492) );
  AND2_X1 U17311 ( .A1(n17497), .A2(n17498), .ZN(n17495) );
  OR2_X1 U17312 ( .A1(n17499), .A2(n17500), .ZN(n17498) );
  INV_X1 U17313 ( .A(n17501), .ZN(n17500) );
  OR2_X1 U17314 ( .A1(n17501), .A2(n17502), .ZN(n17497) );
  INV_X1 U17315 ( .A(n17499), .ZN(n17502) );
  OR2_X1 U17316 ( .A1(n15106), .A2(n14801), .ZN(n17068) );
  OR2_X1 U17317 ( .A1(n17079), .A2(n17076), .ZN(n17396) );
  OR2_X1 U17318 ( .A1(n17503), .A2(n17504), .ZN(n17076) );
  INV_X1 U17319 ( .A(n17505), .ZN(n17504) );
  OR2_X1 U17320 ( .A1(n17506), .A2(n17507), .ZN(n17505) );
  AND2_X1 U17321 ( .A1(n17507), .A2(n17506), .ZN(n17503) );
  AND2_X1 U17322 ( .A1(n17508), .A2(n17509), .ZN(n17506) );
  OR2_X1 U17323 ( .A1(n17510), .A2(n17511), .ZN(n17509) );
  INV_X1 U17324 ( .A(n17512), .ZN(n17511) );
  OR2_X1 U17325 ( .A1(n17512), .A2(n17513), .ZN(n17508) );
  INV_X1 U17326 ( .A(n17510), .ZN(n17513) );
  OR2_X1 U17327 ( .A1(n15140), .A2(n14801), .ZN(n17079) );
  OR2_X1 U17328 ( .A1(n17090), .A2(n17087), .ZN(n17393) );
  OR2_X1 U17329 ( .A1(n17514), .A2(n17515), .ZN(n17087) );
  INV_X1 U17330 ( .A(n17516), .ZN(n17515) );
  OR2_X1 U17331 ( .A1(n17517), .A2(n17518), .ZN(n17516) );
  AND2_X1 U17332 ( .A1(n17518), .A2(n17517), .ZN(n17514) );
  AND2_X1 U17333 ( .A1(n17519), .A2(n17520), .ZN(n17517) );
  OR2_X1 U17334 ( .A1(n17521), .A2(n17522), .ZN(n17520) );
  INV_X1 U17335 ( .A(n17523), .ZN(n17522) );
  OR2_X1 U17336 ( .A1(n17523), .A2(n17524), .ZN(n17519) );
  INV_X1 U17337 ( .A(n17521), .ZN(n17524) );
  OR2_X1 U17338 ( .A1(n15174), .A2(n14801), .ZN(n17090) );
  OR2_X1 U17339 ( .A1(n17101), .A2(n17098), .ZN(n17390) );
  OR2_X1 U17340 ( .A1(n17525), .A2(n17526), .ZN(n17098) );
  INV_X1 U17341 ( .A(n17527), .ZN(n17526) );
  OR2_X1 U17342 ( .A1(n17528), .A2(n17529), .ZN(n17527) );
  AND2_X1 U17343 ( .A1(n17529), .A2(n17528), .ZN(n17525) );
  AND2_X1 U17344 ( .A1(n17530), .A2(n17531), .ZN(n17528) );
  OR2_X1 U17345 ( .A1(n17532), .A2(n17533), .ZN(n17531) );
  INV_X1 U17346 ( .A(n17534), .ZN(n17533) );
  OR2_X1 U17347 ( .A1(n17534), .A2(n17535), .ZN(n17530) );
  INV_X1 U17348 ( .A(n17532), .ZN(n17535) );
  OR2_X1 U17349 ( .A1(n15208), .A2(n14801), .ZN(n17101) );
  OR2_X1 U17350 ( .A1(n17112), .A2(n17109), .ZN(n17387) );
  OR2_X1 U17351 ( .A1(n17536), .A2(n17537), .ZN(n17109) );
  INV_X1 U17352 ( .A(n17538), .ZN(n17537) );
  OR2_X1 U17353 ( .A1(n17539), .A2(n17540), .ZN(n17538) );
  AND2_X1 U17354 ( .A1(n17540), .A2(n17539), .ZN(n17536) );
  AND2_X1 U17355 ( .A1(n17541), .A2(n17542), .ZN(n17539) );
  OR2_X1 U17356 ( .A1(n17543), .A2(n17544), .ZN(n17542) );
  INV_X1 U17357 ( .A(n17545), .ZN(n17544) );
  OR2_X1 U17358 ( .A1(n17545), .A2(n17546), .ZN(n17541) );
  INV_X1 U17359 ( .A(n17543), .ZN(n17546) );
  OR2_X1 U17360 ( .A1(n15242), .A2(n14801), .ZN(n17112) );
  OR2_X1 U17361 ( .A1(n17123), .A2(n17120), .ZN(n17384) );
  OR2_X1 U17362 ( .A1(n17547), .A2(n17548), .ZN(n17120) );
  INV_X1 U17363 ( .A(n17549), .ZN(n17548) );
  OR2_X1 U17364 ( .A1(n17550), .A2(n17551), .ZN(n17549) );
  AND2_X1 U17365 ( .A1(n17551), .A2(n17550), .ZN(n17547) );
  AND2_X1 U17366 ( .A1(n17552), .A2(n17553), .ZN(n17550) );
  OR2_X1 U17367 ( .A1(n17554), .A2(n17555), .ZN(n17553) );
  INV_X1 U17368 ( .A(n17556), .ZN(n17555) );
  OR2_X1 U17369 ( .A1(n17556), .A2(n17557), .ZN(n17552) );
  INV_X1 U17370 ( .A(n17554), .ZN(n17557) );
  OR2_X1 U17371 ( .A1(n15287), .A2(n14801), .ZN(n17123) );
  OR2_X1 U17372 ( .A1(n17134), .A2(n17131), .ZN(n17381) );
  OR2_X1 U17373 ( .A1(n17558), .A2(n17559), .ZN(n17131) );
  INV_X1 U17374 ( .A(n17560), .ZN(n17559) );
  OR2_X1 U17375 ( .A1(n17561), .A2(n17562), .ZN(n17560) );
  AND2_X1 U17376 ( .A1(n17562), .A2(n17561), .ZN(n17558) );
  AND2_X1 U17377 ( .A1(n17563), .A2(n17564), .ZN(n17561) );
  OR2_X1 U17378 ( .A1(n17565), .A2(n17566), .ZN(n17564) );
  INV_X1 U17379 ( .A(n17567), .ZN(n17566) );
  OR2_X1 U17380 ( .A1(n17567), .A2(n17568), .ZN(n17563) );
  INV_X1 U17381 ( .A(n17565), .ZN(n17568) );
  OR2_X1 U17382 ( .A1(n15321), .A2(n14801), .ZN(n17134) );
  OR2_X1 U17383 ( .A1(n17145), .A2(n17142), .ZN(n17378) );
  OR2_X1 U17384 ( .A1(n17569), .A2(n17570), .ZN(n17142) );
  INV_X1 U17385 ( .A(n17571), .ZN(n17570) );
  OR2_X1 U17386 ( .A1(n17572), .A2(n17573), .ZN(n17571) );
  AND2_X1 U17387 ( .A1(n17573), .A2(n17572), .ZN(n17569) );
  AND2_X1 U17388 ( .A1(n17574), .A2(n17575), .ZN(n17572) );
  OR2_X1 U17389 ( .A1(n17576), .A2(n17577), .ZN(n17575) );
  INV_X1 U17390 ( .A(n17578), .ZN(n17577) );
  OR2_X1 U17391 ( .A1(n17578), .A2(n17579), .ZN(n17574) );
  INV_X1 U17392 ( .A(n17576), .ZN(n17579) );
  OR2_X1 U17393 ( .A1(n15355), .A2(n14801), .ZN(n17145) );
  OR2_X1 U17394 ( .A1(n17156), .A2(n17153), .ZN(n17375) );
  OR2_X1 U17395 ( .A1(n17580), .A2(n17581), .ZN(n17153) );
  INV_X1 U17396 ( .A(n17582), .ZN(n17581) );
  OR2_X1 U17397 ( .A1(n17583), .A2(n17584), .ZN(n17582) );
  AND2_X1 U17398 ( .A1(n17584), .A2(n17583), .ZN(n17580) );
  AND2_X1 U17399 ( .A1(n17585), .A2(n17586), .ZN(n17583) );
  OR2_X1 U17400 ( .A1(n17587), .A2(n17588), .ZN(n17586) );
  INV_X1 U17401 ( .A(n17589), .ZN(n17588) );
  OR2_X1 U17402 ( .A1(n17589), .A2(n17590), .ZN(n17585) );
  INV_X1 U17403 ( .A(n17587), .ZN(n17590) );
  OR2_X1 U17404 ( .A1(n15389), .A2(n14801), .ZN(n17156) );
  OR2_X1 U17405 ( .A1(n17167), .A2(n17164), .ZN(n17372) );
  OR2_X1 U17406 ( .A1(n17591), .A2(n17592), .ZN(n17164) );
  INV_X1 U17407 ( .A(n17593), .ZN(n17592) );
  OR2_X1 U17408 ( .A1(n17594), .A2(n17595), .ZN(n17593) );
  AND2_X1 U17409 ( .A1(n17595), .A2(n17594), .ZN(n17591) );
  AND2_X1 U17410 ( .A1(n17596), .A2(n17597), .ZN(n17594) );
  OR2_X1 U17411 ( .A1(n17598), .A2(n17599), .ZN(n17597) );
  INV_X1 U17412 ( .A(n17600), .ZN(n17599) );
  OR2_X1 U17413 ( .A1(n17600), .A2(n17601), .ZN(n17596) );
  INV_X1 U17414 ( .A(n17598), .ZN(n17601) );
  OR2_X1 U17415 ( .A1(n15423), .A2(n14801), .ZN(n17167) );
  OR2_X1 U17416 ( .A1(n17178), .A2(n17175), .ZN(n17369) );
  OR2_X1 U17417 ( .A1(n17602), .A2(n17603), .ZN(n17175) );
  INV_X1 U17418 ( .A(n17604), .ZN(n17603) );
  OR2_X1 U17419 ( .A1(n17605), .A2(n17606), .ZN(n17604) );
  AND2_X1 U17420 ( .A1(n17606), .A2(n17605), .ZN(n17602) );
  AND2_X1 U17421 ( .A1(n17607), .A2(n17608), .ZN(n17605) );
  OR2_X1 U17422 ( .A1(n17609), .A2(n17610), .ZN(n17608) );
  INV_X1 U17423 ( .A(n17611), .ZN(n17610) );
  OR2_X1 U17424 ( .A1(n17611), .A2(n17612), .ZN(n17607) );
  INV_X1 U17425 ( .A(n17609), .ZN(n17612) );
  OR2_X1 U17426 ( .A1(n15457), .A2(n14801), .ZN(n17178) );
  OR2_X1 U17427 ( .A1(n17189), .A2(n17186), .ZN(n17366) );
  OR2_X1 U17428 ( .A1(n17613), .A2(n17614), .ZN(n17186) );
  INV_X1 U17429 ( .A(n17615), .ZN(n17614) );
  OR2_X1 U17430 ( .A1(n17616), .A2(n17617), .ZN(n17615) );
  AND2_X1 U17431 ( .A1(n17617), .A2(n17616), .ZN(n17613) );
  AND2_X1 U17432 ( .A1(n17618), .A2(n17619), .ZN(n17616) );
  OR2_X1 U17433 ( .A1(n17620), .A2(n17621), .ZN(n17619) );
  INV_X1 U17434 ( .A(n17622), .ZN(n17621) );
  OR2_X1 U17435 ( .A1(n17622), .A2(n17623), .ZN(n17618) );
  INV_X1 U17436 ( .A(n17620), .ZN(n17623) );
  OR2_X1 U17437 ( .A1(n15491), .A2(n14801), .ZN(n17189) );
  OR2_X1 U17438 ( .A1(n17200), .A2(n17197), .ZN(n17363) );
  OR2_X1 U17439 ( .A1(n17624), .A2(n17625), .ZN(n17197) );
  INV_X1 U17440 ( .A(n17626), .ZN(n17625) );
  OR2_X1 U17441 ( .A1(n17627), .A2(n17628), .ZN(n17626) );
  AND2_X1 U17442 ( .A1(n17628), .A2(n17627), .ZN(n17624) );
  AND2_X1 U17443 ( .A1(n17629), .A2(n17630), .ZN(n17627) );
  OR2_X1 U17444 ( .A1(n17631), .A2(n17632), .ZN(n17630) );
  INV_X1 U17445 ( .A(n17633), .ZN(n17632) );
  OR2_X1 U17446 ( .A1(n17633), .A2(n17634), .ZN(n17629) );
  INV_X1 U17447 ( .A(n17631), .ZN(n17634) );
  OR2_X1 U17448 ( .A1(n15525), .A2(n14801), .ZN(n17200) );
  OR2_X1 U17449 ( .A1(n17211), .A2(n17208), .ZN(n17360) );
  OR2_X1 U17450 ( .A1(n17635), .A2(n17636), .ZN(n17208) );
  INV_X1 U17451 ( .A(n17637), .ZN(n17636) );
  OR2_X1 U17452 ( .A1(n17638), .A2(n17639), .ZN(n17637) );
  AND2_X1 U17453 ( .A1(n17639), .A2(n17638), .ZN(n17635) );
  AND2_X1 U17454 ( .A1(n17640), .A2(n17641), .ZN(n17638) );
  OR2_X1 U17455 ( .A1(n17642), .A2(n17643), .ZN(n17641) );
  INV_X1 U17456 ( .A(n17644), .ZN(n17643) );
  OR2_X1 U17457 ( .A1(n17644), .A2(n17645), .ZN(n17640) );
  INV_X1 U17458 ( .A(n17642), .ZN(n17645) );
  OR2_X1 U17459 ( .A1(n15559), .A2(n14801), .ZN(n17211) );
  OR2_X1 U17460 ( .A1(n17222), .A2(n17219), .ZN(n17357) );
  OR2_X1 U17461 ( .A1(n17646), .A2(n17647), .ZN(n17219) );
  INV_X1 U17462 ( .A(n17648), .ZN(n17647) );
  OR2_X1 U17463 ( .A1(n17649), .A2(n17650), .ZN(n17648) );
  AND2_X1 U17464 ( .A1(n17650), .A2(n17649), .ZN(n17646) );
  AND2_X1 U17465 ( .A1(n17651), .A2(n17652), .ZN(n17649) );
  OR2_X1 U17466 ( .A1(n17653), .A2(n17654), .ZN(n17652) );
  INV_X1 U17467 ( .A(n17655), .ZN(n17654) );
  OR2_X1 U17468 ( .A1(n17655), .A2(n17656), .ZN(n17651) );
  INV_X1 U17469 ( .A(n17653), .ZN(n17656) );
  OR2_X1 U17470 ( .A1(n15593), .A2(n14801), .ZN(n17222) );
  OR2_X1 U17471 ( .A1(n17233), .A2(n17230), .ZN(n17354) );
  OR2_X1 U17472 ( .A1(n17657), .A2(n17658), .ZN(n17230) );
  INV_X1 U17473 ( .A(n17659), .ZN(n17658) );
  OR2_X1 U17474 ( .A1(n17660), .A2(n17661), .ZN(n17659) );
  AND2_X1 U17475 ( .A1(n17661), .A2(n17660), .ZN(n17657) );
  AND2_X1 U17476 ( .A1(n17662), .A2(n17663), .ZN(n17660) );
  OR2_X1 U17477 ( .A1(n17664), .A2(n17665), .ZN(n17663) );
  INV_X1 U17478 ( .A(n17666), .ZN(n17665) );
  OR2_X1 U17479 ( .A1(n17666), .A2(n17667), .ZN(n17662) );
  INV_X1 U17480 ( .A(n17664), .ZN(n17667) );
  OR2_X1 U17481 ( .A1(n15638), .A2(n14801), .ZN(n17233) );
  OR2_X1 U17482 ( .A1(n17244), .A2(n17241), .ZN(n17351) );
  OR2_X1 U17483 ( .A1(n17668), .A2(n17669), .ZN(n17241) );
  INV_X1 U17484 ( .A(n17670), .ZN(n17669) );
  OR2_X1 U17485 ( .A1(n17671), .A2(n17672), .ZN(n17670) );
  AND2_X1 U17486 ( .A1(n17672), .A2(n17671), .ZN(n17668) );
  AND2_X1 U17487 ( .A1(n17673), .A2(n17674), .ZN(n17671) );
  OR2_X1 U17488 ( .A1(n17675), .A2(n17676), .ZN(n17674) );
  INV_X1 U17489 ( .A(n17677), .ZN(n17676) );
  OR2_X1 U17490 ( .A1(n17677), .A2(n17678), .ZN(n17673) );
  INV_X1 U17491 ( .A(n17675), .ZN(n17678) );
  OR2_X1 U17492 ( .A1(n15672), .A2(n14801), .ZN(n17244) );
  OR2_X1 U17493 ( .A1(n17255), .A2(n17252), .ZN(n17348) );
  OR2_X1 U17494 ( .A1(n17679), .A2(n17680), .ZN(n17252) );
  INV_X1 U17495 ( .A(n17681), .ZN(n17680) );
  OR2_X1 U17496 ( .A1(n17682), .A2(n17683), .ZN(n17681) );
  AND2_X1 U17497 ( .A1(n17683), .A2(n17682), .ZN(n17679) );
  AND2_X1 U17498 ( .A1(n17684), .A2(n17685), .ZN(n17682) );
  OR2_X1 U17499 ( .A1(n17686), .A2(n17687), .ZN(n17685) );
  INV_X1 U17500 ( .A(n17688), .ZN(n17687) );
  OR2_X1 U17501 ( .A1(n17688), .A2(n17689), .ZN(n17684) );
  INV_X1 U17502 ( .A(n17686), .ZN(n17689) );
  OR2_X1 U17503 ( .A1(n15706), .A2(n14801), .ZN(n17255) );
  OR2_X1 U17504 ( .A1(n17266), .A2(n17263), .ZN(n17345) );
  OR2_X1 U17505 ( .A1(n17690), .A2(n17691), .ZN(n17263) );
  INV_X1 U17506 ( .A(n17692), .ZN(n17691) );
  OR2_X1 U17507 ( .A1(n17693), .A2(n17694), .ZN(n17692) );
  AND2_X1 U17508 ( .A1(n17694), .A2(n17693), .ZN(n17690) );
  AND2_X1 U17509 ( .A1(n17695), .A2(n17696), .ZN(n17693) );
  OR2_X1 U17510 ( .A1(n17697), .A2(n17698), .ZN(n17696) );
  INV_X1 U17511 ( .A(n17699), .ZN(n17698) );
  OR2_X1 U17512 ( .A1(n17699), .A2(n17700), .ZN(n17695) );
  INV_X1 U17513 ( .A(n17697), .ZN(n17700) );
  OR2_X1 U17514 ( .A1(n15740), .A2(n14801), .ZN(n17266) );
  OR2_X1 U17515 ( .A1(n17277), .A2(n17274), .ZN(n17342) );
  OR2_X1 U17516 ( .A1(n17701), .A2(n17702), .ZN(n17274) );
  INV_X1 U17517 ( .A(n17703), .ZN(n17702) );
  OR2_X1 U17518 ( .A1(n17704), .A2(n17705), .ZN(n17703) );
  AND2_X1 U17519 ( .A1(n17705), .A2(n17704), .ZN(n17701) );
  AND2_X1 U17520 ( .A1(n17706), .A2(n17707), .ZN(n17704) );
  OR2_X1 U17521 ( .A1(n17708), .A2(n17709), .ZN(n17707) );
  INV_X1 U17522 ( .A(n17710), .ZN(n17709) );
  OR2_X1 U17523 ( .A1(n17710), .A2(n17711), .ZN(n17706) );
  INV_X1 U17524 ( .A(n17708), .ZN(n17711) );
  OR2_X1 U17525 ( .A1(n15774), .A2(n14801), .ZN(n17277) );
  OR2_X1 U17526 ( .A1(n17288), .A2(n17285), .ZN(n17339) );
  OR2_X1 U17527 ( .A1(n17712), .A2(n17713), .ZN(n17285) );
  INV_X1 U17528 ( .A(n17714), .ZN(n17713) );
  OR2_X1 U17529 ( .A1(n17715), .A2(n17716), .ZN(n17714) );
  AND2_X1 U17530 ( .A1(n17716), .A2(n17715), .ZN(n17712) );
  AND2_X1 U17531 ( .A1(n17717), .A2(n17718), .ZN(n17715) );
  OR2_X1 U17532 ( .A1(n17719), .A2(n17720), .ZN(n17718) );
  INV_X1 U17533 ( .A(n17721), .ZN(n17720) );
  OR2_X1 U17534 ( .A1(n17721), .A2(n17722), .ZN(n17717) );
  INV_X1 U17535 ( .A(n17719), .ZN(n17722) );
  OR2_X1 U17536 ( .A1(n15808), .A2(n14801), .ZN(n17288) );
  OR2_X1 U17537 ( .A1(n17299), .A2(n17296), .ZN(n17336) );
  OR2_X1 U17538 ( .A1(n17723), .A2(n17724), .ZN(n17296) );
  INV_X1 U17539 ( .A(n17725), .ZN(n17724) );
  OR2_X1 U17540 ( .A1(n17726), .A2(n17727), .ZN(n17725) );
  AND2_X1 U17541 ( .A1(n17727), .A2(n17726), .ZN(n17723) );
  AND2_X1 U17542 ( .A1(n17728), .A2(n17729), .ZN(n17726) );
  OR2_X1 U17543 ( .A1(n17730), .A2(n17731), .ZN(n17729) );
  INV_X1 U17544 ( .A(n17732), .ZN(n17731) );
  OR2_X1 U17545 ( .A1(n17732), .A2(n17733), .ZN(n17728) );
  INV_X1 U17546 ( .A(n17730), .ZN(n17733) );
  OR2_X1 U17547 ( .A1(n15842), .A2(n14801), .ZN(n17299) );
  INV_X1 U17548 ( .A(b_30_), .ZN(n14801) );
  OR2_X1 U17549 ( .A1(n17734), .A2(n17735), .ZN(n17324) );
  INV_X1 U17550 ( .A(n17736), .ZN(n17735) );
  OR2_X1 U17551 ( .A1(n17737), .A2(n17738), .ZN(n17736) );
  AND2_X1 U17552 ( .A1(n17738), .A2(n17737), .ZN(n17734) );
  AND2_X1 U17553 ( .A1(n17739), .A2(n17740), .ZN(n17737) );
  OR2_X1 U17554 ( .A1(n17741), .A2(n17742), .ZN(n17740) );
  INV_X1 U17555 ( .A(n17743), .ZN(n17742) );
  OR2_X1 U17556 ( .A1(n17743), .A2(n17744), .ZN(n17739) );
  INV_X1 U17557 ( .A(n17741), .ZN(n17744) );
  AND3_X1 U17558 ( .A1(n16875), .A2(n16877), .A3(n16876), .ZN(n16011) );
  INV_X1 U17559 ( .A(n16885), .ZN(n16876) );
  OR2_X1 U17560 ( .A1(n17745), .A2(n17746), .ZN(n16885) );
  AND2_X1 U17561 ( .A1(n17315), .A2(n17313), .ZN(n17746) );
  AND2_X1 U17562 ( .A1(n17311), .A2(n17747), .ZN(n17745) );
  OR2_X1 U17563 ( .A1(n17315), .A2(n17313), .ZN(n17747) );
  OR2_X1 U17564 ( .A1(n17748), .A2(n17749), .ZN(n17313) );
  AND2_X1 U17565 ( .A1(n17741), .A2(n17743), .ZN(n17749) );
  AND2_X1 U17566 ( .A1(n17738), .A2(n17750), .ZN(n17748) );
  OR2_X1 U17567 ( .A1(n17741), .A2(n17743), .ZN(n17750) );
  OR2_X1 U17568 ( .A1(n17751), .A2(n17752), .ZN(n17743) );
  AND2_X1 U17569 ( .A1(n17730), .A2(n17732), .ZN(n17752) );
  AND2_X1 U17570 ( .A1(n17727), .A2(n17753), .ZN(n17751) );
  OR2_X1 U17571 ( .A1(n17730), .A2(n17732), .ZN(n17753) );
  OR2_X1 U17572 ( .A1(n17754), .A2(n17755), .ZN(n17732) );
  AND2_X1 U17573 ( .A1(n17719), .A2(n17721), .ZN(n17755) );
  AND2_X1 U17574 ( .A1(n17716), .A2(n17756), .ZN(n17754) );
  OR2_X1 U17575 ( .A1(n17719), .A2(n17721), .ZN(n17756) );
  OR2_X1 U17576 ( .A1(n17757), .A2(n17758), .ZN(n17721) );
  AND2_X1 U17577 ( .A1(n17708), .A2(n17710), .ZN(n17758) );
  AND2_X1 U17578 ( .A1(n17705), .A2(n17759), .ZN(n17757) );
  OR2_X1 U17579 ( .A1(n17708), .A2(n17710), .ZN(n17759) );
  OR2_X1 U17580 ( .A1(n17760), .A2(n17761), .ZN(n17710) );
  AND2_X1 U17581 ( .A1(n17697), .A2(n17699), .ZN(n17761) );
  AND2_X1 U17582 ( .A1(n17694), .A2(n17762), .ZN(n17760) );
  OR2_X1 U17583 ( .A1(n17697), .A2(n17699), .ZN(n17762) );
  OR2_X1 U17584 ( .A1(n17763), .A2(n17764), .ZN(n17699) );
  AND2_X1 U17585 ( .A1(n17686), .A2(n17688), .ZN(n17764) );
  AND2_X1 U17586 ( .A1(n17683), .A2(n17765), .ZN(n17763) );
  OR2_X1 U17587 ( .A1(n17686), .A2(n17688), .ZN(n17765) );
  OR2_X1 U17588 ( .A1(n17766), .A2(n17767), .ZN(n17688) );
  AND2_X1 U17589 ( .A1(n17675), .A2(n17677), .ZN(n17767) );
  AND2_X1 U17590 ( .A1(n17672), .A2(n17768), .ZN(n17766) );
  OR2_X1 U17591 ( .A1(n17675), .A2(n17677), .ZN(n17768) );
  OR2_X1 U17592 ( .A1(n17769), .A2(n17770), .ZN(n17677) );
  AND2_X1 U17593 ( .A1(n17664), .A2(n17666), .ZN(n17770) );
  AND2_X1 U17594 ( .A1(n17661), .A2(n17771), .ZN(n17769) );
  OR2_X1 U17595 ( .A1(n17664), .A2(n17666), .ZN(n17771) );
  OR2_X1 U17596 ( .A1(n17772), .A2(n17773), .ZN(n17666) );
  AND2_X1 U17597 ( .A1(n17653), .A2(n17655), .ZN(n17773) );
  AND2_X1 U17598 ( .A1(n17650), .A2(n17774), .ZN(n17772) );
  OR2_X1 U17599 ( .A1(n17653), .A2(n17655), .ZN(n17774) );
  OR2_X1 U17600 ( .A1(n17775), .A2(n17776), .ZN(n17655) );
  AND2_X1 U17601 ( .A1(n17642), .A2(n17644), .ZN(n17776) );
  AND2_X1 U17602 ( .A1(n17639), .A2(n17777), .ZN(n17775) );
  OR2_X1 U17603 ( .A1(n17642), .A2(n17644), .ZN(n17777) );
  OR2_X1 U17604 ( .A1(n17778), .A2(n17779), .ZN(n17644) );
  AND2_X1 U17605 ( .A1(n17631), .A2(n17633), .ZN(n17779) );
  AND2_X1 U17606 ( .A1(n17628), .A2(n17780), .ZN(n17778) );
  OR2_X1 U17607 ( .A1(n17631), .A2(n17633), .ZN(n17780) );
  OR2_X1 U17608 ( .A1(n17781), .A2(n17782), .ZN(n17633) );
  AND2_X1 U17609 ( .A1(n17620), .A2(n17622), .ZN(n17782) );
  AND2_X1 U17610 ( .A1(n17617), .A2(n17783), .ZN(n17781) );
  OR2_X1 U17611 ( .A1(n17620), .A2(n17622), .ZN(n17783) );
  OR2_X1 U17612 ( .A1(n17784), .A2(n17785), .ZN(n17622) );
  AND2_X1 U17613 ( .A1(n17609), .A2(n17611), .ZN(n17785) );
  AND2_X1 U17614 ( .A1(n17606), .A2(n17786), .ZN(n17784) );
  OR2_X1 U17615 ( .A1(n17609), .A2(n17611), .ZN(n17786) );
  OR2_X1 U17616 ( .A1(n17787), .A2(n17788), .ZN(n17611) );
  AND2_X1 U17617 ( .A1(n17598), .A2(n17600), .ZN(n17788) );
  AND2_X1 U17618 ( .A1(n17595), .A2(n17789), .ZN(n17787) );
  OR2_X1 U17619 ( .A1(n17598), .A2(n17600), .ZN(n17789) );
  OR2_X1 U17620 ( .A1(n17790), .A2(n17791), .ZN(n17600) );
  AND2_X1 U17621 ( .A1(n17587), .A2(n17589), .ZN(n17791) );
  AND2_X1 U17622 ( .A1(n17584), .A2(n17792), .ZN(n17790) );
  OR2_X1 U17623 ( .A1(n17587), .A2(n17589), .ZN(n17792) );
  OR2_X1 U17624 ( .A1(n17793), .A2(n17794), .ZN(n17589) );
  AND2_X1 U17625 ( .A1(n17576), .A2(n17578), .ZN(n17794) );
  AND2_X1 U17626 ( .A1(n17573), .A2(n17795), .ZN(n17793) );
  OR2_X1 U17627 ( .A1(n17576), .A2(n17578), .ZN(n17795) );
  OR2_X1 U17628 ( .A1(n17796), .A2(n17797), .ZN(n17578) );
  AND2_X1 U17629 ( .A1(n17565), .A2(n17567), .ZN(n17797) );
  AND2_X1 U17630 ( .A1(n17562), .A2(n17798), .ZN(n17796) );
  OR2_X1 U17631 ( .A1(n17565), .A2(n17567), .ZN(n17798) );
  OR2_X1 U17632 ( .A1(n17799), .A2(n17800), .ZN(n17567) );
  AND2_X1 U17633 ( .A1(n17554), .A2(n17556), .ZN(n17800) );
  AND2_X1 U17634 ( .A1(n17551), .A2(n17801), .ZN(n17799) );
  OR2_X1 U17635 ( .A1(n17554), .A2(n17556), .ZN(n17801) );
  OR2_X1 U17636 ( .A1(n17802), .A2(n17803), .ZN(n17556) );
  AND2_X1 U17637 ( .A1(n17543), .A2(n17545), .ZN(n17803) );
  AND2_X1 U17638 ( .A1(n17540), .A2(n17804), .ZN(n17802) );
  OR2_X1 U17639 ( .A1(n17543), .A2(n17545), .ZN(n17804) );
  OR2_X1 U17640 ( .A1(n17805), .A2(n17806), .ZN(n17545) );
  AND2_X1 U17641 ( .A1(n17532), .A2(n17534), .ZN(n17806) );
  AND2_X1 U17642 ( .A1(n17529), .A2(n17807), .ZN(n17805) );
  OR2_X1 U17643 ( .A1(n17532), .A2(n17534), .ZN(n17807) );
  OR2_X1 U17644 ( .A1(n17808), .A2(n17809), .ZN(n17534) );
  AND2_X1 U17645 ( .A1(n17521), .A2(n17523), .ZN(n17809) );
  AND2_X1 U17646 ( .A1(n17518), .A2(n17810), .ZN(n17808) );
  OR2_X1 U17647 ( .A1(n17521), .A2(n17523), .ZN(n17810) );
  OR2_X1 U17648 ( .A1(n17811), .A2(n17812), .ZN(n17523) );
  AND2_X1 U17649 ( .A1(n17510), .A2(n17512), .ZN(n17812) );
  AND2_X1 U17650 ( .A1(n17507), .A2(n17813), .ZN(n17811) );
  OR2_X1 U17651 ( .A1(n17510), .A2(n17512), .ZN(n17813) );
  OR2_X1 U17652 ( .A1(n17814), .A2(n17815), .ZN(n17512) );
  AND2_X1 U17653 ( .A1(n17499), .A2(n17501), .ZN(n17815) );
  AND2_X1 U17654 ( .A1(n17496), .A2(n17816), .ZN(n17814) );
  OR2_X1 U17655 ( .A1(n17499), .A2(n17501), .ZN(n17816) );
  OR2_X1 U17656 ( .A1(n17817), .A2(n17818), .ZN(n17501) );
  AND2_X1 U17657 ( .A1(n17488), .A2(n17490), .ZN(n17818) );
  AND2_X1 U17658 ( .A1(n17485), .A2(n17819), .ZN(n17817) );
  OR2_X1 U17659 ( .A1(n17488), .A2(n17490), .ZN(n17819) );
  OR2_X1 U17660 ( .A1(n17820), .A2(n17821), .ZN(n17490) );
  AND2_X1 U17661 ( .A1(n17477), .A2(n17479), .ZN(n17821) );
  AND2_X1 U17662 ( .A1(n17474), .A2(n17822), .ZN(n17820) );
  OR2_X1 U17663 ( .A1(n17477), .A2(n17479), .ZN(n17822) );
  OR2_X1 U17664 ( .A1(n17823), .A2(n17824), .ZN(n17479) );
  AND2_X1 U17665 ( .A1(n17466), .A2(n17468), .ZN(n17824) );
  AND2_X1 U17666 ( .A1(n17463), .A2(n17825), .ZN(n17823) );
  OR2_X1 U17667 ( .A1(n17466), .A2(n17468), .ZN(n17825) );
  OR2_X1 U17668 ( .A1(n17826), .A2(n17827), .ZN(n17468) );
  AND2_X1 U17669 ( .A1(n17455), .A2(n17457), .ZN(n17827) );
  AND2_X1 U17670 ( .A1(n17452), .A2(n17828), .ZN(n17826) );
  OR2_X1 U17671 ( .A1(n17455), .A2(n17457), .ZN(n17828) );
  OR2_X1 U17672 ( .A1(n17829), .A2(n17830), .ZN(n17457) );
  AND2_X1 U17673 ( .A1(n17444), .A2(n17446), .ZN(n17830) );
  AND2_X1 U17674 ( .A1(n17441), .A2(n17831), .ZN(n17829) );
  OR2_X1 U17675 ( .A1(n17444), .A2(n17446), .ZN(n17831) );
  OR2_X1 U17676 ( .A1(n17832), .A2(n17833), .ZN(n17446) );
  AND2_X1 U17677 ( .A1(n15954), .A2(n17434), .ZN(n17833) );
  AND2_X1 U17678 ( .A1(n17433), .A2(n17834), .ZN(n17832) );
  OR2_X1 U17679 ( .A1(n15954), .A2(n17434), .ZN(n17834) );
  INV_X1 U17680 ( .A(n17435), .ZN(n17434) );
  AND3_X1 U17681 ( .A1(b_29_), .A2(b_28_), .A3(n15957), .ZN(n17435) );
  OR2_X1 U17682 ( .A1(n14857), .A2(n14856), .ZN(n15954) );
  INV_X1 U17683 ( .A(n17436), .ZN(n17433) );
  OR2_X1 U17684 ( .A1(n17835), .A2(n17836), .ZN(n17436) );
  AND2_X1 U17685 ( .A1(b_28_), .A2(n17837), .ZN(n17836) );
  OR2_X1 U17686 ( .A1(n17838), .A2(n16981), .ZN(n17837) );
  AND2_X1 U17687 ( .A1(a_30_), .A2(n14935), .ZN(n17838) );
  AND2_X1 U17688 ( .A1(b_27_), .A2(n17839), .ZN(n17835) );
  OR2_X1 U17689 ( .A1(n17840), .A2(n14817), .ZN(n17839) );
  AND2_X1 U17690 ( .A1(a_31_), .A2(n14890), .ZN(n17840) );
  OR2_X1 U17691 ( .A1(n14891), .A2(n14856), .ZN(n17444) );
  OR2_X1 U17692 ( .A1(n17841), .A2(n17842), .ZN(n17441) );
  AND2_X1 U17693 ( .A1(n17843), .A2(n17844), .ZN(n17842) );
  INV_X1 U17694 ( .A(n17845), .ZN(n17841) );
  OR2_X1 U17695 ( .A1(n17843), .A2(n17844), .ZN(n17845) );
  OR2_X1 U17696 ( .A1(n17846), .A2(n17847), .ZN(n17843) );
  AND2_X1 U17697 ( .A1(n17848), .A2(n17849), .ZN(n17847) );
  AND2_X1 U17698 ( .A1(n17850), .A2(n17851), .ZN(n17846) );
  OR2_X1 U17699 ( .A1(n14936), .A2(n14856), .ZN(n17455) );
  OR2_X1 U17700 ( .A1(n17852), .A2(n17853), .ZN(n17452) );
  INV_X1 U17701 ( .A(n17854), .ZN(n17853) );
  OR2_X1 U17702 ( .A1(n17855), .A2(n17856), .ZN(n17854) );
  AND2_X1 U17703 ( .A1(n17856), .A2(n17855), .ZN(n17852) );
  AND2_X1 U17704 ( .A1(n17857), .A2(n17858), .ZN(n17855) );
  OR2_X1 U17705 ( .A1(n15951), .A2(n17859), .ZN(n17858) );
  INV_X1 U17706 ( .A(n17860), .ZN(n17859) );
  OR2_X1 U17707 ( .A1(n17860), .A2(n17861), .ZN(n17857) );
  INV_X1 U17708 ( .A(n15951), .ZN(n17861) );
  OR2_X1 U17709 ( .A1(n14970), .A2(n14856), .ZN(n17466) );
  OR2_X1 U17710 ( .A1(n17862), .A2(n17863), .ZN(n17463) );
  INV_X1 U17711 ( .A(n17864), .ZN(n17863) );
  OR2_X1 U17712 ( .A1(n17865), .A2(n17866), .ZN(n17864) );
  AND2_X1 U17713 ( .A1(n17866), .A2(n17865), .ZN(n17862) );
  AND2_X1 U17714 ( .A1(n17867), .A2(n17868), .ZN(n17865) );
  OR2_X1 U17715 ( .A1(n17869), .A2(n17870), .ZN(n17868) );
  INV_X1 U17716 ( .A(n17871), .ZN(n17870) );
  OR2_X1 U17717 ( .A1(n17871), .A2(n17872), .ZN(n17867) );
  INV_X1 U17718 ( .A(n17869), .ZN(n17872) );
  OR2_X1 U17719 ( .A1(n15004), .A2(n14856), .ZN(n17477) );
  OR2_X1 U17720 ( .A1(n17873), .A2(n17874), .ZN(n17474) );
  INV_X1 U17721 ( .A(n17875), .ZN(n17874) );
  OR2_X1 U17722 ( .A1(n17876), .A2(n17877), .ZN(n17875) );
  AND2_X1 U17723 ( .A1(n17877), .A2(n17876), .ZN(n17873) );
  AND2_X1 U17724 ( .A1(n17878), .A2(n17879), .ZN(n17876) );
  OR2_X1 U17725 ( .A1(n17880), .A2(n17881), .ZN(n17879) );
  INV_X1 U17726 ( .A(n17882), .ZN(n17881) );
  OR2_X1 U17727 ( .A1(n17882), .A2(n17883), .ZN(n17878) );
  INV_X1 U17728 ( .A(n17880), .ZN(n17883) );
  OR2_X1 U17729 ( .A1(n15038), .A2(n14856), .ZN(n17488) );
  OR2_X1 U17730 ( .A1(n17884), .A2(n17885), .ZN(n17485) );
  INV_X1 U17731 ( .A(n17886), .ZN(n17885) );
  OR2_X1 U17732 ( .A1(n17887), .A2(n17888), .ZN(n17886) );
  AND2_X1 U17733 ( .A1(n17888), .A2(n17887), .ZN(n17884) );
  AND2_X1 U17734 ( .A1(n17889), .A2(n17890), .ZN(n17887) );
  OR2_X1 U17735 ( .A1(n17891), .A2(n17892), .ZN(n17890) );
  INV_X1 U17736 ( .A(n17893), .ZN(n17892) );
  OR2_X1 U17737 ( .A1(n17893), .A2(n17894), .ZN(n17889) );
  INV_X1 U17738 ( .A(n17891), .ZN(n17894) );
  OR2_X1 U17739 ( .A1(n15072), .A2(n14856), .ZN(n17499) );
  OR2_X1 U17740 ( .A1(n17895), .A2(n17896), .ZN(n17496) );
  INV_X1 U17741 ( .A(n17897), .ZN(n17896) );
  OR2_X1 U17742 ( .A1(n17898), .A2(n17899), .ZN(n17897) );
  AND2_X1 U17743 ( .A1(n17899), .A2(n17898), .ZN(n17895) );
  AND2_X1 U17744 ( .A1(n17900), .A2(n17901), .ZN(n17898) );
  OR2_X1 U17745 ( .A1(n17902), .A2(n17903), .ZN(n17901) );
  INV_X1 U17746 ( .A(n17904), .ZN(n17903) );
  OR2_X1 U17747 ( .A1(n17904), .A2(n17905), .ZN(n17900) );
  INV_X1 U17748 ( .A(n17902), .ZN(n17905) );
  OR2_X1 U17749 ( .A1(n15106), .A2(n14856), .ZN(n17510) );
  OR2_X1 U17750 ( .A1(n17906), .A2(n17907), .ZN(n17507) );
  INV_X1 U17751 ( .A(n17908), .ZN(n17907) );
  OR2_X1 U17752 ( .A1(n17909), .A2(n17910), .ZN(n17908) );
  AND2_X1 U17753 ( .A1(n17910), .A2(n17909), .ZN(n17906) );
  AND2_X1 U17754 ( .A1(n17911), .A2(n17912), .ZN(n17909) );
  OR2_X1 U17755 ( .A1(n17913), .A2(n17914), .ZN(n17912) );
  INV_X1 U17756 ( .A(n17915), .ZN(n17914) );
  OR2_X1 U17757 ( .A1(n17915), .A2(n17916), .ZN(n17911) );
  INV_X1 U17758 ( .A(n17913), .ZN(n17916) );
  OR2_X1 U17759 ( .A1(n15140), .A2(n14856), .ZN(n17521) );
  OR2_X1 U17760 ( .A1(n17917), .A2(n17918), .ZN(n17518) );
  INV_X1 U17761 ( .A(n17919), .ZN(n17918) );
  OR2_X1 U17762 ( .A1(n17920), .A2(n17921), .ZN(n17919) );
  AND2_X1 U17763 ( .A1(n17921), .A2(n17920), .ZN(n17917) );
  AND2_X1 U17764 ( .A1(n17922), .A2(n17923), .ZN(n17920) );
  OR2_X1 U17765 ( .A1(n17924), .A2(n17925), .ZN(n17923) );
  INV_X1 U17766 ( .A(n17926), .ZN(n17925) );
  OR2_X1 U17767 ( .A1(n17926), .A2(n17927), .ZN(n17922) );
  INV_X1 U17768 ( .A(n17924), .ZN(n17927) );
  OR2_X1 U17769 ( .A1(n15174), .A2(n14856), .ZN(n17532) );
  OR2_X1 U17770 ( .A1(n17928), .A2(n17929), .ZN(n17529) );
  INV_X1 U17771 ( .A(n17930), .ZN(n17929) );
  OR2_X1 U17772 ( .A1(n17931), .A2(n17932), .ZN(n17930) );
  AND2_X1 U17773 ( .A1(n17932), .A2(n17931), .ZN(n17928) );
  AND2_X1 U17774 ( .A1(n17933), .A2(n17934), .ZN(n17931) );
  OR2_X1 U17775 ( .A1(n17935), .A2(n17936), .ZN(n17934) );
  INV_X1 U17776 ( .A(n17937), .ZN(n17936) );
  OR2_X1 U17777 ( .A1(n17937), .A2(n17938), .ZN(n17933) );
  INV_X1 U17778 ( .A(n17935), .ZN(n17938) );
  OR2_X1 U17779 ( .A1(n15208), .A2(n14856), .ZN(n17543) );
  OR2_X1 U17780 ( .A1(n17939), .A2(n17940), .ZN(n17540) );
  INV_X1 U17781 ( .A(n17941), .ZN(n17940) );
  OR2_X1 U17782 ( .A1(n17942), .A2(n17943), .ZN(n17941) );
  AND2_X1 U17783 ( .A1(n17943), .A2(n17942), .ZN(n17939) );
  AND2_X1 U17784 ( .A1(n17944), .A2(n17945), .ZN(n17942) );
  OR2_X1 U17785 ( .A1(n17946), .A2(n17947), .ZN(n17945) );
  INV_X1 U17786 ( .A(n17948), .ZN(n17947) );
  OR2_X1 U17787 ( .A1(n17948), .A2(n17949), .ZN(n17944) );
  INV_X1 U17788 ( .A(n17946), .ZN(n17949) );
  OR2_X1 U17789 ( .A1(n15242), .A2(n14856), .ZN(n17554) );
  OR2_X1 U17790 ( .A1(n17950), .A2(n17951), .ZN(n17551) );
  INV_X1 U17791 ( .A(n17952), .ZN(n17951) );
  OR2_X1 U17792 ( .A1(n17953), .A2(n17954), .ZN(n17952) );
  AND2_X1 U17793 ( .A1(n17954), .A2(n17953), .ZN(n17950) );
  AND2_X1 U17794 ( .A1(n17955), .A2(n17956), .ZN(n17953) );
  OR2_X1 U17795 ( .A1(n17957), .A2(n17958), .ZN(n17956) );
  INV_X1 U17796 ( .A(n17959), .ZN(n17958) );
  OR2_X1 U17797 ( .A1(n17959), .A2(n17960), .ZN(n17955) );
  INV_X1 U17798 ( .A(n17957), .ZN(n17960) );
  OR2_X1 U17799 ( .A1(n15287), .A2(n14856), .ZN(n17565) );
  OR2_X1 U17800 ( .A1(n17961), .A2(n17962), .ZN(n17562) );
  INV_X1 U17801 ( .A(n17963), .ZN(n17962) );
  OR2_X1 U17802 ( .A1(n17964), .A2(n17965), .ZN(n17963) );
  AND2_X1 U17803 ( .A1(n17965), .A2(n17964), .ZN(n17961) );
  AND2_X1 U17804 ( .A1(n17966), .A2(n17967), .ZN(n17964) );
  OR2_X1 U17805 ( .A1(n17968), .A2(n17969), .ZN(n17967) );
  INV_X1 U17806 ( .A(n17970), .ZN(n17969) );
  OR2_X1 U17807 ( .A1(n17970), .A2(n17971), .ZN(n17966) );
  INV_X1 U17808 ( .A(n17968), .ZN(n17971) );
  OR2_X1 U17809 ( .A1(n15321), .A2(n14856), .ZN(n17576) );
  OR2_X1 U17810 ( .A1(n17972), .A2(n17973), .ZN(n17573) );
  INV_X1 U17811 ( .A(n17974), .ZN(n17973) );
  OR2_X1 U17812 ( .A1(n17975), .A2(n17976), .ZN(n17974) );
  AND2_X1 U17813 ( .A1(n17976), .A2(n17975), .ZN(n17972) );
  AND2_X1 U17814 ( .A1(n17977), .A2(n17978), .ZN(n17975) );
  OR2_X1 U17815 ( .A1(n17979), .A2(n17980), .ZN(n17978) );
  INV_X1 U17816 ( .A(n17981), .ZN(n17980) );
  OR2_X1 U17817 ( .A1(n17981), .A2(n17982), .ZN(n17977) );
  INV_X1 U17818 ( .A(n17979), .ZN(n17982) );
  OR2_X1 U17819 ( .A1(n15355), .A2(n14856), .ZN(n17587) );
  OR2_X1 U17820 ( .A1(n17983), .A2(n17984), .ZN(n17584) );
  INV_X1 U17821 ( .A(n17985), .ZN(n17984) );
  OR2_X1 U17822 ( .A1(n17986), .A2(n17987), .ZN(n17985) );
  AND2_X1 U17823 ( .A1(n17987), .A2(n17986), .ZN(n17983) );
  AND2_X1 U17824 ( .A1(n17988), .A2(n17989), .ZN(n17986) );
  OR2_X1 U17825 ( .A1(n17990), .A2(n17991), .ZN(n17989) );
  INV_X1 U17826 ( .A(n17992), .ZN(n17991) );
  OR2_X1 U17827 ( .A1(n17992), .A2(n17993), .ZN(n17988) );
  INV_X1 U17828 ( .A(n17990), .ZN(n17993) );
  OR2_X1 U17829 ( .A1(n15389), .A2(n14856), .ZN(n17598) );
  OR2_X1 U17830 ( .A1(n17994), .A2(n17995), .ZN(n17595) );
  INV_X1 U17831 ( .A(n17996), .ZN(n17995) );
  OR2_X1 U17832 ( .A1(n17997), .A2(n17998), .ZN(n17996) );
  AND2_X1 U17833 ( .A1(n17998), .A2(n17997), .ZN(n17994) );
  AND2_X1 U17834 ( .A1(n17999), .A2(n18000), .ZN(n17997) );
  OR2_X1 U17835 ( .A1(n18001), .A2(n18002), .ZN(n18000) );
  INV_X1 U17836 ( .A(n18003), .ZN(n18002) );
  OR2_X1 U17837 ( .A1(n18003), .A2(n18004), .ZN(n17999) );
  INV_X1 U17838 ( .A(n18001), .ZN(n18004) );
  OR2_X1 U17839 ( .A1(n15423), .A2(n14856), .ZN(n17609) );
  OR2_X1 U17840 ( .A1(n18005), .A2(n18006), .ZN(n17606) );
  INV_X1 U17841 ( .A(n18007), .ZN(n18006) );
  OR2_X1 U17842 ( .A1(n18008), .A2(n18009), .ZN(n18007) );
  AND2_X1 U17843 ( .A1(n18009), .A2(n18008), .ZN(n18005) );
  AND2_X1 U17844 ( .A1(n18010), .A2(n18011), .ZN(n18008) );
  OR2_X1 U17845 ( .A1(n18012), .A2(n18013), .ZN(n18011) );
  INV_X1 U17846 ( .A(n18014), .ZN(n18013) );
  OR2_X1 U17847 ( .A1(n18014), .A2(n18015), .ZN(n18010) );
  INV_X1 U17848 ( .A(n18012), .ZN(n18015) );
  OR2_X1 U17849 ( .A1(n15457), .A2(n14856), .ZN(n17620) );
  OR2_X1 U17850 ( .A1(n18016), .A2(n18017), .ZN(n17617) );
  INV_X1 U17851 ( .A(n18018), .ZN(n18017) );
  OR2_X1 U17852 ( .A1(n18019), .A2(n18020), .ZN(n18018) );
  AND2_X1 U17853 ( .A1(n18020), .A2(n18019), .ZN(n18016) );
  AND2_X1 U17854 ( .A1(n18021), .A2(n18022), .ZN(n18019) );
  OR2_X1 U17855 ( .A1(n18023), .A2(n18024), .ZN(n18022) );
  INV_X1 U17856 ( .A(n18025), .ZN(n18024) );
  OR2_X1 U17857 ( .A1(n18025), .A2(n18026), .ZN(n18021) );
  INV_X1 U17858 ( .A(n18023), .ZN(n18026) );
  OR2_X1 U17859 ( .A1(n15491), .A2(n14856), .ZN(n17631) );
  OR2_X1 U17860 ( .A1(n18027), .A2(n18028), .ZN(n17628) );
  INV_X1 U17861 ( .A(n18029), .ZN(n18028) );
  OR2_X1 U17862 ( .A1(n18030), .A2(n18031), .ZN(n18029) );
  AND2_X1 U17863 ( .A1(n18031), .A2(n18030), .ZN(n18027) );
  AND2_X1 U17864 ( .A1(n18032), .A2(n18033), .ZN(n18030) );
  OR2_X1 U17865 ( .A1(n18034), .A2(n18035), .ZN(n18033) );
  INV_X1 U17866 ( .A(n18036), .ZN(n18035) );
  OR2_X1 U17867 ( .A1(n18036), .A2(n18037), .ZN(n18032) );
  INV_X1 U17868 ( .A(n18034), .ZN(n18037) );
  OR2_X1 U17869 ( .A1(n15525), .A2(n14856), .ZN(n17642) );
  OR2_X1 U17870 ( .A1(n18038), .A2(n18039), .ZN(n17639) );
  INV_X1 U17871 ( .A(n18040), .ZN(n18039) );
  OR2_X1 U17872 ( .A1(n18041), .A2(n18042), .ZN(n18040) );
  AND2_X1 U17873 ( .A1(n18042), .A2(n18041), .ZN(n18038) );
  AND2_X1 U17874 ( .A1(n18043), .A2(n18044), .ZN(n18041) );
  OR2_X1 U17875 ( .A1(n18045), .A2(n18046), .ZN(n18044) );
  INV_X1 U17876 ( .A(n18047), .ZN(n18046) );
  OR2_X1 U17877 ( .A1(n18047), .A2(n18048), .ZN(n18043) );
  INV_X1 U17878 ( .A(n18045), .ZN(n18048) );
  OR2_X1 U17879 ( .A1(n15559), .A2(n14856), .ZN(n17653) );
  OR2_X1 U17880 ( .A1(n18049), .A2(n18050), .ZN(n17650) );
  INV_X1 U17881 ( .A(n18051), .ZN(n18050) );
  OR2_X1 U17882 ( .A1(n18052), .A2(n18053), .ZN(n18051) );
  AND2_X1 U17883 ( .A1(n18053), .A2(n18052), .ZN(n18049) );
  AND2_X1 U17884 ( .A1(n18054), .A2(n18055), .ZN(n18052) );
  OR2_X1 U17885 ( .A1(n18056), .A2(n18057), .ZN(n18055) );
  INV_X1 U17886 ( .A(n18058), .ZN(n18057) );
  OR2_X1 U17887 ( .A1(n18058), .A2(n18059), .ZN(n18054) );
  INV_X1 U17888 ( .A(n18056), .ZN(n18059) );
  OR2_X1 U17889 ( .A1(n15593), .A2(n14856), .ZN(n17664) );
  OR2_X1 U17890 ( .A1(n18060), .A2(n18061), .ZN(n17661) );
  INV_X1 U17891 ( .A(n18062), .ZN(n18061) );
  OR2_X1 U17892 ( .A1(n18063), .A2(n18064), .ZN(n18062) );
  AND2_X1 U17893 ( .A1(n18064), .A2(n18063), .ZN(n18060) );
  AND2_X1 U17894 ( .A1(n18065), .A2(n18066), .ZN(n18063) );
  OR2_X1 U17895 ( .A1(n18067), .A2(n18068), .ZN(n18066) );
  INV_X1 U17896 ( .A(n18069), .ZN(n18068) );
  OR2_X1 U17897 ( .A1(n18069), .A2(n18070), .ZN(n18065) );
  INV_X1 U17898 ( .A(n18067), .ZN(n18070) );
  OR2_X1 U17899 ( .A1(n15638), .A2(n14856), .ZN(n17675) );
  OR2_X1 U17900 ( .A1(n18071), .A2(n18072), .ZN(n17672) );
  INV_X1 U17901 ( .A(n18073), .ZN(n18072) );
  OR2_X1 U17902 ( .A1(n18074), .A2(n18075), .ZN(n18073) );
  AND2_X1 U17903 ( .A1(n18075), .A2(n18074), .ZN(n18071) );
  AND2_X1 U17904 ( .A1(n18076), .A2(n18077), .ZN(n18074) );
  OR2_X1 U17905 ( .A1(n18078), .A2(n18079), .ZN(n18077) );
  INV_X1 U17906 ( .A(n18080), .ZN(n18079) );
  OR2_X1 U17907 ( .A1(n18080), .A2(n18081), .ZN(n18076) );
  INV_X1 U17908 ( .A(n18078), .ZN(n18081) );
  OR2_X1 U17909 ( .A1(n15672), .A2(n14856), .ZN(n17686) );
  OR2_X1 U17910 ( .A1(n18082), .A2(n18083), .ZN(n17683) );
  INV_X1 U17911 ( .A(n18084), .ZN(n18083) );
  OR2_X1 U17912 ( .A1(n18085), .A2(n18086), .ZN(n18084) );
  AND2_X1 U17913 ( .A1(n18086), .A2(n18085), .ZN(n18082) );
  AND2_X1 U17914 ( .A1(n18087), .A2(n18088), .ZN(n18085) );
  OR2_X1 U17915 ( .A1(n18089), .A2(n18090), .ZN(n18088) );
  INV_X1 U17916 ( .A(n18091), .ZN(n18090) );
  OR2_X1 U17917 ( .A1(n18091), .A2(n18092), .ZN(n18087) );
  INV_X1 U17918 ( .A(n18089), .ZN(n18092) );
  OR2_X1 U17919 ( .A1(n15706), .A2(n14856), .ZN(n17697) );
  OR2_X1 U17920 ( .A1(n18093), .A2(n18094), .ZN(n17694) );
  INV_X1 U17921 ( .A(n18095), .ZN(n18094) );
  OR2_X1 U17922 ( .A1(n18096), .A2(n18097), .ZN(n18095) );
  AND2_X1 U17923 ( .A1(n18097), .A2(n18096), .ZN(n18093) );
  AND2_X1 U17924 ( .A1(n18098), .A2(n18099), .ZN(n18096) );
  OR2_X1 U17925 ( .A1(n18100), .A2(n18101), .ZN(n18099) );
  INV_X1 U17926 ( .A(n18102), .ZN(n18101) );
  OR2_X1 U17927 ( .A1(n18102), .A2(n18103), .ZN(n18098) );
  INV_X1 U17928 ( .A(n18100), .ZN(n18103) );
  OR2_X1 U17929 ( .A1(n15740), .A2(n14856), .ZN(n17708) );
  OR2_X1 U17930 ( .A1(n18104), .A2(n18105), .ZN(n17705) );
  INV_X1 U17931 ( .A(n18106), .ZN(n18105) );
  OR2_X1 U17932 ( .A1(n18107), .A2(n18108), .ZN(n18106) );
  AND2_X1 U17933 ( .A1(n18108), .A2(n18107), .ZN(n18104) );
  AND2_X1 U17934 ( .A1(n18109), .A2(n18110), .ZN(n18107) );
  OR2_X1 U17935 ( .A1(n18111), .A2(n18112), .ZN(n18110) );
  INV_X1 U17936 ( .A(n18113), .ZN(n18112) );
  OR2_X1 U17937 ( .A1(n18113), .A2(n18114), .ZN(n18109) );
  INV_X1 U17938 ( .A(n18111), .ZN(n18114) );
  OR2_X1 U17939 ( .A1(n15774), .A2(n14856), .ZN(n17719) );
  OR2_X1 U17940 ( .A1(n18115), .A2(n18116), .ZN(n17716) );
  INV_X1 U17941 ( .A(n18117), .ZN(n18116) );
  OR2_X1 U17942 ( .A1(n18118), .A2(n18119), .ZN(n18117) );
  AND2_X1 U17943 ( .A1(n18119), .A2(n18118), .ZN(n18115) );
  AND2_X1 U17944 ( .A1(n18120), .A2(n18121), .ZN(n18118) );
  OR2_X1 U17945 ( .A1(n18122), .A2(n18123), .ZN(n18121) );
  INV_X1 U17946 ( .A(n18124), .ZN(n18123) );
  OR2_X1 U17947 ( .A1(n18124), .A2(n18125), .ZN(n18120) );
  INV_X1 U17948 ( .A(n18122), .ZN(n18125) );
  OR2_X1 U17949 ( .A1(n15808), .A2(n14856), .ZN(n17730) );
  OR2_X1 U17950 ( .A1(n18126), .A2(n18127), .ZN(n17727) );
  INV_X1 U17951 ( .A(n18128), .ZN(n18127) );
  OR2_X1 U17952 ( .A1(n18129), .A2(n18130), .ZN(n18128) );
  AND2_X1 U17953 ( .A1(n18130), .A2(n18129), .ZN(n18126) );
  AND2_X1 U17954 ( .A1(n18131), .A2(n18132), .ZN(n18129) );
  OR2_X1 U17955 ( .A1(n18133), .A2(n18134), .ZN(n18132) );
  INV_X1 U17956 ( .A(n18135), .ZN(n18134) );
  OR2_X1 U17957 ( .A1(n18135), .A2(n18136), .ZN(n18131) );
  INV_X1 U17958 ( .A(n18133), .ZN(n18136) );
  OR2_X1 U17959 ( .A1(n15842), .A2(n14856), .ZN(n17741) );
  OR2_X1 U17960 ( .A1(n18137), .A2(n18138), .ZN(n17738) );
  INV_X1 U17961 ( .A(n18139), .ZN(n18138) );
  OR2_X1 U17962 ( .A1(n18140), .A2(n18141), .ZN(n18139) );
  AND2_X1 U17963 ( .A1(n18141), .A2(n18140), .ZN(n18137) );
  AND2_X1 U17964 ( .A1(n18142), .A2(n18143), .ZN(n18140) );
  OR2_X1 U17965 ( .A1(n18144), .A2(n18145), .ZN(n18143) );
  INV_X1 U17966 ( .A(n18146), .ZN(n18145) );
  OR2_X1 U17967 ( .A1(n18146), .A2(n18147), .ZN(n18142) );
  INV_X1 U17968 ( .A(n18144), .ZN(n18147) );
  OR2_X1 U17969 ( .A1(n16512), .A2(n14856), .ZN(n17315) );
  INV_X1 U17970 ( .A(b_29_), .ZN(n14856) );
  INV_X1 U17971 ( .A(n17317), .ZN(n17311) );
  AND2_X1 U17972 ( .A1(n18148), .A2(n18149), .ZN(n17317) );
  OR2_X1 U17973 ( .A1(n18150), .A2(n18151), .ZN(n18149) );
  INV_X1 U17974 ( .A(n18152), .ZN(n18148) );
  AND2_X1 U17975 ( .A1(n18151), .A2(n18150), .ZN(n18152) );
  AND2_X1 U17976 ( .A1(n18153), .A2(n18154), .ZN(n18150) );
  INV_X1 U17977 ( .A(n18155), .ZN(n18154) );
  AND2_X1 U17978 ( .A1(n18156), .A2(n18157), .ZN(n18155) );
  OR2_X1 U17979 ( .A1(n18157), .A2(n18156), .ZN(n18153) );
  INV_X1 U17980 ( .A(n18158), .ZN(n18156) );
  INV_X1 U17981 ( .A(n16886), .ZN(n16877) );
  AND2_X1 U17982 ( .A1(n18159), .A2(n18160), .ZN(n16886) );
  INV_X1 U17983 ( .A(n18161), .ZN(n18160) );
  AND2_X1 U17984 ( .A1(n18162), .A2(n18163), .ZN(n18161) );
  OR2_X1 U17985 ( .A1(n18163), .A2(n18162), .ZN(n18159) );
  OR2_X1 U17986 ( .A1(n18164), .A2(n18165), .ZN(n18162) );
  AND2_X1 U17987 ( .A1(n18166), .A2(n18167), .ZN(n18165) );
  INV_X1 U17988 ( .A(n18168), .ZN(n18166) );
  AND2_X1 U17989 ( .A1(n18169), .A2(n18168), .ZN(n18164) );
  INV_X1 U17990 ( .A(n18167), .ZN(n18169) );
  OR2_X1 U17991 ( .A1(n18170), .A2(n18171), .ZN(n16875) );
  AND2_X1 U17992 ( .A1(n18172), .A2(n18173), .ZN(n18171) );
  AND2_X1 U17993 ( .A1(n18174), .A2(n18175), .ZN(n18170) );
  AND2_X1 U17994 ( .A1(n16873), .A2(n16872), .ZN(n16020) );
  AND2_X1 U17995 ( .A1(n18172), .A2(n18175), .ZN(n16872) );
  INV_X1 U17996 ( .A(n18173), .ZN(n18175) );
  OR2_X1 U17997 ( .A1(n18176), .A2(n18177), .ZN(n18173) );
  AND2_X1 U17998 ( .A1(n18168), .A2(n18167), .ZN(n18177) );
  AND2_X1 U17999 ( .A1(n18163), .A2(n18178), .ZN(n18176) );
  OR2_X1 U18000 ( .A1(n18168), .A2(n18167), .ZN(n18178) );
  OR2_X1 U18001 ( .A1(n18179), .A2(n18180), .ZN(n18167) );
  AND2_X1 U18002 ( .A1(n18158), .A2(n18157), .ZN(n18180) );
  AND2_X1 U18003 ( .A1(n18151), .A2(n18181), .ZN(n18179) );
  OR2_X1 U18004 ( .A1(n18158), .A2(n18157), .ZN(n18181) );
  OR2_X1 U18005 ( .A1(n18182), .A2(n18183), .ZN(n18157) );
  AND2_X1 U18006 ( .A1(n18144), .A2(n18146), .ZN(n18183) );
  AND2_X1 U18007 ( .A1(n18141), .A2(n18184), .ZN(n18182) );
  OR2_X1 U18008 ( .A1(n18144), .A2(n18146), .ZN(n18184) );
  OR2_X1 U18009 ( .A1(n18185), .A2(n18186), .ZN(n18146) );
  AND2_X1 U18010 ( .A1(n18133), .A2(n18135), .ZN(n18186) );
  AND2_X1 U18011 ( .A1(n18130), .A2(n18187), .ZN(n18185) );
  OR2_X1 U18012 ( .A1(n18133), .A2(n18135), .ZN(n18187) );
  OR2_X1 U18013 ( .A1(n18188), .A2(n18189), .ZN(n18135) );
  AND2_X1 U18014 ( .A1(n18122), .A2(n18124), .ZN(n18189) );
  AND2_X1 U18015 ( .A1(n18119), .A2(n18190), .ZN(n18188) );
  OR2_X1 U18016 ( .A1(n18122), .A2(n18124), .ZN(n18190) );
  OR2_X1 U18017 ( .A1(n18191), .A2(n18192), .ZN(n18124) );
  AND2_X1 U18018 ( .A1(n18111), .A2(n18113), .ZN(n18192) );
  AND2_X1 U18019 ( .A1(n18108), .A2(n18193), .ZN(n18191) );
  OR2_X1 U18020 ( .A1(n18111), .A2(n18113), .ZN(n18193) );
  OR2_X1 U18021 ( .A1(n18194), .A2(n18195), .ZN(n18113) );
  AND2_X1 U18022 ( .A1(n18100), .A2(n18102), .ZN(n18195) );
  AND2_X1 U18023 ( .A1(n18097), .A2(n18196), .ZN(n18194) );
  OR2_X1 U18024 ( .A1(n18100), .A2(n18102), .ZN(n18196) );
  OR2_X1 U18025 ( .A1(n18197), .A2(n18198), .ZN(n18102) );
  AND2_X1 U18026 ( .A1(n18089), .A2(n18091), .ZN(n18198) );
  AND2_X1 U18027 ( .A1(n18086), .A2(n18199), .ZN(n18197) );
  OR2_X1 U18028 ( .A1(n18089), .A2(n18091), .ZN(n18199) );
  OR2_X1 U18029 ( .A1(n18200), .A2(n18201), .ZN(n18091) );
  AND2_X1 U18030 ( .A1(n18078), .A2(n18080), .ZN(n18201) );
  AND2_X1 U18031 ( .A1(n18075), .A2(n18202), .ZN(n18200) );
  OR2_X1 U18032 ( .A1(n18078), .A2(n18080), .ZN(n18202) );
  OR2_X1 U18033 ( .A1(n18203), .A2(n18204), .ZN(n18080) );
  AND2_X1 U18034 ( .A1(n18067), .A2(n18069), .ZN(n18204) );
  AND2_X1 U18035 ( .A1(n18064), .A2(n18205), .ZN(n18203) );
  OR2_X1 U18036 ( .A1(n18067), .A2(n18069), .ZN(n18205) );
  OR2_X1 U18037 ( .A1(n18206), .A2(n18207), .ZN(n18069) );
  AND2_X1 U18038 ( .A1(n18056), .A2(n18058), .ZN(n18207) );
  AND2_X1 U18039 ( .A1(n18053), .A2(n18208), .ZN(n18206) );
  OR2_X1 U18040 ( .A1(n18056), .A2(n18058), .ZN(n18208) );
  OR2_X1 U18041 ( .A1(n18209), .A2(n18210), .ZN(n18058) );
  AND2_X1 U18042 ( .A1(n18045), .A2(n18047), .ZN(n18210) );
  AND2_X1 U18043 ( .A1(n18042), .A2(n18211), .ZN(n18209) );
  OR2_X1 U18044 ( .A1(n18045), .A2(n18047), .ZN(n18211) );
  OR2_X1 U18045 ( .A1(n18212), .A2(n18213), .ZN(n18047) );
  AND2_X1 U18046 ( .A1(n18034), .A2(n18036), .ZN(n18213) );
  AND2_X1 U18047 ( .A1(n18031), .A2(n18214), .ZN(n18212) );
  OR2_X1 U18048 ( .A1(n18034), .A2(n18036), .ZN(n18214) );
  OR2_X1 U18049 ( .A1(n18215), .A2(n18216), .ZN(n18036) );
  AND2_X1 U18050 ( .A1(n18023), .A2(n18025), .ZN(n18216) );
  AND2_X1 U18051 ( .A1(n18020), .A2(n18217), .ZN(n18215) );
  OR2_X1 U18052 ( .A1(n18023), .A2(n18025), .ZN(n18217) );
  OR2_X1 U18053 ( .A1(n18218), .A2(n18219), .ZN(n18025) );
  AND2_X1 U18054 ( .A1(n18012), .A2(n18014), .ZN(n18219) );
  AND2_X1 U18055 ( .A1(n18009), .A2(n18220), .ZN(n18218) );
  OR2_X1 U18056 ( .A1(n18012), .A2(n18014), .ZN(n18220) );
  OR2_X1 U18057 ( .A1(n18221), .A2(n18222), .ZN(n18014) );
  AND2_X1 U18058 ( .A1(n18001), .A2(n18003), .ZN(n18222) );
  AND2_X1 U18059 ( .A1(n17998), .A2(n18223), .ZN(n18221) );
  OR2_X1 U18060 ( .A1(n18001), .A2(n18003), .ZN(n18223) );
  OR2_X1 U18061 ( .A1(n18224), .A2(n18225), .ZN(n18003) );
  AND2_X1 U18062 ( .A1(n17990), .A2(n17992), .ZN(n18225) );
  AND2_X1 U18063 ( .A1(n17987), .A2(n18226), .ZN(n18224) );
  OR2_X1 U18064 ( .A1(n17990), .A2(n17992), .ZN(n18226) );
  OR2_X1 U18065 ( .A1(n18227), .A2(n18228), .ZN(n17992) );
  AND2_X1 U18066 ( .A1(n17979), .A2(n17981), .ZN(n18228) );
  AND2_X1 U18067 ( .A1(n17976), .A2(n18229), .ZN(n18227) );
  OR2_X1 U18068 ( .A1(n17979), .A2(n17981), .ZN(n18229) );
  OR2_X1 U18069 ( .A1(n18230), .A2(n18231), .ZN(n17981) );
  AND2_X1 U18070 ( .A1(n17968), .A2(n17970), .ZN(n18231) );
  AND2_X1 U18071 ( .A1(n17965), .A2(n18232), .ZN(n18230) );
  OR2_X1 U18072 ( .A1(n17968), .A2(n17970), .ZN(n18232) );
  OR2_X1 U18073 ( .A1(n18233), .A2(n18234), .ZN(n17970) );
  AND2_X1 U18074 ( .A1(n17957), .A2(n17959), .ZN(n18234) );
  AND2_X1 U18075 ( .A1(n17954), .A2(n18235), .ZN(n18233) );
  OR2_X1 U18076 ( .A1(n17957), .A2(n17959), .ZN(n18235) );
  OR2_X1 U18077 ( .A1(n18236), .A2(n18237), .ZN(n17959) );
  AND2_X1 U18078 ( .A1(n17946), .A2(n17948), .ZN(n18237) );
  AND2_X1 U18079 ( .A1(n17943), .A2(n18238), .ZN(n18236) );
  OR2_X1 U18080 ( .A1(n17946), .A2(n17948), .ZN(n18238) );
  OR2_X1 U18081 ( .A1(n18239), .A2(n18240), .ZN(n17948) );
  AND2_X1 U18082 ( .A1(n17935), .A2(n17937), .ZN(n18240) );
  AND2_X1 U18083 ( .A1(n17932), .A2(n18241), .ZN(n18239) );
  OR2_X1 U18084 ( .A1(n17935), .A2(n17937), .ZN(n18241) );
  OR2_X1 U18085 ( .A1(n18242), .A2(n18243), .ZN(n17937) );
  AND2_X1 U18086 ( .A1(n17924), .A2(n17926), .ZN(n18243) );
  AND2_X1 U18087 ( .A1(n17921), .A2(n18244), .ZN(n18242) );
  OR2_X1 U18088 ( .A1(n17924), .A2(n17926), .ZN(n18244) );
  OR2_X1 U18089 ( .A1(n18245), .A2(n18246), .ZN(n17926) );
  AND2_X1 U18090 ( .A1(n17913), .A2(n17915), .ZN(n18246) );
  AND2_X1 U18091 ( .A1(n17910), .A2(n18247), .ZN(n18245) );
  OR2_X1 U18092 ( .A1(n17913), .A2(n17915), .ZN(n18247) );
  OR2_X1 U18093 ( .A1(n18248), .A2(n18249), .ZN(n17915) );
  AND2_X1 U18094 ( .A1(n17902), .A2(n17904), .ZN(n18249) );
  AND2_X1 U18095 ( .A1(n17899), .A2(n18250), .ZN(n18248) );
  OR2_X1 U18096 ( .A1(n17902), .A2(n17904), .ZN(n18250) );
  OR2_X1 U18097 ( .A1(n18251), .A2(n18252), .ZN(n17904) );
  AND2_X1 U18098 ( .A1(n17891), .A2(n17893), .ZN(n18252) );
  AND2_X1 U18099 ( .A1(n17888), .A2(n18253), .ZN(n18251) );
  OR2_X1 U18100 ( .A1(n17891), .A2(n17893), .ZN(n18253) );
  OR2_X1 U18101 ( .A1(n18254), .A2(n18255), .ZN(n17893) );
  AND2_X1 U18102 ( .A1(n17880), .A2(n17882), .ZN(n18255) );
  AND2_X1 U18103 ( .A1(n17877), .A2(n18256), .ZN(n18254) );
  OR2_X1 U18104 ( .A1(n17880), .A2(n17882), .ZN(n18256) );
  OR2_X1 U18105 ( .A1(n18257), .A2(n18258), .ZN(n17882) );
  AND2_X1 U18106 ( .A1(n17869), .A2(n17871), .ZN(n18258) );
  AND2_X1 U18107 ( .A1(n17866), .A2(n18259), .ZN(n18257) );
  OR2_X1 U18108 ( .A1(n17869), .A2(n17871), .ZN(n18259) );
  OR2_X1 U18109 ( .A1(n18260), .A2(n18261), .ZN(n17871) );
  AND2_X1 U18110 ( .A1(n15951), .A2(n17860), .ZN(n18261) );
  AND2_X1 U18111 ( .A1(n17856), .A2(n18262), .ZN(n18260) );
  OR2_X1 U18112 ( .A1(n15951), .A2(n17860), .ZN(n18262) );
  OR2_X1 U18113 ( .A1(n18263), .A2(n18264), .ZN(n17860) );
  AND2_X1 U18114 ( .A1(n17844), .A2(n17849), .ZN(n18264) );
  AND2_X1 U18115 ( .A1(n17848), .A2(n18265), .ZN(n18263) );
  OR2_X1 U18116 ( .A1(n17844), .A2(n17849), .ZN(n18265) );
  INV_X1 U18117 ( .A(n17850), .ZN(n17849) );
  AND3_X1 U18118 ( .A1(b_28_), .A2(b_27_), .A3(n15957), .ZN(n17850) );
  OR2_X1 U18119 ( .A1(n14857), .A2(n14890), .ZN(n17844) );
  INV_X1 U18120 ( .A(n17851), .ZN(n17848) );
  OR2_X1 U18121 ( .A1(n18266), .A2(n18267), .ZN(n17851) );
  AND2_X1 U18122 ( .A1(b_27_), .A2(n18268), .ZN(n18267) );
  OR2_X1 U18123 ( .A1(n18269), .A2(n16981), .ZN(n18268) );
  AND2_X1 U18124 ( .A1(a_30_), .A2(n14969), .ZN(n18269) );
  AND2_X1 U18125 ( .A1(b_26_), .A2(n18270), .ZN(n18266) );
  OR2_X1 U18126 ( .A1(n18271), .A2(n14817), .ZN(n18270) );
  AND2_X1 U18127 ( .A1(a_31_), .A2(n14935), .ZN(n18271) );
  OR2_X1 U18128 ( .A1(n14891), .A2(n14890), .ZN(n15951) );
  OR2_X1 U18129 ( .A1(n18272), .A2(n18273), .ZN(n17856) );
  AND2_X1 U18130 ( .A1(n18274), .A2(n18275), .ZN(n18273) );
  INV_X1 U18131 ( .A(n18276), .ZN(n18272) );
  OR2_X1 U18132 ( .A1(n18274), .A2(n18275), .ZN(n18276) );
  OR2_X1 U18133 ( .A1(n18277), .A2(n18278), .ZN(n18274) );
  AND2_X1 U18134 ( .A1(n18279), .A2(n18280), .ZN(n18278) );
  AND2_X1 U18135 ( .A1(n18281), .A2(n18282), .ZN(n18277) );
  OR2_X1 U18136 ( .A1(n14936), .A2(n14890), .ZN(n17869) );
  OR2_X1 U18137 ( .A1(n18283), .A2(n18284), .ZN(n17866) );
  INV_X1 U18138 ( .A(n18285), .ZN(n18284) );
  OR2_X1 U18139 ( .A1(n18286), .A2(n18287), .ZN(n18285) );
  AND2_X1 U18140 ( .A1(n18287), .A2(n18286), .ZN(n18283) );
  AND2_X1 U18141 ( .A1(n18288), .A2(n18289), .ZN(n18286) );
  OR2_X1 U18142 ( .A1(n18290), .A2(n18291), .ZN(n18289) );
  INV_X1 U18143 ( .A(n18292), .ZN(n18291) );
  OR2_X1 U18144 ( .A1(n18292), .A2(n18293), .ZN(n18288) );
  INV_X1 U18145 ( .A(n18290), .ZN(n18293) );
  OR2_X1 U18146 ( .A1(n14970), .A2(n14890), .ZN(n17880) );
  OR2_X1 U18147 ( .A1(n18294), .A2(n18295), .ZN(n17877) );
  INV_X1 U18148 ( .A(n18296), .ZN(n18295) );
  OR2_X1 U18149 ( .A1(n18297), .A2(n18298), .ZN(n18296) );
  AND2_X1 U18150 ( .A1(n18298), .A2(n18297), .ZN(n18294) );
  AND2_X1 U18151 ( .A1(n18299), .A2(n18300), .ZN(n18297) );
  OR2_X1 U18152 ( .A1(n15948), .A2(n18301), .ZN(n18300) );
  INV_X1 U18153 ( .A(n18302), .ZN(n18301) );
  OR2_X1 U18154 ( .A1(n18302), .A2(n18303), .ZN(n18299) );
  INV_X1 U18155 ( .A(n15948), .ZN(n18303) );
  OR2_X1 U18156 ( .A1(n15004), .A2(n14890), .ZN(n17891) );
  OR2_X1 U18157 ( .A1(n18304), .A2(n18305), .ZN(n17888) );
  INV_X1 U18158 ( .A(n18306), .ZN(n18305) );
  OR2_X1 U18159 ( .A1(n18307), .A2(n18308), .ZN(n18306) );
  AND2_X1 U18160 ( .A1(n18308), .A2(n18307), .ZN(n18304) );
  AND2_X1 U18161 ( .A1(n18309), .A2(n18310), .ZN(n18307) );
  OR2_X1 U18162 ( .A1(n18311), .A2(n18312), .ZN(n18310) );
  INV_X1 U18163 ( .A(n18313), .ZN(n18312) );
  OR2_X1 U18164 ( .A1(n18313), .A2(n18314), .ZN(n18309) );
  INV_X1 U18165 ( .A(n18311), .ZN(n18314) );
  OR2_X1 U18166 ( .A1(n15038), .A2(n14890), .ZN(n17902) );
  OR2_X1 U18167 ( .A1(n18315), .A2(n18316), .ZN(n17899) );
  INV_X1 U18168 ( .A(n18317), .ZN(n18316) );
  OR2_X1 U18169 ( .A1(n18318), .A2(n18319), .ZN(n18317) );
  AND2_X1 U18170 ( .A1(n18319), .A2(n18318), .ZN(n18315) );
  AND2_X1 U18171 ( .A1(n18320), .A2(n18321), .ZN(n18318) );
  OR2_X1 U18172 ( .A1(n18322), .A2(n18323), .ZN(n18321) );
  INV_X1 U18173 ( .A(n18324), .ZN(n18323) );
  OR2_X1 U18174 ( .A1(n18324), .A2(n18325), .ZN(n18320) );
  INV_X1 U18175 ( .A(n18322), .ZN(n18325) );
  OR2_X1 U18176 ( .A1(n15072), .A2(n14890), .ZN(n17913) );
  OR2_X1 U18177 ( .A1(n18326), .A2(n18327), .ZN(n17910) );
  INV_X1 U18178 ( .A(n18328), .ZN(n18327) );
  OR2_X1 U18179 ( .A1(n18329), .A2(n18330), .ZN(n18328) );
  AND2_X1 U18180 ( .A1(n18330), .A2(n18329), .ZN(n18326) );
  AND2_X1 U18181 ( .A1(n18331), .A2(n18332), .ZN(n18329) );
  OR2_X1 U18182 ( .A1(n18333), .A2(n18334), .ZN(n18332) );
  INV_X1 U18183 ( .A(n18335), .ZN(n18334) );
  OR2_X1 U18184 ( .A1(n18335), .A2(n18336), .ZN(n18331) );
  INV_X1 U18185 ( .A(n18333), .ZN(n18336) );
  OR2_X1 U18186 ( .A1(n15106), .A2(n14890), .ZN(n17924) );
  OR2_X1 U18187 ( .A1(n18337), .A2(n18338), .ZN(n17921) );
  INV_X1 U18188 ( .A(n18339), .ZN(n18338) );
  OR2_X1 U18189 ( .A1(n18340), .A2(n18341), .ZN(n18339) );
  AND2_X1 U18190 ( .A1(n18341), .A2(n18340), .ZN(n18337) );
  AND2_X1 U18191 ( .A1(n18342), .A2(n18343), .ZN(n18340) );
  OR2_X1 U18192 ( .A1(n18344), .A2(n18345), .ZN(n18343) );
  INV_X1 U18193 ( .A(n18346), .ZN(n18345) );
  OR2_X1 U18194 ( .A1(n18346), .A2(n18347), .ZN(n18342) );
  INV_X1 U18195 ( .A(n18344), .ZN(n18347) );
  OR2_X1 U18196 ( .A1(n15140), .A2(n14890), .ZN(n17935) );
  OR2_X1 U18197 ( .A1(n18348), .A2(n18349), .ZN(n17932) );
  INV_X1 U18198 ( .A(n18350), .ZN(n18349) );
  OR2_X1 U18199 ( .A1(n18351), .A2(n18352), .ZN(n18350) );
  AND2_X1 U18200 ( .A1(n18352), .A2(n18351), .ZN(n18348) );
  AND2_X1 U18201 ( .A1(n18353), .A2(n18354), .ZN(n18351) );
  OR2_X1 U18202 ( .A1(n18355), .A2(n18356), .ZN(n18354) );
  INV_X1 U18203 ( .A(n18357), .ZN(n18356) );
  OR2_X1 U18204 ( .A1(n18357), .A2(n18358), .ZN(n18353) );
  INV_X1 U18205 ( .A(n18355), .ZN(n18358) );
  OR2_X1 U18206 ( .A1(n15174), .A2(n14890), .ZN(n17946) );
  OR2_X1 U18207 ( .A1(n18359), .A2(n18360), .ZN(n17943) );
  INV_X1 U18208 ( .A(n18361), .ZN(n18360) );
  OR2_X1 U18209 ( .A1(n18362), .A2(n18363), .ZN(n18361) );
  AND2_X1 U18210 ( .A1(n18363), .A2(n18362), .ZN(n18359) );
  AND2_X1 U18211 ( .A1(n18364), .A2(n18365), .ZN(n18362) );
  OR2_X1 U18212 ( .A1(n18366), .A2(n18367), .ZN(n18365) );
  INV_X1 U18213 ( .A(n18368), .ZN(n18367) );
  OR2_X1 U18214 ( .A1(n18368), .A2(n18369), .ZN(n18364) );
  INV_X1 U18215 ( .A(n18366), .ZN(n18369) );
  OR2_X1 U18216 ( .A1(n15208), .A2(n14890), .ZN(n17957) );
  OR2_X1 U18217 ( .A1(n18370), .A2(n18371), .ZN(n17954) );
  INV_X1 U18218 ( .A(n18372), .ZN(n18371) );
  OR2_X1 U18219 ( .A1(n18373), .A2(n18374), .ZN(n18372) );
  AND2_X1 U18220 ( .A1(n18374), .A2(n18373), .ZN(n18370) );
  AND2_X1 U18221 ( .A1(n18375), .A2(n18376), .ZN(n18373) );
  OR2_X1 U18222 ( .A1(n18377), .A2(n18378), .ZN(n18376) );
  INV_X1 U18223 ( .A(n18379), .ZN(n18378) );
  OR2_X1 U18224 ( .A1(n18379), .A2(n18380), .ZN(n18375) );
  INV_X1 U18225 ( .A(n18377), .ZN(n18380) );
  OR2_X1 U18226 ( .A1(n15242), .A2(n14890), .ZN(n17968) );
  OR2_X1 U18227 ( .A1(n18381), .A2(n18382), .ZN(n17965) );
  INV_X1 U18228 ( .A(n18383), .ZN(n18382) );
  OR2_X1 U18229 ( .A1(n18384), .A2(n18385), .ZN(n18383) );
  AND2_X1 U18230 ( .A1(n18385), .A2(n18384), .ZN(n18381) );
  AND2_X1 U18231 ( .A1(n18386), .A2(n18387), .ZN(n18384) );
  OR2_X1 U18232 ( .A1(n18388), .A2(n18389), .ZN(n18387) );
  INV_X1 U18233 ( .A(n18390), .ZN(n18389) );
  OR2_X1 U18234 ( .A1(n18390), .A2(n18391), .ZN(n18386) );
  INV_X1 U18235 ( .A(n18388), .ZN(n18391) );
  OR2_X1 U18236 ( .A1(n15287), .A2(n14890), .ZN(n17979) );
  OR2_X1 U18237 ( .A1(n18392), .A2(n18393), .ZN(n17976) );
  INV_X1 U18238 ( .A(n18394), .ZN(n18393) );
  OR2_X1 U18239 ( .A1(n18395), .A2(n18396), .ZN(n18394) );
  AND2_X1 U18240 ( .A1(n18396), .A2(n18395), .ZN(n18392) );
  AND2_X1 U18241 ( .A1(n18397), .A2(n18398), .ZN(n18395) );
  OR2_X1 U18242 ( .A1(n18399), .A2(n18400), .ZN(n18398) );
  INV_X1 U18243 ( .A(n18401), .ZN(n18400) );
  OR2_X1 U18244 ( .A1(n18401), .A2(n18402), .ZN(n18397) );
  INV_X1 U18245 ( .A(n18399), .ZN(n18402) );
  OR2_X1 U18246 ( .A1(n15321), .A2(n14890), .ZN(n17990) );
  OR2_X1 U18247 ( .A1(n18403), .A2(n18404), .ZN(n17987) );
  INV_X1 U18248 ( .A(n18405), .ZN(n18404) );
  OR2_X1 U18249 ( .A1(n18406), .A2(n18407), .ZN(n18405) );
  AND2_X1 U18250 ( .A1(n18407), .A2(n18406), .ZN(n18403) );
  AND2_X1 U18251 ( .A1(n18408), .A2(n18409), .ZN(n18406) );
  OR2_X1 U18252 ( .A1(n18410), .A2(n18411), .ZN(n18409) );
  INV_X1 U18253 ( .A(n18412), .ZN(n18411) );
  OR2_X1 U18254 ( .A1(n18412), .A2(n18413), .ZN(n18408) );
  INV_X1 U18255 ( .A(n18410), .ZN(n18413) );
  OR2_X1 U18256 ( .A1(n15355), .A2(n14890), .ZN(n18001) );
  OR2_X1 U18257 ( .A1(n18414), .A2(n18415), .ZN(n17998) );
  INV_X1 U18258 ( .A(n18416), .ZN(n18415) );
  OR2_X1 U18259 ( .A1(n18417), .A2(n18418), .ZN(n18416) );
  AND2_X1 U18260 ( .A1(n18418), .A2(n18417), .ZN(n18414) );
  AND2_X1 U18261 ( .A1(n18419), .A2(n18420), .ZN(n18417) );
  OR2_X1 U18262 ( .A1(n18421), .A2(n18422), .ZN(n18420) );
  INV_X1 U18263 ( .A(n18423), .ZN(n18422) );
  OR2_X1 U18264 ( .A1(n18423), .A2(n18424), .ZN(n18419) );
  INV_X1 U18265 ( .A(n18421), .ZN(n18424) );
  OR2_X1 U18266 ( .A1(n15389), .A2(n14890), .ZN(n18012) );
  OR2_X1 U18267 ( .A1(n18425), .A2(n18426), .ZN(n18009) );
  INV_X1 U18268 ( .A(n18427), .ZN(n18426) );
  OR2_X1 U18269 ( .A1(n18428), .A2(n18429), .ZN(n18427) );
  AND2_X1 U18270 ( .A1(n18429), .A2(n18428), .ZN(n18425) );
  AND2_X1 U18271 ( .A1(n18430), .A2(n18431), .ZN(n18428) );
  OR2_X1 U18272 ( .A1(n18432), .A2(n18433), .ZN(n18431) );
  INV_X1 U18273 ( .A(n18434), .ZN(n18433) );
  OR2_X1 U18274 ( .A1(n18434), .A2(n18435), .ZN(n18430) );
  INV_X1 U18275 ( .A(n18432), .ZN(n18435) );
  OR2_X1 U18276 ( .A1(n15423), .A2(n14890), .ZN(n18023) );
  OR2_X1 U18277 ( .A1(n18436), .A2(n18437), .ZN(n18020) );
  INV_X1 U18278 ( .A(n18438), .ZN(n18437) );
  OR2_X1 U18279 ( .A1(n18439), .A2(n18440), .ZN(n18438) );
  AND2_X1 U18280 ( .A1(n18440), .A2(n18439), .ZN(n18436) );
  AND2_X1 U18281 ( .A1(n18441), .A2(n18442), .ZN(n18439) );
  OR2_X1 U18282 ( .A1(n18443), .A2(n18444), .ZN(n18442) );
  INV_X1 U18283 ( .A(n18445), .ZN(n18444) );
  OR2_X1 U18284 ( .A1(n18445), .A2(n18446), .ZN(n18441) );
  INV_X1 U18285 ( .A(n18443), .ZN(n18446) );
  OR2_X1 U18286 ( .A1(n15457), .A2(n14890), .ZN(n18034) );
  OR2_X1 U18287 ( .A1(n18447), .A2(n18448), .ZN(n18031) );
  INV_X1 U18288 ( .A(n18449), .ZN(n18448) );
  OR2_X1 U18289 ( .A1(n18450), .A2(n18451), .ZN(n18449) );
  AND2_X1 U18290 ( .A1(n18451), .A2(n18450), .ZN(n18447) );
  AND2_X1 U18291 ( .A1(n18452), .A2(n18453), .ZN(n18450) );
  OR2_X1 U18292 ( .A1(n18454), .A2(n18455), .ZN(n18453) );
  INV_X1 U18293 ( .A(n18456), .ZN(n18455) );
  OR2_X1 U18294 ( .A1(n18456), .A2(n18457), .ZN(n18452) );
  INV_X1 U18295 ( .A(n18454), .ZN(n18457) );
  OR2_X1 U18296 ( .A1(n15491), .A2(n14890), .ZN(n18045) );
  OR2_X1 U18297 ( .A1(n18458), .A2(n18459), .ZN(n18042) );
  INV_X1 U18298 ( .A(n18460), .ZN(n18459) );
  OR2_X1 U18299 ( .A1(n18461), .A2(n18462), .ZN(n18460) );
  AND2_X1 U18300 ( .A1(n18462), .A2(n18461), .ZN(n18458) );
  AND2_X1 U18301 ( .A1(n18463), .A2(n18464), .ZN(n18461) );
  OR2_X1 U18302 ( .A1(n18465), .A2(n18466), .ZN(n18464) );
  INV_X1 U18303 ( .A(n18467), .ZN(n18466) );
  OR2_X1 U18304 ( .A1(n18467), .A2(n18468), .ZN(n18463) );
  INV_X1 U18305 ( .A(n18465), .ZN(n18468) );
  OR2_X1 U18306 ( .A1(n15525), .A2(n14890), .ZN(n18056) );
  OR2_X1 U18307 ( .A1(n18469), .A2(n18470), .ZN(n18053) );
  INV_X1 U18308 ( .A(n18471), .ZN(n18470) );
  OR2_X1 U18309 ( .A1(n18472), .A2(n18473), .ZN(n18471) );
  AND2_X1 U18310 ( .A1(n18473), .A2(n18472), .ZN(n18469) );
  AND2_X1 U18311 ( .A1(n18474), .A2(n18475), .ZN(n18472) );
  OR2_X1 U18312 ( .A1(n18476), .A2(n18477), .ZN(n18475) );
  INV_X1 U18313 ( .A(n18478), .ZN(n18477) );
  OR2_X1 U18314 ( .A1(n18478), .A2(n18479), .ZN(n18474) );
  INV_X1 U18315 ( .A(n18476), .ZN(n18479) );
  OR2_X1 U18316 ( .A1(n15559), .A2(n14890), .ZN(n18067) );
  OR2_X1 U18317 ( .A1(n18480), .A2(n18481), .ZN(n18064) );
  INV_X1 U18318 ( .A(n18482), .ZN(n18481) );
  OR2_X1 U18319 ( .A1(n18483), .A2(n18484), .ZN(n18482) );
  AND2_X1 U18320 ( .A1(n18484), .A2(n18483), .ZN(n18480) );
  AND2_X1 U18321 ( .A1(n18485), .A2(n18486), .ZN(n18483) );
  OR2_X1 U18322 ( .A1(n18487), .A2(n18488), .ZN(n18486) );
  INV_X1 U18323 ( .A(n18489), .ZN(n18488) );
  OR2_X1 U18324 ( .A1(n18489), .A2(n18490), .ZN(n18485) );
  INV_X1 U18325 ( .A(n18487), .ZN(n18490) );
  OR2_X1 U18326 ( .A1(n15593), .A2(n14890), .ZN(n18078) );
  OR2_X1 U18327 ( .A1(n18491), .A2(n18492), .ZN(n18075) );
  INV_X1 U18328 ( .A(n18493), .ZN(n18492) );
  OR2_X1 U18329 ( .A1(n18494), .A2(n18495), .ZN(n18493) );
  AND2_X1 U18330 ( .A1(n18495), .A2(n18494), .ZN(n18491) );
  AND2_X1 U18331 ( .A1(n18496), .A2(n18497), .ZN(n18494) );
  OR2_X1 U18332 ( .A1(n18498), .A2(n18499), .ZN(n18497) );
  INV_X1 U18333 ( .A(n18500), .ZN(n18499) );
  OR2_X1 U18334 ( .A1(n18500), .A2(n18501), .ZN(n18496) );
  INV_X1 U18335 ( .A(n18498), .ZN(n18501) );
  OR2_X1 U18336 ( .A1(n15638), .A2(n14890), .ZN(n18089) );
  OR2_X1 U18337 ( .A1(n18502), .A2(n18503), .ZN(n18086) );
  INV_X1 U18338 ( .A(n18504), .ZN(n18503) );
  OR2_X1 U18339 ( .A1(n18505), .A2(n18506), .ZN(n18504) );
  AND2_X1 U18340 ( .A1(n18506), .A2(n18505), .ZN(n18502) );
  AND2_X1 U18341 ( .A1(n18507), .A2(n18508), .ZN(n18505) );
  OR2_X1 U18342 ( .A1(n18509), .A2(n18510), .ZN(n18508) );
  INV_X1 U18343 ( .A(n18511), .ZN(n18510) );
  OR2_X1 U18344 ( .A1(n18511), .A2(n18512), .ZN(n18507) );
  INV_X1 U18345 ( .A(n18509), .ZN(n18512) );
  OR2_X1 U18346 ( .A1(n15672), .A2(n14890), .ZN(n18100) );
  OR2_X1 U18347 ( .A1(n18513), .A2(n18514), .ZN(n18097) );
  INV_X1 U18348 ( .A(n18515), .ZN(n18514) );
  OR2_X1 U18349 ( .A1(n18516), .A2(n18517), .ZN(n18515) );
  AND2_X1 U18350 ( .A1(n18517), .A2(n18516), .ZN(n18513) );
  AND2_X1 U18351 ( .A1(n18518), .A2(n18519), .ZN(n18516) );
  OR2_X1 U18352 ( .A1(n18520), .A2(n18521), .ZN(n18519) );
  INV_X1 U18353 ( .A(n18522), .ZN(n18521) );
  OR2_X1 U18354 ( .A1(n18522), .A2(n18523), .ZN(n18518) );
  INV_X1 U18355 ( .A(n18520), .ZN(n18523) );
  OR2_X1 U18356 ( .A1(n15706), .A2(n14890), .ZN(n18111) );
  OR2_X1 U18357 ( .A1(n18524), .A2(n18525), .ZN(n18108) );
  INV_X1 U18358 ( .A(n18526), .ZN(n18525) );
  OR2_X1 U18359 ( .A1(n18527), .A2(n18528), .ZN(n18526) );
  AND2_X1 U18360 ( .A1(n18528), .A2(n18527), .ZN(n18524) );
  AND2_X1 U18361 ( .A1(n18529), .A2(n18530), .ZN(n18527) );
  OR2_X1 U18362 ( .A1(n18531), .A2(n18532), .ZN(n18530) );
  INV_X1 U18363 ( .A(n18533), .ZN(n18532) );
  OR2_X1 U18364 ( .A1(n18533), .A2(n18534), .ZN(n18529) );
  INV_X1 U18365 ( .A(n18531), .ZN(n18534) );
  OR2_X1 U18366 ( .A1(n15740), .A2(n14890), .ZN(n18122) );
  OR2_X1 U18367 ( .A1(n18535), .A2(n18536), .ZN(n18119) );
  INV_X1 U18368 ( .A(n18537), .ZN(n18536) );
  OR2_X1 U18369 ( .A1(n18538), .A2(n18539), .ZN(n18537) );
  AND2_X1 U18370 ( .A1(n18539), .A2(n18538), .ZN(n18535) );
  AND2_X1 U18371 ( .A1(n18540), .A2(n18541), .ZN(n18538) );
  OR2_X1 U18372 ( .A1(n18542), .A2(n18543), .ZN(n18541) );
  INV_X1 U18373 ( .A(n18544), .ZN(n18543) );
  OR2_X1 U18374 ( .A1(n18544), .A2(n18545), .ZN(n18540) );
  INV_X1 U18375 ( .A(n18542), .ZN(n18545) );
  OR2_X1 U18376 ( .A1(n15774), .A2(n14890), .ZN(n18133) );
  OR2_X1 U18377 ( .A1(n18546), .A2(n18547), .ZN(n18130) );
  INV_X1 U18378 ( .A(n18548), .ZN(n18547) );
  OR2_X1 U18379 ( .A1(n18549), .A2(n18550), .ZN(n18548) );
  AND2_X1 U18380 ( .A1(n18550), .A2(n18549), .ZN(n18546) );
  AND2_X1 U18381 ( .A1(n18551), .A2(n18552), .ZN(n18549) );
  OR2_X1 U18382 ( .A1(n18553), .A2(n18554), .ZN(n18552) );
  INV_X1 U18383 ( .A(n18555), .ZN(n18554) );
  OR2_X1 U18384 ( .A1(n18555), .A2(n18556), .ZN(n18551) );
  INV_X1 U18385 ( .A(n18553), .ZN(n18556) );
  OR2_X1 U18386 ( .A1(n15808), .A2(n14890), .ZN(n18144) );
  OR2_X1 U18387 ( .A1(n18557), .A2(n18558), .ZN(n18141) );
  INV_X1 U18388 ( .A(n18559), .ZN(n18558) );
  OR2_X1 U18389 ( .A1(n18560), .A2(n18561), .ZN(n18559) );
  AND2_X1 U18390 ( .A1(n18561), .A2(n18560), .ZN(n18557) );
  AND2_X1 U18391 ( .A1(n18562), .A2(n18563), .ZN(n18560) );
  OR2_X1 U18392 ( .A1(n18564), .A2(n18565), .ZN(n18563) );
  INV_X1 U18393 ( .A(n18566), .ZN(n18565) );
  OR2_X1 U18394 ( .A1(n18566), .A2(n18567), .ZN(n18562) );
  INV_X1 U18395 ( .A(n18564), .ZN(n18567) );
  OR2_X1 U18396 ( .A1(n15842), .A2(n14890), .ZN(n18158) );
  OR2_X1 U18397 ( .A1(n18568), .A2(n18569), .ZN(n18151) );
  INV_X1 U18398 ( .A(n18570), .ZN(n18569) );
  OR2_X1 U18399 ( .A1(n18571), .A2(n18572), .ZN(n18570) );
  AND2_X1 U18400 ( .A1(n18572), .A2(n18571), .ZN(n18568) );
  AND2_X1 U18401 ( .A1(n18573), .A2(n18574), .ZN(n18571) );
  INV_X1 U18402 ( .A(n18575), .ZN(n18574) );
  AND2_X1 U18403 ( .A1(n18576), .A2(n18577), .ZN(n18575) );
  OR2_X1 U18404 ( .A1(n18577), .A2(n18576), .ZN(n18573) );
  INV_X1 U18405 ( .A(n18578), .ZN(n18576) );
  OR2_X1 U18406 ( .A1(n16512), .A2(n14890), .ZN(n18168) );
  INV_X1 U18407 ( .A(b_28_), .ZN(n14890) );
  AND2_X1 U18408 ( .A1(n18579), .A2(n18580), .ZN(n18163) );
  INV_X1 U18409 ( .A(n18581), .ZN(n18580) );
  AND2_X1 U18410 ( .A1(n18582), .A2(n18583), .ZN(n18581) );
  OR2_X1 U18411 ( .A1(n18583), .A2(n18582), .ZN(n18579) );
  OR2_X1 U18412 ( .A1(n18584), .A2(n18585), .ZN(n18582) );
  AND2_X1 U18413 ( .A1(n18586), .A2(n18587), .ZN(n18585) );
  INV_X1 U18414 ( .A(n18588), .ZN(n18586) );
  AND2_X1 U18415 ( .A1(n18589), .A2(n18588), .ZN(n18584) );
  INV_X1 U18416 ( .A(n18587), .ZN(n18589) );
  INV_X1 U18417 ( .A(n18174), .ZN(n18172) );
  AND2_X1 U18418 ( .A1(n18590), .A2(n18591), .ZN(n18174) );
  INV_X1 U18419 ( .A(n18592), .ZN(n18591) );
  AND2_X1 U18420 ( .A1(n18593), .A2(n18594), .ZN(n18592) );
  OR2_X1 U18421 ( .A1(n18594), .A2(n18593), .ZN(n18590) );
  OR2_X1 U18422 ( .A1(n18595), .A2(n18596), .ZN(n18593) );
  AND2_X1 U18423 ( .A1(n18597), .A2(n18598), .ZN(n18596) );
  INV_X1 U18424 ( .A(n18599), .ZN(n18597) );
  AND2_X1 U18425 ( .A1(n18600), .A2(n18599), .ZN(n18595) );
  INV_X1 U18426 ( .A(n18598), .ZN(n18600) );
  OR2_X1 U18427 ( .A1(n18601), .A2(n18602), .ZN(n16873) );
  AND2_X1 U18428 ( .A1(n16818), .A2(n18603), .ZN(n18602) );
  AND2_X1 U18429 ( .A1(n18604), .A2(n16819), .ZN(n18601) );
  INV_X1 U18430 ( .A(n18603), .ZN(n16819) );
  OR2_X1 U18431 ( .A1(n18605), .A2(n18606), .ZN(n18603) );
  AND2_X1 U18432 ( .A1(n18599), .A2(n18598), .ZN(n18606) );
  AND2_X1 U18433 ( .A1(n18594), .A2(n18607), .ZN(n18605) );
  OR2_X1 U18434 ( .A1(n18599), .A2(n18598), .ZN(n18607) );
  OR2_X1 U18435 ( .A1(n18608), .A2(n18609), .ZN(n18598) );
  AND2_X1 U18436 ( .A1(n18588), .A2(n18587), .ZN(n18609) );
  AND2_X1 U18437 ( .A1(n18583), .A2(n18610), .ZN(n18608) );
  OR2_X1 U18438 ( .A1(n18588), .A2(n18587), .ZN(n18610) );
  OR2_X1 U18439 ( .A1(n18611), .A2(n18612), .ZN(n18587) );
  AND2_X1 U18440 ( .A1(n18578), .A2(n18577), .ZN(n18612) );
  AND2_X1 U18441 ( .A1(n18572), .A2(n18613), .ZN(n18611) );
  OR2_X1 U18442 ( .A1(n18578), .A2(n18577), .ZN(n18613) );
  OR2_X1 U18443 ( .A1(n18614), .A2(n18615), .ZN(n18577) );
  AND2_X1 U18444 ( .A1(n18564), .A2(n18566), .ZN(n18615) );
  AND2_X1 U18445 ( .A1(n18561), .A2(n18616), .ZN(n18614) );
  OR2_X1 U18446 ( .A1(n18564), .A2(n18566), .ZN(n18616) );
  OR2_X1 U18447 ( .A1(n18617), .A2(n18618), .ZN(n18566) );
  AND2_X1 U18448 ( .A1(n18553), .A2(n18555), .ZN(n18618) );
  AND2_X1 U18449 ( .A1(n18550), .A2(n18619), .ZN(n18617) );
  OR2_X1 U18450 ( .A1(n18553), .A2(n18555), .ZN(n18619) );
  OR2_X1 U18451 ( .A1(n18620), .A2(n18621), .ZN(n18555) );
  AND2_X1 U18452 ( .A1(n18542), .A2(n18544), .ZN(n18621) );
  AND2_X1 U18453 ( .A1(n18539), .A2(n18622), .ZN(n18620) );
  OR2_X1 U18454 ( .A1(n18542), .A2(n18544), .ZN(n18622) );
  OR2_X1 U18455 ( .A1(n18623), .A2(n18624), .ZN(n18544) );
  AND2_X1 U18456 ( .A1(n18531), .A2(n18533), .ZN(n18624) );
  AND2_X1 U18457 ( .A1(n18528), .A2(n18625), .ZN(n18623) );
  OR2_X1 U18458 ( .A1(n18531), .A2(n18533), .ZN(n18625) );
  OR2_X1 U18459 ( .A1(n18626), .A2(n18627), .ZN(n18533) );
  AND2_X1 U18460 ( .A1(n18520), .A2(n18522), .ZN(n18627) );
  AND2_X1 U18461 ( .A1(n18517), .A2(n18628), .ZN(n18626) );
  OR2_X1 U18462 ( .A1(n18520), .A2(n18522), .ZN(n18628) );
  OR2_X1 U18463 ( .A1(n18629), .A2(n18630), .ZN(n18522) );
  AND2_X1 U18464 ( .A1(n18509), .A2(n18511), .ZN(n18630) );
  AND2_X1 U18465 ( .A1(n18506), .A2(n18631), .ZN(n18629) );
  OR2_X1 U18466 ( .A1(n18509), .A2(n18511), .ZN(n18631) );
  OR2_X1 U18467 ( .A1(n18632), .A2(n18633), .ZN(n18511) );
  AND2_X1 U18468 ( .A1(n18498), .A2(n18500), .ZN(n18633) );
  AND2_X1 U18469 ( .A1(n18495), .A2(n18634), .ZN(n18632) );
  OR2_X1 U18470 ( .A1(n18498), .A2(n18500), .ZN(n18634) );
  OR2_X1 U18471 ( .A1(n18635), .A2(n18636), .ZN(n18500) );
  AND2_X1 U18472 ( .A1(n18487), .A2(n18489), .ZN(n18636) );
  AND2_X1 U18473 ( .A1(n18484), .A2(n18637), .ZN(n18635) );
  OR2_X1 U18474 ( .A1(n18487), .A2(n18489), .ZN(n18637) );
  OR2_X1 U18475 ( .A1(n18638), .A2(n18639), .ZN(n18489) );
  AND2_X1 U18476 ( .A1(n18476), .A2(n18478), .ZN(n18639) );
  AND2_X1 U18477 ( .A1(n18473), .A2(n18640), .ZN(n18638) );
  OR2_X1 U18478 ( .A1(n18476), .A2(n18478), .ZN(n18640) );
  OR2_X1 U18479 ( .A1(n18641), .A2(n18642), .ZN(n18478) );
  AND2_X1 U18480 ( .A1(n18465), .A2(n18467), .ZN(n18642) );
  AND2_X1 U18481 ( .A1(n18462), .A2(n18643), .ZN(n18641) );
  OR2_X1 U18482 ( .A1(n18465), .A2(n18467), .ZN(n18643) );
  OR2_X1 U18483 ( .A1(n18644), .A2(n18645), .ZN(n18467) );
  AND2_X1 U18484 ( .A1(n18454), .A2(n18456), .ZN(n18645) );
  AND2_X1 U18485 ( .A1(n18451), .A2(n18646), .ZN(n18644) );
  OR2_X1 U18486 ( .A1(n18454), .A2(n18456), .ZN(n18646) );
  OR2_X1 U18487 ( .A1(n18647), .A2(n18648), .ZN(n18456) );
  AND2_X1 U18488 ( .A1(n18443), .A2(n18445), .ZN(n18648) );
  AND2_X1 U18489 ( .A1(n18440), .A2(n18649), .ZN(n18647) );
  OR2_X1 U18490 ( .A1(n18443), .A2(n18445), .ZN(n18649) );
  OR2_X1 U18491 ( .A1(n18650), .A2(n18651), .ZN(n18445) );
  AND2_X1 U18492 ( .A1(n18432), .A2(n18434), .ZN(n18651) );
  AND2_X1 U18493 ( .A1(n18429), .A2(n18652), .ZN(n18650) );
  OR2_X1 U18494 ( .A1(n18432), .A2(n18434), .ZN(n18652) );
  OR2_X1 U18495 ( .A1(n18653), .A2(n18654), .ZN(n18434) );
  AND2_X1 U18496 ( .A1(n18421), .A2(n18423), .ZN(n18654) );
  AND2_X1 U18497 ( .A1(n18418), .A2(n18655), .ZN(n18653) );
  OR2_X1 U18498 ( .A1(n18421), .A2(n18423), .ZN(n18655) );
  OR2_X1 U18499 ( .A1(n18656), .A2(n18657), .ZN(n18423) );
  AND2_X1 U18500 ( .A1(n18410), .A2(n18412), .ZN(n18657) );
  AND2_X1 U18501 ( .A1(n18407), .A2(n18658), .ZN(n18656) );
  OR2_X1 U18502 ( .A1(n18410), .A2(n18412), .ZN(n18658) );
  OR2_X1 U18503 ( .A1(n18659), .A2(n18660), .ZN(n18412) );
  AND2_X1 U18504 ( .A1(n18399), .A2(n18401), .ZN(n18660) );
  AND2_X1 U18505 ( .A1(n18396), .A2(n18661), .ZN(n18659) );
  OR2_X1 U18506 ( .A1(n18399), .A2(n18401), .ZN(n18661) );
  OR2_X1 U18507 ( .A1(n18662), .A2(n18663), .ZN(n18401) );
  AND2_X1 U18508 ( .A1(n18388), .A2(n18390), .ZN(n18663) );
  AND2_X1 U18509 ( .A1(n18385), .A2(n18664), .ZN(n18662) );
  OR2_X1 U18510 ( .A1(n18388), .A2(n18390), .ZN(n18664) );
  OR2_X1 U18511 ( .A1(n18665), .A2(n18666), .ZN(n18390) );
  AND2_X1 U18512 ( .A1(n18377), .A2(n18379), .ZN(n18666) );
  AND2_X1 U18513 ( .A1(n18374), .A2(n18667), .ZN(n18665) );
  OR2_X1 U18514 ( .A1(n18377), .A2(n18379), .ZN(n18667) );
  OR2_X1 U18515 ( .A1(n18668), .A2(n18669), .ZN(n18379) );
  AND2_X1 U18516 ( .A1(n18366), .A2(n18368), .ZN(n18669) );
  AND2_X1 U18517 ( .A1(n18363), .A2(n18670), .ZN(n18668) );
  OR2_X1 U18518 ( .A1(n18366), .A2(n18368), .ZN(n18670) );
  OR2_X1 U18519 ( .A1(n18671), .A2(n18672), .ZN(n18368) );
  AND2_X1 U18520 ( .A1(n18355), .A2(n18357), .ZN(n18672) );
  AND2_X1 U18521 ( .A1(n18352), .A2(n18673), .ZN(n18671) );
  OR2_X1 U18522 ( .A1(n18355), .A2(n18357), .ZN(n18673) );
  OR2_X1 U18523 ( .A1(n18674), .A2(n18675), .ZN(n18357) );
  AND2_X1 U18524 ( .A1(n18344), .A2(n18346), .ZN(n18675) );
  AND2_X1 U18525 ( .A1(n18341), .A2(n18676), .ZN(n18674) );
  OR2_X1 U18526 ( .A1(n18344), .A2(n18346), .ZN(n18676) );
  OR2_X1 U18527 ( .A1(n18677), .A2(n18678), .ZN(n18346) );
  AND2_X1 U18528 ( .A1(n18333), .A2(n18335), .ZN(n18678) );
  AND2_X1 U18529 ( .A1(n18330), .A2(n18679), .ZN(n18677) );
  OR2_X1 U18530 ( .A1(n18333), .A2(n18335), .ZN(n18679) );
  OR2_X1 U18531 ( .A1(n18680), .A2(n18681), .ZN(n18335) );
  AND2_X1 U18532 ( .A1(n18322), .A2(n18324), .ZN(n18681) );
  AND2_X1 U18533 ( .A1(n18319), .A2(n18682), .ZN(n18680) );
  OR2_X1 U18534 ( .A1(n18322), .A2(n18324), .ZN(n18682) );
  OR2_X1 U18535 ( .A1(n18683), .A2(n18684), .ZN(n18324) );
  AND2_X1 U18536 ( .A1(n18311), .A2(n18313), .ZN(n18684) );
  AND2_X1 U18537 ( .A1(n18308), .A2(n18685), .ZN(n18683) );
  OR2_X1 U18538 ( .A1(n18311), .A2(n18313), .ZN(n18685) );
  OR2_X1 U18539 ( .A1(n18686), .A2(n18687), .ZN(n18313) );
  AND2_X1 U18540 ( .A1(n15948), .A2(n18302), .ZN(n18687) );
  AND2_X1 U18541 ( .A1(n18298), .A2(n18688), .ZN(n18686) );
  OR2_X1 U18542 ( .A1(n15948), .A2(n18302), .ZN(n18688) );
  OR2_X1 U18543 ( .A1(n18689), .A2(n18690), .ZN(n18302) );
  AND2_X1 U18544 ( .A1(n18290), .A2(n18292), .ZN(n18690) );
  AND2_X1 U18545 ( .A1(n18287), .A2(n18691), .ZN(n18689) );
  OR2_X1 U18546 ( .A1(n18290), .A2(n18292), .ZN(n18691) );
  OR2_X1 U18547 ( .A1(n18692), .A2(n18693), .ZN(n18292) );
  AND2_X1 U18548 ( .A1(n18275), .A2(n18280), .ZN(n18693) );
  AND2_X1 U18549 ( .A1(n18279), .A2(n18694), .ZN(n18692) );
  OR2_X1 U18550 ( .A1(n18275), .A2(n18280), .ZN(n18694) );
  INV_X1 U18551 ( .A(n18281), .ZN(n18280) );
  AND3_X1 U18552 ( .A1(b_27_), .A2(b_26_), .A3(n15957), .ZN(n18281) );
  OR2_X1 U18553 ( .A1(n14857), .A2(n14935), .ZN(n18275) );
  INV_X1 U18554 ( .A(n18282), .ZN(n18279) );
  OR2_X1 U18555 ( .A1(n18695), .A2(n18696), .ZN(n18282) );
  AND2_X1 U18556 ( .A1(b_26_), .A2(n18697), .ZN(n18696) );
  OR2_X1 U18557 ( .A1(n18698), .A2(n16981), .ZN(n18697) );
  AND2_X1 U18558 ( .A1(a_30_), .A2(n15003), .ZN(n18698) );
  AND2_X1 U18559 ( .A1(b_25_), .A2(n18699), .ZN(n18695) );
  OR2_X1 U18560 ( .A1(n18700), .A2(n14817), .ZN(n18699) );
  AND2_X1 U18561 ( .A1(a_31_), .A2(n14969), .ZN(n18700) );
  OR2_X1 U18562 ( .A1(n14891), .A2(n14935), .ZN(n18290) );
  OR2_X1 U18563 ( .A1(n18701), .A2(n18702), .ZN(n18287) );
  AND2_X1 U18564 ( .A1(n18703), .A2(n18704), .ZN(n18702) );
  INV_X1 U18565 ( .A(n18705), .ZN(n18701) );
  OR2_X1 U18566 ( .A1(n18703), .A2(n18704), .ZN(n18705) );
  OR2_X1 U18567 ( .A1(n18706), .A2(n18707), .ZN(n18703) );
  AND2_X1 U18568 ( .A1(n18708), .A2(n18709), .ZN(n18707) );
  AND2_X1 U18569 ( .A1(n18710), .A2(n18711), .ZN(n18706) );
  OR2_X1 U18570 ( .A1(n14936), .A2(n14935), .ZN(n15948) );
  OR2_X1 U18571 ( .A1(n18712), .A2(n18713), .ZN(n18298) );
  INV_X1 U18572 ( .A(n18714), .ZN(n18713) );
  OR2_X1 U18573 ( .A1(n18715), .A2(n18716), .ZN(n18714) );
  AND2_X1 U18574 ( .A1(n18716), .A2(n18715), .ZN(n18712) );
  AND2_X1 U18575 ( .A1(n18717), .A2(n18718), .ZN(n18715) );
  OR2_X1 U18576 ( .A1(n18719), .A2(n18720), .ZN(n18718) );
  INV_X1 U18577 ( .A(n18721), .ZN(n18720) );
  OR2_X1 U18578 ( .A1(n18721), .A2(n18722), .ZN(n18717) );
  INV_X1 U18579 ( .A(n18719), .ZN(n18722) );
  OR2_X1 U18580 ( .A1(n14970), .A2(n14935), .ZN(n18311) );
  OR2_X1 U18581 ( .A1(n18723), .A2(n18724), .ZN(n18308) );
  INV_X1 U18582 ( .A(n18725), .ZN(n18724) );
  OR2_X1 U18583 ( .A1(n18726), .A2(n18727), .ZN(n18725) );
  AND2_X1 U18584 ( .A1(n18727), .A2(n18726), .ZN(n18723) );
  AND2_X1 U18585 ( .A1(n18728), .A2(n18729), .ZN(n18726) );
  OR2_X1 U18586 ( .A1(n18730), .A2(n18731), .ZN(n18729) );
  INV_X1 U18587 ( .A(n18732), .ZN(n18731) );
  OR2_X1 U18588 ( .A1(n18732), .A2(n18733), .ZN(n18728) );
  INV_X1 U18589 ( .A(n18730), .ZN(n18733) );
  OR2_X1 U18590 ( .A1(n15004), .A2(n14935), .ZN(n18322) );
  OR2_X1 U18591 ( .A1(n18734), .A2(n18735), .ZN(n18319) );
  INV_X1 U18592 ( .A(n18736), .ZN(n18735) );
  OR2_X1 U18593 ( .A1(n18737), .A2(n18738), .ZN(n18736) );
  AND2_X1 U18594 ( .A1(n18738), .A2(n18737), .ZN(n18734) );
  AND2_X1 U18595 ( .A1(n18739), .A2(n18740), .ZN(n18737) );
  OR2_X1 U18596 ( .A1(n15945), .A2(n18741), .ZN(n18740) );
  INV_X1 U18597 ( .A(n18742), .ZN(n18741) );
  OR2_X1 U18598 ( .A1(n18742), .A2(n18743), .ZN(n18739) );
  INV_X1 U18599 ( .A(n15945), .ZN(n18743) );
  OR2_X1 U18600 ( .A1(n15038), .A2(n14935), .ZN(n18333) );
  OR2_X1 U18601 ( .A1(n18744), .A2(n18745), .ZN(n18330) );
  INV_X1 U18602 ( .A(n18746), .ZN(n18745) );
  OR2_X1 U18603 ( .A1(n18747), .A2(n18748), .ZN(n18746) );
  AND2_X1 U18604 ( .A1(n18748), .A2(n18747), .ZN(n18744) );
  AND2_X1 U18605 ( .A1(n18749), .A2(n18750), .ZN(n18747) );
  OR2_X1 U18606 ( .A1(n18751), .A2(n18752), .ZN(n18750) );
  INV_X1 U18607 ( .A(n18753), .ZN(n18752) );
  OR2_X1 U18608 ( .A1(n18753), .A2(n18754), .ZN(n18749) );
  INV_X1 U18609 ( .A(n18751), .ZN(n18754) );
  OR2_X1 U18610 ( .A1(n15072), .A2(n14935), .ZN(n18344) );
  OR2_X1 U18611 ( .A1(n18755), .A2(n18756), .ZN(n18341) );
  INV_X1 U18612 ( .A(n18757), .ZN(n18756) );
  OR2_X1 U18613 ( .A1(n18758), .A2(n18759), .ZN(n18757) );
  AND2_X1 U18614 ( .A1(n18759), .A2(n18758), .ZN(n18755) );
  AND2_X1 U18615 ( .A1(n18760), .A2(n18761), .ZN(n18758) );
  OR2_X1 U18616 ( .A1(n18762), .A2(n18763), .ZN(n18761) );
  INV_X1 U18617 ( .A(n18764), .ZN(n18763) );
  OR2_X1 U18618 ( .A1(n18764), .A2(n18765), .ZN(n18760) );
  INV_X1 U18619 ( .A(n18762), .ZN(n18765) );
  OR2_X1 U18620 ( .A1(n15106), .A2(n14935), .ZN(n18355) );
  OR2_X1 U18621 ( .A1(n18766), .A2(n18767), .ZN(n18352) );
  INV_X1 U18622 ( .A(n18768), .ZN(n18767) );
  OR2_X1 U18623 ( .A1(n18769), .A2(n18770), .ZN(n18768) );
  AND2_X1 U18624 ( .A1(n18770), .A2(n18769), .ZN(n18766) );
  AND2_X1 U18625 ( .A1(n18771), .A2(n18772), .ZN(n18769) );
  OR2_X1 U18626 ( .A1(n18773), .A2(n18774), .ZN(n18772) );
  INV_X1 U18627 ( .A(n18775), .ZN(n18774) );
  OR2_X1 U18628 ( .A1(n18775), .A2(n18776), .ZN(n18771) );
  INV_X1 U18629 ( .A(n18773), .ZN(n18776) );
  OR2_X1 U18630 ( .A1(n15140), .A2(n14935), .ZN(n18366) );
  OR2_X1 U18631 ( .A1(n18777), .A2(n18778), .ZN(n18363) );
  INV_X1 U18632 ( .A(n18779), .ZN(n18778) );
  OR2_X1 U18633 ( .A1(n18780), .A2(n18781), .ZN(n18779) );
  AND2_X1 U18634 ( .A1(n18781), .A2(n18780), .ZN(n18777) );
  AND2_X1 U18635 ( .A1(n18782), .A2(n18783), .ZN(n18780) );
  OR2_X1 U18636 ( .A1(n18784), .A2(n18785), .ZN(n18783) );
  INV_X1 U18637 ( .A(n18786), .ZN(n18785) );
  OR2_X1 U18638 ( .A1(n18786), .A2(n18787), .ZN(n18782) );
  INV_X1 U18639 ( .A(n18784), .ZN(n18787) );
  OR2_X1 U18640 ( .A1(n15174), .A2(n14935), .ZN(n18377) );
  OR2_X1 U18641 ( .A1(n18788), .A2(n18789), .ZN(n18374) );
  INV_X1 U18642 ( .A(n18790), .ZN(n18789) );
  OR2_X1 U18643 ( .A1(n18791), .A2(n18792), .ZN(n18790) );
  AND2_X1 U18644 ( .A1(n18792), .A2(n18791), .ZN(n18788) );
  AND2_X1 U18645 ( .A1(n18793), .A2(n18794), .ZN(n18791) );
  OR2_X1 U18646 ( .A1(n18795), .A2(n18796), .ZN(n18794) );
  INV_X1 U18647 ( .A(n18797), .ZN(n18796) );
  OR2_X1 U18648 ( .A1(n18797), .A2(n18798), .ZN(n18793) );
  INV_X1 U18649 ( .A(n18795), .ZN(n18798) );
  OR2_X1 U18650 ( .A1(n15208), .A2(n14935), .ZN(n18388) );
  OR2_X1 U18651 ( .A1(n18799), .A2(n18800), .ZN(n18385) );
  INV_X1 U18652 ( .A(n18801), .ZN(n18800) );
  OR2_X1 U18653 ( .A1(n18802), .A2(n18803), .ZN(n18801) );
  AND2_X1 U18654 ( .A1(n18803), .A2(n18802), .ZN(n18799) );
  AND2_X1 U18655 ( .A1(n18804), .A2(n18805), .ZN(n18802) );
  OR2_X1 U18656 ( .A1(n18806), .A2(n18807), .ZN(n18805) );
  INV_X1 U18657 ( .A(n18808), .ZN(n18807) );
  OR2_X1 U18658 ( .A1(n18808), .A2(n18809), .ZN(n18804) );
  INV_X1 U18659 ( .A(n18806), .ZN(n18809) );
  OR2_X1 U18660 ( .A1(n15242), .A2(n14935), .ZN(n18399) );
  OR2_X1 U18661 ( .A1(n18810), .A2(n18811), .ZN(n18396) );
  INV_X1 U18662 ( .A(n18812), .ZN(n18811) );
  OR2_X1 U18663 ( .A1(n18813), .A2(n18814), .ZN(n18812) );
  AND2_X1 U18664 ( .A1(n18814), .A2(n18813), .ZN(n18810) );
  AND2_X1 U18665 ( .A1(n18815), .A2(n18816), .ZN(n18813) );
  OR2_X1 U18666 ( .A1(n18817), .A2(n18818), .ZN(n18816) );
  INV_X1 U18667 ( .A(n18819), .ZN(n18818) );
  OR2_X1 U18668 ( .A1(n18819), .A2(n18820), .ZN(n18815) );
  INV_X1 U18669 ( .A(n18817), .ZN(n18820) );
  OR2_X1 U18670 ( .A1(n15287), .A2(n14935), .ZN(n18410) );
  OR2_X1 U18671 ( .A1(n18821), .A2(n18822), .ZN(n18407) );
  INV_X1 U18672 ( .A(n18823), .ZN(n18822) );
  OR2_X1 U18673 ( .A1(n18824), .A2(n18825), .ZN(n18823) );
  AND2_X1 U18674 ( .A1(n18825), .A2(n18824), .ZN(n18821) );
  AND2_X1 U18675 ( .A1(n18826), .A2(n18827), .ZN(n18824) );
  OR2_X1 U18676 ( .A1(n18828), .A2(n18829), .ZN(n18827) );
  INV_X1 U18677 ( .A(n18830), .ZN(n18829) );
  OR2_X1 U18678 ( .A1(n18830), .A2(n18831), .ZN(n18826) );
  INV_X1 U18679 ( .A(n18828), .ZN(n18831) );
  OR2_X1 U18680 ( .A1(n15321), .A2(n14935), .ZN(n18421) );
  OR2_X1 U18681 ( .A1(n18832), .A2(n18833), .ZN(n18418) );
  INV_X1 U18682 ( .A(n18834), .ZN(n18833) );
  OR2_X1 U18683 ( .A1(n18835), .A2(n18836), .ZN(n18834) );
  AND2_X1 U18684 ( .A1(n18836), .A2(n18835), .ZN(n18832) );
  AND2_X1 U18685 ( .A1(n18837), .A2(n18838), .ZN(n18835) );
  OR2_X1 U18686 ( .A1(n18839), .A2(n18840), .ZN(n18838) );
  INV_X1 U18687 ( .A(n18841), .ZN(n18840) );
  OR2_X1 U18688 ( .A1(n18841), .A2(n18842), .ZN(n18837) );
  INV_X1 U18689 ( .A(n18839), .ZN(n18842) );
  OR2_X1 U18690 ( .A1(n15355), .A2(n14935), .ZN(n18432) );
  OR2_X1 U18691 ( .A1(n18843), .A2(n18844), .ZN(n18429) );
  INV_X1 U18692 ( .A(n18845), .ZN(n18844) );
  OR2_X1 U18693 ( .A1(n18846), .A2(n18847), .ZN(n18845) );
  AND2_X1 U18694 ( .A1(n18847), .A2(n18846), .ZN(n18843) );
  AND2_X1 U18695 ( .A1(n18848), .A2(n18849), .ZN(n18846) );
  OR2_X1 U18696 ( .A1(n18850), .A2(n18851), .ZN(n18849) );
  INV_X1 U18697 ( .A(n18852), .ZN(n18851) );
  OR2_X1 U18698 ( .A1(n18852), .A2(n18853), .ZN(n18848) );
  INV_X1 U18699 ( .A(n18850), .ZN(n18853) );
  OR2_X1 U18700 ( .A1(n15389), .A2(n14935), .ZN(n18443) );
  OR2_X1 U18701 ( .A1(n18854), .A2(n18855), .ZN(n18440) );
  INV_X1 U18702 ( .A(n18856), .ZN(n18855) );
  OR2_X1 U18703 ( .A1(n18857), .A2(n18858), .ZN(n18856) );
  AND2_X1 U18704 ( .A1(n18858), .A2(n18857), .ZN(n18854) );
  AND2_X1 U18705 ( .A1(n18859), .A2(n18860), .ZN(n18857) );
  OR2_X1 U18706 ( .A1(n18861), .A2(n18862), .ZN(n18860) );
  INV_X1 U18707 ( .A(n18863), .ZN(n18862) );
  OR2_X1 U18708 ( .A1(n18863), .A2(n18864), .ZN(n18859) );
  INV_X1 U18709 ( .A(n18861), .ZN(n18864) );
  OR2_X1 U18710 ( .A1(n15423), .A2(n14935), .ZN(n18454) );
  OR2_X1 U18711 ( .A1(n18865), .A2(n18866), .ZN(n18451) );
  INV_X1 U18712 ( .A(n18867), .ZN(n18866) );
  OR2_X1 U18713 ( .A1(n18868), .A2(n18869), .ZN(n18867) );
  AND2_X1 U18714 ( .A1(n18869), .A2(n18868), .ZN(n18865) );
  AND2_X1 U18715 ( .A1(n18870), .A2(n18871), .ZN(n18868) );
  OR2_X1 U18716 ( .A1(n18872), .A2(n18873), .ZN(n18871) );
  INV_X1 U18717 ( .A(n18874), .ZN(n18873) );
  OR2_X1 U18718 ( .A1(n18874), .A2(n18875), .ZN(n18870) );
  INV_X1 U18719 ( .A(n18872), .ZN(n18875) );
  OR2_X1 U18720 ( .A1(n15457), .A2(n14935), .ZN(n18465) );
  OR2_X1 U18721 ( .A1(n18876), .A2(n18877), .ZN(n18462) );
  INV_X1 U18722 ( .A(n18878), .ZN(n18877) );
  OR2_X1 U18723 ( .A1(n18879), .A2(n18880), .ZN(n18878) );
  AND2_X1 U18724 ( .A1(n18880), .A2(n18879), .ZN(n18876) );
  AND2_X1 U18725 ( .A1(n18881), .A2(n18882), .ZN(n18879) );
  OR2_X1 U18726 ( .A1(n18883), .A2(n18884), .ZN(n18882) );
  INV_X1 U18727 ( .A(n18885), .ZN(n18884) );
  OR2_X1 U18728 ( .A1(n18885), .A2(n18886), .ZN(n18881) );
  INV_X1 U18729 ( .A(n18883), .ZN(n18886) );
  OR2_X1 U18730 ( .A1(n15491), .A2(n14935), .ZN(n18476) );
  OR2_X1 U18731 ( .A1(n18887), .A2(n18888), .ZN(n18473) );
  INV_X1 U18732 ( .A(n18889), .ZN(n18888) );
  OR2_X1 U18733 ( .A1(n18890), .A2(n18891), .ZN(n18889) );
  AND2_X1 U18734 ( .A1(n18891), .A2(n18890), .ZN(n18887) );
  AND2_X1 U18735 ( .A1(n18892), .A2(n18893), .ZN(n18890) );
  OR2_X1 U18736 ( .A1(n18894), .A2(n18895), .ZN(n18893) );
  INV_X1 U18737 ( .A(n18896), .ZN(n18895) );
  OR2_X1 U18738 ( .A1(n18896), .A2(n18897), .ZN(n18892) );
  INV_X1 U18739 ( .A(n18894), .ZN(n18897) );
  OR2_X1 U18740 ( .A1(n15525), .A2(n14935), .ZN(n18487) );
  OR2_X1 U18741 ( .A1(n18898), .A2(n18899), .ZN(n18484) );
  INV_X1 U18742 ( .A(n18900), .ZN(n18899) );
  OR2_X1 U18743 ( .A1(n18901), .A2(n18902), .ZN(n18900) );
  AND2_X1 U18744 ( .A1(n18902), .A2(n18901), .ZN(n18898) );
  AND2_X1 U18745 ( .A1(n18903), .A2(n18904), .ZN(n18901) );
  OR2_X1 U18746 ( .A1(n18905), .A2(n18906), .ZN(n18904) );
  INV_X1 U18747 ( .A(n18907), .ZN(n18906) );
  OR2_X1 U18748 ( .A1(n18907), .A2(n18908), .ZN(n18903) );
  INV_X1 U18749 ( .A(n18905), .ZN(n18908) );
  OR2_X1 U18750 ( .A1(n15559), .A2(n14935), .ZN(n18498) );
  OR2_X1 U18751 ( .A1(n18909), .A2(n18910), .ZN(n18495) );
  INV_X1 U18752 ( .A(n18911), .ZN(n18910) );
  OR2_X1 U18753 ( .A1(n18912), .A2(n18913), .ZN(n18911) );
  AND2_X1 U18754 ( .A1(n18913), .A2(n18912), .ZN(n18909) );
  AND2_X1 U18755 ( .A1(n18914), .A2(n18915), .ZN(n18912) );
  OR2_X1 U18756 ( .A1(n18916), .A2(n18917), .ZN(n18915) );
  INV_X1 U18757 ( .A(n18918), .ZN(n18917) );
  OR2_X1 U18758 ( .A1(n18918), .A2(n18919), .ZN(n18914) );
  INV_X1 U18759 ( .A(n18916), .ZN(n18919) );
  OR2_X1 U18760 ( .A1(n15593), .A2(n14935), .ZN(n18509) );
  OR2_X1 U18761 ( .A1(n18920), .A2(n18921), .ZN(n18506) );
  INV_X1 U18762 ( .A(n18922), .ZN(n18921) );
  OR2_X1 U18763 ( .A1(n18923), .A2(n18924), .ZN(n18922) );
  AND2_X1 U18764 ( .A1(n18924), .A2(n18923), .ZN(n18920) );
  AND2_X1 U18765 ( .A1(n18925), .A2(n18926), .ZN(n18923) );
  OR2_X1 U18766 ( .A1(n18927), .A2(n18928), .ZN(n18926) );
  INV_X1 U18767 ( .A(n18929), .ZN(n18928) );
  OR2_X1 U18768 ( .A1(n18929), .A2(n18930), .ZN(n18925) );
  INV_X1 U18769 ( .A(n18927), .ZN(n18930) );
  OR2_X1 U18770 ( .A1(n15638), .A2(n14935), .ZN(n18520) );
  OR2_X1 U18771 ( .A1(n18931), .A2(n18932), .ZN(n18517) );
  INV_X1 U18772 ( .A(n18933), .ZN(n18932) );
  OR2_X1 U18773 ( .A1(n18934), .A2(n18935), .ZN(n18933) );
  AND2_X1 U18774 ( .A1(n18935), .A2(n18934), .ZN(n18931) );
  AND2_X1 U18775 ( .A1(n18936), .A2(n18937), .ZN(n18934) );
  OR2_X1 U18776 ( .A1(n18938), .A2(n18939), .ZN(n18937) );
  INV_X1 U18777 ( .A(n18940), .ZN(n18939) );
  OR2_X1 U18778 ( .A1(n18940), .A2(n18941), .ZN(n18936) );
  INV_X1 U18779 ( .A(n18938), .ZN(n18941) );
  OR2_X1 U18780 ( .A1(n15672), .A2(n14935), .ZN(n18531) );
  OR2_X1 U18781 ( .A1(n18942), .A2(n18943), .ZN(n18528) );
  INV_X1 U18782 ( .A(n18944), .ZN(n18943) );
  OR2_X1 U18783 ( .A1(n18945), .A2(n18946), .ZN(n18944) );
  AND2_X1 U18784 ( .A1(n18946), .A2(n18945), .ZN(n18942) );
  AND2_X1 U18785 ( .A1(n18947), .A2(n18948), .ZN(n18945) );
  OR2_X1 U18786 ( .A1(n18949), .A2(n18950), .ZN(n18948) );
  INV_X1 U18787 ( .A(n18951), .ZN(n18950) );
  OR2_X1 U18788 ( .A1(n18951), .A2(n18952), .ZN(n18947) );
  INV_X1 U18789 ( .A(n18949), .ZN(n18952) );
  OR2_X1 U18790 ( .A1(n15706), .A2(n14935), .ZN(n18542) );
  OR2_X1 U18791 ( .A1(n18953), .A2(n18954), .ZN(n18539) );
  INV_X1 U18792 ( .A(n18955), .ZN(n18954) );
  OR2_X1 U18793 ( .A1(n18956), .A2(n18957), .ZN(n18955) );
  AND2_X1 U18794 ( .A1(n18957), .A2(n18956), .ZN(n18953) );
  AND2_X1 U18795 ( .A1(n18958), .A2(n18959), .ZN(n18956) );
  OR2_X1 U18796 ( .A1(n18960), .A2(n18961), .ZN(n18959) );
  INV_X1 U18797 ( .A(n18962), .ZN(n18961) );
  OR2_X1 U18798 ( .A1(n18962), .A2(n18963), .ZN(n18958) );
  INV_X1 U18799 ( .A(n18960), .ZN(n18963) );
  OR2_X1 U18800 ( .A1(n15740), .A2(n14935), .ZN(n18553) );
  OR2_X1 U18801 ( .A1(n18964), .A2(n18965), .ZN(n18550) );
  INV_X1 U18802 ( .A(n18966), .ZN(n18965) );
  OR2_X1 U18803 ( .A1(n18967), .A2(n18968), .ZN(n18966) );
  AND2_X1 U18804 ( .A1(n18968), .A2(n18967), .ZN(n18964) );
  AND2_X1 U18805 ( .A1(n18969), .A2(n18970), .ZN(n18967) );
  OR2_X1 U18806 ( .A1(n18971), .A2(n18972), .ZN(n18970) );
  INV_X1 U18807 ( .A(n18973), .ZN(n18972) );
  OR2_X1 U18808 ( .A1(n18973), .A2(n18974), .ZN(n18969) );
  INV_X1 U18809 ( .A(n18971), .ZN(n18974) );
  OR2_X1 U18810 ( .A1(n15774), .A2(n14935), .ZN(n18564) );
  OR2_X1 U18811 ( .A1(n18975), .A2(n18976), .ZN(n18561) );
  INV_X1 U18812 ( .A(n18977), .ZN(n18976) );
  OR2_X1 U18813 ( .A1(n18978), .A2(n18979), .ZN(n18977) );
  AND2_X1 U18814 ( .A1(n18979), .A2(n18978), .ZN(n18975) );
  AND2_X1 U18815 ( .A1(n18980), .A2(n18981), .ZN(n18978) );
  OR2_X1 U18816 ( .A1(n18982), .A2(n18983), .ZN(n18981) );
  INV_X1 U18817 ( .A(n18984), .ZN(n18983) );
  OR2_X1 U18818 ( .A1(n18984), .A2(n18985), .ZN(n18980) );
  INV_X1 U18819 ( .A(n18982), .ZN(n18985) );
  OR2_X1 U18820 ( .A1(n15808), .A2(n14935), .ZN(n18578) );
  OR2_X1 U18821 ( .A1(n18986), .A2(n18987), .ZN(n18572) );
  INV_X1 U18822 ( .A(n18988), .ZN(n18987) );
  OR2_X1 U18823 ( .A1(n18989), .A2(n18990), .ZN(n18988) );
  AND2_X1 U18824 ( .A1(n18990), .A2(n18989), .ZN(n18986) );
  AND2_X1 U18825 ( .A1(n18991), .A2(n18992), .ZN(n18989) );
  INV_X1 U18826 ( .A(n18993), .ZN(n18992) );
  AND2_X1 U18827 ( .A1(n18994), .A2(n18995), .ZN(n18993) );
  OR2_X1 U18828 ( .A1(n18995), .A2(n18994), .ZN(n18991) );
  INV_X1 U18829 ( .A(n18996), .ZN(n18994) );
  OR2_X1 U18830 ( .A1(n15842), .A2(n14935), .ZN(n18588) );
  AND2_X1 U18831 ( .A1(n18997), .A2(n18998), .ZN(n18583) );
  INV_X1 U18832 ( .A(n18999), .ZN(n18998) );
  AND2_X1 U18833 ( .A1(n19000), .A2(n19001), .ZN(n18999) );
  OR2_X1 U18834 ( .A1(n19001), .A2(n19000), .ZN(n18997) );
  OR2_X1 U18835 ( .A1(n19002), .A2(n19003), .ZN(n19000) );
  AND2_X1 U18836 ( .A1(n19004), .A2(n19005), .ZN(n19003) );
  INV_X1 U18837 ( .A(n19006), .ZN(n19004) );
  AND2_X1 U18838 ( .A1(n19007), .A2(n19006), .ZN(n19002) );
  INV_X1 U18839 ( .A(n19005), .ZN(n19007) );
  OR2_X1 U18840 ( .A1(n16512), .A2(n14935), .ZN(n18599) );
  INV_X1 U18841 ( .A(b_27_), .ZN(n14935) );
  AND2_X1 U18842 ( .A1(n19008), .A2(n19009), .ZN(n18594) );
  INV_X1 U18843 ( .A(n19010), .ZN(n19009) );
  AND2_X1 U18844 ( .A1(n19011), .A2(n19012), .ZN(n19010) );
  OR2_X1 U18845 ( .A1(n19012), .A2(n19011), .ZN(n19008) );
  OR2_X1 U18846 ( .A1(n19013), .A2(n19014), .ZN(n19011) );
  AND2_X1 U18847 ( .A1(n19015), .A2(n19016), .ZN(n19014) );
  INV_X1 U18848 ( .A(n19017), .ZN(n19015) );
  AND2_X1 U18849 ( .A1(n19018), .A2(n19017), .ZN(n19013) );
  INV_X1 U18850 ( .A(n19016), .ZN(n19018) );
  INV_X1 U18851 ( .A(n16818), .ZN(n18604) );
  OR2_X1 U18852 ( .A1(n19019), .A2(n19020), .ZN(n16818) );
  AND2_X1 U18853 ( .A1(n19021), .A2(n16831), .ZN(n19020) );
  INV_X1 U18854 ( .A(n19022), .ZN(n19019) );
  OR2_X1 U18855 ( .A1(n16831), .A2(n19021), .ZN(n19022) );
  OR2_X1 U18856 ( .A1(n19023), .A2(n19024), .ZN(n19021) );
  AND2_X1 U18857 ( .A1(n19025), .A2(n16830), .ZN(n19024) );
  INV_X1 U18858 ( .A(n16829), .ZN(n19025) );
  AND2_X1 U18859 ( .A1(n19026), .A2(n16829), .ZN(n19023) );
  OR2_X1 U18860 ( .A1(n16512), .A2(n14969), .ZN(n16829) );
  INV_X1 U18861 ( .A(n16830), .ZN(n19026) );
  OR2_X1 U18862 ( .A1(n19027), .A2(n19028), .ZN(n16830) );
  AND2_X1 U18863 ( .A1(n19017), .A2(n19016), .ZN(n19028) );
  AND2_X1 U18864 ( .A1(n19012), .A2(n19029), .ZN(n19027) );
  OR2_X1 U18865 ( .A1(n19017), .A2(n19016), .ZN(n19029) );
  OR2_X1 U18866 ( .A1(n19030), .A2(n19031), .ZN(n19016) );
  AND2_X1 U18867 ( .A1(n19006), .A2(n19005), .ZN(n19031) );
  AND2_X1 U18868 ( .A1(n19001), .A2(n19032), .ZN(n19030) );
  OR2_X1 U18869 ( .A1(n19006), .A2(n19005), .ZN(n19032) );
  OR2_X1 U18870 ( .A1(n19033), .A2(n19034), .ZN(n19005) );
  AND2_X1 U18871 ( .A1(n18996), .A2(n18995), .ZN(n19034) );
  AND2_X1 U18872 ( .A1(n18990), .A2(n19035), .ZN(n19033) );
  OR2_X1 U18873 ( .A1(n18996), .A2(n18995), .ZN(n19035) );
  OR2_X1 U18874 ( .A1(n19036), .A2(n19037), .ZN(n18995) );
  AND2_X1 U18875 ( .A1(n18982), .A2(n18984), .ZN(n19037) );
  AND2_X1 U18876 ( .A1(n18979), .A2(n19038), .ZN(n19036) );
  OR2_X1 U18877 ( .A1(n18982), .A2(n18984), .ZN(n19038) );
  OR2_X1 U18878 ( .A1(n19039), .A2(n19040), .ZN(n18984) );
  AND2_X1 U18879 ( .A1(n18971), .A2(n18973), .ZN(n19040) );
  AND2_X1 U18880 ( .A1(n18968), .A2(n19041), .ZN(n19039) );
  OR2_X1 U18881 ( .A1(n18971), .A2(n18973), .ZN(n19041) );
  OR2_X1 U18882 ( .A1(n19042), .A2(n19043), .ZN(n18973) );
  AND2_X1 U18883 ( .A1(n18960), .A2(n18962), .ZN(n19043) );
  AND2_X1 U18884 ( .A1(n18957), .A2(n19044), .ZN(n19042) );
  OR2_X1 U18885 ( .A1(n18960), .A2(n18962), .ZN(n19044) );
  OR2_X1 U18886 ( .A1(n19045), .A2(n19046), .ZN(n18962) );
  AND2_X1 U18887 ( .A1(n18949), .A2(n18951), .ZN(n19046) );
  AND2_X1 U18888 ( .A1(n18946), .A2(n19047), .ZN(n19045) );
  OR2_X1 U18889 ( .A1(n18949), .A2(n18951), .ZN(n19047) );
  OR2_X1 U18890 ( .A1(n19048), .A2(n19049), .ZN(n18951) );
  AND2_X1 U18891 ( .A1(n18938), .A2(n18940), .ZN(n19049) );
  AND2_X1 U18892 ( .A1(n18935), .A2(n19050), .ZN(n19048) );
  OR2_X1 U18893 ( .A1(n18938), .A2(n18940), .ZN(n19050) );
  OR2_X1 U18894 ( .A1(n19051), .A2(n19052), .ZN(n18940) );
  AND2_X1 U18895 ( .A1(n18927), .A2(n18929), .ZN(n19052) );
  AND2_X1 U18896 ( .A1(n18924), .A2(n19053), .ZN(n19051) );
  OR2_X1 U18897 ( .A1(n18927), .A2(n18929), .ZN(n19053) );
  OR2_X1 U18898 ( .A1(n19054), .A2(n19055), .ZN(n18929) );
  AND2_X1 U18899 ( .A1(n18916), .A2(n18918), .ZN(n19055) );
  AND2_X1 U18900 ( .A1(n18913), .A2(n19056), .ZN(n19054) );
  OR2_X1 U18901 ( .A1(n18916), .A2(n18918), .ZN(n19056) );
  OR2_X1 U18902 ( .A1(n19057), .A2(n19058), .ZN(n18918) );
  AND2_X1 U18903 ( .A1(n18905), .A2(n18907), .ZN(n19058) );
  AND2_X1 U18904 ( .A1(n18902), .A2(n19059), .ZN(n19057) );
  OR2_X1 U18905 ( .A1(n18905), .A2(n18907), .ZN(n19059) );
  OR2_X1 U18906 ( .A1(n19060), .A2(n19061), .ZN(n18907) );
  AND2_X1 U18907 ( .A1(n18894), .A2(n18896), .ZN(n19061) );
  AND2_X1 U18908 ( .A1(n18891), .A2(n19062), .ZN(n19060) );
  OR2_X1 U18909 ( .A1(n18894), .A2(n18896), .ZN(n19062) );
  OR2_X1 U18910 ( .A1(n19063), .A2(n19064), .ZN(n18896) );
  AND2_X1 U18911 ( .A1(n18883), .A2(n18885), .ZN(n19064) );
  AND2_X1 U18912 ( .A1(n18880), .A2(n19065), .ZN(n19063) );
  OR2_X1 U18913 ( .A1(n18883), .A2(n18885), .ZN(n19065) );
  OR2_X1 U18914 ( .A1(n19066), .A2(n19067), .ZN(n18885) );
  AND2_X1 U18915 ( .A1(n18872), .A2(n18874), .ZN(n19067) );
  AND2_X1 U18916 ( .A1(n18869), .A2(n19068), .ZN(n19066) );
  OR2_X1 U18917 ( .A1(n18872), .A2(n18874), .ZN(n19068) );
  OR2_X1 U18918 ( .A1(n19069), .A2(n19070), .ZN(n18874) );
  AND2_X1 U18919 ( .A1(n18861), .A2(n18863), .ZN(n19070) );
  AND2_X1 U18920 ( .A1(n18858), .A2(n19071), .ZN(n19069) );
  OR2_X1 U18921 ( .A1(n18861), .A2(n18863), .ZN(n19071) );
  OR2_X1 U18922 ( .A1(n19072), .A2(n19073), .ZN(n18863) );
  AND2_X1 U18923 ( .A1(n18850), .A2(n18852), .ZN(n19073) );
  AND2_X1 U18924 ( .A1(n18847), .A2(n19074), .ZN(n19072) );
  OR2_X1 U18925 ( .A1(n18850), .A2(n18852), .ZN(n19074) );
  OR2_X1 U18926 ( .A1(n19075), .A2(n19076), .ZN(n18852) );
  AND2_X1 U18927 ( .A1(n18839), .A2(n18841), .ZN(n19076) );
  AND2_X1 U18928 ( .A1(n18836), .A2(n19077), .ZN(n19075) );
  OR2_X1 U18929 ( .A1(n18839), .A2(n18841), .ZN(n19077) );
  OR2_X1 U18930 ( .A1(n19078), .A2(n19079), .ZN(n18841) );
  AND2_X1 U18931 ( .A1(n18828), .A2(n18830), .ZN(n19079) );
  AND2_X1 U18932 ( .A1(n18825), .A2(n19080), .ZN(n19078) );
  OR2_X1 U18933 ( .A1(n18828), .A2(n18830), .ZN(n19080) );
  OR2_X1 U18934 ( .A1(n19081), .A2(n19082), .ZN(n18830) );
  AND2_X1 U18935 ( .A1(n18817), .A2(n18819), .ZN(n19082) );
  AND2_X1 U18936 ( .A1(n18814), .A2(n19083), .ZN(n19081) );
  OR2_X1 U18937 ( .A1(n18817), .A2(n18819), .ZN(n19083) );
  OR2_X1 U18938 ( .A1(n19084), .A2(n19085), .ZN(n18819) );
  AND2_X1 U18939 ( .A1(n18806), .A2(n18808), .ZN(n19085) );
  AND2_X1 U18940 ( .A1(n18803), .A2(n19086), .ZN(n19084) );
  OR2_X1 U18941 ( .A1(n18806), .A2(n18808), .ZN(n19086) );
  OR2_X1 U18942 ( .A1(n19087), .A2(n19088), .ZN(n18808) );
  AND2_X1 U18943 ( .A1(n18795), .A2(n18797), .ZN(n19088) );
  AND2_X1 U18944 ( .A1(n18792), .A2(n19089), .ZN(n19087) );
  OR2_X1 U18945 ( .A1(n18795), .A2(n18797), .ZN(n19089) );
  OR2_X1 U18946 ( .A1(n19090), .A2(n19091), .ZN(n18797) );
  AND2_X1 U18947 ( .A1(n18784), .A2(n18786), .ZN(n19091) );
  AND2_X1 U18948 ( .A1(n18781), .A2(n19092), .ZN(n19090) );
  OR2_X1 U18949 ( .A1(n18784), .A2(n18786), .ZN(n19092) );
  OR2_X1 U18950 ( .A1(n19093), .A2(n19094), .ZN(n18786) );
  AND2_X1 U18951 ( .A1(n18773), .A2(n18775), .ZN(n19094) );
  AND2_X1 U18952 ( .A1(n18770), .A2(n19095), .ZN(n19093) );
  OR2_X1 U18953 ( .A1(n18773), .A2(n18775), .ZN(n19095) );
  OR2_X1 U18954 ( .A1(n19096), .A2(n19097), .ZN(n18775) );
  AND2_X1 U18955 ( .A1(n18762), .A2(n18764), .ZN(n19097) );
  AND2_X1 U18956 ( .A1(n18759), .A2(n19098), .ZN(n19096) );
  OR2_X1 U18957 ( .A1(n18762), .A2(n18764), .ZN(n19098) );
  OR2_X1 U18958 ( .A1(n19099), .A2(n19100), .ZN(n18764) );
  AND2_X1 U18959 ( .A1(n18751), .A2(n18753), .ZN(n19100) );
  AND2_X1 U18960 ( .A1(n18748), .A2(n19101), .ZN(n19099) );
  OR2_X1 U18961 ( .A1(n18751), .A2(n18753), .ZN(n19101) );
  OR2_X1 U18962 ( .A1(n19102), .A2(n19103), .ZN(n18753) );
  AND2_X1 U18963 ( .A1(n15945), .A2(n18742), .ZN(n19103) );
  AND2_X1 U18964 ( .A1(n18738), .A2(n19104), .ZN(n19102) );
  OR2_X1 U18965 ( .A1(n15945), .A2(n18742), .ZN(n19104) );
  OR2_X1 U18966 ( .A1(n19105), .A2(n19106), .ZN(n18742) );
  AND2_X1 U18967 ( .A1(n18730), .A2(n18732), .ZN(n19106) );
  AND2_X1 U18968 ( .A1(n18727), .A2(n19107), .ZN(n19105) );
  OR2_X1 U18969 ( .A1(n18730), .A2(n18732), .ZN(n19107) );
  OR2_X1 U18970 ( .A1(n19108), .A2(n19109), .ZN(n18732) );
  AND2_X1 U18971 ( .A1(n18719), .A2(n18721), .ZN(n19109) );
  AND2_X1 U18972 ( .A1(n18716), .A2(n19110), .ZN(n19108) );
  OR2_X1 U18973 ( .A1(n18719), .A2(n18721), .ZN(n19110) );
  OR2_X1 U18974 ( .A1(n19111), .A2(n19112), .ZN(n18721) );
  AND2_X1 U18975 ( .A1(n18704), .A2(n18709), .ZN(n19112) );
  AND2_X1 U18976 ( .A1(n18708), .A2(n19113), .ZN(n19111) );
  OR2_X1 U18977 ( .A1(n18704), .A2(n18709), .ZN(n19113) );
  INV_X1 U18978 ( .A(n18710), .ZN(n18709) );
  AND3_X1 U18979 ( .A1(b_26_), .A2(b_25_), .A3(n15957), .ZN(n18710) );
  OR2_X1 U18980 ( .A1(n14857), .A2(n14969), .ZN(n18704) );
  INV_X1 U18981 ( .A(n18711), .ZN(n18708) );
  OR2_X1 U18982 ( .A1(n19114), .A2(n19115), .ZN(n18711) );
  AND2_X1 U18983 ( .A1(b_25_), .A2(n19116), .ZN(n19115) );
  OR2_X1 U18984 ( .A1(n19117), .A2(n16981), .ZN(n19116) );
  AND2_X1 U18985 ( .A1(a_30_), .A2(n15037), .ZN(n19117) );
  AND2_X1 U18986 ( .A1(b_24_), .A2(n19118), .ZN(n19114) );
  OR2_X1 U18987 ( .A1(n19119), .A2(n14817), .ZN(n19118) );
  AND2_X1 U18988 ( .A1(a_31_), .A2(n15003), .ZN(n19119) );
  OR2_X1 U18989 ( .A1(n14891), .A2(n14969), .ZN(n18719) );
  OR2_X1 U18990 ( .A1(n19120), .A2(n19121), .ZN(n18716) );
  AND2_X1 U18991 ( .A1(n19122), .A2(n19123), .ZN(n19121) );
  INV_X1 U18992 ( .A(n19124), .ZN(n19120) );
  OR2_X1 U18993 ( .A1(n19122), .A2(n19123), .ZN(n19124) );
  OR2_X1 U18994 ( .A1(n19125), .A2(n19126), .ZN(n19122) );
  AND2_X1 U18995 ( .A1(n19127), .A2(n19128), .ZN(n19126) );
  AND2_X1 U18996 ( .A1(n19129), .A2(n19130), .ZN(n19125) );
  OR2_X1 U18997 ( .A1(n14936), .A2(n14969), .ZN(n18730) );
  OR2_X1 U18998 ( .A1(n19131), .A2(n19132), .ZN(n18727) );
  INV_X1 U18999 ( .A(n19133), .ZN(n19132) );
  OR2_X1 U19000 ( .A1(n19134), .A2(n19135), .ZN(n19133) );
  AND2_X1 U19001 ( .A1(n19135), .A2(n19134), .ZN(n19131) );
  AND2_X1 U19002 ( .A1(n19136), .A2(n19137), .ZN(n19134) );
  OR2_X1 U19003 ( .A1(n19138), .A2(n19139), .ZN(n19137) );
  INV_X1 U19004 ( .A(n19140), .ZN(n19139) );
  OR2_X1 U19005 ( .A1(n19140), .A2(n19141), .ZN(n19136) );
  INV_X1 U19006 ( .A(n19138), .ZN(n19141) );
  OR2_X1 U19007 ( .A1(n14970), .A2(n14969), .ZN(n15945) );
  OR2_X1 U19008 ( .A1(n19142), .A2(n19143), .ZN(n18738) );
  INV_X1 U19009 ( .A(n19144), .ZN(n19143) );
  OR2_X1 U19010 ( .A1(n19145), .A2(n19146), .ZN(n19144) );
  AND2_X1 U19011 ( .A1(n19146), .A2(n19145), .ZN(n19142) );
  AND2_X1 U19012 ( .A1(n19147), .A2(n19148), .ZN(n19145) );
  OR2_X1 U19013 ( .A1(n19149), .A2(n19150), .ZN(n19148) );
  INV_X1 U19014 ( .A(n19151), .ZN(n19150) );
  OR2_X1 U19015 ( .A1(n19151), .A2(n19152), .ZN(n19147) );
  INV_X1 U19016 ( .A(n19149), .ZN(n19152) );
  OR2_X1 U19017 ( .A1(n15004), .A2(n14969), .ZN(n18751) );
  OR2_X1 U19018 ( .A1(n19153), .A2(n19154), .ZN(n18748) );
  INV_X1 U19019 ( .A(n19155), .ZN(n19154) );
  OR2_X1 U19020 ( .A1(n19156), .A2(n19157), .ZN(n19155) );
  AND2_X1 U19021 ( .A1(n19157), .A2(n19156), .ZN(n19153) );
  AND2_X1 U19022 ( .A1(n19158), .A2(n19159), .ZN(n19156) );
  OR2_X1 U19023 ( .A1(n19160), .A2(n19161), .ZN(n19159) );
  INV_X1 U19024 ( .A(n19162), .ZN(n19161) );
  OR2_X1 U19025 ( .A1(n19162), .A2(n19163), .ZN(n19158) );
  INV_X1 U19026 ( .A(n19160), .ZN(n19163) );
  OR2_X1 U19027 ( .A1(n15038), .A2(n14969), .ZN(n18762) );
  OR2_X1 U19028 ( .A1(n19164), .A2(n19165), .ZN(n18759) );
  INV_X1 U19029 ( .A(n19166), .ZN(n19165) );
  OR2_X1 U19030 ( .A1(n19167), .A2(n19168), .ZN(n19166) );
  AND2_X1 U19031 ( .A1(n19168), .A2(n19167), .ZN(n19164) );
  AND2_X1 U19032 ( .A1(n19169), .A2(n19170), .ZN(n19167) );
  OR2_X1 U19033 ( .A1(n15942), .A2(n19171), .ZN(n19170) );
  INV_X1 U19034 ( .A(n19172), .ZN(n19171) );
  OR2_X1 U19035 ( .A1(n19172), .A2(n19173), .ZN(n19169) );
  INV_X1 U19036 ( .A(n15942), .ZN(n19173) );
  OR2_X1 U19037 ( .A1(n15072), .A2(n14969), .ZN(n18773) );
  OR2_X1 U19038 ( .A1(n19174), .A2(n19175), .ZN(n18770) );
  INV_X1 U19039 ( .A(n19176), .ZN(n19175) );
  OR2_X1 U19040 ( .A1(n19177), .A2(n19178), .ZN(n19176) );
  AND2_X1 U19041 ( .A1(n19178), .A2(n19177), .ZN(n19174) );
  AND2_X1 U19042 ( .A1(n19179), .A2(n19180), .ZN(n19177) );
  OR2_X1 U19043 ( .A1(n19181), .A2(n19182), .ZN(n19180) );
  INV_X1 U19044 ( .A(n19183), .ZN(n19182) );
  OR2_X1 U19045 ( .A1(n19183), .A2(n19184), .ZN(n19179) );
  INV_X1 U19046 ( .A(n19181), .ZN(n19184) );
  OR2_X1 U19047 ( .A1(n15106), .A2(n14969), .ZN(n18784) );
  OR2_X1 U19048 ( .A1(n19185), .A2(n19186), .ZN(n18781) );
  INV_X1 U19049 ( .A(n19187), .ZN(n19186) );
  OR2_X1 U19050 ( .A1(n19188), .A2(n19189), .ZN(n19187) );
  AND2_X1 U19051 ( .A1(n19189), .A2(n19188), .ZN(n19185) );
  AND2_X1 U19052 ( .A1(n19190), .A2(n19191), .ZN(n19188) );
  OR2_X1 U19053 ( .A1(n19192), .A2(n19193), .ZN(n19191) );
  INV_X1 U19054 ( .A(n19194), .ZN(n19193) );
  OR2_X1 U19055 ( .A1(n19194), .A2(n19195), .ZN(n19190) );
  INV_X1 U19056 ( .A(n19192), .ZN(n19195) );
  OR2_X1 U19057 ( .A1(n15140), .A2(n14969), .ZN(n18795) );
  OR2_X1 U19058 ( .A1(n19196), .A2(n19197), .ZN(n18792) );
  INV_X1 U19059 ( .A(n19198), .ZN(n19197) );
  OR2_X1 U19060 ( .A1(n19199), .A2(n19200), .ZN(n19198) );
  AND2_X1 U19061 ( .A1(n19200), .A2(n19199), .ZN(n19196) );
  AND2_X1 U19062 ( .A1(n19201), .A2(n19202), .ZN(n19199) );
  OR2_X1 U19063 ( .A1(n19203), .A2(n19204), .ZN(n19202) );
  INV_X1 U19064 ( .A(n19205), .ZN(n19204) );
  OR2_X1 U19065 ( .A1(n19205), .A2(n19206), .ZN(n19201) );
  INV_X1 U19066 ( .A(n19203), .ZN(n19206) );
  OR2_X1 U19067 ( .A1(n15174), .A2(n14969), .ZN(n18806) );
  OR2_X1 U19068 ( .A1(n19207), .A2(n19208), .ZN(n18803) );
  INV_X1 U19069 ( .A(n19209), .ZN(n19208) );
  OR2_X1 U19070 ( .A1(n19210), .A2(n19211), .ZN(n19209) );
  AND2_X1 U19071 ( .A1(n19211), .A2(n19210), .ZN(n19207) );
  AND2_X1 U19072 ( .A1(n19212), .A2(n19213), .ZN(n19210) );
  OR2_X1 U19073 ( .A1(n19214), .A2(n19215), .ZN(n19213) );
  INV_X1 U19074 ( .A(n19216), .ZN(n19215) );
  OR2_X1 U19075 ( .A1(n19216), .A2(n19217), .ZN(n19212) );
  INV_X1 U19076 ( .A(n19214), .ZN(n19217) );
  OR2_X1 U19077 ( .A1(n15208), .A2(n14969), .ZN(n18817) );
  OR2_X1 U19078 ( .A1(n19218), .A2(n19219), .ZN(n18814) );
  INV_X1 U19079 ( .A(n19220), .ZN(n19219) );
  OR2_X1 U19080 ( .A1(n19221), .A2(n19222), .ZN(n19220) );
  AND2_X1 U19081 ( .A1(n19222), .A2(n19221), .ZN(n19218) );
  AND2_X1 U19082 ( .A1(n19223), .A2(n19224), .ZN(n19221) );
  OR2_X1 U19083 ( .A1(n19225), .A2(n19226), .ZN(n19224) );
  INV_X1 U19084 ( .A(n19227), .ZN(n19226) );
  OR2_X1 U19085 ( .A1(n19227), .A2(n19228), .ZN(n19223) );
  INV_X1 U19086 ( .A(n19225), .ZN(n19228) );
  OR2_X1 U19087 ( .A1(n15242), .A2(n14969), .ZN(n18828) );
  OR2_X1 U19088 ( .A1(n19229), .A2(n19230), .ZN(n18825) );
  INV_X1 U19089 ( .A(n19231), .ZN(n19230) );
  OR2_X1 U19090 ( .A1(n19232), .A2(n19233), .ZN(n19231) );
  AND2_X1 U19091 ( .A1(n19233), .A2(n19232), .ZN(n19229) );
  AND2_X1 U19092 ( .A1(n19234), .A2(n19235), .ZN(n19232) );
  OR2_X1 U19093 ( .A1(n19236), .A2(n19237), .ZN(n19235) );
  INV_X1 U19094 ( .A(n19238), .ZN(n19237) );
  OR2_X1 U19095 ( .A1(n19238), .A2(n19239), .ZN(n19234) );
  INV_X1 U19096 ( .A(n19236), .ZN(n19239) );
  OR2_X1 U19097 ( .A1(n15287), .A2(n14969), .ZN(n18839) );
  OR2_X1 U19098 ( .A1(n19240), .A2(n19241), .ZN(n18836) );
  INV_X1 U19099 ( .A(n19242), .ZN(n19241) );
  OR2_X1 U19100 ( .A1(n19243), .A2(n19244), .ZN(n19242) );
  AND2_X1 U19101 ( .A1(n19244), .A2(n19243), .ZN(n19240) );
  AND2_X1 U19102 ( .A1(n19245), .A2(n19246), .ZN(n19243) );
  OR2_X1 U19103 ( .A1(n19247), .A2(n19248), .ZN(n19246) );
  INV_X1 U19104 ( .A(n19249), .ZN(n19248) );
  OR2_X1 U19105 ( .A1(n19249), .A2(n19250), .ZN(n19245) );
  INV_X1 U19106 ( .A(n19247), .ZN(n19250) );
  OR2_X1 U19107 ( .A1(n15321), .A2(n14969), .ZN(n18850) );
  OR2_X1 U19108 ( .A1(n19251), .A2(n19252), .ZN(n18847) );
  INV_X1 U19109 ( .A(n19253), .ZN(n19252) );
  OR2_X1 U19110 ( .A1(n19254), .A2(n19255), .ZN(n19253) );
  AND2_X1 U19111 ( .A1(n19255), .A2(n19254), .ZN(n19251) );
  AND2_X1 U19112 ( .A1(n19256), .A2(n19257), .ZN(n19254) );
  OR2_X1 U19113 ( .A1(n19258), .A2(n19259), .ZN(n19257) );
  INV_X1 U19114 ( .A(n19260), .ZN(n19259) );
  OR2_X1 U19115 ( .A1(n19260), .A2(n19261), .ZN(n19256) );
  INV_X1 U19116 ( .A(n19258), .ZN(n19261) );
  OR2_X1 U19117 ( .A1(n15355), .A2(n14969), .ZN(n18861) );
  OR2_X1 U19118 ( .A1(n19262), .A2(n19263), .ZN(n18858) );
  INV_X1 U19119 ( .A(n19264), .ZN(n19263) );
  OR2_X1 U19120 ( .A1(n19265), .A2(n19266), .ZN(n19264) );
  AND2_X1 U19121 ( .A1(n19266), .A2(n19265), .ZN(n19262) );
  AND2_X1 U19122 ( .A1(n19267), .A2(n19268), .ZN(n19265) );
  OR2_X1 U19123 ( .A1(n19269), .A2(n19270), .ZN(n19268) );
  INV_X1 U19124 ( .A(n19271), .ZN(n19270) );
  OR2_X1 U19125 ( .A1(n19271), .A2(n19272), .ZN(n19267) );
  INV_X1 U19126 ( .A(n19269), .ZN(n19272) );
  OR2_X1 U19127 ( .A1(n15389), .A2(n14969), .ZN(n18872) );
  OR2_X1 U19128 ( .A1(n19273), .A2(n19274), .ZN(n18869) );
  INV_X1 U19129 ( .A(n19275), .ZN(n19274) );
  OR2_X1 U19130 ( .A1(n19276), .A2(n19277), .ZN(n19275) );
  AND2_X1 U19131 ( .A1(n19277), .A2(n19276), .ZN(n19273) );
  AND2_X1 U19132 ( .A1(n19278), .A2(n19279), .ZN(n19276) );
  OR2_X1 U19133 ( .A1(n19280), .A2(n19281), .ZN(n19279) );
  INV_X1 U19134 ( .A(n19282), .ZN(n19281) );
  OR2_X1 U19135 ( .A1(n19282), .A2(n19283), .ZN(n19278) );
  INV_X1 U19136 ( .A(n19280), .ZN(n19283) );
  OR2_X1 U19137 ( .A1(n15423), .A2(n14969), .ZN(n18883) );
  OR2_X1 U19138 ( .A1(n19284), .A2(n19285), .ZN(n18880) );
  INV_X1 U19139 ( .A(n19286), .ZN(n19285) );
  OR2_X1 U19140 ( .A1(n19287), .A2(n19288), .ZN(n19286) );
  AND2_X1 U19141 ( .A1(n19288), .A2(n19287), .ZN(n19284) );
  AND2_X1 U19142 ( .A1(n19289), .A2(n19290), .ZN(n19287) );
  OR2_X1 U19143 ( .A1(n19291), .A2(n19292), .ZN(n19290) );
  INV_X1 U19144 ( .A(n19293), .ZN(n19292) );
  OR2_X1 U19145 ( .A1(n19293), .A2(n19294), .ZN(n19289) );
  INV_X1 U19146 ( .A(n19291), .ZN(n19294) );
  OR2_X1 U19147 ( .A1(n15457), .A2(n14969), .ZN(n18894) );
  OR2_X1 U19148 ( .A1(n19295), .A2(n19296), .ZN(n18891) );
  INV_X1 U19149 ( .A(n19297), .ZN(n19296) );
  OR2_X1 U19150 ( .A1(n19298), .A2(n19299), .ZN(n19297) );
  AND2_X1 U19151 ( .A1(n19299), .A2(n19298), .ZN(n19295) );
  AND2_X1 U19152 ( .A1(n19300), .A2(n19301), .ZN(n19298) );
  OR2_X1 U19153 ( .A1(n19302), .A2(n19303), .ZN(n19301) );
  INV_X1 U19154 ( .A(n19304), .ZN(n19303) );
  OR2_X1 U19155 ( .A1(n19304), .A2(n19305), .ZN(n19300) );
  INV_X1 U19156 ( .A(n19302), .ZN(n19305) );
  OR2_X1 U19157 ( .A1(n15491), .A2(n14969), .ZN(n18905) );
  OR2_X1 U19158 ( .A1(n19306), .A2(n19307), .ZN(n18902) );
  INV_X1 U19159 ( .A(n19308), .ZN(n19307) );
  OR2_X1 U19160 ( .A1(n19309), .A2(n19310), .ZN(n19308) );
  AND2_X1 U19161 ( .A1(n19310), .A2(n19309), .ZN(n19306) );
  AND2_X1 U19162 ( .A1(n19311), .A2(n19312), .ZN(n19309) );
  OR2_X1 U19163 ( .A1(n19313), .A2(n19314), .ZN(n19312) );
  INV_X1 U19164 ( .A(n19315), .ZN(n19314) );
  OR2_X1 U19165 ( .A1(n19315), .A2(n19316), .ZN(n19311) );
  INV_X1 U19166 ( .A(n19313), .ZN(n19316) );
  OR2_X1 U19167 ( .A1(n15525), .A2(n14969), .ZN(n18916) );
  OR2_X1 U19168 ( .A1(n19317), .A2(n19318), .ZN(n18913) );
  INV_X1 U19169 ( .A(n19319), .ZN(n19318) );
  OR2_X1 U19170 ( .A1(n19320), .A2(n19321), .ZN(n19319) );
  AND2_X1 U19171 ( .A1(n19321), .A2(n19320), .ZN(n19317) );
  AND2_X1 U19172 ( .A1(n19322), .A2(n19323), .ZN(n19320) );
  OR2_X1 U19173 ( .A1(n19324), .A2(n19325), .ZN(n19323) );
  INV_X1 U19174 ( .A(n19326), .ZN(n19325) );
  OR2_X1 U19175 ( .A1(n19326), .A2(n19327), .ZN(n19322) );
  INV_X1 U19176 ( .A(n19324), .ZN(n19327) );
  OR2_X1 U19177 ( .A1(n15559), .A2(n14969), .ZN(n18927) );
  OR2_X1 U19178 ( .A1(n19328), .A2(n19329), .ZN(n18924) );
  INV_X1 U19179 ( .A(n19330), .ZN(n19329) );
  OR2_X1 U19180 ( .A1(n19331), .A2(n19332), .ZN(n19330) );
  AND2_X1 U19181 ( .A1(n19332), .A2(n19331), .ZN(n19328) );
  AND2_X1 U19182 ( .A1(n19333), .A2(n19334), .ZN(n19331) );
  OR2_X1 U19183 ( .A1(n19335), .A2(n19336), .ZN(n19334) );
  INV_X1 U19184 ( .A(n19337), .ZN(n19336) );
  OR2_X1 U19185 ( .A1(n19337), .A2(n19338), .ZN(n19333) );
  INV_X1 U19186 ( .A(n19335), .ZN(n19338) );
  OR2_X1 U19187 ( .A1(n15593), .A2(n14969), .ZN(n18938) );
  OR2_X1 U19188 ( .A1(n19339), .A2(n19340), .ZN(n18935) );
  INV_X1 U19189 ( .A(n19341), .ZN(n19340) );
  OR2_X1 U19190 ( .A1(n19342), .A2(n19343), .ZN(n19341) );
  AND2_X1 U19191 ( .A1(n19343), .A2(n19342), .ZN(n19339) );
  AND2_X1 U19192 ( .A1(n19344), .A2(n19345), .ZN(n19342) );
  OR2_X1 U19193 ( .A1(n19346), .A2(n19347), .ZN(n19345) );
  INV_X1 U19194 ( .A(n19348), .ZN(n19347) );
  OR2_X1 U19195 ( .A1(n19348), .A2(n19349), .ZN(n19344) );
  INV_X1 U19196 ( .A(n19346), .ZN(n19349) );
  OR2_X1 U19197 ( .A1(n15638), .A2(n14969), .ZN(n18949) );
  OR2_X1 U19198 ( .A1(n19350), .A2(n19351), .ZN(n18946) );
  INV_X1 U19199 ( .A(n19352), .ZN(n19351) );
  OR2_X1 U19200 ( .A1(n19353), .A2(n19354), .ZN(n19352) );
  AND2_X1 U19201 ( .A1(n19354), .A2(n19353), .ZN(n19350) );
  AND2_X1 U19202 ( .A1(n19355), .A2(n19356), .ZN(n19353) );
  OR2_X1 U19203 ( .A1(n19357), .A2(n19358), .ZN(n19356) );
  INV_X1 U19204 ( .A(n19359), .ZN(n19358) );
  OR2_X1 U19205 ( .A1(n19359), .A2(n19360), .ZN(n19355) );
  INV_X1 U19206 ( .A(n19357), .ZN(n19360) );
  OR2_X1 U19207 ( .A1(n15672), .A2(n14969), .ZN(n18960) );
  OR2_X1 U19208 ( .A1(n19361), .A2(n19362), .ZN(n18957) );
  INV_X1 U19209 ( .A(n19363), .ZN(n19362) );
  OR2_X1 U19210 ( .A1(n19364), .A2(n19365), .ZN(n19363) );
  AND2_X1 U19211 ( .A1(n19365), .A2(n19364), .ZN(n19361) );
  AND2_X1 U19212 ( .A1(n19366), .A2(n19367), .ZN(n19364) );
  OR2_X1 U19213 ( .A1(n19368), .A2(n19369), .ZN(n19367) );
  INV_X1 U19214 ( .A(n19370), .ZN(n19369) );
  OR2_X1 U19215 ( .A1(n19370), .A2(n19371), .ZN(n19366) );
  INV_X1 U19216 ( .A(n19368), .ZN(n19371) );
  OR2_X1 U19217 ( .A1(n15706), .A2(n14969), .ZN(n18971) );
  OR2_X1 U19218 ( .A1(n19372), .A2(n19373), .ZN(n18968) );
  INV_X1 U19219 ( .A(n19374), .ZN(n19373) );
  OR2_X1 U19220 ( .A1(n19375), .A2(n19376), .ZN(n19374) );
  AND2_X1 U19221 ( .A1(n19376), .A2(n19375), .ZN(n19372) );
  AND2_X1 U19222 ( .A1(n19377), .A2(n19378), .ZN(n19375) );
  OR2_X1 U19223 ( .A1(n19379), .A2(n19380), .ZN(n19378) );
  INV_X1 U19224 ( .A(n19381), .ZN(n19380) );
  OR2_X1 U19225 ( .A1(n19381), .A2(n19382), .ZN(n19377) );
  INV_X1 U19226 ( .A(n19379), .ZN(n19382) );
  OR2_X1 U19227 ( .A1(n15740), .A2(n14969), .ZN(n18982) );
  OR2_X1 U19228 ( .A1(n19383), .A2(n19384), .ZN(n18979) );
  INV_X1 U19229 ( .A(n19385), .ZN(n19384) );
  OR2_X1 U19230 ( .A1(n19386), .A2(n19387), .ZN(n19385) );
  AND2_X1 U19231 ( .A1(n19387), .A2(n19386), .ZN(n19383) );
  AND2_X1 U19232 ( .A1(n19388), .A2(n19389), .ZN(n19386) );
  OR2_X1 U19233 ( .A1(n19390), .A2(n19391), .ZN(n19389) );
  INV_X1 U19234 ( .A(n19392), .ZN(n19391) );
  OR2_X1 U19235 ( .A1(n19392), .A2(n19393), .ZN(n19388) );
  INV_X1 U19236 ( .A(n19390), .ZN(n19393) );
  OR2_X1 U19237 ( .A1(n15774), .A2(n14969), .ZN(n18996) );
  OR2_X1 U19238 ( .A1(n19394), .A2(n19395), .ZN(n18990) );
  INV_X1 U19239 ( .A(n19396), .ZN(n19395) );
  OR2_X1 U19240 ( .A1(n19397), .A2(n19398), .ZN(n19396) );
  AND2_X1 U19241 ( .A1(n19398), .A2(n19397), .ZN(n19394) );
  AND2_X1 U19242 ( .A1(n19399), .A2(n19400), .ZN(n19397) );
  INV_X1 U19243 ( .A(n19401), .ZN(n19400) );
  AND2_X1 U19244 ( .A1(n19402), .A2(n19403), .ZN(n19401) );
  OR2_X1 U19245 ( .A1(n19403), .A2(n19402), .ZN(n19399) );
  INV_X1 U19246 ( .A(n19404), .ZN(n19402) );
  OR2_X1 U19247 ( .A1(n15808), .A2(n14969), .ZN(n19006) );
  AND2_X1 U19248 ( .A1(n19405), .A2(n19406), .ZN(n19001) );
  INV_X1 U19249 ( .A(n19407), .ZN(n19406) );
  AND2_X1 U19250 ( .A1(n19408), .A2(n19409), .ZN(n19407) );
  OR2_X1 U19251 ( .A1(n19409), .A2(n19408), .ZN(n19405) );
  OR2_X1 U19252 ( .A1(n19410), .A2(n19411), .ZN(n19408) );
  AND2_X1 U19253 ( .A1(n19412), .A2(n19413), .ZN(n19411) );
  INV_X1 U19254 ( .A(n19414), .ZN(n19412) );
  AND2_X1 U19255 ( .A1(n19415), .A2(n19414), .ZN(n19410) );
  INV_X1 U19256 ( .A(n19413), .ZN(n19415) );
  OR2_X1 U19257 ( .A1(n15842), .A2(n14969), .ZN(n19017) );
  INV_X1 U19258 ( .A(b_26_), .ZN(n14969) );
  AND2_X1 U19259 ( .A1(n19416), .A2(n19417), .ZN(n19012) );
  INV_X1 U19260 ( .A(n19418), .ZN(n19417) );
  AND2_X1 U19261 ( .A1(n19419), .A2(n19420), .ZN(n19418) );
  OR2_X1 U19262 ( .A1(n19420), .A2(n19419), .ZN(n19416) );
  OR2_X1 U19263 ( .A1(n19421), .A2(n19422), .ZN(n19419) );
  AND2_X1 U19264 ( .A1(n19423), .A2(n19424), .ZN(n19422) );
  INV_X1 U19265 ( .A(n19425), .ZN(n19423) );
  AND2_X1 U19266 ( .A1(n19426), .A2(n19425), .ZN(n19421) );
  INV_X1 U19267 ( .A(n19424), .ZN(n19426) );
  AND2_X1 U19268 ( .A1(n19427), .A2(n19428), .ZN(n16831) );
  INV_X1 U19269 ( .A(n19429), .ZN(n19428) );
  AND2_X1 U19270 ( .A1(n19430), .A2(n16845), .ZN(n19429) );
  OR2_X1 U19271 ( .A1(n16845), .A2(n19430), .ZN(n19427) );
  OR2_X1 U19272 ( .A1(n19431), .A2(n19432), .ZN(n19430) );
  AND2_X1 U19273 ( .A1(n19433), .A2(n16844), .ZN(n19432) );
  INV_X1 U19274 ( .A(n16843), .ZN(n19433) );
  AND2_X1 U19275 ( .A1(n19434), .A2(n16843), .ZN(n19431) );
  OR2_X1 U19276 ( .A1(n15842), .A2(n15003), .ZN(n16843) );
  INV_X1 U19277 ( .A(n16844), .ZN(n19434) );
  OR2_X1 U19278 ( .A1(n19435), .A2(n19436), .ZN(n16844) );
  AND2_X1 U19279 ( .A1(n19425), .A2(n19424), .ZN(n19436) );
  AND2_X1 U19280 ( .A1(n19420), .A2(n19437), .ZN(n19435) );
  OR2_X1 U19281 ( .A1(n19425), .A2(n19424), .ZN(n19437) );
  OR2_X1 U19282 ( .A1(n19438), .A2(n19439), .ZN(n19424) );
  AND2_X1 U19283 ( .A1(n19414), .A2(n19413), .ZN(n19439) );
  AND2_X1 U19284 ( .A1(n19409), .A2(n19440), .ZN(n19438) );
  OR2_X1 U19285 ( .A1(n19414), .A2(n19413), .ZN(n19440) );
  OR2_X1 U19286 ( .A1(n19441), .A2(n19442), .ZN(n19413) );
  AND2_X1 U19287 ( .A1(n19404), .A2(n19403), .ZN(n19442) );
  AND2_X1 U19288 ( .A1(n19398), .A2(n19443), .ZN(n19441) );
  OR2_X1 U19289 ( .A1(n19404), .A2(n19403), .ZN(n19443) );
  OR2_X1 U19290 ( .A1(n19444), .A2(n19445), .ZN(n19403) );
  AND2_X1 U19291 ( .A1(n19390), .A2(n19392), .ZN(n19445) );
  AND2_X1 U19292 ( .A1(n19387), .A2(n19446), .ZN(n19444) );
  OR2_X1 U19293 ( .A1(n19390), .A2(n19392), .ZN(n19446) );
  OR2_X1 U19294 ( .A1(n19447), .A2(n19448), .ZN(n19392) );
  AND2_X1 U19295 ( .A1(n19379), .A2(n19381), .ZN(n19448) );
  AND2_X1 U19296 ( .A1(n19376), .A2(n19449), .ZN(n19447) );
  OR2_X1 U19297 ( .A1(n19379), .A2(n19381), .ZN(n19449) );
  OR2_X1 U19298 ( .A1(n19450), .A2(n19451), .ZN(n19381) );
  AND2_X1 U19299 ( .A1(n19368), .A2(n19370), .ZN(n19451) );
  AND2_X1 U19300 ( .A1(n19365), .A2(n19452), .ZN(n19450) );
  OR2_X1 U19301 ( .A1(n19368), .A2(n19370), .ZN(n19452) );
  OR2_X1 U19302 ( .A1(n19453), .A2(n19454), .ZN(n19370) );
  AND2_X1 U19303 ( .A1(n19357), .A2(n19359), .ZN(n19454) );
  AND2_X1 U19304 ( .A1(n19354), .A2(n19455), .ZN(n19453) );
  OR2_X1 U19305 ( .A1(n19357), .A2(n19359), .ZN(n19455) );
  OR2_X1 U19306 ( .A1(n19456), .A2(n19457), .ZN(n19359) );
  AND2_X1 U19307 ( .A1(n19346), .A2(n19348), .ZN(n19457) );
  AND2_X1 U19308 ( .A1(n19343), .A2(n19458), .ZN(n19456) );
  OR2_X1 U19309 ( .A1(n19346), .A2(n19348), .ZN(n19458) );
  OR2_X1 U19310 ( .A1(n19459), .A2(n19460), .ZN(n19348) );
  AND2_X1 U19311 ( .A1(n19335), .A2(n19337), .ZN(n19460) );
  AND2_X1 U19312 ( .A1(n19332), .A2(n19461), .ZN(n19459) );
  OR2_X1 U19313 ( .A1(n19335), .A2(n19337), .ZN(n19461) );
  OR2_X1 U19314 ( .A1(n19462), .A2(n19463), .ZN(n19337) );
  AND2_X1 U19315 ( .A1(n19324), .A2(n19326), .ZN(n19463) );
  AND2_X1 U19316 ( .A1(n19321), .A2(n19464), .ZN(n19462) );
  OR2_X1 U19317 ( .A1(n19324), .A2(n19326), .ZN(n19464) );
  OR2_X1 U19318 ( .A1(n19465), .A2(n19466), .ZN(n19326) );
  AND2_X1 U19319 ( .A1(n19313), .A2(n19315), .ZN(n19466) );
  AND2_X1 U19320 ( .A1(n19310), .A2(n19467), .ZN(n19465) );
  OR2_X1 U19321 ( .A1(n19313), .A2(n19315), .ZN(n19467) );
  OR2_X1 U19322 ( .A1(n19468), .A2(n19469), .ZN(n19315) );
  AND2_X1 U19323 ( .A1(n19302), .A2(n19304), .ZN(n19469) );
  AND2_X1 U19324 ( .A1(n19299), .A2(n19470), .ZN(n19468) );
  OR2_X1 U19325 ( .A1(n19302), .A2(n19304), .ZN(n19470) );
  OR2_X1 U19326 ( .A1(n19471), .A2(n19472), .ZN(n19304) );
  AND2_X1 U19327 ( .A1(n19291), .A2(n19293), .ZN(n19472) );
  AND2_X1 U19328 ( .A1(n19288), .A2(n19473), .ZN(n19471) );
  OR2_X1 U19329 ( .A1(n19291), .A2(n19293), .ZN(n19473) );
  OR2_X1 U19330 ( .A1(n19474), .A2(n19475), .ZN(n19293) );
  AND2_X1 U19331 ( .A1(n19280), .A2(n19282), .ZN(n19475) );
  AND2_X1 U19332 ( .A1(n19277), .A2(n19476), .ZN(n19474) );
  OR2_X1 U19333 ( .A1(n19280), .A2(n19282), .ZN(n19476) );
  OR2_X1 U19334 ( .A1(n19477), .A2(n19478), .ZN(n19282) );
  AND2_X1 U19335 ( .A1(n19269), .A2(n19271), .ZN(n19478) );
  AND2_X1 U19336 ( .A1(n19266), .A2(n19479), .ZN(n19477) );
  OR2_X1 U19337 ( .A1(n19269), .A2(n19271), .ZN(n19479) );
  OR2_X1 U19338 ( .A1(n19480), .A2(n19481), .ZN(n19271) );
  AND2_X1 U19339 ( .A1(n19258), .A2(n19260), .ZN(n19481) );
  AND2_X1 U19340 ( .A1(n19255), .A2(n19482), .ZN(n19480) );
  OR2_X1 U19341 ( .A1(n19258), .A2(n19260), .ZN(n19482) );
  OR2_X1 U19342 ( .A1(n19483), .A2(n19484), .ZN(n19260) );
  AND2_X1 U19343 ( .A1(n19247), .A2(n19249), .ZN(n19484) );
  AND2_X1 U19344 ( .A1(n19244), .A2(n19485), .ZN(n19483) );
  OR2_X1 U19345 ( .A1(n19247), .A2(n19249), .ZN(n19485) );
  OR2_X1 U19346 ( .A1(n19486), .A2(n19487), .ZN(n19249) );
  AND2_X1 U19347 ( .A1(n19236), .A2(n19238), .ZN(n19487) );
  AND2_X1 U19348 ( .A1(n19233), .A2(n19488), .ZN(n19486) );
  OR2_X1 U19349 ( .A1(n19236), .A2(n19238), .ZN(n19488) );
  OR2_X1 U19350 ( .A1(n19489), .A2(n19490), .ZN(n19238) );
  AND2_X1 U19351 ( .A1(n19225), .A2(n19227), .ZN(n19490) );
  AND2_X1 U19352 ( .A1(n19222), .A2(n19491), .ZN(n19489) );
  OR2_X1 U19353 ( .A1(n19225), .A2(n19227), .ZN(n19491) );
  OR2_X1 U19354 ( .A1(n19492), .A2(n19493), .ZN(n19227) );
  AND2_X1 U19355 ( .A1(n19214), .A2(n19216), .ZN(n19493) );
  AND2_X1 U19356 ( .A1(n19211), .A2(n19494), .ZN(n19492) );
  OR2_X1 U19357 ( .A1(n19214), .A2(n19216), .ZN(n19494) );
  OR2_X1 U19358 ( .A1(n19495), .A2(n19496), .ZN(n19216) );
  AND2_X1 U19359 ( .A1(n19203), .A2(n19205), .ZN(n19496) );
  AND2_X1 U19360 ( .A1(n19200), .A2(n19497), .ZN(n19495) );
  OR2_X1 U19361 ( .A1(n19203), .A2(n19205), .ZN(n19497) );
  OR2_X1 U19362 ( .A1(n19498), .A2(n19499), .ZN(n19205) );
  AND2_X1 U19363 ( .A1(n19192), .A2(n19194), .ZN(n19499) );
  AND2_X1 U19364 ( .A1(n19189), .A2(n19500), .ZN(n19498) );
  OR2_X1 U19365 ( .A1(n19192), .A2(n19194), .ZN(n19500) );
  OR2_X1 U19366 ( .A1(n19501), .A2(n19502), .ZN(n19194) );
  AND2_X1 U19367 ( .A1(n19181), .A2(n19183), .ZN(n19502) );
  AND2_X1 U19368 ( .A1(n19178), .A2(n19503), .ZN(n19501) );
  OR2_X1 U19369 ( .A1(n19181), .A2(n19183), .ZN(n19503) );
  OR2_X1 U19370 ( .A1(n19504), .A2(n19505), .ZN(n19183) );
  AND2_X1 U19371 ( .A1(n15942), .A2(n19172), .ZN(n19505) );
  AND2_X1 U19372 ( .A1(n19168), .A2(n19506), .ZN(n19504) );
  OR2_X1 U19373 ( .A1(n15942), .A2(n19172), .ZN(n19506) );
  OR2_X1 U19374 ( .A1(n19507), .A2(n19508), .ZN(n19172) );
  AND2_X1 U19375 ( .A1(n19160), .A2(n19162), .ZN(n19508) );
  AND2_X1 U19376 ( .A1(n19157), .A2(n19509), .ZN(n19507) );
  OR2_X1 U19377 ( .A1(n19160), .A2(n19162), .ZN(n19509) );
  OR2_X1 U19378 ( .A1(n19510), .A2(n19511), .ZN(n19162) );
  AND2_X1 U19379 ( .A1(n19149), .A2(n19151), .ZN(n19511) );
  AND2_X1 U19380 ( .A1(n19146), .A2(n19512), .ZN(n19510) );
  OR2_X1 U19381 ( .A1(n19149), .A2(n19151), .ZN(n19512) );
  OR2_X1 U19382 ( .A1(n19513), .A2(n19514), .ZN(n19151) );
  AND2_X1 U19383 ( .A1(n19138), .A2(n19140), .ZN(n19514) );
  AND2_X1 U19384 ( .A1(n19135), .A2(n19515), .ZN(n19513) );
  OR2_X1 U19385 ( .A1(n19138), .A2(n19140), .ZN(n19515) );
  OR2_X1 U19386 ( .A1(n19516), .A2(n19517), .ZN(n19140) );
  AND2_X1 U19387 ( .A1(n19123), .A2(n19128), .ZN(n19517) );
  AND2_X1 U19388 ( .A1(n19127), .A2(n19518), .ZN(n19516) );
  OR2_X1 U19389 ( .A1(n19123), .A2(n19128), .ZN(n19518) );
  INV_X1 U19390 ( .A(n19129), .ZN(n19128) );
  AND3_X1 U19391 ( .A1(b_25_), .A2(b_24_), .A3(n15957), .ZN(n19129) );
  OR2_X1 U19392 ( .A1(n14857), .A2(n15003), .ZN(n19123) );
  INV_X1 U19393 ( .A(n19130), .ZN(n19127) );
  OR2_X1 U19394 ( .A1(n19519), .A2(n19520), .ZN(n19130) );
  AND2_X1 U19395 ( .A1(b_24_), .A2(n19521), .ZN(n19520) );
  OR2_X1 U19396 ( .A1(n19522), .A2(n16981), .ZN(n19521) );
  AND2_X1 U19397 ( .A1(a_30_), .A2(n15071), .ZN(n19522) );
  AND2_X1 U19398 ( .A1(b_23_), .A2(n19523), .ZN(n19519) );
  OR2_X1 U19399 ( .A1(n19524), .A2(n14817), .ZN(n19523) );
  AND2_X1 U19400 ( .A1(a_31_), .A2(n15037), .ZN(n19524) );
  OR2_X1 U19401 ( .A1(n14891), .A2(n15003), .ZN(n19138) );
  OR2_X1 U19402 ( .A1(n19525), .A2(n19526), .ZN(n19135) );
  AND2_X1 U19403 ( .A1(n19527), .A2(n19528), .ZN(n19526) );
  INV_X1 U19404 ( .A(n19529), .ZN(n19525) );
  OR2_X1 U19405 ( .A1(n19527), .A2(n19528), .ZN(n19529) );
  OR2_X1 U19406 ( .A1(n19530), .A2(n19531), .ZN(n19527) );
  AND2_X1 U19407 ( .A1(n19532), .A2(n19533), .ZN(n19531) );
  AND2_X1 U19408 ( .A1(n19534), .A2(n19535), .ZN(n19530) );
  OR2_X1 U19409 ( .A1(n14936), .A2(n15003), .ZN(n19149) );
  OR2_X1 U19410 ( .A1(n19536), .A2(n19537), .ZN(n19146) );
  INV_X1 U19411 ( .A(n19538), .ZN(n19537) );
  OR2_X1 U19412 ( .A1(n19539), .A2(n19540), .ZN(n19538) );
  AND2_X1 U19413 ( .A1(n19540), .A2(n19539), .ZN(n19536) );
  AND2_X1 U19414 ( .A1(n19541), .A2(n19542), .ZN(n19539) );
  OR2_X1 U19415 ( .A1(n19543), .A2(n19544), .ZN(n19542) );
  INV_X1 U19416 ( .A(n19545), .ZN(n19544) );
  OR2_X1 U19417 ( .A1(n19545), .A2(n19546), .ZN(n19541) );
  INV_X1 U19418 ( .A(n19543), .ZN(n19546) );
  OR2_X1 U19419 ( .A1(n14970), .A2(n15003), .ZN(n19160) );
  OR2_X1 U19420 ( .A1(n19547), .A2(n19548), .ZN(n19157) );
  INV_X1 U19421 ( .A(n19549), .ZN(n19548) );
  OR2_X1 U19422 ( .A1(n19550), .A2(n19551), .ZN(n19549) );
  AND2_X1 U19423 ( .A1(n19551), .A2(n19550), .ZN(n19547) );
  AND2_X1 U19424 ( .A1(n19552), .A2(n19553), .ZN(n19550) );
  OR2_X1 U19425 ( .A1(n19554), .A2(n19555), .ZN(n19553) );
  INV_X1 U19426 ( .A(n19556), .ZN(n19555) );
  OR2_X1 U19427 ( .A1(n19556), .A2(n19557), .ZN(n19552) );
  INV_X1 U19428 ( .A(n19554), .ZN(n19557) );
  OR2_X1 U19429 ( .A1(n15004), .A2(n15003), .ZN(n15942) );
  OR2_X1 U19430 ( .A1(n19558), .A2(n19559), .ZN(n19168) );
  INV_X1 U19431 ( .A(n19560), .ZN(n19559) );
  OR2_X1 U19432 ( .A1(n19561), .A2(n19562), .ZN(n19560) );
  AND2_X1 U19433 ( .A1(n19562), .A2(n19561), .ZN(n19558) );
  AND2_X1 U19434 ( .A1(n19563), .A2(n19564), .ZN(n19561) );
  OR2_X1 U19435 ( .A1(n19565), .A2(n19566), .ZN(n19564) );
  INV_X1 U19436 ( .A(n19567), .ZN(n19566) );
  OR2_X1 U19437 ( .A1(n19567), .A2(n19568), .ZN(n19563) );
  INV_X1 U19438 ( .A(n19565), .ZN(n19568) );
  OR2_X1 U19439 ( .A1(n15038), .A2(n15003), .ZN(n19181) );
  OR2_X1 U19440 ( .A1(n19569), .A2(n19570), .ZN(n19178) );
  INV_X1 U19441 ( .A(n19571), .ZN(n19570) );
  OR2_X1 U19442 ( .A1(n19572), .A2(n19573), .ZN(n19571) );
  AND2_X1 U19443 ( .A1(n19573), .A2(n19572), .ZN(n19569) );
  AND2_X1 U19444 ( .A1(n19574), .A2(n19575), .ZN(n19572) );
  OR2_X1 U19445 ( .A1(n19576), .A2(n19577), .ZN(n19575) );
  INV_X1 U19446 ( .A(n19578), .ZN(n19577) );
  OR2_X1 U19447 ( .A1(n19578), .A2(n19579), .ZN(n19574) );
  INV_X1 U19448 ( .A(n19576), .ZN(n19579) );
  OR2_X1 U19449 ( .A1(n15072), .A2(n15003), .ZN(n19192) );
  OR2_X1 U19450 ( .A1(n19580), .A2(n19581), .ZN(n19189) );
  INV_X1 U19451 ( .A(n19582), .ZN(n19581) );
  OR2_X1 U19452 ( .A1(n19583), .A2(n19584), .ZN(n19582) );
  AND2_X1 U19453 ( .A1(n19584), .A2(n19583), .ZN(n19580) );
  AND2_X1 U19454 ( .A1(n19585), .A2(n19586), .ZN(n19583) );
  OR2_X1 U19455 ( .A1(n15939), .A2(n19587), .ZN(n19586) );
  INV_X1 U19456 ( .A(n19588), .ZN(n19587) );
  OR2_X1 U19457 ( .A1(n19588), .A2(n19589), .ZN(n19585) );
  INV_X1 U19458 ( .A(n15939), .ZN(n19589) );
  OR2_X1 U19459 ( .A1(n15106), .A2(n15003), .ZN(n19203) );
  OR2_X1 U19460 ( .A1(n19590), .A2(n19591), .ZN(n19200) );
  INV_X1 U19461 ( .A(n19592), .ZN(n19591) );
  OR2_X1 U19462 ( .A1(n19593), .A2(n19594), .ZN(n19592) );
  AND2_X1 U19463 ( .A1(n19594), .A2(n19593), .ZN(n19590) );
  AND2_X1 U19464 ( .A1(n19595), .A2(n19596), .ZN(n19593) );
  OR2_X1 U19465 ( .A1(n19597), .A2(n19598), .ZN(n19596) );
  INV_X1 U19466 ( .A(n19599), .ZN(n19598) );
  OR2_X1 U19467 ( .A1(n19599), .A2(n19600), .ZN(n19595) );
  INV_X1 U19468 ( .A(n19597), .ZN(n19600) );
  OR2_X1 U19469 ( .A1(n15140), .A2(n15003), .ZN(n19214) );
  OR2_X1 U19470 ( .A1(n19601), .A2(n19602), .ZN(n19211) );
  INV_X1 U19471 ( .A(n19603), .ZN(n19602) );
  OR2_X1 U19472 ( .A1(n19604), .A2(n19605), .ZN(n19603) );
  AND2_X1 U19473 ( .A1(n19605), .A2(n19604), .ZN(n19601) );
  AND2_X1 U19474 ( .A1(n19606), .A2(n19607), .ZN(n19604) );
  OR2_X1 U19475 ( .A1(n19608), .A2(n19609), .ZN(n19607) );
  INV_X1 U19476 ( .A(n19610), .ZN(n19609) );
  OR2_X1 U19477 ( .A1(n19610), .A2(n19611), .ZN(n19606) );
  INV_X1 U19478 ( .A(n19608), .ZN(n19611) );
  OR2_X1 U19479 ( .A1(n15174), .A2(n15003), .ZN(n19225) );
  OR2_X1 U19480 ( .A1(n19612), .A2(n19613), .ZN(n19222) );
  INV_X1 U19481 ( .A(n19614), .ZN(n19613) );
  OR2_X1 U19482 ( .A1(n19615), .A2(n19616), .ZN(n19614) );
  AND2_X1 U19483 ( .A1(n19616), .A2(n19615), .ZN(n19612) );
  AND2_X1 U19484 ( .A1(n19617), .A2(n19618), .ZN(n19615) );
  OR2_X1 U19485 ( .A1(n19619), .A2(n19620), .ZN(n19618) );
  INV_X1 U19486 ( .A(n19621), .ZN(n19620) );
  OR2_X1 U19487 ( .A1(n19621), .A2(n19622), .ZN(n19617) );
  INV_X1 U19488 ( .A(n19619), .ZN(n19622) );
  OR2_X1 U19489 ( .A1(n15208), .A2(n15003), .ZN(n19236) );
  OR2_X1 U19490 ( .A1(n19623), .A2(n19624), .ZN(n19233) );
  INV_X1 U19491 ( .A(n19625), .ZN(n19624) );
  OR2_X1 U19492 ( .A1(n19626), .A2(n19627), .ZN(n19625) );
  AND2_X1 U19493 ( .A1(n19627), .A2(n19626), .ZN(n19623) );
  AND2_X1 U19494 ( .A1(n19628), .A2(n19629), .ZN(n19626) );
  OR2_X1 U19495 ( .A1(n19630), .A2(n19631), .ZN(n19629) );
  INV_X1 U19496 ( .A(n19632), .ZN(n19631) );
  OR2_X1 U19497 ( .A1(n19632), .A2(n19633), .ZN(n19628) );
  INV_X1 U19498 ( .A(n19630), .ZN(n19633) );
  OR2_X1 U19499 ( .A1(n15242), .A2(n15003), .ZN(n19247) );
  OR2_X1 U19500 ( .A1(n19634), .A2(n19635), .ZN(n19244) );
  INV_X1 U19501 ( .A(n19636), .ZN(n19635) );
  OR2_X1 U19502 ( .A1(n19637), .A2(n19638), .ZN(n19636) );
  AND2_X1 U19503 ( .A1(n19638), .A2(n19637), .ZN(n19634) );
  AND2_X1 U19504 ( .A1(n19639), .A2(n19640), .ZN(n19637) );
  OR2_X1 U19505 ( .A1(n19641), .A2(n19642), .ZN(n19640) );
  INV_X1 U19506 ( .A(n19643), .ZN(n19642) );
  OR2_X1 U19507 ( .A1(n19643), .A2(n19644), .ZN(n19639) );
  INV_X1 U19508 ( .A(n19641), .ZN(n19644) );
  OR2_X1 U19509 ( .A1(n15287), .A2(n15003), .ZN(n19258) );
  OR2_X1 U19510 ( .A1(n19645), .A2(n19646), .ZN(n19255) );
  INV_X1 U19511 ( .A(n19647), .ZN(n19646) );
  OR2_X1 U19512 ( .A1(n19648), .A2(n19649), .ZN(n19647) );
  AND2_X1 U19513 ( .A1(n19649), .A2(n19648), .ZN(n19645) );
  AND2_X1 U19514 ( .A1(n19650), .A2(n19651), .ZN(n19648) );
  OR2_X1 U19515 ( .A1(n19652), .A2(n19653), .ZN(n19651) );
  INV_X1 U19516 ( .A(n19654), .ZN(n19653) );
  OR2_X1 U19517 ( .A1(n19654), .A2(n19655), .ZN(n19650) );
  INV_X1 U19518 ( .A(n19652), .ZN(n19655) );
  OR2_X1 U19519 ( .A1(n15321), .A2(n15003), .ZN(n19269) );
  OR2_X1 U19520 ( .A1(n19656), .A2(n19657), .ZN(n19266) );
  INV_X1 U19521 ( .A(n19658), .ZN(n19657) );
  OR2_X1 U19522 ( .A1(n19659), .A2(n19660), .ZN(n19658) );
  AND2_X1 U19523 ( .A1(n19660), .A2(n19659), .ZN(n19656) );
  AND2_X1 U19524 ( .A1(n19661), .A2(n19662), .ZN(n19659) );
  OR2_X1 U19525 ( .A1(n19663), .A2(n19664), .ZN(n19662) );
  INV_X1 U19526 ( .A(n19665), .ZN(n19664) );
  OR2_X1 U19527 ( .A1(n19665), .A2(n19666), .ZN(n19661) );
  INV_X1 U19528 ( .A(n19663), .ZN(n19666) );
  OR2_X1 U19529 ( .A1(n15355), .A2(n15003), .ZN(n19280) );
  OR2_X1 U19530 ( .A1(n19667), .A2(n19668), .ZN(n19277) );
  INV_X1 U19531 ( .A(n19669), .ZN(n19668) );
  OR2_X1 U19532 ( .A1(n19670), .A2(n19671), .ZN(n19669) );
  AND2_X1 U19533 ( .A1(n19671), .A2(n19670), .ZN(n19667) );
  AND2_X1 U19534 ( .A1(n19672), .A2(n19673), .ZN(n19670) );
  OR2_X1 U19535 ( .A1(n19674), .A2(n19675), .ZN(n19673) );
  INV_X1 U19536 ( .A(n19676), .ZN(n19675) );
  OR2_X1 U19537 ( .A1(n19676), .A2(n19677), .ZN(n19672) );
  INV_X1 U19538 ( .A(n19674), .ZN(n19677) );
  OR2_X1 U19539 ( .A1(n15389), .A2(n15003), .ZN(n19291) );
  OR2_X1 U19540 ( .A1(n19678), .A2(n19679), .ZN(n19288) );
  INV_X1 U19541 ( .A(n19680), .ZN(n19679) );
  OR2_X1 U19542 ( .A1(n19681), .A2(n19682), .ZN(n19680) );
  AND2_X1 U19543 ( .A1(n19682), .A2(n19681), .ZN(n19678) );
  AND2_X1 U19544 ( .A1(n19683), .A2(n19684), .ZN(n19681) );
  OR2_X1 U19545 ( .A1(n19685), .A2(n19686), .ZN(n19684) );
  INV_X1 U19546 ( .A(n19687), .ZN(n19686) );
  OR2_X1 U19547 ( .A1(n19687), .A2(n19688), .ZN(n19683) );
  INV_X1 U19548 ( .A(n19685), .ZN(n19688) );
  OR2_X1 U19549 ( .A1(n15423), .A2(n15003), .ZN(n19302) );
  OR2_X1 U19550 ( .A1(n19689), .A2(n19690), .ZN(n19299) );
  INV_X1 U19551 ( .A(n19691), .ZN(n19690) );
  OR2_X1 U19552 ( .A1(n19692), .A2(n19693), .ZN(n19691) );
  AND2_X1 U19553 ( .A1(n19693), .A2(n19692), .ZN(n19689) );
  AND2_X1 U19554 ( .A1(n19694), .A2(n19695), .ZN(n19692) );
  OR2_X1 U19555 ( .A1(n19696), .A2(n19697), .ZN(n19695) );
  INV_X1 U19556 ( .A(n19698), .ZN(n19697) );
  OR2_X1 U19557 ( .A1(n19698), .A2(n19699), .ZN(n19694) );
  INV_X1 U19558 ( .A(n19696), .ZN(n19699) );
  OR2_X1 U19559 ( .A1(n15457), .A2(n15003), .ZN(n19313) );
  OR2_X1 U19560 ( .A1(n19700), .A2(n19701), .ZN(n19310) );
  INV_X1 U19561 ( .A(n19702), .ZN(n19701) );
  OR2_X1 U19562 ( .A1(n19703), .A2(n19704), .ZN(n19702) );
  AND2_X1 U19563 ( .A1(n19704), .A2(n19703), .ZN(n19700) );
  AND2_X1 U19564 ( .A1(n19705), .A2(n19706), .ZN(n19703) );
  OR2_X1 U19565 ( .A1(n19707), .A2(n19708), .ZN(n19706) );
  INV_X1 U19566 ( .A(n19709), .ZN(n19708) );
  OR2_X1 U19567 ( .A1(n19709), .A2(n19710), .ZN(n19705) );
  INV_X1 U19568 ( .A(n19707), .ZN(n19710) );
  OR2_X1 U19569 ( .A1(n15491), .A2(n15003), .ZN(n19324) );
  OR2_X1 U19570 ( .A1(n19711), .A2(n19712), .ZN(n19321) );
  INV_X1 U19571 ( .A(n19713), .ZN(n19712) );
  OR2_X1 U19572 ( .A1(n19714), .A2(n19715), .ZN(n19713) );
  AND2_X1 U19573 ( .A1(n19715), .A2(n19714), .ZN(n19711) );
  AND2_X1 U19574 ( .A1(n19716), .A2(n19717), .ZN(n19714) );
  OR2_X1 U19575 ( .A1(n19718), .A2(n19719), .ZN(n19717) );
  INV_X1 U19576 ( .A(n19720), .ZN(n19719) );
  OR2_X1 U19577 ( .A1(n19720), .A2(n19721), .ZN(n19716) );
  INV_X1 U19578 ( .A(n19718), .ZN(n19721) );
  OR2_X1 U19579 ( .A1(n15525), .A2(n15003), .ZN(n19335) );
  OR2_X1 U19580 ( .A1(n19722), .A2(n19723), .ZN(n19332) );
  INV_X1 U19581 ( .A(n19724), .ZN(n19723) );
  OR2_X1 U19582 ( .A1(n19725), .A2(n19726), .ZN(n19724) );
  AND2_X1 U19583 ( .A1(n19726), .A2(n19725), .ZN(n19722) );
  AND2_X1 U19584 ( .A1(n19727), .A2(n19728), .ZN(n19725) );
  OR2_X1 U19585 ( .A1(n19729), .A2(n19730), .ZN(n19728) );
  INV_X1 U19586 ( .A(n19731), .ZN(n19730) );
  OR2_X1 U19587 ( .A1(n19731), .A2(n19732), .ZN(n19727) );
  INV_X1 U19588 ( .A(n19729), .ZN(n19732) );
  OR2_X1 U19589 ( .A1(n15559), .A2(n15003), .ZN(n19346) );
  OR2_X1 U19590 ( .A1(n19733), .A2(n19734), .ZN(n19343) );
  INV_X1 U19591 ( .A(n19735), .ZN(n19734) );
  OR2_X1 U19592 ( .A1(n19736), .A2(n19737), .ZN(n19735) );
  AND2_X1 U19593 ( .A1(n19737), .A2(n19736), .ZN(n19733) );
  AND2_X1 U19594 ( .A1(n19738), .A2(n19739), .ZN(n19736) );
  OR2_X1 U19595 ( .A1(n19740), .A2(n19741), .ZN(n19739) );
  INV_X1 U19596 ( .A(n19742), .ZN(n19741) );
  OR2_X1 U19597 ( .A1(n19742), .A2(n19743), .ZN(n19738) );
  INV_X1 U19598 ( .A(n19740), .ZN(n19743) );
  OR2_X1 U19599 ( .A1(n15593), .A2(n15003), .ZN(n19357) );
  OR2_X1 U19600 ( .A1(n19744), .A2(n19745), .ZN(n19354) );
  INV_X1 U19601 ( .A(n19746), .ZN(n19745) );
  OR2_X1 U19602 ( .A1(n19747), .A2(n19748), .ZN(n19746) );
  AND2_X1 U19603 ( .A1(n19748), .A2(n19747), .ZN(n19744) );
  AND2_X1 U19604 ( .A1(n19749), .A2(n19750), .ZN(n19747) );
  OR2_X1 U19605 ( .A1(n19751), .A2(n19752), .ZN(n19750) );
  INV_X1 U19606 ( .A(n19753), .ZN(n19752) );
  OR2_X1 U19607 ( .A1(n19753), .A2(n19754), .ZN(n19749) );
  INV_X1 U19608 ( .A(n19751), .ZN(n19754) );
  OR2_X1 U19609 ( .A1(n15638), .A2(n15003), .ZN(n19368) );
  OR2_X1 U19610 ( .A1(n19755), .A2(n19756), .ZN(n19365) );
  INV_X1 U19611 ( .A(n19757), .ZN(n19756) );
  OR2_X1 U19612 ( .A1(n19758), .A2(n19759), .ZN(n19757) );
  AND2_X1 U19613 ( .A1(n19759), .A2(n19758), .ZN(n19755) );
  AND2_X1 U19614 ( .A1(n19760), .A2(n19761), .ZN(n19758) );
  OR2_X1 U19615 ( .A1(n19762), .A2(n19763), .ZN(n19761) );
  INV_X1 U19616 ( .A(n19764), .ZN(n19763) );
  OR2_X1 U19617 ( .A1(n19764), .A2(n19765), .ZN(n19760) );
  INV_X1 U19618 ( .A(n19762), .ZN(n19765) );
  OR2_X1 U19619 ( .A1(n15672), .A2(n15003), .ZN(n19379) );
  OR2_X1 U19620 ( .A1(n19766), .A2(n19767), .ZN(n19376) );
  INV_X1 U19621 ( .A(n19768), .ZN(n19767) );
  OR2_X1 U19622 ( .A1(n19769), .A2(n19770), .ZN(n19768) );
  AND2_X1 U19623 ( .A1(n19770), .A2(n19769), .ZN(n19766) );
  AND2_X1 U19624 ( .A1(n19771), .A2(n19772), .ZN(n19769) );
  OR2_X1 U19625 ( .A1(n19773), .A2(n19774), .ZN(n19772) );
  INV_X1 U19626 ( .A(n19775), .ZN(n19774) );
  OR2_X1 U19627 ( .A1(n19775), .A2(n19776), .ZN(n19771) );
  INV_X1 U19628 ( .A(n19773), .ZN(n19776) );
  OR2_X1 U19629 ( .A1(n15706), .A2(n15003), .ZN(n19390) );
  OR2_X1 U19630 ( .A1(n19777), .A2(n19778), .ZN(n19387) );
  INV_X1 U19631 ( .A(n19779), .ZN(n19778) );
  OR2_X1 U19632 ( .A1(n19780), .A2(n19781), .ZN(n19779) );
  AND2_X1 U19633 ( .A1(n19781), .A2(n19780), .ZN(n19777) );
  AND2_X1 U19634 ( .A1(n19782), .A2(n19783), .ZN(n19780) );
  OR2_X1 U19635 ( .A1(n19784), .A2(n19785), .ZN(n19783) );
  INV_X1 U19636 ( .A(n19786), .ZN(n19785) );
  OR2_X1 U19637 ( .A1(n19786), .A2(n19787), .ZN(n19782) );
  INV_X1 U19638 ( .A(n19784), .ZN(n19787) );
  OR2_X1 U19639 ( .A1(n15740), .A2(n15003), .ZN(n19404) );
  OR2_X1 U19640 ( .A1(n19788), .A2(n19789), .ZN(n19398) );
  INV_X1 U19641 ( .A(n19790), .ZN(n19789) );
  OR2_X1 U19642 ( .A1(n19791), .A2(n19792), .ZN(n19790) );
  AND2_X1 U19643 ( .A1(n19792), .A2(n19791), .ZN(n19788) );
  AND2_X1 U19644 ( .A1(n19793), .A2(n19794), .ZN(n19791) );
  INV_X1 U19645 ( .A(n19795), .ZN(n19794) );
  AND2_X1 U19646 ( .A1(n19796), .A2(n19797), .ZN(n19795) );
  OR2_X1 U19647 ( .A1(n19797), .A2(n19796), .ZN(n19793) );
  INV_X1 U19648 ( .A(n19798), .ZN(n19796) );
  OR2_X1 U19649 ( .A1(n15774), .A2(n15003), .ZN(n19414) );
  AND2_X1 U19650 ( .A1(n19799), .A2(n19800), .ZN(n19409) );
  INV_X1 U19651 ( .A(n19801), .ZN(n19800) );
  AND2_X1 U19652 ( .A1(n19802), .A2(n19803), .ZN(n19801) );
  OR2_X1 U19653 ( .A1(n19803), .A2(n19802), .ZN(n19799) );
  OR2_X1 U19654 ( .A1(n19804), .A2(n19805), .ZN(n19802) );
  AND2_X1 U19655 ( .A1(n19806), .A2(n19807), .ZN(n19805) );
  INV_X1 U19656 ( .A(n19808), .ZN(n19806) );
  AND2_X1 U19657 ( .A1(n19809), .A2(n19808), .ZN(n19804) );
  INV_X1 U19658 ( .A(n19807), .ZN(n19809) );
  OR2_X1 U19659 ( .A1(n15808), .A2(n15003), .ZN(n19425) );
  INV_X1 U19660 ( .A(b_25_), .ZN(n15003) );
  AND2_X1 U19661 ( .A1(n19810), .A2(n19811), .ZN(n19420) );
  INV_X1 U19662 ( .A(n19812), .ZN(n19811) );
  AND2_X1 U19663 ( .A1(n19813), .A2(n19814), .ZN(n19812) );
  OR2_X1 U19664 ( .A1(n19814), .A2(n19813), .ZN(n19810) );
  OR2_X1 U19665 ( .A1(n19815), .A2(n19816), .ZN(n19813) );
  AND2_X1 U19666 ( .A1(n19817), .A2(n19818), .ZN(n19816) );
  INV_X1 U19667 ( .A(n19819), .ZN(n19817) );
  AND2_X1 U19668 ( .A1(n19820), .A2(n19819), .ZN(n19815) );
  INV_X1 U19669 ( .A(n19818), .ZN(n19820) );
  AND2_X1 U19670 ( .A1(n19821), .A2(n19822), .ZN(n16845) );
  INV_X1 U19671 ( .A(n19823), .ZN(n19822) );
  AND2_X1 U19672 ( .A1(n19824), .A2(n16859), .ZN(n19823) );
  OR2_X1 U19673 ( .A1(n16859), .A2(n19824), .ZN(n19821) );
  OR2_X1 U19674 ( .A1(n19825), .A2(n19826), .ZN(n19824) );
  AND2_X1 U19675 ( .A1(n19827), .A2(n16858), .ZN(n19826) );
  INV_X1 U19676 ( .A(n16857), .ZN(n19827) );
  AND2_X1 U19677 ( .A1(n19828), .A2(n16857), .ZN(n19825) );
  OR2_X1 U19678 ( .A1(n15808), .A2(n15037), .ZN(n16857) );
  INV_X1 U19679 ( .A(n16858), .ZN(n19828) );
  OR2_X1 U19680 ( .A1(n19829), .A2(n19830), .ZN(n16858) );
  AND2_X1 U19681 ( .A1(n19819), .A2(n19818), .ZN(n19830) );
  AND2_X1 U19682 ( .A1(n19814), .A2(n19831), .ZN(n19829) );
  OR2_X1 U19683 ( .A1(n19819), .A2(n19818), .ZN(n19831) );
  OR2_X1 U19684 ( .A1(n19832), .A2(n19833), .ZN(n19818) );
  AND2_X1 U19685 ( .A1(n19808), .A2(n19807), .ZN(n19833) );
  AND2_X1 U19686 ( .A1(n19803), .A2(n19834), .ZN(n19832) );
  OR2_X1 U19687 ( .A1(n19808), .A2(n19807), .ZN(n19834) );
  OR2_X1 U19688 ( .A1(n19835), .A2(n19836), .ZN(n19807) );
  AND2_X1 U19689 ( .A1(n19798), .A2(n19797), .ZN(n19836) );
  AND2_X1 U19690 ( .A1(n19792), .A2(n19837), .ZN(n19835) );
  OR2_X1 U19691 ( .A1(n19798), .A2(n19797), .ZN(n19837) );
  OR2_X1 U19692 ( .A1(n19838), .A2(n19839), .ZN(n19797) );
  AND2_X1 U19693 ( .A1(n19784), .A2(n19786), .ZN(n19839) );
  AND2_X1 U19694 ( .A1(n19781), .A2(n19840), .ZN(n19838) );
  OR2_X1 U19695 ( .A1(n19784), .A2(n19786), .ZN(n19840) );
  OR2_X1 U19696 ( .A1(n19841), .A2(n19842), .ZN(n19786) );
  AND2_X1 U19697 ( .A1(n19773), .A2(n19775), .ZN(n19842) );
  AND2_X1 U19698 ( .A1(n19770), .A2(n19843), .ZN(n19841) );
  OR2_X1 U19699 ( .A1(n19773), .A2(n19775), .ZN(n19843) );
  OR2_X1 U19700 ( .A1(n19844), .A2(n19845), .ZN(n19775) );
  AND2_X1 U19701 ( .A1(n19762), .A2(n19764), .ZN(n19845) );
  AND2_X1 U19702 ( .A1(n19759), .A2(n19846), .ZN(n19844) );
  OR2_X1 U19703 ( .A1(n19762), .A2(n19764), .ZN(n19846) );
  OR2_X1 U19704 ( .A1(n19847), .A2(n19848), .ZN(n19764) );
  AND2_X1 U19705 ( .A1(n19751), .A2(n19753), .ZN(n19848) );
  AND2_X1 U19706 ( .A1(n19748), .A2(n19849), .ZN(n19847) );
  OR2_X1 U19707 ( .A1(n19751), .A2(n19753), .ZN(n19849) );
  OR2_X1 U19708 ( .A1(n19850), .A2(n19851), .ZN(n19753) );
  AND2_X1 U19709 ( .A1(n19740), .A2(n19742), .ZN(n19851) );
  AND2_X1 U19710 ( .A1(n19737), .A2(n19852), .ZN(n19850) );
  OR2_X1 U19711 ( .A1(n19740), .A2(n19742), .ZN(n19852) );
  OR2_X1 U19712 ( .A1(n19853), .A2(n19854), .ZN(n19742) );
  AND2_X1 U19713 ( .A1(n19729), .A2(n19731), .ZN(n19854) );
  AND2_X1 U19714 ( .A1(n19726), .A2(n19855), .ZN(n19853) );
  OR2_X1 U19715 ( .A1(n19729), .A2(n19731), .ZN(n19855) );
  OR2_X1 U19716 ( .A1(n19856), .A2(n19857), .ZN(n19731) );
  AND2_X1 U19717 ( .A1(n19718), .A2(n19720), .ZN(n19857) );
  AND2_X1 U19718 ( .A1(n19715), .A2(n19858), .ZN(n19856) );
  OR2_X1 U19719 ( .A1(n19718), .A2(n19720), .ZN(n19858) );
  OR2_X1 U19720 ( .A1(n19859), .A2(n19860), .ZN(n19720) );
  AND2_X1 U19721 ( .A1(n19707), .A2(n19709), .ZN(n19860) );
  AND2_X1 U19722 ( .A1(n19704), .A2(n19861), .ZN(n19859) );
  OR2_X1 U19723 ( .A1(n19707), .A2(n19709), .ZN(n19861) );
  OR2_X1 U19724 ( .A1(n19862), .A2(n19863), .ZN(n19709) );
  AND2_X1 U19725 ( .A1(n19696), .A2(n19698), .ZN(n19863) );
  AND2_X1 U19726 ( .A1(n19693), .A2(n19864), .ZN(n19862) );
  OR2_X1 U19727 ( .A1(n19696), .A2(n19698), .ZN(n19864) );
  OR2_X1 U19728 ( .A1(n19865), .A2(n19866), .ZN(n19698) );
  AND2_X1 U19729 ( .A1(n19685), .A2(n19687), .ZN(n19866) );
  AND2_X1 U19730 ( .A1(n19682), .A2(n19867), .ZN(n19865) );
  OR2_X1 U19731 ( .A1(n19685), .A2(n19687), .ZN(n19867) );
  OR2_X1 U19732 ( .A1(n19868), .A2(n19869), .ZN(n19687) );
  AND2_X1 U19733 ( .A1(n19674), .A2(n19676), .ZN(n19869) );
  AND2_X1 U19734 ( .A1(n19671), .A2(n19870), .ZN(n19868) );
  OR2_X1 U19735 ( .A1(n19674), .A2(n19676), .ZN(n19870) );
  OR2_X1 U19736 ( .A1(n19871), .A2(n19872), .ZN(n19676) );
  AND2_X1 U19737 ( .A1(n19663), .A2(n19665), .ZN(n19872) );
  AND2_X1 U19738 ( .A1(n19660), .A2(n19873), .ZN(n19871) );
  OR2_X1 U19739 ( .A1(n19663), .A2(n19665), .ZN(n19873) );
  OR2_X1 U19740 ( .A1(n19874), .A2(n19875), .ZN(n19665) );
  AND2_X1 U19741 ( .A1(n19652), .A2(n19654), .ZN(n19875) );
  AND2_X1 U19742 ( .A1(n19649), .A2(n19876), .ZN(n19874) );
  OR2_X1 U19743 ( .A1(n19652), .A2(n19654), .ZN(n19876) );
  OR2_X1 U19744 ( .A1(n19877), .A2(n19878), .ZN(n19654) );
  AND2_X1 U19745 ( .A1(n19641), .A2(n19643), .ZN(n19878) );
  AND2_X1 U19746 ( .A1(n19638), .A2(n19879), .ZN(n19877) );
  OR2_X1 U19747 ( .A1(n19641), .A2(n19643), .ZN(n19879) );
  OR2_X1 U19748 ( .A1(n19880), .A2(n19881), .ZN(n19643) );
  AND2_X1 U19749 ( .A1(n19630), .A2(n19632), .ZN(n19881) );
  AND2_X1 U19750 ( .A1(n19627), .A2(n19882), .ZN(n19880) );
  OR2_X1 U19751 ( .A1(n19630), .A2(n19632), .ZN(n19882) );
  OR2_X1 U19752 ( .A1(n19883), .A2(n19884), .ZN(n19632) );
  AND2_X1 U19753 ( .A1(n19619), .A2(n19621), .ZN(n19884) );
  AND2_X1 U19754 ( .A1(n19616), .A2(n19885), .ZN(n19883) );
  OR2_X1 U19755 ( .A1(n19619), .A2(n19621), .ZN(n19885) );
  OR2_X1 U19756 ( .A1(n19886), .A2(n19887), .ZN(n19621) );
  AND2_X1 U19757 ( .A1(n19608), .A2(n19610), .ZN(n19887) );
  AND2_X1 U19758 ( .A1(n19605), .A2(n19888), .ZN(n19886) );
  OR2_X1 U19759 ( .A1(n19608), .A2(n19610), .ZN(n19888) );
  OR2_X1 U19760 ( .A1(n19889), .A2(n19890), .ZN(n19610) );
  AND2_X1 U19761 ( .A1(n19597), .A2(n19599), .ZN(n19890) );
  AND2_X1 U19762 ( .A1(n19594), .A2(n19891), .ZN(n19889) );
  OR2_X1 U19763 ( .A1(n19597), .A2(n19599), .ZN(n19891) );
  OR2_X1 U19764 ( .A1(n19892), .A2(n19893), .ZN(n19599) );
  AND2_X1 U19765 ( .A1(n15939), .A2(n19588), .ZN(n19893) );
  AND2_X1 U19766 ( .A1(n19584), .A2(n19894), .ZN(n19892) );
  OR2_X1 U19767 ( .A1(n15939), .A2(n19588), .ZN(n19894) );
  OR2_X1 U19768 ( .A1(n19895), .A2(n19896), .ZN(n19588) );
  AND2_X1 U19769 ( .A1(n19576), .A2(n19578), .ZN(n19896) );
  AND2_X1 U19770 ( .A1(n19573), .A2(n19897), .ZN(n19895) );
  OR2_X1 U19771 ( .A1(n19576), .A2(n19578), .ZN(n19897) );
  OR2_X1 U19772 ( .A1(n19898), .A2(n19899), .ZN(n19578) );
  AND2_X1 U19773 ( .A1(n19565), .A2(n19567), .ZN(n19899) );
  AND2_X1 U19774 ( .A1(n19562), .A2(n19900), .ZN(n19898) );
  OR2_X1 U19775 ( .A1(n19565), .A2(n19567), .ZN(n19900) );
  OR2_X1 U19776 ( .A1(n19901), .A2(n19902), .ZN(n19567) );
  AND2_X1 U19777 ( .A1(n19554), .A2(n19556), .ZN(n19902) );
  AND2_X1 U19778 ( .A1(n19551), .A2(n19903), .ZN(n19901) );
  OR2_X1 U19779 ( .A1(n19554), .A2(n19556), .ZN(n19903) );
  OR2_X1 U19780 ( .A1(n19904), .A2(n19905), .ZN(n19556) );
  AND2_X1 U19781 ( .A1(n19543), .A2(n19545), .ZN(n19905) );
  AND2_X1 U19782 ( .A1(n19540), .A2(n19906), .ZN(n19904) );
  OR2_X1 U19783 ( .A1(n19543), .A2(n19545), .ZN(n19906) );
  OR2_X1 U19784 ( .A1(n19907), .A2(n19908), .ZN(n19545) );
  AND2_X1 U19785 ( .A1(n19528), .A2(n19533), .ZN(n19908) );
  AND2_X1 U19786 ( .A1(n19532), .A2(n19909), .ZN(n19907) );
  OR2_X1 U19787 ( .A1(n19528), .A2(n19533), .ZN(n19909) );
  INV_X1 U19788 ( .A(n19534), .ZN(n19533) );
  AND3_X1 U19789 ( .A1(b_24_), .A2(b_23_), .A3(n15957), .ZN(n19534) );
  OR2_X1 U19790 ( .A1(n14857), .A2(n15037), .ZN(n19528) );
  INV_X1 U19791 ( .A(n19535), .ZN(n19532) );
  OR2_X1 U19792 ( .A1(n19910), .A2(n19911), .ZN(n19535) );
  AND2_X1 U19793 ( .A1(b_23_), .A2(n19912), .ZN(n19911) );
  OR2_X1 U19794 ( .A1(n19913), .A2(n16981), .ZN(n19912) );
  AND2_X1 U19795 ( .A1(a_30_), .A2(n15105), .ZN(n19913) );
  AND2_X1 U19796 ( .A1(b_22_), .A2(n19914), .ZN(n19910) );
  OR2_X1 U19797 ( .A1(n19915), .A2(n14817), .ZN(n19914) );
  AND2_X1 U19798 ( .A1(a_31_), .A2(n15071), .ZN(n19915) );
  OR2_X1 U19799 ( .A1(n14891), .A2(n15037), .ZN(n19543) );
  OR2_X1 U19800 ( .A1(n19916), .A2(n19917), .ZN(n19540) );
  AND2_X1 U19801 ( .A1(n19918), .A2(n19919), .ZN(n19917) );
  INV_X1 U19802 ( .A(n19920), .ZN(n19916) );
  OR2_X1 U19803 ( .A1(n19918), .A2(n19919), .ZN(n19920) );
  OR2_X1 U19804 ( .A1(n19921), .A2(n19922), .ZN(n19918) );
  AND2_X1 U19805 ( .A1(n19923), .A2(n19924), .ZN(n19922) );
  AND2_X1 U19806 ( .A1(n19925), .A2(n19926), .ZN(n19921) );
  OR2_X1 U19807 ( .A1(n14936), .A2(n15037), .ZN(n19554) );
  OR2_X1 U19808 ( .A1(n19927), .A2(n19928), .ZN(n19551) );
  INV_X1 U19809 ( .A(n19929), .ZN(n19928) );
  OR2_X1 U19810 ( .A1(n19930), .A2(n19931), .ZN(n19929) );
  AND2_X1 U19811 ( .A1(n19931), .A2(n19930), .ZN(n19927) );
  AND2_X1 U19812 ( .A1(n19932), .A2(n19933), .ZN(n19930) );
  OR2_X1 U19813 ( .A1(n19934), .A2(n19935), .ZN(n19933) );
  INV_X1 U19814 ( .A(n19936), .ZN(n19935) );
  OR2_X1 U19815 ( .A1(n19936), .A2(n19937), .ZN(n19932) );
  INV_X1 U19816 ( .A(n19934), .ZN(n19937) );
  OR2_X1 U19817 ( .A1(n14970), .A2(n15037), .ZN(n19565) );
  OR2_X1 U19818 ( .A1(n19938), .A2(n19939), .ZN(n19562) );
  INV_X1 U19819 ( .A(n19940), .ZN(n19939) );
  OR2_X1 U19820 ( .A1(n19941), .A2(n19942), .ZN(n19940) );
  AND2_X1 U19821 ( .A1(n19942), .A2(n19941), .ZN(n19938) );
  AND2_X1 U19822 ( .A1(n19943), .A2(n19944), .ZN(n19941) );
  OR2_X1 U19823 ( .A1(n19945), .A2(n19946), .ZN(n19944) );
  INV_X1 U19824 ( .A(n19947), .ZN(n19946) );
  OR2_X1 U19825 ( .A1(n19947), .A2(n19948), .ZN(n19943) );
  INV_X1 U19826 ( .A(n19945), .ZN(n19948) );
  OR2_X1 U19827 ( .A1(n15004), .A2(n15037), .ZN(n19576) );
  OR2_X1 U19828 ( .A1(n19949), .A2(n19950), .ZN(n19573) );
  INV_X1 U19829 ( .A(n19951), .ZN(n19950) );
  OR2_X1 U19830 ( .A1(n19952), .A2(n19953), .ZN(n19951) );
  AND2_X1 U19831 ( .A1(n19953), .A2(n19952), .ZN(n19949) );
  AND2_X1 U19832 ( .A1(n19954), .A2(n19955), .ZN(n19952) );
  OR2_X1 U19833 ( .A1(n19956), .A2(n19957), .ZN(n19955) );
  INV_X1 U19834 ( .A(n19958), .ZN(n19957) );
  OR2_X1 U19835 ( .A1(n19958), .A2(n19959), .ZN(n19954) );
  INV_X1 U19836 ( .A(n19956), .ZN(n19959) );
  OR2_X1 U19837 ( .A1(n15038), .A2(n15037), .ZN(n15939) );
  OR2_X1 U19838 ( .A1(n19960), .A2(n19961), .ZN(n19584) );
  INV_X1 U19839 ( .A(n19962), .ZN(n19961) );
  OR2_X1 U19840 ( .A1(n19963), .A2(n19964), .ZN(n19962) );
  AND2_X1 U19841 ( .A1(n19964), .A2(n19963), .ZN(n19960) );
  AND2_X1 U19842 ( .A1(n19965), .A2(n19966), .ZN(n19963) );
  OR2_X1 U19843 ( .A1(n19967), .A2(n19968), .ZN(n19966) );
  INV_X1 U19844 ( .A(n19969), .ZN(n19968) );
  OR2_X1 U19845 ( .A1(n19969), .A2(n19970), .ZN(n19965) );
  INV_X1 U19846 ( .A(n19967), .ZN(n19970) );
  OR2_X1 U19847 ( .A1(n15072), .A2(n15037), .ZN(n19597) );
  OR2_X1 U19848 ( .A1(n19971), .A2(n19972), .ZN(n19594) );
  INV_X1 U19849 ( .A(n19973), .ZN(n19972) );
  OR2_X1 U19850 ( .A1(n19974), .A2(n19975), .ZN(n19973) );
  AND2_X1 U19851 ( .A1(n19975), .A2(n19974), .ZN(n19971) );
  AND2_X1 U19852 ( .A1(n19976), .A2(n19977), .ZN(n19974) );
  OR2_X1 U19853 ( .A1(n19978), .A2(n19979), .ZN(n19977) );
  INV_X1 U19854 ( .A(n19980), .ZN(n19979) );
  OR2_X1 U19855 ( .A1(n19980), .A2(n19981), .ZN(n19976) );
  INV_X1 U19856 ( .A(n19978), .ZN(n19981) );
  OR2_X1 U19857 ( .A1(n15106), .A2(n15037), .ZN(n19608) );
  OR2_X1 U19858 ( .A1(n19982), .A2(n19983), .ZN(n19605) );
  INV_X1 U19859 ( .A(n19984), .ZN(n19983) );
  OR2_X1 U19860 ( .A1(n19985), .A2(n19986), .ZN(n19984) );
  AND2_X1 U19861 ( .A1(n19986), .A2(n19985), .ZN(n19982) );
  AND2_X1 U19862 ( .A1(n19987), .A2(n19988), .ZN(n19985) );
  OR2_X1 U19863 ( .A1(n15936), .A2(n19989), .ZN(n19988) );
  INV_X1 U19864 ( .A(n19990), .ZN(n19989) );
  OR2_X1 U19865 ( .A1(n19990), .A2(n19991), .ZN(n19987) );
  INV_X1 U19866 ( .A(n15936), .ZN(n19991) );
  OR2_X1 U19867 ( .A1(n15140), .A2(n15037), .ZN(n19619) );
  OR2_X1 U19868 ( .A1(n19992), .A2(n19993), .ZN(n19616) );
  INV_X1 U19869 ( .A(n19994), .ZN(n19993) );
  OR2_X1 U19870 ( .A1(n19995), .A2(n19996), .ZN(n19994) );
  AND2_X1 U19871 ( .A1(n19996), .A2(n19995), .ZN(n19992) );
  AND2_X1 U19872 ( .A1(n19997), .A2(n19998), .ZN(n19995) );
  OR2_X1 U19873 ( .A1(n19999), .A2(n20000), .ZN(n19998) );
  INV_X1 U19874 ( .A(n20001), .ZN(n20000) );
  OR2_X1 U19875 ( .A1(n20001), .A2(n20002), .ZN(n19997) );
  INV_X1 U19876 ( .A(n19999), .ZN(n20002) );
  OR2_X1 U19877 ( .A1(n15174), .A2(n15037), .ZN(n19630) );
  OR2_X1 U19878 ( .A1(n20003), .A2(n20004), .ZN(n19627) );
  INV_X1 U19879 ( .A(n20005), .ZN(n20004) );
  OR2_X1 U19880 ( .A1(n20006), .A2(n20007), .ZN(n20005) );
  AND2_X1 U19881 ( .A1(n20007), .A2(n20006), .ZN(n20003) );
  AND2_X1 U19882 ( .A1(n20008), .A2(n20009), .ZN(n20006) );
  OR2_X1 U19883 ( .A1(n20010), .A2(n20011), .ZN(n20009) );
  INV_X1 U19884 ( .A(n20012), .ZN(n20011) );
  OR2_X1 U19885 ( .A1(n20012), .A2(n20013), .ZN(n20008) );
  INV_X1 U19886 ( .A(n20010), .ZN(n20013) );
  OR2_X1 U19887 ( .A1(n15208), .A2(n15037), .ZN(n19641) );
  OR2_X1 U19888 ( .A1(n20014), .A2(n20015), .ZN(n19638) );
  INV_X1 U19889 ( .A(n20016), .ZN(n20015) );
  OR2_X1 U19890 ( .A1(n20017), .A2(n20018), .ZN(n20016) );
  AND2_X1 U19891 ( .A1(n20018), .A2(n20017), .ZN(n20014) );
  AND2_X1 U19892 ( .A1(n20019), .A2(n20020), .ZN(n20017) );
  OR2_X1 U19893 ( .A1(n20021), .A2(n20022), .ZN(n20020) );
  INV_X1 U19894 ( .A(n20023), .ZN(n20022) );
  OR2_X1 U19895 ( .A1(n20023), .A2(n20024), .ZN(n20019) );
  INV_X1 U19896 ( .A(n20021), .ZN(n20024) );
  OR2_X1 U19897 ( .A1(n15242), .A2(n15037), .ZN(n19652) );
  OR2_X1 U19898 ( .A1(n20025), .A2(n20026), .ZN(n19649) );
  INV_X1 U19899 ( .A(n20027), .ZN(n20026) );
  OR2_X1 U19900 ( .A1(n20028), .A2(n20029), .ZN(n20027) );
  AND2_X1 U19901 ( .A1(n20029), .A2(n20028), .ZN(n20025) );
  AND2_X1 U19902 ( .A1(n20030), .A2(n20031), .ZN(n20028) );
  OR2_X1 U19903 ( .A1(n20032), .A2(n20033), .ZN(n20031) );
  INV_X1 U19904 ( .A(n20034), .ZN(n20033) );
  OR2_X1 U19905 ( .A1(n20034), .A2(n20035), .ZN(n20030) );
  INV_X1 U19906 ( .A(n20032), .ZN(n20035) );
  OR2_X1 U19907 ( .A1(n15287), .A2(n15037), .ZN(n19663) );
  OR2_X1 U19908 ( .A1(n20036), .A2(n20037), .ZN(n19660) );
  INV_X1 U19909 ( .A(n20038), .ZN(n20037) );
  OR2_X1 U19910 ( .A1(n20039), .A2(n20040), .ZN(n20038) );
  AND2_X1 U19911 ( .A1(n20040), .A2(n20039), .ZN(n20036) );
  AND2_X1 U19912 ( .A1(n20041), .A2(n20042), .ZN(n20039) );
  OR2_X1 U19913 ( .A1(n20043), .A2(n20044), .ZN(n20042) );
  INV_X1 U19914 ( .A(n20045), .ZN(n20044) );
  OR2_X1 U19915 ( .A1(n20045), .A2(n20046), .ZN(n20041) );
  INV_X1 U19916 ( .A(n20043), .ZN(n20046) );
  OR2_X1 U19917 ( .A1(n15321), .A2(n15037), .ZN(n19674) );
  OR2_X1 U19918 ( .A1(n20047), .A2(n20048), .ZN(n19671) );
  INV_X1 U19919 ( .A(n20049), .ZN(n20048) );
  OR2_X1 U19920 ( .A1(n20050), .A2(n20051), .ZN(n20049) );
  AND2_X1 U19921 ( .A1(n20051), .A2(n20050), .ZN(n20047) );
  AND2_X1 U19922 ( .A1(n20052), .A2(n20053), .ZN(n20050) );
  OR2_X1 U19923 ( .A1(n20054), .A2(n20055), .ZN(n20053) );
  INV_X1 U19924 ( .A(n20056), .ZN(n20055) );
  OR2_X1 U19925 ( .A1(n20056), .A2(n20057), .ZN(n20052) );
  INV_X1 U19926 ( .A(n20054), .ZN(n20057) );
  OR2_X1 U19927 ( .A1(n15355), .A2(n15037), .ZN(n19685) );
  OR2_X1 U19928 ( .A1(n20058), .A2(n20059), .ZN(n19682) );
  INV_X1 U19929 ( .A(n20060), .ZN(n20059) );
  OR2_X1 U19930 ( .A1(n20061), .A2(n20062), .ZN(n20060) );
  AND2_X1 U19931 ( .A1(n20062), .A2(n20061), .ZN(n20058) );
  AND2_X1 U19932 ( .A1(n20063), .A2(n20064), .ZN(n20061) );
  OR2_X1 U19933 ( .A1(n20065), .A2(n20066), .ZN(n20064) );
  INV_X1 U19934 ( .A(n20067), .ZN(n20066) );
  OR2_X1 U19935 ( .A1(n20067), .A2(n20068), .ZN(n20063) );
  INV_X1 U19936 ( .A(n20065), .ZN(n20068) );
  OR2_X1 U19937 ( .A1(n15389), .A2(n15037), .ZN(n19696) );
  OR2_X1 U19938 ( .A1(n20069), .A2(n20070), .ZN(n19693) );
  INV_X1 U19939 ( .A(n20071), .ZN(n20070) );
  OR2_X1 U19940 ( .A1(n20072), .A2(n20073), .ZN(n20071) );
  AND2_X1 U19941 ( .A1(n20073), .A2(n20072), .ZN(n20069) );
  AND2_X1 U19942 ( .A1(n20074), .A2(n20075), .ZN(n20072) );
  OR2_X1 U19943 ( .A1(n20076), .A2(n20077), .ZN(n20075) );
  INV_X1 U19944 ( .A(n20078), .ZN(n20077) );
  OR2_X1 U19945 ( .A1(n20078), .A2(n20079), .ZN(n20074) );
  INV_X1 U19946 ( .A(n20076), .ZN(n20079) );
  OR2_X1 U19947 ( .A1(n15423), .A2(n15037), .ZN(n19707) );
  OR2_X1 U19948 ( .A1(n20080), .A2(n20081), .ZN(n19704) );
  INV_X1 U19949 ( .A(n20082), .ZN(n20081) );
  OR2_X1 U19950 ( .A1(n20083), .A2(n20084), .ZN(n20082) );
  AND2_X1 U19951 ( .A1(n20084), .A2(n20083), .ZN(n20080) );
  AND2_X1 U19952 ( .A1(n20085), .A2(n20086), .ZN(n20083) );
  OR2_X1 U19953 ( .A1(n20087), .A2(n20088), .ZN(n20086) );
  INV_X1 U19954 ( .A(n20089), .ZN(n20088) );
  OR2_X1 U19955 ( .A1(n20089), .A2(n20090), .ZN(n20085) );
  INV_X1 U19956 ( .A(n20087), .ZN(n20090) );
  OR2_X1 U19957 ( .A1(n15457), .A2(n15037), .ZN(n19718) );
  OR2_X1 U19958 ( .A1(n20091), .A2(n20092), .ZN(n19715) );
  INV_X1 U19959 ( .A(n20093), .ZN(n20092) );
  OR2_X1 U19960 ( .A1(n20094), .A2(n20095), .ZN(n20093) );
  AND2_X1 U19961 ( .A1(n20095), .A2(n20094), .ZN(n20091) );
  AND2_X1 U19962 ( .A1(n20096), .A2(n20097), .ZN(n20094) );
  OR2_X1 U19963 ( .A1(n20098), .A2(n20099), .ZN(n20097) );
  INV_X1 U19964 ( .A(n20100), .ZN(n20099) );
  OR2_X1 U19965 ( .A1(n20100), .A2(n20101), .ZN(n20096) );
  INV_X1 U19966 ( .A(n20098), .ZN(n20101) );
  OR2_X1 U19967 ( .A1(n15491), .A2(n15037), .ZN(n19729) );
  OR2_X1 U19968 ( .A1(n20102), .A2(n20103), .ZN(n19726) );
  INV_X1 U19969 ( .A(n20104), .ZN(n20103) );
  OR2_X1 U19970 ( .A1(n20105), .A2(n20106), .ZN(n20104) );
  AND2_X1 U19971 ( .A1(n20106), .A2(n20105), .ZN(n20102) );
  AND2_X1 U19972 ( .A1(n20107), .A2(n20108), .ZN(n20105) );
  OR2_X1 U19973 ( .A1(n20109), .A2(n20110), .ZN(n20108) );
  INV_X1 U19974 ( .A(n20111), .ZN(n20110) );
  OR2_X1 U19975 ( .A1(n20111), .A2(n20112), .ZN(n20107) );
  INV_X1 U19976 ( .A(n20109), .ZN(n20112) );
  OR2_X1 U19977 ( .A1(n15525), .A2(n15037), .ZN(n19740) );
  OR2_X1 U19978 ( .A1(n20113), .A2(n20114), .ZN(n19737) );
  INV_X1 U19979 ( .A(n20115), .ZN(n20114) );
  OR2_X1 U19980 ( .A1(n20116), .A2(n20117), .ZN(n20115) );
  AND2_X1 U19981 ( .A1(n20117), .A2(n20116), .ZN(n20113) );
  AND2_X1 U19982 ( .A1(n20118), .A2(n20119), .ZN(n20116) );
  OR2_X1 U19983 ( .A1(n20120), .A2(n20121), .ZN(n20119) );
  INV_X1 U19984 ( .A(n20122), .ZN(n20121) );
  OR2_X1 U19985 ( .A1(n20122), .A2(n20123), .ZN(n20118) );
  INV_X1 U19986 ( .A(n20120), .ZN(n20123) );
  OR2_X1 U19987 ( .A1(n15559), .A2(n15037), .ZN(n19751) );
  OR2_X1 U19988 ( .A1(n20124), .A2(n20125), .ZN(n19748) );
  INV_X1 U19989 ( .A(n20126), .ZN(n20125) );
  OR2_X1 U19990 ( .A1(n20127), .A2(n20128), .ZN(n20126) );
  AND2_X1 U19991 ( .A1(n20128), .A2(n20127), .ZN(n20124) );
  AND2_X1 U19992 ( .A1(n20129), .A2(n20130), .ZN(n20127) );
  OR2_X1 U19993 ( .A1(n20131), .A2(n20132), .ZN(n20130) );
  INV_X1 U19994 ( .A(n20133), .ZN(n20132) );
  OR2_X1 U19995 ( .A1(n20133), .A2(n20134), .ZN(n20129) );
  INV_X1 U19996 ( .A(n20131), .ZN(n20134) );
  OR2_X1 U19997 ( .A1(n15593), .A2(n15037), .ZN(n19762) );
  OR2_X1 U19998 ( .A1(n20135), .A2(n20136), .ZN(n19759) );
  INV_X1 U19999 ( .A(n20137), .ZN(n20136) );
  OR2_X1 U20000 ( .A1(n20138), .A2(n20139), .ZN(n20137) );
  AND2_X1 U20001 ( .A1(n20139), .A2(n20138), .ZN(n20135) );
  AND2_X1 U20002 ( .A1(n20140), .A2(n20141), .ZN(n20138) );
  OR2_X1 U20003 ( .A1(n20142), .A2(n20143), .ZN(n20141) );
  INV_X1 U20004 ( .A(n20144), .ZN(n20143) );
  OR2_X1 U20005 ( .A1(n20144), .A2(n20145), .ZN(n20140) );
  INV_X1 U20006 ( .A(n20142), .ZN(n20145) );
  OR2_X1 U20007 ( .A1(n15638), .A2(n15037), .ZN(n19773) );
  OR2_X1 U20008 ( .A1(n20146), .A2(n20147), .ZN(n19770) );
  INV_X1 U20009 ( .A(n20148), .ZN(n20147) );
  OR2_X1 U20010 ( .A1(n20149), .A2(n20150), .ZN(n20148) );
  AND2_X1 U20011 ( .A1(n20150), .A2(n20149), .ZN(n20146) );
  AND2_X1 U20012 ( .A1(n20151), .A2(n20152), .ZN(n20149) );
  OR2_X1 U20013 ( .A1(n20153), .A2(n20154), .ZN(n20152) );
  INV_X1 U20014 ( .A(n20155), .ZN(n20154) );
  OR2_X1 U20015 ( .A1(n20155), .A2(n20156), .ZN(n20151) );
  INV_X1 U20016 ( .A(n20153), .ZN(n20156) );
  OR2_X1 U20017 ( .A1(n15672), .A2(n15037), .ZN(n19784) );
  OR2_X1 U20018 ( .A1(n20157), .A2(n20158), .ZN(n19781) );
  INV_X1 U20019 ( .A(n20159), .ZN(n20158) );
  OR2_X1 U20020 ( .A1(n20160), .A2(n20161), .ZN(n20159) );
  AND2_X1 U20021 ( .A1(n20161), .A2(n20160), .ZN(n20157) );
  AND2_X1 U20022 ( .A1(n20162), .A2(n20163), .ZN(n20160) );
  OR2_X1 U20023 ( .A1(n20164), .A2(n20165), .ZN(n20163) );
  INV_X1 U20024 ( .A(n20166), .ZN(n20165) );
  OR2_X1 U20025 ( .A1(n20166), .A2(n20167), .ZN(n20162) );
  INV_X1 U20026 ( .A(n20164), .ZN(n20167) );
  OR2_X1 U20027 ( .A1(n15706), .A2(n15037), .ZN(n19798) );
  OR2_X1 U20028 ( .A1(n20168), .A2(n20169), .ZN(n19792) );
  INV_X1 U20029 ( .A(n20170), .ZN(n20169) );
  OR2_X1 U20030 ( .A1(n20171), .A2(n20172), .ZN(n20170) );
  AND2_X1 U20031 ( .A1(n20172), .A2(n20171), .ZN(n20168) );
  AND2_X1 U20032 ( .A1(n20173), .A2(n20174), .ZN(n20171) );
  INV_X1 U20033 ( .A(n20175), .ZN(n20174) );
  AND2_X1 U20034 ( .A1(n20176), .A2(n20177), .ZN(n20175) );
  OR2_X1 U20035 ( .A1(n20177), .A2(n20176), .ZN(n20173) );
  INV_X1 U20036 ( .A(n20178), .ZN(n20176) );
  OR2_X1 U20037 ( .A1(n15740), .A2(n15037), .ZN(n19808) );
  AND2_X1 U20038 ( .A1(n20179), .A2(n20180), .ZN(n19803) );
  INV_X1 U20039 ( .A(n20181), .ZN(n20180) );
  AND2_X1 U20040 ( .A1(n20182), .A2(n20183), .ZN(n20181) );
  OR2_X1 U20041 ( .A1(n20183), .A2(n20182), .ZN(n20179) );
  OR2_X1 U20042 ( .A1(n20184), .A2(n20185), .ZN(n20182) );
  AND2_X1 U20043 ( .A1(n20186), .A2(n20187), .ZN(n20185) );
  INV_X1 U20044 ( .A(n20188), .ZN(n20186) );
  AND2_X1 U20045 ( .A1(n20189), .A2(n20188), .ZN(n20184) );
  INV_X1 U20046 ( .A(n20187), .ZN(n20189) );
  OR2_X1 U20047 ( .A1(n15774), .A2(n15037), .ZN(n19819) );
  INV_X1 U20048 ( .A(b_24_), .ZN(n15037) );
  AND2_X1 U20049 ( .A1(n20190), .A2(n20191), .ZN(n19814) );
  INV_X1 U20050 ( .A(n20192), .ZN(n20191) );
  AND2_X1 U20051 ( .A1(n20193), .A2(n20194), .ZN(n20192) );
  OR2_X1 U20052 ( .A1(n20194), .A2(n20193), .ZN(n20190) );
  OR2_X1 U20053 ( .A1(n20195), .A2(n20196), .ZN(n20193) );
  AND2_X1 U20054 ( .A1(n20197), .A2(n20198), .ZN(n20196) );
  INV_X1 U20055 ( .A(n20199), .ZN(n20197) );
  AND2_X1 U20056 ( .A1(n20200), .A2(n20199), .ZN(n20195) );
  INV_X1 U20057 ( .A(n20198), .ZN(n20200) );
  AND2_X1 U20058 ( .A1(n20201), .A2(n20202), .ZN(n16859) );
  INV_X1 U20059 ( .A(n20203), .ZN(n20202) );
  AND2_X1 U20060 ( .A1(n20204), .A2(n20205), .ZN(n20203) );
  OR2_X1 U20061 ( .A1(n20205), .A2(n20204), .ZN(n20201) );
  OR2_X1 U20062 ( .A1(n20206), .A2(n20207), .ZN(n20204) );
  AND2_X1 U20063 ( .A1(n20208), .A2(n20209), .ZN(n20207) );
  INV_X1 U20064 ( .A(n20210), .ZN(n20208) );
  AND2_X1 U20065 ( .A1(n20211), .A2(n20210), .ZN(n20206) );
  INV_X1 U20066 ( .A(n20209), .ZN(n20211) );
  OR2_X1 U20067 ( .A1(n20212), .A2(n16743), .ZN(n16062) );
  OR2_X1 U20068 ( .A1(n20213), .A2(n20214), .ZN(n16743) );
  AND2_X1 U20069 ( .A1(n16703), .A2(n20215), .ZN(n20214) );
  INV_X1 U20070 ( .A(n20216), .ZN(n16703) );
  AND2_X1 U20071 ( .A1(n20216), .A2(n16705), .ZN(n20213) );
  INV_X1 U20072 ( .A(n20215), .ZN(n16705) );
  OR2_X1 U20073 ( .A1(n20217), .A2(n20218), .ZN(n20215) );
  AND2_X1 U20074 ( .A1(n20219), .A2(n20220), .ZN(n20218) );
  AND2_X1 U20075 ( .A1(n20221), .A2(n20222), .ZN(n20217) );
  OR2_X1 U20076 ( .A1(n20220), .A2(n20219), .ZN(n20222) );
  AND2_X1 U20077 ( .A1(n20223), .A2(n20224), .ZN(n20216) );
  INV_X1 U20078 ( .A(n20225), .ZN(n20224) );
  AND2_X1 U20079 ( .A1(n20226), .A2(n16715), .ZN(n20225) );
  OR2_X1 U20080 ( .A1(n16715), .A2(n20226), .ZN(n20223) );
  OR2_X1 U20081 ( .A1(n20227), .A2(n20228), .ZN(n20226) );
  AND2_X1 U20082 ( .A1(n20229), .A2(n16714), .ZN(n20228) );
  INV_X1 U20083 ( .A(n16713), .ZN(n20229) );
  AND2_X1 U20084 ( .A1(n20230), .A2(n16713), .ZN(n20227) );
  OR2_X1 U20085 ( .A1(n16512), .A2(n15139), .ZN(n16713) );
  INV_X1 U20086 ( .A(n16714), .ZN(n20230) );
  OR2_X1 U20087 ( .A1(n20231), .A2(n20232), .ZN(n16714) );
  AND2_X1 U20088 ( .A1(n20233), .A2(n20234), .ZN(n20232) );
  AND2_X1 U20089 ( .A1(n20235), .A2(n20236), .ZN(n20231) );
  OR2_X1 U20090 ( .A1(n20233), .A2(n20234), .ZN(n20236) );
  AND2_X1 U20091 ( .A1(n20237), .A2(n20238), .ZN(n16715) );
  INV_X1 U20092 ( .A(n20239), .ZN(n20238) );
  AND2_X1 U20093 ( .A1(n20240), .A2(n16729), .ZN(n20239) );
  OR2_X1 U20094 ( .A1(n16729), .A2(n20240), .ZN(n20237) );
  OR2_X1 U20095 ( .A1(n20241), .A2(n20242), .ZN(n20240) );
  AND2_X1 U20096 ( .A1(n20243), .A2(n16728), .ZN(n20242) );
  INV_X1 U20097 ( .A(n16727), .ZN(n20243) );
  AND2_X1 U20098 ( .A1(n20244), .A2(n16727), .ZN(n20241) );
  OR2_X1 U20099 ( .A1(n15842), .A2(n15173), .ZN(n16727) );
  INV_X1 U20100 ( .A(n16728), .ZN(n20244) );
  OR2_X1 U20101 ( .A1(n20245), .A2(n20246), .ZN(n16728) );
  AND2_X1 U20102 ( .A1(n20247), .A2(n20248), .ZN(n20246) );
  AND2_X1 U20103 ( .A1(n20249), .A2(n20250), .ZN(n20245) );
  OR2_X1 U20104 ( .A1(n20247), .A2(n20248), .ZN(n20250) );
  AND2_X1 U20105 ( .A1(n20251), .A2(n20252), .ZN(n16729) );
  INV_X1 U20106 ( .A(n20253), .ZN(n20252) );
  AND2_X1 U20107 ( .A1(n20254), .A2(n20255), .ZN(n20253) );
  OR2_X1 U20108 ( .A1(n20255), .A2(n20254), .ZN(n20251) );
  OR2_X1 U20109 ( .A1(n20256), .A2(n20257), .ZN(n20254) );
  AND2_X1 U20110 ( .A1(n20258), .A2(n20259), .ZN(n20257) );
  INV_X1 U20111 ( .A(n20260), .ZN(n20258) );
  AND2_X1 U20112 ( .A1(n20261), .A2(n20260), .ZN(n20256) );
  INV_X1 U20113 ( .A(n20259), .ZN(n20261) );
  AND2_X1 U20114 ( .A1(n16744), .A2(n16742), .ZN(n20212) );
  INV_X1 U20115 ( .A(n16753), .ZN(n16742) );
  AND2_X1 U20116 ( .A1(n20262), .A2(n20263), .ZN(n16753) );
  INV_X1 U20117 ( .A(n20264), .ZN(n20263) );
  AND2_X1 U20118 ( .A1(n20265), .A2(n20221), .ZN(n20264) );
  OR2_X1 U20119 ( .A1(n20221), .A2(n20265), .ZN(n20262) );
  OR2_X1 U20120 ( .A1(n20266), .A2(n20267), .ZN(n20265) );
  AND2_X1 U20121 ( .A1(n20268), .A2(n20220), .ZN(n20267) );
  INV_X1 U20122 ( .A(n20219), .ZN(n20268) );
  AND2_X1 U20123 ( .A1(n20269), .A2(n20219), .ZN(n20266) );
  OR2_X1 U20124 ( .A1(n16512), .A2(n15105), .ZN(n20219) );
  INV_X1 U20125 ( .A(n20220), .ZN(n20269) );
  OR2_X1 U20126 ( .A1(n20270), .A2(n20271), .ZN(n20220) );
  AND2_X1 U20127 ( .A1(n20272), .A2(n20273), .ZN(n20271) );
  AND2_X1 U20128 ( .A1(n20274), .A2(n20275), .ZN(n20270) );
  OR2_X1 U20129 ( .A1(n20273), .A2(n20272), .ZN(n20275) );
  AND2_X1 U20130 ( .A1(n20276), .A2(n20277), .ZN(n20221) );
  INV_X1 U20131 ( .A(n20278), .ZN(n20277) );
  AND2_X1 U20132 ( .A1(n20279), .A2(n20235), .ZN(n20278) );
  OR2_X1 U20133 ( .A1(n20235), .A2(n20279), .ZN(n20276) );
  OR2_X1 U20134 ( .A1(n20280), .A2(n20281), .ZN(n20279) );
  AND2_X1 U20135 ( .A1(n20282), .A2(n20234), .ZN(n20281) );
  INV_X1 U20136 ( .A(n20233), .ZN(n20282) );
  AND2_X1 U20137 ( .A1(n20283), .A2(n20233), .ZN(n20280) );
  OR2_X1 U20138 ( .A1(n15842), .A2(n15139), .ZN(n20233) );
  INV_X1 U20139 ( .A(n20234), .ZN(n20283) );
  OR2_X1 U20140 ( .A1(n20284), .A2(n20285), .ZN(n20234) );
  AND2_X1 U20141 ( .A1(n20286), .A2(n20287), .ZN(n20285) );
  AND2_X1 U20142 ( .A1(n20288), .A2(n20289), .ZN(n20284) );
  OR2_X1 U20143 ( .A1(n20286), .A2(n20287), .ZN(n20289) );
  AND2_X1 U20144 ( .A1(n20290), .A2(n20291), .ZN(n20235) );
  INV_X1 U20145 ( .A(n20292), .ZN(n20291) );
  AND2_X1 U20146 ( .A1(n20293), .A2(n20249), .ZN(n20292) );
  OR2_X1 U20147 ( .A1(n20249), .A2(n20293), .ZN(n20290) );
  OR2_X1 U20148 ( .A1(n20294), .A2(n20295), .ZN(n20293) );
  AND2_X1 U20149 ( .A1(n20296), .A2(n20248), .ZN(n20295) );
  INV_X1 U20150 ( .A(n20247), .ZN(n20296) );
  AND2_X1 U20151 ( .A1(n20297), .A2(n20247), .ZN(n20294) );
  OR2_X1 U20152 ( .A1(n15808), .A2(n15173), .ZN(n20247) );
  INV_X1 U20153 ( .A(n20248), .ZN(n20297) );
  OR2_X1 U20154 ( .A1(n20298), .A2(n20299), .ZN(n20248) );
  AND2_X1 U20155 ( .A1(n20300), .A2(n20301), .ZN(n20299) );
  AND2_X1 U20156 ( .A1(n20302), .A2(n20303), .ZN(n20298) );
  OR2_X1 U20157 ( .A1(n20300), .A2(n20301), .ZN(n20303) );
  AND2_X1 U20158 ( .A1(n20304), .A2(n20305), .ZN(n20249) );
  INV_X1 U20159 ( .A(n20306), .ZN(n20305) );
  AND2_X1 U20160 ( .A1(n20307), .A2(n20308), .ZN(n20306) );
  OR2_X1 U20161 ( .A1(n20308), .A2(n20307), .ZN(n20304) );
  OR2_X1 U20162 ( .A1(n20309), .A2(n20310), .ZN(n20307) );
  AND2_X1 U20163 ( .A1(n20311), .A2(n20312), .ZN(n20310) );
  INV_X1 U20164 ( .A(n20313), .ZN(n20311) );
  AND2_X1 U20165 ( .A1(n20314), .A2(n20313), .ZN(n20309) );
  INV_X1 U20166 ( .A(n20312), .ZN(n20314) );
  INV_X1 U20167 ( .A(n16752), .ZN(n16744) );
  OR2_X1 U20168 ( .A1(n20315), .A2(n20316), .ZN(n16752) );
  AND2_X1 U20169 ( .A1(n16778), .A2(n16777), .ZN(n20316) );
  AND2_X1 U20170 ( .A1(n16773), .A2(n20317), .ZN(n20315) );
  OR2_X1 U20171 ( .A1(n16778), .A2(n16777), .ZN(n20317) );
  OR2_X1 U20172 ( .A1(n20318), .A2(n20319), .ZN(n16777) );
  AND2_X1 U20173 ( .A1(n16815), .A2(n16814), .ZN(n20319) );
  AND2_X1 U20174 ( .A1(n16810), .A2(n20320), .ZN(n20318) );
  OR2_X1 U20175 ( .A1(n16815), .A2(n16814), .ZN(n20320) );
  OR2_X1 U20176 ( .A1(n20321), .A2(n20322), .ZN(n16814) );
  AND2_X1 U20177 ( .A1(n16870), .A2(n16869), .ZN(n20322) );
  AND2_X1 U20178 ( .A1(n16865), .A2(n20323), .ZN(n20321) );
  OR2_X1 U20179 ( .A1(n16870), .A2(n16869), .ZN(n20323) );
  OR2_X1 U20180 ( .A1(n20324), .A2(n20325), .ZN(n16869) );
  AND2_X1 U20181 ( .A1(n20210), .A2(n20209), .ZN(n20325) );
  AND2_X1 U20182 ( .A1(n20205), .A2(n20326), .ZN(n20324) );
  OR2_X1 U20183 ( .A1(n20210), .A2(n20209), .ZN(n20326) );
  OR2_X1 U20184 ( .A1(n20327), .A2(n20328), .ZN(n20209) );
  AND2_X1 U20185 ( .A1(n20199), .A2(n20198), .ZN(n20328) );
  AND2_X1 U20186 ( .A1(n20194), .A2(n20329), .ZN(n20327) );
  OR2_X1 U20187 ( .A1(n20199), .A2(n20198), .ZN(n20329) );
  OR2_X1 U20188 ( .A1(n20330), .A2(n20331), .ZN(n20198) );
  AND2_X1 U20189 ( .A1(n20188), .A2(n20187), .ZN(n20331) );
  AND2_X1 U20190 ( .A1(n20183), .A2(n20332), .ZN(n20330) );
  OR2_X1 U20191 ( .A1(n20188), .A2(n20187), .ZN(n20332) );
  OR2_X1 U20192 ( .A1(n20333), .A2(n20334), .ZN(n20187) );
  AND2_X1 U20193 ( .A1(n20178), .A2(n20177), .ZN(n20334) );
  AND2_X1 U20194 ( .A1(n20172), .A2(n20335), .ZN(n20333) );
  OR2_X1 U20195 ( .A1(n20178), .A2(n20177), .ZN(n20335) );
  OR2_X1 U20196 ( .A1(n20336), .A2(n20337), .ZN(n20177) );
  AND2_X1 U20197 ( .A1(n20164), .A2(n20166), .ZN(n20337) );
  AND2_X1 U20198 ( .A1(n20161), .A2(n20338), .ZN(n20336) );
  OR2_X1 U20199 ( .A1(n20164), .A2(n20166), .ZN(n20338) );
  OR2_X1 U20200 ( .A1(n20339), .A2(n20340), .ZN(n20166) );
  AND2_X1 U20201 ( .A1(n20153), .A2(n20155), .ZN(n20340) );
  AND2_X1 U20202 ( .A1(n20150), .A2(n20341), .ZN(n20339) );
  OR2_X1 U20203 ( .A1(n20153), .A2(n20155), .ZN(n20341) );
  OR2_X1 U20204 ( .A1(n20342), .A2(n20343), .ZN(n20155) );
  AND2_X1 U20205 ( .A1(n20142), .A2(n20144), .ZN(n20343) );
  AND2_X1 U20206 ( .A1(n20139), .A2(n20344), .ZN(n20342) );
  OR2_X1 U20207 ( .A1(n20142), .A2(n20144), .ZN(n20344) );
  OR2_X1 U20208 ( .A1(n20345), .A2(n20346), .ZN(n20144) );
  AND2_X1 U20209 ( .A1(n20131), .A2(n20133), .ZN(n20346) );
  AND2_X1 U20210 ( .A1(n20128), .A2(n20347), .ZN(n20345) );
  OR2_X1 U20211 ( .A1(n20131), .A2(n20133), .ZN(n20347) );
  OR2_X1 U20212 ( .A1(n20348), .A2(n20349), .ZN(n20133) );
  AND2_X1 U20213 ( .A1(n20120), .A2(n20122), .ZN(n20349) );
  AND2_X1 U20214 ( .A1(n20117), .A2(n20350), .ZN(n20348) );
  OR2_X1 U20215 ( .A1(n20120), .A2(n20122), .ZN(n20350) );
  OR2_X1 U20216 ( .A1(n20351), .A2(n20352), .ZN(n20122) );
  AND2_X1 U20217 ( .A1(n20109), .A2(n20111), .ZN(n20352) );
  AND2_X1 U20218 ( .A1(n20106), .A2(n20353), .ZN(n20351) );
  OR2_X1 U20219 ( .A1(n20109), .A2(n20111), .ZN(n20353) );
  OR2_X1 U20220 ( .A1(n20354), .A2(n20355), .ZN(n20111) );
  AND2_X1 U20221 ( .A1(n20098), .A2(n20100), .ZN(n20355) );
  AND2_X1 U20222 ( .A1(n20095), .A2(n20356), .ZN(n20354) );
  OR2_X1 U20223 ( .A1(n20098), .A2(n20100), .ZN(n20356) );
  OR2_X1 U20224 ( .A1(n20357), .A2(n20358), .ZN(n20100) );
  AND2_X1 U20225 ( .A1(n20087), .A2(n20089), .ZN(n20358) );
  AND2_X1 U20226 ( .A1(n20084), .A2(n20359), .ZN(n20357) );
  OR2_X1 U20227 ( .A1(n20087), .A2(n20089), .ZN(n20359) );
  OR2_X1 U20228 ( .A1(n20360), .A2(n20361), .ZN(n20089) );
  AND2_X1 U20229 ( .A1(n20076), .A2(n20078), .ZN(n20361) );
  AND2_X1 U20230 ( .A1(n20073), .A2(n20362), .ZN(n20360) );
  OR2_X1 U20231 ( .A1(n20076), .A2(n20078), .ZN(n20362) );
  OR2_X1 U20232 ( .A1(n20363), .A2(n20364), .ZN(n20078) );
  AND2_X1 U20233 ( .A1(n20065), .A2(n20067), .ZN(n20364) );
  AND2_X1 U20234 ( .A1(n20062), .A2(n20365), .ZN(n20363) );
  OR2_X1 U20235 ( .A1(n20065), .A2(n20067), .ZN(n20365) );
  OR2_X1 U20236 ( .A1(n20366), .A2(n20367), .ZN(n20067) );
  AND2_X1 U20237 ( .A1(n20054), .A2(n20056), .ZN(n20367) );
  AND2_X1 U20238 ( .A1(n20051), .A2(n20368), .ZN(n20366) );
  OR2_X1 U20239 ( .A1(n20054), .A2(n20056), .ZN(n20368) );
  OR2_X1 U20240 ( .A1(n20369), .A2(n20370), .ZN(n20056) );
  AND2_X1 U20241 ( .A1(n20043), .A2(n20045), .ZN(n20370) );
  AND2_X1 U20242 ( .A1(n20040), .A2(n20371), .ZN(n20369) );
  OR2_X1 U20243 ( .A1(n20043), .A2(n20045), .ZN(n20371) );
  OR2_X1 U20244 ( .A1(n20372), .A2(n20373), .ZN(n20045) );
  AND2_X1 U20245 ( .A1(n20032), .A2(n20034), .ZN(n20373) );
  AND2_X1 U20246 ( .A1(n20029), .A2(n20374), .ZN(n20372) );
  OR2_X1 U20247 ( .A1(n20032), .A2(n20034), .ZN(n20374) );
  OR2_X1 U20248 ( .A1(n20375), .A2(n20376), .ZN(n20034) );
  AND2_X1 U20249 ( .A1(n20021), .A2(n20023), .ZN(n20376) );
  AND2_X1 U20250 ( .A1(n20018), .A2(n20377), .ZN(n20375) );
  OR2_X1 U20251 ( .A1(n20021), .A2(n20023), .ZN(n20377) );
  OR2_X1 U20252 ( .A1(n20378), .A2(n20379), .ZN(n20023) );
  AND2_X1 U20253 ( .A1(n20010), .A2(n20012), .ZN(n20379) );
  AND2_X1 U20254 ( .A1(n20007), .A2(n20380), .ZN(n20378) );
  OR2_X1 U20255 ( .A1(n20010), .A2(n20012), .ZN(n20380) );
  OR2_X1 U20256 ( .A1(n20381), .A2(n20382), .ZN(n20012) );
  AND2_X1 U20257 ( .A1(n19999), .A2(n20001), .ZN(n20382) );
  AND2_X1 U20258 ( .A1(n19996), .A2(n20383), .ZN(n20381) );
  OR2_X1 U20259 ( .A1(n19999), .A2(n20001), .ZN(n20383) );
  OR2_X1 U20260 ( .A1(n20384), .A2(n20385), .ZN(n20001) );
  AND2_X1 U20261 ( .A1(n15936), .A2(n19990), .ZN(n20385) );
  AND2_X1 U20262 ( .A1(n19986), .A2(n20386), .ZN(n20384) );
  OR2_X1 U20263 ( .A1(n15936), .A2(n19990), .ZN(n20386) );
  OR2_X1 U20264 ( .A1(n20387), .A2(n20388), .ZN(n19990) );
  AND2_X1 U20265 ( .A1(n19978), .A2(n19980), .ZN(n20388) );
  AND2_X1 U20266 ( .A1(n19975), .A2(n20389), .ZN(n20387) );
  OR2_X1 U20267 ( .A1(n19978), .A2(n19980), .ZN(n20389) );
  OR2_X1 U20268 ( .A1(n20390), .A2(n20391), .ZN(n19980) );
  AND2_X1 U20269 ( .A1(n19967), .A2(n19969), .ZN(n20391) );
  AND2_X1 U20270 ( .A1(n19964), .A2(n20392), .ZN(n20390) );
  OR2_X1 U20271 ( .A1(n19967), .A2(n19969), .ZN(n20392) );
  OR2_X1 U20272 ( .A1(n20393), .A2(n20394), .ZN(n19969) );
  AND2_X1 U20273 ( .A1(n19956), .A2(n19958), .ZN(n20394) );
  AND2_X1 U20274 ( .A1(n19953), .A2(n20395), .ZN(n20393) );
  OR2_X1 U20275 ( .A1(n19956), .A2(n19958), .ZN(n20395) );
  OR2_X1 U20276 ( .A1(n20396), .A2(n20397), .ZN(n19958) );
  AND2_X1 U20277 ( .A1(n19945), .A2(n19947), .ZN(n20397) );
  AND2_X1 U20278 ( .A1(n19942), .A2(n20398), .ZN(n20396) );
  OR2_X1 U20279 ( .A1(n19945), .A2(n19947), .ZN(n20398) );
  OR2_X1 U20280 ( .A1(n20399), .A2(n20400), .ZN(n19947) );
  AND2_X1 U20281 ( .A1(n19934), .A2(n19936), .ZN(n20400) );
  AND2_X1 U20282 ( .A1(n19931), .A2(n20401), .ZN(n20399) );
  OR2_X1 U20283 ( .A1(n19934), .A2(n19936), .ZN(n20401) );
  OR2_X1 U20284 ( .A1(n20402), .A2(n20403), .ZN(n19936) );
  AND2_X1 U20285 ( .A1(n19919), .A2(n19924), .ZN(n20403) );
  AND2_X1 U20286 ( .A1(n19923), .A2(n20404), .ZN(n20402) );
  OR2_X1 U20287 ( .A1(n19919), .A2(n19924), .ZN(n20404) );
  INV_X1 U20288 ( .A(n19925), .ZN(n19924) );
  AND3_X1 U20289 ( .A1(b_23_), .A2(b_22_), .A3(n15957), .ZN(n19925) );
  OR2_X1 U20290 ( .A1(n14857), .A2(n15071), .ZN(n19919) );
  INV_X1 U20291 ( .A(n19926), .ZN(n19923) );
  OR2_X1 U20292 ( .A1(n20405), .A2(n20406), .ZN(n19926) );
  AND2_X1 U20293 ( .A1(b_22_), .A2(n20407), .ZN(n20406) );
  OR2_X1 U20294 ( .A1(n20408), .A2(n16981), .ZN(n20407) );
  AND2_X1 U20295 ( .A1(a_30_), .A2(n15139), .ZN(n20408) );
  AND2_X1 U20296 ( .A1(b_21_), .A2(n20409), .ZN(n20405) );
  OR2_X1 U20297 ( .A1(n20410), .A2(n14817), .ZN(n20409) );
  AND2_X1 U20298 ( .A1(a_31_), .A2(n15105), .ZN(n20410) );
  OR2_X1 U20299 ( .A1(n14891), .A2(n15071), .ZN(n19934) );
  OR2_X1 U20300 ( .A1(n20411), .A2(n20412), .ZN(n19931) );
  AND2_X1 U20301 ( .A1(n20413), .A2(n20414), .ZN(n20412) );
  INV_X1 U20302 ( .A(n20415), .ZN(n20411) );
  OR2_X1 U20303 ( .A1(n20413), .A2(n20414), .ZN(n20415) );
  OR2_X1 U20304 ( .A1(n20416), .A2(n20417), .ZN(n20413) );
  AND2_X1 U20305 ( .A1(n20418), .A2(n20419), .ZN(n20417) );
  AND2_X1 U20306 ( .A1(n20420), .A2(n20421), .ZN(n20416) );
  OR2_X1 U20307 ( .A1(n14936), .A2(n15071), .ZN(n19945) );
  OR2_X1 U20308 ( .A1(n20422), .A2(n20423), .ZN(n19942) );
  INV_X1 U20309 ( .A(n20424), .ZN(n20423) );
  OR2_X1 U20310 ( .A1(n20425), .A2(n20426), .ZN(n20424) );
  AND2_X1 U20311 ( .A1(n20426), .A2(n20425), .ZN(n20422) );
  AND2_X1 U20312 ( .A1(n20427), .A2(n20428), .ZN(n20425) );
  OR2_X1 U20313 ( .A1(n20429), .A2(n20430), .ZN(n20428) );
  INV_X1 U20314 ( .A(n20431), .ZN(n20430) );
  OR2_X1 U20315 ( .A1(n20431), .A2(n20432), .ZN(n20427) );
  INV_X1 U20316 ( .A(n20429), .ZN(n20432) );
  OR2_X1 U20317 ( .A1(n14970), .A2(n15071), .ZN(n19956) );
  OR2_X1 U20318 ( .A1(n20433), .A2(n20434), .ZN(n19953) );
  INV_X1 U20319 ( .A(n20435), .ZN(n20434) );
  OR2_X1 U20320 ( .A1(n20436), .A2(n20437), .ZN(n20435) );
  AND2_X1 U20321 ( .A1(n20437), .A2(n20436), .ZN(n20433) );
  AND2_X1 U20322 ( .A1(n20438), .A2(n20439), .ZN(n20436) );
  OR2_X1 U20323 ( .A1(n20440), .A2(n20441), .ZN(n20439) );
  INV_X1 U20324 ( .A(n20442), .ZN(n20441) );
  OR2_X1 U20325 ( .A1(n20442), .A2(n20443), .ZN(n20438) );
  INV_X1 U20326 ( .A(n20440), .ZN(n20443) );
  OR2_X1 U20327 ( .A1(n15004), .A2(n15071), .ZN(n19967) );
  OR2_X1 U20328 ( .A1(n20444), .A2(n20445), .ZN(n19964) );
  INV_X1 U20329 ( .A(n20446), .ZN(n20445) );
  OR2_X1 U20330 ( .A1(n20447), .A2(n20448), .ZN(n20446) );
  AND2_X1 U20331 ( .A1(n20448), .A2(n20447), .ZN(n20444) );
  AND2_X1 U20332 ( .A1(n20449), .A2(n20450), .ZN(n20447) );
  OR2_X1 U20333 ( .A1(n20451), .A2(n20452), .ZN(n20450) );
  INV_X1 U20334 ( .A(n20453), .ZN(n20452) );
  OR2_X1 U20335 ( .A1(n20453), .A2(n20454), .ZN(n20449) );
  INV_X1 U20336 ( .A(n20451), .ZN(n20454) );
  OR2_X1 U20337 ( .A1(n15038), .A2(n15071), .ZN(n19978) );
  OR2_X1 U20338 ( .A1(n20455), .A2(n20456), .ZN(n19975) );
  INV_X1 U20339 ( .A(n20457), .ZN(n20456) );
  OR2_X1 U20340 ( .A1(n20458), .A2(n20459), .ZN(n20457) );
  AND2_X1 U20341 ( .A1(n20459), .A2(n20458), .ZN(n20455) );
  AND2_X1 U20342 ( .A1(n20460), .A2(n20461), .ZN(n20458) );
  OR2_X1 U20343 ( .A1(n20462), .A2(n20463), .ZN(n20461) );
  INV_X1 U20344 ( .A(n20464), .ZN(n20463) );
  OR2_X1 U20345 ( .A1(n20464), .A2(n20465), .ZN(n20460) );
  INV_X1 U20346 ( .A(n20462), .ZN(n20465) );
  OR2_X1 U20347 ( .A1(n15072), .A2(n15071), .ZN(n15936) );
  OR2_X1 U20348 ( .A1(n20466), .A2(n20467), .ZN(n19986) );
  INV_X1 U20349 ( .A(n20468), .ZN(n20467) );
  OR2_X1 U20350 ( .A1(n20469), .A2(n20470), .ZN(n20468) );
  AND2_X1 U20351 ( .A1(n20470), .A2(n20469), .ZN(n20466) );
  AND2_X1 U20352 ( .A1(n20471), .A2(n20472), .ZN(n20469) );
  OR2_X1 U20353 ( .A1(n20473), .A2(n20474), .ZN(n20472) );
  INV_X1 U20354 ( .A(n20475), .ZN(n20474) );
  OR2_X1 U20355 ( .A1(n20475), .A2(n20476), .ZN(n20471) );
  INV_X1 U20356 ( .A(n20473), .ZN(n20476) );
  OR2_X1 U20357 ( .A1(n15106), .A2(n15071), .ZN(n19999) );
  OR2_X1 U20358 ( .A1(n20477), .A2(n20478), .ZN(n19996) );
  INV_X1 U20359 ( .A(n20479), .ZN(n20478) );
  OR2_X1 U20360 ( .A1(n20480), .A2(n20481), .ZN(n20479) );
  AND2_X1 U20361 ( .A1(n20481), .A2(n20480), .ZN(n20477) );
  AND2_X1 U20362 ( .A1(n20482), .A2(n20483), .ZN(n20480) );
  OR2_X1 U20363 ( .A1(n20484), .A2(n20485), .ZN(n20483) );
  INV_X1 U20364 ( .A(n20486), .ZN(n20485) );
  OR2_X1 U20365 ( .A1(n20486), .A2(n20487), .ZN(n20482) );
  INV_X1 U20366 ( .A(n20484), .ZN(n20487) );
  OR2_X1 U20367 ( .A1(n15140), .A2(n15071), .ZN(n20010) );
  OR2_X1 U20368 ( .A1(n20488), .A2(n20489), .ZN(n20007) );
  INV_X1 U20369 ( .A(n20490), .ZN(n20489) );
  OR2_X1 U20370 ( .A1(n20491), .A2(n20492), .ZN(n20490) );
  AND2_X1 U20371 ( .A1(n20492), .A2(n20491), .ZN(n20488) );
  AND2_X1 U20372 ( .A1(n20493), .A2(n20494), .ZN(n20491) );
  OR2_X1 U20373 ( .A1(n15933), .A2(n20495), .ZN(n20494) );
  INV_X1 U20374 ( .A(n20496), .ZN(n20495) );
  OR2_X1 U20375 ( .A1(n20496), .A2(n20497), .ZN(n20493) );
  INV_X1 U20376 ( .A(n15933), .ZN(n20497) );
  OR2_X1 U20377 ( .A1(n15174), .A2(n15071), .ZN(n20021) );
  OR2_X1 U20378 ( .A1(n20498), .A2(n20499), .ZN(n20018) );
  INV_X1 U20379 ( .A(n20500), .ZN(n20499) );
  OR2_X1 U20380 ( .A1(n20501), .A2(n20502), .ZN(n20500) );
  AND2_X1 U20381 ( .A1(n20502), .A2(n20501), .ZN(n20498) );
  AND2_X1 U20382 ( .A1(n20503), .A2(n20504), .ZN(n20501) );
  OR2_X1 U20383 ( .A1(n20505), .A2(n20506), .ZN(n20504) );
  INV_X1 U20384 ( .A(n20507), .ZN(n20506) );
  OR2_X1 U20385 ( .A1(n20507), .A2(n20508), .ZN(n20503) );
  INV_X1 U20386 ( .A(n20505), .ZN(n20508) );
  OR2_X1 U20387 ( .A1(n15208), .A2(n15071), .ZN(n20032) );
  OR2_X1 U20388 ( .A1(n20509), .A2(n20510), .ZN(n20029) );
  INV_X1 U20389 ( .A(n20511), .ZN(n20510) );
  OR2_X1 U20390 ( .A1(n20512), .A2(n20513), .ZN(n20511) );
  AND2_X1 U20391 ( .A1(n20513), .A2(n20512), .ZN(n20509) );
  AND2_X1 U20392 ( .A1(n20514), .A2(n20515), .ZN(n20512) );
  OR2_X1 U20393 ( .A1(n20516), .A2(n20517), .ZN(n20515) );
  INV_X1 U20394 ( .A(n20518), .ZN(n20517) );
  OR2_X1 U20395 ( .A1(n20518), .A2(n20519), .ZN(n20514) );
  INV_X1 U20396 ( .A(n20516), .ZN(n20519) );
  OR2_X1 U20397 ( .A1(n15242), .A2(n15071), .ZN(n20043) );
  OR2_X1 U20398 ( .A1(n20520), .A2(n20521), .ZN(n20040) );
  INV_X1 U20399 ( .A(n20522), .ZN(n20521) );
  OR2_X1 U20400 ( .A1(n20523), .A2(n20524), .ZN(n20522) );
  AND2_X1 U20401 ( .A1(n20524), .A2(n20523), .ZN(n20520) );
  AND2_X1 U20402 ( .A1(n20525), .A2(n20526), .ZN(n20523) );
  OR2_X1 U20403 ( .A1(n20527), .A2(n20528), .ZN(n20526) );
  INV_X1 U20404 ( .A(n20529), .ZN(n20528) );
  OR2_X1 U20405 ( .A1(n20529), .A2(n20530), .ZN(n20525) );
  INV_X1 U20406 ( .A(n20527), .ZN(n20530) );
  OR2_X1 U20407 ( .A1(n15287), .A2(n15071), .ZN(n20054) );
  OR2_X1 U20408 ( .A1(n20531), .A2(n20532), .ZN(n20051) );
  INV_X1 U20409 ( .A(n20533), .ZN(n20532) );
  OR2_X1 U20410 ( .A1(n20534), .A2(n20535), .ZN(n20533) );
  AND2_X1 U20411 ( .A1(n20535), .A2(n20534), .ZN(n20531) );
  AND2_X1 U20412 ( .A1(n20536), .A2(n20537), .ZN(n20534) );
  OR2_X1 U20413 ( .A1(n20538), .A2(n20539), .ZN(n20537) );
  INV_X1 U20414 ( .A(n20540), .ZN(n20539) );
  OR2_X1 U20415 ( .A1(n20540), .A2(n20541), .ZN(n20536) );
  INV_X1 U20416 ( .A(n20538), .ZN(n20541) );
  OR2_X1 U20417 ( .A1(n15321), .A2(n15071), .ZN(n20065) );
  OR2_X1 U20418 ( .A1(n20542), .A2(n20543), .ZN(n20062) );
  INV_X1 U20419 ( .A(n20544), .ZN(n20543) );
  OR2_X1 U20420 ( .A1(n20545), .A2(n20546), .ZN(n20544) );
  AND2_X1 U20421 ( .A1(n20546), .A2(n20545), .ZN(n20542) );
  AND2_X1 U20422 ( .A1(n20547), .A2(n20548), .ZN(n20545) );
  OR2_X1 U20423 ( .A1(n20549), .A2(n20550), .ZN(n20548) );
  INV_X1 U20424 ( .A(n20551), .ZN(n20550) );
  OR2_X1 U20425 ( .A1(n20551), .A2(n20552), .ZN(n20547) );
  INV_X1 U20426 ( .A(n20549), .ZN(n20552) );
  OR2_X1 U20427 ( .A1(n15355), .A2(n15071), .ZN(n20076) );
  OR2_X1 U20428 ( .A1(n20553), .A2(n20554), .ZN(n20073) );
  INV_X1 U20429 ( .A(n20555), .ZN(n20554) );
  OR2_X1 U20430 ( .A1(n20556), .A2(n20557), .ZN(n20555) );
  AND2_X1 U20431 ( .A1(n20557), .A2(n20556), .ZN(n20553) );
  AND2_X1 U20432 ( .A1(n20558), .A2(n20559), .ZN(n20556) );
  OR2_X1 U20433 ( .A1(n20560), .A2(n20561), .ZN(n20559) );
  INV_X1 U20434 ( .A(n20562), .ZN(n20561) );
  OR2_X1 U20435 ( .A1(n20562), .A2(n20563), .ZN(n20558) );
  INV_X1 U20436 ( .A(n20560), .ZN(n20563) );
  OR2_X1 U20437 ( .A1(n15389), .A2(n15071), .ZN(n20087) );
  OR2_X1 U20438 ( .A1(n20564), .A2(n20565), .ZN(n20084) );
  INV_X1 U20439 ( .A(n20566), .ZN(n20565) );
  OR2_X1 U20440 ( .A1(n20567), .A2(n20568), .ZN(n20566) );
  AND2_X1 U20441 ( .A1(n20568), .A2(n20567), .ZN(n20564) );
  AND2_X1 U20442 ( .A1(n20569), .A2(n20570), .ZN(n20567) );
  OR2_X1 U20443 ( .A1(n20571), .A2(n20572), .ZN(n20570) );
  INV_X1 U20444 ( .A(n20573), .ZN(n20572) );
  OR2_X1 U20445 ( .A1(n20573), .A2(n20574), .ZN(n20569) );
  INV_X1 U20446 ( .A(n20571), .ZN(n20574) );
  OR2_X1 U20447 ( .A1(n15423), .A2(n15071), .ZN(n20098) );
  OR2_X1 U20448 ( .A1(n20575), .A2(n20576), .ZN(n20095) );
  INV_X1 U20449 ( .A(n20577), .ZN(n20576) );
  OR2_X1 U20450 ( .A1(n20578), .A2(n20579), .ZN(n20577) );
  AND2_X1 U20451 ( .A1(n20579), .A2(n20578), .ZN(n20575) );
  AND2_X1 U20452 ( .A1(n20580), .A2(n20581), .ZN(n20578) );
  OR2_X1 U20453 ( .A1(n20582), .A2(n20583), .ZN(n20581) );
  INV_X1 U20454 ( .A(n20584), .ZN(n20583) );
  OR2_X1 U20455 ( .A1(n20584), .A2(n20585), .ZN(n20580) );
  INV_X1 U20456 ( .A(n20582), .ZN(n20585) );
  OR2_X1 U20457 ( .A1(n15457), .A2(n15071), .ZN(n20109) );
  OR2_X1 U20458 ( .A1(n20586), .A2(n20587), .ZN(n20106) );
  INV_X1 U20459 ( .A(n20588), .ZN(n20587) );
  OR2_X1 U20460 ( .A1(n20589), .A2(n20590), .ZN(n20588) );
  AND2_X1 U20461 ( .A1(n20590), .A2(n20589), .ZN(n20586) );
  AND2_X1 U20462 ( .A1(n20591), .A2(n20592), .ZN(n20589) );
  OR2_X1 U20463 ( .A1(n20593), .A2(n20594), .ZN(n20592) );
  INV_X1 U20464 ( .A(n20595), .ZN(n20594) );
  OR2_X1 U20465 ( .A1(n20595), .A2(n20596), .ZN(n20591) );
  INV_X1 U20466 ( .A(n20593), .ZN(n20596) );
  OR2_X1 U20467 ( .A1(n15491), .A2(n15071), .ZN(n20120) );
  OR2_X1 U20468 ( .A1(n20597), .A2(n20598), .ZN(n20117) );
  INV_X1 U20469 ( .A(n20599), .ZN(n20598) );
  OR2_X1 U20470 ( .A1(n20600), .A2(n20601), .ZN(n20599) );
  AND2_X1 U20471 ( .A1(n20601), .A2(n20600), .ZN(n20597) );
  AND2_X1 U20472 ( .A1(n20602), .A2(n20603), .ZN(n20600) );
  OR2_X1 U20473 ( .A1(n20604), .A2(n20605), .ZN(n20603) );
  INV_X1 U20474 ( .A(n20606), .ZN(n20605) );
  OR2_X1 U20475 ( .A1(n20606), .A2(n20607), .ZN(n20602) );
  INV_X1 U20476 ( .A(n20604), .ZN(n20607) );
  OR2_X1 U20477 ( .A1(n15525), .A2(n15071), .ZN(n20131) );
  OR2_X1 U20478 ( .A1(n20608), .A2(n20609), .ZN(n20128) );
  INV_X1 U20479 ( .A(n20610), .ZN(n20609) );
  OR2_X1 U20480 ( .A1(n20611), .A2(n20612), .ZN(n20610) );
  AND2_X1 U20481 ( .A1(n20612), .A2(n20611), .ZN(n20608) );
  AND2_X1 U20482 ( .A1(n20613), .A2(n20614), .ZN(n20611) );
  OR2_X1 U20483 ( .A1(n20615), .A2(n20616), .ZN(n20614) );
  INV_X1 U20484 ( .A(n20617), .ZN(n20616) );
  OR2_X1 U20485 ( .A1(n20617), .A2(n20618), .ZN(n20613) );
  INV_X1 U20486 ( .A(n20615), .ZN(n20618) );
  OR2_X1 U20487 ( .A1(n15559), .A2(n15071), .ZN(n20142) );
  OR2_X1 U20488 ( .A1(n20619), .A2(n20620), .ZN(n20139) );
  INV_X1 U20489 ( .A(n20621), .ZN(n20620) );
  OR2_X1 U20490 ( .A1(n20622), .A2(n20623), .ZN(n20621) );
  AND2_X1 U20491 ( .A1(n20623), .A2(n20622), .ZN(n20619) );
  AND2_X1 U20492 ( .A1(n20624), .A2(n20625), .ZN(n20622) );
  OR2_X1 U20493 ( .A1(n20626), .A2(n20627), .ZN(n20625) );
  INV_X1 U20494 ( .A(n20628), .ZN(n20627) );
  OR2_X1 U20495 ( .A1(n20628), .A2(n20629), .ZN(n20624) );
  INV_X1 U20496 ( .A(n20626), .ZN(n20629) );
  OR2_X1 U20497 ( .A1(n15593), .A2(n15071), .ZN(n20153) );
  OR2_X1 U20498 ( .A1(n20630), .A2(n20631), .ZN(n20150) );
  INV_X1 U20499 ( .A(n20632), .ZN(n20631) );
  OR2_X1 U20500 ( .A1(n20633), .A2(n20634), .ZN(n20632) );
  AND2_X1 U20501 ( .A1(n20634), .A2(n20633), .ZN(n20630) );
  AND2_X1 U20502 ( .A1(n20635), .A2(n20636), .ZN(n20633) );
  OR2_X1 U20503 ( .A1(n20637), .A2(n20638), .ZN(n20636) );
  INV_X1 U20504 ( .A(n20639), .ZN(n20638) );
  OR2_X1 U20505 ( .A1(n20639), .A2(n20640), .ZN(n20635) );
  INV_X1 U20506 ( .A(n20637), .ZN(n20640) );
  OR2_X1 U20507 ( .A1(n15638), .A2(n15071), .ZN(n20164) );
  OR2_X1 U20508 ( .A1(n20641), .A2(n20642), .ZN(n20161) );
  INV_X1 U20509 ( .A(n20643), .ZN(n20642) );
  OR2_X1 U20510 ( .A1(n20644), .A2(n20645), .ZN(n20643) );
  AND2_X1 U20511 ( .A1(n20645), .A2(n20644), .ZN(n20641) );
  AND2_X1 U20512 ( .A1(n20646), .A2(n20647), .ZN(n20644) );
  OR2_X1 U20513 ( .A1(n20648), .A2(n20649), .ZN(n20647) );
  INV_X1 U20514 ( .A(n20650), .ZN(n20649) );
  OR2_X1 U20515 ( .A1(n20650), .A2(n20651), .ZN(n20646) );
  INV_X1 U20516 ( .A(n20648), .ZN(n20651) );
  OR2_X1 U20517 ( .A1(n15672), .A2(n15071), .ZN(n20178) );
  OR2_X1 U20518 ( .A1(n20652), .A2(n20653), .ZN(n20172) );
  INV_X1 U20519 ( .A(n20654), .ZN(n20653) );
  OR2_X1 U20520 ( .A1(n20655), .A2(n20656), .ZN(n20654) );
  AND2_X1 U20521 ( .A1(n20656), .A2(n20655), .ZN(n20652) );
  AND2_X1 U20522 ( .A1(n20657), .A2(n20658), .ZN(n20655) );
  INV_X1 U20523 ( .A(n20659), .ZN(n20658) );
  AND2_X1 U20524 ( .A1(n20660), .A2(n20661), .ZN(n20659) );
  OR2_X1 U20525 ( .A1(n20661), .A2(n20660), .ZN(n20657) );
  INV_X1 U20526 ( .A(n20662), .ZN(n20660) );
  OR2_X1 U20527 ( .A1(n15706), .A2(n15071), .ZN(n20188) );
  AND2_X1 U20528 ( .A1(n20663), .A2(n20664), .ZN(n20183) );
  INV_X1 U20529 ( .A(n20665), .ZN(n20664) );
  AND2_X1 U20530 ( .A1(n20666), .A2(n20667), .ZN(n20665) );
  OR2_X1 U20531 ( .A1(n20667), .A2(n20666), .ZN(n20663) );
  OR2_X1 U20532 ( .A1(n20668), .A2(n20669), .ZN(n20666) );
  AND2_X1 U20533 ( .A1(n20670), .A2(n20671), .ZN(n20669) );
  INV_X1 U20534 ( .A(n20672), .ZN(n20670) );
  AND2_X1 U20535 ( .A1(n20673), .A2(n20672), .ZN(n20668) );
  INV_X1 U20536 ( .A(n20671), .ZN(n20673) );
  OR2_X1 U20537 ( .A1(n15740), .A2(n15071), .ZN(n20199) );
  AND2_X1 U20538 ( .A1(n20674), .A2(n20675), .ZN(n20194) );
  INV_X1 U20539 ( .A(n20676), .ZN(n20675) );
  AND2_X1 U20540 ( .A1(n20677), .A2(n20678), .ZN(n20676) );
  OR2_X1 U20541 ( .A1(n20678), .A2(n20677), .ZN(n20674) );
  OR2_X1 U20542 ( .A1(n20679), .A2(n20680), .ZN(n20677) );
  AND2_X1 U20543 ( .A1(n20681), .A2(n20682), .ZN(n20680) );
  INV_X1 U20544 ( .A(n20683), .ZN(n20681) );
  AND2_X1 U20545 ( .A1(n20684), .A2(n20683), .ZN(n20679) );
  INV_X1 U20546 ( .A(n20682), .ZN(n20684) );
  OR2_X1 U20547 ( .A1(n15774), .A2(n15071), .ZN(n20210) );
  AND2_X1 U20548 ( .A1(n20685), .A2(n20686), .ZN(n20205) );
  INV_X1 U20549 ( .A(n20687), .ZN(n20686) );
  AND2_X1 U20550 ( .A1(n20688), .A2(n20689), .ZN(n20687) );
  OR2_X1 U20551 ( .A1(n20689), .A2(n20688), .ZN(n20685) );
  OR2_X1 U20552 ( .A1(n20690), .A2(n20691), .ZN(n20688) );
  AND2_X1 U20553 ( .A1(n20692), .A2(n20693), .ZN(n20691) );
  INV_X1 U20554 ( .A(n20694), .ZN(n20692) );
  AND2_X1 U20555 ( .A1(n20695), .A2(n20694), .ZN(n20690) );
  INV_X1 U20556 ( .A(n20693), .ZN(n20695) );
  OR2_X1 U20557 ( .A1(n15808), .A2(n15071), .ZN(n16870) );
  AND2_X1 U20558 ( .A1(n20696), .A2(n20697), .ZN(n16865) );
  INV_X1 U20559 ( .A(n20698), .ZN(n20697) );
  AND2_X1 U20560 ( .A1(n20699), .A2(n20700), .ZN(n20698) );
  OR2_X1 U20561 ( .A1(n20700), .A2(n20699), .ZN(n20696) );
  OR2_X1 U20562 ( .A1(n20701), .A2(n20702), .ZN(n20699) );
  AND2_X1 U20563 ( .A1(n20703), .A2(n20704), .ZN(n20702) );
  INV_X1 U20564 ( .A(n20705), .ZN(n20703) );
  AND2_X1 U20565 ( .A1(n20706), .A2(n20705), .ZN(n20701) );
  INV_X1 U20566 ( .A(n20704), .ZN(n20706) );
  OR2_X1 U20567 ( .A1(n15842), .A2(n15071), .ZN(n16815) );
  AND2_X1 U20568 ( .A1(n20707), .A2(n20708), .ZN(n16810) );
  INV_X1 U20569 ( .A(n20709), .ZN(n20708) );
  AND2_X1 U20570 ( .A1(n20710), .A2(n20711), .ZN(n20709) );
  OR2_X1 U20571 ( .A1(n20711), .A2(n20710), .ZN(n20707) );
  OR2_X1 U20572 ( .A1(n20712), .A2(n20713), .ZN(n20710) );
  AND2_X1 U20573 ( .A1(n20714), .A2(n20715), .ZN(n20713) );
  INV_X1 U20574 ( .A(n20716), .ZN(n20714) );
  AND2_X1 U20575 ( .A1(n20717), .A2(n20716), .ZN(n20712) );
  INV_X1 U20576 ( .A(n20715), .ZN(n20717) );
  OR2_X1 U20577 ( .A1(n16512), .A2(n15071), .ZN(n16778) );
  INV_X1 U20578 ( .A(b_23_), .ZN(n15071) );
  AND2_X1 U20579 ( .A1(n20718), .A2(n20719), .ZN(n16773) );
  INV_X1 U20580 ( .A(n20720), .ZN(n20719) );
  AND2_X1 U20581 ( .A1(n20721), .A2(n20274), .ZN(n20720) );
  OR2_X1 U20582 ( .A1(n20274), .A2(n20721), .ZN(n20718) );
  OR2_X1 U20583 ( .A1(n20722), .A2(n20723), .ZN(n20721) );
  AND2_X1 U20584 ( .A1(n20724), .A2(n20273), .ZN(n20723) );
  INV_X1 U20585 ( .A(n20272), .ZN(n20724) );
  AND2_X1 U20586 ( .A1(n20725), .A2(n20272), .ZN(n20722) );
  OR2_X1 U20587 ( .A1(n15842), .A2(n15105), .ZN(n20272) );
  INV_X1 U20588 ( .A(n20273), .ZN(n20725) );
  OR2_X1 U20589 ( .A1(n20726), .A2(n20727), .ZN(n20273) );
  AND2_X1 U20590 ( .A1(n20716), .A2(n20715), .ZN(n20727) );
  AND2_X1 U20591 ( .A1(n20711), .A2(n20728), .ZN(n20726) );
  OR2_X1 U20592 ( .A1(n20715), .A2(n20716), .ZN(n20728) );
  OR2_X1 U20593 ( .A1(n15808), .A2(n15105), .ZN(n20716) );
  OR2_X1 U20594 ( .A1(n20729), .A2(n20730), .ZN(n20715) );
  AND2_X1 U20595 ( .A1(n20705), .A2(n20704), .ZN(n20730) );
  AND2_X1 U20596 ( .A1(n20700), .A2(n20731), .ZN(n20729) );
  OR2_X1 U20597 ( .A1(n20704), .A2(n20705), .ZN(n20731) );
  OR2_X1 U20598 ( .A1(n15774), .A2(n15105), .ZN(n20705) );
  OR2_X1 U20599 ( .A1(n20732), .A2(n20733), .ZN(n20704) );
  AND2_X1 U20600 ( .A1(n20694), .A2(n20693), .ZN(n20733) );
  AND2_X1 U20601 ( .A1(n20689), .A2(n20734), .ZN(n20732) );
  OR2_X1 U20602 ( .A1(n20693), .A2(n20694), .ZN(n20734) );
  OR2_X1 U20603 ( .A1(n15740), .A2(n15105), .ZN(n20694) );
  OR2_X1 U20604 ( .A1(n20735), .A2(n20736), .ZN(n20693) );
  AND2_X1 U20605 ( .A1(n20683), .A2(n20682), .ZN(n20736) );
  AND2_X1 U20606 ( .A1(n20678), .A2(n20737), .ZN(n20735) );
  OR2_X1 U20607 ( .A1(n20682), .A2(n20683), .ZN(n20737) );
  OR2_X1 U20608 ( .A1(n15706), .A2(n15105), .ZN(n20683) );
  OR2_X1 U20609 ( .A1(n20738), .A2(n20739), .ZN(n20682) );
  AND2_X1 U20610 ( .A1(n20672), .A2(n20671), .ZN(n20739) );
  AND2_X1 U20611 ( .A1(n20667), .A2(n20740), .ZN(n20738) );
  OR2_X1 U20612 ( .A1(n20671), .A2(n20672), .ZN(n20740) );
  OR2_X1 U20613 ( .A1(n15672), .A2(n15105), .ZN(n20672) );
  OR2_X1 U20614 ( .A1(n20741), .A2(n20742), .ZN(n20671) );
  AND2_X1 U20615 ( .A1(n20662), .A2(n20661), .ZN(n20742) );
  AND2_X1 U20616 ( .A1(n20656), .A2(n20743), .ZN(n20741) );
  OR2_X1 U20617 ( .A1(n20661), .A2(n20662), .ZN(n20743) );
  OR2_X1 U20618 ( .A1(n15638), .A2(n15105), .ZN(n20662) );
  OR2_X1 U20619 ( .A1(n20744), .A2(n20745), .ZN(n20661) );
  AND2_X1 U20620 ( .A1(n20648), .A2(n20650), .ZN(n20745) );
  AND2_X1 U20621 ( .A1(n20645), .A2(n20746), .ZN(n20744) );
  OR2_X1 U20622 ( .A1(n20650), .A2(n20648), .ZN(n20746) );
  OR2_X1 U20623 ( .A1(n15593), .A2(n15105), .ZN(n20648) );
  OR2_X1 U20624 ( .A1(n20747), .A2(n20748), .ZN(n20650) );
  AND2_X1 U20625 ( .A1(n20637), .A2(n20639), .ZN(n20748) );
  AND2_X1 U20626 ( .A1(n20634), .A2(n20749), .ZN(n20747) );
  OR2_X1 U20627 ( .A1(n20639), .A2(n20637), .ZN(n20749) );
  OR2_X1 U20628 ( .A1(n15559), .A2(n15105), .ZN(n20637) );
  OR2_X1 U20629 ( .A1(n20750), .A2(n20751), .ZN(n20639) );
  AND2_X1 U20630 ( .A1(n20626), .A2(n20628), .ZN(n20751) );
  AND2_X1 U20631 ( .A1(n20623), .A2(n20752), .ZN(n20750) );
  OR2_X1 U20632 ( .A1(n20628), .A2(n20626), .ZN(n20752) );
  OR2_X1 U20633 ( .A1(n15525), .A2(n15105), .ZN(n20626) );
  OR2_X1 U20634 ( .A1(n20753), .A2(n20754), .ZN(n20628) );
  AND2_X1 U20635 ( .A1(n20615), .A2(n20617), .ZN(n20754) );
  AND2_X1 U20636 ( .A1(n20612), .A2(n20755), .ZN(n20753) );
  OR2_X1 U20637 ( .A1(n20617), .A2(n20615), .ZN(n20755) );
  OR2_X1 U20638 ( .A1(n15491), .A2(n15105), .ZN(n20615) );
  OR2_X1 U20639 ( .A1(n20756), .A2(n20757), .ZN(n20617) );
  AND2_X1 U20640 ( .A1(n20604), .A2(n20606), .ZN(n20757) );
  AND2_X1 U20641 ( .A1(n20601), .A2(n20758), .ZN(n20756) );
  OR2_X1 U20642 ( .A1(n20606), .A2(n20604), .ZN(n20758) );
  OR2_X1 U20643 ( .A1(n15457), .A2(n15105), .ZN(n20604) );
  OR2_X1 U20644 ( .A1(n20759), .A2(n20760), .ZN(n20606) );
  AND2_X1 U20645 ( .A1(n20593), .A2(n20595), .ZN(n20760) );
  AND2_X1 U20646 ( .A1(n20590), .A2(n20761), .ZN(n20759) );
  OR2_X1 U20647 ( .A1(n20595), .A2(n20593), .ZN(n20761) );
  OR2_X1 U20648 ( .A1(n15423), .A2(n15105), .ZN(n20593) );
  OR2_X1 U20649 ( .A1(n20762), .A2(n20763), .ZN(n20595) );
  AND2_X1 U20650 ( .A1(n20582), .A2(n20584), .ZN(n20763) );
  AND2_X1 U20651 ( .A1(n20579), .A2(n20764), .ZN(n20762) );
  OR2_X1 U20652 ( .A1(n20584), .A2(n20582), .ZN(n20764) );
  OR2_X1 U20653 ( .A1(n15389), .A2(n15105), .ZN(n20582) );
  OR2_X1 U20654 ( .A1(n20765), .A2(n20766), .ZN(n20584) );
  AND2_X1 U20655 ( .A1(n20571), .A2(n20573), .ZN(n20766) );
  AND2_X1 U20656 ( .A1(n20568), .A2(n20767), .ZN(n20765) );
  OR2_X1 U20657 ( .A1(n20573), .A2(n20571), .ZN(n20767) );
  OR2_X1 U20658 ( .A1(n15355), .A2(n15105), .ZN(n20571) );
  OR2_X1 U20659 ( .A1(n20768), .A2(n20769), .ZN(n20573) );
  AND2_X1 U20660 ( .A1(n20560), .A2(n20562), .ZN(n20769) );
  AND2_X1 U20661 ( .A1(n20557), .A2(n20770), .ZN(n20768) );
  OR2_X1 U20662 ( .A1(n20562), .A2(n20560), .ZN(n20770) );
  OR2_X1 U20663 ( .A1(n15321), .A2(n15105), .ZN(n20560) );
  OR2_X1 U20664 ( .A1(n20771), .A2(n20772), .ZN(n20562) );
  AND2_X1 U20665 ( .A1(n20549), .A2(n20551), .ZN(n20772) );
  AND2_X1 U20666 ( .A1(n20546), .A2(n20773), .ZN(n20771) );
  OR2_X1 U20667 ( .A1(n20551), .A2(n20549), .ZN(n20773) );
  OR2_X1 U20668 ( .A1(n15287), .A2(n15105), .ZN(n20549) );
  OR2_X1 U20669 ( .A1(n20774), .A2(n20775), .ZN(n20551) );
  AND2_X1 U20670 ( .A1(n20538), .A2(n20540), .ZN(n20775) );
  AND2_X1 U20671 ( .A1(n20535), .A2(n20776), .ZN(n20774) );
  OR2_X1 U20672 ( .A1(n20540), .A2(n20538), .ZN(n20776) );
  OR2_X1 U20673 ( .A1(n15242), .A2(n15105), .ZN(n20538) );
  OR2_X1 U20674 ( .A1(n20777), .A2(n20778), .ZN(n20540) );
  AND2_X1 U20675 ( .A1(n20527), .A2(n20529), .ZN(n20778) );
  AND2_X1 U20676 ( .A1(n20524), .A2(n20779), .ZN(n20777) );
  OR2_X1 U20677 ( .A1(n20529), .A2(n20527), .ZN(n20779) );
  OR2_X1 U20678 ( .A1(n15208), .A2(n15105), .ZN(n20527) );
  OR2_X1 U20679 ( .A1(n20780), .A2(n20781), .ZN(n20529) );
  AND2_X1 U20680 ( .A1(n20516), .A2(n20518), .ZN(n20781) );
  AND2_X1 U20681 ( .A1(n20513), .A2(n20782), .ZN(n20780) );
  OR2_X1 U20682 ( .A1(n20518), .A2(n20516), .ZN(n20782) );
  OR2_X1 U20683 ( .A1(n15174), .A2(n15105), .ZN(n20516) );
  OR2_X1 U20684 ( .A1(n20783), .A2(n20784), .ZN(n20518) );
  AND2_X1 U20685 ( .A1(n20505), .A2(n20507), .ZN(n20784) );
  AND2_X1 U20686 ( .A1(n20502), .A2(n20785), .ZN(n20783) );
  OR2_X1 U20687 ( .A1(n20507), .A2(n20505), .ZN(n20785) );
  OR2_X1 U20688 ( .A1(n15140), .A2(n15105), .ZN(n20505) );
  OR2_X1 U20689 ( .A1(n20786), .A2(n20787), .ZN(n20507) );
  AND2_X1 U20690 ( .A1(n15933), .A2(n20496), .ZN(n20787) );
  AND2_X1 U20691 ( .A1(n20492), .A2(n20788), .ZN(n20786) );
  OR2_X1 U20692 ( .A1(n20496), .A2(n15933), .ZN(n20788) );
  OR2_X1 U20693 ( .A1(n15106), .A2(n15105), .ZN(n15933) );
  OR2_X1 U20694 ( .A1(n20789), .A2(n20790), .ZN(n20496) );
  AND2_X1 U20695 ( .A1(n20484), .A2(n20486), .ZN(n20790) );
  AND2_X1 U20696 ( .A1(n20481), .A2(n20791), .ZN(n20789) );
  OR2_X1 U20697 ( .A1(n20486), .A2(n20484), .ZN(n20791) );
  OR2_X1 U20698 ( .A1(n15072), .A2(n15105), .ZN(n20484) );
  OR2_X1 U20699 ( .A1(n20792), .A2(n20793), .ZN(n20486) );
  AND2_X1 U20700 ( .A1(n20473), .A2(n20475), .ZN(n20793) );
  AND2_X1 U20701 ( .A1(n20470), .A2(n20794), .ZN(n20792) );
  OR2_X1 U20702 ( .A1(n20475), .A2(n20473), .ZN(n20794) );
  OR2_X1 U20703 ( .A1(n15038), .A2(n15105), .ZN(n20473) );
  OR2_X1 U20704 ( .A1(n20795), .A2(n20796), .ZN(n20475) );
  AND2_X1 U20705 ( .A1(n20462), .A2(n20464), .ZN(n20796) );
  AND2_X1 U20706 ( .A1(n20459), .A2(n20797), .ZN(n20795) );
  OR2_X1 U20707 ( .A1(n20464), .A2(n20462), .ZN(n20797) );
  OR2_X1 U20708 ( .A1(n15004), .A2(n15105), .ZN(n20462) );
  OR2_X1 U20709 ( .A1(n20798), .A2(n20799), .ZN(n20464) );
  AND2_X1 U20710 ( .A1(n20451), .A2(n20453), .ZN(n20799) );
  AND2_X1 U20711 ( .A1(n20448), .A2(n20800), .ZN(n20798) );
  OR2_X1 U20712 ( .A1(n20453), .A2(n20451), .ZN(n20800) );
  OR2_X1 U20713 ( .A1(n14970), .A2(n15105), .ZN(n20451) );
  OR2_X1 U20714 ( .A1(n20801), .A2(n20802), .ZN(n20453) );
  AND2_X1 U20715 ( .A1(n20440), .A2(n20442), .ZN(n20802) );
  AND2_X1 U20716 ( .A1(n20437), .A2(n20803), .ZN(n20801) );
  OR2_X1 U20717 ( .A1(n20442), .A2(n20440), .ZN(n20803) );
  OR2_X1 U20718 ( .A1(n14936), .A2(n15105), .ZN(n20440) );
  OR2_X1 U20719 ( .A1(n20804), .A2(n20805), .ZN(n20442) );
  AND2_X1 U20720 ( .A1(n20429), .A2(n20431), .ZN(n20805) );
  AND2_X1 U20721 ( .A1(n20426), .A2(n20806), .ZN(n20804) );
  OR2_X1 U20722 ( .A1(n20431), .A2(n20429), .ZN(n20806) );
  OR2_X1 U20723 ( .A1(n14891), .A2(n15105), .ZN(n20429) );
  OR2_X1 U20724 ( .A1(n20807), .A2(n20808), .ZN(n20431) );
  AND2_X1 U20725 ( .A1(n20414), .A2(n20419), .ZN(n20808) );
  AND2_X1 U20726 ( .A1(n20418), .A2(n20809), .ZN(n20807) );
  OR2_X1 U20727 ( .A1(n20419), .A2(n20414), .ZN(n20809) );
  OR2_X1 U20728 ( .A1(n14857), .A2(n15105), .ZN(n20414) );
  INV_X1 U20729 ( .A(b_22_), .ZN(n15105) );
  INV_X1 U20730 ( .A(n20420), .ZN(n20419) );
  AND3_X1 U20731 ( .A1(b_22_), .A2(b_21_), .A3(n15957), .ZN(n20420) );
  INV_X1 U20732 ( .A(n20421), .ZN(n20418) );
  OR2_X1 U20733 ( .A1(n20810), .A2(n20811), .ZN(n20421) );
  AND2_X1 U20734 ( .A1(b_21_), .A2(n20812), .ZN(n20811) );
  OR2_X1 U20735 ( .A1(n20813), .A2(n16981), .ZN(n20812) );
  AND2_X1 U20736 ( .A1(a_30_), .A2(n15173), .ZN(n20813) );
  AND2_X1 U20737 ( .A1(b_20_), .A2(n20814), .ZN(n20810) );
  OR2_X1 U20738 ( .A1(n20815), .A2(n14817), .ZN(n20814) );
  AND2_X1 U20739 ( .A1(a_31_), .A2(n15139), .ZN(n20815) );
  OR2_X1 U20740 ( .A1(n20816), .A2(n20817), .ZN(n20426) );
  AND2_X1 U20741 ( .A1(n20818), .A2(n20819), .ZN(n20817) );
  INV_X1 U20742 ( .A(n20820), .ZN(n20816) );
  OR2_X1 U20743 ( .A1(n20818), .A2(n20819), .ZN(n20820) );
  OR2_X1 U20744 ( .A1(n20821), .A2(n20822), .ZN(n20818) );
  AND2_X1 U20745 ( .A1(n20823), .A2(n20824), .ZN(n20822) );
  AND2_X1 U20746 ( .A1(n20825), .A2(n20826), .ZN(n20821) );
  OR2_X1 U20747 ( .A1(n20827), .A2(n20828), .ZN(n20437) );
  INV_X1 U20748 ( .A(n20829), .ZN(n20828) );
  OR2_X1 U20749 ( .A1(n20830), .A2(n20831), .ZN(n20829) );
  AND2_X1 U20750 ( .A1(n20831), .A2(n20830), .ZN(n20827) );
  AND2_X1 U20751 ( .A1(n20832), .A2(n20833), .ZN(n20830) );
  OR2_X1 U20752 ( .A1(n20834), .A2(n20835), .ZN(n20833) );
  INV_X1 U20753 ( .A(n20836), .ZN(n20835) );
  OR2_X1 U20754 ( .A1(n20836), .A2(n20837), .ZN(n20832) );
  INV_X1 U20755 ( .A(n20834), .ZN(n20837) );
  OR2_X1 U20756 ( .A1(n20838), .A2(n20839), .ZN(n20448) );
  INV_X1 U20757 ( .A(n20840), .ZN(n20839) );
  OR2_X1 U20758 ( .A1(n20841), .A2(n20842), .ZN(n20840) );
  AND2_X1 U20759 ( .A1(n20842), .A2(n20841), .ZN(n20838) );
  AND2_X1 U20760 ( .A1(n20843), .A2(n20844), .ZN(n20841) );
  OR2_X1 U20761 ( .A1(n20845), .A2(n20846), .ZN(n20844) );
  INV_X1 U20762 ( .A(n20847), .ZN(n20846) );
  OR2_X1 U20763 ( .A1(n20847), .A2(n20848), .ZN(n20843) );
  INV_X1 U20764 ( .A(n20845), .ZN(n20848) );
  OR2_X1 U20765 ( .A1(n20849), .A2(n20850), .ZN(n20459) );
  INV_X1 U20766 ( .A(n20851), .ZN(n20850) );
  OR2_X1 U20767 ( .A1(n20852), .A2(n20853), .ZN(n20851) );
  AND2_X1 U20768 ( .A1(n20853), .A2(n20852), .ZN(n20849) );
  AND2_X1 U20769 ( .A1(n20854), .A2(n20855), .ZN(n20852) );
  OR2_X1 U20770 ( .A1(n20856), .A2(n20857), .ZN(n20855) );
  INV_X1 U20771 ( .A(n20858), .ZN(n20857) );
  OR2_X1 U20772 ( .A1(n20858), .A2(n20859), .ZN(n20854) );
  INV_X1 U20773 ( .A(n20856), .ZN(n20859) );
  OR2_X1 U20774 ( .A1(n20860), .A2(n20861), .ZN(n20470) );
  INV_X1 U20775 ( .A(n20862), .ZN(n20861) );
  OR2_X1 U20776 ( .A1(n20863), .A2(n20864), .ZN(n20862) );
  AND2_X1 U20777 ( .A1(n20864), .A2(n20863), .ZN(n20860) );
  AND2_X1 U20778 ( .A1(n20865), .A2(n20866), .ZN(n20863) );
  OR2_X1 U20779 ( .A1(n20867), .A2(n20868), .ZN(n20866) );
  INV_X1 U20780 ( .A(n20869), .ZN(n20868) );
  OR2_X1 U20781 ( .A1(n20869), .A2(n20870), .ZN(n20865) );
  INV_X1 U20782 ( .A(n20867), .ZN(n20870) );
  OR2_X1 U20783 ( .A1(n20871), .A2(n20872), .ZN(n20481) );
  INV_X1 U20784 ( .A(n20873), .ZN(n20872) );
  OR2_X1 U20785 ( .A1(n20874), .A2(n20875), .ZN(n20873) );
  AND2_X1 U20786 ( .A1(n20875), .A2(n20874), .ZN(n20871) );
  AND2_X1 U20787 ( .A1(n20876), .A2(n20877), .ZN(n20874) );
  OR2_X1 U20788 ( .A1(n20878), .A2(n20879), .ZN(n20877) );
  INV_X1 U20789 ( .A(n20880), .ZN(n20879) );
  OR2_X1 U20790 ( .A1(n20880), .A2(n20881), .ZN(n20876) );
  INV_X1 U20791 ( .A(n20878), .ZN(n20881) );
  OR2_X1 U20792 ( .A1(n20882), .A2(n20883), .ZN(n20492) );
  INV_X1 U20793 ( .A(n20884), .ZN(n20883) );
  OR2_X1 U20794 ( .A1(n20885), .A2(n20886), .ZN(n20884) );
  AND2_X1 U20795 ( .A1(n20886), .A2(n20885), .ZN(n20882) );
  AND2_X1 U20796 ( .A1(n20887), .A2(n20888), .ZN(n20885) );
  OR2_X1 U20797 ( .A1(n20889), .A2(n20890), .ZN(n20888) );
  INV_X1 U20798 ( .A(n20891), .ZN(n20890) );
  OR2_X1 U20799 ( .A1(n20891), .A2(n20892), .ZN(n20887) );
  INV_X1 U20800 ( .A(n20889), .ZN(n20892) );
  OR2_X1 U20801 ( .A1(n20893), .A2(n20894), .ZN(n20502) );
  INV_X1 U20802 ( .A(n20895), .ZN(n20894) );
  OR2_X1 U20803 ( .A1(n20896), .A2(n20897), .ZN(n20895) );
  AND2_X1 U20804 ( .A1(n20897), .A2(n20896), .ZN(n20893) );
  AND2_X1 U20805 ( .A1(n20898), .A2(n20899), .ZN(n20896) );
  OR2_X1 U20806 ( .A1(n20900), .A2(n20901), .ZN(n20899) );
  INV_X1 U20807 ( .A(n20902), .ZN(n20901) );
  OR2_X1 U20808 ( .A1(n20902), .A2(n20903), .ZN(n20898) );
  INV_X1 U20809 ( .A(n20900), .ZN(n20903) );
  OR2_X1 U20810 ( .A1(n20904), .A2(n20905), .ZN(n20513) );
  INV_X1 U20811 ( .A(n20906), .ZN(n20905) );
  OR2_X1 U20812 ( .A1(n20907), .A2(n20908), .ZN(n20906) );
  AND2_X1 U20813 ( .A1(n20908), .A2(n20907), .ZN(n20904) );
  AND2_X1 U20814 ( .A1(n20909), .A2(n20910), .ZN(n20907) );
  OR2_X1 U20815 ( .A1(n15930), .A2(n20911), .ZN(n20910) );
  INV_X1 U20816 ( .A(n20912), .ZN(n20911) );
  OR2_X1 U20817 ( .A1(n20912), .A2(n20913), .ZN(n20909) );
  INV_X1 U20818 ( .A(n15930), .ZN(n20913) );
  OR2_X1 U20819 ( .A1(n20914), .A2(n20915), .ZN(n20524) );
  INV_X1 U20820 ( .A(n20916), .ZN(n20915) );
  OR2_X1 U20821 ( .A1(n20917), .A2(n20918), .ZN(n20916) );
  AND2_X1 U20822 ( .A1(n20918), .A2(n20917), .ZN(n20914) );
  AND2_X1 U20823 ( .A1(n20919), .A2(n20920), .ZN(n20917) );
  OR2_X1 U20824 ( .A1(n20921), .A2(n20922), .ZN(n20920) );
  INV_X1 U20825 ( .A(n20923), .ZN(n20922) );
  OR2_X1 U20826 ( .A1(n20923), .A2(n20924), .ZN(n20919) );
  INV_X1 U20827 ( .A(n20921), .ZN(n20924) );
  OR2_X1 U20828 ( .A1(n20925), .A2(n20926), .ZN(n20535) );
  INV_X1 U20829 ( .A(n20927), .ZN(n20926) );
  OR2_X1 U20830 ( .A1(n20928), .A2(n20929), .ZN(n20927) );
  AND2_X1 U20831 ( .A1(n20929), .A2(n20928), .ZN(n20925) );
  AND2_X1 U20832 ( .A1(n20930), .A2(n20931), .ZN(n20928) );
  OR2_X1 U20833 ( .A1(n20932), .A2(n20933), .ZN(n20931) );
  INV_X1 U20834 ( .A(n20934), .ZN(n20933) );
  OR2_X1 U20835 ( .A1(n20934), .A2(n20935), .ZN(n20930) );
  INV_X1 U20836 ( .A(n20932), .ZN(n20935) );
  OR2_X1 U20837 ( .A1(n20936), .A2(n20937), .ZN(n20546) );
  INV_X1 U20838 ( .A(n20938), .ZN(n20937) );
  OR2_X1 U20839 ( .A1(n20939), .A2(n20940), .ZN(n20938) );
  AND2_X1 U20840 ( .A1(n20940), .A2(n20939), .ZN(n20936) );
  AND2_X1 U20841 ( .A1(n20941), .A2(n20942), .ZN(n20939) );
  OR2_X1 U20842 ( .A1(n20943), .A2(n20944), .ZN(n20942) );
  INV_X1 U20843 ( .A(n20945), .ZN(n20944) );
  OR2_X1 U20844 ( .A1(n20945), .A2(n20946), .ZN(n20941) );
  INV_X1 U20845 ( .A(n20943), .ZN(n20946) );
  OR2_X1 U20846 ( .A1(n20947), .A2(n20948), .ZN(n20557) );
  INV_X1 U20847 ( .A(n20949), .ZN(n20948) );
  OR2_X1 U20848 ( .A1(n20950), .A2(n20951), .ZN(n20949) );
  AND2_X1 U20849 ( .A1(n20951), .A2(n20950), .ZN(n20947) );
  AND2_X1 U20850 ( .A1(n20952), .A2(n20953), .ZN(n20950) );
  OR2_X1 U20851 ( .A1(n20954), .A2(n20955), .ZN(n20953) );
  INV_X1 U20852 ( .A(n20956), .ZN(n20955) );
  OR2_X1 U20853 ( .A1(n20956), .A2(n20957), .ZN(n20952) );
  INV_X1 U20854 ( .A(n20954), .ZN(n20957) );
  OR2_X1 U20855 ( .A1(n20958), .A2(n20959), .ZN(n20568) );
  INV_X1 U20856 ( .A(n20960), .ZN(n20959) );
  OR2_X1 U20857 ( .A1(n20961), .A2(n20962), .ZN(n20960) );
  AND2_X1 U20858 ( .A1(n20962), .A2(n20961), .ZN(n20958) );
  AND2_X1 U20859 ( .A1(n20963), .A2(n20964), .ZN(n20961) );
  OR2_X1 U20860 ( .A1(n20965), .A2(n20966), .ZN(n20964) );
  INV_X1 U20861 ( .A(n20967), .ZN(n20966) );
  OR2_X1 U20862 ( .A1(n20967), .A2(n20968), .ZN(n20963) );
  INV_X1 U20863 ( .A(n20965), .ZN(n20968) );
  OR2_X1 U20864 ( .A1(n20969), .A2(n20970), .ZN(n20579) );
  INV_X1 U20865 ( .A(n20971), .ZN(n20970) );
  OR2_X1 U20866 ( .A1(n20972), .A2(n20973), .ZN(n20971) );
  AND2_X1 U20867 ( .A1(n20973), .A2(n20972), .ZN(n20969) );
  AND2_X1 U20868 ( .A1(n20974), .A2(n20975), .ZN(n20972) );
  OR2_X1 U20869 ( .A1(n20976), .A2(n20977), .ZN(n20975) );
  INV_X1 U20870 ( .A(n20978), .ZN(n20977) );
  OR2_X1 U20871 ( .A1(n20978), .A2(n20979), .ZN(n20974) );
  INV_X1 U20872 ( .A(n20976), .ZN(n20979) );
  OR2_X1 U20873 ( .A1(n20980), .A2(n20981), .ZN(n20590) );
  INV_X1 U20874 ( .A(n20982), .ZN(n20981) );
  OR2_X1 U20875 ( .A1(n20983), .A2(n20984), .ZN(n20982) );
  AND2_X1 U20876 ( .A1(n20984), .A2(n20983), .ZN(n20980) );
  AND2_X1 U20877 ( .A1(n20985), .A2(n20986), .ZN(n20983) );
  OR2_X1 U20878 ( .A1(n20987), .A2(n20988), .ZN(n20986) );
  INV_X1 U20879 ( .A(n20989), .ZN(n20988) );
  OR2_X1 U20880 ( .A1(n20989), .A2(n20990), .ZN(n20985) );
  INV_X1 U20881 ( .A(n20987), .ZN(n20990) );
  OR2_X1 U20882 ( .A1(n20991), .A2(n20992), .ZN(n20601) );
  INV_X1 U20883 ( .A(n20993), .ZN(n20992) );
  OR2_X1 U20884 ( .A1(n20994), .A2(n20995), .ZN(n20993) );
  AND2_X1 U20885 ( .A1(n20995), .A2(n20994), .ZN(n20991) );
  AND2_X1 U20886 ( .A1(n20996), .A2(n20997), .ZN(n20994) );
  OR2_X1 U20887 ( .A1(n20998), .A2(n20999), .ZN(n20997) );
  INV_X1 U20888 ( .A(n21000), .ZN(n20999) );
  OR2_X1 U20889 ( .A1(n21000), .A2(n21001), .ZN(n20996) );
  INV_X1 U20890 ( .A(n20998), .ZN(n21001) );
  OR2_X1 U20891 ( .A1(n21002), .A2(n21003), .ZN(n20612) );
  INV_X1 U20892 ( .A(n21004), .ZN(n21003) );
  OR2_X1 U20893 ( .A1(n21005), .A2(n21006), .ZN(n21004) );
  AND2_X1 U20894 ( .A1(n21006), .A2(n21005), .ZN(n21002) );
  AND2_X1 U20895 ( .A1(n21007), .A2(n21008), .ZN(n21005) );
  OR2_X1 U20896 ( .A1(n21009), .A2(n21010), .ZN(n21008) );
  INV_X1 U20897 ( .A(n21011), .ZN(n21010) );
  OR2_X1 U20898 ( .A1(n21011), .A2(n21012), .ZN(n21007) );
  INV_X1 U20899 ( .A(n21009), .ZN(n21012) );
  OR2_X1 U20900 ( .A1(n21013), .A2(n21014), .ZN(n20623) );
  INV_X1 U20901 ( .A(n21015), .ZN(n21014) );
  OR2_X1 U20902 ( .A1(n21016), .A2(n21017), .ZN(n21015) );
  AND2_X1 U20903 ( .A1(n21017), .A2(n21016), .ZN(n21013) );
  AND2_X1 U20904 ( .A1(n21018), .A2(n21019), .ZN(n21016) );
  OR2_X1 U20905 ( .A1(n21020), .A2(n21021), .ZN(n21019) );
  INV_X1 U20906 ( .A(n21022), .ZN(n21021) );
  OR2_X1 U20907 ( .A1(n21022), .A2(n21023), .ZN(n21018) );
  INV_X1 U20908 ( .A(n21020), .ZN(n21023) );
  OR2_X1 U20909 ( .A1(n21024), .A2(n21025), .ZN(n20634) );
  INV_X1 U20910 ( .A(n21026), .ZN(n21025) );
  OR2_X1 U20911 ( .A1(n21027), .A2(n21028), .ZN(n21026) );
  AND2_X1 U20912 ( .A1(n21028), .A2(n21027), .ZN(n21024) );
  AND2_X1 U20913 ( .A1(n21029), .A2(n21030), .ZN(n21027) );
  OR2_X1 U20914 ( .A1(n21031), .A2(n21032), .ZN(n21030) );
  INV_X1 U20915 ( .A(n21033), .ZN(n21032) );
  OR2_X1 U20916 ( .A1(n21033), .A2(n21034), .ZN(n21029) );
  INV_X1 U20917 ( .A(n21031), .ZN(n21034) );
  OR2_X1 U20918 ( .A1(n21035), .A2(n21036), .ZN(n20645) );
  INV_X1 U20919 ( .A(n21037), .ZN(n21036) );
  OR2_X1 U20920 ( .A1(n21038), .A2(n21039), .ZN(n21037) );
  AND2_X1 U20921 ( .A1(n21039), .A2(n21038), .ZN(n21035) );
  AND2_X1 U20922 ( .A1(n21040), .A2(n21041), .ZN(n21038) );
  OR2_X1 U20923 ( .A1(n21042), .A2(n21043), .ZN(n21041) );
  INV_X1 U20924 ( .A(n21044), .ZN(n21043) );
  OR2_X1 U20925 ( .A1(n21044), .A2(n21045), .ZN(n21040) );
  INV_X1 U20926 ( .A(n21042), .ZN(n21045) );
  OR2_X1 U20927 ( .A1(n21046), .A2(n21047), .ZN(n20656) );
  INV_X1 U20928 ( .A(n21048), .ZN(n21047) );
  OR2_X1 U20929 ( .A1(n21049), .A2(n21050), .ZN(n21048) );
  AND2_X1 U20930 ( .A1(n21050), .A2(n21049), .ZN(n21046) );
  AND2_X1 U20931 ( .A1(n21051), .A2(n21052), .ZN(n21049) );
  INV_X1 U20932 ( .A(n21053), .ZN(n21052) );
  AND2_X1 U20933 ( .A1(n21054), .A2(n21055), .ZN(n21053) );
  OR2_X1 U20934 ( .A1(n21055), .A2(n21054), .ZN(n21051) );
  INV_X1 U20935 ( .A(n21056), .ZN(n21054) );
  AND2_X1 U20936 ( .A1(n21057), .A2(n21058), .ZN(n20667) );
  INV_X1 U20937 ( .A(n21059), .ZN(n21058) );
  AND2_X1 U20938 ( .A1(n21060), .A2(n21061), .ZN(n21059) );
  OR2_X1 U20939 ( .A1(n21061), .A2(n21060), .ZN(n21057) );
  OR2_X1 U20940 ( .A1(n21062), .A2(n21063), .ZN(n21060) );
  AND2_X1 U20941 ( .A1(n21064), .A2(n21065), .ZN(n21063) );
  INV_X1 U20942 ( .A(n21066), .ZN(n21064) );
  AND2_X1 U20943 ( .A1(n21067), .A2(n21066), .ZN(n21062) );
  INV_X1 U20944 ( .A(n21065), .ZN(n21067) );
  AND2_X1 U20945 ( .A1(n21068), .A2(n21069), .ZN(n20678) );
  INV_X1 U20946 ( .A(n21070), .ZN(n21069) );
  AND2_X1 U20947 ( .A1(n21071), .A2(n21072), .ZN(n21070) );
  OR2_X1 U20948 ( .A1(n21072), .A2(n21071), .ZN(n21068) );
  OR2_X1 U20949 ( .A1(n21073), .A2(n21074), .ZN(n21071) );
  AND2_X1 U20950 ( .A1(n21075), .A2(n21076), .ZN(n21074) );
  INV_X1 U20951 ( .A(n21077), .ZN(n21075) );
  AND2_X1 U20952 ( .A1(n21078), .A2(n21077), .ZN(n21073) );
  INV_X1 U20953 ( .A(n21076), .ZN(n21078) );
  AND2_X1 U20954 ( .A1(n21079), .A2(n21080), .ZN(n20689) );
  INV_X1 U20955 ( .A(n21081), .ZN(n21080) );
  AND2_X1 U20956 ( .A1(n21082), .A2(n21083), .ZN(n21081) );
  OR2_X1 U20957 ( .A1(n21083), .A2(n21082), .ZN(n21079) );
  OR2_X1 U20958 ( .A1(n21084), .A2(n21085), .ZN(n21082) );
  AND2_X1 U20959 ( .A1(n21086), .A2(n21087), .ZN(n21085) );
  INV_X1 U20960 ( .A(n21088), .ZN(n21086) );
  AND2_X1 U20961 ( .A1(n21089), .A2(n21088), .ZN(n21084) );
  INV_X1 U20962 ( .A(n21087), .ZN(n21089) );
  AND2_X1 U20963 ( .A1(n21090), .A2(n21091), .ZN(n20700) );
  INV_X1 U20964 ( .A(n21092), .ZN(n21091) );
  AND2_X1 U20965 ( .A1(n21093), .A2(n21094), .ZN(n21092) );
  OR2_X1 U20966 ( .A1(n21094), .A2(n21093), .ZN(n21090) );
  OR2_X1 U20967 ( .A1(n21095), .A2(n21096), .ZN(n21093) );
  AND2_X1 U20968 ( .A1(n21097), .A2(n21098), .ZN(n21096) );
  INV_X1 U20969 ( .A(n21099), .ZN(n21097) );
  AND2_X1 U20970 ( .A1(n21100), .A2(n21099), .ZN(n21095) );
  INV_X1 U20971 ( .A(n21098), .ZN(n21100) );
  AND2_X1 U20972 ( .A1(n21101), .A2(n21102), .ZN(n20711) );
  INV_X1 U20973 ( .A(n21103), .ZN(n21102) );
  AND2_X1 U20974 ( .A1(n21104), .A2(n21105), .ZN(n21103) );
  OR2_X1 U20975 ( .A1(n21105), .A2(n21104), .ZN(n21101) );
  OR2_X1 U20976 ( .A1(n21106), .A2(n21107), .ZN(n21104) );
  AND2_X1 U20977 ( .A1(n21108), .A2(n21109), .ZN(n21107) );
  INV_X1 U20978 ( .A(n21110), .ZN(n21108) );
  AND2_X1 U20979 ( .A1(n21111), .A2(n21110), .ZN(n21106) );
  INV_X1 U20980 ( .A(n21109), .ZN(n21111) );
  AND2_X1 U20981 ( .A1(n21112), .A2(n21113), .ZN(n20274) );
  INV_X1 U20982 ( .A(n21114), .ZN(n21113) );
  AND2_X1 U20983 ( .A1(n21115), .A2(n20288), .ZN(n21114) );
  OR2_X1 U20984 ( .A1(n20288), .A2(n21115), .ZN(n21112) );
  OR2_X1 U20985 ( .A1(n21116), .A2(n21117), .ZN(n21115) );
  AND2_X1 U20986 ( .A1(n21118), .A2(n20287), .ZN(n21117) );
  INV_X1 U20987 ( .A(n20286), .ZN(n21118) );
  AND2_X1 U20988 ( .A1(n21119), .A2(n20286), .ZN(n21116) );
  OR2_X1 U20989 ( .A1(n15808), .A2(n15139), .ZN(n20286) );
  INV_X1 U20990 ( .A(n20287), .ZN(n21119) );
  OR2_X1 U20991 ( .A1(n21120), .A2(n21121), .ZN(n20287) );
  AND2_X1 U20992 ( .A1(n21110), .A2(n21109), .ZN(n21121) );
  AND2_X1 U20993 ( .A1(n21105), .A2(n21122), .ZN(n21120) );
  OR2_X1 U20994 ( .A1(n21110), .A2(n21109), .ZN(n21122) );
  OR2_X1 U20995 ( .A1(n21123), .A2(n21124), .ZN(n21109) );
  AND2_X1 U20996 ( .A1(n21099), .A2(n21098), .ZN(n21124) );
  AND2_X1 U20997 ( .A1(n21094), .A2(n21125), .ZN(n21123) );
  OR2_X1 U20998 ( .A1(n21099), .A2(n21098), .ZN(n21125) );
  OR2_X1 U20999 ( .A1(n21126), .A2(n21127), .ZN(n21098) );
  AND2_X1 U21000 ( .A1(n21088), .A2(n21087), .ZN(n21127) );
  AND2_X1 U21001 ( .A1(n21083), .A2(n21128), .ZN(n21126) );
  OR2_X1 U21002 ( .A1(n21088), .A2(n21087), .ZN(n21128) );
  OR2_X1 U21003 ( .A1(n21129), .A2(n21130), .ZN(n21087) );
  AND2_X1 U21004 ( .A1(n21077), .A2(n21076), .ZN(n21130) );
  AND2_X1 U21005 ( .A1(n21072), .A2(n21131), .ZN(n21129) );
  OR2_X1 U21006 ( .A1(n21077), .A2(n21076), .ZN(n21131) );
  OR2_X1 U21007 ( .A1(n21132), .A2(n21133), .ZN(n21076) );
  AND2_X1 U21008 ( .A1(n21066), .A2(n21065), .ZN(n21133) );
  AND2_X1 U21009 ( .A1(n21061), .A2(n21134), .ZN(n21132) );
  OR2_X1 U21010 ( .A1(n21066), .A2(n21065), .ZN(n21134) );
  OR2_X1 U21011 ( .A1(n21135), .A2(n21136), .ZN(n21065) );
  AND2_X1 U21012 ( .A1(n21056), .A2(n21055), .ZN(n21136) );
  AND2_X1 U21013 ( .A1(n21050), .A2(n21137), .ZN(n21135) );
  OR2_X1 U21014 ( .A1(n21056), .A2(n21055), .ZN(n21137) );
  OR2_X1 U21015 ( .A1(n21138), .A2(n21139), .ZN(n21055) );
  AND2_X1 U21016 ( .A1(n21042), .A2(n21044), .ZN(n21139) );
  AND2_X1 U21017 ( .A1(n21039), .A2(n21140), .ZN(n21138) );
  OR2_X1 U21018 ( .A1(n21042), .A2(n21044), .ZN(n21140) );
  OR2_X1 U21019 ( .A1(n21141), .A2(n21142), .ZN(n21044) );
  AND2_X1 U21020 ( .A1(n21031), .A2(n21033), .ZN(n21142) );
  AND2_X1 U21021 ( .A1(n21028), .A2(n21143), .ZN(n21141) );
  OR2_X1 U21022 ( .A1(n21031), .A2(n21033), .ZN(n21143) );
  OR2_X1 U21023 ( .A1(n21144), .A2(n21145), .ZN(n21033) );
  AND2_X1 U21024 ( .A1(n21020), .A2(n21022), .ZN(n21145) );
  AND2_X1 U21025 ( .A1(n21017), .A2(n21146), .ZN(n21144) );
  OR2_X1 U21026 ( .A1(n21020), .A2(n21022), .ZN(n21146) );
  OR2_X1 U21027 ( .A1(n21147), .A2(n21148), .ZN(n21022) );
  AND2_X1 U21028 ( .A1(n21009), .A2(n21011), .ZN(n21148) );
  AND2_X1 U21029 ( .A1(n21006), .A2(n21149), .ZN(n21147) );
  OR2_X1 U21030 ( .A1(n21009), .A2(n21011), .ZN(n21149) );
  OR2_X1 U21031 ( .A1(n21150), .A2(n21151), .ZN(n21011) );
  AND2_X1 U21032 ( .A1(n20998), .A2(n21000), .ZN(n21151) );
  AND2_X1 U21033 ( .A1(n20995), .A2(n21152), .ZN(n21150) );
  OR2_X1 U21034 ( .A1(n20998), .A2(n21000), .ZN(n21152) );
  OR2_X1 U21035 ( .A1(n21153), .A2(n21154), .ZN(n21000) );
  AND2_X1 U21036 ( .A1(n20987), .A2(n20989), .ZN(n21154) );
  AND2_X1 U21037 ( .A1(n20984), .A2(n21155), .ZN(n21153) );
  OR2_X1 U21038 ( .A1(n20987), .A2(n20989), .ZN(n21155) );
  OR2_X1 U21039 ( .A1(n21156), .A2(n21157), .ZN(n20989) );
  AND2_X1 U21040 ( .A1(n20976), .A2(n20978), .ZN(n21157) );
  AND2_X1 U21041 ( .A1(n20973), .A2(n21158), .ZN(n21156) );
  OR2_X1 U21042 ( .A1(n20976), .A2(n20978), .ZN(n21158) );
  OR2_X1 U21043 ( .A1(n21159), .A2(n21160), .ZN(n20978) );
  AND2_X1 U21044 ( .A1(n20965), .A2(n20967), .ZN(n21160) );
  AND2_X1 U21045 ( .A1(n20962), .A2(n21161), .ZN(n21159) );
  OR2_X1 U21046 ( .A1(n20965), .A2(n20967), .ZN(n21161) );
  OR2_X1 U21047 ( .A1(n21162), .A2(n21163), .ZN(n20967) );
  AND2_X1 U21048 ( .A1(n20954), .A2(n20956), .ZN(n21163) );
  AND2_X1 U21049 ( .A1(n20951), .A2(n21164), .ZN(n21162) );
  OR2_X1 U21050 ( .A1(n20954), .A2(n20956), .ZN(n21164) );
  OR2_X1 U21051 ( .A1(n21165), .A2(n21166), .ZN(n20956) );
  AND2_X1 U21052 ( .A1(n20943), .A2(n20945), .ZN(n21166) );
  AND2_X1 U21053 ( .A1(n20940), .A2(n21167), .ZN(n21165) );
  OR2_X1 U21054 ( .A1(n20943), .A2(n20945), .ZN(n21167) );
  OR2_X1 U21055 ( .A1(n21168), .A2(n21169), .ZN(n20945) );
  AND2_X1 U21056 ( .A1(n20932), .A2(n20934), .ZN(n21169) );
  AND2_X1 U21057 ( .A1(n20929), .A2(n21170), .ZN(n21168) );
  OR2_X1 U21058 ( .A1(n20932), .A2(n20934), .ZN(n21170) );
  OR2_X1 U21059 ( .A1(n21171), .A2(n21172), .ZN(n20934) );
  AND2_X1 U21060 ( .A1(n20921), .A2(n20923), .ZN(n21172) );
  AND2_X1 U21061 ( .A1(n20918), .A2(n21173), .ZN(n21171) );
  OR2_X1 U21062 ( .A1(n20921), .A2(n20923), .ZN(n21173) );
  OR2_X1 U21063 ( .A1(n21174), .A2(n21175), .ZN(n20923) );
  AND2_X1 U21064 ( .A1(n15930), .A2(n20912), .ZN(n21175) );
  AND2_X1 U21065 ( .A1(n20908), .A2(n21176), .ZN(n21174) );
  OR2_X1 U21066 ( .A1(n15930), .A2(n20912), .ZN(n21176) );
  OR2_X1 U21067 ( .A1(n21177), .A2(n21178), .ZN(n20912) );
  AND2_X1 U21068 ( .A1(n20900), .A2(n20902), .ZN(n21178) );
  AND2_X1 U21069 ( .A1(n20897), .A2(n21179), .ZN(n21177) );
  OR2_X1 U21070 ( .A1(n20900), .A2(n20902), .ZN(n21179) );
  OR2_X1 U21071 ( .A1(n21180), .A2(n21181), .ZN(n20902) );
  AND2_X1 U21072 ( .A1(n20889), .A2(n20891), .ZN(n21181) );
  AND2_X1 U21073 ( .A1(n20886), .A2(n21182), .ZN(n21180) );
  OR2_X1 U21074 ( .A1(n20889), .A2(n20891), .ZN(n21182) );
  OR2_X1 U21075 ( .A1(n21183), .A2(n21184), .ZN(n20891) );
  AND2_X1 U21076 ( .A1(n20878), .A2(n20880), .ZN(n21184) );
  AND2_X1 U21077 ( .A1(n20875), .A2(n21185), .ZN(n21183) );
  OR2_X1 U21078 ( .A1(n20878), .A2(n20880), .ZN(n21185) );
  OR2_X1 U21079 ( .A1(n21186), .A2(n21187), .ZN(n20880) );
  AND2_X1 U21080 ( .A1(n20867), .A2(n20869), .ZN(n21187) );
  AND2_X1 U21081 ( .A1(n20864), .A2(n21188), .ZN(n21186) );
  OR2_X1 U21082 ( .A1(n20867), .A2(n20869), .ZN(n21188) );
  OR2_X1 U21083 ( .A1(n21189), .A2(n21190), .ZN(n20869) );
  AND2_X1 U21084 ( .A1(n20856), .A2(n20858), .ZN(n21190) );
  AND2_X1 U21085 ( .A1(n20853), .A2(n21191), .ZN(n21189) );
  OR2_X1 U21086 ( .A1(n20856), .A2(n20858), .ZN(n21191) );
  OR2_X1 U21087 ( .A1(n21192), .A2(n21193), .ZN(n20858) );
  AND2_X1 U21088 ( .A1(n20845), .A2(n20847), .ZN(n21193) );
  AND2_X1 U21089 ( .A1(n20842), .A2(n21194), .ZN(n21192) );
  OR2_X1 U21090 ( .A1(n20845), .A2(n20847), .ZN(n21194) );
  OR2_X1 U21091 ( .A1(n21195), .A2(n21196), .ZN(n20847) );
  AND2_X1 U21092 ( .A1(n20834), .A2(n20836), .ZN(n21196) );
  AND2_X1 U21093 ( .A1(n20831), .A2(n21197), .ZN(n21195) );
  OR2_X1 U21094 ( .A1(n20834), .A2(n20836), .ZN(n21197) );
  OR2_X1 U21095 ( .A1(n21198), .A2(n21199), .ZN(n20836) );
  AND2_X1 U21096 ( .A1(n20819), .A2(n20824), .ZN(n21199) );
  AND2_X1 U21097 ( .A1(n20823), .A2(n21200), .ZN(n21198) );
  OR2_X1 U21098 ( .A1(n20819), .A2(n20824), .ZN(n21200) );
  INV_X1 U21099 ( .A(n20825), .ZN(n20824) );
  AND3_X1 U21100 ( .A1(b_21_), .A2(b_20_), .A3(n15957), .ZN(n20825) );
  OR2_X1 U21101 ( .A1(n14857), .A2(n15139), .ZN(n20819) );
  INV_X1 U21102 ( .A(n20826), .ZN(n20823) );
  OR2_X1 U21103 ( .A1(n21201), .A2(n21202), .ZN(n20826) );
  AND2_X1 U21104 ( .A1(b_20_), .A2(n21203), .ZN(n21202) );
  OR2_X1 U21105 ( .A1(n21204), .A2(n16981), .ZN(n21203) );
  AND2_X1 U21106 ( .A1(a_30_), .A2(n15207), .ZN(n21204) );
  AND2_X1 U21107 ( .A1(b_19_), .A2(n21205), .ZN(n21201) );
  OR2_X1 U21108 ( .A1(n21206), .A2(n14817), .ZN(n21205) );
  AND2_X1 U21109 ( .A1(a_31_), .A2(n15173), .ZN(n21206) );
  OR2_X1 U21110 ( .A1(n14891), .A2(n15139), .ZN(n20834) );
  OR2_X1 U21111 ( .A1(n21207), .A2(n21208), .ZN(n20831) );
  AND2_X1 U21112 ( .A1(n21209), .A2(n21210), .ZN(n21208) );
  INV_X1 U21113 ( .A(n21211), .ZN(n21207) );
  OR2_X1 U21114 ( .A1(n21209), .A2(n21210), .ZN(n21211) );
  OR2_X1 U21115 ( .A1(n21212), .A2(n21213), .ZN(n21209) );
  AND2_X1 U21116 ( .A1(n21214), .A2(n21215), .ZN(n21213) );
  AND2_X1 U21117 ( .A1(n21216), .A2(n21217), .ZN(n21212) );
  OR2_X1 U21118 ( .A1(n14936), .A2(n15139), .ZN(n20845) );
  OR2_X1 U21119 ( .A1(n21218), .A2(n21219), .ZN(n20842) );
  INV_X1 U21120 ( .A(n21220), .ZN(n21219) );
  OR2_X1 U21121 ( .A1(n21221), .A2(n21222), .ZN(n21220) );
  AND2_X1 U21122 ( .A1(n21222), .A2(n21221), .ZN(n21218) );
  AND2_X1 U21123 ( .A1(n21223), .A2(n21224), .ZN(n21221) );
  OR2_X1 U21124 ( .A1(n21225), .A2(n21226), .ZN(n21224) );
  INV_X1 U21125 ( .A(n21227), .ZN(n21226) );
  OR2_X1 U21126 ( .A1(n21227), .A2(n21228), .ZN(n21223) );
  INV_X1 U21127 ( .A(n21225), .ZN(n21228) );
  OR2_X1 U21128 ( .A1(n14970), .A2(n15139), .ZN(n20856) );
  OR2_X1 U21129 ( .A1(n21229), .A2(n21230), .ZN(n20853) );
  INV_X1 U21130 ( .A(n21231), .ZN(n21230) );
  OR2_X1 U21131 ( .A1(n21232), .A2(n21233), .ZN(n21231) );
  AND2_X1 U21132 ( .A1(n21233), .A2(n21232), .ZN(n21229) );
  AND2_X1 U21133 ( .A1(n21234), .A2(n21235), .ZN(n21232) );
  OR2_X1 U21134 ( .A1(n21236), .A2(n21237), .ZN(n21235) );
  INV_X1 U21135 ( .A(n21238), .ZN(n21237) );
  OR2_X1 U21136 ( .A1(n21238), .A2(n21239), .ZN(n21234) );
  INV_X1 U21137 ( .A(n21236), .ZN(n21239) );
  OR2_X1 U21138 ( .A1(n15004), .A2(n15139), .ZN(n20867) );
  OR2_X1 U21139 ( .A1(n21240), .A2(n21241), .ZN(n20864) );
  INV_X1 U21140 ( .A(n21242), .ZN(n21241) );
  OR2_X1 U21141 ( .A1(n21243), .A2(n21244), .ZN(n21242) );
  AND2_X1 U21142 ( .A1(n21244), .A2(n21243), .ZN(n21240) );
  AND2_X1 U21143 ( .A1(n21245), .A2(n21246), .ZN(n21243) );
  OR2_X1 U21144 ( .A1(n21247), .A2(n21248), .ZN(n21246) );
  INV_X1 U21145 ( .A(n21249), .ZN(n21248) );
  OR2_X1 U21146 ( .A1(n21249), .A2(n21250), .ZN(n21245) );
  INV_X1 U21147 ( .A(n21247), .ZN(n21250) );
  OR2_X1 U21148 ( .A1(n15038), .A2(n15139), .ZN(n20878) );
  OR2_X1 U21149 ( .A1(n21251), .A2(n21252), .ZN(n20875) );
  INV_X1 U21150 ( .A(n21253), .ZN(n21252) );
  OR2_X1 U21151 ( .A1(n21254), .A2(n21255), .ZN(n21253) );
  AND2_X1 U21152 ( .A1(n21255), .A2(n21254), .ZN(n21251) );
  AND2_X1 U21153 ( .A1(n21256), .A2(n21257), .ZN(n21254) );
  OR2_X1 U21154 ( .A1(n21258), .A2(n21259), .ZN(n21257) );
  INV_X1 U21155 ( .A(n21260), .ZN(n21259) );
  OR2_X1 U21156 ( .A1(n21260), .A2(n21261), .ZN(n21256) );
  INV_X1 U21157 ( .A(n21258), .ZN(n21261) );
  OR2_X1 U21158 ( .A1(n15072), .A2(n15139), .ZN(n20889) );
  OR2_X1 U21159 ( .A1(n21262), .A2(n21263), .ZN(n20886) );
  INV_X1 U21160 ( .A(n21264), .ZN(n21263) );
  OR2_X1 U21161 ( .A1(n21265), .A2(n21266), .ZN(n21264) );
  AND2_X1 U21162 ( .A1(n21266), .A2(n21265), .ZN(n21262) );
  AND2_X1 U21163 ( .A1(n21267), .A2(n21268), .ZN(n21265) );
  OR2_X1 U21164 ( .A1(n21269), .A2(n21270), .ZN(n21268) );
  INV_X1 U21165 ( .A(n21271), .ZN(n21270) );
  OR2_X1 U21166 ( .A1(n21271), .A2(n21272), .ZN(n21267) );
  INV_X1 U21167 ( .A(n21269), .ZN(n21272) );
  OR2_X1 U21168 ( .A1(n15106), .A2(n15139), .ZN(n20900) );
  OR2_X1 U21169 ( .A1(n21273), .A2(n21274), .ZN(n20897) );
  INV_X1 U21170 ( .A(n21275), .ZN(n21274) );
  OR2_X1 U21171 ( .A1(n21276), .A2(n21277), .ZN(n21275) );
  AND2_X1 U21172 ( .A1(n21277), .A2(n21276), .ZN(n21273) );
  AND2_X1 U21173 ( .A1(n21278), .A2(n21279), .ZN(n21276) );
  OR2_X1 U21174 ( .A1(n21280), .A2(n21281), .ZN(n21279) );
  INV_X1 U21175 ( .A(n21282), .ZN(n21281) );
  OR2_X1 U21176 ( .A1(n21282), .A2(n21283), .ZN(n21278) );
  INV_X1 U21177 ( .A(n21280), .ZN(n21283) );
  OR2_X1 U21178 ( .A1(n15140), .A2(n15139), .ZN(n15930) );
  OR2_X1 U21179 ( .A1(n21284), .A2(n21285), .ZN(n20908) );
  INV_X1 U21180 ( .A(n21286), .ZN(n21285) );
  OR2_X1 U21181 ( .A1(n21287), .A2(n21288), .ZN(n21286) );
  AND2_X1 U21182 ( .A1(n21288), .A2(n21287), .ZN(n21284) );
  AND2_X1 U21183 ( .A1(n21289), .A2(n21290), .ZN(n21287) );
  OR2_X1 U21184 ( .A1(n21291), .A2(n21292), .ZN(n21290) );
  INV_X1 U21185 ( .A(n21293), .ZN(n21292) );
  OR2_X1 U21186 ( .A1(n21293), .A2(n21294), .ZN(n21289) );
  INV_X1 U21187 ( .A(n21291), .ZN(n21294) );
  OR2_X1 U21188 ( .A1(n15174), .A2(n15139), .ZN(n20921) );
  OR2_X1 U21189 ( .A1(n21295), .A2(n21296), .ZN(n20918) );
  INV_X1 U21190 ( .A(n21297), .ZN(n21296) );
  OR2_X1 U21191 ( .A1(n21298), .A2(n21299), .ZN(n21297) );
  AND2_X1 U21192 ( .A1(n21299), .A2(n21298), .ZN(n21295) );
  AND2_X1 U21193 ( .A1(n21300), .A2(n21301), .ZN(n21298) );
  OR2_X1 U21194 ( .A1(n21302), .A2(n21303), .ZN(n21301) );
  INV_X1 U21195 ( .A(n21304), .ZN(n21303) );
  OR2_X1 U21196 ( .A1(n21304), .A2(n21305), .ZN(n21300) );
  INV_X1 U21197 ( .A(n21302), .ZN(n21305) );
  OR2_X1 U21198 ( .A1(n15208), .A2(n15139), .ZN(n20932) );
  OR2_X1 U21199 ( .A1(n21306), .A2(n21307), .ZN(n20929) );
  INV_X1 U21200 ( .A(n21308), .ZN(n21307) );
  OR2_X1 U21201 ( .A1(n21309), .A2(n21310), .ZN(n21308) );
  AND2_X1 U21202 ( .A1(n21310), .A2(n21309), .ZN(n21306) );
  AND2_X1 U21203 ( .A1(n21311), .A2(n21312), .ZN(n21309) );
  OR2_X1 U21204 ( .A1(n15927), .A2(n21313), .ZN(n21312) );
  INV_X1 U21205 ( .A(n21314), .ZN(n21313) );
  OR2_X1 U21206 ( .A1(n21314), .A2(n21315), .ZN(n21311) );
  INV_X1 U21207 ( .A(n15927), .ZN(n21315) );
  OR2_X1 U21208 ( .A1(n15242), .A2(n15139), .ZN(n20943) );
  OR2_X1 U21209 ( .A1(n21316), .A2(n21317), .ZN(n20940) );
  INV_X1 U21210 ( .A(n21318), .ZN(n21317) );
  OR2_X1 U21211 ( .A1(n21319), .A2(n21320), .ZN(n21318) );
  AND2_X1 U21212 ( .A1(n21320), .A2(n21319), .ZN(n21316) );
  AND2_X1 U21213 ( .A1(n21321), .A2(n21322), .ZN(n21319) );
  OR2_X1 U21214 ( .A1(n21323), .A2(n21324), .ZN(n21322) );
  INV_X1 U21215 ( .A(n21325), .ZN(n21324) );
  OR2_X1 U21216 ( .A1(n21325), .A2(n21326), .ZN(n21321) );
  INV_X1 U21217 ( .A(n21323), .ZN(n21326) );
  OR2_X1 U21218 ( .A1(n15287), .A2(n15139), .ZN(n20954) );
  OR2_X1 U21219 ( .A1(n21327), .A2(n21328), .ZN(n20951) );
  INV_X1 U21220 ( .A(n21329), .ZN(n21328) );
  OR2_X1 U21221 ( .A1(n21330), .A2(n21331), .ZN(n21329) );
  AND2_X1 U21222 ( .A1(n21331), .A2(n21330), .ZN(n21327) );
  AND2_X1 U21223 ( .A1(n21332), .A2(n21333), .ZN(n21330) );
  OR2_X1 U21224 ( .A1(n21334), .A2(n21335), .ZN(n21333) );
  INV_X1 U21225 ( .A(n21336), .ZN(n21335) );
  OR2_X1 U21226 ( .A1(n21336), .A2(n21337), .ZN(n21332) );
  INV_X1 U21227 ( .A(n21334), .ZN(n21337) );
  OR2_X1 U21228 ( .A1(n15321), .A2(n15139), .ZN(n20965) );
  OR2_X1 U21229 ( .A1(n21338), .A2(n21339), .ZN(n20962) );
  INV_X1 U21230 ( .A(n21340), .ZN(n21339) );
  OR2_X1 U21231 ( .A1(n21341), .A2(n21342), .ZN(n21340) );
  AND2_X1 U21232 ( .A1(n21342), .A2(n21341), .ZN(n21338) );
  AND2_X1 U21233 ( .A1(n21343), .A2(n21344), .ZN(n21341) );
  OR2_X1 U21234 ( .A1(n21345), .A2(n21346), .ZN(n21344) );
  INV_X1 U21235 ( .A(n21347), .ZN(n21346) );
  OR2_X1 U21236 ( .A1(n21347), .A2(n21348), .ZN(n21343) );
  INV_X1 U21237 ( .A(n21345), .ZN(n21348) );
  OR2_X1 U21238 ( .A1(n15355), .A2(n15139), .ZN(n20976) );
  OR2_X1 U21239 ( .A1(n21349), .A2(n21350), .ZN(n20973) );
  INV_X1 U21240 ( .A(n21351), .ZN(n21350) );
  OR2_X1 U21241 ( .A1(n21352), .A2(n21353), .ZN(n21351) );
  AND2_X1 U21242 ( .A1(n21353), .A2(n21352), .ZN(n21349) );
  AND2_X1 U21243 ( .A1(n21354), .A2(n21355), .ZN(n21352) );
  OR2_X1 U21244 ( .A1(n21356), .A2(n21357), .ZN(n21355) );
  INV_X1 U21245 ( .A(n21358), .ZN(n21357) );
  OR2_X1 U21246 ( .A1(n21358), .A2(n21359), .ZN(n21354) );
  INV_X1 U21247 ( .A(n21356), .ZN(n21359) );
  OR2_X1 U21248 ( .A1(n15389), .A2(n15139), .ZN(n20987) );
  OR2_X1 U21249 ( .A1(n21360), .A2(n21361), .ZN(n20984) );
  INV_X1 U21250 ( .A(n21362), .ZN(n21361) );
  OR2_X1 U21251 ( .A1(n21363), .A2(n21364), .ZN(n21362) );
  AND2_X1 U21252 ( .A1(n21364), .A2(n21363), .ZN(n21360) );
  AND2_X1 U21253 ( .A1(n21365), .A2(n21366), .ZN(n21363) );
  OR2_X1 U21254 ( .A1(n21367), .A2(n21368), .ZN(n21366) );
  INV_X1 U21255 ( .A(n21369), .ZN(n21368) );
  OR2_X1 U21256 ( .A1(n21369), .A2(n21370), .ZN(n21365) );
  INV_X1 U21257 ( .A(n21367), .ZN(n21370) );
  OR2_X1 U21258 ( .A1(n15423), .A2(n15139), .ZN(n20998) );
  OR2_X1 U21259 ( .A1(n21371), .A2(n21372), .ZN(n20995) );
  INV_X1 U21260 ( .A(n21373), .ZN(n21372) );
  OR2_X1 U21261 ( .A1(n21374), .A2(n21375), .ZN(n21373) );
  AND2_X1 U21262 ( .A1(n21375), .A2(n21374), .ZN(n21371) );
  AND2_X1 U21263 ( .A1(n21376), .A2(n21377), .ZN(n21374) );
  OR2_X1 U21264 ( .A1(n21378), .A2(n21379), .ZN(n21377) );
  INV_X1 U21265 ( .A(n21380), .ZN(n21379) );
  OR2_X1 U21266 ( .A1(n21380), .A2(n21381), .ZN(n21376) );
  INV_X1 U21267 ( .A(n21378), .ZN(n21381) );
  OR2_X1 U21268 ( .A1(n15457), .A2(n15139), .ZN(n21009) );
  OR2_X1 U21269 ( .A1(n21382), .A2(n21383), .ZN(n21006) );
  INV_X1 U21270 ( .A(n21384), .ZN(n21383) );
  OR2_X1 U21271 ( .A1(n21385), .A2(n21386), .ZN(n21384) );
  AND2_X1 U21272 ( .A1(n21386), .A2(n21385), .ZN(n21382) );
  AND2_X1 U21273 ( .A1(n21387), .A2(n21388), .ZN(n21385) );
  OR2_X1 U21274 ( .A1(n21389), .A2(n21390), .ZN(n21388) );
  INV_X1 U21275 ( .A(n21391), .ZN(n21390) );
  OR2_X1 U21276 ( .A1(n21391), .A2(n21392), .ZN(n21387) );
  INV_X1 U21277 ( .A(n21389), .ZN(n21392) );
  OR2_X1 U21278 ( .A1(n15491), .A2(n15139), .ZN(n21020) );
  OR2_X1 U21279 ( .A1(n21393), .A2(n21394), .ZN(n21017) );
  INV_X1 U21280 ( .A(n21395), .ZN(n21394) );
  OR2_X1 U21281 ( .A1(n21396), .A2(n21397), .ZN(n21395) );
  AND2_X1 U21282 ( .A1(n21397), .A2(n21396), .ZN(n21393) );
  AND2_X1 U21283 ( .A1(n21398), .A2(n21399), .ZN(n21396) );
  OR2_X1 U21284 ( .A1(n21400), .A2(n21401), .ZN(n21399) );
  INV_X1 U21285 ( .A(n21402), .ZN(n21401) );
  OR2_X1 U21286 ( .A1(n21402), .A2(n21403), .ZN(n21398) );
  INV_X1 U21287 ( .A(n21400), .ZN(n21403) );
  OR2_X1 U21288 ( .A1(n15525), .A2(n15139), .ZN(n21031) );
  OR2_X1 U21289 ( .A1(n21404), .A2(n21405), .ZN(n21028) );
  INV_X1 U21290 ( .A(n21406), .ZN(n21405) );
  OR2_X1 U21291 ( .A1(n21407), .A2(n21408), .ZN(n21406) );
  AND2_X1 U21292 ( .A1(n21408), .A2(n21407), .ZN(n21404) );
  AND2_X1 U21293 ( .A1(n21409), .A2(n21410), .ZN(n21407) );
  OR2_X1 U21294 ( .A1(n21411), .A2(n21412), .ZN(n21410) );
  INV_X1 U21295 ( .A(n21413), .ZN(n21412) );
  OR2_X1 U21296 ( .A1(n21413), .A2(n21414), .ZN(n21409) );
  INV_X1 U21297 ( .A(n21411), .ZN(n21414) );
  OR2_X1 U21298 ( .A1(n15559), .A2(n15139), .ZN(n21042) );
  OR2_X1 U21299 ( .A1(n21415), .A2(n21416), .ZN(n21039) );
  INV_X1 U21300 ( .A(n21417), .ZN(n21416) );
  OR2_X1 U21301 ( .A1(n21418), .A2(n21419), .ZN(n21417) );
  AND2_X1 U21302 ( .A1(n21419), .A2(n21418), .ZN(n21415) );
  AND2_X1 U21303 ( .A1(n21420), .A2(n21421), .ZN(n21418) );
  OR2_X1 U21304 ( .A1(n21422), .A2(n21423), .ZN(n21421) );
  INV_X1 U21305 ( .A(n21424), .ZN(n21423) );
  OR2_X1 U21306 ( .A1(n21424), .A2(n21425), .ZN(n21420) );
  INV_X1 U21307 ( .A(n21422), .ZN(n21425) );
  OR2_X1 U21308 ( .A1(n15593), .A2(n15139), .ZN(n21056) );
  OR2_X1 U21309 ( .A1(n21426), .A2(n21427), .ZN(n21050) );
  INV_X1 U21310 ( .A(n21428), .ZN(n21427) );
  OR2_X1 U21311 ( .A1(n21429), .A2(n21430), .ZN(n21428) );
  AND2_X1 U21312 ( .A1(n21430), .A2(n21429), .ZN(n21426) );
  AND2_X1 U21313 ( .A1(n21431), .A2(n21432), .ZN(n21429) );
  INV_X1 U21314 ( .A(n21433), .ZN(n21432) );
  AND2_X1 U21315 ( .A1(n21434), .A2(n21435), .ZN(n21433) );
  OR2_X1 U21316 ( .A1(n21435), .A2(n21434), .ZN(n21431) );
  INV_X1 U21317 ( .A(n21436), .ZN(n21434) );
  OR2_X1 U21318 ( .A1(n15638), .A2(n15139), .ZN(n21066) );
  AND2_X1 U21319 ( .A1(n21437), .A2(n21438), .ZN(n21061) );
  INV_X1 U21320 ( .A(n21439), .ZN(n21438) );
  AND2_X1 U21321 ( .A1(n21440), .A2(n21441), .ZN(n21439) );
  OR2_X1 U21322 ( .A1(n21441), .A2(n21440), .ZN(n21437) );
  OR2_X1 U21323 ( .A1(n21442), .A2(n21443), .ZN(n21440) );
  AND2_X1 U21324 ( .A1(n21444), .A2(n21445), .ZN(n21443) );
  INV_X1 U21325 ( .A(n21446), .ZN(n21444) );
  AND2_X1 U21326 ( .A1(n21447), .A2(n21446), .ZN(n21442) );
  INV_X1 U21327 ( .A(n21445), .ZN(n21447) );
  OR2_X1 U21328 ( .A1(n15672), .A2(n15139), .ZN(n21077) );
  AND2_X1 U21329 ( .A1(n21448), .A2(n21449), .ZN(n21072) );
  INV_X1 U21330 ( .A(n21450), .ZN(n21449) );
  AND2_X1 U21331 ( .A1(n21451), .A2(n21452), .ZN(n21450) );
  OR2_X1 U21332 ( .A1(n21452), .A2(n21451), .ZN(n21448) );
  OR2_X1 U21333 ( .A1(n21453), .A2(n21454), .ZN(n21451) );
  AND2_X1 U21334 ( .A1(n21455), .A2(n21456), .ZN(n21454) );
  INV_X1 U21335 ( .A(n21457), .ZN(n21455) );
  AND2_X1 U21336 ( .A1(n21458), .A2(n21457), .ZN(n21453) );
  INV_X1 U21337 ( .A(n21456), .ZN(n21458) );
  OR2_X1 U21338 ( .A1(n15706), .A2(n15139), .ZN(n21088) );
  AND2_X1 U21339 ( .A1(n21459), .A2(n21460), .ZN(n21083) );
  INV_X1 U21340 ( .A(n21461), .ZN(n21460) );
  AND2_X1 U21341 ( .A1(n21462), .A2(n21463), .ZN(n21461) );
  OR2_X1 U21342 ( .A1(n21463), .A2(n21462), .ZN(n21459) );
  OR2_X1 U21343 ( .A1(n21464), .A2(n21465), .ZN(n21462) );
  AND2_X1 U21344 ( .A1(n21466), .A2(n21467), .ZN(n21465) );
  INV_X1 U21345 ( .A(n21468), .ZN(n21466) );
  AND2_X1 U21346 ( .A1(n21469), .A2(n21468), .ZN(n21464) );
  INV_X1 U21347 ( .A(n21467), .ZN(n21469) );
  OR2_X1 U21348 ( .A1(n15740), .A2(n15139), .ZN(n21099) );
  AND2_X1 U21349 ( .A1(n21470), .A2(n21471), .ZN(n21094) );
  INV_X1 U21350 ( .A(n21472), .ZN(n21471) );
  AND2_X1 U21351 ( .A1(n21473), .A2(n21474), .ZN(n21472) );
  OR2_X1 U21352 ( .A1(n21474), .A2(n21473), .ZN(n21470) );
  OR2_X1 U21353 ( .A1(n21475), .A2(n21476), .ZN(n21473) );
  AND2_X1 U21354 ( .A1(n21477), .A2(n21478), .ZN(n21476) );
  INV_X1 U21355 ( .A(n21479), .ZN(n21477) );
  AND2_X1 U21356 ( .A1(n21480), .A2(n21479), .ZN(n21475) );
  INV_X1 U21357 ( .A(n21478), .ZN(n21480) );
  OR2_X1 U21358 ( .A1(n15774), .A2(n15139), .ZN(n21110) );
  INV_X1 U21359 ( .A(b_21_), .ZN(n15139) );
  AND2_X1 U21360 ( .A1(n21481), .A2(n21482), .ZN(n21105) );
  INV_X1 U21361 ( .A(n21483), .ZN(n21482) );
  AND2_X1 U21362 ( .A1(n21484), .A2(n21485), .ZN(n21483) );
  OR2_X1 U21363 ( .A1(n21485), .A2(n21484), .ZN(n21481) );
  OR2_X1 U21364 ( .A1(n21486), .A2(n21487), .ZN(n21484) );
  AND2_X1 U21365 ( .A1(n21488), .A2(n21489), .ZN(n21487) );
  INV_X1 U21366 ( .A(n21490), .ZN(n21488) );
  AND2_X1 U21367 ( .A1(n21491), .A2(n21490), .ZN(n21486) );
  INV_X1 U21368 ( .A(n21489), .ZN(n21491) );
  AND2_X1 U21369 ( .A1(n21492), .A2(n21493), .ZN(n20288) );
  INV_X1 U21370 ( .A(n21494), .ZN(n21493) );
  AND2_X1 U21371 ( .A1(n21495), .A2(n20302), .ZN(n21494) );
  OR2_X1 U21372 ( .A1(n20302), .A2(n21495), .ZN(n21492) );
  OR2_X1 U21373 ( .A1(n21496), .A2(n21497), .ZN(n21495) );
  AND2_X1 U21374 ( .A1(n21498), .A2(n20301), .ZN(n21497) );
  INV_X1 U21375 ( .A(n20300), .ZN(n21498) );
  AND2_X1 U21376 ( .A1(n21499), .A2(n20300), .ZN(n21496) );
  OR2_X1 U21377 ( .A1(n15774), .A2(n15173), .ZN(n20300) );
  INV_X1 U21378 ( .A(n20301), .ZN(n21499) );
  OR2_X1 U21379 ( .A1(n21500), .A2(n21501), .ZN(n20301) );
  AND2_X1 U21380 ( .A1(n21490), .A2(n21489), .ZN(n21501) );
  AND2_X1 U21381 ( .A1(n21485), .A2(n21502), .ZN(n21500) );
  OR2_X1 U21382 ( .A1(n21490), .A2(n21489), .ZN(n21502) );
  OR2_X1 U21383 ( .A1(n21503), .A2(n21504), .ZN(n21489) );
  AND2_X1 U21384 ( .A1(n21479), .A2(n21478), .ZN(n21504) );
  AND2_X1 U21385 ( .A1(n21474), .A2(n21505), .ZN(n21503) );
  OR2_X1 U21386 ( .A1(n21479), .A2(n21478), .ZN(n21505) );
  OR2_X1 U21387 ( .A1(n21506), .A2(n21507), .ZN(n21478) );
  AND2_X1 U21388 ( .A1(n21468), .A2(n21467), .ZN(n21507) );
  AND2_X1 U21389 ( .A1(n21463), .A2(n21508), .ZN(n21506) );
  OR2_X1 U21390 ( .A1(n21468), .A2(n21467), .ZN(n21508) );
  OR2_X1 U21391 ( .A1(n21509), .A2(n21510), .ZN(n21467) );
  AND2_X1 U21392 ( .A1(n21457), .A2(n21456), .ZN(n21510) );
  AND2_X1 U21393 ( .A1(n21452), .A2(n21511), .ZN(n21509) );
  OR2_X1 U21394 ( .A1(n21457), .A2(n21456), .ZN(n21511) );
  OR2_X1 U21395 ( .A1(n21512), .A2(n21513), .ZN(n21456) );
  AND2_X1 U21396 ( .A1(n21446), .A2(n21445), .ZN(n21513) );
  AND2_X1 U21397 ( .A1(n21441), .A2(n21514), .ZN(n21512) );
  OR2_X1 U21398 ( .A1(n21446), .A2(n21445), .ZN(n21514) );
  OR2_X1 U21399 ( .A1(n21515), .A2(n21516), .ZN(n21445) );
  AND2_X1 U21400 ( .A1(n21436), .A2(n21435), .ZN(n21516) );
  AND2_X1 U21401 ( .A1(n21430), .A2(n21517), .ZN(n21515) );
  OR2_X1 U21402 ( .A1(n21436), .A2(n21435), .ZN(n21517) );
  OR2_X1 U21403 ( .A1(n21518), .A2(n21519), .ZN(n21435) );
  AND2_X1 U21404 ( .A1(n21422), .A2(n21424), .ZN(n21519) );
  AND2_X1 U21405 ( .A1(n21419), .A2(n21520), .ZN(n21518) );
  OR2_X1 U21406 ( .A1(n21422), .A2(n21424), .ZN(n21520) );
  OR2_X1 U21407 ( .A1(n21521), .A2(n21522), .ZN(n21424) );
  AND2_X1 U21408 ( .A1(n21411), .A2(n21413), .ZN(n21522) );
  AND2_X1 U21409 ( .A1(n21408), .A2(n21523), .ZN(n21521) );
  OR2_X1 U21410 ( .A1(n21411), .A2(n21413), .ZN(n21523) );
  OR2_X1 U21411 ( .A1(n21524), .A2(n21525), .ZN(n21413) );
  AND2_X1 U21412 ( .A1(n21400), .A2(n21402), .ZN(n21525) );
  AND2_X1 U21413 ( .A1(n21397), .A2(n21526), .ZN(n21524) );
  OR2_X1 U21414 ( .A1(n21400), .A2(n21402), .ZN(n21526) );
  OR2_X1 U21415 ( .A1(n21527), .A2(n21528), .ZN(n21402) );
  AND2_X1 U21416 ( .A1(n21389), .A2(n21391), .ZN(n21528) );
  AND2_X1 U21417 ( .A1(n21386), .A2(n21529), .ZN(n21527) );
  OR2_X1 U21418 ( .A1(n21389), .A2(n21391), .ZN(n21529) );
  OR2_X1 U21419 ( .A1(n21530), .A2(n21531), .ZN(n21391) );
  AND2_X1 U21420 ( .A1(n21378), .A2(n21380), .ZN(n21531) );
  AND2_X1 U21421 ( .A1(n21375), .A2(n21532), .ZN(n21530) );
  OR2_X1 U21422 ( .A1(n21378), .A2(n21380), .ZN(n21532) );
  OR2_X1 U21423 ( .A1(n21533), .A2(n21534), .ZN(n21380) );
  AND2_X1 U21424 ( .A1(n21367), .A2(n21369), .ZN(n21534) );
  AND2_X1 U21425 ( .A1(n21364), .A2(n21535), .ZN(n21533) );
  OR2_X1 U21426 ( .A1(n21367), .A2(n21369), .ZN(n21535) );
  OR2_X1 U21427 ( .A1(n21536), .A2(n21537), .ZN(n21369) );
  AND2_X1 U21428 ( .A1(n21356), .A2(n21358), .ZN(n21537) );
  AND2_X1 U21429 ( .A1(n21353), .A2(n21538), .ZN(n21536) );
  OR2_X1 U21430 ( .A1(n21356), .A2(n21358), .ZN(n21538) );
  OR2_X1 U21431 ( .A1(n21539), .A2(n21540), .ZN(n21358) );
  AND2_X1 U21432 ( .A1(n21345), .A2(n21347), .ZN(n21540) );
  AND2_X1 U21433 ( .A1(n21342), .A2(n21541), .ZN(n21539) );
  OR2_X1 U21434 ( .A1(n21345), .A2(n21347), .ZN(n21541) );
  OR2_X1 U21435 ( .A1(n21542), .A2(n21543), .ZN(n21347) );
  AND2_X1 U21436 ( .A1(n21334), .A2(n21336), .ZN(n21543) );
  AND2_X1 U21437 ( .A1(n21331), .A2(n21544), .ZN(n21542) );
  OR2_X1 U21438 ( .A1(n21334), .A2(n21336), .ZN(n21544) );
  OR2_X1 U21439 ( .A1(n21545), .A2(n21546), .ZN(n21336) );
  AND2_X1 U21440 ( .A1(n21323), .A2(n21325), .ZN(n21546) );
  AND2_X1 U21441 ( .A1(n21320), .A2(n21547), .ZN(n21545) );
  OR2_X1 U21442 ( .A1(n21323), .A2(n21325), .ZN(n21547) );
  OR2_X1 U21443 ( .A1(n21548), .A2(n21549), .ZN(n21325) );
  AND2_X1 U21444 ( .A1(n15927), .A2(n21314), .ZN(n21549) );
  AND2_X1 U21445 ( .A1(n21310), .A2(n21550), .ZN(n21548) );
  OR2_X1 U21446 ( .A1(n15927), .A2(n21314), .ZN(n21550) );
  OR2_X1 U21447 ( .A1(n21551), .A2(n21552), .ZN(n21314) );
  AND2_X1 U21448 ( .A1(n21302), .A2(n21304), .ZN(n21552) );
  AND2_X1 U21449 ( .A1(n21299), .A2(n21553), .ZN(n21551) );
  OR2_X1 U21450 ( .A1(n21302), .A2(n21304), .ZN(n21553) );
  OR2_X1 U21451 ( .A1(n21554), .A2(n21555), .ZN(n21304) );
  AND2_X1 U21452 ( .A1(n21291), .A2(n21293), .ZN(n21555) );
  AND2_X1 U21453 ( .A1(n21288), .A2(n21556), .ZN(n21554) );
  OR2_X1 U21454 ( .A1(n21291), .A2(n21293), .ZN(n21556) );
  OR2_X1 U21455 ( .A1(n21557), .A2(n21558), .ZN(n21293) );
  AND2_X1 U21456 ( .A1(n21280), .A2(n21282), .ZN(n21558) );
  AND2_X1 U21457 ( .A1(n21277), .A2(n21559), .ZN(n21557) );
  OR2_X1 U21458 ( .A1(n21280), .A2(n21282), .ZN(n21559) );
  OR2_X1 U21459 ( .A1(n21560), .A2(n21561), .ZN(n21282) );
  AND2_X1 U21460 ( .A1(n21269), .A2(n21271), .ZN(n21561) );
  AND2_X1 U21461 ( .A1(n21266), .A2(n21562), .ZN(n21560) );
  OR2_X1 U21462 ( .A1(n21269), .A2(n21271), .ZN(n21562) );
  OR2_X1 U21463 ( .A1(n21563), .A2(n21564), .ZN(n21271) );
  AND2_X1 U21464 ( .A1(n21258), .A2(n21260), .ZN(n21564) );
  AND2_X1 U21465 ( .A1(n21255), .A2(n21565), .ZN(n21563) );
  OR2_X1 U21466 ( .A1(n21258), .A2(n21260), .ZN(n21565) );
  OR2_X1 U21467 ( .A1(n21566), .A2(n21567), .ZN(n21260) );
  AND2_X1 U21468 ( .A1(n21247), .A2(n21249), .ZN(n21567) );
  AND2_X1 U21469 ( .A1(n21244), .A2(n21568), .ZN(n21566) );
  OR2_X1 U21470 ( .A1(n21247), .A2(n21249), .ZN(n21568) );
  OR2_X1 U21471 ( .A1(n21569), .A2(n21570), .ZN(n21249) );
  AND2_X1 U21472 ( .A1(n21236), .A2(n21238), .ZN(n21570) );
  AND2_X1 U21473 ( .A1(n21233), .A2(n21571), .ZN(n21569) );
  OR2_X1 U21474 ( .A1(n21236), .A2(n21238), .ZN(n21571) );
  OR2_X1 U21475 ( .A1(n21572), .A2(n21573), .ZN(n21238) );
  AND2_X1 U21476 ( .A1(n21225), .A2(n21227), .ZN(n21573) );
  AND2_X1 U21477 ( .A1(n21222), .A2(n21574), .ZN(n21572) );
  OR2_X1 U21478 ( .A1(n21225), .A2(n21227), .ZN(n21574) );
  OR2_X1 U21479 ( .A1(n21575), .A2(n21576), .ZN(n21227) );
  AND2_X1 U21480 ( .A1(n21210), .A2(n21215), .ZN(n21576) );
  AND2_X1 U21481 ( .A1(n21214), .A2(n21577), .ZN(n21575) );
  OR2_X1 U21482 ( .A1(n21210), .A2(n21215), .ZN(n21577) );
  INV_X1 U21483 ( .A(n21216), .ZN(n21215) );
  AND3_X1 U21484 ( .A1(b_20_), .A2(b_19_), .A3(n15957), .ZN(n21216) );
  OR2_X1 U21485 ( .A1(n14857), .A2(n15173), .ZN(n21210) );
  INV_X1 U21486 ( .A(n21217), .ZN(n21214) );
  OR2_X1 U21487 ( .A1(n21578), .A2(n21579), .ZN(n21217) );
  AND2_X1 U21488 ( .A1(b_19_), .A2(n21580), .ZN(n21579) );
  OR2_X1 U21489 ( .A1(n21581), .A2(n16981), .ZN(n21580) );
  AND2_X1 U21490 ( .A1(a_30_), .A2(n15241), .ZN(n21581) );
  AND2_X1 U21491 ( .A1(b_18_), .A2(n21582), .ZN(n21578) );
  OR2_X1 U21492 ( .A1(n21583), .A2(n14817), .ZN(n21582) );
  AND2_X1 U21493 ( .A1(a_31_), .A2(n15207), .ZN(n21583) );
  OR2_X1 U21494 ( .A1(n14891), .A2(n15173), .ZN(n21225) );
  OR2_X1 U21495 ( .A1(n21584), .A2(n21585), .ZN(n21222) );
  AND2_X1 U21496 ( .A1(n21586), .A2(n21587), .ZN(n21585) );
  INV_X1 U21497 ( .A(n21588), .ZN(n21584) );
  OR2_X1 U21498 ( .A1(n21586), .A2(n21587), .ZN(n21588) );
  OR2_X1 U21499 ( .A1(n21589), .A2(n21590), .ZN(n21586) );
  AND2_X1 U21500 ( .A1(n21591), .A2(n21592), .ZN(n21590) );
  AND2_X1 U21501 ( .A1(n21593), .A2(n21594), .ZN(n21589) );
  OR2_X1 U21502 ( .A1(n14936), .A2(n15173), .ZN(n21236) );
  OR2_X1 U21503 ( .A1(n21595), .A2(n21596), .ZN(n21233) );
  INV_X1 U21504 ( .A(n21597), .ZN(n21596) );
  OR2_X1 U21505 ( .A1(n21598), .A2(n21599), .ZN(n21597) );
  AND2_X1 U21506 ( .A1(n21599), .A2(n21598), .ZN(n21595) );
  AND2_X1 U21507 ( .A1(n21600), .A2(n21601), .ZN(n21598) );
  OR2_X1 U21508 ( .A1(n21602), .A2(n21603), .ZN(n21601) );
  INV_X1 U21509 ( .A(n21604), .ZN(n21603) );
  OR2_X1 U21510 ( .A1(n21604), .A2(n21605), .ZN(n21600) );
  INV_X1 U21511 ( .A(n21602), .ZN(n21605) );
  OR2_X1 U21512 ( .A1(n14970), .A2(n15173), .ZN(n21247) );
  OR2_X1 U21513 ( .A1(n21606), .A2(n21607), .ZN(n21244) );
  INV_X1 U21514 ( .A(n21608), .ZN(n21607) );
  OR2_X1 U21515 ( .A1(n21609), .A2(n21610), .ZN(n21608) );
  AND2_X1 U21516 ( .A1(n21610), .A2(n21609), .ZN(n21606) );
  AND2_X1 U21517 ( .A1(n21611), .A2(n21612), .ZN(n21609) );
  OR2_X1 U21518 ( .A1(n21613), .A2(n21614), .ZN(n21612) );
  INV_X1 U21519 ( .A(n21615), .ZN(n21614) );
  OR2_X1 U21520 ( .A1(n21615), .A2(n21616), .ZN(n21611) );
  INV_X1 U21521 ( .A(n21613), .ZN(n21616) );
  OR2_X1 U21522 ( .A1(n15004), .A2(n15173), .ZN(n21258) );
  OR2_X1 U21523 ( .A1(n21617), .A2(n21618), .ZN(n21255) );
  INV_X1 U21524 ( .A(n21619), .ZN(n21618) );
  OR2_X1 U21525 ( .A1(n21620), .A2(n21621), .ZN(n21619) );
  AND2_X1 U21526 ( .A1(n21621), .A2(n21620), .ZN(n21617) );
  AND2_X1 U21527 ( .A1(n21622), .A2(n21623), .ZN(n21620) );
  OR2_X1 U21528 ( .A1(n21624), .A2(n21625), .ZN(n21623) );
  INV_X1 U21529 ( .A(n21626), .ZN(n21625) );
  OR2_X1 U21530 ( .A1(n21626), .A2(n21627), .ZN(n21622) );
  INV_X1 U21531 ( .A(n21624), .ZN(n21627) );
  OR2_X1 U21532 ( .A1(n15038), .A2(n15173), .ZN(n21269) );
  OR2_X1 U21533 ( .A1(n21628), .A2(n21629), .ZN(n21266) );
  INV_X1 U21534 ( .A(n21630), .ZN(n21629) );
  OR2_X1 U21535 ( .A1(n21631), .A2(n21632), .ZN(n21630) );
  AND2_X1 U21536 ( .A1(n21632), .A2(n21631), .ZN(n21628) );
  AND2_X1 U21537 ( .A1(n21633), .A2(n21634), .ZN(n21631) );
  OR2_X1 U21538 ( .A1(n21635), .A2(n21636), .ZN(n21634) );
  INV_X1 U21539 ( .A(n21637), .ZN(n21636) );
  OR2_X1 U21540 ( .A1(n21637), .A2(n21638), .ZN(n21633) );
  INV_X1 U21541 ( .A(n21635), .ZN(n21638) );
  OR2_X1 U21542 ( .A1(n15072), .A2(n15173), .ZN(n21280) );
  OR2_X1 U21543 ( .A1(n21639), .A2(n21640), .ZN(n21277) );
  INV_X1 U21544 ( .A(n21641), .ZN(n21640) );
  OR2_X1 U21545 ( .A1(n21642), .A2(n21643), .ZN(n21641) );
  AND2_X1 U21546 ( .A1(n21643), .A2(n21642), .ZN(n21639) );
  AND2_X1 U21547 ( .A1(n21644), .A2(n21645), .ZN(n21642) );
  OR2_X1 U21548 ( .A1(n21646), .A2(n21647), .ZN(n21645) );
  INV_X1 U21549 ( .A(n21648), .ZN(n21647) );
  OR2_X1 U21550 ( .A1(n21648), .A2(n21649), .ZN(n21644) );
  INV_X1 U21551 ( .A(n21646), .ZN(n21649) );
  OR2_X1 U21552 ( .A1(n15106), .A2(n15173), .ZN(n21291) );
  OR2_X1 U21553 ( .A1(n21650), .A2(n21651), .ZN(n21288) );
  INV_X1 U21554 ( .A(n21652), .ZN(n21651) );
  OR2_X1 U21555 ( .A1(n21653), .A2(n21654), .ZN(n21652) );
  AND2_X1 U21556 ( .A1(n21654), .A2(n21653), .ZN(n21650) );
  AND2_X1 U21557 ( .A1(n21655), .A2(n21656), .ZN(n21653) );
  OR2_X1 U21558 ( .A1(n21657), .A2(n21658), .ZN(n21656) );
  INV_X1 U21559 ( .A(n21659), .ZN(n21658) );
  OR2_X1 U21560 ( .A1(n21659), .A2(n21660), .ZN(n21655) );
  INV_X1 U21561 ( .A(n21657), .ZN(n21660) );
  OR2_X1 U21562 ( .A1(n15140), .A2(n15173), .ZN(n21302) );
  OR2_X1 U21563 ( .A1(n21661), .A2(n21662), .ZN(n21299) );
  INV_X1 U21564 ( .A(n21663), .ZN(n21662) );
  OR2_X1 U21565 ( .A1(n21664), .A2(n21665), .ZN(n21663) );
  AND2_X1 U21566 ( .A1(n21665), .A2(n21664), .ZN(n21661) );
  AND2_X1 U21567 ( .A1(n21666), .A2(n21667), .ZN(n21664) );
  OR2_X1 U21568 ( .A1(n21668), .A2(n21669), .ZN(n21667) );
  INV_X1 U21569 ( .A(n21670), .ZN(n21669) );
  OR2_X1 U21570 ( .A1(n21670), .A2(n21671), .ZN(n21666) );
  INV_X1 U21571 ( .A(n21668), .ZN(n21671) );
  OR2_X1 U21572 ( .A1(n15174), .A2(n15173), .ZN(n15927) );
  OR2_X1 U21573 ( .A1(n21672), .A2(n21673), .ZN(n21310) );
  INV_X1 U21574 ( .A(n21674), .ZN(n21673) );
  OR2_X1 U21575 ( .A1(n21675), .A2(n21676), .ZN(n21674) );
  AND2_X1 U21576 ( .A1(n21676), .A2(n21675), .ZN(n21672) );
  AND2_X1 U21577 ( .A1(n21677), .A2(n21678), .ZN(n21675) );
  OR2_X1 U21578 ( .A1(n21679), .A2(n21680), .ZN(n21678) );
  INV_X1 U21579 ( .A(n21681), .ZN(n21680) );
  OR2_X1 U21580 ( .A1(n21681), .A2(n21682), .ZN(n21677) );
  INV_X1 U21581 ( .A(n21679), .ZN(n21682) );
  OR2_X1 U21582 ( .A1(n15208), .A2(n15173), .ZN(n21323) );
  OR2_X1 U21583 ( .A1(n21683), .A2(n21684), .ZN(n21320) );
  INV_X1 U21584 ( .A(n21685), .ZN(n21684) );
  OR2_X1 U21585 ( .A1(n21686), .A2(n21687), .ZN(n21685) );
  AND2_X1 U21586 ( .A1(n21687), .A2(n21686), .ZN(n21683) );
  AND2_X1 U21587 ( .A1(n21688), .A2(n21689), .ZN(n21686) );
  OR2_X1 U21588 ( .A1(n21690), .A2(n21691), .ZN(n21689) );
  INV_X1 U21589 ( .A(n21692), .ZN(n21691) );
  OR2_X1 U21590 ( .A1(n21692), .A2(n21693), .ZN(n21688) );
  INV_X1 U21591 ( .A(n21690), .ZN(n21693) );
  OR2_X1 U21592 ( .A1(n15242), .A2(n15173), .ZN(n21334) );
  OR2_X1 U21593 ( .A1(n21694), .A2(n21695), .ZN(n21331) );
  INV_X1 U21594 ( .A(n21696), .ZN(n21695) );
  OR2_X1 U21595 ( .A1(n21697), .A2(n21698), .ZN(n21696) );
  AND2_X1 U21596 ( .A1(n21698), .A2(n21697), .ZN(n21694) );
  AND2_X1 U21597 ( .A1(n21699), .A2(n21700), .ZN(n21697) );
  OR2_X1 U21598 ( .A1(n15924), .A2(n21701), .ZN(n21700) );
  INV_X1 U21599 ( .A(n21702), .ZN(n21701) );
  OR2_X1 U21600 ( .A1(n21702), .A2(n21703), .ZN(n21699) );
  INV_X1 U21601 ( .A(n15924), .ZN(n21703) );
  OR2_X1 U21602 ( .A1(n15287), .A2(n15173), .ZN(n21345) );
  OR2_X1 U21603 ( .A1(n21704), .A2(n21705), .ZN(n21342) );
  INV_X1 U21604 ( .A(n21706), .ZN(n21705) );
  OR2_X1 U21605 ( .A1(n21707), .A2(n21708), .ZN(n21706) );
  AND2_X1 U21606 ( .A1(n21708), .A2(n21707), .ZN(n21704) );
  AND2_X1 U21607 ( .A1(n21709), .A2(n21710), .ZN(n21707) );
  OR2_X1 U21608 ( .A1(n21711), .A2(n21712), .ZN(n21710) );
  INV_X1 U21609 ( .A(n21713), .ZN(n21712) );
  OR2_X1 U21610 ( .A1(n21713), .A2(n21714), .ZN(n21709) );
  INV_X1 U21611 ( .A(n21711), .ZN(n21714) );
  OR2_X1 U21612 ( .A1(n15321), .A2(n15173), .ZN(n21356) );
  OR2_X1 U21613 ( .A1(n21715), .A2(n21716), .ZN(n21353) );
  INV_X1 U21614 ( .A(n21717), .ZN(n21716) );
  OR2_X1 U21615 ( .A1(n21718), .A2(n21719), .ZN(n21717) );
  AND2_X1 U21616 ( .A1(n21719), .A2(n21718), .ZN(n21715) );
  AND2_X1 U21617 ( .A1(n21720), .A2(n21721), .ZN(n21718) );
  OR2_X1 U21618 ( .A1(n21722), .A2(n21723), .ZN(n21721) );
  INV_X1 U21619 ( .A(n21724), .ZN(n21723) );
  OR2_X1 U21620 ( .A1(n21724), .A2(n21725), .ZN(n21720) );
  INV_X1 U21621 ( .A(n21722), .ZN(n21725) );
  OR2_X1 U21622 ( .A1(n15355), .A2(n15173), .ZN(n21367) );
  OR2_X1 U21623 ( .A1(n21726), .A2(n21727), .ZN(n21364) );
  INV_X1 U21624 ( .A(n21728), .ZN(n21727) );
  OR2_X1 U21625 ( .A1(n21729), .A2(n21730), .ZN(n21728) );
  AND2_X1 U21626 ( .A1(n21730), .A2(n21729), .ZN(n21726) );
  AND2_X1 U21627 ( .A1(n21731), .A2(n21732), .ZN(n21729) );
  OR2_X1 U21628 ( .A1(n21733), .A2(n21734), .ZN(n21732) );
  INV_X1 U21629 ( .A(n21735), .ZN(n21734) );
  OR2_X1 U21630 ( .A1(n21735), .A2(n21736), .ZN(n21731) );
  INV_X1 U21631 ( .A(n21733), .ZN(n21736) );
  OR2_X1 U21632 ( .A1(n15389), .A2(n15173), .ZN(n21378) );
  OR2_X1 U21633 ( .A1(n21737), .A2(n21738), .ZN(n21375) );
  INV_X1 U21634 ( .A(n21739), .ZN(n21738) );
  OR2_X1 U21635 ( .A1(n21740), .A2(n21741), .ZN(n21739) );
  AND2_X1 U21636 ( .A1(n21741), .A2(n21740), .ZN(n21737) );
  AND2_X1 U21637 ( .A1(n21742), .A2(n21743), .ZN(n21740) );
  OR2_X1 U21638 ( .A1(n21744), .A2(n21745), .ZN(n21743) );
  INV_X1 U21639 ( .A(n21746), .ZN(n21745) );
  OR2_X1 U21640 ( .A1(n21746), .A2(n21747), .ZN(n21742) );
  INV_X1 U21641 ( .A(n21744), .ZN(n21747) );
  OR2_X1 U21642 ( .A1(n15423), .A2(n15173), .ZN(n21389) );
  OR2_X1 U21643 ( .A1(n21748), .A2(n21749), .ZN(n21386) );
  INV_X1 U21644 ( .A(n21750), .ZN(n21749) );
  OR2_X1 U21645 ( .A1(n21751), .A2(n21752), .ZN(n21750) );
  AND2_X1 U21646 ( .A1(n21752), .A2(n21751), .ZN(n21748) );
  AND2_X1 U21647 ( .A1(n21753), .A2(n21754), .ZN(n21751) );
  OR2_X1 U21648 ( .A1(n21755), .A2(n21756), .ZN(n21754) );
  INV_X1 U21649 ( .A(n21757), .ZN(n21756) );
  OR2_X1 U21650 ( .A1(n21757), .A2(n21758), .ZN(n21753) );
  INV_X1 U21651 ( .A(n21755), .ZN(n21758) );
  OR2_X1 U21652 ( .A1(n15457), .A2(n15173), .ZN(n21400) );
  OR2_X1 U21653 ( .A1(n21759), .A2(n21760), .ZN(n21397) );
  INV_X1 U21654 ( .A(n21761), .ZN(n21760) );
  OR2_X1 U21655 ( .A1(n21762), .A2(n21763), .ZN(n21761) );
  AND2_X1 U21656 ( .A1(n21763), .A2(n21762), .ZN(n21759) );
  AND2_X1 U21657 ( .A1(n21764), .A2(n21765), .ZN(n21762) );
  OR2_X1 U21658 ( .A1(n21766), .A2(n21767), .ZN(n21765) );
  INV_X1 U21659 ( .A(n21768), .ZN(n21767) );
  OR2_X1 U21660 ( .A1(n21768), .A2(n21769), .ZN(n21764) );
  INV_X1 U21661 ( .A(n21766), .ZN(n21769) );
  OR2_X1 U21662 ( .A1(n15491), .A2(n15173), .ZN(n21411) );
  OR2_X1 U21663 ( .A1(n21770), .A2(n21771), .ZN(n21408) );
  INV_X1 U21664 ( .A(n21772), .ZN(n21771) );
  OR2_X1 U21665 ( .A1(n21773), .A2(n21774), .ZN(n21772) );
  AND2_X1 U21666 ( .A1(n21774), .A2(n21773), .ZN(n21770) );
  AND2_X1 U21667 ( .A1(n21775), .A2(n21776), .ZN(n21773) );
  OR2_X1 U21668 ( .A1(n21777), .A2(n21778), .ZN(n21776) );
  INV_X1 U21669 ( .A(n21779), .ZN(n21778) );
  OR2_X1 U21670 ( .A1(n21779), .A2(n21780), .ZN(n21775) );
  INV_X1 U21671 ( .A(n21777), .ZN(n21780) );
  OR2_X1 U21672 ( .A1(n15525), .A2(n15173), .ZN(n21422) );
  OR2_X1 U21673 ( .A1(n21781), .A2(n21782), .ZN(n21419) );
  INV_X1 U21674 ( .A(n21783), .ZN(n21782) );
  OR2_X1 U21675 ( .A1(n21784), .A2(n21785), .ZN(n21783) );
  AND2_X1 U21676 ( .A1(n21785), .A2(n21784), .ZN(n21781) );
  AND2_X1 U21677 ( .A1(n21786), .A2(n21787), .ZN(n21784) );
  OR2_X1 U21678 ( .A1(n21788), .A2(n21789), .ZN(n21787) );
  INV_X1 U21679 ( .A(n21790), .ZN(n21789) );
  OR2_X1 U21680 ( .A1(n21790), .A2(n21791), .ZN(n21786) );
  INV_X1 U21681 ( .A(n21788), .ZN(n21791) );
  OR2_X1 U21682 ( .A1(n15559), .A2(n15173), .ZN(n21436) );
  OR2_X1 U21683 ( .A1(n21792), .A2(n21793), .ZN(n21430) );
  INV_X1 U21684 ( .A(n21794), .ZN(n21793) );
  OR2_X1 U21685 ( .A1(n21795), .A2(n21796), .ZN(n21794) );
  AND2_X1 U21686 ( .A1(n21796), .A2(n21795), .ZN(n21792) );
  AND2_X1 U21687 ( .A1(n21797), .A2(n21798), .ZN(n21795) );
  INV_X1 U21688 ( .A(n21799), .ZN(n21798) );
  AND2_X1 U21689 ( .A1(n21800), .A2(n21801), .ZN(n21799) );
  OR2_X1 U21690 ( .A1(n21801), .A2(n21800), .ZN(n21797) );
  INV_X1 U21691 ( .A(n21802), .ZN(n21800) );
  OR2_X1 U21692 ( .A1(n15593), .A2(n15173), .ZN(n21446) );
  AND2_X1 U21693 ( .A1(n21803), .A2(n21804), .ZN(n21441) );
  INV_X1 U21694 ( .A(n21805), .ZN(n21804) );
  AND2_X1 U21695 ( .A1(n21806), .A2(n21807), .ZN(n21805) );
  OR2_X1 U21696 ( .A1(n21807), .A2(n21806), .ZN(n21803) );
  OR2_X1 U21697 ( .A1(n21808), .A2(n21809), .ZN(n21806) );
  AND2_X1 U21698 ( .A1(n21810), .A2(n21811), .ZN(n21809) );
  INV_X1 U21699 ( .A(n21812), .ZN(n21810) );
  AND2_X1 U21700 ( .A1(n21813), .A2(n21812), .ZN(n21808) );
  INV_X1 U21701 ( .A(n21811), .ZN(n21813) );
  OR2_X1 U21702 ( .A1(n15638), .A2(n15173), .ZN(n21457) );
  AND2_X1 U21703 ( .A1(n21814), .A2(n21815), .ZN(n21452) );
  INV_X1 U21704 ( .A(n21816), .ZN(n21815) );
  AND2_X1 U21705 ( .A1(n21817), .A2(n21818), .ZN(n21816) );
  OR2_X1 U21706 ( .A1(n21818), .A2(n21817), .ZN(n21814) );
  OR2_X1 U21707 ( .A1(n21819), .A2(n21820), .ZN(n21817) );
  AND2_X1 U21708 ( .A1(n21821), .A2(n21822), .ZN(n21820) );
  INV_X1 U21709 ( .A(n21823), .ZN(n21821) );
  AND2_X1 U21710 ( .A1(n21824), .A2(n21823), .ZN(n21819) );
  INV_X1 U21711 ( .A(n21822), .ZN(n21824) );
  OR2_X1 U21712 ( .A1(n15672), .A2(n15173), .ZN(n21468) );
  AND2_X1 U21713 ( .A1(n21825), .A2(n21826), .ZN(n21463) );
  INV_X1 U21714 ( .A(n21827), .ZN(n21826) );
  AND2_X1 U21715 ( .A1(n21828), .A2(n21829), .ZN(n21827) );
  OR2_X1 U21716 ( .A1(n21829), .A2(n21828), .ZN(n21825) );
  OR2_X1 U21717 ( .A1(n21830), .A2(n21831), .ZN(n21828) );
  AND2_X1 U21718 ( .A1(n21832), .A2(n21833), .ZN(n21831) );
  INV_X1 U21719 ( .A(n21834), .ZN(n21832) );
  AND2_X1 U21720 ( .A1(n21835), .A2(n21834), .ZN(n21830) );
  INV_X1 U21721 ( .A(n21833), .ZN(n21835) );
  OR2_X1 U21722 ( .A1(n15706), .A2(n15173), .ZN(n21479) );
  AND2_X1 U21723 ( .A1(n21836), .A2(n21837), .ZN(n21474) );
  INV_X1 U21724 ( .A(n21838), .ZN(n21837) );
  AND2_X1 U21725 ( .A1(n21839), .A2(n21840), .ZN(n21838) );
  OR2_X1 U21726 ( .A1(n21840), .A2(n21839), .ZN(n21836) );
  OR2_X1 U21727 ( .A1(n21841), .A2(n21842), .ZN(n21839) );
  AND2_X1 U21728 ( .A1(n21843), .A2(n21844), .ZN(n21842) );
  INV_X1 U21729 ( .A(n21845), .ZN(n21843) );
  AND2_X1 U21730 ( .A1(n21846), .A2(n21845), .ZN(n21841) );
  INV_X1 U21731 ( .A(n21844), .ZN(n21846) );
  OR2_X1 U21732 ( .A1(n15740), .A2(n15173), .ZN(n21490) );
  INV_X1 U21733 ( .A(b_20_), .ZN(n15173) );
  AND2_X1 U21734 ( .A1(n21847), .A2(n21848), .ZN(n21485) );
  INV_X1 U21735 ( .A(n21849), .ZN(n21848) );
  AND2_X1 U21736 ( .A1(n21850), .A2(n21851), .ZN(n21849) );
  OR2_X1 U21737 ( .A1(n21851), .A2(n21850), .ZN(n21847) );
  OR2_X1 U21738 ( .A1(n21852), .A2(n21853), .ZN(n21850) );
  AND2_X1 U21739 ( .A1(n21854), .A2(n21855), .ZN(n21853) );
  INV_X1 U21740 ( .A(n21856), .ZN(n21854) );
  AND2_X1 U21741 ( .A1(n21857), .A2(n21856), .ZN(n21852) );
  INV_X1 U21742 ( .A(n21855), .ZN(n21857) );
  AND2_X1 U21743 ( .A1(n21858), .A2(n21859), .ZN(n20302) );
  INV_X1 U21744 ( .A(n21860), .ZN(n21859) );
  AND2_X1 U21745 ( .A1(n21861), .A2(n21862), .ZN(n21860) );
  OR2_X1 U21746 ( .A1(n21862), .A2(n21861), .ZN(n21858) );
  OR2_X1 U21747 ( .A1(n21863), .A2(n21864), .ZN(n21861) );
  AND2_X1 U21748 ( .A1(n21865), .A2(n21866), .ZN(n21864) );
  INV_X1 U21749 ( .A(n21867), .ZN(n21865) );
  AND2_X1 U21750 ( .A1(n21868), .A2(n21867), .ZN(n21863) );
  INV_X1 U21751 ( .A(n21866), .ZN(n21868) );
  OR2_X1 U21752 ( .A1(n21869), .A2(n16665), .ZN(n16109) );
  OR2_X1 U21753 ( .A1(n21870), .A2(n21871), .ZN(n16665) );
  AND2_X1 U21754 ( .A1(n21872), .A2(n16656), .ZN(n21871) );
  INV_X1 U21755 ( .A(n16655), .ZN(n21872) );
  AND2_X1 U21756 ( .A1(n16655), .A2(n21873), .ZN(n21870) );
  INV_X1 U21757 ( .A(n16656), .ZN(n21873) );
  OR2_X1 U21758 ( .A1(n21874), .A2(n21875), .ZN(n16656) );
  AND2_X1 U21759 ( .A1(n21876), .A2(n21877), .ZN(n21875) );
  AND2_X1 U21760 ( .A1(n21878), .A2(n21879), .ZN(n21874) );
  OR2_X1 U21761 ( .A1(n21876), .A2(n21877), .ZN(n21879) );
  AND2_X1 U21762 ( .A1(n21880), .A2(n21881), .ZN(n16655) );
  INV_X1 U21763 ( .A(n21882), .ZN(n21881) );
  AND2_X1 U21764 ( .A1(n21883), .A2(n21884), .ZN(n21882) );
  OR2_X1 U21765 ( .A1(n21884), .A2(n21883), .ZN(n21880) );
  OR2_X1 U21766 ( .A1(n21885), .A2(n21886), .ZN(n21883) );
  AND2_X1 U21767 ( .A1(n21887), .A2(n21888), .ZN(n21886) );
  INV_X1 U21768 ( .A(n21889), .ZN(n21887) );
  AND2_X1 U21769 ( .A1(n21890), .A2(n21889), .ZN(n21885) );
  INV_X1 U21770 ( .A(n21888), .ZN(n21890) );
  AND2_X1 U21771 ( .A1(n16666), .A2(n16664), .ZN(n21869) );
  INV_X1 U21772 ( .A(n16676), .ZN(n16664) );
  AND2_X1 U21773 ( .A1(n21891), .A2(n21892), .ZN(n16676) );
  INV_X1 U21774 ( .A(n21893), .ZN(n21892) );
  AND2_X1 U21775 ( .A1(n21894), .A2(n21878), .ZN(n21893) );
  OR2_X1 U21776 ( .A1(n21878), .A2(n21894), .ZN(n21891) );
  OR2_X1 U21777 ( .A1(n21895), .A2(n21896), .ZN(n21894) );
  AND2_X1 U21778 ( .A1(n21897), .A2(n21877), .ZN(n21896) );
  INV_X1 U21779 ( .A(n21876), .ZN(n21897) );
  AND2_X1 U21780 ( .A1(n21898), .A2(n21876), .ZN(n21895) );
  OR2_X1 U21781 ( .A1(n16512), .A2(n15241), .ZN(n21876) );
  INV_X1 U21782 ( .A(n21877), .ZN(n21898) );
  OR2_X1 U21783 ( .A1(n21899), .A2(n21900), .ZN(n21877) );
  AND2_X1 U21784 ( .A1(n21901), .A2(n21902), .ZN(n21900) );
  AND2_X1 U21785 ( .A1(n21903), .A2(n21904), .ZN(n21899) );
  OR2_X1 U21786 ( .A1(n21901), .A2(n21902), .ZN(n21904) );
  AND2_X1 U21787 ( .A1(n21905), .A2(n21906), .ZN(n21878) );
  INV_X1 U21788 ( .A(n21907), .ZN(n21906) );
  AND2_X1 U21789 ( .A1(n21908), .A2(n21909), .ZN(n21907) );
  OR2_X1 U21790 ( .A1(n21909), .A2(n21908), .ZN(n21905) );
  OR2_X1 U21791 ( .A1(n21910), .A2(n21911), .ZN(n21908) );
  AND2_X1 U21792 ( .A1(n21912), .A2(n21913), .ZN(n21911) );
  INV_X1 U21793 ( .A(n21914), .ZN(n21912) );
  AND2_X1 U21794 ( .A1(n21915), .A2(n21914), .ZN(n21910) );
  INV_X1 U21795 ( .A(n21913), .ZN(n21915) );
  INV_X1 U21796 ( .A(n16675), .ZN(n16666) );
  OR2_X1 U21797 ( .A1(n21916), .A2(n21917), .ZN(n16675) );
  AND2_X1 U21798 ( .A1(n16701), .A2(n16700), .ZN(n21917) );
  AND2_X1 U21799 ( .A1(n16696), .A2(n21918), .ZN(n21916) );
  OR2_X1 U21800 ( .A1(n16701), .A2(n16700), .ZN(n21918) );
  OR2_X1 U21801 ( .A1(n21919), .A2(n21920), .ZN(n16700) );
  AND2_X1 U21802 ( .A1(n16740), .A2(n16739), .ZN(n21920) );
  AND2_X1 U21803 ( .A1(n16735), .A2(n21921), .ZN(n21919) );
  OR2_X1 U21804 ( .A1(n16740), .A2(n16739), .ZN(n21921) );
  OR2_X1 U21805 ( .A1(n21922), .A2(n21923), .ZN(n16739) );
  AND2_X1 U21806 ( .A1(n20260), .A2(n20259), .ZN(n21923) );
  AND2_X1 U21807 ( .A1(n20255), .A2(n21924), .ZN(n21922) );
  OR2_X1 U21808 ( .A1(n20260), .A2(n20259), .ZN(n21924) );
  OR2_X1 U21809 ( .A1(n21925), .A2(n21926), .ZN(n20259) );
  AND2_X1 U21810 ( .A1(n20313), .A2(n20312), .ZN(n21926) );
  AND2_X1 U21811 ( .A1(n20308), .A2(n21927), .ZN(n21925) );
  OR2_X1 U21812 ( .A1(n20313), .A2(n20312), .ZN(n21927) );
  OR2_X1 U21813 ( .A1(n21928), .A2(n21929), .ZN(n20312) );
  AND2_X1 U21814 ( .A1(n21867), .A2(n21866), .ZN(n21929) );
  AND2_X1 U21815 ( .A1(n21862), .A2(n21930), .ZN(n21928) );
  OR2_X1 U21816 ( .A1(n21867), .A2(n21866), .ZN(n21930) );
  OR2_X1 U21817 ( .A1(n21931), .A2(n21932), .ZN(n21866) );
  AND2_X1 U21818 ( .A1(n21856), .A2(n21855), .ZN(n21932) );
  AND2_X1 U21819 ( .A1(n21851), .A2(n21933), .ZN(n21931) );
  OR2_X1 U21820 ( .A1(n21856), .A2(n21855), .ZN(n21933) );
  OR2_X1 U21821 ( .A1(n21934), .A2(n21935), .ZN(n21855) );
  AND2_X1 U21822 ( .A1(n21845), .A2(n21844), .ZN(n21935) );
  AND2_X1 U21823 ( .A1(n21840), .A2(n21936), .ZN(n21934) );
  OR2_X1 U21824 ( .A1(n21845), .A2(n21844), .ZN(n21936) );
  OR2_X1 U21825 ( .A1(n21937), .A2(n21938), .ZN(n21844) );
  AND2_X1 U21826 ( .A1(n21834), .A2(n21833), .ZN(n21938) );
  AND2_X1 U21827 ( .A1(n21829), .A2(n21939), .ZN(n21937) );
  OR2_X1 U21828 ( .A1(n21834), .A2(n21833), .ZN(n21939) );
  OR2_X1 U21829 ( .A1(n21940), .A2(n21941), .ZN(n21833) );
  AND2_X1 U21830 ( .A1(n21823), .A2(n21822), .ZN(n21941) );
  AND2_X1 U21831 ( .A1(n21818), .A2(n21942), .ZN(n21940) );
  OR2_X1 U21832 ( .A1(n21823), .A2(n21822), .ZN(n21942) );
  OR2_X1 U21833 ( .A1(n21943), .A2(n21944), .ZN(n21822) );
  AND2_X1 U21834 ( .A1(n21812), .A2(n21811), .ZN(n21944) );
  AND2_X1 U21835 ( .A1(n21807), .A2(n21945), .ZN(n21943) );
  OR2_X1 U21836 ( .A1(n21812), .A2(n21811), .ZN(n21945) );
  OR2_X1 U21837 ( .A1(n21946), .A2(n21947), .ZN(n21811) );
  AND2_X1 U21838 ( .A1(n21802), .A2(n21801), .ZN(n21947) );
  AND2_X1 U21839 ( .A1(n21796), .A2(n21948), .ZN(n21946) );
  OR2_X1 U21840 ( .A1(n21802), .A2(n21801), .ZN(n21948) );
  OR2_X1 U21841 ( .A1(n21949), .A2(n21950), .ZN(n21801) );
  AND2_X1 U21842 ( .A1(n21788), .A2(n21790), .ZN(n21950) );
  AND2_X1 U21843 ( .A1(n21785), .A2(n21951), .ZN(n21949) );
  OR2_X1 U21844 ( .A1(n21788), .A2(n21790), .ZN(n21951) );
  OR2_X1 U21845 ( .A1(n21952), .A2(n21953), .ZN(n21790) );
  AND2_X1 U21846 ( .A1(n21777), .A2(n21779), .ZN(n21953) );
  AND2_X1 U21847 ( .A1(n21774), .A2(n21954), .ZN(n21952) );
  OR2_X1 U21848 ( .A1(n21777), .A2(n21779), .ZN(n21954) );
  OR2_X1 U21849 ( .A1(n21955), .A2(n21956), .ZN(n21779) );
  AND2_X1 U21850 ( .A1(n21766), .A2(n21768), .ZN(n21956) );
  AND2_X1 U21851 ( .A1(n21763), .A2(n21957), .ZN(n21955) );
  OR2_X1 U21852 ( .A1(n21766), .A2(n21768), .ZN(n21957) );
  OR2_X1 U21853 ( .A1(n21958), .A2(n21959), .ZN(n21768) );
  AND2_X1 U21854 ( .A1(n21755), .A2(n21757), .ZN(n21959) );
  AND2_X1 U21855 ( .A1(n21752), .A2(n21960), .ZN(n21958) );
  OR2_X1 U21856 ( .A1(n21755), .A2(n21757), .ZN(n21960) );
  OR2_X1 U21857 ( .A1(n21961), .A2(n21962), .ZN(n21757) );
  AND2_X1 U21858 ( .A1(n21744), .A2(n21746), .ZN(n21962) );
  AND2_X1 U21859 ( .A1(n21741), .A2(n21963), .ZN(n21961) );
  OR2_X1 U21860 ( .A1(n21744), .A2(n21746), .ZN(n21963) );
  OR2_X1 U21861 ( .A1(n21964), .A2(n21965), .ZN(n21746) );
  AND2_X1 U21862 ( .A1(n21733), .A2(n21735), .ZN(n21965) );
  AND2_X1 U21863 ( .A1(n21730), .A2(n21966), .ZN(n21964) );
  OR2_X1 U21864 ( .A1(n21733), .A2(n21735), .ZN(n21966) );
  OR2_X1 U21865 ( .A1(n21967), .A2(n21968), .ZN(n21735) );
  AND2_X1 U21866 ( .A1(n21722), .A2(n21724), .ZN(n21968) );
  AND2_X1 U21867 ( .A1(n21719), .A2(n21969), .ZN(n21967) );
  OR2_X1 U21868 ( .A1(n21722), .A2(n21724), .ZN(n21969) );
  OR2_X1 U21869 ( .A1(n21970), .A2(n21971), .ZN(n21724) );
  AND2_X1 U21870 ( .A1(n21711), .A2(n21713), .ZN(n21971) );
  AND2_X1 U21871 ( .A1(n21708), .A2(n21972), .ZN(n21970) );
  OR2_X1 U21872 ( .A1(n21711), .A2(n21713), .ZN(n21972) );
  OR2_X1 U21873 ( .A1(n21973), .A2(n21974), .ZN(n21713) );
  AND2_X1 U21874 ( .A1(n15924), .A2(n21702), .ZN(n21974) );
  AND2_X1 U21875 ( .A1(n21698), .A2(n21975), .ZN(n21973) );
  OR2_X1 U21876 ( .A1(n15924), .A2(n21702), .ZN(n21975) );
  OR2_X1 U21877 ( .A1(n21976), .A2(n21977), .ZN(n21702) );
  AND2_X1 U21878 ( .A1(n21690), .A2(n21692), .ZN(n21977) );
  AND2_X1 U21879 ( .A1(n21687), .A2(n21978), .ZN(n21976) );
  OR2_X1 U21880 ( .A1(n21690), .A2(n21692), .ZN(n21978) );
  OR2_X1 U21881 ( .A1(n21979), .A2(n21980), .ZN(n21692) );
  AND2_X1 U21882 ( .A1(n21679), .A2(n21681), .ZN(n21980) );
  AND2_X1 U21883 ( .A1(n21676), .A2(n21981), .ZN(n21979) );
  OR2_X1 U21884 ( .A1(n21679), .A2(n21681), .ZN(n21981) );
  OR2_X1 U21885 ( .A1(n21982), .A2(n21983), .ZN(n21681) );
  AND2_X1 U21886 ( .A1(n21668), .A2(n21670), .ZN(n21983) );
  AND2_X1 U21887 ( .A1(n21665), .A2(n21984), .ZN(n21982) );
  OR2_X1 U21888 ( .A1(n21668), .A2(n21670), .ZN(n21984) );
  OR2_X1 U21889 ( .A1(n21985), .A2(n21986), .ZN(n21670) );
  AND2_X1 U21890 ( .A1(n21657), .A2(n21659), .ZN(n21986) );
  AND2_X1 U21891 ( .A1(n21654), .A2(n21987), .ZN(n21985) );
  OR2_X1 U21892 ( .A1(n21657), .A2(n21659), .ZN(n21987) );
  OR2_X1 U21893 ( .A1(n21988), .A2(n21989), .ZN(n21659) );
  AND2_X1 U21894 ( .A1(n21646), .A2(n21648), .ZN(n21989) );
  AND2_X1 U21895 ( .A1(n21643), .A2(n21990), .ZN(n21988) );
  OR2_X1 U21896 ( .A1(n21646), .A2(n21648), .ZN(n21990) );
  OR2_X1 U21897 ( .A1(n21991), .A2(n21992), .ZN(n21648) );
  AND2_X1 U21898 ( .A1(n21635), .A2(n21637), .ZN(n21992) );
  AND2_X1 U21899 ( .A1(n21632), .A2(n21993), .ZN(n21991) );
  OR2_X1 U21900 ( .A1(n21635), .A2(n21637), .ZN(n21993) );
  OR2_X1 U21901 ( .A1(n21994), .A2(n21995), .ZN(n21637) );
  AND2_X1 U21902 ( .A1(n21624), .A2(n21626), .ZN(n21995) );
  AND2_X1 U21903 ( .A1(n21621), .A2(n21996), .ZN(n21994) );
  OR2_X1 U21904 ( .A1(n21624), .A2(n21626), .ZN(n21996) );
  OR2_X1 U21905 ( .A1(n21997), .A2(n21998), .ZN(n21626) );
  AND2_X1 U21906 ( .A1(n21613), .A2(n21615), .ZN(n21998) );
  AND2_X1 U21907 ( .A1(n21610), .A2(n21999), .ZN(n21997) );
  OR2_X1 U21908 ( .A1(n21613), .A2(n21615), .ZN(n21999) );
  OR2_X1 U21909 ( .A1(n22000), .A2(n22001), .ZN(n21615) );
  AND2_X1 U21910 ( .A1(n21602), .A2(n21604), .ZN(n22001) );
  AND2_X1 U21911 ( .A1(n21599), .A2(n22002), .ZN(n22000) );
  OR2_X1 U21912 ( .A1(n21602), .A2(n21604), .ZN(n22002) );
  OR2_X1 U21913 ( .A1(n22003), .A2(n22004), .ZN(n21604) );
  AND2_X1 U21914 ( .A1(n21587), .A2(n21592), .ZN(n22004) );
  AND2_X1 U21915 ( .A1(n21591), .A2(n22005), .ZN(n22003) );
  OR2_X1 U21916 ( .A1(n21587), .A2(n21592), .ZN(n22005) );
  INV_X1 U21917 ( .A(n21593), .ZN(n21592) );
  AND3_X1 U21918 ( .A1(b_19_), .A2(b_18_), .A3(n15957), .ZN(n21593) );
  OR2_X1 U21919 ( .A1(n14857), .A2(n15207), .ZN(n21587) );
  INV_X1 U21920 ( .A(n21594), .ZN(n21591) );
  OR2_X1 U21921 ( .A1(n22006), .A2(n22007), .ZN(n21594) );
  AND2_X1 U21922 ( .A1(b_18_), .A2(n22008), .ZN(n22007) );
  OR2_X1 U21923 ( .A1(n22009), .A2(n16981), .ZN(n22008) );
  AND2_X1 U21924 ( .A1(a_30_), .A2(n15286), .ZN(n22009) );
  AND2_X1 U21925 ( .A1(b_17_), .A2(n22010), .ZN(n22006) );
  OR2_X1 U21926 ( .A1(n22011), .A2(n14817), .ZN(n22010) );
  AND2_X1 U21927 ( .A1(a_31_), .A2(n15241), .ZN(n22011) );
  OR2_X1 U21928 ( .A1(n14891), .A2(n15207), .ZN(n21602) );
  OR2_X1 U21929 ( .A1(n22012), .A2(n22013), .ZN(n21599) );
  AND2_X1 U21930 ( .A1(n22014), .A2(n22015), .ZN(n22013) );
  INV_X1 U21931 ( .A(n22016), .ZN(n22012) );
  OR2_X1 U21932 ( .A1(n22014), .A2(n22015), .ZN(n22016) );
  OR2_X1 U21933 ( .A1(n22017), .A2(n22018), .ZN(n22014) );
  AND2_X1 U21934 ( .A1(n22019), .A2(n22020), .ZN(n22018) );
  AND2_X1 U21935 ( .A1(n22021), .A2(n22022), .ZN(n22017) );
  OR2_X1 U21936 ( .A1(n14936), .A2(n15207), .ZN(n21613) );
  OR2_X1 U21937 ( .A1(n22023), .A2(n22024), .ZN(n21610) );
  INV_X1 U21938 ( .A(n22025), .ZN(n22024) );
  OR2_X1 U21939 ( .A1(n22026), .A2(n22027), .ZN(n22025) );
  AND2_X1 U21940 ( .A1(n22027), .A2(n22026), .ZN(n22023) );
  AND2_X1 U21941 ( .A1(n22028), .A2(n22029), .ZN(n22026) );
  OR2_X1 U21942 ( .A1(n22030), .A2(n22031), .ZN(n22029) );
  INV_X1 U21943 ( .A(n22032), .ZN(n22031) );
  OR2_X1 U21944 ( .A1(n22032), .A2(n22033), .ZN(n22028) );
  INV_X1 U21945 ( .A(n22030), .ZN(n22033) );
  OR2_X1 U21946 ( .A1(n14970), .A2(n15207), .ZN(n21624) );
  OR2_X1 U21947 ( .A1(n22034), .A2(n22035), .ZN(n21621) );
  INV_X1 U21948 ( .A(n22036), .ZN(n22035) );
  OR2_X1 U21949 ( .A1(n22037), .A2(n22038), .ZN(n22036) );
  AND2_X1 U21950 ( .A1(n22038), .A2(n22037), .ZN(n22034) );
  AND2_X1 U21951 ( .A1(n22039), .A2(n22040), .ZN(n22037) );
  OR2_X1 U21952 ( .A1(n22041), .A2(n22042), .ZN(n22040) );
  INV_X1 U21953 ( .A(n22043), .ZN(n22042) );
  OR2_X1 U21954 ( .A1(n22043), .A2(n22044), .ZN(n22039) );
  INV_X1 U21955 ( .A(n22041), .ZN(n22044) );
  OR2_X1 U21956 ( .A1(n15004), .A2(n15207), .ZN(n21635) );
  OR2_X1 U21957 ( .A1(n22045), .A2(n22046), .ZN(n21632) );
  INV_X1 U21958 ( .A(n22047), .ZN(n22046) );
  OR2_X1 U21959 ( .A1(n22048), .A2(n22049), .ZN(n22047) );
  AND2_X1 U21960 ( .A1(n22049), .A2(n22048), .ZN(n22045) );
  AND2_X1 U21961 ( .A1(n22050), .A2(n22051), .ZN(n22048) );
  OR2_X1 U21962 ( .A1(n22052), .A2(n22053), .ZN(n22051) );
  INV_X1 U21963 ( .A(n22054), .ZN(n22053) );
  OR2_X1 U21964 ( .A1(n22054), .A2(n22055), .ZN(n22050) );
  INV_X1 U21965 ( .A(n22052), .ZN(n22055) );
  OR2_X1 U21966 ( .A1(n15038), .A2(n15207), .ZN(n21646) );
  OR2_X1 U21967 ( .A1(n22056), .A2(n22057), .ZN(n21643) );
  INV_X1 U21968 ( .A(n22058), .ZN(n22057) );
  OR2_X1 U21969 ( .A1(n22059), .A2(n22060), .ZN(n22058) );
  AND2_X1 U21970 ( .A1(n22060), .A2(n22059), .ZN(n22056) );
  AND2_X1 U21971 ( .A1(n22061), .A2(n22062), .ZN(n22059) );
  OR2_X1 U21972 ( .A1(n22063), .A2(n22064), .ZN(n22062) );
  INV_X1 U21973 ( .A(n22065), .ZN(n22064) );
  OR2_X1 U21974 ( .A1(n22065), .A2(n22066), .ZN(n22061) );
  INV_X1 U21975 ( .A(n22063), .ZN(n22066) );
  OR2_X1 U21976 ( .A1(n15072), .A2(n15207), .ZN(n21657) );
  OR2_X1 U21977 ( .A1(n22067), .A2(n22068), .ZN(n21654) );
  INV_X1 U21978 ( .A(n22069), .ZN(n22068) );
  OR2_X1 U21979 ( .A1(n22070), .A2(n22071), .ZN(n22069) );
  AND2_X1 U21980 ( .A1(n22071), .A2(n22070), .ZN(n22067) );
  AND2_X1 U21981 ( .A1(n22072), .A2(n22073), .ZN(n22070) );
  OR2_X1 U21982 ( .A1(n22074), .A2(n22075), .ZN(n22073) );
  INV_X1 U21983 ( .A(n22076), .ZN(n22075) );
  OR2_X1 U21984 ( .A1(n22076), .A2(n22077), .ZN(n22072) );
  INV_X1 U21985 ( .A(n22074), .ZN(n22077) );
  OR2_X1 U21986 ( .A1(n15106), .A2(n15207), .ZN(n21668) );
  OR2_X1 U21987 ( .A1(n22078), .A2(n22079), .ZN(n21665) );
  INV_X1 U21988 ( .A(n22080), .ZN(n22079) );
  OR2_X1 U21989 ( .A1(n22081), .A2(n22082), .ZN(n22080) );
  AND2_X1 U21990 ( .A1(n22082), .A2(n22081), .ZN(n22078) );
  AND2_X1 U21991 ( .A1(n22083), .A2(n22084), .ZN(n22081) );
  OR2_X1 U21992 ( .A1(n22085), .A2(n22086), .ZN(n22084) );
  INV_X1 U21993 ( .A(n22087), .ZN(n22086) );
  OR2_X1 U21994 ( .A1(n22087), .A2(n22088), .ZN(n22083) );
  INV_X1 U21995 ( .A(n22085), .ZN(n22088) );
  OR2_X1 U21996 ( .A1(n15140), .A2(n15207), .ZN(n21679) );
  OR2_X1 U21997 ( .A1(n22089), .A2(n22090), .ZN(n21676) );
  INV_X1 U21998 ( .A(n22091), .ZN(n22090) );
  OR2_X1 U21999 ( .A1(n22092), .A2(n22093), .ZN(n22091) );
  AND2_X1 U22000 ( .A1(n22093), .A2(n22092), .ZN(n22089) );
  AND2_X1 U22001 ( .A1(n22094), .A2(n22095), .ZN(n22092) );
  OR2_X1 U22002 ( .A1(n22096), .A2(n22097), .ZN(n22095) );
  INV_X1 U22003 ( .A(n22098), .ZN(n22097) );
  OR2_X1 U22004 ( .A1(n22098), .A2(n22099), .ZN(n22094) );
  INV_X1 U22005 ( .A(n22096), .ZN(n22099) );
  OR2_X1 U22006 ( .A1(n15174), .A2(n15207), .ZN(n21690) );
  OR2_X1 U22007 ( .A1(n22100), .A2(n22101), .ZN(n21687) );
  INV_X1 U22008 ( .A(n22102), .ZN(n22101) );
  OR2_X1 U22009 ( .A1(n22103), .A2(n22104), .ZN(n22102) );
  AND2_X1 U22010 ( .A1(n22104), .A2(n22103), .ZN(n22100) );
  AND2_X1 U22011 ( .A1(n22105), .A2(n22106), .ZN(n22103) );
  OR2_X1 U22012 ( .A1(n22107), .A2(n22108), .ZN(n22106) );
  INV_X1 U22013 ( .A(n22109), .ZN(n22108) );
  OR2_X1 U22014 ( .A1(n22109), .A2(n22110), .ZN(n22105) );
  INV_X1 U22015 ( .A(n22107), .ZN(n22110) );
  OR2_X1 U22016 ( .A1(n15208), .A2(n15207), .ZN(n15924) );
  OR2_X1 U22017 ( .A1(n22111), .A2(n22112), .ZN(n21698) );
  INV_X1 U22018 ( .A(n22113), .ZN(n22112) );
  OR2_X1 U22019 ( .A1(n22114), .A2(n22115), .ZN(n22113) );
  AND2_X1 U22020 ( .A1(n22115), .A2(n22114), .ZN(n22111) );
  AND2_X1 U22021 ( .A1(n22116), .A2(n22117), .ZN(n22114) );
  OR2_X1 U22022 ( .A1(n22118), .A2(n22119), .ZN(n22117) );
  INV_X1 U22023 ( .A(n22120), .ZN(n22119) );
  OR2_X1 U22024 ( .A1(n22120), .A2(n22121), .ZN(n22116) );
  INV_X1 U22025 ( .A(n22118), .ZN(n22121) );
  OR2_X1 U22026 ( .A1(n15242), .A2(n15207), .ZN(n21711) );
  OR2_X1 U22027 ( .A1(n22122), .A2(n22123), .ZN(n21708) );
  INV_X1 U22028 ( .A(n22124), .ZN(n22123) );
  OR2_X1 U22029 ( .A1(n22125), .A2(n22126), .ZN(n22124) );
  AND2_X1 U22030 ( .A1(n22126), .A2(n22125), .ZN(n22122) );
  AND2_X1 U22031 ( .A1(n22127), .A2(n22128), .ZN(n22125) );
  OR2_X1 U22032 ( .A1(n22129), .A2(n22130), .ZN(n22128) );
  INV_X1 U22033 ( .A(n22131), .ZN(n22130) );
  OR2_X1 U22034 ( .A1(n22131), .A2(n22132), .ZN(n22127) );
  INV_X1 U22035 ( .A(n22129), .ZN(n22132) );
  OR2_X1 U22036 ( .A1(n15287), .A2(n15207), .ZN(n21722) );
  OR2_X1 U22037 ( .A1(n22133), .A2(n22134), .ZN(n21719) );
  INV_X1 U22038 ( .A(n22135), .ZN(n22134) );
  OR2_X1 U22039 ( .A1(n22136), .A2(n22137), .ZN(n22135) );
  AND2_X1 U22040 ( .A1(n22137), .A2(n22136), .ZN(n22133) );
  AND2_X1 U22041 ( .A1(n22138), .A2(n22139), .ZN(n22136) );
  OR2_X1 U22042 ( .A1(n15921), .A2(n22140), .ZN(n22139) );
  INV_X1 U22043 ( .A(n22141), .ZN(n22140) );
  OR2_X1 U22044 ( .A1(n22141), .A2(n22142), .ZN(n22138) );
  INV_X1 U22045 ( .A(n15921), .ZN(n22142) );
  OR2_X1 U22046 ( .A1(n15321), .A2(n15207), .ZN(n21733) );
  OR2_X1 U22047 ( .A1(n22143), .A2(n22144), .ZN(n21730) );
  INV_X1 U22048 ( .A(n22145), .ZN(n22144) );
  OR2_X1 U22049 ( .A1(n22146), .A2(n22147), .ZN(n22145) );
  AND2_X1 U22050 ( .A1(n22147), .A2(n22146), .ZN(n22143) );
  AND2_X1 U22051 ( .A1(n22148), .A2(n22149), .ZN(n22146) );
  OR2_X1 U22052 ( .A1(n22150), .A2(n22151), .ZN(n22149) );
  INV_X1 U22053 ( .A(n22152), .ZN(n22151) );
  OR2_X1 U22054 ( .A1(n22152), .A2(n22153), .ZN(n22148) );
  INV_X1 U22055 ( .A(n22150), .ZN(n22153) );
  OR2_X1 U22056 ( .A1(n15355), .A2(n15207), .ZN(n21744) );
  OR2_X1 U22057 ( .A1(n22154), .A2(n22155), .ZN(n21741) );
  INV_X1 U22058 ( .A(n22156), .ZN(n22155) );
  OR2_X1 U22059 ( .A1(n22157), .A2(n22158), .ZN(n22156) );
  AND2_X1 U22060 ( .A1(n22158), .A2(n22157), .ZN(n22154) );
  AND2_X1 U22061 ( .A1(n22159), .A2(n22160), .ZN(n22157) );
  OR2_X1 U22062 ( .A1(n22161), .A2(n22162), .ZN(n22160) );
  INV_X1 U22063 ( .A(n22163), .ZN(n22162) );
  OR2_X1 U22064 ( .A1(n22163), .A2(n22164), .ZN(n22159) );
  INV_X1 U22065 ( .A(n22161), .ZN(n22164) );
  OR2_X1 U22066 ( .A1(n15389), .A2(n15207), .ZN(n21755) );
  OR2_X1 U22067 ( .A1(n22165), .A2(n22166), .ZN(n21752) );
  INV_X1 U22068 ( .A(n22167), .ZN(n22166) );
  OR2_X1 U22069 ( .A1(n22168), .A2(n22169), .ZN(n22167) );
  AND2_X1 U22070 ( .A1(n22169), .A2(n22168), .ZN(n22165) );
  AND2_X1 U22071 ( .A1(n22170), .A2(n22171), .ZN(n22168) );
  OR2_X1 U22072 ( .A1(n22172), .A2(n22173), .ZN(n22171) );
  INV_X1 U22073 ( .A(n22174), .ZN(n22173) );
  OR2_X1 U22074 ( .A1(n22174), .A2(n22175), .ZN(n22170) );
  INV_X1 U22075 ( .A(n22172), .ZN(n22175) );
  OR2_X1 U22076 ( .A1(n15423), .A2(n15207), .ZN(n21766) );
  OR2_X1 U22077 ( .A1(n22176), .A2(n22177), .ZN(n21763) );
  INV_X1 U22078 ( .A(n22178), .ZN(n22177) );
  OR2_X1 U22079 ( .A1(n22179), .A2(n22180), .ZN(n22178) );
  AND2_X1 U22080 ( .A1(n22180), .A2(n22179), .ZN(n22176) );
  AND2_X1 U22081 ( .A1(n22181), .A2(n22182), .ZN(n22179) );
  OR2_X1 U22082 ( .A1(n22183), .A2(n22184), .ZN(n22182) );
  INV_X1 U22083 ( .A(n22185), .ZN(n22184) );
  OR2_X1 U22084 ( .A1(n22185), .A2(n22186), .ZN(n22181) );
  INV_X1 U22085 ( .A(n22183), .ZN(n22186) );
  OR2_X1 U22086 ( .A1(n15457), .A2(n15207), .ZN(n21777) );
  OR2_X1 U22087 ( .A1(n22187), .A2(n22188), .ZN(n21774) );
  INV_X1 U22088 ( .A(n22189), .ZN(n22188) );
  OR2_X1 U22089 ( .A1(n22190), .A2(n22191), .ZN(n22189) );
  AND2_X1 U22090 ( .A1(n22191), .A2(n22190), .ZN(n22187) );
  AND2_X1 U22091 ( .A1(n22192), .A2(n22193), .ZN(n22190) );
  OR2_X1 U22092 ( .A1(n22194), .A2(n22195), .ZN(n22193) );
  INV_X1 U22093 ( .A(n22196), .ZN(n22195) );
  OR2_X1 U22094 ( .A1(n22196), .A2(n22197), .ZN(n22192) );
  INV_X1 U22095 ( .A(n22194), .ZN(n22197) );
  OR2_X1 U22096 ( .A1(n15491), .A2(n15207), .ZN(n21788) );
  OR2_X1 U22097 ( .A1(n22198), .A2(n22199), .ZN(n21785) );
  INV_X1 U22098 ( .A(n22200), .ZN(n22199) );
  OR2_X1 U22099 ( .A1(n22201), .A2(n22202), .ZN(n22200) );
  AND2_X1 U22100 ( .A1(n22202), .A2(n22201), .ZN(n22198) );
  AND2_X1 U22101 ( .A1(n22203), .A2(n22204), .ZN(n22201) );
  OR2_X1 U22102 ( .A1(n22205), .A2(n22206), .ZN(n22204) );
  INV_X1 U22103 ( .A(n22207), .ZN(n22206) );
  OR2_X1 U22104 ( .A1(n22207), .A2(n22208), .ZN(n22203) );
  INV_X1 U22105 ( .A(n22205), .ZN(n22208) );
  OR2_X1 U22106 ( .A1(n15525), .A2(n15207), .ZN(n21802) );
  OR2_X1 U22107 ( .A1(n22209), .A2(n22210), .ZN(n21796) );
  INV_X1 U22108 ( .A(n22211), .ZN(n22210) );
  OR2_X1 U22109 ( .A1(n22212), .A2(n22213), .ZN(n22211) );
  AND2_X1 U22110 ( .A1(n22213), .A2(n22212), .ZN(n22209) );
  AND2_X1 U22111 ( .A1(n22214), .A2(n22215), .ZN(n22212) );
  INV_X1 U22112 ( .A(n22216), .ZN(n22215) );
  AND2_X1 U22113 ( .A1(n22217), .A2(n22218), .ZN(n22216) );
  OR2_X1 U22114 ( .A1(n22218), .A2(n22217), .ZN(n22214) );
  INV_X1 U22115 ( .A(n22219), .ZN(n22217) );
  OR2_X1 U22116 ( .A1(n15559), .A2(n15207), .ZN(n21812) );
  AND2_X1 U22117 ( .A1(n22220), .A2(n22221), .ZN(n21807) );
  INV_X1 U22118 ( .A(n22222), .ZN(n22221) );
  AND2_X1 U22119 ( .A1(n22223), .A2(n22224), .ZN(n22222) );
  OR2_X1 U22120 ( .A1(n22224), .A2(n22223), .ZN(n22220) );
  OR2_X1 U22121 ( .A1(n22225), .A2(n22226), .ZN(n22223) );
  AND2_X1 U22122 ( .A1(n22227), .A2(n22228), .ZN(n22226) );
  INV_X1 U22123 ( .A(n22229), .ZN(n22227) );
  AND2_X1 U22124 ( .A1(n22230), .A2(n22229), .ZN(n22225) );
  INV_X1 U22125 ( .A(n22228), .ZN(n22230) );
  OR2_X1 U22126 ( .A1(n15593), .A2(n15207), .ZN(n21823) );
  AND2_X1 U22127 ( .A1(n22231), .A2(n22232), .ZN(n21818) );
  INV_X1 U22128 ( .A(n22233), .ZN(n22232) );
  AND2_X1 U22129 ( .A1(n22234), .A2(n22235), .ZN(n22233) );
  OR2_X1 U22130 ( .A1(n22235), .A2(n22234), .ZN(n22231) );
  OR2_X1 U22131 ( .A1(n22236), .A2(n22237), .ZN(n22234) );
  AND2_X1 U22132 ( .A1(n22238), .A2(n22239), .ZN(n22237) );
  INV_X1 U22133 ( .A(n22240), .ZN(n22238) );
  AND2_X1 U22134 ( .A1(n22241), .A2(n22240), .ZN(n22236) );
  INV_X1 U22135 ( .A(n22239), .ZN(n22241) );
  OR2_X1 U22136 ( .A1(n15638), .A2(n15207), .ZN(n21834) );
  AND2_X1 U22137 ( .A1(n22242), .A2(n22243), .ZN(n21829) );
  INV_X1 U22138 ( .A(n22244), .ZN(n22243) );
  AND2_X1 U22139 ( .A1(n22245), .A2(n22246), .ZN(n22244) );
  OR2_X1 U22140 ( .A1(n22246), .A2(n22245), .ZN(n22242) );
  OR2_X1 U22141 ( .A1(n22247), .A2(n22248), .ZN(n22245) );
  AND2_X1 U22142 ( .A1(n22249), .A2(n22250), .ZN(n22248) );
  INV_X1 U22143 ( .A(n22251), .ZN(n22249) );
  AND2_X1 U22144 ( .A1(n22252), .A2(n22251), .ZN(n22247) );
  INV_X1 U22145 ( .A(n22250), .ZN(n22252) );
  OR2_X1 U22146 ( .A1(n15672), .A2(n15207), .ZN(n21845) );
  AND2_X1 U22147 ( .A1(n22253), .A2(n22254), .ZN(n21840) );
  INV_X1 U22148 ( .A(n22255), .ZN(n22254) );
  AND2_X1 U22149 ( .A1(n22256), .A2(n22257), .ZN(n22255) );
  OR2_X1 U22150 ( .A1(n22257), .A2(n22256), .ZN(n22253) );
  OR2_X1 U22151 ( .A1(n22258), .A2(n22259), .ZN(n22256) );
  AND2_X1 U22152 ( .A1(n22260), .A2(n22261), .ZN(n22259) );
  INV_X1 U22153 ( .A(n22262), .ZN(n22260) );
  AND2_X1 U22154 ( .A1(n22263), .A2(n22262), .ZN(n22258) );
  INV_X1 U22155 ( .A(n22261), .ZN(n22263) );
  OR2_X1 U22156 ( .A1(n15706), .A2(n15207), .ZN(n21856) );
  AND2_X1 U22157 ( .A1(n22264), .A2(n22265), .ZN(n21851) );
  INV_X1 U22158 ( .A(n22266), .ZN(n22265) );
  AND2_X1 U22159 ( .A1(n22267), .A2(n22268), .ZN(n22266) );
  OR2_X1 U22160 ( .A1(n22268), .A2(n22267), .ZN(n22264) );
  OR2_X1 U22161 ( .A1(n22269), .A2(n22270), .ZN(n22267) );
  AND2_X1 U22162 ( .A1(n22271), .A2(n22272), .ZN(n22270) );
  INV_X1 U22163 ( .A(n22273), .ZN(n22271) );
  AND2_X1 U22164 ( .A1(n22274), .A2(n22273), .ZN(n22269) );
  INV_X1 U22165 ( .A(n22272), .ZN(n22274) );
  OR2_X1 U22166 ( .A1(n15740), .A2(n15207), .ZN(n21867) );
  AND2_X1 U22167 ( .A1(n22275), .A2(n22276), .ZN(n21862) );
  INV_X1 U22168 ( .A(n22277), .ZN(n22276) );
  AND2_X1 U22169 ( .A1(n22278), .A2(n22279), .ZN(n22277) );
  OR2_X1 U22170 ( .A1(n22279), .A2(n22278), .ZN(n22275) );
  OR2_X1 U22171 ( .A1(n22280), .A2(n22281), .ZN(n22278) );
  AND2_X1 U22172 ( .A1(n22282), .A2(n22283), .ZN(n22281) );
  INV_X1 U22173 ( .A(n22284), .ZN(n22282) );
  AND2_X1 U22174 ( .A1(n22285), .A2(n22284), .ZN(n22280) );
  INV_X1 U22175 ( .A(n22283), .ZN(n22285) );
  OR2_X1 U22176 ( .A1(n15774), .A2(n15207), .ZN(n20313) );
  AND2_X1 U22177 ( .A1(n22286), .A2(n22287), .ZN(n20308) );
  INV_X1 U22178 ( .A(n22288), .ZN(n22287) );
  AND2_X1 U22179 ( .A1(n22289), .A2(n22290), .ZN(n22288) );
  OR2_X1 U22180 ( .A1(n22290), .A2(n22289), .ZN(n22286) );
  OR2_X1 U22181 ( .A1(n22291), .A2(n22292), .ZN(n22289) );
  AND2_X1 U22182 ( .A1(n22293), .A2(n22294), .ZN(n22292) );
  INV_X1 U22183 ( .A(n22295), .ZN(n22293) );
  AND2_X1 U22184 ( .A1(n22296), .A2(n22295), .ZN(n22291) );
  INV_X1 U22185 ( .A(n22294), .ZN(n22296) );
  OR2_X1 U22186 ( .A1(n15808), .A2(n15207), .ZN(n20260) );
  AND2_X1 U22187 ( .A1(n22297), .A2(n22298), .ZN(n20255) );
  INV_X1 U22188 ( .A(n22299), .ZN(n22298) );
  AND2_X1 U22189 ( .A1(n22300), .A2(n22301), .ZN(n22299) );
  OR2_X1 U22190 ( .A1(n22301), .A2(n22300), .ZN(n22297) );
  OR2_X1 U22191 ( .A1(n22302), .A2(n22303), .ZN(n22300) );
  AND2_X1 U22192 ( .A1(n22304), .A2(n22305), .ZN(n22303) );
  INV_X1 U22193 ( .A(n22306), .ZN(n22304) );
  AND2_X1 U22194 ( .A1(n22307), .A2(n22306), .ZN(n22302) );
  INV_X1 U22195 ( .A(n22305), .ZN(n22307) );
  OR2_X1 U22196 ( .A1(n15842), .A2(n15207), .ZN(n16740) );
  AND2_X1 U22197 ( .A1(n22308), .A2(n22309), .ZN(n16735) );
  INV_X1 U22198 ( .A(n22310), .ZN(n22309) );
  AND2_X1 U22199 ( .A1(n22311), .A2(n22312), .ZN(n22310) );
  OR2_X1 U22200 ( .A1(n22312), .A2(n22311), .ZN(n22308) );
  OR2_X1 U22201 ( .A1(n22313), .A2(n22314), .ZN(n22311) );
  AND2_X1 U22202 ( .A1(n22315), .A2(n22316), .ZN(n22314) );
  INV_X1 U22203 ( .A(n22317), .ZN(n22315) );
  AND2_X1 U22204 ( .A1(n22318), .A2(n22317), .ZN(n22313) );
  INV_X1 U22205 ( .A(n22316), .ZN(n22318) );
  OR2_X1 U22206 ( .A1(n16512), .A2(n15207), .ZN(n16701) );
  INV_X1 U22207 ( .A(b_19_), .ZN(n15207) );
  AND2_X1 U22208 ( .A1(n22319), .A2(n22320), .ZN(n16696) );
  INV_X1 U22209 ( .A(n22321), .ZN(n22320) );
  AND2_X1 U22210 ( .A1(n22322), .A2(n21903), .ZN(n22321) );
  OR2_X1 U22211 ( .A1(n21903), .A2(n22322), .ZN(n22319) );
  OR2_X1 U22212 ( .A1(n22323), .A2(n22324), .ZN(n22322) );
  AND2_X1 U22213 ( .A1(n22325), .A2(n21902), .ZN(n22324) );
  INV_X1 U22214 ( .A(n21901), .ZN(n22325) );
  AND2_X1 U22215 ( .A1(n22326), .A2(n21901), .ZN(n22323) );
  OR2_X1 U22216 ( .A1(n15842), .A2(n15241), .ZN(n21901) );
  INV_X1 U22217 ( .A(n21902), .ZN(n22326) );
  OR2_X1 U22218 ( .A1(n22327), .A2(n22328), .ZN(n21902) );
  AND2_X1 U22219 ( .A1(n22317), .A2(n22316), .ZN(n22328) );
  AND2_X1 U22220 ( .A1(n22312), .A2(n22329), .ZN(n22327) );
  OR2_X1 U22221 ( .A1(n22317), .A2(n22316), .ZN(n22329) );
  OR2_X1 U22222 ( .A1(n22330), .A2(n22331), .ZN(n22316) );
  AND2_X1 U22223 ( .A1(n22306), .A2(n22305), .ZN(n22331) );
  AND2_X1 U22224 ( .A1(n22301), .A2(n22332), .ZN(n22330) );
  OR2_X1 U22225 ( .A1(n22306), .A2(n22305), .ZN(n22332) );
  OR2_X1 U22226 ( .A1(n22333), .A2(n22334), .ZN(n22305) );
  AND2_X1 U22227 ( .A1(n22295), .A2(n22294), .ZN(n22334) );
  AND2_X1 U22228 ( .A1(n22290), .A2(n22335), .ZN(n22333) );
  OR2_X1 U22229 ( .A1(n22295), .A2(n22294), .ZN(n22335) );
  OR2_X1 U22230 ( .A1(n22336), .A2(n22337), .ZN(n22294) );
  AND2_X1 U22231 ( .A1(n22284), .A2(n22283), .ZN(n22337) );
  AND2_X1 U22232 ( .A1(n22279), .A2(n22338), .ZN(n22336) );
  OR2_X1 U22233 ( .A1(n22284), .A2(n22283), .ZN(n22338) );
  OR2_X1 U22234 ( .A1(n22339), .A2(n22340), .ZN(n22283) );
  AND2_X1 U22235 ( .A1(n22273), .A2(n22272), .ZN(n22340) );
  AND2_X1 U22236 ( .A1(n22268), .A2(n22341), .ZN(n22339) );
  OR2_X1 U22237 ( .A1(n22273), .A2(n22272), .ZN(n22341) );
  OR2_X1 U22238 ( .A1(n22342), .A2(n22343), .ZN(n22272) );
  AND2_X1 U22239 ( .A1(n22262), .A2(n22261), .ZN(n22343) );
  AND2_X1 U22240 ( .A1(n22257), .A2(n22344), .ZN(n22342) );
  OR2_X1 U22241 ( .A1(n22262), .A2(n22261), .ZN(n22344) );
  OR2_X1 U22242 ( .A1(n22345), .A2(n22346), .ZN(n22261) );
  AND2_X1 U22243 ( .A1(n22251), .A2(n22250), .ZN(n22346) );
  AND2_X1 U22244 ( .A1(n22246), .A2(n22347), .ZN(n22345) );
  OR2_X1 U22245 ( .A1(n22251), .A2(n22250), .ZN(n22347) );
  OR2_X1 U22246 ( .A1(n22348), .A2(n22349), .ZN(n22250) );
  AND2_X1 U22247 ( .A1(n22240), .A2(n22239), .ZN(n22349) );
  AND2_X1 U22248 ( .A1(n22235), .A2(n22350), .ZN(n22348) );
  OR2_X1 U22249 ( .A1(n22240), .A2(n22239), .ZN(n22350) );
  OR2_X1 U22250 ( .A1(n22351), .A2(n22352), .ZN(n22239) );
  AND2_X1 U22251 ( .A1(n22229), .A2(n22228), .ZN(n22352) );
  AND2_X1 U22252 ( .A1(n22224), .A2(n22353), .ZN(n22351) );
  OR2_X1 U22253 ( .A1(n22229), .A2(n22228), .ZN(n22353) );
  OR2_X1 U22254 ( .A1(n22354), .A2(n22355), .ZN(n22228) );
  AND2_X1 U22255 ( .A1(n22219), .A2(n22218), .ZN(n22355) );
  AND2_X1 U22256 ( .A1(n22213), .A2(n22356), .ZN(n22354) );
  OR2_X1 U22257 ( .A1(n22219), .A2(n22218), .ZN(n22356) );
  OR2_X1 U22258 ( .A1(n22357), .A2(n22358), .ZN(n22218) );
  AND2_X1 U22259 ( .A1(n22205), .A2(n22207), .ZN(n22358) );
  AND2_X1 U22260 ( .A1(n22202), .A2(n22359), .ZN(n22357) );
  OR2_X1 U22261 ( .A1(n22205), .A2(n22207), .ZN(n22359) );
  OR2_X1 U22262 ( .A1(n22360), .A2(n22361), .ZN(n22207) );
  AND2_X1 U22263 ( .A1(n22194), .A2(n22196), .ZN(n22361) );
  AND2_X1 U22264 ( .A1(n22191), .A2(n22362), .ZN(n22360) );
  OR2_X1 U22265 ( .A1(n22194), .A2(n22196), .ZN(n22362) );
  OR2_X1 U22266 ( .A1(n22363), .A2(n22364), .ZN(n22196) );
  AND2_X1 U22267 ( .A1(n22183), .A2(n22185), .ZN(n22364) );
  AND2_X1 U22268 ( .A1(n22180), .A2(n22365), .ZN(n22363) );
  OR2_X1 U22269 ( .A1(n22183), .A2(n22185), .ZN(n22365) );
  OR2_X1 U22270 ( .A1(n22366), .A2(n22367), .ZN(n22185) );
  AND2_X1 U22271 ( .A1(n22172), .A2(n22174), .ZN(n22367) );
  AND2_X1 U22272 ( .A1(n22169), .A2(n22368), .ZN(n22366) );
  OR2_X1 U22273 ( .A1(n22172), .A2(n22174), .ZN(n22368) );
  OR2_X1 U22274 ( .A1(n22369), .A2(n22370), .ZN(n22174) );
  AND2_X1 U22275 ( .A1(n22161), .A2(n22163), .ZN(n22370) );
  AND2_X1 U22276 ( .A1(n22158), .A2(n22371), .ZN(n22369) );
  OR2_X1 U22277 ( .A1(n22161), .A2(n22163), .ZN(n22371) );
  OR2_X1 U22278 ( .A1(n22372), .A2(n22373), .ZN(n22163) );
  AND2_X1 U22279 ( .A1(n22150), .A2(n22152), .ZN(n22373) );
  AND2_X1 U22280 ( .A1(n22147), .A2(n22374), .ZN(n22372) );
  OR2_X1 U22281 ( .A1(n22150), .A2(n22152), .ZN(n22374) );
  OR2_X1 U22282 ( .A1(n22375), .A2(n22376), .ZN(n22152) );
  AND2_X1 U22283 ( .A1(n15921), .A2(n22141), .ZN(n22376) );
  AND2_X1 U22284 ( .A1(n22137), .A2(n22377), .ZN(n22375) );
  OR2_X1 U22285 ( .A1(n15921), .A2(n22141), .ZN(n22377) );
  OR2_X1 U22286 ( .A1(n22378), .A2(n22379), .ZN(n22141) );
  AND2_X1 U22287 ( .A1(n22129), .A2(n22131), .ZN(n22379) );
  AND2_X1 U22288 ( .A1(n22126), .A2(n22380), .ZN(n22378) );
  OR2_X1 U22289 ( .A1(n22129), .A2(n22131), .ZN(n22380) );
  OR2_X1 U22290 ( .A1(n22381), .A2(n22382), .ZN(n22131) );
  AND2_X1 U22291 ( .A1(n22118), .A2(n22120), .ZN(n22382) );
  AND2_X1 U22292 ( .A1(n22115), .A2(n22383), .ZN(n22381) );
  OR2_X1 U22293 ( .A1(n22118), .A2(n22120), .ZN(n22383) );
  OR2_X1 U22294 ( .A1(n22384), .A2(n22385), .ZN(n22120) );
  AND2_X1 U22295 ( .A1(n22107), .A2(n22109), .ZN(n22385) );
  AND2_X1 U22296 ( .A1(n22104), .A2(n22386), .ZN(n22384) );
  OR2_X1 U22297 ( .A1(n22107), .A2(n22109), .ZN(n22386) );
  OR2_X1 U22298 ( .A1(n22387), .A2(n22388), .ZN(n22109) );
  AND2_X1 U22299 ( .A1(n22096), .A2(n22098), .ZN(n22388) );
  AND2_X1 U22300 ( .A1(n22093), .A2(n22389), .ZN(n22387) );
  OR2_X1 U22301 ( .A1(n22096), .A2(n22098), .ZN(n22389) );
  OR2_X1 U22302 ( .A1(n22390), .A2(n22391), .ZN(n22098) );
  AND2_X1 U22303 ( .A1(n22085), .A2(n22087), .ZN(n22391) );
  AND2_X1 U22304 ( .A1(n22082), .A2(n22392), .ZN(n22390) );
  OR2_X1 U22305 ( .A1(n22085), .A2(n22087), .ZN(n22392) );
  OR2_X1 U22306 ( .A1(n22393), .A2(n22394), .ZN(n22087) );
  AND2_X1 U22307 ( .A1(n22074), .A2(n22076), .ZN(n22394) );
  AND2_X1 U22308 ( .A1(n22071), .A2(n22395), .ZN(n22393) );
  OR2_X1 U22309 ( .A1(n22074), .A2(n22076), .ZN(n22395) );
  OR2_X1 U22310 ( .A1(n22396), .A2(n22397), .ZN(n22076) );
  AND2_X1 U22311 ( .A1(n22063), .A2(n22065), .ZN(n22397) );
  AND2_X1 U22312 ( .A1(n22060), .A2(n22398), .ZN(n22396) );
  OR2_X1 U22313 ( .A1(n22063), .A2(n22065), .ZN(n22398) );
  OR2_X1 U22314 ( .A1(n22399), .A2(n22400), .ZN(n22065) );
  AND2_X1 U22315 ( .A1(n22052), .A2(n22054), .ZN(n22400) );
  AND2_X1 U22316 ( .A1(n22049), .A2(n22401), .ZN(n22399) );
  OR2_X1 U22317 ( .A1(n22052), .A2(n22054), .ZN(n22401) );
  OR2_X1 U22318 ( .A1(n22402), .A2(n22403), .ZN(n22054) );
  AND2_X1 U22319 ( .A1(n22041), .A2(n22043), .ZN(n22403) );
  AND2_X1 U22320 ( .A1(n22038), .A2(n22404), .ZN(n22402) );
  OR2_X1 U22321 ( .A1(n22041), .A2(n22043), .ZN(n22404) );
  OR2_X1 U22322 ( .A1(n22405), .A2(n22406), .ZN(n22043) );
  AND2_X1 U22323 ( .A1(n22030), .A2(n22032), .ZN(n22406) );
  AND2_X1 U22324 ( .A1(n22027), .A2(n22407), .ZN(n22405) );
  OR2_X1 U22325 ( .A1(n22030), .A2(n22032), .ZN(n22407) );
  OR2_X1 U22326 ( .A1(n22408), .A2(n22409), .ZN(n22032) );
  AND2_X1 U22327 ( .A1(n22015), .A2(n22020), .ZN(n22409) );
  AND2_X1 U22328 ( .A1(n22019), .A2(n22410), .ZN(n22408) );
  OR2_X1 U22329 ( .A1(n22015), .A2(n22020), .ZN(n22410) );
  INV_X1 U22330 ( .A(n22021), .ZN(n22020) );
  AND3_X1 U22331 ( .A1(b_18_), .A2(b_17_), .A3(n15957), .ZN(n22021) );
  OR2_X1 U22332 ( .A1(n14857), .A2(n15241), .ZN(n22015) );
  INV_X1 U22333 ( .A(n22022), .ZN(n22019) );
  OR2_X1 U22334 ( .A1(n22411), .A2(n22412), .ZN(n22022) );
  AND2_X1 U22335 ( .A1(b_17_), .A2(n22413), .ZN(n22412) );
  OR2_X1 U22336 ( .A1(n22414), .A2(n16981), .ZN(n22413) );
  AND2_X1 U22337 ( .A1(a_30_), .A2(n15320), .ZN(n22414) );
  AND2_X1 U22338 ( .A1(b_16_), .A2(n22415), .ZN(n22411) );
  OR2_X1 U22339 ( .A1(n22416), .A2(n14817), .ZN(n22415) );
  AND2_X1 U22340 ( .A1(a_31_), .A2(n15286), .ZN(n22416) );
  OR2_X1 U22341 ( .A1(n14891), .A2(n15241), .ZN(n22030) );
  OR2_X1 U22342 ( .A1(n22417), .A2(n22418), .ZN(n22027) );
  AND2_X1 U22343 ( .A1(n22419), .A2(n22420), .ZN(n22418) );
  INV_X1 U22344 ( .A(n22421), .ZN(n22417) );
  OR2_X1 U22345 ( .A1(n22419), .A2(n22420), .ZN(n22421) );
  OR2_X1 U22346 ( .A1(n22422), .A2(n22423), .ZN(n22419) );
  AND2_X1 U22347 ( .A1(n22424), .A2(n22425), .ZN(n22423) );
  AND2_X1 U22348 ( .A1(n22426), .A2(n22427), .ZN(n22422) );
  OR2_X1 U22349 ( .A1(n14936), .A2(n15241), .ZN(n22041) );
  OR2_X1 U22350 ( .A1(n22428), .A2(n22429), .ZN(n22038) );
  INV_X1 U22351 ( .A(n22430), .ZN(n22429) );
  OR2_X1 U22352 ( .A1(n22431), .A2(n22432), .ZN(n22430) );
  AND2_X1 U22353 ( .A1(n22432), .A2(n22431), .ZN(n22428) );
  AND2_X1 U22354 ( .A1(n22433), .A2(n22434), .ZN(n22431) );
  OR2_X1 U22355 ( .A1(n22435), .A2(n22436), .ZN(n22434) );
  INV_X1 U22356 ( .A(n22437), .ZN(n22436) );
  OR2_X1 U22357 ( .A1(n22437), .A2(n22438), .ZN(n22433) );
  INV_X1 U22358 ( .A(n22435), .ZN(n22438) );
  OR2_X1 U22359 ( .A1(n14970), .A2(n15241), .ZN(n22052) );
  OR2_X1 U22360 ( .A1(n22439), .A2(n22440), .ZN(n22049) );
  INV_X1 U22361 ( .A(n22441), .ZN(n22440) );
  OR2_X1 U22362 ( .A1(n22442), .A2(n22443), .ZN(n22441) );
  AND2_X1 U22363 ( .A1(n22443), .A2(n22442), .ZN(n22439) );
  AND2_X1 U22364 ( .A1(n22444), .A2(n22445), .ZN(n22442) );
  OR2_X1 U22365 ( .A1(n22446), .A2(n22447), .ZN(n22445) );
  INV_X1 U22366 ( .A(n22448), .ZN(n22447) );
  OR2_X1 U22367 ( .A1(n22448), .A2(n22449), .ZN(n22444) );
  INV_X1 U22368 ( .A(n22446), .ZN(n22449) );
  OR2_X1 U22369 ( .A1(n15004), .A2(n15241), .ZN(n22063) );
  OR2_X1 U22370 ( .A1(n22450), .A2(n22451), .ZN(n22060) );
  INV_X1 U22371 ( .A(n22452), .ZN(n22451) );
  OR2_X1 U22372 ( .A1(n22453), .A2(n22454), .ZN(n22452) );
  AND2_X1 U22373 ( .A1(n22454), .A2(n22453), .ZN(n22450) );
  AND2_X1 U22374 ( .A1(n22455), .A2(n22456), .ZN(n22453) );
  OR2_X1 U22375 ( .A1(n22457), .A2(n22458), .ZN(n22456) );
  INV_X1 U22376 ( .A(n22459), .ZN(n22458) );
  OR2_X1 U22377 ( .A1(n22459), .A2(n22460), .ZN(n22455) );
  INV_X1 U22378 ( .A(n22457), .ZN(n22460) );
  OR2_X1 U22379 ( .A1(n15038), .A2(n15241), .ZN(n22074) );
  OR2_X1 U22380 ( .A1(n22461), .A2(n22462), .ZN(n22071) );
  INV_X1 U22381 ( .A(n22463), .ZN(n22462) );
  OR2_X1 U22382 ( .A1(n22464), .A2(n22465), .ZN(n22463) );
  AND2_X1 U22383 ( .A1(n22465), .A2(n22464), .ZN(n22461) );
  AND2_X1 U22384 ( .A1(n22466), .A2(n22467), .ZN(n22464) );
  OR2_X1 U22385 ( .A1(n22468), .A2(n22469), .ZN(n22467) );
  INV_X1 U22386 ( .A(n22470), .ZN(n22469) );
  OR2_X1 U22387 ( .A1(n22470), .A2(n22471), .ZN(n22466) );
  INV_X1 U22388 ( .A(n22468), .ZN(n22471) );
  OR2_X1 U22389 ( .A1(n15072), .A2(n15241), .ZN(n22085) );
  OR2_X1 U22390 ( .A1(n22472), .A2(n22473), .ZN(n22082) );
  INV_X1 U22391 ( .A(n22474), .ZN(n22473) );
  OR2_X1 U22392 ( .A1(n22475), .A2(n22476), .ZN(n22474) );
  AND2_X1 U22393 ( .A1(n22476), .A2(n22475), .ZN(n22472) );
  AND2_X1 U22394 ( .A1(n22477), .A2(n22478), .ZN(n22475) );
  OR2_X1 U22395 ( .A1(n22479), .A2(n22480), .ZN(n22478) );
  INV_X1 U22396 ( .A(n22481), .ZN(n22480) );
  OR2_X1 U22397 ( .A1(n22481), .A2(n22482), .ZN(n22477) );
  INV_X1 U22398 ( .A(n22479), .ZN(n22482) );
  OR2_X1 U22399 ( .A1(n15106), .A2(n15241), .ZN(n22096) );
  OR2_X1 U22400 ( .A1(n22483), .A2(n22484), .ZN(n22093) );
  INV_X1 U22401 ( .A(n22485), .ZN(n22484) );
  OR2_X1 U22402 ( .A1(n22486), .A2(n22487), .ZN(n22485) );
  AND2_X1 U22403 ( .A1(n22487), .A2(n22486), .ZN(n22483) );
  AND2_X1 U22404 ( .A1(n22488), .A2(n22489), .ZN(n22486) );
  OR2_X1 U22405 ( .A1(n22490), .A2(n22491), .ZN(n22489) );
  INV_X1 U22406 ( .A(n22492), .ZN(n22491) );
  OR2_X1 U22407 ( .A1(n22492), .A2(n22493), .ZN(n22488) );
  INV_X1 U22408 ( .A(n22490), .ZN(n22493) );
  OR2_X1 U22409 ( .A1(n15140), .A2(n15241), .ZN(n22107) );
  OR2_X1 U22410 ( .A1(n22494), .A2(n22495), .ZN(n22104) );
  INV_X1 U22411 ( .A(n22496), .ZN(n22495) );
  OR2_X1 U22412 ( .A1(n22497), .A2(n22498), .ZN(n22496) );
  AND2_X1 U22413 ( .A1(n22498), .A2(n22497), .ZN(n22494) );
  AND2_X1 U22414 ( .A1(n22499), .A2(n22500), .ZN(n22497) );
  OR2_X1 U22415 ( .A1(n22501), .A2(n22502), .ZN(n22500) );
  INV_X1 U22416 ( .A(n22503), .ZN(n22502) );
  OR2_X1 U22417 ( .A1(n22503), .A2(n22504), .ZN(n22499) );
  INV_X1 U22418 ( .A(n22501), .ZN(n22504) );
  OR2_X1 U22419 ( .A1(n15174), .A2(n15241), .ZN(n22118) );
  OR2_X1 U22420 ( .A1(n22505), .A2(n22506), .ZN(n22115) );
  INV_X1 U22421 ( .A(n22507), .ZN(n22506) );
  OR2_X1 U22422 ( .A1(n22508), .A2(n22509), .ZN(n22507) );
  AND2_X1 U22423 ( .A1(n22509), .A2(n22508), .ZN(n22505) );
  AND2_X1 U22424 ( .A1(n22510), .A2(n22511), .ZN(n22508) );
  OR2_X1 U22425 ( .A1(n22512), .A2(n22513), .ZN(n22511) );
  INV_X1 U22426 ( .A(n22514), .ZN(n22513) );
  OR2_X1 U22427 ( .A1(n22514), .A2(n22515), .ZN(n22510) );
  INV_X1 U22428 ( .A(n22512), .ZN(n22515) );
  OR2_X1 U22429 ( .A1(n15208), .A2(n15241), .ZN(n22129) );
  OR2_X1 U22430 ( .A1(n22516), .A2(n22517), .ZN(n22126) );
  INV_X1 U22431 ( .A(n22518), .ZN(n22517) );
  OR2_X1 U22432 ( .A1(n22519), .A2(n22520), .ZN(n22518) );
  AND2_X1 U22433 ( .A1(n22520), .A2(n22519), .ZN(n22516) );
  AND2_X1 U22434 ( .A1(n22521), .A2(n22522), .ZN(n22519) );
  OR2_X1 U22435 ( .A1(n22523), .A2(n22524), .ZN(n22522) );
  INV_X1 U22436 ( .A(n22525), .ZN(n22524) );
  OR2_X1 U22437 ( .A1(n22525), .A2(n22526), .ZN(n22521) );
  INV_X1 U22438 ( .A(n22523), .ZN(n22526) );
  OR2_X1 U22439 ( .A1(n15242), .A2(n15241), .ZN(n15921) );
  OR2_X1 U22440 ( .A1(n22527), .A2(n22528), .ZN(n22137) );
  INV_X1 U22441 ( .A(n22529), .ZN(n22528) );
  OR2_X1 U22442 ( .A1(n22530), .A2(n22531), .ZN(n22529) );
  AND2_X1 U22443 ( .A1(n22531), .A2(n22530), .ZN(n22527) );
  AND2_X1 U22444 ( .A1(n22532), .A2(n22533), .ZN(n22530) );
  OR2_X1 U22445 ( .A1(n22534), .A2(n22535), .ZN(n22533) );
  INV_X1 U22446 ( .A(n22536), .ZN(n22535) );
  OR2_X1 U22447 ( .A1(n22536), .A2(n22537), .ZN(n22532) );
  INV_X1 U22448 ( .A(n22534), .ZN(n22537) );
  OR2_X1 U22449 ( .A1(n15287), .A2(n15241), .ZN(n22150) );
  OR2_X1 U22450 ( .A1(n22538), .A2(n22539), .ZN(n22147) );
  INV_X1 U22451 ( .A(n22540), .ZN(n22539) );
  OR2_X1 U22452 ( .A1(n22541), .A2(n22542), .ZN(n22540) );
  AND2_X1 U22453 ( .A1(n22542), .A2(n22541), .ZN(n22538) );
  AND2_X1 U22454 ( .A1(n22543), .A2(n22544), .ZN(n22541) );
  OR2_X1 U22455 ( .A1(n22545), .A2(n22546), .ZN(n22544) );
  INV_X1 U22456 ( .A(n22547), .ZN(n22546) );
  OR2_X1 U22457 ( .A1(n22547), .A2(n22548), .ZN(n22543) );
  INV_X1 U22458 ( .A(n22545), .ZN(n22548) );
  OR2_X1 U22459 ( .A1(n15321), .A2(n15241), .ZN(n22161) );
  OR2_X1 U22460 ( .A1(n22549), .A2(n22550), .ZN(n22158) );
  INV_X1 U22461 ( .A(n22551), .ZN(n22550) );
  OR2_X1 U22462 ( .A1(n22552), .A2(n22553), .ZN(n22551) );
  AND2_X1 U22463 ( .A1(n22553), .A2(n22552), .ZN(n22549) );
  AND2_X1 U22464 ( .A1(n22554), .A2(n22555), .ZN(n22552) );
  OR2_X1 U22465 ( .A1(n15918), .A2(n22556), .ZN(n22555) );
  INV_X1 U22466 ( .A(n22557), .ZN(n22556) );
  OR2_X1 U22467 ( .A1(n22557), .A2(n22558), .ZN(n22554) );
  INV_X1 U22468 ( .A(n15918), .ZN(n22558) );
  OR2_X1 U22469 ( .A1(n15355), .A2(n15241), .ZN(n22172) );
  OR2_X1 U22470 ( .A1(n22559), .A2(n22560), .ZN(n22169) );
  INV_X1 U22471 ( .A(n22561), .ZN(n22560) );
  OR2_X1 U22472 ( .A1(n22562), .A2(n22563), .ZN(n22561) );
  AND2_X1 U22473 ( .A1(n22563), .A2(n22562), .ZN(n22559) );
  AND2_X1 U22474 ( .A1(n22564), .A2(n22565), .ZN(n22562) );
  OR2_X1 U22475 ( .A1(n22566), .A2(n22567), .ZN(n22565) );
  INV_X1 U22476 ( .A(n22568), .ZN(n22567) );
  OR2_X1 U22477 ( .A1(n22568), .A2(n22569), .ZN(n22564) );
  INV_X1 U22478 ( .A(n22566), .ZN(n22569) );
  OR2_X1 U22479 ( .A1(n15389), .A2(n15241), .ZN(n22183) );
  OR2_X1 U22480 ( .A1(n22570), .A2(n22571), .ZN(n22180) );
  INV_X1 U22481 ( .A(n22572), .ZN(n22571) );
  OR2_X1 U22482 ( .A1(n22573), .A2(n22574), .ZN(n22572) );
  AND2_X1 U22483 ( .A1(n22574), .A2(n22573), .ZN(n22570) );
  AND2_X1 U22484 ( .A1(n22575), .A2(n22576), .ZN(n22573) );
  OR2_X1 U22485 ( .A1(n22577), .A2(n22578), .ZN(n22576) );
  INV_X1 U22486 ( .A(n22579), .ZN(n22578) );
  OR2_X1 U22487 ( .A1(n22579), .A2(n22580), .ZN(n22575) );
  INV_X1 U22488 ( .A(n22577), .ZN(n22580) );
  OR2_X1 U22489 ( .A1(n15423), .A2(n15241), .ZN(n22194) );
  OR2_X1 U22490 ( .A1(n22581), .A2(n22582), .ZN(n22191) );
  INV_X1 U22491 ( .A(n22583), .ZN(n22582) );
  OR2_X1 U22492 ( .A1(n22584), .A2(n22585), .ZN(n22583) );
  AND2_X1 U22493 ( .A1(n22585), .A2(n22584), .ZN(n22581) );
  AND2_X1 U22494 ( .A1(n22586), .A2(n22587), .ZN(n22584) );
  OR2_X1 U22495 ( .A1(n22588), .A2(n22589), .ZN(n22587) );
  INV_X1 U22496 ( .A(n22590), .ZN(n22589) );
  OR2_X1 U22497 ( .A1(n22590), .A2(n22591), .ZN(n22586) );
  INV_X1 U22498 ( .A(n22588), .ZN(n22591) );
  OR2_X1 U22499 ( .A1(n15457), .A2(n15241), .ZN(n22205) );
  OR2_X1 U22500 ( .A1(n22592), .A2(n22593), .ZN(n22202) );
  INV_X1 U22501 ( .A(n22594), .ZN(n22593) );
  OR2_X1 U22502 ( .A1(n22595), .A2(n22596), .ZN(n22594) );
  AND2_X1 U22503 ( .A1(n22596), .A2(n22595), .ZN(n22592) );
  AND2_X1 U22504 ( .A1(n22597), .A2(n22598), .ZN(n22595) );
  OR2_X1 U22505 ( .A1(n22599), .A2(n22600), .ZN(n22598) );
  INV_X1 U22506 ( .A(n22601), .ZN(n22600) );
  OR2_X1 U22507 ( .A1(n22601), .A2(n22602), .ZN(n22597) );
  INV_X1 U22508 ( .A(n22599), .ZN(n22602) );
  OR2_X1 U22509 ( .A1(n15491), .A2(n15241), .ZN(n22219) );
  OR2_X1 U22510 ( .A1(n22603), .A2(n22604), .ZN(n22213) );
  INV_X1 U22511 ( .A(n22605), .ZN(n22604) );
  OR2_X1 U22512 ( .A1(n22606), .A2(n22607), .ZN(n22605) );
  AND2_X1 U22513 ( .A1(n22607), .A2(n22606), .ZN(n22603) );
  AND2_X1 U22514 ( .A1(n22608), .A2(n22609), .ZN(n22606) );
  INV_X1 U22515 ( .A(n22610), .ZN(n22609) );
  AND2_X1 U22516 ( .A1(n22611), .A2(n22612), .ZN(n22610) );
  OR2_X1 U22517 ( .A1(n22612), .A2(n22611), .ZN(n22608) );
  INV_X1 U22518 ( .A(n22613), .ZN(n22611) );
  OR2_X1 U22519 ( .A1(n15525), .A2(n15241), .ZN(n22229) );
  AND2_X1 U22520 ( .A1(n22614), .A2(n22615), .ZN(n22224) );
  INV_X1 U22521 ( .A(n22616), .ZN(n22615) );
  AND2_X1 U22522 ( .A1(n22617), .A2(n22618), .ZN(n22616) );
  OR2_X1 U22523 ( .A1(n22618), .A2(n22617), .ZN(n22614) );
  OR2_X1 U22524 ( .A1(n22619), .A2(n22620), .ZN(n22617) );
  AND2_X1 U22525 ( .A1(n22621), .A2(n22622), .ZN(n22620) );
  INV_X1 U22526 ( .A(n22623), .ZN(n22621) );
  AND2_X1 U22527 ( .A1(n22624), .A2(n22623), .ZN(n22619) );
  INV_X1 U22528 ( .A(n22622), .ZN(n22624) );
  OR2_X1 U22529 ( .A1(n15559), .A2(n15241), .ZN(n22240) );
  AND2_X1 U22530 ( .A1(n22625), .A2(n22626), .ZN(n22235) );
  INV_X1 U22531 ( .A(n22627), .ZN(n22626) );
  AND2_X1 U22532 ( .A1(n22628), .A2(n22629), .ZN(n22627) );
  OR2_X1 U22533 ( .A1(n22629), .A2(n22628), .ZN(n22625) );
  OR2_X1 U22534 ( .A1(n22630), .A2(n22631), .ZN(n22628) );
  AND2_X1 U22535 ( .A1(n22632), .A2(n22633), .ZN(n22631) );
  INV_X1 U22536 ( .A(n22634), .ZN(n22632) );
  AND2_X1 U22537 ( .A1(n22635), .A2(n22634), .ZN(n22630) );
  INV_X1 U22538 ( .A(n22633), .ZN(n22635) );
  OR2_X1 U22539 ( .A1(n15593), .A2(n15241), .ZN(n22251) );
  AND2_X1 U22540 ( .A1(n22636), .A2(n22637), .ZN(n22246) );
  INV_X1 U22541 ( .A(n22638), .ZN(n22637) );
  AND2_X1 U22542 ( .A1(n22639), .A2(n22640), .ZN(n22638) );
  OR2_X1 U22543 ( .A1(n22640), .A2(n22639), .ZN(n22636) );
  OR2_X1 U22544 ( .A1(n22641), .A2(n22642), .ZN(n22639) );
  AND2_X1 U22545 ( .A1(n22643), .A2(n22644), .ZN(n22642) );
  INV_X1 U22546 ( .A(n22645), .ZN(n22643) );
  AND2_X1 U22547 ( .A1(n22646), .A2(n22645), .ZN(n22641) );
  INV_X1 U22548 ( .A(n22644), .ZN(n22646) );
  OR2_X1 U22549 ( .A1(n15638), .A2(n15241), .ZN(n22262) );
  AND2_X1 U22550 ( .A1(n22647), .A2(n22648), .ZN(n22257) );
  INV_X1 U22551 ( .A(n22649), .ZN(n22648) );
  AND2_X1 U22552 ( .A1(n22650), .A2(n22651), .ZN(n22649) );
  OR2_X1 U22553 ( .A1(n22651), .A2(n22650), .ZN(n22647) );
  OR2_X1 U22554 ( .A1(n22652), .A2(n22653), .ZN(n22650) );
  AND2_X1 U22555 ( .A1(n22654), .A2(n22655), .ZN(n22653) );
  INV_X1 U22556 ( .A(n22656), .ZN(n22654) );
  AND2_X1 U22557 ( .A1(n22657), .A2(n22656), .ZN(n22652) );
  INV_X1 U22558 ( .A(n22655), .ZN(n22657) );
  OR2_X1 U22559 ( .A1(n15672), .A2(n15241), .ZN(n22273) );
  AND2_X1 U22560 ( .A1(n22658), .A2(n22659), .ZN(n22268) );
  INV_X1 U22561 ( .A(n22660), .ZN(n22659) );
  AND2_X1 U22562 ( .A1(n22661), .A2(n22662), .ZN(n22660) );
  OR2_X1 U22563 ( .A1(n22662), .A2(n22661), .ZN(n22658) );
  OR2_X1 U22564 ( .A1(n22663), .A2(n22664), .ZN(n22661) );
  AND2_X1 U22565 ( .A1(n22665), .A2(n22666), .ZN(n22664) );
  INV_X1 U22566 ( .A(n22667), .ZN(n22665) );
  AND2_X1 U22567 ( .A1(n22668), .A2(n22667), .ZN(n22663) );
  INV_X1 U22568 ( .A(n22666), .ZN(n22668) );
  OR2_X1 U22569 ( .A1(n15706), .A2(n15241), .ZN(n22284) );
  AND2_X1 U22570 ( .A1(n22669), .A2(n22670), .ZN(n22279) );
  INV_X1 U22571 ( .A(n22671), .ZN(n22670) );
  AND2_X1 U22572 ( .A1(n22672), .A2(n22673), .ZN(n22671) );
  OR2_X1 U22573 ( .A1(n22673), .A2(n22672), .ZN(n22669) );
  OR2_X1 U22574 ( .A1(n22674), .A2(n22675), .ZN(n22672) );
  AND2_X1 U22575 ( .A1(n22676), .A2(n22677), .ZN(n22675) );
  INV_X1 U22576 ( .A(n22678), .ZN(n22676) );
  AND2_X1 U22577 ( .A1(n22679), .A2(n22678), .ZN(n22674) );
  INV_X1 U22578 ( .A(n22677), .ZN(n22679) );
  OR2_X1 U22579 ( .A1(n15740), .A2(n15241), .ZN(n22295) );
  AND2_X1 U22580 ( .A1(n22680), .A2(n22681), .ZN(n22290) );
  INV_X1 U22581 ( .A(n22682), .ZN(n22681) );
  AND2_X1 U22582 ( .A1(n22683), .A2(n22684), .ZN(n22682) );
  OR2_X1 U22583 ( .A1(n22684), .A2(n22683), .ZN(n22680) );
  OR2_X1 U22584 ( .A1(n22685), .A2(n22686), .ZN(n22683) );
  AND2_X1 U22585 ( .A1(n22687), .A2(n22688), .ZN(n22686) );
  INV_X1 U22586 ( .A(n22689), .ZN(n22687) );
  AND2_X1 U22587 ( .A1(n22690), .A2(n22689), .ZN(n22685) );
  INV_X1 U22588 ( .A(n22688), .ZN(n22690) );
  OR2_X1 U22589 ( .A1(n15774), .A2(n15241), .ZN(n22306) );
  AND2_X1 U22590 ( .A1(n22691), .A2(n22692), .ZN(n22301) );
  INV_X1 U22591 ( .A(n22693), .ZN(n22692) );
  AND2_X1 U22592 ( .A1(n22694), .A2(n22695), .ZN(n22693) );
  OR2_X1 U22593 ( .A1(n22695), .A2(n22694), .ZN(n22691) );
  OR2_X1 U22594 ( .A1(n22696), .A2(n22697), .ZN(n22694) );
  AND2_X1 U22595 ( .A1(n22698), .A2(n22699), .ZN(n22697) );
  INV_X1 U22596 ( .A(n22700), .ZN(n22698) );
  AND2_X1 U22597 ( .A1(n22701), .A2(n22700), .ZN(n22696) );
  INV_X1 U22598 ( .A(n22699), .ZN(n22701) );
  OR2_X1 U22599 ( .A1(n15808), .A2(n15241), .ZN(n22317) );
  INV_X1 U22600 ( .A(b_18_), .ZN(n15241) );
  AND2_X1 U22601 ( .A1(n22702), .A2(n22703), .ZN(n22312) );
  INV_X1 U22602 ( .A(n22704), .ZN(n22703) );
  AND2_X1 U22603 ( .A1(n22705), .A2(n22706), .ZN(n22704) );
  OR2_X1 U22604 ( .A1(n22706), .A2(n22705), .ZN(n22702) );
  OR2_X1 U22605 ( .A1(n22707), .A2(n22708), .ZN(n22705) );
  AND2_X1 U22606 ( .A1(n22709), .A2(n22710), .ZN(n22708) );
  INV_X1 U22607 ( .A(n22711), .ZN(n22709) );
  AND2_X1 U22608 ( .A1(n22712), .A2(n22711), .ZN(n22707) );
  INV_X1 U22609 ( .A(n22710), .ZN(n22712) );
  AND2_X1 U22610 ( .A1(n22713), .A2(n22714), .ZN(n21903) );
  INV_X1 U22611 ( .A(n22715), .ZN(n22714) );
  AND2_X1 U22612 ( .A1(n22716), .A2(n22717), .ZN(n22715) );
  OR2_X1 U22613 ( .A1(n22717), .A2(n22716), .ZN(n22713) );
  OR2_X1 U22614 ( .A1(n22718), .A2(n22719), .ZN(n22716) );
  AND2_X1 U22615 ( .A1(n22720), .A2(n22721), .ZN(n22719) );
  INV_X1 U22616 ( .A(n22722), .ZN(n22720) );
  AND2_X1 U22617 ( .A1(n22723), .A2(n22722), .ZN(n22718) );
  INV_X1 U22618 ( .A(n22721), .ZN(n22723) );
  AND2_X1 U22619 ( .A1(n16128), .A2(n16129), .ZN(n16127) );
  INV_X1 U22620 ( .A(n22724), .ZN(n16129) );
  OR2_X1 U22621 ( .A1(n16662), .A2(n16661), .ZN(n22724) );
  OR2_X1 U22622 ( .A1(n22725), .A2(n22726), .ZN(n16661) );
  AND2_X1 U22623 ( .A1(n21889), .A2(n21888), .ZN(n22726) );
  AND2_X1 U22624 ( .A1(n21884), .A2(n22727), .ZN(n22725) );
  OR2_X1 U22625 ( .A1(n21889), .A2(n21888), .ZN(n22727) );
  OR2_X1 U22626 ( .A1(n22728), .A2(n22729), .ZN(n21888) );
  AND2_X1 U22627 ( .A1(n21914), .A2(n21913), .ZN(n22729) );
  AND2_X1 U22628 ( .A1(n21909), .A2(n22730), .ZN(n22728) );
  OR2_X1 U22629 ( .A1(n21914), .A2(n21913), .ZN(n22730) );
  OR2_X1 U22630 ( .A1(n22731), .A2(n22732), .ZN(n21913) );
  AND2_X1 U22631 ( .A1(n22722), .A2(n22721), .ZN(n22732) );
  AND2_X1 U22632 ( .A1(n22717), .A2(n22733), .ZN(n22731) );
  OR2_X1 U22633 ( .A1(n22722), .A2(n22721), .ZN(n22733) );
  OR2_X1 U22634 ( .A1(n22734), .A2(n22735), .ZN(n22721) );
  AND2_X1 U22635 ( .A1(n22711), .A2(n22710), .ZN(n22735) );
  AND2_X1 U22636 ( .A1(n22706), .A2(n22736), .ZN(n22734) );
  OR2_X1 U22637 ( .A1(n22711), .A2(n22710), .ZN(n22736) );
  OR2_X1 U22638 ( .A1(n22737), .A2(n22738), .ZN(n22710) );
  AND2_X1 U22639 ( .A1(n22700), .A2(n22699), .ZN(n22738) );
  AND2_X1 U22640 ( .A1(n22695), .A2(n22739), .ZN(n22737) );
  OR2_X1 U22641 ( .A1(n22700), .A2(n22699), .ZN(n22739) );
  OR2_X1 U22642 ( .A1(n22740), .A2(n22741), .ZN(n22699) );
  AND2_X1 U22643 ( .A1(n22689), .A2(n22688), .ZN(n22741) );
  AND2_X1 U22644 ( .A1(n22684), .A2(n22742), .ZN(n22740) );
  OR2_X1 U22645 ( .A1(n22689), .A2(n22688), .ZN(n22742) );
  OR2_X1 U22646 ( .A1(n22743), .A2(n22744), .ZN(n22688) );
  AND2_X1 U22647 ( .A1(n22678), .A2(n22677), .ZN(n22744) );
  AND2_X1 U22648 ( .A1(n22673), .A2(n22745), .ZN(n22743) );
  OR2_X1 U22649 ( .A1(n22678), .A2(n22677), .ZN(n22745) );
  OR2_X1 U22650 ( .A1(n22746), .A2(n22747), .ZN(n22677) );
  AND2_X1 U22651 ( .A1(n22667), .A2(n22666), .ZN(n22747) );
  AND2_X1 U22652 ( .A1(n22662), .A2(n22748), .ZN(n22746) );
  OR2_X1 U22653 ( .A1(n22667), .A2(n22666), .ZN(n22748) );
  OR2_X1 U22654 ( .A1(n22749), .A2(n22750), .ZN(n22666) );
  AND2_X1 U22655 ( .A1(n22656), .A2(n22655), .ZN(n22750) );
  AND2_X1 U22656 ( .A1(n22651), .A2(n22751), .ZN(n22749) );
  OR2_X1 U22657 ( .A1(n22656), .A2(n22655), .ZN(n22751) );
  OR2_X1 U22658 ( .A1(n22752), .A2(n22753), .ZN(n22655) );
  AND2_X1 U22659 ( .A1(n22645), .A2(n22644), .ZN(n22753) );
  AND2_X1 U22660 ( .A1(n22640), .A2(n22754), .ZN(n22752) );
  OR2_X1 U22661 ( .A1(n22645), .A2(n22644), .ZN(n22754) );
  OR2_X1 U22662 ( .A1(n22755), .A2(n22756), .ZN(n22644) );
  AND2_X1 U22663 ( .A1(n22634), .A2(n22633), .ZN(n22756) );
  AND2_X1 U22664 ( .A1(n22629), .A2(n22757), .ZN(n22755) );
  OR2_X1 U22665 ( .A1(n22634), .A2(n22633), .ZN(n22757) );
  OR2_X1 U22666 ( .A1(n22758), .A2(n22759), .ZN(n22633) );
  AND2_X1 U22667 ( .A1(n22623), .A2(n22622), .ZN(n22759) );
  AND2_X1 U22668 ( .A1(n22618), .A2(n22760), .ZN(n22758) );
  OR2_X1 U22669 ( .A1(n22623), .A2(n22622), .ZN(n22760) );
  OR2_X1 U22670 ( .A1(n22761), .A2(n22762), .ZN(n22622) );
  AND2_X1 U22671 ( .A1(n22613), .A2(n22612), .ZN(n22762) );
  AND2_X1 U22672 ( .A1(n22607), .A2(n22763), .ZN(n22761) );
  OR2_X1 U22673 ( .A1(n22613), .A2(n22612), .ZN(n22763) );
  OR2_X1 U22674 ( .A1(n22764), .A2(n22765), .ZN(n22612) );
  AND2_X1 U22675 ( .A1(n22599), .A2(n22601), .ZN(n22765) );
  AND2_X1 U22676 ( .A1(n22596), .A2(n22766), .ZN(n22764) );
  OR2_X1 U22677 ( .A1(n22599), .A2(n22601), .ZN(n22766) );
  OR2_X1 U22678 ( .A1(n22767), .A2(n22768), .ZN(n22601) );
  AND2_X1 U22679 ( .A1(n22588), .A2(n22590), .ZN(n22768) );
  AND2_X1 U22680 ( .A1(n22585), .A2(n22769), .ZN(n22767) );
  OR2_X1 U22681 ( .A1(n22588), .A2(n22590), .ZN(n22769) );
  OR2_X1 U22682 ( .A1(n22770), .A2(n22771), .ZN(n22590) );
  AND2_X1 U22683 ( .A1(n22577), .A2(n22579), .ZN(n22771) );
  AND2_X1 U22684 ( .A1(n22574), .A2(n22772), .ZN(n22770) );
  OR2_X1 U22685 ( .A1(n22577), .A2(n22579), .ZN(n22772) );
  OR2_X1 U22686 ( .A1(n22773), .A2(n22774), .ZN(n22579) );
  AND2_X1 U22687 ( .A1(n22566), .A2(n22568), .ZN(n22774) );
  AND2_X1 U22688 ( .A1(n22563), .A2(n22775), .ZN(n22773) );
  OR2_X1 U22689 ( .A1(n22566), .A2(n22568), .ZN(n22775) );
  OR2_X1 U22690 ( .A1(n22776), .A2(n22777), .ZN(n22568) );
  AND2_X1 U22691 ( .A1(n15918), .A2(n22557), .ZN(n22777) );
  AND2_X1 U22692 ( .A1(n22553), .A2(n22778), .ZN(n22776) );
  OR2_X1 U22693 ( .A1(n15918), .A2(n22557), .ZN(n22778) );
  OR2_X1 U22694 ( .A1(n22779), .A2(n22780), .ZN(n22557) );
  AND2_X1 U22695 ( .A1(n22545), .A2(n22547), .ZN(n22780) );
  AND2_X1 U22696 ( .A1(n22542), .A2(n22781), .ZN(n22779) );
  OR2_X1 U22697 ( .A1(n22545), .A2(n22547), .ZN(n22781) );
  OR2_X1 U22698 ( .A1(n22782), .A2(n22783), .ZN(n22547) );
  AND2_X1 U22699 ( .A1(n22534), .A2(n22536), .ZN(n22783) );
  AND2_X1 U22700 ( .A1(n22531), .A2(n22784), .ZN(n22782) );
  OR2_X1 U22701 ( .A1(n22534), .A2(n22536), .ZN(n22784) );
  OR2_X1 U22702 ( .A1(n22785), .A2(n22786), .ZN(n22536) );
  AND2_X1 U22703 ( .A1(n22523), .A2(n22525), .ZN(n22786) );
  AND2_X1 U22704 ( .A1(n22520), .A2(n22787), .ZN(n22785) );
  OR2_X1 U22705 ( .A1(n22523), .A2(n22525), .ZN(n22787) );
  OR2_X1 U22706 ( .A1(n22788), .A2(n22789), .ZN(n22525) );
  AND2_X1 U22707 ( .A1(n22512), .A2(n22514), .ZN(n22789) );
  AND2_X1 U22708 ( .A1(n22509), .A2(n22790), .ZN(n22788) );
  OR2_X1 U22709 ( .A1(n22512), .A2(n22514), .ZN(n22790) );
  OR2_X1 U22710 ( .A1(n22791), .A2(n22792), .ZN(n22514) );
  AND2_X1 U22711 ( .A1(n22501), .A2(n22503), .ZN(n22792) );
  AND2_X1 U22712 ( .A1(n22498), .A2(n22793), .ZN(n22791) );
  OR2_X1 U22713 ( .A1(n22501), .A2(n22503), .ZN(n22793) );
  OR2_X1 U22714 ( .A1(n22794), .A2(n22795), .ZN(n22503) );
  AND2_X1 U22715 ( .A1(n22490), .A2(n22492), .ZN(n22795) );
  AND2_X1 U22716 ( .A1(n22487), .A2(n22796), .ZN(n22794) );
  OR2_X1 U22717 ( .A1(n22490), .A2(n22492), .ZN(n22796) );
  OR2_X1 U22718 ( .A1(n22797), .A2(n22798), .ZN(n22492) );
  AND2_X1 U22719 ( .A1(n22479), .A2(n22481), .ZN(n22798) );
  AND2_X1 U22720 ( .A1(n22476), .A2(n22799), .ZN(n22797) );
  OR2_X1 U22721 ( .A1(n22479), .A2(n22481), .ZN(n22799) );
  OR2_X1 U22722 ( .A1(n22800), .A2(n22801), .ZN(n22481) );
  AND2_X1 U22723 ( .A1(n22468), .A2(n22470), .ZN(n22801) );
  AND2_X1 U22724 ( .A1(n22465), .A2(n22802), .ZN(n22800) );
  OR2_X1 U22725 ( .A1(n22468), .A2(n22470), .ZN(n22802) );
  OR2_X1 U22726 ( .A1(n22803), .A2(n22804), .ZN(n22470) );
  AND2_X1 U22727 ( .A1(n22457), .A2(n22459), .ZN(n22804) );
  AND2_X1 U22728 ( .A1(n22454), .A2(n22805), .ZN(n22803) );
  OR2_X1 U22729 ( .A1(n22457), .A2(n22459), .ZN(n22805) );
  OR2_X1 U22730 ( .A1(n22806), .A2(n22807), .ZN(n22459) );
  AND2_X1 U22731 ( .A1(n22446), .A2(n22448), .ZN(n22807) );
  AND2_X1 U22732 ( .A1(n22443), .A2(n22808), .ZN(n22806) );
  OR2_X1 U22733 ( .A1(n22446), .A2(n22448), .ZN(n22808) );
  OR2_X1 U22734 ( .A1(n22809), .A2(n22810), .ZN(n22448) );
  AND2_X1 U22735 ( .A1(n22435), .A2(n22437), .ZN(n22810) );
  AND2_X1 U22736 ( .A1(n22432), .A2(n22811), .ZN(n22809) );
  OR2_X1 U22737 ( .A1(n22435), .A2(n22437), .ZN(n22811) );
  OR2_X1 U22738 ( .A1(n22812), .A2(n22813), .ZN(n22437) );
  AND2_X1 U22739 ( .A1(n22420), .A2(n22425), .ZN(n22813) );
  AND2_X1 U22740 ( .A1(n22424), .A2(n22814), .ZN(n22812) );
  OR2_X1 U22741 ( .A1(n22420), .A2(n22425), .ZN(n22814) );
  INV_X1 U22742 ( .A(n22426), .ZN(n22425) );
  AND3_X1 U22743 ( .A1(b_17_), .A2(b_16_), .A3(n15957), .ZN(n22426) );
  OR2_X1 U22744 ( .A1(n14857), .A2(n15286), .ZN(n22420) );
  INV_X1 U22745 ( .A(n22427), .ZN(n22424) );
  OR2_X1 U22746 ( .A1(n22815), .A2(n22816), .ZN(n22427) );
  AND2_X1 U22747 ( .A1(b_16_), .A2(n22817), .ZN(n22816) );
  OR2_X1 U22748 ( .A1(n22818), .A2(n16981), .ZN(n22817) );
  AND2_X1 U22749 ( .A1(a_30_), .A2(n15354), .ZN(n22818) );
  AND2_X1 U22750 ( .A1(b_15_), .A2(n22819), .ZN(n22815) );
  OR2_X1 U22751 ( .A1(n22820), .A2(n14817), .ZN(n22819) );
  AND2_X1 U22752 ( .A1(a_31_), .A2(n15320), .ZN(n22820) );
  OR2_X1 U22753 ( .A1(n14891), .A2(n15286), .ZN(n22435) );
  OR2_X1 U22754 ( .A1(n22821), .A2(n22822), .ZN(n22432) );
  AND2_X1 U22755 ( .A1(n22823), .A2(n22824), .ZN(n22822) );
  INV_X1 U22756 ( .A(n22825), .ZN(n22821) );
  OR2_X1 U22757 ( .A1(n22823), .A2(n22824), .ZN(n22825) );
  OR2_X1 U22758 ( .A1(n22826), .A2(n22827), .ZN(n22823) );
  AND2_X1 U22759 ( .A1(n22828), .A2(n22829), .ZN(n22827) );
  AND2_X1 U22760 ( .A1(n22830), .A2(n22831), .ZN(n22826) );
  OR2_X1 U22761 ( .A1(n14936), .A2(n15286), .ZN(n22446) );
  OR2_X1 U22762 ( .A1(n22832), .A2(n22833), .ZN(n22443) );
  INV_X1 U22763 ( .A(n22834), .ZN(n22833) );
  OR2_X1 U22764 ( .A1(n22835), .A2(n22836), .ZN(n22834) );
  AND2_X1 U22765 ( .A1(n22836), .A2(n22835), .ZN(n22832) );
  AND2_X1 U22766 ( .A1(n22837), .A2(n22838), .ZN(n22835) );
  OR2_X1 U22767 ( .A1(n22839), .A2(n22840), .ZN(n22838) );
  INV_X1 U22768 ( .A(n22841), .ZN(n22840) );
  OR2_X1 U22769 ( .A1(n22841), .A2(n22842), .ZN(n22837) );
  INV_X1 U22770 ( .A(n22839), .ZN(n22842) );
  OR2_X1 U22771 ( .A1(n14970), .A2(n15286), .ZN(n22457) );
  OR2_X1 U22772 ( .A1(n22843), .A2(n22844), .ZN(n22454) );
  INV_X1 U22773 ( .A(n22845), .ZN(n22844) );
  OR2_X1 U22774 ( .A1(n22846), .A2(n22847), .ZN(n22845) );
  AND2_X1 U22775 ( .A1(n22847), .A2(n22846), .ZN(n22843) );
  AND2_X1 U22776 ( .A1(n22848), .A2(n22849), .ZN(n22846) );
  OR2_X1 U22777 ( .A1(n22850), .A2(n22851), .ZN(n22849) );
  INV_X1 U22778 ( .A(n22852), .ZN(n22851) );
  OR2_X1 U22779 ( .A1(n22852), .A2(n22853), .ZN(n22848) );
  INV_X1 U22780 ( .A(n22850), .ZN(n22853) );
  OR2_X1 U22781 ( .A1(n15004), .A2(n15286), .ZN(n22468) );
  OR2_X1 U22782 ( .A1(n22854), .A2(n22855), .ZN(n22465) );
  INV_X1 U22783 ( .A(n22856), .ZN(n22855) );
  OR2_X1 U22784 ( .A1(n22857), .A2(n22858), .ZN(n22856) );
  AND2_X1 U22785 ( .A1(n22858), .A2(n22857), .ZN(n22854) );
  AND2_X1 U22786 ( .A1(n22859), .A2(n22860), .ZN(n22857) );
  OR2_X1 U22787 ( .A1(n22861), .A2(n22862), .ZN(n22860) );
  INV_X1 U22788 ( .A(n22863), .ZN(n22862) );
  OR2_X1 U22789 ( .A1(n22863), .A2(n22864), .ZN(n22859) );
  INV_X1 U22790 ( .A(n22861), .ZN(n22864) );
  OR2_X1 U22791 ( .A1(n15038), .A2(n15286), .ZN(n22479) );
  OR2_X1 U22792 ( .A1(n22865), .A2(n22866), .ZN(n22476) );
  INV_X1 U22793 ( .A(n22867), .ZN(n22866) );
  OR2_X1 U22794 ( .A1(n22868), .A2(n22869), .ZN(n22867) );
  AND2_X1 U22795 ( .A1(n22869), .A2(n22868), .ZN(n22865) );
  AND2_X1 U22796 ( .A1(n22870), .A2(n22871), .ZN(n22868) );
  OR2_X1 U22797 ( .A1(n22872), .A2(n22873), .ZN(n22871) );
  INV_X1 U22798 ( .A(n22874), .ZN(n22873) );
  OR2_X1 U22799 ( .A1(n22874), .A2(n22875), .ZN(n22870) );
  INV_X1 U22800 ( .A(n22872), .ZN(n22875) );
  OR2_X1 U22801 ( .A1(n15072), .A2(n15286), .ZN(n22490) );
  OR2_X1 U22802 ( .A1(n22876), .A2(n22877), .ZN(n22487) );
  INV_X1 U22803 ( .A(n22878), .ZN(n22877) );
  OR2_X1 U22804 ( .A1(n22879), .A2(n22880), .ZN(n22878) );
  AND2_X1 U22805 ( .A1(n22880), .A2(n22879), .ZN(n22876) );
  AND2_X1 U22806 ( .A1(n22881), .A2(n22882), .ZN(n22879) );
  OR2_X1 U22807 ( .A1(n22883), .A2(n22884), .ZN(n22882) );
  INV_X1 U22808 ( .A(n22885), .ZN(n22884) );
  OR2_X1 U22809 ( .A1(n22885), .A2(n22886), .ZN(n22881) );
  INV_X1 U22810 ( .A(n22883), .ZN(n22886) );
  OR2_X1 U22811 ( .A1(n15106), .A2(n15286), .ZN(n22501) );
  OR2_X1 U22812 ( .A1(n22887), .A2(n22888), .ZN(n22498) );
  INV_X1 U22813 ( .A(n22889), .ZN(n22888) );
  OR2_X1 U22814 ( .A1(n22890), .A2(n22891), .ZN(n22889) );
  AND2_X1 U22815 ( .A1(n22891), .A2(n22890), .ZN(n22887) );
  AND2_X1 U22816 ( .A1(n22892), .A2(n22893), .ZN(n22890) );
  OR2_X1 U22817 ( .A1(n22894), .A2(n22895), .ZN(n22893) );
  INV_X1 U22818 ( .A(n22896), .ZN(n22895) );
  OR2_X1 U22819 ( .A1(n22896), .A2(n22897), .ZN(n22892) );
  INV_X1 U22820 ( .A(n22894), .ZN(n22897) );
  OR2_X1 U22821 ( .A1(n15140), .A2(n15286), .ZN(n22512) );
  OR2_X1 U22822 ( .A1(n22898), .A2(n22899), .ZN(n22509) );
  INV_X1 U22823 ( .A(n22900), .ZN(n22899) );
  OR2_X1 U22824 ( .A1(n22901), .A2(n22902), .ZN(n22900) );
  AND2_X1 U22825 ( .A1(n22902), .A2(n22901), .ZN(n22898) );
  AND2_X1 U22826 ( .A1(n22903), .A2(n22904), .ZN(n22901) );
  OR2_X1 U22827 ( .A1(n22905), .A2(n22906), .ZN(n22904) );
  INV_X1 U22828 ( .A(n22907), .ZN(n22906) );
  OR2_X1 U22829 ( .A1(n22907), .A2(n22908), .ZN(n22903) );
  INV_X1 U22830 ( .A(n22905), .ZN(n22908) );
  OR2_X1 U22831 ( .A1(n15174), .A2(n15286), .ZN(n22523) );
  OR2_X1 U22832 ( .A1(n22909), .A2(n22910), .ZN(n22520) );
  INV_X1 U22833 ( .A(n22911), .ZN(n22910) );
  OR2_X1 U22834 ( .A1(n22912), .A2(n22913), .ZN(n22911) );
  AND2_X1 U22835 ( .A1(n22913), .A2(n22912), .ZN(n22909) );
  AND2_X1 U22836 ( .A1(n22914), .A2(n22915), .ZN(n22912) );
  OR2_X1 U22837 ( .A1(n22916), .A2(n22917), .ZN(n22915) );
  INV_X1 U22838 ( .A(n22918), .ZN(n22917) );
  OR2_X1 U22839 ( .A1(n22918), .A2(n22919), .ZN(n22914) );
  INV_X1 U22840 ( .A(n22916), .ZN(n22919) );
  OR2_X1 U22841 ( .A1(n15208), .A2(n15286), .ZN(n22534) );
  OR2_X1 U22842 ( .A1(n22920), .A2(n22921), .ZN(n22531) );
  INV_X1 U22843 ( .A(n22922), .ZN(n22921) );
  OR2_X1 U22844 ( .A1(n22923), .A2(n22924), .ZN(n22922) );
  AND2_X1 U22845 ( .A1(n22924), .A2(n22923), .ZN(n22920) );
  AND2_X1 U22846 ( .A1(n22925), .A2(n22926), .ZN(n22923) );
  OR2_X1 U22847 ( .A1(n22927), .A2(n22928), .ZN(n22926) );
  INV_X1 U22848 ( .A(n22929), .ZN(n22928) );
  OR2_X1 U22849 ( .A1(n22929), .A2(n22930), .ZN(n22925) );
  INV_X1 U22850 ( .A(n22927), .ZN(n22930) );
  OR2_X1 U22851 ( .A1(n15242), .A2(n15286), .ZN(n22545) );
  OR2_X1 U22852 ( .A1(n22931), .A2(n22932), .ZN(n22542) );
  INV_X1 U22853 ( .A(n22933), .ZN(n22932) );
  OR2_X1 U22854 ( .A1(n22934), .A2(n22935), .ZN(n22933) );
  AND2_X1 U22855 ( .A1(n22935), .A2(n22934), .ZN(n22931) );
  AND2_X1 U22856 ( .A1(n22936), .A2(n22937), .ZN(n22934) );
  OR2_X1 U22857 ( .A1(n22938), .A2(n22939), .ZN(n22937) );
  INV_X1 U22858 ( .A(n22940), .ZN(n22939) );
  OR2_X1 U22859 ( .A1(n22940), .A2(n22941), .ZN(n22936) );
  INV_X1 U22860 ( .A(n22938), .ZN(n22941) );
  OR2_X1 U22861 ( .A1(n15287), .A2(n15286), .ZN(n15918) );
  OR2_X1 U22862 ( .A1(n22942), .A2(n22943), .ZN(n22553) );
  INV_X1 U22863 ( .A(n22944), .ZN(n22943) );
  OR2_X1 U22864 ( .A1(n22945), .A2(n22946), .ZN(n22944) );
  AND2_X1 U22865 ( .A1(n22946), .A2(n22945), .ZN(n22942) );
  AND2_X1 U22866 ( .A1(n22947), .A2(n22948), .ZN(n22945) );
  OR2_X1 U22867 ( .A1(n22949), .A2(n22950), .ZN(n22948) );
  INV_X1 U22868 ( .A(n22951), .ZN(n22950) );
  OR2_X1 U22869 ( .A1(n22951), .A2(n22952), .ZN(n22947) );
  INV_X1 U22870 ( .A(n22949), .ZN(n22952) );
  OR2_X1 U22871 ( .A1(n15321), .A2(n15286), .ZN(n22566) );
  OR2_X1 U22872 ( .A1(n22953), .A2(n22954), .ZN(n22563) );
  INV_X1 U22873 ( .A(n22955), .ZN(n22954) );
  OR2_X1 U22874 ( .A1(n22956), .A2(n22957), .ZN(n22955) );
  AND2_X1 U22875 ( .A1(n22957), .A2(n22956), .ZN(n22953) );
  AND2_X1 U22876 ( .A1(n22958), .A2(n22959), .ZN(n22956) );
  OR2_X1 U22877 ( .A1(n22960), .A2(n22961), .ZN(n22959) );
  INV_X1 U22878 ( .A(n22962), .ZN(n22961) );
  OR2_X1 U22879 ( .A1(n22962), .A2(n22963), .ZN(n22958) );
  INV_X1 U22880 ( .A(n22960), .ZN(n22963) );
  OR2_X1 U22881 ( .A1(n15355), .A2(n15286), .ZN(n22577) );
  OR2_X1 U22882 ( .A1(n22964), .A2(n22965), .ZN(n22574) );
  INV_X1 U22883 ( .A(n22966), .ZN(n22965) );
  OR2_X1 U22884 ( .A1(n22967), .A2(n22968), .ZN(n22966) );
  AND2_X1 U22885 ( .A1(n22968), .A2(n22967), .ZN(n22964) );
  AND2_X1 U22886 ( .A1(n22969), .A2(n22970), .ZN(n22967) );
  OR2_X1 U22887 ( .A1(n15915), .A2(n22971), .ZN(n22970) );
  INV_X1 U22888 ( .A(n22972), .ZN(n22971) );
  OR2_X1 U22889 ( .A1(n22972), .A2(n22973), .ZN(n22969) );
  INV_X1 U22890 ( .A(n15915), .ZN(n22973) );
  OR2_X1 U22891 ( .A1(n15389), .A2(n15286), .ZN(n22588) );
  OR2_X1 U22892 ( .A1(n22974), .A2(n22975), .ZN(n22585) );
  INV_X1 U22893 ( .A(n22976), .ZN(n22975) );
  OR2_X1 U22894 ( .A1(n22977), .A2(n22978), .ZN(n22976) );
  AND2_X1 U22895 ( .A1(n22978), .A2(n22977), .ZN(n22974) );
  AND2_X1 U22896 ( .A1(n22979), .A2(n22980), .ZN(n22977) );
  OR2_X1 U22897 ( .A1(n22981), .A2(n22982), .ZN(n22980) );
  INV_X1 U22898 ( .A(n22983), .ZN(n22982) );
  OR2_X1 U22899 ( .A1(n22983), .A2(n22984), .ZN(n22979) );
  INV_X1 U22900 ( .A(n22981), .ZN(n22984) );
  OR2_X1 U22901 ( .A1(n15423), .A2(n15286), .ZN(n22599) );
  OR2_X1 U22902 ( .A1(n22985), .A2(n22986), .ZN(n22596) );
  INV_X1 U22903 ( .A(n22987), .ZN(n22986) );
  OR2_X1 U22904 ( .A1(n22988), .A2(n22989), .ZN(n22987) );
  AND2_X1 U22905 ( .A1(n22989), .A2(n22988), .ZN(n22985) );
  AND2_X1 U22906 ( .A1(n22990), .A2(n22991), .ZN(n22988) );
  OR2_X1 U22907 ( .A1(n22992), .A2(n22993), .ZN(n22991) );
  INV_X1 U22908 ( .A(n22994), .ZN(n22993) );
  OR2_X1 U22909 ( .A1(n22994), .A2(n22995), .ZN(n22990) );
  INV_X1 U22910 ( .A(n22992), .ZN(n22995) );
  OR2_X1 U22911 ( .A1(n15457), .A2(n15286), .ZN(n22613) );
  OR2_X1 U22912 ( .A1(n22996), .A2(n22997), .ZN(n22607) );
  INV_X1 U22913 ( .A(n22998), .ZN(n22997) );
  OR2_X1 U22914 ( .A1(n22999), .A2(n23000), .ZN(n22998) );
  AND2_X1 U22915 ( .A1(n23000), .A2(n22999), .ZN(n22996) );
  AND2_X1 U22916 ( .A1(n23001), .A2(n23002), .ZN(n22999) );
  INV_X1 U22917 ( .A(n23003), .ZN(n23002) );
  AND2_X1 U22918 ( .A1(n23004), .A2(n23005), .ZN(n23003) );
  OR2_X1 U22919 ( .A1(n23005), .A2(n23004), .ZN(n23001) );
  INV_X1 U22920 ( .A(n23006), .ZN(n23004) );
  OR2_X1 U22921 ( .A1(n15491), .A2(n15286), .ZN(n22623) );
  AND2_X1 U22922 ( .A1(n23007), .A2(n23008), .ZN(n22618) );
  INV_X1 U22923 ( .A(n23009), .ZN(n23008) );
  AND2_X1 U22924 ( .A1(n23010), .A2(n23011), .ZN(n23009) );
  OR2_X1 U22925 ( .A1(n23011), .A2(n23010), .ZN(n23007) );
  OR2_X1 U22926 ( .A1(n23012), .A2(n23013), .ZN(n23010) );
  AND2_X1 U22927 ( .A1(n23014), .A2(n23015), .ZN(n23013) );
  INV_X1 U22928 ( .A(n23016), .ZN(n23014) );
  AND2_X1 U22929 ( .A1(n23017), .A2(n23016), .ZN(n23012) );
  INV_X1 U22930 ( .A(n23015), .ZN(n23017) );
  OR2_X1 U22931 ( .A1(n15525), .A2(n15286), .ZN(n22634) );
  AND2_X1 U22932 ( .A1(n23018), .A2(n23019), .ZN(n22629) );
  INV_X1 U22933 ( .A(n23020), .ZN(n23019) );
  AND2_X1 U22934 ( .A1(n23021), .A2(n23022), .ZN(n23020) );
  OR2_X1 U22935 ( .A1(n23022), .A2(n23021), .ZN(n23018) );
  OR2_X1 U22936 ( .A1(n23023), .A2(n23024), .ZN(n23021) );
  AND2_X1 U22937 ( .A1(n23025), .A2(n23026), .ZN(n23024) );
  INV_X1 U22938 ( .A(n23027), .ZN(n23025) );
  AND2_X1 U22939 ( .A1(n23028), .A2(n23027), .ZN(n23023) );
  INV_X1 U22940 ( .A(n23026), .ZN(n23028) );
  OR2_X1 U22941 ( .A1(n15559), .A2(n15286), .ZN(n22645) );
  AND2_X1 U22942 ( .A1(n23029), .A2(n23030), .ZN(n22640) );
  INV_X1 U22943 ( .A(n23031), .ZN(n23030) );
  AND2_X1 U22944 ( .A1(n23032), .A2(n23033), .ZN(n23031) );
  OR2_X1 U22945 ( .A1(n23033), .A2(n23032), .ZN(n23029) );
  OR2_X1 U22946 ( .A1(n23034), .A2(n23035), .ZN(n23032) );
  AND2_X1 U22947 ( .A1(n23036), .A2(n23037), .ZN(n23035) );
  INV_X1 U22948 ( .A(n23038), .ZN(n23036) );
  AND2_X1 U22949 ( .A1(n23039), .A2(n23038), .ZN(n23034) );
  INV_X1 U22950 ( .A(n23037), .ZN(n23039) );
  OR2_X1 U22951 ( .A1(n15593), .A2(n15286), .ZN(n22656) );
  AND2_X1 U22952 ( .A1(n23040), .A2(n23041), .ZN(n22651) );
  INV_X1 U22953 ( .A(n23042), .ZN(n23041) );
  AND2_X1 U22954 ( .A1(n23043), .A2(n23044), .ZN(n23042) );
  OR2_X1 U22955 ( .A1(n23044), .A2(n23043), .ZN(n23040) );
  OR2_X1 U22956 ( .A1(n23045), .A2(n23046), .ZN(n23043) );
  AND2_X1 U22957 ( .A1(n23047), .A2(n23048), .ZN(n23046) );
  INV_X1 U22958 ( .A(n23049), .ZN(n23047) );
  AND2_X1 U22959 ( .A1(n23050), .A2(n23049), .ZN(n23045) );
  INV_X1 U22960 ( .A(n23048), .ZN(n23050) );
  OR2_X1 U22961 ( .A1(n15638), .A2(n15286), .ZN(n22667) );
  AND2_X1 U22962 ( .A1(n23051), .A2(n23052), .ZN(n22662) );
  INV_X1 U22963 ( .A(n23053), .ZN(n23052) );
  AND2_X1 U22964 ( .A1(n23054), .A2(n23055), .ZN(n23053) );
  OR2_X1 U22965 ( .A1(n23055), .A2(n23054), .ZN(n23051) );
  OR2_X1 U22966 ( .A1(n23056), .A2(n23057), .ZN(n23054) );
  AND2_X1 U22967 ( .A1(n23058), .A2(n23059), .ZN(n23057) );
  INV_X1 U22968 ( .A(n23060), .ZN(n23058) );
  AND2_X1 U22969 ( .A1(n23061), .A2(n23060), .ZN(n23056) );
  INV_X1 U22970 ( .A(n23059), .ZN(n23061) );
  OR2_X1 U22971 ( .A1(n15672), .A2(n15286), .ZN(n22678) );
  AND2_X1 U22972 ( .A1(n23062), .A2(n23063), .ZN(n22673) );
  INV_X1 U22973 ( .A(n23064), .ZN(n23063) );
  AND2_X1 U22974 ( .A1(n23065), .A2(n23066), .ZN(n23064) );
  OR2_X1 U22975 ( .A1(n23066), .A2(n23065), .ZN(n23062) );
  OR2_X1 U22976 ( .A1(n23067), .A2(n23068), .ZN(n23065) );
  AND2_X1 U22977 ( .A1(n23069), .A2(n23070), .ZN(n23068) );
  INV_X1 U22978 ( .A(n23071), .ZN(n23069) );
  AND2_X1 U22979 ( .A1(n23072), .A2(n23071), .ZN(n23067) );
  INV_X1 U22980 ( .A(n23070), .ZN(n23072) );
  OR2_X1 U22981 ( .A1(n15706), .A2(n15286), .ZN(n22689) );
  AND2_X1 U22982 ( .A1(n23073), .A2(n23074), .ZN(n22684) );
  INV_X1 U22983 ( .A(n23075), .ZN(n23074) );
  AND2_X1 U22984 ( .A1(n23076), .A2(n23077), .ZN(n23075) );
  OR2_X1 U22985 ( .A1(n23077), .A2(n23076), .ZN(n23073) );
  OR2_X1 U22986 ( .A1(n23078), .A2(n23079), .ZN(n23076) );
  AND2_X1 U22987 ( .A1(n23080), .A2(n23081), .ZN(n23079) );
  INV_X1 U22988 ( .A(n23082), .ZN(n23080) );
  AND2_X1 U22989 ( .A1(n23083), .A2(n23082), .ZN(n23078) );
  INV_X1 U22990 ( .A(n23081), .ZN(n23083) );
  OR2_X1 U22991 ( .A1(n15740), .A2(n15286), .ZN(n22700) );
  AND2_X1 U22992 ( .A1(n23084), .A2(n23085), .ZN(n22695) );
  INV_X1 U22993 ( .A(n23086), .ZN(n23085) );
  AND2_X1 U22994 ( .A1(n23087), .A2(n23088), .ZN(n23086) );
  OR2_X1 U22995 ( .A1(n23088), .A2(n23087), .ZN(n23084) );
  OR2_X1 U22996 ( .A1(n23089), .A2(n23090), .ZN(n23087) );
  AND2_X1 U22997 ( .A1(n23091), .A2(n23092), .ZN(n23090) );
  INV_X1 U22998 ( .A(n23093), .ZN(n23091) );
  AND2_X1 U22999 ( .A1(n23094), .A2(n23093), .ZN(n23089) );
  INV_X1 U23000 ( .A(n23092), .ZN(n23094) );
  OR2_X1 U23001 ( .A1(n15774), .A2(n15286), .ZN(n22711) );
  AND2_X1 U23002 ( .A1(n23095), .A2(n23096), .ZN(n22706) );
  INV_X1 U23003 ( .A(n23097), .ZN(n23096) );
  AND2_X1 U23004 ( .A1(n23098), .A2(n23099), .ZN(n23097) );
  OR2_X1 U23005 ( .A1(n23099), .A2(n23098), .ZN(n23095) );
  OR2_X1 U23006 ( .A1(n23100), .A2(n23101), .ZN(n23098) );
  AND2_X1 U23007 ( .A1(n23102), .A2(n23103), .ZN(n23101) );
  INV_X1 U23008 ( .A(n23104), .ZN(n23102) );
  AND2_X1 U23009 ( .A1(n23105), .A2(n23104), .ZN(n23100) );
  INV_X1 U23010 ( .A(n23103), .ZN(n23105) );
  OR2_X1 U23011 ( .A1(n15808), .A2(n15286), .ZN(n22722) );
  AND2_X1 U23012 ( .A1(n23106), .A2(n23107), .ZN(n22717) );
  INV_X1 U23013 ( .A(n23108), .ZN(n23107) );
  AND2_X1 U23014 ( .A1(n23109), .A2(n23110), .ZN(n23108) );
  OR2_X1 U23015 ( .A1(n23110), .A2(n23109), .ZN(n23106) );
  OR2_X1 U23016 ( .A1(n23111), .A2(n23112), .ZN(n23109) );
  AND2_X1 U23017 ( .A1(n23113), .A2(n23114), .ZN(n23112) );
  INV_X1 U23018 ( .A(n23115), .ZN(n23113) );
  AND2_X1 U23019 ( .A1(n23116), .A2(n23115), .ZN(n23111) );
  INV_X1 U23020 ( .A(n23114), .ZN(n23116) );
  OR2_X1 U23021 ( .A1(n15842), .A2(n15286), .ZN(n21914) );
  AND2_X1 U23022 ( .A1(n23117), .A2(n23118), .ZN(n21909) );
  INV_X1 U23023 ( .A(n23119), .ZN(n23118) );
  AND2_X1 U23024 ( .A1(n23120), .A2(n23121), .ZN(n23119) );
  OR2_X1 U23025 ( .A1(n23121), .A2(n23120), .ZN(n23117) );
  OR2_X1 U23026 ( .A1(n23122), .A2(n23123), .ZN(n23120) );
  AND2_X1 U23027 ( .A1(n23124), .A2(n23125), .ZN(n23123) );
  INV_X1 U23028 ( .A(n23126), .ZN(n23124) );
  AND2_X1 U23029 ( .A1(n23127), .A2(n23126), .ZN(n23122) );
  INV_X1 U23030 ( .A(n23125), .ZN(n23127) );
  OR2_X1 U23031 ( .A1(n16512), .A2(n15286), .ZN(n21889) );
  INV_X1 U23032 ( .A(b_17_), .ZN(n15286) );
  AND2_X1 U23033 ( .A1(n23128), .A2(n23129), .ZN(n21884) );
  INV_X1 U23034 ( .A(n23130), .ZN(n23129) );
  AND2_X1 U23035 ( .A1(n23131), .A2(n23132), .ZN(n23130) );
  OR2_X1 U23036 ( .A1(n23132), .A2(n23131), .ZN(n23128) );
  OR2_X1 U23037 ( .A1(n23133), .A2(n23134), .ZN(n23131) );
  AND2_X1 U23038 ( .A1(n23135), .A2(n23136), .ZN(n23134) );
  INV_X1 U23039 ( .A(n23137), .ZN(n23135) );
  AND2_X1 U23040 ( .A1(n23138), .A2(n23137), .ZN(n23133) );
  INV_X1 U23041 ( .A(n23136), .ZN(n23138) );
  AND2_X1 U23042 ( .A1(n23139), .A2(n23140), .ZN(n16662) );
  INV_X1 U23043 ( .A(n23141), .ZN(n23140) );
  AND2_X1 U23044 ( .A1(n23142), .A2(n23143), .ZN(n23141) );
  OR2_X1 U23045 ( .A1(n23143), .A2(n23142), .ZN(n23139) );
  OR2_X1 U23046 ( .A1(n23144), .A2(n23145), .ZN(n23142) );
  AND2_X1 U23047 ( .A1(n23146), .A2(n23147), .ZN(n23145) );
  INV_X1 U23048 ( .A(n23148), .ZN(n23146) );
  AND2_X1 U23049 ( .A1(n23149), .A2(n23148), .ZN(n23144) );
  INV_X1 U23050 ( .A(n23147), .ZN(n23149) );
  AND2_X1 U23051 ( .A1(n23150), .A2(n16139), .ZN(n16128) );
  INV_X1 U23052 ( .A(n23151), .ZN(n23150) );
  AND2_X1 U23053 ( .A1(n23152), .A2(n23153), .ZN(n23151) );
  OR2_X1 U23054 ( .A1(n16139), .A2(n16140), .ZN(n16137) );
  OR2_X1 U23055 ( .A1(n23154), .A2(n23155), .ZN(n16140) );
  INV_X1 U23056 ( .A(n16150), .ZN(n23155) );
  OR2_X1 U23057 ( .A1(n23156), .A2(n23157), .ZN(n16150) );
  AND2_X1 U23058 ( .A1(n23156), .A2(n23157), .ZN(n23154) );
  OR2_X1 U23059 ( .A1(n23158), .A2(n23159), .ZN(n23157) );
  AND2_X1 U23060 ( .A1(n23160), .A2(n23161), .ZN(n23159) );
  AND2_X1 U23061 ( .A1(n23162), .A2(n23163), .ZN(n23158) );
  OR2_X1 U23062 ( .A1(n23160), .A2(n23161), .ZN(n23163) );
  AND2_X1 U23063 ( .A1(n23164), .A2(n23165), .ZN(n23156) );
  INV_X1 U23064 ( .A(n23166), .ZN(n23165) );
  AND2_X1 U23065 ( .A1(n23167), .A2(n23168), .ZN(n23166) );
  OR2_X1 U23066 ( .A1(n23168), .A2(n23167), .ZN(n23164) );
  OR2_X1 U23067 ( .A1(n23169), .A2(n23170), .ZN(n23167) );
  AND2_X1 U23068 ( .A1(n23171), .A2(n23172), .ZN(n23170) );
  INV_X1 U23069 ( .A(n23173), .ZN(n23171) );
  AND2_X1 U23070 ( .A1(n23174), .A2(n23173), .ZN(n23169) );
  INV_X1 U23071 ( .A(n23172), .ZN(n23174) );
  OR2_X1 U23072 ( .A1(n23152), .A2(n23153), .ZN(n16139) );
  OR2_X1 U23073 ( .A1(n23175), .A2(n23176), .ZN(n23153) );
  AND2_X1 U23074 ( .A1(n23148), .A2(n23147), .ZN(n23176) );
  AND2_X1 U23075 ( .A1(n23143), .A2(n23177), .ZN(n23175) );
  OR2_X1 U23076 ( .A1(n23148), .A2(n23147), .ZN(n23177) );
  OR2_X1 U23077 ( .A1(n23178), .A2(n23179), .ZN(n23147) );
  AND2_X1 U23078 ( .A1(n23137), .A2(n23136), .ZN(n23179) );
  AND2_X1 U23079 ( .A1(n23132), .A2(n23180), .ZN(n23178) );
  OR2_X1 U23080 ( .A1(n23137), .A2(n23136), .ZN(n23180) );
  OR2_X1 U23081 ( .A1(n23181), .A2(n23182), .ZN(n23136) );
  AND2_X1 U23082 ( .A1(n23126), .A2(n23125), .ZN(n23182) );
  AND2_X1 U23083 ( .A1(n23121), .A2(n23183), .ZN(n23181) );
  OR2_X1 U23084 ( .A1(n23126), .A2(n23125), .ZN(n23183) );
  OR2_X1 U23085 ( .A1(n23184), .A2(n23185), .ZN(n23125) );
  AND2_X1 U23086 ( .A1(n23115), .A2(n23114), .ZN(n23185) );
  AND2_X1 U23087 ( .A1(n23110), .A2(n23186), .ZN(n23184) );
  OR2_X1 U23088 ( .A1(n23115), .A2(n23114), .ZN(n23186) );
  OR2_X1 U23089 ( .A1(n23187), .A2(n23188), .ZN(n23114) );
  AND2_X1 U23090 ( .A1(n23104), .A2(n23103), .ZN(n23188) );
  AND2_X1 U23091 ( .A1(n23099), .A2(n23189), .ZN(n23187) );
  OR2_X1 U23092 ( .A1(n23104), .A2(n23103), .ZN(n23189) );
  OR2_X1 U23093 ( .A1(n23190), .A2(n23191), .ZN(n23103) );
  AND2_X1 U23094 ( .A1(n23093), .A2(n23092), .ZN(n23191) );
  AND2_X1 U23095 ( .A1(n23088), .A2(n23192), .ZN(n23190) );
  OR2_X1 U23096 ( .A1(n23093), .A2(n23092), .ZN(n23192) );
  OR2_X1 U23097 ( .A1(n23193), .A2(n23194), .ZN(n23092) );
  AND2_X1 U23098 ( .A1(n23082), .A2(n23081), .ZN(n23194) );
  AND2_X1 U23099 ( .A1(n23077), .A2(n23195), .ZN(n23193) );
  OR2_X1 U23100 ( .A1(n23082), .A2(n23081), .ZN(n23195) );
  OR2_X1 U23101 ( .A1(n23196), .A2(n23197), .ZN(n23081) );
  AND2_X1 U23102 ( .A1(n23071), .A2(n23070), .ZN(n23197) );
  AND2_X1 U23103 ( .A1(n23066), .A2(n23198), .ZN(n23196) );
  OR2_X1 U23104 ( .A1(n23071), .A2(n23070), .ZN(n23198) );
  OR2_X1 U23105 ( .A1(n23199), .A2(n23200), .ZN(n23070) );
  AND2_X1 U23106 ( .A1(n23060), .A2(n23059), .ZN(n23200) );
  AND2_X1 U23107 ( .A1(n23055), .A2(n23201), .ZN(n23199) );
  OR2_X1 U23108 ( .A1(n23060), .A2(n23059), .ZN(n23201) );
  OR2_X1 U23109 ( .A1(n23202), .A2(n23203), .ZN(n23059) );
  AND2_X1 U23110 ( .A1(n23049), .A2(n23048), .ZN(n23203) );
  AND2_X1 U23111 ( .A1(n23044), .A2(n23204), .ZN(n23202) );
  OR2_X1 U23112 ( .A1(n23049), .A2(n23048), .ZN(n23204) );
  OR2_X1 U23113 ( .A1(n23205), .A2(n23206), .ZN(n23048) );
  AND2_X1 U23114 ( .A1(n23038), .A2(n23037), .ZN(n23206) );
  AND2_X1 U23115 ( .A1(n23033), .A2(n23207), .ZN(n23205) );
  OR2_X1 U23116 ( .A1(n23038), .A2(n23037), .ZN(n23207) );
  OR2_X1 U23117 ( .A1(n23208), .A2(n23209), .ZN(n23037) );
  AND2_X1 U23118 ( .A1(n23027), .A2(n23026), .ZN(n23209) );
  AND2_X1 U23119 ( .A1(n23022), .A2(n23210), .ZN(n23208) );
  OR2_X1 U23120 ( .A1(n23027), .A2(n23026), .ZN(n23210) );
  OR2_X1 U23121 ( .A1(n23211), .A2(n23212), .ZN(n23026) );
  AND2_X1 U23122 ( .A1(n23016), .A2(n23015), .ZN(n23212) );
  AND2_X1 U23123 ( .A1(n23011), .A2(n23213), .ZN(n23211) );
  OR2_X1 U23124 ( .A1(n23016), .A2(n23015), .ZN(n23213) );
  OR2_X1 U23125 ( .A1(n23214), .A2(n23215), .ZN(n23015) );
  AND2_X1 U23126 ( .A1(n23000), .A2(n23006), .ZN(n23215) );
  AND2_X1 U23127 ( .A1(n23216), .A2(n23005), .ZN(n23214) );
  OR2_X1 U23128 ( .A1(n23217), .A2(n23218), .ZN(n23005) );
  AND2_X1 U23129 ( .A1(n22992), .A2(n22994), .ZN(n23218) );
  AND2_X1 U23130 ( .A1(n22989), .A2(n23219), .ZN(n23217) );
  OR2_X1 U23131 ( .A1(n22992), .A2(n22994), .ZN(n23219) );
  OR2_X1 U23132 ( .A1(n23220), .A2(n23221), .ZN(n22994) );
  AND2_X1 U23133 ( .A1(n22978), .A2(n22981), .ZN(n23221) );
  AND2_X1 U23134 ( .A1(n23222), .A2(n22983), .ZN(n23220) );
  OR2_X1 U23135 ( .A1(n23223), .A2(n23224), .ZN(n22983) );
  AND2_X1 U23136 ( .A1(n22968), .A2(n15915), .ZN(n23224) );
  AND2_X1 U23137 ( .A1(n23225), .A2(n22972), .ZN(n23223) );
  OR2_X1 U23138 ( .A1(n23226), .A2(n23227), .ZN(n22972) );
  AND2_X1 U23139 ( .A1(n22957), .A2(n22960), .ZN(n23227) );
  AND2_X1 U23140 ( .A1(n23228), .A2(n22962), .ZN(n23226) );
  OR2_X1 U23141 ( .A1(n23229), .A2(n23230), .ZN(n22962) );
  AND2_X1 U23142 ( .A1(n22946), .A2(n22949), .ZN(n23230) );
  AND2_X1 U23143 ( .A1(n23231), .A2(n22951), .ZN(n23229) );
  OR2_X1 U23144 ( .A1(n23232), .A2(n23233), .ZN(n22951) );
  AND2_X1 U23145 ( .A1(n22935), .A2(n22938), .ZN(n23233) );
  AND2_X1 U23146 ( .A1(n23234), .A2(n22940), .ZN(n23232) );
  OR2_X1 U23147 ( .A1(n23235), .A2(n23236), .ZN(n22940) );
  AND2_X1 U23148 ( .A1(n22924), .A2(n22927), .ZN(n23236) );
  AND2_X1 U23149 ( .A1(n23237), .A2(n22929), .ZN(n23235) );
  OR2_X1 U23150 ( .A1(n23238), .A2(n23239), .ZN(n22929) );
  AND2_X1 U23151 ( .A1(n22913), .A2(n22916), .ZN(n23239) );
  AND2_X1 U23152 ( .A1(n23240), .A2(n22918), .ZN(n23238) );
  OR2_X1 U23153 ( .A1(n23241), .A2(n23242), .ZN(n22918) );
  AND2_X1 U23154 ( .A1(n22902), .A2(n22905), .ZN(n23242) );
  AND2_X1 U23155 ( .A1(n23243), .A2(n22907), .ZN(n23241) );
  OR2_X1 U23156 ( .A1(n23244), .A2(n23245), .ZN(n22907) );
  AND2_X1 U23157 ( .A1(n22891), .A2(n22894), .ZN(n23245) );
  AND2_X1 U23158 ( .A1(n23246), .A2(n22896), .ZN(n23244) );
  OR2_X1 U23159 ( .A1(n23247), .A2(n23248), .ZN(n22896) );
  AND2_X1 U23160 ( .A1(n22880), .A2(n22883), .ZN(n23248) );
  AND2_X1 U23161 ( .A1(n23249), .A2(n22885), .ZN(n23247) );
  OR2_X1 U23162 ( .A1(n23250), .A2(n23251), .ZN(n22885) );
  AND2_X1 U23163 ( .A1(n22869), .A2(n22872), .ZN(n23251) );
  AND2_X1 U23164 ( .A1(n23252), .A2(n22874), .ZN(n23250) );
  OR2_X1 U23165 ( .A1(n23253), .A2(n23254), .ZN(n22874) );
  AND2_X1 U23166 ( .A1(n22858), .A2(n22861), .ZN(n23254) );
  AND2_X1 U23167 ( .A1(n23255), .A2(n22863), .ZN(n23253) );
  OR2_X1 U23168 ( .A1(n23256), .A2(n23257), .ZN(n22863) );
  AND2_X1 U23169 ( .A1(n22847), .A2(n22850), .ZN(n23257) );
  AND2_X1 U23170 ( .A1(n23258), .A2(n22852), .ZN(n23256) );
  OR2_X1 U23171 ( .A1(n23259), .A2(n23260), .ZN(n22852) );
  AND2_X1 U23172 ( .A1(n22836), .A2(n22839), .ZN(n23260) );
  AND2_X1 U23173 ( .A1(n23261), .A2(n22841), .ZN(n23259) );
  OR2_X1 U23174 ( .A1(n23262), .A2(n23263), .ZN(n22841) );
  AND2_X1 U23175 ( .A1(n22824), .A2(n22829), .ZN(n23263) );
  AND2_X1 U23176 ( .A1(n22828), .A2(n23264), .ZN(n23262) );
  OR2_X1 U23177 ( .A1(n22824), .A2(n22829), .ZN(n23264) );
  INV_X1 U23178 ( .A(n22830), .ZN(n22829) );
  AND3_X1 U23179 ( .A1(b_16_), .A2(b_15_), .A3(n15957), .ZN(n22830) );
  OR2_X1 U23180 ( .A1(n14857), .A2(n15320), .ZN(n22824) );
  INV_X1 U23181 ( .A(n22831), .ZN(n22828) );
  OR2_X1 U23182 ( .A1(n23265), .A2(n23266), .ZN(n22831) );
  AND2_X1 U23183 ( .A1(b_15_), .A2(n23267), .ZN(n23266) );
  OR2_X1 U23184 ( .A1(n23268), .A2(n16981), .ZN(n23267) );
  AND2_X1 U23185 ( .A1(a_30_), .A2(n15388), .ZN(n23268) );
  AND2_X1 U23186 ( .A1(b_14_), .A2(n23269), .ZN(n23265) );
  OR2_X1 U23187 ( .A1(n23270), .A2(n14817), .ZN(n23269) );
  AND2_X1 U23188 ( .A1(a_31_), .A2(n15354), .ZN(n23270) );
  OR2_X1 U23189 ( .A1(n22836), .A2(n22839), .ZN(n23261) );
  OR2_X1 U23190 ( .A1(n14891), .A2(n15320), .ZN(n22839) );
  OR2_X1 U23191 ( .A1(n23271), .A2(n23272), .ZN(n22836) );
  AND2_X1 U23192 ( .A1(n23273), .A2(n23274), .ZN(n23272) );
  INV_X1 U23193 ( .A(n23275), .ZN(n23271) );
  OR2_X1 U23194 ( .A1(n23273), .A2(n23274), .ZN(n23275) );
  OR2_X1 U23195 ( .A1(n23276), .A2(n23277), .ZN(n23273) );
  AND2_X1 U23196 ( .A1(n23278), .A2(n23279), .ZN(n23277) );
  AND2_X1 U23197 ( .A1(n23280), .A2(n23281), .ZN(n23276) );
  OR2_X1 U23198 ( .A1(n22847), .A2(n22850), .ZN(n23258) );
  OR2_X1 U23199 ( .A1(n14936), .A2(n15320), .ZN(n22850) );
  OR2_X1 U23200 ( .A1(n23282), .A2(n23283), .ZN(n22847) );
  INV_X1 U23201 ( .A(n23284), .ZN(n23283) );
  OR2_X1 U23202 ( .A1(n23285), .A2(n23286), .ZN(n23284) );
  AND2_X1 U23203 ( .A1(n23286), .A2(n23285), .ZN(n23282) );
  AND2_X1 U23204 ( .A1(n23287), .A2(n23288), .ZN(n23285) );
  OR2_X1 U23205 ( .A1(n23289), .A2(n23290), .ZN(n23288) );
  INV_X1 U23206 ( .A(n23291), .ZN(n23290) );
  OR2_X1 U23207 ( .A1(n23291), .A2(n23292), .ZN(n23287) );
  INV_X1 U23208 ( .A(n23289), .ZN(n23292) );
  OR2_X1 U23209 ( .A1(n22858), .A2(n22861), .ZN(n23255) );
  OR2_X1 U23210 ( .A1(n14970), .A2(n15320), .ZN(n22861) );
  OR2_X1 U23211 ( .A1(n23293), .A2(n23294), .ZN(n22858) );
  INV_X1 U23212 ( .A(n23295), .ZN(n23294) );
  OR2_X1 U23213 ( .A1(n23296), .A2(n23297), .ZN(n23295) );
  AND2_X1 U23214 ( .A1(n23297), .A2(n23296), .ZN(n23293) );
  AND2_X1 U23215 ( .A1(n23298), .A2(n23299), .ZN(n23296) );
  OR2_X1 U23216 ( .A1(n23300), .A2(n23301), .ZN(n23299) );
  INV_X1 U23217 ( .A(n23302), .ZN(n23301) );
  OR2_X1 U23218 ( .A1(n23302), .A2(n23303), .ZN(n23298) );
  INV_X1 U23219 ( .A(n23300), .ZN(n23303) );
  OR2_X1 U23220 ( .A1(n22869), .A2(n22872), .ZN(n23252) );
  OR2_X1 U23221 ( .A1(n15004), .A2(n15320), .ZN(n22872) );
  OR2_X1 U23222 ( .A1(n23304), .A2(n23305), .ZN(n22869) );
  INV_X1 U23223 ( .A(n23306), .ZN(n23305) );
  OR2_X1 U23224 ( .A1(n23307), .A2(n23308), .ZN(n23306) );
  AND2_X1 U23225 ( .A1(n23308), .A2(n23307), .ZN(n23304) );
  AND2_X1 U23226 ( .A1(n23309), .A2(n23310), .ZN(n23307) );
  OR2_X1 U23227 ( .A1(n23311), .A2(n23312), .ZN(n23310) );
  INV_X1 U23228 ( .A(n23313), .ZN(n23312) );
  OR2_X1 U23229 ( .A1(n23313), .A2(n23314), .ZN(n23309) );
  INV_X1 U23230 ( .A(n23311), .ZN(n23314) );
  OR2_X1 U23231 ( .A1(n22880), .A2(n22883), .ZN(n23249) );
  OR2_X1 U23232 ( .A1(n15038), .A2(n15320), .ZN(n22883) );
  OR2_X1 U23233 ( .A1(n23315), .A2(n23316), .ZN(n22880) );
  INV_X1 U23234 ( .A(n23317), .ZN(n23316) );
  OR2_X1 U23235 ( .A1(n23318), .A2(n23319), .ZN(n23317) );
  AND2_X1 U23236 ( .A1(n23319), .A2(n23318), .ZN(n23315) );
  AND2_X1 U23237 ( .A1(n23320), .A2(n23321), .ZN(n23318) );
  OR2_X1 U23238 ( .A1(n23322), .A2(n23323), .ZN(n23321) );
  INV_X1 U23239 ( .A(n23324), .ZN(n23323) );
  OR2_X1 U23240 ( .A1(n23324), .A2(n23325), .ZN(n23320) );
  INV_X1 U23241 ( .A(n23322), .ZN(n23325) );
  OR2_X1 U23242 ( .A1(n22891), .A2(n22894), .ZN(n23246) );
  OR2_X1 U23243 ( .A1(n15072), .A2(n15320), .ZN(n22894) );
  OR2_X1 U23244 ( .A1(n23326), .A2(n23327), .ZN(n22891) );
  INV_X1 U23245 ( .A(n23328), .ZN(n23327) );
  OR2_X1 U23246 ( .A1(n23329), .A2(n23330), .ZN(n23328) );
  AND2_X1 U23247 ( .A1(n23330), .A2(n23329), .ZN(n23326) );
  AND2_X1 U23248 ( .A1(n23331), .A2(n23332), .ZN(n23329) );
  OR2_X1 U23249 ( .A1(n23333), .A2(n23334), .ZN(n23332) );
  INV_X1 U23250 ( .A(n23335), .ZN(n23334) );
  OR2_X1 U23251 ( .A1(n23335), .A2(n23336), .ZN(n23331) );
  INV_X1 U23252 ( .A(n23333), .ZN(n23336) );
  OR2_X1 U23253 ( .A1(n22902), .A2(n22905), .ZN(n23243) );
  OR2_X1 U23254 ( .A1(n15106), .A2(n15320), .ZN(n22905) );
  OR2_X1 U23255 ( .A1(n23337), .A2(n23338), .ZN(n22902) );
  INV_X1 U23256 ( .A(n23339), .ZN(n23338) );
  OR2_X1 U23257 ( .A1(n23340), .A2(n23341), .ZN(n23339) );
  AND2_X1 U23258 ( .A1(n23341), .A2(n23340), .ZN(n23337) );
  AND2_X1 U23259 ( .A1(n23342), .A2(n23343), .ZN(n23340) );
  OR2_X1 U23260 ( .A1(n23344), .A2(n23345), .ZN(n23343) );
  INV_X1 U23261 ( .A(n23346), .ZN(n23345) );
  OR2_X1 U23262 ( .A1(n23346), .A2(n23347), .ZN(n23342) );
  INV_X1 U23263 ( .A(n23344), .ZN(n23347) );
  OR2_X1 U23264 ( .A1(n22913), .A2(n22916), .ZN(n23240) );
  OR2_X1 U23265 ( .A1(n15140), .A2(n15320), .ZN(n22916) );
  OR2_X1 U23266 ( .A1(n23348), .A2(n23349), .ZN(n22913) );
  INV_X1 U23267 ( .A(n23350), .ZN(n23349) );
  OR2_X1 U23268 ( .A1(n23351), .A2(n23352), .ZN(n23350) );
  AND2_X1 U23269 ( .A1(n23352), .A2(n23351), .ZN(n23348) );
  AND2_X1 U23270 ( .A1(n23353), .A2(n23354), .ZN(n23351) );
  OR2_X1 U23271 ( .A1(n23355), .A2(n23356), .ZN(n23354) );
  INV_X1 U23272 ( .A(n23357), .ZN(n23356) );
  OR2_X1 U23273 ( .A1(n23357), .A2(n23358), .ZN(n23353) );
  INV_X1 U23274 ( .A(n23355), .ZN(n23358) );
  OR2_X1 U23275 ( .A1(n22924), .A2(n22927), .ZN(n23237) );
  OR2_X1 U23276 ( .A1(n15174), .A2(n15320), .ZN(n22927) );
  OR2_X1 U23277 ( .A1(n23359), .A2(n23360), .ZN(n22924) );
  INV_X1 U23278 ( .A(n23361), .ZN(n23360) );
  OR2_X1 U23279 ( .A1(n23362), .A2(n23363), .ZN(n23361) );
  AND2_X1 U23280 ( .A1(n23363), .A2(n23362), .ZN(n23359) );
  AND2_X1 U23281 ( .A1(n23364), .A2(n23365), .ZN(n23362) );
  OR2_X1 U23282 ( .A1(n23366), .A2(n23367), .ZN(n23365) );
  INV_X1 U23283 ( .A(n23368), .ZN(n23367) );
  OR2_X1 U23284 ( .A1(n23368), .A2(n23369), .ZN(n23364) );
  INV_X1 U23285 ( .A(n23366), .ZN(n23369) );
  OR2_X1 U23286 ( .A1(n22935), .A2(n22938), .ZN(n23234) );
  OR2_X1 U23287 ( .A1(n15208), .A2(n15320), .ZN(n22938) );
  OR2_X1 U23288 ( .A1(n23370), .A2(n23371), .ZN(n22935) );
  INV_X1 U23289 ( .A(n23372), .ZN(n23371) );
  OR2_X1 U23290 ( .A1(n23373), .A2(n23374), .ZN(n23372) );
  AND2_X1 U23291 ( .A1(n23374), .A2(n23373), .ZN(n23370) );
  AND2_X1 U23292 ( .A1(n23375), .A2(n23376), .ZN(n23373) );
  OR2_X1 U23293 ( .A1(n23377), .A2(n23378), .ZN(n23376) );
  INV_X1 U23294 ( .A(n23379), .ZN(n23378) );
  OR2_X1 U23295 ( .A1(n23379), .A2(n23380), .ZN(n23375) );
  INV_X1 U23296 ( .A(n23377), .ZN(n23380) );
  OR2_X1 U23297 ( .A1(n22946), .A2(n22949), .ZN(n23231) );
  OR2_X1 U23298 ( .A1(n15242), .A2(n15320), .ZN(n22949) );
  OR2_X1 U23299 ( .A1(n23381), .A2(n23382), .ZN(n22946) );
  INV_X1 U23300 ( .A(n23383), .ZN(n23382) );
  OR2_X1 U23301 ( .A1(n23384), .A2(n23385), .ZN(n23383) );
  AND2_X1 U23302 ( .A1(n23385), .A2(n23384), .ZN(n23381) );
  AND2_X1 U23303 ( .A1(n23386), .A2(n23387), .ZN(n23384) );
  OR2_X1 U23304 ( .A1(n23388), .A2(n23389), .ZN(n23387) );
  INV_X1 U23305 ( .A(n23390), .ZN(n23389) );
  OR2_X1 U23306 ( .A1(n23390), .A2(n23391), .ZN(n23386) );
  INV_X1 U23307 ( .A(n23388), .ZN(n23391) );
  OR2_X1 U23308 ( .A1(n22957), .A2(n22960), .ZN(n23228) );
  OR2_X1 U23309 ( .A1(n15287), .A2(n15320), .ZN(n22960) );
  OR2_X1 U23310 ( .A1(n23392), .A2(n23393), .ZN(n22957) );
  INV_X1 U23311 ( .A(n23394), .ZN(n23393) );
  OR2_X1 U23312 ( .A1(n23395), .A2(n23396), .ZN(n23394) );
  AND2_X1 U23313 ( .A1(n23396), .A2(n23395), .ZN(n23392) );
  AND2_X1 U23314 ( .A1(n23397), .A2(n23398), .ZN(n23395) );
  OR2_X1 U23315 ( .A1(n23399), .A2(n23400), .ZN(n23398) );
  INV_X1 U23316 ( .A(n23401), .ZN(n23400) );
  OR2_X1 U23317 ( .A1(n23401), .A2(n23402), .ZN(n23397) );
  INV_X1 U23318 ( .A(n23399), .ZN(n23402) );
  OR2_X1 U23319 ( .A1(n22968), .A2(n15915), .ZN(n23225) );
  OR2_X1 U23320 ( .A1(n15321), .A2(n15320), .ZN(n15915) );
  OR2_X1 U23321 ( .A1(n23403), .A2(n23404), .ZN(n22968) );
  INV_X1 U23322 ( .A(n23405), .ZN(n23404) );
  OR2_X1 U23323 ( .A1(n23406), .A2(n23407), .ZN(n23405) );
  AND2_X1 U23324 ( .A1(n23407), .A2(n23406), .ZN(n23403) );
  AND2_X1 U23325 ( .A1(n23408), .A2(n23409), .ZN(n23406) );
  OR2_X1 U23326 ( .A1(n23410), .A2(n23411), .ZN(n23409) );
  INV_X1 U23327 ( .A(n23412), .ZN(n23411) );
  OR2_X1 U23328 ( .A1(n23412), .A2(n23413), .ZN(n23408) );
  INV_X1 U23329 ( .A(n23410), .ZN(n23413) );
  OR2_X1 U23330 ( .A1(n22978), .A2(n22981), .ZN(n23222) );
  OR2_X1 U23331 ( .A1(n15355), .A2(n15320), .ZN(n22981) );
  OR2_X1 U23332 ( .A1(n23414), .A2(n23415), .ZN(n22978) );
  INV_X1 U23333 ( .A(n23416), .ZN(n23415) );
  OR2_X1 U23334 ( .A1(n23417), .A2(n23418), .ZN(n23416) );
  AND2_X1 U23335 ( .A1(n23418), .A2(n23417), .ZN(n23414) );
  AND2_X1 U23336 ( .A1(n23419), .A2(n23420), .ZN(n23417) );
  OR2_X1 U23337 ( .A1(n23421), .A2(n23422), .ZN(n23420) );
  INV_X1 U23338 ( .A(n23423), .ZN(n23422) );
  OR2_X1 U23339 ( .A1(n23423), .A2(n23424), .ZN(n23419) );
  INV_X1 U23340 ( .A(n23421), .ZN(n23424) );
  OR2_X1 U23341 ( .A1(n15389), .A2(n15320), .ZN(n22992) );
  OR2_X1 U23342 ( .A1(n23425), .A2(n23426), .ZN(n22989) );
  INV_X1 U23343 ( .A(n23427), .ZN(n23426) );
  OR2_X1 U23344 ( .A1(n23428), .A2(n23429), .ZN(n23427) );
  AND2_X1 U23345 ( .A1(n23429), .A2(n23428), .ZN(n23425) );
  AND2_X1 U23346 ( .A1(n23430), .A2(n23431), .ZN(n23428) );
  OR2_X1 U23347 ( .A1(n15912), .A2(n23432), .ZN(n23431) );
  INV_X1 U23348 ( .A(n23433), .ZN(n23432) );
  OR2_X1 U23349 ( .A1(n23433), .A2(n23434), .ZN(n23430) );
  INV_X1 U23350 ( .A(n15912), .ZN(n23434) );
  OR2_X1 U23351 ( .A1(n23000), .A2(n23006), .ZN(n23216) );
  OR2_X1 U23352 ( .A1(n15423), .A2(n15320), .ZN(n23006) );
  OR2_X1 U23353 ( .A1(n23435), .A2(n23436), .ZN(n23000) );
  INV_X1 U23354 ( .A(n23437), .ZN(n23436) );
  OR2_X1 U23355 ( .A1(n23438), .A2(n23439), .ZN(n23437) );
  AND2_X1 U23356 ( .A1(n23439), .A2(n23438), .ZN(n23435) );
  AND2_X1 U23357 ( .A1(n23440), .A2(n23441), .ZN(n23438) );
  INV_X1 U23358 ( .A(n23442), .ZN(n23441) );
  AND2_X1 U23359 ( .A1(n23443), .A2(n23444), .ZN(n23442) );
  OR2_X1 U23360 ( .A1(n23444), .A2(n23443), .ZN(n23440) );
  INV_X1 U23361 ( .A(n23445), .ZN(n23443) );
  OR2_X1 U23362 ( .A1(n15457), .A2(n15320), .ZN(n23016) );
  AND2_X1 U23363 ( .A1(n23446), .A2(n23447), .ZN(n23011) );
  INV_X1 U23364 ( .A(n23448), .ZN(n23447) );
  AND2_X1 U23365 ( .A1(n23449), .A2(n23450), .ZN(n23448) );
  OR2_X1 U23366 ( .A1(n23450), .A2(n23449), .ZN(n23446) );
  OR2_X1 U23367 ( .A1(n23451), .A2(n23452), .ZN(n23449) );
  AND2_X1 U23368 ( .A1(n23453), .A2(n23454), .ZN(n23452) );
  INV_X1 U23369 ( .A(n23455), .ZN(n23453) );
  AND2_X1 U23370 ( .A1(n23456), .A2(n23455), .ZN(n23451) );
  INV_X1 U23371 ( .A(n23454), .ZN(n23456) );
  OR2_X1 U23372 ( .A1(n15491), .A2(n15320), .ZN(n23027) );
  AND2_X1 U23373 ( .A1(n23457), .A2(n23458), .ZN(n23022) );
  INV_X1 U23374 ( .A(n23459), .ZN(n23458) );
  AND2_X1 U23375 ( .A1(n23460), .A2(n23461), .ZN(n23459) );
  OR2_X1 U23376 ( .A1(n23461), .A2(n23460), .ZN(n23457) );
  OR2_X1 U23377 ( .A1(n23462), .A2(n23463), .ZN(n23460) );
  AND2_X1 U23378 ( .A1(n23464), .A2(n23465), .ZN(n23463) );
  INV_X1 U23379 ( .A(n23466), .ZN(n23464) );
  AND2_X1 U23380 ( .A1(n23467), .A2(n23466), .ZN(n23462) );
  INV_X1 U23381 ( .A(n23465), .ZN(n23467) );
  OR2_X1 U23382 ( .A1(n15525), .A2(n15320), .ZN(n23038) );
  AND2_X1 U23383 ( .A1(n23468), .A2(n23469), .ZN(n23033) );
  INV_X1 U23384 ( .A(n23470), .ZN(n23469) );
  AND2_X1 U23385 ( .A1(n23471), .A2(n23472), .ZN(n23470) );
  OR2_X1 U23386 ( .A1(n23472), .A2(n23471), .ZN(n23468) );
  OR2_X1 U23387 ( .A1(n23473), .A2(n23474), .ZN(n23471) );
  AND2_X1 U23388 ( .A1(n23475), .A2(n23476), .ZN(n23474) );
  INV_X1 U23389 ( .A(n23477), .ZN(n23475) );
  AND2_X1 U23390 ( .A1(n23478), .A2(n23477), .ZN(n23473) );
  INV_X1 U23391 ( .A(n23476), .ZN(n23478) );
  OR2_X1 U23392 ( .A1(n15559), .A2(n15320), .ZN(n23049) );
  AND2_X1 U23393 ( .A1(n23479), .A2(n23480), .ZN(n23044) );
  INV_X1 U23394 ( .A(n23481), .ZN(n23480) );
  AND2_X1 U23395 ( .A1(n23482), .A2(n23483), .ZN(n23481) );
  OR2_X1 U23396 ( .A1(n23483), .A2(n23482), .ZN(n23479) );
  OR2_X1 U23397 ( .A1(n23484), .A2(n23485), .ZN(n23482) );
  AND2_X1 U23398 ( .A1(n23486), .A2(n23487), .ZN(n23485) );
  INV_X1 U23399 ( .A(n23488), .ZN(n23486) );
  AND2_X1 U23400 ( .A1(n23489), .A2(n23488), .ZN(n23484) );
  INV_X1 U23401 ( .A(n23487), .ZN(n23489) );
  OR2_X1 U23402 ( .A1(n15593), .A2(n15320), .ZN(n23060) );
  AND2_X1 U23403 ( .A1(n23490), .A2(n23491), .ZN(n23055) );
  INV_X1 U23404 ( .A(n23492), .ZN(n23491) );
  AND2_X1 U23405 ( .A1(n23493), .A2(n23494), .ZN(n23492) );
  OR2_X1 U23406 ( .A1(n23494), .A2(n23493), .ZN(n23490) );
  OR2_X1 U23407 ( .A1(n23495), .A2(n23496), .ZN(n23493) );
  AND2_X1 U23408 ( .A1(n23497), .A2(n23498), .ZN(n23496) );
  INV_X1 U23409 ( .A(n23499), .ZN(n23497) );
  AND2_X1 U23410 ( .A1(n23500), .A2(n23499), .ZN(n23495) );
  INV_X1 U23411 ( .A(n23498), .ZN(n23500) );
  OR2_X1 U23412 ( .A1(n15638), .A2(n15320), .ZN(n23071) );
  AND2_X1 U23413 ( .A1(n23501), .A2(n23502), .ZN(n23066) );
  INV_X1 U23414 ( .A(n23503), .ZN(n23502) );
  AND2_X1 U23415 ( .A1(n23504), .A2(n23505), .ZN(n23503) );
  OR2_X1 U23416 ( .A1(n23505), .A2(n23504), .ZN(n23501) );
  OR2_X1 U23417 ( .A1(n23506), .A2(n23507), .ZN(n23504) );
  AND2_X1 U23418 ( .A1(n23508), .A2(n23509), .ZN(n23507) );
  INV_X1 U23419 ( .A(n23510), .ZN(n23508) );
  AND2_X1 U23420 ( .A1(n23511), .A2(n23510), .ZN(n23506) );
  INV_X1 U23421 ( .A(n23509), .ZN(n23511) );
  OR2_X1 U23422 ( .A1(n15672), .A2(n15320), .ZN(n23082) );
  AND2_X1 U23423 ( .A1(n23512), .A2(n23513), .ZN(n23077) );
  INV_X1 U23424 ( .A(n23514), .ZN(n23513) );
  AND2_X1 U23425 ( .A1(n23515), .A2(n23516), .ZN(n23514) );
  OR2_X1 U23426 ( .A1(n23516), .A2(n23515), .ZN(n23512) );
  OR2_X1 U23427 ( .A1(n23517), .A2(n23518), .ZN(n23515) );
  AND2_X1 U23428 ( .A1(n23519), .A2(n23520), .ZN(n23518) );
  INV_X1 U23429 ( .A(n23521), .ZN(n23519) );
  AND2_X1 U23430 ( .A1(n23522), .A2(n23521), .ZN(n23517) );
  INV_X1 U23431 ( .A(n23520), .ZN(n23522) );
  OR2_X1 U23432 ( .A1(n15706), .A2(n15320), .ZN(n23093) );
  AND2_X1 U23433 ( .A1(n23523), .A2(n23524), .ZN(n23088) );
  INV_X1 U23434 ( .A(n23525), .ZN(n23524) );
  AND2_X1 U23435 ( .A1(n23526), .A2(n23527), .ZN(n23525) );
  OR2_X1 U23436 ( .A1(n23527), .A2(n23526), .ZN(n23523) );
  OR2_X1 U23437 ( .A1(n23528), .A2(n23529), .ZN(n23526) );
  AND2_X1 U23438 ( .A1(n23530), .A2(n23531), .ZN(n23529) );
  INV_X1 U23439 ( .A(n23532), .ZN(n23530) );
  AND2_X1 U23440 ( .A1(n23533), .A2(n23532), .ZN(n23528) );
  INV_X1 U23441 ( .A(n23531), .ZN(n23533) );
  OR2_X1 U23442 ( .A1(n15740), .A2(n15320), .ZN(n23104) );
  AND2_X1 U23443 ( .A1(n23534), .A2(n23535), .ZN(n23099) );
  INV_X1 U23444 ( .A(n23536), .ZN(n23535) );
  AND2_X1 U23445 ( .A1(n23537), .A2(n23538), .ZN(n23536) );
  OR2_X1 U23446 ( .A1(n23538), .A2(n23537), .ZN(n23534) );
  OR2_X1 U23447 ( .A1(n23539), .A2(n23540), .ZN(n23537) );
  AND2_X1 U23448 ( .A1(n23541), .A2(n23542), .ZN(n23540) );
  INV_X1 U23449 ( .A(n23543), .ZN(n23541) );
  AND2_X1 U23450 ( .A1(n23544), .A2(n23543), .ZN(n23539) );
  INV_X1 U23451 ( .A(n23542), .ZN(n23544) );
  OR2_X1 U23452 ( .A1(n15774), .A2(n15320), .ZN(n23115) );
  AND2_X1 U23453 ( .A1(n23545), .A2(n23546), .ZN(n23110) );
  INV_X1 U23454 ( .A(n23547), .ZN(n23546) );
  AND2_X1 U23455 ( .A1(n23548), .A2(n23549), .ZN(n23547) );
  OR2_X1 U23456 ( .A1(n23549), .A2(n23548), .ZN(n23545) );
  OR2_X1 U23457 ( .A1(n23550), .A2(n23551), .ZN(n23548) );
  AND2_X1 U23458 ( .A1(n23552), .A2(n23553), .ZN(n23551) );
  INV_X1 U23459 ( .A(n23554), .ZN(n23552) );
  AND2_X1 U23460 ( .A1(n23555), .A2(n23554), .ZN(n23550) );
  INV_X1 U23461 ( .A(n23553), .ZN(n23555) );
  OR2_X1 U23462 ( .A1(n15808), .A2(n15320), .ZN(n23126) );
  AND2_X1 U23463 ( .A1(n23556), .A2(n23557), .ZN(n23121) );
  INV_X1 U23464 ( .A(n23558), .ZN(n23557) );
  AND2_X1 U23465 ( .A1(n23559), .A2(n23560), .ZN(n23558) );
  OR2_X1 U23466 ( .A1(n23560), .A2(n23559), .ZN(n23556) );
  OR2_X1 U23467 ( .A1(n23561), .A2(n23562), .ZN(n23559) );
  AND2_X1 U23468 ( .A1(n23563), .A2(n23564), .ZN(n23562) );
  INV_X1 U23469 ( .A(n23565), .ZN(n23563) );
  AND2_X1 U23470 ( .A1(n23566), .A2(n23565), .ZN(n23561) );
  INV_X1 U23471 ( .A(n23564), .ZN(n23566) );
  OR2_X1 U23472 ( .A1(n15842), .A2(n15320), .ZN(n23137) );
  AND2_X1 U23473 ( .A1(n23567), .A2(n23568), .ZN(n23132) );
  INV_X1 U23474 ( .A(n23569), .ZN(n23568) );
  AND2_X1 U23475 ( .A1(n23570), .A2(n23571), .ZN(n23569) );
  OR2_X1 U23476 ( .A1(n23571), .A2(n23570), .ZN(n23567) );
  OR2_X1 U23477 ( .A1(n23572), .A2(n23573), .ZN(n23570) );
  AND2_X1 U23478 ( .A1(n23574), .A2(n23575), .ZN(n23573) );
  INV_X1 U23479 ( .A(n23576), .ZN(n23574) );
  AND2_X1 U23480 ( .A1(n23577), .A2(n23576), .ZN(n23572) );
  INV_X1 U23481 ( .A(n23575), .ZN(n23577) );
  OR2_X1 U23482 ( .A1(n16512), .A2(n15320), .ZN(n23148) );
  INV_X1 U23483 ( .A(b_16_), .ZN(n15320) );
  AND2_X1 U23484 ( .A1(n23578), .A2(n23579), .ZN(n23143) );
  INV_X1 U23485 ( .A(n23580), .ZN(n23579) );
  AND2_X1 U23486 ( .A1(n23581), .A2(n23582), .ZN(n23580) );
  OR2_X1 U23487 ( .A1(n23582), .A2(n23581), .ZN(n23578) );
  OR2_X1 U23488 ( .A1(n23583), .A2(n23584), .ZN(n23581) );
  AND2_X1 U23489 ( .A1(n23585), .A2(n23586), .ZN(n23584) );
  INV_X1 U23490 ( .A(n23587), .ZN(n23585) );
  AND2_X1 U23491 ( .A1(n23588), .A2(n23587), .ZN(n23583) );
  INV_X1 U23492 ( .A(n23586), .ZN(n23588) );
  AND2_X1 U23493 ( .A1(n23589), .A2(n23590), .ZN(n23152) );
  INV_X1 U23494 ( .A(n23591), .ZN(n23590) );
  AND2_X1 U23495 ( .A1(n23592), .A2(n23162), .ZN(n23591) );
  OR2_X1 U23496 ( .A1(n23162), .A2(n23592), .ZN(n23589) );
  OR2_X1 U23497 ( .A1(n23593), .A2(n23594), .ZN(n23592) );
  AND2_X1 U23498 ( .A1(n23595), .A2(n23161), .ZN(n23594) );
  INV_X1 U23499 ( .A(n23160), .ZN(n23595) );
  AND2_X1 U23500 ( .A1(n23596), .A2(n23160), .ZN(n23593) );
  OR2_X1 U23501 ( .A1(n16512), .A2(n15354), .ZN(n23160) );
  INV_X1 U23502 ( .A(n23161), .ZN(n23596) );
  OR2_X1 U23503 ( .A1(n23597), .A2(n23598), .ZN(n23161) );
  AND2_X1 U23504 ( .A1(n23587), .A2(n23586), .ZN(n23598) );
  AND2_X1 U23505 ( .A1(n23582), .A2(n23599), .ZN(n23597) );
  OR2_X1 U23506 ( .A1(n23587), .A2(n23586), .ZN(n23599) );
  OR2_X1 U23507 ( .A1(n23600), .A2(n23601), .ZN(n23586) );
  AND2_X1 U23508 ( .A1(n23576), .A2(n23575), .ZN(n23601) );
  AND2_X1 U23509 ( .A1(n23571), .A2(n23602), .ZN(n23600) );
  OR2_X1 U23510 ( .A1(n23576), .A2(n23575), .ZN(n23602) );
  OR2_X1 U23511 ( .A1(n23603), .A2(n23604), .ZN(n23575) );
  AND2_X1 U23512 ( .A1(n23565), .A2(n23564), .ZN(n23604) );
  AND2_X1 U23513 ( .A1(n23560), .A2(n23605), .ZN(n23603) );
  OR2_X1 U23514 ( .A1(n23565), .A2(n23564), .ZN(n23605) );
  OR2_X1 U23515 ( .A1(n23606), .A2(n23607), .ZN(n23564) );
  AND2_X1 U23516 ( .A1(n23554), .A2(n23553), .ZN(n23607) );
  AND2_X1 U23517 ( .A1(n23549), .A2(n23608), .ZN(n23606) );
  OR2_X1 U23518 ( .A1(n23554), .A2(n23553), .ZN(n23608) );
  OR2_X1 U23519 ( .A1(n23609), .A2(n23610), .ZN(n23553) );
  AND2_X1 U23520 ( .A1(n23543), .A2(n23542), .ZN(n23610) );
  AND2_X1 U23521 ( .A1(n23538), .A2(n23611), .ZN(n23609) );
  OR2_X1 U23522 ( .A1(n23543), .A2(n23542), .ZN(n23611) );
  OR2_X1 U23523 ( .A1(n23612), .A2(n23613), .ZN(n23542) );
  AND2_X1 U23524 ( .A1(n23532), .A2(n23531), .ZN(n23613) );
  AND2_X1 U23525 ( .A1(n23527), .A2(n23614), .ZN(n23612) );
  OR2_X1 U23526 ( .A1(n23532), .A2(n23531), .ZN(n23614) );
  OR2_X1 U23527 ( .A1(n23615), .A2(n23616), .ZN(n23531) );
  AND2_X1 U23528 ( .A1(n23521), .A2(n23520), .ZN(n23616) );
  AND2_X1 U23529 ( .A1(n23516), .A2(n23617), .ZN(n23615) );
  OR2_X1 U23530 ( .A1(n23521), .A2(n23520), .ZN(n23617) );
  OR2_X1 U23531 ( .A1(n23618), .A2(n23619), .ZN(n23520) );
  AND2_X1 U23532 ( .A1(n23510), .A2(n23509), .ZN(n23619) );
  AND2_X1 U23533 ( .A1(n23505), .A2(n23620), .ZN(n23618) );
  OR2_X1 U23534 ( .A1(n23510), .A2(n23509), .ZN(n23620) );
  OR2_X1 U23535 ( .A1(n23621), .A2(n23622), .ZN(n23509) );
  AND2_X1 U23536 ( .A1(n23499), .A2(n23498), .ZN(n23622) );
  AND2_X1 U23537 ( .A1(n23494), .A2(n23623), .ZN(n23621) );
  OR2_X1 U23538 ( .A1(n23499), .A2(n23498), .ZN(n23623) );
  OR2_X1 U23539 ( .A1(n23624), .A2(n23625), .ZN(n23498) );
  AND2_X1 U23540 ( .A1(n23488), .A2(n23487), .ZN(n23625) );
  AND2_X1 U23541 ( .A1(n23483), .A2(n23626), .ZN(n23624) );
  OR2_X1 U23542 ( .A1(n23488), .A2(n23487), .ZN(n23626) );
  OR2_X1 U23543 ( .A1(n23627), .A2(n23628), .ZN(n23487) );
  AND2_X1 U23544 ( .A1(n23477), .A2(n23476), .ZN(n23628) );
  AND2_X1 U23545 ( .A1(n23472), .A2(n23629), .ZN(n23627) );
  OR2_X1 U23546 ( .A1(n23477), .A2(n23476), .ZN(n23629) );
  OR2_X1 U23547 ( .A1(n23630), .A2(n23631), .ZN(n23476) );
  AND2_X1 U23548 ( .A1(n23466), .A2(n23465), .ZN(n23631) );
  AND2_X1 U23549 ( .A1(n23461), .A2(n23632), .ZN(n23630) );
  OR2_X1 U23550 ( .A1(n23466), .A2(n23465), .ZN(n23632) );
  OR2_X1 U23551 ( .A1(n23633), .A2(n23634), .ZN(n23465) );
  AND2_X1 U23552 ( .A1(n23455), .A2(n23454), .ZN(n23634) );
  AND2_X1 U23553 ( .A1(n23450), .A2(n23635), .ZN(n23633) );
  OR2_X1 U23554 ( .A1(n23455), .A2(n23454), .ZN(n23635) );
  OR2_X1 U23555 ( .A1(n23636), .A2(n23637), .ZN(n23454) );
  AND2_X1 U23556 ( .A1(n23445), .A2(n23444), .ZN(n23637) );
  AND2_X1 U23557 ( .A1(n23439), .A2(n23638), .ZN(n23636) );
  OR2_X1 U23558 ( .A1(n23445), .A2(n23444), .ZN(n23638) );
  OR2_X1 U23559 ( .A1(n23639), .A2(n23640), .ZN(n23444) );
  AND2_X1 U23560 ( .A1(n15912), .A2(n23433), .ZN(n23640) );
  AND2_X1 U23561 ( .A1(n23429), .A2(n23641), .ZN(n23639) );
  OR2_X1 U23562 ( .A1(n15912), .A2(n23433), .ZN(n23641) );
  OR2_X1 U23563 ( .A1(n23642), .A2(n23643), .ZN(n23433) );
  AND2_X1 U23564 ( .A1(n23421), .A2(n23423), .ZN(n23643) );
  AND2_X1 U23565 ( .A1(n23418), .A2(n23644), .ZN(n23642) );
  OR2_X1 U23566 ( .A1(n23421), .A2(n23423), .ZN(n23644) );
  OR2_X1 U23567 ( .A1(n23645), .A2(n23646), .ZN(n23423) );
  AND2_X1 U23568 ( .A1(n23410), .A2(n23412), .ZN(n23646) );
  AND2_X1 U23569 ( .A1(n23407), .A2(n23647), .ZN(n23645) );
  OR2_X1 U23570 ( .A1(n23410), .A2(n23412), .ZN(n23647) );
  OR2_X1 U23571 ( .A1(n23648), .A2(n23649), .ZN(n23412) );
  AND2_X1 U23572 ( .A1(n23399), .A2(n23401), .ZN(n23649) );
  AND2_X1 U23573 ( .A1(n23396), .A2(n23650), .ZN(n23648) );
  OR2_X1 U23574 ( .A1(n23399), .A2(n23401), .ZN(n23650) );
  OR2_X1 U23575 ( .A1(n23651), .A2(n23652), .ZN(n23401) );
  AND2_X1 U23576 ( .A1(n23388), .A2(n23390), .ZN(n23652) );
  AND2_X1 U23577 ( .A1(n23385), .A2(n23653), .ZN(n23651) );
  OR2_X1 U23578 ( .A1(n23388), .A2(n23390), .ZN(n23653) );
  OR2_X1 U23579 ( .A1(n23654), .A2(n23655), .ZN(n23390) );
  AND2_X1 U23580 ( .A1(n23377), .A2(n23379), .ZN(n23655) );
  AND2_X1 U23581 ( .A1(n23374), .A2(n23656), .ZN(n23654) );
  OR2_X1 U23582 ( .A1(n23377), .A2(n23379), .ZN(n23656) );
  OR2_X1 U23583 ( .A1(n23657), .A2(n23658), .ZN(n23379) );
  AND2_X1 U23584 ( .A1(n23366), .A2(n23368), .ZN(n23658) );
  AND2_X1 U23585 ( .A1(n23363), .A2(n23659), .ZN(n23657) );
  OR2_X1 U23586 ( .A1(n23366), .A2(n23368), .ZN(n23659) );
  OR2_X1 U23587 ( .A1(n23660), .A2(n23661), .ZN(n23368) );
  AND2_X1 U23588 ( .A1(n23355), .A2(n23357), .ZN(n23661) );
  AND2_X1 U23589 ( .A1(n23352), .A2(n23662), .ZN(n23660) );
  OR2_X1 U23590 ( .A1(n23355), .A2(n23357), .ZN(n23662) );
  OR2_X1 U23591 ( .A1(n23663), .A2(n23664), .ZN(n23357) );
  AND2_X1 U23592 ( .A1(n23344), .A2(n23346), .ZN(n23664) );
  AND2_X1 U23593 ( .A1(n23341), .A2(n23665), .ZN(n23663) );
  OR2_X1 U23594 ( .A1(n23344), .A2(n23346), .ZN(n23665) );
  OR2_X1 U23595 ( .A1(n23666), .A2(n23667), .ZN(n23346) );
  AND2_X1 U23596 ( .A1(n23333), .A2(n23335), .ZN(n23667) );
  AND2_X1 U23597 ( .A1(n23330), .A2(n23668), .ZN(n23666) );
  OR2_X1 U23598 ( .A1(n23333), .A2(n23335), .ZN(n23668) );
  OR2_X1 U23599 ( .A1(n23669), .A2(n23670), .ZN(n23335) );
  AND2_X1 U23600 ( .A1(n23322), .A2(n23324), .ZN(n23670) );
  AND2_X1 U23601 ( .A1(n23319), .A2(n23671), .ZN(n23669) );
  OR2_X1 U23602 ( .A1(n23322), .A2(n23324), .ZN(n23671) );
  OR2_X1 U23603 ( .A1(n23672), .A2(n23673), .ZN(n23324) );
  AND2_X1 U23604 ( .A1(n23311), .A2(n23313), .ZN(n23673) );
  AND2_X1 U23605 ( .A1(n23308), .A2(n23674), .ZN(n23672) );
  OR2_X1 U23606 ( .A1(n23311), .A2(n23313), .ZN(n23674) );
  OR2_X1 U23607 ( .A1(n23675), .A2(n23676), .ZN(n23313) );
  AND2_X1 U23608 ( .A1(n23300), .A2(n23302), .ZN(n23676) );
  AND2_X1 U23609 ( .A1(n23297), .A2(n23677), .ZN(n23675) );
  OR2_X1 U23610 ( .A1(n23300), .A2(n23302), .ZN(n23677) );
  OR2_X1 U23611 ( .A1(n23678), .A2(n23679), .ZN(n23302) );
  AND2_X1 U23612 ( .A1(n23289), .A2(n23291), .ZN(n23679) );
  AND2_X1 U23613 ( .A1(n23286), .A2(n23680), .ZN(n23678) );
  OR2_X1 U23614 ( .A1(n23289), .A2(n23291), .ZN(n23680) );
  OR2_X1 U23615 ( .A1(n23681), .A2(n23682), .ZN(n23291) );
  AND2_X1 U23616 ( .A1(n23274), .A2(n23279), .ZN(n23682) );
  AND2_X1 U23617 ( .A1(n23278), .A2(n23683), .ZN(n23681) );
  OR2_X1 U23618 ( .A1(n23274), .A2(n23279), .ZN(n23683) );
  INV_X1 U23619 ( .A(n23280), .ZN(n23279) );
  AND3_X1 U23620 ( .A1(b_15_), .A2(b_14_), .A3(n15957), .ZN(n23280) );
  OR2_X1 U23621 ( .A1(n14857), .A2(n15354), .ZN(n23274) );
  INV_X1 U23622 ( .A(n23281), .ZN(n23278) );
  OR2_X1 U23623 ( .A1(n23684), .A2(n23685), .ZN(n23281) );
  AND2_X1 U23624 ( .A1(b_14_), .A2(n23686), .ZN(n23685) );
  OR2_X1 U23625 ( .A1(n23687), .A2(n16981), .ZN(n23686) );
  AND2_X1 U23626 ( .A1(a_30_), .A2(n15422), .ZN(n23687) );
  AND2_X1 U23627 ( .A1(b_13_), .A2(n23688), .ZN(n23684) );
  OR2_X1 U23628 ( .A1(n23689), .A2(n14817), .ZN(n23688) );
  AND2_X1 U23629 ( .A1(a_31_), .A2(n15388), .ZN(n23689) );
  OR2_X1 U23630 ( .A1(n14891), .A2(n15354), .ZN(n23289) );
  OR2_X1 U23631 ( .A1(n23690), .A2(n23691), .ZN(n23286) );
  AND2_X1 U23632 ( .A1(n23692), .A2(n23693), .ZN(n23691) );
  INV_X1 U23633 ( .A(n23694), .ZN(n23690) );
  OR2_X1 U23634 ( .A1(n23692), .A2(n23693), .ZN(n23694) );
  OR2_X1 U23635 ( .A1(n23695), .A2(n23696), .ZN(n23692) );
  AND2_X1 U23636 ( .A1(n23697), .A2(n23698), .ZN(n23696) );
  AND2_X1 U23637 ( .A1(n23699), .A2(n23700), .ZN(n23695) );
  OR2_X1 U23638 ( .A1(n14936), .A2(n15354), .ZN(n23300) );
  OR2_X1 U23639 ( .A1(n23701), .A2(n23702), .ZN(n23297) );
  INV_X1 U23640 ( .A(n23703), .ZN(n23702) );
  OR2_X1 U23641 ( .A1(n23704), .A2(n23705), .ZN(n23703) );
  AND2_X1 U23642 ( .A1(n23705), .A2(n23704), .ZN(n23701) );
  AND2_X1 U23643 ( .A1(n23706), .A2(n23707), .ZN(n23704) );
  OR2_X1 U23644 ( .A1(n23708), .A2(n23709), .ZN(n23707) );
  INV_X1 U23645 ( .A(n23710), .ZN(n23709) );
  OR2_X1 U23646 ( .A1(n23710), .A2(n23711), .ZN(n23706) );
  INV_X1 U23647 ( .A(n23708), .ZN(n23711) );
  OR2_X1 U23648 ( .A1(n14970), .A2(n15354), .ZN(n23311) );
  OR2_X1 U23649 ( .A1(n23712), .A2(n23713), .ZN(n23308) );
  INV_X1 U23650 ( .A(n23714), .ZN(n23713) );
  OR2_X1 U23651 ( .A1(n23715), .A2(n23716), .ZN(n23714) );
  AND2_X1 U23652 ( .A1(n23716), .A2(n23715), .ZN(n23712) );
  AND2_X1 U23653 ( .A1(n23717), .A2(n23718), .ZN(n23715) );
  OR2_X1 U23654 ( .A1(n23719), .A2(n23720), .ZN(n23718) );
  INV_X1 U23655 ( .A(n23721), .ZN(n23720) );
  OR2_X1 U23656 ( .A1(n23721), .A2(n23722), .ZN(n23717) );
  INV_X1 U23657 ( .A(n23719), .ZN(n23722) );
  OR2_X1 U23658 ( .A1(n15004), .A2(n15354), .ZN(n23322) );
  OR2_X1 U23659 ( .A1(n23723), .A2(n23724), .ZN(n23319) );
  INV_X1 U23660 ( .A(n23725), .ZN(n23724) );
  OR2_X1 U23661 ( .A1(n23726), .A2(n23727), .ZN(n23725) );
  AND2_X1 U23662 ( .A1(n23727), .A2(n23726), .ZN(n23723) );
  AND2_X1 U23663 ( .A1(n23728), .A2(n23729), .ZN(n23726) );
  OR2_X1 U23664 ( .A1(n23730), .A2(n23731), .ZN(n23729) );
  INV_X1 U23665 ( .A(n23732), .ZN(n23731) );
  OR2_X1 U23666 ( .A1(n23732), .A2(n23733), .ZN(n23728) );
  INV_X1 U23667 ( .A(n23730), .ZN(n23733) );
  OR2_X1 U23668 ( .A1(n15038), .A2(n15354), .ZN(n23333) );
  OR2_X1 U23669 ( .A1(n23734), .A2(n23735), .ZN(n23330) );
  INV_X1 U23670 ( .A(n23736), .ZN(n23735) );
  OR2_X1 U23671 ( .A1(n23737), .A2(n23738), .ZN(n23736) );
  AND2_X1 U23672 ( .A1(n23738), .A2(n23737), .ZN(n23734) );
  AND2_X1 U23673 ( .A1(n23739), .A2(n23740), .ZN(n23737) );
  OR2_X1 U23674 ( .A1(n23741), .A2(n23742), .ZN(n23740) );
  INV_X1 U23675 ( .A(n23743), .ZN(n23742) );
  OR2_X1 U23676 ( .A1(n23743), .A2(n23744), .ZN(n23739) );
  INV_X1 U23677 ( .A(n23741), .ZN(n23744) );
  OR2_X1 U23678 ( .A1(n15072), .A2(n15354), .ZN(n23344) );
  OR2_X1 U23679 ( .A1(n23745), .A2(n23746), .ZN(n23341) );
  INV_X1 U23680 ( .A(n23747), .ZN(n23746) );
  OR2_X1 U23681 ( .A1(n23748), .A2(n23749), .ZN(n23747) );
  AND2_X1 U23682 ( .A1(n23749), .A2(n23748), .ZN(n23745) );
  AND2_X1 U23683 ( .A1(n23750), .A2(n23751), .ZN(n23748) );
  OR2_X1 U23684 ( .A1(n23752), .A2(n23753), .ZN(n23751) );
  INV_X1 U23685 ( .A(n23754), .ZN(n23753) );
  OR2_X1 U23686 ( .A1(n23754), .A2(n23755), .ZN(n23750) );
  INV_X1 U23687 ( .A(n23752), .ZN(n23755) );
  OR2_X1 U23688 ( .A1(n15106), .A2(n15354), .ZN(n23355) );
  OR2_X1 U23689 ( .A1(n23756), .A2(n23757), .ZN(n23352) );
  INV_X1 U23690 ( .A(n23758), .ZN(n23757) );
  OR2_X1 U23691 ( .A1(n23759), .A2(n23760), .ZN(n23758) );
  AND2_X1 U23692 ( .A1(n23760), .A2(n23759), .ZN(n23756) );
  AND2_X1 U23693 ( .A1(n23761), .A2(n23762), .ZN(n23759) );
  OR2_X1 U23694 ( .A1(n23763), .A2(n23764), .ZN(n23762) );
  INV_X1 U23695 ( .A(n23765), .ZN(n23764) );
  OR2_X1 U23696 ( .A1(n23765), .A2(n23766), .ZN(n23761) );
  INV_X1 U23697 ( .A(n23763), .ZN(n23766) );
  OR2_X1 U23698 ( .A1(n15140), .A2(n15354), .ZN(n23366) );
  OR2_X1 U23699 ( .A1(n23767), .A2(n23768), .ZN(n23363) );
  INV_X1 U23700 ( .A(n23769), .ZN(n23768) );
  OR2_X1 U23701 ( .A1(n23770), .A2(n23771), .ZN(n23769) );
  AND2_X1 U23702 ( .A1(n23771), .A2(n23770), .ZN(n23767) );
  AND2_X1 U23703 ( .A1(n23772), .A2(n23773), .ZN(n23770) );
  OR2_X1 U23704 ( .A1(n23774), .A2(n23775), .ZN(n23773) );
  INV_X1 U23705 ( .A(n23776), .ZN(n23775) );
  OR2_X1 U23706 ( .A1(n23776), .A2(n23777), .ZN(n23772) );
  INV_X1 U23707 ( .A(n23774), .ZN(n23777) );
  OR2_X1 U23708 ( .A1(n15174), .A2(n15354), .ZN(n23377) );
  OR2_X1 U23709 ( .A1(n23778), .A2(n23779), .ZN(n23374) );
  INV_X1 U23710 ( .A(n23780), .ZN(n23779) );
  OR2_X1 U23711 ( .A1(n23781), .A2(n23782), .ZN(n23780) );
  AND2_X1 U23712 ( .A1(n23782), .A2(n23781), .ZN(n23778) );
  AND2_X1 U23713 ( .A1(n23783), .A2(n23784), .ZN(n23781) );
  OR2_X1 U23714 ( .A1(n23785), .A2(n23786), .ZN(n23784) );
  INV_X1 U23715 ( .A(n23787), .ZN(n23786) );
  OR2_X1 U23716 ( .A1(n23787), .A2(n23788), .ZN(n23783) );
  INV_X1 U23717 ( .A(n23785), .ZN(n23788) );
  OR2_X1 U23718 ( .A1(n15208), .A2(n15354), .ZN(n23388) );
  OR2_X1 U23719 ( .A1(n23789), .A2(n23790), .ZN(n23385) );
  INV_X1 U23720 ( .A(n23791), .ZN(n23790) );
  OR2_X1 U23721 ( .A1(n23792), .A2(n23793), .ZN(n23791) );
  AND2_X1 U23722 ( .A1(n23793), .A2(n23792), .ZN(n23789) );
  AND2_X1 U23723 ( .A1(n23794), .A2(n23795), .ZN(n23792) );
  OR2_X1 U23724 ( .A1(n23796), .A2(n23797), .ZN(n23795) );
  INV_X1 U23725 ( .A(n23798), .ZN(n23797) );
  OR2_X1 U23726 ( .A1(n23798), .A2(n23799), .ZN(n23794) );
  INV_X1 U23727 ( .A(n23796), .ZN(n23799) );
  OR2_X1 U23728 ( .A1(n15242), .A2(n15354), .ZN(n23399) );
  OR2_X1 U23729 ( .A1(n23800), .A2(n23801), .ZN(n23396) );
  INV_X1 U23730 ( .A(n23802), .ZN(n23801) );
  OR2_X1 U23731 ( .A1(n23803), .A2(n23804), .ZN(n23802) );
  AND2_X1 U23732 ( .A1(n23804), .A2(n23803), .ZN(n23800) );
  AND2_X1 U23733 ( .A1(n23805), .A2(n23806), .ZN(n23803) );
  OR2_X1 U23734 ( .A1(n23807), .A2(n23808), .ZN(n23806) );
  INV_X1 U23735 ( .A(n23809), .ZN(n23808) );
  OR2_X1 U23736 ( .A1(n23809), .A2(n23810), .ZN(n23805) );
  INV_X1 U23737 ( .A(n23807), .ZN(n23810) );
  OR2_X1 U23738 ( .A1(n15287), .A2(n15354), .ZN(n23410) );
  OR2_X1 U23739 ( .A1(n23811), .A2(n23812), .ZN(n23407) );
  INV_X1 U23740 ( .A(n23813), .ZN(n23812) );
  OR2_X1 U23741 ( .A1(n23814), .A2(n23815), .ZN(n23813) );
  AND2_X1 U23742 ( .A1(n23815), .A2(n23814), .ZN(n23811) );
  AND2_X1 U23743 ( .A1(n23816), .A2(n23817), .ZN(n23814) );
  OR2_X1 U23744 ( .A1(n23818), .A2(n23819), .ZN(n23817) );
  INV_X1 U23745 ( .A(n23820), .ZN(n23819) );
  OR2_X1 U23746 ( .A1(n23820), .A2(n23821), .ZN(n23816) );
  INV_X1 U23747 ( .A(n23818), .ZN(n23821) );
  OR2_X1 U23748 ( .A1(n15321), .A2(n15354), .ZN(n23421) );
  OR2_X1 U23749 ( .A1(n23822), .A2(n23823), .ZN(n23418) );
  INV_X1 U23750 ( .A(n23824), .ZN(n23823) );
  OR2_X1 U23751 ( .A1(n23825), .A2(n23826), .ZN(n23824) );
  AND2_X1 U23752 ( .A1(n23826), .A2(n23825), .ZN(n23822) );
  AND2_X1 U23753 ( .A1(n23827), .A2(n23828), .ZN(n23825) );
  OR2_X1 U23754 ( .A1(n23829), .A2(n23830), .ZN(n23828) );
  INV_X1 U23755 ( .A(n23831), .ZN(n23830) );
  OR2_X1 U23756 ( .A1(n23831), .A2(n23832), .ZN(n23827) );
  INV_X1 U23757 ( .A(n23829), .ZN(n23832) );
  OR2_X1 U23758 ( .A1(n15355), .A2(n15354), .ZN(n15912) );
  OR2_X1 U23759 ( .A1(n23833), .A2(n23834), .ZN(n23429) );
  INV_X1 U23760 ( .A(n23835), .ZN(n23834) );
  OR2_X1 U23761 ( .A1(n23836), .A2(n23837), .ZN(n23835) );
  AND2_X1 U23762 ( .A1(n23837), .A2(n23836), .ZN(n23833) );
  AND2_X1 U23763 ( .A1(n23838), .A2(n23839), .ZN(n23836) );
  OR2_X1 U23764 ( .A1(n23840), .A2(n23841), .ZN(n23839) );
  INV_X1 U23765 ( .A(n23842), .ZN(n23841) );
  OR2_X1 U23766 ( .A1(n23842), .A2(n23843), .ZN(n23838) );
  INV_X1 U23767 ( .A(n23840), .ZN(n23843) );
  OR2_X1 U23768 ( .A1(n15389), .A2(n15354), .ZN(n23445) );
  OR2_X1 U23769 ( .A1(n23844), .A2(n23845), .ZN(n23439) );
  INV_X1 U23770 ( .A(n23846), .ZN(n23845) );
  OR2_X1 U23771 ( .A1(n23847), .A2(n23848), .ZN(n23846) );
  AND2_X1 U23772 ( .A1(n23848), .A2(n23847), .ZN(n23844) );
  AND2_X1 U23773 ( .A1(n23849), .A2(n23850), .ZN(n23847) );
  INV_X1 U23774 ( .A(n23851), .ZN(n23850) );
  AND2_X1 U23775 ( .A1(n23852), .A2(n23853), .ZN(n23851) );
  OR2_X1 U23776 ( .A1(n23853), .A2(n23852), .ZN(n23849) );
  INV_X1 U23777 ( .A(n23854), .ZN(n23852) );
  OR2_X1 U23778 ( .A1(n15423), .A2(n15354), .ZN(n23455) );
  AND2_X1 U23779 ( .A1(n23855), .A2(n23856), .ZN(n23450) );
  INV_X1 U23780 ( .A(n23857), .ZN(n23856) );
  AND2_X1 U23781 ( .A1(n23858), .A2(n23859), .ZN(n23857) );
  OR2_X1 U23782 ( .A1(n23859), .A2(n23858), .ZN(n23855) );
  OR2_X1 U23783 ( .A1(n23860), .A2(n23861), .ZN(n23858) );
  AND2_X1 U23784 ( .A1(n23862), .A2(n23863), .ZN(n23861) );
  INV_X1 U23785 ( .A(n15909), .ZN(n23862) );
  AND2_X1 U23786 ( .A1(n23864), .A2(n15909), .ZN(n23860) );
  INV_X1 U23787 ( .A(n23863), .ZN(n23864) );
  OR2_X1 U23788 ( .A1(n15457), .A2(n15354), .ZN(n23466) );
  AND2_X1 U23789 ( .A1(n23865), .A2(n23866), .ZN(n23461) );
  INV_X1 U23790 ( .A(n23867), .ZN(n23866) );
  AND2_X1 U23791 ( .A1(n23868), .A2(n23869), .ZN(n23867) );
  OR2_X1 U23792 ( .A1(n23869), .A2(n23868), .ZN(n23865) );
  OR2_X1 U23793 ( .A1(n23870), .A2(n23871), .ZN(n23868) );
  AND2_X1 U23794 ( .A1(n23872), .A2(n23873), .ZN(n23871) );
  INV_X1 U23795 ( .A(n23874), .ZN(n23872) );
  AND2_X1 U23796 ( .A1(n23875), .A2(n23874), .ZN(n23870) );
  INV_X1 U23797 ( .A(n23873), .ZN(n23875) );
  OR2_X1 U23798 ( .A1(n15491), .A2(n15354), .ZN(n23477) );
  AND2_X1 U23799 ( .A1(n23876), .A2(n23877), .ZN(n23472) );
  INV_X1 U23800 ( .A(n23878), .ZN(n23877) );
  AND2_X1 U23801 ( .A1(n23879), .A2(n23880), .ZN(n23878) );
  OR2_X1 U23802 ( .A1(n23880), .A2(n23879), .ZN(n23876) );
  OR2_X1 U23803 ( .A1(n23881), .A2(n23882), .ZN(n23879) );
  AND2_X1 U23804 ( .A1(n23883), .A2(n23884), .ZN(n23882) );
  INV_X1 U23805 ( .A(n23885), .ZN(n23883) );
  AND2_X1 U23806 ( .A1(n23886), .A2(n23885), .ZN(n23881) );
  INV_X1 U23807 ( .A(n23884), .ZN(n23886) );
  OR2_X1 U23808 ( .A1(n15525), .A2(n15354), .ZN(n23488) );
  AND2_X1 U23809 ( .A1(n23887), .A2(n23888), .ZN(n23483) );
  INV_X1 U23810 ( .A(n23889), .ZN(n23888) );
  AND2_X1 U23811 ( .A1(n23890), .A2(n23891), .ZN(n23889) );
  OR2_X1 U23812 ( .A1(n23891), .A2(n23890), .ZN(n23887) );
  OR2_X1 U23813 ( .A1(n23892), .A2(n23893), .ZN(n23890) );
  AND2_X1 U23814 ( .A1(n23894), .A2(n23895), .ZN(n23893) );
  INV_X1 U23815 ( .A(n23896), .ZN(n23894) );
  AND2_X1 U23816 ( .A1(n23897), .A2(n23896), .ZN(n23892) );
  INV_X1 U23817 ( .A(n23895), .ZN(n23897) );
  OR2_X1 U23818 ( .A1(n15559), .A2(n15354), .ZN(n23499) );
  AND2_X1 U23819 ( .A1(n23898), .A2(n23899), .ZN(n23494) );
  INV_X1 U23820 ( .A(n23900), .ZN(n23899) );
  AND2_X1 U23821 ( .A1(n23901), .A2(n23902), .ZN(n23900) );
  OR2_X1 U23822 ( .A1(n23902), .A2(n23901), .ZN(n23898) );
  OR2_X1 U23823 ( .A1(n23903), .A2(n23904), .ZN(n23901) );
  AND2_X1 U23824 ( .A1(n23905), .A2(n23906), .ZN(n23904) );
  INV_X1 U23825 ( .A(n23907), .ZN(n23905) );
  AND2_X1 U23826 ( .A1(n23908), .A2(n23907), .ZN(n23903) );
  INV_X1 U23827 ( .A(n23906), .ZN(n23908) );
  OR2_X1 U23828 ( .A1(n15593), .A2(n15354), .ZN(n23510) );
  AND2_X1 U23829 ( .A1(n23909), .A2(n23910), .ZN(n23505) );
  INV_X1 U23830 ( .A(n23911), .ZN(n23910) );
  AND2_X1 U23831 ( .A1(n23912), .A2(n23913), .ZN(n23911) );
  OR2_X1 U23832 ( .A1(n23913), .A2(n23912), .ZN(n23909) );
  OR2_X1 U23833 ( .A1(n23914), .A2(n23915), .ZN(n23912) );
  AND2_X1 U23834 ( .A1(n23916), .A2(n23917), .ZN(n23915) );
  INV_X1 U23835 ( .A(n23918), .ZN(n23916) );
  AND2_X1 U23836 ( .A1(n23919), .A2(n23918), .ZN(n23914) );
  INV_X1 U23837 ( .A(n23917), .ZN(n23919) );
  OR2_X1 U23838 ( .A1(n15638), .A2(n15354), .ZN(n23521) );
  AND2_X1 U23839 ( .A1(n23920), .A2(n23921), .ZN(n23516) );
  INV_X1 U23840 ( .A(n23922), .ZN(n23921) );
  AND2_X1 U23841 ( .A1(n23923), .A2(n23924), .ZN(n23922) );
  OR2_X1 U23842 ( .A1(n23924), .A2(n23923), .ZN(n23920) );
  OR2_X1 U23843 ( .A1(n23925), .A2(n23926), .ZN(n23923) );
  AND2_X1 U23844 ( .A1(n23927), .A2(n23928), .ZN(n23926) );
  INV_X1 U23845 ( .A(n23929), .ZN(n23927) );
  AND2_X1 U23846 ( .A1(n23930), .A2(n23929), .ZN(n23925) );
  INV_X1 U23847 ( .A(n23928), .ZN(n23930) );
  OR2_X1 U23848 ( .A1(n15672), .A2(n15354), .ZN(n23532) );
  AND2_X1 U23849 ( .A1(n23931), .A2(n23932), .ZN(n23527) );
  INV_X1 U23850 ( .A(n23933), .ZN(n23932) );
  AND2_X1 U23851 ( .A1(n23934), .A2(n23935), .ZN(n23933) );
  OR2_X1 U23852 ( .A1(n23935), .A2(n23934), .ZN(n23931) );
  OR2_X1 U23853 ( .A1(n23936), .A2(n23937), .ZN(n23934) );
  AND2_X1 U23854 ( .A1(n23938), .A2(n23939), .ZN(n23937) );
  INV_X1 U23855 ( .A(n23940), .ZN(n23938) );
  AND2_X1 U23856 ( .A1(n23941), .A2(n23940), .ZN(n23936) );
  INV_X1 U23857 ( .A(n23939), .ZN(n23941) );
  OR2_X1 U23858 ( .A1(n15706), .A2(n15354), .ZN(n23543) );
  AND2_X1 U23859 ( .A1(n23942), .A2(n23943), .ZN(n23538) );
  INV_X1 U23860 ( .A(n23944), .ZN(n23943) );
  AND2_X1 U23861 ( .A1(n23945), .A2(n23946), .ZN(n23944) );
  OR2_X1 U23862 ( .A1(n23946), .A2(n23945), .ZN(n23942) );
  OR2_X1 U23863 ( .A1(n23947), .A2(n23948), .ZN(n23945) );
  AND2_X1 U23864 ( .A1(n23949), .A2(n23950), .ZN(n23948) );
  INV_X1 U23865 ( .A(n23951), .ZN(n23949) );
  AND2_X1 U23866 ( .A1(n23952), .A2(n23951), .ZN(n23947) );
  INV_X1 U23867 ( .A(n23950), .ZN(n23952) );
  OR2_X1 U23868 ( .A1(n15740), .A2(n15354), .ZN(n23554) );
  AND2_X1 U23869 ( .A1(n23953), .A2(n23954), .ZN(n23549) );
  INV_X1 U23870 ( .A(n23955), .ZN(n23954) );
  AND2_X1 U23871 ( .A1(n23956), .A2(n23957), .ZN(n23955) );
  OR2_X1 U23872 ( .A1(n23957), .A2(n23956), .ZN(n23953) );
  OR2_X1 U23873 ( .A1(n23958), .A2(n23959), .ZN(n23956) );
  AND2_X1 U23874 ( .A1(n23960), .A2(n23961), .ZN(n23959) );
  INV_X1 U23875 ( .A(n23962), .ZN(n23960) );
  AND2_X1 U23876 ( .A1(n23963), .A2(n23962), .ZN(n23958) );
  INV_X1 U23877 ( .A(n23961), .ZN(n23963) );
  OR2_X1 U23878 ( .A1(n15774), .A2(n15354), .ZN(n23565) );
  AND2_X1 U23879 ( .A1(n23964), .A2(n23965), .ZN(n23560) );
  INV_X1 U23880 ( .A(n23966), .ZN(n23965) );
  AND2_X1 U23881 ( .A1(n23967), .A2(n23968), .ZN(n23966) );
  OR2_X1 U23882 ( .A1(n23968), .A2(n23967), .ZN(n23964) );
  OR2_X1 U23883 ( .A1(n23969), .A2(n23970), .ZN(n23967) );
  AND2_X1 U23884 ( .A1(n23971), .A2(n23972), .ZN(n23970) );
  INV_X1 U23885 ( .A(n23973), .ZN(n23971) );
  AND2_X1 U23886 ( .A1(n23974), .A2(n23973), .ZN(n23969) );
  INV_X1 U23887 ( .A(n23972), .ZN(n23974) );
  OR2_X1 U23888 ( .A1(n15808), .A2(n15354), .ZN(n23576) );
  AND2_X1 U23889 ( .A1(n23975), .A2(n23976), .ZN(n23571) );
  INV_X1 U23890 ( .A(n23977), .ZN(n23976) );
  AND2_X1 U23891 ( .A1(n23978), .A2(n23979), .ZN(n23977) );
  OR2_X1 U23892 ( .A1(n23979), .A2(n23978), .ZN(n23975) );
  OR2_X1 U23893 ( .A1(n23980), .A2(n23981), .ZN(n23978) );
  AND2_X1 U23894 ( .A1(n23982), .A2(n23983), .ZN(n23981) );
  INV_X1 U23895 ( .A(n23984), .ZN(n23982) );
  AND2_X1 U23896 ( .A1(n23985), .A2(n23984), .ZN(n23980) );
  INV_X1 U23897 ( .A(n23983), .ZN(n23985) );
  OR2_X1 U23898 ( .A1(n15842), .A2(n15354), .ZN(n23587) );
  INV_X1 U23899 ( .A(b_15_), .ZN(n15354) );
  AND2_X1 U23900 ( .A1(n23986), .A2(n23987), .ZN(n23582) );
  INV_X1 U23901 ( .A(n23988), .ZN(n23987) );
  AND2_X1 U23902 ( .A1(n23989), .A2(n23990), .ZN(n23988) );
  OR2_X1 U23903 ( .A1(n23990), .A2(n23989), .ZN(n23986) );
  OR2_X1 U23904 ( .A1(n23991), .A2(n23992), .ZN(n23989) );
  AND2_X1 U23905 ( .A1(n23993), .A2(n23994), .ZN(n23992) );
  INV_X1 U23906 ( .A(n23995), .ZN(n23993) );
  AND2_X1 U23907 ( .A1(n23996), .A2(n23995), .ZN(n23991) );
  INV_X1 U23908 ( .A(n23994), .ZN(n23996) );
  AND2_X1 U23909 ( .A1(n23997), .A2(n23998), .ZN(n23162) );
  INV_X1 U23910 ( .A(n23999), .ZN(n23998) );
  AND2_X1 U23911 ( .A1(n24000), .A2(n24001), .ZN(n23999) );
  OR2_X1 U23912 ( .A1(n24001), .A2(n24000), .ZN(n23997) );
  OR2_X1 U23913 ( .A1(n24002), .A2(n24003), .ZN(n24000) );
  AND2_X1 U23914 ( .A1(n24004), .A2(n24005), .ZN(n24003) );
  INV_X1 U23915 ( .A(n24006), .ZN(n24004) );
  AND2_X1 U23916 ( .A1(n24007), .A2(n24006), .ZN(n24002) );
  INV_X1 U23917 ( .A(n24005), .ZN(n24007) );
  AND2_X1 U23918 ( .A1(n24008), .A2(n24009), .ZN(n16149) );
  INV_X1 U23919 ( .A(n24010), .ZN(n24009) );
  AND2_X1 U23920 ( .A1(n16646), .A2(n16648), .ZN(n24010) );
  OR2_X1 U23921 ( .A1(n16646), .A2(n16648), .ZN(n24008) );
  OR2_X1 U23922 ( .A1(n24011), .A2(n24012), .ZN(n16648) );
  AND2_X1 U23923 ( .A1(n23173), .A2(n23172), .ZN(n24012) );
  AND2_X1 U23924 ( .A1(n23168), .A2(n24013), .ZN(n24011) );
  OR2_X1 U23925 ( .A1(n23172), .A2(n23173), .ZN(n24013) );
  OR2_X1 U23926 ( .A1(n16512), .A2(n15388), .ZN(n23173) );
  OR2_X1 U23927 ( .A1(n24014), .A2(n24015), .ZN(n23172) );
  AND2_X1 U23928 ( .A1(n24006), .A2(n24005), .ZN(n24015) );
  AND2_X1 U23929 ( .A1(n24001), .A2(n24016), .ZN(n24014) );
  OR2_X1 U23930 ( .A1(n24005), .A2(n24006), .ZN(n24016) );
  OR2_X1 U23931 ( .A1(n15842), .A2(n15388), .ZN(n24006) );
  OR2_X1 U23932 ( .A1(n24017), .A2(n24018), .ZN(n24005) );
  AND2_X1 U23933 ( .A1(n23995), .A2(n23994), .ZN(n24018) );
  AND2_X1 U23934 ( .A1(n23990), .A2(n24019), .ZN(n24017) );
  OR2_X1 U23935 ( .A1(n23994), .A2(n23995), .ZN(n24019) );
  OR2_X1 U23936 ( .A1(n15808), .A2(n15388), .ZN(n23995) );
  OR2_X1 U23937 ( .A1(n24020), .A2(n24021), .ZN(n23994) );
  AND2_X1 U23938 ( .A1(n23984), .A2(n23983), .ZN(n24021) );
  AND2_X1 U23939 ( .A1(n23979), .A2(n24022), .ZN(n24020) );
  OR2_X1 U23940 ( .A1(n23983), .A2(n23984), .ZN(n24022) );
  OR2_X1 U23941 ( .A1(n15774), .A2(n15388), .ZN(n23984) );
  OR2_X1 U23942 ( .A1(n24023), .A2(n24024), .ZN(n23983) );
  AND2_X1 U23943 ( .A1(n23973), .A2(n23972), .ZN(n24024) );
  AND2_X1 U23944 ( .A1(n23968), .A2(n24025), .ZN(n24023) );
  OR2_X1 U23945 ( .A1(n23972), .A2(n23973), .ZN(n24025) );
  OR2_X1 U23946 ( .A1(n15740), .A2(n15388), .ZN(n23973) );
  OR2_X1 U23947 ( .A1(n24026), .A2(n24027), .ZN(n23972) );
  AND2_X1 U23948 ( .A1(n23962), .A2(n23961), .ZN(n24027) );
  AND2_X1 U23949 ( .A1(n23957), .A2(n24028), .ZN(n24026) );
  OR2_X1 U23950 ( .A1(n23961), .A2(n23962), .ZN(n24028) );
  OR2_X1 U23951 ( .A1(n15706), .A2(n15388), .ZN(n23962) );
  OR2_X1 U23952 ( .A1(n24029), .A2(n24030), .ZN(n23961) );
  AND2_X1 U23953 ( .A1(n23951), .A2(n23950), .ZN(n24030) );
  AND2_X1 U23954 ( .A1(n23946), .A2(n24031), .ZN(n24029) );
  OR2_X1 U23955 ( .A1(n23950), .A2(n23951), .ZN(n24031) );
  OR2_X1 U23956 ( .A1(n15672), .A2(n15388), .ZN(n23951) );
  OR2_X1 U23957 ( .A1(n24032), .A2(n24033), .ZN(n23950) );
  AND2_X1 U23958 ( .A1(n23940), .A2(n23939), .ZN(n24033) );
  AND2_X1 U23959 ( .A1(n23935), .A2(n24034), .ZN(n24032) );
  OR2_X1 U23960 ( .A1(n23939), .A2(n23940), .ZN(n24034) );
  OR2_X1 U23961 ( .A1(n15638), .A2(n15388), .ZN(n23940) );
  OR2_X1 U23962 ( .A1(n24035), .A2(n24036), .ZN(n23939) );
  AND2_X1 U23963 ( .A1(n23929), .A2(n23928), .ZN(n24036) );
  AND2_X1 U23964 ( .A1(n23924), .A2(n24037), .ZN(n24035) );
  OR2_X1 U23965 ( .A1(n23928), .A2(n23929), .ZN(n24037) );
  OR2_X1 U23966 ( .A1(n15593), .A2(n15388), .ZN(n23929) );
  OR2_X1 U23967 ( .A1(n24038), .A2(n24039), .ZN(n23928) );
  AND2_X1 U23968 ( .A1(n23918), .A2(n23917), .ZN(n24039) );
  AND2_X1 U23969 ( .A1(n23913), .A2(n24040), .ZN(n24038) );
  OR2_X1 U23970 ( .A1(n23917), .A2(n23918), .ZN(n24040) );
  OR2_X1 U23971 ( .A1(n15559), .A2(n15388), .ZN(n23918) );
  OR2_X1 U23972 ( .A1(n24041), .A2(n24042), .ZN(n23917) );
  AND2_X1 U23973 ( .A1(n23907), .A2(n23906), .ZN(n24042) );
  AND2_X1 U23974 ( .A1(n23902), .A2(n24043), .ZN(n24041) );
  OR2_X1 U23975 ( .A1(n23906), .A2(n23907), .ZN(n24043) );
  OR2_X1 U23976 ( .A1(n15525), .A2(n15388), .ZN(n23907) );
  OR2_X1 U23977 ( .A1(n24044), .A2(n24045), .ZN(n23906) );
  AND2_X1 U23978 ( .A1(n23896), .A2(n23895), .ZN(n24045) );
  AND2_X1 U23979 ( .A1(n23891), .A2(n24046), .ZN(n24044) );
  OR2_X1 U23980 ( .A1(n23895), .A2(n23896), .ZN(n24046) );
  OR2_X1 U23981 ( .A1(n15491), .A2(n15388), .ZN(n23896) );
  OR2_X1 U23982 ( .A1(n24047), .A2(n24048), .ZN(n23895) );
  AND2_X1 U23983 ( .A1(n23885), .A2(n23884), .ZN(n24048) );
  AND2_X1 U23984 ( .A1(n23880), .A2(n24049), .ZN(n24047) );
  OR2_X1 U23985 ( .A1(n23884), .A2(n23885), .ZN(n24049) );
  OR2_X1 U23986 ( .A1(n15457), .A2(n15388), .ZN(n23885) );
  OR2_X1 U23987 ( .A1(n24050), .A2(n24051), .ZN(n23884) );
  AND2_X1 U23988 ( .A1(n23874), .A2(n23873), .ZN(n24051) );
  AND2_X1 U23989 ( .A1(n23869), .A2(n24052), .ZN(n24050) );
  OR2_X1 U23990 ( .A1(n23873), .A2(n23874), .ZN(n24052) );
  OR2_X1 U23991 ( .A1(n15423), .A2(n15388), .ZN(n23874) );
  OR2_X1 U23992 ( .A1(n24053), .A2(n24054), .ZN(n23873) );
  AND2_X1 U23993 ( .A1(n15909), .A2(n23863), .ZN(n24054) );
  AND2_X1 U23994 ( .A1(n23859), .A2(n24055), .ZN(n24053) );
  OR2_X1 U23995 ( .A1(n23863), .A2(n15909), .ZN(n24055) );
  OR2_X1 U23996 ( .A1(n15389), .A2(n15388), .ZN(n15909) );
  OR2_X1 U23997 ( .A1(n24056), .A2(n24057), .ZN(n23863) );
  AND2_X1 U23998 ( .A1(n23854), .A2(n23853), .ZN(n24057) );
  AND2_X1 U23999 ( .A1(n23848), .A2(n24058), .ZN(n24056) );
  OR2_X1 U24000 ( .A1(n23853), .A2(n23854), .ZN(n24058) );
  OR2_X1 U24001 ( .A1(n15355), .A2(n15388), .ZN(n23854) );
  OR2_X1 U24002 ( .A1(n24059), .A2(n24060), .ZN(n23853) );
  AND2_X1 U24003 ( .A1(n23840), .A2(n23842), .ZN(n24060) );
  AND2_X1 U24004 ( .A1(n23837), .A2(n24061), .ZN(n24059) );
  OR2_X1 U24005 ( .A1(n23842), .A2(n23840), .ZN(n24061) );
  OR2_X1 U24006 ( .A1(n15321), .A2(n15388), .ZN(n23840) );
  OR2_X1 U24007 ( .A1(n24062), .A2(n24063), .ZN(n23842) );
  AND2_X1 U24008 ( .A1(n23829), .A2(n23831), .ZN(n24063) );
  AND2_X1 U24009 ( .A1(n23826), .A2(n24064), .ZN(n24062) );
  OR2_X1 U24010 ( .A1(n23831), .A2(n23829), .ZN(n24064) );
  OR2_X1 U24011 ( .A1(n15287), .A2(n15388), .ZN(n23829) );
  OR2_X1 U24012 ( .A1(n24065), .A2(n24066), .ZN(n23831) );
  AND2_X1 U24013 ( .A1(n23818), .A2(n23820), .ZN(n24066) );
  AND2_X1 U24014 ( .A1(n23815), .A2(n24067), .ZN(n24065) );
  OR2_X1 U24015 ( .A1(n23820), .A2(n23818), .ZN(n24067) );
  OR2_X1 U24016 ( .A1(n15242), .A2(n15388), .ZN(n23818) );
  OR2_X1 U24017 ( .A1(n24068), .A2(n24069), .ZN(n23820) );
  AND2_X1 U24018 ( .A1(n23807), .A2(n23809), .ZN(n24069) );
  AND2_X1 U24019 ( .A1(n23804), .A2(n24070), .ZN(n24068) );
  OR2_X1 U24020 ( .A1(n23809), .A2(n23807), .ZN(n24070) );
  OR2_X1 U24021 ( .A1(n15208), .A2(n15388), .ZN(n23807) );
  OR2_X1 U24022 ( .A1(n24071), .A2(n24072), .ZN(n23809) );
  AND2_X1 U24023 ( .A1(n23796), .A2(n23798), .ZN(n24072) );
  AND2_X1 U24024 ( .A1(n23793), .A2(n24073), .ZN(n24071) );
  OR2_X1 U24025 ( .A1(n23798), .A2(n23796), .ZN(n24073) );
  OR2_X1 U24026 ( .A1(n15174), .A2(n15388), .ZN(n23796) );
  OR2_X1 U24027 ( .A1(n24074), .A2(n24075), .ZN(n23798) );
  AND2_X1 U24028 ( .A1(n23785), .A2(n23787), .ZN(n24075) );
  AND2_X1 U24029 ( .A1(n23782), .A2(n24076), .ZN(n24074) );
  OR2_X1 U24030 ( .A1(n23787), .A2(n23785), .ZN(n24076) );
  OR2_X1 U24031 ( .A1(n15140), .A2(n15388), .ZN(n23785) );
  OR2_X1 U24032 ( .A1(n24077), .A2(n24078), .ZN(n23787) );
  AND2_X1 U24033 ( .A1(n23774), .A2(n23776), .ZN(n24078) );
  AND2_X1 U24034 ( .A1(n23771), .A2(n24079), .ZN(n24077) );
  OR2_X1 U24035 ( .A1(n23776), .A2(n23774), .ZN(n24079) );
  OR2_X1 U24036 ( .A1(n15106), .A2(n15388), .ZN(n23774) );
  OR2_X1 U24037 ( .A1(n24080), .A2(n24081), .ZN(n23776) );
  AND2_X1 U24038 ( .A1(n23763), .A2(n23765), .ZN(n24081) );
  AND2_X1 U24039 ( .A1(n23760), .A2(n24082), .ZN(n24080) );
  OR2_X1 U24040 ( .A1(n23765), .A2(n23763), .ZN(n24082) );
  OR2_X1 U24041 ( .A1(n15072), .A2(n15388), .ZN(n23763) );
  OR2_X1 U24042 ( .A1(n24083), .A2(n24084), .ZN(n23765) );
  AND2_X1 U24043 ( .A1(n23752), .A2(n23754), .ZN(n24084) );
  AND2_X1 U24044 ( .A1(n23749), .A2(n24085), .ZN(n24083) );
  OR2_X1 U24045 ( .A1(n23754), .A2(n23752), .ZN(n24085) );
  OR2_X1 U24046 ( .A1(n15038), .A2(n15388), .ZN(n23752) );
  OR2_X1 U24047 ( .A1(n24086), .A2(n24087), .ZN(n23754) );
  AND2_X1 U24048 ( .A1(n23741), .A2(n23743), .ZN(n24087) );
  AND2_X1 U24049 ( .A1(n23738), .A2(n24088), .ZN(n24086) );
  OR2_X1 U24050 ( .A1(n23743), .A2(n23741), .ZN(n24088) );
  OR2_X1 U24051 ( .A1(n15004), .A2(n15388), .ZN(n23741) );
  OR2_X1 U24052 ( .A1(n24089), .A2(n24090), .ZN(n23743) );
  AND2_X1 U24053 ( .A1(n23730), .A2(n23732), .ZN(n24090) );
  AND2_X1 U24054 ( .A1(n23727), .A2(n24091), .ZN(n24089) );
  OR2_X1 U24055 ( .A1(n23732), .A2(n23730), .ZN(n24091) );
  OR2_X1 U24056 ( .A1(n14970), .A2(n15388), .ZN(n23730) );
  OR2_X1 U24057 ( .A1(n24092), .A2(n24093), .ZN(n23732) );
  AND2_X1 U24058 ( .A1(n23719), .A2(n23721), .ZN(n24093) );
  AND2_X1 U24059 ( .A1(n23716), .A2(n24094), .ZN(n24092) );
  OR2_X1 U24060 ( .A1(n23721), .A2(n23719), .ZN(n24094) );
  OR2_X1 U24061 ( .A1(n14936), .A2(n15388), .ZN(n23719) );
  OR2_X1 U24062 ( .A1(n24095), .A2(n24096), .ZN(n23721) );
  AND2_X1 U24063 ( .A1(n23708), .A2(n23710), .ZN(n24096) );
  AND2_X1 U24064 ( .A1(n23705), .A2(n24097), .ZN(n24095) );
  OR2_X1 U24065 ( .A1(n23710), .A2(n23708), .ZN(n24097) );
  OR2_X1 U24066 ( .A1(n14891), .A2(n15388), .ZN(n23708) );
  OR2_X1 U24067 ( .A1(n24098), .A2(n24099), .ZN(n23710) );
  AND2_X1 U24068 ( .A1(n23693), .A2(n23698), .ZN(n24099) );
  AND2_X1 U24069 ( .A1(n23697), .A2(n24100), .ZN(n24098) );
  OR2_X1 U24070 ( .A1(n23698), .A2(n23693), .ZN(n24100) );
  OR2_X1 U24071 ( .A1(n14857), .A2(n15388), .ZN(n23693) );
  INV_X1 U24072 ( .A(b_14_), .ZN(n15388) );
  INV_X1 U24073 ( .A(n23699), .ZN(n23698) );
  AND3_X1 U24074 ( .A1(b_14_), .A2(b_13_), .A3(n15957), .ZN(n23699) );
  INV_X1 U24075 ( .A(n23700), .ZN(n23697) );
  OR2_X1 U24076 ( .A1(n24101), .A2(n24102), .ZN(n23700) );
  AND2_X1 U24077 ( .A1(b_13_), .A2(n24103), .ZN(n24102) );
  OR2_X1 U24078 ( .A1(n24104), .A2(n16981), .ZN(n24103) );
  AND2_X1 U24079 ( .A1(a_30_), .A2(n15456), .ZN(n24104) );
  AND2_X1 U24080 ( .A1(b_12_), .A2(n24105), .ZN(n24101) );
  OR2_X1 U24081 ( .A1(n24106), .A2(n14817), .ZN(n24105) );
  AND2_X1 U24082 ( .A1(a_31_), .A2(n15422), .ZN(n24106) );
  OR2_X1 U24083 ( .A1(n24107), .A2(n24108), .ZN(n23705) );
  AND2_X1 U24084 ( .A1(n24109), .A2(n24110), .ZN(n24108) );
  INV_X1 U24085 ( .A(n24111), .ZN(n24107) );
  OR2_X1 U24086 ( .A1(n24109), .A2(n24110), .ZN(n24111) );
  OR2_X1 U24087 ( .A1(n24112), .A2(n24113), .ZN(n24109) );
  AND2_X1 U24088 ( .A1(n24114), .A2(n24115), .ZN(n24113) );
  AND2_X1 U24089 ( .A1(n24116), .A2(n24117), .ZN(n24112) );
  OR2_X1 U24090 ( .A1(n24118), .A2(n24119), .ZN(n23716) );
  INV_X1 U24091 ( .A(n24120), .ZN(n24119) );
  OR2_X1 U24092 ( .A1(n24121), .A2(n24122), .ZN(n24120) );
  AND2_X1 U24093 ( .A1(n24122), .A2(n24121), .ZN(n24118) );
  AND2_X1 U24094 ( .A1(n24123), .A2(n24124), .ZN(n24121) );
  OR2_X1 U24095 ( .A1(n24125), .A2(n24126), .ZN(n24124) );
  INV_X1 U24096 ( .A(n24127), .ZN(n24126) );
  OR2_X1 U24097 ( .A1(n24127), .A2(n24128), .ZN(n24123) );
  INV_X1 U24098 ( .A(n24125), .ZN(n24128) );
  OR2_X1 U24099 ( .A1(n24129), .A2(n24130), .ZN(n23727) );
  INV_X1 U24100 ( .A(n24131), .ZN(n24130) );
  OR2_X1 U24101 ( .A1(n24132), .A2(n24133), .ZN(n24131) );
  AND2_X1 U24102 ( .A1(n24133), .A2(n24132), .ZN(n24129) );
  AND2_X1 U24103 ( .A1(n24134), .A2(n24135), .ZN(n24132) );
  OR2_X1 U24104 ( .A1(n24136), .A2(n24137), .ZN(n24135) );
  INV_X1 U24105 ( .A(n24138), .ZN(n24137) );
  OR2_X1 U24106 ( .A1(n24138), .A2(n24139), .ZN(n24134) );
  INV_X1 U24107 ( .A(n24136), .ZN(n24139) );
  OR2_X1 U24108 ( .A1(n24140), .A2(n24141), .ZN(n23738) );
  INV_X1 U24109 ( .A(n24142), .ZN(n24141) );
  OR2_X1 U24110 ( .A1(n24143), .A2(n24144), .ZN(n24142) );
  AND2_X1 U24111 ( .A1(n24144), .A2(n24143), .ZN(n24140) );
  AND2_X1 U24112 ( .A1(n24145), .A2(n24146), .ZN(n24143) );
  OR2_X1 U24113 ( .A1(n24147), .A2(n24148), .ZN(n24146) );
  INV_X1 U24114 ( .A(n24149), .ZN(n24148) );
  OR2_X1 U24115 ( .A1(n24149), .A2(n24150), .ZN(n24145) );
  INV_X1 U24116 ( .A(n24147), .ZN(n24150) );
  OR2_X1 U24117 ( .A1(n24151), .A2(n24152), .ZN(n23749) );
  INV_X1 U24118 ( .A(n24153), .ZN(n24152) );
  OR2_X1 U24119 ( .A1(n24154), .A2(n24155), .ZN(n24153) );
  AND2_X1 U24120 ( .A1(n24155), .A2(n24154), .ZN(n24151) );
  AND2_X1 U24121 ( .A1(n24156), .A2(n24157), .ZN(n24154) );
  OR2_X1 U24122 ( .A1(n24158), .A2(n24159), .ZN(n24157) );
  INV_X1 U24123 ( .A(n24160), .ZN(n24159) );
  OR2_X1 U24124 ( .A1(n24160), .A2(n24161), .ZN(n24156) );
  INV_X1 U24125 ( .A(n24158), .ZN(n24161) );
  OR2_X1 U24126 ( .A1(n24162), .A2(n24163), .ZN(n23760) );
  INV_X1 U24127 ( .A(n24164), .ZN(n24163) );
  OR2_X1 U24128 ( .A1(n24165), .A2(n24166), .ZN(n24164) );
  AND2_X1 U24129 ( .A1(n24166), .A2(n24165), .ZN(n24162) );
  AND2_X1 U24130 ( .A1(n24167), .A2(n24168), .ZN(n24165) );
  OR2_X1 U24131 ( .A1(n24169), .A2(n24170), .ZN(n24168) );
  INV_X1 U24132 ( .A(n24171), .ZN(n24170) );
  OR2_X1 U24133 ( .A1(n24171), .A2(n24172), .ZN(n24167) );
  INV_X1 U24134 ( .A(n24169), .ZN(n24172) );
  OR2_X1 U24135 ( .A1(n24173), .A2(n24174), .ZN(n23771) );
  INV_X1 U24136 ( .A(n24175), .ZN(n24174) );
  OR2_X1 U24137 ( .A1(n24176), .A2(n24177), .ZN(n24175) );
  AND2_X1 U24138 ( .A1(n24177), .A2(n24176), .ZN(n24173) );
  AND2_X1 U24139 ( .A1(n24178), .A2(n24179), .ZN(n24176) );
  OR2_X1 U24140 ( .A1(n24180), .A2(n24181), .ZN(n24179) );
  INV_X1 U24141 ( .A(n24182), .ZN(n24181) );
  OR2_X1 U24142 ( .A1(n24182), .A2(n24183), .ZN(n24178) );
  INV_X1 U24143 ( .A(n24180), .ZN(n24183) );
  OR2_X1 U24144 ( .A1(n24184), .A2(n24185), .ZN(n23782) );
  INV_X1 U24145 ( .A(n24186), .ZN(n24185) );
  OR2_X1 U24146 ( .A1(n24187), .A2(n24188), .ZN(n24186) );
  AND2_X1 U24147 ( .A1(n24188), .A2(n24187), .ZN(n24184) );
  AND2_X1 U24148 ( .A1(n24189), .A2(n24190), .ZN(n24187) );
  OR2_X1 U24149 ( .A1(n24191), .A2(n24192), .ZN(n24190) );
  INV_X1 U24150 ( .A(n24193), .ZN(n24192) );
  OR2_X1 U24151 ( .A1(n24193), .A2(n24194), .ZN(n24189) );
  INV_X1 U24152 ( .A(n24191), .ZN(n24194) );
  OR2_X1 U24153 ( .A1(n24195), .A2(n24196), .ZN(n23793) );
  INV_X1 U24154 ( .A(n24197), .ZN(n24196) );
  OR2_X1 U24155 ( .A1(n24198), .A2(n24199), .ZN(n24197) );
  AND2_X1 U24156 ( .A1(n24199), .A2(n24198), .ZN(n24195) );
  AND2_X1 U24157 ( .A1(n24200), .A2(n24201), .ZN(n24198) );
  OR2_X1 U24158 ( .A1(n24202), .A2(n24203), .ZN(n24201) );
  INV_X1 U24159 ( .A(n24204), .ZN(n24203) );
  OR2_X1 U24160 ( .A1(n24204), .A2(n24205), .ZN(n24200) );
  INV_X1 U24161 ( .A(n24202), .ZN(n24205) );
  OR2_X1 U24162 ( .A1(n24206), .A2(n24207), .ZN(n23804) );
  INV_X1 U24163 ( .A(n24208), .ZN(n24207) );
  OR2_X1 U24164 ( .A1(n24209), .A2(n24210), .ZN(n24208) );
  AND2_X1 U24165 ( .A1(n24210), .A2(n24209), .ZN(n24206) );
  AND2_X1 U24166 ( .A1(n24211), .A2(n24212), .ZN(n24209) );
  OR2_X1 U24167 ( .A1(n24213), .A2(n24214), .ZN(n24212) );
  INV_X1 U24168 ( .A(n24215), .ZN(n24214) );
  OR2_X1 U24169 ( .A1(n24215), .A2(n24216), .ZN(n24211) );
  INV_X1 U24170 ( .A(n24213), .ZN(n24216) );
  OR2_X1 U24171 ( .A1(n24217), .A2(n24218), .ZN(n23815) );
  INV_X1 U24172 ( .A(n24219), .ZN(n24218) );
  OR2_X1 U24173 ( .A1(n24220), .A2(n24221), .ZN(n24219) );
  AND2_X1 U24174 ( .A1(n24221), .A2(n24220), .ZN(n24217) );
  AND2_X1 U24175 ( .A1(n24222), .A2(n24223), .ZN(n24220) );
  OR2_X1 U24176 ( .A1(n24224), .A2(n24225), .ZN(n24223) );
  INV_X1 U24177 ( .A(n24226), .ZN(n24225) );
  OR2_X1 U24178 ( .A1(n24226), .A2(n24227), .ZN(n24222) );
  INV_X1 U24179 ( .A(n24224), .ZN(n24227) );
  OR2_X1 U24180 ( .A1(n24228), .A2(n24229), .ZN(n23826) );
  INV_X1 U24181 ( .A(n24230), .ZN(n24229) );
  OR2_X1 U24182 ( .A1(n24231), .A2(n24232), .ZN(n24230) );
  AND2_X1 U24183 ( .A1(n24232), .A2(n24231), .ZN(n24228) );
  AND2_X1 U24184 ( .A1(n24233), .A2(n24234), .ZN(n24231) );
  OR2_X1 U24185 ( .A1(n24235), .A2(n24236), .ZN(n24234) );
  INV_X1 U24186 ( .A(n24237), .ZN(n24236) );
  OR2_X1 U24187 ( .A1(n24237), .A2(n24238), .ZN(n24233) );
  INV_X1 U24188 ( .A(n24235), .ZN(n24238) );
  OR2_X1 U24189 ( .A1(n24239), .A2(n24240), .ZN(n23837) );
  INV_X1 U24190 ( .A(n24241), .ZN(n24240) );
  OR2_X1 U24191 ( .A1(n24242), .A2(n24243), .ZN(n24241) );
  AND2_X1 U24192 ( .A1(n24243), .A2(n24242), .ZN(n24239) );
  AND2_X1 U24193 ( .A1(n24244), .A2(n24245), .ZN(n24242) );
  OR2_X1 U24194 ( .A1(n24246), .A2(n24247), .ZN(n24245) );
  INV_X1 U24195 ( .A(n24248), .ZN(n24247) );
  OR2_X1 U24196 ( .A1(n24248), .A2(n24249), .ZN(n24244) );
  INV_X1 U24197 ( .A(n24246), .ZN(n24249) );
  OR2_X1 U24198 ( .A1(n24250), .A2(n24251), .ZN(n23848) );
  INV_X1 U24199 ( .A(n24252), .ZN(n24251) );
  OR2_X1 U24200 ( .A1(n24253), .A2(n24254), .ZN(n24252) );
  AND2_X1 U24201 ( .A1(n24254), .A2(n24253), .ZN(n24250) );
  AND2_X1 U24202 ( .A1(n24255), .A2(n24256), .ZN(n24253) );
  INV_X1 U24203 ( .A(n24257), .ZN(n24256) );
  AND2_X1 U24204 ( .A1(n24258), .A2(n24259), .ZN(n24257) );
  OR2_X1 U24205 ( .A1(n24259), .A2(n24258), .ZN(n24255) );
  INV_X1 U24206 ( .A(n24260), .ZN(n24258) );
  AND2_X1 U24207 ( .A1(n24261), .A2(n24262), .ZN(n23859) );
  INV_X1 U24208 ( .A(n24263), .ZN(n24262) );
  AND2_X1 U24209 ( .A1(n24264), .A2(n24265), .ZN(n24263) );
  OR2_X1 U24210 ( .A1(n24265), .A2(n24264), .ZN(n24261) );
  OR2_X1 U24211 ( .A1(n24266), .A2(n24267), .ZN(n24264) );
  AND2_X1 U24212 ( .A1(n24268), .A2(n24269), .ZN(n24267) );
  INV_X1 U24213 ( .A(n24270), .ZN(n24268) );
  AND2_X1 U24214 ( .A1(n24271), .A2(n24270), .ZN(n24266) );
  INV_X1 U24215 ( .A(n24269), .ZN(n24271) );
  AND2_X1 U24216 ( .A1(n24272), .A2(n24273), .ZN(n23869) );
  INV_X1 U24217 ( .A(n24274), .ZN(n24273) );
  AND2_X1 U24218 ( .A1(n24275), .A2(n24276), .ZN(n24274) );
  OR2_X1 U24219 ( .A1(n24276), .A2(n24275), .ZN(n24272) );
  OR2_X1 U24220 ( .A1(n24277), .A2(n24278), .ZN(n24275) );
  AND2_X1 U24221 ( .A1(n24279), .A2(n24280), .ZN(n24278) );
  INV_X1 U24222 ( .A(n24281), .ZN(n24279) );
  AND2_X1 U24223 ( .A1(n24282), .A2(n24281), .ZN(n24277) );
  INV_X1 U24224 ( .A(n24280), .ZN(n24282) );
  AND2_X1 U24225 ( .A1(n24283), .A2(n24284), .ZN(n23880) );
  INV_X1 U24226 ( .A(n24285), .ZN(n24284) );
  AND2_X1 U24227 ( .A1(n24286), .A2(n24287), .ZN(n24285) );
  OR2_X1 U24228 ( .A1(n24287), .A2(n24286), .ZN(n24283) );
  OR2_X1 U24229 ( .A1(n24288), .A2(n24289), .ZN(n24286) );
  AND2_X1 U24230 ( .A1(n24290), .A2(n24291), .ZN(n24289) );
  INV_X1 U24231 ( .A(n15906), .ZN(n24290) );
  AND2_X1 U24232 ( .A1(n24292), .A2(n15906), .ZN(n24288) );
  INV_X1 U24233 ( .A(n24291), .ZN(n24292) );
  AND2_X1 U24234 ( .A1(n24293), .A2(n24294), .ZN(n23891) );
  INV_X1 U24235 ( .A(n24295), .ZN(n24294) );
  AND2_X1 U24236 ( .A1(n24296), .A2(n24297), .ZN(n24295) );
  OR2_X1 U24237 ( .A1(n24297), .A2(n24296), .ZN(n24293) );
  OR2_X1 U24238 ( .A1(n24298), .A2(n24299), .ZN(n24296) );
  AND2_X1 U24239 ( .A1(n24300), .A2(n24301), .ZN(n24299) );
  INV_X1 U24240 ( .A(n24302), .ZN(n24300) );
  AND2_X1 U24241 ( .A1(n24303), .A2(n24302), .ZN(n24298) );
  INV_X1 U24242 ( .A(n24301), .ZN(n24303) );
  AND2_X1 U24243 ( .A1(n24304), .A2(n24305), .ZN(n23902) );
  INV_X1 U24244 ( .A(n24306), .ZN(n24305) );
  AND2_X1 U24245 ( .A1(n24307), .A2(n24308), .ZN(n24306) );
  OR2_X1 U24246 ( .A1(n24308), .A2(n24307), .ZN(n24304) );
  OR2_X1 U24247 ( .A1(n24309), .A2(n24310), .ZN(n24307) );
  AND2_X1 U24248 ( .A1(n24311), .A2(n24312), .ZN(n24310) );
  INV_X1 U24249 ( .A(n24313), .ZN(n24311) );
  AND2_X1 U24250 ( .A1(n24314), .A2(n24313), .ZN(n24309) );
  INV_X1 U24251 ( .A(n24312), .ZN(n24314) );
  AND2_X1 U24252 ( .A1(n24315), .A2(n24316), .ZN(n23913) );
  INV_X1 U24253 ( .A(n24317), .ZN(n24316) );
  AND2_X1 U24254 ( .A1(n24318), .A2(n24319), .ZN(n24317) );
  OR2_X1 U24255 ( .A1(n24319), .A2(n24318), .ZN(n24315) );
  OR2_X1 U24256 ( .A1(n24320), .A2(n24321), .ZN(n24318) );
  AND2_X1 U24257 ( .A1(n24322), .A2(n24323), .ZN(n24321) );
  INV_X1 U24258 ( .A(n24324), .ZN(n24322) );
  AND2_X1 U24259 ( .A1(n24325), .A2(n24324), .ZN(n24320) );
  INV_X1 U24260 ( .A(n24323), .ZN(n24325) );
  AND2_X1 U24261 ( .A1(n24326), .A2(n24327), .ZN(n23924) );
  INV_X1 U24262 ( .A(n24328), .ZN(n24327) );
  AND2_X1 U24263 ( .A1(n24329), .A2(n24330), .ZN(n24328) );
  OR2_X1 U24264 ( .A1(n24330), .A2(n24329), .ZN(n24326) );
  OR2_X1 U24265 ( .A1(n24331), .A2(n24332), .ZN(n24329) );
  AND2_X1 U24266 ( .A1(n24333), .A2(n24334), .ZN(n24332) );
  INV_X1 U24267 ( .A(n24335), .ZN(n24333) );
  AND2_X1 U24268 ( .A1(n24336), .A2(n24335), .ZN(n24331) );
  INV_X1 U24269 ( .A(n24334), .ZN(n24336) );
  AND2_X1 U24270 ( .A1(n24337), .A2(n24338), .ZN(n23935) );
  INV_X1 U24271 ( .A(n24339), .ZN(n24338) );
  AND2_X1 U24272 ( .A1(n24340), .A2(n24341), .ZN(n24339) );
  OR2_X1 U24273 ( .A1(n24341), .A2(n24340), .ZN(n24337) );
  OR2_X1 U24274 ( .A1(n24342), .A2(n24343), .ZN(n24340) );
  AND2_X1 U24275 ( .A1(n24344), .A2(n24345), .ZN(n24343) );
  INV_X1 U24276 ( .A(n24346), .ZN(n24344) );
  AND2_X1 U24277 ( .A1(n24347), .A2(n24346), .ZN(n24342) );
  INV_X1 U24278 ( .A(n24345), .ZN(n24347) );
  AND2_X1 U24279 ( .A1(n24348), .A2(n24349), .ZN(n23946) );
  INV_X1 U24280 ( .A(n24350), .ZN(n24349) );
  AND2_X1 U24281 ( .A1(n24351), .A2(n24352), .ZN(n24350) );
  OR2_X1 U24282 ( .A1(n24352), .A2(n24351), .ZN(n24348) );
  OR2_X1 U24283 ( .A1(n24353), .A2(n24354), .ZN(n24351) );
  AND2_X1 U24284 ( .A1(n24355), .A2(n24356), .ZN(n24354) );
  INV_X1 U24285 ( .A(n24357), .ZN(n24355) );
  AND2_X1 U24286 ( .A1(n24358), .A2(n24357), .ZN(n24353) );
  INV_X1 U24287 ( .A(n24356), .ZN(n24358) );
  AND2_X1 U24288 ( .A1(n24359), .A2(n24360), .ZN(n23957) );
  INV_X1 U24289 ( .A(n24361), .ZN(n24360) );
  AND2_X1 U24290 ( .A1(n24362), .A2(n24363), .ZN(n24361) );
  OR2_X1 U24291 ( .A1(n24363), .A2(n24362), .ZN(n24359) );
  OR2_X1 U24292 ( .A1(n24364), .A2(n24365), .ZN(n24362) );
  AND2_X1 U24293 ( .A1(n24366), .A2(n24367), .ZN(n24365) );
  INV_X1 U24294 ( .A(n24368), .ZN(n24366) );
  AND2_X1 U24295 ( .A1(n24369), .A2(n24368), .ZN(n24364) );
  INV_X1 U24296 ( .A(n24367), .ZN(n24369) );
  AND2_X1 U24297 ( .A1(n24370), .A2(n24371), .ZN(n23968) );
  INV_X1 U24298 ( .A(n24372), .ZN(n24371) );
  AND2_X1 U24299 ( .A1(n24373), .A2(n24374), .ZN(n24372) );
  OR2_X1 U24300 ( .A1(n24374), .A2(n24373), .ZN(n24370) );
  OR2_X1 U24301 ( .A1(n24375), .A2(n24376), .ZN(n24373) );
  AND2_X1 U24302 ( .A1(n24377), .A2(n24378), .ZN(n24376) );
  INV_X1 U24303 ( .A(n24379), .ZN(n24377) );
  AND2_X1 U24304 ( .A1(n24380), .A2(n24379), .ZN(n24375) );
  INV_X1 U24305 ( .A(n24378), .ZN(n24380) );
  AND2_X1 U24306 ( .A1(n24381), .A2(n24382), .ZN(n23979) );
  INV_X1 U24307 ( .A(n24383), .ZN(n24382) );
  AND2_X1 U24308 ( .A1(n24384), .A2(n24385), .ZN(n24383) );
  OR2_X1 U24309 ( .A1(n24385), .A2(n24384), .ZN(n24381) );
  OR2_X1 U24310 ( .A1(n24386), .A2(n24387), .ZN(n24384) );
  AND2_X1 U24311 ( .A1(n24388), .A2(n24389), .ZN(n24387) );
  INV_X1 U24312 ( .A(n24390), .ZN(n24388) );
  AND2_X1 U24313 ( .A1(n24391), .A2(n24390), .ZN(n24386) );
  INV_X1 U24314 ( .A(n24389), .ZN(n24391) );
  AND2_X1 U24315 ( .A1(n24392), .A2(n24393), .ZN(n23990) );
  INV_X1 U24316 ( .A(n24394), .ZN(n24393) );
  AND2_X1 U24317 ( .A1(n24395), .A2(n24396), .ZN(n24394) );
  OR2_X1 U24318 ( .A1(n24396), .A2(n24395), .ZN(n24392) );
  OR2_X1 U24319 ( .A1(n24397), .A2(n24398), .ZN(n24395) );
  AND2_X1 U24320 ( .A1(n24399), .A2(n24400), .ZN(n24398) );
  INV_X1 U24321 ( .A(n24401), .ZN(n24399) );
  AND2_X1 U24322 ( .A1(n24402), .A2(n24401), .ZN(n24397) );
  INV_X1 U24323 ( .A(n24400), .ZN(n24402) );
  AND2_X1 U24324 ( .A1(n24403), .A2(n24404), .ZN(n24001) );
  INV_X1 U24325 ( .A(n24405), .ZN(n24404) );
  AND2_X1 U24326 ( .A1(n24406), .A2(n24407), .ZN(n24405) );
  OR2_X1 U24327 ( .A1(n24407), .A2(n24406), .ZN(n24403) );
  OR2_X1 U24328 ( .A1(n24408), .A2(n24409), .ZN(n24406) );
  AND2_X1 U24329 ( .A1(n24410), .A2(n24411), .ZN(n24409) );
  INV_X1 U24330 ( .A(n24412), .ZN(n24410) );
  AND2_X1 U24331 ( .A1(n24413), .A2(n24412), .ZN(n24408) );
  INV_X1 U24332 ( .A(n24411), .ZN(n24413) );
  AND2_X1 U24333 ( .A1(n24414), .A2(n24415), .ZN(n23168) );
  INV_X1 U24334 ( .A(n24416), .ZN(n24415) );
  AND2_X1 U24335 ( .A1(n24417), .A2(n24418), .ZN(n24416) );
  OR2_X1 U24336 ( .A1(n24418), .A2(n24417), .ZN(n24414) );
  OR2_X1 U24337 ( .A1(n24419), .A2(n24420), .ZN(n24417) );
  AND2_X1 U24338 ( .A1(n24421), .A2(n24422), .ZN(n24420) );
  INV_X1 U24339 ( .A(n24423), .ZN(n24421) );
  AND2_X1 U24340 ( .A1(n24424), .A2(n24423), .ZN(n24419) );
  INV_X1 U24341 ( .A(n24422), .ZN(n24424) );
  OR2_X1 U24342 ( .A1(n24425), .A2(n24426), .ZN(n16646) );
  AND2_X1 U24343 ( .A1(n24427), .A2(n16591), .ZN(n24426) );
  INV_X1 U24344 ( .A(n24428), .ZN(n24425) );
  OR2_X1 U24345 ( .A1(n16591), .A2(n24427), .ZN(n24428) );
  OR2_X1 U24346 ( .A1(n24429), .A2(n24430), .ZN(n24427) );
  AND2_X1 U24347 ( .A1(n24431), .A2(n16590), .ZN(n24430) );
  INV_X1 U24348 ( .A(n16589), .ZN(n24431) );
  AND2_X1 U24349 ( .A1(n24432), .A2(n16589), .ZN(n24429) );
  OR2_X1 U24350 ( .A1(n16512), .A2(n15422), .ZN(n16589) );
  INV_X1 U24351 ( .A(n16590), .ZN(n24432) );
  OR2_X1 U24352 ( .A1(n24433), .A2(n24434), .ZN(n16590) );
  AND2_X1 U24353 ( .A1(n24423), .A2(n24422), .ZN(n24434) );
  AND2_X1 U24354 ( .A1(n24418), .A2(n24435), .ZN(n24433) );
  OR2_X1 U24355 ( .A1(n24423), .A2(n24422), .ZN(n24435) );
  OR2_X1 U24356 ( .A1(n24436), .A2(n24437), .ZN(n24422) );
  AND2_X1 U24357 ( .A1(n24412), .A2(n24411), .ZN(n24437) );
  AND2_X1 U24358 ( .A1(n24407), .A2(n24438), .ZN(n24436) );
  OR2_X1 U24359 ( .A1(n24412), .A2(n24411), .ZN(n24438) );
  OR2_X1 U24360 ( .A1(n24439), .A2(n24440), .ZN(n24411) );
  AND2_X1 U24361 ( .A1(n24401), .A2(n24400), .ZN(n24440) );
  AND2_X1 U24362 ( .A1(n24396), .A2(n24441), .ZN(n24439) );
  OR2_X1 U24363 ( .A1(n24401), .A2(n24400), .ZN(n24441) );
  OR2_X1 U24364 ( .A1(n24442), .A2(n24443), .ZN(n24400) );
  AND2_X1 U24365 ( .A1(n24390), .A2(n24389), .ZN(n24443) );
  AND2_X1 U24366 ( .A1(n24385), .A2(n24444), .ZN(n24442) );
  OR2_X1 U24367 ( .A1(n24390), .A2(n24389), .ZN(n24444) );
  OR2_X1 U24368 ( .A1(n24445), .A2(n24446), .ZN(n24389) );
  AND2_X1 U24369 ( .A1(n24379), .A2(n24378), .ZN(n24446) );
  AND2_X1 U24370 ( .A1(n24374), .A2(n24447), .ZN(n24445) );
  OR2_X1 U24371 ( .A1(n24379), .A2(n24378), .ZN(n24447) );
  OR2_X1 U24372 ( .A1(n24448), .A2(n24449), .ZN(n24378) );
  AND2_X1 U24373 ( .A1(n24368), .A2(n24367), .ZN(n24449) );
  AND2_X1 U24374 ( .A1(n24363), .A2(n24450), .ZN(n24448) );
  OR2_X1 U24375 ( .A1(n24368), .A2(n24367), .ZN(n24450) );
  OR2_X1 U24376 ( .A1(n24451), .A2(n24452), .ZN(n24367) );
  AND2_X1 U24377 ( .A1(n24357), .A2(n24356), .ZN(n24452) );
  AND2_X1 U24378 ( .A1(n24352), .A2(n24453), .ZN(n24451) );
  OR2_X1 U24379 ( .A1(n24357), .A2(n24356), .ZN(n24453) );
  OR2_X1 U24380 ( .A1(n24454), .A2(n24455), .ZN(n24356) );
  AND2_X1 U24381 ( .A1(n24346), .A2(n24345), .ZN(n24455) );
  AND2_X1 U24382 ( .A1(n24341), .A2(n24456), .ZN(n24454) );
  OR2_X1 U24383 ( .A1(n24346), .A2(n24345), .ZN(n24456) );
  OR2_X1 U24384 ( .A1(n24457), .A2(n24458), .ZN(n24345) );
  AND2_X1 U24385 ( .A1(n24335), .A2(n24334), .ZN(n24458) );
  AND2_X1 U24386 ( .A1(n24330), .A2(n24459), .ZN(n24457) );
  OR2_X1 U24387 ( .A1(n24335), .A2(n24334), .ZN(n24459) );
  OR2_X1 U24388 ( .A1(n24460), .A2(n24461), .ZN(n24334) );
  AND2_X1 U24389 ( .A1(n24324), .A2(n24323), .ZN(n24461) );
  AND2_X1 U24390 ( .A1(n24319), .A2(n24462), .ZN(n24460) );
  OR2_X1 U24391 ( .A1(n24324), .A2(n24323), .ZN(n24462) );
  OR2_X1 U24392 ( .A1(n24463), .A2(n24464), .ZN(n24323) );
  AND2_X1 U24393 ( .A1(n24313), .A2(n24312), .ZN(n24464) );
  AND2_X1 U24394 ( .A1(n24308), .A2(n24465), .ZN(n24463) );
  OR2_X1 U24395 ( .A1(n24313), .A2(n24312), .ZN(n24465) );
  OR2_X1 U24396 ( .A1(n24466), .A2(n24467), .ZN(n24312) );
  AND2_X1 U24397 ( .A1(n24302), .A2(n24301), .ZN(n24467) );
  AND2_X1 U24398 ( .A1(n24297), .A2(n24468), .ZN(n24466) );
  OR2_X1 U24399 ( .A1(n24302), .A2(n24301), .ZN(n24468) );
  OR2_X1 U24400 ( .A1(n24469), .A2(n24470), .ZN(n24301) );
  AND2_X1 U24401 ( .A1(n15906), .A2(n24291), .ZN(n24470) );
  AND2_X1 U24402 ( .A1(n24287), .A2(n24471), .ZN(n24469) );
  OR2_X1 U24403 ( .A1(n15906), .A2(n24291), .ZN(n24471) );
  OR2_X1 U24404 ( .A1(n24472), .A2(n24473), .ZN(n24291) );
  AND2_X1 U24405 ( .A1(n24281), .A2(n24280), .ZN(n24473) );
  AND2_X1 U24406 ( .A1(n24276), .A2(n24474), .ZN(n24472) );
  OR2_X1 U24407 ( .A1(n24281), .A2(n24280), .ZN(n24474) );
  OR2_X1 U24408 ( .A1(n24475), .A2(n24476), .ZN(n24280) );
  AND2_X1 U24409 ( .A1(n24270), .A2(n24269), .ZN(n24476) );
  AND2_X1 U24410 ( .A1(n24265), .A2(n24477), .ZN(n24475) );
  OR2_X1 U24411 ( .A1(n24270), .A2(n24269), .ZN(n24477) );
  OR2_X1 U24412 ( .A1(n24478), .A2(n24479), .ZN(n24269) );
  AND2_X1 U24413 ( .A1(n24260), .A2(n24259), .ZN(n24479) );
  AND2_X1 U24414 ( .A1(n24254), .A2(n24480), .ZN(n24478) );
  OR2_X1 U24415 ( .A1(n24260), .A2(n24259), .ZN(n24480) );
  OR2_X1 U24416 ( .A1(n24481), .A2(n24482), .ZN(n24259) );
  AND2_X1 U24417 ( .A1(n24246), .A2(n24248), .ZN(n24482) );
  AND2_X1 U24418 ( .A1(n24243), .A2(n24483), .ZN(n24481) );
  OR2_X1 U24419 ( .A1(n24246), .A2(n24248), .ZN(n24483) );
  OR2_X1 U24420 ( .A1(n24484), .A2(n24485), .ZN(n24248) );
  AND2_X1 U24421 ( .A1(n24235), .A2(n24237), .ZN(n24485) );
  AND2_X1 U24422 ( .A1(n24232), .A2(n24486), .ZN(n24484) );
  OR2_X1 U24423 ( .A1(n24235), .A2(n24237), .ZN(n24486) );
  OR2_X1 U24424 ( .A1(n24487), .A2(n24488), .ZN(n24237) );
  AND2_X1 U24425 ( .A1(n24224), .A2(n24226), .ZN(n24488) );
  AND2_X1 U24426 ( .A1(n24221), .A2(n24489), .ZN(n24487) );
  OR2_X1 U24427 ( .A1(n24224), .A2(n24226), .ZN(n24489) );
  OR2_X1 U24428 ( .A1(n24490), .A2(n24491), .ZN(n24226) );
  AND2_X1 U24429 ( .A1(n24213), .A2(n24215), .ZN(n24491) );
  AND2_X1 U24430 ( .A1(n24210), .A2(n24492), .ZN(n24490) );
  OR2_X1 U24431 ( .A1(n24213), .A2(n24215), .ZN(n24492) );
  OR2_X1 U24432 ( .A1(n24493), .A2(n24494), .ZN(n24215) );
  AND2_X1 U24433 ( .A1(n24202), .A2(n24204), .ZN(n24494) );
  AND2_X1 U24434 ( .A1(n24199), .A2(n24495), .ZN(n24493) );
  OR2_X1 U24435 ( .A1(n24202), .A2(n24204), .ZN(n24495) );
  OR2_X1 U24436 ( .A1(n24496), .A2(n24497), .ZN(n24204) );
  AND2_X1 U24437 ( .A1(n24191), .A2(n24193), .ZN(n24497) );
  AND2_X1 U24438 ( .A1(n24188), .A2(n24498), .ZN(n24496) );
  OR2_X1 U24439 ( .A1(n24191), .A2(n24193), .ZN(n24498) );
  OR2_X1 U24440 ( .A1(n24499), .A2(n24500), .ZN(n24193) );
  AND2_X1 U24441 ( .A1(n24180), .A2(n24182), .ZN(n24500) );
  AND2_X1 U24442 ( .A1(n24177), .A2(n24501), .ZN(n24499) );
  OR2_X1 U24443 ( .A1(n24180), .A2(n24182), .ZN(n24501) );
  OR2_X1 U24444 ( .A1(n24502), .A2(n24503), .ZN(n24182) );
  AND2_X1 U24445 ( .A1(n24169), .A2(n24171), .ZN(n24503) );
  AND2_X1 U24446 ( .A1(n24166), .A2(n24504), .ZN(n24502) );
  OR2_X1 U24447 ( .A1(n24169), .A2(n24171), .ZN(n24504) );
  OR2_X1 U24448 ( .A1(n24505), .A2(n24506), .ZN(n24171) );
  AND2_X1 U24449 ( .A1(n24158), .A2(n24160), .ZN(n24506) );
  AND2_X1 U24450 ( .A1(n24155), .A2(n24507), .ZN(n24505) );
  OR2_X1 U24451 ( .A1(n24158), .A2(n24160), .ZN(n24507) );
  OR2_X1 U24452 ( .A1(n24508), .A2(n24509), .ZN(n24160) );
  AND2_X1 U24453 ( .A1(n24147), .A2(n24149), .ZN(n24509) );
  AND2_X1 U24454 ( .A1(n24144), .A2(n24510), .ZN(n24508) );
  OR2_X1 U24455 ( .A1(n24147), .A2(n24149), .ZN(n24510) );
  OR2_X1 U24456 ( .A1(n24511), .A2(n24512), .ZN(n24149) );
  AND2_X1 U24457 ( .A1(n24136), .A2(n24138), .ZN(n24512) );
  AND2_X1 U24458 ( .A1(n24133), .A2(n24513), .ZN(n24511) );
  OR2_X1 U24459 ( .A1(n24136), .A2(n24138), .ZN(n24513) );
  OR2_X1 U24460 ( .A1(n24514), .A2(n24515), .ZN(n24138) );
  AND2_X1 U24461 ( .A1(n24125), .A2(n24127), .ZN(n24515) );
  AND2_X1 U24462 ( .A1(n24122), .A2(n24516), .ZN(n24514) );
  OR2_X1 U24463 ( .A1(n24125), .A2(n24127), .ZN(n24516) );
  OR2_X1 U24464 ( .A1(n24517), .A2(n24518), .ZN(n24127) );
  AND2_X1 U24465 ( .A1(n24110), .A2(n24115), .ZN(n24518) );
  AND2_X1 U24466 ( .A1(n24114), .A2(n24519), .ZN(n24517) );
  OR2_X1 U24467 ( .A1(n24110), .A2(n24115), .ZN(n24519) );
  INV_X1 U24468 ( .A(n24116), .ZN(n24115) );
  AND3_X1 U24469 ( .A1(b_13_), .A2(b_12_), .A3(n15957), .ZN(n24116) );
  OR2_X1 U24470 ( .A1(n14857), .A2(n15422), .ZN(n24110) );
  INV_X1 U24471 ( .A(n24117), .ZN(n24114) );
  OR2_X1 U24472 ( .A1(n24520), .A2(n24521), .ZN(n24117) );
  AND2_X1 U24473 ( .A1(b_12_), .A2(n24522), .ZN(n24521) );
  OR2_X1 U24474 ( .A1(n24523), .A2(n16981), .ZN(n24522) );
  AND2_X1 U24475 ( .A1(a_30_), .A2(n15490), .ZN(n24523) );
  AND2_X1 U24476 ( .A1(b_11_), .A2(n24524), .ZN(n24520) );
  OR2_X1 U24477 ( .A1(n24525), .A2(n14817), .ZN(n24524) );
  AND2_X1 U24478 ( .A1(a_31_), .A2(n15456), .ZN(n24525) );
  OR2_X1 U24479 ( .A1(n14891), .A2(n15422), .ZN(n24125) );
  OR2_X1 U24480 ( .A1(n24526), .A2(n24527), .ZN(n24122) );
  AND2_X1 U24481 ( .A1(n24528), .A2(n24529), .ZN(n24527) );
  INV_X1 U24482 ( .A(n24530), .ZN(n24526) );
  OR2_X1 U24483 ( .A1(n24528), .A2(n24529), .ZN(n24530) );
  OR2_X1 U24484 ( .A1(n24531), .A2(n24532), .ZN(n24528) );
  AND2_X1 U24485 ( .A1(n24533), .A2(n24534), .ZN(n24532) );
  AND2_X1 U24486 ( .A1(n24535), .A2(n24536), .ZN(n24531) );
  OR2_X1 U24487 ( .A1(n14936), .A2(n15422), .ZN(n24136) );
  OR2_X1 U24488 ( .A1(n24537), .A2(n24538), .ZN(n24133) );
  INV_X1 U24489 ( .A(n24539), .ZN(n24538) );
  OR2_X1 U24490 ( .A1(n24540), .A2(n24541), .ZN(n24539) );
  AND2_X1 U24491 ( .A1(n24541), .A2(n24540), .ZN(n24537) );
  AND2_X1 U24492 ( .A1(n24542), .A2(n24543), .ZN(n24540) );
  OR2_X1 U24493 ( .A1(n24544), .A2(n24545), .ZN(n24543) );
  INV_X1 U24494 ( .A(n24546), .ZN(n24545) );
  OR2_X1 U24495 ( .A1(n24546), .A2(n24547), .ZN(n24542) );
  INV_X1 U24496 ( .A(n24544), .ZN(n24547) );
  OR2_X1 U24497 ( .A1(n14970), .A2(n15422), .ZN(n24147) );
  OR2_X1 U24498 ( .A1(n24548), .A2(n24549), .ZN(n24144) );
  INV_X1 U24499 ( .A(n24550), .ZN(n24549) );
  OR2_X1 U24500 ( .A1(n24551), .A2(n24552), .ZN(n24550) );
  AND2_X1 U24501 ( .A1(n24552), .A2(n24551), .ZN(n24548) );
  AND2_X1 U24502 ( .A1(n24553), .A2(n24554), .ZN(n24551) );
  OR2_X1 U24503 ( .A1(n24555), .A2(n24556), .ZN(n24554) );
  INV_X1 U24504 ( .A(n24557), .ZN(n24556) );
  OR2_X1 U24505 ( .A1(n24557), .A2(n24558), .ZN(n24553) );
  INV_X1 U24506 ( .A(n24555), .ZN(n24558) );
  OR2_X1 U24507 ( .A1(n15004), .A2(n15422), .ZN(n24158) );
  OR2_X1 U24508 ( .A1(n24559), .A2(n24560), .ZN(n24155) );
  INV_X1 U24509 ( .A(n24561), .ZN(n24560) );
  OR2_X1 U24510 ( .A1(n24562), .A2(n24563), .ZN(n24561) );
  AND2_X1 U24511 ( .A1(n24563), .A2(n24562), .ZN(n24559) );
  AND2_X1 U24512 ( .A1(n24564), .A2(n24565), .ZN(n24562) );
  OR2_X1 U24513 ( .A1(n24566), .A2(n24567), .ZN(n24565) );
  INV_X1 U24514 ( .A(n24568), .ZN(n24567) );
  OR2_X1 U24515 ( .A1(n24568), .A2(n24569), .ZN(n24564) );
  INV_X1 U24516 ( .A(n24566), .ZN(n24569) );
  OR2_X1 U24517 ( .A1(n15038), .A2(n15422), .ZN(n24169) );
  OR2_X1 U24518 ( .A1(n24570), .A2(n24571), .ZN(n24166) );
  INV_X1 U24519 ( .A(n24572), .ZN(n24571) );
  OR2_X1 U24520 ( .A1(n24573), .A2(n24574), .ZN(n24572) );
  AND2_X1 U24521 ( .A1(n24574), .A2(n24573), .ZN(n24570) );
  AND2_X1 U24522 ( .A1(n24575), .A2(n24576), .ZN(n24573) );
  OR2_X1 U24523 ( .A1(n24577), .A2(n24578), .ZN(n24576) );
  INV_X1 U24524 ( .A(n24579), .ZN(n24578) );
  OR2_X1 U24525 ( .A1(n24579), .A2(n24580), .ZN(n24575) );
  INV_X1 U24526 ( .A(n24577), .ZN(n24580) );
  OR2_X1 U24527 ( .A1(n15072), .A2(n15422), .ZN(n24180) );
  OR2_X1 U24528 ( .A1(n24581), .A2(n24582), .ZN(n24177) );
  INV_X1 U24529 ( .A(n24583), .ZN(n24582) );
  OR2_X1 U24530 ( .A1(n24584), .A2(n24585), .ZN(n24583) );
  AND2_X1 U24531 ( .A1(n24585), .A2(n24584), .ZN(n24581) );
  AND2_X1 U24532 ( .A1(n24586), .A2(n24587), .ZN(n24584) );
  OR2_X1 U24533 ( .A1(n24588), .A2(n24589), .ZN(n24587) );
  INV_X1 U24534 ( .A(n24590), .ZN(n24589) );
  OR2_X1 U24535 ( .A1(n24590), .A2(n24591), .ZN(n24586) );
  INV_X1 U24536 ( .A(n24588), .ZN(n24591) );
  OR2_X1 U24537 ( .A1(n15106), .A2(n15422), .ZN(n24191) );
  OR2_X1 U24538 ( .A1(n24592), .A2(n24593), .ZN(n24188) );
  INV_X1 U24539 ( .A(n24594), .ZN(n24593) );
  OR2_X1 U24540 ( .A1(n24595), .A2(n24596), .ZN(n24594) );
  AND2_X1 U24541 ( .A1(n24596), .A2(n24595), .ZN(n24592) );
  AND2_X1 U24542 ( .A1(n24597), .A2(n24598), .ZN(n24595) );
  OR2_X1 U24543 ( .A1(n24599), .A2(n24600), .ZN(n24598) );
  INV_X1 U24544 ( .A(n24601), .ZN(n24600) );
  OR2_X1 U24545 ( .A1(n24601), .A2(n24602), .ZN(n24597) );
  INV_X1 U24546 ( .A(n24599), .ZN(n24602) );
  OR2_X1 U24547 ( .A1(n15140), .A2(n15422), .ZN(n24202) );
  OR2_X1 U24548 ( .A1(n24603), .A2(n24604), .ZN(n24199) );
  INV_X1 U24549 ( .A(n24605), .ZN(n24604) );
  OR2_X1 U24550 ( .A1(n24606), .A2(n24607), .ZN(n24605) );
  AND2_X1 U24551 ( .A1(n24607), .A2(n24606), .ZN(n24603) );
  AND2_X1 U24552 ( .A1(n24608), .A2(n24609), .ZN(n24606) );
  OR2_X1 U24553 ( .A1(n24610), .A2(n24611), .ZN(n24609) );
  INV_X1 U24554 ( .A(n24612), .ZN(n24611) );
  OR2_X1 U24555 ( .A1(n24612), .A2(n24613), .ZN(n24608) );
  INV_X1 U24556 ( .A(n24610), .ZN(n24613) );
  OR2_X1 U24557 ( .A1(n15174), .A2(n15422), .ZN(n24213) );
  OR2_X1 U24558 ( .A1(n24614), .A2(n24615), .ZN(n24210) );
  INV_X1 U24559 ( .A(n24616), .ZN(n24615) );
  OR2_X1 U24560 ( .A1(n24617), .A2(n24618), .ZN(n24616) );
  AND2_X1 U24561 ( .A1(n24618), .A2(n24617), .ZN(n24614) );
  AND2_X1 U24562 ( .A1(n24619), .A2(n24620), .ZN(n24617) );
  OR2_X1 U24563 ( .A1(n24621), .A2(n24622), .ZN(n24620) );
  INV_X1 U24564 ( .A(n24623), .ZN(n24622) );
  OR2_X1 U24565 ( .A1(n24623), .A2(n24624), .ZN(n24619) );
  INV_X1 U24566 ( .A(n24621), .ZN(n24624) );
  OR2_X1 U24567 ( .A1(n15208), .A2(n15422), .ZN(n24224) );
  OR2_X1 U24568 ( .A1(n24625), .A2(n24626), .ZN(n24221) );
  INV_X1 U24569 ( .A(n24627), .ZN(n24626) );
  OR2_X1 U24570 ( .A1(n24628), .A2(n24629), .ZN(n24627) );
  AND2_X1 U24571 ( .A1(n24629), .A2(n24628), .ZN(n24625) );
  AND2_X1 U24572 ( .A1(n24630), .A2(n24631), .ZN(n24628) );
  OR2_X1 U24573 ( .A1(n24632), .A2(n24633), .ZN(n24631) );
  INV_X1 U24574 ( .A(n24634), .ZN(n24633) );
  OR2_X1 U24575 ( .A1(n24634), .A2(n24635), .ZN(n24630) );
  INV_X1 U24576 ( .A(n24632), .ZN(n24635) );
  OR2_X1 U24577 ( .A1(n15242), .A2(n15422), .ZN(n24235) );
  OR2_X1 U24578 ( .A1(n24636), .A2(n24637), .ZN(n24232) );
  INV_X1 U24579 ( .A(n24638), .ZN(n24637) );
  OR2_X1 U24580 ( .A1(n24639), .A2(n24640), .ZN(n24638) );
  AND2_X1 U24581 ( .A1(n24640), .A2(n24639), .ZN(n24636) );
  AND2_X1 U24582 ( .A1(n24641), .A2(n24642), .ZN(n24639) );
  OR2_X1 U24583 ( .A1(n24643), .A2(n24644), .ZN(n24642) );
  INV_X1 U24584 ( .A(n24645), .ZN(n24644) );
  OR2_X1 U24585 ( .A1(n24645), .A2(n24646), .ZN(n24641) );
  INV_X1 U24586 ( .A(n24643), .ZN(n24646) );
  OR2_X1 U24587 ( .A1(n15287), .A2(n15422), .ZN(n24246) );
  OR2_X1 U24588 ( .A1(n24647), .A2(n24648), .ZN(n24243) );
  INV_X1 U24589 ( .A(n24649), .ZN(n24648) );
  OR2_X1 U24590 ( .A1(n24650), .A2(n24651), .ZN(n24649) );
  AND2_X1 U24591 ( .A1(n24651), .A2(n24650), .ZN(n24647) );
  AND2_X1 U24592 ( .A1(n24652), .A2(n24653), .ZN(n24650) );
  OR2_X1 U24593 ( .A1(n24654), .A2(n24655), .ZN(n24653) );
  INV_X1 U24594 ( .A(n24656), .ZN(n24655) );
  OR2_X1 U24595 ( .A1(n24656), .A2(n24657), .ZN(n24652) );
  INV_X1 U24596 ( .A(n24654), .ZN(n24657) );
  OR2_X1 U24597 ( .A1(n15321), .A2(n15422), .ZN(n24260) );
  OR2_X1 U24598 ( .A1(n24658), .A2(n24659), .ZN(n24254) );
  INV_X1 U24599 ( .A(n24660), .ZN(n24659) );
  OR2_X1 U24600 ( .A1(n24661), .A2(n24662), .ZN(n24660) );
  AND2_X1 U24601 ( .A1(n24662), .A2(n24661), .ZN(n24658) );
  AND2_X1 U24602 ( .A1(n24663), .A2(n24664), .ZN(n24661) );
  INV_X1 U24603 ( .A(n24665), .ZN(n24664) );
  AND2_X1 U24604 ( .A1(n24666), .A2(n24667), .ZN(n24665) );
  OR2_X1 U24605 ( .A1(n24667), .A2(n24666), .ZN(n24663) );
  INV_X1 U24606 ( .A(n24668), .ZN(n24666) );
  OR2_X1 U24607 ( .A1(n15355), .A2(n15422), .ZN(n24270) );
  AND2_X1 U24608 ( .A1(n24669), .A2(n24670), .ZN(n24265) );
  INV_X1 U24609 ( .A(n24671), .ZN(n24670) );
  AND2_X1 U24610 ( .A1(n24672), .A2(n24673), .ZN(n24671) );
  OR2_X1 U24611 ( .A1(n24673), .A2(n24672), .ZN(n24669) );
  OR2_X1 U24612 ( .A1(n24674), .A2(n24675), .ZN(n24672) );
  AND2_X1 U24613 ( .A1(n24676), .A2(n24677), .ZN(n24675) );
  INV_X1 U24614 ( .A(n24678), .ZN(n24676) );
  AND2_X1 U24615 ( .A1(n24679), .A2(n24678), .ZN(n24674) );
  INV_X1 U24616 ( .A(n24677), .ZN(n24679) );
  OR2_X1 U24617 ( .A1(n15389), .A2(n15422), .ZN(n24281) );
  AND2_X1 U24618 ( .A1(n24680), .A2(n24681), .ZN(n24276) );
  INV_X1 U24619 ( .A(n24682), .ZN(n24681) );
  AND2_X1 U24620 ( .A1(n24683), .A2(n24684), .ZN(n24682) );
  OR2_X1 U24621 ( .A1(n24684), .A2(n24683), .ZN(n24680) );
  OR2_X1 U24622 ( .A1(n24685), .A2(n24686), .ZN(n24683) );
  AND2_X1 U24623 ( .A1(n24687), .A2(n24688), .ZN(n24686) );
  INV_X1 U24624 ( .A(n24689), .ZN(n24687) );
  AND2_X1 U24625 ( .A1(n24690), .A2(n24689), .ZN(n24685) );
  INV_X1 U24626 ( .A(n24688), .ZN(n24690) );
  OR2_X1 U24627 ( .A1(n15423), .A2(n15422), .ZN(n15906) );
  AND2_X1 U24628 ( .A1(n24691), .A2(n24692), .ZN(n24287) );
  INV_X1 U24629 ( .A(n24693), .ZN(n24692) );
  AND2_X1 U24630 ( .A1(n24694), .A2(n24695), .ZN(n24693) );
  OR2_X1 U24631 ( .A1(n24695), .A2(n24694), .ZN(n24691) );
  OR2_X1 U24632 ( .A1(n24696), .A2(n24697), .ZN(n24694) );
  AND2_X1 U24633 ( .A1(n24698), .A2(n24699), .ZN(n24697) );
  INV_X1 U24634 ( .A(n24700), .ZN(n24698) );
  AND2_X1 U24635 ( .A1(n24701), .A2(n24700), .ZN(n24696) );
  INV_X1 U24636 ( .A(n24699), .ZN(n24701) );
  OR2_X1 U24637 ( .A1(n15457), .A2(n15422), .ZN(n24302) );
  AND2_X1 U24638 ( .A1(n24702), .A2(n24703), .ZN(n24297) );
  INV_X1 U24639 ( .A(n24704), .ZN(n24703) );
  AND2_X1 U24640 ( .A1(n24705), .A2(n24706), .ZN(n24704) );
  OR2_X1 U24641 ( .A1(n24706), .A2(n24705), .ZN(n24702) );
  OR2_X1 U24642 ( .A1(n24707), .A2(n24708), .ZN(n24705) );
  AND2_X1 U24643 ( .A1(n24709), .A2(n24710), .ZN(n24708) );
  INV_X1 U24644 ( .A(n24711), .ZN(n24709) );
  AND2_X1 U24645 ( .A1(n24712), .A2(n24711), .ZN(n24707) );
  INV_X1 U24646 ( .A(n24710), .ZN(n24712) );
  OR2_X1 U24647 ( .A1(n15491), .A2(n15422), .ZN(n24313) );
  AND2_X1 U24648 ( .A1(n24713), .A2(n24714), .ZN(n24308) );
  INV_X1 U24649 ( .A(n24715), .ZN(n24714) );
  AND2_X1 U24650 ( .A1(n24716), .A2(n24717), .ZN(n24715) );
  OR2_X1 U24651 ( .A1(n24717), .A2(n24716), .ZN(n24713) );
  OR2_X1 U24652 ( .A1(n24718), .A2(n24719), .ZN(n24716) );
  AND2_X1 U24653 ( .A1(n24720), .A2(n24721), .ZN(n24719) );
  INV_X1 U24654 ( .A(n15903), .ZN(n24720) );
  AND2_X1 U24655 ( .A1(n24722), .A2(n15903), .ZN(n24718) );
  INV_X1 U24656 ( .A(n24721), .ZN(n24722) );
  OR2_X1 U24657 ( .A1(n15525), .A2(n15422), .ZN(n24324) );
  AND2_X1 U24658 ( .A1(n24723), .A2(n24724), .ZN(n24319) );
  INV_X1 U24659 ( .A(n24725), .ZN(n24724) );
  AND2_X1 U24660 ( .A1(n24726), .A2(n24727), .ZN(n24725) );
  OR2_X1 U24661 ( .A1(n24727), .A2(n24726), .ZN(n24723) );
  OR2_X1 U24662 ( .A1(n24728), .A2(n24729), .ZN(n24726) );
  AND2_X1 U24663 ( .A1(n24730), .A2(n24731), .ZN(n24729) );
  INV_X1 U24664 ( .A(n24732), .ZN(n24730) );
  AND2_X1 U24665 ( .A1(n24733), .A2(n24732), .ZN(n24728) );
  INV_X1 U24666 ( .A(n24731), .ZN(n24733) );
  OR2_X1 U24667 ( .A1(n15559), .A2(n15422), .ZN(n24335) );
  AND2_X1 U24668 ( .A1(n24734), .A2(n24735), .ZN(n24330) );
  INV_X1 U24669 ( .A(n24736), .ZN(n24735) );
  AND2_X1 U24670 ( .A1(n24737), .A2(n24738), .ZN(n24736) );
  OR2_X1 U24671 ( .A1(n24738), .A2(n24737), .ZN(n24734) );
  OR2_X1 U24672 ( .A1(n24739), .A2(n24740), .ZN(n24737) );
  AND2_X1 U24673 ( .A1(n24741), .A2(n24742), .ZN(n24740) );
  INV_X1 U24674 ( .A(n24743), .ZN(n24741) );
  AND2_X1 U24675 ( .A1(n24744), .A2(n24743), .ZN(n24739) );
  INV_X1 U24676 ( .A(n24742), .ZN(n24744) );
  OR2_X1 U24677 ( .A1(n15593), .A2(n15422), .ZN(n24346) );
  AND2_X1 U24678 ( .A1(n24745), .A2(n24746), .ZN(n24341) );
  INV_X1 U24679 ( .A(n24747), .ZN(n24746) );
  AND2_X1 U24680 ( .A1(n24748), .A2(n24749), .ZN(n24747) );
  OR2_X1 U24681 ( .A1(n24749), .A2(n24748), .ZN(n24745) );
  OR2_X1 U24682 ( .A1(n24750), .A2(n24751), .ZN(n24748) );
  AND2_X1 U24683 ( .A1(n24752), .A2(n24753), .ZN(n24751) );
  INV_X1 U24684 ( .A(n24754), .ZN(n24752) );
  AND2_X1 U24685 ( .A1(n24755), .A2(n24754), .ZN(n24750) );
  INV_X1 U24686 ( .A(n24753), .ZN(n24755) );
  OR2_X1 U24687 ( .A1(n15638), .A2(n15422), .ZN(n24357) );
  AND2_X1 U24688 ( .A1(n24756), .A2(n24757), .ZN(n24352) );
  INV_X1 U24689 ( .A(n24758), .ZN(n24757) );
  AND2_X1 U24690 ( .A1(n24759), .A2(n24760), .ZN(n24758) );
  OR2_X1 U24691 ( .A1(n24760), .A2(n24759), .ZN(n24756) );
  OR2_X1 U24692 ( .A1(n24761), .A2(n24762), .ZN(n24759) );
  AND2_X1 U24693 ( .A1(n24763), .A2(n24764), .ZN(n24762) );
  INV_X1 U24694 ( .A(n24765), .ZN(n24763) );
  AND2_X1 U24695 ( .A1(n24766), .A2(n24765), .ZN(n24761) );
  INV_X1 U24696 ( .A(n24764), .ZN(n24766) );
  OR2_X1 U24697 ( .A1(n15672), .A2(n15422), .ZN(n24368) );
  AND2_X1 U24698 ( .A1(n24767), .A2(n24768), .ZN(n24363) );
  INV_X1 U24699 ( .A(n24769), .ZN(n24768) );
  AND2_X1 U24700 ( .A1(n24770), .A2(n24771), .ZN(n24769) );
  OR2_X1 U24701 ( .A1(n24771), .A2(n24770), .ZN(n24767) );
  OR2_X1 U24702 ( .A1(n24772), .A2(n24773), .ZN(n24770) );
  AND2_X1 U24703 ( .A1(n24774), .A2(n24775), .ZN(n24773) );
  INV_X1 U24704 ( .A(n24776), .ZN(n24774) );
  AND2_X1 U24705 ( .A1(n24777), .A2(n24776), .ZN(n24772) );
  INV_X1 U24706 ( .A(n24775), .ZN(n24777) );
  OR2_X1 U24707 ( .A1(n15706), .A2(n15422), .ZN(n24379) );
  AND2_X1 U24708 ( .A1(n24778), .A2(n24779), .ZN(n24374) );
  INV_X1 U24709 ( .A(n24780), .ZN(n24779) );
  AND2_X1 U24710 ( .A1(n24781), .A2(n24782), .ZN(n24780) );
  OR2_X1 U24711 ( .A1(n24782), .A2(n24781), .ZN(n24778) );
  OR2_X1 U24712 ( .A1(n24783), .A2(n24784), .ZN(n24781) );
  AND2_X1 U24713 ( .A1(n24785), .A2(n24786), .ZN(n24784) );
  INV_X1 U24714 ( .A(n24787), .ZN(n24785) );
  AND2_X1 U24715 ( .A1(n24788), .A2(n24787), .ZN(n24783) );
  INV_X1 U24716 ( .A(n24786), .ZN(n24788) );
  OR2_X1 U24717 ( .A1(n15740), .A2(n15422), .ZN(n24390) );
  AND2_X1 U24718 ( .A1(n24789), .A2(n24790), .ZN(n24385) );
  INV_X1 U24719 ( .A(n24791), .ZN(n24790) );
  AND2_X1 U24720 ( .A1(n24792), .A2(n24793), .ZN(n24791) );
  OR2_X1 U24721 ( .A1(n24793), .A2(n24792), .ZN(n24789) );
  OR2_X1 U24722 ( .A1(n24794), .A2(n24795), .ZN(n24792) );
  AND2_X1 U24723 ( .A1(n24796), .A2(n24797), .ZN(n24795) );
  INV_X1 U24724 ( .A(n24798), .ZN(n24796) );
  AND2_X1 U24725 ( .A1(n24799), .A2(n24798), .ZN(n24794) );
  INV_X1 U24726 ( .A(n24797), .ZN(n24799) );
  OR2_X1 U24727 ( .A1(n15774), .A2(n15422), .ZN(n24401) );
  AND2_X1 U24728 ( .A1(n24800), .A2(n24801), .ZN(n24396) );
  INV_X1 U24729 ( .A(n24802), .ZN(n24801) );
  AND2_X1 U24730 ( .A1(n24803), .A2(n24804), .ZN(n24802) );
  OR2_X1 U24731 ( .A1(n24804), .A2(n24803), .ZN(n24800) );
  OR2_X1 U24732 ( .A1(n24805), .A2(n24806), .ZN(n24803) );
  AND2_X1 U24733 ( .A1(n24807), .A2(n24808), .ZN(n24806) );
  INV_X1 U24734 ( .A(n24809), .ZN(n24807) );
  AND2_X1 U24735 ( .A1(n24810), .A2(n24809), .ZN(n24805) );
  INV_X1 U24736 ( .A(n24808), .ZN(n24810) );
  OR2_X1 U24737 ( .A1(n15808), .A2(n15422), .ZN(n24412) );
  AND2_X1 U24738 ( .A1(n24811), .A2(n24812), .ZN(n24407) );
  INV_X1 U24739 ( .A(n24813), .ZN(n24812) );
  AND2_X1 U24740 ( .A1(n24814), .A2(n24815), .ZN(n24813) );
  OR2_X1 U24741 ( .A1(n24815), .A2(n24814), .ZN(n24811) );
  OR2_X1 U24742 ( .A1(n24816), .A2(n24817), .ZN(n24814) );
  AND2_X1 U24743 ( .A1(n24818), .A2(n24819), .ZN(n24817) );
  INV_X1 U24744 ( .A(n24820), .ZN(n24818) );
  AND2_X1 U24745 ( .A1(n24821), .A2(n24820), .ZN(n24816) );
  INV_X1 U24746 ( .A(n24819), .ZN(n24821) );
  OR2_X1 U24747 ( .A1(n15842), .A2(n15422), .ZN(n24423) );
  INV_X1 U24748 ( .A(b_13_), .ZN(n15422) );
  AND2_X1 U24749 ( .A1(n24822), .A2(n24823), .ZN(n24418) );
  INV_X1 U24750 ( .A(n24824), .ZN(n24823) );
  AND2_X1 U24751 ( .A1(n24825), .A2(n24826), .ZN(n24824) );
  OR2_X1 U24752 ( .A1(n24826), .A2(n24825), .ZN(n24822) );
  OR2_X1 U24753 ( .A1(n24827), .A2(n24828), .ZN(n24825) );
  AND2_X1 U24754 ( .A1(n24829), .A2(n24830), .ZN(n24828) );
  INV_X1 U24755 ( .A(n24831), .ZN(n24829) );
  AND2_X1 U24756 ( .A1(n24832), .A2(n24831), .ZN(n24827) );
  INV_X1 U24757 ( .A(n24830), .ZN(n24832) );
  AND2_X1 U24758 ( .A1(n24833), .A2(n24834), .ZN(n16591) );
  INV_X1 U24759 ( .A(n24835), .ZN(n24834) );
  AND2_X1 U24760 ( .A1(n24836), .A2(n16605), .ZN(n24835) );
  OR2_X1 U24761 ( .A1(n16605), .A2(n24836), .ZN(n24833) );
  OR2_X1 U24762 ( .A1(n24837), .A2(n24838), .ZN(n24836) );
  AND2_X1 U24763 ( .A1(n24839), .A2(n16604), .ZN(n24838) );
  INV_X1 U24764 ( .A(n16603), .ZN(n24839) );
  AND2_X1 U24765 ( .A1(n24840), .A2(n16603), .ZN(n24837) );
  OR2_X1 U24766 ( .A1(n15842), .A2(n15456), .ZN(n16603) );
  INV_X1 U24767 ( .A(n16604), .ZN(n24840) );
  OR2_X1 U24768 ( .A1(n24841), .A2(n24842), .ZN(n16604) );
  AND2_X1 U24769 ( .A1(n24831), .A2(n24830), .ZN(n24842) );
  AND2_X1 U24770 ( .A1(n24826), .A2(n24843), .ZN(n24841) );
  OR2_X1 U24771 ( .A1(n24830), .A2(n24831), .ZN(n24843) );
  OR2_X1 U24772 ( .A1(n15808), .A2(n15456), .ZN(n24831) );
  OR2_X1 U24773 ( .A1(n24844), .A2(n24845), .ZN(n24830) );
  AND2_X1 U24774 ( .A1(n24820), .A2(n24819), .ZN(n24845) );
  AND2_X1 U24775 ( .A1(n24815), .A2(n24846), .ZN(n24844) );
  OR2_X1 U24776 ( .A1(n24819), .A2(n24820), .ZN(n24846) );
  OR2_X1 U24777 ( .A1(n15774), .A2(n15456), .ZN(n24820) );
  OR2_X1 U24778 ( .A1(n24847), .A2(n24848), .ZN(n24819) );
  AND2_X1 U24779 ( .A1(n24809), .A2(n24808), .ZN(n24848) );
  AND2_X1 U24780 ( .A1(n24804), .A2(n24849), .ZN(n24847) );
  OR2_X1 U24781 ( .A1(n24808), .A2(n24809), .ZN(n24849) );
  OR2_X1 U24782 ( .A1(n15740), .A2(n15456), .ZN(n24809) );
  OR2_X1 U24783 ( .A1(n24850), .A2(n24851), .ZN(n24808) );
  AND2_X1 U24784 ( .A1(n24798), .A2(n24797), .ZN(n24851) );
  AND2_X1 U24785 ( .A1(n24793), .A2(n24852), .ZN(n24850) );
  OR2_X1 U24786 ( .A1(n24797), .A2(n24798), .ZN(n24852) );
  OR2_X1 U24787 ( .A1(n15706), .A2(n15456), .ZN(n24798) );
  OR2_X1 U24788 ( .A1(n24853), .A2(n24854), .ZN(n24797) );
  AND2_X1 U24789 ( .A1(n24787), .A2(n24786), .ZN(n24854) );
  AND2_X1 U24790 ( .A1(n24782), .A2(n24855), .ZN(n24853) );
  OR2_X1 U24791 ( .A1(n24786), .A2(n24787), .ZN(n24855) );
  OR2_X1 U24792 ( .A1(n15672), .A2(n15456), .ZN(n24787) );
  OR2_X1 U24793 ( .A1(n24856), .A2(n24857), .ZN(n24786) );
  AND2_X1 U24794 ( .A1(n24776), .A2(n24775), .ZN(n24857) );
  AND2_X1 U24795 ( .A1(n24771), .A2(n24858), .ZN(n24856) );
  OR2_X1 U24796 ( .A1(n24775), .A2(n24776), .ZN(n24858) );
  OR2_X1 U24797 ( .A1(n15638), .A2(n15456), .ZN(n24776) );
  OR2_X1 U24798 ( .A1(n24859), .A2(n24860), .ZN(n24775) );
  AND2_X1 U24799 ( .A1(n24765), .A2(n24764), .ZN(n24860) );
  AND2_X1 U24800 ( .A1(n24760), .A2(n24861), .ZN(n24859) );
  OR2_X1 U24801 ( .A1(n24764), .A2(n24765), .ZN(n24861) );
  OR2_X1 U24802 ( .A1(n15593), .A2(n15456), .ZN(n24765) );
  OR2_X1 U24803 ( .A1(n24862), .A2(n24863), .ZN(n24764) );
  AND2_X1 U24804 ( .A1(n24754), .A2(n24753), .ZN(n24863) );
  AND2_X1 U24805 ( .A1(n24749), .A2(n24864), .ZN(n24862) );
  OR2_X1 U24806 ( .A1(n24753), .A2(n24754), .ZN(n24864) );
  OR2_X1 U24807 ( .A1(n15559), .A2(n15456), .ZN(n24754) );
  OR2_X1 U24808 ( .A1(n24865), .A2(n24866), .ZN(n24753) );
  AND2_X1 U24809 ( .A1(n24743), .A2(n24742), .ZN(n24866) );
  AND2_X1 U24810 ( .A1(n24738), .A2(n24867), .ZN(n24865) );
  OR2_X1 U24811 ( .A1(n24742), .A2(n24743), .ZN(n24867) );
  OR2_X1 U24812 ( .A1(n15525), .A2(n15456), .ZN(n24743) );
  OR2_X1 U24813 ( .A1(n24868), .A2(n24869), .ZN(n24742) );
  AND2_X1 U24814 ( .A1(n24732), .A2(n24731), .ZN(n24869) );
  AND2_X1 U24815 ( .A1(n24727), .A2(n24870), .ZN(n24868) );
  OR2_X1 U24816 ( .A1(n24731), .A2(n24732), .ZN(n24870) );
  OR2_X1 U24817 ( .A1(n15491), .A2(n15456), .ZN(n24732) );
  OR2_X1 U24818 ( .A1(n24871), .A2(n24872), .ZN(n24731) );
  AND2_X1 U24819 ( .A1(n15903), .A2(n24721), .ZN(n24872) );
  AND2_X1 U24820 ( .A1(n24717), .A2(n24873), .ZN(n24871) );
  OR2_X1 U24821 ( .A1(n24721), .A2(n15903), .ZN(n24873) );
  OR2_X1 U24822 ( .A1(n15457), .A2(n15456), .ZN(n15903) );
  OR2_X1 U24823 ( .A1(n24874), .A2(n24875), .ZN(n24721) );
  AND2_X1 U24824 ( .A1(n24711), .A2(n24710), .ZN(n24875) );
  AND2_X1 U24825 ( .A1(n24706), .A2(n24876), .ZN(n24874) );
  OR2_X1 U24826 ( .A1(n24710), .A2(n24711), .ZN(n24876) );
  OR2_X1 U24827 ( .A1(n15423), .A2(n15456), .ZN(n24711) );
  OR2_X1 U24828 ( .A1(n24877), .A2(n24878), .ZN(n24710) );
  AND2_X1 U24829 ( .A1(n24700), .A2(n24699), .ZN(n24878) );
  AND2_X1 U24830 ( .A1(n24695), .A2(n24879), .ZN(n24877) );
  OR2_X1 U24831 ( .A1(n24699), .A2(n24700), .ZN(n24879) );
  OR2_X1 U24832 ( .A1(n15389), .A2(n15456), .ZN(n24700) );
  OR2_X1 U24833 ( .A1(n24880), .A2(n24881), .ZN(n24699) );
  AND2_X1 U24834 ( .A1(n24689), .A2(n24688), .ZN(n24881) );
  AND2_X1 U24835 ( .A1(n24684), .A2(n24882), .ZN(n24880) );
  OR2_X1 U24836 ( .A1(n24688), .A2(n24689), .ZN(n24882) );
  OR2_X1 U24837 ( .A1(n15355), .A2(n15456), .ZN(n24689) );
  OR2_X1 U24838 ( .A1(n24883), .A2(n24884), .ZN(n24688) );
  AND2_X1 U24839 ( .A1(n24678), .A2(n24677), .ZN(n24884) );
  AND2_X1 U24840 ( .A1(n24673), .A2(n24885), .ZN(n24883) );
  OR2_X1 U24841 ( .A1(n24677), .A2(n24678), .ZN(n24885) );
  OR2_X1 U24842 ( .A1(n15321), .A2(n15456), .ZN(n24678) );
  OR2_X1 U24843 ( .A1(n24886), .A2(n24887), .ZN(n24677) );
  AND2_X1 U24844 ( .A1(n24668), .A2(n24667), .ZN(n24887) );
  AND2_X1 U24845 ( .A1(n24662), .A2(n24888), .ZN(n24886) );
  OR2_X1 U24846 ( .A1(n24667), .A2(n24668), .ZN(n24888) );
  OR2_X1 U24847 ( .A1(n15287), .A2(n15456), .ZN(n24668) );
  OR2_X1 U24848 ( .A1(n24889), .A2(n24890), .ZN(n24667) );
  AND2_X1 U24849 ( .A1(n24654), .A2(n24656), .ZN(n24890) );
  AND2_X1 U24850 ( .A1(n24651), .A2(n24891), .ZN(n24889) );
  OR2_X1 U24851 ( .A1(n24656), .A2(n24654), .ZN(n24891) );
  OR2_X1 U24852 ( .A1(n15242), .A2(n15456), .ZN(n24654) );
  OR2_X1 U24853 ( .A1(n24892), .A2(n24893), .ZN(n24656) );
  AND2_X1 U24854 ( .A1(n24643), .A2(n24645), .ZN(n24893) );
  AND2_X1 U24855 ( .A1(n24640), .A2(n24894), .ZN(n24892) );
  OR2_X1 U24856 ( .A1(n24645), .A2(n24643), .ZN(n24894) );
  OR2_X1 U24857 ( .A1(n15208), .A2(n15456), .ZN(n24643) );
  OR2_X1 U24858 ( .A1(n24895), .A2(n24896), .ZN(n24645) );
  AND2_X1 U24859 ( .A1(n24632), .A2(n24634), .ZN(n24896) );
  AND2_X1 U24860 ( .A1(n24629), .A2(n24897), .ZN(n24895) );
  OR2_X1 U24861 ( .A1(n24634), .A2(n24632), .ZN(n24897) );
  OR2_X1 U24862 ( .A1(n15174), .A2(n15456), .ZN(n24632) );
  OR2_X1 U24863 ( .A1(n24898), .A2(n24899), .ZN(n24634) );
  AND2_X1 U24864 ( .A1(n24621), .A2(n24623), .ZN(n24899) );
  AND2_X1 U24865 ( .A1(n24618), .A2(n24900), .ZN(n24898) );
  OR2_X1 U24866 ( .A1(n24623), .A2(n24621), .ZN(n24900) );
  OR2_X1 U24867 ( .A1(n15140), .A2(n15456), .ZN(n24621) );
  OR2_X1 U24868 ( .A1(n24901), .A2(n24902), .ZN(n24623) );
  AND2_X1 U24869 ( .A1(n24610), .A2(n24612), .ZN(n24902) );
  AND2_X1 U24870 ( .A1(n24607), .A2(n24903), .ZN(n24901) );
  OR2_X1 U24871 ( .A1(n24612), .A2(n24610), .ZN(n24903) );
  OR2_X1 U24872 ( .A1(n15106), .A2(n15456), .ZN(n24610) );
  OR2_X1 U24873 ( .A1(n24904), .A2(n24905), .ZN(n24612) );
  AND2_X1 U24874 ( .A1(n24599), .A2(n24601), .ZN(n24905) );
  AND2_X1 U24875 ( .A1(n24596), .A2(n24906), .ZN(n24904) );
  OR2_X1 U24876 ( .A1(n24601), .A2(n24599), .ZN(n24906) );
  OR2_X1 U24877 ( .A1(n15072), .A2(n15456), .ZN(n24599) );
  OR2_X1 U24878 ( .A1(n24907), .A2(n24908), .ZN(n24601) );
  AND2_X1 U24879 ( .A1(n24588), .A2(n24590), .ZN(n24908) );
  AND2_X1 U24880 ( .A1(n24585), .A2(n24909), .ZN(n24907) );
  OR2_X1 U24881 ( .A1(n24590), .A2(n24588), .ZN(n24909) );
  OR2_X1 U24882 ( .A1(n15038), .A2(n15456), .ZN(n24588) );
  OR2_X1 U24883 ( .A1(n24910), .A2(n24911), .ZN(n24590) );
  AND2_X1 U24884 ( .A1(n24577), .A2(n24579), .ZN(n24911) );
  AND2_X1 U24885 ( .A1(n24574), .A2(n24912), .ZN(n24910) );
  OR2_X1 U24886 ( .A1(n24579), .A2(n24577), .ZN(n24912) );
  OR2_X1 U24887 ( .A1(n15004), .A2(n15456), .ZN(n24577) );
  OR2_X1 U24888 ( .A1(n24913), .A2(n24914), .ZN(n24579) );
  AND2_X1 U24889 ( .A1(n24566), .A2(n24568), .ZN(n24914) );
  AND2_X1 U24890 ( .A1(n24563), .A2(n24915), .ZN(n24913) );
  OR2_X1 U24891 ( .A1(n24568), .A2(n24566), .ZN(n24915) );
  OR2_X1 U24892 ( .A1(n14970), .A2(n15456), .ZN(n24566) );
  OR2_X1 U24893 ( .A1(n24916), .A2(n24917), .ZN(n24568) );
  AND2_X1 U24894 ( .A1(n24555), .A2(n24557), .ZN(n24917) );
  AND2_X1 U24895 ( .A1(n24552), .A2(n24918), .ZN(n24916) );
  OR2_X1 U24896 ( .A1(n24557), .A2(n24555), .ZN(n24918) );
  OR2_X1 U24897 ( .A1(n14936), .A2(n15456), .ZN(n24555) );
  OR2_X1 U24898 ( .A1(n24919), .A2(n24920), .ZN(n24557) );
  AND2_X1 U24899 ( .A1(n24544), .A2(n24546), .ZN(n24920) );
  AND2_X1 U24900 ( .A1(n24541), .A2(n24921), .ZN(n24919) );
  OR2_X1 U24901 ( .A1(n24546), .A2(n24544), .ZN(n24921) );
  OR2_X1 U24902 ( .A1(n14891), .A2(n15456), .ZN(n24544) );
  OR2_X1 U24903 ( .A1(n24922), .A2(n24923), .ZN(n24546) );
  AND2_X1 U24904 ( .A1(n24529), .A2(n24534), .ZN(n24923) );
  AND2_X1 U24905 ( .A1(n24533), .A2(n24924), .ZN(n24922) );
  OR2_X1 U24906 ( .A1(n24534), .A2(n24529), .ZN(n24924) );
  OR2_X1 U24907 ( .A1(n14857), .A2(n15456), .ZN(n24529) );
  INV_X1 U24908 ( .A(b_12_), .ZN(n15456) );
  INV_X1 U24909 ( .A(n24535), .ZN(n24534) );
  AND3_X1 U24910 ( .A1(b_12_), .A2(b_11_), .A3(n15957), .ZN(n24535) );
  INV_X1 U24911 ( .A(n24536), .ZN(n24533) );
  OR2_X1 U24912 ( .A1(n24925), .A2(n24926), .ZN(n24536) );
  AND2_X1 U24913 ( .A1(b_11_), .A2(n24927), .ZN(n24926) );
  OR2_X1 U24914 ( .A1(n24928), .A2(n16981), .ZN(n24927) );
  AND2_X1 U24915 ( .A1(a_30_), .A2(n15524), .ZN(n24928) );
  AND2_X1 U24916 ( .A1(b_10_), .A2(n24929), .ZN(n24925) );
  OR2_X1 U24917 ( .A1(n24930), .A2(n14817), .ZN(n24929) );
  AND2_X1 U24918 ( .A1(a_31_), .A2(n15490), .ZN(n24930) );
  OR2_X1 U24919 ( .A1(n24931), .A2(n24932), .ZN(n24541) );
  AND2_X1 U24920 ( .A1(n24933), .A2(n24934), .ZN(n24932) );
  INV_X1 U24921 ( .A(n24935), .ZN(n24931) );
  OR2_X1 U24922 ( .A1(n24933), .A2(n24934), .ZN(n24935) );
  OR2_X1 U24923 ( .A1(n24936), .A2(n24937), .ZN(n24933) );
  AND2_X1 U24924 ( .A1(n24938), .A2(n24939), .ZN(n24937) );
  AND2_X1 U24925 ( .A1(n24940), .A2(n24941), .ZN(n24936) );
  OR2_X1 U24926 ( .A1(n24942), .A2(n24943), .ZN(n24552) );
  INV_X1 U24927 ( .A(n24944), .ZN(n24943) );
  OR2_X1 U24928 ( .A1(n24945), .A2(n24946), .ZN(n24944) );
  AND2_X1 U24929 ( .A1(n24946), .A2(n24945), .ZN(n24942) );
  AND2_X1 U24930 ( .A1(n24947), .A2(n24948), .ZN(n24945) );
  OR2_X1 U24931 ( .A1(n24949), .A2(n24950), .ZN(n24948) );
  INV_X1 U24932 ( .A(n24951), .ZN(n24950) );
  OR2_X1 U24933 ( .A1(n24951), .A2(n24952), .ZN(n24947) );
  INV_X1 U24934 ( .A(n24949), .ZN(n24952) );
  OR2_X1 U24935 ( .A1(n24953), .A2(n24954), .ZN(n24563) );
  INV_X1 U24936 ( .A(n24955), .ZN(n24954) );
  OR2_X1 U24937 ( .A1(n24956), .A2(n24957), .ZN(n24955) );
  AND2_X1 U24938 ( .A1(n24957), .A2(n24956), .ZN(n24953) );
  AND2_X1 U24939 ( .A1(n24958), .A2(n24959), .ZN(n24956) );
  OR2_X1 U24940 ( .A1(n24960), .A2(n24961), .ZN(n24959) );
  INV_X1 U24941 ( .A(n24962), .ZN(n24961) );
  OR2_X1 U24942 ( .A1(n24962), .A2(n24963), .ZN(n24958) );
  INV_X1 U24943 ( .A(n24960), .ZN(n24963) );
  OR2_X1 U24944 ( .A1(n24964), .A2(n24965), .ZN(n24574) );
  INV_X1 U24945 ( .A(n24966), .ZN(n24965) );
  OR2_X1 U24946 ( .A1(n24967), .A2(n24968), .ZN(n24966) );
  AND2_X1 U24947 ( .A1(n24968), .A2(n24967), .ZN(n24964) );
  AND2_X1 U24948 ( .A1(n24969), .A2(n24970), .ZN(n24967) );
  OR2_X1 U24949 ( .A1(n24971), .A2(n24972), .ZN(n24970) );
  INV_X1 U24950 ( .A(n24973), .ZN(n24972) );
  OR2_X1 U24951 ( .A1(n24973), .A2(n24974), .ZN(n24969) );
  INV_X1 U24952 ( .A(n24971), .ZN(n24974) );
  OR2_X1 U24953 ( .A1(n24975), .A2(n24976), .ZN(n24585) );
  INV_X1 U24954 ( .A(n24977), .ZN(n24976) );
  OR2_X1 U24955 ( .A1(n24978), .A2(n24979), .ZN(n24977) );
  AND2_X1 U24956 ( .A1(n24979), .A2(n24978), .ZN(n24975) );
  AND2_X1 U24957 ( .A1(n24980), .A2(n24981), .ZN(n24978) );
  OR2_X1 U24958 ( .A1(n24982), .A2(n24983), .ZN(n24981) );
  INV_X1 U24959 ( .A(n24984), .ZN(n24983) );
  OR2_X1 U24960 ( .A1(n24984), .A2(n24985), .ZN(n24980) );
  INV_X1 U24961 ( .A(n24982), .ZN(n24985) );
  OR2_X1 U24962 ( .A1(n24986), .A2(n24987), .ZN(n24596) );
  INV_X1 U24963 ( .A(n24988), .ZN(n24987) );
  OR2_X1 U24964 ( .A1(n24989), .A2(n24990), .ZN(n24988) );
  AND2_X1 U24965 ( .A1(n24990), .A2(n24989), .ZN(n24986) );
  AND2_X1 U24966 ( .A1(n24991), .A2(n24992), .ZN(n24989) );
  OR2_X1 U24967 ( .A1(n24993), .A2(n24994), .ZN(n24992) );
  INV_X1 U24968 ( .A(n24995), .ZN(n24994) );
  OR2_X1 U24969 ( .A1(n24995), .A2(n24996), .ZN(n24991) );
  INV_X1 U24970 ( .A(n24993), .ZN(n24996) );
  OR2_X1 U24971 ( .A1(n24997), .A2(n24998), .ZN(n24607) );
  INV_X1 U24972 ( .A(n24999), .ZN(n24998) );
  OR2_X1 U24973 ( .A1(n25000), .A2(n25001), .ZN(n24999) );
  AND2_X1 U24974 ( .A1(n25001), .A2(n25000), .ZN(n24997) );
  AND2_X1 U24975 ( .A1(n25002), .A2(n25003), .ZN(n25000) );
  OR2_X1 U24976 ( .A1(n25004), .A2(n25005), .ZN(n25003) );
  INV_X1 U24977 ( .A(n25006), .ZN(n25005) );
  OR2_X1 U24978 ( .A1(n25006), .A2(n25007), .ZN(n25002) );
  INV_X1 U24979 ( .A(n25004), .ZN(n25007) );
  OR2_X1 U24980 ( .A1(n25008), .A2(n25009), .ZN(n24618) );
  INV_X1 U24981 ( .A(n25010), .ZN(n25009) );
  OR2_X1 U24982 ( .A1(n25011), .A2(n25012), .ZN(n25010) );
  AND2_X1 U24983 ( .A1(n25012), .A2(n25011), .ZN(n25008) );
  AND2_X1 U24984 ( .A1(n25013), .A2(n25014), .ZN(n25011) );
  OR2_X1 U24985 ( .A1(n25015), .A2(n25016), .ZN(n25014) );
  INV_X1 U24986 ( .A(n25017), .ZN(n25016) );
  OR2_X1 U24987 ( .A1(n25017), .A2(n25018), .ZN(n25013) );
  INV_X1 U24988 ( .A(n25015), .ZN(n25018) );
  OR2_X1 U24989 ( .A1(n25019), .A2(n25020), .ZN(n24629) );
  INV_X1 U24990 ( .A(n25021), .ZN(n25020) );
  OR2_X1 U24991 ( .A1(n25022), .A2(n25023), .ZN(n25021) );
  AND2_X1 U24992 ( .A1(n25023), .A2(n25022), .ZN(n25019) );
  AND2_X1 U24993 ( .A1(n25024), .A2(n25025), .ZN(n25022) );
  OR2_X1 U24994 ( .A1(n25026), .A2(n25027), .ZN(n25025) );
  INV_X1 U24995 ( .A(n25028), .ZN(n25027) );
  OR2_X1 U24996 ( .A1(n25028), .A2(n25029), .ZN(n25024) );
  INV_X1 U24997 ( .A(n25026), .ZN(n25029) );
  OR2_X1 U24998 ( .A1(n25030), .A2(n25031), .ZN(n24640) );
  INV_X1 U24999 ( .A(n25032), .ZN(n25031) );
  OR2_X1 U25000 ( .A1(n25033), .A2(n25034), .ZN(n25032) );
  AND2_X1 U25001 ( .A1(n25034), .A2(n25033), .ZN(n25030) );
  AND2_X1 U25002 ( .A1(n25035), .A2(n25036), .ZN(n25033) );
  OR2_X1 U25003 ( .A1(n25037), .A2(n25038), .ZN(n25036) );
  INV_X1 U25004 ( .A(n25039), .ZN(n25038) );
  OR2_X1 U25005 ( .A1(n25039), .A2(n25040), .ZN(n25035) );
  INV_X1 U25006 ( .A(n25037), .ZN(n25040) );
  OR2_X1 U25007 ( .A1(n25041), .A2(n25042), .ZN(n24651) );
  INV_X1 U25008 ( .A(n25043), .ZN(n25042) );
  OR2_X1 U25009 ( .A1(n25044), .A2(n25045), .ZN(n25043) );
  AND2_X1 U25010 ( .A1(n25045), .A2(n25044), .ZN(n25041) );
  AND2_X1 U25011 ( .A1(n25046), .A2(n25047), .ZN(n25044) );
  OR2_X1 U25012 ( .A1(n25048), .A2(n25049), .ZN(n25047) );
  INV_X1 U25013 ( .A(n25050), .ZN(n25049) );
  OR2_X1 U25014 ( .A1(n25050), .A2(n25051), .ZN(n25046) );
  INV_X1 U25015 ( .A(n25048), .ZN(n25051) );
  OR2_X1 U25016 ( .A1(n25052), .A2(n25053), .ZN(n24662) );
  INV_X1 U25017 ( .A(n25054), .ZN(n25053) );
  OR2_X1 U25018 ( .A1(n25055), .A2(n25056), .ZN(n25054) );
  AND2_X1 U25019 ( .A1(n25056), .A2(n25055), .ZN(n25052) );
  AND2_X1 U25020 ( .A1(n25057), .A2(n25058), .ZN(n25055) );
  INV_X1 U25021 ( .A(n25059), .ZN(n25058) );
  AND2_X1 U25022 ( .A1(n25060), .A2(n25061), .ZN(n25059) );
  OR2_X1 U25023 ( .A1(n25061), .A2(n25060), .ZN(n25057) );
  INV_X1 U25024 ( .A(n25062), .ZN(n25060) );
  AND2_X1 U25025 ( .A1(n25063), .A2(n25064), .ZN(n24673) );
  INV_X1 U25026 ( .A(n25065), .ZN(n25064) );
  AND2_X1 U25027 ( .A1(n25066), .A2(n25067), .ZN(n25065) );
  OR2_X1 U25028 ( .A1(n25067), .A2(n25066), .ZN(n25063) );
  OR2_X1 U25029 ( .A1(n25068), .A2(n25069), .ZN(n25066) );
  AND2_X1 U25030 ( .A1(n25070), .A2(n25071), .ZN(n25069) );
  INV_X1 U25031 ( .A(n25072), .ZN(n25070) );
  AND2_X1 U25032 ( .A1(n25073), .A2(n25072), .ZN(n25068) );
  INV_X1 U25033 ( .A(n25071), .ZN(n25073) );
  AND2_X1 U25034 ( .A1(n25074), .A2(n25075), .ZN(n24684) );
  INV_X1 U25035 ( .A(n25076), .ZN(n25075) );
  AND2_X1 U25036 ( .A1(n25077), .A2(n25078), .ZN(n25076) );
  OR2_X1 U25037 ( .A1(n25078), .A2(n25077), .ZN(n25074) );
  OR2_X1 U25038 ( .A1(n25079), .A2(n25080), .ZN(n25077) );
  AND2_X1 U25039 ( .A1(n25081), .A2(n25082), .ZN(n25080) );
  INV_X1 U25040 ( .A(n25083), .ZN(n25081) );
  AND2_X1 U25041 ( .A1(n25084), .A2(n25083), .ZN(n25079) );
  INV_X1 U25042 ( .A(n25082), .ZN(n25084) );
  AND2_X1 U25043 ( .A1(n25085), .A2(n25086), .ZN(n24695) );
  INV_X1 U25044 ( .A(n25087), .ZN(n25086) );
  AND2_X1 U25045 ( .A1(n25088), .A2(n25089), .ZN(n25087) );
  OR2_X1 U25046 ( .A1(n25089), .A2(n25088), .ZN(n25085) );
  OR2_X1 U25047 ( .A1(n25090), .A2(n25091), .ZN(n25088) );
  AND2_X1 U25048 ( .A1(n25092), .A2(n25093), .ZN(n25091) );
  INV_X1 U25049 ( .A(n25094), .ZN(n25092) );
  AND2_X1 U25050 ( .A1(n25095), .A2(n25094), .ZN(n25090) );
  INV_X1 U25051 ( .A(n25093), .ZN(n25095) );
  AND2_X1 U25052 ( .A1(n25096), .A2(n25097), .ZN(n24706) );
  INV_X1 U25053 ( .A(n25098), .ZN(n25097) );
  AND2_X1 U25054 ( .A1(n25099), .A2(n25100), .ZN(n25098) );
  OR2_X1 U25055 ( .A1(n25100), .A2(n25099), .ZN(n25096) );
  OR2_X1 U25056 ( .A1(n25101), .A2(n25102), .ZN(n25099) );
  AND2_X1 U25057 ( .A1(n25103), .A2(n25104), .ZN(n25102) );
  INV_X1 U25058 ( .A(n25105), .ZN(n25103) );
  AND2_X1 U25059 ( .A1(n25106), .A2(n25105), .ZN(n25101) );
  INV_X1 U25060 ( .A(n25104), .ZN(n25106) );
  AND2_X1 U25061 ( .A1(n25107), .A2(n25108), .ZN(n24717) );
  INV_X1 U25062 ( .A(n25109), .ZN(n25108) );
  AND2_X1 U25063 ( .A1(n25110), .A2(n25111), .ZN(n25109) );
  OR2_X1 U25064 ( .A1(n25111), .A2(n25110), .ZN(n25107) );
  OR2_X1 U25065 ( .A1(n25112), .A2(n25113), .ZN(n25110) );
  AND2_X1 U25066 ( .A1(n25114), .A2(n25115), .ZN(n25113) );
  INV_X1 U25067 ( .A(n25116), .ZN(n25114) );
  AND2_X1 U25068 ( .A1(n25117), .A2(n25116), .ZN(n25112) );
  INV_X1 U25069 ( .A(n25115), .ZN(n25117) );
  AND2_X1 U25070 ( .A1(n25118), .A2(n25119), .ZN(n24727) );
  INV_X1 U25071 ( .A(n25120), .ZN(n25119) );
  AND2_X1 U25072 ( .A1(n25121), .A2(n25122), .ZN(n25120) );
  OR2_X1 U25073 ( .A1(n25122), .A2(n25121), .ZN(n25118) );
  OR2_X1 U25074 ( .A1(n25123), .A2(n25124), .ZN(n25121) );
  AND2_X1 U25075 ( .A1(n25125), .A2(n25126), .ZN(n25124) );
  INV_X1 U25076 ( .A(n25127), .ZN(n25125) );
  AND2_X1 U25077 ( .A1(n25128), .A2(n25127), .ZN(n25123) );
  INV_X1 U25078 ( .A(n25126), .ZN(n25128) );
  AND2_X1 U25079 ( .A1(n25129), .A2(n25130), .ZN(n24738) );
  INV_X1 U25080 ( .A(n25131), .ZN(n25130) );
  AND2_X1 U25081 ( .A1(n25132), .A2(n25133), .ZN(n25131) );
  OR2_X1 U25082 ( .A1(n25133), .A2(n25132), .ZN(n25129) );
  OR2_X1 U25083 ( .A1(n25134), .A2(n25135), .ZN(n25132) );
  AND2_X1 U25084 ( .A1(n25136), .A2(n25137), .ZN(n25135) );
  INV_X1 U25085 ( .A(n15900), .ZN(n25136) );
  AND2_X1 U25086 ( .A1(n25138), .A2(n15900), .ZN(n25134) );
  INV_X1 U25087 ( .A(n25137), .ZN(n25138) );
  AND2_X1 U25088 ( .A1(n25139), .A2(n25140), .ZN(n24749) );
  INV_X1 U25089 ( .A(n25141), .ZN(n25140) );
  AND2_X1 U25090 ( .A1(n25142), .A2(n25143), .ZN(n25141) );
  OR2_X1 U25091 ( .A1(n25143), .A2(n25142), .ZN(n25139) );
  OR2_X1 U25092 ( .A1(n25144), .A2(n25145), .ZN(n25142) );
  AND2_X1 U25093 ( .A1(n25146), .A2(n25147), .ZN(n25145) );
  INV_X1 U25094 ( .A(n25148), .ZN(n25146) );
  AND2_X1 U25095 ( .A1(n25149), .A2(n25148), .ZN(n25144) );
  INV_X1 U25096 ( .A(n25147), .ZN(n25149) );
  AND2_X1 U25097 ( .A1(n25150), .A2(n25151), .ZN(n24760) );
  INV_X1 U25098 ( .A(n25152), .ZN(n25151) );
  AND2_X1 U25099 ( .A1(n25153), .A2(n25154), .ZN(n25152) );
  OR2_X1 U25100 ( .A1(n25154), .A2(n25153), .ZN(n25150) );
  OR2_X1 U25101 ( .A1(n25155), .A2(n25156), .ZN(n25153) );
  AND2_X1 U25102 ( .A1(n25157), .A2(n25158), .ZN(n25156) );
  INV_X1 U25103 ( .A(n25159), .ZN(n25157) );
  AND2_X1 U25104 ( .A1(n25160), .A2(n25159), .ZN(n25155) );
  INV_X1 U25105 ( .A(n25158), .ZN(n25160) );
  AND2_X1 U25106 ( .A1(n25161), .A2(n25162), .ZN(n24771) );
  INV_X1 U25107 ( .A(n25163), .ZN(n25162) );
  AND2_X1 U25108 ( .A1(n25164), .A2(n25165), .ZN(n25163) );
  OR2_X1 U25109 ( .A1(n25165), .A2(n25164), .ZN(n25161) );
  OR2_X1 U25110 ( .A1(n25166), .A2(n25167), .ZN(n25164) );
  AND2_X1 U25111 ( .A1(n25168), .A2(n25169), .ZN(n25167) );
  INV_X1 U25112 ( .A(n25170), .ZN(n25168) );
  AND2_X1 U25113 ( .A1(n25171), .A2(n25170), .ZN(n25166) );
  INV_X1 U25114 ( .A(n25169), .ZN(n25171) );
  AND2_X1 U25115 ( .A1(n25172), .A2(n25173), .ZN(n24782) );
  INV_X1 U25116 ( .A(n25174), .ZN(n25173) );
  AND2_X1 U25117 ( .A1(n25175), .A2(n25176), .ZN(n25174) );
  OR2_X1 U25118 ( .A1(n25176), .A2(n25175), .ZN(n25172) );
  OR2_X1 U25119 ( .A1(n25177), .A2(n25178), .ZN(n25175) );
  AND2_X1 U25120 ( .A1(n25179), .A2(n25180), .ZN(n25178) );
  INV_X1 U25121 ( .A(n25181), .ZN(n25179) );
  AND2_X1 U25122 ( .A1(n25182), .A2(n25181), .ZN(n25177) );
  INV_X1 U25123 ( .A(n25180), .ZN(n25182) );
  AND2_X1 U25124 ( .A1(n25183), .A2(n25184), .ZN(n24793) );
  INV_X1 U25125 ( .A(n25185), .ZN(n25184) );
  AND2_X1 U25126 ( .A1(n25186), .A2(n25187), .ZN(n25185) );
  OR2_X1 U25127 ( .A1(n25187), .A2(n25186), .ZN(n25183) );
  OR2_X1 U25128 ( .A1(n25188), .A2(n25189), .ZN(n25186) );
  AND2_X1 U25129 ( .A1(n25190), .A2(n25191), .ZN(n25189) );
  INV_X1 U25130 ( .A(n25192), .ZN(n25190) );
  AND2_X1 U25131 ( .A1(n25193), .A2(n25192), .ZN(n25188) );
  INV_X1 U25132 ( .A(n25191), .ZN(n25193) );
  AND2_X1 U25133 ( .A1(n25194), .A2(n25195), .ZN(n24804) );
  INV_X1 U25134 ( .A(n25196), .ZN(n25195) );
  AND2_X1 U25135 ( .A1(n25197), .A2(n25198), .ZN(n25196) );
  OR2_X1 U25136 ( .A1(n25198), .A2(n25197), .ZN(n25194) );
  OR2_X1 U25137 ( .A1(n25199), .A2(n25200), .ZN(n25197) );
  AND2_X1 U25138 ( .A1(n25201), .A2(n25202), .ZN(n25200) );
  INV_X1 U25139 ( .A(n25203), .ZN(n25201) );
  AND2_X1 U25140 ( .A1(n25204), .A2(n25203), .ZN(n25199) );
  INV_X1 U25141 ( .A(n25202), .ZN(n25204) );
  AND2_X1 U25142 ( .A1(n25205), .A2(n25206), .ZN(n24815) );
  INV_X1 U25143 ( .A(n25207), .ZN(n25206) );
  AND2_X1 U25144 ( .A1(n25208), .A2(n25209), .ZN(n25207) );
  OR2_X1 U25145 ( .A1(n25209), .A2(n25208), .ZN(n25205) );
  OR2_X1 U25146 ( .A1(n25210), .A2(n25211), .ZN(n25208) );
  AND2_X1 U25147 ( .A1(n25212), .A2(n25213), .ZN(n25211) );
  INV_X1 U25148 ( .A(n25214), .ZN(n25212) );
  AND2_X1 U25149 ( .A1(n25215), .A2(n25214), .ZN(n25210) );
  INV_X1 U25150 ( .A(n25213), .ZN(n25215) );
  AND2_X1 U25151 ( .A1(n25216), .A2(n25217), .ZN(n24826) );
  INV_X1 U25152 ( .A(n25218), .ZN(n25217) );
  AND2_X1 U25153 ( .A1(n25219), .A2(n25220), .ZN(n25218) );
  OR2_X1 U25154 ( .A1(n25220), .A2(n25219), .ZN(n25216) );
  OR2_X1 U25155 ( .A1(n25221), .A2(n25222), .ZN(n25219) );
  AND2_X1 U25156 ( .A1(n25223), .A2(n25224), .ZN(n25222) );
  INV_X1 U25157 ( .A(n25225), .ZN(n25223) );
  AND2_X1 U25158 ( .A1(n25226), .A2(n25225), .ZN(n25221) );
  INV_X1 U25159 ( .A(n25224), .ZN(n25226) );
  AND2_X1 U25160 ( .A1(n25227), .A2(n25228), .ZN(n16605) );
  INV_X1 U25161 ( .A(n25229), .ZN(n25228) );
  AND2_X1 U25162 ( .A1(n25230), .A2(n16619), .ZN(n25229) );
  OR2_X1 U25163 ( .A1(n16619), .A2(n25230), .ZN(n25227) );
  OR2_X1 U25164 ( .A1(n25231), .A2(n25232), .ZN(n25230) );
  AND2_X1 U25165 ( .A1(n25233), .A2(n16618), .ZN(n25232) );
  INV_X1 U25166 ( .A(n16617), .ZN(n25233) );
  AND2_X1 U25167 ( .A1(n25234), .A2(n16617), .ZN(n25231) );
  OR2_X1 U25168 ( .A1(n15808), .A2(n15490), .ZN(n16617) );
  INV_X1 U25169 ( .A(n16618), .ZN(n25234) );
  OR2_X1 U25170 ( .A1(n25235), .A2(n25236), .ZN(n16618) );
  AND2_X1 U25171 ( .A1(n25225), .A2(n25224), .ZN(n25236) );
  AND2_X1 U25172 ( .A1(n25220), .A2(n25237), .ZN(n25235) );
  OR2_X1 U25173 ( .A1(n25225), .A2(n25224), .ZN(n25237) );
  OR2_X1 U25174 ( .A1(n25238), .A2(n25239), .ZN(n25224) );
  AND2_X1 U25175 ( .A1(n25214), .A2(n25213), .ZN(n25239) );
  AND2_X1 U25176 ( .A1(n25209), .A2(n25240), .ZN(n25238) );
  OR2_X1 U25177 ( .A1(n25214), .A2(n25213), .ZN(n25240) );
  OR2_X1 U25178 ( .A1(n25241), .A2(n25242), .ZN(n25213) );
  AND2_X1 U25179 ( .A1(n25203), .A2(n25202), .ZN(n25242) );
  AND2_X1 U25180 ( .A1(n25198), .A2(n25243), .ZN(n25241) );
  OR2_X1 U25181 ( .A1(n25203), .A2(n25202), .ZN(n25243) );
  OR2_X1 U25182 ( .A1(n25244), .A2(n25245), .ZN(n25202) );
  AND2_X1 U25183 ( .A1(n25192), .A2(n25191), .ZN(n25245) );
  AND2_X1 U25184 ( .A1(n25187), .A2(n25246), .ZN(n25244) );
  OR2_X1 U25185 ( .A1(n25192), .A2(n25191), .ZN(n25246) );
  OR2_X1 U25186 ( .A1(n25247), .A2(n25248), .ZN(n25191) );
  AND2_X1 U25187 ( .A1(n25181), .A2(n25180), .ZN(n25248) );
  AND2_X1 U25188 ( .A1(n25176), .A2(n25249), .ZN(n25247) );
  OR2_X1 U25189 ( .A1(n25181), .A2(n25180), .ZN(n25249) );
  OR2_X1 U25190 ( .A1(n25250), .A2(n25251), .ZN(n25180) );
  AND2_X1 U25191 ( .A1(n25170), .A2(n25169), .ZN(n25251) );
  AND2_X1 U25192 ( .A1(n25165), .A2(n25252), .ZN(n25250) );
  OR2_X1 U25193 ( .A1(n25170), .A2(n25169), .ZN(n25252) );
  OR2_X1 U25194 ( .A1(n25253), .A2(n25254), .ZN(n25169) );
  AND2_X1 U25195 ( .A1(n25159), .A2(n25158), .ZN(n25254) );
  AND2_X1 U25196 ( .A1(n25154), .A2(n25255), .ZN(n25253) );
  OR2_X1 U25197 ( .A1(n25159), .A2(n25158), .ZN(n25255) );
  OR2_X1 U25198 ( .A1(n25256), .A2(n25257), .ZN(n25158) );
  AND2_X1 U25199 ( .A1(n25148), .A2(n25147), .ZN(n25257) );
  AND2_X1 U25200 ( .A1(n25143), .A2(n25258), .ZN(n25256) );
  OR2_X1 U25201 ( .A1(n25148), .A2(n25147), .ZN(n25258) );
  OR2_X1 U25202 ( .A1(n25259), .A2(n25260), .ZN(n25147) );
  AND2_X1 U25203 ( .A1(n15900), .A2(n25137), .ZN(n25260) );
  AND2_X1 U25204 ( .A1(n25133), .A2(n25261), .ZN(n25259) );
  OR2_X1 U25205 ( .A1(n15900), .A2(n25137), .ZN(n25261) );
  OR2_X1 U25206 ( .A1(n25262), .A2(n25263), .ZN(n25137) );
  AND2_X1 U25207 ( .A1(n25127), .A2(n25126), .ZN(n25263) );
  AND2_X1 U25208 ( .A1(n25122), .A2(n25264), .ZN(n25262) );
  OR2_X1 U25209 ( .A1(n25127), .A2(n25126), .ZN(n25264) );
  OR2_X1 U25210 ( .A1(n25265), .A2(n25266), .ZN(n25126) );
  AND2_X1 U25211 ( .A1(n25116), .A2(n25115), .ZN(n25266) );
  AND2_X1 U25212 ( .A1(n25111), .A2(n25267), .ZN(n25265) );
  OR2_X1 U25213 ( .A1(n25116), .A2(n25115), .ZN(n25267) );
  OR2_X1 U25214 ( .A1(n25268), .A2(n25269), .ZN(n25115) );
  AND2_X1 U25215 ( .A1(n25105), .A2(n25104), .ZN(n25269) );
  AND2_X1 U25216 ( .A1(n25100), .A2(n25270), .ZN(n25268) );
  OR2_X1 U25217 ( .A1(n25105), .A2(n25104), .ZN(n25270) );
  OR2_X1 U25218 ( .A1(n25271), .A2(n25272), .ZN(n25104) );
  AND2_X1 U25219 ( .A1(n25094), .A2(n25093), .ZN(n25272) );
  AND2_X1 U25220 ( .A1(n25089), .A2(n25273), .ZN(n25271) );
  OR2_X1 U25221 ( .A1(n25094), .A2(n25093), .ZN(n25273) );
  OR2_X1 U25222 ( .A1(n25274), .A2(n25275), .ZN(n25093) );
  AND2_X1 U25223 ( .A1(n25083), .A2(n25082), .ZN(n25275) );
  AND2_X1 U25224 ( .A1(n25078), .A2(n25276), .ZN(n25274) );
  OR2_X1 U25225 ( .A1(n25083), .A2(n25082), .ZN(n25276) );
  OR2_X1 U25226 ( .A1(n25277), .A2(n25278), .ZN(n25082) );
  AND2_X1 U25227 ( .A1(n25072), .A2(n25071), .ZN(n25278) );
  AND2_X1 U25228 ( .A1(n25067), .A2(n25279), .ZN(n25277) );
  OR2_X1 U25229 ( .A1(n25072), .A2(n25071), .ZN(n25279) );
  OR2_X1 U25230 ( .A1(n25280), .A2(n25281), .ZN(n25071) );
  AND2_X1 U25231 ( .A1(n25062), .A2(n25061), .ZN(n25281) );
  AND2_X1 U25232 ( .A1(n25056), .A2(n25282), .ZN(n25280) );
  OR2_X1 U25233 ( .A1(n25062), .A2(n25061), .ZN(n25282) );
  OR2_X1 U25234 ( .A1(n25283), .A2(n25284), .ZN(n25061) );
  AND2_X1 U25235 ( .A1(n25048), .A2(n25050), .ZN(n25284) );
  AND2_X1 U25236 ( .A1(n25045), .A2(n25285), .ZN(n25283) );
  OR2_X1 U25237 ( .A1(n25048), .A2(n25050), .ZN(n25285) );
  OR2_X1 U25238 ( .A1(n25286), .A2(n25287), .ZN(n25050) );
  AND2_X1 U25239 ( .A1(n25037), .A2(n25039), .ZN(n25287) );
  AND2_X1 U25240 ( .A1(n25034), .A2(n25288), .ZN(n25286) );
  OR2_X1 U25241 ( .A1(n25037), .A2(n25039), .ZN(n25288) );
  OR2_X1 U25242 ( .A1(n25289), .A2(n25290), .ZN(n25039) );
  AND2_X1 U25243 ( .A1(n25026), .A2(n25028), .ZN(n25290) );
  AND2_X1 U25244 ( .A1(n25023), .A2(n25291), .ZN(n25289) );
  OR2_X1 U25245 ( .A1(n25026), .A2(n25028), .ZN(n25291) );
  OR2_X1 U25246 ( .A1(n25292), .A2(n25293), .ZN(n25028) );
  AND2_X1 U25247 ( .A1(n25015), .A2(n25017), .ZN(n25293) );
  AND2_X1 U25248 ( .A1(n25012), .A2(n25294), .ZN(n25292) );
  OR2_X1 U25249 ( .A1(n25015), .A2(n25017), .ZN(n25294) );
  OR2_X1 U25250 ( .A1(n25295), .A2(n25296), .ZN(n25017) );
  AND2_X1 U25251 ( .A1(n25004), .A2(n25006), .ZN(n25296) );
  AND2_X1 U25252 ( .A1(n25001), .A2(n25297), .ZN(n25295) );
  OR2_X1 U25253 ( .A1(n25004), .A2(n25006), .ZN(n25297) );
  OR2_X1 U25254 ( .A1(n25298), .A2(n25299), .ZN(n25006) );
  AND2_X1 U25255 ( .A1(n24993), .A2(n24995), .ZN(n25299) );
  AND2_X1 U25256 ( .A1(n24990), .A2(n25300), .ZN(n25298) );
  OR2_X1 U25257 ( .A1(n24993), .A2(n24995), .ZN(n25300) );
  OR2_X1 U25258 ( .A1(n25301), .A2(n25302), .ZN(n24995) );
  AND2_X1 U25259 ( .A1(n24982), .A2(n24984), .ZN(n25302) );
  AND2_X1 U25260 ( .A1(n24979), .A2(n25303), .ZN(n25301) );
  OR2_X1 U25261 ( .A1(n24982), .A2(n24984), .ZN(n25303) );
  OR2_X1 U25262 ( .A1(n25304), .A2(n25305), .ZN(n24984) );
  AND2_X1 U25263 ( .A1(n24971), .A2(n24973), .ZN(n25305) );
  AND2_X1 U25264 ( .A1(n24968), .A2(n25306), .ZN(n25304) );
  OR2_X1 U25265 ( .A1(n24971), .A2(n24973), .ZN(n25306) );
  OR2_X1 U25266 ( .A1(n25307), .A2(n25308), .ZN(n24973) );
  AND2_X1 U25267 ( .A1(n24960), .A2(n24962), .ZN(n25308) );
  AND2_X1 U25268 ( .A1(n24957), .A2(n25309), .ZN(n25307) );
  OR2_X1 U25269 ( .A1(n24960), .A2(n24962), .ZN(n25309) );
  OR2_X1 U25270 ( .A1(n25310), .A2(n25311), .ZN(n24962) );
  AND2_X1 U25271 ( .A1(n24949), .A2(n24951), .ZN(n25311) );
  AND2_X1 U25272 ( .A1(n24946), .A2(n25312), .ZN(n25310) );
  OR2_X1 U25273 ( .A1(n24949), .A2(n24951), .ZN(n25312) );
  OR2_X1 U25274 ( .A1(n25313), .A2(n25314), .ZN(n24951) );
  AND2_X1 U25275 ( .A1(n24934), .A2(n24939), .ZN(n25314) );
  AND2_X1 U25276 ( .A1(n24938), .A2(n25315), .ZN(n25313) );
  OR2_X1 U25277 ( .A1(n24934), .A2(n24939), .ZN(n25315) );
  INV_X1 U25278 ( .A(n24940), .ZN(n24939) );
  AND3_X1 U25279 ( .A1(b_11_), .A2(b_10_), .A3(n15957), .ZN(n24940) );
  OR2_X1 U25280 ( .A1(n14857), .A2(n15490), .ZN(n24934) );
  INV_X1 U25281 ( .A(n24941), .ZN(n24938) );
  OR2_X1 U25282 ( .A1(n25316), .A2(n25317), .ZN(n24941) );
  AND2_X1 U25283 ( .A1(b_9_), .A2(n25318), .ZN(n25317) );
  OR2_X1 U25284 ( .A1(n25319), .A2(n14817), .ZN(n25318) );
  AND2_X1 U25285 ( .A1(a_31_), .A2(n15524), .ZN(n25319) );
  AND2_X1 U25286 ( .A1(b_10_), .A2(n25320), .ZN(n25316) );
  OR2_X1 U25287 ( .A1(n25321), .A2(n16981), .ZN(n25320) );
  AND2_X1 U25288 ( .A1(a_30_), .A2(n15558), .ZN(n25321) );
  OR2_X1 U25289 ( .A1(n14891), .A2(n15490), .ZN(n24949) );
  OR2_X1 U25290 ( .A1(n25322), .A2(n25323), .ZN(n24946) );
  AND2_X1 U25291 ( .A1(n25324), .A2(n25325), .ZN(n25323) );
  INV_X1 U25292 ( .A(n25326), .ZN(n25322) );
  OR2_X1 U25293 ( .A1(n25324), .A2(n25325), .ZN(n25326) );
  OR2_X1 U25294 ( .A1(n25327), .A2(n25328), .ZN(n25324) );
  AND2_X1 U25295 ( .A1(n25329), .A2(n25330), .ZN(n25328) );
  AND2_X1 U25296 ( .A1(n25331), .A2(n25332), .ZN(n25327) );
  OR2_X1 U25297 ( .A1(n14936), .A2(n15490), .ZN(n24960) );
  OR2_X1 U25298 ( .A1(n25333), .A2(n25334), .ZN(n24957) );
  INV_X1 U25299 ( .A(n25335), .ZN(n25334) );
  OR2_X1 U25300 ( .A1(n25336), .A2(n25337), .ZN(n25335) );
  AND2_X1 U25301 ( .A1(n25337), .A2(n25336), .ZN(n25333) );
  AND2_X1 U25302 ( .A1(n25338), .A2(n25339), .ZN(n25336) );
  OR2_X1 U25303 ( .A1(n25340), .A2(n25341), .ZN(n25339) );
  INV_X1 U25304 ( .A(n25342), .ZN(n25341) );
  OR2_X1 U25305 ( .A1(n25342), .A2(n25343), .ZN(n25338) );
  INV_X1 U25306 ( .A(n25340), .ZN(n25343) );
  OR2_X1 U25307 ( .A1(n14970), .A2(n15490), .ZN(n24971) );
  OR2_X1 U25308 ( .A1(n25344), .A2(n25345), .ZN(n24968) );
  INV_X1 U25309 ( .A(n25346), .ZN(n25345) );
  OR2_X1 U25310 ( .A1(n25347), .A2(n25348), .ZN(n25346) );
  AND2_X1 U25311 ( .A1(n25348), .A2(n25347), .ZN(n25344) );
  AND2_X1 U25312 ( .A1(n25349), .A2(n25350), .ZN(n25347) );
  OR2_X1 U25313 ( .A1(n25351), .A2(n25352), .ZN(n25350) );
  INV_X1 U25314 ( .A(n25353), .ZN(n25352) );
  OR2_X1 U25315 ( .A1(n25353), .A2(n25354), .ZN(n25349) );
  INV_X1 U25316 ( .A(n25351), .ZN(n25354) );
  OR2_X1 U25317 ( .A1(n15004), .A2(n15490), .ZN(n24982) );
  OR2_X1 U25318 ( .A1(n25355), .A2(n25356), .ZN(n24979) );
  INV_X1 U25319 ( .A(n25357), .ZN(n25356) );
  OR2_X1 U25320 ( .A1(n25358), .A2(n25359), .ZN(n25357) );
  AND2_X1 U25321 ( .A1(n25359), .A2(n25358), .ZN(n25355) );
  AND2_X1 U25322 ( .A1(n25360), .A2(n25361), .ZN(n25358) );
  OR2_X1 U25323 ( .A1(n25362), .A2(n25363), .ZN(n25361) );
  INV_X1 U25324 ( .A(n25364), .ZN(n25363) );
  OR2_X1 U25325 ( .A1(n25364), .A2(n25365), .ZN(n25360) );
  INV_X1 U25326 ( .A(n25362), .ZN(n25365) );
  OR2_X1 U25327 ( .A1(n15038), .A2(n15490), .ZN(n24993) );
  OR2_X1 U25328 ( .A1(n25366), .A2(n25367), .ZN(n24990) );
  INV_X1 U25329 ( .A(n25368), .ZN(n25367) );
  OR2_X1 U25330 ( .A1(n25369), .A2(n25370), .ZN(n25368) );
  AND2_X1 U25331 ( .A1(n25370), .A2(n25369), .ZN(n25366) );
  AND2_X1 U25332 ( .A1(n25371), .A2(n25372), .ZN(n25369) );
  OR2_X1 U25333 ( .A1(n25373), .A2(n25374), .ZN(n25372) );
  INV_X1 U25334 ( .A(n25375), .ZN(n25374) );
  OR2_X1 U25335 ( .A1(n25375), .A2(n25376), .ZN(n25371) );
  INV_X1 U25336 ( .A(n25373), .ZN(n25376) );
  OR2_X1 U25337 ( .A1(n15072), .A2(n15490), .ZN(n25004) );
  OR2_X1 U25338 ( .A1(n25377), .A2(n25378), .ZN(n25001) );
  INV_X1 U25339 ( .A(n25379), .ZN(n25378) );
  OR2_X1 U25340 ( .A1(n25380), .A2(n25381), .ZN(n25379) );
  AND2_X1 U25341 ( .A1(n25381), .A2(n25380), .ZN(n25377) );
  AND2_X1 U25342 ( .A1(n25382), .A2(n25383), .ZN(n25380) );
  OR2_X1 U25343 ( .A1(n25384), .A2(n25385), .ZN(n25383) );
  INV_X1 U25344 ( .A(n25386), .ZN(n25385) );
  OR2_X1 U25345 ( .A1(n25386), .A2(n25387), .ZN(n25382) );
  INV_X1 U25346 ( .A(n25384), .ZN(n25387) );
  OR2_X1 U25347 ( .A1(n15106), .A2(n15490), .ZN(n25015) );
  OR2_X1 U25348 ( .A1(n25388), .A2(n25389), .ZN(n25012) );
  INV_X1 U25349 ( .A(n25390), .ZN(n25389) );
  OR2_X1 U25350 ( .A1(n25391), .A2(n25392), .ZN(n25390) );
  AND2_X1 U25351 ( .A1(n25392), .A2(n25391), .ZN(n25388) );
  AND2_X1 U25352 ( .A1(n25393), .A2(n25394), .ZN(n25391) );
  OR2_X1 U25353 ( .A1(n25395), .A2(n25396), .ZN(n25394) );
  INV_X1 U25354 ( .A(n25397), .ZN(n25396) );
  OR2_X1 U25355 ( .A1(n25397), .A2(n25398), .ZN(n25393) );
  INV_X1 U25356 ( .A(n25395), .ZN(n25398) );
  OR2_X1 U25357 ( .A1(n15140), .A2(n15490), .ZN(n25026) );
  OR2_X1 U25358 ( .A1(n25399), .A2(n25400), .ZN(n25023) );
  INV_X1 U25359 ( .A(n25401), .ZN(n25400) );
  OR2_X1 U25360 ( .A1(n25402), .A2(n25403), .ZN(n25401) );
  AND2_X1 U25361 ( .A1(n25403), .A2(n25402), .ZN(n25399) );
  AND2_X1 U25362 ( .A1(n25404), .A2(n25405), .ZN(n25402) );
  OR2_X1 U25363 ( .A1(n25406), .A2(n25407), .ZN(n25405) );
  INV_X1 U25364 ( .A(n25408), .ZN(n25407) );
  OR2_X1 U25365 ( .A1(n25408), .A2(n25409), .ZN(n25404) );
  INV_X1 U25366 ( .A(n25406), .ZN(n25409) );
  OR2_X1 U25367 ( .A1(n15174), .A2(n15490), .ZN(n25037) );
  OR2_X1 U25368 ( .A1(n25410), .A2(n25411), .ZN(n25034) );
  INV_X1 U25369 ( .A(n25412), .ZN(n25411) );
  OR2_X1 U25370 ( .A1(n25413), .A2(n25414), .ZN(n25412) );
  AND2_X1 U25371 ( .A1(n25414), .A2(n25413), .ZN(n25410) );
  AND2_X1 U25372 ( .A1(n25415), .A2(n25416), .ZN(n25413) );
  OR2_X1 U25373 ( .A1(n25417), .A2(n25418), .ZN(n25416) );
  INV_X1 U25374 ( .A(n25419), .ZN(n25418) );
  OR2_X1 U25375 ( .A1(n25419), .A2(n25420), .ZN(n25415) );
  INV_X1 U25376 ( .A(n25417), .ZN(n25420) );
  OR2_X1 U25377 ( .A1(n15208), .A2(n15490), .ZN(n25048) );
  OR2_X1 U25378 ( .A1(n25421), .A2(n25422), .ZN(n25045) );
  INV_X1 U25379 ( .A(n25423), .ZN(n25422) );
  OR2_X1 U25380 ( .A1(n25424), .A2(n25425), .ZN(n25423) );
  AND2_X1 U25381 ( .A1(n25425), .A2(n25424), .ZN(n25421) );
  AND2_X1 U25382 ( .A1(n25426), .A2(n25427), .ZN(n25424) );
  OR2_X1 U25383 ( .A1(n25428), .A2(n25429), .ZN(n25427) );
  INV_X1 U25384 ( .A(n25430), .ZN(n25429) );
  OR2_X1 U25385 ( .A1(n25430), .A2(n25431), .ZN(n25426) );
  INV_X1 U25386 ( .A(n25428), .ZN(n25431) );
  OR2_X1 U25387 ( .A1(n15242), .A2(n15490), .ZN(n25062) );
  OR2_X1 U25388 ( .A1(n25432), .A2(n25433), .ZN(n25056) );
  INV_X1 U25389 ( .A(n25434), .ZN(n25433) );
  OR2_X1 U25390 ( .A1(n25435), .A2(n25436), .ZN(n25434) );
  AND2_X1 U25391 ( .A1(n25436), .A2(n25435), .ZN(n25432) );
  AND2_X1 U25392 ( .A1(n25437), .A2(n25438), .ZN(n25435) );
  INV_X1 U25393 ( .A(n25439), .ZN(n25438) );
  AND2_X1 U25394 ( .A1(n25440), .A2(n25441), .ZN(n25439) );
  OR2_X1 U25395 ( .A1(n25441), .A2(n25440), .ZN(n25437) );
  INV_X1 U25396 ( .A(n25442), .ZN(n25440) );
  OR2_X1 U25397 ( .A1(n15287), .A2(n15490), .ZN(n25072) );
  AND2_X1 U25398 ( .A1(n25443), .A2(n25444), .ZN(n25067) );
  INV_X1 U25399 ( .A(n25445), .ZN(n25444) );
  AND2_X1 U25400 ( .A1(n25446), .A2(n25447), .ZN(n25445) );
  OR2_X1 U25401 ( .A1(n25447), .A2(n25446), .ZN(n25443) );
  OR2_X1 U25402 ( .A1(n25448), .A2(n25449), .ZN(n25446) );
  AND2_X1 U25403 ( .A1(n25450), .A2(n25451), .ZN(n25449) );
  INV_X1 U25404 ( .A(n25452), .ZN(n25450) );
  AND2_X1 U25405 ( .A1(n25453), .A2(n25452), .ZN(n25448) );
  INV_X1 U25406 ( .A(n25451), .ZN(n25453) );
  OR2_X1 U25407 ( .A1(n15321), .A2(n15490), .ZN(n25083) );
  AND2_X1 U25408 ( .A1(n25454), .A2(n25455), .ZN(n25078) );
  INV_X1 U25409 ( .A(n25456), .ZN(n25455) );
  AND2_X1 U25410 ( .A1(n25457), .A2(n25458), .ZN(n25456) );
  OR2_X1 U25411 ( .A1(n25458), .A2(n25457), .ZN(n25454) );
  OR2_X1 U25412 ( .A1(n25459), .A2(n25460), .ZN(n25457) );
  AND2_X1 U25413 ( .A1(n25461), .A2(n25462), .ZN(n25460) );
  INV_X1 U25414 ( .A(n25463), .ZN(n25461) );
  AND2_X1 U25415 ( .A1(n25464), .A2(n25463), .ZN(n25459) );
  INV_X1 U25416 ( .A(n25462), .ZN(n25464) );
  OR2_X1 U25417 ( .A1(n15355), .A2(n15490), .ZN(n25094) );
  AND2_X1 U25418 ( .A1(n25465), .A2(n25466), .ZN(n25089) );
  INV_X1 U25419 ( .A(n25467), .ZN(n25466) );
  AND2_X1 U25420 ( .A1(n25468), .A2(n25469), .ZN(n25467) );
  OR2_X1 U25421 ( .A1(n25469), .A2(n25468), .ZN(n25465) );
  OR2_X1 U25422 ( .A1(n25470), .A2(n25471), .ZN(n25468) );
  AND2_X1 U25423 ( .A1(n25472), .A2(n25473), .ZN(n25471) );
  INV_X1 U25424 ( .A(n25474), .ZN(n25472) );
  AND2_X1 U25425 ( .A1(n25475), .A2(n25474), .ZN(n25470) );
  INV_X1 U25426 ( .A(n25473), .ZN(n25475) );
  OR2_X1 U25427 ( .A1(n15389), .A2(n15490), .ZN(n25105) );
  AND2_X1 U25428 ( .A1(n25476), .A2(n25477), .ZN(n25100) );
  INV_X1 U25429 ( .A(n25478), .ZN(n25477) );
  AND2_X1 U25430 ( .A1(n25479), .A2(n25480), .ZN(n25478) );
  OR2_X1 U25431 ( .A1(n25480), .A2(n25479), .ZN(n25476) );
  OR2_X1 U25432 ( .A1(n25481), .A2(n25482), .ZN(n25479) );
  AND2_X1 U25433 ( .A1(n25483), .A2(n25484), .ZN(n25482) );
  INV_X1 U25434 ( .A(n25485), .ZN(n25483) );
  AND2_X1 U25435 ( .A1(n25486), .A2(n25485), .ZN(n25481) );
  INV_X1 U25436 ( .A(n25484), .ZN(n25486) );
  OR2_X1 U25437 ( .A1(n15423), .A2(n15490), .ZN(n25116) );
  AND2_X1 U25438 ( .A1(n25487), .A2(n25488), .ZN(n25111) );
  INV_X1 U25439 ( .A(n25489), .ZN(n25488) );
  AND2_X1 U25440 ( .A1(n25490), .A2(n25491), .ZN(n25489) );
  OR2_X1 U25441 ( .A1(n25491), .A2(n25490), .ZN(n25487) );
  OR2_X1 U25442 ( .A1(n25492), .A2(n25493), .ZN(n25490) );
  AND2_X1 U25443 ( .A1(n25494), .A2(n25495), .ZN(n25493) );
  INV_X1 U25444 ( .A(n25496), .ZN(n25494) );
  AND2_X1 U25445 ( .A1(n25497), .A2(n25496), .ZN(n25492) );
  INV_X1 U25446 ( .A(n25495), .ZN(n25497) );
  OR2_X1 U25447 ( .A1(n15457), .A2(n15490), .ZN(n25127) );
  AND2_X1 U25448 ( .A1(n25498), .A2(n25499), .ZN(n25122) );
  INV_X1 U25449 ( .A(n25500), .ZN(n25499) );
  AND2_X1 U25450 ( .A1(n25501), .A2(n25502), .ZN(n25500) );
  OR2_X1 U25451 ( .A1(n25502), .A2(n25501), .ZN(n25498) );
  OR2_X1 U25452 ( .A1(n25503), .A2(n25504), .ZN(n25501) );
  AND2_X1 U25453 ( .A1(n25505), .A2(n25506), .ZN(n25504) );
  INV_X1 U25454 ( .A(n25507), .ZN(n25505) );
  AND2_X1 U25455 ( .A1(n25508), .A2(n25507), .ZN(n25503) );
  INV_X1 U25456 ( .A(n25506), .ZN(n25508) );
  OR2_X1 U25457 ( .A1(n15491), .A2(n15490), .ZN(n15900) );
  AND2_X1 U25458 ( .A1(n25509), .A2(n25510), .ZN(n25133) );
  INV_X1 U25459 ( .A(n25511), .ZN(n25510) );
  AND2_X1 U25460 ( .A1(n25512), .A2(n25513), .ZN(n25511) );
  OR2_X1 U25461 ( .A1(n25513), .A2(n25512), .ZN(n25509) );
  OR2_X1 U25462 ( .A1(n25514), .A2(n25515), .ZN(n25512) );
  AND2_X1 U25463 ( .A1(n25516), .A2(n25517), .ZN(n25515) );
  INV_X1 U25464 ( .A(n25518), .ZN(n25516) );
  AND2_X1 U25465 ( .A1(n25519), .A2(n25518), .ZN(n25514) );
  INV_X1 U25466 ( .A(n25517), .ZN(n25519) );
  OR2_X1 U25467 ( .A1(n15525), .A2(n15490), .ZN(n25148) );
  AND2_X1 U25468 ( .A1(n25520), .A2(n25521), .ZN(n25143) );
  INV_X1 U25469 ( .A(n25522), .ZN(n25521) );
  AND2_X1 U25470 ( .A1(n25523), .A2(n25524), .ZN(n25522) );
  OR2_X1 U25471 ( .A1(n25524), .A2(n25523), .ZN(n25520) );
  OR2_X1 U25472 ( .A1(n25525), .A2(n25526), .ZN(n25523) );
  AND2_X1 U25473 ( .A1(n25527), .A2(n25528), .ZN(n25526) );
  INV_X1 U25474 ( .A(n25529), .ZN(n25527) );
  AND2_X1 U25475 ( .A1(n25530), .A2(n25529), .ZN(n25525) );
  INV_X1 U25476 ( .A(n25528), .ZN(n25530) );
  OR2_X1 U25477 ( .A1(n15559), .A2(n15490), .ZN(n25159) );
  AND2_X1 U25478 ( .A1(n25531), .A2(n25532), .ZN(n25154) );
  INV_X1 U25479 ( .A(n25533), .ZN(n25532) );
  AND2_X1 U25480 ( .A1(n25534), .A2(n25535), .ZN(n25533) );
  OR2_X1 U25481 ( .A1(n25535), .A2(n25534), .ZN(n25531) );
  OR2_X1 U25482 ( .A1(n25536), .A2(n25537), .ZN(n25534) );
  AND2_X1 U25483 ( .A1(n25538), .A2(n25539), .ZN(n25537) );
  INV_X1 U25484 ( .A(n15897), .ZN(n25538) );
  AND2_X1 U25485 ( .A1(n25540), .A2(n15897), .ZN(n25536) );
  INV_X1 U25486 ( .A(n25539), .ZN(n25540) );
  OR2_X1 U25487 ( .A1(n15593), .A2(n15490), .ZN(n25170) );
  AND2_X1 U25488 ( .A1(n25541), .A2(n25542), .ZN(n25165) );
  INV_X1 U25489 ( .A(n25543), .ZN(n25542) );
  AND2_X1 U25490 ( .A1(n25544), .A2(n25545), .ZN(n25543) );
  OR2_X1 U25491 ( .A1(n25545), .A2(n25544), .ZN(n25541) );
  OR2_X1 U25492 ( .A1(n25546), .A2(n25547), .ZN(n25544) );
  AND2_X1 U25493 ( .A1(n25548), .A2(n25549), .ZN(n25547) );
  INV_X1 U25494 ( .A(n25550), .ZN(n25548) );
  AND2_X1 U25495 ( .A1(n25551), .A2(n25550), .ZN(n25546) );
  INV_X1 U25496 ( .A(n25549), .ZN(n25551) );
  OR2_X1 U25497 ( .A1(n15638), .A2(n15490), .ZN(n25181) );
  AND2_X1 U25498 ( .A1(n25552), .A2(n25553), .ZN(n25176) );
  INV_X1 U25499 ( .A(n25554), .ZN(n25553) );
  AND2_X1 U25500 ( .A1(n25555), .A2(n25556), .ZN(n25554) );
  OR2_X1 U25501 ( .A1(n25556), .A2(n25555), .ZN(n25552) );
  OR2_X1 U25502 ( .A1(n25557), .A2(n25558), .ZN(n25555) );
  AND2_X1 U25503 ( .A1(n25559), .A2(n25560), .ZN(n25558) );
  INV_X1 U25504 ( .A(n25561), .ZN(n25559) );
  AND2_X1 U25505 ( .A1(n25562), .A2(n25561), .ZN(n25557) );
  INV_X1 U25506 ( .A(n25560), .ZN(n25562) );
  OR2_X1 U25507 ( .A1(n15672), .A2(n15490), .ZN(n25192) );
  AND2_X1 U25508 ( .A1(n25563), .A2(n25564), .ZN(n25187) );
  INV_X1 U25509 ( .A(n25565), .ZN(n25564) );
  AND2_X1 U25510 ( .A1(n25566), .A2(n25567), .ZN(n25565) );
  OR2_X1 U25511 ( .A1(n25567), .A2(n25566), .ZN(n25563) );
  OR2_X1 U25512 ( .A1(n25568), .A2(n25569), .ZN(n25566) );
  AND2_X1 U25513 ( .A1(n25570), .A2(n25571), .ZN(n25569) );
  INV_X1 U25514 ( .A(n25572), .ZN(n25570) );
  AND2_X1 U25515 ( .A1(n25573), .A2(n25572), .ZN(n25568) );
  INV_X1 U25516 ( .A(n25571), .ZN(n25573) );
  OR2_X1 U25517 ( .A1(n15706), .A2(n15490), .ZN(n25203) );
  AND2_X1 U25518 ( .A1(n25574), .A2(n25575), .ZN(n25198) );
  INV_X1 U25519 ( .A(n25576), .ZN(n25575) );
  AND2_X1 U25520 ( .A1(n25577), .A2(n25578), .ZN(n25576) );
  OR2_X1 U25521 ( .A1(n25578), .A2(n25577), .ZN(n25574) );
  OR2_X1 U25522 ( .A1(n25579), .A2(n25580), .ZN(n25577) );
  AND2_X1 U25523 ( .A1(n25581), .A2(n25582), .ZN(n25580) );
  INV_X1 U25524 ( .A(n25583), .ZN(n25581) );
  AND2_X1 U25525 ( .A1(n25584), .A2(n25583), .ZN(n25579) );
  INV_X1 U25526 ( .A(n25582), .ZN(n25584) );
  OR2_X1 U25527 ( .A1(n15740), .A2(n15490), .ZN(n25214) );
  AND2_X1 U25528 ( .A1(n25585), .A2(n25586), .ZN(n25209) );
  INV_X1 U25529 ( .A(n25587), .ZN(n25586) );
  AND2_X1 U25530 ( .A1(n25588), .A2(n25589), .ZN(n25587) );
  OR2_X1 U25531 ( .A1(n25589), .A2(n25588), .ZN(n25585) );
  OR2_X1 U25532 ( .A1(n25590), .A2(n25591), .ZN(n25588) );
  AND2_X1 U25533 ( .A1(n25592), .A2(n25593), .ZN(n25591) );
  INV_X1 U25534 ( .A(n25594), .ZN(n25592) );
  AND2_X1 U25535 ( .A1(n25595), .A2(n25594), .ZN(n25590) );
  INV_X1 U25536 ( .A(n25593), .ZN(n25595) );
  OR2_X1 U25537 ( .A1(n15774), .A2(n15490), .ZN(n25225) );
  INV_X1 U25538 ( .A(b_11_), .ZN(n15490) );
  AND2_X1 U25539 ( .A1(n25596), .A2(n25597), .ZN(n25220) );
  INV_X1 U25540 ( .A(n25598), .ZN(n25597) );
  AND2_X1 U25541 ( .A1(n25599), .A2(n25600), .ZN(n25598) );
  OR2_X1 U25542 ( .A1(n25600), .A2(n25599), .ZN(n25596) );
  OR2_X1 U25543 ( .A1(n25601), .A2(n25602), .ZN(n25599) );
  AND2_X1 U25544 ( .A1(n25603), .A2(n25604), .ZN(n25602) );
  INV_X1 U25545 ( .A(n25605), .ZN(n25603) );
  AND2_X1 U25546 ( .A1(n25606), .A2(n25605), .ZN(n25601) );
  INV_X1 U25547 ( .A(n25604), .ZN(n25606) );
  AND2_X1 U25548 ( .A1(n25607), .A2(n25608), .ZN(n16619) );
  INV_X1 U25549 ( .A(n25609), .ZN(n25608) );
  AND2_X1 U25550 ( .A1(n25610), .A2(n16633), .ZN(n25609) );
  OR2_X1 U25551 ( .A1(n16633), .A2(n25610), .ZN(n25607) );
  OR2_X1 U25552 ( .A1(n25611), .A2(n25612), .ZN(n25610) );
  AND2_X1 U25553 ( .A1(n25613), .A2(n16632), .ZN(n25612) );
  INV_X1 U25554 ( .A(n16631), .ZN(n25613) );
  AND2_X1 U25555 ( .A1(n25614), .A2(n16631), .ZN(n25611) );
  OR2_X1 U25556 ( .A1(n15774), .A2(n15524), .ZN(n16631) );
  INV_X1 U25557 ( .A(n16632), .ZN(n25614) );
  OR2_X1 U25558 ( .A1(n25615), .A2(n25616), .ZN(n16632) );
  AND2_X1 U25559 ( .A1(n25605), .A2(n25604), .ZN(n25616) );
  AND2_X1 U25560 ( .A1(n25600), .A2(n25617), .ZN(n25615) );
  OR2_X1 U25561 ( .A1(n25605), .A2(n25604), .ZN(n25617) );
  OR2_X1 U25562 ( .A1(n25618), .A2(n25619), .ZN(n25604) );
  AND2_X1 U25563 ( .A1(n25594), .A2(n25593), .ZN(n25619) );
  AND2_X1 U25564 ( .A1(n25589), .A2(n25620), .ZN(n25618) );
  OR2_X1 U25565 ( .A1(n25594), .A2(n25593), .ZN(n25620) );
  OR2_X1 U25566 ( .A1(n25621), .A2(n25622), .ZN(n25593) );
  AND2_X1 U25567 ( .A1(n25583), .A2(n25582), .ZN(n25622) );
  AND2_X1 U25568 ( .A1(n25578), .A2(n25623), .ZN(n25621) );
  OR2_X1 U25569 ( .A1(n25583), .A2(n25582), .ZN(n25623) );
  OR2_X1 U25570 ( .A1(n25624), .A2(n25625), .ZN(n25582) );
  AND2_X1 U25571 ( .A1(n25572), .A2(n25571), .ZN(n25625) );
  AND2_X1 U25572 ( .A1(n25567), .A2(n25626), .ZN(n25624) );
  OR2_X1 U25573 ( .A1(n25572), .A2(n25571), .ZN(n25626) );
  OR2_X1 U25574 ( .A1(n25627), .A2(n25628), .ZN(n25571) );
  AND2_X1 U25575 ( .A1(n25561), .A2(n25560), .ZN(n25628) );
  AND2_X1 U25576 ( .A1(n25556), .A2(n25629), .ZN(n25627) );
  OR2_X1 U25577 ( .A1(n25561), .A2(n25560), .ZN(n25629) );
  OR2_X1 U25578 ( .A1(n25630), .A2(n25631), .ZN(n25560) );
  AND2_X1 U25579 ( .A1(n25550), .A2(n25549), .ZN(n25631) );
  AND2_X1 U25580 ( .A1(n25545), .A2(n25632), .ZN(n25630) );
  OR2_X1 U25581 ( .A1(n25550), .A2(n25549), .ZN(n25632) );
  OR2_X1 U25582 ( .A1(n25633), .A2(n25634), .ZN(n25549) );
  AND2_X1 U25583 ( .A1(n15897), .A2(n25539), .ZN(n25634) );
  AND2_X1 U25584 ( .A1(n25535), .A2(n25635), .ZN(n25633) );
  OR2_X1 U25585 ( .A1(n15897), .A2(n25539), .ZN(n25635) );
  OR2_X1 U25586 ( .A1(n25636), .A2(n25637), .ZN(n25539) );
  AND2_X1 U25587 ( .A1(n25529), .A2(n25528), .ZN(n25637) );
  AND2_X1 U25588 ( .A1(n25524), .A2(n25638), .ZN(n25636) );
  OR2_X1 U25589 ( .A1(n25529), .A2(n25528), .ZN(n25638) );
  OR2_X1 U25590 ( .A1(n25639), .A2(n25640), .ZN(n25528) );
  AND2_X1 U25591 ( .A1(n25518), .A2(n25517), .ZN(n25640) );
  AND2_X1 U25592 ( .A1(n25513), .A2(n25641), .ZN(n25639) );
  OR2_X1 U25593 ( .A1(n25518), .A2(n25517), .ZN(n25641) );
  OR2_X1 U25594 ( .A1(n25642), .A2(n25643), .ZN(n25517) );
  AND2_X1 U25595 ( .A1(n25507), .A2(n25506), .ZN(n25643) );
  AND2_X1 U25596 ( .A1(n25502), .A2(n25644), .ZN(n25642) );
  OR2_X1 U25597 ( .A1(n25507), .A2(n25506), .ZN(n25644) );
  OR2_X1 U25598 ( .A1(n25645), .A2(n25646), .ZN(n25506) );
  AND2_X1 U25599 ( .A1(n25496), .A2(n25495), .ZN(n25646) );
  AND2_X1 U25600 ( .A1(n25491), .A2(n25647), .ZN(n25645) );
  OR2_X1 U25601 ( .A1(n25496), .A2(n25495), .ZN(n25647) );
  OR2_X1 U25602 ( .A1(n25648), .A2(n25649), .ZN(n25495) );
  AND2_X1 U25603 ( .A1(n25485), .A2(n25484), .ZN(n25649) );
  AND2_X1 U25604 ( .A1(n25480), .A2(n25650), .ZN(n25648) );
  OR2_X1 U25605 ( .A1(n25485), .A2(n25484), .ZN(n25650) );
  OR2_X1 U25606 ( .A1(n25651), .A2(n25652), .ZN(n25484) );
  AND2_X1 U25607 ( .A1(n25474), .A2(n25473), .ZN(n25652) );
  AND2_X1 U25608 ( .A1(n25469), .A2(n25653), .ZN(n25651) );
  OR2_X1 U25609 ( .A1(n25474), .A2(n25473), .ZN(n25653) );
  OR2_X1 U25610 ( .A1(n25654), .A2(n25655), .ZN(n25473) );
  AND2_X1 U25611 ( .A1(n25463), .A2(n25462), .ZN(n25655) );
  AND2_X1 U25612 ( .A1(n25458), .A2(n25656), .ZN(n25654) );
  OR2_X1 U25613 ( .A1(n25463), .A2(n25462), .ZN(n25656) );
  OR2_X1 U25614 ( .A1(n25657), .A2(n25658), .ZN(n25462) );
  AND2_X1 U25615 ( .A1(n25452), .A2(n25451), .ZN(n25658) );
  AND2_X1 U25616 ( .A1(n25447), .A2(n25659), .ZN(n25657) );
  OR2_X1 U25617 ( .A1(n25452), .A2(n25451), .ZN(n25659) );
  OR2_X1 U25618 ( .A1(n25660), .A2(n25661), .ZN(n25451) );
  AND2_X1 U25619 ( .A1(n25436), .A2(n25442), .ZN(n25661) );
  AND2_X1 U25620 ( .A1(n25662), .A2(n25441), .ZN(n25660) );
  OR2_X1 U25621 ( .A1(n25663), .A2(n25664), .ZN(n25441) );
  AND2_X1 U25622 ( .A1(n25428), .A2(n25430), .ZN(n25664) );
  AND2_X1 U25623 ( .A1(n25425), .A2(n25665), .ZN(n25663) );
  OR2_X1 U25624 ( .A1(n25428), .A2(n25430), .ZN(n25665) );
  OR2_X1 U25625 ( .A1(n25666), .A2(n25667), .ZN(n25430) );
  AND2_X1 U25626 ( .A1(n25414), .A2(n25417), .ZN(n25667) );
  AND2_X1 U25627 ( .A1(n25668), .A2(n25419), .ZN(n25666) );
  OR2_X1 U25628 ( .A1(n25669), .A2(n25670), .ZN(n25419) );
  AND2_X1 U25629 ( .A1(n25403), .A2(n25406), .ZN(n25670) );
  AND2_X1 U25630 ( .A1(n25671), .A2(n25408), .ZN(n25669) );
  OR2_X1 U25631 ( .A1(n25672), .A2(n25673), .ZN(n25408) );
  AND2_X1 U25632 ( .A1(n25392), .A2(n25395), .ZN(n25673) );
  AND2_X1 U25633 ( .A1(n25674), .A2(n25397), .ZN(n25672) );
  OR2_X1 U25634 ( .A1(n25675), .A2(n25676), .ZN(n25397) );
  AND2_X1 U25635 ( .A1(n25381), .A2(n25384), .ZN(n25676) );
  AND2_X1 U25636 ( .A1(n25677), .A2(n25386), .ZN(n25675) );
  OR2_X1 U25637 ( .A1(n25678), .A2(n25679), .ZN(n25386) );
  AND2_X1 U25638 ( .A1(n25370), .A2(n25373), .ZN(n25679) );
  AND2_X1 U25639 ( .A1(n25680), .A2(n25375), .ZN(n25678) );
  OR2_X1 U25640 ( .A1(n25681), .A2(n25682), .ZN(n25375) );
  AND2_X1 U25641 ( .A1(n25359), .A2(n25362), .ZN(n25682) );
  AND2_X1 U25642 ( .A1(n25683), .A2(n25364), .ZN(n25681) );
  OR2_X1 U25643 ( .A1(n25684), .A2(n25685), .ZN(n25364) );
  AND2_X1 U25644 ( .A1(n25348), .A2(n25351), .ZN(n25685) );
  AND2_X1 U25645 ( .A1(n25686), .A2(n25353), .ZN(n25684) );
  OR2_X1 U25646 ( .A1(n25687), .A2(n25688), .ZN(n25353) );
  AND2_X1 U25647 ( .A1(n25337), .A2(n25340), .ZN(n25688) );
  AND2_X1 U25648 ( .A1(n25689), .A2(n25342), .ZN(n25687) );
  OR2_X1 U25649 ( .A1(n25690), .A2(n25691), .ZN(n25342) );
  AND2_X1 U25650 ( .A1(n25325), .A2(n25330), .ZN(n25691) );
  AND2_X1 U25651 ( .A1(n25329), .A2(n25692), .ZN(n25690) );
  OR2_X1 U25652 ( .A1(n25325), .A2(n25330), .ZN(n25692) );
  INV_X1 U25653 ( .A(n25331), .ZN(n25330) );
  AND3_X1 U25654 ( .A1(b_10_), .A2(b_9_), .A3(n15957), .ZN(n25331) );
  OR2_X1 U25655 ( .A1(n14857), .A2(n15524), .ZN(n25325) );
  INV_X1 U25656 ( .A(n25332), .ZN(n25329) );
  OR2_X1 U25657 ( .A1(n25693), .A2(n25694), .ZN(n25332) );
  AND2_X1 U25658 ( .A1(b_9_), .A2(n25695), .ZN(n25694) );
  OR2_X1 U25659 ( .A1(n25696), .A2(n16981), .ZN(n25695) );
  AND2_X1 U25660 ( .A1(a_30_), .A2(n15592), .ZN(n25696) );
  AND2_X1 U25661 ( .A1(b_8_), .A2(n25697), .ZN(n25693) );
  OR2_X1 U25662 ( .A1(n25698), .A2(n14817), .ZN(n25697) );
  AND2_X1 U25663 ( .A1(a_31_), .A2(n15558), .ZN(n25698) );
  OR2_X1 U25664 ( .A1(n25337), .A2(n25340), .ZN(n25689) );
  OR2_X1 U25665 ( .A1(n14891), .A2(n15524), .ZN(n25340) );
  OR2_X1 U25666 ( .A1(n25699), .A2(n25700), .ZN(n25337) );
  AND2_X1 U25667 ( .A1(n25701), .A2(n25702), .ZN(n25700) );
  INV_X1 U25668 ( .A(n25703), .ZN(n25699) );
  OR2_X1 U25669 ( .A1(n25701), .A2(n25702), .ZN(n25703) );
  OR2_X1 U25670 ( .A1(n25704), .A2(n25705), .ZN(n25701) );
  AND2_X1 U25671 ( .A1(n25706), .A2(n25707), .ZN(n25705) );
  AND2_X1 U25672 ( .A1(n25708), .A2(n25709), .ZN(n25704) );
  OR2_X1 U25673 ( .A1(n25348), .A2(n25351), .ZN(n25686) );
  OR2_X1 U25674 ( .A1(n14936), .A2(n15524), .ZN(n25351) );
  OR2_X1 U25675 ( .A1(n25710), .A2(n25711), .ZN(n25348) );
  INV_X1 U25676 ( .A(n25712), .ZN(n25711) );
  OR2_X1 U25677 ( .A1(n25713), .A2(n25714), .ZN(n25712) );
  AND2_X1 U25678 ( .A1(n25714), .A2(n25713), .ZN(n25710) );
  AND2_X1 U25679 ( .A1(n25715), .A2(n25716), .ZN(n25713) );
  OR2_X1 U25680 ( .A1(n25717), .A2(n25718), .ZN(n25716) );
  INV_X1 U25681 ( .A(n25719), .ZN(n25718) );
  OR2_X1 U25682 ( .A1(n25719), .A2(n25720), .ZN(n25715) );
  INV_X1 U25683 ( .A(n25717), .ZN(n25720) );
  OR2_X1 U25684 ( .A1(n25359), .A2(n25362), .ZN(n25683) );
  OR2_X1 U25685 ( .A1(n14970), .A2(n15524), .ZN(n25362) );
  OR2_X1 U25686 ( .A1(n25721), .A2(n25722), .ZN(n25359) );
  INV_X1 U25687 ( .A(n25723), .ZN(n25722) );
  OR2_X1 U25688 ( .A1(n25724), .A2(n25725), .ZN(n25723) );
  AND2_X1 U25689 ( .A1(n25725), .A2(n25724), .ZN(n25721) );
  AND2_X1 U25690 ( .A1(n25726), .A2(n25727), .ZN(n25724) );
  OR2_X1 U25691 ( .A1(n25728), .A2(n25729), .ZN(n25727) );
  INV_X1 U25692 ( .A(n25730), .ZN(n25729) );
  OR2_X1 U25693 ( .A1(n25730), .A2(n25731), .ZN(n25726) );
  INV_X1 U25694 ( .A(n25728), .ZN(n25731) );
  OR2_X1 U25695 ( .A1(n25370), .A2(n25373), .ZN(n25680) );
  OR2_X1 U25696 ( .A1(n15004), .A2(n15524), .ZN(n25373) );
  OR2_X1 U25697 ( .A1(n25732), .A2(n25733), .ZN(n25370) );
  INV_X1 U25698 ( .A(n25734), .ZN(n25733) );
  OR2_X1 U25699 ( .A1(n25735), .A2(n25736), .ZN(n25734) );
  AND2_X1 U25700 ( .A1(n25736), .A2(n25735), .ZN(n25732) );
  AND2_X1 U25701 ( .A1(n25737), .A2(n25738), .ZN(n25735) );
  OR2_X1 U25702 ( .A1(n25739), .A2(n25740), .ZN(n25738) );
  INV_X1 U25703 ( .A(n25741), .ZN(n25740) );
  OR2_X1 U25704 ( .A1(n25741), .A2(n25742), .ZN(n25737) );
  INV_X1 U25705 ( .A(n25739), .ZN(n25742) );
  OR2_X1 U25706 ( .A1(n25381), .A2(n25384), .ZN(n25677) );
  OR2_X1 U25707 ( .A1(n15038), .A2(n15524), .ZN(n25384) );
  OR2_X1 U25708 ( .A1(n25743), .A2(n25744), .ZN(n25381) );
  INV_X1 U25709 ( .A(n25745), .ZN(n25744) );
  OR2_X1 U25710 ( .A1(n25746), .A2(n25747), .ZN(n25745) );
  AND2_X1 U25711 ( .A1(n25747), .A2(n25746), .ZN(n25743) );
  AND2_X1 U25712 ( .A1(n25748), .A2(n25749), .ZN(n25746) );
  OR2_X1 U25713 ( .A1(n25750), .A2(n25751), .ZN(n25749) );
  INV_X1 U25714 ( .A(n25752), .ZN(n25751) );
  OR2_X1 U25715 ( .A1(n25752), .A2(n25753), .ZN(n25748) );
  INV_X1 U25716 ( .A(n25750), .ZN(n25753) );
  OR2_X1 U25717 ( .A1(n25392), .A2(n25395), .ZN(n25674) );
  OR2_X1 U25718 ( .A1(n15072), .A2(n15524), .ZN(n25395) );
  OR2_X1 U25719 ( .A1(n25754), .A2(n25755), .ZN(n25392) );
  INV_X1 U25720 ( .A(n25756), .ZN(n25755) );
  OR2_X1 U25721 ( .A1(n25757), .A2(n25758), .ZN(n25756) );
  AND2_X1 U25722 ( .A1(n25758), .A2(n25757), .ZN(n25754) );
  AND2_X1 U25723 ( .A1(n25759), .A2(n25760), .ZN(n25757) );
  OR2_X1 U25724 ( .A1(n25761), .A2(n25762), .ZN(n25760) );
  INV_X1 U25725 ( .A(n25763), .ZN(n25762) );
  OR2_X1 U25726 ( .A1(n25763), .A2(n25764), .ZN(n25759) );
  INV_X1 U25727 ( .A(n25761), .ZN(n25764) );
  OR2_X1 U25728 ( .A1(n25403), .A2(n25406), .ZN(n25671) );
  OR2_X1 U25729 ( .A1(n15106), .A2(n15524), .ZN(n25406) );
  OR2_X1 U25730 ( .A1(n25765), .A2(n25766), .ZN(n25403) );
  INV_X1 U25731 ( .A(n25767), .ZN(n25766) );
  OR2_X1 U25732 ( .A1(n25768), .A2(n25769), .ZN(n25767) );
  AND2_X1 U25733 ( .A1(n25769), .A2(n25768), .ZN(n25765) );
  AND2_X1 U25734 ( .A1(n25770), .A2(n25771), .ZN(n25768) );
  OR2_X1 U25735 ( .A1(n25772), .A2(n25773), .ZN(n25771) );
  INV_X1 U25736 ( .A(n25774), .ZN(n25773) );
  OR2_X1 U25737 ( .A1(n25774), .A2(n25775), .ZN(n25770) );
  INV_X1 U25738 ( .A(n25772), .ZN(n25775) );
  OR2_X1 U25739 ( .A1(n25414), .A2(n25417), .ZN(n25668) );
  OR2_X1 U25740 ( .A1(n15140), .A2(n15524), .ZN(n25417) );
  OR2_X1 U25741 ( .A1(n25776), .A2(n25777), .ZN(n25414) );
  INV_X1 U25742 ( .A(n25778), .ZN(n25777) );
  OR2_X1 U25743 ( .A1(n25779), .A2(n25780), .ZN(n25778) );
  AND2_X1 U25744 ( .A1(n25780), .A2(n25779), .ZN(n25776) );
  AND2_X1 U25745 ( .A1(n25781), .A2(n25782), .ZN(n25779) );
  OR2_X1 U25746 ( .A1(n25783), .A2(n25784), .ZN(n25782) );
  INV_X1 U25747 ( .A(n25785), .ZN(n25784) );
  OR2_X1 U25748 ( .A1(n25785), .A2(n25786), .ZN(n25781) );
  INV_X1 U25749 ( .A(n25783), .ZN(n25786) );
  OR2_X1 U25750 ( .A1(n15174), .A2(n15524), .ZN(n25428) );
  OR2_X1 U25751 ( .A1(n25787), .A2(n25788), .ZN(n25425) );
  INV_X1 U25752 ( .A(n25789), .ZN(n25788) );
  OR2_X1 U25753 ( .A1(n25790), .A2(n25791), .ZN(n25789) );
  AND2_X1 U25754 ( .A1(n25791), .A2(n25790), .ZN(n25787) );
  AND2_X1 U25755 ( .A1(n25792), .A2(n25793), .ZN(n25790) );
  OR2_X1 U25756 ( .A1(n25794), .A2(n25795), .ZN(n25793) );
  INV_X1 U25757 ( .A(n25796), .ZN(n25795) );
  OR2_X1 U25758 ( .A1(n25796), .A2(n25797), .ZN(n25792) );
  INV_X1 U25759 ( .A(n25794), .ZN(n25797) );
  OR2_X1 U25760 ( .A1(n25436), .A2(n25442), .ZN(n25662) );
  OR2_X1 U25761 ( .A1(n15208), .A2(n15524), .ZN(n25442) );
  OR2_X1 U25762 ( .A1(n25798), .A2(n25799), .ZN(n25436) );
  INV_X1 U25763 ( .A(n25800), .ZN(n25799) );
  OR2_X1 U25764 ( .A1(n25801), .A2(n25802), .ZN(n25800) );
  AND2_X1 U25765 ( .A1(n25802), .A2(n25801), .ZN(n25798) );
  AND2_X1 U25766 ( .A1(n25803), .A2(n25804), .ZN(n25801) );
  INV_X1 U25767 ( .A(n25805), .ZN(n25804) );
  AND2_X1 U25768 ( .A1(n25806), .A2(n25807), .ZN(n25805) );
  OR2_X1 U25769 ( .A1(n25807), .A2(n25806), .ZN(n25803) );
  INV_X1 U25770 ( .A(n25808), .ZN(n25806) );
  OR2_X1 U25771 ( .A1(n15242), .A2(n15524), .ZN(n25452) );
  AND2_X1 U25772 ( .A1(n25809), .A2(n25810), .ZN(n25447) );
  INV_X1 U25773 ( .A(n25811), .ZN(n25810) );
  AND2_X1 U25774 ( .A1(n25812), .A2(n25813), .ZN(n25811) );
  OR2_X1 U25775 ( .A1(n25813), .A2(n25812), .ZN(n25809) );
  OR2_X1 U25776 ( .A1(n25814), .A2(n25815), .ZN(n25812) );
  AND2_X1 U25777 ( .A1(n25816), .A2(n25817), .ZN(n25815) );
  INV_X1 U25778 ( .A(n25818), .ZN(n25816) );
  AND2_X1 U25779 ( .A1(n25819), .A2(n25818), .ZN(n25814) );
  INV_X1 U25780 ( .A(n25817), .ZN(n25819) );
  OR2_X1 U25781 ( .A1(n15287), .A2(n15524), .ZN(n25463) );
  AND2_X1 U25782 ( .A1(n25820), .A2(n25821), .ZN(n25458) );
  INV_X1 U25783 ( .A(n25822), .ZN(n25821) );
  AND2_X1 U25784 ( .A1(n25823), .A2(n25824), .ZN(n25822) );
  OR2_X1 U25785 ( .A1(n25824), .A2(n25823), .ZN(n25820) );
  OR2_X1 U25786 ( .A1(n25825), .A2(n25826), .ZN(n25823) );
  AND2_X1 U25787 ( .A1(n25827), .A2(n25828), .ZN(n25826) );
  INV_X1 U25788 ( .A(n25829), .ZN(n25827) );
  AND2_X1 U25789 ( .A1(n25830), .A2(n25829), .ZN(n25825) );
  INV_X1 U25790 ( .A(n25828), .ZN(n25830) );
  OR2_X1 U25791 ( .A1(n15321), .A2(n15524), .ZN(n25474) );
  AND2_X1 U25792 ( .A1(n25831), .A2(n25832), .ZN(n25469) );
  INV_X1 U25793 ( .A(n25833), .ZN(n25832) );
  AND2_X1 U25794 ( .A1(n25834), .A2(n25835), .ZN(n25833) );
  OR2_X1 U25795 ( .A1(n25835), .A2(n25834), .ZN(n25831) );
  OR2_X1 U25796 ( .A1(n25836), .A2(n25837), .ZN(n25834) );
  AND2_X1 U25797 ( .A1(n25838), .A2(n25839), .ZN(n25837) );
  INV_X1 U25798 ( .A(n25840), .ZN(n25838) );
  AND2_X1 U25799 ( .A1(n25841), .A2(n25840), .ZN(n25836) );
  INV_X1 U25800 ( .A(n25839), .ZN(n25841) );
  OR2_X1 U25801 ( .A1(n15355), .A2(n15524), .ZN(n25485) );
  AND2_X1 U25802 ( .A1(n25842), .A2(n25843), .ZN(n25480) );
  INV_X1 U25803 ( .A(n25844), .ZN(n25843) );
  AND2_X1 U25804 ( .A1(n25845), .A2(n25846), .ZN(n25844) );
  OR2_X1 U25805 ( .A1(n25846), .A2(n25845), .ZN(n25842) );
  OR2_X1 U25806 ( .A1(n25847), .A2(n25848), .ZN(n25845) );
  AND2_X1 U25807 ( .A1(n25849), .A2(n25850), .ZN(n25848) );
  INV_X1 U25808 ( .A(n25851), .ZN(n25849) );
  AND2_X1 U25809 ( .A1(n25852), .A2(n25851), .ZN(n25847) );
  INV_X1 U25810 ( .A(n25850), .ZN(n25852) );
  OR2_X1 U25811 ( .A1(n15389), .A2(n15524), .ZN(n25496) );
  AND2_X1 U25812 ( .A1(n25853), .A2(n25854), .ZN(n25491) );
  INV_X1 U25813 ( .A(n25855), .ZN(n25854) );
  AND2_X1 U25814 ( .A1(n25856), .A2(n25857), .ZN(n25855) );
  OR2_X1 U25815 ( .A1(n25857), .A2(n25856), .ZN(n25853) );
  OR2_X1 U25816 ( .A1(n25858), .A2(n25859), .ZN(n25856) );
  AND2_X1 U25817 ( .A1(n25860), .A2(n25861), .ZN(n25859) );
  INV_X1 U25818 ( .A(n25862), .ZN(n25860) );
  AND2_X1 U25819 ( .A1(n25863), .A2(n25862), .ZN(n25858) );
  INV_X1 U25820 ( .A(n25861), .ZN(n25863) );
  OR2_X1 U25821 ( .A1(n15423), .A2(n15524), .ZN(n25507) );
  AND2_X1 U25822 ( .A1(n25864), .A2(n25865), .ZN(n25502) );
  INV_X1 U25823 ( .A(n25866), .ZN(n25865) );
  AND2_X1 U25824 ( .A1(n25867), .A2(n25868), .ZN(n25866) );
  OR2_X1 U25825 ( .A1(n25868), .A2(n25867), .ZN(n25864) );
  OR2_X1 U25826 ( .A1(n25869), .A2(n25870), .ZN(n25867) );
  AND2_X1 U25827 ( .A1(n25871), .A2(n25872), .ZN(n25870) );
  INV_X1 U25828 ( .A(n25873), .ZN(n25871) );
  AND2_X1 U25829 ( .A1(n25874), .A2(n25873), .ZN(n25869) );
  INV_X1 U25830 ( .A(n25872), .ZN(n25874) );
  OR2_X1 U25831 ( .A1(n15457), .A2(n15524), .ZN(n25518) );
  AND2_X1 U25832 ( .A1(n25875), .A2(n25876), .ZN(n25513) );
  INV_X1 U25833 ( .A(n25877), .ZN(n25876) );
  AND2_X1 U25834 ( .A1(n25878), .A2(n25879), .ZN(n25877) );
  OR2_X1 U25835 ( .A1(n25879), .A2(n25878), .ZN(n25875) );
  OR2_X1 U25836 ( .A1(n25880), .A2(n25881), .ZN(n25878) );
  AND2_X1 U25837 ( .A1(n25882), .A2(n25883), .ZN(n25881) );
  INV_X1 U25838 ( .A(n25884), .ZN(n25882) );
  AND2_X1 U25839 ( .A1(n25885), .A2(n25884), .ZN(n25880) );
  INV_X1 U25840 ( .A(n25883), .ZN(n25885) );
  OR2_X1 U25841 ( .A1(n15491), .A2(n15524), .ZN(n25529) );
  AND2_X1 U25842 ( .A1(n25886), .A2(n25887), .ZN(n25524) );
  INV_X1 U25843 ( .A(n25888), .ZN(n25887) );
  AND2_X1 U25844 ( .A1(n25889), .A2(n25890), .ZN(n25888) );
  OR2_X1 U25845 ( .A1(n25890), .A2(n25889), .ZN(n25886) );
  OR2_X1 U25846 ( .A1(n25891), .A2(n25892), .ZN(n25889) );
  AND2_X1 U25847 ( .A1(n25893), .A2(n25894), .ZN(n25892) );
  INV_X1 U25848 ( .A(n25895), .ZN(n25893) );
  AND2_X1 U25849 ( .A1(n25896), .A2(n25895), .ZN(n25891) );
  INV_X1 U25850 ( .A(n25894), .ZN(n25896) );
  OR2_X1 U25851 ( .A1(n15525), .A2(n15524), .ZN(n15897) );
  AND2_X1 U25852 ( .A1(n25897), .A2(n25898), .ZN(n25535) );
  INV_X1 U25853 ( .A(n25899), .ZN(n25898) );
  AND2_X1 U25854 ( .A1(n25900), .A2(n25901), .ZN(n25899) );
  OR2_X1 U25855 ( .A1(n25901), .A2(n25900), .ZN(n25897) );
  OR2_X1 U25856 ( .A1(n25902), .A2(n25903), .ZN(n25900) );
  AND2_X1 U25857 ( .A1(n25904), .A2(n25905), .ZN(n25903) );
  INV_X1 U25858 ( .A(n25906), .ZN(n25904) );
  AND2_X1 U25859 ( .A1(n25907), .A2(n25906), .ZN(n25902) );
  INV_X1 U25860 ( .A(n25905), .ZN(n25907) );
  OR2_X1 U25861 ( .A1(n15559), .A2(n15524), .ZN(n25550) );
  AND2_X1 U25862 ( .A1(n25908), .A2(n25909), .ZN(n25545) );
  INV_X1 U25863 ( .A(n25910), .ZN(n25909) );
  AND2_X1 U25864 ( .A1(n25911), .A2(n25912), .ZN(n25910) );
  OR2_X1 U25865 ( .A1(n25912), .A2(n25911), .ZN(n25908) );
  OR2_X1 U25866 ( .A1(n25913), .A2(n25914), .ZN(n25911) );
  AND2_X1 U25867 ( .A1(n25915), .A2(n25916), .ZN(n25914) );
  INV_X1 U25868 ( .A(n25917), .ZN(n25915) );
  AND2_X1 U25869 ( .A1(n25918), .A2(n25917), .ZN(n25913) );
  INV_X1 U25870 ( .A(n25916), .ZN(n25918) );
  OR2_X1 U25871 ( .A1(n15593), .A2(n15524), .ZN(n25561) );
  AND2_X1 U25872 ( .A1(n25919), .A2(n25920), .ZN(n25556) );
  INV_X1 U25873 ( .A(n25921), .ZN(n25920) );
  AND2_X1 U25874 ( .A1(n25922), .A2(n25923), .ZN(n25921) );
  OR2_X1 U25875 ( .A1(n25923), .A2(n25922), .ZN(n25919) );
  OR2_X1 U25876 ( .A1(n25924), .A2(n25925), .ZN(n25922) );
  AND2_X1 U25877 ( .A1(n25926), .A2(n25927), .ZN(n25925) );
  INV_X1 U25878 ( .A(n15894), .ZN(n25926) );
  AND2_X1 U25879 ( .A1(n25928), .A2(n15894), .ZN(n25924) );
  INV_X1 U25880 ( .A(n25927), .ZN(n25928) );
  OR2_X1 U25881 ( .A1(n15638), .A2(n15524), .ZN(n25572) );
  AND2_X1 U25882 ( .A1(n25929), .A2(n25930), .ZN(n25567) );
  INV_X1 U25883 ( .A(n25931), .ZN(n25930) );
  AND2_X1 U25884 ( .A1(n25932), .A2(n25933), .ZN(n25931) );
  OR2_X1 U25885 ( .A1(n25933), .A2(n25932), .ZN(n25929) );
  OR2_X1 U25886 ( .A1(n25934), .A2(n25935), .ZN(n25932) );
  AND2_X1 U25887 ( .A1(n25936), .A2(n25937), .ZN(n25935) );
  INV_X1 U25888 ( .A(n25938), .ZN(n25936) );
  AND2_X1 U25889 ( .A1(n25939), .A2(n25938), .ZN(n25934) );
  INV_X1 U25890 ( .A(n25937), .ZN(n25939) );
  OR2_X1 U25891 ( .A1(n15672), .A2(n15524), .ZN(n25583) );
  AND2_X1 U25892 ( .A1(n25940), .A2(n25941), .ZN(n25578) );
  INV_X1 U25893 ( .A(n25942), .ZN(n25941) );
  AND2_X1 U25894 ( .A1(n25943), .A2(n25944), .ZN(n25942) );
  OR2_X1 U25895 ( .A1(n25944), .A2(n25943), .ZN(n25940) );
  OR2_X1 U25896 ( .A1(n25945), .A2(n25946), .ZN(n25943) );
  AND2_X1 U25897 ( .A1(n25947), .A2(n25948), .ZN(n25946) );
  INV_X1 U25898 ( .A(n25949), .ZN(n25947) );
  AND2_X1 U25899 ( .A1(n25950), .A2(n25949), .ZN(n25945) );
  INV_X1 U25900 ( .A(n25948), .ZN(n25950) );
  OR2_X1 U25901 ( .A1(n15706), .A2(n15524), .ZN(n25594) );
  AND2_X1 U25902 ( .A1(n25951), .A2(n25952), .ZN(n25589) );
  INV_X1 U25903 ( .A(n25953), .ZN(n25952) );
  AND2_X1 U25904 ( .A1(n25954), .A2(n25955), .ZN(n25953) );
  OR2_X1 U25905 ( .A1(n25955), .A2(n25954), .ZN(n25951) );
  OR2_X1 U25906 ( .A1(n25956), .A2(n25957), .ZN(n25954) );
  AND2_X1 U25907 ( .A1(n25958), .A2(n25959), .ZN(n25957) );
  INV_X1 U25908 ( .A(n25960), .ZN(n25958) );
  AND2_X1 U25909 ( .A1(n25961), .A2(n25960), .ZN(n25956) );
  INV_X1 U25910 ( .A(n25959), .ZN(n25961) );
  OR2_X1 U25911 ( .A1(n15740), .A2(n15524), .ZN(n25605) );
  INV_X1 U25912 ( .A(b_10_), .ZN(n15524) );
  AND2_X1 U25913 ( .A1(n25962), .A2(n25963), .ZN(n25600) );
  INV_X1 U25914 ( .A(n25964), .ZN(n25963) );
  AND2_X1 U25915 ( .A1(n25965), .A2(n25966), .ZN(n25964) );
  OR2_X1 U25916 ( .A1(n25966), .A2(n25965), .ZN(n25962) );
  OR2_X1 U25917 ( .A1(n25967), .A2(n25968), .ZN(n25965) );
  AND2_X1 U25918 ( .A1(n25969), .A2(n25970), .ZN(n25968) );
  INV_X1 U25919 ( .A(n25971), .ZN(n25969) );
  AND2_X1 U25920 ( .A1(n25972), .A2(n25971), .ZN(n25967) );
  INV_X1 U25921 ( .A(n25970), .ZN(n25972) );
  AND2_X1 U25922 ( .A1(n25973), .A2(n25974), .ZN(n16633) );
  INV_X1 U25923 ( .A(n25975), .ZN(n25974) );
  AND2_X1 U25924 ( .A1(n25976), .A2(n25977), .ZN(n25975) );
  OR2_X1 U25925 ( .A1(n25977), .A2(n25976), .ZN(n25973) );
  OR2_X1 U25926 ( .A1(n25978), .A2(n25979), .ZN(n25976) );
  AND2_X1 U25927 ( .A1(n25980), .A2(n25981), .ZN(n25979) );
  INV_X1 U25928 ( .A(n25982), .ZN(n25980) );
  AND2_X1 U25929 ( .A1(n25983), .A2(n25982), .ZN(n25978) );
  INV_X1 U25930 ( .A(n25981), .ZN(n25983) );
  OR2_X1 U25931 ( .A1(n16471), .A2(n16472), .ZN(n14761) );
  OR2_X1 U25932 ( .A1(n25984), .A2(n25985), .ZN(n16472) );
  AND2_X1 U25933 ( .A1(n16492), .A2(n16491), .ZN(n25985) );
  AND2_X1 U25934 ( .A1(n16487), .A2(n25986), .ZN(n25984) );
  OR2_X1 U25935 ( .A1(n16491), .A2(n16492), .ZN(n25986) );
  OR2_X1 U25936 ( .A1(n16512), .A2(n15558), .ZN(n16492) );
  OR2_X1 U25937 ( .A1(n25987), .A2(n25988), .ZN(n16491) );
  AND2_X1 U25938 ( .A1(n16528), .A2(n16527), .ZN(n25988) );
  AND2_X1 U25939 ( .A1(n16523), .A2(n25989), .ZN(n25987) );
  OR2_X1 U25940 ( .A1(n16527), .A2(n16528), .ZN(n25989) );
  OR2_X1 U25941 ( .A1(n15842), .A2(n15558), .ZN(n16528) );
  OR2_X1 U25942 ( .A1(n25990), .A2(n25991), .ZN(n16527) );
  AND2_X1 U25943 ( .A1(n16581), .A2(n16580), .ZN(n25991) );
  AND2_X1 U25944 ( .A1(n16576), .A2(n25992), .ZN(n25990) );
  OR2_X1 U25945 ( .A1(n16580), .A2(n16581), .ZN(n25992) );
  OR2_X1 U25946 ( .A1(n15808), .A2(n15558), .ZN(n16581) );
  OR2_X1 U25947 ( .A1(n25993), .A2(n25994), .ZN(n16580) );
  AND2_X1 U25948 ( .A1(n16644), .A2(n16643), .ZN(n25994) );
  AND2_X1 U25949 ( .A1(n16639), .A2(n25995), .ZN(n25993) );
  OR2_X1 U25950 ( .A1(n16643), .A2(n16644), .ZN(n25995) );
  OR2_X1 U25951 ( .A1(n15774), .A2(n15558), .ZN(n16644) );
  OR2_X1 U25952 ( .A1(n25996), .A2(n25997), .ZN(n16643) );
  AND2_X1 U25953 ( .A1(n25982), .A2(n25981), .ZN(n25997) );
  AND2_X1 U25954 ( .A1(n25977), .A2(n25998), .ZN(n25996) );
  OR2_X1 U25955 ( .A1(n25981), .A2(n25982), .ZN(n25998) );
  OR2_X1 U25956 ( .A1(n15740), .A2(n15558), .ZN(n25982) );
  OR2_X1 U25957 ( .A1(n25999), .A2(n26000), .ZN(n25981) );
  AND2_X1 U25958 ( .A1(n25971), .A2(n25970), .ZN(n26000) );
  AND2_X1 U25959 ( .A1(n25966), .A2(n26001), .ZN(n25999) );
  OR2_X1 U25960 ( .A1(n25970), .A2(n25971), .ZN(n26001) );
  OR2_X1 U25961 ( .A1(n15706), .A2(n15558), .ZN(n25971) );
  OR2_X1 U25962 ( .A1(n26002), .A2(n26003), .ZN(n25970) );
  AND2_X1 U25963 ( .A1(n25960), .A2(n25959), .ZN(n26003) );
  AND2_X1 U25964 ( .A1(n25955), .A2(n26004), .ZN(n26002) );
  OR2_X1 U25965 ( .A1(n25959), .A2(n25960), .ZN(n26004) );
  OR2_X1 U25966 ( .A1(n15672), .A2(n15558), .ZN(n25960) );
  OR2_X1 U25967 ( .A1(n26005), .A2(n26006), .ZN(n25959) );
  AND2_X1 U25968 ( .A1(n25949), .A2(n25948), .ZN(n26006) );
  AND2_X1 U25969 ( .A1(n25944), .A2(n26007), .ZN(n26005) );
  OR2_X1 U25970 ( .A1(n25948), .A2(n25949), .ZN(n26007) );
  OR2_X1 U25971 ( .A1(n15638), .A2(n15558), .ZN(n25949) );
  OR2_X1 U25972 ( .A1(n26008), .A2(n26009), .ZN(n25948) );
  AND2_X1 U25973 ( .A1(n25938), .A2(n25937), .ZN(n26009) );
  AND2_X1 U25974 ( .A1(n25933), .A2(n26010), .ZN(n26008) );
  OR2_X1 U25975 ( .A1(n25937), .A2(n25938), .ZN(n26010) );
  OR2_X1 U25976 ( .A1(n15593), .A2(n15558), .ZN(n25938) );
  OR2_X1 U25977 ( .A1(n26011), .A2(n26012), .ZN(n25937) );
  AND2_X1 U25978 ( .A1(n15894), .A2(n25927), .ZN(n26012) );
  AND2_X1 U25979 ( .A1(n25923), .A2(n26013), .ZN(n26011) );
  OR2_X1 U25980 ( .A1(n25927), .A2(n15894), .ZN(n26013) );
  OR2_X1 U25981 ( .A1(n15559), .A2(n15558), .ZN(n15894) );
  OR2_X1 U25982 ( .A1(n26014), .A2(n26015), .ZN(n25927) );
  AND2_X1 U25983 ( .A1(n25917), .A2(n25916), .ZN(n26015) );
  AND2_X1 U25984 ( .A1(n25912), .A2(n26016), .ZN(n26014) );
  OR2_X1 U25985 ( .A1(n25916), .A2(n25917), .ZN(n26016) );
  OR2_X1 U25986 ( .A1(n15525), .A2(n15558), .ZN(n25917) );
  OR2_X1 U25987 ( .A1(n26017), .A2(n26018), .ZN(n25916) );
  AND2_X1 U25988 ( .A1(n25906), .A2(n25905), .ZN(n26018) );
  AND2_X1 U25989 ( .A1(n25901), .A2(n26019), .ZN(n26017) );
  OR2_X1 U25990 ( .A1(n25905), .A2(n25906), .ZN(n26019) );
  OR2_X1 U25991 ( .A1(n15491), .A2(n15558), .ZN(n25906) );
  OR2_X1 U25992 ( .A1(n26020), .A2(n26021), .ZN(n25905) );
  AND2_X1 U25993 ( .A1(n25895), .A2(n25894), .ZN(n26021) );
  AND2_X1 U25994 ( .A1(n25890), .A2(n26022), .ZN(n26020) );
  OR2_X1 U25995 ( .A1(n25894), .A2(n25895), .ZN(n26022) );
  OR2_X1 U25996 ( .A1(n15457), .A2(n15558), .ZN(n25895) );
  OR2_X1 U25997 ( .A1(n26023), .A2(n26024), .ZN(n25894) );
  AND2_X1 U25998 ( .A1(n25884), .A2(n25883), .ZN(n26024) );
  AND2_X1 U25999 ( .A1(n25879), .A2(n26025), .ZN(n26023) );
  OR2_X1 U26000 ( .A1(n25883), .A2(n25884), .ZN(n26025) );
  OR2_X1 U26001 ( .A1(n15423), .A2(n15558), .ZN(n25884) );
  OR2_X1 U26002 ( .A1(n26026), .A2(n26027), .ZN(n25883) );
  AND2_X1 U26003 ( .A1(n25873), .A2(n25872), .ZN(n26027) );
  AND2_X1 U26004 ( .A1(n25868), .A2(n26028), .ZN(n26026) );
  OR2_X1 U26005 ( .A1(n25872), .A2(n25873), .ZN(n26028) );
  OR2_X1 U26006 ( .A1(n15389), .A2(n15558), .ZN(n25873) );
  OR2_X1 U26007 ( .A1(n26029), .A2(n26030), .ZN(n25872) );
  AND2_X1 U26008 ( .A1(n25862), .A2(n25861), .ZN(n26030) );
  AND2_X1 U26009 ( .A1(n25857), .A2(n26031), .ZN(n26029) );
  OR2_X1 U26010 ( .A1(n25861), .A2(n25862), .ZN(n26031) );
  OR2_X1 U26011 ( .A1(n15355), .A2(n15558), .ZN(n25862) );
  OR2_X1 U26012 ( .A1(n26032), .A2(n26033), .ZN(n25861) );
  AND2_X1 U26013 ( .A1(n25851), .A2(n25850), .ZN(n26033) );
  AND2_X1 U26014 ( .A1(n25846), .A2(n26034), .ZN(n26032) );
  OR2_X1 U26015 ( .A1(n25850), .A2(n25851), .ZN(n26034) );
  OR2_X1 U26016 ( .A1(n15321), .A2(n15558), .ZN(n25851) );
  OR2_X1 U26017 ( .A1(n26035), .A2(n26036), .ZN(n25850) );
  AND2_X1 U26018 ( .A1(n25840), .A2(n25839), .ZN(n26036) );
  AND2_X1 U26019 ( .A1(n25835), .A2(n26037), .ZN(n26035) );
  OR2_X1 U26020 ( .A1(n25839), .A2(n25840), .ZN(n26037) );
  OR2_X1 U26021 ( .A1(n15287), .A2(n15558), .ZN(n25840) );
  OR2_X1 U26022 ( .A1(n26038), .A2(n26039), .ZN(n25839) );
  AND2_X1 U26023 ( .A1(n25829), .A2(n25828), .ZN(n26039) );
  AND2_X1 U26024 ( .A1(n25824), .A2(n26040), .ZN(n26038) );
  OR2_X1 U26025 ( .A1(n25828), .A2(n25829), .ZN(n26040) );
  OR2_X1 U26026 ( .A1(n15242), .A2(n15558), .ZN(n25829) );
  OR2_X1 U26027 ( .A1(n26041), .A2(n26042), .ZN(n25828) );
  AND2_X1 U26028 ( .A1(n25818), .A2(n25817), .ZN(n26042) );
  AND2_X1 U26029 ( .A1(n25813), .A2(n26043), .ZN(n26041) );
  OR2_X1 U26030 ( .A1(n25817), .A2(n25818), .ZN(n26043) );
  OR2_X1 U26031 ( .A1(n15208), .A2(n15558), .ZN(n25818) );
  OR2_X1 U26032 ( .A1(n26044), .A2(n26045), .ZN(n25817) );
  AND2_X1 U26033 ( .A1(n25802), .A2(n25808), .ZN(n26045) );
  AND2_X1 U26034 ( .A1(n26046), .A2(n25807), .ZN(n26044) );
  OR2_X1 U26035 ( .A1(n26047), .A2(n26048), .ZN(n25807) );
  AND2_X1 U26036 ( .A1(n25794), .A2(n25796), .ZN(n26048) );
  AND2_X1 U26037 ( .A1(n25791), .A2(n26049), .ZN(n26047) );
  OR2_X1 U26038 ( .A1(n25796), .A2(n25794), .ZN(n26049) );
  OR2_X1 U26039 ( .A1(n15140), .A2(n15558), .ZN(n25794) );
  OR2_X1 U26040 ( .A1(n26050), .A2(n26051), .ZN(n25796) );
  AND2_X1 U26041 ( .A1(n25780), .A2(n25783), .ZN(n26051) );
  AND2_X1 U26042 ( .A1(n26052), .A2(n25785), .ZN(n26050) );
  OR2_X1 U26043 ( .A1(n26053), .A2(n26054), .ZN(n25785) );
  AND2_X1 U26044 ( .A1(n25769), .A2(n25772), .ZN(n26054) );
  AND2_X1 U26045 ( .A1(n26055), .A2(n25774), .ZN(n26053) );
  OR2_X1 U26046 ( .A1(n26056), .A2(n26057), .ZN(n25774) );
  AND2_X1 U26047 ( .A1(n25758), .A2(n25761), .ZN(n26057) );
  AND2_X1 U26048 ( .A1(n26058), .A2(n25763), .ZN(n26056) );
  OR2_X1 U26049 ( .A1(n26059), .A2(n26060), .ZN(n25763) );
  AND2_X1 U26050 ( .A1(n25747), .A2(n25750), .ZN(n26060) );
  AND2_X1 U26051 ( .A1(n26061), .A2(n25752), .ZN(n26059) );
  OR2_X1 U26052 ( .A1(n26062), .A2(n26063), .ZN(n25752) );
  AND2_X1 U26053 ( .A1(n25736), .A2(n25739), .ZN(n26063) );
  AND2_X1 U26054 ( .A1(n26064), .A2(n25741), .ZN(n26062) );
  OR2_X1 U26055 ( .A1(n26065), .A2(n26066), .ZN(n25741) );
  AND2_X1 U26056 ( .A1(n25725), .A2(n25728), .ZN(n26066) );
  AND2_X1 U26057 ( .A1(n26067), .A2(n25730), .ZN(n26065) );
  OR2_X1 U26058 ( .A1(n26068), .A2(n26069), .ZN(n25730) );
  AND2_X1 U26059 ( .A1(n25714), .A2(n25717), .ZN(n26069) );
  AND2_X1 U26060 ( .A1(n26070), .A2(n25719), .ZN(n26068) );
  OR2_X1 U26061 ( .A1(n26071), .A2(n26072), .ZN(n25719) );
  AND2_X1 U26062 ( .A1(n25702), .A2(n25707), .ZN(n26072) );
  AND2_X1 U26063 ( .A1(n25706), .A2(n26073), .ZN(n26071) );
  OR2_X1 U26064 ( .A1(n25707), .A2(n25702), .ZN(n26073) );
  OR2_X1 U26065 ( .A1(n14857), .A2(n15558), .ZN(n25702) );
  INV_X1 U26066 ( .A(n25708), .ZN(n25707) );
  AND3_X1 U26067 ( .A1(b_9_), .A2(b_8_), .A3(n15957), .ZN(n25708) );
  INV_X1 U26068 ( .A(n25709), .ZN(n25706) );
  OR2_X1 U26069 ( .A1(n26074), .A2(n26075), .ZN(n25709) );
  AND2_X1 U26070 ( .A1(b_8_), .A2(n26076), .ZN(n26075) );
  OR2_X1 U26071 ( .A1(n26077), .A2(n16981), .ZN(n26076) );
  AND2_X1 U26072 ( .A1(a_30_), .A2(n15637), .ZN(n26077) );
  AND2_X1 U26073 ( .A1(b_7_), .A2(n26078), .ZN(n26074) );
  OR2_X1 U26074 ( .A1(n26079), .A2(n14817), .ZN(n26078) );
  AND2_X1 U26075 ( .A1(a_31_), .A2(n15592), .ZN(n26079) );
  OR2_X1 U26076 ( .A1(n25717), .A2(n25714), .ZN(n26070) );
  OR2_X1 U26077 ( .A1(n26080), .A2(n26081), .ZN(n25714) );
  AND2_X1 U26078 ( .A1(n26082), .A2(n26083), .ZN(n26081) );
  INV_X1 U26079 ( .A(n26084), .ZN(n26080) );
  OR2_X1 U26080 ( .A1(n26082), .A2(n26083), .ZN(n26084) );
  OR2_X1 U26081 ( .A1(n26085), .A2(n26086), .ZN(n26082) );
  AND2_X1 U26082 ( .A1(n26087), .A2(n26088), .ZN(n26086) );
  AND2_X1 U26083 ( .A1(n26089), .A2(n26090), .ZN(n26085) );
  OR2_X1 U26084 ( .A1(n14891), .A2(n15558), .ZN(n25717) );
  OR2_X1 U26085 ( .A1(n25728), .A2(n25725), .ZN(n26067) );
  OR2_X1 U26086 ( .A1(n26091), .A2(n26092), .ZN(n25725) );
  INV_X1 U26087 ( .A(n26093), .ZN(n26092) );
  OR2_X1 U26088 ( .A1(n26094), .A2(n26095), .ZN(n26093) );
  AND2_X1 U26089 ( .A1(n26095), .A2(n26094), .ZN(n26091) );
  AND2_X1 U26090 ( .A1(n26096), .A2(n26097), .ZN(n26094) );
  OR2_X1 U26091 ( .A1(n26098), .A2(n26099), .ZN(n26097) );
  INV_X1 U26092 ( .A(n26100), .ZN(n26099) );
  OR2_X1 U26093 ( .A1(n26100), .A2(n26101), .ZN(n26096) );
  INV_X1 U26094 ( .A(n26098), .ZN(n26101) );
  OR2_X1 U26095 ( .A1(n14936), .A2(n15558), .ZN(n25728) );
  OR2_X1 U26096 ( .A1(n25739), .A2(n25736), .ZN(n26064) );
  OR2_X1 U26097 ( .A1(n26102), .A2(n26103), .ZN(n25736) );
  INV_X1 U26098 ( .A(n26104), .ZN(n26103) );
  OR2_X1 U26099 ( .A1(n26105), .A2(n26106), .ZN(n26104) );
  AND2_X1 U26100 ( .A1(n26106), .A2(n26105), .ZN(n26102) );
  AND2_X1 U26101 ( .A1(n26107), .A2(n26108), .ZN(n26105) );
  OR2_X1 U26102 ( .A1(n26109), .A2(n26110), .ZN(n26108) );
  INV_X1 U26103 ( .A(n26111), .ZN(n26110) );
  OR2_X1 U26104 ( .A1(n26111), .A2(n26112), .ZN(n26107) );
  INV_X1 U26105 ( .A(n26109), .ZN(n26112) );
  OR2_X1 U26106 ( .A1(n14970), .A2(n15558), .ZN(n25739) );
  OR2_X1 U26107 ( .A1(n25750), .A2(n25747), .ZN(n26061) );
  OR2_X1 U26108 ( .A1(n26113), .A2(n26114), .ZN(n25747) );
  INV_X1 U26109 ( .A(n26115), .ZN(n26114) );
  OR2_X1 U26110 ( .A1(n26116), .A2(n26117), .ZN(n26115) );
  AND2_X1 U26111 ( .A1(n26117), .A2(n26116), .ZN(n26113) );
  AND2_X1 U26112 ( .A1(n26118), .A2(n26119), .ZN(n26116) );
  OR2_X1 U26113 ( .A1(n26120), .A2(n26121), .ZN(n26119) );
  INV_X1 U26114 ( .A(n26122), .ZN(n26121) );
  OR2_X1 U26115 ( .A1(n26122), .A2(n26123), .ZN(n26118) );
  INV_X1 U26116 ( .A(n26120), .ZN(n26123) );
  OR2_X1 U26117 ( .A1(n15004), .A2(n15558), .ZN(n25750) );
  OR2_X1 U26118 ( .A1(n25761), .A2(n25758), .ZN(n26058) );
  OR2_X1 U26119 ( .A1(n26124), .A2(n26125), .ZN(n25758) );
  INV_X1 U26120 ( .A(n26126), .ZN(n26125) );
  OR2_X1 U26121 ( .A1(n26127), .A2(n26128), .ZN(n26126) );
  AND2_X1 U26122 ( .A1(n26128), .A2(n26127), .ZN(n26124) );
  AND2_X1 U26123 ( .A1(n26129), .A2(n26130), .ZN(n26127) );
  OR2_X1 U26124 ( .A1(n26131), .A2(n26132), .ZN(n26130) );
  INV_X1 U26125 ( .A(n26133), .ZN(n26132) );
  OR2_X1 U26126 ( .A1(n26133), .A2(n26134), .ZN(n26129) );
  INV_X1 U26127 ( .A(n26131), .ZN(n26134) );
  OR2_X1 U26128 ( .A1(n15038), .A2(n15558), .ZN(n25761) );
  OR2_X1 U26129 ( .A1(n25772), .A2(n25769), .ZN(n26055) );
  OR2_X1 U26130 ( .A1(n26135), .A2(n26136), .ZN(n25769) );
  INV_X1 U26131 ( .A(n26137), .ZN(n26136) );
  OR2_X1 U26132 ( .A1(n26138), .A2(n26139), .ZN(n26137) );
  AND2_X1 U26133 ( .A1(n26139), .A2(n26138), .ZN(n26135) );
  AND2_X1 U26134 ( .A1(n26140), .A2(n26141), .ZN(n26138) );
  OR2_X1 U26135 ( .A1(n26142), .A2(n26143), .ZN(n26141) );
  INV_X1 U26136 ( .A(n26144), .ZN(n26143) );
  OR2_X1 U26137 ( .A1(n26144), .A2(n26145), .ZN(n26140) );
  INV_X1 U26138 ( .A(n26142), .ZN(n26145) );
  OR2_X1 U26139 ( .A1(n15072), .A2(n15558), .ZN(n25772) );
  OR2_X1 U26140 ( .A1(n25783), .A2(n25780), .ZN(n26052) );
  OR2_X1 U26141 ( .A1(n26146), .A2(n26147), .ZN(n25780) );
  INV_X1 U26142 ( .A(n26148), .ZN(n26147) );
  OR2_X1 U26143 ( .A1(n26149), .A2(n26150), .ZN(n26148) );
  AND2_X1 U26144 ( .A1(n26150), .A2(n26149), .ZN(n26146) );
  AND2_X1 U26145 ( .A1(n26151), .A2(n26152), .ZN(n26149) );
  OR2_X1 U26146 ( .A1(n26153), .A2(n26154), .ZN(n26152) );
  INV_X1 U26147 ( .A(n26155), .ZN(n26154) );
  OR2_X1 U26148 ( .A1(n26155), .A2(n26156), .ZN(n26151) );
  INV_X1 U26149 ( .A(n26153), .ZN(n26156) );
  OR2_X1 U26150 ( .A1(n15106), .A2(n15558), .ZN(n25783) );
  OR2_X1 U26151 ( .A1(n26157), .A2(n26158), .ZN(n25791) );
  INV_X1 U26152 ( .A(n26159), .ZN(n26158) );
  OR2_X1 U26153 ( .A1(n26160), .A2(n26161), .ZN(n26159) );
  AND2_X1 U26154 ( .A1(n26161), .A2(n26160), .ZN(n26157) );
  AND2_X1 U26155 ( .A1(n26162), .A2(n26163), .ZN(n26160) );
  OR2_X1 U26156 ( .A1(n26164), .A2(n26165), .ZN(n26163) );
  INV_X1 U26157 ( .A(n26166), .ZN(n26165) );
  OR2_X1 U26158 ( .A1(n26166), .A2(n26167), .ZN(n26162) );
  INV_X1 U26159 ( .A(n26164), .ZN(n26167) );
  OR2_X1 U26160 ( .A1(n25808), .A2(n25802), .ZN(n26046) );
  OR2_X1 U26161 ( .A1(n26168), .A2(n26169), .ZN(n25802) );
  INV_X1 U26162 ( .A(n26170), .ZN(n26169) );
  OR2_X1 U26163 ( .A1(n26171), .A2(n26172), .ZN(n26170) );
  AND2_X1 U26164 ( .A1(n26172), .A2(n26171), .ZN(n26168) );
  AND2_X1 U26165 ( .A1(n26173), .A2(n26174), .ZN(n26171) );
  INV_X1 U26166 ( .A(n26175), .ZN(n26174) );
  AND2_X1 U26167 ( .A1(n26176), .A2(n26177), .ZN(n26175) );
  OR2_X1 U26168 ( .A1(n26177), .A2(n26176), .ZN(n26173) );
  INV_X1 U26169 ( .A(n26178), .ZN(n26176) );
  OR2_X1 U26170 ( .A1(n15174), .A2(n15558), .ZN(n25808) );
  INV_X1 U26171 ( .A(b_9_), .ZN(n15558) );
  AND2_X1 U26172 ( .A1(n26179), .A2(n26180), .ZN(n25813) );
  INV_X1 U26173 ( .A(n26181), .ZN(n26180) );
  AND2_X1 U26174 ( .A1(n26182), .A2(n26183), .ZN(n26181) );
  OR2_X1 U26175 ( .A1(n26183), .A2(n26182), .ZN(n26179) );
  OR2_X1 U26176 ( .A1(n26184), .A2(n26185), .ZN(n26182) );
  AND2_X1 U26177 ( .A1(n26186), .A2(n26187), .ZN(n26185) );
  INV_X1 U26178 ( .A(n26188), .ZN(n26186) );
  AND2_X1 U26179 ( .A1(n26189), .A2(n26188), .ZN(n26184) );
  INV_X1 U26180 ( .A(n26187), .ZN(n26189) );
  AND2_X1 U26181 ( .A1(n26190), .A2(n26191), .ZN(n25824) );
  INV_X1 U26182 ( .A(n26192), .ZN(n26191) );
  AND2_X1 U26183 ( .A1(n26193), .A2(n26194), .ZN(n26192) );
  OR2_X1 U26184 ( .A1(n26194), .A2(n26193), .ZN(n26190) );
  OR2_X1 U26185 ( .A1(n26195), .A2(n26196), .ZN(n26193) );
  AND2_X1 U26186 ( .A1(n26197), .A2(n26198), .ZN(n26196) );
  INV_X1 U26187 ( .A(n26199), .ZN(n26197) );
  AND2_X1 U26188 ( .A1(n26200), .A2(n26199), .ZN(n26195) );
  INV_X1 U26189 ( .A(n26198), .ZN(n26200) );
  AND2_X1 U26190 ( .A1(n26201), .A2(n26202), .ZN(n25835) );
  INV_X1 U26191 ( .A(n26203), .ZN(n26202) );
  AND2_X1 U26192 ( .A1(n26204), .A2(n26205), .ZN(n26203) );
  OR2_X1 U26193 ( .A1(n26205), .A2(n26204), .ZN(n26201) );
  OR2_X1 U26194 ( .A1(n26206), .A2(n26207), .ZN(n26204) );
  AND2_X1 U26195 ( .A1(n26208), .A2(n26209), .ZN(n26207) );
  INV_X1 U26196 ( .A(n26210), .ZN(n26208) );
  AND2_X1 U26197 ( .A1(n26211), .A2(n26210), .ZN(n26206) );
  INV_X1 U26198 ( .A(n26209), .ZN(n26211) );
  AND2_X1 U26199 ( .A1(n26212), .A2(n26213), .ZN(n25846) );
  INV_X1 U26200 ( .A(n26214), .ZN(n26213) );
  AND2_X1 U26201 ( .A1(n26215), .A2(n26216), .ZN(n26214) );
  OR2_X1 U26202 ( .A1(n26216), .A2(n26215), .ZN(n26212) );
  OR2_X1 U26203 ( .A1(n26217), .A2(n26218), .ZN(n26215) );
  AND2_X1 U26204 ( .A1(n26219), .A2(n26220), .ZN(n26218) );
  INV_X1 U26205 ( .A(n26221), .ZN(n26219) );
  AND2_X1 U26206 ( .A1(n26222), .A2(n26221), .ZN(n26217) );
  INV_X1 U26207 ( .A(n26220), .ZN(n26222) );
  AND2_X1 U26208 ( .A1(n26223), .A2(n26224), .ZN(n25857) );
  INV_X1 U26209 ( .A(n26225), .ZN(n26224) );
  AND2_X1 U26210 ( .A1(n26226), .A2(n26227), .ZN(n26225) );
  OR2_X1 U26211 ( .A1(n26227), .A2(n26226), .ZN(n26223) );
  OR2_X1 U26212 ( .A1(n26228), .A2(n26229), .ZN(n26226) );
  AND2_X1 U26213 ( .A1(n26230), .A2(n26231), .ZN(n26229) );
  INV_X1 U26214 ( .A(n26232), .ZN(n26230) );
  AND2_X1 U26215 ( .A1(n26233), .A2(n26232), .ZN(n26228) );
  INV_X1 U26216 ( .A(n26231), .ZN(n26233) );
  AND2_X1 U26217 ( .A1(n26234), .A2(n26235), .ZN(n25868) );
  INV_X1 U26218 ( .A(n26236), .ZN(n26235) );
  AND2_X1 U26219 ( .A1(n26237), .A2(n26238), .ZN(n26236) );
  OR2_X1 U26220 ( .A1(n26238), .A2(n26237), .ZN(n26234) );
  OR2_X1 U26221 ( .A1(n26239), .A2(n26240), .ZN(n26237) );
  AND2_X1 U26222 ( .A1(n26241), .A2(n26242), .ZN(n26240) );
  INV_X1 U26223 ( .A(n26243), .ZN(n26241) );
  AND2_X1 U26224 ( .A1(n26244), .A2(n26243), .ZN(n26239) );
  INV_X1 U26225 ( .A(n26242), .ZN(n26244) );
  AND2_X1 U26226 ( .A1(n26245), .A2(n26246), .ZN(n25879) );
  INV_X1 U26227 ( .A(n26247), .ZN(n26246) );
  AND2_X1 U26228 ( .A1(n26248), .A2(n26249), .ZN(n26247) );
  OR2_X1 U26229 ( .A1(n26249), .A2(n26248), .ZN(n26245) );
  OR2_X1 U26230 ( .A1(n26250), .A2(n26251), .ZN(n26248) );
  AND2_X1 U26231 ( .A1(n26252), .A2(n26253), .ZN(n26251) );
  INV_X1 U26232 ( .A(n26254), .ZN(n26252) );
  AND2_X1 U26233 ( .A1(n26255), .A2(n26254), .ZN(n26250) );
  INV_X1 U26234 ( .A(n26253), .ZN(n26255) );
  AND2_X1 U26235 ( .A1(n26256), .A2(n26257), .ZN(n25890) );
  INV_X1 U26236 ( .A(n26258), .ZN(n26257) );
  AND2_X1 U26237 ( .A1(n26259), .A2(n26260), .ZN(n26258) );
  OR2_X1 U26238 ( .A1(n26260), .A2(n26259), .ZN(n26256) );
  OR2_X1 U26239 ( .A1(n26261), .A2(n26262), .ZN(n26259) );
  AND2_X1 U26240 ( .A1(n26263), .A2(n26264), .ZN(n26262) );
  INV_X1 U26241 ( .A(n26265), .ZN(n26263) );
  AND2_X1 U26242 ( .A1(n26266), .A2(n26265), .ZN(n26261) );
  INV_X1 U26243 ( .A(n26264), .ZN(n26266) );
  AND2_X1 U26244 ( .A1(n26267), .A2(n26268), .ZN(n25901) );
  INV_X1 U26245 ( .A(n26269), .ZN(n26268) );
  AND2_X1 U26246 ( .A1(n26270), .A2(n26271), .ZN(n26269) );
  OR2_X1 U26247 ( .A1(n26271), .A2(n26270), .ZN(n26267) );
  OR2_X1 U26248 ( .A1(n26272), .A2(n26273), .ZN(n26270) );
  AND2_X1 U26249 ( .A1(n26274), .A2(n26275), .ZN(n26273) );
  INV_X1 U26250 ( .A(n26276), .ZN(n26274) );
  AND2_X1 U26251 ( .A1(n26277), .A2(n26276), .ZN(n26272) );
  INV_X1 U26252 ( .A(n26275), .ZN(n26277) );
  AND2_X1 U26253 ( .A1(n26278), .A2(n26279), .ZN(n25912) );
  INV_X1 U26254 ( .A(n26280), .ZN(n26279) );
  AND2_X1 U26255 ( .A1(n26281), .A2(n26282), .ZN(n26280) );
  OR2_X1 U26256 ( .A1(n26282), .A2(n26281), .ZN(n26278) );
  OR2_X1 U26257 ( .A1(n26283), .A2(n26284), .ZN(n26281) );
  AND2_X1 U26258 ( .A1(n26285), .A2(n26286), .ZN(n26284) );
  INV_X1 U26259 ( .A(n26287), .ZN(n26285) );
  AND2_X1 U26260 ( .A1(n26288), .A2(n26287), .ZN(n26283) );
  INV_X1 U26261 ( .A(n26286), .ZN(n26288) );
  AND2_X1 U26262 ( .A1(n26289), .A2(n26290), .ZN(n25923) );
  INV_X1 U26263 ( .A(n26291), .ZN(n26290) );
  AND2_X1 U26264 ( .A1(n26292), .A2(n26293), .ZN(n26291) );
  OR2_X1 U26265 ( .A1(n26293), .A2(n26292), .ZN(n26289) );
  OR2_X1 U26266 ( .A1(n26294), .A2(n26295), .ZN(n26292) );
  AND2_X1 U26267 ( .A1(n26296), .A2(n26297), .ZN(n26295) );
  INV_X1 U26268 ( .A(n26298), .ZN(n26296) );
  AND2_X1 U26269 ( .A1(n26299), .A2(n26298), .ZN(n26294) );
  INV_X1 U26270 ( .A(n26297), .ZN(n26299) );
  AND2_X1 U26271 ( .A1(n26300), .A2(n26301), .ZN(n25933) );
  INV_X1 U26272 ( .A(n26302), .ZN(n26301) );
  AND2_X1 U26273 ( .A1(n26303), .A2(n26304), .ZN(n26302) );
  OR2_X1 U26274 ( .A1(n26304), .A2(n26303), .ZN(n26300) );
  OR2_X1 U26275 ( .A1(n26305), .A2(n26306), .ZN(n26303) );
  AND2_X1 U26276 ( .A1(n26307), .A2(n26308), .ZN(n26306) );
  INV_X1 U26277 ( .A(n26309), .ZN(n26307) );
  AND2_X1 U26278 ( .A1(n26310), .A2(n26309), .ZN(n26305) );
  INV_X1 U26279 ( .A(n26308), .ZN(n26310) );
  AND2_X1 U26280 ( .A1(n26311), .A2(n26312), .ZN(n25944) );
  INV_X1 U26281 ( .A(n26313), .ZN(n26312) );
  AND2_X1 U26282 ( .A1(n26314), .A2(n26315), .ZN(n26313) );
  OR2_X1 U26283 ( .A1(n26315), .A2(n26314), .ZN(n26311) );
  OR2_X1 U26284 ( .A1(n26316), .A2(n26317), .ZN(n26314) );
  AND2_X1 U26285 ( .A1(n26318), .A2(n26319), .ZN(n26317) );
  INV_X1 U26286 ( .A(n15891), .ZN(n26318) );
  AND2_X1 U26287 ( .A1(n26320), .A2(n15891), .ZN(n26316) );
  INV_X1 U26288 ( .A(n26319), .ZN(n26320) );
  AND2_X1 U26289 ( .A1(n26321), .A2(n26322), .ZN(n25955) );
  INV_X1 U26290 ( .A(n26323), .ZN(n26322) );
  AND2_X1 U26291 ( .A1(n26324), .A2(n26325), .ZN(n26323) );
  OR2_X1 U26292 ( .A1(n26325), .A2(n26324), .ZN(n26321) );
  OR2_X1 U26293 ( .A1(n26326), .A2(n26327), .ZN(n26324) );
  AND2_X1 U26294 ( .A1(n26328), .A2(n26329), .ZN(n26327) );
  INV_X1 U26295 ( .A(n26330), .ZN(n26328) );
  AND2_X1 U26296 ( .A1(n26331), .A2(n26330), .ZN(n26326) );
  INV_X1 U26297 ( .A(n26329), .ZN(n26331) );
  AND2_X1 U26298 ( .A1(n26332), .A2(n26333), .ZN(n25966) );
  INV_X1 U26299 ( .A(n26334), .ZN(n26333) );
  AND2_X1 U26300 ( .A1(n26335), .A2(n26336), .ZN(n26334) );
  OR2_X1 U26301 ( .A1(n26336), .A2(n26335), .ZN(n26332) );
  OR2_X1 U26302 ( .A1(n26337), .A2(n26338), .ZN(n26335) );
  AND2_X1 U26303 ( .A1(n26339), .A2(n26340), .ZN(n26338) );
  INV_X1 U26304 ( .A(n26341), .ZN(n26339) );
  AND2_X1 U26305 ( .A1(n26342), .A2(n26341), .ZN(n26337) );
  INV_X1 U26306 ( .A(n26340), .ZN(n26342) );
  AND2_X1 U26307 ( .A1(n26343), .A2(n26344), .ZN(n25977) );
  INV_X1 U26308 ( .A(n26345), .ZN(n26344) );
  AND2_X1 U26309 ( .A1(n26346), .A2(n26347), .ZN(n26345) );
  OR2_X1 U26310 ( .A1(n26347), .A2(n26346), .ZN(n26343) );
  OR2_X1 U26311 ( .A1(n26348), .A2(n26349), .ZN(n26346) );
  AND2_X1 U26312 ( .A1(n26350), .A2(n26351), .ZN(n26349) );
  INV_X1 U26313 ( .A(n26352), .ZN(n26350) );
  AND2_X1 U26314 ( .A1(n26353), .A2(n26352), .ZN(n26348) );
  INV_X1 U26315 ( .A(n26351), .ZN(n26353) );
  AND2_X1 U26316 ( .A1(n26354), .A2(n26355), .ZN(n16639) );
  INV_X1 U26317 ( .A(n26356), .ZN(n26355) );
  AND2_X1 U26318 ( .A1(n26357), .A2(n26358), .ZN(n26356) );
  OR2_X1 U26319 ( .A1(n26358), .A2(n26357), .ZN(n26354) );
  OR2_X1 U26320 ( .A1(n26359), .A2(n26360), .ZN(n26357) );
  AND2_X1 U26321 ( .A1(n26361), .A2(n26362), .ZN(n26360) );
  INV_X1 U26322 ( .A(n26363), .ZN(n26361) );
  AND2_X1 U26323 ( .A1(n26364), .A2(n26363), .ZN(n26359) );
  INV_X1 U26324 ( .A(n26362), .ZN(n26364) );
  AND2_X1 U26325 ( .A1(n26365), .A2(n26366), .ZN(n16576) );
  INV_X1 U26326 ( .A(n26367), .ZN(n26366) );
  AND2_X1 U26327 ( .A1(n26368), .A2(n26369), .ZN(n26367) );
  OR2_X1 U26328 ( .A1(n26369), .A2(n26368), .ZN(n26365) );
  OR2_X1 U26329 ( .A1(n26370), .A2(n26371), .ZN(n26368) );
  AND2_X1 U26330 ( .A1(n26372), .A2(n26373), .ZN(n26371) );
  INV_X1 U26331 ( .A(n26374), .ZN(n26372) );
  AND2_X1 U26332 ( .A1(n26375), .A2(n26374), .ZN(n26370) );
  INV_X1 U26333 ( .A(n26373), .ZN(n26375) );
  AND2_X1 U26334 ( .A1(n26376), .A2(n26377), .ZN(n16523) );
  INV_X1 U26335 ( .A(n26378), .ZN(n26377) );
  AND2_X1 U26336 ( .A1(n26379), .A2(n26380), .ZN(n26378) );
  OR2_X1 U26337 ( .A1(n26380), .A2(n26379), .ZN(n26376) );
  OR2_X1 U26338 ( .A1(n26381), .A2(n26382), .ZN(n26379) );
  AND2_X1 U26339 ( .A1(n26383), .A2(n26384), .ZN(n26382) );
  INV_X1 U26340 ( .A(n26385), .ZN(n26383) );
  AND2_X1 U26341 ( .A1(n26386), .A2(n26385), .ZN(n26381) );
  INV_X1 U26342 ( .A(n26384), .ZN(n26386) );
  AND2_X1 U26343 ( .A1(n26387), .A2(n26388), .ZN(n16487) );
  INV_X1 U26344 ( .A(n26389), .ZN(n26388) );
  AND2_X1 U26345 ( .A1(n26390), .A2(n26391), .ZN(n26389) );
  OR2_X1 U26346 ( .A1(n26391), .A2(n26390), .ZN(n26387) );
  OR2_X1 U26347 ( .A1(n26392), .A2(n26393), .ZN(n26390) );
  AND2_X1 U26348 ( .A1(n26394), .A2(n26395), .ZN(n26393) );
  INV_X1 U26349 ( .A(n26396), .ZN(n26394) );
  AND2_X1 U26350 ( .A1(n26397), .A2(n26396), .ZN(n26392) );
  INV_X1 U26351 ( .A(n26395), .ZN(n26397) );
  AND2_X1 U26352 ( .A1(n26398), .A2(n26399), .ZN(n16471) );
  INV_X1 U26353 ( .A(n26400), .ZN(n26399) );
  AND2_X1 U26354 ( .A1(n26401), .A2(n16456), .ZN(n26400) );
  OR2_X1 U26355 ( .A1(n16456), .A2(n26401), .ZN(n26398) );
  OR2_X1 U26356 ( .A1(n26402), .A2(n26403), .ZN(n26401) );
  AND2_X1 U26357 ( .A1(n26404), .A2(n16455), .ZN(n26403) );
  INV_X1 U26358 ( .A(n16454), .ZN(n26404) );
  AND2_X1 U26359 ( .A1(n26405), .A2(n16454), .ZN(n26402) );
  OR2_X1 U26360 ( .A1(n16512), .A2(n15592), .ZN(n16454) );
  INV_X1 U26361 ( .A(n16455), .ZN(n26405) );
  OR2_X1 U26362 ( .A1(n26406), .A2(n26407), .ZN(n16455) );
  AND2_X1 U26363 ( .A1(n26396), .A2(n26395), .ZN(n26407) );
  AND2_X1 U26364 ( .A1(n26391), .A2(n26408), .ZN(n26406) );
  OR2_X1 U26365 ( .A1(n26395), .A2(n26396), .ZN(n26408) );
  OR2_X1 U26366 ( .A1(n15842), .A2(n15592), .ZN(n26396) );
  OR2_X1 U26367 ( .A1(n26409), .A2(n26410), .ZN(n26395) );
  AND2_X1 U26368 ( .A1(n26385), .A2(n26384), .ZN(n26410) );
  AND2_X1 U26369 ( .A1(n26380), .A2(n26411), .ZN(n26409) );
  OR2_X1 U26370 ( .A1(n26384), .A2(n26385), .ZN(n26411) );
  OR2_X1 U26371 ( .A1(n15808), .A2(n15592), .ZN(n26385) );
  OR2_X1 U26372 ( .A1(n26412), .A2(n26413), .ZN(n26384) );
  AND2_X1 U26373 ( .A1(n26374), .A2(n26373), .ZN(n26413) );
  AND2_X1 U26374 ( .A1(n26369), .A2(n26414), .ZN(n26412) );
  OR2_X1 U26375 ( .A1(n26373), .A2(n26374), .ZN(n26414) );
  OR2_X1 U26376 ( .A1(n15774), .A2(n15592), .ZN(n26374) );
  OR2_X1 U26377 ( .A1(n26415), .A2(n26416), .ZN(n26373) );
  AND2_X1 U26378 ( .A1(n26363), .A2(n26362), .ZN(n26416) );
  AND2_X1 U26379 ( .A1(n26358), .A2(n26417), .ZN(n26415) );
  OR2_X1 U26380 ( .A1(n26362), .A2(n26363), .ZN(n26417) );
  OR2_X1 U26381 ( .A1(n15740), .A2(n15592), .ZN(n26363) );
  OR2_X1 U26382 ( .A1(n26418), .A2(n26419), .ZN(n26362) );
  AND2_X1 U26383 ( .A1(n26352), .A2(n26351), .ZN(n26419) );
  AND2_X1 U26384 ( .A1(n26347), .A2(n26420), .ZN(n26418) );
  OR2_X1 U26385 ( .A1(n26351), .A2(n26352), .ZN(n26420) );
  OR2_X1 U26386 ( .A1(n15706), .A2(n15592), .ZN(n26352) );
  OR2_X1 U26387 ( .A1(n26421), .A2(n26422), .ZN(n26351) );
  AND2_X1 U26388 ( .A1(n26341), .A2(n26340), .ZN(n26422) );
  AND2_X1 U26389 ( .A1(n26336), .A2(n26423), .ZN(n26421) );
  OR2_X1 U26390 ( .A1(n26340), .A2(n26341), .ZN(n26423) );
  OR2_X1 U26391 ( .A1(n15672), .A2(n15592), .ZN(n26341) );
  OR2_X1 U26392 ( .A1(n26424), .A2(n26425), .ZN(n26340) );
  AND2_X1 U26393 ( .A1(n26330), .A2(n26329), .ZN(n26425) );
  AND2_X1 U26394 ( .A1(n26325), .A2(n26426), .ZN(n26424) );
  OR2_X1 U26395 ( .A1(n26329), .A2(n26330), .ZN(n26426) );
  OR2_X1 U26396 ( .A1(n15638), .A2(n15592), .ZN(n26330) );
  OR2_X1 U26397 ( .A1(n26427), .A2(n26428), .ZN(n26329) );
  AND2_X1 U26398 ( .A1(n15891), .A2(n26319), .ZN(n26428) );
  AND2_X1 U26399 ( .A1(n26315), .A2(n26429), .ZN(n26427) );
  OR2_X1 U26400 ( .A1(n26319), .A2(n15891), .ZN(n26429) );
  OR2_X1 U26401 ( .A1(n15593), .A2(n15592), .ZN(n15891) );
  OR2_X1 U26402 ( .A1(n26430), .A2(n26431), .ZN(n26319) );
  AND2_X1 U26403 ( .A1(n26309), .A2(n26308), .ZN(n26431) );
  AND2_X1 U26404 ( .A1(n26304), .A2(n26432), .ZN(n26430) );
  OR2_X1 U26405 ( .A1(n26308), .A2(n26309), .ZN(n26432) );
  OR2_X1 U26406 ( .A1(n15559), .A2(n15592), .ZN(n26309) );
  OR2_X1 U26407 ( .A1(n26433), .A2(n26434), .ZN(n26308) );
  AND2_X1 U26408 ( .A1(n26298), .A2(n26297), .ZN(n26434) );
  AND2_X1 U26409 ( .A1(n26293), .A2(n26435), .ZN(n26433) );
  OR2_X1 U26410 ( .A1(n26297), .A2(n26298), .ZN(n26435) );
  OR2_X1 U26411 ( .A1(n15525), .A2(n15592), .ZN(n26298) );
  OR2_X1 U26412 ( .A1(n26436), .A2(n26437), .ZN(n26297) );
  AND2_X1 U26413 ( .A1(n26287), .A2(n26286), .ZN(n26437) );
  AND2_X1 U26414 ( .A1(n26282), .A2(n26438), .ZN(n26436) );
  OR2_X1 U26415 ( .A1(n26286), .A2(n26287), .ZN(n26438) );
  OR2_X1 U26416 ( .A1(n15491), .A2(n15592), .ZN(n26287) );
  OR2_X1 U26417 ( .A1(n26439), .A2(n26440), .ZN(n26286) );
  AND2_X1 U26418 ( .A1(n26276), .A2(n26275), .ZN(n26440) );
  AND2_X1 U26419 ( .A1(n26271), .A2(n26441), .ZN(n26439) );
  OR2_X1 U26420 ( .A1(n26275), .A2(n26276), .ZN(n26441) );
  OR2_X1 U26421 ( .A1(n15457), .A2(n15592), .ZN(n26276) );
  OR2_X1 U26422 ( .A1(n26442), .A2(n26443), .ZN(n26275) );
  AND2_X1 U26423 ( .A1(n26265), .A2(n26264), .ZN(n26443) );
  AND2_X1 U26424 ( .A1(n26260), .A2(n26444), .ZN(n26442) );
  OR2_X1 U26425 ( .A1(n26264), .A2(n26265), .ZN(n26444) );
  OR2_X1 U26426 ( .A1(n15423), .A2(n15592), .ZN(n26265) );
  OR2_X1 U26427 ( .A1(n26445), .A2(n26446), .ZN(n26264) );
  AND2_X1 U26428 ( .A1(n26254), .A2(n26253), .ZN(n26446) );
  AND2_X1 U26429 ( .A1(n26249), .A2(n26447), .ZN(n26445) );
  OR2_X1 U26430 ( .A1(n26253), .A2(n26254), .ZN(n26447) );
  OR2_X1 U26431 ( .A1(n15389), .A2(n15592), .ZN(n26254) );
  OR2_X1 U26432 ( .A1(n26448), .A2(n26449), .ZN(n26253) );
  AND2_X1 U26433 ( .A1(n26243), .A2(n26242), .ZN(n26449) );
  AND2_X1 U26434 ( .A1(n26238), .A2(n26450), .ZN(n26448) );
  OR2_X1 U26435 ( .A1(n26242), .A2(n26243), .ZN(n26450) );
  OR2_X1 U26436 ( .A1(n15355), .A2(n15592), .ZN(n26243) );
  OR2_X1 U26437 ( .A1(n26451), .A2(n26452), .ZN(n26242) );
  AND2_X1 U26438 ( .A1(n26232), .A2(n26231), .ZN(n26452) );
  AND2_X1 U26439 ( .A1(n26227), .A2(n26453), .ZN(n26451) );
  OR2_X1 U26440 ( .A1(n26231), .A2(n26232), .ZN(n26453) );
  OR2_X1 U26441 ( .A1(n15321), .A2(n15592), .ZN(n26232) );
  OR2_X1 U26442 ( .A1(n26454), .A2(n26455), .ZN(n26231) );
  AND2_X1 U26443 ( .A1(n26221), .A2(n26220), .ZN(n26455) );
  AND2_X1 U26444 ( .A1(n26216), .A2(n26456), .ZN(n26454) );
  OR2_X1 U26445 ( .A1(n26220), .A2(n26221), .ZN(n26456) );
  OR2_X1 U26446 ( .A1(n15287), .A2(n15592), .ZN(n26221) );
  OR2_X1 U26447 ( .A1(n26457), .A2(n26458), .ZN(n26220) );
  AND2_X1 U26448 ( .A1(n26210), .A2(n26209), .ZN(n26458) );
  AND2_X1 U26449 ( .A1(n26205), .A2(n26459), .ZN(n26457) );
  OR2_X1 U26450 ( .A1(n26209), .A2(n26210), .ZN(n26459) );
  OR2_X1 U26451 ( .A1(n15242), .A2(n15592), .ZN(n26210) );
  OR2_X1 U26452 ( .A1(n26460), .A2(n26461), .ZN(n26209) );
  AND2_X1 U26453 ( .A1(n26199), .A2(n26198), .ZN(n26461) );
  AND2_X1 U26454 ( .A1(n26194), .A2(n26462), .ZN(n26460) );
  OR2_X1 U26455 ( .A1(n26198), .A2(n26199), .ZN(n26462) );
  OR2_X1 U26456 ( .A1(n15208), .A2(n15592), .ZN(n26199) );
  OR2_X1 U26457 ( .A1(n26463), .A2(n26464), .ZN(n26198) );
  AND2_X1 U26458 ( .A1(n26188), .A2(n26187), .ZN(n26464) );
  AND2_X1 U26459 ( .A1(n26183), .A2(n26465), .ZN(n26463) );
  OR2_X1 U26460 ( .A1(n26187), .A2(n26188), .ZN(n26465) );
  OR2_X1 U26461 ( .A1(n15174), .A2(n15592), .ZN(n26188) );
  OR2_X1 U26462 ( .A1(n26466), .A2(n26467), .ZN(n26187) );
  AND2_X1 U26463 ( .A1(n26172), .A2(n26178), .ZN(n26467) );
  AND2_X1 U26464 ( .A1(n26468), .A2(n26177), .ZN(n26466) );
  OR2_X1 U26465 ( .A1(n26469), .A2(n26470), .ZN(n26177) );
  AND2_X1 U26466 ( .A1(n26164), .A2(n26166), .ZN(n26470) );
  AND2_X1 U26467 ( .A1(n26161), .A2(n26471), .ZN(n26469) );
  OR2_X1 U26468 ( .A1(n26166), .A2(n26164), .ZN(n26471) );
  OR2_X1 U26469 ( .A1(n15106), .A2(n15592), .ZN(n26164) );
  OR2_X1 U26470 ( .A1(n26472), .A2(n26473), .ZN(n26166) );
  AND2_X1 U26471 ( .A1(n26150), .A2(n26153), .ZN(n26473) );
  AND2_X1 U26472 ( .A1(n26474), .A2(n26155), .ZN(n26472) );
  OR2_X1 U26473 ( .A1(n26475), .A2(n26476), .ZN(n26155) );
  AND2_X1 U26474 ( .A1(n26139), .A2(n26142), .ZN(n26476) );
  AND2_X1 U26475 ( .A1(n26477), .A2(n26144), .ZN(n26475) );
  OR2_X1 U26476 ( .A1(n26478), .A2(n26479), .ZN(n26144) );
  AND2_X1 U26477 ( .A1(n26128), .A2(n26131), .ZN(n26479) );
  AND2_X1 U26478 ( .A1(n26480), .A2(n26133), .ZN(n26478) );
  OR2_X1 U26479 ( .A1(n26481), .A2(n26482), .ZN(n26133) );
  AND2_X1 U26480 ( .A1(n26117), .A2(n26120), .ZN(n26482) );
  AND2_X1 U26481 ( .A1(n26483), .A2(n26122), .ZN(n26481) );
  OR2_X1 U26482 ( .A1(n26484), .A2(n26485), .ZN(n26122) );
  AND2_X1 U26483 ( .A1(n26106), .A2(n26109), .ZN(n26485) );
  AND2_X1 U26484 ( .A1(n26486), .A2(n26111), .ZN(n26484) );
  OR2_X1 U26485 ( .A1(n26487), .A2(n26488), .ZN(n26111) );
  AND2_X1 U26486 ( .A1(n26095), .A2(n26098), .ZN(n26488) );
  AND2_X1 U26487 ( .A1(n26489), .A2(n26100), .ZN(n26487) );
  OR2_X1 U26488 ( .A1(n26490), .A2(n26491), .ZN(n26100) );
  AND2_X1 U26489 ( .A1(n26083), .A2(n26088), .ZN(n26491) );
  AND2_X1 U26490 ( .A1(n26087), .A2(n26492), .ZN(n26490) );
  OR2_X1 U26491 ( .A1(n26088), .A2(n26083), .ZN(n26492) );
  OR2_X1 U26492 ( .A1(n14857), .A2(n15592), .ZN(n26083) );
  INV_X1 U26493 ( .A(n26089), .ZN(n26088) );
  AND3_X1 U26494 ( .A1(b_8_), .A2(b_7_), .A3(n15957), .ZN(n26089) );
  INV_X1 U26495 ( .A(n26090), .ZN(n26087) );
  OR2_X1 U26496 ( .A1(n26493), .A2(n26494), .ZN(n26090) );
  AND2_X1 U26497 ( .A1(b_7_), .A2(n26495), .ZN(n26494) );
  OR2_X1 U26498 ( .A1(n26496), .A2(n16981), .ZN(n26495) );
  AND2_X1 U26499 ( .A1(a_30_), .A2(n15671), .ZN(n26496) );
  AND2_X1 U26500 ( .A1(b_6_), .A2(n26497), .ZN(n26493) );
  OR2_X1 U26501 ( .A1(n26498), .A2(n14817), .ZN(n26497) );
  AND2_X1 U26502 ( .A1(a_31_), .A2(n15637), .ZN(n26498) );
  OR2_X1 U26503 ( .A1(n26098), .A2(n26095), .ZN(n26489) );
  OR2_X1 U26504 ( .A1(n26499), .A2(n26500), .ZN(n26095) );
  AND2_X1 U26505 ( .A1(n26501), .A2(n26502), .ZN(n26500) );
  INV_X1 U26506 ( .A(n26503), .ZN(n26499) );
  OR2_X1 U26507 ( .A1(n26501), .A2(n26502), .ZN(n26503) );
  OR2_X1 U26508 ( .A1(n26504), .A2(n26505), .ZN(n26501) );
  AND2_X1 U26509 ( .A1(n26506), .A2(n26507), .ZN(n26505) );
  AND2_X1 U26510 ( .A1(n26508), .A2(n26509), .ZN(n26504) );
  OR2_X1 U26511 ( .A1(n14891), .A2(n15592), .ZN(n26098) );
  OR2_X1 U26512 ( .A1(n26109), .A2(n26106), .ZN(n26486) );
  OR2_X1 U26513 ( .A1(n26510), .A2(n26511), .ZN(n26106) );
  INV_X1 U26514 ( .A(n26512), .ZN(n26511) );
  OR2_X1 U26515 ( .A1(n26513), .A2(n26514), .ZN(n26512) );
  AND2_X1 U26516 ( .A1(n26514), .A2(n26513), .ZN(n26510) );
  AND2_X1 U26517 ( .A1(n26515), .A2(n26516), .ZN(n26513) );
  OR2_X1 U26518 ( .A1(n26517), .A2(n26518), .ZN(n26516) );
  INV_X1 U26519 ( .A(n26519), .ZN(n26518) );
  OR2_X1 U26520 ( .A1(n26519), .A2(n26520), .ZN(n26515) );
  INV_X1 U26521 ( .A(n26517), .ZN(n26520) );
  OR2_X1 U26522 ( .A1(n14936), .A2(n15592), .ZN(n26109) );
  OR2_X1 U26523 ( .A1(n26120), .A2(n26117), .ZN(n26483) );
  OR2_X1 U26524 ( .A1(n26521), .A2(n26522), .ZN(n26117) );
  INV_X1 U26525 ( .A(n26523), .ZN(n26522) );
  OR2_X1 U26526 ( .A1(n26524), .A2(n26525), .ZN(n26523) );
  AND2_X1 U26527 ( .A1(n26525), .A2(n26524), .ZN(n26521) );
  AND2_X1 U26528 ( .A1(n26526), .A2(n26527), .ZN(n26524) );
  OR2_X1 U26529 ( .A1(n26528), .A2(n26529), .ZN(n26527) );
  INV_X1 U26530 ( .A(n26530), .ZN(n26529) );
  OR2_X1 U26531 ( .A1(n26530), .A2(n26531), .ZN(n26526) );
  INV_X1 U26532 ( .A(n26528), .ZN(n26531) );
  OR2_X1 U26533 ( .A1(n14970), .A2(n15592), .ZN(n26120) );
  OR2_X1 U26534 ( .A1(n26131), .A2(n26128), .ZN(n26480) );
  OR2_X1 U26535 ( .A1(n26532), .A2(n26533), .ZN(n26128) );
  INV_X1 U26536 ( .A(n26534), .ZN(n26533) );
  OR2_X1 U26537 ( .A1(n26535), .A2(n26536), .ZN(n26534) );
  AND2_X1 U26538 ( .A1(n26536), .A2(n26535), .ZN(n26532) );
  AND2_X1 U26539 ( .A1(n26537), .A2(n26538), .ZN(n26535) );
  OR2_X1 U26540 ( .A1(n26539), .A2(n26540), .ZN(n26538) );
  INV_X1 U26541 ( .A(n26541), .ZN(n26540) );
  OR2_X1 U26542 ( .A1(n26541), .A2(n26542), .ZN(n26537) );
  INV_X1 U26543 ( .A(n26539), .ZN(n26542) );
  OR2_X1 U26544 ( .A1(n15004), .A2(n15592), .ZN(n26131) );
  OR2_X1 U26545 ( .A1(n26142), .A2(n26139), .ZN(n26477) );
  OR2_X1 U26546 ( .A1(n26543), .A2(n26544), .ZN(n26139) );
  INV_X1 U26547 ( .A(n26545), .ZN(n26544) );
  OR2_X1 U26548 ( .A1(n26546), .A2(n26547), .ZN(n26545) );
  AND2_X1 U26549 ( .A1(n26547), .A2(n26546), .ZN(n26543) );
  AND2_X1 U26550 ( .A1(n26548), .A2(n26549), .ZN(n26546) );
  OR2_X1 U26551 ( .A1(n26550), .A2(n26551), .ZN(n26549) );
  INV_X1 U26552 ( .A(n26552), .ZN(n26551) );
  OR2_X1 U26553 ( .A1(n26552), .A2(n26553), .ZN(n26548) );
  INV_X1 U26554 ( .A(n26550), .ZN(n26553) );
  OR2_X1 U26555 ( .A1(n15038), .A2(n15592), .ZN(n26142) );
  OR2_X1 U26556 ( .A1(n26153), .A2(n26150), .ZN(n26474) );
  OR2_X1 U26557 ( .A1(n26554), .A2(n26555), .ZN(n26150) );
  INV_X1 U26558 ( .A(n26556), .ZN(n26555) );
  OR2_X1 U26559 ( .A1(n26557), .A2(n26558), .ZN(n26556) );
  AND2_X1 U26560 ( .A1(n26558), .A2(n26557), .ZN(n26554) );
  AND2_X1 U26561 ( .A1(n26559), .A2(n26560), .ZN(n26557) );
  OR2_X1 U26562 ( .A1(n26561), .A2(n26562), .ZN(n26560) );
  INV_X1 U26563 ( .A(n26563), .ZN(n26562) );
  OR2_X1 U26564 ( .A1(n26563), .A2(n26564), .ZN(n26559) );
  INV_X1 U26565 ( .A(n26561), .ZN(n26564) );
  OR2_X1 U26566 ( .A1(n15072), .A2(n15592), .ZN(n26153) );
  OR2_X1 U26567 ( .A1(n26565), .A2(n26566), .ZN(n26161) );
  INV_X1 U26568 ( .A(n26567), .ZN(n26566) );
  OR2_X1 U26569 ( .A1(n26568), .A2(n26569), .ZN(n26567) );
  AND2_X1 U26570 ( .A1(n26569), .A2(n26568), .ZN(n26565) );
  AND2_X1 U26571 ( .A1(n26570), .A2(n26571), .ZN(n26568) );
  OR2_X1 U26572 ( .A1(n26572), .A2(n26573), .ZN(n26571) );
  INV_X1 U26573 ( .A(n26574), .ZN(n26573) );
  OR2_X1 U26574 ( .A1(n26574), .A2(n26575), .ZN(n26570) );
  INV_X1 U26575 ( .A(n26572), .ZN(n26575) );
  OR2_X1 U26576 ( .A1(n26178), .A2(n26172), .ZN(n26468) );
  OR2_X1 U26577 ( .A1(n26576), .A2(n26577), .ZN(n26172) );
  INV_X1 U26578 ( .A(n26578), .ZN(n26577) );
  OR2_X1 U26579 ( .A1(n26579), .A2(n26580), .ZN(n26578) );
  AND2_X1 U26580 ( .A1(n26580), .A2(n26579), .ZN(n26576) );
  AND2_X1 U26581 ( .A1(n26581), .A2(n26582), .ZN(n26579) );
  INV_X1 U26582 ( .A(n26583), .ZN(n26582) );
  AND2_X1 U26583 ( .A1(n26584), .A2(n26585), .ZN(n26583) );
  OR2_X1 U26584 ( .A1(n26585), .A2(n26584), .ZN(n26581) );
  INV_X1 U26585 ( .A(n26586), .ZN(n26584) );
  OR2_X1 U26586 ( .A1(n15140), .A2(n15592), .ZN(n26178) );
  INV_X1 U26587 ( .A(b_8_), .ZN(n15592) );
  AND2_X1 U26588 ( .A1(n26587), .A2(n26588), .ZN(n26183) );
  INV_X1 U26589 ( .A(n26589), .ZN(n26588) );
  AND2_X1 U26590 ( .A1(n26590), .A2(n26591), .ZN(n26589) );
  OR2_X1 U26591 ( .A1(n26591), .A2(n26590), .ZN(n26587) );
  OR2_X1 U26592 ( .A1(n26592), .A2(n26593), .ZN(n26590) );
  AND2_X1 U26593 ( .A1(n26594), .A2(n26595), .ZN(n26593) );
  INV_X1 U26594 ( .A(n26596), .ZN(n26594) );
  AND2_X1 U26595 ( .A1(n26597), .A2(n26596), .ZN(n26592) );
  INV_X1 U26596 ( .A(n26595), .ZN(n26597) );
  AND2_X1 U26597 ( .A1(n26598), .A2(n26599), .ZN(n26194) );
  INV_X1 U26598 ( .A(n26600), .ZN(n26599) );
  AND2_X1 U26599 ( .A1(n26601), .A2(n26602), .ZN(n26600) );
  OR2_X1 U26600 ( .A1(n26602), .A2(n26601), .ZN(n26598) );
  OR2_X1 U26601 ( .A1(n26603), .A2(n26604), .ZN(n26601) );
  AND2_X1 U26602 ( .A1(n26605), .A2(n26606), .ZN(n26604) );
  INV_X1 U26603 ( .A(n26607), .ZN(n26605) );
  AND2_X1 U26604 ( .A1(n26608), .A2(n26607), .ZN(n26603) );
  INV_X1 U26605 ( .A(n26606), .ZN(n26608) );
  AND2_X1 U26606 ( .A1(n26609), .A2(n26610), .ZN(n26205) );
  INV_X1 U26607 ( .A(n26611), .ZN(n26610) );
  AND2_X1 U26608 ( .A1(n26612), .A2(n26613), .ZN(n26611) );
  OR2_X1 U26609 ( .A1(n26613), .A2(n26612), .ZN(n26609) );
  OR2_X1 U26610 ( .A1(n26614), .A2(n26615), .ZN(n26612) );
  AND2_X1 U26611 ( .A1(n26616), .A2(n26617), .ZN(n26615) );
  INV_X1 U26612 ( .A(n26618), .ZN(n26616) );
  AND2_X1 U26613 ( .A1(n26619), .A2(n26618), .ZN(n26614) );
  INV_X1 U26614 ( .A(n26617), .ZN(n26619) );
  AND2_X1 U26615 ( .A1(n26620), .A2(n26621), .ZN(n26216) );
  INV_X1 U26616 ( .A(n26622), .ZN(n26621) );
  AND2_X1 U26617 ( .A1(n26623), .A2(n26624), .ZN(n26622) );
  OR2_X1 U26618 ( .A1(n26624), .A2(n26623), .ZN(n26620) );
  OR2_X1 U26619 ( .A1(n26625), .A2(n26626), .ZN(n26623) );
  AND2_X1 U26620 ( .A1(n26627), .A2(n26628), .ZN(n26626) );
  INV_X1 U26621 ( .A(n26629), .ZN(n26627) );
  AND2_X1 U26622 ( .A1(n26630), .A2(n26629), .ZN(n26625) );
  INV_X1 U26623 ( .A(n26628), .ZN(n26630) );
  AND2_X1 U26624 ( .A1(n26631), .A2(n26632), .ZN(n26227) );
  INV_X1 U26625 ( .A(n26633), .ZN(n26632) );
  AND2_X1 U26626 ( .A1(n26634), .A2(n26635), .ZN(n26633) );
  OR2_X1 U26627 ( .A1(n26635), .A2(n26634), .ZN(n26631) );
  OR2_X1 U26628 ( .A1(n26636), .A2(n26637), .ZN(n26634) );
  AND2_X1 U26629 ( .A1(n26638), .A2(n26639), .ZN(n26637) );
  INV_X1 U26630 ( .A(n26640), .ZN(n26638) );
  AND2_X1 U26631 ( .A1(n26641), .A2(n26640), .ZN(n26636) );
  INV_X1 U26632 ( .A(n26639), .ZN(n26641) );
  AND2_X1 U26633 ( .A1(n26642), .A2(n26643), .ZN(n26238) );
  INV_X1 U26634 ( .A(n26644), .ZN(n26643) );
  AND2_X1 U26635 ( .A1(n26645), .A2(n26646), .ZN(n26644) );
  OR2_X1 U26636 ( .A1(n26646), .A2(n26645), .ZN(n26642) );
  OR2_X1 U26637 ( .A1(n26647), .A2(n26648), .ZN(n26645) );
  AND2_X1 U26638 ( .A1(n26649), .A2(n26650), .ZN(n26648) );
  INV_X1 U26639 ( .A(n26651), .ZN(n26649) );
  AND2_X1 U26640 ( .A1(n26652), .A2(n26651), .ZN(n26647) );
  INV_X1 U26641 ( .A(n26650), .ZN(n26652) );
  AND2_X1 U26642 ( .A1(n26653), .A2(n26654), .ZN(n26249) );
  INV_X1 U26643 ( .A(n26655), .ZN(n26654) );
  AND2_X1 U26644 ( .A1(n26656), .A2(n26657), .ZN(n26655) );
  OR2_X1 U26645 ( .A1(n26657), .A2(n26656), .ZN(n26653) );
  OR2_X1 U26646 ( .A1(n26658), .A2(n26659), .ZN(n26656) );
  AND2_X1 U26647 ( .A1(n26660), .A2(n26661), .ZN(n26659) );
  INV_X1 U26648 ( .A(n26662), .ZN(n26660) );
  AND2_X1 U26649 ( .A1(n26663), .A2(n26662), .ZN(n26658) );
  INV_X1 U26650 ( .A(n26661), .ZN(n26663) );
  AND2_X1 U26651 ( .A1(n26664), .A2(n26665), .ZN(n26260) );
  INV_X1 U26652 ( .A(n26666), .ZN(n26665) );
  AND2_X1 U26653 ( .A1(n26667), .A2(n26668), .ZN(n26666) );
  OR2_X1 U26654 ( .A1(n26668), .A2(n26667), .ZN(n26664) );
  OR2_X1 U26655 ( .A1(n26669), .A2(n26670), .ZN(n26667) );
  AND2_X1 U26656 ( .A1(n26671), .A2(n26672), .ZN(n26670) );
  INV_X1 U26657 ( .A(n26673), .ZN(n26671) );
  AND2_X1 U26658 ( .A1(n26674), .A2(n26673), .ZN(n26669) );
  INV_X1 U26659 ( .A(n26672), .ZN(n26674) );
  AND2_X1 U26660 ( .A1(n26675), .A2(n26676), .ZN(n26271) );
  INV_X1 U26661 ( .A(n26677), .ZN(n26676) );
  AND2_X1 U26662 ( .A1(n26678), .A2(n26679), .ZN(n26677) );
  OR2_X1 U26663 ( .A1(n26679), .A2(n26678), .ZN(n26675) );
  OR2_X1 U26664 ( .A1(n26680), .A2(n26681), .ZN(n26678) );
  AND2_X1 U26665 ( .A1(n26682), .A2(n26683), .ZN(n26681) );
  INV_X1 U26666 ( .A(n26684), .ZN(n26682) );
  AND2_X1 U26667 ( .A1(n26685), .A2(n26684), .ZN(n26680) );
  INV_X1 U26668 ( .A(n26683), .ZN(n26685) );
  AND2_X1 U26669 ( .A1(n26686), .A2(n26687), .ZN(n26282) );
  INV_X1 U26670 ( .A(n26688), .ZN(n26687) );
  AND2_X1 U26671 ( .A1(n26689), .A2(n26690), .ZN(n26688) );
  OR2_X1 U26672 ( .A1(n26690), .A2(n26689), .ZN(n26686) );
  OR2_X1 U26673 ( .A1(n26691), .A2(n26692), .ZN(n26689) );
  AND2_X1 U26674 ( .A1(n26693), .A2(n26694), .ZN(n26692) );
  INV_X1 U26675 ( .A(n26695), .ZN(n26693) );
  AND2_X1 U26676 ( .A1(n26696), .A2(n26695), .ZN(n26691) );
  INV_X1 U26677 ( .A(n26694), .ZN(n26696) );
  AND2_X1 U26678 ( .A1(n26697), .A2(n26698), .ZN(n26293) );
  INV_X1 U26679 ( .A(n26699), .ZN(n26698) );
  AND2_X1 U26680 ( .A1(n26700), .A2(n26701), .ZN(n26699) );
  OR2_X1 U26681 ( .A1(n26701), .A2(n26700), .ZN(n26697) );
  OR2_X1 U26682 ( .A1(n26702), .A2(n26703), .ZN(n26700) );
  AND2_X1 U26683 ( .A1(n26704), .A2(n26705), .ZN(n26703) );
  INV_X1 U26684 ( .A(n26706), .ZN(n26704) );
  AND2_X1 U26685 ( .A1(n26707), .A2(n26706), .ZN(n26702) );
  INV_X1 U26686 ( .A(n26705), .ZN(n26707) );
  AND2_X1 U26687 ( .A1(n26708), .A2(n26709), .ZN(n26304) );
  INV_X1 U26688 ( .A(n26710), .ZN(n26709) );
  AND2_X1 U26689 ( .A1(n26711), .A2(n26712), .ZN(n26710) );
  OR2_X1 U26690 ( .A1(n26712), .A2(n26711), .ZN(n26708) );
  OR2_X1 U26691 ( .A1(n26713), .A2(n26714), .ZN(n26711) );
  AND2_X1 U26692 ( .A1(n26715), .A2(n26716), .ZN(n26714) );
  INV_X1 U26693 ( .A(n26717), .ZN(n26715) );
  AND2_X1 U26694 ( .A1(n26718), .A2(n26717), .ZN(n26713) );
  INV_X1 U26695 ( .A(n26716), .ZN(n26718) );
  AND2_X1 U26696 ( .A1(n26719), .A2(n26720), .ZN(n26315) );
  INV_X1 U26697 ( .A(n26721), .ZN(n26720) );
  AND2_X1 U26698 ( .A1(n26722), .A2(n26723), .ZN(n26721) );
  OR2_X1 U26699 ( .A1(n26723), .A2(n26722), .ZN(n26719) );
  OR2_X1 U26700 ( .A1(n26724), .A2(n26725), .ZN(n26722) );
  AND2_X1 U26701 ( .A1(n26726), .A2(n26727), .ZN(n26725) );
  INV_X1 U26702 ( .A(n26728), .ZN(n26726) );
  AND2_X1 U26703 ( .A1(n26729), .A2(n26728), .ZN(n26724) );
  INV_X1 U26704 ( .A(n26727), .ZN(n26729) );
  AND2_X1 U26705 ( .A1(n26730), .A2(n26731), .ZN(n26325) );
  INV_X1 U26706 ( .A(n26732), .ZN(n26731) );
  AND2_X1 U26707 ( .A1(n26733), .A2(n26734), .ZN(n26732) );
  OR2_X1 U26708 ( .A1(n26734), .A2(n26733), .ZN(n26730) );
  OR2_X1 U26709 ( .A1(n26735), .A2(n26736), .ZN(n26733) );
  AND2_X1 U26710 ( .A1(n26737), .A2(n26738), .ZN(n26736) );
  INV_X1 U26711 ( .A(n26739), .ZN(n26737) );
  AND2_X1 U26712 ( .A1(n26740), .A2(n26739), .ZN(n26735) );
  INV_X1 U26713 ( .A(n26738), .ZN(n26740) );
  AND2_X1 U26714 ( .A1(n26741), .A2(n26742), .ZN(n26336) );
  INV_X1 U26715 ( .A(n26743), .ZN(n26742) );
  AND2_X1 U26716 ( .A1(n26744), .A2(n26745), .ZN(n26743) );
  OR2_X1 U26717 ( .A1(n26745), .A2(n26744), .ZN(n26741) );
  OR2_X1 U26718 ( .A1(n26746), .A2(n26747), .ZN(n26744) );
  AND2_X1 U26719 ( .A1(n26748), .A2(n26749), .ZN(n26747) );
  INV_X1 U26720 ( .A(n15888), .ZN(n26748) );
  AND2_X1 U26721 ( .A1(n26750), .A2(n15888), .ZN(n26746) );
  INV_X1 U26722 ( .A(n26749), .ZN(n26750) );
  AND2_X1 U26723 ( .A1(n26751), .A2(n26752), .ZN(n26347) );
  INV_X1 U26724 ( .A(n26753), .ZN(n26752) );
  AND2_X1 U26725 ( .A1(n26754), .A2(n26755), .ZN(n26753) );
  OR2_X1 U26726 ( .A1(n26755), .A2(n26754), .ZN(n26751) );
  OR2_X1 U26727 ( .A1(n26756), .A2(n26757), .ZN(n26754) );
  AND2_X1 U26728 ( .A1(n26758), .A2(n26759), .ZN(n26757) );
  INV_X1 U26729 ( .A(n26760), .ZN(n26758) );
  AND2_X1 U26730 ( .A1(n26761), .A2(n26760), .ZN(n26756) );
  INV_X1 U26731 ( .A(n26759), .ZN(n26761) );
  AND2_X1 U26732 ( .A1(n26762), .A2(n26763), .ZN(n26358) );
  INV_X1 U26733 ( .A(n26764), .ZN(n26763) );
  AND2_X1 U26734 ( .A1(n26765), .A2(n26766), .ZN(n26764) );
  OR2_X1 U26735 ( .A1(n26766), .A2(n26765), .ZN(n26762) );
  OR2_X1 U26736 ( .A1(n26767), .A2(n26768), .ZN(n26765) );
  AND2_X1 U26737 ( .A1(n26769), .A2(n26770), .ZN(n26768) );
  INV_X1 U26738 ( .A(n26771), .ZN(n26769) );
  AND2_X1 U26739 ( .A1(n26772), .A2(n26771), .ZN(n26767) );
  INV_X1 U26740 ( .A(n26770), .ZN(n26772) );
  AND2_X1 U26741 ( .A1(n26773), .A2(n26774), .ZN(n26369) );
  INV_X1 U26742 ( .A(n26775), .ZN(n26774) );
  AND2_X1 U26743 ( .A1(n26776), .A2(n26777), .ZN(n26775) );
  OR2_X1 U26744 ( .A1(n26777), .A2(n26776), .ZN(n26773) );
  OR2_X1 U26745 ( .A1(n26778), .A2(n26779), .ZN(n26776) );
  AND2_X1 U26746 ( .A1(n26780), .A2(n26781), .ZN(n26779) );
  INV_X1 U26747 ( .A(n26782), .ZN(n26780) );
  AND2_X1 U26748 ( .A1(n26783), .A2(n26782), .ZN(n26778) );
  INV_X1 U26749 ( .A(n26781), .ZN(n26783) );
  AND2_X1 U26750 ( .A1(n26784), .A2(n26785), .ZN(n26380) );
  INV_X1 U26751 ( .A(n26786), .ZN(n26785) );
  AND2_X1 U26752 ( .A1(n26787), .A2(n26788), .ZN(n26786) );
  OR2_X1 U26753 ( .A1(n26788), .A2(n26787), .ZN(n26784) );
  OR2_X1 U26754 ( .A1(n26789), .A2(n26790), .ZN(n26787) );
  AND2_X1 U26755 ( .A1(n26791), .A2(n26792), .ZN(n26790) );
  INV_X1 U26756 ( .A(n26793), .ZN(n26791) );
  AND2_X1 U26757 ( .A1(n26794), .A2(n26793), .ZN(n26789) );
  INV_X1 U26758 ( .A(n26792), .ZN(n26794) );
  AND2_X1 U26759 ( .A1(n26795), .A2(n26796), .ZN(n26391) );
  INV_X1 U26760 ( .A(n26797), .ZN(n26796) );
  AND2_X1 U26761 ( .A1(n26798), .A2(n26799), .ZN(n26797) );
  OR2_X1 U26762 ( .A1(n26799), .A2(n26798), .ZN(n26795) );
  OR2_X1 U26763 ( .A1(n26800), .A2(n26801), .ZN(n26798) );
  AND2_X1 U26764 ( .A1(n26802), .A2(n26803), .ZN(n26801) );
  INV_X1 U26765 ( .A(n26804), .ZN(n26802) );
  AND2_X1 U26766 ( .A1(n26805), .A2(n26804), .ZN(n26800) );
  INV_X1 U26767 ( .A(n26803), .ZN(n26805) );
  AND2_X1 U26768 ( .A1(n26806), .A2(n26807), .ZN(n16456) );
  INV_X1 U26769 ( .A(n26808), .ZN(n26807) );
  AND2_X1 U26770 ( .A1(n26809), .A2(n26810), .ZN(n26808) );
  OR2_X1 U26771 ( .A1(n26810), .A2(n26809), .ZN(n26806) );
  OR2_X1 U26772 ( .A1(n26811), .A2(n26812), .ZN(n26809) );
  AND2_X1 U26773 ( .A1(n26813), .A2(n26814), .ZN(n26812) );
  INV_X1 U26774 ( .A(n26815), .ZN(n26813) );
  AND2_X1 U26775 ( .A1(n26816), .A2(n26815), .ZN(n26811) );
  INV_X1 U26776 ( .A(n26814), .ZN(n26816) );
  OR2_X1 U26777 ( .A1(n16446), .A2(n16447), .ZN(n14783) );
  OR2_X1 U26778 ( .A1(n26817), .A2(n26818), .ZN(n16447) );
  AND2_X1 U26779 ( .A1(n16467), .A2(n16466), .ZN(n26818) );
  AND2_X1 U26780 ( .A1(n16462), .A2(n26819), .ZN(n26817) );
  OR2_X1 U26781 ( .A1(n16466), .A2(n16467), .ZN(n26819) );
  OR2_X1 U26782 ( .A1(n16512), .A2(n15637), .ZN(n16467) );
  OR2_X1 U26783 ( .A1(n26820), .A2(n26821), .ZN(n16466) );
  AND2_X1 U26784 ( .A1(n26815), .A2(n26814), .ZN(n26821) );
  AND2_X1 U26785 ( .A1(n26810), .A2(n26822), .ZN(n26820) );
  OR2_X1 U26786 ( .A1(n26814), .A2(n26815), .ZN(n26822) );
  OR2_X1 U26787 ( .A1(n15842), .A2(n15637), .ZN(n26815) );
  OR2_X1 U26788 ( .A1(n26823), .A2(n26824), .ZN(n26814) );
  AND2_X1 U26789 ( .A1(n26804), .A2(n26803), .ZN(n26824) );
  AND2_X1 U26790 ( .A1(n26799), .A2(n26825), .ZN(n26823) );
  OR2_X1 U26791 ( .A1(n26803), .A2(n26804), .ZN(n26825) );
  OR2_X1 U26792 ( .A1(n15808), .A2(n15637), .ZN(n26804) );
  OR2_X1 U26793 ( .A1(n26826), .A2(n26827), .ZN(n26803) );
  AND2_X1 U26794 ( .A1(n26793), .A2(n26792), .ZN(n26827) );
  AND2_X1 U26795 ( .A1(n26788), .A2(n26828), .ZN(n26826) );
  OR2_X1 U26796 ( .A1(n26792), .A2(n26793), .ZN(n26828) );
  OR2_X1 U26797 ( .A1(n15774), .A2(n15637), .ZN(n26793) );
  OR2_X1 U26798 ( .A1(n26829), .A2(n26830), .ZN(n26792) );
  AND2_X1 U26799 ( .A1(n26782), .A2(n26781), .ZN(n26830) );
  AND2_X1 U26800 ( .A1(n26777), .A2(n26831), .ZN(n26829) );
  OR2_X1 U26801 ( .A1(n26781), .A2(n26782), .ZN(n26831) );
  OR2_X1 U26802 ( .A1(n15740), .A2(n15637), .ZN(n26782) );
  OR2_X1 U26803 ( .A1(n26832), .A2(n26833), .ZN(n26781) );
  AND2_X1 U26804 ( .A1(n26771), .A2(n26770), .ZN(n26833) );
  AND2_X1 U26805 ( .A1(n26766), .A2(n26834), .ZN(n26832) );
  OR2_X1 U26806 ( .A1(n26770), .A2(n26771), .ZN(n26834) );
  OR2_X1 U26807 ( .A1(n15706), .A2(n15637), .ZN(n26771) );
  OR2_X1 U26808 ( .A1(n26835), .A2(n26836), .ZN(n26770) );
  AND2_X1 U26809 ( .A1(n26760), .A2(n26759), .ZN(n26836) );
  AND2_X1 U26810 ( .A1(n26755), .A2(n26837), .ZN(n26835) );
  OR2_X1 U26811 ( .A1(n26759), .A2(n26760), .ZN(n26837) );
  OR2_X1 U26812 ( .A1(n15672), .A2(n15637), .ZN(n26760) );
  OR2_X1 U26813 ( .A1(n26838), .A2(n26839), .ZN(n26759) );
  AND2_X1 U26814 ( .A1(n15888), .A2(n26749), .ZN(n26839) );
  AND2_X1 U26815 ( .A1(n26745), .A2(n26840), .ZN(n26838) );
  OR2_X1 U26816 ( .A1(n26749), .A2(n15888), .ZN(n26840) );
  OR2_X1 U26817 ( .A1(n15638), .A2(n15637), .ZN(n15888) );
  OR2_X1 U26818 ( .A1(n26841), .A2(n26842), .ZN(n26749) );
  AND2_X1 U26819 ( .A1(n26739), .A2(n26738), .ZN(n26842) );
  AND2_X1 U26820 ( .A1(n26734), .A2(n26843), .ZN(n26841) );
  OR2_X1 U26821 ( .A1(n26738), .A2(n26739), .ZN(n26843) );
  OR2_X1 U26822 ( .A1(n15593), .A2(n15637), .ZN(n26739) );
  OR2_X1 U26823 ( .A1(n26844), .A2(n26845), .ZN(n26738) );
  AND2_X1 U26824 ( .A1(n26728), .A2(n26727), .ZN(n26845) );
  AND2_X1 U26825 ( .A1(n26723), .A2(n26846), .ZN(n26844) );
  OR2_X1 U26826 ( .A1(n26727), .A2(n26728), .ZN(n26846) );
  OR2_X1 U26827 ( .A1(n15559), .A2(n15637), .ZN(n26728) );
  OR2_X1 U26828 ( .A1(n26847), .A2(n26848), .ZN(n26727) );
  AND2_X1 U26829 ( .A1(n26717), .A2(n26716), .ZN(n26848) );
  AND2_X1 U26830 ( .A1(n26712), .A2(n26849), .ZN(n26847) );
  OR2_X1 U26831 ( .A1(n26716), .A2(n26717), .ZN(n26849) );
  OR2_X1 U26832 ( .A1(n15525), .A2(n15637), .ZN(n26717) );
  OR2_X1 U26833 ( .A1(n26850), .A2(n26851), .ZN(n26716) );
  AND2_X1 U26834 ( .A1(n26706), .A2(n26705), .ZN(n26851) );
  AND2_X1 U26835 ( .A1(n26701), .A2(n26852), .ZN(n26850) );
  OR2_X1 U26836 ( .A1(n26705), .A2(n26706), .ZN(n26852) );
  OR2_X1 U26837 ( .A1(n15491), .A2(n15637), .ZN(n26706) );
  OR2_X1 U26838 ( .A1(n26853), .A2(n26854), .ZN(n26705) );
  AND2_X1 U26839 ( .A1(n26695), .A2(n26694), .ZN(n26854) );
  AND2_X1 U26840 ( .A1(n26690), .A2(n26855), .ZN(n26853) );
  OR2_X1 U26841 ( .A1(n26694), .A2(n26695), .ZN(n26855) );
  OR2_X1 U26842 ( .A1(n15457), .A2(n15637), .ZN(n26695) );
  OR2_X1 U26843 ( .A1(n26856), .A2(n26857), .ZN(n26694) );
  AND2_X1 U26844 ( .A1(n26684), .A2(n26683), .ZN(n26857) );
  AND2_X1 U26845 ( .A1(n26679), .A2(n26858), .ZN(n26856) );
  OR2_X1 U26846 ( .A1(n26683), .A2(n26684), .ZN(n26858) );
  OR2_X1 U26847 ( .A1(n15423), .A2(n15637), .ZN(n26684) );
  OR2_X1 U26848 ( .A1(n26859), .A2(n26860), .ZN(n26683) );
  AND2_X1 U26849 ( .A1(n26673), .A2(n26672), .ZN(n26860) );
  AND2_X1 U26850 ( .A1(n26668), .A2(n26861), .ZN(n26859) );
  OR2_X1 U26851 ( .A1(n26672), .A2(n26673), .ZN(n26861) );
  OR2_X1 U26852 ( .A1(n15389), .A2(n15637), .ZN(n26673) );
  OR2_X1 U26853 ( .A1(n26862), .A2(n26863), .ZN(n26672) );
  AND2_X1 U26854 ( .A1(n26662), .A2(n26661), .ZN(n26863) );
  AND2_X1 U26855 ( .A1(n26657), .A2(n26864), .ZN(n26862) );
  OR2_X1 U26856 ( .A1(n26661), .A2(n26662), .ZN(n26864) );
  OR2_X1 U26857 ( .A1(n15355), .A2(n15637), .ZN(n26662) );
  OR2_X1 U26858 ( .A1(n26865), .A2(n26866), .ZN(n26661) );
  AND2_X1 U26859 ( .A1(n26651), .A2(n26650), .ZN(n26866) );
  AND2_X1 U26860 ( .A1(n26646), .A2(n26867), .ZN(n26865) );
  OR2_X1 U26861 ( .A1(n26650), .A2(n26651), .ZN(n26867) );
  OR2_X1 U26862 ( .A1(n15321), .A2(n15637), .ZN(n26651) );
  OR2_X1 U26863 ( .A1(n26868), .A2(n26869), .ZN(n26650) );
  AND2_X1 U26864 ( .A1(n26640), .A2(n26639), .ZN(n26869) );
  AND2_X1 U26865 ( .A1(n26635), .A2(n26870), .ZN(n26868) );
  OR2_X1 U26866 ( .A1(n26639), .A2(n26640), .ZN(n26870) );
  OR2_X1 U26867 ( .A1(n15287), .A2(n15637), .ZN(n26640) );
  OR2_X1 U26868 ( .A1(n26871), .A2(n26872), .ZN(n26639) );
  AND2_X1 U26869 ( .A1(n26629), .A2(n26628), .ZN(n26872) );
  AND2_X1 U26870 ( .A1(n26624), .A2(n26873), .ZN(n26871) );
  OR2_X1 U26871 ( .A1(n26628), .A2(n26629), .ZN(n26873) );
  OR2_X1 U26872 ( .A1(n15242), .A2(n15637), .ZN(n26629) );
  OR2_X1 U26873 ( .A1(n26874), .A2(n26875), .ZN(n26628) );
  AND2_X1 U26874 ( .A1(n26618), .A2(n26617), .ZN(n26875) );
  AND2_X1 U26875 ( .A1(n26613), .A2(n26876), .ZN(n26874) );
  OR2_X1 U26876 ( .A1(n26617), .A2(n26618), .ZN(n26876) );
  OR2_X1 U26877 ( .A1(n15208), .A2(n15637), .ZN(n26618) );
  OR2_X1 U26878 ( .A1(n26877), .A2(n26878), .ZN(n26617) );
  AND2_X1 U26879 ( .A1(n26607), .A2(n26606), .ZN(n26878) );
  AND2_X1 U26880 ( .A1(n26602), .A2(n26879), .ZN(n26877) );
  OR2_X1 U26881 ( .A1(n26606), .A2(n26607), .ZN(n26879) );
  OR2_X1 U26882 ( .A1(n15174), .A2(n15637), .ZN(n26607) );
  OR2_X1 U26883 ( .A1(n26880), .A2(n26881), .ZN(n26606) );
  AND2_X1 U26884 ( .A1(n26596), .A2(n26595), .ZN(n26881) );
  AND2_X1 U26885 ( .A1(n26591), .A2(n26882), .ZN(n26880) );
  OR2_X1 U26886 ( .A1(n26595), .A2(n26596), .ZN(n26882) );
  OR2_X1 U26887 ( .A1(n15140), .A2(n15637), .ZN(n26596) );
  OR2_X1 U26888 ( .A1(n26883), .A2(n26884), .ZN(n26595) );
  AND2_X1 U26889 ( .A1(n26580), .A2(n26586), .ZN(n26884) );
  AND2_X1 U26890 ( .A1(n26885), .A2(n26585), .ZN(n26883) );
  OR2_X1 U26891 ( .A1(n26886), .A2(n26887), .ZN(n26585) );
  AND2_X1 U26892 ( .A1(n26572), .A2(n26574), .ZN(n26887) );
  AND2_X1 U26893 ( .A1(n26569), .A2(n26888), .ZN(n26886) );
  OR2_X1 U26894 ( .A1(n26574), .A2(n26572), .ZN(n26888) );
  OR2_X1 U26895 ( .A1(n15072), .A2(n15637), .ZN(n26572) );
  OR2_X1 U26896 ( .A1(n26889), .A2(n26890), .ZN(n26574) );
  AND2_X1 U26897 ( .A1(n26558), .A2(n26561), .ZN(n26890) );
  AND2_X1 U26898 ( .A1(n26891), .A2(n26563), .ZN(n26889) );
  OR2_X1 U26899 ( .A1(n26892), .A2(n26893), .ZN(n26563) );
  AND2_X1 U26900 ( .A1(n26547), .A2(n26550), .ZN(n26893) );
  AND2_X1 U26901 ( .A1(n26894), .A2(n26552), .ZN(n26892) );
  OR2_X1 U26902 ( .A1(n26895), .A2(n26896), .ZN(n26552) );
  AND2_X1 U26903 ( .A1(n26536), .A2(n26539), .ZN(n26896) );
  AND2_X1 U26904 ( .A1(n26897), .A2(n26541), .ZN(n26895) );
  OR2_X1 U26905 ( .A1(n26898), .A2(n26899), .ZN(n26541) );
  AND2_X1 U26906 ( .A1(n26525), .A2(n26528), .ZN(n26899) );
  AND2_X1 U26907 ( .A1(n26900), .A2(n26530), .ZN(n26898) );
  OR2_X1 U26908 ( .A1(n26901), .A2(n26902), .ZN(n26530) );
  AND2_X1 U26909 ( .A1(n26514), .A2(n26517), .ZN(n26902) );
  AND2_X1 U26910 ( .A1(n26903), .A2(n26519), .ZN(n26901) );
  OR2_X1 U26911 ( .A1(n26904), .A2(n26905), .ZN(n26519) );
  AND2_X1 U26912 ( .A1(n26502), .A2(n26507), .ZN(n26905) );
  AND2_X1 U26913 ( .A1(n26506), .A2(n26906), .ZN(n26904) );
  OR2_X1 U26914 ( .A1(n26507), .A2(n26502), .ZN(n26906) );
  OR2_X1 U26915 ( .A1(n14857), .A2(n15637), .ZN(n26502) );
  INV_X1 U26916 ( .A(n26508), .ZN(n26507) );
  AND3_X1 U26917 ( .A1(b_7_), .A2(b_6_), .A3(n15957), .ZN(n26508) );
  INV_X1 U26918 ( .A(n26509), .ZN(n26506) );
  OR2_X1 U26919 ( .A1(n26907), .A2(n26908), .ZN(n26509) );
  AND2_X1 U26920 ( .A1(b_6_), .A2(n26909), .ZN(n26908) );
  OR2_X1 U26921 ( .A1(n26910), .A2(n16981), .ZN(n26909) );
  AND2_X1 U26922 ( .A1(a_30_), .A2(n15705), .ZN(n26910) );
  AND2_X1 U26923 ( .A1(b_5_), .A2(n26911), .ZN(n26907) );
  OR2_X1 U26924 ( .A1(n26912), .A2(n14817), .ZN(n26911) );
  AND2_X1 U26925 ( .A1(a_31_), .A2(n15671), .ZN(n26912) );
  OR2_X1 U26926 ( .A1(n26517), .A2(n26514), .ZN(n26903) );
  OR2_X1 U26927 ( .A1(n26913), .A2(n26914), .ZN(n26514) );
  AND2_X1 U26928 ( .A1(n26915), .A2(n26916), .ZN(n26914) );
  INV_X1 U26929 ( .A(n26917), .ZN(n26913) );
  OR2_X1 U26930 ( .A1(n26915), .A2(n26916), .ZN(n26917) );
  OR2_X1 U26931 ( .A1(n26918), .A2(n26919), .ZN(n26915) );
  AND2_X1 U26932 ( .A1(n26920), .A2(n26921), .ZN(n26919) );
  AND2_X1 U26933 ( .A1(n26922), .A2(n26923), .ZN(n26918) );
  OR2_X1 U26934 ( .A1(n14891), .A2(n15637), .ZN(n26517) );
  OR2_X1 U26935 ( .A1(n26528), .A2(n26525), .ZN(n26900) );
  OR2_X1 U26936 ( .A1(n26924), .A2(n26925), .ZN(n26525) );
  INV_X1 U26937 ( .A(n26926), .ZN(n26925) );
  OR2_X1 U26938 ( .A1(n26927), .A2(n26928), .ZN(n26926) );
  AND2_X1 U26939 ( .A1(n26928), .A2(n26927), .ZN(n26924) );
  AND2_X1 U26940 ( .A1(n26929), .A2(n26930), .ZN(n26927) );
  OR2_X1 U26941 ( .A1(n26931), .A2(n26932), .ZN(n26930) );
  INV_X1 U26942 ( .A(n26933), .ZN(n26932) );
  OR2_X1 U26943 ( .A1(n26933), .A2(n26934), .ZN(n26929) );
  INV_X1 U26944 ( .A(n26931), .ZN(n26934) );
  OR2_X1 U26945 ( .A1(n14936), .A2(n15637), .ZN(n26528) );
  OR2_X1 U26946 ( .A1(n26539), .A2(n26536), .ZN(n26897) );
  OR2_X1 U26947 ( .A1(n26935), .A2(n26936), .ZN(n26536) );
  INV_X1 U26948 ( .A(n26937), .ZN(n26936) );
  OR2_X1 U26949 ( .A1(n26938), .A2(n26939), .ZN(n26937) );
  AND2_X1 U26950 ( .A1(n26939), .A2(n26938), .ZN(n26935) );
  AND2_X1 U26951 ( .A1(n26940), .A2(n26941), .ZN(n26938) );
  OR2_X1 U26952 ( .A1(n26942), .A2(n26943), .ZN(n26941) );
  INV_X1 U26953 ( .A(n26944), .ZN(n26943) );
  OR2_X1 U26954 ( .A1(n26944), .A2(n26945), .ZN(n26940) );
  INV_X1 U26955 ( .A(n26942), .ZN(n26945) );
  OR2_X1 U26956 ( .A1(n14970), .A2(n15637), .ZN(n26539) );
  OR2_X1 U26957 ( .A1(n26550), .A2(n26547), .ZN(n26894) );
  OR2_X1 U26958 ( .A1(n26946), .A2(n26947), .ZN(n26547) );
  INV_X1 U26959 ( .A(n26948), .ZN(n26947) );
  OR2_X1 U26960 ( .A1(n26949), .A2(n26950), .ZN(n26948) );
  AND2_X1 U26961 ( .A1(n26950), .A2(n26949), .ZN(n26946) );
  AND2_X1 U26962 ( .A1(n26951), .A2(n26952), .ZN(n26949) );
  OR2_X1 U26963 ( .A1(n26953), .A2(n26954), .ZN(n26952) );
  INV_X1 U26964 ( .A(n26955), .ZN(n26954) );
  OR2_X1 U26965 ( .A1(n26955), .A2(n26956), .ZN(n26951) );
  INV_X1 U26966 ( .A(n26953), .ZN(n26956) );
  OR2_X1 U26967 ( .A1(n15004), .A2(n15637), .ZN(n26550) );
  OR2_X1 U26968 ( .A1(n26561), .A2(n26558), .ZN(n26891) );
  OR2_X1 U26969 ( .A1(n26957), .A2(n26958), .ZN(n26558) );
  INV_X1 U26970 ( .A(n26959), .ZN(n26958) );
  OR2_X1 U26971 ( .A1(n26960), .A2(n26961), .ZN(n26959) );
  AND2_X1 U26972 ( .A1(n26961), .A2(n26960), .ZN(n26957) );
  AND2_X1 U26973 ( .A1(n26962), .A2(n26963), .ZN(n26960) );
  OR2_X1 U26974 ( .A1(n26964), .A2(n26965), .ZN(n26963) );
  INV_X1 U26975 ( .A(n26966), .ZN(n26965) );
  OR2_X1 U26976 ( .A1(n26966), .A2(n26967), .ZN(n26962) );
  INV_X1 U26977 ( .A(n26964), .ZN(n26967) );
  OR2_X1 U26978 ( .A1(n15038), .A2(n15637), .ZN(n26561) );
  OR2_X1 U26979 ( .A1(n26968), .A2(n26969), .ZN(n26569) );
  INV_X1 U26980 ( .A(n26970), .ZN(n26969) );
  OR2_X1 U26981 ( .A1(n26971), .A2(n26972), .ZN(n26970) );
  AND2_X1 U26982 ( .A1(n26972), .A2(n26971), .ZN(n26968) );
  AND2_X1 U26983 ( .A1(n26973), .A2(n26974), .ZN(n26971) );
  OR2_X1 U26984 ( .A1(n26975), .A2(n26976), .ZN(n26974) );
  INV_X1 U26985 ( .A(n26977), .ZN(n26976) );
  OR2_X1 U26986 ( .A1(n26977), .A2(n26978), .ZN(n26973) );
  INV_X1 U26987 ( .A(n26975), .ZN(n26978) );
  OR2_X1 U26988 ( .A1(n26586), .A2(n26580), .ZN(n26885) );
  OR2_X1 U26989 ( .A1(n26979), .A2(n26980), .ZN(n26580) );
  INV_X1 U26990 ( .A(n26981), .ZN(n26980) );
  OR2_X1 U26991 ( .A1(n26982), .A2(n26983), .ZN(n26981) );
  AND2_X1 U26992 ( .A1(n26983), .A2(n26982), .ZN(n26979) );
  AND2_X1 U26993 ( .A1(n26984), .A2(n26985), .ZN(n26982) );
  INV_X1 U26994 ( .A(n26986), .ZN(n26985) );
  AND2_X1 U26995 ( .A1(n26987), .A2(n26988), .ZN(n26986) );
  OR2_X1 U26996 ( .A1(n26988), .A2(n26987), .ZN(n26984) );
  INV_X1 U26997 ( .A(n26989), .ZN(n26987) );
  OR2_X1 U26998 ( .A1(n15106), .A2(n15637), .ZN(n26586) );
  INV_X1 U26999 ( .A(b_7_), .ZN(n15637) );
  AND2_X1 U27000 ( .A1(n26990), .A2(n26991), .ZN(n26591) );
  INV_X1 U27001 ( .A(n26992), .ZN(n26991) );
  AND2_X1 U27002 ( .A1(n26993), .A2(n26994), .ZN(n26992) );
  OR2_X1 U27003 ( .A1(n26994), .A2(n26993), .ZN(n26990) );
  OR2_X1 U27004 ( .A1(n26995), .A2(n26996), .ZN(n26993) );
  AND2_X1 U27005 ( .A1(n26997), .A2(n26998), .ZN(n26996) );
  INV_X1 U27006 ( .A(n26999), .ZN(n26997) );
  AND2_X1 U27007 ( .A1(n27000), .A2(n26999), .ZN(n26995) );
  INV_X1 U27008 ( .A(n26998), .ZN(n27000) );
  AND2_X1 U27009 ( .A1(n27001), .A2(n27002), .ZN(n26602) );
  INV_X1 U27010 ( .A(n27003), .ZN(n27002) );
  AND2_X1 U27011 ( .A1(n27004), .A2(n27005), .ZN(n27003) );
  OR2_X1 U27012 ( .A1(n27005), .A2(n27004), .ZN(n27001) );
  OR2_X1 U27013 ( .A1(n27006), .A2(n27007), .ZN(n27004) );
  AND2_X1 U27014 ( .A1(n27008), .A2(n27009), .ZN(n27007) );
  INV_X1 U27015 ( .A(n27010), .ZN(n27008) );
  AND2_X1 U27016 ( .A1(n27011), .A2(n27010), .ZN(n27006) );
  INV_X1 U27017 ( .A(n27009), .ZN(n27011) );
  AND2_X1 U27018 ( .A1(n27012), .A2(n27013), .ZN(n26613) );
  INV_X1 U27019 ( .A(n27014), .ZN(n27013) );
  AND2_X1 U27020 ( .A1(n27015), .A2(n27016), .ZN(n27014) );
  OR2_X1 U27021 ( .A1(n27016), .A2(n27015), .ZN(n27012) );
  OR2_X1 U27022 ( .A1(n27017), .A2(n27018), .ZN(n27015) );
  AND2_X1 U27023 ( .A1(n27019), .A2(n27020), .ZN(n27018) );
  INV_X1 U27024 ( .A(n27021), .ZN(n27019) );
  AND2_X1 U27025 ( .A1(n27022), .A2(n27021), .ZN(n27017) );
  INV_X1 U27026 ( .A(n27020), .ZN(n27022) );
  AND2_X1 U27027 ( .A1(n27023), .A2(n27024), .ZN(n26624) );
  INV_X1 U27028 ( .A(n27025), .ZN(n27024) );
  AND2_X1 U27029 ( .A1(n27026), .A2(n27027), .ZN(n27025) );
  OR2_X1 U27030 ( .A1(n27027), .A2(n27026), .ZN(n27023) );
  OR2_X1 U27031 ( .A1(n27028), .A2(n27029), .ZN(n27026) );
  AND2_X1 U27032 ( .A1(n27030), .A2(n27031), .ZN(n27029) );
  INV_X1 U27033 ( .A(n27032), .ZN(n27030) );
  AND2_X1 U27034 ( .A1(n27033), .A2(n27032), .ZN(n27028) );
  INV_X1 U27035 ( .A(n27031), .ZN(n27033) );
  AND2_X1 U27036 ( .A1(n27034), .A2(n27035), .ZN(n26635) );
  INV_X1 U27037 ( .A(n27036), .ZN(n27035) );
  AND2_X1 U27038 ( .A1(n27037), .A2(n27038), .ZN(n27036) );
  OR2_X1 U27039 ( .A1(n27038), .A2(n27037), .ZN(n27034) );
  OR2_X1 U27040 ( .A1(n27039), .A2(n27040), .ZN(n27037) );
  AND2_X1 U27041 ( .A1(n27041), .A2(n27042), .ZN(n27040) );
  INV_X1 U27042 ( .A(n27043), .ZN(n27041) );
  AND2_X1 U27043 ( .A1(n27044), .A2(n27043), .ZN(n27039) );
  INV_X1 U27044 ( .A(n27042), .ZN(n27044) );
  AND2_X1 U27045 ( .A1(n27045), .A2(n27046), .ZN(n26646) );
  INV_X1 U27046 ( .A(n27047), .ZN(n27046) );
  AND2_X1 U27047 ( .A1(n27048), .A2(n27049), .ZN(n27047) );
  OR2_X1 U27048 ( .A1(n27049), .A2(n27048), .ZN(n27045) );
  OR2_X1 U27049 ( .A1(n27050), .A2(n27051), .ZN(n27048) );
  AND2_X1 U27050 ( .A1(n27052), .A2(n27053), .ZN(n27051) );
  INV_X1 U27051 ( .A(n27054), .ZN(n27052) );
  AND2_X1 U27052 ( .A1(n27055), .A2(n27054), .ZN(n27050) );
  INV_X1 U27053 ( .A(n27053), .ZN(n27055) );
  AND2_X1 U27054 ( .A1(n27056), .A2(n27057), .ZN(n26657) );
  INV_X1 U27055 ( .A(n27058), .ZN(n27057) );
  AND2_X1 U27056 ( .A1(n27059), .A2(n27060), .ZN(n27058) );
  OR2_X1 U27057 ( .A1(n27060), .A2(n27059), .ZN(n27056) );
  OR2_X1 U27058 ( .A1(n27061), .A2(n27062), .ZN(n27059) );
  AND2_X1 U27059 ( .A1(n27063), .A2(n27064), .ZN(n27062) );
  INV_X1 U27060 ( .A(n27065), .ZN(n27063) );
  AND2_X1 U27061 ( .A1(n27066), .A2(n27065), .ZN(n27061) );
  INV_X1 U27062 ( .A(n27064), .ZN(n27066) );
  AND2_X1 U27063 ( .A1(n27067), .A2(n27068), .ZN(n26668) );
  INV_X1 U27064 ( .A(n27069), .ZN(n27068) );
  AND2_X1 U27065 ( .A1(n27070), .A2(n27071), .ZN(n27069) );
  OR2_X1 U27066 ( .A1(n27071), .A2(n27070), .ZN(n27067) );
  OR2_X1 U27067 ( .A1(n27072), .A2(n27073), .ZN(n27070) );
  AND2_X1 U27068 ( .A1(n27074), .A2(n27075), .ZN(n27073) );
  INV_X1 U27069 ( .A(n27076), .ZN(n27074) );
  AND2_X1 U27070 ( .A1(n27077), .A2(n27076), .ZN(n27072) );
  INV_X1 U27071 ( .A(n27075), .ZN(n27077) );
  AND2_X1 U27072 ( .A1(n27078), .A2(n27079), .ZN(n26679) );
  INV_X1 U27073 ( .A(n27080), .ZN(n27079) );
  AND2_X1 U27074 ( .A1(n27081), .A2(n27082), .ZN(n27080) );
  OR2_X1 U27075 ( .A1(n27082), .A2(n27081), .ZN(n27078) );
  OR2_X1 U27076 ( .A1(n27083), .A2(n27084), .ZN(n27081) );
  AND2_X1 U27077 ( .A1(n27085), .A2(n27086), .ZN(n27084) );
  INV_X1 U27078 ( .A(n27087), .ZN(n27085) );
  AND2_X1 U27079 ( .A1(n27088), .A2(n27087), .ZN(n27083) );
  INV_X1 U27080 ( .A(n27086), .ZN(n27088) );
  AND2_X1 U27081 ( .A1(n27089), .A2(n27090), .ZN(n26690) );
  INV_X1 U27082 ( .A(n27091), .ZN(n27090) );
  AND2_X1 U27083 ( .A1(n27092), .A2(n27093), .ZN(n27091) );
  OR2_X1 U27084 ( .A1(n27093), .A2(n27092), .ZN(n27089) );
  OR2_X1 U27085 ( .A1(n27094), .A2(n27095), .ZN(n27092) );
  AND2_X1 U27086 ( .A1(n27096), .A2(n27097), .ZN(n27095) );
  INV_X1 U27087 ( .A(n27098), .ZN(n27096) );
  AND2_X1 U27088 ( .A1(n27099), .A2(n27098), .ZN(n27094) );
  INV_X1 U27089 ( .A(n27097), .ZN(n27099) );
  AND2_X1 U27090 ( .A1(n27100), .A2(n27101), .ZN(n26701) );
  INV_X1 U27091 ( .A(n27102), .ZN(n27101) );
  AND2_X1 U27092 ( .A1(n27103), .A2(n27104), .ZN(n27102) );
  OR2_X1 U27093 ( .A1(n27104), .A2(n27103), .ZN(n27100) );
  OR2_X1 U27094 ( .A1(n27105), .A2(n27106), .ZN(n27103) );
  AND2_X1 U27095 ( .A1(n27107), .A2(n27108), .ZN(n27106) );
  INV_X1 U27096 ( .A(n27109), .ZN(n27107) );
  AND2_X1 U27097 ( .A1(n27110), .A2(n27109), .ZN(n27105) );
  INV_X1 U27098 ( .A(n27108), .ZN(n27110) );
  AND2_X1 U27099 ( .A1(n27111), .A2(n27112), .ZN(n26712) );
  INV_X1 U27100 ( .A(n27113), .ZN(n27112) );
  AND2_X1 U27101 ( .A1(n27114), .A2(n27115), .ZN(n27113) );
  OR2_X1 U27102 ( .A1(n27115), .A2(n27114), .ZN(n27111) );
  OR2_X1 U27103 ( .A1(n27116), .A2(n27117), .ZN(n27114) );
  AND2_X1 U27104 ( .A1(n27118), .A2(n27119), .ZN(n27117) );
  INV_X1 U27105 ( .A(n27120), .ZN(n27118) );
  AND2_X1 U27106 ( .A1(n27121), .A2(n27120), .ZN(n27116) );
  INV_X1 U27107 ( .A(n27119), .ZN(n27121) );
  AND2_X1 U27108 ( .A1(n27122), .A2(n27123), .ZN(n26723) );
  INV_X1 U27109 ( .A(n27124), .ZN(n27123) );
  AND2_X1 U27110 ( .A1(n27125), .A2(n27126), .ZN(n27124) );
  OR2_X1 U27111 ( .A1(n27126), .A2(n27125), .ZN(n27122) );
  OR2_X1 U27112 ( .A1(n27127), .A2(n27128), .ZN(n27125) );
  AND2_X1 U27113 ( .A1(n27129), .A2(n27130), .ZN(n27128) );
  INV_X1 U27114 ( .A(n27131), .ZN(n27129) );
  AND2_X1 U27115 ( .A1(n27132), .A2(n27131), .ZN(n27127) );
  INV_X1 U27116 ( .A(n27130), .ZN(n27132) );
  AND2_X1 U27117 ( .A1(n27133), .A2(n27134), .ZN(n26734) );
  INV_X1 U27118 ( .A(n27135), .ZN(n27134) );
  AND2_X1 U27119 ( .A1(n27136), .A2(n27137), .ZN(n27135) );
  OR2_X1 U27120 ( .A1(n27137), .A2(n27136), .ZN(n27133) );
  OR2_X1 U27121 ( .A1(n27138), .A2(n27139), .ZN(n27136) );
  AND2_X1 U27122 ( .A1(n27140), .A2(n27141), .ZN(n27139) );
  INV_X1 U27123 ( .A(n27142), .ZN(n27140) );
  AND2_X1 U27124 ( .A1(n27143), .A2(n27142), .ZN(n27138) );
  INV_X1 U27125 ( .A(n27141), .ZN(n27143) );
  AND2_X1 U27126 ( .A1(n27144), .A2(n27145), .ZN(n26745) );
  INV_X1 U27127 ( .A(n27146), .ZN(n27145) );
  AND2_X1 U27128 ( .A1(n27147), .A2(n27148), .ZN(n27146) );
  OR2_X1 U27129 ( .A1(n27148), .A2(n27147), .ZN(n27144) );
  OR2_X1 U27130 ( .A1(n27149), .A2(n27150), .ZN(n27147) );
  AND2_X1 U27131 ( .A1(n27151), .A2(n27152), .ZN(n27150) );
  INV_X1 U27132 ( .A(n27153), .ZN(n27151) );
  AND2_X1 U27133 ( .A1(n27154), .A2(n27153), .ZN(n27149) );
  INV_X1 U27134 ( .A(n27152), .ZN(n27154) );
  AND2_X1 U27135 ( .A1(n27155), .A2(n27156), .ZN(n26755) );
  INV_X1 U27136 ( .A(n27157), .ZN(n27156) );
  AND2_X1 U27137 ( .A1(n27158), .A2(n27159), .ZN(n27157) );
  OR2_X1 U27138 ( .A1(n27159), .A2(n27158), .ZN(n27155) );
  OR2_X1 U27139 ( .A1(n27160), .A2(n27161), .ZN(n27158) );
  AND2_X1 U27140 ( .A1(n27162), .A2(n27163), .ZN(n27161) );
  INV_X1 U27141 ( .A(n27164), .ZN(n27162) );
  AND2_X1 U27142 ( .A1(n27165), .A2(n27164), .ZN(n27160) );
  INV_X1 U27143 ( .A(n27163), .ZN(n27165) );
  AND2_X1 U27144 ( .A1(n27166), .A2(n27167), .ZN(n26766) );
  INV_X1 U27145 ( .A(n27168), .ZN(n27167) );
  AND2_X1 U27146 ( .A1(n27169), .A2(n27170), .ZN(n27168) );
  OR2_X1 U27147 ( .A1(n27170), .A2(n27169), .ZN(n27166) );
  OR2_X1 U27148 ( .A1(n27171), .A2(n27172), .ZN(n27169) );
  AND2_X1 U27149 ( .A1(n27173), .A2(n27174), .ZN(n27172) );
  INV_X1 U27150 ( .A(n15885), .ZN(n27173) );
  AND2_X1 U27151 ( .A1(n27175), .A2(n15885), .ZN(n27171) );
  INV_X1 U27152 ( .A(n27174), .ZN(n27175) );
  AND2_X1 U27153 ( .A1(n27176), .A2(n27177), .ZN(n26777) );
  INV_X1 U27154 ( .A(n27178), .ZN(n27177) );
  AND2_X1 U27155 ( .A1(n27179), .A2(n27180), .ZN(n27178) );
  OR2_X1 U27156 ( .A1(n27180), .A2(n27179), .ZN(n27176) );
  OR2_X1 U27157 ( .A1(n27181), .A2(n27182), .ZN(n27179) );
  AND2_X1 U27158 ( .A1(n27183), .A2(n27184), .ZN(n27182) );
  INV_X1 U27159 ( .A(n27185), .ZN(n27183) );
  AND2_X1 U27160 ( .A1(n27186), .A2(n27185), .ZN(n27181) );
  INV_X1 U27161 ( .A(n27184), .ZN(n27186) );
  AND2_X1 U27162 ( .A1(n27187), .A2(n27188), .ZN(n26788) );
  INV_X1 U27163 ( .A(n27189), .ZN(n27188) );
  AND2_X1 U27164 ( .A1(n27190), .A2(n27191), .ZN(n27189) );
  OR2_X1 U27165 ( .A1(n27191), .A2(n27190), .ZN(n27187) );
  OR2_X1 U27166 ( .A1(n27192), .A2(n27193), .ZN(n27190) );
  AND2_X1 U27167 ( .A1(n27194), .A2(n27195), .ZN(n27193) );
  INV_X1 U27168 ( .A(n27196), .ZN(n27194) );
  AND2_X1 U27169 ( .A1(n27197), .A2(n27196), .ZN(n27192) );
  INV_X1 U27170 ( .A(n27195), .ZN(n27197) );
  AND2_X1 U27171 ( .A1(n27198), .A2(n27199), .ZN(n26799) );
  INV_X1 U27172 ( .A(n27200), .ZN(n27199) );
  AND2_X1 U27173 ( .A1(n27201), .A2(n27202), .ZN(n27200) );
  OR2_X1 U27174 ( .A1(n27202), .A2(n27201), .ZN(n27198) );
  OR2_X1 U27175 ( .A1(n27203), .A2(n27204), .ZN(n27201) );
  AND2_X1 U27176 ( .A1(n27205), .A2(n27206), .ZN(n27204) );
  INV_X1 U27177 ( .A(n27207), .ZN(n27205) );
  AND2_X1 U27178 ( .A1(n27208), .A2(n27207), .ZN(n27203) );
  INV_X1 U27179 ( .A(n27206), .ZN(n27208) );
  AND2_X1 U27180 ( .A1(n27209), .A2(n27210), .ZN(n26810) );
  INV_X1 U27181 ( .A(n27211), .ZN(n27210) );
  AND2_X1 U27182 ( .A1(n27212), .A2(n27213), .ZN(n27211) );
  OR2_X1 U27183 ( .A1(n27213), .A2(n27212), .ZN(n27209) );
  OR2_X1 U27184 ( .A1(n27214), .A2(n27215), .ZN(n27212) );
  AND2_X1 U27185 ( .A1(n27216), .A2(n27217), .ZN(n27215) );
  INV_X1 U27186 ( .A(n27218), .ZN(n27216) );
  AND2_X1 U27187 ( .A1(n27219), .A2(n27218), .ZN(n27214) );
  INV_X1 U27188 ( .A(n27217), .ZN(n27219) );
  AND2_X1 U27189 ( .A1(n27220), .A2(n27221), .ZN(n16462) );
  INV_X1 U27190 ( .A(n27222), .ZN(n27221) );
  AND2_X1 U27191 ( .A1(n27223), .A2(n27224), .ZN(n27222) );
  OR2_X1 U27192 ( .A1(n27224), .A2(n27223), .ZN(n27220) );
  OR2_X1 U27193 ( .A1(n27225), .A2(n27226), .ZN(n27223) );
  AND2_X1 U27194 ( .A1(n27227), .A2(n27228), .ZN(n27226) );
  INV_X1 U27195 ( .A(n27229), .ZN(n27227) );
  AND2_X1 U27196 ( .A1(n27230), .A2(n27229), .ZN(n27225) );
  INV_X1 U27197 ( .A(n27228), .ZN(n27230) );
  AND2_X1 U27198 ( .A1(n27231), .A2(n27232), .ZN(n16446) );
  INV_X1 U27199 ( .A(n27233), .ZN(n27232) );
  AND2_X1 U27200 ( .A1(n27234), .A2(n16431), .ZN(n27233) );
  OR2_X1 U27201 ( .A1(n16431), .A2(n27234), .ZN(n27231) );
  OR2_X1 U27202 ( .A1(n27235), .A2(n27236), .ZN(n27234) );
  AND2_X1 U27203 ( .A1(n27237), .A2(n16430), .ZN(n27236) );
  INV_X1 U27204 ( .A(n16429), .ZN(n27237) );
  AND2_X1 U27205 ( .A1(n27238), .A2(n16429), .ZN(n27235) );
  OR2_X1 U27206 ( .A1(n16512), .A2(n15671), .ZN(n16429) );
  INV_X1 U27207 ( .A(n16430), .ZN(n27238) );
  OR2_X1 U27208 ( .A1(n27239), .A2(n27240), .ZN(n16430) );
  AND2_X1 U27209 ( .A1(n27229), .A2(n27228), .ZN(n27240) );
  AND2_X1 U27210 ( .A1(n27224), .A2(n27241), .ZN(n27239) );
  OR2_X1 U27211 ( .A1(n27228), .A2(n27229), .ZN(n27241) );
  OR2_X1 U27212 ( .A1(n15842), .A2(n15671), .ZN(n27229) );
  OR2_X1 U27213 ( .A1(n27242), .A2(n27243), .ZN(n27228) );
  AND2_X1 U27214 ( .A1(n27218), .A2(n27217), .ZN(n27243) );
  AND2_X1 U27215 ( .A1(n27213), .A2(n27244), .ZN(n27242) );
  OR2_X1 U27216 ( .A1(n27217), .A2(n27218), .ZN(n27244) );
  OR2_X1 U27217 ( .A1(n15808), .A2(n15671), .ZN(n27218) );
  OR2_X1 U27218 ( .A1(n27245), .A2(n27246), .ZN(n27217) );
  AND2_X1 U27219 ( .A1(n27207), .A2(n27206), .ZN(n27246) );
  AND2_X1 U27220 ( .A1(n27202), .A2(n27247), .ZN(n27245) );
  OR2_X1 U27221 ( .A1(n27206), .A2(n27207), .ZN(n27247) );
  OR2_X1 U27222 ( .A1(n15774), .A2(n15671), .ZN(n27207) );
  OR2_X1 U27223 ( .A1(n27248), .A2(n27249), .ZN(n27206) );
  AND2_X1 U27224 ( .A1(n27196), .A2(n27195), .ZN(n27249) );
  AND2_X1 U27225 ( .A1(n27191), .A2(n27250), .ZN(n27248) );
  OR2_X1 U27226 ( .A1(n27195), .A2(n27196), .ZN(n27250) );
  OR2_X1 U27227 ( .A1(n15740), .A2(n15671), .ZN(n27196) );
  OR2_X1 U27228 ( .A1(n27251), .A2(n27252), .ZN(n27195) );
  AND2_X1 U27229 ( .A1(n27185), .A2(n27184), .ZN(n27252) );
  AND2_X1 U27230 ( .A1(n27180), .A2(n27253), .ZN(n27251) );
  OR2_X1 U27231 ( .A1(n27184), .A2(n27185), .ZN(n27253) );
  OR2_X1 U27232 ( .A1(n15706), .A2(n15671), .ZN(n27185) );
  OR2_X1 U27233 ( .A1(n27254), .A2(n27255), .ZN(n27184) );
  AND2_X1 U27234 ( .A1(n15885), .A2(n27174), .ZN(n27255) );
  AND2_X1 U27235 ( .A1(n27170), .A2(n27256), .ZN(n27254) );
  OR2_X1 U27236 ( .A1(n27174), .A2(n15885), .ZN(n27256) );
  OR2_X1 U27237 ( .A1(n15672), .A2(n15671), .ZN(n15885) );
  OR2_X1 U27238 ( .A1(n27257), .A2(n27258), .ZN(n27174) );
  AND2_X1 U27239 ( .A1(n27164), .A2(n27163), .ZN(n27258) );
  AND2_X1 U27240 ( .A1(n27159), .A2(n27259), .ZN(n27257) );
  OR2_X1 U27241 ( .A1(n27163), .A2(n27164), .ZN(n27259) );
  OR2_X1 U27242 ( .A1(n15638), .A2(n15671), .ZN(n27164) );
  OR2_X1 U27243 ( .A1(n27260), .A2(n27261), .ZN(n27163) );
  AND2_X1 U27244 ( .A1(n27153), .A2(n27152), .ZN(n27261) );
  AND2_X1 U27245 ( .A1(n27148), .A2(n27262), .ZN(n27260) );
  OR2_X1 U27246 ( .A1(n27152), .A2(n27153), .ZN(n27262) );
  OR2_X1 U27247 ( .A1(n15593), .A2(n15671), .ZN(n27153) );
  OR2_X1 U27248 ( .A1(n27263), .A2(n27264), .ZN(n27152) );
  AND2_X1 U27249 ( .A1(n27142), .A2(n27141), .ZN(n27264) );
  AND2_X1 U27250 ( .A1(n27137), .A2(n27265), .ZN(n27263) );
  OR2_X1 U27251 ( .A1(n27141), .A2(n27142), .ZN(n27265) );
  OR2_X1 U27252 ( .A1(n15559), .A2(n15671), .ZN(n27142) );
  OR2_X1 U27253 ( .A1(n27266), .A2(n27267), .ZN(n27141) );
  AND2_X1 U27254 ( .A1(n27131), .A2(n27130), .ZN(n27267) );
  AND2_X1 U27255 ( .A1(n27126), .A2(n27268), .ZN(n27266) );
  OR2_X1 U27256 ( .A1(n27130), .A2(n27131), .ZN(n27268) );
  OR2_X1 U27257 ( .A1(n15525), .A2(n15671), .ZN(n27131) );
  OR2_X1 U27258 ( .A1(n27269), .A2(n27270), .ZN(n27130) );
  AND2_X1 U27259 ( .A1(n27120), .A2(n27119), .ZN(n27270) );
  AND2_X1 U27260 ( .A1(n27115), .A2(n27271), .ZN(n27269) );
  OR2_X1 U27261 ( .A1(n27119), .A2(n27120), .ZN(n27271) );
  OR2_X1 U27262 ( .A1(n15491), .A2(n15671), .ZN(n27120) );
  OR2_X1 U27263 ( .A1(n27272), .A2(n27273), .ZN(n27119) );
  AND2_X1 U27264 ( .A1(n27109), .A2(n27108), .ZN(n27273) );
  AND2_X1 U27265 ( .A1(n27104), .A2(n27274), .ZN(n27272) );
  OR2_X1 U27266 ( .A1(n27108), .A2(n27109), .ZN(n27274) );
  OR2_X1 U27267 ( .A1(n15457), .A2(n15671), .ZN(n27109) );
  OR2_X1 U27268 ( .A1(n27275), .A2(n27276), .ZN(n27108) );
  AND2_X1 U27269 ( .A1(n27098), .A2(n27097), .ZN(n27276) );
  AND2_X1 U27270 ( .A1(n27093), .A2(n27277), .ZN(n27275) );
  OR2_X1 U27271 ( .A1(n27097), .A2(n27098), .ZN(n27277) );
  OR2_X1 U27272 ( .A1(n15423), .A2(n15671), .ZN(n27098) );
  OR2_X1 U27273 ( .A1(n27278), .A2(n27279), .ZN(n27097) );
  AND2_X1 U27274 ( .A1(n27087), .A2(n27086), .ZN(n27279) );
  AND2_X1 U27275 ( .A1(n27082), .A2(n27280), .ZN(n27278) );
  OR2_X1 U27276 ( .A1(n27086), .A2(n27087), .ZN(n27280) );
  OR2_X1 U27277 ( .A1(n15389), .A2(n15671), .ZN(n27087) );
  OR2_X1 U27278 ( .A1(n27281), .A2(n27282), .ZN(n27086) );
  AND2_X1 U27279 ( .A1(n27076), .A2(n27075), .ZN(n27282) );
  AND2_X1 U27280 ( .A1(n27071), .A2(n27283), .ZN(n27281) );
  OR2_X1 U27281 ( .A1(n27075), .A2(n27076), .ZN(n27283) );
  OR2_X1 U27282 ( .A1(n15355), .A2(n15671), .ZN(n27076) );
  OR2_X1 U27283 ( .A1(n27284), .A2(n27285), .ZN(n27075) );
  AND2_X1 U27284 ( .A1(n27065), .A2(n27064), .ZN(n27285) );
  AND2_X1 U27285 ( .A1(n27060), .A2(n27286), .ZN(n27284) );
  OR2_X1 U27286 ( .A1(n27064), .A2(n27065), .ZN(n27286) );
  OR2_X1 U27287 ( .A1(n15321), .A2(n15671), .ZN(n27065) );
  OR2_X1 U27288 ( .A1(n27287), .A2(n27288), .ZN(n27064) );
  AND2_X1 U27289 ( .A1(n27054), .A2(n27053), .ZN(n27288) );
  AND2_X1 U27290 ( .A1(n27049), .A2(n27289), .ZN(n27287) );
  OR2_X1 U27291 ( .A1(n27053), .A2(n27054), .ZN(n27289) );
  OR2_X1 U27292 ( .A1(n15287), .A2(n15671), .ZN(n27054) );
  OR2_X1 U27293 ( .A1(n27290), .A2(n27291), .ZN(n27053) );
  AND2_X1 U27294 ( .A1(n27043), .A2(n27042), .ZN(n27291) );
  AND2_X1 U27295 ( .A1(n27038), .A2(n27292), .ZN(n27290) );
  OR2_X1 U27296 ( .A1(n27042), .A2(n27043), .ZN(n27292) );
  OR2_X1 U27297 ( .A1(n15242), .A2(n15671), .ZN(n27043) );
  OR2_X1 U27298 ( .A1(n27293), .A2(n27294), .ZN(n27042) );
  AND2_X1 U27299 ( .A1(n27032), .A2(n27031), .ZN(n27294) );
  AND2_X1 U27300 ( .A1(n27027), .A2(n27295), .ZN(n27293) );
  OR2_X1 U27301 ( .A1(n27031), .A2(n27032), .ZN(n27295) );
  OR2_X1 U27302 ( .A1(n15208), .A2(n15671), .ZN(n27032) );
  OR2_X1 U27303 ( .A1(n27296), .A2(n27297), .ZN(n27031) );
  AND2_X1 U27304 ( .A1(n27021), .A2(n27020), .ZN(n27297) );
  AND2_X1 U27305 ( .A1(n27016), .A2(n27298), .ZN(n27296) );
  OR2_X1 U27306 ( .A1(n27020), .A2(n27021), .ZN(n27298) );
  OR2_X1 U27307 ( .A1(n15174), .A2(n15671), .ZN(n27021) );
  OR2_X1 U27308 ( .A1(n27299), .A2(n27300), .ZN(n27020) );
  AND2_X1 U27309 ( .A1(n27010), .A2(n27009), .ZN(n27300) );
  AND2_X1 U27310 ( .A1(n27005), .A2(n27301), .ZN(n27299) );
  OR2_X1 U27311 ( .A1(n27009), .A2(n27010), .ZN(n27301) );
  OR2_X1 U27312 ( .A1(n15140), .A2(n15671), .ZN(n27010) );
  OR2_X1 U27313 ( .A1(n27302), .A2(n27303), .ZN(n27009) );
  AND2_X1 U27314 ( .A1(n26999), .A2(n26998), .ZN(n27303) );
  AND2_X1 U27315 ( .A1(n26994), .A2(n27304), .ZN(n27302) );
  OR2_X1 U27316 ( .A1(n26998), .A2(n26999), .ZN(n27304) );
  OR2_X1 U27317 ( .A1(n15106), .A2(n15671), .ZN(n26999) );
  OR2_X1 U27318 ( .A1(n27305), .A2(n27306), .ZN(n26998) );
  AND2_X1 U27319 ( .A1(n26983), .A2(n26989), .ZN(n27306) );
  AND2_X1 U27320 ( .A1(n27307), .A2(n26988), .ZN(n27305) );
  OR2_X1 U27321 ( .A1(n27308), .A2(n27309), .ZN(n26988) );
  AND2_X1 U27322 ( .A1(n26975), .A2(n26977), .ZN(n27309) );
  AND2_X1 U27323 ( .A1(n26972), .A2(n27310), .ZN(n27308) );
  OR2_X1 U27324 ( .A1(n26977), .A2(n26975), .ZN(n27310) );
  OR2_X1 U27325 ( .A1(n15038), .A2(n15671), .ZN(n26975) );
  OR2_X1 U27326 ( .A1(n27311), .A2(n27312), .ZN(n26977) );
  AND2_X1 U27327 ( .A1(n26961), .A2(n26964), .ZN(n27312) );
  AND2_X1 U27328 ( .A1(n27313), .A2(n26966), .ZN(n27311) );
  OR2_X1 U27329 ( .A1(n27314), .A2(n27315), .ZN(n26966) );
  AND2_X1 U27330 ( .A1(n26950), .A2(n26953), .ZN(n27315) );
  AND2_X1 U27331 ( .A1(n27316), .A2(n26955), .ZN(n27314) );
  OR2_X1 U27332 ( .A1(n27317), .A2(n27318), .ZN(n26955) );
  AND2_X1 U27333 ( .A1(n26939), .A2(n26942), .ZN(n27318) );
  AND2_X1 U27334 ( .A1(n27319), .A2(n26944), .ZN(n27317) );
  OR2_X1 U27335 ( .A1(n27320), .A2(n27321), .ZN(n26944) );
  AND2_X1 U27336 ( .A1(n26928), .A2(n26931), .ZN(n27321) );
  AND2_X1 U27337 ( .A1(n27322), .A2(n26933), .ZN(n27320) );
  OR2_X1 U27338 ( .A1(n27323), .A2(n27324), .ZN(n26933) );
  AND2_X1 U27339 ( .A1(n26916), .A2(n26921), .ZN(n27324) );
  AND2_X1 U27340 ( .A1(n26920), .A2(n27325), .ZN(n27323) );
  OR2_X1 U27341 ( .A1(n26921), .A2(n26916), .ZN(n27325) );
  OR2_X1 U27342 ( .A1(n14857), .A2(n15671), .ZN(n26916) );
  INV_X1 U27343 ( .A(n26922), .ZN(n26921) );
  AND3_X1 U27344 ( .A1(b_6_), .A2(b_5_), .A3(n15957), .ZN(n26922) );
  INV_X1 U27345 ( .A(n26923), .ZN(n26920) );
  OR2_X1 U27346 ( .A1(n27326), .A2(n27327), .ZN(n26923) );
  AND2_X1 U27347 ( .A1(b_5_), .A2(n27328), .ZN(n27327) );
  OR2_X1 U27348 ( .A1(n27329), .A2(n16981), .ZN(n27328) );
  AND2_X1 U27349 ( .A1(a_30_), .A2(n15739), .ZN(n27329) );
  AND2_X1 U27350 ( .A1(b_4_), .A2(n27330), .ZN(n27326) );
  OR2_X1 U27351 ( .A1(n27331), .A2(n14817), .ZN(n27330) );
  AND2_X1 U27352 ( .A1(a_31_), .A2(n15705), .ZN(n27331) );
  OR2_X1 U27353 ( .A1(n26931), .A2(n26928), .ZN(n27322) );
  OR2_X1 U27354 ( .A1(n27332), .A2(n27333), .ZN(n26928) );
  AND2_X1 U27355 ( .A1(n27334), .A2(n27335), .ZN(n27333) );
  INV_X1 U27356 ( .A(n27336), .ZN(n27332) );
  OR2_X1 U27357 ( .A1(n27334), .A2(n27335), .ZN(n27336) );
  OR2_X1 U27358 ( .A1(n27337), .A2(n27338), .ZN(n27334) );
  AND2_X1 U27359 ( .A1(n27339), .A2(n27340), .ZN(n27338) );
  AND2_X1 U27360 ( .A1(n27341), .A2(n27342), .ZN(n27337) );
  OR2_X1 U27361 ( .A1(n14891), .A2(n15671), .ZN(n26931) );
  OR2_X1 U27362 ( .A1(n26942), .A2(n26939), .ZN(n27319) );
  OR2_X1 U27363 ( .A1(n27343), .A2(n27344), .ZN(n26939) );
  INV_X1 U27364 ( .A(n27345), .ZN(n27344) );
  OR2_X1 U27365 ( .A1(n27346), .A2(n27347), .ZN(n27345) );
  AND2_X1 U27366 ( .A1(n27347), .A2(n27346), .ZN(n27343) );
  AND2_X1 U27367 ( .A1(n27348), .A2(n27349), .ZN(n27346) );
  OR2_X1 U27368 ( .A1(n27350), .A2(n27351), .ZN(n27349) );
  INV_X1 U27369 ( .A(n27352), .ZN(n27351) );
  OR2_X1 U27370 ( .A1(n27352), .A2(n27353), .ZN(n27348) );
  INV_X1 U27371 ( .A(n27350), .ZN(n27353) );
  OR2_X1 U27372 ( .A1(n14936), .A2(n15671), .ZN(n26942) );
  OR2_X1 U27373 ( .A1(n26953), .A2(n26950), .ZN(n27316) );
  OR2_X1 U27374 ( .A1(n27354), .A2(n27355), .ZN(n26950) );
  INV_X1 U27375 ( .A(n27356), .ZN(n27355) );
  OR2_X1 U27376 ( .A1(n27357), .A2(n27358), .ZN(n27356) );
  AND2_X1 U27377 ( .A1(n27358), .A2(n27357), .ZN(n27354) );
  AND2_X1 U27378 ( .A1(n27359), .A2(n27360), .ZN(n27357) );
  OR2_X1 U27379 ( .A1(n27361), .A2(n27362), .ZN(n27360) );
  INV_X1 U27380 ( .A(n27363), .ZN(n27362) );
  OR2_X1 U27381 ( .A1(n27363), .A2(n27364), .ZN(n27359) );
  INV_X1 U27382 ( .A(n27361), .ZN(n27364) );
  OR2_X1 U27383 ( .A1(n14970), .A2(n15671), .ZN(n26953) );
  OR2_X1 U27384 ( .A1(n26964), .A2(n26961), .ZN(n27313) );
  OR2_X1 U27385 ( .A1(n27365), .A2(n27366), .ZN(n26961) );
  INV_X1 U27386 ( .A(n27367), .ZN(n27366) );
  OR2_X1 U27387 ( .A1(n27368), .A2(n27369), .ZN(n27367) );
  AND2_X1 U27388 ( .A1(n27369), .A2(n27368), .ZN(n27365) );
  AND2_X1 U27389 ( .A1(n27370), .A2(n27371), .ZN(n27368) );
  OR2_X1 U27390 ( .A1(n27372), .A2(n27373), .ZN(n27371) );
  INV_X1 U27391 ( .A(n27374), .ZN(n27373) );
  OR2_X1 U27392 ( .A1(n27374), .A2(n27375), .ZN(n27370) );
  INV_X1 U27393 ( .A(n27372), .ZN(n27375) );
  OR2_X1 U27394 ( .A1(n15004), .A2(n15671), .ZN(n26964) );
  OR2_X1 U27395 ( .A1(n27376), .A2(n27377), .ZN(n26972) );
  INV_X1 U27396 ( .A(n27378), .ZN(n27377) );
  OR2_X1 U27397 ( .A1(n27379), .A2(n27380), .ZN(n27378) );
  AND2_X1 U27398 ( .A1(n27380), .A2(n27379), .ZN(n27376) );
  AND2_X1 U27399 ( .A1(n27381), .A2(n27382), .ZN(n27379) );
  OR2_X1 U27400 ( .A1(n27383), .A2(n27384), .ZN(n27382) );
  INV_X1 U27401 ( .A(n27385), .ZN(n27384) );
  OR2_X1 U27402 ( .A1(n27385), .A2(n27386), .ZN(n27381) );
  INV_X1 U27403 ( .A(n27383), .ZN(n27386) );
  OR2_X1 U27404 ( .A1(n26989), .A2(n26983), .ZN(n27307) );
  OR2_X1 U27405 ( .A1(n27387), .A2(n27388), .ZN(n26983) );
  INV_X1 U27406 ( .A(n27389), .ZN(n27388) );
  OR2_X1 U27407 ( .A1(n27390), .A2(n27391), .ZN(n27389) );
  AND2_X1 U27408 ( .A1(n27391), .A2(n27390), .ZN(n27387) );
  AND2_X1 U27409 ( .A1(n27392), .A2(n27393), .ZN(n27390) );
  INV_X1 U27410 ( .A(n27394), .ZN(n27393) );
  AND2_X1 U27411 ( .A1(n27395), .A2(n27396), .ZN(n27394) );
  OR2_X1 U27412 ( .A1(n27396), .A2(n27395), .ZN(n27392) );
  INV_X1 U27413 ( .A(n27397), .ZN(n27395) );
  OR2_X1 U27414 ( .A1(n15072), .A2(n15671), .ZN(n26989) );
  INV_X1 U27415 ( .A(b_6_), .ZN(n15671) );
  AND2_X1 U27416 ( .A1(n27398), .A2(n27399), .ZN(n26994) );
  INV_X1 U27417 ( .A(n27400), .ZN(n27399) );
  AND2_X1 U27418 ( .A1(n27401), .A2(n27402), .ZN(n27400) );
  OR2_X1 U27419 ( .A1(n27402), .A2(n27401), .ZN(n27398) );
  OR2_X1 U27420 ( .A1(n27403), .A2(n27404), .ZN(n27401) );
  AND2_X1 U27421 ( .A1(n27405), .A2(n27406), .ZN(n27404) );
  INV_X1 U27422 ( .A(n27407), .ZN(n27405) );
  AND2_X1 U27423 ( .A1(n27408), .A2(n27407), .ZN(n27403) );
  INV_X1 U27424 ( .A(n27406), .ZN(n27408) );
  AND2_X1 U27425 ( .A1(n27409), .A2(n27410), .ZN(n27005) );
  INV_X1 U27426 ( .A(n27411), .ZN(n27410) );
  AND2_X1 U27427 ( .A1(n27412), .A2(n27413), .ZN(n27411) );
  OR2_X1 U27428 ( .A1(n27413), .A2(n27412), .ZN(n27409) );
  OR2_X1 U27429 ( .A1(n27414), .A2(n27415), .ZN(n27412) );
  AND2_X1 U27430 ( .A1(n27416), .A2(n27417), .ZN(n27415) );
  INV_X1 U27431 ( .A(n27418), .ZN(n27416) );
  AND2_X1 U27432 ( .A1(n27419), .A2(n27418), .ZN(n27414) );
  INV_X1 U27433 ( .A(n27417), .ZN(n27419) );
  AND2_X1 U27434 ( .A1(n27420), .A2(n27421), .ZN(n27016) );
  INV_X1 U27435 ( .A(n27422), .ZN(n27421) );
  AND2_X1 U27436 ( .A1(n27423), .A2(n27424), .ZN(n27422) );
  OR2_X1 U27437 ( .A1(n27424), .A2(n27423), .ZN(n27420) );
  OR2_X1 U27438 ( .A1(n27425), .A2(n27426), .ZN(n27423) );
  AND2_X1 U27439 ( .A1(n27427), .A2(n27428), .ZN(n27426) );
  INV_X1 U27440 ( .A(n27429), .ZN(n27427) );
  AND2_X1 U27441 ( .A1(n27430), .A2(n27429), .ZN(n27425) );
  INV_X1 U27442 ( .A(n27428), .ZN(n27430) );
  AND2_X1 U27443 ( .A1(n27431), .A2(n27432), .ZN(n27027) );
  INV_X1 U27444 ( .A(n27433), .ZN(n27432) );
  AND2_X1 U27445 ( .A1(n27434), .A2(n27435), .ZN(n27433) );
  OR2_X1 U27446 ( .A1(n27435), .A2(n27434), .ZN(n27431) );
  OR2_X1 U27447 ( .A1(n27436), .A2(n27437), .ZN(n27434) );
  AND2_X1 U27448 ( .A1(n27438), .A2(n27439), .ZN(n27437) );
  INV_X1 U27449 ( .A(n27440), .ZN(n27438) );
  AND2_X1 U27450 ( .A1(n27441), .A2(n27440), .ZN(n27436) );
  INV_X1 U27451 ( .A(n27439), .ZN(n27441) );
  AND2_X1 U27452 ( .A1(n27442), .A2(n27443), .ZN(n27038) );
  INV_X1 U27453 ( .A(n27444), .ZN(n27443) );
  AND2_X1 U27454 ( .A1(n27445), .A2(n27446), .ZN(n27444) );
  OR2_X1 U27455 ( .A1(n27446), .A2(n27445), .ZN(n27442) );
  OR2_X1 U27456 ( .A1(n27447), .A2(n27448), .ZN(n27445) );
  AND2_X1 U27457 ( .A1(n27449), .A2(n27450), .ZN(n27448) );
  INV_X1 U27458 ( .A(n27451), .ZN(n27449) );
  AND2_X1 U27459 ( .A1(n27452), .A2(n27451), .ZN(n27447) );
  INV_X1 U27460 ( .A(n27450), .ZN(n27452) );
  AND2_X1 U27461 ( .A1(n27453), .A2(n27454), .ZN(n27049) );
  INV_X1 U27462 ( .A(n27455), .ZN(n27454) );
  AND2_X1 U27463 ( .A1(n27456), .A2(n27457), .ZN(n27455) );
  OR2_X1 U27464 ( .A1(n27457), .A2(n27456), .ZN(n27453) );
  OR2_X1 U27465 ( .A1(n27458), .A2(n27459), .ZN(n27456) );
  AND2_X1 U27466 ( .A1(n27460), .A2(n27461), .ZN(n27459) );
  INV_X1 U27467 ( .A(n27462), .ZN(n27460) );
  AND2_X1 U27468 ( .A1(n27463), .A2(n27462), .ZN(n27458) );
  INV_X1 U27469 ( .A(n27461), .ZN(n27463) );
  AND2_X1 U27470 ( .A1(n27464), .A2(n27465), .ZN(n27060) );
  INV_X1 U27471 ( .A(n27466), .ZN(n27465) );
  AND2_X1 U27472 ( .A1(n27467), .A2(n27468), .ZN(n27466) );
  OR2_X1 U27473 ( .A1(n27468), .A2(n27467), .ZN(n27464) );
  OR2_X1 U27474 ( .A1(n27469), .A2(n27470), .ZN(n27467) );
  AND2_X1 U27475 ( .A1(n27471), .A2(n27472), .ZN(n27470) );
  INV_X1 U27476 ( .A(n27473), .ZN(n27471) );
  AND2_X1 U27477 ( .A1(n27474), .A2(n27473), .ZN(n27469) );
  INV_X1 U27478 ( .A(n27472), .ZN(n27474) );
  AND2_X1 U27479 ( .A1(n27475), .A2(n27476), .ZN(n27071) );
  INV_X1 U27480 ( .A(n27477), .ZN(n27476) );
  AND2_X1 U27481 ( .A1(n27478), .A2(n27479), .ZN(n27477) );
  OR2_X1 U27482 ( .A1(n27479), .A2(n27478), .ZN(n27475) );
  OR2_X1 U27483 ( .A1(n27480), .A2(n27481), .ZN(n27478) );
  AND2_X1 U27484 ( .A1(n27482), .A2(n27483), .ZN(n27481) );
  INV_X1 U27485 ( .A(n27484), .ZN(n27482) );
  AND2_X1 U27486 ( .A1(n27485), .A2(n27484), .ZN(n27480) );
  INV_X1 U27487 ( .A(n27483), .ZN(n27485) );
  AND2_X1 U27488 ( .A1(n27486), .A2(n27487), .ZN(n27082) );
  INV_X1 U27489 ( .A(n27488), .ZN(n27487) );
  AND2_X1 U27490 ( .A1(n27489), .A2(n27490), .ZN(n27488) );
  OR2_X1 U27491 ( .A1(n27490), .A2(n27489), .ZN(n27486) );
  OR2_X1 U27492 ( .A1(n27491), .A2(n27492), .ZN(n27489) );
  AND2_X1 U27493 ( .A1(n27493), .A2(n27494), .ZN(n27492) );
  INV_X1 U27494 ( .A(n27495), .ZN(n27493) );
  AND2_X1 U27495 ( .A1(n27496), .A2(n27495), .ZN(n27491) );
  INV_X1 U27496 ( .A(n27494), .ZN(n27496) );
  AND2_X1 U27497 ( .A1(n27497), .A2(n27498), .ZN(n27093) );
  INV_X1 U27498 ( .A(n27499), .ZN(n27498) );
  AND2_X1 U27499 ( .A1(n27500), .A2(n27501), .ZN(n27499) );
  OR2_X1 U27500 ( .A1(n27501), .A2(n27500), .ZN(n27497) );
  OR2_X1 U27501 ( .A1(n27502), .A2(n27503), .ZN(n27500) );
  AND2_X1 U27502 ( .A1(n27504), .A2(n27505), .ZN(n27503) );
  INV_X1 U27503 ( .A(n27506), .ZN(n27504) );
  AND2_X1 U27504 ( .A1(n27507), .A2(n27506), .ZN(n27502) );
  INV_X1 U27505 ( .A(n27505), .ZN(n27507) );
  AND2_X1 U27506 ( .A1(n27508), .A2(n27509), .ZN(n27104) );
  INV_X1 U27507 ( .A(n27510), .ZN(n27509) );
  AND2_X1 U27508 ( .A1(n27511), .A2(n27512), .ZN(n27510) );
  OR2_X1 U27509 ( .A1(n27512), .A2(n27511), .ZN(n27508) );
  OR2_X1 U27510 ( .A1(n27513), .A2(n27514), .ZN(n27511) );
  AND2_X1 U27511 ( .A1(n27515), .A2(n27516), .ZN(n27514) );
  INV_X1 U27512 ( .A(n27517), .ZN(n27515) );
  AND2_X1 U27513 ( .A1(n27518), .A2(n27517), .ZN(n27513) );
  INV_X1 U27514 ( .A(n27516), .ZN(n27518) );
  AND2_X1 U27515 ( .A1(n27519), .A2(n27520), .ZN(n27115) );
  INV_X1 U27516 ( .A(n27521), .ZN(n27520) );
  AND2_X1 U27517 ( .A1(n27522), .A2(n27523), .ZN(n27521) );
  OR2_X1 U27518 ( .A1(n27523), .A2(n27522), .ZN(n27519) );
  OR2_X1 U27519 ( .A1(n27524), .A2(n27525), .ZN(n27522) );
  AND2_X1 U27520 ( .A1(n27526), .A2(n27527), .ZN(n27525) );
  INV_X1 U27521 ( .A(n27528), .ZN(n27526) );
  AND2_X1 U27522 ( .A1(n27529), .A2(n27528), .ZN(n27524) );
  INV_X1 U27523 ( .A(n27527), .ZN(n27529) );
  AND2_X1 U27524 ( .A1(n27530), .A2(n27531), .ZN(n27126) );
  INV_X1 U27525 ( .A(n27532), .ZN(n27531) );
  AND2_X1 U27526 ( .A1(n27533), .A2(n27534), .ZN(n27532) );
  OR2_X1 U27527 ( .A1(n27534), .A2(n27533), .ZN(n27530) );
  OR2_X1 U27528 ( .A1(n27535), .A2(n27536), .ZN(n27533) );
  AND2_X1 U27529 ( .A1(n27537), .A2(n27538), .ZN(n27536) );
  INV_X1 U27530 ( .A(n27539), .ZN(n27537) );
  AND2_X1 U27531 ( .A1(n27540), .A2(n27539), .ZN(n27535) );
  INV_X1 U27532 ( .A(n27538), .ZN(n27540) );
  AND2_X1 U27533 ( .A1(n27541), .A2(n27542), .ZN(n27137) );
  INV_X1 U27534 ( .A(n27543), .ZN(n27542) );
  AND2_X1 U27535 ( .A1(n27544), .A2(n27545), .ZN(n27543) );
  OR2_X1 U27536 ( .A1(n27545), .A2(n27544), .ZN(n27541) );
  OR2_X1 U27537 ( .A1(n27546), .A2(n27547), .ZN(n27544) );
  AND2_X1 U27538 ( .A1(n27548), .A2(n27549), .ZN(n27547) );
  INV_X1 U27539 ( .A(n27550), .ZN(n27548) );
  AND2_X1 U27540 ( .A1(n27551), .A2(n27550), .ZN(n27546) );
  INV_X1 U27541 ( .A(n27549), .ZN(n27551) );
  AND2_X1 U27542 ( .A1(n27552), .A2(n27553), .ZN(n27148) );
  INV_X1 U27543 ( .A(n27554), .ZN(n27553) );
  AND2_X1 U27544 ( .A1(n27555), .A2(n27556), .ZN(n27554) );
  OR2_X1 U27545 ( .A1(n27556), .A2(n27555), .ZN(n27552) );
  OR2_X1 U27546 ( .A1(n27557), .A2(n27558), .ZN(n27555) );
  AND2_X1 U27547 ( .A1(n27559), .A2(n27560), .ZN(n27558) );
  INV_X1 U27548 ( .A(n27561), .ZN(n27559) );
  AND2_X1 U27549 ( .A1(n27562), .A2(n27561), .ZN(n27557) );
  INV_X1 U27550 ( .A(n27560), .ZN(n27562) );
  AND2_X1 U27551 ( .A1(n27563), .A2(n27564), .ZN(n27159) );
  INV_X1 U27552 ( .A(n27565), .ZN(n27564) );
  AND2_X1 U27553 ( .A1(n27566), .A2(n27567), .ZN(n27565) );
  OR2_X1 U27554 ( .A1(n27567), .A2(n27566), .ZN(n27563) );
  OR2_X1 U27555 ( .A1(n27568), .A2(n27569), .ZN(n27566) );
  AND2_X1 U27556 ( .A1(n27570), .A2(n27571), .ZN(n27569) );
  INV_X1 U27557 ( .A(n27572), .ZN(n27570) );
  AND2_X1 U27558 ( .A1(n27573), .A2(n27572), .ZN(n27568) );
  INV_X1 U27559 ( .A(n27571), .ZN(n27573) );
  AND2_X1 U27560 ( .A1(n27574), .A2(n27575), .ZN(n27170) );
  INV_X1 U27561 ( .A(n27576), .ZN(n27575) );
  AND2_X1 U27562 ( .A1(n27577), .A2(n27578), .ZN(n27576) );
  OR2_X1 U27563 ( .A1(n27578), .A2(n27577), .ZN(n27574) );
  OR2_X1 U27564 ( .A1(n27579), .A2(n27580), .ZN(n27577) );
  AND2_X1 U27565 ( .A1(n27581), .A2(n27582), .ZN(n27580) );
  INV_X1 U27566 ( .A(n27583), .ZN(n27581) );
  AND2_X1 U27567 ( .A1(n27584), .A2(n27583), .ZN(n27579) );
  INV_X1 U27568 ( .A(n27582), .ZN(n27584) );
  AND2_X1 U27569 ( .A1(n27585), .A2(n27586), .ZN(n27180) );
  INV_X1 U27570 ( .A(n27587), .ZN(n27586) );
  AND2_X1 U27571 ( .A1(n27588), .A2(n27589), .ZN(n27587) );
  OR2_X1 U27572 ( .A1(n27589), .A2(n27588), .ZN(n27585) );
  OR2_X1 U27573 ( .A1(n27590), .A2(n27591), .ZN(n27588) );
  AND2_X1 U27574 ( .A1(n27592), .A2(n27593), .ZN(n27591) );
  INV_X1 U27575 ( .A(n27594), .ZN(n27592) );
  AND2_X1 U27576 ( .A1(n27595), .A2(n27594), .ZN(n27590) );
  INV_X1 U27577 ( .A(n27593), .ZN(n27595) );
  AND2_X1 U27578 ( .A1(n27596), .A2(n27597), .ZN(n27191) );
  INV_X1 U27579 ( .A(n27598), .ZN(n27597) );
  AND2_X1 U27580 ( .A1(n27599), .A2(n27600), .ZN(n27598) );
  OR2_X1 U27581 ( .A1(n27600), .A2(n27599), .ZN(n27596) );
  OR2_X1 U27582 ( .A1(n27601), .A2(n27602), .ZN(n27599) );
  AND2_X1 U27583 ( .A1(n27603), .A2(n27604), .ZN(n27602) );
  INV_X1 U27584 ( .A(n15882), .ZN(n27603) );
  AND2_X1 U27585 ( .A1(n27605), .A2(n15882), .ZN(n27601) );
  INV_X1 U27586 ( .A(n27604), .ZN(n27605) );
  AND2_X1 U27587 ( .A1(n27606), .A2(n27607), .ZN(n27202) );
  INV_X1 U27588 ( .A(n27608), .ZN(n27607) );
  AND2_X1 U27589 ( .A1(n27609), .A2(n27610), .ZN(n27608) );
  OR2_X1 U27590 ( .A1(n27610), .A2(n27609), .ZN(n27606) );
  OR2_X1 U27591 ( .A1(n27611), .A2(n27612), .ZN(n27609) );
  AND2_X1 U27592 ( .A1(n27613), .A2(n27614), .ZN(n27612) );
  INV_X1 U27593 ( .A(n27615), .ZN(n27613) );
  AND2_X1 U27594 ( .A1(n27616), .A2(n27615), .ZN(n27611) );
  INV_X1 U27595 ( .A(n27614), .ZN(n27616) );
  AND2_X1 U27596 ( .A1(n27617), .A2(n27618), .ZN(n27213) );
  INV_X1 U27597 ( .A(n27619), .ZN(n27618) );
  AND2_X1 U27598 ( .A1(n27620), .A2(n27621), .ZN(n27619) );
  OR2_X1 U27599 ( .A1(n27621), .A2(n27620), .ZN(n27617) );
  OR2_X1 U27600 ( .A1(n27622), .A2(n27623), .ZN(n27620) );
  AND2_X1 U27601 ( .A1(n27624), .A2(n27625), .ZN(n27623) );
  INV_X1 U27602 ( .A(n27626), .ZN(n27624) );
  AND2_X1 U27603 ( .A1(n27627), .A2(n27626), .ZN(n27622) );
  INV_X1 U27604 ( .A(n27625), .ZN(n27627) );
  AND2_X1 U27605 ( .A1(n27628), .A2(n27629), .ZN(n27224) );
  INV_X1 U27606 ( .A(n27630), .ZN(n27629) );
  AND2_X1 U27607 ( .A1(n27631), .A2(n27632), .ZN(n27630) );
  OR2_X1 U27608 ( .A1(n27632), .A2(n27631), .ZN(n27628) );
  OR2_X1 U27609 ( .A1(n27633), .A2(n27634), .ZN(n27631) );
  AND2_X1 U27610 ( .A1(n27635), .A2(n27636), .ZN(n27634) );
  INV_X1 U27611 ( .A(n27637), .ZN(n27635) );
  AND2_X1 U27612 ( .A1(n27638), .A2(n27637), .ZN(n27633) );
  INV_X1 U27613 ( .A(n27636), .ZN(n27638) );
  AND2_X1 U27614 ( .A1(n27639), .A2(n27640), .ZN(n16431) );
  INV_X1 U27615 ( .A(n27641), .ZN(n27640) );
  AND2_X1 U27616 ( .A1(n27642), .A2(n27643), .ZN(n27641) );
  OR2_X1 U27617 ( .A1(n27643), .A2(n27642), .ZN(n27639) );
  OR2_X1 U27618 ( .A1(n27644), .A2(n27645), .ZN(n27642) );
  AND2_X1 U27619 ( .A1(n27646), .A2(n27647), .ZN(n27645) );
  INV_X1 U27620 ( .A(n27648), .ZN(n27646) );
  AND2_X1 U27621 ( .A1(n27649), .A2(n27648), .ZN(n27644) );
  INV_X1 U27622 ( .A(n27647), .ZN(n27649) );
  OR2_X1 U27623 ( .A1(n16421), .A2(n16422), .ZN(n15251) );
  OR2_X1 U27624 ( .A1(n27650), .A2(n27651), .ZN(n16422) );
  AND2_X1 U27625 ( .A1(n16442), .A2(n16441), .ZN(n27651) );
  AND2_X1 U27626 ( .A1(n16437), .A2(n27652), .ZN(n27650) );
  OR2_X1 U27627 ( .A1(n16441), .A2(n16442), .ZN(n27652) );
  OR2_X1 U27628 ( .A1(n16512), .A2(n15705), .ZN(n16442) );
  OR2_X1 U27629 ( .A1(n27653), .A2(n27654), .ZN(n16441) );
  AND2_X1 U27630 ( .A1(n27648), .A2(n27647), .ZN(n27654) );
  AND2_X1 U27631 ( .A1(n27643), .A2(n27655), .ZN(n27653) );
  OR2_X1 U27632 ( .A1(n27647), .A2(n27648), .ZN(n27655) );
  OR2_X1 U27633 ( .A1(n15842), .A2(n15705), .ZN(n27648) );
  OR2_X1 U27634 ( .A1(n27656), .A2(n27657), .ZN(n27647) );
  AND2_X1 U27635 ( .A1(n27637), .A2(n27636), .ZN(n27657) );
  AND2_X1 U27636 ( .A1(n27632), .A2(n27658), .ZN(n27656) );
  OR2_X1 U27637 ( .A1(n27636), .A2(n27637), .ZN(n27658) );
  OR2_X1 U27638 ( .A1(n15808), .A2(n15705), .ZN(n27637) );
  OR2_X1 U27639 ( .A1(n27659), .A2(n27660), .ZN(n27636) );
  AND2_X1 U27640 ( .A1(n27626), .A2(n27625), .ZN(n27660) );
  AND2_X1 U27641 ( .A1(n27621), .A2(n27661), .ZN(n27659) );
  OR2_X1 U27642 ( .A1(n27625), .A2(n27626), .ZN(n27661) );
  OR2_X1 U27643 ( .A1(n15774), .A2(n15705), .ZN(n27626) );
  OR2_X1 U27644 ( .A1(n27662), .A2(n27663), .ZN(n27625) );
  AND2_X1 U27645 ( .A1(n27615), .A2(n27614), .ZN(n27663) );
  AND2_X1 U27646 ( .A1(n27610), .A2(n27664), .ZN(n27662) );
  OR2_X1 U27647 ( .A1(n27614), .A2(n27615), .ZN(n27664) );
  OR2_X1 U27648 ( .A1(n15740), .A2(n15705), .ZN(n27615) );
  OR2_X1 U27649 ( .A1(n27665), .A2(n27666), .ZN(n27614) );
  AND2_X1 U27650 ( .A1(n15882), .A2(n27604), .ZN(n27666) );
  AND2_X1 U27651 ( .A1(n27600), .A2(n27667), .ZN(n27665) );
  OR2_X1 U27652 ( .A1(n27604), .A2(n15882), .ZN(n27667) );
  OR2_X1 U27653 ( .A1(n15706), .A2(n15705), .ZN(n15882) );
  OR2_X1 U27654 ( .A1(n27668), .A2(n27669), .ZN(n27604) );
  AND2_X1 U27655 ( .A1(n27594), .A2(n27593), .ZN(n27669) );
  AND2_X1 U27656 ( .A1(n27589), .A2(n27670), .ZN(n27668) );
  OR2_X1 U27657 ( .A1(n27593), .A2(n27594), .ZN(n27670) );
  OR2_X1 U27658 ( .A1(n15672), .A2(n15705), .ZN(n27594) );
  OR2_X1 U27659 ( .A1(n27671), .A2(n27672), .ZN(n27593) );
  AND2_X1 U27660 ( .A1(n27583), .A2(n27582), .ZN(n27672) );
  AND2_X1 U27661 ( .A1(n27578), .A2(n27673), .ZN(n27671) );
  OR2_X1 U27662 ( .A1(n27582), .A2(n27583), .ZN(n27673) );
  OR2_X1 U27663 ( .A1(n15638), .A2(n15705), .ZN(n27583) );
  OR2_X1 U27664 ( .A1(n27674), .A2(n27675), .ZN(n27582) );
  AND2_X1 U27665 ( .A1(n27572), .A2(n27571), .ZN(n27675) );
  AND2_X1 U27666 ( .A1(n27567), .A2(n27676), .ZN(n27674) );
  OR2_X1 U27667 ( .A1(n27571), .A2(n27572), .ZN(n27676) );
  OR2_X1 U27668 ( .A1(n15593), .A2(n15705), .ZN(n27572) );
  OR2_X1 U27669 ( .A1(n27677), .A2(n27678), .ZN(n27571) );
  AND2_X1 U27670 ( .A1(n27561), .A2(n27560), .ZN(n27678) );
  AND2_X1 U27671 ( .A1(n27556), .A2(n27679), .ZN(n27677) );
  OR2_X1 U27672 ( .A1(n27560), .A2(n27561), .ZN(n27679) );
  OR2_X1 U27673 ( .A1(n15559), .A2(n15705), .ZN(n27561) );
  OR2_X1 U27674 ( .A1(n27680), .A2(n27681), .ZN(n27560) );
  AND2_X1 U27675 ( .A1(n27550), .A2(n27549), .ZN(n27681) );
  AND2_X1 U27676 ( .A1(n27545), .A2(n27682), .ZN(n27680) );
  OR2_X1 U27677 ( .A1(n27549), .A2(n27550), .ZN(n27682) );
  OR2_X1 U27678 ( .A1(n15525), .A2(n15705), .ZN(n27550) );
  OR2_X1 U27679 ( .A1(n27683), .A2(n27684), .ZN(n27549) );
  AND2_X1 U27680 ( .A1(n27539), .A2(n27538), .ZN(n27684) );
  AND2_X1 U27681 ( .A1(n27534), .A2(n27685), .ZN(n27683) );
  OR2_X1 U27682 ( .A1(n27538), .A2(n27539), .ZN(n27685) );
  OR2_X1 U27683 ( .A1(n15491), .A2(n15705), .ZN(n27539) );
  OR2_X1 U27684 ( .A1(n27686), .A2(n27687), .ZN(n27538) );
  AND2_X1 U27685 ( .A1(n27528), .A2(n27527), .ZN(n27687) );
  AND2_X1 U27686 ( .A1(n27523), .A2(n27688), .ZN(n27686) );
  OR2_X1 U27687 ( .A1(n27527), .A2(n27528), .ZN(n27688) );
  OR2_X1 U27688 ( .A1(n15457), .A2(n15705), .ZN(n27528) );
  OR2_X1 U27689 ( .A1(n27689), .A2(n27690), .ZN(n27527) );
  AND2_X1 U27690 ( .A1(n27517), .A2(n27516), .ZN(n27690) );
  AND2_X1 U27691 ( .A1(n27512), .A2(n27691), .ZN(n27689) );
  OR2_X1 U27692 ( .A1(n27516), .A2(n27517), .ZN(n27691) );
  OR2_X1 U27693 ( .A1(n15423), .A2(n15705), .ZN(n27517) );
  OR2_X1 U27694 ( .A1(n27692), .A2(n27693), .ZN(n27516) );
  AND2_X1 U27695 ( .A1(n27506), .A2(n27505), .ZN(n27693) );
  AND2_X1 U27696 ( .A1(n27501), .A2(n27694), .ZN(n27692) );
  OR2_X1 U27697 ( .A1(n27505), .A2(n27506), .ZN(n27694) );
  OR2_X1 U27698 ( .A1(n15389), .A2(n15705), .ZN(n27506) );
  OR2_X1 U27699 ( .A1(n27695), .A2(n27696), .ZN(n27505) );
  AND2_X1 U27700 ( .A1(n27495), .A2(n27494), .ZN(n27696) );
  AND2_X1 U27701 ( .A1(n27490), .A2(n27697), .ZN(n27695) );
  OR2_X1 U27702 ( .A1(n27494), .A2(n27495), .ZN(n27697) );
  OR2_X1 U27703 ( .A1(n15355), .A2(n15705), .ZN(n27495) );
  OR2_X1 U27704 ( .A1(n27698), .A2(n27699), .ZN(n27494) );
  AND2_X1 U27705 ( .A1(n27484), .A2(n27483), .ZN(n27699) );
  AND2_X1 U27706 ( .A1(n27479), .A2(n27700), .ZN(n27698) );
  OR2_X1 U27707 ( .A1(n27483), .A2(n27484), .ZN(n27700) );
  OR2_X1 U27708 ( .A1(n15321), .A2(n15705), .ZN(n27484) );
  OR2_X1 U27709 ( .A1(n27701), .A2(n27702), .ZN(n27483) );
  AND2_X1 U27710 ( .A1(n27473), .A2(n27472), .ZN(n27702) );
  AND2_X1 U27711 ( .A1(n27468), .A2(n27703), .ZN(n27701) );
  OR2_X1 U27712 ( .A1(n27472), .A2(n27473), .ZN(n27703) );
  OR2_X1 U27713 ( .A1(n15287), .A2(n15705), .ZN(n27473) );
  OR2_X1 U27714 ( .A1(n27704), .A2(n27705), .ZN(n27472) );
  AND2_X1 U27715 ( .A1(n27462), .A2(n27461), .ZN(n27705) );
  AND2_X1 U27716 ( .A1(n27457), .A2(n27706), .ZN(n27704) );
  OR2_X1 U27717 ( .A1(n27461), .A2(n27462), .ZN(n27706) );
  OR2_X1 U27718 ( .A1(n15242), .A2(n15705), .ZN(n27462) );
  OR2_X1 U27719 ( .A1(n27707), .A2(n27708), .ZN(n27461) );
  AND2_X1 U27720 ( .A1(n27451), .A2(n27450), .ZN(n27708) );
  AND2_X1 U27721 ( .A1(n27446), .A2(n27709), .ZN(n27707) );
  OR2_X1 U27722 ( .A1(n27450), .A2(n27451), .ZN(n27709) );
  OR2_X1 U27723 ( .A1(n15208), .A2(n15705), .ZN(n27451) );
  OR2_X1 U27724 ( .A1(n27710), .A2(n27711), .ZN(n27450) );
  AND2_X1 U27725 ( .A1(n27440), .A2(n27439), .ZN(n27711) );
  AND2_X1 U27726 ( .A1(n27435), .A2(n27712), .ZN(n27710) );
  OR2_X1 U27727 ( .A1(n27439), .A2(n27440), .ZN(n27712) );
  OR2_X1 U27728 ( .A1(n15174), .A2(n15705), .ZN(n27440) );
  OR2_X1 U27729 ( .A1(n27713), .A2(n27714), .ZN(n27439) );
  AND2_X1 U27730 ( .A1(n27429), .A2(n27428), .ZN(n27714) );
  AND2_X1 U27731 ( .A1(n27424), .A2(n27715), .ZN(n27713) );
  OR2_X1 U27732 ( .A1(n27428), .A2(n27429), .ZN(n27715) );
  OR2_X1 U27733 ( .A1(n15140), .A2(n15705), .ZN(n27429) );
  OR2_X1 U27734 ( .A1(n27716), .A2(n27717), .ZN(n27428) );
  AND2_X1 U27735 ( .A1(n27418), .A2(n27417), .ZN(n27717) );
  AND2_X1 U27736 ( .A1(n27413), .A2(n27718), .ZN(n27716) );
  OR2_X1 U27737 ( .A1(n27417), .A2(n27418), .ZN(n27718) );
  OR2_X1 U27738 ( .A1(n15106), .A2(n15705), .ZN(n27418) );
  OR2_X1 U27739 ( .A1(n27719), .A2(n27720), .ZN(n27417) );
  AND2_X1 U27740 ( .A1(n27407), .A2(n27406), .ZN(n27720) );
  AND2_X1 U27741 ( .A1(n27402), .A2(n27721), .ZN(n27719) );
  OR2_X1 U27742 ( .A1(n27406), .A2(n27407), .ZN(n27721) );
  OR2_X1 U27743 ( .A1(n15072), .A2(n15705), .ZN(n27407) );
  OR2_X1 U27744 ( .A1(n27722), .A2(n27723), .ZN(n27406) );
  AND2_X1 U27745 ( .A1(n27391), .A2(n27397), .ZN(n27723) );
  AND2_X1 U27746 ( .A1(n27724), .A2(n27396), .ZN(n27722) );
  OR2_X1 U27747 ( .A1(n27725), .A2(n27726), .ZN(n27396) );
  AND2_X1 U27748 ( .A1(n27383), .A2(n27385), .ZN(n27726) );
  AND2_X1 U27749 ( .A1(n27380), .A2(n27727), .ZN(n27725) );
  OR2_X1 U27750 ( .A1(n27385), .A2(n27383), .ZN(n27727) );
  OR2_X1 U27751 ( .A1(n15004), .A2(n15705), .ZN(n27383) );
  OR2_X1 U27752 ( .A1(n27728), .A2(n27729), .ZN(n27385) );
  AND2_X1 U27753 ( .A1(n27369), .A2(n27372), .ZN(n27729) );
  AND2_X1 U27754 ( .A1(n27730), .A2(n27374), .ZN(n27728) );
  OR2_X1 U27755 ( .A1(n27731), .A2(n27732), .ZN(n27374) );
  AND2_X1 U27756 ( .A1(n27358), .A2(n27361), .ZN(n27732) );
  AND2_X1 U27757 ( .A1(n27733), .A2(n27363), .ZN(n27731) );
  OR2_X1 U27758 ( .A1(n27734), .A2(n27735), .ZN(n27363) );
  AND2_X1 U27759 ( .A1(n27347), .A2(n27350), .ZN(n27735) );
  AND2_X1 U27760 ( .A1(n27736), .A2(n27352), .ZN(n27734) );
  OR2_X1 U27761 ( .A1(n27737), .A2(n27738), .ZN(n27352) );
  AND2_X1 U27762 ( .A1(n27335), .A2(n27340), .ZN(n27738) );
  AND2_X1 U27763 ( .A1(n27339), .A2(n27739), .ZN(n27737) );
  OR2_X1 U27764 ( .A1(n27340), .A2(n27335), .ZN(n27739) );
  OR2_X1 U27765 ( .A1(n14857), .A2(n15705), .ZN(n27335) );
  INV_X1 U27766 ( .A(n27341), .ZN(n27340) );
  AND3_X1 U27767 ( .A1(b_5_), .A2(b_4_), .A3(n15957), .ZN(n27341) );
  INV_X1 U27768 ( .A(n27342), .ZN(n27339) );
  OR2_X1 U27769 ( .A1(n27740), .A2(n27741), .ZN(n27342) );
  AND2_X1 U27770 ( .A1(b_4_), .A2(n27742), .ZN(n27741) );
  OR2_X1 U27771 ( .A1(n27743), .A2(n16981), .ZN(n27742) );
  AND2_X1 U27772 ( .A1(a_30_), .A2(n15773), .ZN(n27743) );
  AND2_X1 U27773 ( .A1(b_3_), .A2(n27744), .ZN(n27740) );
  OR2_X1 U27774 ( .A1(n27745), .A2(n14817), .ZN(n27744) );
  AND2_X1 U27775 ( .A1(a_31_), .A2(n15739), .ZN(n27745) );
  OR2_X1 U27776 ( .A1(n27350), .A2(n27347), .ZN(n27736) );
  OR2_X1 U27777 ( .A1(n27746), .A2(n27747), .ZN(n27347) );
  AND2_X1 U27778 ( .A1(n27748), .A2(n27749), .ZN(n27747) );
  INV_X1 U27779 ( .A(n27750), .ZN(n27746) );
  OR2_X1 U27780 ( .A1(n27748), .A2(n27749), .ZN(n27750) );
  OR2_X1 U27781 ( .A1(n27751), .A2(n27752), .ZN(n27748) );
  AND2_X1 U27782 ( .A1(n27753), .A2(n27754), .ZN(n27752) );
  AND2_X1 U27783 ( .A1(n27755), .A2(n27756), .ZN(n27751) );
  OR2_X1 U27784 ( .A1(n14891), .A2(n15705), .ZN(n27350) );
  OR2_X1 U27785 ( .A1(n27361), .A2(n27358), .ZN(n27733) );
  OR2_X1 U27786 ( .A1(n27757), .A2(n27758), .ZN(n27358) );
  INV_X1 U27787 ( .A(n27759), .ZN(n27758) );
  OR2_X1 U27788 ( .A1(n27760), .A2(n27761), .ZN(n27759) );
  AND2_X1 U27789 ( .A1(n27761), .A2(n27760), .ZN(n27757) );
  AND2_X1 U27790 ( .A1(n27762), .A2(n27763), .ZN(n27760) );
  OR2_X1 U27791 ( .A1(n27764), .A2(n27765), .ZN(n27763) );
  INV_X1 U27792 ( .A(n27766), .ZN(n27765) );
  OR2_X1 U27793 ( .A1(n27766), .A2(n27767), .ZN(n27762) );
  INV_X1 U27794 ( .A(n27764), .ZN(n27767) );
  OR2_X1 U27795 ( .A1(n14936), .A2(n15705), .ZN(n27361) );
  OR2_X1 U27796 ( .A1(n27372), .A2(n27369), .ZN(n27730) );
  OR2_X1 U27797 ( .A1(n27768), .A2(n27769), .ZN(n27369) );
  INV_X1 U27798 ( .A(n27770), .ZN(n27769) );
  OR2_X1 U27799 ( .A1(n27771), .A2(n27772), .ZN(n27770) );
  AND2_X1 U27800 ( .A1(n27772), .A2(n27771), .ZN(n27768) );
  AND2_X1 U27801 ( .A1(n27773), .A2(n27774), .ZN(n27771) );
  OR2_X1 U27802 ( .A1(n27775), .A2(n27776), .ZN(n27774) );
  INV_X1 U27803 ( .A(n27777), .ZN(n27776) );
  OR2_X1 U27804 ( .A1(n27777), .A2(n27778), .ZN(n27773) );
  INV_X1 U27805 ( .A(n27775), .ZN(n27778) );
  OR2_X1 U27806 ( .A1(n14970), .A2(n15705), .ZN(n27372) );
  OR2_X1 U27807 ( .A1(n27779), .A2(n27780), .ZN(n27380) );
  INV_X1 U27808 ( .A(n27781), .ZN(n27780) );
  OR2_X1 U27809 ( .A1(n27782), .A2(n27783), .ZN(n27781) );
  AND2_X1 U27810 ( .A1(n27783), .A2(n27782), .ZN(n27779) );
  AND2_X1 U27811 ( .A1(n27784), .A2(n27785), .ZN(n27782) );
  OR2_X1 U27812 ( .A1(n27786), .A2(n27787), .ZN(n27785) );
  INV_X1 U27813 ( .A(n27788), .ZN(n27787) );
  OR2_X1 U27814 ( .A1(n27788), .A2(n27789), .ZN(n27784) );
  INV_X1 U27815 ( .A(n27786), .ZN(n27789) );
  OR2_X1 U27816 ( .A1(n27397), .A2(n27391), .ZN(n27724) );
  OR2_X1 U27817 ( .A1(n27790), .A2(n27791), .ZN(n27391) );
  INV_X1 U27818 ( .A(n27792), .ZN(n27791) );
  OR2_X1 U27819 ( .A1(n27793), .A2(n27794), .ZN(n27792) );
  AND2_X1 U27820 ( .A1(n27794), .A2(n27793), .ZN(n27790) );
  AND2_X1 U27821 ( .A1(n27795), .A2(n27796), .ZN(n27793) );
  INV_X1 U27822 ( .A(n27797), .ZN(n27796) );
  AND2_X1 U27823 ( .A1(n27798), .A2(n27799), .ZN(n27797) );
  OR2_X1 U27824 ( .A1(n27799), .A2(n27798), .ZN(n27795) );
  INV_X1 U27825 ( .A(n27800), .ZN(n27798) );
  OR2_X1 U27826 ( .A1(n15038), .A2(n15705), .ZN(n27397) );
  INV_X1 U27827 ( .A(b_5_), .ZN(n15705) );
  AND2_X1 U27828 ( .A1(n27801), .A2(n27802), .ZN(n27402) );
  INV_X1 U27829 ( .A(n27803), .ZN(n27802) );
  AND2_X1 U27830 ( .A1(n27804), .A2(n27805), .ZN(n27803) );
  OR2_X1 U27831 ( .A1(n27805), .A2(n27804), .ZN(n27801) );
  OR2_X1 U27832 ( .A1(n27806), .A2(n27807), .ZN(n27804) );
  AND2_X1 U27833 ( .A1(n27808), .A2(n27809), .ZN(n27807) );
  INV_X1 U27834 ( .A(n27810), .ZN(n27808) );
  AND2_X1 U27835 ( .A1(n27811), .A2(n27810), .ZN(n27806) );
  INV_X1 U27836 ( .A(n27809), .ZN(n27811) );
  AND2_X1 U27837 ( .A1(n27812), .A2(n27813), .ZN(n27413) );
  INV_X1 U27838 ( .A(n27814), .ZN(n27813) );
  AND2_X1 U27839 ( .A1(n27815), .A2(n27816), .ZN(n27814) );
  OR2_X1 U27840 ( .A1(n27816), .A2(n27815), .ZN(n27812) );
  OR2_X1 U27841 ( .A1(n27817), .A2(n27818), .ZN(n27815) );
  AND2_X1 U27842 ( .A1(n27819), .A2(n27820), .ZN(n27818) );
  INV_X1 U27843 ( .A(n27821), .ZN(n27819) );
  AND2_X1 U27844 ( .A1(n27822), .A2(n27821), .ZN(n27817) );
  INV_X1 U27845 ( .A(n27820), .ZN(n27822) );
  AND2_X1 U27846 ( .A1(n27823), .A2(n27824), .ZN(n27424) );
  INV_X1 U27847 ( .A(n27825), .ZN(n27824) );
  AND2_X1 U27848 ( .A1(n27826), .A2(n27827), .ZN(n27825) );
  OR2_X1 U27849 ( .A1(n27827), .A2(n27826), .ZN(n27823) );
  OR2_X1 U27850 ( .A1(n27828), .A2(n27829), .ZN(n27826) );
  AND2_X1 U27851 ( .A1(n27830), .A2(n27831), .ZN(n27829) );
  INV_X1 U27852 ( .A(n27832), .ZN(n27830) );
  AND2_X1 U27853 ( .A1(n27833), .A2(n27832), .ZN(n27828) );
  INV_X1 U27854 ( .A(n27831), .ZN(n27833) );
  AND2_X1 U27855 ( .A1(n27834), .A2(n27835), .ZN(n27435) );
  INV_X1 U27856 ( .A(n27836), .ZN(n27835) );
  AND2_X1 U27857 ( .A1(n27837), .A2(n27838), .ZN(n27836) );
  OR2_X1 U27858 ( .A1(n27838), .A2(n27837), .ZN(n27834) );
  OR2_X1 U27859 ( .A1(n27839), .A2(n27840), .ZN(n27837) );
  AND2_X1 U27860 ( .A1(n27841), .A2(n27842), .ZN(n27840) );
  INV_X1 U27861 ( .A(n27843), .ZN(n27841) );
  AND2_X1 U27862 ( .A1(n27844), .A2(n27843), .ZN(n27839) );
  INV_X1 U27863 ( .A(n27842), .ZN(n27844) );
  AND2_X1 U27864 ( .A1(n27845), .A2(n27846), .ZN(n27446) );
  INV_X1 U27865 ( .A(n27847), .ZN(n27846) );
  AND2_X1 U27866 ( .A1(n27848), .A2(n27849), .ZN(n27847) );
  OR2_X1 U27867 ( .A1(n27849), .A2(n27848), .ZN(n27845) );
  OR2_X1 U27868 ( .A1(n27850), .A2(n27851), .ZN(n27848) );
  AND2_X1 U27869 ( .A1(n27852), .A2(n27853), .ZN(n27851) );
  INV_X1 U27870 ( .A(n27854), .ZN(n27852) );
  AND2_X1 U27871 ( .A1(n27855), .A2(n27854), .ZN(n27850) );
  INV_X1 U27872 ( .A(n27853), .ZN(n27855) );
  AND2_X1 U27873 ( .A1(n27856), .A2(n27857), .ZN(n27457) );
  INV_X1 U27874 ( .A(n27858), .ZN(n27857) );
  AND2_X1 U27875 ( .A1(n27859), .A2(n27860), .ZN(n27858) );
  OR2_X1 U27876 ( .A1(n27860), .A2(n27859), .ZN(n27856) );
  OR2_X1 U27877 ( .A1(n27861), .A2(n27862), .ZN(n27859) );
  AND2_X1 U27878 ( .A1(n27863), .A2(n27864), .ZN(n27862) );
  INV_X1 U27879 ( .A(n27865), .ZN(n27863) );
  AND2_X1 U27880 ( .A1(n27866), .A2(n27865), .ZN(n27861) );
  INV_X1 U27881 ( .A(n27864), .ZN(n27866) );
  AND2_X1 U27882 ( .A1(n27867), .A2(n27868), .ZN(n27468) );
  INV_X1 U27883 ( .A(n27869), .ZN(n27868) );
  AND2_X1 U27884 ( .A1(n27870), .A2(n27871), .ZN(n27869) );
  OR2_X1 U27885 ( .A1(n27871), .A2(n27870), .ZN(n27867) );
  OR2_X1 U27886 ( .A1(n27872), .A2(n27873), .ZN(n27870) );
  AND2_X1 U27887 ( .A1(n27874), .A2(n27875), .ZN(n27873) );
  INV_X1 U27888 ( .A(n27876), .ZN(n27874) );
  AND2_X1 U27889 ( .A1(n27877), .A2(n27876), .ZN(n27872) );
  INV_X1 U27890 ( .A(n27875), .ZN(n27877) );
  AND2_X1 U27891 ( .A1(n27878), .A2(n27879), .ZN(n27479) );
  INV_X1 U27892 ( .A(n27880), .ZN(n27879) );
  AND2_X1 U27893 ( .A1(n27881), .A2(n27882), .ZN(n27880) );
  OR2_X1 U27894 ( .A1(n27882), .A2(n27881), .ZN(n27878) );
  OR2_X1 U27895 ( .A1(n27883), .A2(n27884), .ZN(n27881) );
  AND2_X1 U27896 ( .A1(n27885), .A2(n27886), .ZN(n27884) );
  INV_X1 U27897 ( .A(n27887), .ZN(n27885) );
  AND2_X1 U27898 ( .A1(n27888), .A2(n27887), .ZN(n27883) );
  INV_X1 U27899 ( .A(n27886), .ZN(n27888) );
  AND2_X1 U27900 ( .A1(n27889), .A2(n27890), .ZN(n27490) );
  INV_X1 U27901 ( .A(n27891), .ZN(n27890) );
  AND2_X1 U27902 ( .A1(n27892), .A2(n27893), .ZN(n27891) );
  OR2_X1 U27903 ( .A1(n27893), .A2(n27892), .ZN(n27889) );
  OR2_X1 U27904 ( .A1(n27894), .A2(n27895), .ZN(n27892) );
  AND2_X1 U27905 ( .A1(n27896), .A2(n27897), .ZN(n27895) );
  INV_X1 U27906 ( .A(n27898), .ZN(n27896) );
  AND2_X1 U27907 ( .A1(n27899), .A2(n27898), .ZN(n27894) );
  INV_X1 U27908 ( .A(n27897), .ZN(n27899) );
  AND2_X1 U27909 ( .A1(n27900), .A2(n27901), .ZN(n27501) );
  INV_X1 U27910 ( .A(n27902), .ZN(n27901) );
  AND2_X1 U27911 ( .A1(n27903), .A2(n27904), .ZN(n27902) );
  OR2_X1 U27912 ( .A1(n27904), .A2(n27903), .ZN(n27900) );
  OR2_X1 U27913 ( .A1(n27905), .A2(n27906), .ZN(n27903) );
  AND2_X1 U27914 ( .A1(n27907), .A2(n27908), .ZN(n27906) );
  INV_X1 U27915 ( .A(n27909), .ZN(n27907) );
  AND2_X1 U27916 ( .A1(n27910), .A2(n27909), .ZN(n27905) );
  INV_X1 U27917 ( .A(n27908), .ZN(n27910) );
  AND2_X1 U27918 ( .A1(n27911), .A2(n27912), .ZN(n27512) );
  INV_X1 U27919 ( .A(n27913), .ZN(n27912) );
  AND2_X1 U27920 ( .A1(n27914), .A2(n27915), .ZN(n27913) );
  OR2_X1 U27921 ( .A1(n27915), .A2(n27914), .ZN(n27911) );
  OR2_X1 U27922 ( .A1(n27916), .A2(n27917), .ZN(n27914) );
  AND2_X1 U27923 ( .A1(n27918), .A2(n27919), .ZN(n27917) );
  INV_X1 U27924 ( .A(n27920), .ZN(n27918) );
  AND2_X1 U27925 ( .A1(n27921), .A2(n27920), .ZN(n27916) );
  INV_X1 U27926 ( .A(n27919), .ZN(n27921) );
  AND2_X1 U27927 ( .A1(n27922), .A2(n27923), .ZN(n27523) );
  INV_X1 U27928 ( .A(n27924), .ZN(n27923) );
  AND2_X1 U27929 ( .A1(n27925), .A2(n27926), .ZN(n27924) );
  OR2_X1 U27930 ( .A1(n27926), .A2(n27925), .ZN(n27922) );
  OR2_X1 U27931 ( .A1(n27927), .A2(n27928), .ZN(n27925) );
  AND2_X1 U27932 ( .A1(n27929), .A2(n27930), .ZN(n27928) );
  INV_X1 U27933 ( .A(n27931), .ZN(n27929) );
  AND2_X1 U27934 ( .A1(n27932), .A2(n27931), .ZN(n27927) );
  INV_X1 U27935 ( .A(n27930), .ZN(n27932) );
  AND2_X1 U27936 ( .A1(n27933), .A2(n27934), .ZN(n27534) );
  INV_X1 U27937 ( .A(n27935), .ZN(n27934) );
  AND2_X1 U27938 ( .A1(n27936), .A2(n27937), .ZN(n27935) );
  OR2_X1 U27939 ( .A1(n27937), .A2(n27936), .ZN(n27933) );
  OR2_X1 U27940 ( .A1(n27938), .A2(n27939), .ZN(n27936) );
  AND2_X1 U27941 ( .A1(n27940), .A2(n27941), .ZN(n27939) );
  INV_X1 U27942 ( .A(n27942), .ZN(n27940) );
  AND2_X1 U27943 ( .A1(n27943), .A2(n27942), .ZN(n27938) );
  INV_X1 U27944 ( .A(n27941), .ZN(n27943) );
  AND2_X1 U27945 ( .A1(n27944), .A2(n27945), .ZN(n27545) );
  INV_X1 U27946 ( .A(n27946), .ZN(n27945) );
  AND2_X1 U27947 ( .A1(n27947), .A2(n27948), .ZN(n27946) );
  OR2_X1 U27948 ( .A1(n27948), .A2(n27947), .ZN(n27944) );
  OR2_X1 U27949 ( .A1(n27949), .A2(n27950), .ZN(n27947) );
  AND2_X1 U27950 ( .A1(n27951), .A2(n27952), .ZN(n27950) );
  INV_X1 U27951 ( .A(n27953), .ZN(n27951) );
  AND2_X1 U27952 ( .A1(n27954), .A2(n27953), .ZN(n27949) );
  INV_X1 U27953 ( .A(n27952), .ZN(n27954) );
  AND2_X1 U27954 ( .A1(n27955), .A2(n27956), .ZN(n27556) );
  INV_X1 U27955 ( .A(n27957), .ZN(n27956) );
  AND2_X1 U27956 ( .A1(n27958), .A2(n27959), .ZN(n27957) );
  OR2_X1 U27957 ( .A1(n27959), .A2(n27958), .ZN(n27955) );
  OR2_X1 U27958 ( .A1(n27960), .A2(n27961), .ZN(n27958) );
  AND2_X1 U27959 ( .A1(n27962), .A2(n27963), .ZN(n27961) );
  INV_X1 U27960 ( .A(n27964), .ZN(n27962) );
  AND2_X1 U27961 ( .A1(n27965), .A2(n27964), .ZN(n27960) );
  INV_X1 U27962 ( .A(n27963), .ZN(n27965) );
  AND2_X1 U27963 ( .A1(n27966), .A2(n27967), .ZN(n27567) );
  INV_X1 U27964 ( .A(n27968), .ZN(n27967) );
  AND2_X1 U27965 ( .A1(n27969), .A2(n27970), .ZN(n27968) );
  OR2_X1 U27966 ( .A1(n27970), .A2(n27969), .ZN(n27966) );
  OR2_X1 U27967 ( .A1(n27971), .A2(n27972), .ZN(n27969) );
  AND2_X1 U27968 ( .A1(n27973), .A2(n27974), .ZN(n27972) );
  INV_X1 U27969 ( .A(n27975), .ZN(n27973) );
  AND2_X1 U27970 ( .A1(n27976), .A2(n27975), .ZN(n27971) );
  INV_X1 U27971 ( .A(n27974), .ZN(n27976) );
  AND2_X1 U27972 ( .A1(n27977), .A2(n27978), .ZN(n27578) );
  INV_X1 U27973 ( .A(n27979), .ZN(n27978) );
  AND2_X1 U27974 ( .A1(n27980), .A2(n27981), .ZN(n27979) );
  OR2_X1 U27975 ( .A1(n27981), .A2(n27980), .ZN(n27977) );
  OR2_X1 U27976 ( .A1(n27982), .A2(n27983), .ZN(n27980) );
  AND2_X1 U27977 ( .A1(n27984), .A2(n27985), .ZN(n27983) );
  INV_X1 U27978 ( .A(n27986), .ZN(n27984) );
  AND2_X1 U27979 ( .A1(n27987), .A2(n27986), .ZN(n27982) );
  INV_X1 U27980 ( .A(n27985), .ZN(n27987) );
  AND2_X1 U27981 ( .A1(n27988), .A2(n27989), .ZN(n27589) );
  INV_X1 U27982 ( .A(n27990), .ZN(n27989) );
  AND2_X1 U27983 ( .A1(n27991), .A2(n27992), .ZN(n27990) );
  OR2_X1 U27984 ( .A1(n27992), .A2(n27991), .ZN(n27988) );
  OR2_X1 U27985 ( .A1(n27993), .A2(n27994), .ZN(n27991) );
  AND2_X1 U27986 ( .A1(n27995), .A2(n27996), .ZN(n27994) );
  INV_X1 U27987 ( .A(n27997), .ZN(n27995) );
  AND2_X1 U27988 ( .A1(n27998), .A2(n27997), .ZN(n27993) );
  INV_X1 U27989 ( .A(n27996), .ZN(n27998) );
  AND2_X1 U27990 ( .A1(n27999), .A2(n28000), .ZN(n27600) );
  INV_X1 U27991 ( .A(n28001), .ZN(n28000) );
  AND2_X1 U27992 ( .A1(n28002), .A2(n28003), .ZN(n28001) );
  OR2_X1 U27993 ( .A1(n28003), .A2(n28002), .ZN(n27999) );
  OR2_X1 U27994 ( .A1(n28004), .A2(n28005), .ZN(n28002) );
  AND2_X1 U27995 ( .A1(n28006), .A2(n28007), .ZN(n28005) );
  INV_X1 U27996 ( .A(n28008), .ZN(n28006) );
  AND2_X1 U27997 ( .A1(n28009), .A2(n28008), .ZN(n28004) );
  INV_X1 U27998 ( .A(n28007), .ZN(n28009) );
  AND2_X1 U27999 ( .A1(n28010), .A2(n28011), .ZN(n27610) );
  INV_X1 U28000 ( .A(n28012), .ZN(n28011) );
  AND2_X1 U28001 ( .A1(n28013), .A2(n28014), .ZN(n28012) );
  OR2_X1 U28002 ( .A1(n28014), .A2(n28013), .ZN(n28010) );
  OR2_X1 U28003 ( .A1(n28015), .A2(n28016), .ZN(n28013) );
  AND2_X1 U28004 ( .A1(n28017), .A2(n28018), .ZN(n28016) );
  INV_X1 U28005 ( .A(n28019), .ZN(n28017) );
  AND2_X1 U28006 ( .A1(n28020), .A2(n28019), .ZN(n28015) );
  INV_X1 U28007 ( .A(n28018), .ZN(n28020) );
  AND2_X1 U28008 ( .A1(n28021), .A2(n28022), .ZN(n27621) );
  INV_X1 U28009 ( .A(n28023), .ZN(n28022) );
  AND2_X1 U28010 ( .A1(n28024), .A2(n28025), .ZN(n28023) );
  OR2_X1 U28011 ( .A1(n28025), .A2(n28024), .ZN(n28021) );
  OR2_X1 U28012 ( .A1(n28026), .A2(n28027), .ZN(n28024) );
  AND2_X1 U28013 ( .A1(n28028), .A2(n28029), .ZN(n28027) );
  INV_X1 U28014 ( .A(n15879), .ZN(n28028) );
  AND2_X1 U28015 ( .A1(n28030), .A2(n15879), .ZN(n28026) );
  INV_X1 U28016 ( .A(n28029), .ZN(n28030) );
  AND2_X1 U28017 ( .A1(n28031), .A2(n28032), .ZN(n27632) );
  INV_X1 U28018 ( .A(n28033), .ZN(n28032) );
  AND2_X1 U28019 ( .A1(n28034), .A2(n28035), .ZN(n28033) );
  OR2_X1 U28020 ( .A1(n28035), .A2(n28034), .ZN(n28031) );
  OR2_X1 U28021 ( .A1(n28036), .A2(n28037), .ZN(n28034) );
  AND2_X1 U28022 ( .A1(n28038), .A2(n28039), .ZN(n28037) );
  INV_X1 U28023 ( .A(n28040), .ZN(n28038) );
  AND2_X1 U28024 ( .A1(n28041), .A2(n28040), .ZN(n28036) );
  INV_X1 U28025 ( .A(n28039), .ZN(n28041) );
  AND2_X1 U28026 ( .A1(n28042), .A2(n28043), .ZN(n27643) );
  INV_X1 U28027 ( .A(n28044), .ZN(n28043) );
  AND2_X1 U28028 ( .A1(n28045), .A2(n28046), .ZN(n28044) );
  OR2_X1 U28029 ( .A1(n28046), .A2(n28045), .ZN(n28042) );
  OR2_X1 U28030 ( .A1(n28047), .A2(n28048), .ZN(n28045) );
  AND2_X1 U28031 ( .A1(n28049), .A2(n28050), .ZN(n28048) );
  INV_X1 U28032 ( .A(n28051), .ZN(n28049) );
  AND2_X1 U28033 ( .A1(n28052), .A2(n28051), .ZN(n28047) );
  INV_X1 U28034 ( .A(n28050), .ZN(n28052) );
  AND2_X1 U28035 ( .A1(n28053), .A2(n28054), .ZN(n16437) );
  INV_X1 U28036 ( .A(n28055), .ZN(n28054) );
  AND2_X1 U28037 ( .A1(n28056), .A2(n28057), .ZN(n28055) );
  OR2_X1 U28038 ( .A1(n28057), .A2(n28056), .ZN(n28053) );
  OR2_X1 U28039 ( .A1(n28058), .A2(n28059), .ZN(n28056) );
  AND2_X1 U28040 ( .A1(n28060), .A2(n28061), .ZN(n28059) );
  INV_X1 U28041 ( .A(n28062), .ZN(n28060) );
  AND2_X1 U28042 ( .A1(n28063), .A2(n28062), .ZN(n28058) );
  INV_X1 U28043 ( .A(n28061), .ZN(n28063) );
  AND2_X1 U28044 ( .A1(n28064), .A2(n28065), .ZN(n16421) );
  INV_X1 U28045 ( .A(n28066), .ZN(n28065) );
  AND2_X1 U28046 ( .A1(n28067), .A2(n16406), .ZN(n28066) );
  OR2_X1 U28047 ( .A1(n16406), .A2(n28067), .ZN(n28064) );
  OR2_X1 U28048 ( .A1(n28068), .A2(n28069), .ZN(n28067) );
  AND2_X1 U28049 ( .A1(n28070), .A2(n16405), .ZN(n28069) );
  INV_X1 U28050 ( .A(n16404), .ZN(n28070) );
  AND2_X1 U28051 ( .A1(n28071), .A2(n16404), .ZN(n28068) );
  OR2_X1 U28052 ( .A1(n16512), .A2(n15739), .ZN(n16404) );
  INV_X1 U28053 ( .A(n16405), .ZN(n28071) );
  OR2_X1 U28054 ( .A1(n28072), .A2(n28073), .ZN(n16405) );
  AND2_X1 U28055 ( .A1(n28062), .A2(n28061), .ZN(n28073) );
  AND2_X1 U28056 ( .A1(n28057), .A2(n28074), .ZN(n28072) );
  OR2_X1 U28057 ( .A1(n28061), .A2(n28062), .ZN(n28074) );
  OR2_X1 U28058 ( .A1(n15842), .A2(n15739), .ZN(n28062) );
  OR2_X1 U28059 ( .A1(n28075), .A2(n28076), .ZN(n28061) );
  AND2_X1 U28060 ( .A1(n28051), .A2(n28050), .ZN(n28076) );
  AND2_X1 U28061 ( .A1(n28046), .A2(n28077), .ZN(n28075) );
  OR2_X1 U28062 ( .A1(n28050), .A2(n28051), .ZN(n28077) );
  OR2_X1 U28063 ( .A1(n15808), .A2(n15739), .ZN(n28051) );
  OR2_X1 U28064 ( .A1(n28078), .A2(n28079), .ZN(n28050) );
  AND2_X1 U28065 ( .A1(n28040), .A2(n28039), .ZN(n28079) );
  AND2_X1 U28066 ( .A1(n28035), .A2(n28080), .ZN(n28078) );
  OR2_X1 U28067 ( .A1(n28039), .A2(n28040), .ZN(n28080) );
  OR2_X1 U28068 ( .A1(n15774), .A2(n15739), .ZN(n28040) );
  OR2_X1 U28069 ( .A1(n28081), .A2(n28082), .ZN(n28039) );
  AND2_X1 U28070 ( .A1(n15879), .A2(n28029), .ZN(n28082) );
  AND2_X1 U28071 ( .A1(n28025), .A2(n28083), .ZN(n28081) );
  OR2_X1 U28072 ( .A1(n28029), .A2(n15879), .ZN(n28083) );
  OR2_X1 U28073 ( .A1(n15740), .A2(n15739), .ZN(n15879) );
  OR2_X1 U28074 ( .A1(n28084), .A2(n28085), .ZN(n28029) );
  AND2_X1 U28075 ( .A1(n28019), .A2(n28018), .ZN(n28085) );
  AND2_X1 U28076 ( .A1(n28014), .A2(n28086), .ZN(n28084) );
  OR2_X1 U28077 ( .A1(n28018), .A2(n28019), .ZN(n28086) );
  OR2_X1 U28078 ( .A1(n15706), .A2(n15739), .ZN(n28019) );
  OR2_X1 U28079 ( .A1(n28087), .A2(n28088), .ZN(n28018) );
  AND2_X1 U28080 ( .A1(n28008), .A2(n28007), .ZN(n28088) );
  AND2_X1 U28081 ( .A1(n28003), .A2(n28089), .ZN(n28087) );
  OR2_X1 U28082 ( .A1(n28007), .A2(n28008), .ZN(n28089) );
  OR2_X1 U28083 ( .A1(n15672), .A2(n15739), .ZN(n28008) );
  OR2_X1 U28084 ( .A1(n28090), .A2(n28091), .ZN(n28007) );
  AND2_X1 U28085 ( .A1(n27997), .A2(n27996), .ZN(n28091) );
  AND2_X1 U28086 ( .A1(n27992), .A2(n28092), .ZN(n28090) );
  OR2_X1 U28087 ( .A1(n27996), .A2(n27997), .ZN(n28092) );
  OR2_X1 U28088 ( .A1(n15638), .A2(n15739), .ZN(n27997) );
  OR2_X1 U28089 ( .A1(n28093), .A2(n28094), .ZN(n27996) );
  AND2_X1 U28090 ( .A1(n27986), .A2(n27985), .ZN(n28094) );
  AND2_X1 U28091 ( .A1(n27981), .A2(n28095), .ZN(n28093) );
  OR2_X1 U28092 ( .A1(n27985), .A2(n27986), .ZN(n28095) );
  OR2_X1 U28093 ( .A1(n15593), .A2(n15739), .ZN(n27986) );
  OR2_X1 U28094 ( .A1(n28096), .A2(n28097), .ZN(n27985) );
  AND2_X1 U28095 ( .A1(n27975), .A2(n27974), .ZN(n28097) );
  AND2_X1 U28096 ( .A1(n27970), .A2(n28098), .ZN(n28096) );
  OR2_X1 U28097 ( .A1(n27974), .A2(n27975), .ZN(n28098) );
  OR2_X1 U28098 ( .A1(n15559), .A2(n15739), .ZN(n27975) );
  OR2_X1 U28099 ( .A1(n28099), .A2(n28100), .ZN(n27974) );
  AND2_X1 U28100 ( .A1(n27964), .A2(n27963), .ZN(n28100) );
  AND2_X1 U28101 ( .A1(n27959), .A2(n28101), .ZN(n28099) );
  OR2_X1 U28102 ( .A1(n27963), .A2(n27964), .ZN(n28101) );
  OR2_X1 U28103 ( .A1(n15525), .A2(n15739), .ZN(n27964) );
  OR2_X1 U28104 ( .A1(n28102), .A2(n28103), .ZN(n27963) );
  AND2_X1 U28105 ( .A1(n27953), .A2(n27952), .ZN(n28103) );
  AND2_X1 U28106 ( .A1(n27948), .A2(n28104), .ZN(n28102) );
  OR2_X1 U28107 ( .A1(n27952), .A2(n27953), .ZN(n28104) );
  OR2_X1 U28108 ( .A1(n15491), .A2(n15739), .ZN(n27953) );
  OR2_X1 U28109 ( .A1(n28105), .A2(n28106), .ZN(n27952) );
  AND2_X1 U28110 ( .A1(n27942), .A2(n27941), .ZN(n28106) );
  AND2_X1 U28111 ( .A1(n27937), .A2(n28107), .ZN(n28105) );
  OR2_X1 U28112 ( .A1(n27941), .A2(n27942), .ZN(n28107) );
  OR2_X1 U28113 ( .A1(n15457), .A2(n15739), .ZN(n27942) );
  OR2_X1 U28114 ( .A1(n28108), .A2(n28109), .ZN(n27941) );
  AND2_X1 U28115 ( .A1(n27931), .A2(n27930), .ZN(n28109) );
  AND2_X1 U28116 ( .A1(n27926), .A2(n28110), .ZN(n28108) );
  OR2_X1 U28117 ( .A1(n27930), .A2(n27931), .ZN(n28110) );
  OR2_X1 U28118 ( .A1(n15423), .A2(n15739), .ZN(n27931) );
  OR2_X1 U28119 ( .A1(n28111), .A2(n28112), .ZN(n27930) );
  AND2_X1 U28120 ( .A1(n27920), .A2(n27919), .ZN(n28112) );
  AND2_X1 U28121 ( .A1(n27915), .A2(n28113), .ZN(n28111) );
  OR2_X1 U28122 ( .A1(n27919), .A2(n27920), .ZN(n28113) );
  OR2_X1 U28123 ( .A1(n15389), .A2(n15739), .ZN(n27920) );
  OR2_X1 U28124 ( .A1(n28114), .A2(n28115), .ZN(n27919) );
  AND2_X1 U28125 ( .A1(n27909), .A2(n27908), .ZN(n28115) );
  AND2_X1 U28126 ( .A1(n27904), .A2(n28116), .ZN(n28114) );
  OR2_X1 U28127 ( .A1(n27908), .A2(n27909), .ZN(n28116) );
  OR2_X1 U28128 ( .A1(n15355), .A2(n15739), .ZN(n27909) );
  OR2_X1 U28129 ( .A1(n28117), .A2(n28118), .ZN(n27908) );
  AND2_X1 U28130 ( .A1(n27898), .A2(n27897), .ZN(n28118) );
  AND2_X1 U28131 ( .A1(n27893), .A2(n28119), .ZN(n28117) );
  OR2_X1 U28132 ( .A1(n27897), .A2(n27898), .ZN(n28119) );
  OR2_X1 U28133 ( .A1(n15321), .A2(n15739), .ZN(n27898) );
  OR2_X1 U28134 ( .A1(n28120), .A2(n28121), .ZN(n27897) );
  AND2_X1 U28135 ( .A1(n27887), .A2(n27886), .ZN(n28121) );
  AND2_X1 U28136 ( .A1(n27882), .A2(n28122), .ZN(n28120) );
  OR2_X1 U28137 ( .A1(n27886), .A2(n27887), .ZN(n28122) );
  OR2_X1 U28138 ( .A1(n15287), .A2(n15739), .ZN(n27887) );
  OR2_X1 U28139 ( .A1(n28123), .A2(n28124), .ZN(n27886) );
  AND2_X1 U28140 ( .A1(n27876), .A2(n27875), .ZN(n28124) );
  AND2_X1 U28141 ( .A1(n27871), .A2(n28125), .ZN(n28123) );
  OR2_X1 U28142 ( .A1(n27875), .A2(n27876), .ZN(n28125) );
  OR2_X1 U28143 ( .A1(n15242), .A2(n15739), .ZN(n27876) );
  OR2_X1 U28144 ( .A1(n28126), .A2(n28127), .ZN(n27875) );
  AND2_X1 U28145 ( .A1(n27865), .A2(n27864), .ZN(n28127) );
  AND2_X1 U28146 ( .A1(n27860), .A2(n28128), .ZN(n28126) );
  OR2_X1 U28147 ( .A1(n27864), .A2(n27865), .ZN(n28128) );
  OR2_X1 U28148 ( .A1(n15208), .A2(n15739), .ZN(n27865) );
  OR2_X1 U28149 ( .A1(n28129), .A2(n28130), .ZN(n27864) );
  AND2_X1 U28150 ( .A1(n27854), .A2(n27853), .ZN(n28130) );
  AND2_X1 U28151 ( .A1(n27849), .A2(n28131), .ZN(n28129) );
  OR2_X1 U28152 ( .A1(n27853), .A2(n27854), .ZN(n28131) );
  OR2_X1 U28153 ( .A1(n15174), .A2(n15739), .ZN(n27854) );
  OR2_X1 U28154 ( .A1(n28132), .A2(n28133), .ZN(n27853) );
  AND2_X1 U28155 ( .A1(n27843), .A2(n27842), .ZN(n28133) );
  AND2_X1 U28156 ( .A1(n27838), .A2(n28134), .ZN(n28132) );
  OR2_X1 U28157 ( .A1(n27842), .A2(n27843), .ZN(n28134) );
  OR2_X1 U28158 ( .A1(n15140), .A2(n15739), .ZN(n27843) );
  OR2_X1 U28159 ( .A1(n28135), .A2(n28136), .ZN(n27842) );
  AND2_X1 U28160 ( .A1(n27832), .A2(n27831), .ZN(n28136) );
  AND2_X1 U28161 ( .A1(n27827), .A2(n28137), .ZN(n28135) );
  OR2_X1 U28162 ( .A1(n27831), .A2(n27832), .ZN(n28137) );
  OR2_X1 U28163 ( .A1(n15106), .A2(n15739), .ZN(n27832) );
  OR2_X1 U28164 ( .A1(n28138), .A2(n28139), .ZN(n27831) );
  AND2_X1 U28165 ( .A1(n27821), .A2(n27820), .ZN(n28139) );
  AND2_X1 U28166 ( .A1(n27816), .A2(n28140), .ZN(n28138) );
  OR2_X1 U28167 ( .A1(n27820), .A2(n27821), .ZN(n28140) );
  OR2_X1 U28168 ( .A1(n15072), .A2(n15739), .ZN(n27821) );
  OR2_X1 U28169 ( .A1(n28141), .A2(n28142), .ZN(n27820) );
  AND2_X1 U28170 ( .A1(n27810), .A2(n27809), .ZN(n28142) );
  AND2_X1 U28171 ( .A1(n27805), .A2(n28143), .ZN(n28141) );
  OR2_X1 U28172 ( .A1(n27809), .A2(n27810), .ZN(n28143) );
  OR2_X1 U28173 ( .A1(n15038), .A2(n15739), .ZN(n27810) );
  OR2_X1 U28174 ( .A1(n28144), .A2(n28145), .ZN(n27809) );
  AND2_X1 U28175 ( .A1(n27794), .A2(n27800), .ZN(n28145) );
  AND2_X1 U28176 ( .A1(n28146), .A2(n27799), .ZN(n28144) );
  OR2_X1 U28177 ( .A1(n28147), .A2(n28148), .ZN(n27799) );
  AND2_X1 U28178 ( .A1(n27786), .A2(n27788), .ZN(n28148) );
  AND2_X1 U28179 ( .A1(n27783), .A2(n28149), .ZN(n28147) );
  OR2_X1 U28180 ( .A1(n27788), .A2(n27786), .ZN(n28149) );
  OR2_X1 U28181 ( .A1(n14970), .A2(n15739), .ZN(n27786) );
  OR2_X1 U28182 ( .A1(n28150), .A2(n28151), .ZN(n27788) );
  AND2_X1 U28183 ( .A1(n27772), .A2(n27775), .ZN(n28151) );
  AND2_X1 U28184 ( .A1(n28152), .A2(n27777), .ZN(n28150) );
  OR2_X1 U28185 ( .A1(n28153), .A2(n28154), .ZN(n27777) );
  AND2_X1 U28186 ( .A1(n27761), .A2(n27764), .ZN(n28154) );
  AND2_X1 U28187 ( .A1(n28155), .A2(n27766), .ZN(n28153) );
  OR2_X1 U28188 ( .A1(n28156), .A2(n28157), .ZN(n27766) );
  AND2_X1 U28189 ( .A1(n27749), .A2(n27754), .ZN(n28157) );
  AND2_X1 U28190 ( .A1(n27753), .A2(n28158), .ZN(n28156) );
  OR2_X1 U28191 ( .A1(n27754), .A2(n27749), .ZN(n28158) );
  OR2_X1 U28192 ( .A1(n14857), .A2(n15739), .ZN(n27749) );
  INV_X1 U28193 ( .A(n27755), .ZN(n27754) );
  AND3_X1 U28194 ( .A1(b_4_), .A2(b_3_), .A3(n15957), .ZN(n27755) );
  INV_X1 U28195 ( .A(n27756), .ZN(n27753) );
  OR2_X1 U28196 ( .A1(n28159), .A2(n28160), .ZN(n27756) );
  AND2_X1 U28197 ( .A1(b_3_), .A2(n28161), .ZN(n28160) );
  OR2_X1 U28198 ( .A1(n28162), .A2(n16981), .ZN(n28161) );
  AND2_X1 U28199 ( .A1(a_30_), .A2(n15807), .ZN(n28162) );
  AND2_X1 U28200 ( .A1(b_2_), .A2(n28163), .ZN(n28159) );
  OR2_X1 U28201 ( .A1(n28164), .A2(n14817), .ZN(n28163) );
  AND2_X1 U28202 ( .A1(a_31_), .A2(n15773), .ZN(n28164) );
  OR2_X1 U28203 ( .A1(n27764), .A2(n27761), .ZN(n28155) );
  OR2_X1 U28204 ( .A1(n28165), .A2(n28166), .ZN(n27761) );
  AND2_X1 U28205 ( .A1(n28167), .A2(n28168), .ZN(n28166) );
  INV_X1 U28206 ( .A(n28169), .ZN(n28165) );
  OR2_X1 U28207 ( .A1(n28167), .A2(n28168), .ZN(n28169) );
  OR2_X1 U28208 ( .A1(n28170), .A2(n28171), .ZN(n28167) );
  AND2_X1 U28209 ( .A1(n28172), .A2(n28173), .ZN(n28171) );
  AND2_X1 U28210 ( .A1(n28174), .A2(n28175), .ZN(n28170) );
  OR2_X1 U28211 ( .A1(n14891), .A2(n15739), .ZN(n27764) );
  OR2_X1 U28212 ( .A1(n27775), .A2(n27772), .ZN(n28152) );
  OR2_X1 U28213 ( .A1(n28176), .A2(n28177), .ZN(n27772) );
  INV_X1 U28214 ( .A(n28178), .ZN(n28177) );
  OR2_X1 U28215 ( .A1(n28179), .A2(n28180), .ZN(n28178) );
  AND2_X1 U28216 ( .A1(n28180), .A2(n28179), .ZN(n28176) );
  AND2_X1 U28217 ( .A1(n28181), .A2(n28182), .ZN(n28179) );
  OR2_X1 U28218 ( .A1(n28183), .A2(n28184), .ZN(n28182) );
  INV_X1 U28219 ( .A(n28185), .ZN(n28184) );
  OR2_X1 U28220 ( .A1(n28185), .A2(n28186), .ZN(n28181) );
  INV_X1 U28221 ( .A(n28183), .ZN(n28186) );
  OR2_X1 U28222 ( .A1(n14936), .A2(n15739), .ZN(n27775) );
  OR2_X1 U28223 ( .A1(n28187), .A2(n28188), .ZN(n27783) );
  INV_X1 U28224 ( .A(n28189), .ZN(n28188) );
  OR2_X1 U28225 ( .A1(n28190), .A2(n28191), .ZN(n28189) );
  AND2_X1 U28226 ( .A1(n28191), .A2(n28190), .ZN(n28187) );
  AND2_X1 U28227 ( .A1(n28192), .A2(n28193), .ZN(n28190) );
  OR2_X1 U28228 ( .A1(n28194), .A2(n28195), .ZN(n28193) );
  INV_X1 U28229 ( .A(n28196), .ZN(n28195) );
  OR2_X1 U28230 ( .A1(n28196), .A2(n28197), .ZN(n28192) );
  INV_X1 U28231 ( .A(n28194), .ZN(n28197) );
  OR2_X1 U28232 ( .A1(n27800), .A2(n27794), .ZN(n28146) );
  OR2_X1 U28233 ( .A1(n28198), .A2(n28199), .ZN(n27794) );
  INV_X1 U28234 ( .A(n28200), .ZN(n28199) );
  OR2_X1 U28235 ( .A1(n28201), .A2(n28202), .ZN(n28200) );
  AND2_X1 U28236 ( .A1(n28202), .A2(n28201), .ZN(n28198) );
  AND2_X1 U28237 ( .A1(n28203), .A2(n28204), .ZN(n28201) );
  INV_X1 U28238 ( .A(n28205), .ZN(n28204) );
  AND2_X1 U28239 ( .A1(n28206), .A2(n28207), .ZN(n28205) );
  OR2_X1 U28240 ( .A1(n28207), .A2(n28206), .ZN(n28203) );
  INV_X1 U28241 ( .A(n28208), .ZN(n28206) );
  OR2_X1 U28242 ( .A1(n15004), .A2(n15739), .ZN(n27800) );
  INV_X1 U28243 ( .A(b_4_), .ZN(n15739) );
  AND2_X1 U28244 ( .A1(n28209), .A2(n28210), .ZN(n27805) );
  INV_X1 U28245 ( .A(n28211), .ZN(n28210) );
  AND2_X1 U28246 ( .A1(n28212), .A2(n28213), .ZN(n28211) );
  OR2_X1 U28247 ( .A1(n28213), .A2(n28212), .ZN(n28209) );
  OR2_X1 U28248 ( .A1(n28214), .A2(n28215), .ZN(n28212) );
  AND2_X1 U28249 ( .A1(n28216), .A2(n28217), .ZN(n28215) );
  INV_X1 U28250 ( .A(n28218), .ZN(n28216) );
  AND2_X1 U28251 ( .A1(n28219), .A2(n28218), .ZN(n28214) );
  INV_X1 U28252 ( .A(n28217), .ZN(n28219) );
  AND2_X1 U28253 ( .A1(n28220), .A2(n28221), .ZN(n27816) );
  INV_X1 U28254 ( .A(n28222), .ZN(n28221) );
  AND2_X1 U28255 ( .A1(n28223), .A2(n28224), .ZN(n28222) );
  OR2_X1 U28256 ( .A1(n28224), .A2(n28223), .ZN(n28220) );
  OR2_X1 U28257 ( .A1(n28225), .A2(n28226), .ZN(n28223) );
  AND2_X1 U28258 ( .A1(n28227), .A2(n28228), .ZN(n28226) );
  INV_X1 U28259 ( .A(n28229), .ZN(n28227) );
  AND2_X1 U28260 ( .A1(n28230), .A2(n28229), .ZN(n28225) );
  INV_X1 U28261 ( .A(n28228), .ZN(n28230) );
  AND2_X1 U28262 ( .A1(n28231), .A2(n28232), .ZN(n27827) );
  INV_X1 U28263 ( .A(n28233), .ZN(n28232) );
  AND2_X1 U28264 ( .A1(n28234), .A2(n28235), .ZN(n28233) );
  OR2_X1 U28265 ( .A1(n28235), .A2(n28234), .ZN(n28231) );
  OR2_X1 U28266 ( .A1(n28236), .A2(n28237), .ZN(n28234) );
  AND2_X1 U28267 ( .A1(n28238), .A2(n28239), .ZN(n28237) );
  INV_X1 U28268 ( .A(n28240), .ZN(n28238) );
  AND2_X1 U28269 ( .A1(n28241), .A2(n28240), .ZN(n28236) );
  INV_X1 U28270 ( .A(n28239), .ZN(n28241) );
  AND2_X1 U28271 ( .A1(n28242), .A2(n28243), .ZN(n27838) );
  INV_X1 U28272 ( .A(n28244), .ZN(n28243) );
  AND2_X1 U28273 ( .A1(n28245), .A2(n28246), .ZN(n28244) );
  OR2_X1 U28274 ( .A1(n28246), .A2(n28245), .ZN(n28242) );
  OR2_X1 U28275 ( .A1(n28247), .A2(n28248), .ZN(n28245) );
  AND2_X1 U28276 ( .A1(n28249), .A2(n28250), .ZN(n28248) );
  INV_X1 U28277 ( .A(n28251), .ZN(n28249) );
  AND2_X1 U28278 ( .A1(n28252), .A2(n28251), .ZN(n28247) );
  INV_X1 U28279 ( .A(n28250), .ZN(n28252) );
  AND2_X1 U28280 ( .A1(n28253), .A2(n28254), .ZN(n27849) );
  INV_X1 U28281 ( .A(n28255), .ZN(n28254) );
  AND2_X1 U28282 ( .A1(n28256), .A2(n28257), .ZN(n28255) );
  OR2_X1 U28283 ( .A1(n28257), .A2(n28256), .ZN(n28253) );
  OR2_X1 U28284 ( .A1(n28258), .A2(n28259), .ZN(n28256) );
  AND2_X1 U28285 ( .A1(n28260), .A2(n28261), .ZN(n28259) );
  INV_X1 U28286 ( .A(n28262), .ZN(n28260) );
  AND2_X1 U28287 ( .A1(n28263), .A2(n28262), .ZN(n28258) );
  INV_X1 U28288 ( .A(n28261), .ZN(n28263) );
  AND2_X1 U28289 ( .A1(n28264), .A2(n28265), .ZN(n27860) );
  INV_X1 U28290 ( .A(n28266), .ZN(n28265) );
  AND2_X1 U28291 ( .A1(n28267), .A2(n28268), .ZN(n28266) );
  OR2_X1 U28292 ( .A1(n28268), .A2(n28267), .ZN(n28264) );
  OR2_X1 U28293 ( .A1(n28269), .A2(n28270), .ZN(n28267) );
  AND2_X1 U28294 ( .A1(n28271), .A2(n28272), .ZN(n28270) );
  INV_X1 U28295 ( .A(n28273), .ZN(n28271) );
  AND2_X1 U28296 ( .A1(n28274), .A2(n28273), .ZN(n28269) );
  INV_X1 U28297 ( .A(n28272), .ZN(n28274) );
  AND2_X1 U28298 ( .A1(n28275), .A2(n28276), .ZN(n27871) );
  INV_X1 U28299 ( .A(n28277), .ZN(n28276) );
  AND2_X1 U28300 ( .A1(n28278), .A2(n28279), .ZN(n28277) );
  OR2_X1 U28301 ( .A1(n28279), .A2(n28278), .ZN(n28275) );
  OR2_X1 U28302 ( .A1(n28280), .A2(n28281), .ZN(n28278) );
  AND2_X1 U28303 ( .A1(n28282), .A2(n28283), .ZN(n28281) );
  INV_X1 U28304 ( .A(n28284), .ZN(n28282) );
  AND2_X1 U28305 ( .A1(n28285), .A2(n28284), .ZN(n28280) );
  INV_X1 U28306 ( .A(n28283), .ZN(n28285) );
  AND2_X1 U28307 ( .A1(n28286), .A2(n28287), .ZN(n27882) );
  INV_X1 U28308 ( .A(n28288), .ZN(n28287) );
  AND2_X1 U28309 ( .A1(n28289), .A2(n28290), .ZN(n28288) );
  OR2_X1 U28310 ( .A1(n28290), .A2(n28289), .ZN(n28286) );
  OR2_X1 U28311 ( .A1(n28291), .A2(n28292), .ZN(n28289) );
  AND2_X1 U28312 ( .A1(n28293), .A2(n28294), .ZN(n28292) );
  INV_X1 U28313 ( .A(n28295), .ZN(n28293) );
  AND2_X1 U28314 ( .A1(n28296), .A2(n28295), .ZN(n28291) );
  INV_X1 U28315 ( .A(n28294), .ZN(n28296) );
  AND2_X1 U28316 ( .A1(n28297), .A2(n28298), .ZN(n27893) );
  INV_X1 U28317 ( .A(n28299), .ZN(n28298) );
  AND2_X1 U28318 ( .A1(n28300), .A2(n28301), .ZN(n28299) );
  OR2_X1 U28319 ( .A1(n28301), .A2(n28300), .ZN(n28297) );
  OR2_X1 U28320 ( .A1(n28302), .A2(n28303), .ZN(n28300) );
  AND2_X1 U28321 ( .A1(n28304), .A2(n28305), .ZN(n28303) );
  INV_X1 U28322 ( .A(n28306), .ZN(n28304) );
  AND2_X1 U28323 ( .A1(n28307), .A2(n28306), .ZN(n28302) );
  INV_X1 U28324 ( .A(n28305), .ZN(n28307) );
  AND2_X1 U28325 ( .A1(n28308), .A2(n28309), .ZN(n27904) );
  INV_X1 U28326 ( .A(n28310), .ZN(n28309) );
  AND2_X1 U28327 ( .A1(n28311), .A2(n28312), .ZN(n28310) );
  OR2_X1 U28328 ( .A1(n28312), .A2(n28311), .ZN(n28308) );
  OR2_X1 U28329 ( .A1(n28313), .A2(n28314), .ZN(n28311) );
  AND2_X1 U28330 ( .A1(n28315), .A2(n28316), .ZN(n28314) );
  INV_X1 U28331 ( .A(n28317), .ZN(n28315) );
  AND2_X1 U28332 ( .A1(n28318), .A2(n28317), .ZN(n28313) );
  INV_X1 U28333 ( .A(n28316), .ZN(n28318) );
  AND2_X1 U28334 ( .A1(n28319), .A2(n28320), .ZN(n27915) );
  INV_X1 U28335 ( .A(n28321), .ZN(n28320) );
  AND2_X1 U28336 ( .A1(n28322), .A2(n28323), .ZN(n28321) );
  OR2_X1 U28337 ( .A1(n28323), .A2(n28322), .ZN(n28319) );
  OR2_X1 U28338 ( .A1(n28324), .A2(n28325), .ZN(n28322) );
  AND2_X1 U28339 ( .A1(n28326), .A2(n28327), .ZN(n28325) );
  INV_X1 U28340 ( .A(n28328), .ZN(n28326) );
  AND2_X1 U28341 ( .A1(n28329), .A2(n28328), .ZN(n28324) );
  INV_X1 U28342 ( .A(n28327), .ZN(n28329) );
  AND2_X1 U28343 ( .A1(n28330), .A2(n28331), .ZN(n27926) );
  INV_X1 U28344 ( .A(n28332), .ZN(n28331) );
  AND2_X1 U28345 ( .A1(n28333), .A2(n28334), .ZN(n28332) );
  OR2_X1 U28346 ( .A1(n28334), .A2(n28333), .ZN(n28330) );
  OR2_X1 U28347 ( .A1(n28335), .A2(n28336), .ZN(n28333) );
  AND2_X1 U28348 ( .A1(n28337), .A2(n28338), .ZN(n28336) );
  INV_X1 U28349 ( .A(n28339), .ZN(n28337) );
  AND2_X1 U28350 ( .A1(n28340), .A2(n28339), .ZN(n28335) );
  INV_X1 U28351 ( .A(n28338), .ZN(n28340) );
  AND2_X1 U28352 ( .A1(n28341), .A2(n28342), .ZN(n27937) );
  INV_X1 U28353 ( .A(n28343), .ZN(n28342) );
  AND2_X1 U28354 ( .A1(n28344), .A2(n28345), .ZN(n28343) );
  OR2_X1 U28355 ( .A1(n28345), .A2(n28344), .ZN(n28341) );
  OR2_X1 U28356 ( .A1(n28346), .A2(n28347), .ZN(n28344) );
  AND2_X1 U28357 ( .A1(n28348), .A2(n28349), .ZN(n28347) );
  INV_X1 U28358 ( .A(n28350), .ZN(n28348) );
  AND2_X1 U28359 ( .A1(n28351), .A2(n28350), .ZN(n28346) );
  INV_X1 U28360 ( .A(n28349), .ZN(n28351) );
  AND2_X1 U28361 ( .A1(n28352), .A2(n28353), .ZN(n27948) );
  INV_X1 U28362 ( .A(n28354), .ZN(n28353) );
  AND2_X1 U28363 ( .A1(n28355), .A2(n28356), .ZN(n28354) );
  OR2_X1 U28364 ( .A1(n28356), .A2(n28355), .ZN(n28352) );
  OR2_X1 U28365 ( .A1(n28357), .A2(n28358), .ZN(n28355) );
  AND2_X1 U28366 ( .A1(n28359), .A2(n28360), .ZN(n28358) );
  INV_X1 U28367 ( .A(n28361), .ZN(n28359) );
  AND2_X1 U28368 ( .A1(n28362), .A2(n28361), .ZN(n28357) );
  INV_X1 U28369 ( .A(n28360), .ZN(n28362) );
  AND2_X1 U28370 ( .A1(n28363), .A2(n28364), .ZN(n27959) );
  INV_X1 U28371 ( .A(n28365), .ZN(n28364) );
  AND2_X1 U28372 ( .A1(n28366), .A2(n28367), .ZN(n28365) );
  OR2_X1 U28373 ( .A1(n28367), .A2(n28366), .ZN(n28363) );
  OR2_X1 U28374 ( .A1(n28368), .A2(n28369), .ZN(n28366) );
  AND2_X1 U28375 ( .A1(n28370), .A2(n28371), .ZN(n28369) );
  INV_X1 U28376 ( .A(n28372), .ZN(n28370) );
  AND2_X1 U28377 ( .A1(n28373), .A2(n28372), .ZN(n28368) );
  INV_X1 U28378 ( .A(n28371), .ZN(n28373) );
  AND2_X1 U28379 ( .A1(n28374), .A2(n28375), .ZN(n27970) );
  INV_X1 U28380 ( .A(n28376), .ZN(n28375) );
  AND2_X1 U28381 ( .A1(n28377), .A2(n28378), .ZN(n28376) );
  OR2_X1 U28382 ( .A1(n28378), .A2(n28377), .ZN(n28374) );
  OR2_X1 U28383 ( .A1(n28379), .A2(n28380), .ZN(n28377) );
  AND2_X1 U28384 ( .A1(n28381), .A2(n28382), .ZN(n28380) );
  INV_X1 U28385 ( .A(n28383), .ZN(n28381) );
  AND2_X1 U28386 ( .A1(n28384), .A2(n28383), .ZN(n28379) );
  INV_X1 U28387 ( .A(n28382), .ZN(n28384) );
  AND2_X1 U28388 ( .A1(n28385), .A2(n28386), .ZN(n27981) );
  INV_X1 U28389 ( .A(n28387), .ZN(n28386) );
  AND2_X1 U28390 ( .A1(n28388), .A2(n28389), .ZN(n28387) );
  OR2_X1 U28391 ( .A1(n28389), .A2(n28388), .ZN(n28385) );
  OR2_X1 U28392 ( .A1(n28390), .A2(n28391), .ZN(n28388) );
  AND2_X1 U28393 ( .A1(n28392), .A2(n28393), .ZN(n28391) );
  INV_X1 U28394 ( .A(n28394), .ZN(n28392) );
  AND2_X1 U28395 ( .A1(n28395), .A2(n28394), .ZN(n28390) );
  INV_X1 U28396 ( .A(n28393), .ZN(n28395) );
  AND2_X1 U28397 ( .A1(n28396), .A2(n28397), .ZN(n27992) );
  INV_X1 U28398 ( .A(n28398), .ZN(n28397) );
  AND2_X1 U28399 ( .A1(n28399), .A2(n28400), .ZN(n28398) );
  OR2_X1 U28400 ( .A1(n28400), .A2(n28399), .ZN(n28396) );
  OR2_X1 U28401 ( .A1(n28401), .A2(n28402), .ZN(n28399) );
  AND2_X1 U28402 ( .A1(n28403), .A2(n28404), .ZN(n28402) );
  INV_X1 U28403 ( .A(n28405), .ZN(n28403) );
  AND2_X1 U28404 ( .A1(n28406), .A2(n28405), .ZN(n28401) );
  INV_X1 U28405 ( .A(n28404), .ZN(n28406) );
  AND2_X1 U28406 ( .A1(n28407), .A2(n28408), .ZN(n28003) );
  INV_X1 U28407 ( .A(n28409), .ZN(n28408) );
  AND2_X1 U28408 ( .A1(n28410), .A2(n28411), .ZN(n28409) );
  OR2_X1 U28409 ( .A1(n28411), .A2(n28410), .ZN(n28407) );
  OR2_X1 U28410 ( .A1(n28412), .A2(n28413), .ZN(n28410) );
  AND2_X1 U28411 ( .A1(n28414), .A2(n28415), .ZN(n28413) );
  INV_X1 U28412 ( .A(n28416), .ZN(n28414) );
  AND2_X1 U28413 ( .A1(n28417), .A2(n28416), .ZN(n28412) );
  INV_X1 U28414 ( .A(n28415), .ZN(n28417) );
  AND2_X1 U28415 ( .A1(n28418), .A2(n28419), .ZN(n28014) );
  INV_X1 U28416 ( .A(n28420), .ZN(n28419) );
  AND2_X1 U28417 ( .A1(n28421), .A2(n28422), .ZN(n28420) );
  OR2_X1 U28418 ( .A1(n28422), .A2(n28421), .ZN(n28418) );
  OR2_X1 U28419 ( .A1(n28423), .A2(n28424), .ZN(n28421) );
  AND2_X1 U28420 ( .A1(n28425), .A2(n28426), .ZN(n28424) );
  INV_X1 U28421 ( .A(n28427), .ZN(n28425) );
  AND2_X1 U28422 ( .A1(n28428), .A2(n28427), .ZN(n28423) );
  INV_X1 U28423 ( .A(n28426), .ZN(n28428) );
  AND2_X1 U28424 ( .A1(n28429), .A2(n28430), .ZN(n28025) );
  INV_X1 U28425 ( .A(n28431), .ZN(n28430) );
  AND2_X1 U28426 ( .A1(n28432), .A2(n28433), .ZN(n28431) );
  OR2_X1 U28427 ( .A1(n28433), .A2(n28432), .ZN(n28429) );
  OR2_X1 U28428 ( .A1(n28434), .A2(n28435), .ZN(n28432) );
  AND2_X1 U28429 ( .A1(n28436), .A2(n28437), .ZN(n28435) );
  INV_X1 U28430 ( .A(n28438), .ZN(n28436) );
  AND2_X1 U28431 ( .A1(n28439), .A2(n28438), .ZN(n28434) );
  INV_X1 U28432 ( .A(n28437), .ZN(n28439) );
  AND2_X1 U28433 ( .A1(n28440), .A2(n28441), .ZN(n28035) );
  INV_X1 U28434 ( .A(n28442), .ZN(n28441) );
  AND2_X1 U28435 ( .A1(n28443), .A2(n28444), .ZN(n28442) );
  OR2_X1 U28436 ( .A1(n28444), .A2(n28443), .ZN(n28440) );
  OR2_X1 U28437 ( .A1(n28445), .A2(n28446), .ZN(n28443) );
  AND2_X1 U28438 ( .A1(n28447), .A2(n28448), .ZN(n28446) );
  INV_X1 U28439 ( .A(n28449), .ZN(n28447) );
  AND2_X1 U28440 ( .A1(n28450), .A2(n28449), .ZN(n28445) );
  INV_X1 U28441 ( .A(n28448), .ZN(n28450) );
  AND2_X1 U28442 ( .A1(n28451), .A2(n28452), .ZN(n28046) );
  INV_X1 U28443 ( .A(n28453), .ZN(n28452) );
  AND2_X1 U28444 ( .A1(n28454), .A2(n28455), .ZN(n28453) );
  OR2_X1 U28445 ( .A1(n28455), .A2(n28454), .ZN(n28451) );
  OR2_X1 U28446 ( .A1(n28456), .A2(n28457), .ZN(n28454) );
  AND2_X1 U28447 ( .A1(n28458), .A2(n28459), .ZN(n28457) );
  INV_X1 U28448 ( .A(n15876), .ZN(n28458) );
  AND2_X1 U28449 ( .A1(n28460), .A2(n15876), .ZN(n28456) );
  INV_X1 U28450 ( .A(n28459), .ZN(n28460) );
  AND2_X1 U28451 ( .A1(n28461), .A2(n28462), .ZN(n28057) );
  INV_X1 U28452 ( .A(n28463), .ZN(n28462) );
  AND2_X1 U28453 ( .A1(n28464), .A2(n28465), .ZN(n28463) );
  OR2_X1 U28454 ( .A1(n28465), .A2(n28464), .ZN(n28461) );
  OR2_X1 U28455 ( .A1(n28466), .A2(n28467), .ZN(n28464) );
  AND2_X1 U28456 ( .A1(n28468), .A2(n28469), .ZN(n28467) );
  INV_X1 U28457 ( .A(n28470), .ZN(n28468) );
  AND2_X1 U28458 ( .A1(n28471), .A2(n28470), .ZN(n28466) );
  INV_X1 U28459 ( .A(n28469), .ZN(n28471) );
  AND2_X1 U28460 ( .A1(n28472), .A2(n28473), .ZN(n16406) );
  INV_X1 U28461 ( .A(n28474), .ZN(n28473) );
  AND2_X1 U28462 ( .A1(n28475), .A2(n28476), .ZN(n28474) );
  OR2_X1 U28463 ( .A1(n28476), .A2(n28475), .ZN(n28472) );
  OR2_X1 U28464 ( .A1(n28477), .A2(n28478), .ZN(n28475) );
  AND2_X1 U28465 ( .A1(n28479), .A2(n28480), .ZN(n28478) );
  INV_X1 U28466 ( .A(n28481), .ZN(n28479) );
  AND2_X1 U28467 ( .A1(n28482), .A2(n28481), .ZN(n28477) );
  INV_X1 U28468 ( .A(n28480), .ZN(n28482) );
  OR2_X1 U28469 ( .A1(n16396), .A2(n16397), .ZN(n15991) );
  OR2_X1 U28470 ( .A1(n28483), .A2(n28484), .ZN(n16397) );
  AND2_X1 U28471 ( .A1(n16417), .A2(n16416), .ZN(n28484) );
  AND2_X1 U28472 ( .A1(n16412), .A2(n28485), .ZN(n28483) );
  OR2_X1 U28473 ( .A1(n16416), .A2(n16417), .ZN(n28485) );
  OR2_X1 U28474 ( .A1(n16512), .A2(n15773), .ZN(n16417) );
  OR2_X1 U28475 ( .A1(n28486), .A2(n28487), .ZN(n16416) );
  AND2_X1 U28476 ( .A1(n28481), .A2(n28480), .ZN(n28487) );
  AND2_X1 U28477 ( .A1(n28476), .A2(n28488), .ZN(n28486) );
  OR2_X1 U28478 ( .A1(n28480), .A2(n28481), .ZN(n28488) );
  OR2_X1 U28479 ( .A1(n15842), .A2(n15773), .ZN(n28481) );
  OR2_X1 U28480 ( .A1(n28489), .A2(n28490), .ZN(n28480) );
  AND2_X1 U28481 ( .A1(n28470), .A2(n28469), .ZN(n28490) );
  AND2_X1 U28482 ( .A1(n28465), .A2(n28491), .ZN(n28489) );
  OR2_X1 U28483 ( .A1(n28469), .A2(n28470), .ZN(n28491) );
  OR2_X1 U28484 ( .A1(n15808), .A2(n15773), .ZN(n28470) );
  OR2_X1 U28485 ( .A1(n28492), .A2(n28493), .ZN(n28469) );
  AND2_X1 U28486 ( .A1(n15876), .A2(n28459), .ZN(n28493) );
  AND2_X1 U28487 ( .A1(n28455), .A2(n28494), .ZN(n28492) );
  OR2_X1 U28488 ( .A1(n28459), .A2(n15876), .ZN(n28494) );
  OR2_X1 U28489 ( .A1(n15774), .A2(n15773), .ZN(n15876) );
  OR2_X1 U28490 ( .A1(n28495), .A2(n28496), .ZN(n28459) );
  AND2_X1 U28491 ( .A1(n28449), .A2(n28448), .ZN(n28496) );
  AND2_X1 U28492 ( .A1(n28444), .A2(n28497), .ZN(n28495) );
  OR2_X1 U28493 ( .A1(n28448), .A2(n28449), .ZN(n28497) );
  OR2_X1 U28494 ( .A1(n15740), .A2(n15773), .ZN(n28449) );
  OR2_X1 U28495 ( .A1(n28498), .A2(n28499), .ZN(n28448) );
  AND2_X1 U28496 ( .A1(n28438), .A2(n28437), .ZN(n28499) );
  AND2_X1 U28497 ( .A1(n28433), .A2(n28500), .ZN(n28498) );
  OR2_X1 U28498 ( .A1(n28437), .A2(n28438), .ZN(n28500) );
  OR2_X1 U28499 ( .A1(n15706), .A2(n15773), .ZN(n28438) );
  OR2_X1 U28500 ( .A1(n28501), .A2(n28502), .ZN(n28437) );
  AND2_X1 U28501 ( .A1(n28427), .A2(n28426), .ZN(n28502) );
  AND2_X1 U28502 ( .A1(n28422), .A2(n28503), .ZN(n28501) );
  OR2_X1 U28503 ( .A1(n28426), .A2(n28427), .ZN(n28503) );
  OR2_X1 U28504 ( .A1(n15672), .A2(n15773), .ZN(n28427) );
  OR2_X1 U28505 ( .A1(n28504), .A2(n28505), .ZN(n28426) );
  AND2_X1 U28506 ( .A1(n28416), .A2(n28415), .ZN(n28505) );
  AND2_X1 U28507 ( .A1(n28411), .A2(n28506), .ZN(n28504) );
  OR2_X1 U28508 ( .A1(n28415), .A2(n28416), .ZN(n28506) );
  OR2_X1 U28509 ( .A1(n15638), .A2(n15773), .ZN(n28416) );
  OR2_X1 U28510 ( .A1(n28507), .A2(n28508), .ZN(n28415) );
  AND2_X1 U28511 ( .A1(n28405), .A2(n28404), .ZN(n28508) );
  AND2_X1 U28512 ( .A1(n28400), .A2(n28509), .ZN(n28507) );
  OR2_X1 U28513 ( .A1(n28404), .A2(n28405), .ZN(n28509) );
  OR2_X1 U28514 ( .A1(n15593), .A2(n15773), .ZN(n28405) );
  OR2_X1 U28515 ( .A1(n28510), .A2(n28511), .ZN(n28404) );
  AND2_X1 U28516 ( .A1(n28394), .A2(n28393), .ZN(n28511) );
  AND2_X1 U28517 ( .A1(n28389), .A2(n28512), .ZN(n28510) );
  OR2_X1 U28518 ( .A1(n28393), .A2(n28394), .ZN(n28512) );
  OR2_X1 U28519 ( .A1(n15559), .A2(n15773), .ZN(n28394) );
  OR2_X1 U28520 ( .A1(n28513), .A2(n28514), .ZN(n28393) );
  AND2_X1 U28521 ( .A1(n28383), .A2(n28382), .ZN(n28514) );
  AND2_X1 U28522 ( .A1(n28378), .A2(n28515), .ZN(n28513) );
  OR2_X1 U28523 ( .A1(n28382), .A2(n28383), .ZN(n28515) );
  OR2_X1 U28524 ( .A1(n15525), .A2(n15773), .ZN(n28383) );
  OR2_X1 U28525 ( .A1(n28516), .A2(n28517), .ZN(n28382) );
  AND2_X1 U28526 ( .A1(n28372), .A2(n28371), .ZN(n28517) );
  AND2_X1 U28527 ( .A1(n28367), .A2(n28518), .ZN(n28516) );
  OR2_X1 U28528 ( .A1(n28371), .A2(n28372), .ZN(n28518) );
  OR2_X1 U28529 ( .A1(n15491), .A2(n15773), .ZN(n28372) );
  OR2_X1 U28530 ( .A1(n28519), .A2(n28520), .ZN(n28371) );
  AND2_X1 U28531 ( .A1(n28361), .A2(n28360), .ZN(n28520) );
  AND2_X1 U28532 ( .A1(n28356), .A2(n28521), .ZN(n28519) );
  OR2_X1 U28533 ( .A1(n28360), .A2(n28361), .ZN(n28521) );
  OR2_X1 U28534 ( .A1(n15457), .A2(n15773), .ZN(n28361) );
  OR2_X1 U28535 ( .A1(n28522), .A2(n28523), .ZN(n28360) );
  AND2_X1 U28536 ( .A1(n28350), .A2(n28349), .ZN(n28523) );
  AND2_X1 U28537 ( .A1(n28345), .A2(n28524), .ZN(n28522) );
  OR2_X1 U28538 ( .A1(n28349), .A2(n28350), .ZN(n28524) );
  OR2_X1 U28539 ( .A1(n15423), .A2(n15773), .ZN(n28350) );
  OR2_X1 U28540 ( .A1(n28525), .A2(n28526), .ZN(n28349) );
  AND2_X1 U28541 ( .A1(n28339), .A2(n28338), .ZN(n28526) );
  AND2_X1 U28542 ( .A1(n28334), .A2(n28527), .ZN(n28525) );
  OR2_X1 U28543 ( .A1(n28338), .A2(n28339), .ZN(n28527) );
  OR2_X1 U28544 ( .A1(n15389), .A2(n15773), .ZN(n28339) );
  OR2_X1 U28545 ( .A1(n28528), .A2(n28529), .ZN(n28338) );
  AND2_X1 U28546 ( .A1(n28328), .A2(n28327), .ZN(n28529) );
  AND2_X1 U28547 ( .A1(n28323), .A2(n28530), .ZN(n28528) );
  OR2_X1 U28548 ( .A1(n28327), .A2(n28328), .ZN(n28530) );
  OR2_X1 U28549 ( .A1(n15355), .A2(n15773), .ZN(n28328) );
  OR2_X1 U28550 ( .A1(n28531), .A2(n28532), .ZN(n28327) );
  AND2_X1 U28551 ( .A1(n28317), .A2(n28316), .ZN(n28532) );
  AND2_X1 U28552 ( .A1(n28312), .A2(n28533), .ZN(n28531) );
  OR2_X1 U28553 ( .A1(n28316), .A2(n28317), .ZN(n28533) );
  OR2_X1 U28554 ( .A1(n15321), .A2(n15773), .ZN(n28317) );
  OR2_X1 U28555 ( .A1(n28534), .A2(n28535), .ZN(n28316) );
  AND2_X1 U28556 ( .A1(n28306), .A2(n28305), .ZN(n28535) );
  AND2_X1 U28557 ( .A1(n28301), .A2(n28536), .ZN(n28534) );
  OR2_X1 U28558 ( .A1(n28305), .A2(n28306), .ZN(n28536) );
  OR2_X1 U28559 ( .A1(n15287), .A2(n15773), .ZN(n28306) );
  OR2_X1 U28560 ( .A1(n28537), .A2(n28538), .ZN(n28305) );
  AND2_X1 U28561 ( .A1(n28295), .A2(n28294), .ZN(n28538) );
  AND2_X1 U28562 ( .A1(n28290), .A2(n28539), .ZN(n28537) );
  OR2_X1 U28563 ( .A1(n28294), .A2(n28295), .ZN(n28539) );
  OR2_X1 U28564 ( .A1(n15242), .A2(n15773), .ZN(n28295) );
  OR2_X1 U28565 ( .A1(n28540), .A2(n28541), .ZN(n28294) );
  AND2_X1 U28566 ( .A1(n28284), .A2(n28283), .ZN(n28541) );
  AND2_X1 U28567 ( .A1(n28279), .A2(n28542), .ZN(n28540) );
  OR2_X1 U28568 ( .A1(n28283), .A2(n28284), .ZN(n28542) );
  OR2_X1 U28569 ( .A1(n15208), .A2(n15773), .ZN(n28284) );
  OR2_X1 U28570 ( .A1(n28543), .A2(n28544), .ZN(n28283) );
  AND2_X1 U28571 ( .A1(n28273), .A2(n28272), .ZN(n28544) );
  AND2_X1 U28572 ( .A1(n28268), .A2(n28545), .ZN(n28543) );
  OR2_X1 U28573 ( .A1(n28272), .A2(n28273), .ZN(n28545) );
  OR2_X1 U28574 ( .A1(n15174), .A2(n15773), .ZN(n28273) );
  OR2_X1 U28575 ( .A1(n28546), .A2(n28547), .ZN(n28272) );
  AND2_X1 U28576 ( .A1(n28262), .A2(n28261), .ZN(n28547) );
  AND2_X1 U28577 ( .A1(n28257), .A2(n28548), .ZN(n28546) );
  OR2_X1 U28578 ( .A1(n28261), .A2(n28262), .ZN(n28548) );
  OR2_X1 U28579 ( .A1(n15140), .A2(n15773), .ZN(n28262) );
  OR2_X1 U28580 ( .A1(n28549), .A2(n28550), .ZN(n28261) );
  AND2_X1 U28581 ( .A1(n28251), .A2(n28250), .ZN(n28550) );
  AND2_X1 U28582 ( .A1(n28246), .A2(n28551), .ZN(n28549) );
  OR2_X1 U28583 ( .A1(n28250), .A2(n28251), .ZN(n28551) );
  OR2_X1 U28584 ( .A1(n15106), .A2(n15773), .ZN(n28251) );
  OR2_X1 U28585 ( .A1(n28552), .A2(n28553), .ZN(n28250) );
  AND2_X1 U28586 ( .A1(n28240), .A2(n28239), .ZN(n28553) );
  AND2_X1 U28587 ( .A1(n28235), .A2(n28554), .ZN(n28552) );
  OR2_X1 U28588 ( .A1(n28239), .A2(n28240), .ZN(n28554) );
  OR2_X1 U28589 ( .A1(n15072), .A2(n15773), .ZN(n28240) );
  OR2_X1 U28590 ( .A1(n28555), .A2(n28556), .ZN(n28239) );
  AND2_X1 U28591 ( .A1(n28229), .A2(n28228), .ZN(n28556) );
  AND2_X1 U28592 ( .A1(n28224), .A2(n28557), .ZN(n28555) );
  OR2_X1 U28593 ( .A1(n28228), .A2(n28229), .ZN(n28557) );
  OR2_X1 U28594 ( .A1(n15038), .A2(n15773), .ZN(n28229) );
  OR2_X1 U28595 ( .A1(n28558), .A2(n28559), .ZN(n28228) );
  AND2_X1 U28596 ( .A1(n28218), .A2(n28217), .ZN(n28559) );
  AND2_X1 U28597 ( .A1(n28213), .A2(n28560), .ZN(n28558) );
  OR2_X1 U28598 ( .A1(n28217), .A2(n28218), .ZN(n28560) );
  OR2_X1 U28599 ( .A1(n15004), .A2(n15773), .ZN(n28218) );
  OR2_X1 U28600 ( .A1(n28561), .A2(n28562), .ZN(n28217) );
  AND2_X1 U28601 ( .A1(n28202), .A2(n28208), .ZN(n28562) );
  AND2_X1 U28602 ( .A1(n28563), .A2(n28207), .ZN(n28561) );
  OR2_X1 U28603 ( .A1(n28564), .A2(n28565), .ZN(n28207) );
  AND2_X1 U28604 ( .A1(n28194), .A2(n28196), .ZN(n28565) );
  AND2_X1 U28605 ( .A1(n28191), .A2(n28566), .ZN(n28564) );
  OR2_X1 U28606 ( .A1(n28196), .A2(n28194), .ZN(n28566) );
  OR2_X1 U28607 ( .A1(n14936), .A2(n15773), .ZN(n28194) );
  OR2_X1 U28608 ( .A1(n28567), .A2(n28568), .ZN(n28196) );
  AND2_X1 U28609 ( .A1(n28180), .A2(n28183), .ZN(n28568) );
  AND2_X1 U28610 ( .A1(n28569), .A2(n28185), .ZN(n28567) );
  OR2_X1 U28611 ( .A1(n28570), .A2(n28571), .ZN(n28185) );
  AND2_X1 U28612 ( .A1(n28168), .A2(n28173), .ZN(n28571) );
  AND2_X1 U28613 ( .A1(n28172), .A2(n28572), .ZN(n28570) );
  OR2_X1 U28614 ( .A1(n28173), .A2(n28168), .ZN(n28572) );
  OR2_X1 U28615 ( .A1(n14857), .A2(n15773), .ZN(n28168) );
  INV_X1 U28616 ( .A(n28174), .ZN(n28173) );
  AND3_X1 U28617 ( .A1(b_3_), .A2(b_2_), .A3(n15957), .ZN(n28174) );
  INV_X1 U28618 ( .A(n28175), .ZN(n28172) );
  OR2_X1 U28619 ( .A1(n28573), .A2(n28574), .ZN(n28175) );
  AND2_X1 U28620 ( .A1(b_2_), .A2(n28575), .ZN(n28574) );
  OR2_X1 U28621 ( .A1(n28576), .A2(n16981), .ZN(n28575) );
  AND2_X1 U28622 ( .A1(a_30_), .A2(n15841), .ZN(n28576) );
  AND2_X1 U28623 ( .A1(b_1_), .A2(n28577), .ZN(n28573) );
  OR2_X1 U28624 ( .A1(n28578), .A2(n14817), .ZN(n28577) );
  AND2_X1 U28625 ( .A1(a_31_), .A2(n15807), .ZN(n28578) );
  OR2_X1 U28626 ( .A1(n28183), .A2(n28180), .ZN(n28569) );
  OR2_X1 U28627 ( .A1(n28579), .A2(n28580), .ZN(n28180) );
  AND2_X1 U28628 ( .A1(n28581), .A2(n28582), .ZN(n28580) );
  INV_X1 U28629 ( .A(n28583), .ZN(n28579) );
  OR2_X1 U28630 ( .A1(n28581), .A2(n28582), .ZN(n28583) );
  OR2_X1 U28631 ( .A1(n28584), .A2(n28585), .ZN(n28581) );
  AND2_X1 U28632 ( .A1(n28586), .A2(n28587), .ZN(n28585) );
  AND2_X1 U28633 ( .A1(n28588), .A2(n28589), .ZN(n28584) );
  OR2_X1 U28634 ( .A1(n14891), .A2(n15773), .ZN(n28183) );
  OR2_X1 U28635 ( .A1(n28590), .A2(n28591), .ZN(n28191) );
  INV_X1 U28636 ( .A(n28592), .ZN(n28591) );
  OR2_X1 U28637 ( .A1(n28593), .A2(n28594), .ZN(n28592) );
  AND2_X1 U28638 ( .A1(n28594), .A2(n28593), .ZN(n28590) );
  AND2_X1 U28639 ( .A1(n28595), .A2(n28596), .ZN(n28593) );
  OR2_X1 U28640 ( .A1(n28597), .A2(n28598), .ZN(n28596) );
  INV_X1 U28641 ( .A(n28599), .ZN(n28598) );
  OR2_X1 U28642 ( .A1(n28599), .A2(n28600), .ZN(n28595) );
  INV_X1 U28643 ( .A(n28597), .ZN(n28600) );
  OR2_X1 U28644 ( .A1(n28208), .A2(n28202), .ZN(n28563) );
  OR2_X1 U28645 ( .A1(n28601), .A2(n28602), .ZN(n28202) );
  INV_X1 U28646 ( .A(n28603), .ZN(n28602) );
  OR2_X1 U28647 ( .A1(n28604), .A2(n28605), .ZN(n28603) );
  AND2_X1 U28648 ( .A1(n28605), .A2(n28604), .ZN(n28601) );
  AND2_X1 U28649 ( .A1(n28606), .A2(n28607), .ZN(n28604) );
  INV_X1 U28650 ( .A(n28608), .ZN(n28607) );
  AND2_X1 U28651 ( .A1(n28609), .A2(n28610), .ZN(n28608) );
  OR2_X1 U28652 ( .A1(n28610), .A2(n28609), .ZN(n28606) );
  INV_X1 U28653 ( .A(n28611), .ZN(n28609) );
  OR2_X1 U28654 ( .A1(n14970), .A2(n15773), .ZN(n28208) );
  INV_X1 U28655 ( .A(b_3_), .ZN(n15773) );
  AND2_X1 U28656 ( .A1(n28612), .A2(n28613), .ZN(n28213) );
  INV_X1 U28657 ( .A(n28614), .ZN(n28613) );
  AND2_X1 U28658 ( .A1(n28615), .A2(n28616), .ZN(n28614) );
  OR2_X1 U28659 ( .A1(n28616), .A2(n28615), .ZN(n28612) );
  OR2_X1 U28660 ( .A1(n28617), .A2(n28618), .ZN(n28615) );
  AND2_X1 U28661 ( .A1(n28619), .A2(n28620), .ZN(n28618) );
  INV_X1 U28662 ( .A(n28621), .ZN(n28619) );
  AND2_X1 U28663 ( .A1(n28622), .A2(n28621), .ZN(n28617) );
  INV_X1 U28664 ( .A(n28620), .ZN(n28622) );
  AND2_X1 U28665 ( .A1(n28623), .A2(n28624), .ZN(n28224) );
  INV_X1 U28666 ( .A(n28625), .ZN(n28624) );
  AND2_X1 U28667 ( .A1(n28626), .A2(n28627), .ZN(n28625) );
  OR2_X1 U28668 ( .A1(n28627), .A2(n28626), .ZN(n28623) );
  OR2_X1 U28669 ( .A1(n28628), .A2(n28629), .ZN(n28626) );
  AND2_X1 U28670 ( .A1(n28630), .A2(n28631), .ZN(n28629) );
  INV_X1 U28671 ( .A(n28632), .ZN(n28630) );
  AND2_X1 U28672 ( .A1(n28633), .A2(n28632), .ZN(n28628) );
  INV_X1 U28673 ( .A(n28631), .ZN(n28633) );
  AND2_X1 U28674 ( .A1(n28634), .A2(n28635), .ZN(n28235) );
  INV_X1 U28675 ( .A(n28636), .ZN(n28635) );
  AND2_X1 U28676 ( .A1(n28637), .A2(n28638), .ZN(n28636) );
  OR2_X1 U28677 ( .A1(n28638), .A2(n28637), .ZN(n28634) );
  OR2_X1 U28678 ( .A1(n28639), .A2(n28640), .ZN(n28637) );
  AND2_X1 U28679 ( .A1(n28641), .A2(n28642), .ZN(n28640) );
  INV_X1 U28680 ( .A(n28643), .ZN(n28641) );
  AND2_X1 U28681 ( .A1(n28644), .A2(n28643), .ZN(n28639) );
  INV_X1 U28682 ( .A(n28642), .ZN(n28644) );
  AND2_X1 U28683 ( .A1(n28645), .A2(n28646), .ZN(n28246) );
  INV_X1 U28684 ( .A(n28647), .ZN(n28646) );
  AND2_X1 U28685 ( .A1(n28648), .A2(n28649), .ZN(n28647) );
  OR2_X1 U28686 ( .A1(n28649), .A2(n28648), .ZN(n28645) );
  OR2_X1 U28687 ( .A1(n28650), .A2(n28651), .ZN(n28648) );
  AND2_X1 U28688 ( .A1(n28652), .A2(n28653), .ZN(n28651) );
  INV_X1 U28689 ( .A(n28654), .ZN(n28652) );
  AND2_X1 U28690 ( .A1(n28655), .A2(n28654), .ZN(n28650) );
  INV_X1 U28691 ( .A(n28653), .ZN(n28655) );
  AND2_X1 U28692 ( .A1(n28656), .A2(n28657), .ZN(n28257) );
  INV_X1 U28693 ( .A(n28658), .ZN(n28657) );
  AND2_X1 U28694 ( .A1(n28659), .A2(n28660), .ZN(n28658) );
  OR2_X1 U28695 ( .A1(n28660), .A2(n28659), .ZN(n28656) );
  OR2_X1 U28696 ( .A1(n28661), .A2(n28662), .ZN(n28659) );
  AND2_X1 U28697 ( .A1(n28663), .A2(n28664), .ZN(n28662) );
  INV_X1 U28698 ( .A(n28665), .ZN(n28663) );
  AND2_X1 U28699 ( .A1(n28666), .A2(n28665), .ZN(n28661) );
  INV_X1 U28700 ( .A(n28664), .ZN(n28666) );
  AND2_X1 U28701 ( .A1(n28667), .A2(n28668), .ZN(n28268) );
  INV_X1 U28702 ( .A(n28669), .ZN(n28668) );
  AND2_X1 U28703 ( .A1(n28670), .A2(n28671), .ZN(n28669) );
  OR2_X1 U28704 ( .A1(n28671), .A2(n28670), .ZN(n28667) );
  OR2_X1 U28705 ( .A1(n28672), .A2(n28673), .ZN(n28670) );
  AND2_X1 U28706 ( .A1(n28674), .A2(n28675), .ZN(n28673) );
  INV_X1 U28707 ( .A(n28676), .ZN(n28674) );
  AND2_X1 U28708 ( .A1(n28677), .A2(n28676), .ZN(n28672) );
  INV_X1 U28709 ( .A(n28675), .ZN(n28677) );
  AND2_X1 U28710 ( .A1(n28678), .A2(n28679), .ZN(n28279) );
  INV_X1 U28711 ( .A(n28680), .ZN(n28679) );
  AND2_X1 U28712 ( .A1(n28681), .A2(n28682), .ZN(n28680) );
  OR2_X1 U28713 ( .A1(n28682), .A2(n28681), .ZN(n28678) );
  OR2_X1 U28714 ( .A1(n28683), .A2(n28684), .ZN(n28681) );
  AND2_X1 U28715 ( .A1(n28685), .A2(n28686), .ZN(n28684) );
  INV_X1 U28716 ( .A(n28687), .ZN(n28685) );
  AND2_X1 U28717 ( .A1(n28688), .A2(n28687), .ZN(n28683) );
  INV_X1 U28718 ( .A(n28686), .ZN(n28688) );
  AND2_X1 U28719 ( .A1(n28689), .A2(n28690), .ZN(n28290) );
  INV_X1 U28720 ( .A(n28691), .ZN(n28690) );
  AND2_X1 U28721 ( .A1(n28692), .A2(n28693), .ZN(n28691) );
  OR2_X1 U28722 ( .A1(n28693), .A2(n28692), .ZN(n28689) );
  OR2_X1 U28723 ( .A1(n28694), .A2(n28695), .ZN(n28692) );
  AND2_X1 U28724 ( .A1(n28696), .A2(n28697), .ZN(n28695) );
  INV_X1 U28725 ( .A(n28698), .ZN(n28696) );
  AND2_X1 U28726 ( .A1(n28699), .A2(n28698), .ZN(n28694) );
  INV_X1 U28727 ( .A(n28697), .ZN(n28699) );
  AND2_X1 U28728 ( .A1(n28700), .A2(n28701), .ZN(n28301) );
  INV_X1 U28729 ( .A(n28702), .ZN(n28701) );
  AND2_X1 U28730 ( .A1(n28703), .A2(n28704), .ZN(n28702) );
  OR2_X1 U28731 ( .A1(n28704), .A2(n28703), .ZN(n28700) );
  OR2_X1 U28732 ( .A1(n28705), .A2(n28706), .ZN(n28703) );
  AND2_X1 U28733 ( .A1(n28707), .A2(n28708), .ZN(n28706) );
  INV_X1 U28734 ( .A(n28709), .ZN(n28707) );
  AND2_X1 U28735 ( .A1(n28710), .A2(n28709), .ZN(n28705) );
  INV_X1 U28736 ( .A(n28708), .ZN(n28710) );
  AND2_X1 U28737 ( .A1(n28711), .A2(n28712), .ZN(n28312) );
  INV_X1 U28738 ( .A(n28713), .ZN(n28712) );
  AND2_X1 U28739 ( .A1(n28714), .A2(n28715), .ZN(n28713) );
  OR2_X1 U28740 ( .A1(n28715), .A2(n28714), .ZN(n28711) );
  OR2_X1 U28741 ( .A1(n28716), .A2(n28717), .ZN(n28714) );
  AND2_X1 U28742 ( .A1(n28718), .A2(n28719), .ZN(n28717) );
  INV_X1 U28743 ( .A(n28720), .ZN(n28718) );
  AND2_X1 U28744 ( .A1(n28721), .A2(n28720), .ZN(n28716) );
  INV_X1 U28745 ( .A(n28719), .ZN(n28721) );
  AND2_X1 U28746 ( .A1(n28722), .A2(n28723), .ZN(n28323) );
  INV_X1 U28747 ( .A(n28724), .ZN(n28723) );
  AND2_X1 U28748 ( .A1(n28725), .A2(n28726), .ZN(n28724) );
  OR2_X1 U28749 ( .A1(n28726), .A2(n28725), .ZN(n28722) );
  OR2_X1 U28750 ( .A1(n28727), .A2(n28728), .ZN(n28725) );
  AND2_X1 U28751 ( .A1(n28729), .A2(n28730), .ZN(n28728) );
  INV_X1 U28752 ( .A(n28731), .ZN(n28729) );
  AND2_X1 U28753 ( .A1(n28732), .A2(n28731), .ZN(n28727) );
  INV_X1 U28754 ( .A(n28730), .ZN(n28732) );
  AND2_X1 U28755 ( .A1(n28733), .A2(n28734), .ZN(n28334) );
  INV_X1 U28756 ( .A(n28735), .ZN(n28734) );
  AND2_X1 U28757 ( .A1(n28736), .A2(n28737), .ZN(n28735) );
  OR2_X1 U28758 ( .A1(n28737), .A2(n28736), .ZN(n28733) );
  OR2_X1 U28759 ( .A1(n28738), .A2(n28739), .ZN(n28736) );
  AND2_X1 U28760 ( .A1(n28740), .A2(n28741), .ZN(n28739) );
  INV_X1 U28761 ( .A(n28742), .ZN(n28740) );
  AND2_X1 U28762 ( .A1(n28743), .A2(n28742), .ZN(n28738) );
  INV_X1 U28763 ( .A(n28741), .ZN(n28743) );
  AND2_X1 U28764 ( .A1(n28744), .A2(n28745), .ZN(n28345) );
  INV_X1 U28765 ( .A(n28746), .ZN(n28745) );
  AND2_X1 U28766 ( .A1(n28747), .A2(n28748), .ZN(n28746) );
  OR2_X1 U28767 ( .A1(n28748), .A2(n28747), .ZN(n28744) );
  OR2_X1 U28768 ( .A1(n28749), .A2(n28750), .ZN(n28747) );
  AND2_X1 U28769 ( .A1(n28751), .A2(n28752), .ZN(n28750) );
  INV_X1 U28770 ( .A(n28753), .ZN(n28751) );
  AND2_X1 U28771 ( .A1(n28754), .A2(n28753), .ZN(n28749) );
  INV_X1 U28772 ( .A(n28752), .ZN(n28754) );
  AND2_X1 U28773 ( .A1(n28755), .A2(n28756), .ZN(n28356) );
  INV_X1 U28774 ( .A(n28757), .ZN(n28756) );
  AND2_X1 U28775 ( .A1(n28758), .A2(n28759), .ZN(n28757) );
  OR2_X1 U28776 ( .A1(n28759), .A2(n28758), .ZN(n28755) );
  OR2_X1 U28777 ( .A1(n28760), .A2(n28761), .ZN(n28758) );
  AND2_X1 U28778 ( .A1(n28762), .A2(n28763), .ZN(n28761) );
  INV_X1 U28779 ( .A(n28764), .ZN(n28762) );
  AND2_X1 U28780 ( .A1(n28765), .A2(n28764), .ZN(n28760) );
  INV_X1 U28781 ( .A(n28763), .ZN(n28765) );
  AND2_X1 U28782 ( .A1(n28766), .A2(n28767), .ZN(n28367) );
  INV_X1 U28783 ( .A(n28768), .ZN(n28767) );
  AND2_X1 U28784 ( .A1(n28769), .A2(n28770), .ZN(n28768) );
  OR2_X1 U28785 ( .A1(n28770), .A2(n28769), .ZN(n28766) );
  OR2_X1 U28786 ( .A1(n28771), .A2(n28772), .ZN(n28769) );
  AND2_X1 U28787 ( .A1(n28773), .A2(n28774), .ZN(n28772) );
  INV_X1 U28788 ( .A(n28775), .ZN(n28773) );
  AND2_X1 U28789 ( .A1(n28776), .A2(n28775), .ZN(n28771) );
  INV_X1 U28790 ( .A(n28774), .ZN(n28776) );
  AND2_X1 U28791 ( .A1(n28777), .A2(n28778), .ZN(n28378) );
  INV_X1 U28792 ( .A(n28779), .ZN(n28778) );
  AND2_X1 U28793 ( .A1(n28780), .A2(n28781), .ZN(n28779) );
  OR2_X1 U28794 ( .A1(n28781), .A2(n28780), .ZN(n28777) );
  OR2_X1 U28795 ( .A1(n28782), .A2(n28783), .ZN(n28780) );
  AND2_X1 U28796 ( .A1(n28784), .A2(n28785), .ZN(n28783) );
  INV_X1 U28797 ( .A(n28786), .ZN(n28784) );
  AND2_X1 U28798 ( .A1(n28787), .A2(n28786), .ZN(n28782) );
  INV_X1 U28799 ( .A(n28785), .ZN(n28787) );
  AND2_X1 U28800 ( .A1(n28788), .A2(n28789), .ZN(n28389) );
  INV_X1 U28801 ( .A(n28790), .ZN(n28789) );
  AND2_X1 U28802 ( .A1(n28791), .A2(n28792), .ZN(n28790) );
  OR2_X1 U28803 ( .A1(n28792), .A2(n28791), .ZN(n28788) );
  OR2_X1 U28804 ( .A1(n28793), .A2(n28794), .ZN(n28791) );
  AND2_X1 U28805 ( .A1(n28795), .A2(n28796), .ZN(n28794) );
  INV_X1 U28806 ( .A(n28797), .ZN(n28795) );
  AND2_X1 U28807 ( .A1(n28798), .A2(n28797), .ZN(n28793) );
  INV_X1 U28808 ( .A(n28796), .ZN(n28798) );
  AND2_X1 U28809 ( .A1(n28799), .A2(n28800), .ZN(n28400) );
  INV_X1 U28810 ( .A(n28801), .ZN(n28800) );
  AND2_X1 U28811 ( .A1(n28802), .A2(n28803), .ZN(n28801) );
  OR2_X1 U28812 ( .A1(n28803), .A2(n28802), .ZN(n28799) );
  OR2_X1 U28813 ( .A1(n28804), .A2(n28805), .ZN(n28802) );
  AND2_X1 U28814 ( .A1(n28806), .A2(n28807), .ZN(n28805) );
  INV_X1 U28815 ( .A(n28808), .ZN(n28806) );
  AND2_X1 U28816 ( .A1(n28809), .A2(n28808), .ZN(n28804) );
  INV_X1 U28817 ( .A(n28807), .ZN(n28809) );
  AND2_X1 U28818 ( .A1(n28810), .A2(n28811), .ZN(n28411) );
  INV_X1 U28819 ( .A(n28812), .ZN(n28811) );
  AND2_X1 U28820 ( .A1(n28813), .A2(n28814), .ZN(n28812) );
  OR2_X1 U28821 ( .A1(n28814), .A2(n28813), .ZN(n28810) );
  OR2_X1 U28822 ( .A1(n28815), .A2(n28816), .ZN(n28813) );
  AND2_X1 U28823 ( .A1(n28817), .A2(n28818), .ZN(n28816) );
  INV_X1 U28824 ( .A(n28819), .ZN(n28817) );
  AND2_X1 U28825 ( .A1(n28820), .A2(n28819), .ZN(n28815) );
  INV_X1 U28826 ( .A(n28818), .ZN(n28820) );
  AND2_X1 U28827 ( .A1(n28821), .A2(n28822), .ZN(n28422) );
  INV_X1 U28828 ( .A(n28823), .ZN(n28822) );
  AND2_X1 U28829 ( .A1(n28824), .A2(n28825), .ZN(n28823) );
  OR2_X1 U28830 ( .A1(n28825), .A2(n28824), .ZN(n28821) );
  OR2_X1 U28831 ( .A1(n28826), .A2(n28827), .ZN(n28824) );
  AND2_X1 U28832 ( .A1(n28828), .A2(n28829), .ZN(n28827) );
  INV_X1 U28833 ( .A(n28830), .ZN(n28828) );
  AND2_X1 U28834 ( .A1(n28831), .A2(n28830), .ZN(n28826) );
  INV_X1 U28835 ( .A(n28829), .ZN(n28831) );
  AND2_X1 U28836 ( .A1(n28832), .A2(n28833), .ZN(n28433) );
  INV_X1 U28837 ( .A(n28834), .ZN(n28833) );
  AND2_X1 U28838 ( .A1(n28835), .A2(n28836), .ZN(n28834) );
  OR2_X1 U28839 ( .A1(n28836), .A2(n28835), .ZN(n28832) );
  OR2_X1 U28840 ( .A1(n28837), .A2(n28838), .ZN(n28835) );
  AND2_X1 U28841 ( .A1(n28839), .A2(n28840), .ZN(n28838) );
  INV_X1 U28842 ( .A(n28841), .ZN(n28839) );
  AND2_X1 U28843 ( .A1(n28842), .A2(n28841), .ZN(n28837) );
  INV_X1 U28844 ( .A(n28840), .ZN(n28842) );
  AND2_X1 U28845 ( .A1(n28843), .A2(n28844), .ZN(n28444) );
  INV_X1 U28846 ( .A(n28845), .ZN(n28844) );
  AND2_X1 U28847 ( .A1(n28846), .A2(n28847), .ZN(n28845) );
  OR2_X1 U28848 ( .A1(n28847), .A2(n28846), .ZN(n28843) );
  OR2_X1 U28849 ( .A1(n28848), .A2(n28849), .ZN(n28846) );
  AND2_X1 U28850 ( .A1(n28850), .A2(n28851), .ZN(n28849) );
  INV_X1 U28851 ( .A(n28852), .ZN(n28850) );
  AND2_X1 U28852 ( .A1(n28853), .A2(n28852), .ZN(n28848) );
  INV_X1 U28853 ( .A(n28851), .ZN(n28853) );
  AND2_X1 U28854 ( .A1(n28854), .A2(n28855), .ZN(n28455) );
  INV_X1 U28855 ( .A(n28856), .ZN(n28855) );
  AND2_X1 U28856 ( .A1(n28857), .A2(n28858), .ZN(n28856) );
  OR2_X1 U28857 ( .A1(n28858), .A2(n28857), .ZN(n28854) );
  OR2_X1 U28858 ( .A1(n28859), .A2(n28860), .ZN(n28857) );
  AND2_X1 U28859 ( .A1(n28861), .A2(n28862), .ZN(n28860) );
  INV_X1 U28860 ( .A(n28863), .ZN(n28861) );
  AND2_X1 U28861 ( .A1(n28864), .A2(n28863), .ZN(n28859) );
  INV_X1 U28862 ( .A(n28862), .ZN(n28864) );
  AND2_X1 U28863 ( .A1(n28865), .A2(n28866), .ZN(n28465) );
  INV_X1 U28864 ( .A(n28867), .ZN(n28866) );
  AND2_X1 U28865 ( .A1(n28868), .A2(n28869), .ZN(n28867) );
  OR2_X1 U28866 ( .A1(n28869), .A2(n28868), .ZN(n28865) );
  OR2_X1 U28867 ( .A1(n28870), .A2(n28871), .ZN(n28868) );
  AND2_X1 U28868 ( .A1(n28872), .A2(n28873), .ZN(n28871) );
  INV_X1 U28869 ( .A(n28874), .ZN(n28872) );
  AND2_X1 U28870 ( .A1(n28875), .A2(n28874), .ZN(n28870) );
  INV_X1 U28871 ( .A(n28873), .ZN(n28875) );
  AND2_X1 U28872 ( .A1(n28876), .A2(n28877), .ZN(n28476) );
  INV_X1 U28873 ( .A(n28878), .ZN(n28877) );
  AND2_X1 U28874 ( .A1(n28879), .A2(n28880), .ZN(n28878) );
  OR2_X1 U28875 ( .A1(n28880), .A2(n28879), .ZN(n28876) );
  OR2_X1 U28876 ( .A1(n28881), .A2(n28882), .ZN(n28879) );
  AND2_X1 U28877 ( .A1(n28883), .A2(n28884), .ZN(n28882) );
  INV_X1 U28878 ( .A(n15873), .ZN(n28883) );
  AND2_X1 U28879 ( .A1(n28885), .A2(n15873), .ZN(n28881) );
  INV_X1 U28880 ( .A(n28884), .ZN(n28885) );
  AND2_X1 U28881 ( .A1(n28886), .A2(n28887), .ZN(n16412) );
  INV_X1 U28882 ( .A(n28888), .ZN(n28887) );
  AND2_X1 U28883 ( .A1(n28889), .A2(n28890), .ZN(n28888) );
  OR2_X1 U28884 ( .A1(n28890), .A2(n28889), .ZN(n28886) );
  OR2_X1 U28885 ( .A1(n28891), .A2(n28892), .ZN(n28889) );
  AND2_X1 U28886 ( .A1(n28893), .A2(n28894), .ZN(n28892) );
  INV_X1 U28887 ( .A(n28895), .ZN(n28893) );
  AND2_X1 U28888 ( .A1(n28896), .A2(n28895), .ZN(n28891) );
  INV_X1 U28889 ( .A(n28894), .ZN(n28896) );
  AND2_X1 U28890 ( .A1(n28897), .A2(n28898), .ZN(n16396) );
  INV_X1 U28891 ( .A(n28899), .ZN(n28898) );
  AND2_X1 U28892 ( .A1(n28900), .A2(n28901), .ZN(n28899) );
  OR2_X1 U28893 ( .A1(n28901), .A2(n28900), .ZN(n28897) );
  OR2_X1 U28894 ( .A1(n28902), .A2(n28903), .ZN(n28900) );
  AND2_X1 U28895 ( .A1(n28904), .A2(n28905), .ZN(n28903) );
  INV_X1 U28896 ( .A(n28906), .ZN(n28904) );
  AND2_X1 U28897 ( .A1(n28907), .A2(n28906), .ZN(n28902) );
  INV_X1 U28898 ( .A(n28905), .ZN(n28907) );
  AND2_X1 U28899 ( .A1(n16093), .A2(n16090), .ZN(n16386) );
  INV_X1 U28900 ( .A(n16092), .ZN(n16090) );
  AND2_X1 U28901 ( .A1(n28908), .A2(n28909), .ZN(n16092) );
  OR2_X1 U28902 ( .A1(n28910), .A2(n16389), .ZN(n28909) );
  INV_X1 U28903 ( .A(n28911), .ZN(n16389) );
  INV_X1 U28904 ( .A(n28912), .ZN(n28910) );
  OR2_X1 U28905 ( .A1(n28911), .A2(n28912), .ZN(n28908) );
  AND2_X1 U28906 ( .A1(b_0_), .A2(a_0_), .ZN(n28912) );
  OR2_X1 U28907 ( .A1(n28913), .A2(n28914), .ZN(n28911) );
  AND2_X1 U28908 ( .A1(n28915), .A2(n28916), .ZN(n28914) );
  AND2_X1 U28909 ( .A1(n28917), .A2(n28918), .ZN(n28913) );
  OR2_X1 U28910 ( .A1(n28916), .A2(n28915), .ZN(n28917) );
  INV_X1 U28911 ( .A(n16091), .ZN(n16093) );
  OR2_X1 U28912 ( .A1(n16392), .A2(n16393), .ZN(n16091) );
  OR2_X1 U28913 ( .A1(n28919), .A2(n28920), .ZN(n16393) );
  AND2_X1 U28914 ( .A1(n28906), .A2(n28905), .ZN(n28920) );
  AND2_X1 U28915 ( .A1(n28901), .A2(n28921), .ZN(n28919) );
  OR2_X1 U28916 ( .A1(n28905), .A2(n28906), .ZN(n28921) );
  OR2_X1 U28917 ( .A1(n16512), .A2(n15807), .ZN(n28906) );
  OR2_X1 U28918 ( .A1(n28922), .A2(n28923), .ZN(n28905) );
  AND2_X1 U28919 ( .A1(n28895), .A2(n28894), .ZN(n28923) );
  AND2_X1 U28920 ( .A1(n28890), .A2(n28924), .ZN(n28922) );
  OR2_X1 U28921 ( .A1(n28894), .A2(n28895), .ZN(n28924) );
  OR2_X1 U28922 ( .A1(n15842), .A2(n15807), .ZN(n28895) );
  INV_X1 U28923 ( .A(a_1_), .ZN(n15842) );
  OR2_X1 U28924 ( .A1(n28925), .A2(n28926), .ZN(n28894) );
  AND2_X1 U28925 ( .A1(n15873), .A2(n28884), .ZN(n28926) );
  AND2_X1 U28926 ( .A1(n28880), .A2(n28927), .ZN(n28925) );
  OR2_X1 U28927 ( .A1(n28884), .A2(n15873), .ZN(n28927) );
  OR2_X1 U28928 ( .A1(n15808), .A2(n15807), .ZN(n15873) );
  OR2_X1 U28929 ( .A1(n28928), .A2(n28929), .ZN(n28884) );
  AND2_X1 U28930 ( .A1(n28874), .A2(n28873), .ZN(n28929) );
  AND2_X1 U28931 ( .A1(n28869), .A2(n28930), .ZN(n28928) );
  OR2_X1 U28932 ( .A1(n28873), .A2(n28874), .ZN(n28930) );
  OR2_X1 U28933 ( .A1(n15774), .A2(n15807), .ZN(n28874) );
  OR2_X1 U28934 ( .A1(n28931), .A2(n28932), .ZN(n28873) );
  AND2_X1 U28935 ( .A1(n28863), .A2(n28862), .ZN(n28932) );
  AND2_X1 U28936 ( .A1(n28858), .A2(n28933), .ZN(n28931) );
  OR2_X1 U28937 ( .A1(n28862), .A2(n28863), .ZN(n28933) );
  OR2_X1 U28938 ( .A1(n15740), .A2(n15807), .ZN(n28863) );
  OR2_X1 U28939 ( .A1(n28934), .A2(n28935), .ZN(n28862) );
  AND2_X1 U28940 ( .A1(n28852), .A2(n28851), .ZN(n28935) );
  AND2_X1 U28941 ( .A1(n28847), .A2(n28936), .ZN(n28934) );
  OR2_X1 U28942 ( .A1(n28851), .A2(n28852), .ZN(n28936) );
  OR2_X1 U28943 ( .A1(n15706), .A2(n15807), .ZN(n28852) );
  OR2_X1 U28944 ( .A1(n28937), .A2(n28938), .ZN(n28851) );
  AND2_X1 U28945 ( .A1(n28841), .A2(n28840), .ZN(n28938) );
  AND2_X1 U28946 ( .A1(n28836), .A2(n28939), .ZN(n28937) );
  OR2_X1 U28947 ( .A1(n28840), .A2(n28841), .ZN(n28939) );
  OR2_X1 U28948 ( .A1(n15672), .A2(n15807), .ZN(n28841) );
  OR2_X1 U28949 ( .A1(n28940), .A2(n28941), .ZN(n28840) );
  AND2_X1 U28950 ( .A1(n28830), .A2(n28829), .ZN(n28941) );
  AND2_X1 U28951 ( .A1(n28825), .A2(n28942), .ZN(n28940) );
  OR2_X1 U28952 ( .A1(n28829), .A2(n28830), .ZN(n28942) );
  OR2_X1 U28953 ( .A1(n15638), .A2(n15807), .ZN(n28830) );
  OR2_X1 U28954 ( .A1(n28943), .A2(n28944), .ZN(n28829) );
  AND2_X1 U28955 ( .A1(n28819), .A2(n28818), .ZN(n28944) );
  AND2_X1 U28956 ( .A1(n28814), .A2(n28945), .ZN(n28943) );
  OR2_X1 U28957 ( .A1(n28818), .A2(n28819), .ZN(n28945) );
  OR2_X1 U28958 ( .A1(n15593), .A2(n15807), .ZN(n28819) );
  OR2_X1 U28959 ( .A1(n28946), .A2(n28947), .ZN(n28818) );
  AND2_X1 U28960 ( .A1(n28808), .A2(n28807), .ZN(n28947) );
  AND2_X1 U28961 ( .A1(n28803), .A2(n28948), .ZN(n28946) );
  OR2_X1 U28962 ( .A1(n28807), .A2(n28808), .ZN(n28948) );
  OR2_X1 U28963 ( .A1(n15559), .A2(n15807), .ZN(n28808) );
  INV_X1 U28964 ( .A(a_9_), .ZN(n15559) );
  OR2_X1 U28965 ( .A1(n28949), .A2(n28950), .ZN(n28807) );
  AND2_X1 U28966 ( .A1(n28797), .A2(n28796), .ZN(n28950) );
  AND2_X1 U28967 ( .A1(n28792), .A2(n28951), .ZN(n28949) );
  OR2_X1 U28968 ( .A1(n28796), .A2(n28797), .ZN(n28951) );
  OR2_X1 U28969 ( .A1(n15525), .A2(n15807), .ZN(n28797) );
  OR2_X1 U28970 ( .A1(n28952), .A2(n28953), .ZN(n28796) );
  AND2_X1 U28971 ( .A1(n28786), .A2(n28785), .ZN(n28953) );
  AND2_X1 U28972 ( .A1(n28781), .A2(n28954), .ZN(n28952) );
  OR2_X1 U28973 ( .A1(n28785), .A2(n28786), .ZN(n28954) );
  OR2_X1 U28974 ( .A1(n15491), .A2(n15807), .ZN(n28786) );
  OR2_X1 U28975 ( .A1(n28955), .A2(n28956), .ZN(n28785) );
  AND2_X1 U28976 ( .A1(n28775), .A2(n28774), .ZN(n28956) );
  AND2_X1 U28977 ( .A1(n28770), .A2(n28957), .ZN(n28955) );
  OR2_X1 U28978 ( .A1(n28774), .A2(n28775), .ZN(n28957) );
  OR2_X1 U28979 ( .A1(n15457), .A2(n15807), .ZN(n28775) );
  OR2_X1 U28980 ( .A1(n28958), .A2(n28959), .ZN(n28774) );
  AND2_X1 U28981 ( .A1(n28764), .A2(n28763), .ZN(n28959) );
  AND2_X1 U28982 ( .A1(n28759), .A2(n28960), .ZN(n28958) );
  OR2_X1 U28983 ( .A1(n28763), .A2(n28764), .ZN(n28960) );
  OR2_X1 U28984 ( .A1(n15423), .A2(n15807), .ZN(n28764) );
  OR2_X1 U28985 ( .A1(n28961), .A2(n28962), .ZN(n28763) );
  AND2_X1 U28986 ( .A1(n28753), .A2(n28752), .ZN(n28962) );
  AND2_X1 U28987 ( .A1(n28748), .A2(n28963), .ZN(n28961) );
  OR2_X1 U28988 ( .A1(n28752), .A2(n28753), .ZN(n28963) );
  OR2_X1 U28989 ( .A1(n15389), .A2(n15807), .ZN(n28753) );
  OR2_X1 U28990 ( .A1(n28964), .A2(n28965), .ZN(n28752) );
  AND2_X1 U28991 ( .A1(n28742), .A2(n28741), .ZN(n28965) );
  AND2_X1 U28992 ( .A1(n28737), .A2(n28966), .ZN(n28964) );
  OR2_X1 U28993 ( .A1(n28741), .A2(n28742), .ZN(n28966) );
  OR2_X1 U28994 ( .A1(n15355), .A2(n15807), .ZN(n28742) );
  OR2_X1 U28995 ( .A1(n28967), .A2(n28968), .ZN(n28741) );
  AND2_X1 U28996 ( .A1(n28731), .A2(n28730), .ZN(n28968) );
  AND2_X1 U28997 ( .A1(n28726), .A2(n28969), .ZN(n28967) );
  OR2_X1 U28998 ( .A1(n28730), .A2(n28731), .ZN(n28969) );
  OR2_X1 U28999 ( .A1(n15321), .A2(n15807), .ZN(n28731) );
  OR2_X1 U29000 ( .A1(n28970), .A2(n28971), .ZN(n28730) );
  AND2_X1 U29001 ( .A1(n28720), .A2(n28719), .ZN(n28971) );
  AND2_X1 U29002 ( .A1(n28715), .A2(n28972), .ZN(n28970) );
  OR2_X1 U29003 ( .A1(n28719), .A2(n28720), .ZN(n28972) );
  OR2_X1 U29004 ( .A1(n15287), .A2(n15807), .ZN(n28720) );
  OR2_X1 U29005 ( .A1(n28973), .A2(n28974), .ZN(n28719) );
  AND2_X1 U29006 ( .A1(n28709), .A2(n28708), .ZN(n28974) );
  AND2_X1 U29007 ( .A1(n28704), .A2(n28975), .ZN(n28973) );
  OR2_X1 U29008 ( .A1(n28708), .A2(n28709), .ZN(n28975) );
  OR2_X1 U29009 ( .A1(n15242), .A2(n15807), .ZN(n28709) );
  OR2_X1 U29010 ( .A1(n28976), .A2(n28977), .ZN(n28708) );
  AND2_X1 U29011 ( .A1(n28698), .A2(n28697), .ZN(n28977) );
  AND2_X1 U29012 ( .A1(n28693), .A2(n28978), .ZN(n28976) );
  OR2_X1 U29013 ( .A1(n28697), .A2(n28698), .ZN(n28978) );
  OR2_X1 U29014 ( .A1(n15208), .A2(n15807), .ZN(n28698) );
  OR2_X1 U29015 ( .A1(n28979), .A2(n28980), .ZN(n28697) );
  AND2_X1 U29016 ( .A1(n28687), .A2(n28686), .ZN(n28980) );
  AND2_X1 U29017 ( .A1(n28682), .A2(n28981), .ZN(n28979) );
  OR2_X1 U29018 ( .A1(n28686), .A2(n28687), .ZN(n28981) );
  OR2_X1 U29019 ( .A1(n15174), .A2(n15807), .ZN(n28687) );
  OR2_X1 U29020 ( .A1(n28982), .A2(n28983), .ZN(n28686) );
  AND2_X1 U29021 ( .A1(n28676), .A2(n28675), .ZN(n28983) );
  AND2_X1 U29022 ( .A1(n28671), .A2(n28984), .ZN(n28982) );
  OR2_X1 U29023 ( .A1(n28675), .A2(n28676), .ZN(n28984) );
  OR2_X1 U29024 ( .A1(n15140), .A2(n15807), .ZN(n28676) );
  OR2_X1 U29025 ( .A1(n28985), .A2(n28986), .ZN(n28675) );
  AND2_X1 U29026 ( .A1(n28665), .A2(n28664), .ZN(n28986) );
  AND2_X1 U29027 ( .A1(n28660), .A2(n28987), .ZN(n28985) );
  OR2_X1 U29028 ( .A1(n28664), .A2(n28665), .ZN(n28987) );
  OR2_X1 U29029 ( .A1(n15106), .A2(n15807), .ZN(n28665) );
  OR2_X1 U29030 ( .A1(n28988), .A2(n28989), .ZN(n28664) );
  AND2_X1 U29031 ( .A1(n28654), .A2(n28653), .ZN(n28989) );
  AND2_X1 U29032 ( .A1(n28649), .A2(n28990), .ZN(n28988) );
  OR2_X1 U29033 ( .A1(n28653), .A2(n28654), .ZN(n28990) );
  OR2_X1 U29034 ( .A1(n15072), .A2(n15807), .ZN(n28654) );
  OR2_X1 U29035 ( .A1(n28991), .A2(n28992), .ZN(n28653) );
  AND2_X1 U29036 ( .A1(n28643), .A2(n28642), .ZN(n28992) );
  AND2_X1 U29037 ( .A1(n28638), .A2(n28993), .ZN(n28991) );
  OR2_X1 U29038 ( .A1(n28642), .A2(n28643), .ZN(n28993) );
  OR2_X1 U29039 ( .A1(n15038), .A2(n15807), .ZN(n28643) );
  OR2_X1 U29040 ( .A1(n28994), .A2(n28995), .ZN(n28642) );
  AND2_X1 U29041 ( .A1(n28632), .A2(n28631), .ZN(n28995) );
  AND2_X1 U29042 ( .A1(n28627), .A2(n28996), .ZN(n28994) );
  OR2_X1 U29043 ( .A1(n28631), .A2(n28632), .ZN(n28996) );
  OR2_X1 U29044 ( .A1(n15004), .A2(n15807), .ZN(n28632) );
  OR2_X1 U29045 ( .A1(n28997), .A2(n28998), .ZN(n28631) );
  AND2_X1 U29046 ( .A1(n28621), .A2(n28620), .ZN(n28998) );
  AND2_X1 U29047 ( .A1(n28616), .A2(n28999), .ZN(n28997) );
  OR2_X1 U29048 ( .A1(n28620), .A2(n28621), .ZN(n28999) );
  OR2_X1 U29049 ( .A1(n14970), .A2(n15807), .ZN(n28621) );
  OR2_X1 U29050 ( .A1(n29000), .A2(n29001), .ZN(n28620) );
  AND2_X1 U29051 ( .A1(n28605), .A2(n28611), .ZN(n29001) );
  AND2_X1 U29052 ( .A1(n29002), .A2(n28610), .ZN(n29000) );
  OR2_X1 U29053 ( .A1(n29003), .A2(n29004), .ZN(n28610) );
  AND2_X1 U29054 ( .A1(n28597), .A2(n28599), .ZN(n29004) );
  AND2_X1 U29055 ( .A1(n28594), .A2(n29005), .ZN(n29003) );
  OR2_X1 U29056 ( .A1(n28599), .A2(n28597), .ZN(n29005) );
  OR2_X1 U29057 ( .A1(n14891), .A2(n15807), .ZN(n28597) );
  OR2_X1 U29058 ( .A1(n29006), .A2(n29007), .ZN(n28599) );
  AND2_X1 U29059 ( .A1(n28582), .A2(n28587), .ZN(n29007) );
  AND2_X1 U29060 ( .A1(n28586), .A2(n29008), .ZN(n29006) );
  OR2_X1 U29061 ( .A1(n28587), .A2(n28582), .ZN(n29008) );
  OR2_X1 U29062 ( .A1(n14857), .A2(n15807), .ZN(n28582) );
  INV_X1 U29063 ( .A(n28588), .ZN(n28587) );
  AND3_X1 U29064 ( .A1(b_2_), .A2(b_1_), .A3(n15957), .ZN(n28588) );
  INV_X1 U29065 ( .A(n28589), .ZN(n28586) );
  OR2_X1 U29066 ( .A1(n29009), .A2(n29010), .ZN(n28589) );
  AND2_X1 U29067 ( .A1(b_1_), .A2(n29011), .ZN(n29010) );
  OR2_X1 U29068 ( .A1(n29012), .A2(n16981), .ZN(n29011) );
  AND2_X1 U29069 ( .A1(n15958), .A2(a_30_), .ZN(n16981) );
  INV_X1 U29070 ( .A(a_31_), .ZN(n15958) );
  AND2_X1 U29071 ( .A1(a_30_), .A2(n16294), .ZN(n29012) );
  AND2_X1 U29072 ( .A1(b_0_), .A2(n29013), .ZN(n29009) );
  OR2_X1 U29073 ( .A1(n29014), .A2(n14817), .ZN(n29013) );
  AND2_X1 U29074 ( .A1(n14806), .A2(a_31_), .ZN(n14817) );
  AND2_X1 U29075 ( .A1(a_31_), .A2(n15841), .ZN(n29014) );
  OR2_X1 U29076 ( .A1(n29015), .A2(n29016), .ZN(n28594) );
  INV_X1 U29077 ( .A(n29017), .ZN(n29016) );
  OR2_X1 U29078 ( .A1(n29018), .A2(n29019), .ZN(n29017) );
  AND2_X1 U29079 ( .A1(n29019), .A2(n29018), .ZN(n29015) );
  OR2_X1 U29080 ( .A1(n29020), .A2(n29021), .ZN(n29018) );
  AND3_X1 U29081 ( .A1(a_29_), .A2(n29022), .A3(b_1_), .ZN(n29021) );
  OR2_X1 U29082 ( .A1(n16294), .A2(n14806), .ZN(n29022) );
  INV_X1 U29083 ( .A(a_30_), .ZN(n14806) );
  AND3_X1 U29084 ( .A1(b_0_), .A2(n29023), .A3(a_30_), .ZN(n29020) );
  OR2_X1 U29085 ( .A1(n14857), .A2(n15841), .ZN(n29023) );
  OR2_X1 U29086 ( .A1(n28611), .A2(n28605), .ZN(n29002) );
  OR2_X1 U29087 ( .A1(n29024), .A2(n29025), .ZN(n28605) );
  AND2_X1 U29088 ( .A1(n29026), .A2(n29027), .ZN(n29025) );
  INV_X1 U29089 ( .A(n29028), .ZN(n29026) );
  AND2_X1 U29090 ( .A1(n29028), .A2(n29029), .ZN(n29024) );
  AND2_X1 U29091 ( .A1(n29030), .A2(n29031), .ZN(n29028) );
  OR2_X1 U29092 ( .A1(n29032), .A2(n29033), .ZN(n29031) );
  INV_X1 U29093 ( .A(n29034), .ZN(n29030) );
  AND2_X1 U29094 ( .A1(n29033), .A2(n29032), .ZN(n29034) );
  OR2_X1 U29095 ( .A1(n14936), .A2(n15807), .ZN(n28611) );
  INV_X1 U29096 ( .A(b_2_), .ZN(n15807) );
  AND2_X1 U29097 ( .A1(n29035), .A2(n29036), .ZN(n28616) );
  INV_X1 U29098 ( .A(n29037), .ZN(n29036) );
  AND2_X1 U29099 ( .A1(n29038), .A2(n29039), .ZN(n29037) );
  OR2_X1 U29100 ( .A1(n29038), .A2(n29039), .ZN(n29035) );
  OR2_X1 U29101 ( .A1(n29040), .A2(n29041), .ZN(n29038) );
  AND2_X1 U29102 ( .A1(n29042), .A2(n29043), .ZN(n29041) );
  AND2_X1 U29103 ( .A1(n29044), .A2(n29045), .ZN(n29040) );
  INV_X1 U29104 ( .A(n29043), .ZN(n29044) );
  AND2_X1 U29105 ( .A1(n29046), .A2(n29047), .ZN(n28627) );
  INV_X1 U29106 ( .A(n29048), .ZN(n29047) );
  AND2_X1 U29107 ( .A1(n29049), .A2(n29050), .ZN(n29048) );
  OR2_X1 U29108 ( .A1(n29049), .A2(n29050), .ZN(n29046) );
  OR2_X1 U29109 ( .A1(n29051), .A2(n29052), .ZN(n29049) );
  AND2_X1 U29110 ( .A1(n29053), .A2(n29054), .ZN(n29052) );
  AND2_X1 U29111 ( .A1(n29055), .A2(n29056), .ZN(n29051) );
  INV_X1 U29112 ( .A(n29054), .ZN(n29055) );
  AND2_X1 U29113 ( .A1(n29057), .A2(n29058), .ZN(n28638) );
  INV_X1 U29114 ( .A(n29059), .ZN(n29058) );
  AND2_X1 U29115 ( .A1(n29060), .A2(n29061), .ZN(n29059) );
  OR2_X1 U29116 ( .A1(n29060), .A2(n29061), .ZN(n29057) );
  OR2_X1 U29117 ( .A1(n29062), .A2(n29063), .ZN(n29060) );
  AND2_X1 U29118 ( .A1(n29064), .A2(n29065), .ZN(n29063) );
  AND2_X1 U29119 ( .A1(n29066), .A2(n29067), .ZN(n29062) );
  INV_X1 U29120 ( .A(n29065), .ZN(n29066) );
  AND2_X1 U29121 ( .A1(n29068), .A2(n29069), .ZN(n28649) );
  INV_X1 U29122 ( .A(n29070), .ZN(n29069) );
  AND2_X1 U29123 ( .A1(n29071), .A2(n29072), .ZN(n29070) );
  OR2_X1 U29124 ( .A1(n29071), .A2(n29072), .ZN(n29068) );
  OR2_X1 U29125 ( .A1(n29073), .A2(n29074), .ZN(n29071) );
  AND2_X1 U29126 ( .A1(n29075), .A2(n29076), .ZN(n29074) );
  AND2_X1 U29127 ( .A1(n29077), .A2(n29078), .ZN(n29073) );
  INV_X1 U29128 ( .A(n29076), .ZN(n29077) );
  AND2_X1 U29129 ( .A1(n29079), .A2(n29080), .ZN(n28660) );
  INV_X1 U29130 ( .A(n29081), .ZN(n29080) );
  AND2_X1 U29131 ( .A1(n29082), .A2(n29083), .ZN(n29081) );
  OR2_X1 U29132 ( .A1(n29082), .A2(n29083), .ZN(n29079) );
  OR2_X1 U29133 ( .A1(n29084), .A2(n29085), .ZN(n29082) );
  AND2_X1 U29134 ( .A1(n29086), .A2(n29087), .ZN(n29085) );
  AND2_X1 U29135 ( .A1(n29088), .A2(n29089), .ZN(n29084) );
  INV_X1 U29136 ( .A(n29087), .ZN(n29088) );
  AND2_X1 U29137 ( .A1(n29090), .A2(n29091), .ZN(n28671) );
  INV_X1 U29138 ( .A(n29092), .ZN(n29091) );
  AND2_X1 U29139 ( .A1(n29093), .A2(n29094), .ZN(n29092) );
  OR2_X1 U29140 ( .A1(n29093), .A2(n29094), .ZN(n29090) );
  OR2_X1 U29141 ( .A1(n29095), .A2(n29096), .ZN(n29093) );
  AND2_X1 U29142 ( .A1(n29097), .A2(n29098), .ZN(n29096) );
  AND2_X1 U29143 ( .A1(n29099), .A2(n29100), .ZN(n29095) );
  INV_X1 U29144 ( .A(n29098), .ZN(n29099) );
  AND2_X1 U29145 ( .A1(n29101), .A2(n29102), .ZN(n28682) );
  INV_X1 U29146 ( .A(n29103), .ZN(n29102) );
  AND2_X1 U29147 ( .A1(n29104), .A2(n29105), .ZN(n29103) );
  OR2_X1 U29148 ( .A1(n29104), .A2(n29105), .ZN(n29101) );
  OR2_X1 U29149 ( .A1(n29106), .A2(n29107), .ZN(n29104) );
  AND2_X1 U29150 ( .A1(n29108), .A2(n29109), .ZN(n29107) );
  AND2_X1 U29151 ( .A1(n29110), .A2(n29111), .ZN(n29106) );
  INV_X1 U29152 ( .A(n29109), .ZN(n29110) );
  AND2_X1 U29153 ( .A1(n29112), .A2(n29113), .ZN(n28693) );
  INV_X1 U29154 ( .A(n29114), .ZN(n29113) );
  AND2_X1 U29155 ( .A1(n29115), .A2(n29116), .ZN(n29114) );
  OR2_X1 U29156 ( .A1(n29115), .A2(n29116), .ZN(n29112) );
  OR2_X1 U29157 ( .A1(n29117), .A2(n29118), .ZN(n29115) );
  AND2_X1 U29158 ( .A1(n29119), .A2(n29120), .ZN(n29118) );
  AND2_X1 U29159 ( .A1(n29121), .A2(n29122), .ZN(n29117) );
  INV_X1 U29160 ( .A(n29120), .ZN(n29121) );
  AND2_X1 U29161 ( .A1(n29123), .A2(n29124), .ZN(n28704) );
  INV_X1 U29162 ( .A(n29125), .ZN(n29124) );
  AND2_X1 U29163 ( .A1(n29126), .A2(n29127), .ZN(n29125) );
  OR2_X1 U29164 ( .A1(n29126), .A2(n29127), .ZN(n29123) );
  OR2_X1 U29165 ( .A1(n29128), .A2(n29129), .ZN(n29126) );
  AND2_X1 U29166 ( .A1(n29130), .A2(n29131), .ZN(n29129) );
  AND2_X1 U29167 ( .A1(n29132), .A2(n29133), .ZN(n29128) );
  INV_X1 U29168 ( .A(n29131), .ZN(n29132) );
  AND2_X1 U29169 ( .A1(n29134), .A2(n29135), .ZN(n28715) );
  INV_X1 U29170 ( .A(n29136), .ZN(n29135) );
  AND2_X1 U29171 ( .A1(n29137), .A2(n29138), .ZN(n29136) );
  OR2_X1 U29172 ( .A1(n29137), .A2(n29138), .ZN(n29134) );
  OR2_X1 U29173 ( .A1(n29139), .A2(n29140), .ZN(n29137) );
  AND2_X1 U29174 ( .A1(n29141), .A2(n29142), .ZN(n29140) );
  AND2_X1 U29175 ( .A1(n29143), .A2(n29144), .ZN(n29139) );
  INV_X1 U29176 ( .A(n29142), .ZN(n29143) );
  AND2_X1 U29177 ( .A1(n29145), .A2(n29146), .ZN(n28726) );
  INV_X1 U29178 ( .A(n29147), .ZN(n29146) );
  AND2_X1 U29179 ( .A1(n29148), .A2(n29149), .ZN(n29147) );
  OR2_X1 U29180 ( .A1(n29148), .A2(n29149), .ZN(n29145) );
  OR2_X1 U29181 ( .A1(n29150), .A2(n29151), .ZN(n29148) );
  AND2_X1 U29182 ( .A1(n29152), .A2(n29153), .ZN(n29151) );
  AND2_X1 U29183 ( .A1(n29154), .A2(n29155), .ZN(n29150) );
  INV_X1 U29184 ( .A(n29153), .ZN(n29154) );
  AND2_X1 U29185 ( .A1(n29156), .A2(n29157), .ZN(n28737) );
  INV_X1 U29186 ( .A(n29158), .ZN(n29157) );
  AND2_X1 U29187 ( .A1(n29159), .A2(n29160), .ZN(n29158) );
  OR2_X1 U29188 ( .A1(n29159), .A2(n29160), .ZN(n29156) );
  OR2_X1 U29189 ( .A1(n29161), .A2(n29162), .ZN(n29159) );
  AND2_X1 U29190 ( .A1(n29163), .A2(n29164), .ZN(n29162) );
  AND2_X1 U29191 ( .A1(n29165), .A2(n29166), .ZN(n29161) );
  INV_X1 U29192 ( .A(n29164), .ZN(n29165) );
  AND2_X1 U29193 ( .A1(n29167), .A2(n29168), .ZN(n28748) );
  INV_X1 U29194 ( .A(n29169), .ZN(n29168) );
  AND2_X1 U29195 ( .A1(n29170), .A2(n29171), .ZN(n29169) );
  OR2_X1 U29196 ( .A1(n29170), .A2(n29171), .ZN(n29167) );
  OR2_X1 U29197 ( .A1(n29172), .A2(n29173), .ZN(n29170) );
  AND2_X1 U29198 ( .A1(n29174), .A2(n29175), .ZN(n29173) );
  AND2_X1 U29199 ( .A1(n29176), .A2(n29177), .ZN(n29172) );
  INV_X1 U29200 ( .A(n29175), .ZN(n29176) );
  AND2_X1 U29201 ( .A1(n29178), .A2(n29179), .ZN(n28759) );
  INV_X1 U29202 ( .A(n29180), .ZN(n29179) );
  AND2_X1 U29203 ( .A1(n29181), .A2(n29182), .ZN(n29180) );
  OR2_X1 U29204 ( .A1(n29181), .A2(n29182), .ZN(n29178) );
  OR2_X1 U29205 ( .A1(n29183), .A2(n29184), .ZN(n29181) );
  AND2_X1 U29206 ( .A1(n29185), .A2(n29186), .ZN(n29184) );
  AND2_X1 U29207 ( .A1(n29187), .A2(n29188), .ZN(n29183) );
  INV_X1 U29208 ( .A(n29186), .ZN(n29187) );
  AND2_X1 U29209 ( .A1(n29189), .A2(n29190), .ZN(n28770) );
  INV_X1 U29210 ( .A(n29191), .ZN(n29190) );
  AND2_X1 U29211 ( .A1(n29192), .A2(n29193), .ZN(n29191) );
  OR2_X1 U29212 ( .A1(n29192), .A2(n29193), .ZN(n29189) );
  OR2_X1 U29213 ( .A1(n29194), .A2(n29195), .ZN(n29192) );
  AND2_X1 U29214 ( .A1(n29196), .A2(n29197), .ZN(n29195) );
  AND2_X1 U29215 ( .A1(n29198), .A2(n29199), .ZN(n29194) );
  INV_X1 U29216 ( .A(n29197), .ZN(n29198) );
  AND2_X1 U29217 ( .A1(n29200), .A2(n29201), .ZN(n28781) );
  INV_X1 U29218 ( .A(n29202), .ZN(n29201) );
  AND2_X1 U29219 ( .A1(n29203), .A2(n29204), .ZN(n29202) );
  OR2_X1 U29220 ( .A1(n29203), .A2(n29204), .ZN(n29200) );
  OR2_X1 U29221 ( .A1(n29205), .A2(n29206), .ZN(n29203) );
  AND2_X1 U29222 ( .A1(n29207), .A2(n29208), .ZN(n29206) );
  AND2_X1 U29223 ( .A1(n29209), .A2(n29210), .ZN(n29205) );
  INV_X1 U29224 ( .A(n29208), .ZN(n29209) );
  AND2_X1 U29225 ( .A1(n29211), .A2(n29212), .ZN(n28792) );
  INV_X1 U29226 ( .A(n29213), .ZN(n29212) );
  AND2_X1 U29227 ( .A1(n29214), .A2(n29215), .ZN(n29213) );
  OR2_X1 U29228 ( .A1(n29214), .A2(n29215), .ZN(n29211) );
  OR2_X1 U29229 ( .A1(n29216), .A2(n29217), .ZN(n29214) );
  AND2_X1 U29230 ( .A1(n29218), .A2(n29219), .ZN(n29217) );
  AND2_X1 U29231 ( .A1(n29220), .A2(n29221), .ZN(n29216) );
  INV_X1 U29232 ( .A(n29219), .ZN(n29220) );
  AND2_X1 U29233 ( .A1(n29222), .A2(n29223), .ZN(n28803) );
  INV_X1 U29234 ( .A(n29224), .ZN(n29223) );
  AND2_X1 U29235 ( .A1(n29225), .A2(n29226), .ZN(n29224) );
  OR2_X1 U29236 ( .A1(n29225), .A2(n29226), .ZN(n29222) );
  OR2_X1 U29237 ( .A1(n29227), .A2(n29228), .ZN(n29225) );
  AND2_X1 U29238 ( .A1(n29229), .A2(n29230), .ZN(n29228) );
  AND2_X1 U29239 ( .A1(n29231), .A2(n29232), .ZN(n29227) );
  INV_X1 U29240 ( .A(n29230), .ZN(n29231) );
  AND2_X1 U29241 ( .A1(n29233), .A2(n29234), .ZN(n28814) );
  INV_X1 U29242 ( .A(n29235), .ZN(n29234) );
  AND2_X1 U29243 ( .A1(n29236), .A2(n29237), .ZN(n29235) );
  OR2_X1 U29244 ( .A1(n29236), .A2(n29237), .ZN(n29233) );
  OR2_X1 U29245 ( .A1(n29238), .A2(n29239), .ZN(n29236) );
  AND2_X1 U29246 ( .A1(n29240), .A2(n29241), .ZN(n29239) );
  AND2_X1 U29247 ( .A1(n29242), .A2(n29243), .ZN(n29238) );
  INV_X1 U29248 ( .A(n29241), .ZN(n29242) );
  AND2_X1 U29249 ( .A1(n29244), .A2(n29245), .ZN(n28825) );
  INV_X1 U29250 ( .A(n29246), .ZN(n29245) );
  AND2_X1 U29251 ( .A1(n29247), .A2(n29248), .ZN(n29246) );
  OR2_X1 U29252 ( .A1(n29247), .A2(n29248), .ZN(n29244) );
  OR2_X1 U29253 ( .A1(n29249), .A2(n29250), .ZN(n29247) );
  INV_X1 U29254 ( .A(n29251), .ZN(n29250) );
  OR2_X1 U29255 ( .A1(n29252), .A2(n29253), .ZN(n29251) );
  AND2_X1 U29256 ( .A1(n29253), .A2(n29252), .ZN(n29249) );
  AND2_X1 U29257 ( .A1(n29254), .A2(n29255), .ZN(n28836) );
  INV_X1 U29258 ( .A(n29256), .ZN(n29255) );
  AND2_X1 U29259 ( .A1(n29257), .A2(n29258), .ZN(n29256) );
  OR2_X1 U29260 ( .A1(n29257), .A2(n29258), .ZN(n29254) );
  OR2_X1 U29261 ( .A1(n29259), .A2(n29260), .ZN(n29257) );
  INV_X1 U29262 ( .A(n29261), .ZN(n29260) );
  OR2_X1 U29263 ( .A1(n29262), .A2(n29263), .ZN(n29261) );
  AND2_X1 U29264 ( .A1(n29263), .A2(n29262), .ZN(n29259) );
  AND2_X1 U29265 ( .A1(n29264), .A2(n29265), .ZN(n28847) );
  INV_X1 U29266 ( .A(n29266), .ZN(n29265) );
  AND2_X1 U29267 ( .A1(n29267), .A2(n29268), .ZN(n29266) );
  OR2_X1 U29268 ( .A1(n29267), .A2(n29268), .ZN(n29264) );
  OR2_X1 U29269 ( .A1(n29269), .A2(n29270), .ZN(n29267) );
  INV_X1 U29270 ( .A(n29271), .ZN(n29270) );
  OR2_X1 U29271 ( .A1(n29272), .A2(n29273), .ZN(n29271) );
  AND2_X1 U29272 ( .A1(n29273), .A2(n29272), .ZN(n29269) );
  AND2_X1 U29273 ( .A1(n29274), .A2(n29275), .ZN(n28858) );
  INV_X1 U29274 ( .A(n29276), .ZN(n29275) );
  AND2_X1 U29275 ( .A1(n29277), .A2(n29278), .ZN(n29276) );
  OR2_X1 U29276 ( .A1(n29277), .A2(n29278), .ZN(n29274) );
  OR2_X1 U29277 ( .A1(n29279), .A2(n29280), .ZN(n29277) );
  INV_X1 U29278 ( .A(n29281), .ZN(n29280) );
  OR2_X1 U29279 ( .A1(n29282), .A2(n29283), .ZN(n29281) );
  AND2_X1 U29280 ( .A1(n29283), .A2(n29282), .ZN(n29279) );
  AND2_X1 U29281 ( .A1(n29284), .A2(n29285), .ZN(n28869) );
  INV_X1 U29282 ( .A(n29286), .ZN(n29285) );
  AND2_X1 U29283 ( .A1(n29287), .A2(n29288), .ZN(n29286) );
  OR2_X1 U29284 ( .A1(n29287), .A2(n29288), .ZN(n29284) );
  OR2_X1 U29285 ( .A1(n29289), .A2(n29290), .ZN(n29287) );
  INV_X1 U29286 ( .A(n29291), .ZN(n29290) );
  OR2_X1 U29287 ( .A1(n29292), .A2(n29293), .ZN(n29291) );
  AND2_X1 U29288 ( .A1(n29293), .A2(n29292), .ZN(n29289) );
  AND2_X1 U29289 ( .A1(n29294), .A2(n29295), .ZN(n28880) );
  INV_X1 U29290 ( .A(n29296), .ZN(n29295) );
  AND2_X1 U29291 ( .A1(n29297), .A2(n29298), .ZN(n29296) );
  OR2_X1 U29292 ( .A1(n29297), .A2(n29298), .ZN(n29294) );
  OR2_X1 U29293 ( .A1(n29299), .A2(n29300), .ZN(n29297) );
  INV_X1 U29294 ( .A(n29301), .ZN(n29300) );
  OR2_X1 U29295 ( .A1(n29302), .A2(n29303), .ZN(n29301) );
  AND2_X1 U29296 ( .A1(n29303), .A2(n29302), .ZN(n29299) );
  AND2_X1 U29297 ( .A1(n29304), .A2(n29305), .ZN(n28890) );
  INV_X1 U29298 ( .A(n29306), .ZN(n29305) );
  AND2_X1 U29299 ( .A1(n29307), .A2(n29308), .ZN(n29306) );
  OR2_X1 U29300 ( .A1(n29307), .A2(n29308), .ZN(n29304) );
  OR2_X1 U29301 ( .A1(n29309), .A2(n29310), .ZN(n29307) );
  INV_X1 U29302 ( .A(n29311), .ZN(n29310) );
  OR2_X1 U29303 ( .A1(n29312), .A2(n29313), .ZN(n29311) );
  AND2_X1 U29304 ( .A1(n29313), .A2(n29312), .ZN(n29309) );
  AND2_X1 U29305 ( .A1(n29314), .A2(n29315), .ZN(n28901) );
  INV_X1 U29306 ( .A(n29316), .ZN(n29315) );
  AND2_X1 U29307 ( .A1(n29317), .A2(n29318), .ZN(n29316) );
  OR2_X1 U29308 ( .A1(n29317), .A2(n29318), .ZN(n29314) );
  OR2_X1 U29309 ( .A1(n29319), .A2(n29320), .ZN(n29317) );
  INV_X1 U29310 ( .A(n29321), .ZN(n29320) );
  OR2_X1 U29311 ( .A1(n29322), .A2(n29323), .ZN(n29321) );
  AND2_X1 U29312 ( .A1(n29323), .A2(n29322), .ZN(n29319) );
  AND2_X1 U29313 ( .A1(n29324), .A2(n29325), .ZN(n16392) );
  INV_X1 U29314 ( .A(n29326), .ZN(n29325) );
  AND2_X1 U29315 ( .A1(n29327), .A2(n28915), .ZN(n29326) );
  OR2_X1 U29316 ( .A1(n29327), .A2(n28915), .ZN(n29324) );
  OR2_X1 U29317 ( .A1(n29328), .A2(n29329), .ZN(n28915) );
  AND2_X1 U29318 ( .A1(n29318), .A2(n29322), .ZN(n29329) );
  AND2_X1 U29319 ( .A1(n29330), .A2(n15870), .ZN(n29328) );
  INV_X1 U29320 ( .A(n29323), .ZN(n15870) );
  AND2_X1 U29321 ( .A1(a_1_), .A2(b_1_), .ZN(n29323) );
  OR2_X1 U29322 ( .A1(n29322), .A2(n29318), .ZN(n29330) );
  OR2_X1 U29323 ( .A1(n16294), .A2(n15808), .ZN(n29318) );
  OR2_X1 U29324 ( .A1(n29331), .A2(n29332), .ZN(n29322) );
  AND2_X1 U29325 ( .A1(n29308), .A2(n29312), .ZN(n29332) );
  AND2_X1 U29326 ( .A1(n29333), .A2(n29334), .ZN(n29331) );
  INV_X1 U29327 ( .A(n29313), .ZN(n29334) );
  AND2_X1 U29328 ( .A1(b_0_), .A2(a_3_), .ZN(n29313) );
  OR2_X1 U29329 ( .A1(n29312), .A2(n29308), .ZN(n29333) );
  OR2_X1 U29330 ( .A1(n15808), .A2(n15841), .ZN(n29308) );
  OR2_X1 U29331 ( .A1(n29335), .A2(n29336), .ZN(n29312) );
  AND2_X1 U29332 ( .A1(n29298), .A2(n29302), .ZN(n29336) );
  AND2_X1 U29333 ( .A1(n29337), .A2(n29338), .ZN(n29335) );
  INV_X1 U29334 ( .A(n29303), .ZN(n29338) );
  AND2_X1 U29335 ( .A1(b_0_), .A2(a_4_), .ZN(n29303) );
  OR2_X1 U29336 ( .A1(n29302), .A2(n29298), .ZN(n29337) );
  OR2_X1 U29337 ( .A1(n15774), .A2(n15841), .ZN(n29298) );
  INV_X1 U29338 ( .A(a_3_), .ZN(n15774) );
  OR2_X1 U29339 ( .A1(n29339), .A2(n29340), .ZN(n29302) );
  AND2_X1 U29340 ( .A1(n29288), .A2(n29292), .ZN(n29340) );
  AND2_X1 U29341 ( .A1(n29341), .A2(n29342), .ZN(n29339) );
  INV_X1 U29342 ( .A(n29293), .ZN(n29342) );
  AND2_X1 U29343 ( .A1(b_0_), .A2(a_5_), .ZN(n29293) );
  OR2_X1 U29344 ( .A1(n29292), .A2(n29288), .ZN(n29341) );
  OR2_X1 U29345 ( .A1(n15740), .A2(n15841), .ZN(n29288) );
  INV_X1 U29346 ( .A(a_4_), .ZN(n15740) );
  OR2_X1 U29347 ( .A1(n29343), .A2(n29344), .ZN(n29292) );
  AND2_X1 U29348 ( .A1(n29278), .A2(n29282), .ZN(n29344) );
  AND2_X1 U29349 ( .A1(n29345), .A2(n29346), .ZN(n29343) );
  INV_X1 U29350 ( .A(n29283), .ZN(n29346) );
  AND2_X1 U29351 ( .A1(b_0_), .A2(a_6_), .ZN(n29283) );
  OR2_X1 U29352 ( .A1(n29282), .A2(n29278), .ZN(n29345) );
  OR2_X1 U29353 ( .A1(n15706), .A2(n15841), .ZN(n29278) );
  INV_X1 U29354 ( .A(a_5_), .ZN(n15706) );
  OR2_X1 U29355 ( .A1(n29347), .A2(n29348), .ZN(n29282) );
  AND2_X1 U29356 ( .A1(n29268), .A2(n29272), .ZN(n29348) );
  AND2_X1 U29357 ( .A1(n29349), .A2(n29350), .ZN(n29347) );
  INV_X1 U29358 ( .A(n29273), .ZN(n29350) );
  AND2_X1 U29359 ( .A1(b_0_), .A2(a_7_), .ZN(n29273) );
  OR2_X1 U29360 ( .A1(n29272), .A2(n29268), .ZN(n29349) );
  OR2_X1 U29361 ( .A1(n15672), .A2(n15841), .ZN(n29268) );
  INV_X1 U29362 ( .A(a_6_), .ZN(n15672) );
  OR2_X1 U29363 ( .A1(n29351), .A2(n29352), .ZN(n29272) );
  AND2_X1 U29364 ( .A1(n29258), .A2(n29262), .ZN(n29352) );
  AND2_X1 U29365 ( .A1(n29353), .A2(n29354), .ZN(n29351) );
  INV_X1 U29366 ( .A(n29263), .ZN(n29354) );
  AND2_X1 U29367 ( .A1(b_0_), .A2(a_8_), .ZN(n29263) );
  OR2_X1 U29368 ( .A1(n29262), .A2(n29258), .ZN(n29353) );
  OR2_X1 U29369 ( .A1(n15638), .A2(n15841), .ZN(n29258) );
  INV_X1 U29370 ( .A(a_7_), .ZN(n15638) );
  OR2_X1 U29371 ( .A1(n29355), .A2(n29356), .ZN(n29262) );
  AND2_X1 U29372 ( .A1(n29248), .A2(n29252), .ZN(n29356) );
  AND2_X1 U29373 ( .A1(n29357), .A2(n29358), .ZN(n29355) );
  INV_X1 U29374 ( .A(n29253), .ZN(n29358) );
  AND2_X1 U29375 ( .A1(b_0_), .A2(a_9_), .ZN(n29253) );
  OR2_X1 U29376 ( .A1(n29252), .A2(n29248), .ZN(n29357) );
  OR2_X1 U29377 ( .A1(n15593), .A2(n15841), .ZN(n29248) );
  INV_X1 U29378 ( .A(a_8_), .ZN(n15593) );
  OR2_X1 U29379 ( .A1(n29359), .A2(n29360), .ZN(n29252) );
  AND2_X1 U29380 ( .A1(n29237), .A2(n29243), .ZN(n29360) );
  AND2_X1 U29381 ( .A1(n29361), .A2(n29241), .ZN(n29359) );
  OR2_X1 U29382 ( .A1(n16294), .A2(n15525), .ZN(n29241) );
  INV_X1 U29383 ( .A(a_10_), .ZN(n15525) );
  OR2_X1 U29384 ( .A1(n29243), .A2(n29237), .ZN(n29361) );
  OR2_X1 U29385 ( .A1(n29362), .A2(n29363), .ZN(n29237) );
  AND2_X1 U29386 ( .A1(n29226), .A2(n29232), .ZN(n29363) );
  AND2_X1 U29387 ( .A1(n29364), .A2(n29230), .ZN(n29362) );
  OR2_X1 U29388 ( .A1(n16294), .A2(n15491), .ZN(n29230) );
  INV_X1 U29389 ( .A(a_11_), .ZN(n15491) );
  OR2_X1 U29390 ( .A1(n29232), .A2(n29226), .ZN(n29364) );
  OR2_X1 U29391 ( .A1(n29365), .A2(n29366), .ZN(n29226) );
  AND2_X1 U29392 ( .A1(n29215), .A2(n29221), .ZN(n29366) );
  AND2_X1 U29393 ( .A1(n29367), .A2(n29219), .ZN(n29365) );
  OR2_X1 U29394 ( .A1(n16294), .A2(n15457), .ZN(n29219) );
  INV_X1 U29395 ( .A(a_12_), .ZN(n15457) );
  OR2_X1 U29396 ( .A1(n29221), .A2(n29215), .ZN(n29367) );
  OR2_X1 U29397 ( .A1(n29368), .A2(n29369), .ZN(n29215) );
  AND2_X1 U29398 ( .A1(n29204), .A2(n29210), .ZN(n29369) );
  AND2_X1 U29399 ( .A1(n29370), .A2(n29208), .ZN(n29368) );
  OR2_X1 U29400 ( .A1(n16294), .A2(n15423), .ZN(n29208) );
  INV_X1 U29401 ( .A(a_13_), .ZN(n15423) );
  OR2_X1 U29402 ( .A1(n29210), .A2(n29204), .ZN(n29370) );
  OR2_X1 U29403 ( .A1(n29371), .A2(n29372), .ZN(n29204) );
  AND2_X1 U29404 ( .A1(n29193), .A2(n29199), .ZN(n29372) );
  AND2_X1 U29405 ( .A1(n29373), .A2(n29197), .ZN(n29371) );
  OR2_X1 U29406 ( .A1(n16294), .A2(n15389), .ZN(n29197) );
  INV_X1 U29407 ( .A(a_14_), .ZN(n15389) );
  OR2_X1 U29408 ( .A1(n29199), .A2(n29193), .ZN(n29373) );
  OR2_X1 U29409 ( .A1(n29374), .A2(n29375), .ZN(n29193) );
  AND2_X1 U29410 ( .A1(n29182), .A2(n29188), .ZN(n29375) );
  AND2_X1 U29411 ( .A1(n29376), .A2(n29186), .ZN(n29374) );
  OR2_X1 U29412 ( .A1(n16294), .A2(n15355), .ZN(n29186) );
  INV_X1 U29413 ( .A(a_15_), .ZN(n15355) );
  OR2_X1 U29414 ( .A1(n29188), .A2(n29182), .ZN(n29376) );
  OR2_X1 U29415 ( .A1(n29377), .A2(n29378), .ZN(n29182) );
  AND2_X1 U29416 ( .A1(n29171), .A2(n29177), .ZN(n29378) );
  AND2_X1 U29417 ( .A1(n29379), .A2(n29175), .ZN(n29377) );
  OR2_X1 U29418 ( .A1(n16294), .A2(n15321), .ZN(n29175) );
  INV_X1 U29419 ( .A(a_16_), .ZN(n15321) );
  OR2_X1 U29420 ( .A1(n29177), .A2(n29171), .ZN(n29379) );
  OR2_X1 U29421 ( .A1(n29380), .A2(n29381), .ZN(n29171) );
  AND2_X1 U29422 ( .A1(n29160), .A2(n29166), .ZN(n29381) );
  AND2_X1 U29423 ( .A1(n29382), .A2(n29164), .ZN(n29380) );
  OR2_X1 U29424 ( .A1(n16294), .A2(n15287), .ZN(n29164) );
  INV_X1 U29425 ( .A(a_17_), .ZN(n15287) );
  OR2_X1 U29426 ( .A1(n29166), .A2(n29160), .ZN(n29382) );
  OR2_X1 U29427 ( .A1(n29383), .A2(n29384), .ZN(n29160) );
  AND2_X1 U29428 ( .A1(n29149), .A2(n29155), .ZN(n29384) );
  AND2_X1 U29429 ( .A1(n29385), .A2(n29153), .ZN(n29383) );
  OR2_X1 U29430 ( .A1(n16294), .A2(n15242), .ZN(n29153) );
  INV_X1 U29431 ( .A(a_18_), .ZN(n15242) );
  OR2_X1 U29432 ( .A1(n29155), .A2(n29149), .ZN(n29385) );
  OR2_X1 U29433 ( .A1(n29386), .A2(n29387), .ZN(n29149) );
  AND2_X1 U29434 ( .A1(n29138), .A2(n29144), .ZN(n29387) );
  AND2_X1 U29435 ( .A1(n29388), .A2(n29142), .ZN(n29386) );
  OR2_X1 U29436 ( .A1(n16294), .A2(n15208), .ZN(n29142) );
  INV_X1 U29437 ( .A(a_19_), .ZN(n15208) );
  OR2_X1 U29438 ( .A1(n29144), .A2(n29138), .ZN(n29388) );
  OR2_X1 U29439 ( .A1(n29389), .A2(n29390), .ZN(n29138) );
  AND2_X1 U29440 ( .A1(n29127), .A2(n29133), .ZN(n29390) );
  AND2_X1 U29441 ( .A1(n29391), .A2(n29131), .ZN(n29389) );
  OR2_X1 U29442 ( .A1(n16294), .A2(n15174), .ZN(n29131) );
  INV_X1 U29443 ( .A(a_20_), .ZN(n15174) );
  OR2_X1 U29444 ( .A1(n29133), .A2(n29127), .ZN(n29391) );
  OR2_X1 U29445 ( .A1(n29392), .A2(n29393), .ZN(n29127) );
  AND2_X1 U29446 ( .A1(n29116), .A2(n29122), .ZN(n29393) );
  AND2_X1 U29447 ( .A1(n29394), .A2(n29120), .ZN(n29392) );
  OR2_X1 U29448 ( .A1(n16294), .A2(n15140), .ZN(n29120) );
  INV_X1 U29449 ( .A(a_21_), .ZN(n15140) );
  OR2_X1 U29450 ( .A1(n29122), .A2(n29116), .ZN(n29394) );
  OR2_X1 U29451 ( .A1(n29395), .A2(n29396), .ZN(n29116) );
  AND2_X1 U29452 ( .A1(n29105), .A2(n29111), .ZN(n29396) );
  AND2_X1 U29453 ( .A1(n29397), .A2(n29109), .ZN(n29395) );
  OR2_X1 U29454 ( .A1(n16294), .A2(n15106), .ZN(n29109) );
  INV_X1 U29455 ( .A(a_22_), .ZN(n15106) );
  OR2_X1 U29456 ( .A1(n29111), .A2(n29105), .ZN(n29397) );
  OR2_X1 U29457 ( .A1(n29398), .A2(n29399), .ZN(n29105) );
  AND2_X1 U29458 ( .A1(n29094), .A2(n29100), .ZN(n29399) );
  AND2_X1 U29459 ( .A1(n29400), .A2(n29098), .ZN(n29398) );
  OR2_X1 U29460 ( .A1(n16294), .A2(n15072), .ZN(n29098) );
  INV_X1 U29461 ( .A(a_23_), .ZN(n15072) );
  OR2_X1 U29462 ( .A1(n29100), .A2(n29094), .ZN(n29400) );
  OR2_X1 U29463 ( .A1(n29401), .A2(n29402), .ZN(n29094) );
  AND2_X1 U29464 ( .A1(n29083), .A2(n29089), .ZN(n29402) );
  AND2_X1 U29465 ( .A1(n29403), .A2(n29087), .ZN(n29401) );
  OR2_X1 U29466 ( .A1(n16294), .A2(n15038), .ZN(n29087) );
  INV_X1 U29467 ( .A(a_24_), .ZN(n15038) );
  OR2_X1 U29468 ( .A1(n29089), .A2(n29083), .ZN(n29403) );
  OR2_X1 U29469 ( .A1(n29404), .A2(n29405), .ZN(n29083) );
  AND2_X1 U29470 ( .A1(n29072), .A2(n29078), .ZN(n29405) );
  AND2_X1 U29471 ( .A1(n29406), .A2(n29076), .ZN(n29404) );
  OR2_X1 U29472 ( .A1(n16294), .A2(n15004), .ZN(n29076) );
  INV_X1 U29473 ( .A(a_25_), .ZN(n15004) );
  OR2_X1 U29474 ( .A1(n29078), .A2(n29072), .ZN(n29406) );
  OR2_X1 U29475 ( .A1(n29407), .A2(n29408), .ZN(n29072) );
  AND2_X1 U29476 ( .A1(n29061), .A2(n29067), .ZN(n29408) );
  AND2_X1 U29477 ( .A1(n29409), .A2(n29065), .ZN(n29407) );
  OR2_X1 U29478 ( .A1(n16294), .A2(n14970), .ZN(n29065) );
  INV_X1 U29479 ( .A(a_26_), .ZN(n14970) );
  OR2_X1 U29480 ( .A1(n29067), .A2(n29061), .ZN(n29409) );
  OR2_X1 U29481 ( .A1(n29410), .A2(n29411), .ZN(n29061) );
  AND2_X1 U29482 ( .A1(n29050), .A2(n29056), .ZN(n29411) );
  AND2_X1 U29483 ( .A1(n29412), .A2(n29054), .ZN(n29410) );
  OR2_X1 U29484 ( .A1(n16294), .A2(n14936), .ZN(n29054) );
  INV_X1 U29485 ( .A(a_27_), .ZN(n14936) );
  OR2_X1 U29486 ( .A1(n29056), .A2(n29050), .ZN(n29412) );
  OR2_X1 U29487 ( .A1(n29413), .A2(n29414), .ZN(n29050) );
  AND2_X1 U29488 ( .A1(n29039), .A2(n29045), .ZN(n29414) );
  AND2_X1 U29489 ( .A1(n29415), .A2(n29043), .ZN(n29413) );
  OR2_X1 U29490 ( .A1(n16294), .A2(n14891), .ZN(n29043) );
  OR2_X1 U29491 ( .A1(n29045), .A2(n29039), .ZN(n29415) );
  OR2_X1 U29492 ( .A1(n29416), .A2(n29417), .ZN(n29039) );
  AND2_X1 U29493 ( .A1(n29032), .A2(n29418), .ZN(n29417) );
  AND2_X1 U29494 ( .A1(n29029), .A2(n29419), .ZN(n29416) );
  OR2_X1 U29495 ( .A1(n29418), .A2(n29032), .ZN(n29419) );
  OR2_X1 U29496 ( .A1(n14891), .A2(n15841), .ZN(n29032) );
  INV_X1 U29497 ( .A(n29027), .ZN(n29029) );
  OR2_X1 U29498 ( .A1(n29420), .A2(n29019), .ZN(n29027) );
  AND3_X1 U29499 ( .A1(b_0_), .A2(b_1_), .A3(n15957), .ZN(n29019) );
  AND2_X1 U29500 ( .A1(a_31_), .A2(a_30_), .ZN(n15957) );
  AND3_X1 U29501 ( .A1(b_1_), .A2(a_30_), .A3(n29033), .ZN(n29420) );
  INV_X1 U29502 ( .A(n29418), .ZN(n29033) );
  OR2_X1 U29503 ( .A1(n16294), .A2(n14857), .ZN(n29418) );
  INV_X1 U29504 ( .A(a_29_), .ZN(n14857) );
  INV_X1 U29505 ( .A(b_0_), .ZN(n16294) );
  INV_X1 U29506 ( .A(n29042), .ZN(n29045) );
  AND2_X1 U29507 ( .A1(a_27_), .A2(b_1_), .ZN(n29042) );
  INV_X1 U29508 ( .A(n29053), .ZN(n29056) );
  AND2_X1 U29509 ( .A1(a_26_), .A2(b_1_), .ZN(n29053) );
  INV_X1 U29510 ( .A(n29064), .ZN(n29067) );
  AND2_X1 U29511 ( .A1(a_25_), .A2(b_1_), .ZN(n29064) );
  INV_X1 U29512 ( .A(n29075), .ZN(n29078) );
  AND2_X1 U29513 ( .A1(a_24_), .A2(b_1_), .ZN(n29075) );
  INV_X1 U29514 ( .A(n29086), .ZN(n29089) );
  AND2_X1 U29515 ( .A1(a_23_), .A2(b_1_), .ZN(n29086) );
  INV_X1 U29516 ( .A(n29097), .ZN(n29100) );
  AND2_X1 U29517 ( .A1(a_22_), .A2(b_1_), .ZN(n29097) );
  INV_X1 U29518 ( .A(n29108), .ZN(n29111) );
  AND2_X1 U29519 ( .A1(a_21_), .A2(b_1_), .ZN(n29108) );
  INV_X1 U29520 ( .A(n29119), .ZN(n29122) );
  AND2_X1 U29521 ( .A1(a_20_), .A2(b_1_), .ZN(n29119) );
  INV_X1 U29522 ( .A(n29130), .ZN(n29133) );
  AND2_X1 U29523 ( .A1(a_19_), .A2(b_1_), .ZN(n29130) );
  INV_X1 U29524 ( .A(n29141), .ZN(n29144) );
  AND2_X1 U29525 ( .A1(a_18_), .A2(b_1_), .ZN(n29141) );
  INV_X1 U29526 ( .A(n29152), .ZN(n29155) );
  AND2_X1 U29527 ( .A1(a_17_), .A2(b_1_), .ZN(n29152) );
  INV_X1 U29528 ( .A(n29163), .ZN(n29166) );
  AND2_X1 U29529 ( .A1(a_16_), .A2(b_1_), .ZN(n29163) );
  INV_X1 U29530 ( .A(n29174), .ZN(n29177) );
  AND2_X1 U29531 ( .A1(a_15_), .A2(b_1_), .ZN(n29174) );
  INV_X1 U29532 ( .A(n29185), .ZN(n29188) );
  AND2_X1 U29533 ( .A1(a_14_), .A2(b_1_), .ZN(n29185) );
  INV_X1 U29534 ( .A(n29196), .ZN(n29199) );
  AND2_X1 U29535 ( .A1(a_13_), .A2(b_1_), .ZN(n29196) );
  INV_X1 U29536 ( .A(n29207), .ZN(n29210) );
  AND2_X1 U29537 ( .A1(a_12_), .A2(b_1_), .ZN(n29207) );
  INV_X1 U29538 ( .A(n29218), .ZN(n29221) );
  AND2_X1 U29539 ( .A1(a_11_), .A2(b_1_), .ZN(n29218) );
  INV_X1 U29540 ( .A(n29229), .ZN(n29232) );
  AND2_X1 U29541 ( .A1(a_10_), .A2(b_1_), .ZN(n29229) );
  INV_X1 U29542 ( .A(n29240), .ZN(n29243) );
  AND2_X1 U29543 ( .A1(a_9_), .A2(b_1_), .ZN(n29240) );
  OR2_X1 U29544 ( .A1(n29421), .A2(n29422), .ZN(n29327) );
  AND2_X1 U29545 ( .A1(n29423), .A2(n28918), .ZN(n29422) );
  AND2_X1 U29546 ( .A1(n29424), .A2(n28916), .ZN(n29421) );
  INV_X1 U29547 ( .A(n29423), .ZN(n28916) );
  AND2_X1 U29548 ( .A1(b_0_), .A2(a_1_), .ZN(n29423) );
  INV_X1 U29549 ( .A(n28918), .ZN(n29424) );
  OR2_X1 U29550 ( .A1(n16512), .A2(n15841), .ZN(n28918) );
  INV_X1 U29551 ( .A(b_1_), .ZN(n15841) );
  INV_X1 U29552 ( .A(a_0_), .ZN(n16512) );
endmodule

