module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n641_, new_n339_, new_n365_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n456_, new_n246_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n642_, new_n211_, new_n552_, new_n342_, new_n649_, new_n462_, new_n603_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n257_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n297_, new_n361_, new_n565_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n524_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n346_, new_n396_, new_n198_, new_n208_, new_n632_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n562_, new_n485_, new_n578_, new_n525_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n605_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n662_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n151_, N75 );
nand g001 ( new_n152_, N29, N42 );
nor g002 ( N388, new_n152_, new_n151_ );
not g003 ( new_n154_, N80 );
nand g004 ( new_n155_, N29, N36 );
nor g005 ( N389, new_n155_, new_n154_ );
not g006 ( new_n157_, N42 );
nor g007 ( N390, new_n155_, new_n157_ );
and g008 ( N391, N85, N86 );
not g009 ( new_n160_, N13 );
nand g010 ( new_n161_, N1, N8 );
nor g011 ( new_n162_, new_n161_, new_n160_ );
and g012 ( N418, new_n162_, N17 );
not g013 ( new_n164_, N390 );
nand g014 ( new_n165_, N1, N26 );
nand g015 ( new_n166_, N13, N17 );
nor g016 ( new_n167_, new_n165_, new_n166_ );
nand g017 ( N419, new_n164_, new_n167_ );
and g018 ( new_n169_, N59, N75 );
nand g019 ( N420, new_n169_, N80 );
and g020 ( new_n171_, N36, N59 );
nand g021 ( N421, new_n171_, N80 );
nand g022 ( N422, new_n171_, N42 );
not g023 ( new_n174_, N90 );
nor g024 ( new_n175_, N87, N88 );
nor g025 ( N423, new_n175_, new_n174_ );
nand g026 ( N446, new_n167_, N390 );
not g027 ( new_n178_, N51 );
nor g028 ( new_n179_, new_n165_, new_n178_ );
xnor g029 ( N447, new_n179_, keyIn_0_0 );
nand g030 ( new_n181_, new_n162_, N55 );
nand g031 ( new_n182_, N29, N68 );
nor g032 ( N448, new_n181_, new_n182_ );
and g033 ( new_n184_, N59, N68 );
nand g034 ( new_n185_, new_n184_, N74 );
nor g035 ( N449, new_n181_, new_n185_ );
not g036 ( new_n187_, N89 );
nor g037 ( N450, new_n175_, new_n187_ );
xor g038 ( new_n189_, N111, N116 );
xnor g039 ( new_n190_, N121, N126 );
xnor g040 ( new_n191_, new_n189_, new_n190_ );
xnor g041 ( new_n192_, new_n191_, N135 );
xnor g042 ( new_n193_, N91, N96 );
xnor g043 ( new_n194_, N101, N106 );
xnor g044 ( new_n195_, new_n193_, new_n194_ );
xnor g045 ( new_n196_, new_n195_, N130 );
xnor g046 ( N767, new_n192_, new_n196_ );
xor g047 ( new_n198_, N183, N189 );
xnor g048 ( new_n199_, N195, N201 );
xnor g049 ( new_n200_, new_n198_, new_n199_ );
xnor g050 ( new_n201_, new_n200_, N207 );
xnor g051 ( new_n202_, N159, N165 );
xnor g052 ( new_n203_, N171, N177 );
xnor g053 ( new_n204_, new_n202_, new_n203_ );
xnor g054 ( new_n205_, new_n204_, N130 );
xnor g055 ( N768, new_n201_, new_n205_ );
not g056 ( new_n207_, N261 );
not g057 ( new_n208_, N201 );
not g058 ( new_n209_, keyIn_0_37 );
not g059 ( new_n210_, keyIn_0_31 );
not g060 ( new_n211_, keyIn_0_19 );
not g061 ( new_n212_, keyIn_0_8 );
and g062 ( new_n213_, N1, N26 );
nand g063 ( new_n214_, new_n213_, N51 );
nand g064 ( new_n215_, new_n214_, keyIn_0_0 );
not g065 ( new_n216_, keyIn_0_0 );
nand g066 ( new_n217_, new_n179_, new_n216_ );
nand g067 ( new_n218_, new_n215_, new_n217_ );
nand g068 ( new_n219_, new_n218_, new_n212_ );
nand g069 ( new_n220_, N447, keyIn_0_8 );
nand g070 ( new_n221_, new_n220_, new_n219_ );
nand g071 ( new_n222_, new_n221_, keyIn_0_14 );
not g072 ( new_n223_, keyIn_0_14 );
xnor g073 ( new_n224_, new_n218_, keyIn_0_8 );
nand g074 ( new_n225_, new_n224_, new_n223_ );
nand g075 ( new_n226_, new_n225_, new_n222_ );
not g076 ( new_n227_, keyIn_0_13 );
nor g077 ( new_n228_, N17, N42 );
xnor g078 ( new_n229_, new_n228_, keyIn_0_6 );
nand g079 ( new_n230_, N17, N42 );
xnor g080 ( new_n231_, new_n230_, keyIn_0_7 );
nand g081 ( new_n232_, new_n229_, new_n231_ );
nor g082 ( new_n233_, new_n232_, new_n227_ );
nand g083 ( new_n234_, N59, N156 );
not g084 ( new_n235_, new_n234_ );
nand g085 ( new_n236_, new_n232_, new_n227_ );
nand g086 ( new_n237_, new_n236_, new_n235_ );
nor g087 ( new_n238_, new_n237_, new_n233_ );
nand g088 ( new_n239_, new_n226_, new_n238_ );
nor g089 ( new_n240_, new_n239_, new_n211_ );
not g090 ( new_n241_, new_n240_ );
nand g091 ( new_n242_, new_n239_, new_n211_ );
not g092 ( new_n243_, keyIn_0_9 );
not g093 ( new_n244_, keyIn_0_1 );
nand g094 ( new_n245_, N17, N51 );
nor g095 ( new_n246_, new_n161_, new_n245_ );
xnor g096 ( new_n247_, new_n246_, new_n244_ );
xnor g097 ( new_n248_, new_n247_, new_n243_ );
not g098 ( new_n249_, keyIn_0_11 );
not g099 ( new_n250_, keyIn_0_3 );
nand g100 ( new_n251_, N42, N59 );
nor g101 ( new_n252_, new_n251_, new_n151_ );
xnor g102 ( new_n253_, new_n252_, new_n250_ );
xnor g103 ( new_n254_, new_n253_, new_n249_ );
nand g104 ( new_n255_, new_n248_, new_n254_ );
nand g105 ( new_n256_, new_n255_, keyIn_0_15 );
not g106 ( new_n257_, keyIn_0_15 );
xnor g107 ( new_n258_, new_n247_, keyIn_0_9 );
xnor g108 ( new_n259_, new_n253_, keyIn_0_11 );
nor g109 ( new_n260_, new_n258_, new_n259_ );
nand g110 ( new_n261_, new_n260_, new_n257_ );
nand g111 ( new_n262_, new_n261_, new_n256_ );
and g112 ( new_n263_, new_n242_, new_n262_ );
nand g113 ( new_n264_, new_n263_, new_n241_ );
nand g114 ( new_n265_, new_n264_, keyIn_0_21 );
not g115 ( new_n266_, keyIn_0_21 );
nand g116 ( new_n267_, new_n242_, new_n262_ );
nor g117 ( new_n268_, new_n267_, new_n240_ );
nand g118 ( new_n269_, new_n268_, new_n266_ );
nand g119 ( new_n270_, new_n265_, new_n269_ );
nand g120 ( new_n271_, new_n270_, N126 );
nor g121 ( new_n272_, new_n271_, new_n210_ );
nand g122 ( new_n273_, new_n271_, new_n210_ );
not g123 ( new_n274_, keyIn_0_24 );
not g124 ( new_n275_, keyIn_0_20 );
not g125 ( new_n276_, N17 );
xor g126 ( new_n277_, new_n234_, keyIn_0_5 );
nor g127 ( new_n278_, new_n277_, new_n276_ );
nand g128 ( new_n279_, new_n226_, new_n278_ );
nor g129 ( new_n280_, new_n279_, new_n275_ );
nand g130 ( new_n281_, new_n279_, new_n275_ );
nand g131 ( new_n282_, new_n281_, N1 );
nor g132 ( new_n283_, new_n282_, new_n280_ );
xnor g133 ( new_n284_, new_n283_, new_n274_ );
nand g134 ( new_n285_, new_n284_, N153 );
nand g135 ( new_n286_, new_n273_, new_n285_ );
nor g136 ( new_n287_, new_n286_, new_n272_ );
xnor g137 ( new_n288_, new_n287_, new_n209_ );
not g138 ( new_n289_, N55 );
nand g139 ( new_n290_, N29, N75 );
nor g140 ( new_n291_, new_n290_, new_n154_ );
xnor g141 ( new_n292_, new_n291_, keyIn_0_2 );
nand g142 ( new_n293_, new_n226_, new_n292_ );
nor g143 ( new_n294_, new_n293_, new_n289_ );
nand g144 ( new_n295_, new_n294_, keyIn_0_18 );
xnor g145 ( new_n296_, keyIn_0_4, N268 );
xnor g146 ( new_n297_, new_n296_, keyIn_0_12 );
nor g147 ( new_n298_, new_n294_, keyIn_0_18 );
nor g148 ( new_n299_, new_n298_, new_n297_ );
nand g149 ( new_n300_, new_n299_, new_n295_ );
xor g150 ( new_n301_, new_n300_, keyIn_0_28 );
not g151 ( new_n302_, new_n301_ );
nand g152 ( new_n303_, new_n288_, new_n302_ );
nand g153 ( new_n304_, new_n303_, keyIn_0_43 );
not g154 ( new_n305_, keyIn_0_43 );
xnor g155 ( new_n306_, new_n287_, keyIn_0_37 );
nor g156 ( new_n307_, new_n306_, new_n301_ );
nand g157 ( new_n308_, new_n307_, new_n305_ );
nand g158 ( new_n309_, new_n308_, new_n304_ );
nand g159 ( new_n310_, new_n309_, new_n208_ );
nor g160 ( new_n311_, new_n309_, new_n208_ );
not g161 ( new_n312_, new_n311_ );
nand g162 ( new_n313_, new_n312_, new_n310_ );
and g163 ( new_n314_, new_n313_, new_n207_ );
and g164 ( new_n315_, new_n310_, N261 );
nand g165 ( new_n316_, new_n315_, new_n312_ );
nand g166 ( new_n317_, new_n316_, N219 );
nor g167 ( new_n318_, new_n317_, new_n314_ );
not g168 ( new_n319_, N228 );
or g169 ( new_n320_, new_n313_, new_n319_ );
not g170 ( new_n321_, N237 );
nor g171 ( new_n322_, new_n312_, new_n321_ );
not g172 ( new_n323_, N246 );
or g173 ( new_n324_, new_n309_, new_n323_ );
and g174 ( new_n325_, N42, N72 );
nand g175 ( new_n326_, new_n184_, new_n325_ );
nor g176 ( new_n327_, new_n181_, new_n326_ );
nor g177 ( new_n328_, new_n327_, keyIn_0_10 );
nand g178 ( new_n329_, new_n327_, keyIn_0_10 );
nand g179 ( new_n330_, new_n329_, N73 );
nor g180 ( new_n331_, new_n330_, new_n328_ );
and g181 ( new_n332_, new_n331_, N201 );
nand g182 ( new_n333_, N255, N267 );
nand g183 ( new_n334_, N121, N210 );
nand g184 ( new_n335_, new_n333_, new_n334_ );
nor g185 ( new_n336_, new_n332_, new_n335_ );
nand g186 ( new_n337_, new_n324_, new_n336_ );
nor g187 ( new_n338_, new_n322_, new_n337_ );
nand g188 ( new_n339_, new_n320_, new_n338_ );
nor g189 ( new_n340_, new_n318_, new_n339_ );
xor g190 ( N850, new_n340_, keyIn_0_52 );
nand g191 ( new_n342_, new_n284_, N143 );
nand g192 ( new_n343_, new_n270_, N111 );
nand g193 ( new_n344_, new_n342_, new_n343_ );
xnor g194 ( new_n345_, new_n344_, keyIn_0_34 );
xor g195 ( new_n346_, new_n300_, keyIn_0_25 );
nand g196 ( new_n347_, new_n345_, new_n346_ );
xnor g197 ( new_n348_, new_n347_, keyIn_0_40 );
nand g198 ( new_n349_, new_n348_, N183 );
not g199 ( new_n350_, new_n349_ );
not g200 ( new_n351_, keyIn_0_46 );
not g201 ( new_n352_, N195 );
not g202 ( new_n353_, keyIn_0_42 );
not g203 ( new_n354_, keyIn_0_36 );
nand g204 ( new_n355_, new_n270_, N121 );
nand g205 ( new_n356_, new_n284_, N149 );
nand g206 ( new_n357_, new_n356_, new_n355_ );
nor g207 ( new_n358_, new_n357_, new_n354_ );
not g208 ( new_n359_, new_n358_ );
xnor g209 ( new_n360_, new_n300_, keyIn_0_27 );
nand g210 ( new_n361_, new_n357_, new_n354_ );
and g211 ( new_n362_, new_n361_, new_n360_ );
nand g212 ( new_n363_, new_n362_, new_n359_ );
nand g213 ( new_n364_, new_n363_, new_n353_ );
nand g214 ( new_n365_, new_n361_, new_n360_ );
nor g215 ( new_n366_, new_n365_, new_n358_ );
nand g216 ( new_n367_, new_n366_, keyIn_0_42 );
nand g217 ( new_n368_, new_n364_, new_n367_ );
nand g218 ( new_n369_, new_n368_, new_n352_ );
not g219 ( new_n370_, N189 );
not g220 ( new_n371_, keyIn_0_41 );
nand g221 ( new_n372_, new_n270_, N116 );
nand g222 ( new_n373_, new_n284_, N146 );
nand g223 ( new_n374_, new_n373_, new_n372_ );
nor g224 ( new_n375_, new_n374_, keyIn_0_35 );
not g225 ( new_n376_, new_n375_ );
xor g226 ( new_n377_, new_n300_, keyIn_0_26 );
nand g227 ( new_n378_, new_n374_, keyIn_0_35 );
and g228 ( new_n379_, new_n378_, new_n377_ );
nand g229 ( new_n380_, new_n379_, new_n376_ );
nand g230 ( new_n381_, new_n380_, new_n371_ );
nand g231 ( new_n382_, new_n378_, new_n377_ );
nor g232 ( new_n383_, new_n382_, new_n375_ );
nand g233 ( new_n384_, new_n383_, keyIn_0_41 );
nand g234 ( new_n385_, new_n381_, new_n384_ );
nand g235 ( new_n386_, new_n385_, new_n370_ );
nand g236 ( new_n387_, new_n369_, new_n386_ );
not g237 ( new_n388_, new_n387_ );
nand g238 ( new_n389_, new_n311_, new_n388_ );
nor g239 ( new_n390_, new_n389_, new_n351_ );
nand g240 ( new_n391_, new_n389_, new_n351_ );
not g241 ( new_n392_, keyIn_0_45 );
nor g242 ( new_n393_, new_n368_, new_n352_ );
nand g243 ( new_n394_, new_n393_, new_n386_ );
nor g244 ( new_n395_, new_n394_, new_n392_ );
not g245 ( new_n396_, new_n385_ );
nand g246 ( new_n397_, new_n396_, N189 );
nand g247 ( new_n398_, new_n394_, new_n392_ );
nand g248 ( new_n399_, new_n398_, new_n397_ );
nor g249 ( new_n400_, new_n399_, new_n395_ );
nand g250 ( new_n401_, new_n391_, new_n400_ );
nor g251 ( new_n402_, new_n401_, new_n390_ );
not g252 ( new_n403_, keyIn_0_44 );
nand g253 ( new_n404_, new_n310_, N261 );
nor g254 ( new_n405_, new_n404_, new_n387_ );
xnor g255 ( new_n406_, new_n405_, new_n403_ );
nand g256 ( new_n407_, new_n406_, new_n402_ );
nand g257 ( new_n408_, new_n407_, keyIn_0_48 );
not g258 ( new_n409_, keyIn_0_48 );
not g259 ( new_n410_, new_n390_ );
and g260 ( new_n411_, new_n391_, new_n400_ );
nand g261 ( new_n412_, new_n411_, new_n410_ );
nand g262 ( new_n413_, new_n315_, new_n388_ );
nand g263 ( new_n414_, new_n413_, new_n403_ );
nand g264 ( new_n415_, new_n405_, keyIn_0_44 );
nand g265 ( new_n416_, new_n414_, new_n415_ );
nor g266 ( new_n417_, new_n412_, new_n416_ );
nand g267 ( new_n418_, new_n417_, new_n409_ );
nand g268 ( new_n419_, new_n418_, new_n408_ );
nor g269 ( new_n420_, new_n348_, N183 );
not g270 ( new_n421_, new_n420_ );
nand g271 ( new_n422_, new_n419_, new_n421_ );
nor g272 ( new_n423_, new_n422_, new_n350_ );
nor g273 ( new_n424_, new_n350_, new_n420_ );
or g274 ( new_n425_, new_n419_, new_n424_ );
nand g275 ( new_n426_, new_n425_, N219 );
nor g276 ( new_n427_, new_n426_, new_n423_ );
nand g277 ( new_n428_, new_n424_, N228 );
nor g278 ( new_n429_, new_n349_, new_n321_ );
nand g279 ( new_n430_, new_n348_, N246 );
nand g280 ( new_n431_, N106, N210 );
nand g281 ( new_n432_, new_n331_, N183 );
and g282 ( new_n433_, new_n432_, new_n431_ );
nand g283 ( new_n434_, new_n430_, new_n433_ );
nor g284 ( new_n435_, new_n429_, new_n434_ );
nand g285 ( new_n436_, new_n428_, new_n435_ );
nor g286 ( new_n437_, new_n427_, new_n436_ );
xnor g287 ( N863, new_n437_, keyIn_0_57 );
not g288 ( new_n439_, new_n393_ );
nand g289 ( new_n440_, new_n404_, new_n312_ );
nand g290 ( new_n441_, new_n440_, new_n369_ );
nand g291 ( new_n442_, new_n441_, new_n439_ );
xor g292 ( new_n443_, new_n442_, keyIn_0_49 );
nand g293 ( new_n444_, new_n397_, new_n386_ );
nor g294 ( new_n445_, new_n443_, new_n444_ );
nand g295 ( new_n446_, new_n443_, new_n444_ );
nand g296 ( new_n447_, new_n446_, N219 );
nor g297 ( new_n448_, new_n447_, new_n445_ );
or g298 ( new_n449_, new_n444_, new_n319_ );
nor g299 ( new_n450_, new_n397_, new_n321_ );
nand g300 ( new_n451_, new_n396_, N246 );
and g301 ( new_n452_, new_n331_, N189 );
nand g302 ( new_n453_, N255, N259 );
nand g303 ( new_n454_, N111, N210 );
nand g304 ( new_n455_, new_n453_, new_n454_ );
nor g305 ( new_n456_, new_n452_, new_n455_ );
nand g306 ( new_n457_, new_n451_, new_n456_ );
nor g307 ( new_n458_, new_n450_, new_n457_ );
nand g308 ( new_n459_, new_n449_, new_n458_ );
nor g309 ( new_n460_, new_n448_, new_n459_ );
xor g310 ( N864, new_n460_, keyIn_0_58 );
or g311 ( new_n462_, new_n441_, new_n393_ );
not g312 ( new_n463_, N219 );
nand g313 ( new_n464_, new_n439_, new_n369_ );
not g314 ( new_n465_, new_n464_ );
nor g315 ( new_n466_, new_n440_, new_n465_ );
nor g316 ( new_n467_, new_n466_, new_n463_ );
nand g317 ( new_n468_, new_n462_, new_n467_ );
nor g318 ( new_n469_, new_n464_, new_n319_ );
nand g319 ( new_n470_, new_n393_, N237 );
nor g320 ( new_n471_, new_n368_, new_n323_ );
nand g321 ( new_n472_, new_n331_, N195 );
nand g322 ( new_n473_, N255, N260 );
nand g323 ( new_n474_, N116, N210 );
and g324 ( new_n475_, new_n473_, new_n474_ );
nand g325 ( new_n476_, new_n472_, new_n475_ );
nor g326 ( new_n477_, new_n471_, new_n476_ );
nand g327 ( new_n478_, new_n477_, new_n470_ );
nor g328 ( new_n479_, new_n469_, new_n478_ );
nand g329 ( new_n480_, new_n468_, new_n479_ );
xnor g330 ( N865, new_n480_, keyIn_0_59 );
nand g331 ( new_n482_, new_n270_, N91 );
nor g332 ( new_n483_, new_n293_, new_n276_ );
nor g333 ( new_n484_, new_n483_, keyIn_0_17 );
nand g334 ( new_n485_, new_n483_, keyIn_0_17 );
nand g335 ( new_n486_, new_n485_, new_n296_ );
nor g336 ( new_n487_, new_n486_, new_n484_ );
nand g337 ( new_n488_, N8, N138 );
nor g338 ( new_n489_, new_n277_, new_n289_ );
nand g339 ( new_n490_, new_n226_, new_n489_ );
xnor g340 ( new_n491_, new_n490_, keyIn_0_16 );
nand g341 ( new_n492_, new_n491_, N143 );
nand g342 ( new_n493_, new_n492_, new_n488_ );
nor g343 ( new_n494_, new_n493_, new_n487_ );
nand g344 ( new_n495_, new_n482_, new_n494_ );
nand g345 ( new_n496_, new_n495_, N159 );
or g346 ( new_n497_, new_n495_, N159 );
not g347 ( new_n498_, keyIn_0_51 );
not g348 ( new_n499_, keyIn_0_50 );
xnor g349 ( new_n500_, new_n422_, new_n499_ );
nand g350 ( new_n501_, new_n500_, new_n349_ );
nand g351 ( new_n502_, new_n501_, new_n498_ );
xnor g352 ( new_n503_, new_n422_, keyIn_0_50 );
nor g353 ( new_n504_, new_n503_, new_n350_ );
nand g354 ( new_n505_, new_n504_, keyIn_0_51 );
nand g355 ( new_n506_, new_n505_, new_n502_ );
xor g356 ( new_n507_, new_n487_, keyIn_0_22 );
nand g357 ( new_n508_, new_n491_, N149 );
nand g358 ( new_n509_, new_n507_, new_n508_ );
xnor g359 ( new_n510_, new_n509_, keyIn_0_29 );
nand g360 ( new_n511_, new_n270_, N101 );
nand g361 ( new_n512_, N17, N138 );
nand g362 ( new_n513_, new_n511_, new_n512_ );
xnor g363 ( new_n514_, new_n513_, keyIn_0_32 );
nand g364 ( new_n515_, new_n510_, new_n514_ );
xor g365 ( new_n516_, new_n515_, keyIn_0_38 );
nor g366 ( new_n517_, new_n516_, N171 );
nand g367 ( new_n518_, new_n270_, N96 );
nand g368 ( new_n519_, N51, N138 );
nand g369 ( new_n520_, new_n491_, N146 );
nand g370 ( new_n521_, new_n520_, new_n519_ );
nor g371 ( new_n522_, new_n521_, new_n487_ );
nand g372 ( new_n523_, new_n518_, new_n522_ );
nor g373 ( new_n524_, new_n523_, N165 );
nor g374 ( new_n525_, new_n517_, new_n524_ );
not g375 ( new_n526_, new_n525_ );
xnor g376 ( new_n527_, new_n487_, keyIn_0_23 );
nand g377 ( new_n528_, new_n491_, N153 );
nand g378 ( new_n529_, new_n527_, new_n528_ );
xor g379 ( new_n530_, new_n529_, keyIn_0_30 );
nand g380 ( new_n531_, new_n270_, N106 );
nand g381 ( new_n532_, N138, N152 );
nand g382 ( new_n533_, new_n531_, new_n532_ );
xnor g383 ( new_n534_, new_n533_, keyIn_0_33 );
nand g384 ( new_n535_, new_n530_, new_n534_ );
xor g385 ( new_n536_, new_n535_, keyIn_0_39 );
nor g386 ( new_n537_, new_n536_, N177 );
nor g387 ( new_n538_, new_n526_, new_n537_ );
nand g388 ( new_n539_, new_n506_, new_n538_ );
nor g389 ( new_n540_, new_n539_, keyIn_0_54 );
not g390 ( new_n541_, new_n540_ );
nand g391 ( new_n542_, new_n539_, keyIn_0_54 );
nand g392 ( new_n543_, new_n536_, N177 );
nor g393 ( new_n544_, new_n526_, new_n543_ );
nor g394 ( new_n545_, new_n544_, keyIn_0_47 );
nand g395 ( new_n546_, new_n544_, keyIn_0_47 );
nand g396 ( new_n547_, new_n523_, N165 );
not g397 ( new_n548_, new_n547_ );
nand g398 ( new_n549_, new_n516_, N171 );
nor g399 ( new_n550_, new_n549_, new_n524_ );
nor g400 ( new_n551_, new_n550_, new_n548_ );
nand g401 ( new_n552_, new_n546_, new_n551_ );
nor g402 ( new_n553_, new_n552_, new_n545_ );
and g403 ( new_n554_, new_n542_, new_n553_ );
nand g404 ( new_n555_, new_n554_, new_n541_ );
nand g405 ( new_n556_, new_n555_, keyIn_0_55 );
not g406 ( new_n557_, keyIn_0_55 );
nand g407 ( new_n558_, new_n542_, new_n553_ );
nor g408 ( new_n559_, new_n558_, new_n540_ );
nand g409 ( new_n560_, new_n559_, new_n557_ );
nand g410 ( new_n561_, new_n556_, new_n560_ );
not g411 ( new_n562_, new_n561_ );
nand g412 ( new_n563_, new_n562_, new_n497_ );
nand g413 ( N866, new_n563_, new_n496_ );
not g414 ( new_n565_, new_n543_ );
not g415 ( new_n566_, new_n537_ );
nand g416 ( new_n567_, new_n506_, new_n566_ );
nor g417 ( new_n568_, new_n567_, new_n565_ );
nor g418 ( new_n569_, new_n565_, new_n537_ );
or g419 ( new_n570_, new_n506_, new_n569_ );
nand g420 ( new_n571_, new_n570_, N219 );
nor g421 ( new_n572_, new_n571_, new_n568_ );
nand g422 ( new_n573_, new_n569_, N228 );
nor g423 ( new_n574_, new_n543_, new_n321_ );
nand g424 ( new_n575_, new_n536_, N246 );
nand g425 ( new_n576_, N101, N210 );
nand g426 ( new_n577_, new_n331_, N177 );
and g427 ( new_n578_, new_n577_, new_n576_ );
nand g428 ( new_n579_, new_n575_, new_n578_ );
nor g429 ( new_n580_, new_n574_, new_n579_ );
nand g430 ( new_n581_, new_n573_, new_n580_ );
nor g431 ( new_n582_, new_n572_, new_n581_ );
xor g432 ( N874, new_n582_, keyIn_0_60 );
nand g433 ( new_n584_, new_n497_, new_n496_ );
nor g434 ( new_n585_, new_n561_, new_n584_ );
not g435 ( new_n586_, new_n585_ );
nand g436 ( new_n587_, new_n561_, new_n584_ );
and g437 ( new_n588_, new_n587_, N219 );
nand g438 ( new_n589_, new_n588_, new_n586_ );
nor g439 ( new_n590_, new_n584_, new_n319_ );
nor g440 ( new_n591_, new_n496_, new_n321_ );
nand g441 ( new_n592_, new_n495_, N246 );
nand g442 ( new_n593_, new_n297_, N210 );
nand g443 ( new_n594_, new_n331_, N159 );
and g444 ( new_n595_, new_n594_, new_n593_ );
nand g445 ( new_n596_, new_n592_, new_n595_ );
nor g446 ( new_n597_, new_n591_, new_n596_ );
not g447 ( new_n598_, new_n597_ );
nor g448 ( new_n599_, new_n598_, new_n590_ );
nand g449 ( new_n600_, new_n589_, new_n599_ );
nand g450 ( new_n601_, new_n600_, keyIn_0_61 );
not g451 ( new_n602_, keyIn_0_61 );
nand g452 ( new_n603_, new_n587_, N219 );
nor g453 ( new_n604_, new_n603_, new_n585_ );
not g454 ( new_n605_, new_n599_ );
nor g455 ( new_n606_, new_n604_, new_n605_ );
nand g456 ( new_n607_, new_n606_, new_n602_ );
nand g457 ( N878, new_n601_, new_n607_ );
not g458 ( new_n609_, keyIn_0_62 );
not g459 ( new_n610_, keyIn_0_56 );
not g460 ( new_n611_, keyIn_0_53 );
nor g461 ( new_n612_, new_n517_, new_n537_ );
nand g462 ( new_n613_, new_n506_, new_n612_ );
nor g463 ( new_n614_, new_n613_, new_n611_ );
not g464 ( new_n615_, new_n614_ );
nand g465 ( new_n616_, new_n613_, new_n611_ );
not g466 ( new_n617_, new_n549_ );
nor g467 ( new_n618_, new_n517_, new_n543_ );
nor g468 ( new_n619_, new_n618_, new_n617_ );
and g469 ( new_n620_, new_n616_, new_n619_ );
nand g470 ( new_n621_, new_n620_, new_n615_ );
nand g471 ( new_n622_, new_n621_, new_n610_ );
nand g472 ( new_n623_, new_n616_, new_n619_ );
nor g473 ( new_n624_, new_n623_, new_n614_ );
nand g474 ( new_n625_, new_n624_, keyIn_0_56 );
nand g475 ( new_n626_, new_n622_, new_n625_ );
nor g476 ( new_n627_, new_n548_, new_n524_ );
not g477 ( new_n628_, new_n627_ );
nor g478 ( new_n629_, new_n626_, new_n628_ );
not g479 ( new_n630_, new_n629_ );
nand g480 ( new_n631_, new_n626_, new_n628_ );
and g481 ( new_n632_, new_n631_, N219 );
nand g482 ( new_n633_, new_n632_, new_n630_ );
nor g483 ( new_n634_, new_n628_, new_n319_ );
nor g484 ( new_n635_, new_n547_, new_n321_ );
nand g485 ( new_n636_, new_n523_, N246 );
nand g486 ( new_n637_, N91, N210 );
nand g487 ( new_n638_, new_n331_, N165 );
and g488 ( new_n639_, new_n638_, new_n637_ );
nand g489 ( new_n640_, new_n636_, new_n639_ );
nor g490 ( new_n641_, new_n635_, new_n640_ );
not g491 ( new_n642_, new_n641_ );
nor g492 ( new_n643_, new_n634_, new_n642_ );
nand g493 ( new_n644_, new_n633_, new_n643_ );
nand g494 ( new_n645_, new_n644_, new_n609_ );
nand g495 ( new_n646_, new_n631_, N219 );
nor g496 ( new_n647_, new_n646_, new_n629_ );
not g497 ( new_n648_, new_n643_ );
nor g498 ( new_n649_, new_n647_, new_n648_ );
nand g499 ( new_n650_, new_n649_, keyIn_0_62 );
nand g500 ( N879, new_n645_, new_n650_ );
nand g501 ( new_n652_, new_n567_, new_n543_ );
nor g502 ( new_n653_, new_n617_, new_n517_ );
nand g503 ( new_n654_, new_n652_, new_n653_ );
nor g504 ( new_n655_, new_n652_, new_n653_ );
nor g505 ( new_n656_, new_n655_, new_n463_ );
nand g506 ( new_n657_, new_n656_, new_n654_ );
and g507 ( new_n658_, new_n653_, N228 );
nand g508 ( new_n659_, new_n617_, N237 );
and g509 ( new_n660_, new_n516_, N246 );
nand g510 ( new_n661_, N96, N210 );
nand g511 ( new_n662_, new_n331_, N171 );
nand g512 ( new_n663_, new_n662_, new_n661_ );
nor g513 ( new_n664_, new_n660_, new_n663_ );
nand g514 ( new_n665_, new_n664_, new_n659_ );
nor g515 ( new_n666_, new_n658_, new_n665_ );
nand g516 ( new_n667_, new_n657_, new_n666_ );
xor g517 ( N880, new_n667_, keyIn_0_63 );
endmodule