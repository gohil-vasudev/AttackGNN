module add_mul_comp_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212;

  NAND2_X1 U111 ( .A1(n103), .A2(n104), .ZN(Result_7_) );
  NAND2_X1 U112 ( .A1(n105), .A2(n106), .ZN(n104) );
  NAND2_X1 U113 ( .A1(n107), .A2(n108), .ZN(n103) );
  NAND2_X1 U114 ( .A1(n109), .A2(n110), .ZN(n108) );
  NAND2_X1 U115 ( .A1(b_3_), .A2(n111), .ZN(n110) );
  NAND2_X1 U116 ( .A1(n112), .A2(n113), .ZN(Result_6_) );
  NAND2_X1 U117 ( .A1(n114), .A2(n106), .ZN(n113) );
  XNOR2_X1 U118 ( .A(n115), .B(n116), .ZN(n114) );
  NAND2_X1 U119 ( .A1(b_2_), .A2(a_3_), .ZN(n116) );
  NAND2_X1 U120 ( .A1(n117), .A2(n107), .ZN(n112) );
  XOR2_X1 U121 ( .A(n105), .B(n118), .Z(n117) );
  XOR2_X1 U122 ( .A(b_2_), .B(a_2_), .Z(n118) );
  NAND2_X1 U123 ( .A1(n119), .A2(n120), .ZN(Result_5_) );
  NAND2_X1 U124 ( .A1(n107), .A2(n121), .ZN(n120) );
  NAND2_X1 U125 ( .A1(n122), .A2(n123), .ZN(n121) );
  OR2_X1 U126 ( .A1(n124), .A2(n125), .ZN(n123) );
  NOR2_X1 U127 ( .A1(n126), .A2(n127), .ZN(n122) );
  NOR2_X1 U128 ( .A1(b_1_), .A2(n128), .ZN(n127) );
  XOR2_X1 U129 ( .A(a_1_), .B(n125), .Z(n128) );
  NOR2_X1 U130 ( .A1(n129), .A2(n130), .ZN(n126) );
  NAND2_X1 U131 ( .A1(n125), .A2(n131), .ZN(n130) );
  NAND2_X1 U132 ( .A1(n132), .A2(n106), .ZN(n119) );
  XOR2_X1 U133 ( .A(n133), .B(n134), .Z(n132) );
  XOR2_X1 U134 ( .A(n135), .B(n136), .Z(n134) );
  NAND2_X1 U135 ( .A1(n137), .A2(n138), .ZN(Result_4_) );
  NAND2_X1 U136 ( .A1(n139), .A2(n106), .ZN(n138) );
  XOR2_X1 U137 ( .A(n140), .B(n141), .Z(n139) );
  XOR2_X1 U138 ( .A(n142), .B(n143), .Z(n141) );
  NOR2_X1 U139 ( .A1(n144), .A2(n145), .ZN(n143) );
  NAND2_X1 U140 ( .A1(n146), .A2(n107), .ZN(n137) );
  XOR2_X1 U141 ( .A(n147), .B(n148), .Z(n146) );
  NAND2_X1 U142 ( .A1(n149), .A2(n150), .ZN(n148) );
  NAND2_X1 U143 ( .A1(n125), .A2(n124), .ZN(n150) );
  NOR2_X1 U144 ( .A1(n151), .A2(n152), .ZN(n125) );
  AND2_X1 U145 ( .A1(n105), .A2(n153), .ZN(n151) );
  NAND2_X1 U146 ( .A1(n154), .A2(n155), .ZN(n153) );
  NOR2_X1 U147 ( .A1(n145), .A2(n111), .ZN(n105) );
  NAND2_X1 U148 ( .A1(n131), .A2(n129), .ZN(n149) );
  NOR2_X1 U149 ( .A1(n107), .A2(n156), .ZN(Result_3_) );
  XNOR2_X1 U150 ( .A(n157), .B(n158), .ZN(n156) );
  NOR2_X1 U151 ( .A1(n107), .A2(n159), .ZN(Result_2_) );
  XNOR2_X1 U152 ( .A(n160), .B(n161), .ZN(n159) );
  NOR2_X1 U153 ( .A1(n107), .A2(n162), .ZN(Result_1_) );
  XNOR2_X1 U154 ( .A(n163), .B(n164), .ZN(n162) );
  NOR2_X1 U155 ( .A1(n107), .A2(n165), .ZN(Result_0_) );
  NOR2_X1 U156 ( .A1(n166), .A2(n167), .ZN(n165) );
  NAND2_X1 U157 ( .A1(n168), .A2(n169), .ZN(n167) );
  NOR2_X1 U158 ( .A1(n164), .A2(n163), .ZN(n166) );
  NAND2_X1 U159 ( .A1(n168), .A2(n170), .ZN(n163) );
  NAND2_X1 U160 ( .A1(n171), .A2(n172), .ZN(n170) );
  OR2_X1 U161 ( .A1(n172), .A2(n171), .ZN(n168) );
  NAND2_X1 U162 ( .A1(n173), .A2(n174), .ZN(n171) );
  NAND2_X1 U163 ( .A1(b_0_), .A2(n169), .ZN(n172) );
  OR2_X1 U164 ( .A1(n175), .A2(n129), .ZN(n169) );
  NAND2_X1 U165 ( .A1(n160), .A2(n161), .ZN(n164) );
  XOR2_X1 U166 ( .A(n174), .B(n173), .Z(n161) );
  XNOR2_X1 U167 ( .A(n175), .B(n176), .ZN(n173) );
  NOR2_X1 U168 ( .A1(n144), .A2(n177), .ZN(n176) );
  NAND2_X1 U169 ( .A1(b_1_), .A2(n178), .ZN(n177) );
  NAND2_X1 U170 ( .A1(a_1_), .A2(b_0_), .ZN(n175) );
  NAND2_X1 U171 ( .A1(n179), .A2(n180), .ZN(n174) );
  NAND2_X1 U172 ( .A1(b_2_), .A2(n181), .ZN(n180) );
  AND2_X1 U173 ( .A1(n158), .A2(n157), .ZN(n160) );
  NAND2_X1 U174 ( .A1(n142), .A2(n182), .ZN(n157) );
  NAND2_X1 U175 ( .A1(n183), .A2(b_3_), .ZN(n182) );
  NOR2_X1 U176 ( .A1(n140), .A2(n144), .ZN(n183) );
  XNOR2_X1 U177 ( .A(n184), .B(n185), .ZN(n140) );
  XNOR2_X1 U178 ( .A(n186), .B(n187), .ZN(n184) );
  NAND2_X1 U179 ( .A1(b_2_), .A2(a_1_), .ZN(n186) );
  AND2_X1 U180 ( .A1(n188), .A2(n189), .ZN(n142) );
  NAND2_X1 U181 ( .A1(n135), .A2(n190), .ZN(n189) );
  NAND2_X1 U182 ( .A1(n191), .A2(n192), .ZN(n190) );
  AND2_X1 U183 ( .A1(n193), .A2(n115), .ZN(n135) );
  NOR2_X1 U184 ( .A1(n145), .A2(n154), .ZN(n115) );
  NOR2_X1 U185 ( .A1(n111), .A2(n155), .ZN(n193) );
  NAND2_X1 U186 ( .A1(n136), .A2(n133), .ZN(n188) );
  INV_X1 U187 ( .A(n191), .ZN(n133) );
  XNOR2_X1 U188 ( .A(n152), .B(n194), .ZN(n191) );
  INV_X1 U189 ( .A(n192), .ZN(n136) );
  NAND2_X1 U190 ( .A1(b_3_), .A2(a_1_), .ZN(n192) );
  XNOR2_X1 U191 ( .A(n195), .B(n196), .ZN(n158) );
  NOR2_X1 U192 ( .A1(n155), .A2(n144), .ZN(n196) );
  XOR2_X1 U193 ( .A(n181), .B(n179), .Z(n195) );
  AND2_X1 U194 ( .A1(n187), .A2(n197), .ZN(n179) );
  NAND2_X1 U195 ( .A1(n198), .A2(b_2_), .ZN(n197) );
  NOR2_X1 U196 ( .A1(n185), .A2(n131), .ZN(n198) );
  XNOR2_X1 U197 ( .A(n199), .B(n200), .ZN(n185) );
  NOR2_X1 U198 ( .A1(n154), .A2(n129), .ZN(n200) );
  NAND2_X1 U199 ( .A1(n194), .A2(n152), .ZN(n187) );
  NOR2_X1 U200 ( .A1(n155), .A2(n154), .ZN(n152) );
  NOR2_X1 U201 ( .A1(n129), .A2(n111), .ZN(n194) );
  INV_X1 U202 ( .A(a_3_), .ZN(n111) );
  NAND2_X1 U203 ( .A1(n201), .A2(n202), .ZN(n181) );
  NAND2_X1 U204 ( .A1(n199), .A2(a_2_), .ZN(n202) );
  AND2_X1 U205 ( .A1(a_3_), .A2(b_0_), .ZN(n199) );
  XNOR2_X1 U206 ( .A(n124), .B(n178), .ZN(n201) );
  NAND2_X1 U207 ( .A1(a_2_), .A2(b_0_), .ZN(n178) );
  NAND2_X1 U208 ( .A1(b_1_), .A2(a_1_), .ZN(n124) );
  INV_X1 U209 ( .A(n106), .ZN(n107) );
  NAND2_X1 U210 ( .A1(n203), .A2(n204), .ZN(n106) );
  NAND2_X1 U211 ( .A1(n205), .A2(n147), .ZN(n204) );
  NAND2_X1 U212 ( .A1(b_0_), .A2(n144), .ZN(n147) );
  NAND2_X1 U213 ( .A1(n206), .A2(n207), .ZN(n205) );
  NAND2_X1 U214 ( .A1(a_1_), .A2(n129), .ZN(n207) );
  INV_X1 U215 ( .A(b_1_), .ZN(n129) );
  NAND2_X1 U216 ( .A1(n208), .A2(n209), .ZN(n206) );
  NAND2_X1 U217 ( .A1(b_1_), .A2(n131), .ZN(n209) );
  INV_X1 U218 ( .A(a_1_), .ZN(n131) );
  NOR2_X1 U219 ( .A1(n210), .A2(n211), .ZN(n208) );
  AND2_X1 U220 ( .A1(n154), .A2(n109), .ZN(n211) );
  NOR2_X1 U221 ( .A1(n212), .A2(n155), .ZN(n210) );
  INV_X1 U222 ( .A(b_2_), .ZN(n155) );
  NOR2_X1 U223 ( .A1(n109), .A2(n154), .ZN(n212) );
  INV_X1 U224 ( .A(a_2_), .ZN(n154) );
  NAND2_X1 U225 ( .A1(a_3_), .A2(n145), .ZN(n109) );
  INV_X1 U226 ( .A(b_3_), .ZN(n145) );
  OR2_X1 U227 ( .A1(n144), .A2(b_0_), .ZN(n203) );
  INV_X1 U228 ( .A(a_0_), .ZN(n144) );
endmodule

