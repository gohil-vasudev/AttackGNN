module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n701_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n855_, new_n606_, new_n589_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n882_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n851_, new_n878_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n837_, new_n789_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n651_, new_n433_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n904_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, keyIn_0_20 );
not g001 ( new_n107_, keyIn_0_4 );
not g002 ( new_n108_, N69 );
nand g003 ( new_n109_, new_n108_, N65 );
not g004 ( new_n110_, N65 );
nand g005 ( new_n111_, new_n110_, N69 );
nand g006 ( new_n112_, new_n109_, new_n111_ );
not g007 ( new_n113_, N77 );
nand g008 ( new_n114_, new_n113_, N73 );
not g009 ( new_n115_, N73 );
nand g010 ( new_n116_, new_n115_, N77 );
nand g011 ( new_n117_, new_n114_, new_n116_ );
not g012 ( new_n118_, new_n117_ );
nand g013 ( new_n119_, new_n118_, new_n112_ );
nor g014 ( new_n120_, new_n110_, N69 );
nor g015 ( new_n121_, new_n108_, N65 );
nor g016 ( new_n122_, new_n120_, new_n121_ );
nand g017 ( new_n123_, new_n122_, new_n117_ );
nand g018 ( new_n124_, new_n119_, new_n123_ );
nand g019 ( new_n125_, new_n124_, new_n107_ );
not g020 ( new_n126_, new_n124_ );
nand g021 ( new_n127_, new_n126_, keyIn_0_4 );
nand g022 ( new_n128_, new_n127_, new_n125_ );
not g023 ( new_n129_, N89 );
nor g024 ( new_n130_, new_n129_, N93 );
not g025 ( new_n131_, N93 );
nor g026 ( new_n132_, new_n131_, N89 );
nor g027 ( new_n133_, new_n130_, new_n132_ );
not g028 ( new_n134_, N81 );
nor g029 ( new_n135_, new_n134_, N85 );
not g030 ( new_n136_, N85 );
nor g031 ( new_n137_, new_n136_, N81 );
nor g032 ( new_n138_, new_n135_, new_n137_ );
not g033 ( new_n139_, new_n138_ );
nand g034 ( new_n140_, new_n139_, new_n133_ );
not g035 ( new_n141_, new_n133_ );
nand g036 ( new_n142_, new_n141_, new_n138_ );
nand g037 ( new_n143_, new_n140_, new_n142_ );
nand g038 ( new_n144_, new_n143_, keyIn_0_5 );
not g039 ( new_n145_, new_n144_ );
nor g040 ( new_n146_, new_n143_, keyIn_0_5 );
nor g041 ( new_n147_, new_n145_, new_n146_ );
nand g042 ( new_n148_, new_n147_, new_n128_ );
not g043 ( new_n149_, new_n125_ );
nor g044 ( new_n150_, new_n124_, new_n107_ );
nor g045 ( new_n151_, new_n149_, new_n150_ );
not g046 ( new_n152_, new_n146_ );
nand g047 ( new_n153_, new_n152_, new_n144_ );
nand g048 ( new_n154_, new_n153_, new_n151_ );
nand g049 ( new_n155_, new_n148_, new_n154_ );
nand g050 ( new_n156_, new_n155_, new_n106_ );
not g051 ( new_n157_, new_n155_ );
nand g052 ( new_n158_, new_n157_, keyIn_0_20 );
nand g053 ( new_n159_, new_n158_, new_n156_ );
nand g054 ( new_n160_, N129, N137 );
not g055 ( new_n161_, new_n160_ );
nand g056 ( new_n162_, new_n159_, new_n161_ );
not g057 ( new_n163_, new_n156_ );
nor g058 ( new_n164_, new_n155_, new_n106_ );
nor g059 ( new_n165_, new_n163_, new_n164_ );
nand g060 ( new_n166_, new_n165_, new_n160_ );
nand g061 ( new_n167_, new_n166_, new_n162_ );
nand g062 ( new_n168_, new_n167_, keyIn_0_24 );
not g063 ( new_n169_, keyIn_0_24 );
nor g064 ( new_n170_, new_n165_, new_n160_ );
nor g065 ( new_n171_, new_n159_, new_n161_ );
nor g066 ( new_n172_, new_n170_, new_n171_ );
nand g067 ( new_n173_, new_n172_, new_n169_ );
nand g068 ( new_n174_, new_n173_, new_n168_ );
not g069 ( new_n175_, keyIn_0_8 );
not g070 ( new_n176_, N33 );
nor g071 ( new_n177_, new_n176_, N49 );
not g072 ( new_n178_, N49 );
nor g073 ( new_n179_, new_n178_, N33 );
nor g074 ( new_n180_, new_n177_, new_n179_ );
not g075 ( new_n181_, new_n180_ );
not g076 ( new_n182_, N1 );
nor g077 ( new_n183_, new_n182_, N17 );
not g078 ( new_n184_, N17 );
nor g079 ( new_n185_, new_n184_, N1 );
nor g080 ( new_n186_, new_n183_, new_n185_ );
nor g081 ( new_n187_, new_n181_, new_n186_ );
nand g082 ( new_n188_, new_n181_, new_n186_ );
not g083 ( new_n189_, new_n188_ );
nor g084 ( new_n190_, new_n189_, new_n187_ );
not g085 ( new_n191_, new_n190_ );
nand g086 ( new_n192_, new_n191_, new_n175_ );
not g087 ( new_n193_, new_n192_ );
nor g088 ( new_n194_, new_n191_, new_n175_ );
nor g089 ( new_n195_, new_n193_, new_n194_ );
not g090 ( new_n196_, new_n195_ );
nand g091 ( new_n197_, new_n174_, new_n196_ );
not g092 ( new_n198_, new_n168_ );
nor g093 ( new_n199_, new_n167_, keyIn_0_24 );
nor g094 ( new_n200_, new_n198_, new_n199_ );
nand g095 ( new_n201_, new_n200_, new_n195_ );
nand g096 ( new_n202_, new_n201_, new_n197_ );
not g097 ( new_n203_, keyIn_0_7 );
not g098 ( new_n204_, N117 );
nand g099 ( new_n205_, new_n204_, N113 );
not g100 ( new_n206_, N113 );
nand g101 ( new_n207_, new_n206_, N117 );
nand g102 ( new_n208_, new_n205_, new_n207_ );
not g103 ( new_n209_, N125 );
nand g104 ( new_n210_, new_n209_, N121 );
not g105 ( new_n211_, N121 );
nand g106 ( new_n212_, new_n211_, N125 );
nand g107 ( new_n213_, new_n210_, new_n212_ );
not g108 ( new_n214_, new_n213_ );
nand g109 ( new_n215_, new_n214_, new_n208_ );
not g110 ( new_n216_, new_n208_ );
nand g111 ( new_n217_, new_n216_, new_n213_ );
nand g112 ( new_n218_, new_n215_, new_n217_ );
nand g113 ( new_n219_, new_n218_, new_n203_ );
not g114 ( new_n220_, new_n219_ );
nor g115 ( new_n221_, new_n218_, new_n203_ );
nor g116 ( new_n222_, new_n220_, new_n221_ );
not g117 ( new_n223_, N101 );
nand g118 ( new_n224_, new_n223_, N97 );
not g119 ( new_n225_, N97 );
nand g120 ( new_n226_, new_n225_, N101 );
nand g121 ( new_n227_, new_n224_, new_n226_ );
not g122 ( new_n228_, N105 );
nor g123 ( new_n229_, new_n228_, N109 );
not g124 ( new_n230_, N109 );
nor g125 ( new_n231_, new_n230_, N105 );
nor g126 ( new_n232_, new_n229_, new_n231_ );
nand g127 ( new_n233_, new_n232_, new_n227_ );
nor g128 ( new_n234_, new_n225_, N101 );
nor g129 ( new_n235_, new_n223_, N97 );
nor g130 ( new_n236_, new_n234_, new_n235_ );
nand g131 ( new_n237_, new_n230_, N105 );
nand g132 ( new_n238_, new_n228_, N109 );
nand g133 ( new_n239_, new_n237_, new_n238_ );
nand g134 ( new_n240_, new_n236_, new_n239_ );
nand g135 ( new_n241_, new_n233_, new_n240_ );
nand g136 ( new_n242_, new_n241_, keyIn_0_6 );
not g137 ( new_n243_, new_n242_ );
nor g138 ( new_n244_, new_n241_, keyIn_0_6 );
nor g139 ( new_n245_, new_n243_, new_n244_ );
nand g140 ( new_n246_, new_n222_, new_n245_ );
not g141 ( new_n247_, new_n218_ );
nand g142 ( new_n248_, new_n247_, keyIn_0_7 );
nand g143 ( new_n249_, new_n248_, new_n219_ );
not g144 ( new_n250_, keyIn_0_6 );
not g145 ( new_n251_, new_n241_ );
nand g146 ( new_n252_, new_n251_, new_n250_ );
nand g147 ( new_n253_, new_n252_, new_n242_ );
nand g148 ( new_n254_, new_n249_, new_n253_ );
nand g149 ( new_n255_, new_n246_, new_n254_ );
nor g150 ( new_n256_, new_n255_, keyIn_0_21 );
nand g151 ( new_n257_, new_n255_, keyIn_0_21 );
not g152 ( new_n258_, new_n257_ );
nor g153 ( new_n259_, new_n258_, new_n256_ );
nand g154 ( new_n260_, N130, N137 );
not g155 ( new_n261_, new_n260_ );
nor g156 ( new_n262_, new_n259_, new_n261_ );
not g157 ( new_n263_, keyIn_0_21 );
not g158 ( new_n264_, new_n255_ );
nand g159 ( new_n265_, new_n264_, new_n263_ );
nand g160 ( new_n266_, new_n265_, new_n257_ );
nor g161 ( new_n267_, new_n266_, new_n260_ );
nor g162 ( new_n268_, new_n262_, new_n267_ );
nor g163 ( new_n269_, new_n268_, keyIn_0_25 );
not g164 ( new_n270_, keyIn_0_25 );
nand g165 ( new_n271_, new_n266_, new_n260_ );
nand g166 ( new_n272_, new_n259_, new_n261_ );
nand g167 ( new_n273_, new_n272_, new_n271_ );
nor g168 ( new_n274_, new_n273_, new_n270_ );
nor g169 ( new_n275_, new_n269_, new_n274_ );
not g170 ( new_n276_, N37 );
nor g171 ( new_n277_, new_n276_, N53 );
not g172 ( new_n278_, N53 );
nor g173 ( new_n279_, new_n278_, N37 );
nor g174 ( new_n280_, new_n277_, new_n279_ );
not g175 ( new_n281_, new_n280_ );
not g176 ( new_n282_, N5 );
nor g177 ( new_n283_, new_n282_, N21 );
not g178 ( new_n284_, N21 );
nor g179 ( new_n285_, new_n284_, N5 );
nor g180 ( new_n286_, new_n283_, new_n285_ );
nor g181 ( new_n287_, new_n281_, new_n286_ );
nand g182 ( new_n288_, new_n281_, new_n286_ );
not g183 ( new_n289_, new_n288_ );
nor g184 ( new_n290_, new_n289_, new_n287_ );
not g185 ( new_n291_, new_n290_ );
nand g186 ( new_n292_, new_n291_, keyIn_0_9 );
not g187 ( new_n293_, new_n292_ );
nor g188 ( new_n294_, new_n291_, keyIn_0_9 );
nor g189 ( new_n295_, new_n293_, new_n294_ );
nand g190 ( new_n296_, new_n275_, new_n295_ );
nand g191 ( new_n297_, new_n273_, new_n270_ );
nand g192 ( new_n298_, new_n268_, keyIn_0_25 );
nand g193 ( new_n299_, new_n298_, new_n297_ );
not g194 ( new_n300_, new_n295_ );
nand g195 ( new_n301_, new_n299_, new_n300_ );
nand g196 ( new_n302_, new_n296_, new_n301_ );
not g197 ( new_n303_, keyIn_0_26 );
not g198 ( new_n304_, keyIn_0_22 );
nand g199 ( new_n305_, new_n151_, new_n245_ );
nand g200 ( new_n306_, new_n128_, new_n253_ );
nand g201 ( new_n307_, new_n305_, new_n306_ );
nor g202 ( new_n308_, new_n307_, new_n304_ );
nand g203 ( new_n309_, new_n307_, new_n304_ );
not g204 ( new_n310_, new_n309_ );
nor g205 ( new_n311_, new_n310_, new_n308_ );
nand g206 ( new_n312_, N131, N137 );
nor g207 ( new_n313_, new_n311_, new_n312_ );
not g208 ( new_n314_, new_n307_ );
nand g209 ( new_n315_, new_n314_, keyIn_0_22 );
nand g210 ( new_n316_, new_n315_, new_n309_ );
not g211 ( new_n317_, new_n312_ );
nor g212 ( new_n318_, new_n316_, new_n317_ );
nor g213 ( new_n319_, new_n313_, new_n318_ );
nor g214 ( new_n320_, new_n319_, new_n303_ );
nand g215 ( new_n321_, new_n316_, new_n317_ );
nand g216 ( new_n322_, new_n311_, new_n312_ );
nand g217 ( new_n323_, new_n322_, new_n321_ );
nor g218 ( new_n324_, new_n323_, keyIn_0_26 );
nor g219 ( new_n325_, new_n320_, new_n324_ );
not g220 ( new_n326_, keyIn_0_10 );
not g221 ( new_n327_, N41 );
nor g222 ( new_n328_, new_n327_, N57 );
not g223 ( new_n329_, N57 );
nor g224 ( new_n330_, new_n329_, N41 );
nor g225 ( new_n331_, new_n328_, new_n330_ );
not g226 ( new_n332_, new_n331_ );
not g227 ( new_n333_, N9 );
nor g228 ( new_n334_, new_n333_, N25 );
not g229 ( new_n335_, N25 );
nor g230 ( new_n336_, new_n335_, N9 );
nor g231 ( new_n337_, new_n334_, new_n336_ );
nor g232 ( new_n338_, new_n332_, new_n337_ );
nand g233 ( new_n339_, new_n332_, new_n337_ );
not g234 ( new_n340_, new_n339_ );
nor g235 ( new_n341_, new_n340_, new_n338_ );
not g236 ( new_n342_, new_n341_ );
nand g237 ( new_n343_, new_n342_, new_n326_ );
not g238 ( new_n344_, new_n343_ );
nor g239 ( new_n345_, new_n342_, new_n326_ );
nor g240 ( new_n346_, new_n344_, new_n345_ );
not g241 ( new_n347_, new_n346_ );
nand g242 ( new_n348_, new_n325_, new_n347_ );
nand g243 ( new_n349_, new_n323_, keyIn_0_26 );
nand g244 ( new_n350_, new_n319_, new_n303_ );
nand g245 ( new_n351_, new_n350_, new_n349_ );
nand g246 ( new_n352_, new_n351_, new_n346_ );
nand g247 ( new_n353_, new_n348_, new_n352_ );
nor g248 ( new_n354_, new_n302_, new_n353_ );
nand g249 ( new_n355_, new_n354_, new_n202_ );
not g250 ( new_n356_, keyIn_0_27 );
nand g251 ( new_n357_, new_n147_, new_n249_ );
nand g252 ( new_n358_, new_n153_, new_n222_ );
nand g253 ( new_n359_, new_n357_, new_n358_ );
nand g254 ( new_n360_, new_n359_, keyIn_0_23 );
not g255 ( new_n361_, keyIn_0_23 );
not g256 ( new_n362_, new_n359_ );
nand g257 ( new_n363_, new_n362_, new_n361_ );
nand g258 ( new_n364_, new_n363_, new_n360_ );
nand g259 ( new_n365_, N132, N137 );
nand g260 ( new_n366_, new_n364_, new_n365_ );
not g261 ( new_n367_, new_n360_ );
nor g262 ( new_n368_, new_n359_, keyIn_0_23 );
nor g263 ( new_n369_, new_n367_, new_n368_ );
not g264 ( new_n370_, new_n365_ );
nand g265 ( new_n371_, new_n369_, new_n370_ );
nand g266 ( new_n372_, new_n371_, new_n366_ );
nand g267 ( new_n373_, new_n372_, new_n356_ );
not g268 ( new_n374_, new_n373_ );
nor g269 ( new_n375_, new_n372_, new_n356_ );
nor g270 ( new_n376_, new_n374_, new_n375_ );
not g271 ( new_n377_, N45 );
nor g272 ( new_n378_, new_n377_, N61 );
not g273 ( new_n379_, N61 );
nor g274 ( new_n380_, new_n379_, N45 );
nor g275 ( new_n381_, new_n378_, new_n380_ );
not g276 ( new_n382_, new_n381_ );
not g277 ( new_n383_, N13 );
nor g278 ( new_n384_, new_n383_, N29 );
not g279 ( new_n385_, N29 );
nor g280 ( new_n386_, new_n385_, N13 );
nor g281 ( new_n387_, new_n384_, new_n386_ );
nor g282 ( new_n388_, new_n382_, new_n387_ );
nand g283 ( new_n389_, new_n382_, new_n387_ );
not g284 ( new_n390_, new_n389_ );
nor g285 ( new_n391_, new_n390_, new_n388_ );
not g286 ( new_n392_, new_n391_ );
nand g287 ( new_n393_, new_n392_, keyIn_0_11 );
not g288 ( new_n394_, new_n393_ );
nor g289 ( new_n395_, new_n392_, keyIn_0_11 );
nor g290 ( new_n396_, new_n394_, new_n395_ );
not g291 ( new_n397_, new_n396_ );
nand g292 ( new_n398_, new_n376_, new_n397_ );
nor g293 ( new_n399_, new_n369_, new_n370_ );
nor g294 ( new_n400_, new_n364_, new_n365_ );
nor g295 ( new_n401_, new_n399_, new_n400_ );
nand g296 ( new_n402_, new_n401_, keyIn_0_27 );
nand g297 ( new_n403_, new_n402_, new_n373_ );
nand g298 ( new_n404_, new_n403_, new_n396_ );
nand g299 ( new_n405_, new_n398_, new_n404_ );
nor g300 ( new_n406_, new_n355_, new_n405_ );
not g301 ( new_n407_, keyIn_0_0 );
nor g302 ( new_n408_, new_n333_, N13 );
nor g303 ( new_n409_, new_n383_, N9 );
nor g304 ( new_n410_, new_n408_, new_n409_ );
nor g305 ( new_n411_, new_n182_, N5 );
nor g306 ( new_n412_, new_n282_, N1 );
nor g307 ( new_n413_, new_n411_, new_n412_ );
not g308 ( new_n414_, new_n413_ );
nand g309 ( new_n415_, new_n414_, new_n410_ );
not g310 ( new_n416_, new_n410_ );
nand g311 ( new_n417_, new_n416_, new_n413_ );
nand g312 ( new_n418_, new_n415_, new_n417_ );
nand g313 ( new_n419_, new_n418_, new_n407_ );
not g314 ( new_n420_, new_n419_ );
nor g315 ( new_n421_, new_n418_, new_n407_ );
nor g316 ( new_n422_, new_n420_, new_n421_ );
not g317 ( new_n423_, keyIn_0_2 );
nor g318 ( new_n424_, new_n327_, N45 );
nor g319 ( new_n425_, new_n377_, N41 );
nor g320 ( new_n426_, new_n424_, new_n425_ );
nor g321 ( new_n427_, new_n176_, N37 );
nor g322 ( new_n428_, new_n276_, N33 );
nor g323 ( new_n429_, new_n427_, new_n428_ );
not g324 ( new_n430_, new_n429_ );
nand g325 ( new_n431_, new_n430_, new_n426_ );
not g326 ( new_n432_, new_n426_ );
nand g327 ( new_n433_, new_n432_, new_n429_ );
nand g328 ( new_n434_, new_n431_, new_n433_ );
nor g329 ( new_n435_, new_n434_, new_n423_ );
not g330 ( new_n436_, new_n435_ );
nand g331 ( new_n437_, new_n434_, new_n423_ );
nand g332 ( new_n438_, new_n436_, new_n437_ );
nand g333 ( new_n439_, new_n422_, new_n438_ );
not g334 ( new_n440_, new_n421_ );
nand g335 ( new_n441_, new_n440_, new_n419_ );
not g336 ( new_n442_, new_n437_ );
nor g337 ( new_n443_, new_n442_, new_n435_ );
nand g338 ( new_n444_, new_n443_, new_n441_ );
nand g339 ( new_n445_, new_n439_, new_n444_ );
nand g340 ( new_n446_, new_n445_, keyIn_0_18 );
not g341 ( new_n447_, keyIn_0_18 );
not g342 ( new_n448_, new_n445_ );
nand g343 ( new_n449_, new_n448_, new_n447_ );
nand g344 ( new_n450_, new_n449_, new_n446_ );
nand g345 ( new_n451_, N135, N137 );
not g346 ( new_n452_, new_n451_ );
nand g347 ( new_n453_, new_n450_, new_n452_ );
not g348 ( new_n454_, new_n446_ );
nor g349 ( new_n455_, new_n445_, keyIn_0_18 );
nor g350 ( new_n456_, new_n454_, new_n455_ );
nand g351 ( new_n457_, new_n456_, new_n451_ );
nand g352 ( new_n458_, new_n457_, new_n453_ );
nand g353 ( new_n459_, new_n458_, keyIn_0_30 );
not g354 ( new_n460_, keyIn_0_30 );
nor g355 ( new_n461_, new_n456_, new_n451_ );
nor g356 ( new_n462_, new_n450_, new_n452_ );
nor g357 ( new_n463_, new_n461_, new_n462_ );
nand g358 ( new_n464_, new_n463_, new_n460_ );
nand g359 ( new_n465_, new_n464_, new_n459_ );
not g360 ( new_n466_, keyIn_0_14 );
nor g361 ( new_n467_, new_n228_, N121 );
nor g362 ( new_n468_, new_n211_, N105 );
nor g363 ( new_n469_, new_n467_, new_n468_ );
not g364 ( new_n470_, new_n469_ );
nor g365 ( new_n471_, new_n115_, N89 );
nor g366 ( new_n472_, new_n129_, N73 );
nor g367 ( new_n473_, new_n471_, new_n472_ );
nor g368 ( new_n474_, new_n470_, new_n473_ );
nand g369 ( new_n475_, new_n470_, new_n473_ );
not g370 ( new_n476_, new_n475_ );
nor g371 ( new_n477_, new_n476_, new_n474_ );
not g372 ( new_n478_, new_n477_ );
nand g373 ( new_n479_, new_n478_, new_n466_ );
not g374 ( new_n480_, new_n479_ );
nor g375 ( new_n481_, new_n478_, new_n466_ );
nor g376 ( new_n482_, new_n480_, new_n481_ );
not g377 ( new_n483_, new_n482_ );
nand g378 ( new_n484_, new_n465_, new_n483_ );
nor g379 ( new_n485_, new_n463_, new_n460_ );
nor g380 ( new_n486_, new_n458_, keyIn_0_30 );
nor g381 ( new_n487_, new_n485_, new_n486_ );
nand g382 ( new_n488_, new_n487_, new_n482_ );
nand g383 ( new_n489_, new_n488_, new_n484_ );
nor g384 ( new_n490_, new_n329_, N61 );
nor g385 ( new_n491_, new_n379_, N57 );
nor g386 ( new_n492_, new_n490_, new_n491_ );
nor g387 ( new_n493_, new_n178_, N53 );
nor g388 ( new_n494_, new_n278_, N49 );
nor g389 ( new_n495_, new_n493_, new_n494_ );
not g390 ( new_n496_, new_n495_ );
nand g391 ( new_n497_, new_n496_, new_n492_ );
not g392 ( new_n498_, new_n490_ );
not g393 ( new_n499_, new_n491_ );
nand g394 ( new_n500_, new_n498_, new_n499_ );
nand g395 ( new_n501_, new_n500_, new_n495_ );
nand g396 ( new_n502_, new_n497_, new_n501_ );
nand g397 ( new_n503_, new_n502_, keyIn_0_3 );
not g398 ( new_n504_, new_n503_ );
nor g399 ( new_n505_, new_n502_, keyIn_0_3 );
nor g400 ( new_n506_, new_n504_, new_n505_ );
not g401 ( new_n507_, keyIn_0_1 );
nor g402 ( new_n508_, new_n335_, N29 );
nor g403 ( new_n509_, new_n385_, N25 );
nor g404 ( new_n510_, new_n508_, new_n509_ );
nor g405 ( new_n511_, new_n184_, N21 );
nor g406 ( new_n512_, new_n284_, N17 );
nor g407 ( new_n513_, new_n511_, new_n512_ );
not g408 ( new_n514_, new_n513_ );
nand g409 ( new_n515_, new_n514_, new_n510_ );
not g410 ( new_n516_, new_n508_ );
not g411 ( new_n517_, new_n509_ );
nand g412 ( new_n518_, new_n516_, new_n517_ );
nand g413 ( new_n519_, new_n518_, new_n513_ );
nand g414 ( new_n520_, new_n515_, new_n519_ );
nor g415 ( new_n521_, new_n520_, new_n507_ );
not g416 ( new_n522_, new_n521_ );
nand g417 ( new_n523_, new_n520_, new_n507_ );
nand g418 ( new_n524_, new_n522_, new_n523_ );
nand g419 ( new_n525_, new_n506_, new_n524_ );
not g420 ( new_n526_, new_n505_ );
nand g421 ( new_n527_, new_n526_, new_n503_ );
not g422 ( new_n528_, new_n523_ );
nor g423 ( new_n529_, new_n528_, new_n521_ );
nand g424 ( new_n530_, new_n529_, new_n527_ );
nand g425 ( new_n531_, new_n525_, new_n530_ );
nand g426 ( new_n532_, new_n531_, keyIn_0_19 );
not g427 ( new_n533_, keyIn_0_19 );
not g428 ( new_n534_, new_n531_ );
nand g429 ( new_n535_, new_n534_, new_n533_ );
nand g430 ( new_n536_, new_n535_, new_n532_ );
nand g431 ( new_n537_, N136, N137 );
nand g432 ( new_n538_, new_n536_, new_n537_ );
not g433 ( new_n539_, new_n532_ );
nor g434 ( new_n540_, new_n531_, keyIn_0_19 );
nor g435 ( new_n541_, new_n539_, new_n540_ );
not g436 ( new_n542_, new_n537_ );
nand g437 ( new_n543_, new_n541_, new_n542_ );
nand g438 ( new_n544_, new_n543_, new_n538_ );
nand g439 ( new_n545_, new_n544_, keyIn_0_31 );
not g440 ( new_n546_, keyIn_0_31 );
nor g441 ( new_n547_, new_n541_, new_n542_ );
nor g442 ( new_n548_, new_n536_, new_n537_ );
nor g443 ( new_n549_, new_n547_, new_n548_ );
nand g444 ( new_n550_, new_n549_, new_n546_ );
nand g445 ( new_n551_, new_n550_, new_n545_ );
not g446 ( new_n552_, keyIn_0_15 );
nor g447 ( new_n553_, new_n230_, N125 );
nor g448 ( new_n554_, new_n209_, N109 );
nor g449 ( new_n555_, new_n553_, new_n554_ );
not g450 ( new_n556_, new_n555_ );
nor g451 ( new_n557_, new_n113_, N93 );
nor g452 ( new_n558_, new_n131_, N77 );
nor g453 ( new_n559_, new_n557_, new_n558_ );
nor g454 ( new_n560_, new_n556_, new_n559_ );
nand g455 ( new_n561_, new_n556_, new_n559_ );
not g456 ( new_n562_, new_n561_ );
nor g457 ( new_n563_, new_n562_, new_n560_ );
not g458 ( new_n564_, new_n563_ );
nand g459 ( new_n565_, new_n564_, new_n552_ );
not g460 ( new_n566_, new_n565_ );
nor g461 ( new_n567_, new_n564_, new_n552_ );
nor g462 ( new_n568_, new_n566_, new_n567_ );
nor g463 ( new_n569_, new_n551_, new_n568_ );
nor g464 ( new_n570_, new_n549_, new_n546_ );
nor g465 ( new_n571_, new_n544_, keyIn_0_31 );
nor g466 ( new_n572_, new_n570_, new_n571_ );
not g467 ( new_n573_, new_n568_ );
nor g468 ( new_n574_, new_n572_, new_n573_ );
nor g469 ( new_n575_, new_n574_, new_n569_ );
nand g470 ( new_n576_, new_n575_, new_n489_ );
nand g471 ( new_n577_, new_n441_, new_n524_ );
nand g472 ( new_n578_, new_n422_, new_n529_ );
nand g473 ( new_n579_, new_n578_, new_n577_ );
not g474 ( new_n580_, new_n579_ );
nand g475 ( new_n581_, new_n580_, keyIn_0_16 );
not g476 ( new_n582_, keyIn_0_16 );
nand g477 ( new_n583_, new_n579_, new_n582_ );
nand g478 ( new_n584_, new_n581_, new_n583_ );
nand g479 ( new_n585_, N133, N137 );
not g480 ( new_n586_, new_n585_ );
nand g481 ( new_n587_, new_n584_, new_n586_ );
nor g482 ( new_n588_, new_n579_, new_n582_ );
not g483 ( new_n589_, new_n583_ );
nor g484 ( new_n590_, new_n589_, new_n588_ );
nand g485 ( new_n591_, new_n590_, new_n585_ );
nand g486 ( new_n592_, new_n591_, new_n587_ );
nand g487 ( new_n593_, new_n592_, keyIn_0_28 );
not g488 ( new_n594_, keyIn_0_28 );
nor g489 ( new_n595_, new_n590_, new_n585_ );
nor g490 ( new_n596_, new_n584_, new_n586_ );
nor g491 ( new_n597_, new_n595_, new_n596_ );
nand g492 ( new_n598_, new_n597_, new_n594_ );
nand g493 ( new_n599_, new_n598_, new_n593_ );
nor g494 ( new_n600_, new_n225_, N113 );
nor g495 ( new_n601_, new_n206_, N97 );
nor g496 ( new_n602_, new_n600_, new_n601_ );
not g497 ( new_n603_, new_n602_ );
nor g498 ( new_n604_, new_n110_, N81 );
nor g499 ( new_n605_, new_n134_, N65 );
nor g500 ( new_n606_, new_n604_, new_n605_ );
nor g501 ( new_n607_, new_n603_, new_n606_ );
nand g502 ( new_n608_, new_n603_, new_n606_ );
not g503 ( new_n609_, new_n608_ );
nor g504 ( new_n610_, new_n609_, new_n607_ );
not g505 ( new_n611_, new_n610_ );
nand g506 ( new_n612_, new_n611_, keyIn_0_12 );
not g507 ( new_n613_, new_n612_ );
nor g508 ( new_n614_, new_n611_, keyIn_0_12 );
nor g509 ( new_n615_, new_n613_, new_n614_ );
nand g510 ( new_n616_, new_n599_, new_n615_ );
nor g511 ( new_n617_, new_n597_, new_n594_ );
nor g512 ( new_n618_, new_n592_, keyIn_0_28 );
nor g513 ( new_n619_, new_n617_, new_n618_ );
not g514 ( new_n620_, new_n615_ );
nand g515 ( new_n621_, new_n619_, new_n620_ );
nand g516 ( new_n622_, new_n621_, new_n616_ );
not g517 ( new_n623_, keyIn_0_17 );
nand g518 ( new_n624_, new_n438_, new_n527_ );
nand g519 ( new_n625_, new_n443_, new_n506_ );
nand g520 ( new_n626_, new_n625_, new_n624_ );
not g521 ( new_n627_, new_n626_ );
nand g522 ( new_n628_, new_n627_, new_n623_ );
nand g523 ( new_n629_, new_n626_, keyIn_0_17 );
nand g524 ( new_n630_, new_n628_, new_n629_ );
nand g525 ( new_n631_, N134, N137 );
nand g526 ( new_n632_, new_n630_, new_n631_ );
nor g527 ( new_n633_, new_n626_, keyIn_0_17 );
not g528 ( new_n634_, new_n629_ );
nor g529 ( new_n635_, new_n634_, new_n633_ );
not g530 ( new_n636_, new_n631_ );
nand g531 ( new_n637_, new_n635_, new_n636_ );
nand g532 ( new_n638_, new_n637_, new_n632_ );
nand g533 ( new_n639_, new_n638_, keyIn_0_29 );
not g534 ( new_n640_, keyIn_0_29 );
nor g535 ( new_n641_, new_n635_, new_n636_ );
nor g536 ( new_n642_, new_n630_, new_n631_ );
nor g537 ( new_n643_, new_n641_, new_n642_ );
nand g538 ( new_n644_, new_n643_, new_n640_ );
nand g539 ( new_n645_, new_n644_, new_n639_ );
nor g540 ( new_n646_, new_n223_, N117 );
nor g541 ( new_n647_, new_n204_, N101 );
nor g542 ( new_n648_, new_n646_, new_n647_ );
not g543 ( new_n649_, new_n648_ );
nor g544 ( new_n650_, new_n108_, N85 );
nor g545 ( new_n651_, new_n136_, N69 );
nor g546 ( new_n652_, new_n650_, new_n651_ );
nor g547 ( new_n653_, new_n649_, new_n652_ );
nand g548 ( new_n654_, new_n649_, new_n652_ );
not g549 ( new_n655_, new_n654_ );
nor g550 ( new_n656_, new_n655_, new_n653_ );
not g551 ( new_n657_, new_n656_ );
nand g552 ( new_n658_, new_n657_, keyIn_0_13 );
not g553 ( new_n659_, new_n658_ );
nor g554 ( new_n660_, new_n657_, keyIn_0_13 );
nor g555 ( new_n661_, new_n659_, new_n660_ );
not g556 ( new_n662_, new_n661_ );
nor g557 ( new_n663_, new_n645_, new_n662_ );
nor g558 ( new_n664_, new_n643_, new_n640_ );
nor g559 ( new_n665_, new_n638_, keyIn_0_29 );
nor g560 ( new_n666_, new_n664_, new_n665_ );
nor g561 ( new_n667_, new_n666_, new_n661_ );
nor g562 ( new_n668_, new_n667_, new_n663_ );
nand g563 ( new_n669_, new_n668_, new_n622_ );
nor g564 ( new_n670_, new_n576_, new_n669_ );
nand g565 ( new_n671_, new_n406_, new_n670_ );
nand g566 ( new_n672_, new_n671_, N1 );
not g567 ( new_n673_, new_n197_ );
nor g568 ( new_n674_, new_n174_, new_n196_ );
nor g569 ( new_n675_, new_n673_, new_n674_ );
nor g570 ( new_n676_, new_n299_, new_n300_ );
nor g571 ( new_n677_, new_n275_, new_n295_ );
nor g572 ( new_n678_, new_n677_, new_n676_ );
nor g573 ( new_n679_, new_n351_, new_n346_ );
nor g574 ( new_n680_, new_n325_, new_n347_ );
nor g575 ( new_n681_, new_n680_, new_n679_ );
nand g576 ( new_n682_, new_n678_, new_n681_ );
nor g577 ( new_n683_, new_n682_, new_n675_ );
nor g578 ( new_n684_, new_n403_, new_n396_ );
not g579 ( new_n685_, new_n404_ );
nor g580 ( new_n686_, new_n685_, new_n684_ );
nand g581 ( new_n687_, new_n683_, new_n686_ );
nor g582 ( new_n688_, new_n487_, new_n482_ );
nor g583 ( new_n689_, new_n465_, new_n483_ );
nor g584 ( new_n690_, new_n688_, new_n689_ );
nand g585 ( new_n691_, new_n572_, new_n573_ );
nand g586 ( new_n692_, new_n551_, new_n568_ );
nand g587 ( new_n693_, new_n691_, new_n692_ );
nor g588 ( new_n694_, new_n690_, new_n693_ );
nor g589 ( new_n695_, new_n619_, new_n620_ );
nor g590 ( new_n696_, new_n599_, new_n615_ );
nor g591 ( new_n697_, new_n695_, new_n696_ );
nand g592 ( new_n698_, new_n666_, new_n661_ );
nand g593 ( new_n699_, new_n645_, new_n662_ );
nand g594 ( new_n700_, new_n698_, new_n699_ );
nor g595 ( new_n701_, new_n697_, new_n700_ );
nand g596 ( new_n702_, new_n694_, new_n701_ );
nor g597 ( new_n703_, new_n687_, new_n702_ );
nand g598 ( new_n704_, new_n703_, new_n182_ );
nand g599 ( N724, new_n704_, new_n672_ );
nand g600 ( new_n706_, new_n675_, new_n302_ );
nand g601 ( new_n707_, new_n686_, new_n681_ );
nor g602 ( new_n708_, new_n707_, new_n706_ );
nand g603 ( new_n709_, new_n708_, new_n670_ );
nand g604 ( new_n710_, new_n709_, N5 );
nor g605 ( new_n711_, new_n202_, new_n678_ );
nor g606 ( new_n712_, new_n405_, new_n353_ );
nand g607 ( new_n713_, new_n711_, new_n712_ );
nor g608 ( new_n714_, new_n702_, new_n713_ );
nand g609 ( new_n715_, new_n714_, new_n282_ );
nand g610 ( N725, new_n715_, new_n710_ );
nand g611 ( new_n717_, new_n686_, new_n353_ );
nand g612 ( new_n718_, new_n675_, new_n678_ );
nor g613 ( new_n719_, new_n718_, new_n717_ );
nand g614 ( new_n720_, new_n719_, new_n670_ );
nand g615 ( new_n721_, new_n720_, N9 );
nor g616 ( new_n722_, new_n405_, new_n681_ );
nor g617 ( new_n723_, new_n202_, new_n302_ );
nand g618 ( new_n724_, new_n722_, new_n723_ );
nor g619 ( new_n725_, new_n702_, new_n724_ );
nand g620 ( new_n726_, new_n725_, new_n333_ );
nand g621 ( N726, new_n726_, new_n721_ );
nand g622 ( new_n728_, new_n405_, new_n681_ );
nor g623 ( new_n729_, new_n718_, new_n728_ );
nand g624 ( new_n730_, new_n670_, new_n729_ );
nand g625 ( new_n731_, new_n730_, N13 );
not g626 ( new_n732_, new_n728_ );
nand g627 ( new_n733_, new_n732_, new_n723_ );
nor g628 ( new_n734_, new_n702_, new_n733_ );
nand g629 ( new_n735_, new_n734_, new_n383_ );
nand g630 ( N727, new_n735_, new_n731_ );
nand g631 ( new_n737_, new_n690_, new_n693_ );
nor g632 ( new_n738_, new_n737_, new_n669_ );
nand g633 ( new_n739_, new_n406_, new_n738_ );
nand g634 ( new_n740_, new_n739_, N17 );
nor g635 ( new_n741_, new_n575_, new_n489_ );
nand g636 ( new_n742_, new_n701_, new_n741_ );
nor g637 ( new_n743_, new_n687_, new_n742_ );
nand g638 ( new_n744_, new_n743_, new_n184_ );
nand g639 ( N728, new_n744_, new_n740_ );
nand g640 ( new_n746_, new_n708_, new_n738_ );
nand g641 ( new_n747_, new_n746_, N21 );
nor g642 ( new_n748_, new_n742_, new_n713_ );
nand g643 ( new_n749_, new_n748_, new_n284_ );
nand g644 ( N729, new_n749_, new_n747_ );
nand g645 ( new_n751_, new_n719_, new_n738_ );
nand g646 ( new_n752_, new_n751_, N25 );
nor g647 ( new_n753_, new_n742_, new_n724_ );
nand g648 ( new_n754_, new_n753_, new_n335_ );
nand g649 ( N730, new_n754_, new_n752_ );
nand g650 ( new_n756_, new_n738_, new_n729_ );
nand g651 ( new_n757_, new_n756_, N29 );
nor g652 ( new_n758_, new_n742_, new_n733_ );
nand g653 ( new_n759_, new_n758_, new_n385_ );
nand g654 ( N731, new_n759_, new_n757_ );
nand g655 ( new_n761_, new_n697_, new_n700_ );
nor g656 ( new_n762_, new_n576_, new_n761_ );
nand g657 ( new_n763_, new_n406_, new_n762_ );
nand g658 ( new_n764_, new_n763_, N33 );
nor g659 ( new_n765_, new_n668_, new_n622_ );
nand g660 ( new_n766_, new_n694_, new_n765_ );
nor g661 ( new_n767_, new_n687_, new_n766_ );
nand g662 ( new_n768_, new_n767_, new_n176_ );
nand g663 ( N732, new_n768_, new_n764_ );
nand g664 ( new_n770_, new_n708_, new_n762_ );
nand g665 ( new_n771_, new_n770_, N37 );
nor g666 ( new_n772_, new_n766_, new_n713_ );
nand g667 ( new_n773_, new_n772_, new_n276_ );
nand g668 ( N733, new_n773_, new_n771_ );
nand g669 ( new_n775_, new_n719_, new_n762_ );
nand g670 ( new_n776_, new_n775_, N41 );
nor g671 ( new_n777_, new_n766_, new_n724_ );
nand g672 ( new_n778_, new_n777_, new_n327_ );
nand g673 ( N734, new_n778_, new_n776_ );
nand g674 ( new_n780_, new_n762_, new_n729_ );
nand g675 ( new_n781_, new_n780_, N45 );
nor g676 ( new_n782_, new_n766_, new_n733_ );
nand g677 ( new_n783_, new_n782_, new_n377_ );
nand g678 ( N735, new_n783_, new_n781_ );
nor g679 ( new_n785_, new_n737_, new_n761_ );
nand g680 ( new_n786_, new_n406_, new_n785_ );
nand g681 ( new_n787_, new_n786_, N49 );
nand g682 ( new_n788_, new_n741_, new_n765_ );
nor g683 ( new_n789_, new_n687_, new_n788_ );
nand g684 ( new_n790_, new_n789_, new_n178_ );
nand g685 ( N736, new_n790_, new_n787_ );
nand g686 ( new_n792_, new_n708_, new_n785_ );
nand g687 ( new_n793_, new_n792_, N53 );
nor g688 ( new_n794_, new_n788_, new_n713_ );
nand g689 ( new_n795_, new_n794_, new_n278_ );
nand g690 ( N737, new_n795_, new_n793_ );
nand g691 ( new_n797_, new_n719_, new_n785_ );
nand g692 ( new_n798_, new_n797_, N57 );
nor g693 ( new_n799_, new_n788_, new_n724_ );
nand g694 ( new_n800_, new_n799_, new_n329_ );
nand g695 ( N738, new_n800_, new_n798_ );
nand g696 ( new_n802_, new_n785_, new_n729_ );
nand g697 ( new_n803_, new_n802_, N61 );
nor g698 ( new_n804_, new_n788_, new_n733_ );
nand g699 ( new_n805_, new_n804_, new_n379_ );
nand g700 ( N739, new_n805_, new_n803_ );
nand g701 ( new_n807_, new_n690_, new_n575_ );
nor g702 ( new_n808_, new_n807_, new_n669_ );
nand g703 ( new_n809_, new_n202_, new_n678_ );
nor g704 ( new_n810_, new_n717_, new_n809_ );
nand g705 ( new_n811_, new_n808_, new_n810_ );
nand g706 ( new_n812_, new_n811_, N65 );
nor g707 ( new_n813_, new_n489_, new_n693_ );
nand g708 ( new_n814_, new_n701_, new_n813_ );
not g709 ( new_n815_, new_n809_ );
nand g710 ( new_n816_, new_n815_, new_n722_ );
nor g711 ( new_n817_, new_n816_, new_n814_ );
nand g712 ( new_n818_, new_n817_, new_n110_ );
nand g713 ( N740, new_n818_, new_n812_ );
nor g714 ( new_n820_, new_n807_, new_n761_ );
nand g715 ( new_n821_, new_n820_, new_n810_ );
nand g716 ( new_n822_, new_n821_, N69 );
nand g717 ( new_n823_, new_n765_, new_n813_ );
nor g718 ( new_n824_, new_n816_, new_n823_ );
nand g719 ( new_n825_, new_n824_, new_n108_ );
nand g720 ( N741, new_n825_, new_n822_ );
nand g721 ( new_n827_, new_n697_, new_n668_ );
nor g722 ( new_n828_, new_n827_, new_n576_ );
nand g723 ( new_n829_, new_n828_, new_n810_ );
nand g724 ( new_n830_, new_n829_, N73 );
nor g725 ( new_n831_, new_n622_, new_n700_ );
nand g726 ( new_n832_, new_n694_, new_n831_ );
nor g727 ( new_n833_, new_n832_, new_n816_ );
nand g728 ( new_n834_, new_n833_, new_n115_ );
nand g729 ( N742, new_n834_, new_n830_ );
nor g730 ( new_n836_, new_n827_, new_n737_ );
nand g731 ( new_n837_, new_n836_, new_n810_ );
nand g732 ( new_n838_, new_n837_, N77 );
nand g733 ( new_n839_, new_n741_, new_n831_ );
nor g734 ( new_n840_, new_n816_, new_n839_ );
nand g735 ( new_n841_, new_n840_, new_n113_ );
nand g736 ( N743, new_n841_, new_n838_ );
nor g737 ( new_n843_, new_n355_, new_n686_ );
nand g738 ( new_n844_, new_n843_, new_n808_ );
nand g739 ( new_n845_, new_n844_, N81 );
nand g740 ( new_n846_, new_n683_, new_n405_ );
nor g741 ( new_n847_, new_n846_, new_n814_ );
nand g742 ( new_n848_, new_n847_, new_n134_ );
nand g743 ( N744, new_n848_, new_n845_ );
nand g744 ( new_n850_, new_n843_, new_n820_ );
nand g745 ( new_n851_, new_n850_, N85 );
nor g746 ( new_n852_, new_n846_, new_n823_ );
nand g747 ( new_n853_, new_n852_, new_n136_ );
nand g748 ( N745, new_n853_, new_n851_ );
nand g749 ( new_n855_, new_n843_, new_n828_ );
nand g750 ( new_n856_, new_n855_, N89 );
nor g751 ( new_n857_, new_n846_, new_n832_ );
nand g752 ( new_n858_, new_n857_, new_n129_ );
nand g753 ( N746, new_n858_, new_n856_ );
nand g754 ( new_n860_, new_n836_, new_n843_ );
nand g755 ( new_n861_, new_n860_, N93 );
nor g756 ( new_n862_, new_n846_, new_n839_ );
nand g757 ( new_n863_, new_n862_, new_n131_ );
nand g758 ( N747, new_n863_, new_n861_ );
nor g759 ( new_n865_, new_n706_, new_n717_ );
nand g760 ( new_n866_, new_n865_, new_n808_ );
nand g761 ( new_n867_, new_n866_, N97 );
nand g762 ( new_n868_, new_n711_, new_n722_ );
nor g763 ( new_n869_, new_n814_, new_n868_ );
nand g764 ( new_n870_, new_n869_, new_n225_ );
nand g765 ( N748, new_n867_, new_n870_ );
nand g766 ( new_n872_, new_n865_, new_n820_ );
nand g767 ( new_n873_, new_n872_, N101 );
nor g768 ( new_n874_, new_n823_, new_n868_ );
nand g769 ( new_n875_, new_n874_, new_n223_ );
nand g770 ( N749, new_n873_, new_n875_ );
nand g771 ( new_n877_, new_n865_, new_n828_ );
nand g772 ( new_n878_, new_n877_, N105 );
nor g773 ( new_n879_, new_n832_, new_n868_ );
nand g774 ( new_n880_, new_n879_, new_n228_ );
nand g775 ( N750, new_n880_, new_n878_ );
nand g776 ( new_n882_, new_n836_, new_n865_ );
nand g777 ( new_n883_, new_n882_, N109 );
nor g778 ( new_n884_, new_n839_, new_n868_ );
nand g779 ( new_n885_, new_n884_, new_n230_ );
nand g780 ( N751, new_n883_, new_n885_ );
nor g781 ( new_n887_, new_n706_, new_n728_ );
nand g782 ( new_n888_, new_n808_, new_n887_ );
nand g783 ( new_n889_, new_n888_, N113 );
nand g784 ( new_n890_, new_n732_, new_n711_ );
nor g785 ( new_n891_, new_n890_, new_n814_ );
nand g786 ( new_n892_, new_n891_, new_n206_ );
nand g787 ( N752, new_n892_, new_n889_ );
nand g788 ( new_n894_, new_n820_, new_n887_ );
nand g789 ( new_n895_, new_n894_, N117 );
nor g790 ( new_n896_, new_n890_, new_n823_ );
nand g791 ( new_n897_, new_n896_, new_n204_ );
nand g792 ( N753, new_n897_, new_n895_ );
nand g793 ( new_n899_, new_n828_, new_n887_ );
nand g794 ( new_n900_, new_n899_, N121 );
nor g795 ( new_n901_, new_n832_, new_n890_ );
nand g796 ( new_n902_, new_n901_, new_n211_ );
nand g797 ( N754, new_n902_, new_n900_ );
nand g798 ( new_n904_, new_n836_, new_n887_ );
nand g799 ( new_n905_, new_n904_, N125 );
nor g800 ( new_n906_, new_n890_, new_n839_ );
nand g801 ( new_n907_, new_n906_, new_n209_ );
nand g802 ( N755, new_n907_, new_n905_ );
endmodule