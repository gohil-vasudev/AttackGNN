module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n1157_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n170_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n1163_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n1167_, new_n215_, new_n626_, new_n152_, new_n959_, new_n990_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n164_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1151_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1083_, new_n167_, new_n385_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n158_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n1145_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1159_, new_n1113_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n140_, new_n1147_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n1154_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n1090_, new_n457_, new_n161_, new_n553_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n954_, new_n1032_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n1161_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n1096_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n176_, new_n1109_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n1160_, new_n809_, new_n1142_, new_n654_, new_n1166_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n1135_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n138_, new_n749_, new_n861_, new_n1095_, new_n310_, new_n144_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1065_, new_n1118_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n993_, new_n1063_, new_n824_, new_n143_, new_n520_, new_n1001_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n1155_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1069_, new_n651_, new_n433_, new_n1164_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n1165_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g0000 ( new_n138_, keyIn_0_38 );
not g0001 ( new_n139_, keyIn_0_30 );
not g0002 ( new_n140_, keyIn_0_5 );
not g0003 ( new_n141_, N69 );
nand g0004 ( new_n142_, new_n141_, N65 );
not g0005 ( new_n143_, N65 );
nand g0006 ( new_n144_, new_n143_, N69 );
nand g0007 ( new_n145_, new_n142_, new_n144_ );
nand g0008 ( new_n146_, new_n145_, new_n140_ );
not g0009 ( new_n147_, new_n146_ );
nor g0010 ( new_n148_, new_n145_, new_n140_ );
nor g0011 ( new_n149_, new_n147_, new_n148_ );
not g0012 ( new_n150_, N73 );
nor g0013 ( new_n151_, new_n150_, N77 );
not g0014 ( new_n152_, N77 );
nor g0015 ( new_n153_, new_n152_, N73 );
nor g0016 ( new_n154_, new_n151_, new_n153_ );
nor g0017 ( new_n155_, new_n149_, new_n154_ );
not g0018 ( new_n156_, new_n145_ );
nand g0019 ( new_n157_, new_n156_, keyIn_0_5 );
nand g0020 ( new_n158_, new_n157_, new_n146_ );
not g0021 ( new_n159_, new_n154_ );
nor g0022 ( new_n160_, new_n158_, new_n159_ );
nor g0023 ( new_n161_, new_n155_, new_n160_ );
nor g0024 ( new_n162_, new_n161_, keyIn_0_10 );
not g0025 ( new_n163_, keyIn_0_10 );
nand g0026 ( new_n164_, new_n158_, new_n159_ );
nand g0027 ( new_n165_, new_n149_, new_n154_ );
nand g0028 ( new_n166_, new_n165_, new_n164_ );
nor g0029 ( new_n167_, new_n166_, new_n163_ );
nor g0030 ( new_n168_, new_n162_, new_n167_ );
not g0031 ( new_n169_, keyIn_0_11 );
nand g0032 ( new_n170_, N81, N85 );
not g0033 ( new_n171_, new_n170_ );
nor g0034 ( new_n172_, N81, N85 );
nor g0035 ( new_n173_, new_n171_, new_n172_ );
nand g0036 ( new_n174_, N89, N93 );
not g0037 ( new_n175_, new_n174_ );
nor g0038 ( new_n176_, N89, N93 );
nor g0039 ( new_n177_, new_n175_, new_n176_ );
nor g0040 ( new_n178_, new_n173_, new_n177_ );
not g0041 ( new_n179_, new_n178_ );
nand g0042 ( new_n180_, new_n173_, new_n177_ );
nand g0043 ( new_n181_, new_n179_, new_n180_ );
nand g0044 ( new_n182_, new_n181_, new_n169_ );
not g0045 ( new_n183_, new_n182_ );
nor g0046 ( new_n184_, new_n181_, new_n169_ );
nor g0047 ( new_n185_, new_n183_, new_n184_ );
nor g0048 ( new_n186_, new_n168_, new_n185_ );
nand g0049 ( new_n187_, new_n166_, new_n163_ );
nand g0050 ( new_n188_, new_n161_, keyIn_0_10 );
nand g0051 ( new_n189_, new_n188_, new_n187_ );
not g0052 ( new_n190_, new_n181_ );
nand g0053 ( new_n191_, new_n190_, keyIn_0_11 );
nand g0054 ( new_n192_, new_n191_, new_n182_ );
nor g0055 ( new_n193_, new_n189_, new_n192_ );
nor g0056 ( new_n194_, new_n186_, new_n193_ );
nor g0057 ( new_n195_, new_n194_, keyIn_0_26 );
not g0058 ( new_n196_, keyIn_0_26 );
nand g0059 ( new_n197_, new_n189_, new_n192_ );
nand g0060 ( new_n198_, new_n168_, new_n185_ );
nand g0061 ( new_n199_, new_n198_, new_n197_ );
nor g0062 ( new_n200_, new_n199_, new_n196_ );
nor g0063 ( new_n201_, new_n195_, new_n200_ );
nand g0064 ( new_n202_, N129, N137 );
nor g0065 ( new_n203_, new_n201_, new_n202_ );
nand g0066 ( new_n204_, new_n199_, new_n196_ );
nand g0067 ( new_n205_, new_n194_, keyIn_0_26 );
nand g0068 ( new_n206_, new_n205_, new_n204_ );
not g0069 ( new_n207_, new_n202_ );
nor g0070 ( new_n208_, new_n206_, new_n207_ );
nor g0071 ( new_n209_, new_n203_, new_n208_ );
nor g0072 ( new_n210_, new_n209_, new_n139_ );
nand g0073 ( new_n211_, new_n206_, new_n207_ );
nand g0074 ( new_n212_, new_n201_, new_n202_ );
nand g0075 ( new_n213_, new_n212_, new_n211_ );
nor g0076 ( new_n214_, new_n213_, keyIn_0_30 );
nor g0077 ( new_n215_, new_n210_, new_n214_ );
not g0078 ( new_n216_, N1 );
nor g0079 ( new_n217_, new_n216_, N17 );
not g0080 ( new_n218_, N17 );
nor g0081 ( new_n219_, new_n218_, N1 );
nor g0082 ( new_n220_, new_n217_, new_n219_ );
not g0083 ( new_n221_, new_n220_ );
nor g0084 ( new_n222_, N33, N49 );
nand g0085 ( new_n223_, N33, N49 );
not g0086 ( new_n224_, new_n223_ );
nor g0087 ( new_n225_, new_n224_, new_n222_ );
not g0088 ( new_n226_, new_n225_ );
nor g0089 ( new_n227_, new_n221_, new_n226_ );
nor g0090 ( new_n228_, new_n220_, new_n225_ );
nor g0091 ( new_n229_, new_n227_, new_n228_ );
nor g0092 ( new_n230_, new_n229_, keyIn_0_14 );
nand g0093 ( new_n231_, new_n229_, keyIn_0_14 );
not g0094 ( new_n232_, new_n231_ );
nor g0095 ( new_n233_, new_n232_, new_n230_ );
nor g0096 ( new_n234_, new_n215_, new_n233_ );
nand g0097 ( new_n235_, new_n213_, keyIn_0_30 );
nand g0098 ( new_n236_, new_n209_, new_n139_ );
nand g0099 ( new_n237_, new_n236_, new_n235_ );
not g0100 ( new_n238_, new_n233_ );
nor g0101 ( new_n239_, new_n237_, new_n238_ );
nor g0102 ( new_n240_, new_n234_, new_n239_ );
nor g0103 ( new_n241_, new_n240_, new_n138_ );
nand g0104 ( new_n242_, new_n237_, new_n238_ );
nand g0105 ( new_n243_, new_n215_, new_n233_ );
nand g0106 ( new_n244_, new_n243_, new_n242_ );
nor g0107 ( new_n245_, new_n244_, keyIn_0_38 );
nor g0108 ( new_n246_, new_n241_, new_n245_ );
not g0109 ( new_n247_, keyIn_0_56 );
not g0110 ( new_n248_, keyIn_0_54 );
not g0111 ( new_n249_, keyIn_0_41 );
nand g0112 ( new_n250_, N113, N117 );
not g0113 ( new_n251_, new_n250_ );
nor g0114 ( new_n252_, N113, N117 );
nor g0115 ( new_n253_, new_n251_, new_n252_ );
not g0116 ( new_n254_, new_n253_ );
nand g0117 ( new_n255_, N121, N125 );
not g0118 ( new_n256_, new_n255_ );
nor g0119 ( new_n257_, N121, N125 );
nor g0120 ( new_n258_, new_n256_, new_n257_ );
nand g0121 ( new_n259_, new_n254_, new_n258_ );
not g0122 ( new_n260_, new_n258_ );
nand g0123 ( new_n261_, new_n260_, new_n253_ );
nand g0124 ( new_n262_, new_n259_, new_n261_ );
nand g0125 ( new_n263_, new_n262_, keyIn_0_13 );
nor g0126 ( new_n264_, new_n262_, keyIn_0_13 );
not g0127 ( new_n265_, new_n264_ );
nand g0128 ( new_n266_, new_n265_, new_n263_ );
nand g0129 ( new_n267_, new_n185_, new_n266_ );
not g0130 ( new_n268_, new_n263_ );
nor g0131 ( new_n269_, new_n268_, new_n264_ );
nand g0132 ( new_n270_, new_n192_, new_n269_ );
nand g0133 ( new_n271_, new_n267_, new_n270_ );
nand g0134 ( new_n272_, new_n271_, keyIn_0_29 );
nor g0135 ( new_n273_, new_n271_, keyIn_0_29 );
not g0136 ( new_n274_, new_n273_ );
nand g0137 ( new_n275_, new_n274_, new_n272_ );
nand g0138 ( new_n276_, N132, N137 );
not g0139 ( new_n277_, new_n276_ );
nand g0140 ( new_n278_, new_n275_, new_n277_ );
not g0141 ( new_n279_, new_n272_ );
nor g0142 ( new_n280_, new_n279_, new_n273_ );
nand g0143 ( new_n281_, new_n280_, new_n276_ );
nand g0144 ( new_n282_, new_n281_, new_n278_ );
nand g0145 ( new_n283_, new_n282_, keyIn_0_33 );
not g0146 ( new_n284_, new_n283_ );
nor g0147 ( new_n285_, new_n282_, keyIn_0_33 );
nor g0148 ( new_n286_, new_n284_, new_n285_ );
not g0149 ( new_n287_, keyIn_0_17 );
not g0150 ( new_n288_, N13 );
nor g0151 ( new_n289_, new_n288_, N29 );
not g0152 ( new_n290_, N29 );
nor g0153 ( new_n291_, new_n290_, N13 );
nor g0154 ( new_n292_, new_n289_, new_n291_ );
not g0155 ( new_n293_, new_n292_ );
nor g0156 ( new_n294_, N45, N61 );
nand g0157 ( new_n295_, N45, N61 );
not g0158 ( new_n296_, new_n295_ );
nor g0159 ( new_n297_, new_n296_, new_n294_ );
not g0160 ( new_n298_, new_n297_ );
nor g0161 ( new_n299_, new_n293_, new_n298_ );
nor g0162 ( new_n300_, new_n292_, new_n297_ );
nor g0163 ( new_n301_, new_n299_, new_n300_ );
nor g0164 ( new_n302_, new_n301_, new_n287_ );
nand g0165 ( new_n303_, new_n301_, new_n287_ );
not g0166 ( new_n304_, new_n303_ );
nor g0167 ( new_n305_, new_n304_, new_n302_ );
nor g0168 ( new_n306_, new_n286_, new_n305_ );
not g0169 ( new_n307_, keyIn_0_33 );
nor g0170 ( new_n308_, new_n280_, new_n276_ );
nor g0171 ( new_n309_, new_n275_, new_n277_ );
nor g0172 ( new_n310_, new_n308_, new_n309_ );
nand g0173 ( new_n311_, new_n310_, new_n307_ );
nand g0174 ( new_n312_, new_n311_, new_n283_ );
not g0175 ( new_n313_, new_n305_ );
nor g0176 ( new_n314_, new_n312_, new_n313_ );
nor g0177 ( new_n315_, new_n306_, new_n314_ );
nor g0178 ( new_n316_, new_n315_, new_n249_ );
nand g0179 ( new_n317_, new_n312_, new_n313_ );
nand g0180 ( new_n318_, new_n286_, new_n305_ );
nand g0181 ( new_n319_, new_n318_, new_n317_ );
nor g0182 ( new_n320_, new_n319_, keyIn_0_41 );
nor g0183 ( new_n321_, new_n316_, new_n320_ );
not g0184 ( new_n322_, keyIn_0_32 );
not g0185 ( new_n323_, keyIn_0_28 );
nand g0186 ( new_n324_, N97, N101 );
not g0187 ( new_n325_, new_n324_ );
nor g0188 ( new_n326_, N97, N101 );
nor g0189 ( new_n327_, new_n325_, new_n326_ );
not g0190 ( new_n328_, new_n327_ );
nand g0191 ( new_n329_, N105, N109 );
not g0192 ( new_n330_, new_n329_ );
nor g0193 ( new_n331_, N105, N109 );
nor g0194 ( new_n332_, new_n330_, new_n331_ );
not g0195 ( new_n333_, new_n332_ );
nand g0196 ( new_n334_, new_n328_, new_n333_ );
nand g0197 ( new_n335_, new_n327_, new_n332_ );
nand g0198 ( new_n336_, new_n334_, new_n335_ );
nand g0199 ( new_n337_, new_n336_, keyIn_0_12 );
nor g0200 ( new_n338_, new_n336_, keyIn_0_12 );
not g0201 ( new_n339_, new_n338_ );
nand g0202 ( new_n340_, new_n339_, new_n337_ );
nand g0203 ( new_n341_, new_n189_, new_n340_ );
not g0204 ( new_n342_, new_n337_ );
nor g0205 ( new_n343_, new_n342_, new_n338_ );
nand g0206 ( new_n344_, new_n168_, new_n343_ );
nand g0207 ( new_n345_, new_n344_, new_n341_ );
nand g0208 ( new_n346_, new_n345_, new_n323_ );
nor g0209 ( new_n347_, new_n168_, new_n343_ );
nor g0210 ( new_n348_, new_n189_, new_n340_ );
nor g0211 ( new_n349_, new_n347_, new_n348_ );
nand g0212 ( new_n350_, new_n349_, keyIn_0_28 );
nand g0213 ( new_n351_, new_n350_, new_n346_ );
nand g0214 ( new_n352_, N131, N137 );
not g0215 ( new_n353_, new_n352_ );
nand g0216 ( new_n354_, new_n351_, new_n353_ );
nor g0217 ( new_n355_, new_n349_, keyIn_0_28 );
nor g0218 ( new_n356_, new_n345_, new_n323_ );
nor g0219 ( new_n357_, new_n355_, new_n356_ );
nand g0220 ( new_n358_, new_n357_, new_n352_ );
nand g0221 ( new_n359_, new_n358_, new_n354_ );
nand g0222 ( new_n360_, new_n359_, new_n322_ );
nor g0223 ( new_n361_, new_n357_, new_n352_ );
nor g0224 ( new_n362_, new_n351_, new_n353_ );
nor g0225 ( new_n363_, new_n361_, new_n362_ );
nand g0226 ( new_n364_, new_n363_, keyIn_0_32 );
nand g0227 ( new_n365_, new_n364_, new_n360_ );
not g0228 ( new_n366_, N9 );
nor g0229 ( new_n367_, new_n366_, N25 );
not g0230 ( new_n368_, N25 );
nor g0231 ( new_n369_, new_n368_, N9 );
nor g0232 ( new_n370_, new_n367_, new_n369_ );
not g0233 ( new_n371_, new_n370_ );
nor g0234 ( new_n372_, N41, N57 );
nand g0235 ( new_n373_, N41, N57 );
not g0236 ( new_n374_, new_n373_ );
nor g0237 ( new_n375_, new_n374_, new_n372_ );
not g0238 ( new_n376_, new_n375_ );
nor g0239 ( new_n377_, new_n371_, new_n376_ );
nor g0240 ( new_n378_, new_n370_, new_n375_ );
nor g0241 ( new_n379_, new_n377_, new_n378_ );
nor g0242 ( new_n380_, new_n379_, keyIn_0_16 );
nand g0243 ( new_n381_, new_n379_, keyIn_0_16 );
not g0244 ( new_n382_, new_n381_ );
nor g0245 ( new_n383_, new_n382_, new_n380_ );
not g0246 ( new_n384_, new_n383_ );
nand g0247 ( new_n385_, new_n365_, new_n384_ );
nor g0248 ( new_n386_, new_n363_, keyIn_0_32 );
nor g0249 ( new_n387_, new_n359_, new_n322_ );
nor g0250 ( new_n388_, new_n386_, new_n387_ );
nand g0251 ( new_n389_, new_n388_, new_n383_ );
nand g0252 ( new_n390_, new_n389_, new_n385_ );
nand g0253 ( new_n391_, new_n390_, keyIn_0_40 );
not g0254 ( new_n392_, keyIn_0_40 );
nor g0255 ( new_n393_, new_n388_, new_n383_ );
nor g0256 ( new_n394_, new_n365_, new_n384_ );
nor g0257 ( new_n395_, new_n393_, new_n394_ );
nand g0258 ( new_n396_, new_n395_, new_n392_ );
nand g0259 ( new_n397_, new_n396_, new_n391_ );
nand g0260 ( new_n398_, new_n244_, keyIn_0_38 );
nand g0261 ( new_n399_, new_n240_, new_n138_ );
nand g0262 ( new_n400_, new_n399_, new_n398_ );
not g0263 ( new_n401_, keyIn_0_39 );
nand g0264 ( new_n402_, new_n343_, new_n266_ );
nand g0265 ( new_n403_, new_n269_, new_n340_ );
nand g0266 ( new_n404_, new_n402_, new_n403_ );
nand g0267 ( new_n405_, new_n404_, keyIn_0_27 );
not g0268 ( new_n406_, keyIn_0_27 );
not g0269 ( new_n407_, new_n404_ );
nand g0270 ( new_n408_, new_n407_, new_n406_ );
nand g0271 ( new_n409_, new_n408_, new_n405_ );
nand g0272 ( new_n410_, N130, N137 );
not g0273 ( new_n411_, new_n410_ );
nand g0274 ( new_n412_, new_n409_, new_n411_ );
not g0275 ( new_n413_, new_n405_ );
nor g0276 ( new_n414_, new_n404_, keyIn_0_27 );
nor g0277 ( new_n415_, new_n413_, new_n414_ );
nand g0278 ( new_n416_, new_n415_, new_n410_ );
nand g0279 ( new_n417_, new_n416_, new_n412_ );
nand g0280 ( new_n418_, new_n417_, keyIn_0_31 );
not g0281 ( new_n419_, new_n418_ );
nor g0282 ( new_n420_, new_n417_, keyIn_0_31 );
nor g0283 ( new_n421_, new_n419_, new_n420_ );
not g0284 ( new_n422_, keyIn_0_15 );
not g0285 ( new_n423_, N5 );
nor g0286 ( new_n424_, new_n423_, N21 );
not g0287 ( new_n425_, N21 );
nor g0288 ( new_n426_, new_n425_, N5 );
nor g0289 ( new_n427_, new_n424_, new_n426_ );
not g0290 ( new_n428_, new_n427_ );
nor g0291 ( new_n429_, N37, N53 );
nand g0292 ( new_n430_, N37, N53 );
not g0293 ( new_n431_, new_n430_ );
nor g0294 ( new_n432_, new_n431_, new_n429_ );
not g0295 ( new_n433_, new_n432_ );
nor g0296 ( new_n434_, new_n428_, new_n433_ );
nor g0297 ( new_n435_, new_n427_, new_n432_ );
nor g0298 ( new_n436_, new_n434_, new_n435_ );
nor g0299 ( new_n437_, new_n436_, new_n422_ );
nand g0300 ( new_n438_, new_n436_, new_n422_ );
not g0301 ( new_n439_, new_n438_ );
nor g0302 ( new_n440_, new_n439_, new_n437_ );
nand g0303 ( new_n441_, new_n421_, new_n440_ );
not g0304 ( new_n442_, keyIn_0_31 );
nor g0305 ( new_n443_, new_n415_, new_n410_ );
nor g0306 ( new_n444_, new_n409_, new_n411_ );
nor g0307 ( new_n445_, new_n443_, new_n444_ );
nand g0308 ( new_n446_, new_n445_, new_n442_ );
nand g0309 ( new_n447_, new_n446_, new_n418_ );
not g0310 ( new_n448_, new_n440_ );
nand g0311 ( new_n449_, new_n447_, new_n448_ );
nand g0312 ( new_n450_, new_n441_, new_n449_ );
nand g0313 ( new_n451_, new_n450_, new_n401_ );
nor g0314 ( new_n452_, new_n447_, new_n448_ );
not g0315 ( new_n453_, new_n449_ );
nor g0316 ( new_n454_, new_n453_, new_n452_ );
nand g0317 ( new_n455_, new_n454_, keyIn_0_39 );
nand g0318 ( new_n456_, new_n455_, new_n451_ );
nor g0319 ( new_n457_, new_n400_, new_n456_ );
nand g0320 ( new_n458_, new_n457_, new_n397_ );
nor g0321 ( new_n459_, new_n458_, new_n321_ );
nor g0322 ( new_n460_, new_n459_, keyIn_0_49 );
nand g0323 ( new_n461_, new_n459_, keyIn_0_49 );
not g0324 ( new_n462_, new_n461_ );
nor g0325 ( new_n463_, new_n462_, new_n460_ );
not g0326 ( new_n464_, new_n463_ );
nand g0327 ( new_n465_, new_n319_, keyIn_0_41 );
nand g0328 ( new_n466_, new_n315_, new_n249_ );
nand g0329 ( new_n467_, new_n466_, new_n465_ );
nor g0330 ( new_n468_, new_n395_, new_n392_ );
nor g0331 ( new_n469_, new_n390_, keyIn_0_40 );
nor g0332 ( new_n470_, new_n468_, new_n469_ );
nand g0333 ( new_n471_, new_n400_, new_n456_ );
nor g0334 ( new_n472_, new_n471_, new_n470_ );
nand g0335 ( new_n473_, new_n472_, new_n467_ );
nor g0336 ( new_n474_, new_n473_, keyIn_0_48 );
nand g0337 ( new_n475_, new_n473_, keyIn_0_48 );
not g0338 ( new_n476_, new_n475_ );
nor g0339 ( new_n477_, new_n476_, new_n474_ );
not g0340 ( new_n478_, keyIn_0_47 );
nor g0341 ( new_n479_, new_n397_, new_n321_ );
not g0342 ( new_n480_, new_n451_ );
nor g0343 ( new_n481_, new_n450_, new_n401_ );
nor g0344 ( new_n482_, new_n480_, new_n481_ );
nand g0345 ( new_n483_, new_n400_, new_n482_ );
not g0346 ( new_n484_, new_n483_ );
nand g0347 ( new_n485_, new_n484_, new_n479_ );
nand g0348 ( new_n486_, new_n485_, new_n478_ );
nand g0349 ( new_n487_, new_n470_, new_n467_ );
nor g0350 ( new_n488_, new_n487_, new_n483_ );
nand g0351 ( new_n489_, new_n488_, keyIn_0_47 );
nand g0352 ( new_n490_, new_n486_, new_n489_ );
nand g0353 ( new_n491_, new_n321_, new_n482_ );
nor g0354 ( new_n492_, new_n246_, new_n491_ );
nand g0355 ( new_n493_, new_n492_, new_n397_ );
nand g0356 ( new_n494_, new_n493_, keyIn_0_46 );
not g0357 ( new_n495_, keyIn_0_46 );
nor g0358 ( new_n496_, new_n467_, new_n456_ );
nand g0359 ( new_n497_, new_n400_, new_n496_ );
nor g0360 ( new_n498_, new_n497_, new_n470_ );
nand g0361 ( new_n499_, new_n498_, new_n495_ );
nand g0362 ( new_n500_, new_n494_, new_n499_ );
nand g0363 ( new_n501_, new_n490_, new_n500_ );
nor g0364 ( new_n502_, new_n477_, new_n501_ );
nand g0365 ( new_n503_, new_n502_, new_n464_ );
nand g0366 ( new_n504_, new_n503_, new_n248_ );
not g0367 ( new_n505_, new_n474_ );
nand g0368 ( new_n506_, new_n505_, new_n475_ );
not g0369 ( new_n507_, new_n501_ );
nand g0370 ( new_n508_, new_n507_, new_n506_ );
nor g0371 ( new_n509_, new_n508_, new_n463_ );
nand g0372 ( new_n510_, new_n509_, keyIn_0_54 );
nand g0373 ( new_n511_, new_n510_, new_n504_ );
not g0374 ( new_n512_, keyIn_0_37 );
nor g0375 ( new_n513_, N57, N61 );
nand g0376 ( new_n514_, N57, N61 );
not g0377 ( new_n515_, new_n514_ );
nor g0378 ( new_n516_, new_n515_, new_n513_ );
nand g0379 ( new_n517_, new_n516_, keyIn_0_4 );
nor g0380 ( new_n518_, new_n516_, keyIn_0_4 );
not g0381 ( new_n519_, new_n518_ );
nand g0382 ( new_n520_, new_n519_, new_n517_ );
nor g0383 ( new_n521_, N49, N53 );
nand g0384 ( new_n522_, N49, N53 );
not g0385 ( new_n523_, new_n522_ );
nor g0386 ( new_n524_, new_n523_, new_n521_ );
nand g0387 ( new_n525_, new_n524_, keyIn_0_3 );
nor g0388 ( new_n526_, new_n524_, keyIn_0_3 );
not g0389 ( new_n527_, new_n526_ );
nand g0390 ( new_n528_, new_n527_, new_n525_ );
nor g0391 ( new_n529_, new_n520_, new_n528_ );
nand g0392 ( new_n530_, new_n520_, new_n528_ );
not g0393 ( new_n531_, new_n530_ );
nor g0394 ( new_n532_, new_n531_, new_n529_ );
nor g0395 ( new_n533_, new_n532_, keyIn_0_9 );
not g0396 ( new_n534_, keyIn_0_9 );
not g0397 ( new_n535_, new_n529_ );
nand g0398 ( new_n536_, new_n535_, new_n530_ );
nor g0399 ( new_n537_, new_n536_, new_n534_ );
nor g0400 ( new_n538_, new_n537_, new_n533_ );
not g0401 ( new_n539_, keyIn_0_7 );
not g0402 ( new_n540_, keyIn_0_0 );
nor g0403 ( new_n541_, N25, N29 );
nand g0404 ( new_n542_, N25, N29 );
not g0405 ( new_n543_, new_n542_ );
nor g0406 ( new_n544_, new_n543_, new_n541_ );
nor g0407 ( new_n545_, new_n544_, new_n540_ );
not g0408 ( new_n546_, new_n545_ );
nand g0409 ( new_n547_, new_n544_, new_n540_ );
nand g0410 ( new_n548_, new_n546_, new_n547_ );
nor g0411 ( new_n549_, new_n218_, N21 );
nor g0412 ( new_n550_, new_n425_, N17 );
nor g0413 ( new_n551_, new_n549_, new_n550_ );
nand g0414 ( new_n552_, new_n548_, new_n551_ );
nor g0415 ( new_n553_, new_n548_, new_n551_ );
not g0416 ( new_n554_, new_n553_ );
nand g0417 ( new_n555_, new_n554_, new_n552_ );
nand g0418 ( new_n556_, new_n555_, new_n539_ );
not g0419 ( new_n557_, new_n552_ );
nor g0420 ( new_n558_, new_n557_, new_n553_ );
nand g0421 ( new_n559_, new_n558_, keyIn_0_7 );
nand g0422 ( new_n560_, new_n559_, new_n556_ );
nand g0423 ( new_n561_, new_n538_, new_n560_ );
nand g0424 ( new_n562_, new_n536_, new_n534_ );
nand g0425 ( new_n563_, new_n532_, keyIn_0_9 );
nand g0426 ( new_n564_, new_n562_, new_n563_ );
nor g0427 ( new_n565_, new_n558_, keyIn_0_7 );
nor g0428 ( new_n566_, new_n555_, new_n539_ );
nor g0429 ( new_n567_, new_n565_, new_n566_ );
nand g0430 ( new_n568_, new_n567_, new_n564_ );
nand g0431 ( new_n569_, new_n561_, new_n568_ );
nand g0432 ( new_n570_, new_n569_, keyIn_0_25 );
not g0433 ( new_n571_, keyIn_0_25 );
nor g0434 ( new_n572_, new_n567_, new_n564_ );
nor g0435 ( new_n573_, new_n538_, new_n560_ );
nor g0436 ( new_n574_, new_n573_, new_n572_ );
nand g0437 ( new_n575_, new_n574_, new_n571_ );
nand g0438 ( new_n576_, new_n575_, new_n570_ );
nand g0439 ( new_n577_, N136, N137 );
not g0440 ( new_n578_, new_n577_ );
nand g0441 ( new_n579_, new_n576_, new_n578_ );
not g0442 ( new_n580_, new_n570_ );
nor g0443 ( new_n581_, new_n569_, keyIn_0_25 );
nor g0444 ( new_n582_, new_n580_, new_n581_ );
nand g0445 ( new_n583_, new_n582_, new_n577_ );
nand g0446 ( new_n584_, new_n583_, new_n579_ );
nand g0447 ( new_n585_, new_n584_, new_n512_ );
not g0448 ( new_n586_, new_n579_ );
nor g0449 ( new_n587_, new_n576_, new_n578_ );
nor g0450 ( new_n588_, new_n586_, new_n587_ );
nand g0451 ( new_n589_, new_n588_, keyIn_0_37 );
nand g0452 ( new_n590_, new_n589_, new_n585_ );
not g0453 ( new_n591_, keyIn_0_21 );
nor g0454 ( new_n592_, N77, N93 );
nand g0455 ( new_n593_, N77, N93 );
not g0456 ( new_n594_, new_n593_ );
nor g0457 ( new_n595_, new_n594_, new_n592_ );
not g0458 ( new_n596_, new_n595_ );
nor g0459 ( new_n597_, N109, N125 );
nand g0460 ( new_n598_, N109, N125 );
not g0461 ( new_n599_, new_n598_ );
nor g0462 ( new_n600_, new_n599_, new_n597_ );
not g0463 ( new_n601_, new_n600_ );
nor g0464 ( new_n602_, new_n596_, new_n601_ );
nor g0465 ( new_n603_, new_n595_, new_n600_ );
nor g0466 ( new_n604_, new_n602_, new_n603_ );
not g0467 ( new_n605_, new_n604_ );
nand g0468 ( new_n606_, new_n605_, new_n591_ );
not g0469 ( new_n607_, new_n606_ );
nor g0470 ( new_n608_, new_n605_, new_n591_ );
nor g0471 ( new_n609_, new_n607_, new_n608_ );
not g0472 ( new_n610_, new_n609_ );
nand g0473 ( new_n611_, new_n590_, new_n610_ );
not g0474 ( new_n612_, new_n585_ );
nor g0475 ( new_n613_, new_n584_, new_n512_ );
nor g0476 ( new_n614_, new_n612_, new_n613_ );
nand g0477 ( new_n615_, new_n614_, new_n609_ );
nand g0478 ( new_n616_, new_n615_, new_n611_ );
nand g0479 ( new_n617_, new_n616_, keyIn_0_45 );
not g0480 ( new_n618_, keyIn_0_45 );
nor g0481 ( new_n619_, new_n614_, new_n609_ );
nor g0482 ( new_n620_, new_n590_, new_n610_ );
nor g0483 ( new_n621_, new_n619_, new_n620_ );
nand g0484 ( new_n622_, new_n621_, new_n618_ );
nand g0485 ( new_n623_, new_n622_, new_n617_ );
not g0486 ( new_n624_, keyIn_0_44 );
nor g0487 ( new_n625_, keyIn_0_1, N33 );
nand g0488 ( new_n626_, keyIn_0_1, N33 );
not g0489 ( new_n627_, new_n626_ );
nor g0490 ( new_n628_, new_n627_, new_n625_ );
nand g0491 ( new_n629_, new_n628_, N37 );
nor g0492 ( new_n630_, new_n628_, N37 );
not g0493 ( new_n631_, new_n630_ );
nand g0494 ( new_n632_, new_n631_, new_n629_ );
not g0495 ( new_n633_, keyIn_0_2 );
nor g0496 ( new_n634_, N41, N45 );
nand g0497 ( new_n635_, N41, N45 );
not g0498 ( new_n636_, new_n635_ );
nor g0499 ( new_n637_, new_n636_, new_n634_ );
nand g0500 ( new_n638_, new_n637_, new_n633_ );
nor g0501 ( new_n639_, new_n637_, new_n633_ );
not g0502 ( new_n640_, new_n639_ );
nand g0503 ( new_n641_, new_n640_, new_n638_ );
nor g0504 ( new_n642_, new_n632_, new_n641_ );
nand g0505 ( new_n643_, new_n632_, new_n641_ );
not g0506 ( new_n644_, new_n643_ );
nor g0507 ( new_n645_, new_n644_, new_n642_ );
nand g0508 ( new_n646_, new_n645_, keyIn_0_8 );
not g0509 ( new_n647_, keyIn_0_8 );
not g0510 ( new_n648_, new_n642_ );
nand g0511 ( new_n649_, new_n648_, new_n643_ );
nand g0512 ( new_n650_, new_n649_, new_n647_ );
nand g0513 ( new_n651_, new_n650_, new_n646_ );
nor g0514 ( new_n652_, N1, N5 );
nand g0515 ( new_n653_, N1, N5 );
not g0516 ( new_n654_, new_n653_ );
nor g0517 ( new_n655_, new_n654_, new_n652_ );
nand g0518 ( new_n656_, N9, N13 );
not g0519 ( new_n657_, new_n656_ );
nor g0520 ( new_n658_, N9, N13 );
nor g0521 ( new_n659_, new_n657_, new_n658_ );
nand g0522 ( new_n660_, new_n655_, new_n659_ );
not g0523 ( new_n661_, new_n655_ );
not g0524 ( new_n662_, new_n659_ );
nand g0525 ( new_n663_, new_n661_, new_n662_ );
nand g0526 ( new_n664_, new_n663_, new_n660_ );
nand g0527 ( new_n665_, new_n664_, keyIn_0_6 );
not g0528 ( new_n666_, new_n665_ );
nor g0529 ( new_n667_, new_n664_, keyIn_0_6 );
nor g0530 ( new_n668_, new_n666_, new_n667_ );
not g0531 ( new_n669_, new_n668_ );
nand g0532 ( new_n670_, new_n651_, new_n669_ );
nor g0533 ( new_n671_, new_n649_, new_n647_ );
nor g0534 ( new_n672_, new_n645_, keyIn_0_8 );
nor g0535 ( new_n673_, new_n671_, new_n672_ );
nand g0536 ( new_n674_, new_n673_, new_n668_ );
nand g0537 ( new_n675_, new_n674_, new_n670_ );
nand g0538 ( new_n676_, new_n675_, keyIn_0_24 );
not g0539 ( new_n677_, keyIn_0_24 );
not g0540 ( new_n678_, new_n670_ );
nor g0541 ( new_n679_, new_n651_, new_n669_ );
nor g0542 ( new_n680_, new_n678_, new_n679_ );
nand g0543 ( new_n681_, new_n680_, new_n677_ );
nand g0544 ( new_n682_, new_n681_, new_n676_ );
nand g0545 ( new_n683_, N135, N137 );
not g0546 ( new_n684_, new_n683_ );
nand g0547 ( new_n685_, new_n682_, new_n684_ );
not g0548 ( new_n686_, new_n676_ );
nor g0549 ( new_n687_, new_n675_, keyIn_0_24 );
nor g0550 ( new_n688_, new_n686_, new_n687_ );
nand g0551 ( new_n689_, new_n688_, new_n683_ );
nand g0552 ( new_n690_, new_n689_, new_n685_ );
nand g0553 ( new_n691_, new_n690_, keyIn_0_36 );
not g0554 ( new_n692_, keyIn_0_36 );
not g0555 ( new_n693_, new_n685_ );
nor g0556 ( new_n694_, new_n682_, new_n684_ );
nor g0557 ( new_n695_, new_n693_, new_n694_ );
nand g0558 ( new_n696_, new_n695_, new_n692_ );
nand g0559 ( new_n697_, new_n696_, new_n691_ );
not g0560 ( new_n698_, keyIn_0_20 );
nor g0561 ( new_n699_, new_n150_, N89 );
not g0562 ( new_n700_, N89 );
nor g0563 ( new_n701_, new_n700_, N73 );
nor g0564 ( new_n702_, new_n699_, new_n701_ );
not g0565 ( new_n703_, new_n702_ );
nor g0566 ( new_n704_, N105, N121 );
nand g0567 ( new_n705_, N105, N121 );
not g0568 ( new_n706_, new_n705_ );
nor g0569 ( new_n707_, new_n706_, new_n704_ );
not g0570 ( new_n708_, new_n707_ );
nor g0571 ( new_n709_, new_n703_, new_n708_ );
nor g0572 ( new_n710_, new_n702_, new_n707_ );
nor g0573 ( new_n711_, new_n709_, new_n710_ );
nor g0574 ( new_n712_, new_n711_, new_n698_ );
nand g0575 ( new_n713_, new_n711_, new_n698_ );
not g0576 ( new_n714_, new_n713_ );
nor g0577 ( new_n715_, new_n714_, new_n712_ );
not g0578 ( new_n716_, new_n715_ );
nand g0579 ( new_n717_, new_n697_, new_n716_ );
nor g0580 ( new_n718_, new_n695_, new_n692_ );
nor g0581 ( new_n719_, new_n690_, keyIn_0_36 );
nor g0582 ( new_n720_, new_n718_, new_n719_ );
nand g0583 ( new_n721_, new_n720_, new_n715_ );
nand g0584 ( new_n722_, new_n721_, new_n717_ );
nand g0585 ( new_n723_, new_n722_, new_n624_ );
nor g0586 ( new_n724_, new_n720_, new_n715_ );
nor g0587 ( new_n725_, new_n697_, new_n716_ );
nor g0588 ( new_n726_, new_n724_, new_n725_ );
nand g0589 ( new_n727_, new_n726_, keyIn_0_44 );
nand g0590 ( new_n728_, new_n727_, new_n723_ );
nand g0591 ( new_n729_, new_n623_, new_n728_ );
nand g0592 ( new_n730_, new_n538_, new_n673_ );
nand g0593 ( new_n731_, new_n564_, new_n651_ );
nand g0594 ( new_n732_, new_n730_, new_n731_ );
nand g0595 ( new_n733_, new_n732_, keyIn_0_23 );
not g0596 ( new_n734_, keyIn_0_23 );
nor g0597 ( new_n735_, new_n564_, new_n651_ );
not g0598 ( new_n736_, new_n731_ );
nor g0599 ( new_n737_, new_n736_, new_n735_ );
nand g0600 ( new_n738_, new_n737_, new_n734_ );
nand g0601 ( new_n739_, new_n738_, new_n733_ );
nand g0602 ( new_n740_, N134, N137 );
not g0603 ( new_n741_, new_n740_ );
nand g0604 ( new_n742_, new_n739_, new_n741_ );
not g0605 ( new_n743_, new_n733_ );
nor g0606 ( new_n744_, new_n732_, keyIn_0_23 );
nor g0607 ( new_n745_, new_n743_, new_n744_ );
nand g0608 ( new_n746_, new_n745_, new_n740_ );
nand g0609 ( new_n747_, new_n746_, new_n742_ );
nand g0610 ( new_n748_, new_n747_, keyIn_0_35 );
not g0611 ( new_n749_, keyIn_0_35 );
not g0612 ( new_n750_, new_n742_ );
nor g0613 ( new_n751_, new_n739_, new_n741_ );
nor g0614 ( new_n752_, new_n750_, new_n751_ );
nand g0615 ( new_n753_, new_n752_, new_n749_ );
nand g0616 ( new_n754_, new_n753_, new_n748_ );
not g0617 ( new_n755_, keyIn_0_19 );
nor g0618 ( new_n756_, N69, N85 );
nand g0619 ( new_n757_, N69, N85 );
not g0620 ( new_n758_, new_n757_ );
nor g0621 ( new_n759_, new_n758_, new_n756_ );
not g0622 ( new_n760_, new_n759_ );
nor g0623 ( new_n761_, N101, N117 );
nand g0624 ( new_n762_, N101, N117 );
not g0625 ( new_n763_, new_n762_ );
nor g0626 ( new_n764_, new_n763_, new_n761_ );
not g0627 ( new_n765_, new_n764_ );
nor g0628 ( new_n766_, new_n760_, new_n765_ );
nor g0629 ( new_n767_, new_n759_, new_n764_ );
nor g0630 ( new_n768_, new_n766_, new_n767_ );
not g0631 ( new_n769_, new_n768_ );
nand g0632 ( new_n770_, new_n769_, new_n755_ );
not g0633 ( new_n771_, new_n770_ );
nor g0634 ( new_n772_, new_n769_, new_n755_ );
nor g0635 ( new_n773_, new_n771_, new_n772_ );
not g0636 ( new_n774_, new_n773_ );
nand g0637 ( new_n775_, new_n754_, new_n774_ );
nor g0638 ( new_n776_, new_n752_, new_n749_ );
nor g0639 ( new_n777_, new_n747_, keyIn_0_35 );
nor g0640 ( new_n778_, new_n776_, new_n777_ );
nand g0641 ( new_n779_, new_n778_, new_n773_ );
nand g0642 ( new_n780_, new_n779_, new_n775_ );
nand g0643 ( new_n781_, new_n780_, keyIn_0_43 );
not g0644 ( new_n782_, keyIn_0_43 );
nor g0645 ( new_n783_, new_n778_, new_n773_ );
nor g0646 ( new_n784_, new_n754_, new_n774_ );
nor g0647 ( new_n785_, new_n783_, new_n784_ );
nand g0648 ( new_n786_, new_n785_, new_n782_ );
nand g0649 ( new_n787_, new_n786_, new_n781_ );
not g0650 ( new_n788_, keyIn_0_22 );
nand g0651 ( new_n789_, new_n560_, new_n669_ );
nand g0652 ( new_n790_, new_n567_, new_n668_ );
nand g0653 ( new_n791_, new_n790_, new_n789_ );
nand g0654 ( new_n792_, new_n791_, new_n788_ );
not g0655 ( new_n793_, new_n789_ );
nor g0656 ( new_n794_, new_n560_, new_n669_ );
nor g0657 ( new_n795_, new_n793_, new_n794_ );
nand g0658 ( new_n796_, new_n795_, keyIn_0_22 );
nand g0659 ( new_n797_, new_n796_, new_n792_ );
nand g0660 ( new_n798_, N133, N137 );
not g0661 ( new_n799_, new_n798_ );
nand g0662 ( new_n800_, new_n797_, new_n799_ );
nor g0663 ( new_n801_, new_n795_, keyIn_0_22 );
nor g0664 ( new_n802_, new_n791_, new_n788_ );
nor g0665 ( new_n803_, new_n801_, new_n802_ );
nand g0666 ( new_n804_, new_n803_, new_n798_ );
nand g0667 ( new_n805_, new_n804_, new_n800_ );
nand g0668 ( new_n806_, new_n805_, keyIn_0_34 );
not g0669 ( new_n807_, keyIn_0_34 );
nor g0670 ( new_n808_, new_n803_, new_n798_ );
nor g0671 ( new_n809_, new_n797_, new_n799_ );
nor g0672 ( new_n810_, new_n808_, new_n809_ );
nand g0673 ( new_n811_, new_n810_, new_n807_ );
nand g0674 ( new_n812_, new_n811_, new_n806_ );
nor g0675 ( new_n813_, new_n143_, N81 );
not g0676 ( new_n814_, N81 );
nor g0677 ( new_n815_, new_n814_, N65 );
nor g0678 ( new_n816_, new_n813_, new_n815_ );
not g0679 ( new_n817_, new_n816_ );
nor g0680 ( new_n818_, N97, N113 );
nand g0681 ( new_n819_, N97, N113 );
not g0682 ( new_n820_, new_n819_ );
nor g0683 ( new_n821_, new_n820_, new_n818_ );
not g0684 ( new_n822_, new_n821_ );
nor g0685 ( new_n823_, new_n817_, new_n822_ );
nor g0686 ( new_n824_, new_n816_, new_n821_ );
nor g0687 ( new_n825_, new_n823_, new_n824_ );
nor g0688 ( new_n826_, new_n825_, keyIn_0_18 );
nand g0689 ( new_n827_, new_n825_, keyIn_0_18 );
not g0690 ( new_n828_, new_n827_ );
nor g0691 ( new_n829_, new_n828_, new_n826_ );
not g0692 ( new_n830_, new_n829_ );
nand g0693 ( new_n831_, new_n812_, new_n830_ );
nor g0694 ( new_n832_, new_n810_, new_n807_ );
nor g0695 ( new_n833_, new_n805_, keyIn_0_34 );
nor g0696 ( new_n834_, new_n832_, new_n833_ );
nand g0697 ( new_n835_, new_n834_, new_n829_ );
nand g0698 ( new_n836_, new_n835_, new_n831_ );
nor g0699 ( new_n837_, new_n836_, keyIn_0_42 );
not g0700 ( new_n838_, keyIn_0_42 );
nor g0701 ( new_n839_, new_n834_, new_n829_ );
nor g0702 ( new_n840_, new_n812_, new_n830_ );
nor g0703 ( new_n841_, new_n839_, new_n840_ );
nor g0704 ( new_n842_, new_n841_, new_n838_ );
nor g0705 ( new_n843_, new_n842_, new_n837_ );
nand g0706 ( new_n844_, new_n843_, new_n787_ );
nor g0707 ( new_n845_, new_n844_, new_n729_ );
nand g0708 ( new_n846_, new_n511_, new_n845_ );
nand g0709 ( new_n847_, new_n846_, new_n247_ );
nor g0710 ( new_n848_, new_n846_, new_n247_ );
not g0711 ( new_n849_, new_n848_ );
nand g0712 ( new_n850_, new_n849_, new_n847_ );
nand g0713 ( new_n851_, new_n850_, new_n246_ );
nand g0714 ( new_n852_, new_n851_, N1 );
not g0715 ( new_n853_, new_n847_ );
nor g0716 ( new_n854_, new_n853_, new_n848_ );
nor g0717 ( new_n855_, new_n854_, new_n400_ );
nand g0718 ( new_n856_, new_n855_, new_n216_ );
nand g0719 ( N724, new_n856_, new_n852_ );
nand g0720 ( new_n858_, new_n850_, new_n456_ );
nand g0721 ( new_n859_, new_n858_, N5 );
nor g0722 ( new_n860_, new_n854_, new_n482_ );
nand g0723 ( new_n861_, new_n860_, new_n423_ );
nand g0724 ( N725, new_n861_, new_n859_ );
nand g0725 ( new_n863_, new_n850_, new_n470_ );
nand g0726 ( new_n864_, new_n863_, N9 );
nor g0727 ( new_n865_, new_n854_, new_n397_ );
nand g0728 ( new_n866_, new_n865_, new_n366_ );
nand g0729 ( N726, new_n866_, new_n864_ );
nand g0730 ( new_n868_, new_n850_, new_n321_ );
nand g0731 ( new_n869_, new_n868_, N13 );
nor g0732 ( new_n870_, new_n854_, new_n467_ );
nand g0733 ( new_n871_, new_n870_, new_n288_ );
nand g0734 ( N727, new_n871_, new_n869_ );
not g0735 ( new_n873_, keyIn_0_57 );
nor g0736 ( new_n874_, new_n621_, new_n618_ );
nor g0737 ( new_n875_, new_n616_, keyIn_0_45 );
nor g0738 ( new_n876_, new_n874_, new_n875_ );
nor g0739 ( new_n877_, new_n726_, keyIn_0_44 );
nor g0740 ( new_n878_, new_n722_, new_n624_ );
nor g0741 ( new_n879_, new_n877_, new_n878_ );
nand g0742 ( new_n880_, new_n876_, new_n879_ );
nor g0743 ( new_n881_, new_n880_, new_n844_ );
nand g0744 ( new_n882_, new_n511_, new_n881_ );
nand g0745 ( new_n883_, new_n882_, new_n873_ );
nor g0746 ( new_n884_, new_n882_, new_n873_ );
not g0747 ( new_n885_, new_n884_ );
nand g0748 ( new_n886_, new_n885_, new_n883_ );
nand g0749 ( new_n887_, new_n886_, new_n246_ );
nand g0750 ( new_n888_, new_n887_, N17 );
not g0751 ( new_n889_, new_n883_ );
nor g0752 ( new_n890_, new_n889_, new_n884_ );
nor g0753 ( new_n891_, new_n890_, new_n400_ );
nand g0754 ( new_n892_, new_n891_, new_n218_ );
nand g0755 ( N728, new_n892_, new_n888_ );
nand g0756 ( new_n894_, new_n886_, new_n456_ );
nand g0757 ( new_n895_, new_n894_, N21 );
nor g0758 ( new_n896_, new_n890_, new_n482_ );
nand g0759 ( new_n897_, new_n896_, new_n425_ );
nand g0760 ( N729, new_n897_, new_n895_ );
nand g0761 ( new_n899_, new_n886_, new_n470_ );
nand g0762 ( new_n900_, new_n899_, N25 );
nor g0763 ( new_n901_, new_n890_, new_n397_ );
nand g0764 ( new_n902_, new_n901_, new_n368_ );
nand g0765 ( N730, new_n902_, new_n900_ );
nand g0766 ( new_n904_, new_n886_, new_n321_ );
nand g0767 ( new_n905_, new_n904_, N29 );
nor g0768 ( new_n906_, new_n890_, new_n467_ );
nand g0769 ( new_n907_, new_n906_, new_n290_ );
nand g0770 ( N731, new_n907_, new_n905_ );
not g0771 ( new_n909_, keyIn_0_58 );
not g0772 ( new_n910_, new_n781_ );
nor g0773 ( new_n911_, new_n780_, keyIn_0_43 );
nor g0774 ( new_n912_, new_n910_, new_n911_ );
not g0775 ( new_n913_, new_n837_ );
nand g0776 ( new_n914_, new_n836_, keyIn_0_42 );
nand g0777 ( new_n915_, new_n913_, new_n914_ );
nand g0778 ( new_n916_, new_n912_, new_n915_ );
nor g0779 ( new_n917_, new_n916_, new_n729_ );
nand g0780 ( new_n918_, new_n511_, new_n917_ );
nand g0781 ( new_n919_, new_n918_, new_n909_ );
nor g0782 ( new_n920_, new_n918_, new_n909_ );
not g0783 ( new_n921_, new_n920_ );
nand g0784 ( new_n922_, new_n921_, new_n919_ );
nand g0785 ( new_n923_, new_n922_, new_n246_ );
nand g0786 ( new_n924_, new_n923_, N33 );
not g0787 ( new_n925_, N33 );
not g0788 ( new_n926_, new_n919_ );
nor g0789 ( new_n927_, new_n926_, new_n920_ );
nor g0790 ( new_n928_, new_n927_, new_n400_ );
nand g0791 ( new_n929_, new_n928_, new_n925_ );
nand g0792 ( N732, new_n929_, new_n924_ );
nand g0793 ( new_n931_, new_n922_, new_n456_ );
nand g0794 ( new_n932_, new_n931_, N37 );
not g0795 ( new_n933_, N37 );
nor g0796 ( new_n934_, new_n927_, new_n482_ );
nand g0797 ( new_n935_, new_n934_, new_n933_ );
nand g0798 ( N733, new_n935_, new_n932_ );
nand g0799 ( new_n937_, new_n922_, new_n470_ );
nand g0800 ( new_n938_, new_n937_, N41 );
not g0801 ( new_n939_, N41 );
nor g0802 ( new_n940_, new_n927_, new_n397_ );
nand g0803 ( new_n941_, new_n940_, new_n939_ );
nand g0804 ( N734, new_n941_, new_n938_ );
nand g0805 ( new_n943_, new_n922_, new_n321_ );
nand g0806 ( new_n944_, new_n943_, N45 );
not g0807 ( new_n945_, N45 );
nor g0808 ( new_n946_, new_n927_, new_n467_ );
nand g0809 ( new_n947_, new_n946_, new_n945_ );
nand g0810 ( N735, new_n947_, new_n944_ );
not g0811 ( new_n949_, keyIn_0_59 );
nor g0812 ( new_n950_, new_n916_, new_n880_ );
nand g0813 ( new_n951_, new_n511_, new_n950_ );
nand g0814 ( new_n952_, new_n951_, new_n949_ );
nor g0815 ( new_n953_, new_n951_, new_n949_ );
not g0816 ( new_n954_, new_n953_ );
nand g0817 ( new_n955_, new_n954_, new_n952_ );
nand g0818 ( new_n956_, new_n955_, new_n246_ );
nand g0819 ( new_n957_, new_n956_, N49 );
not g0820 ( new_n958_, N49 );
not g0821 ( new_n959_, new_n952_ );
nor g0822 ( new_n960_, new_n959_, new_n953_ );
nor g0823 ( new_n961_, new_n960_, new_n400_ );
nand g0824 ( new_n962_, new_n961_, new_n958_ );
nand g0825 ( N736, new_n962_, new_n957_ );
nand g0826 ( new_n964_, new_n955_, new_n456_ );
nand g0827 ( new_n965_, new_n964_, N53 );
not g0828 ( new_n966_, N53 );
nor g0829 ( new_n967_, new_n960_, new_n482_ );
nand g0830 ( new_n968_, new_n967_, new_n966_ );
nand g0831 ( N737, new_n968_, new_n965_ );
nand g0832 ( new_n970_, new_n955_, new_n470_ );
nand g0833 ( new_n971_, new_n970_, N57 );
not g0834 ( new_n972_, N57 );
nor g0835 ( new_n973_, new_n960_, new_n397_ );
nand g0836 ( new_n974_, new_n973_, new_n972_ );
nand g0837 ( N738, new_n974_, new_n971_ );
nand g0838 ( new_n976_, new_n955_, new_n321_ );
nand g0839 ( new_n977_, new_n976_, N61 );
not g0840 ( new_n978_, N61 );
nor g0841 ( new_n979_, new_n960_, new_n467_ );
nand g0842 ( new_n980_, new_n979_, new_n978_ );
nand g0843 ( N739, new_n980_, new_n977_ );
not g0844 ( new_n982_, keyIn_0_60 );
not g0845 ( new_n983_, keyIn_0_55 );
not g0846 ( new_n984_, keyIn_0_51 );
nand g0847 ( new_n985_, new_n915_, new_n787_ );
nor g0848 ( new_n986_, new_n985_, new_n729_ );
nor g0849 ( new_n987_, new_n986_, new_n984_ );
not g0850 ( new_n988_, new_n729_ );
nor g0851 ( new_n989_, new_n912_, new_n843_ );
nand g0852 ( new_n990_, new_n988_, new_n989_ );
nor g0853 ( new_n991_, new_n990_, keyIn_0_51 );
nor g0854 ( new_n992_, new_n991_, new_n987_ );
nand g0855 ( new_n993_, new_n879_, new_n623_ );
nor g0856 ( new_n994_, new_n993_, new_n844_ );
nand g0857 ( new_n995_, new_n994_, keyIn_0_53 );
not g0858 ( new_n996_, keyIn_0_53 );
nor g0859 ( new_n997_, new_n912_, new_n915_ );
nor g0860 ( new_n998_, new_n876_, new_n728_ );
nand g0861 ( new_n999_, new_n997_, new_n998_ );
nand g0862 ( new_n1000_, new_n999_, new_n996_ );
nand g0863 ( new_n1001_, new_n1000_, new_n995_ );
nor g0864 ( new_n1002_, new_n992_, new_n1001_ );
not g0865 ( new_n1003_, keyIn_0_50 );
nor g0866 ( new_n1004_, new_n623_, new_n728_ );
nand g0867 ( new_n1005_, new_n989_, new_n1004_ );
nand g0868 ( new_n1006_, new_n1005_, new_n1003_ );
nor g0869 ( new_n1007_, new_n880_, new_n985_ );
nand g0870 ( new_n1008_, new_n1007_, keyIn_0_50 );
nand g0871 ( new_n1009_, new_n1006_, new_n1008_ );
not g0872 ( new_n1010_, keyIn_0_52 );
nor g0873 ( new_n1011_, new_n843_, new_n787_ );
nand g0874 ( new_n1012_, new_n998_, new_n1011_ );
nand g0875 ( new_n1013_, new_n1012_, new_n1010_ );
nor g0876 ( new_n1014_, new_n916_, new_n993_ );
nand g0877 ( new_n1015_, new_n1014_, keyIn_0_52 );
nand g0878 ( new_n1016_, new_n1015_, new_n1013_ );
nand g0879 ( new_n1017_, new_n1009_, new_n1016_ );
not g0880 ( new_n1018_, new_n1017_ );
nand g0881 ( new_n1019_, new_n1018_, new_n1002_ );
nand g0882 ( new_n1020_, new_n1019_, new_n983_ );
nand g0883 ( new_n1021_, new_n990_, keyIn_0_51 );
nand g0884 ( new_n1022_, new_n986_, new_n984_ );
nand g0885 ( new_n1023_, new_n1021_, new_n1022_ );
nor g0886 ( new_n1024_, new_n999_, new_n996_ );
nor g0887 ( new_n1025_, new_n994_, keyIn_0_53 );
nor g0888 ( new_n1026_, new_n1024_, new_n1025_ );
nand g0889 ( new_n1027_, new_n1026_, new_n1023_ );
nor g0890 ( new_n1028_, new_n1027_, new_n1017_ );
nand g0891 ( new_n1029_, new_n1028_, keyIn_0_55 );
nand g0892 ( new_n1030_, new_n1020_, new_n1029_ );
not g0893 ( new_n1031_, new_n457_ );
nor g0894 ( new_n1032_, new_n1031_, new_n487_ );
nand g0895 ( new_n1033_, new_n1030_, new_n1032_ );
nand g0896 ( new_n1034_, new_n1033_, new_n982_ );
not g0897 ( new_n1035_, new_n1034_ );
nor g0898 ( new_n1036_, new_n1033_, new_n982_ );
nor g0899 ( new_n1037_, new_n1035_, new_n1036_ );
nand g0900 ( new_n1038_, new_n1037_, new_n843_ );
nand g0901 ( new_n1039_, new_n1038_, N65 );
nor g0902 ( new_n1040_, new_n1028_, keyIn_0_55 );
nor g0903 ( new_n1041_, new_n1019_, new_n983_ );
nor g0904 ( new_n1042_, new_n1041_, new_n1040_ );
not g0905 ( new_n1043_, new_n1032_ );
nor g0906 ( new_n1044_, new_n1042_, new_n1043_ );
nand g0907 ( new_n1045_, new_n1044_, keyIn_0_60 );
nand g0908 ( new_n1046_, new_n1045_, new_n1034_ );
nor g0909 ( new_n1047_, new_n1046_, new_n915_ );
nand g0910 ( new_n1048_, new_n1047_, new_n143_ );
nand g0911 ( N740, new_n1039_, new_n1048_ );
nand g0912 ( new_n1050_, new_n1037_, new_n912_ );
nand g0913 ( new_n1051_, new_n1050_, N69 );
nor g0914 ( new_n1052_, new_n1046_, new_n787_ );
nand g0915 ( new_n1053_, new_n1052_, new_n141_ );
nand g0916 ( N741, new_n1051_, new_n1053_ );
nand g0917 ( new_n1055_, new_n1037_, new_n728_ );
nand g0918 ( new_n1056_, new_n1055_, N73 );
nor g0919 ( new_n1057_, new_n1046_, new_n879_ );
nand g0920 ( new_n1058_, new_n1057_, new_n150_ );
nand g0921 ( N742, new_n1056_, new_n1058_ );
nand g0922 ( new_n1060_, new_n1037_, new_n876_ );
nand g0923 ( new_n1061_, new_n1060_, N77 );
nor g0924 ( new_n1062_, new_n1046_, new_n623_ );
nand g0925 ( new_n1063_, new_n1062_, new_n152_ );
nand g0926 ( N743, new_n1061_, new_n1063_ );
not g0927 ( new_n1065_, keyIn_0_61 );
nor g0928 ( new_n1066_, new_n458_, new_n467_ );
nand g0929 ( new_n1067_, new_n1030_, new_n1066_ );
nand g0930 ( new_n1068_, new_n1067_, new_n1065_ );
not g0931 ( new_n1069_, new_n1068_ );
nor g0932 ( new_n1070_, new_n1067_, new_n1065_ );
nor g0933 ( new_n1071_, new_n1069_, new_n1070_ );
nand g0934 ( new_n1072_, new_n1071_, new_n843_ );
nand g0935 ( new_n1073_, new_n1072_, N81 );
not g0936 ( new_n1074_, new_n1066_ );
nor g0937 ( new_n1075_, new_n1042_, new_n1074_ );
nand g0938 ( new_n1076_, new_n1075_, keyIn_0_61 );
nand g0939 ( new_n1077_, new_n1076_, new_n1068_ );
nor g0940 ( new_n1078_, new_n1077_, new_n915_ );
nand g0941 ( new_n1079_, new_n1078_, new_n814_ );
nand g0942 ( N744, new_n1073_, new_n1079_ );
nand g0943 ( new_n1081_, new_n1071_, new_n912_ );
nand g0944 ( new_n1082_, new_n1081_, N85 );
not g0945 ( new_n1083_, N85 );
nor g0946 ( new_n1084_, new_n1077_, new_n787_ );
nand g0947 ( new_n1085_, new_n1084_, new_n1083_ );
nand g0948 ( N745, new_n1082_, new_n1085_ );
nand g0949 ( new_n1087_, new_n1071_, new_n728_ );
nand g0950 ( new_n1088_, new_n1087_, N89 );
nor g0951 ( new_n1089_, new_n1077_, new_n879_ );
nand g0952 ( new_n1090_, new_n1089_, new_n700_ );
nand g0953 ( N746, new_n1088_, new_n1090_ );
nand g0954 ( new_n1092_, new_n1071_, new_n876_ );
nand g0955 ( new_n1093_, new_n1092_, N93 );
not g0956 ( new_n1094_, N93 );
nor g0957 ( new_n1095_, new_n1077_, new_n623_ );
nand g0958 ( new_n1096_, new_n1095_, new_n1094_ );
nand g0959 ( N747, new_n1093_, new_n1096_ );
not g0960 ( new_n1098_, keyIn_0_62 );
nor g0961 ( new_n1099_, new_n487_, new_n471_ );
nand g0962 ( new_n1100_, new_n1030_, new_n1099_ );
nand g0963 ( new_n1101_, new_n1100_, new_n1098_ );
not g0964 ( new_n1102_, new_n1101_ );
nor g0965 ( new_n1103_, new_n1100_, new_n1098_ );
nor g0966 ( new_n1104_, new_n1102_, new_n1103_ );
nand g0967 ( new_n1105_, new_n1104_, new_n843_ );
nand g0968 ( new_n1106_, new_n1105_, N97 );
not g0969 ( new_n1107_, N97 );
not g0970 ( new_n1108_, new_n1099_ );
nor g0971 ( new_n1109_, new_n1042_, new_n1108_ );
nand g0972 ( new_n1110_, new_n1109_, keyIn_0_62 );
nand g0973 ( new_n1111_, new_n1110_, new_n1101_ );
nor g0974 ( new_n1112_, new_n1111_, new_n915_ );
nand g0975 ( new_n1113_, new_n1112_, new_n1107_ );
nand g0976 ( N748, new_n1106_, new_n1113_ );
nand g0977 ( new_n1115_, new_n1104_, new_n912_ );
nand g0978 ( new_n1116_, new_n1115_, N101 );
not g0979 ( new_n1117_, N101 );
nor g0980 ( new_n1118_, new_n1111_, new_n787_ );
nand g0981 ( new_n1119_, new_n1118_, new_n1117_ );
nand g0982 ( N749, new_n1116_, new_n1119_ );
nand g0983 ( new_n1121_, new_n1104_, new_n728_ );
nand g0984 ( new_n1122_, new_n1121_, N105 );
not g0985 ( new_n1123_, N105 );
nor g0986 ( new_n1124_, new_n1111_, new_n879_ );
nand g0987 ( new_n1125_, new_n1124_, new_n1123_ );
nand g0988 ( N750, new_n1122_, new_n1125_ );
nand g0989 ( new_n1127_, new_n1104_, new_n876_ );
nand g0990 ( new_n1128_, new_n1127_, N109 );
not g0991 ( new_n1129_, N109 );
nor g0992 ( new_n1130_, new_n1111_, new_n623_ );
nand g0993 ( new_n1131_, new_n1130_, new_n1129_ );
nand g0994 ( N751, new_n1128_, new_n1131_ );
not g0995 ( new_n1133_, keyIn_0_63 );
not g0996 ( new_n1134_, new_n472_ );
nor g0997 ( new_n1135_, new_n1134_, new_n467_ );
nand g0998 ( new_n1136_, new_n1030_, new_n1135_ );
nand g0999 ( new_n1137_, new_n1136_, new_n1133_ );
not g1000 ( new_n1138_, new_n1137_ );
nor g1001 ( new_n1139_, new_n1136_, new_n1133_ );
nor g1002 ( new_n1140_, new_n1138_, new_n1139_ );
nand g1003 ( new_n1141_, new_n1140_, new_n843_ );
nand g1004 ( new_n1142_, new_n1141_, N113 );
not g1005 ( new_n1143_, N113 );
not g1006 ( new_n1144_, new_n1135_ );
nor g1007 ( new_n1145_, new_n1042_, new_n1144_ );
nand g1008 ( new_n1146_, new_n1145_, keyIn_0_63 );
nand g1009 ( new_n1147_, new_n1146_, new_n1137_ );
nor g1010 ( new_n1148_, new_n1147_, new_n915_ );
nand g1011 ( new_n1149_, new_n1148_, new_n1143_ );
nand g1012 ( N752, new_n1142_, new_n1149_ );
nand g1013 ( new_n1151_, new_n1140_, new_n912_ );
nand g1014 ( new_n1152_, new_n1151_, N117 );
not g1015 ( new_n1153_, N117 );
nor g1016 ( new_n1154_, new_n1147_, new_n787_ );
nand g1017 ( new_n1155_, new_n1154_, new_n1153_ );
nand g1018 ( N753, new_n1152_, new_n1155_ );
nand g1019 ( new_n1157_, new_n1140_, new_n728_ );
nand g1020 ( new_n1158_, new_n1157_, N121 );
not g1021 ( new_n1159_, N121 );
nor g1022 ( new_n1160_, new_n1147_, new_n879_ );
nand g1023 ( new_n1161_, new_n1160_, new_n1159_ );
nand g1024 ( N754, new_n1158_, new_n1161_ );
nand g1025 ( new_n1163_, new_n1140_, new_n876_ );
nand g1026 ( new_n1164_, new_n1163_, N125 );
not g1027 ( new_n1165_, N125 );
nor g1028 ( new_n1166_, new_n1147_, new_n623_ );
nand g1029 ( new_n1167_, new_n1166_, new_n1165_ );
nand g1030 ( N755, new_n1164_, new_n1167_ );
endmodule