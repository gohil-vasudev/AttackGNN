module add_mul_combine_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_mul_0_, 
        Result_mul_1_, Result_mul_2_, Result_mul_3_, Result_mul_4_, 
        Result_mul_5_, Result_mul_6_, Result_mul_7_, Result_mul_8_, 
        Result_mul_9_, Result_mul_10_, Result_mul_11_, Result_mul_12_, 
        Result_mul_13_, Result_mul_14_, Result_mul_15_, Result_add_0_, 
        Result_add_1_, Result_add_2_, Result_add_3_, Result_add_4_, 
        Result_add_5_, Result_add_6_, Result_add_7_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_;
  wire   n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921;

  XOR2_X1 U480 ( .A(n456), .B(n457), .Z(Result_mul_9_) );
  XNOR2_X1 U481 ( .A(n458), .B(n459), .ZN(n457) );
  NAND2_X1 U482 ( .A1(a_1_), .A2(b_7_), .ZN(n459) );
  XOR2_X1 U483 ( .A(n460), .B(n461), .Z(Result_mul_8_) );
  XNOR2_X1 U484 ( .A(n462), .B(n463), .ZN(n461) );
  XOR2_X1 U485 ( .A(n464), .B(n465), .Z(Result_mul_7_) );
  NOR2_X1 U486 ( .A1(n466), .A2(n467), .ZN(Result_mul_6_) );
  NOR2_X1 U487 ( .A1(n468), .A2(n469), .ZN(n467) );
  NOR2_X1 U488 ( .A1(n465), .A2(n464), .ZN(n468) );
  XNOR2_X1 U489 ( .A(n466), .B(n470), .ZN(Result_mul_5_) );
  NAND2_X1 U490 ( .A1(n471), .A2(n472), .ZN(n470) );
  NAND2_X1 U491 ( .A1(n473), .A2(n474), .ZN(n472) );
  NAND2_X1 U492 ( .A1(n475), .A2(n476), .ZN(n474) );
  INV_X1 U493 ( .A(n477), .ZN(n473) );
  XOR2_X1 U494 ( .A(n478), .B(n479), .Z(Result_mul_4_) );
  XNOR2_X1 U495 ( .A(n480), .B(n481), .ZN(Result_mul_3_) );
  NAND2_X1 U496 ( .A1(n478), .A2(n479), .ZN(n481) );
  NOR2_X1 U497 ( .A1(n482), .A2(n483), .ZN(n480) );
  INV_X1 U498 ( .A(n484), .ZN(n483) );
  NOR2_X1 U499 ( .A1(n485), .A2(n486), .ZN(n482) );
  INV_X1 U500 ( .A(n487), .ZN(n485) );
  NAND2_X1 U501 ( .A1(n488), .A2(n489), .ZN(n487) );
  XOR2_X1 U502 ( .A(n490), .B(n491), .Z(Result_mul_2_) );
  XNOR2_X1 U503 ( .A(n492), .B(n493), .ZN(Result_mul_1_) );
  NAND2_X1 U504 ( .A1(n494), .A2(n495), .ZN(n493) );
  XNOR2_X1 U505 ( .A(n496), .B(n497), .ZN(Result_mul_14_) );
  NAND2_X1 U506 ( .A1(b_7_), .A2(a_6_), .ZN(n497) );
  XOR2_X1 U507 ( .A(n498), .B(n499), .Z(Result_mul_13_) );
  XNOR2_X1 U508 ( .A(n500), .B(n501), .ZN(n499) );
  XNOR2_X1 U509 ( .A(n502), .B(n503), .ZN(Result_mul_12_) );
  NAND2_X1 U510 ( .A1(n504), .A2(n505), .ZN(n502) );
  XOR2_X1 U511 ( .A(n506), .B(n507), .Z(Result_mul_11_) );
  XOR2_X1 U512 ( .A(n508), .B(n509), .Z(n506) );
  NOR2_X1 U513 ( .A1(n510), .A2(n511), .ZN(n509) );
  XOR2_X1 U514 ( .A(n512), .B(n513), .Z(Result_mul_10_) );
  XNOR2_X1 U515 ( .A(n514), .B(n515), .ZN(n513) );
  NAND2_X1 U516 ( .A1(b_7_), .A2(a_2_), .ZN(n515) );
  NAND3_X1 U517 ( .A1(n516), .A2(n494), .A3(n517), .ZN(Result_mul_0_) );
  NAND2_X1 U518 ( .A1(a_0_), .A2(n518), .ZN(n517) );
  INV_X1 U519 ( .A(n519), .ZN(n518) );
  NAND4_X1 U520 ( .A1(n519), .A2(n520), .A3(n521), .A4(n522), .ZN(n494) );
  NAND2_X1 U521 ( .A1(n492), .A2(n495), .ZN(n516) );
  NAND2_X1 U522 ( .A1(n523), .A2(n524), .ZN(n495) );
  NAND2_X1 U523 ( .A1(n521), .A2(n522), .ZN(n524) );
  XOR2_X1 U524 ( .A(n520), .B(n519), .Z(n523) );
  NOR2_X1 U525 ( .A1(n525), .A2(n526), .ZN(n519) );
  INV_X1 U526 ( .A(n527), .ZN(n526) );
  NAND2_X1 U527 ( .A1(n528), .A2(n529), .ZN(n527) );
  NAND2_X1 U528 ( .A1(n530), .A2(n531), .ZN(n528) );
  INV_X1 U529 ( .A(n532), .ZN(n492) );
  NAND2_X1 U530 ( .A1(n491), .A2(n490), .ZN(n532) );
  NAND3_X1 U531 ( .A1(n533), .A2(n484), .A3(n534), .ZN(n490) );
  NAND2_X1 U532 ( .A1(n535), .A2(n536), .ZN(n534) );
  NAND3_X1 U533 ( .A1(n489), .A2(n488), .A3(n486), .ZN(n484) );
  NAND3_X1 U534 ( .A1(n486), .A2(n478), .A3(n479), .ZN(n533) );
  XOR2_X1 U535 ( .A(n488), .B(n489), .Z(n479) );
  XOR2_X1 U536 ( .A(n537), .B(n538), .Z(n489) );
  XOR2_X1 U537 ( .A(n539), .B(n540), .Z(n537) );
  NAND2_X1 U538 ( .A1(n541), .A2(n542), .ZN(n488) );
  NAND2_X1 U539 ( .A1(n543), .A2(n544), .ZN(n542) );
  NAND3_X1 U540 ( .A1(n545), .A2(n471), .A3(n546), .ZN(n478) );
  NAND2_X1 U541 ( .A1(n466), .A2(n477), .ZN(n546) );
  NOR3_X1 U542 ( .A1(n465), .A2(n464), .A3(n547), .ZN(n466) );
  INV_X1 U543 ( .A(n469), .ZN(n547) );
  XOR2_X1 U544 ( .A(n475), .B(n476), .Z(n469) );
  NAND2_X1 U545 ( .A1(n548), .A2(n549), .ZN(n464) );
  NAND2_X1 U546 ( .A1(n460), .A2(n550), .ZN(n549) );
  INV_X1 U547 ( .A(n551), .ZN(n550) );
  NOR2_X1 U548 ( .A1(n463), .A2(n462), .ZN(n551) );
  XNOR2_X1 U549 ( .A(n552), .B(n553), .ZN(n460) );
  XOR2_X1 U550 ( .A(n554), .B(n555), .Z(n552) );
  NOR2_X1 U551 ( .A1(n556), .A2(n531), .ZN(n555) );
  NAND2_X1 U552 ( .A1(n462), .A2(n463), .ZN(n548) );
  NAND2_X1 U553 ( .A1(a_0_), .A2(b_7_), .ZN(n463) );
  NOR2_X1 U554 ( .A1(n557), .A2(n558), .ZN(n462) );
  INV_X1 U555 ( .A(n559), .ZN(n558) );
  NAND3_X1 U556 ( .A1(b_7_), .A2(n560), .A3(a_1_), .ZN(n559) );
  NAND2_X1 U557 ( .A1(n458), .A2(n456), .ZN(n560) );
  NOR2_X1 U558 ( .A1(n456), .A2(n458), .ZN(n557) );
  NOR2_X1 U559 ( .A1(n561), .A2(n562), .ZN(n458) );
  INV_X1 U560 ( .A(n563), .ZN(n562) );
  NAND3_X1 U561 ( .A1(a_2_), .A2(n564), .A3(b_7_), .ZN(n563) );
  NAND2_X1 U562 ( .A1(n514), .A2(n512), .ZN(n564) );
  NOR2_X1 U563 ( .A1(n512), .A2(n514), .ZN(n561) );
  NOR2_X1 U564 ( .A1(n565), .A2(n566), .ZN(n514) );
  NOR3_X1 U565 ( .A1(n510), .A2(n567), .A3(n511), .ZN(n566) );
  NOR2_X1 U566 ( .A1(n508), .A2(n507), .ZN(n567) );
  INV_X1 U567 ( .A(n568), .ZN(n565) );
  NAND2_X1 U568 ( .A1(n507), .A2(n508), .ZN(n568) );
  NAND2_X1 U569 ( .A1(n504), .A2(n569), .ZN(n508) );
  NAND2_X1 U570 ( .A1(n503), .A2(n505), .ZN(n569) );
  NAND2_X1 U571 ( .A1(n570), .A2(n571), .ZN(n505) );
  NAND2_X1 U572 ( .A1(b_7_), .A2(a_4_), .ZN(n571) );
  INV_X1 U573 ( .A(n572), .ZN(n570) );
  XNOR2_X1 U574 ( .A(n573), .B(n574), .ZN(n503) );
  XOR2_X1 U575 ( .A(n575), .B(n576), .Z(n573) );
  NAND2_X1 U576 ( .A1(a_4_), .A2(n572), .ZN(n504) );
  NAND2_X1 U577 ( .A1(n577), .A2(n578), .ZN(n572) );
  INV_X1 U578 ( .A(n579), .ZN(n578) );
  NOR2_X1 U579 ( .A1(n500), .A2(n580), .ZN(n579) );
  NOR2_X1 U580 ( .A1(n498), .A2(n501), .ZN(n580) );
  NAND2_X1 U581 ( .A1(n501), .A2(n498), .ZN(n577) );
  XOR2_X1 U582 ( .A(n581), .B(n582), .Z(n498) );
  NOR2_X1 U583 ( .A1(n583), .A2(n584), .ZN(n582) );
  NOR2_X1 U584 ( .A1(n511), .A2(n585), .ZN(n501) );
  XNOR2_X1 U585 ( .A(n586), .B(n587), .ZN(n507) );
  XNOR2_X1 U586 ( .A(n588), .B(n589), .ZN(n586) );
  XNOR2_X1 U587 ( .A(n590), .B(n591), .ZN(n512) );
  XOR2_X1 U588 ( .A(n592), .B(n593), .Z(n590) );
  XNOR2_X1 U589 ( .A(n594), .B(n595), .ZN(n456) );
  XOR2_X1 U590 ( .A(n596), .B(n597), .Z(n594) );
  XOR2_X1 U591 ( .A(n598), .B(n599), .Z(n465) );
  NAND2_X1 U592 ( .A1(n600), .A2(n601), .ZN(n598) );
  NAND3_X1 U593 ( .A1(n475), .A2(n476), .A3(n477), .ZN(n471) );
  XOR2_X1 U594 ( .A(n602), .B(n603), .Z(n477) );
  NAND2_X1 U595 ( .A1(n600), .A2(n604), .ZN(n476) );
  NAND2_X1 U596 ( .A1(n599), .A2(n601), .ZN(n604) );
  NAND2_X1 U597 ( .A1(n605), .A2(n606), .ZN(n601) );
  NAND2_X1 U598 ( .A1(a_0_), .A2(b_6_), .ZN(n606) );
  XOR2_X1 U599 ( .A(n607), .B(n608), .Z(n599) );
  XNOR2_X1 U600 ( .A(n609), .B(n610), .ZN(n608) );
  NAND2_X1 U601 ( .A1(a_1_), .A2(b_5_), .ZN(n610) );
  NAND2_X1 U602 ( .A1(a_0_), .A2(n611), .ZN(n600) );
  INV_X1 U603 ( .A(n605), .ZN(n611) );
  NOR2_X1 U604 ( .A1(n612), .A2(n613), .ZN(n605) );
  NOR3_X1 U605 ( .A1(n556), .A2(n614), .A3(n531), .ZN(n613) );
  NOR2_X1 U606 ( .A1(n553), .A2(n554), .ZN(n614) );
  INV_X1 U607 ( .A(n615), .ZN(n612) );
  NAND2_X1 U608 ( .A1(n553), .A2(n554), .ZN(n615) );
  NAND2_X1 U609 ( .A1(n616), .A2(n617), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n597), .A2(n618), .ZN(n617) );
  INV_X1 U611 ( .A(n619), .ZN(n618) );
  NOR2_X1 U612 ( .A1(n595), .A2(n596), .ZN(n619) );
  NOR2_X1 U613 ( .A1(n620), .A2(n556), .ZN(n597) );
  NAND2_X1 U614 ( .A1(n595), .A2(n596), .ZN(n616) );
  NAND2_X1 U615 ( .A1(n621), .A2(n622), .ZN(n596) );
  NAND2_X1 U616 ( .A1(n593), .A2(n623), .ZN(n622) );
  INV_X1 U617 ( .A(n624), .ZN(n623) );
  NOR2_X1 U618 ( .A1(n592), .A2(n591), .ZN(n624) );
  NOR2_X1 U619 ( .A1(n556), .A2(n510), .ZN(n593) );
  NAND2_X1 U620 ( .A1(n591), .A2(n592), .ZN(n621) );
  NAND2_X1 U621 ( .A1(n625), .A2(n626), .ZN(n592) );
  NAND2_X1 U622 ( .A1(n589), .A2(n627), .ZN(n626) );
  INV_X1 U623 ( .A(n628), .ZN(n627) );
  NOR2_X1 U624 ( .A1(n587), .A2(n588), .ZN(n628) );
  NOR2_X1 U625 ( .A1(n556), .A2(n629), .ZN(n589) );
  NAND2_X1 U626 ( .A1(n588), .A2(n587), .ZN(n625) );
  XNOR2_X1 U627 ( .A(n630), .B(n631), .ZN(n587) );
  XNOR2_X1 U628 ( .A(n632), .B(n633), .ZN(n631) );
  NOR2_X1 U629 ( .A1(n634), .A2(n635), .ZN(n588) );
  INV_X1 U630 ( .A(n636), .ZN(n635) );
  NAND2_X1 U631 ( .A1(n637), .A2(n576), .ZN(n636) );
  NAND2_X1 U632 ( .A1(n496), .A2(n638), .ZN(n576) );
  NOR2_X1 U633 ( .A1(n556), .A2(n583), .ZN(n496) );
  NAND2_X1 U634 ( .A1(n575), .A2(n574), .ZN(n637) );
  NOR2_X1 U635 ( .A1(n574), .A2(n575), .ZN(n634) );
  NOR2_X1 U636 ( .A1(n556), .A2(n585), .ZN(n575) );
  XOR2_X1 U637 ( .A(n638), .B(n639), .Z(n574) );
  XNOR2_X1 U638 ( .A(n640), .B(n641), .ZN(n591) );
  NAND2_X1 U639 ( .A1(n642), .A2(n643), .ZN(n640) );
  XNOR2_X1 U640 ( .A(n644), .B(n645), .ZN(n595) );
  XOR2_X1 U641 ( .A(n646), .B(n647), .Z(n645) );
  NAND2_X1 U642 ( .A1(a_3_), .A2(b_5_), .ZN(n647) );
  XNOR2_X1 U643 ( .A(n648), .B(n649), .ZN(n553) );
  XNOR2_X1 U644 ( .A(n650), .B(n651), .ZN(n648) );
  NOR2_X1 U645 ( .A1(n584), .A2(n620), .ZN(n651) );
  XNOR2_X1 U646 ( .A(n652), .B(n653), .ZN(n475) );
  XOR2_X1 U647 ( .A(n654), .B(n655), .Z(n652) );
  NAND2_X1 U648 ( .A1(n602), .A2(n603), .ZN(n545) );
  XNOR2_X1 U649 ( .A(n656), .B(n543), .ZN(n603) );
  XNOR2_X1 U650 ( .A(n657), .B(n658), .ZN(n543) );
  XNOR2_X1 U651 ( .A(n659), .B(n660), .ZN(n658) );
  NAND2_X1 U652 ( .A1(n541), .A2(n544), .ZN(n656) );
  NAND2_X1 U653 ( .A1(n661), .A2(n662), .ZN(n544) );
  NAND2_X1 U654 ( .A1(a_0_), .A2(b_4_), .ZN(n662) );
  NAND2_X1 U655 ( .A1(a_0_), .A2(n663), .ZN(n541) );
  INV_X1 U656 ( .A(n661), .ZN(n663) );
  NOR2_X1 U657 ( .A1(n664), .A2(n665), .ZN(n661) );
  INV_X1 U658 ( .A(n666), .ZN(n665) );
  NAND3_X1 U659 ( .A1(b_4_), .A2(n667), .A3(a_1_), .ZN(n666) );
  NAND2_X1 U660 ( .A1(n668), .A2(n669), .ZN(n667) );
  NOR2_X1 U661 ( .A1(n668), .A2(n669), .ZN(n664) );
  INV_X1 U662 ( .A(n670), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n671), .A2(n672), .ZN(n670) );
  NAND2_X1 U664 ( .A1(n653), .A2(n673), .ZN(n672) );
  INV_X1 U665 ( .A(n674), .ZN(n673) );
  NOR2_X1 U666 ( .A1(n655), .A2(n654), .ZN(n674) );
  XOR2_X1 U667 ( .A(n675), .B(n668), .Z(n653) );
  XOR2_X1 U668 ( .A(n676), .B(n677), .Z(n668) );
  XNOR2_X1 U669 ( .A(n678), .B(n679), .ZN(n676) );
  XNOR2_X1 U670 ( .A(n669), .B(n680), .ZN(n675) );
  NOR2_X1 U671 ( .A1(n681), .A2(n531), .ZN(n680) );
  NOR2_X1 U672 ( .A1(n682), .A2(n683), .ZN(n669) );
  INV_X1 U673 ( .A(n684), .ZN(n683) );
  NAND2_X1 U674 ( .A1(n685), .A2(n686), .ZN(n684) );
  NAND2_X1 U675 ( .A1(n687), .A2(n688), .ZN(n686) );
  NOR2_X1 U676 ( .A1(n688), .A2(n687), .ZN(n682) );
  NAND2_X1 U677 ( .A1(n654), .A2(n655), .ZN(n671) );
  NAND2_X1 U678 ( .A1(a_0_), .A2(b_5_), .ZN(n655) );
  NOR2_X1 U679 ( .A1(n689), .A2(n690), .ZN(n654) );
  INV_X1 U680 ( .A(n691), .ZN(n690) );
  NAND3_X1 U681 ( .A1(b_5_), .A2(n692), .A3(a_1_), .ZN(n691) );
  NAND2_X1 U682 ( .A1(n607), .A2(n609), .ZN(n692) );
  NOR2_X1 U683 ( .A1(n607), .A2(n609), .ZN(n689) );
  NOR2_X1 U684 ( .A1(n693), .A2(n694), .ZN(n609) );
  INV_X1 U685 ( .A(n695), .ZN(n694) );
  NAND3_X1 U686 ( .A1(b_5_), .A2(n696), .A3(a_2_), .ZN(n695) );
  NAND2_X1 U687 ( .A1(n650), .A2(n649), .ZN(n696) );
  NOR2_X1 U688 ( .A1(n649), .A2(n650), .ZN(n693) );
  NOR2_X1 U689 ( .A1(n697), .A2(n698), .ZN(n650) );
  NOR3_X1 U690 ( .A1(n584), .A2(n699), .A3(n510), .ZN(n698) );
  NOR2_X1 U691 ( .A1(n646), .A2(n644), .ZN(n699) );
  INV_X1 U692 ( .A(n700), .ZN(n697) );
  NAND2_X1 U693 ( .A1(n644), .A2(n646), .ZN(n700) );
  NAND2_X1 U694 ( .A1(n642), .A2(n701), .ZN(n646) );
  NAND2_X1 U695 ( .A1(n641), .A2(n643), .ZN(n701) );
  NAND2_X1 U696 ( .A1(n702), .A2(n703), .ZN(n643) );
  NAND2_X1 U697 ( .A1(b_5_), .A2(a_4_), .ZN(n703) );
  XNOR2_X1 U698 ( .A(n704), .B(n705), .ZN(n641) );
  NAND2_X1 U699 ( .A1(n706), .A2(n707), .ZN(n704) );
  INV_X1 U700 ( .A(n708), .ZN(n642) );
  NOR2_X1 U701 ( .A1(n702), .A2(n629), .ZN(n708) );
  NAND2_X1 U702 ( .A1(n709), .A2(n710), .ZN(n702) );
  NAND2_X1 U703 ( .A1(n711), .A2(n632), .ZN(n710) );
  NAND2_X1 U704 ( .A1(n638), .A2(n639), .ZN(n632) );
  NOR2_X1 U705 ( .A1(n681), .A2(n583), .ZN(n639) );
  NOR2_X1 U706 ( .A1(n584), .A2(n712), .ZN(n638) );
  NAND2_X1 U707 ( .A1(n633), .A2(n713), .ZN(n711) );
  INV_X1 U708 ( .A(n714), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n630), .A2(n714), .ZN(n709) );
  NAND2_X1 U710 ( .A1(n715), .A2(n716), .ZN(n714) );
  NAND2_X1 U711 ( .A1(n717), .A2(n718), .ZN(n716) );
  XOR2_X1 U712 ( .A(n719), .B(n720), .Z(n644) );
  XNOR2_X1 U713 ( .A(n721), .B(n722), .ZN(n719) );
  XNOR2_X1 U714 ( .A(n723), .B(n724), .ZN(n649) );
  XOR2_X1 U715 ( .A(n725), .B(n726), .Z(n723) );
  XNOR2_X1 U716 ( .A(n688), .B(n727), .ZN(n607) );
  XOR2_X1 U717 ( .A(n687), .B(n685), .Z(n727) );
  NOR2_X1 U718 ( .A1(n620), .A2(n681), .ZN(n685) );
  NOR2_X1 U719 ( .A1(n728), .A2(n729), .ZN(n687) );
  INV_X1 U720 ( .A(n730), .ZN(n729) );
  NAND2_X1 U721 ( .A1(n726), .A2(n731), .ZN(n730) );
  NAND2_X1 U722 ( .A1(n724), .A2(n725), .ZN(n731) );
  NOR2_X1 U723 ( .A1(n510), .A2(n681), .ZN(n726) );
  NOR2_X1 U724 ( .A1(n724), .A2(n725), .ZN(n728) );
  NAND2_X1 U725 ( .A1(n732), .A2(n733), .ZN(n725) );
  NAND2_X1 U726 ( .A1(n734), .A2(n722), .ZN(n733) );
  NAND2_X1 U727 ( .A1(n720), .A2(n721), .ZN(n734) );
  INV_X1 U728 ( .A(n735), .ZN(n732) );
  NOR2_X1 U729 ( .A1(n720), .A2(n721), .ZN(n735) );
  NAND2_X1 U730 ( .A1(n706), .A2(n736), .ZN(n721) );
  NAND2_X1 U731 ( .A1(n705), .A2(n707), .ZN(n736) );
  NAND2_X1 U732 ( .A1(n715), .A2(n737), .ZN(n707) );
  NAND2_X1 U733 ( .A1(b_4_), .A2(a_5_), .ZN(n737) );
  INV_X1 U734 ( .A(n738), .ZN(n715) );
  NOR2_X1 U735 ( .A1(n739), .A2(n740), .ZN(n705) );
  INV_X1 U736 ( .A(n741), .ZN(n740) );
  NAND2_X1 U737 ( .A1(n742), .A2(n743), .ZN(n741) );
  NAND2_X1 U738 ( .A1(n738), .A2(a_5_), .ZN(n706) );
  NOR2_X1 U739 ( .A1(n718), .A2(n717), .ZN(n738) );
  NAND2_X1 U740 ( .A1(b_4_), .A2(a_6_), .ZN(n717) );
  NAND2_X1 U741 ( .A1(a_7_), .A2(b_3_), .ZN(n718) );
  XNOR2_X1 U742 ( .A(n744), .B(n745), .ZN(n720) );
  XNOR2_X1 U743 ( .A(n746), .B(n739), .ZN(n745) );
  XNOR2_X1 U744 ( .A(n747), .B(n748), .ZN(n724) );
  XOR2_X1 U745 ( .A(n749), .B(n750), .Z(n747) );
  XOR2_X1 U746 ( .A(n751), .B(n752), .Z(n688) );
  XNOR2_X1 U747 ( .A(n753), .B(n754), .ZN(n751) );
  XOR2_X1 U748 ( .A(n536), .B(n535), .Z(n486) );
  XNOR2_X1 U749 ( .A(n755), .B(n756), .ZN(n535) );
  NAND2_X1 U750 ( .A1(n757), .A2(n758), .ZN(n755) );
  NAND2_X1 U751 ( .A1(n759), .A2(n760), .ZN(n536) );
  NAND2_X1 U752 ( .A1(n538), .A2(n761), .ZN(n760) );
  NAND2_X1 U753 ( .A1(n540), .A2(n539), .ZN(n761) );
  XNOR2_X1 U754 ( .A(n762), .B(n763), .ZN(n538) );
  XNOR2_X1 U755 ( .A(n764), .B(n765), .ZN(n762) );
  NOR2_X1 U756 ( .A1(n766), .A2(n531), .ZN(n765) );
  INV_X1 U757 ( .A(n767), .ZN(n759) );
  NOR2_X1 U758 ( .A1(n539), .A2(n540), .ZN(n767) );
  NOR2_X1 U759 ( .A1(n768), .A2(n769), .ZN(n540) );
  INV_X1 U760 ( .A(n770), .ZN(n769) );
  NAND2_X1 U761 ( .A1(n657), .A2(n771), .ZN(n770) );
  NAND2_X1 U762 ( .A1(n659), .A2(n660), .ZN(n771) );
  XNOR2_X1 U763 ( .A(n772), .B(n773), .ZN(n657) );
  XNOR2_X1 U764 ( .A(n774), .B(n775), .ZN(n773) );
  NOR2_X1 U765 ( .A1(n660), .A2(n659), .ZN(n768) );
  INV_X1 U766 ( .A(n776), .ZN(n659) );
  NAND2_X1 U767 ( .A1(n777), .A2(n778), .ZN(n776) );
  NAND2_X1 U768 ( .A1(n677), .A2(n779), .ZN(n778) );
  INV_X1 U769 ( .A(n780), .ZN(n779) );
  NOR2_X1 U770 ( .A1(n679), .A2(n678), .ZN(n780) );
  XNOR2_X1 U771 ( .A(n781), .B(n782), .ZN(n677) );
  XOR2_X1 U772 ( .A(n783), .B(n784), .Z(n782) );
  NAND2_X1 U773 ( .A1(n679), .A2(n678), .ZN(n777) );
  NOR2_X1 U774 ( .A1(n785), .A2(n786), .ZN(n678) );
  NOR2_X1 U775 ( .A1(n787), .A2(n754), .ZN(n786) );
  NOR2_X1 U776 ( .A1(n752), .A2(n753), .ZN(n787) );
  INV_X1 U777 ( .A(n788), .ZN(n785) );
  NAND2_X1 U778 ( .A1(n752), .A2(n753), .ZN(n788) );
  NOR2_X1 U779 ( .A1(n789), .A2(n790), .ZN(n753) );
  INV_X1 U780 ( .A(n791), .ZN(n790) );
  NAND2_X1 U781 ( .A1(n748), .A2(n792), .ZN(n791) );
  NAND2_X1 U782 ( .A1(n749), .A2(n750), .ZN(n792) );
  XNOR2_X1 U783 ( .A(n793), .B(n794), .ZN(n748) );
  NAND2_X1 U784 ( .A1(n795), .A2(n796), .ZN(n793) );
  NOR2_X1 U785 ( .A1(n750), .A2(n749), .ZN(n789) );
  NOR2_X1 U786 ( .A1(n797), .A2(n798), .ZN(n749) );
  INV_X1 U787 ( .A(n799), .ZN(n798) );
  NAND2_X1 U788 ( .A1(n739), .A2(n800), .ZN(n799) );
  NAND2_X1 U789 ( .A1(n746), .A2(n744), .ZN(n800) );
  NOR2_X1 U790 ( .A1(n742), .A2(n743), .ZN(n739) );
  NAND2_X1 U791 ( .A1(a_6_), .A2(b_3_), .ZN(n742) );
  NOR2_X1 U792 ( .A1(n744), .A2(n746), .ZN(n797) );
  NAND2_X1 U793 ( .A1(n801), .A2(n802), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n803), .A2(n804), .ZN(n802) );
  NAND2_X1 U795 ( .A1(b_2_), .A2(a_6_), .ZN(n803) );
  NAND2_X1 U796 ( .A1(b_3_), .A2(a_5_), .ZN(n744) );
  NAND2_X1 U797 ( .A1(a_4_), .A2(b_3_), .ZN(n750) );
  XOR2_X1 U798 ( .A(n805), .B(n806), .Z(n752) );
  NAND2_X1 U799 ( .A1(n807), .A2(n808), .ZN(n805) );
  NOR2_X1 U800 ( .A1(n620), .A2(n809), .ZN(n679) );
  NAND2_X1 U801 ( .A1(a_1_), .A2(b_3_), .ZN(n660) );
  NAND2_X1 U802 ( .A1(a_0_), .A2(b_3_), .ZN(n539) );
  XOR2_X1 U803 ( .A(n521), .B(n522), .Z(n491) );
  NAND2_X1 U804 ( .A1(n757), .A2(n810), .ZN(n522) );
  NAND2_X1 U805 ( .A1(n756), .A2(n758), .ZN(n810) );
  NAND2_X1 U806 ( .A1(n811), .A2(n812), .ZN(n758) );
  NAND2_X1 U807 ( .A1(a_0_), .A2(b_2_), .ZN(n812) );
  XOR2_X1 U808 ( .A(n813), .B(n814), .Z(n756) );
  NOR2_X1 U809 ( .A1(n620), .A2(n815), .ZN(n814) );
  XOR2_X1 U810 ( .A(n816), .B(n817), .Z(n813) );
  NAND2_X1 U811 ( .A1(a_0_), .A2(n818), .ZN(n757) );
  INV_X1 U812 ( .A(n811), .ZN(n818) );
  NOR2_X1 U813 ( .A1(n819), .A2(n820), .ZN(n811) );
  NOR3_X1 U814 ( .A1(n766), .A2(n821), .A3(n531), .ZN(n820) );
  NOR2_X1 U815 ( .A1(n763), .A2(n764), .ZN(n821) );
  INV_X1 U816 ( .A(n822), .ZN(n819) );
  NAND2_X1 U817 ( .A1(n763), .A2(n764), .ZN(n822) );
  NOR2_X1 U818 ( .A1(n823), .A2(n824), .ZN(n764) );
  NOR2_X1 U819 ( .A1(n825), .A2(n774), .ZN(n824) );
  NOR2_X1 U820 ( .A1(n772), .A2(n775), .ZN(n825) );
  INV_X1 U821 ( .A(n826), .ZN(n823) );
  NAND2_X1 U822 ( .A1(n772), .A2(n775), .ZN(n826) );
  NAND2_X1 U823 ( .A1(n827), .A2(n828), .ZN(n775) );
  NAND2_X1 U824 ( .A1(n829), .A2(n783), .ZN(n828) );
  NAND2_X1 U825 ( .A1(a_3_), .A2(b_2_), .ZN(n783) );
  NAND2_X1 U826 ( .A1(n781), .A2(n784), .ZN(n829) );
  INV_X1 U827 ( .A(n830), .ZN(n827) );
  NOR2_X1 U828 ( .A1(n784), .A2(n781), .ZN(n830) );
  XOR2_X1 U829 ( .A(n831), .B(n832), .Z(n781) );
  XOR2_X1 U830 ( .A(n833), .B(n834), .Z(n831) );
  NAND2_X1 U831 ( .A1(n807), .A2(n835), .ZN(n784) );
  NAND2_X1 U832 ( .A1(n806), .A2(n808), .ZN(n835) );
  NAND2_X1 U833 ( .A1(n836), .A2(n837), .ZN(n808) );
  NAND2_X1 U834 ( .A1(a_4_), .A2(b_2_), .ZN(n837) );
  INV_X1 U835 ( .A(n838), .ZN(n836) );
  XNOR2_X1 U836 ( .A(n839), .B(n840), .ZN(n806) );
  NOR2_X1 U837 ( .A1(n841), .A2(n842), .ZN(n840) );
  NAND2_X1 U838 ( .A1(a_4_), .A2(n838), .ZN(n807) );
  NAND2_X1 U839 ( .A1(n795), .A2(n843), .ZN(n838) );
  NAND2_X1 U840 ( .A1(n794), .A2(n796), .ZN(n843) );
  NAND2_X1 U841 ( .A1(n801), .A2(n844), .ZN(n796) );
  NAND2_X1 U842 ( .A1(b_2_), .A2(a_5_), .ZN(n844) );
  INV_X1 U843 ( .A(n845), .ZN(n801) );
  XNOR2_X1 U844 ( .A(n846), .B(n847), .ZN(n794) );
  NOR2_X1 U845 ( .A1(n583), .A2(n815), .ZN(n847) );
  NAND2_X1 U846 ( .A1(n845), .A2(a_5_), .ZN(n795) );
  NOR2_X1 U847 ( .A1(n743), .A2(n846), .ZN(n845) );
  NAND2_X1 U848 ( .A1(a_6_), .A2(b_1_), .ZN(n846) );
  NAND2_X1 U849 ( .A1(b_2_), .A2(a_7_), .ZN(n743) );
  XOR2_X1 U850 ( .A(n848), .B(n849), .Z(n772) );
  XNOR2_X1 U851 ( .A(n850), .B(n851), .ZN(n849) );
  XNOR2_X1 U852 ( .A(n852), .B(n853), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n854), .A2(n855), .ZN(n852) );
  NAND2_X1 U854 ( .A1(n856), .A2(n857), .ZN(n855) );
  NAND2_X1 U855 ( .A1(b_0_), .A2(a_3_), .ZN(n856) );
  XOR2_X1 U856 ( .A(n529), .B(n858), .Z(n521) );
  NOR2_X1 U857 ( .A1(n859), .A2(n525), .ZN(n858) );
  NOR3_X1 U858 ( .A1(n815), .A2(n531), .A3(n530), .ZN(n525) );
  NOR2_X1 U859 ( .A1(n860), .A2(n861), .ZN(n859) );
  NOR2_X1 U860 ( .A1(n531), .A2(n815), .ZN(n861) );
  INV_X1 U861 ( .A(n530), .ZN(n860) );
  NAND2_X1 U862 ( .A1(a_0_), .A2(b_1_), .ZN(n530) );
  NAND2_X1 U863 ( .A1(n862), .A2(n863), .ZN(n529) );
  NAND3_X1 U864 ( .A1(a_2_), .A2(n864), .A3(b_0_), .ZN(n863) );
  INV_X1 U865 ( .A(n865), .ZN(n864) );
  NOR2_X1 U866 ( .A1(n816), .A2(n817), .ZN(n865) );
  NAND2_X1 U867 ( .A1(n817), .A2(n816), .ZN(n862) );
  NAND2_X1 U868 ( .A1(n854), .A2(n866), .ZN(n816) );
  NAND2_X1 U869 ( .A1(n867), .A2(n853), .ZN(n866) );
  NAND2_X1 U870 ( .A1(n868), .A2(n869), .ZN(n853) );
  NAND2_X1 U871 ( .A1(n848), .A2(n870), .ZN(n869) );
  NAND2_X1 U872 ( .A1(n850), .A2(n851), .ZN(n870) );
  NOR2_X1 U873 ( .A1(n815), .A2(n629), .ZN(n848) );
  INV_X1 U874 ( .A(n871), .ZN(n868) );
  NOR2_X1 U875 ( .A1(n851), .A2(n850), .ZN(n871) );
  NOR2_X1 U876 ( .A1(n872), .A2(n873), .ZN(n850) );
  INV_X1 U877 ( .A(n874), .ZN(n873) );
  NAND2_X1 U878 ( .A1(n832), .A2(n875), .ZN(n874) );
  NAND2_X1 U879 ( .A1(n834), .A2(n833), .ZN(n875) );
  NOR2_X1 U880 ( .A1(n815), .A2(n585), .ZN(n832) );
  NOR2_X1 U881 ( .A1(n833), .A2(n834), .ZN(n872) );
  NOR2_X1 U882 ( .A1(n876), .A2(n841), .ZN(n834) );
  NOR2_X1 U883 ( .A1(n804), .A2(n842), .ZN(n841) );
  NAND2_X1 U884 ( .A1(b_1_), .A2(a_7_), .ZN(n804) );
  NOR2_X1 U885 ( .A1(n839), .A2(n842), .ZN(n876) );
  NAND2_X1 U886 ( .A1(b_0_), .A2(a_6_), .ZN(n842) );
  NAND2_X1 U887 ( .A1(b_1_), .A2(a_5_), .ZN(n839) );
  NAND2_X1 U888 ( .A1(a_4_), .A2(b_1_), .ZN(n833) );
  NAND2_X1 U889 ( .A1(a_3_), .A2(b_1_), .ZN(n851) );
  NAND2_X1 U890 ( .A1(n857), .A2(n510), .ZN(n867) );
  NAND3_X1 U891 ( .A1(b_0_), .A2(a_3_), .A3(n877), .ZN(n854) );
  INV_X1 U892 ( .A(n857), .ZN(n877) );
  NAND2_X1 U893 ( .A1(a_2_), .A2(b_1_), .ZN(n857) );
  XNOR2_X1 U894 ( .A(n511), .B(a_7_), .ZN(Result_add_7_) );
  NAND3_X1 U895 ( .A1(n878), .A2(n879), .A3(n500), .ZN(Result_add_6_) );
  NAND2_X1 U896 ( .A1(Result_mul_15_), .A2(n581), .ZN(n500) );
  NAND2_X1 U897 ( .A1(n880), .A2(n556), .ZN(n879) );
  XNOR2_X1 U898 ( .A(a_6_), .B(n881), .ZN(n880) );
  NAND3_X1 U899 ( .A1(n881), .A2(n712), .A3(b_6_), .ZN(n878) );
  NAND3_X1 U900 ( .A1(n882), .A2(n883), .A3(n884), .ZN(Result_add_5_) );
  NAND2_X1 U901 ( .A1(n713), .A2(n885), .ZN(n884) );
  INV_X1 U902 ( .A(n630), .ZN(n713) );
  NAND3_X1 U903 ( .A1(n886), .A2(n585), .A3(b_5_), .ZN(n883) );
  NAND2_X1 U904 ( .A1(n887), .A2(n584), .ZN(n882) );
  XNOR2_X1 U905 ( .A(a_5_), .B(n886), .ZN(n887) );
  XNOR2_X1 U906 ( .A(n888), .B(n889), .ZN(Result_add_4_) );
  NAND2_X1 U907 ( .A1(n722), .A2(n890), .ZN(n888) );
  NAND3_X1 U908 ( .A1(n891), .A2(n892), .A3(n893), .ZN(Result_add_3_) );
  NAND2_X1 U909 ( .A1(n754), .A2(n894), .ZN(n893) );
  NAND3_X1 U910 ( .A1(n895), .A2(n510), .A3(b_3_), .ZN(n892) );
  NAND2_X1 U911 ( .A1(n896), .A2(n809), .ZN(n891) );
  XNOR2_X1 U912 ( .A(n894), .B(n510), .ZN(n896) );
  XNOR2_X1 U913 ( .A(n897), .B(n898), .ZN(Result_add_2_) );
  NOR2_X1 U914 ( .A1(n899), .A2(n774), .ZN(n898) );
  NAND2_X1 U915 ( .A1(n900), .A2(n901), .ZN(Result_add_1_) );
  NAND2_X1 U916 ( .A1(n902), .A2(n903), .ZN(n901) );
  INV_X1 U917 ( .A(n904), .ZN(n902) );
  NOR2_X1 U918 ( .A1(n817), .A2(n905), .ZN(n904) );
  NAND2_X1 U919 ( .A1(n906), .A2(n907), .ZN(n900) );
  XNOR2_X1 U920 ( .A(n908), .B(a_1_), .ZN(n906) );
  XOR2_X1 U921 ( .A(n909), .B(n910), .Z(Result_add_0_) );
  NOR2_X1 U922 ( .A1(n911), .A2(n520), .ZN(n910) );
  NOR2_X1 U923 ( .A1(n912), .A2(n815), .ZN(n520) );
  INV_X1 U924 ( .A(b_0_), .ZN(n815) );
  INV_X1 U925 ( .A(a_0_), .ZN(n912) );
  NOR2_X1 U926 ( .A1(b_0_), .A2(a_0_), .ZN(n911) );
  NOR2_X1 U927 ( .A1(n905), .A2(n913), .ZN(n909) );
  NOR2_X1 U928 ( .A1(n817), .A2(n903), .ZN(n913) );
  INV_X1 U929 ( .A(n907), .ZN(n903) );
  NOR2_X1 U930 ( .A1(n774), .A2(n914), .ZN(n907) );
  NOR2_X1 U931 ( .A1(n899), .A2(n897), .ZN(n914) );
  NOR2_X1 U932 ( .A1(n754), .A2(n915), .ZN(n897) );
  NOR2_X1 U933 ( .A1(n916), .A2(n895), .ZN(n915) );
  INV_X1 U934 ( .A(n894), .ZN(n895) );
  NAND2_X1 U935 ( .A1(n722), .A2(n917), .ZN(n894) );
  NAND2_X1 U936 ( .A1(n890), .A2(n889), .ZN(n917) );
  NAND2_X1 U937 ( .A1(n630), .A2(n918), .ZN(n889) );
  NAND2_X1 U938 ( .A1(n919), .A2(n885), .ZN(n918) );
  INV_X1 U939 ( .A(n886), .ZN(n885) );
  NOR2_X1 U940 ( .A1(n581), .A2(n920), .ZN(n886) );
  NOR2_X1 U941 ( .A1(n881), .A2(n921), .ZN(n920) );
  NOR2_X1 U942 ( .A1(b_6_), .A2(a_6_), .ZN(n921) );
  INV_X1 U943 ( .A(Result_mul_15_), .ZN(n881) );
  NOR2_X1 U944 ( .A1(n511), .A2(n583), .ZN(Result_mul_15_) );
  INV_X1 U945 ( .A(a_7_), .ZN(n583) );
  INV_X1 U946 ( .A(b_7_), .ZN(n511) );
  NOR2_X1 U947 ( .A1(n556), .A2(n712), .ZN(n581) );
  INV_X1 U948 ( .A(a_6_), .ZN(n712) );
  INV_X1 U949 ( .A(b_6_), .ZN(n556) );
  NAND2_X1 U950 ( .A1(n584), .A2(n585), .ZN(n919) );
  INV_X1 U951 ( .A(a_5_), .ZN(n585) );
  INV_X1 U952 ( .A(b_5_), .ZN(n584) );
  NAND2_X1 U953 ( .A1(b_5_), .A2(a_5_), .ZN(n630) );
  NAND2_X1 U954 ( .A1(n681), .A2(n629), .ZN(n890) );
  INV_X1 U955 ( .A(a_4_), .ZN(n629) );
  INV_X1 U956 ( .A(b_4_), .ZN(n681) );
  NAND2_X1 U957 ( .A1(b_4_), .A2(a_4_), .ZN(n722) );
  NOR2_X1 U958 ( .A1(b_3_), .A2(a_3_), .ZN(n916) );
  NOR2_X1 U959 ( .A1(n510), .A2(n809), .ZN(n754) );
  INV_X1 U960 ( .A(b_3_), .ZN(n809) );
  INV_X1 U961 ( .A(a_3_), .ZN(n510) );
  NOR2_X1 U962 ( .A1(b_2_), .A2(a_2_), .ZN(n899) );
  NOR2_X1 U963 ( .A1(n620), .A2(n766), .ZN(n774) );
  INV_X1 U964 ( .A(b_2_), .ZN(n766) );
  INV_X1 U965 ( .A(a_2_), .ZN(n620) );
  NOR2_X1 U966 ( .A1(n531), .A2(n908), .ZN(n817) );
  INV_X1 U967 ( .A(b_1_), .ZN(n908) );
  INV_X1 U968 ( .A(a_1_), .ZN(n531) );
  NOR2_X1 U969 ( .A1(b_1_), .A2(a_1_), .ZN(n905) );
endmodule

