module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n702_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n313_, new_n382_, new_n583_, new_n239_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n112_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n651_, new_n433_, new_n435_, new_n109_, new_n265_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n120_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n108_, keyIn_0_26 );
not g001 ( new_n109_, N95 );
and g002 ( new_n110_, keyIn_0_14, N89 );
not g003 ( new_n111_, new_n110_ );
or g004 ( new_n112_, keyIn_0_14, N89 );
and g005 ( new_n113_, new_n111_, new_n112_ );
or g006 ( new_n114_, new_n113_, new_n109_ );
not g007 ( new_n115_, new_n114_ );
and g008 ( new_n116_, new_n115_, new_n108_ );
and g009 ( new_n117_, new_n114_, keyIn_0_26 );
or g010 ( new_n118_, new_n116_, new_n117_ );
not g011 ( new_n119_, keyIn_0_25 );
not g012 ( new_n120_, N82 );
and g013 ( new_n121_, keyIn_0_12, N76 );
not g014 ( new_n122_, new_n121_ );
or g015 ( new_n123_, keyIn_0_12, N76 );
and g016 ( new_n124_, new_n122_, new_n123_ );
or g017 ( new_n125_, new_n124_, new_n120_ );
not g018 ( new_n126_, new_n125_ );
and g019 ( new_n127_, new_n126_, new_n119_ );
and g020 ( new_n128_, new_n125_, keyIn_0_25 );
or g021 ( new_n129_, new_n127_, new_n128_ );
not g022 ( new_n130_, keyIn_0_27 );
or g023 ( new_n131_, keyIn_0_16, N102 );
not g024 ( new_n132_, N108 );
and g025 ( new_n133_, keyIn_0_16, N102 );
or g026 ( new_n134_, new_n133_, new_n132_ );
not g027 ( new_n135_, new_n134_ );
and g028 ( new_n136_, new_n135_, new_n131_ );
not g029 ( new_n137_, new_n136_ );
or g030 ( new_n138_, new_n137_, new_n130_ );
or g031 ( new_n139_, new_n136_, keyIn_0_27 );
and g032 ( new_n140_, new_n138_, new_n139_ );
and g033 ( new_n141_, new_n129_, new_n140_ );
and g034 ( new_n142_, new_n141_, new_n118_ );
not g035 ( new_n143_, keyIn_0_23 );
not g036 ( new_n144_, N56 );
not g037 ( new_n145_, N50 );
and g038 ( new_n146_, new_n145_, keyIn_0_8 );
not g039 ( new_n147_, new_n146_ );
or g040 ( new_n148_, new_n145_, keyIn_0_8 );
and g041 ( new_n149_, new_n147_, new_n148_ );
or g042 ( new_n150_, new_n149_, new_n144_ );
and g043 ( new_n151_, new_n150_, new_n143_ );
not g044 ( new_n152_, new_n150_ );
and g045 ( new_n153_, new_n152_, keyIn_0_23 );
or g046 ( new_n154_, new_n153_, new_n151_ );
not g047 ( new_n155_, keyIn_0_24 );
not g048 ( new_n156_, N69 );
or g049 ( new_n157_, keyIn_0_10, N63 );
and g050 ( new_n158_, keyIn_0_10, N63 );
not g051 ( new_n159_, new_n158_ );
and g052 ( new_n160_, new_n159_, new_n157_ );
or g053 ( new_n161_, new_n160_, new_n156_ );
not g054 ( new_n162_, new_n161_ );
or g055 ( new_n163_, new_n162_, new_n155_ );
or g056 ( new_n164_, new_n161_, keyIn_0_24 );
and g057 ( new_n165_, new_n163_, new_n164_ );
and g058 ( new_n166_, new_n154_, new_n165_ );
not g059 ( new_n167_, keyIn_0_4 );
not g060 ( new_n168_, N24 );
and g061 ( new_n169_, new_n167_, new_n168_ );
and g062 ( new_n170_, keyIn_0_4, N24 );
or g063 ( new_n171_, new_n169_, new_n170_ );
and g064 ( new_n172_, new_n171_, N30 );
or g065 ( new_n173_, new_n172_, keyIn_0_21 );
not g066 ( new_n174_, keyIn_0_21 );
not g067 ( new_n175_, N30 );
or g068 ( new_n176_, keyIn_0_4, N24 );
not g069 ( new_n177_, new_n170_ );
and g070 ( new_n178_, new_n177_, new_n176_ );
or g071 ( new_n179_, new_n178_, new_n175_ );
or g072 ( new_n180_, new_n179_, new_n174_ );
and g073 ( new_n181_, new_n173_, new_n180_ );
not g074 ( new_n182_, keyIn_0_6 );
not g075 ( new_n183_, N37 );
and g076 ( new_n184_, new_n182_, new_n183_ );
and g077 ( new_n185_, keyIn_0_6, N37 );
or g078 ( new_n186_, new_n184_, new_n185_ );
and g079 ( new_n187_, new_n186_, N43 );
or g080 ( new_n188_, new_n187_, keyIn_0_22 );
not g081 ( new_n189_, keyIn_0_22 );
not g082 ( new_n190_, N43 );
or g083 ( new_n191_, keyIn_0_6, N37 );
not g084 ( new_n192_, new_n185_ );
and g085 ( new_n193_, new_n192_, new_n191_ );
or g086 ( new_n194_, new_n193_, new_n190_ );
or g087 ( new_n195_, new_n194_, new_n189_ );
and g088 ( new_n196_, new_n188_, new_n195_ );
and g089 ( new_n197_, new_n181_, new_n196_ );
not g090 ( new_n198_, keyIn_0_18 );
not g091 ( new_n199_, N1 );
and g092 ( new_n200_, new_n199_, keyIn_0_0 );
not g093 ( new_n201_, keyIn_0_0 );
and g094 ( new_n202_, new_n201_, N1 );
or g095 ( new_n203_, new_n200_, new_n202_ );
and g096 ( new_n204_, new_n203_, N4 );
and g097 ( new_n205_, new_n204_, new_n198_ );
not g098 ( new_n206_, N4 );
or g099 ( new_n207_, new_n201_, N1 );
or g100 ( new_n208_, new_n199_, keyIn_0_0 );
and g101 ( new_n209_, new_n207_, new_n208_ );
or g102 ( new_n210_, new_n209_, new_n206_ );
and g103 ( new_n211_, new_n210_, keyIn_0_18 );
or g104 ( new_n212_, new_n211_, new_n205_ );
or g105 ( new_n213_, keyIn_0_2, N11 );
not g106 ( new_n214_, new_n213_ );
not g107 ( new_n215_, N17 );
and g108 ( new_n216_, keyIn_0_2, N11 );
or g109 ( new_n217_, new_n216_, new_n215_ );
or g110 ( new_n218_, new_n217_, new_n214_ );
and g111 ( new_n219_, new_n218_, keyIn_0_20 );
not g112 ( new_n220_, keyIn_0_20 );
not g113 ( new_n221_, new_n218_ );
and g114 ( new_n222_, new_n221_, new_n220_ );
or g115 ( new_n223_, new_n222_, new_n219_ );
and g116 ( new_n224_, new_n212_, new_n223_ );
and g117 ( new_n225_, new_n224_, new_n197_ );
and g118 ( new_n226_, new_n225_, new_n166_ );
and g119 ( new_n227_, new_n226_, new_n142_ );
and g120 ( new_n228_, new_n227_, keyIn_0_36 );
not g121 ( new_n229_, new_n228_ );
or g122 ( new_n230_, new_n227_, keyIn_0_36 );
and g123 ( N223, new_n229_, new_n230_ );
not g124 ( new_n232_, keyIn_0_60 );
not g125 ( new_n233_, keyIn_0_44 );
not g126 ( new_n234_, keyIn_0_37 );
not g127 ( new_n235_, keyIn_0_36 );
not g128 ( new_n236_, new_n227_ );
and g129 ( new_n237_, new_n236_, new_n235_ );
or g130 ( new_n238_, new_n237_, new_n228_ );
and g131 ( new_n239_, new_n238_, new_n234_ );
and g132 ( new_n240_, N223, keyIn_0_37 );
or g133 ( new_n241_, new_n239_, new_n240_ );
and g134 ( new_n242_, new_n241_, new_n129_ );
not g135 ( new_n243_, new_n129_ );
or g136 ( new_n244_, N223, keyIn_0_37 );
or g137 ( new_n245_, new_n238_, new_n234_ );
and g138 ( new_n246_, new_n245_, new_n244_ );
and g139 ( new_n247_, new_n246_, new_n243_ );
or g140 ( new_n248_, new_n242_, new_n247_ );
and g141 ( new_n249_, new_n248_, new_n233_ );
not g142 ( new_n250_, new_n249_ );
or g143 ( new_n251_, new_n248_, new_n233_ );
and g144 ( new_n252_, new_n250_, new_n251_ );
not g145 ( new_n253_, new_n252_ );
not g146 ( new_n254_, keyIn_0_33 );
not g147 ( new_n255_, N86 );
and g148 ( new_n256_, keyIn_0_13, N82 );
not g149 ( new_n257_, new_n256_ );
or g150 ( new_n258_, keyIn_0_13, N82 );
and g151 ( new_n259_, new_n257_, new_n258_ );
and g152 ( new_n260_, new_n259_, new_n255_ );
not g153 ( new_n261_, new_n260_ );
and g154 ( new_n262_, new_n261_, new_n254_ );
and g155 ( new_n263_, new_n260_, keyIn_0_33 );
or g156 ( new_n264_, new_n262_, new_n263_ );
and g157 ( new_n265_, new_n253_, new_n264_ );
not g158 ( new_n266_, new_n265_ );
or g159 ( new_n267_, new_n266_, keyIn_0_53 );
not g160 ( new_n268_, keyIn_0_53 );
or g161 ( new_n269_, new_n265_, new_n268_ );
and g162 ( new_n270_, new_n267_, new_n269_ );
and g163 ( new_n271_, new_n241_, new_n140_ );
not g164 ( new_n272_, new_n271_ );
or g165 ( new_n273_, new_n241_, new_n140_ );
and g166 ( new_n274_, new_n272_, new_n273_ );
or g167 ( new_n275_, new_n274_, keyIn_0_46 );
not g168 ( new_n276_, new_n275_ );
and g169 ( new_n277_, new_n274_, keyIn_0_46 );
or g170 ( new_n278_, new_n276_, new_n277_ );
not g171 ( new_n279_, keyIn_0_35 );
and g172 ( new_n280_, new_n132_, keyIn_0_17 );
not g173 ( new_n281_, new_n280_ );
or g174 ( new_n282_, new_n132_, keyIn_0_17 );
and g175 ( new_n283_, new_n281_, new_n282_ );
not g176 ( new_n284_, new_n283_ );
or g177 ( new_n285_, new_n284_, N112 );
and g178 ( new_n286_, new_n285_, new_n279_ );
not g179 ( new_n287_, new_n286_ );
or g180 ( new_n288_, new_n285_, new_n279_ );
and g181 ( new_n289_, new_n287_, new_n288_ );
and g182 ( new_n290_, new_n278_, new_n289_ );
and g183 ( new_n291_, new_n290_, keyIn_0_55 );
not g184 ( new_n292_, keyIn_0_55 );
not g185 ( new_n293_, new_n277_ );
and g186 ( new_n294_, new_n293_, new_n275_ );
not g187 ( new_n295_, new_n289_ );
or g188 ( new_n296_, new_n294_, new_n295_ );
and g189 ( new_n297_, new_n296_, new_n292_ );
or g190 ( new_n298_, new_n291_, new_n297_ );
not g191 ( new_n299_, keyIn_0_54 );
and g192 ( new_n300_, new_n241_, new_n118_ );
not g193 ( new_n301_, new_n300_ );
or g194 ( new_n302_, new_n241_, new_n118_ );
and g195 ( new_n303_, new_n301_, new_n302_ );
or g196 ( new_n304_, new_n303_, keyIn_0_45 );
not g197 ( new_n305_, new_n304_ );
and g198 ( new_n306_, new_n303_, keyIn_0_45 );
or g199 ( new_n307_, new_n305_, new_n306_ );
not g200 ( new_n308_, N99 );
and g201 ( new_n309_, new_n109_, keyIn_0_15 );
not g202 ( new_n310_, new_n309_ );
or g203 ( new_n311_, new_n109_, keyIn_0_15 );
and g204 ( new_n312_, new_n310_, new_n311_ );
and g205 ( new_n313_, new_n312_, new_n308_ );
not g206 ( new_n314_, new_n313_ );
and g207 ( new_n315_, new_n314_, keyIn_0_34 );
not g208 ( new_n316_, new_n315_ );
or g209 ( new_n317_, new_n314_, keyIn_0_34 );
and g210 ( new_n318_, new_n316_, new_n317_ );
and g211 ( new_n319_, new_n307_, new_n318_ );
and g212 ( new_n320_, new_n319_, new_n299_ );
not g213 ( new_n321_, new_n306_ );
and g214 ( new_n322_, new_n321_, new_n304_ );
not g215 ( new_n323_, new_n318_ );
or g216 ( new_n324_, new_n322_, new_n323_ );
and g217 ( new_n325_, new_n324_, keyIn_0_54 );
or g218 ( new_n326_, new_n320_, new_n325_ );
and g219 ( new_n327_, new_n298_, new_n326_ );
and g220 ( new_n328_, new_n327_, new_n270_ );
not g221 ( new_n329_, keyIn_0_51 );
and g222 ( new_n330_, new_n241_, new_n154_ );
not g223 ( new_n331_, new_n330_ );
or g224 ( new_n332_, new_n241_, new_n154_ );
and g225 ( new_n333_, new_n331_, new_n332_ );
or g226 ( new_n334_, new_n333_, keyIn_0_42 );
and g227 ( new_n335_, new_n333_, keyIn_0_42 );
not g228 ( new_n336_, new_n335_ );
and g229 ( new_n337_, new_n336_, new_n334_ );
not g230 ( new_n338_, keyIn_0_31 );
not g231 ( new_n339_, N60 );
and g232 ( new_n340_, keyIn_0_9, N56 );
not g233 ( new_n341_, new_n340_ );
or g234 ( new_n342_, keyIn_0_9, N56 );
and g235 ( new_n343_, new_n341_, new_n342_ );
and g236 ( new_n344_, new_n343_, new_n339_ );
not g237 ( new_n345_, new_n344_ );
and g238 ( new_n346_, new_n345_, new_n338_ );
and g239 ( new_n347_, new_n344_, keyIn_0_31 );
or g240 ( new_n348_, new_n346_, new_n347_ );
not g241 ( new_n349_, new_n348_ );
and g242 ( new_n350_, new_n337_, new_n349_ );
not g243 ( new_n351_, new_n350_ );
and g244 ( new_n352_, new_n351_, new_n329_ );
and g245 ( new_n353_, new_n350_, keyIn_0_51 );
or g246 ( new_n354_, new_n352_, new_n353_ );
and g247 ( new_n355_, new_n241_, new_n165_ );
not g248 ( new_n356_, new_n355_ );
or g249 ( new_n357_, new_n241_, new_n165_ );
and g250 ( new_n358_, new_n356_, new_n357_ );
or g251 ( new_n359_, new_n358_, keyIn_0_43 );
and g252 ( new_n360_, new_n358_, keyIn_0_43 );
not g253 ( new_n361_, new_n360_ );
and g254 ( new_n362_, new_n361_, new_n359_ );
not g255 ( new_n363_, N73 );
and g256 ( new_n364_, new_n156_, keyIn_0_11 );
not g257 ( new_n365_, new_n364_ );
or g258 ( new_n366_, new_n156_, keyIn_0_11 );
and g259 ( new_n367_, new_n365_, new_n366_ );
not g260 ( new_n368_, new_n367_ );
and g261 ( new_n369_, new_n368_, new_n363_ );
not g262 ( new_n370_, new_n369_ );
and g263 ( new_n371_, new_n370_, keyIn_0_32 );
not g264 ( new_n372_, new_n371_ );
or g265 ( new_n373_, new_n370_, keyIn_0_32 );
and g266 ( new_n374_, new_n372_, new_n373_ );
and g267 ( new_n375_, new_n362_, new_n374_ );
not g268 ( new_n376_, new_n375_ );
and g269 ( new_n377_, new_n376_, keyIn_0_52 );
not g270 ( new_n378_, keyIn_0_52 );
and g271 ( new_n379_, new_n375_, new_n378_ );
or g272 ( new_n380_, new_n377_, new_n379_ );
and g273 ( new_n381_, new_n354_, new_n380_ );
not g274 ( new_n382_, keyIn_0_47 );
and g275 ( new_n383_, new_n241_, new_n212_ );
not g276 ( new_n384_, new_n212_ );
and g277 ( new_n385_, new_n246_, new_n384_ );
or g278 ( new_n386_, new_n383_, new_n385_ );
and g279 ( new_n387_, new_n386_, keyIn_0_38 );
not g280 ( new_n388_, keyIn_0_38 );
or g281 ( new_n389_, new_n246_, new_n384_ );
or g282 ( new_n390_, new_n241_, new_n212_ );
and g283 ( new_n391_, new_n390_, new_n389_ );
and g284 ( new_n392_, new_n391_, new_n388_ );
or g285 ( new_n393_, new_n387_, new_n392_ );
not g286 ( new_n394_, keyIn_0_19 );
and g287 ( new_n395_, keyIn_0_1, N4 );
not g288 ( new_n396_, new_n395_ );
or g289 ( new_n397_, keyIn_0_1, N4 );
and g290 ( new_n398_, new_n396_, new_n397_ );
or g291 ( new_n399_, new_n398_, N8 );
and g292 ( new_n400_, new_n399_, new_n394_ );
not g293 ( new_n401_, new_n400_ );
or g294 ( new_n402_, new_n399_, new_n394_ );
and g295 ( new_n403_, new_n401_, new_n402_ );
or g296 ( new_n404_, new_n393_, new_n403_ );
or g297 ( new_n405_, new_n404_, new_n382_ );
or g298 ( new_n406_, new_n391_, new_n388_ );
or g299 ( new_n407_, new_n386_, keyIn_0_38 );
and g300 ( new_n408_, new_n407_, new_n406_ );
not g301 ( new_n409_, new_n403_ );
and g302 ( new_n410_, new_n408_, new_n409_ );
or g303 ( new_n411_, new_n410_, keyIn_0_47 );
and g304 ( new_n412_, new_n405_, new_n411_ );
not g305 ( new_n413_, keyIn_0_48 );
and g306 ( new_n414_, new_n241_, new_n223_ );
not g307 ( new_n415_, new_n223_ );
and g308 ( new_n416_, new_n246_, new_n415_ );
or g309 ( new_n417_, new_n414_, new_n416_ );
or g310 ( new_n418_, new_n417_, keyIn_0_39 );
not g311 ( new_n419_, keyIn_0_39 );
or g312 ( new_n420_, new_n246_, new_n415_ );
or g313 ( new_n421_, new_n241_, new_n223_ );
and g314 ( new_n422_, new_n421_, new_n420_ );
or g315 ( new_n423_, new_n422_, new_n419_ );
and g316 ( new_n424_, new_n418_, new_n423_ );
and g317 ( new_n425_, new_n215_, keyIn_0_3 );
not g318 ( new_n426_, new_n425_ );
or g319 ( new_n427_, new_n215_, keyIn_0_3 );
and g320 ( new_n428_, new_n426_, new_n427_ );
or g321 ( new_n429_, new_n428_, N21 );
and g322 ( new_n430_, new_n429_, keyIn_0_28 );
not g323 ( new_n431_, new_n430_ );
or g324 ( new_n432_, new_n429_, keyIn_0_28 );
and g325 ( new_n433_, new_n431_, new_n432_ );
not g326 ( new_n434_, new_n433_ );
or g327 ( new_n435_, new_n424_, new_n434_ );
or g328 ( new_n436_, new_n435_, new_n413_ );
and g329 ( new_n437_, new_n422_, new_n419_ );
and g330 ( new_n438_, new_n417_, keyIn_0_39 );
or g331 ( new_n439_, new_n438_, new_n437_ );
and g332 ( new_n440_, new_n439_, new_n433_ );
or g333 ( new_n441_, new_n440_, keyIn_0_48 );
and g334 ( new_n442_, new_n436_, new_n441_ );
and g335 ( new_n443_, new_n412_, new_n442_ );
not g336 ( new_n444_, new_n181_ );
or g337 ( new_n445_, new_n246_, new_n444_ );
or g338 ( new_n446_, new_n241_, new_n181_ );
and g339 ( new_n447_, new_n446_, new_n445_ );
and g340 ( new_n448_, new_n447_, keyIn_0_40 );
not g341 ( new_n449_, keyIn_0_40 );
and g342 ( new_n450_, new_n241_, new_n181_ );
and g343 ( new_n451_, new_n246_, new_n444_ );
or g344 ( new_n452_, new_n450_, new_n451_ );
and g345 ( new_n453_, new_n452_, new_n449_ );
or g346 ( new_n454_, new_n453_, new_n448_ );
not g347 ( new_n455_, N34 );
and g348 ( new_n456_, keyIn_0_5, N30 );
not g349 ( new_n457_, new_n456_ );
or g350 ( new_n458_, keyIn_0_5, N30 );
and g351 ( new_n459_, new_n457_, new_n458_ );
and g352 ( new_n460_, new_n459_, new_n455_ );
not g353 ( new_n461_, new_n460_ );
and g354 ( new_n462_, new_n461_, keyIn_0_29 );
not g355 ( new_n463_, new_n462_ );
or g356 ( new_n464_, new_n461_, keyIn_0_29 );
and g357 ( new_n465_, new_n463_, new_n464_ );
or g358 ( new_n466_, new_n454_, new_n465_ );
or g359 ( new_n467_, new_n466_, keyIn_0_49 );
not g360 ( new_n468_, keyIn_0_49 );
or g361 ( new_n469_, new_n452_, new_n449_ );
or g362 ( new_n470_, new_n447_, keyIn_0_40 );
and g363 ( new_n471_, new_n469_, new_n470_ );
not g364 ( new_n472_, new_n465_ );
and g365 ( new_n473_, new_n471_, new_n472_ );
or g366 ( new_n474_, new_n473_, new_n468_ );
and g367 ( new_n475_, new_n467_, new_n474_ );
and g368 ( new_n476_, new_n241_, new_n196_ );
not g369 ( new_n477_, new_n196_ );
and g370 ( new_n478_, new_n246_, new_n477_ );
or g371 ( new_n479_, new_n476_, new_n478_ );
and g372 ( new_n480_, new_n479_, keyIn_0_41 );
not g373 ( new_n481_, keyIn_0_41 );
or g374 ( new_n482_, new_n246_, new_n477_ );
or g375 ( new_n483_, new_n241_, new_n196_ );
and g376 ( new_n484_, new_n483_, new_n482_ );
and g377 ( new_n485_, new_n484_, new_n481_ );
or g378 ( new_n486_, new_n480_, new_n485_ );
not g379 ( new_n487_, keyIn_0_30 );
not g380 ( new_n488_, N47 );
and g381 ( new_n489_, new_n190_, keyIn_0_7 );
not g382 ( new_n490_, new_n489_ );
or g383 ( new_n491_, new_n190_, keyIn_0_7 );
and g384 ( new_n492_, new_n490_, new_n491_ );
and g385 ( new_n493_, new_n492_, new_n488_ );
not g386 ( new_n494_, new_n493_ );
and g387 ( new_n495_, new_n494_, new_n487_ );
and g388 ( new_n496_, new_n493_, keyIn_0_30 );
or g389 ( new_n497_, new_n495_, new_n496_ );
not g390 ( new_n498_, new_n497_ );
and g391 ( new_n499_, new_n486_, new_n498_ );
or g392 ( new_n500_, new_n499_, keyIn_0_50 );
not g393 ( new_n501_, keyIn_0_50 );
or g394 ( new_n502_, new_n484_, new_n481_ );
or g395 ( new_n503_, new_n479_, keyIn_0_41 );
and g396 ( new_n504_, new_n503_, new_n502_ );
or g397 ( new_n505_, new_n504_, new_n497_ );
or g398 ( new_n506_, new_n505_, new_n501_ );
and g399 ( new_n507_, new_n506_, new_n500_ );
and g400 ( new_n508_, new_n475_, new_n507_ );
and g401 ( new_n509_, new_n443_, new_n508_ );
and g402 ( new_n510_, new_n509_, new_n381_ );
and g403 ( new_n511_, new_n510_, new_n328_ );
and g404 ( new_n512_, new_n511_, new_n232_ );
not g405 ( new_n513_, new_n512_ );
or g406 ( new_n514_, new_n511_, new_n232_ );
and g407 ( N329, new_n513_, new_n514_ );
not g408 ( new_n516_, keyIn_0_62 );
not g409 ( new_n517_, new_n511_ );
and g410 ( new_n518_, new_n517_, keyIn_0_60 );
or g411 ( new_n519_, new_n518_, new_n512_ );
and g412 ( new_n520_, new_n519_, keyIn_0_61 );
not g413 ( new_n521_, keyIn_0_61 );
and g414 ( new_n522_, N329, new_n521_ );
or g415 ( new_n523_, new_n520_, new_n522_ );
or g416 ( new_n524_, new_n523_, new_n442_ );
not g417 ( new_n525_, new_n442_ );
or g418 ( new_n526_, N329, new_n521_ );
or g419 ( new_n527_, new_n519_, keyIn_0_61 );
and g420 ( new_n528_, new_n527_, new_n526_ );
or g421 ( new_n529_, new_n528_, new_n525_ );
and g422 ( new_n530_, new_n524_, new_n529_ );
or g423 ( new_n531_, new_n428_, N27 );
or g424 ( new_n532_, new_n424_, new_n531_ );
or g425 ( new_n533_, new_n530_, new_n532_ );
or g426 ( new_n534_, new_n523_, new_n380_ );
not g427 ( new_n535_, new_n380_ );
or g428 ( new_n536_, new_n528_, new_n535_ );
and g429 ( new_n537_, new_n534_, new_n536_ );
not g430 ( new_n538_, keyIn_0_56 );
not g431 ( new_n539_, N79 );
and g432 ( new_n540_, new_n368_, new_n539_ );
and g433 ( new_n541_, new_n362_, new_n540_ );
not g434 ( new_n542_, new_n541_ );
or g435 ( new_n543_, new_n542_, new_n538_ );
or g436 ( new_n544_, new_n541_, keyIn_0_56 );
and g437 ( new_n545_, new_n543_, new_n544_ );
or g438 ( new_n546_, new_n537_, new_n545_ );
or g439 ( new_n547_, new_n523_, new_n412_ );
not g440 ( new_n548_, new_n412_ );
or g441 ( new_n549_, new_n528_, new_n548_ );
and g442 ( new_n550_, new_n547_, new_n549_ );
or g443 ( new_n551_, new_n398_, N14 );
or g444 ( new_n552_, new_n393_, new_n551_ );
or g445 ( new_n553_, new_n550_, new_n552_ );
and g446 ( new_n554_, new_n546_, new_n553_ );
and g447 ( new_n555_, new_n554_, new_n533_ );
or g448 ( new_n556_, new_n523_, new_n507_ );
not g449 ( new_n557_, new_n507_ );
or g450 ( new_n558_, new_n528_, new_n557_ );
and g451 ( new_n559_, new_n556_, new_n558_ );
not g452 ( new_n560_, new_n492_ );
or g453 ( new_n561_, new_n560_, N53 );
or g454 ( new_n562_, new_n504_, new_n561_ );
or g455 ( new_n563_, new_n559_, new_n562_ );
or g456 ( new_n564_, new_n523_, new_n354_ );
not g457 ( new_n565_, new_n354_ );
or g458 ( new_n566_, new_n528_, new_n565_ );
and g459 ( new_n567_, new_n564_, new_n566_ );
not g460 ( new_n568_, new_n334_ );
or g461 ( new_n569_, new_n568_, new_n335_ );
not g462 ( new_n570_, new_n343_ );
or g463 ( new_n571_, new_n570_, N66 );
or g464 ( new_n572_, new_n569_, new_n571_ );
or g465 ( new_n573_, new_n567_, new_n572_ );
and g466 ( new_n574_, new_n563_, new_n573_ );
or g467 ( new_n575_, new_n523_, new_n326_ );
not g468 ( new_n576_, new_n326_ );
or g469 ( new_n577_, new_n528_, new_n576_ );
and g470 ( new_n578_, new_n575_, new_n577_ );
not g471 ( new_n579_, keyIn_0_58 );
not g472 ( new_n580_, N105 );
and g473 ( new_n581_, new_n312_, new_n580_ );
and g474 ( new_n582_, new_n307_, new_n581_ );
not g475 ( new_n583_, new_n582_ );
and g476 ( new_n584_, new_n583_, new_n579_ );
and g477 ( new_n585_, new_n582_, keyIn_0_58 );
or g478 ( new_n586_, new_n584_, new_n585_ );
or g479 ( new_n587_, new_n578_, new_n586_ );
or g480 ( new_n588_, new_n523_, new_n298_ );
not g481 ( new_n589_, new_n298_ );
or g482 ( new_n590_, new_n528_, new_n589_ );
and g483 ( new_n591_, new_n588_, new_n590_ );
not g484 ( new_n592_, keyIn_0_59 );
or g485 ( new_n593_, new_n284_, N115 );
or g486 ( new_n594_, new_n294_, new_n593_ );
not g487 ( new_n595_, new_n594_ );
and g488 ( new_n596_, new_n595_, new_n592_ );
and g489 ( new_n597_, new_n594_, keyIn_0_59 );
or g490 ( new_n598_, new_n596_, new_n597_ );
or g491 ( new_n599_, new_n591_, new_n598_ );
and g492 ( new_n600_, new_n587_, new_n599_ );
or g493 ( new_n601_, new_n523_, new_n270_ );
not g494 ( new_n602_, new_n270_ );
or g495 ( new_n603_, new_n528_, new_n602_ );
and g496 ( new_n604_, new_n601_, new_n603_ );
not g497 ( new_n605_, N92 );
and g498 ( new_n606_, new_n259_, new_n605_ );
and g499 ( new_n607_, new_n253_, new_n606_ );
not g500 ( new_n608_, new_n607_ );
and g501 ( new_n609_, new_n608_, keyIn_0_57 );
not g502 ( new_n610_, keyIn_0_57 );
and g503 ( new_n611_, new_n607_, new_n610_ );
or g504 ( new_n612_, new_n609_, new_n611_ );
or g505 ( new_n613_, new_n604_, new_n612_ );
or g506 ( new_n614_, new_n523_, new_n475_ );
not g507 ( new_n615_, new_n475_ );
or g508 ( new_n616_, new_n528_, new_n615_ );
and g509 ( new_n617_, new_n614_, new_n616_ );
not g510 ( new_n618_, new_n459_ );
or g511 ( new_n619_, new_n618_, N40 );
or g512 ( new_n620_, new_n454_, new_n619_ );
or g513 ( new_n621_, new_n617_, new_n620_ );
and g514 ( new_n622_, new_n613_, new_n621_ );
and g515 ( new_n623_, new_n600_, new_n622_ );
and g516 ( new_n624_, new_n623_, new_n574_ );
and g517 ( new_n625_, new_n624_, new_n555_ );
and g518 ( new_n626_, new_n625_, new_n516_ );
not g519 ( new_n627_, new_n626_ );
or g520 ( new_n628_, new_n625_, new_n516_ );
and g521 ( N370, new_n627_, new_n628_ );
and g522 ( new_n630_, N370, N27 );
and g523 ( new_n631_, N329, N21 );
and g524 ( new_n632_, N223, N11 );
or g525 ( new_n633_, new_n632_, new_n215_ );
or g526 ( new_n634_, new_n631_, new_n633_ );
or g527 ( new_n635_, new_n630_, new_n634_ );
and g528 ( new_n636_, N370, N40 );
and g529 ( new_n637_, N329, N34 );
and g530 ( new_n638_, N223, N24 );
or g531 ( new_n639_, new_n638_, new_n175_ );
or g532 ( new_n640_, new_n637_, new_n639_ );
or g533 ( new_n641_, new_n636_, new_n640_ );
and g534 ( new_n642_, new_n635_, new_n641_ );
and g535 ( new_n643_, N370, N53 );
and g536 ( new_n644_, N329, N47 );
and g537 ( new_n645_, N223, N37 );
or g538 ( new_n646_, new_n645_, new_n190_ );
or g539 ( new_n647_, new_n644_, new_n646_ );
or g540 ( new_n648_, new_n643_, new_n647_ );
and g541 ( new_n649_, N370, N66 );
and g542 ( new_n650_, N329, N60 );
and g543 ( new_n651_, N223, N50 );
or g544 ( new_n652_, new_n651_, new_n144_ );
or g545 ( new_n653_, new_n650_, new_n652_ );
or g546 ( new_n654_, new_n649_, new_n653_ );
and g547 ( new_n655_, new_n648_, new_n654_ );
and g548 ( new_n656_, new_n642_, new_n655_ );
and g549 ( new_n657_, N370, N79 );
and g550 ( new_n658_, N329, N73 );
and g551 ( new_n659_, N223, N63 );
or g552 ( new_n660_, new_n659_, new_n156_ );
or g553 ( new_n661_, new_n658_, new_n660_ );
or g554 ( new_n662_, new_n657_, new_n661_ );
and g555 ( new_n663_, N370, N92 );
and g556 ( new_n664_, N329, N86 );
and g557 ( new_n665_, N223, N76 );
or g558 ( new_n666_, new_n665_, new_n120_ );
or g559 ( new_n667_, new_n664_, new_n666_ );
or g560 ( new_n668_, new_n663_, new_n667_ );
and g561 ( new_n669_, new_n662_, new_n668_ );
and g562 ( new_n670_, N370, N115 );
and g563 ( new_n671_, N329, N112 );
and g564 ( new_n672_, N223, N102 );
or g565 ( new_n673_, new_n672_, new_n132_ );
or g566 ( new_n674_, new_n671_, new_n673_ );
or g567 ( new_n675_, new_n670_, new_n674_ );
and g568 ( new_n676_, N370, N105 );
and g569 ( new_n677_, N329, N99 );
and g570 ( new_n678_, N223, N89 );
or g571 ( new_n679_, new_n678_, new_n109_ );
or g572 ( new_n680_, new_n677_, new_n679_ );
or g573 ( new_n681_, new_n676_, new_n680_ );
and g574 ( new_n682_, new_n675_, new_n681_ );
and g575 ( new_n683_, new_n669_, new_n682_ );
and g576 ( new_n684_, new_n656_, new_n683_ );
not g577 ( new_n685_, new_n684_ );
and g578 ( new_n686_, new_n685_, keyIn_0_63 );
not g579 ( new_n687_, keyIn_0_63 );
and g580 ( new_n688_, new_n684_, new_n687_ );
or g581 ( new_n689_, new_n686_, new_n688_ );
and g582 ( new_n690_, N370, N14 );
and g583 ( new_n691_, N329, N8 );
and g584 ( new_n692_, N223, N1 );
or g585 ( new_n693_, new_n692_, new_n206_ );
or g586 ( new_n694_, new_n691_, new_n693_ );
or g587 ( new_n695_, new_n690_, new_n694_ );
and g588 ( N421, new_n689_, new_n695_ );
not g589 ( N430, new_n656_ );
not g590 ( new_n698_, new_n642_ );
not g591 ( new_n699_, new_n669_ );
and g592 ( new_n700_, new_n699_, new_n655_ );
or g593 ( N431, new_n700_, new_n698_ );
not g594 ( new_n702_, new_n635_ );
not g595 ( new_n703_, new_n681_ );
and g596 ( new_n704_, new_n703_, new_n668_ );
not g597 ( new_n705_, new_n648_ );
not g598 ( new_n706_, new_n662_ );
and g599 ( new_n707_, new_n706_, new_n654_ );
or g600 ( new_n708_, new_n707_, new_n705_ );
or g601 ( new_n709_, new_n708_, new_n704_ );
and g602 ( new_n710_, new_n709_, new_n641_ );
or g603 ( N432, new_n710_, new_n702_ );
endmodule