module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, 
        test_se, test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, 
        test_si4, test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, 
        test_so7, test_si8, test_so8, test_si9, test_so9, test_si10, test_so10
 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961, test_so1, test_so2, test_so3, test_so4, test_so5,
         test_so6, test_so7, test_so8, test_so9, test_so10;
  wire   g100, g101, g102, g103, g104, g1170, g1173, g1176, g1179, g1182,
         g1185, g1188, g1191, g1194, g1197, g1203, g18, g1960, g1961, g27, g28,
         g29, g30, g31, g41, g42, g43, g44, g45, g46, g47, g48, g5816, g82,
         g83, g84, g85, g8561, g8562, g8563, g8564, g8565, g8566, g86, g87,
         g872, g873, g88, g886, g889, g89, g892, g895, g898, g90, g901, g904,
         g907, g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g9451,
         g95, g96, g99, test_so10, g10722, g10664, g4556, g1289, g8943, g1882,
         n1663, g255, g312, g11257, g452, g7032, g123, g6830, g207, g8920,
         g713, g4340, g1153, n1686, g4239, g1744, g6538, g1558, g8887, g695,
         g11372, g461, n1594, g8260, g940, n1712, g11391, g976, g8432, g709,
         g6088, g1092, g6478, g1574, g6795, g1864, g11320, g369, g6500, g1580,
         g5392, g1736, n1637, g10782, n3065, g6216, g1424, g1737, g10858,
         g1672, g5914, g1077, g7590, g1231, g6656, g4, g6728, g5126, g1104,
         n1658, g7290, g1304, g6841, g243, g8041, g1499, g8766, g1444, n3064,
         g8019, g6545, g1543, g256, g315, g6533, g1534, n1632, g8820, g622,
         n1713, g8941, g1927, g10859, g1660, g6922, g278, g8772, g1436, g8433,
         g718, g6526, n1669, g10793, g554, g11333, g496, n1689, g11392, g981,
         n1720, g794, g829, g6093, g1095, g8889, g704, g7302, g1265, g6525,
         g1786, g8429, g682, g7292, g1296, g6621, n1668, g7134, n3062, g260,
         g327, g6333, g1389, n1603, g6826, g1371, g1955, g1956, g10860, g1675,
         g11483, g354, g6392, g113, g7626, g639, n1692, g10866, g1684, g8193,
         g1639, g6983, g1791, n1702, g6839, g248, n1598, g4076, g1707, g4293,
         g1759, g11482, g351, g6507, g1604, g6096, g1098, g8250, g932, n1591,
         g8282, g1896, g8435, g736, g6924, g1019, g6819, n3061, g746, g745,
         g6244, g1419, n1602, g6627, n1667, g32, n1865, g6071, g1086, g8046,
         g1486, g10707, g1730, g6198, g1504, g8051, g1470, g8024, g822, g10862,
         g1678, g8050, g174, g7133, g1766, g7930, g1801, g6832, g186, g11308,
         g959, g6918, g8769, g1407, g6909, g1868, g4940, g5404, g1718, n1611,
         g11265, g396, g6930, g1015, n1650, g4891, n3059, g6224, g1415, g7586,
         g1227, g10770, g1721, n3058, n3057, g6934, g284, g11256, g426, g6824,
         g219, g1360, n3056, DFF_126_n1, g6126, g806, g8767, g1428, g6546,
         g1564, g4238, g1741, g6823, g225, g6928, g281, g11602, g1308, g9721,
         g611, n1609, g4890, n3055, DFF_136_n1, n1586, g1217, g6524, g1589,
         g8045, g1466, g6469, g1571, g6471, g1861, g6821, n3054, g11514, g1448,
         g4480, g1133, n1706, g11610, g1333, g7843, g153, g11310, g962, g5536,
         g11331, g486, n1621, g11380, g471, n1606, g6838, g1397, n1711, g8288,
         g1950, g755, g756, g4892, n3053, DFF_157_n1, g10855, g1101, g549,
         g10898, g105, g10865, g1669, g6822, g6528, g1531, n1652, g6180, g1458,
         n1703, g10718, g572, g6912, g1011, g10719, n3051, g6234, g1411, g6099,
         g1074, g11259, g444, g8039, g1474, g6059, g1080, g5396, g1713, n1610,
         g262, g333, g6906, g269, g11266, g401, g11294, g1857, n1682, g5421,
         g9, g8649, g664, g11312, g965, g6840, g1400, n1629, g254, g309, g7202,
         g814, g6834, g231, g10795, g557, g875, g869, g6831, g1383, g8060,
         g158, g4893, g627, n1701, g7244, g1023, g6026, g259, n3050, g11608,
         g1327, g7660, g654, g6911, g293, g11640, g1346, g8777, g1633, g4274,
         g1753, g1508, g7297, g1240, g11326, g538, g11269, g416, g11325, g542,
         g10864, g1681, g11290, g374, g10798, g563, g8284, g1914, g11328, g530,
         g10800, g575, g8944, g1936, g7183, n1674, g4465, g1356, g1317, g11484,
         g357, g11263, g386, g6501, g1601, g6757, g166, g11334, g501, n1690,
         g6042, g8384, g1840, g6653, n1666, g257, g318, g5763, g5849, n3048,
         DFF_228_n1, g6929, g302, g11488, g342, g7299, g1250, g4330, g1163,
         g1958, n3047, g7257, g1032, g8775, g1432, g5770, g1453, n1628, g11486,
         g363, g261, g330, g4338, g1157, g4500, n3046, g10721, n3045,
         DFF_242_n1, g8147, g928, n1604, g6038, g11337, g516, n1620, g6045,
         g7191, g826, g861, g8774, g1627, g7293, g1292, g6907, g290, g4903,
         n3044, g6123, g6506, g1583, g11376, g466, n1646, g6542, g1561, g6551,
         g1546, g6901, g287, g10797, g560, g8505, g617, n1645, n1631, g11647,
         g336, g11340, g456, n1641, g253, g305, n1681, g11625, g345, g636, g8,
         g6502, N599, g6049, g8945, g1945, n1697, g4231, g1738, n1640, g8040,
         g1478, n3042, DFF_275_n1, g6155, g1690, n1653, g8043, g1482, g5173,
         g1110, n1677, g6916, g296, g10861, g1663, g8431, g700, g4309, g1762,
         g11485, g360, g6334, g192, g10767, g1657, g8923, g722, n1693, g7189,
         n1673, g10799, g566, g6747, n3041, g6080, g1089, g3381, g5910, g1071,
         g11393, g986, n1722, g11349, g971, g6439, g143, g9266, g1814, n1608,
         g1212, g8940, g1918, g7705, g9269, g1822, n1643, g6820, g237, g8042,
         g1462, g6759, g178, g11487, g366, g802, g837, g9124, g599, n1644,
         g11293, g1854, g11298, g944, g8287, g1941, g8047, g170, g6205, g1520,
         n1710, g8885, g686, n1676, g11305, g953, g5556, n3040, g2478, g1765,
         g10711, g1733, g7303, g5194, g1610, g7541, g1796, n1626, g11607,
         g1324, g6541, g1540, g6827, n3038, g11332, g491, n1691, g4902, n3037,
         DFF_330_n1, g6828, g213, g6516, g1781, n1659, g8938, g1900, n1675,
         g7298, g1245, n3036, g6672, n3035, DFF_336_n1, g8048, g148, g798,
         g833, g8285, g1923, n1718, g8254, g936, n1630, g11604, g1314, g849,
         g11636, g1336, g6910, g272, g8173, g1806, g8245, n1716, g8281, g1887,
         n3034, g11314, g968, g4905, n3033, g4484, g1137, n1597, g8937, g1891,
         n1657, g7300, g1255, g6002, n1588, g874, g9110, g591, n1607, g8926,
         g731, n1696, g8631, g7632, g1218, g9150, g605, n1593, g6531, n1665,
         g6786, g182, g11303, g950, g4477, g1129, n1705, g857, g11258, g448,
         g9272, g1828, n1605, g10773, g1727, g6470, g1592, g5083, g1703, g8286,
         g1932, g8773, g1624, g6054, g11260, g440, g11338, g476, n1599, g5918,
         g119, n1613, g8922, g668, n1662, g8049, g139, g4342, g1149, n1685,
         g10720, n3031, g6755, n3030, DFF_385_n1, g6897, g263, g7709, g818,
         g4255, g1747, g5543, n1622, g6915, g275, g6513, g1524, n1649, g6480,
         g1577, g6733, g810, g11264, g391, g8973, g658, n1615, g6833, g1386,
         g5996, n1587, g4473, g1125, n1708, g5755, g201, n1619, g7295, g1280,
         n1862, g6068, g1083, g7137, g650, n1709, g8779, g1636, g853, g11270,
         g421, g5529, g11306, g956, g11291, g378, g4283, g1756, g841, g6894,
         g1027, g6902, g1003, g8765, g1403, g4498, g1145, n1617, g5148, g1107,
         n1614, g7581, g1223, g11267, g406, g10936, g1811, g10784, n3029,
         g10765, g1654, g6332, g197, n1678, g6479, g1595, g6537, g1537, g8434,
         g727, g6908, g6243, n1717, g11324, g481, g3462, n1647, g11609, g1330,
         g845, g8244, g8194, g1512, n3027, g8052, g1490, g4325, g1166, g11481,
         g348, n3026, DFF_441_n1, g7301, g1260, g6035, g8059, g131, n3025,
         g6015, g258, g11330, g521, n1698, g11605, g1318, g8921, g1872, n1616,
         g8883, g677, n1656, n3024, g6523, g1549, g11300, g947, g9555, g1834,
         n1655, g6481, g1598, g4471, g1121, n1618, g11606, g1321, g11335, g506,
         g10791, g546, g8939, g1909, g6529, g1552, g10776, g1687, g6514, g1586,
         g324, g4490, g1141, n1660, g11639, g1341, g4089, g1710, g10785, n3023,
         g6179, n3022, g8053, g135, g11329, g525, n1695, g6515, g1607, g321,
         g7204, n1672, g11443, g1275, g11603, g8770, g1615, g11292, g382,
         g6331, n3020, g6900, g266, g7294, g1284, n1864, g6829, n3019, g8428,
         g673, g4904, n3018, DFF_489_n1, g8054, g162, g11268, g411, g11262,
         g431, g8283, g1905, g6193, g1515, n1627, g8776, g1630, g7143, n1671,
         g6898, g991, n1871, g7291, g1300, g11478, g339, g6000, g4264, g1750,
         g8768, g1440, g10863, g1666, g6522, g1528, n1635, g11641, g1351,
         n1721, g10780, n3017, g8044, g127, n1704, g11579, g1618, g7296, g1235,
         g6923, g299, g11261, g435, n1878, g6638, n1664, g6534, g1555, g6895,
         g995, g8771, g1621, g4506, n3016, g7441, g643, g8055, g1494, g6468,
         g1567, g8430, g691, g11327, g534, g6508, g1776, n1715, g10717, g569,
         g4334, g1160, n1585, g6679, g1, g11336, g511, n1679, g10771, g1724,
         g5445, g12, g8559, g1878, g7219, g5390, n1654, n1512, n1486, n1485,
         n1545, n1548, n1530, n1420, n1855, n1239, n1472, n1566, n1567, n1479,
         n1858, n1478, n968, n1137, n1195, n1404, n1229, n1262, n1227, n1450,
         n916, n822, n958, n918, n1054, n1116, n1159, n812, n1057, n1056, n817,
         n929, n837, n804, n1016, n1380, n926, n1385, n1391, n1564, n1231,
         n1226, n1232, n1260, n1132, n1107, n1154, n1155, n1093, n1214, n931,
         n962, n902, n1193, n1153, n1125, n1099, n917, n857, n806, n808, n1097,
         n1123, n1151, n1090, n1161, n1162, n967, n921, n898, n1055, n938,
         n1150, n1096, n1098, n1213, n1152, n836, n838, Tg1_OUT1, Tg1_OUT2,
         Tg1_OUT3, Tg1_OUT4, Tg1_OUT5, Tg1_OUT6, Tg1_OUT7, Tg1_OUT8, Tg2_OUT1,
         Tg2_OUT2, Tg2_OUT3, Tg2_OUT4, Tg2_OUT5, Tg2_OUT6, Tg2_OUT7, Tg2_OUT8,
         test_se_NOT, Trigger_select, n3, n11, n16, n18, n20, n28, n34, n36,
         n38, n53, n97, n168, n256, n343, n346, n356, n362, n366, n369, n373,
         n2457, n2458, n2459, n2460, n2461, n2462, n2465, n2467, n2468, n2469,
         n2470, n2472, n2476, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2490, n2491, n2504, n2505, n2507, n2508,
         n2509, n2510, n2511, n2513, n2514, n2515, n2519, n2520, n2521, n2522,
         n2523, n2524, n2526, n2527, n2528, n2529, n2530, n2532, n2533, n2535,
         n2537, n2538, n2544, n2546, n2548, n2550, n2551, n2552, n2554, n2557,
         n2563, n2564, n2565, n2579, n2582, n2593, n2613, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2626, n2627, n2629, n2630,
         n2631, n2632, n2633, n2636, n2638, n2639, n2640, n2641, n2642, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2657, n2658, n2660, n2662, n2663, n2664, n2665, n2667, n2668,
         n2670, n2671, n2672, n2673, n2674, n2675, n2677, n2678, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2690, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2714, n2715, n2716,
         n2717, n2719, n2720, n2721, n2722, n2725, n2726, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3021, n3028, n3032, n3039, n3043,
         n3049, n3052, n3060, n3063, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, U1586_n1, U1754_n1, U1798_n1, U1839_n1,
         U1843_n1, U1877_n1, U1908_n1, U1909_n1, U1987_n1, U2031_n1, U2035_n1,
         U2418_n1, U2468_n1, U2478_n1, U2488_n1, U2533_n1, U2534_n1, U2639_n1,
         U2641_n1, U2654_n1, U2658_n1, U2683_n1, U2699_n1, U2846_n1, U2847_n1,
         U2848_n1, U2859_n1, U2860_n1, U2861_n1, U2867_n1, U2879_n1, U2881_n1,
         U2882_n1, U2883_n1, U2884_n1, U2885_n1, U2886_n1, U2887_n1, U2888_n1,
         U2889_n1, U2890_n1, U2891_n1, U2892_n1, U2893_n1, U2894_n1, U2895_n1,
         U2896_n1, U2897_n1, U2898_n1, U2899_n1, U2900_n1, U2901_n1, U2902_n1,
         U3090_n1, U3092_n1, U3094_n1, U3096_n1, U3098_n1, U3124_n1, U3171_n1;
  assign g11489 = 1'b0;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g4205 = g1170;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4206 = g1197;
  assign g4208 = g1203;
  assign g2355 = g18;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g7744 = g27;
  assign g6285 = g28;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g8271 = g5816;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6920 = g8561;
  assign g6926 = g8562;
  assign g6932 = g8563;
  assign g6942 = g8564;
  assign g6949 = g8565;
  assign g6955 = g8566;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g5101 = g872;
  assign g8061 = g872;
  assign g5105 = g873;
  assign g8062 = g873;
  assign g6270 = g88;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g6271 = g89;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g6272 = g90;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g6273 = g91;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g6274 = g92;
  assign g4204 = g922;
  assign g4196 = g925;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g9961 = g9451;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g8984 = test_so10;

  SDFFX1 DFF_0_Q_reg ( .D(g4556), .SI(test_si1), .SE(n2846), .CLK(n2886), .Q(
        g1289), .QN(n2744) );
  SDFFX1 DFF_1_Q_reg ( .D(g8943), .SI(g1289), .SE(n2827), .CLK(n2895), .Q(
        g1882), .QN(n1663) );
  SDFFX1 DFF_2_Q_reg ( .D(g255), .SI(g1882), .SE(n2833), .CLK(n2892), .Q(g312), 
        .QN(n2683) );
  SDFFX1 DFF_3_Q_reg ( .D(g11257), .SI(g312), .SE(n2829), .CLK(n2894), .Q(g452), .QN(n2642) );
  SDFFX1 DFF_4_Q_reg ( .D(g7032), .SI(g452), .SE(n2836), .CLK(n2890), .Q(g123), 
        .QN(n2488) );
  SDFFX1 DFF_5_Q_reg ( .D(g6830), .SI(g123), .SE(n2836), .CLK(n2890), .Q(g207)
         );
  SDFFX1 DFF_6_Q_reg ( .D(g8920), .SI(g207), .SE(n2816), .CLK(n2900), .Q(g713), 
        .QN(n2515) );
  SDFFX1 DFF_7_Q_reg ( .D(g4340), .SI(g713), .SE(n2816), .CLK(n2900), .Q(g1153), .QN(n1686) );
  SDFFX1 DFF_9_Q_reg ( .D(g4239), .SI(g1153), .SE(n2816), .CLK(n2900), .Q(
        g1744) );
  SDFFX1 DFF_10_Q_reg ( .D(g6538), .SI(g1744), .SE(n2816), .CLK(n2901), .Q(
        g1558), .QN(n2552) );
  SDFFX1 DFF_11_Q_reg ( .D(g8887), .SI(g1558), .SE(n2816), .CLK(n2901), .Q(
        g695), .QN(n2711) );
  SDFFX1 DFF_12_Q_reg ( .D(g11372), .SI(g695), .SE(n2816), .CLK(n2901), .Q(
        g461), .QN(n1594) );
  SDFFX1 DFF_13_Q_reg ( .D(g8260), .SI(g461), .SE(n2831), .CLK(n2893), .Q(g940), .QN(n1712) );
  SDFFX1 DFF_14_Q_reg ( .D(g11391), .SI(g940), .SE(n2831), .CLK(n2893), .Q(
        g976), .QN(n2708) );
  SDFFX1 DFF_15_Q_reg ( .D(g8432), .SI(g976), .SE(n2812), .CLK(n2903), .Q(g709) );
  SDFFX1 DFF_16_Q_reg ( .D(g6088), .SI(g709), .SE(n2815), .CLK(n2901), .Q(
        g1092) );
  SDFFX1 DFF_17_Q_reg ( .D(g6478), .SI(g1092), .SE(n2783), .CLK(n2917), .Q(
        g1574), .QN(n2551) );
  SDFFX1 DFF_18_Q_reg ( .D(g6795), .SI(g1574), .SE(n2783), .CLK(n2917), .Q(
        g1864), .QN(n2730) );
  SDFFX1 DFF_19_Q_reg ( .D(g11320), .SI(g1864), .SE(n2776), .CLK(n2920), .Q(
        g369), .QN(n2616) );
  SDFFX1 DFF_20_Q_reg ( .D(g6500), .SI(g369), .SE(n2815), .CLK(n2901), .Q(
        g1580) );
  SDFFX1 DFF_21_Q_reg ( .D(g5392), .SI(g1580), .SE(n2814), .CLK(n2901), .Q(
        g1736) );
  SDFFX1 DFF_22_Q_reg ( .D(n38), .SI(g1736), .SE(n2814), .CLK(n2901), .Q(n1637), .QN(n4939) );
  SDFFX1 DFF_23_Q_reg ( .D(g10782), .SI(n1637), .SE(n2814), .CLK(n2901), .Q(
        n3065), .QN(n4954) );
  SDFFX1 DFF_24_Q_reg ( .D(g6216), .SI(n3065), .SE(n2814), .CLK(n2902), .Q(
        g1424) );
  SDFFX1 DFF_25_Q_reg ( .D(g1736), .SI(g1424), .SE(n2814), .CLK(n2902), .Q(
        g1737) );
  SDFFX1 DFF_26_Q_reg ( .D(g10858), .SI(g1737), .SE(n2794), .CLK(n2911), .Q(
        g1672) );
  SDFFX1 DFF_27_Q_reg ( .D(g5914), .SI(g1672), .SE(n2837), .CLK(n2890), .Q(
        g1077) );
  SDFFX1 DFF_28_Q_reg ( .D(g7590), .SI(g1077), .SE(n2818), .CLK(n2899), .Q(
        g1231) );
  SDFFX1 DFF_29_Q_reg ( .D(g6656), .SI(g1231), .SE(n2841), .CLK(n2888), .Q(g4)
         );
  SDFFX1 DFF_30_Q_reg ( .D(g6728), .SI(g4), .SE(n2833), .CLK(n2892), .Q(g4177)
         );
  SDFFX1 DFF_31_Q_reg ( .D(g5126), .SI(g4177), .SE(n2793), .CLK(n2912), .Q(
        g1104), .QN(n1658) );
  SDFFX1 DFF_32_Q_reg ( .D(g7290), .SI(g1104), .SE(n2822), .CLK(n2898), .Q(
        g1304) );
  SDFFX1 DFF_33_Q_reg ( .D(g6841), .SI(g1304), .SE(n2802), .CLK(n2908), .Q(
        g243) );
  SDFFX1 DFF_34_Q_reg ( .D(g8041), .SI(g243), .SE(n2842), .CLK(n2888), .Q(
        g1499), .QN(n2673) );
  SDFFX1 DFF_36_Q_reg ( .D(g8766), .SI(g1499), .SE(n2782), .CLK(n2917), .Q(
        g1444), .QN(n2722) );
  SDFFX1 DFF_37_Q_reg ( .D(n11), .SI(g1444), .SE(n2834), .CLK(n2891), .Q(n3064), .QN(n4933) );
  SDFFX1 DFF_38_Q_reg ( .D(g8019), .SI(n3064), .SE(n2788), .CLK(n2915), .Q(
        g4180), .QN(n2524) );
  SDFFX1 DFF_39_Q_reg ( .D(g6545), .SI(g4180), .SE(n2835), .CLK(n2891), .Q(
        g1543), .QN(n2548) );
  SDFFX1 DFF_41_Q_reg ( .D(g256), .SI(g1543), .SE(n2835), .CLK(n2891), .Q(g315), .QN(n2702) );
  SDFFX1 DFF_42_Q_reg ( .D(g6533), .SI(g315), .SE(n2769), .CLK(n2924), .Q(
        g1534), .QN(n1632) );
  SDFFX1 DFF_43_Q_reg ( .D(g8820), .SI(g1534), .SE(n2769), .CLK(n2924), .Q(
        g622), .QN(n1713) );
  SDFFX1 DFF_44_Q_reg ( .D(g8941), .SI(g622), .SE(n2826), .CLK(n2895), .Q(
        g1927), .QN(n2627) );
  SDFFX1 DFF_45_Q_reg ( .D(g10859), .SI(g1927), .SE(n2826), .CLK(n2895), .Q(
        g1660) );
  SDFFX1 DFF_46_Q_reg ( .D(g6922), .SI(g1660), .SE(n2826), .CLK(n2895), .Q(
        g278) );
  SDFFX1 DFF_47_Q_reg ( .D(g8772), .SI(g278), .SE(n2826), .CLK(n2896), .Q(
        g1436), .QN(n2719) );
  SDFFX1 DFF_48_Q_reg ( .D(g8433), .SI(g1436), .SE(n2812), .CLK(n2903), .Q(
        g718) );
  SDFFX1 DFF_49_Q_reg ( .D(g6526), .SI(g718), .SE(n2781), .CLK(n2918), .Q(
        g8985), .QN(n1669) );
  SDFFX1 DFF_50_Q_reg ( .D(g10793), .SI(g8985), .SE(n2781), .CLK(n2918), .Q(
        g554) );
  SDFFX1 DFF_51_Q_reg ( .D(g11333), .SI(g554), .SE(n2838), .CLK(n2890), .Q(
        g496), .QN(n1689) );
  SDFFX1 DFF_52_Q_reg ( .D(g11392), .SI(g496), .SE(n2830), .CLK(n2893), .Q(
        g981), .QN(n1720) );
  SDFFX1 DFF_53_Q_reg ( .D(n28), .SI(g981), .SE(n2834), .CLK(n2892), .Q(g3007)
         );
  SDFFX1 DFF_54_Q_reg ( .D(g1713), .SI(g3007), .SE(n2834), .CLK(n2892), .Q(
        test_so1) );
  SDFFX1 DFF_55_Q_reg ( .D(g794), .SI(test_si2), .SE(n2804), .CLK(n2907), .Q(
        g829) );
  SDFFX1 DFF_56_Q_reg ( .D(g6093), .SI(g829), .SE(n2763), .CLK(n2927), .Q(
        g1095) );
  SDFFX1 DFF_57_Q_reg ( .D(g8889), .SI(g1095), .SE(n2763), .CLK(n2927), .Q(
        g704), .QN(n2682) );
  SDFFX1 DFF_58_Q_reg ( .D(g7302), .SI(g704), .SE(n2822), .CLK(n2897), .Q(
        g1265), .QN(n2633) );
  SDFFX1 DFF_59_Q_reg ( .D(g6525), .SI(g1265), .SE(n2792), .CLK(n2913), .Q(
        g1786), .QN(n2735) );
  SDFFX1 DFF_60_Q_reg ( .D(g8429), .SI(g1786), .SE(n2767), .CLK(n2925), .Q(
        g682) );
  SDFFX1 DFF_61_Q_reg ( .D(g7292), .SI(g682), .SE(n2821), .CLK(n2898), .Q(
        g1296) );
  SDFFX1 DFF_62_Q_reg ( .D(g104), .SI(g1296), .SE(n2821), .CLK(n2898), .Q(
        g2602) );
  SDFFX1 DFF_63_Q_reg ( .D(g6621), .SI(g2602), .SE(n2775), .CLK(n2921), .Q(
        g8977), .QN(n1668) );
  SDFFX1 DFF_64_Q_reg ( .D(g7134), .SI(g8977), .SE(n2767), .CLK(n2925), .Q(
        n3062), .QN(n4940) );
  SDFFX1 DFF_65_Q_reg ( .D(g260), .SI(n3062), .SE(n2767), .CLK(n2925), .Q(g327), .QN(n2664) );
  SDFFX1 DFF_66_Q_reg ( .D(g6333), .SI(g327), .SE(n2806), .CLK(n2905), .Q(
        g1389), .QN(n1603) );
  SDFFX1 DFF_67_Q_reg ( .D(g6826), .SI(g1389), .SE(n2806), .CLK(n2905), .Q(
        g1371), .QN(n2675) );
  SDFFX1 DFF_68_Q_reg ( .D(g1955), .SI(g1371), .SE(n2806), .CLK(n2906), .Q(
        g1956) );
  SDFFX1 DFF_69_Q_reg ( .D(g10860), .SI(g1956), .SE(n2792), .CLK(n2912), .Q(
        g1675) );
  SDFFX1 DFF_70_Q_reg ( .D(g11483), .SI(g1675), .SE(n2801), .CLK(n2908), .Q(
        g354) );
  SDFFX1 DFF_71_Q_reg ( .D(g6392), .SI(g354), .SE(n2801), .CLK(n2908), .Q(g113) );
  SDFFX1 DFF_72_Q_reg ( .D(g7626), .SI(g113), .SE(n2767), .CLK(n2925), .Q(g639), .QN(n1692) );
  SDFFX1 DFF_73_Q_reg ( .D(g10866), .SI(g639), .SE(n2841), .CLK(n2888), .Q(
        g1684) );
  SDFFX1 DFF_74_Q_reg ( .D(g8193), .SI(g1684), .SE(n2841), .CLK(n2888), .Q(
        g1639) );
  SDFFX1 DFF_75_Q_reg ( .D(g6983), .SI(g1639), .SE(n2791), .CLK(n2913), .Q(
        g1791), .QN(n1702) );
  SDFFX1 DFF_76_Q_reg ( .D(g6839), .SI(g1791), .SE(n2773), .CLK(n2922), .Q(
        g248), .QN(n1598) );
  SDFFX1 DFF_77_Q_reg ( .D(g4076), .SI(g248), .SE(n2773), .CLK(n2922), .Q(
        g1707), .QN(n2736) );
  SDFFX1 DFF_78_Q_reg ( .D(g4293), .SI(g1707), .SE(n2791), .CLK(n2913), .Q(
        g1759), .QN(n2717) );
  SDFFX1 DFF_79_Q_reg ( .D(g11482), .SI(g1759), .SE(n2790), .CLK(n2913), .Q(
        g351) );
  SDFFX1 DFF_80_Q_reg ( .D(g1956), .SI(g351), .SE(n2790), .CLK(n2913), .Q(
        g1957) );
  SDFFX1 DFF_81_Q_reg ( .D(g6507), .SI(g1957), .SE(n2790), .CLK(n2913), .Q(
        g1604) );
  SDFFX1 DFF_82_Q_reg ( .D(g6096), .SI(g1604), .SE(n2790), .CLK(n2914), .Q(
        g1098) );
  SDFFX1 DFF_83_Q_reg ( .D(g8250), .SI(g1098), .SE(n2790), .CLK(n2914), .Q(
        g932), .QN(n1591) );
  SDFFX1 DFF_85_Q_reg ( .D(g8282), .SI(g932), .SE(n2765), .CLK(n2926), .Q(
        g1896) );
  SDFFX1 DFF_86_Q_reg ( .D(g8435), .SI(g1896), .SE(n2811), .CLK(n2903), .Q(
        g736), .QN(n2694) );
  SDFFX1 DFF_87_Q_reg ( .D(g6924), .SI(g736), .SE(n2790), .CLK(n2914), .Q(
        g1019), .QN(n2619) );
  SDFFX1 DFF_88_Q_reg ( .D(g6819), .SI(g1019), .SE(n2789), .CLK(n2914), .Q(
        n3061), .QN(n4941) );
  SDFFX1 DFF_89_Q_reg ( .D(g746), .SI(n3061), .SE(n2785), .CLK(n2916), .Q(g745), .QN(n2505) );
  SDFFX1 DFF_90_Q_reg ( .D(g6244), .SI(g745), .SE(n2785), .CLK(n2916), .Q(
        g1419), .QN(n1602) );
  SDFFX1 DFF_91_Q_reg ( .D(g6627), .SI(g1419), .SE(n2775), .CLK(n2921), .Q(
        g8979), .QN(n1667) );
  SDFFX1 DFF_92_Q_reg ( .D(n2747), .SI(g8979), .SE(n2840), .CLK(n2888), .Q(g32), .QN(n4937) );
  SDFFX1 DFF_93_Q_reg ( .D(g3007), .SI(g32), .SE(n2840), .CLK(n2888), .Q(n1865), .QN(n2480) );
  SDFFX1 DFF_94_Q_reg ( .D(g6071), .SI(n1865), .SE(n2800), .CLK(n2908), .Q(
        g1086) );
  SDFFX1 DFF_95_Q_reg ( .D(g8046), .SI(g1086), .SE(n2836), .CLK(n2891), .Q(
        g1486), .QN(n2647) );
  SDFFX1 DFF_96_Q_reg ( .D(g10707), .SI(g1486), .SE(n2799), .CLK(n2909), .Q(
        g1730), .QN(n2467) );
  SDFFX1 DFF_97_Q_reg ( .D(g6198), .SI(g1730), .SE(n2799), .CLK(n2909), .Q(
        g1504), .QN(n2529) );
  SDFFX1 DFF_98_Q_reg ( .D(g8051), .SI(g1504), .SE(n2797), .CLK(n2910), .Q(
        g1470) );
  SDFFX1 DFF_99_Q_reg ( .D(g8024), .SI(g1470), .SE(n2797), .CLK(n2910), .Q(
        g822), .QN(n2740) );
  SDFFX1 DFF_100_Q_reg ( .D(g29), .SI(g822), .SE(n2797), .CLK(n2910), .Q(g2609) );
  SDFFX1 DFF_101_Q_reg ( .D(g10862), .SI(g2609), .SE(n2797), .CLK(n2910), .Q(
        g1678) );
  SDFFX1 DFF_102_Q_reg ( .D(g8050), .SI(g1678), .SE(n2796), .CLK(n2910), .Q(
        g174), .QN(n2741) );
  SDFFX1 DFF_103_Q_reg ( .D(g7133), .SI(g174), .SE(n2796), .CLK(n2910), .Q(
        g1766), .QN(n2728) );
  SDFFX1 DFF_104_Q_reg ( .D(g7930), .SI(g1766), .SE(n2791), .CLK(n2913), .Q(
        g1801), .QN(n2733) );
  SDFFX1 DFF_105_Q_reg ( .D(g6832), .SI(g1801), .SE(n2777), .CLK(n2920), .Q(
        g186), .QN(n2511) );
  SDFFX1 DFF_106_Q_reg ( .D(g11308), .SI(g186), .SE(n2771), .CLK(n2923), .Q(
        g959) );
  SDFFX1 DFF_108_Q_reg ( .D(g6918), .SI(g959), .SE(n2763), .CLK(n2927), .Q(
        test_so2) );
  SDFFX1 DFF_109_Q_reg ( .D(g8769), .SI(test_si3), .SE(n2777), .CLK(n2920), 
        .Q(g1407), .QN(n2532) );
  SDFFX1 DFF_111_Q_reg ( .D(g6909), .SI(g1407), .SE(n2839), .CLK(n2889), .Q(
        g1868) );
  SDFFX1 DFF_112_Q_reg ( .D(g4940), .SI(g1868), .SE(n2839), .CLK(n2889), .Q(
        g4173), .QN(n2521) );
  SDFFX1 DFF_113_Q_reg ( .D(g5404), .SI(g4173), .SE(n2795), .CLK(n2911), .Q(
        g1718), .QN(n1611) );
  SDFFX1 DFF_114_Q_reg ( .D(g11265), .SI(g1718), .SE(n2830), .CLK(n2894), .Q(
        g396) );
  SDFFX1 DFF_115_Q_reg ( .D(g6930), .SI(g396), .SE(n2762), .CLK(n2927), .Q(
        g1015), .QN(n2618) );
  SDFFX1 DFF_116_Q_reg ( .D(n53), .SI(g1015), .SE(n2762), .CLK(n2927), .Q(
        n1650) );
  SDFFX1 DFF_117_Q_reg ( .D(g4891), .SI(n1650), .SE(n2819), .CLK(n2899), .Q(
        n3059) );
  SDFFX1 DFF_118_Q_reg ( .D(g6224), .SI(n3059), .SE(n2784), .CLK(n2917), .Q(
        g1415), .QN(n2527) );
  SDFFX1 DFF_119_Q_reg ( .D(g7586), .SI(g1415), .SE(n2845), .CLK(n2886), .Q(
        g1227), .QN(n2507) );
  SDFFX1 DFF_120_Q_reg ( .D(g10770), .SI(g1227), .SE(n2845), .CLK(n2886), .Q(
        g1721), .QN(n2487) );
  SDFFX1 DFF_121_Q_reg ( .D(g2986), .SI(g1721), .SE(n2831), .CLK(n2893), .Q(
        n3058), .QN(n4934) );
  SDFFX1 DFF_122_Q_reg ( .D(n2753), .SI(n3058), .SE(n2831), .CLK(n2893), .Q(
        n3057) );
  SDFFX1 DFF_123_Q_reg ( .D(g6934), .SI(n3057), .SE(n2843), .CLK(n2887), .Q(
        g284), .QN(n2565) );
  SDFFX1 DFF_124_Q_reg ( .D(g11256), .SI(g284), .SE(n2830), .CLK(n2893), .Q(
        g426), .QN(n2701) );
  SDFFX1 DFF_125_Q_reg ( .D(g6824), .SI(g426), .SE(n2806), .CLK(n2906), .Q(
        g219), .QN(n2514) );
  SDFFX1 DFF_126_Q_reg ( .D(g1360), .SI(g219), .SE(n2794), .CLK(n2912), .Q(
        n3056), .QN(DFF_126_n1) );
  SDFFX1 DFF_127_Q_reg ( .D(g6126), .SI(n3056), .SE(n2782), .CLK(n2918), .Q(
        g806), .QN(n2726) );
  SDFFX1 DFF_128_Q_reg ( .D(g8767), .SI(g806), .SE(n2782), .CLK(n2918), .Q(
        g1428), .QN(n2721) );
  SDFFX1 DFF_129_Q_reg ( .D(g102), .SI(g1428), .SE(n2782), .CLK(n2918), .Q(
        g2605) );
  SDFFX1 DFF_130_Q_reg ( .D(g6546), .SI(g2605), .SE(n2766), .CLK(n2925), .Q(
        g1564), .QN(n2546) );
  SDFFX1 DFF_131_Q_reg ( .D(g4238), .SI(g1564), .SE(n2810), .CLK(n2904), .Q(
        g1741) );
  SDFFX1 DFF_132_Q_reg ( .D(g6823), .SI(g1741), .SE(n2810), .CLK(n2904), .Q(
        g225) );
  SDFFX1 DFF_133_Q_reg ( .D(g6928), .SI(g225), .SE(n2770), .CLK(n2923), .Q(
        g281), .QN(n2564) );
  SDFFX1 DFF_134_Q_reg ( .D(g11602), .SI(g281), .SE(n2770), .CLK(n2923), .Q(
        g1308), .QN(n2479) );
  SDFFX1 DFF_135_Q_reg ( .D(g9721), .SI(g1308), .SE(n2820), .CLK(n2899), .Q(
        g611), .QN(n1609) );
  SDFFX1 DFF_136_Q_reg ( .D(g4890), .SI(g611), .SE(n2820), .CLK(n2899), .Q(
        n3055), .QN(DFF_136_n1) );
  SDFFX1 DFF_137_Q_reg ( .D(n1586), .SI(n3055), .SE(n2820), .CLK(n2899), .Q(
        g1217) );
  SDFFX1 DFF_138_Q_reg ( .D(g6524), .SI(g1217), .SE(n2797), .CLK(n2910), .Q(
        g1589) );
  SDFFX1 DFF_139_Q_reg ( .D(g8045), .SI(g1589), .SE(n2797), .CLK(n2910), .Q(
        g1466), .QN(n2651) );
  SDFFX1 DFF_140_Q_reg ( .D(g6469), .SI(g1466), .SE(n2785), .CLK(n2916), .Q(
        g1571), .QN(n2544) );
  SDFFX1 DFF_141_Q_reg ( .D(g6471), .SI(g1571), .SE(n2785), .CLK(n2916), .Q(
        g1861), .QN(n2732) );
  SDFFX1 DFF_142_Q_reg ( .D(g6821), .SI(g1861), .SE(n2784), .CLK(n2916), .Q(
        n3054), .QN(n4942) );
  SDFFX1 DFF_143_Q_reg ( .D(g11514), .SI(n3054), .SE(n2783), .CLK(n2917), .Q(
        g1448), .QN(n2653) );
  SDFFX1 DFF_145_Q_reg ( .D(g4480), .SI(g1448), .SE(n2783), .CLK(n2917), .Q(
        g1133), .QN(n1706) );
  SDFFX1 DFF_146_Q_reg ( .D(g11610), .SI(g1133), .SE(n2771), .CLK(n2923), .Q(
        g1333), .QN(n2478) );
  SDFFX1 DFF_147_Q_reg ( .D(g7843), .SI(g1333), .SE(n2771), .CLK(n2923), .Q(
        g153), .QN(n2670) );
  SDFFX1 DFF_148_Q_reg ( .D(g11310), .SI(g153), .SE(n2771), .CLK(n2923), .Q(
        g962) );
  SDFFX1 DFF_149_Q_reg ( .D(g5536), .SI(g962), .SE(n2838), .CLK(n2889), .Q(
        g4175) );
  SDFFX1 DFF_150_Q_reg ( .D(g28), .SI(g4175), .SE(n2838), .CLK(n2889), .Q(
        g2603) );
  SDFFX1 DFF_151_Q_reg ( .D(g11331), .SI(g2603), .SE(n2838), .CLK(n2890), .Q(
        g486), .QN(n1621) );
  SDFFX1 DFF_152_Q_reg ( .D(g11380), .SI(g486), .SE(n2786), .CLK(n2915), .Q(
        g471), .QN(n1606) );
  SDFFX1 DFF_153_Q_reg ( .D(g6838), .SI(g471), .SE(n2786), .CLK(n2915), .Q(
        g1397), .QN(n1711) );
  SDFFX1 DFF_154_Q_reg ( .D(g103), .SI(g1397), .SE(n2786), .CLK(n2915), .Q(
        g2606) );
  SDFFX1 DFF_155_Q_reg ( .D(g8288), .SI(g2606), .SE(n2786), .CLK(n2916), .Q(
        g1950), .QN(n2696) );
  SDFFX1 DFF_156_Q_reg ( .D(g755), .SI(g1950), .SE(n2786), .CLK(n2916), .Q(
        g756) );
  SDFFX1 DFF_157_Q_reg ( .D(g4892), .SI(g756), .SE(n2819), .CLK(n2899), .Q(
        n3053), .QN(DFF_157_n1) );
  SDFFX1 DFF_159_Q_reg ( .D(g10855), .SI(g1101), .SE(n2793), .CLK(n2912), .Q(
        g549) );
  SDFFX1 DFF_161_Q_reg ( .D(g10898), .SI(g549), .SE(n2844), .CLK(n2886), .Q(
        g105), .QN(n2483) );
  SDFFX1 DFF_162_Q_reg ( .D(g10865), .SI(g105), .SE(n2844), .CLK(n2886), .Q(
        g1669) );
  SDFFX1 DFF_163_Q_reg ( .D(g6822), .SI(g1669), .SE(n2844), .CLK(n2887), .Q(
        test_so3), .QN(n2674) );
  SDFFX1 DFF_164_Q_reg ( .D(g6528), .SI(test_si4), .SE(n2770), .CLK(n2924), 
        .Q(g1531), .QN(n1652) );
  SDFFX1 DFF_165_Q_reg ( .D(g6180), .SI(g1531), .SE(n2841), .CLK(n2888), .Q(
        g1458), .QN(n1703) );
  SDFFX1 DFF_166_Q_reg ( .D(g10718), .SI(g1458), .SE(n2799), .CLK(n2909), .Q(
        g572) );
  SDFFX1 DFF_167_Q_reg ( .D(g6912), .SI(g572), .SE(n2815), .CLK(n2901), .Q(
        g1011), .QN(n2658) );
  SDFFX1 DFF_168_Q_reg ( .D(g10719), .SI(g1011), .SE(n2815), .CLK(n2901), .Q(
        n3051) );
  SDFFX1 DFF_169_Q_reg ( .D(g6234), .SI(n3051), .SE(n2815), .CLK(n2901), .Q(
        g1411), .QN(n2550) );
  SDFFX1 DFF_170_Q_reg ( .D(g6099), .SI(g1411), .SE(n2763), .CLK(n2927), .Q(
        g1074) );
  SDFFX1 DFF_171_Q_reg ( .D(g11259), .SI(g1074), .SE(n2828), .CLK(n2894), .Q(
        g444), .QN(n2640) );
  SDFFX1 DFF_172_Q_reg ( .D(g8039), .SI(g444), .SE(n2809), .CLK(n2904), .Q(
        g1474) );
  SDFFX1 DFF_173_Q_reg ( .D(g6059), .SI(g1474), .SE(n2772), .CLK(n2922), .Q(
        g1080) );
  SDFFX1 DFF_174_Q_reg ( .D(g5396), .SI(g1080), .SE(n2795), .CLK(n2911), .Q(
        g1713), .QN(n1610) );
  SDFFX1 DFF_175_Q_reg ( .D(g262), .SI(g1713), .SE(n2779), .CLK(n2919), .Q(
        g333), .QN(n2685) );
  SDFFX1 DFF_176_Q_reg ( .D(g6906), .SI(g333), .SE(n2779), .CLK(n2919), .Q(
        g269), .QN(n2563) );
  SDFFX1 DFF_177_Q_reg ( .D(g11266), .SI(g269), .SE(n2830), .CLK(n2894), .Q(
        g401), .QN(n2665) );
  SDFFX1 DFF_178_Q_reg ( .D(g11294), .SI(g401), .SE(n2818), .CLK(n2900), .Q(
        g1857), .QN(n1682) );
  SDFFX1 DFF_179_Q_reg ( .D(g5421), .SI(g1857), .SE(n2817), .CLK(n2900), .Q(g9), .QN(n2623) );
  SDFFX1 DFF_180_Q_reg ( .D(g8649), .SI(g9), .SE(n2817), .CLK(n2900), .Q(g664), 
        .QN(n2621) );
  SDFFX1 DFF_181_Q_reg ( .D(g11312), .SI(g664), .SE(n2802), .CLK(n2908), .Q(
        g965) );
  SDFFX1 DFF_182_Q_reg ( .D(g6840), .SI(g965), .SE(n2802), .CLK(n2908), .Q(
        g1400), .QN(n1629) );
  SDFFX1 DFF_183_Q_reg ( .D(g254), .SI(g1400), .SE(n2788), .CLK(n2914), .Q(
        g309), .QN(n2458) );
  SDFFX1 DFF_184_Q_reg ( .D(g7202), .SI(g309), .SE(n2803), .CLK(n2907), .Q(
        g814), .QN(n2738) );
  SDFFX1 DFF_185_Q_reg ( .D(g6834), .SI(g814), .SE(n2784), .CLK(n2916), .Q(
        g231), .QN(n2677) );
  SDFFX1 DFF_186_Q_reg ( .D(g10795), .SI(g231), .SE(n2777), .CLK(n2920), .Q(
        g557) );
  SDFFX1 DFF_187_Q_reg ( .D(g103), .SI(g557), .SE(n2777), .CLK(n2920), .Q(
        g2612) );
  SDFFX1 DFF_188_Q_reg ( .D(g875), .SI(g2612), .SE(n2778), .CLK(n2920), .Q(
        g869), .QN(n2504) );
  SDFFX1 DFF_189_Q_reg ( .D(g6831), .SI(g869), .SE(n2778), .CLK(n2920), .Q(
        g1383), .QN(n2510) );
  SDFFX1 DFF_190_Q_reg ( .D(g8060), .SI(g1383), .SE(n2808), .CLK(n2904), .Q(
        g158), .QN(n2650) );
  SDFFX1 DFF_191_Q_reg ( .D(g4893), .SI(g158), .SE(n2819), .CLK(n2899), .Q(
        g627), .QN(n1701) );
  SDFFX1 DFF_192_Q_reg ( .D(g7244), .SI(g627), .SE(n2832), .CLK(n2892), .Q(
        g1023), .QN(n2593) );
  SDFFX1 DFF_193_Q_reg ( .D(g6026), .SI(g1023), .SE(n2832), .CLK(n2892), .Q(
        g259) );
  SDFFX1 DFF_194_Q_reg ( .D(g3069), .SI(g259), .SE(n2804), .CLK(n2906), .Q(
        n3050), .QN(n4935) );
  SDFFX1 DFF_195_Q_reg ( .D(g11608), .SI(n3050), .SE(n2791), .CLK(n2913), .Q(
        g1327) );
  SDFFX1 DFF_196_Q_reg ( .D(g7660), .SI(g1327), .SE(n2820), .CLK(n2898), .Q(
        g654), .QN(n2729) );
  SDFFX1 DFF_197_Q_reg ( .D(g6911), .SI(g654), .SE(n2805), .CLK(n2906), .Q(
        g293) );
  SDFFX1 DFF_198_Q_reg ( .D(g11640), .SI(g293), .SE(n2805), .CLK(n2906), .Q(
        g1346), .QN(n2706) );
  SDFFX1 DFF_199_Q_reg ( .D(g8777), .SI(g1346), .SE(n2784), .CLK(n2916), .Q(
        g1633) );
  SDFFX1 DFF_200_Q_reg ( .D(g4274), .SI(g1633), .SE(n2784), .CLK(n2917), .Q(
        g1753), .QN(n2716) );
  SDFFX1 DFF_201_Q_reg ( .D(n2750), .SI(g1753), .SE(n2784), .CLK(n2917), .Q(
        g1508) );
  SDFFX1 DFF_202_Q_reg ( .D(g7297), .SI(g1508), .SE(n2761), .CLK(n2928), .Q(
        g1240), .QN(n2699) );
  SDFFX1 DFF_203_Q_reg ( .D(g11326), .SI(g1240), .SE(n2825), .CLK(n2896), .Q(
        g538) );
  SDFFX1 DFF_204_Q_reg ( .D(g11269), .SI(g538), .SE(n2829), .CLK(n2894), .Q(
        g416), .QN(n2638) );
  SDFFX1 DFF_205_Q_reg ( .D(g11325), .SI(g416), .SE(n2825), .CLK(n2896), .Q(
        g542), .QN(n2693) );
  SDFFX1 DFF_206_Q_reg ( .D(g10864), .SI(g542), .SE(n2794), .CLK(n2911), .Q(
        g1681) );
  SDFFX1 DFF_207_Q_reg ( .D(g11290), .SI(g1681), .SE(n2776), .CLK(n2921), .Q(
        g374), .QN(n2617) );
  SDFFX1 DFF_208_Q_reg ( .D(g10798), .SI(g374), .SE(n2776), .CLK(n2921), .Q(
        g563) );
  SDFFX1 DFF_209_Q_reg ( .D(g8284), .SI(g563), .SE(n2828), .CLK(n2895), .Q(
        g1914) );
  SDFFX1 DFF_210_Q_reg ( .D(g11328), .SI(g1914), .SE(n2824), .CLK(n2896), .Q(
        g530), .QN(n2690) );
  SDFFX1 DFF_211_Q_reg ( .D(g10800), .SI(g530), .SE(n2789), .CLK(n2914), .Q(
        g575) );
  SDFFX1 DFF_212_Q_reg ( .D(g8944), .SI(g575), .SE(n2761), .CLK(n2928), .Q(
        g1936) );
  SDFFX1 DFF_213_Q_reg ( .D(g7183), .SI(g1936), .SE(n2761), .CLK(n2928), .Q(
        g8978), .QN(n1674) );
  SDFFX1 DFF_214_Q_reg ( .D(g4465), .SI(g8978), .SE(n2761), .CLK(n2928), .Q(
        test_so4), .QN(n2755) );
  SDFFX1 DFF_215_Q_reg ( .D(g1356), .SI(test_si5), .SE(n2764), .CLK(n2926), 
        .Q(g1317) );
  SDFFX1 DFF_216_Q_reg ( .D(g11484), .SI(g1317), .SE(n2832), .CLK(n2893), .Q(
        g357) );
  SDFFX1 DFF_217_Q_reg ( .D(g11263), .SI(g357), .SE(n2830), .CLK(n2893), .Q(
        g386), .QN(n2663) );
  SDFFX1 DFF_218_Q_reg ( .D(g6501), .SI(g386), .SE(n2779), .CLK(n2919), .Q(
        g1601) );
  SDFFX1 DFF_220_Q_reg ( .D(g6757), .SI(g1601), .SE(n2779), .CLK(n2919), .Q(
        g166), .QN(n2648) );
  SDFFX1 DFF_221_Q_reg ( .D(g11334), .SI(g166), .SE(n2779), .CLK(n2919), .Q(
        g501), .QN(n1690) );
  SDFFX1 DFF_222_Q_reg ( .D(g6042), .SI(g501), .SE(n2779), .CLK(n2919), .Q(
        g262) );
  SDFFX1 DFF_223_Q_reg ( .D(g8384), .SI(g262), .SE(n2774), .CLK(n2921), .Q(
        g1840), .QN(n2695) );
  SDFFX1 DFF_224_Q_reg ( .D(g6653), .SI(g1840), .SE(n2774), .CLK(n2921), .Q(
        g8983), .QN(n1666) );
  SDFFX1 DFF_225_Q_reg ( .D(g257), .SI(g8983), .SE(n2774), .CLK(n2921), .Q(
        g318), .QN(n2662) );
  SDFFX1 DFF_226_Q_reg ( .D(g5763), .SI(g318), .SE(n2804), .CLK(n2907), .Q(
        g1356) );
  SDFFX1 DFF_227_Q_reg ( .D(g5849), .SI(g1356), .SE(n2804), .CLK(n2907), .Q(
        g794), .QN(n2632) );
  SDFFX1 DFF_228_Q_reg ( .D(g10722), .SI(g794), .SE(n2803), .CLK(n2907), .Q(
        n3048), .QN(DFF_228_n1) );
  SDFFX1 DFF_229_Q_reg ( .D(g6929), .SI(n3048), .SE(n2763), .CLK(n2927), .Q(
        g302) );
  SDFFX1 DFF_230_Q_reg ( .D(g11488), .SI(g302), .SE(n2763), .CLK(n2927), .Q(
        g342) );
  SDFFX1 DFF_231_Q_reg ( .D(g7299), .SI(g342), .SE(n2823), .CLK(n2897), .Q(
        g1250) );
  SDFFX1 DFF_232_Q_reg ( .D(g4330), .SI(g1250), .SE(n2823), .CLK(n2897), .Q(
        g1163) );
  SDFFX1 DFF_233_Q_reg ( .D(g1958), .SI(g1163), .SE(n2810), .CLK(n2903), .Q(
        n3047), .QN(g5816) );
  SDFFX1 DFF_234_Q_reg ( .D(g7257), .SI(n3047), .SE(n2837), .CLK(n2890), .Q(
        g1032) );
  SDFFX1 DFF_235_Q_reg ( .D(g8775), .SI(g1032), .SE(n2783), .CLK(n2917), .Q(
        g1432), .QN(n2654) );
  SDFFX1 DFF_237_Q_reg ( .D(g5770), .SI(g1432), .SE(n2842), .CLK(n2888), .Q(
        g1453), .QN(n1628) );
  SDFFX1 DFF_238_Q_reg ( .D(g11486), .SI(g1453), .SE(n2813), .CLK(n2902), .Q(
        g363) );
  SDFFX1 DFF_239_Q_reg ( .D(g261), .SI(g363), .SE(n2813), .CLK(n2902), .Q(g330), .QN(n2457) );
  SDFFX1 DFF_240_Q_reg ( .D(g4338), .SI(g330), .SE(n2813), .CLK(n2902), .Q(
        g1157) );
  SDFFX1 DFF_241_Q_reg ( .D(g4500), .SI(g1157), .SE(n2813), .CLK(n2902), .Q(
        n3046), .QN(n4951) );
  SDFFX1 DFF_242_Q_reg ( .D(g10721), .SI(n3046), .SE(n2813), .CLK(n2902), .Q(
        n3045), .QN(DFF_242_n1) );
  SDFFX1 DFF_243_Q_reg ( .D(g8147), .SI(n3045), .SE(n2812), .CLK(n2902), .Q(
        g928), .QN(n1604) );
  SDFFX1 DFF_244_Q_reg ( .D(g6038), .SI(g928), .SE(n2789), .CLK(n2914), .Q(
        g261) );
  SDFFX1 DFF_245_Q_reg ( .D(g11337), .SI(g261), .SE(n2825), .CLK(n2896), .Q(
        g516), .QN(n1620) );
  SDFFX1 DFF_246_Q_reg ( .D(g6045), .SI(g516), .SE(n2788), .CLK(n2914), .Q(
        g254) );
  SDFFX1 DFF_247_Q_reg ( .D(g7191), .SI(g254), .SE(n2788), .CLK(n2914), .Q(
        g4178), .QN(n2523) );
  SDFFX1 DFF_248_Q_reg ( .D(g826), .SI(g4178), .SE(n2770), .CLK(n2924), .Q(
        g861), .QN(n2462) );
  SDFFX1 DFF_249_Q_reg ( .D(g8774), .SI(g861), .SE(n2770), .CLK(n2924), .Q(
        g1627), .QN(n2582) );
  SDFFX1 DFF_250_Q_reg ( .D(g7293), .SI(g1627), .SE(n2821), .CLK(n2898), .Q(
        g1292) );
  SDFFX1 DFF_251_Q_reg ( .D(g6907), .SI(g1292), .SE(n2765), .CLK(n2926), .Q(
        g290) );
  SDFFX1 DFF_252_Q_reg ( .D(g4903), .SI(g290), .SE(n2839), .CLK(n2889), .Q(
        n3044) );
  SDFFX1 DFF_253_Q_reg ( .D(g6123), .SI(n3044), .SE(n2833), .CLK(n2892), .Q(
        g4176), .QN(n2522) );
  SDFFX1 DFF_254_Q_reg ( .D(g6506), .SI(g4176), .SE(n2814), .CLK(n2902), .Q(
        g1583) );
  SDFFX1 DFF_255_Q_reg ( .D(g11376), .SI(g1583), .SE(n2813), .CLK(n2902), .Q(
        g466), .QN(n1646) );
  SDFFX1 DFF_256_Q_reg ( .D(g6542), .SI(g466), .SE(n2841), .CLK(n2888), .Q(
        g1561) );
  SDFFX1 DFF_258_Q_reg ( .D(g6551), .SI(g1561), .SE(n2809), .CLK(n2904), .Q(
        g1546) );
  SDFFX1 DFF_259_Q_reg ( .D(g6901), .SI(g1546), .SE(n2809), .CLK(n2904), .Q(
        g287) );
  SDFFX1 DFF_260_Q_reg ( .D(g10797), .SI(g287), .SE(n2808), .CLK(n2904), .Q(
        g560) );
  SDFFX1 DFF_261_Q_reg ( .D(g8505), .SI(g560), .SE(n2811), .CLK(n2903), .Q(
        g617), .QN(n1645) );
  SDFFX1 DFF_262_Q_reg ( .D(n2751), .SI(g617), .SE(n2811), .CLK(n2903), .Q(
        n1631), .QN(n4938) );
  SDFFX1 DFF_263_Q_reg ( .D(g11647), .SI(n1631), .SE(n2845), .CLK(n2886), .Q(
        g336) );
  SDFFX1 DFF_264_Q_reg ( .D(g11340), .SI(g336), .SE(n2773), .CLK(n2922), .Q(
        g456), .QN(n1641) );
  SDFFX1 DFF_265_Q_reg ( .D(g253), .SI(g456), .SE(n2773), .CLK(n2922), .Q(g305), .QN(n1681) );
  SDFFX1 DFF_266_Q_reg ( .D(g11625), .SI(g305), .SE(n2837), .CLK(n2890), .Q(
        g345) );
  SDFFX1 DFF_267_Q_reg ( .D(g636), .SI(g345), .SE(n2842), .CLK(n2887), .Q(g8)
         );
  SDFFX1 DFF_268_Q_reg ( .D(g6502), .SI(g8), .SE(n2792), .CLK(n2912), .Q(
        test_so5) );
  SDFFX1 DFF_269_Q_reg ( .D(N599), .SI(test_si6), .SE(n2833), .CLK(n2892), .Q(
        g2648), .QN(n4936) );
  SDFFX1 DFF_270_Q_reg ( .D(g6049), .SI(g2648), .SE(n2833), .CLK(n2892), .Q(
        g255) );
  SDFFX1 DFF_271_Q_reg ( .D(g8945), .SI(g255), .SE(n2827), .CLK(n2895), .Q(
        g1945), .QN(n1697) );
  SDFFX1 DFF_272_Q_reg ( .D(g4231), .SI(g1945), .SE(n2796), .CLK(n2910), .Q(
        g1738), .QN(n1640) );
  SDFFX1 DFF_273_Q_reg ( .D(g8040), .SI(g1738), .SE(n2809), .CLK(n2904), .Q(
        g1478), .QN(n2725) );
  SDFFX1 DFF_275_Q_reg ( .D(n356), .SI(g1478), .SE(n2809), .CLK(n2904), .Q(
        n3042), .QN(DFF_275_n1) );
  SDFFX1 DFF_276_Q_reg ( .D(g6155), .SI(n3042), .SE(n2773), .CLK(n2922), .Q(
        g1690), .QN(n1653) );
  SDFFX1 DFF_277_Q_reg ( .D(g8043), .SI(g1690), .SE(n2835), .CLK(n2891), .Q(
        g1482), .QN(n2652) );
  SDFFX1 DFF_278_Q_reg ( .D(g5173), .SI(g1482), .SE(n2793), .CLK(n2912), .Q(
        g1110), .QN(n1677) );
  SDFFX1 DFF_279_Q_reg ( .D(g6916), .SI(g1110), .SE(n2764), .CLK(n2926), .Q(
        g296) );
  SDFFX1 DFF_280_Q_reg ( .D(g10861), .SI(g296), .SE(n2812), .CLK(n2902), .Q(
        g1663) );
  SDFFX1 DFF_281_Q_reg ( .D(g8431), .SI(g1663), .SE(n2812), .CLK(n2902), .Q(
        g700), .QN(n2680) );
  SDFFX1 DFF_282_Q_reg ( .D(g4309), .SI(g700), .SE(n2771), .CLK(n2923), .Q(
        g1762), .QN(n2715) );
  SDFFX1 DFF_283_Q_reg ( .D(g11485), .SI(g1762), .SE(n2815), .CLK(n2901), .Q(
        g360) );
  SDFFX1 DFF_284_Q_reg ( .D(g6334), .SI(g360), .SE(n2806), .CLK(n2906), .Q(
        g192) );
  SDFFX1 DFF_285_Q_reg ( .D(g10767), .SI(g192), .SE(n2843), .CLK(n2887), .Q(
        g1657) );
  SDFFX1 DFF_286_Q_reg ( .D(g8923), .SI(g1657), .SE(n2843), .CLK(n2887), .Q(
        g722), .QN(n1693) );
  SDFFX1 DFF_287_Q_reg ( .D(g7189), .SI(g722), .SE(n2775), .CLK(n2921), .Q(
        g8980), .QN(n1673) );
  SDFFX1 DFF_288_Q_reg ( .D(g10799), .SI(g8980), .SE(n2837), .CLK(n2890), .Q(
        g566) );
  SDFFX1 DFF_289_Q_reg ( .D(g6747), .SI(g566), .SE(n2844), .CLK(n2887), .Q(
        n3041), .QN(n4948) );
  SDFFX1 DFF_290_Q_reg ( .D(g6080), .SI(n3041), .SE(n2831), .CLK(n2893), .Q(
        g1089) );
  SDFFX1 DFF_291_Q_reg ( .D(g3381), .SI(g1089), .SE(n2831), .CLK(n2893), .Q(
        g2986), .QN(n2481) );
  SDFFX1 DFF_292_Q_reg ( .D(g5910), .SI(g2986), .SE(n2832), .CLK(n2892), .Q(
        g1071) );
  SDFFX1 DFF_293_Q_reg ( .D(g11393), .SI(g1071), .SE(n2834), .CLK(n2891), .Q(
        g986), .QN(n1722) );
  SDFFX1 DFF_294_Q_reg ( .D(g11349), .SI(g986), .SE(n2834), .CLK(n2891), .Q(
        g971), .QN(n2709) );
  SDFFX1 DFF_295_Q_reg ( .D(g83), .SI(g971), .SE(n2834), .CLK(n2892), .Q(g1955) );
  SDFFX1 DFF_296_Q_reg ( .D(g6439), .SI(g1955), .SE(n2819), .CLK(n2899), .Q(
        g143), .QN(n2671) );
  SDFFX1 DFF_297_Q_reg ( .D(g9266), .SI(g143), .SE(n2818), .CLK(n2899), .Q(
        g1814), .QN(n1608) );
  SDFFX1 DFF_299_Q_reg ( .D(g1217), .SI(g1814), .SE(n2818), .CLK(n2899), .Q(
        g1212), .QN(n2743) );
  SDFFX1 DFF_300_Q_reg ( .D(g8940), .SI(g1212), .SE(n2827), .CLK(n2895), .Q(
        g1918), .QN(n2681) );
  SDFFX1 DFF_301_Q_reg ( .D(g7705), .SI(g1918), .SE(n2788), .CLK(n2915), .Q(
        g4179) );
  SDFFX1 DFF_302_Q_reg ( .D(g9269), .SI(g4179), .SE(n2818), .CLK(n2900), .Q(
        g1822), .QN(n1643) );
  SDFFX1 DFF_303_Q_reg ( .D(g6820), .SI(g1822), .SE(n2789), .CLK(n2914), .Q(
        g237), .QN(n2678) );
  SDFFX1 DFF_304_Q_reg ( .D(g756), .SI(g237), .SE(n2786), .CLK(n2916), .Q(g746), .QN(n2731) );
  SDFFX1 DFF_306_Q_reg ( .D(g8042), .SI(g746), .SE(n2772), .CLK(n2922), .Q(
        g1462) );
  SDFFX1 DFF_307_Q_reg ( .D(g6759), .SI(g1462), .SE(n2772), .CLK(n2922), .Q(
        g178) );
  SDFFX1 DFF_308_Q_reg ( .D(g11487), .SI(g178), .SE(n2772), .CLK(n2923), .Q(
        g366) );
  SDFFX1 DFF_309_Q_reg ( .D(g802), .SI(g366), .SE(n2803), .CLK(n2907), .Q(g837), .QN(n2461) );
  SDFFX1 DFF_310_Q_reg ( .D(g9124), .SI(g837), .SE(n2843), .CLK(n2887), .Q(
        g599), .QN(n1644) );
  SDFFX1 DFF_311_Q_reg ( .D(g11293), .SI(g599), .SE(n2845), .CLK(n2886), .Q(
        g1854) );
  SDFFX1 DFF_312_Q_reg ( .D(g11298), .SI(g1854), .SE(n2845), .CLK(n2886), .Q(
        g944), .QN(n2469) );
  SDFFX1 DFF_313_Q_reg ( .D(g8287), .SI(g944), .SE(n2773), .CLK(n2922), .Q(
        g1941), .QN(n2626) );
  SDFFX1 DFF_314_Q_reg ( .D(g8047), .SI(g1941), .SE(n2837), .CLK(n2890), .Q(
        g170), .QN(n2742) );
  SDFFX1 DFF_315_Q_reg ( .D(g6205), .SI(g170), .SE(n2785), .CLK(n2916), .Q(
        g1520), .QN(n1710) );
  SDFFX1 DFF_316_Q_reg ( .D(g8885), .SI(g1520), .SE(n2811), .CLK(n2903), .Q(
        g686), .QN(n1676) );
  SDFFX1 DFF_317_Q_reg ( .D(g11305), .SI(g686), .SE(n2811), .CLK(n2903), .Q(
        g953), .QN(n2468) );
  SDFFX1 DFF_318_Q_reg ( .D(g5556), .SI(g953), .SE(n2810), .CLK(n2903), .Q(
        g1958) );
  SDFFX1 DFF_319_Q_reg ( .D(g10664), .SI(g1958), .SE(n2810), .CLK(n2903), .Q(
        n3040) );
  SDFFX1 DFF_320_Q_reg ( .D(g2478), .SI(n3040), .SE(n2810), .CLK(n2904), .Q(
        g1765) );
  SDFFX1 DFF_321_Q_reg ( .D(g10711), .SI(g1765), .SE(n2798), .CLK(n2909), .Q(
        g1733), .QN(n2485) );
  SDFFX1 DFF_322_Q_reg ( .D(g7303), .SI(g1733), .SE(n2822), .CLK(n2898), .Q(
        test_so6) );
  SDFFX1 DFF_323_Q_reg ( .D(g5194), .SI(test_si7), .SE(n2799), .CLK(n2909), 
        .Q(g1610) );
  SDFFX1 DFF_324_Q_reg ( .D(g7541), .SI(g1610), .SE(n2791), .CLK(n2913), .Q(
        g1796), .QN(n1626) );
  SDFFX1 DFF_325_Q_reg ( .D(g11607), .SI(g1796), .SE(n2791), .CLK(n2913), .Q(
        g1324), .QN(n2472) );
  SDFFX1 DFF_326_Q_reg ( .D(g6541), .SI(g1324), .SE(n2836), .CLK(n2891), .Q(
        g1540) );
  SDFFX1 DFF_327_Q_reg ( .D(g6827), .SI(g1540), .SE(n2835), .CLK(n2891), .Q(
        n3038), .QN(n4943) );
  SDFFX1 DFF_328_Q_reg ( .D(n2752), .SI(n3038), .SE(n2804), .CLK(n2906), .Q(
        g3069), .QN(n2482) );
  SDFFX1 DFF_329_Q_reg ( .D(g11332), .SI(g3069), .SE(n2838), .CLK(n2890), .Q(
        g491), .QN(n1691) );
  SDFFX1 DFF_330_Q_reg ( .D(g4902), .SI(g491), .SE(n2840), .CLK(n2889), .Q(
        n3037), .QN(DFF_330_n1) );
  SDFFX1 DFF_331_Q_reg ( .D(g6828), .SI(n3037), .SE(n2835), .CLK(n2891), .Q(
        g213), .QN(n2513) );
  SDFFX1 DFF_332_Q_reg ( .D(g6516), .SI(g213), .SE(n2792), .CLK(n2913), .Q(
        g1781), .QN(n1659) );
  SDFFX1 DFF_333_Q_reg ( .D(g8938), .SI(g1781), .SE(n2823), .CLK(n2897), .Q(
        g1900), .QN(n1675) );
  SDFFX1 DFF_334_Q_reg ( .D(g7298), .SI(g1900), .SE(n2823), .CLK(n2897), .Q(
        g1245) );
  SDFFX1 DFF_335_Q_reg ( .D(n3), .SI(g1245), .SE(n2823), .CLK(n2897), .Q(n3036), .QN(n4949) );
  SDFFX1 DFF_336_Q_reg ( .D(g6672), .SI(n3036), .SE(n2819), .CLK(n2899), .Q(
        n3035), .QN(DFF_336_n1) );
  SDFFX1 DFF_337_Q_reg ( .D(g8048), .SI(n3035), .SE(n2819), .CLK(n2899), .Q(
        g148), .QN(n2672) );
  SDFFX1 DFF_338_Q_reg ( .D(g798), .SI(g148), .SE(n2781), .CLK(n2918), .Q(g833), .QN(n2460) );
  SDFFX1 DFF_339_Q_reg ( .D(g8285), .SI(g833), .SE(n2774), .CLK(n2922), .Q(
        g1923), .QN(n1718) );
  SDFFX1 DFF_340_Q_reg ( .D(g8254), .SI(g1923), .SE(n2774), .CLK(n2922), .Q(
        g936), .QN(n1630) );
  SDFFX1 DFF_342_Q_reg ( .D(g11604), .SI(g936), .SE(n2796), .CLK(n2911), .Q(
        g1314) );
  SDFFX1 DFF_343_Q_reg ( .D(g814), .SI(g1314), .SE(n2796), .CLK(n2911), .Q(
        g849), .QN(n2490) );
  SDFFX1 DFF_344_Q_reg ( .D(g11636), .SI(g849), .SE(n2795), .CLK(n2911), .Q(
        g1336), .QN(n2707) );
  SDFFX1 DFF_345_Q_reg ( .D(g6910), .SI(g1336), .SE(n2772), .CLK(n2923), .Q(
        g272), .QN(n2557) );
  SDFFX1 DFF_346_Q_reg ( .D(g8173), .SI(g272), .SE(n2771), .CLK(n2923), .Q(
        g1806), .QN(n2734) );
  SDFFX1 DFF_347_Q_reg ( .D(g8245), .SI(g1806), .SE(n2770), .CLK(n2923), .Q(
        g826), .QN(n1716) );
  SDFFX1 DFF_349_Q_reg ( .D(g8281), .SI(g826), .SE(n2766), .CLK(n2926), .Q(
        g1887) );
  SDFFX1 DFF_350_Q_reg ( .D(n36), .SI(g1887), .SE(n2765), .CLK(n2926), .Q(
        n3034) );
  SDFFX1 DFF_351_Q_reg ( .D(g11314), .SI(n3034), .SE(n2765), .CLK(n2926), .Q(
        g968) );
  SDFFX1 DFF_352_Q_reg ( .D(g4905), .SI(g968), .SE(n2839), .CLK(n2889), .Q(
        n3033), .QN(n4946) );
  SDFFX1 DFF_353_Q_reg ( .D(g4484), .SI(n3033), .SE(n2839), .CLK(n2889), .Q(
        g1137), .QN(n1597) );
  SDFFX1 DFF_354_Q_reg ( .D(g8937), .SI(g1137), .SE(n2827), .CLK(n2895), .Q(
        g1891), .QN(n1657) );
  SDFFX1 DFF_355_Q_reg ( .D(g7300), .SI(g1891), .SE(n2823), .CLK(n2897), .Q(
        g1255), .QN(n2629) );
  SDFFX1 DFF_356_Q_reg ( .D(g6002), .SI(g1255), .SE(n2776), .CLK(n2920), .Q(
        g257) );
  SDFFX1 DFF_357_Q_reg ( .D(n1588), .SI(g257), .SE(n2776), .CLK(n2920), .Q(
        g874) );
  SDFFX1 DFF_358_Q_reg ( .D(g9110), .SI(g874), .SE(n2768), .CLK(n2925), .Q(
        g591), .QN(n1607) );
  SDFFX1 DFF_359_Q_reg ( .D(g8926), .SI(g591), .SE(n2843), .CLK(n2887), .Q(
        g731), .QN(n1696) );
  SDFFX1 DFF_360_Q_reg ( .D(g8631), .SI(g731), .SE(n2842), .CLK(n2887), .Q(
        g636) );
  SDFFX1 DFF_361_Q_reg ( .D(g7632), .SI(g636), .SE(n2846), .CLK(n2886), .Q(
        g1218), .QN(n2508) );
  SDFFX1 DFF_362_Q_reg ( .D(g9150), .SI(g1218), .SE(n2768), .CLK(n2924), .Q(
        g605), .QN(n1593) );
  SDFFX1 DFF_363_Q_reg ( .D(g6531), .SI(g605), .SE(n2768), .CLK(n2924), .Q(
        g8986), .QN(n1665) );
  SDFFX1 DFF_364_Q_reg ( .D(g6786), .SI(g8986), .SE(n2768), .CLK(n2924), .Q(
        g182) );
  SDFFX1 DFF_365_Q_reg ( .D(g11303), .SI(g182), .SE(n2802), .CLK(n2907), .Q(
        g950), .QN(n2470) );
  SDFFX1 DFF_366_Q_reg ( .D(g4477), .SI(g950), .SE(n2802), .CLK(n2907), .Q(
        g1129), .QN(n1705) );
  SDFFX1 DFF_367_Q_reg ( .D(g822), .SI(g1129), .SE(n2802), .CLK(n2907), .Q(
        g857) );
  SDFFX1 DFF_368_Q_reg ( .D(g11258), .SI(g857), .SE(n2829), .CLK(n2894), .Q(
        g448), .QN(n2641) );
  SDFFX1 DFF_369_Q_reg ( .D(g9272), .SI(g448), .SE(n2818), .CLK(n2900), .Q(
        g1828), .QN(n1605) );
  SDFFX1 DFF_370_Q_reg ( .D(g10773), .SI(g1828), .SE(n2765), .CLK(n2926), .Q(
        g1727), .QN(n2486) );
  SDFFX1 DFF_371_Q_reg ( .D(g6470), .SI(g1727), .SE(n2800), .CLK(n2909), .Q(
        g1592), .QN(n2538) );
  SDFFX1 DFF_372_Q_reg ( .D(g5083), .SI(g1592), .SE(n2800), .CLK(n2909), .Q(
        g1703), .QN(n2745) );
  SDFFX1 DFF_373_Q_reg ( .D(g8286), .SI(g1703), .SE(n2774), .CLK(n2922), .Q(
        g1932) );
  SDFFX1 DFF_374_Q_reg ( .D(g8773), .SI(g1932), .SE(n2835), .CLK(n2891), .Q(
        g1624) );
  SDFFX1 DFF_376_Q_reg ( .D(g6054), .SI(g1624), .SE(n2845), .CLK(n2886), .Q(
        test_so7) );
  SDFFX1 DFF_377_Q_reg ( .D(g101), .SI(test_si8), .SE(n2846), .CLK(n2886), .Q(
        g2601) );
  SDFFX1 DFF_378_Q_reg ( .D(g11260), .SI(g2601), .SE(n2828), .CLK(n2894), .Q(
        g440), .QN(n2639) );
  SDFFX1 DFF_379_Q_reg ( .D(g11338), .SI(g440), .SE(n2825), .CLK(n2896), .Q(
        g476), .QN(n1599) );
  SDFFX1 DFF_380_Q_reg ( .D(g5918), .SI(g476), .SE(n2825), .CLK(n2896), .Q(
        g119), .QN(n1613) );
  SDFFX1 DFF_381_Q_reg ( .D(g8922), .SI(g119), .SE(n2817), .CLK(n2900), .Q(
        g668), .QN(n1662) );
  SDFFX1 DFF_382_Q_reg ( .D(g8049), .SI(g668), .SE(n2805), .CLK(n2906), .Q(
        g139), .QN(n2645) );
  SDFFX1 DFF_383_Q_reg ( .D(g4342), .SI(g139), .SE(n2805), .CLK(n2906), .Q(
        g1149), .QN(n1685) );
  SDFFX1 DFF_384_Q_reg ( .D(g10720), .SI(g1149), .SE(n2805), .CLK(n2906), .Q(
        n3031) );
  SDFFX1 DFF_385_Q_reg ( .D(g6755), .SI(n3031), .SE(n2840), .CLK(n2889), .Q(
        n3030), .QN(DFF_385_n1) );
  SDFFX1 DFF_386_Q_reg ( .D(g6897), .SI(n3030), .SE(n2768), .CLK(n2925), .Q(
        g263) );
  SDFFX1 DFF_387_Q_reg ( .D(g7709), .SI(g263), .SE(n2803), .CLK(n2907), .Q(
        g818), .QN(n2739) );
  SDFFX1 DFF_388_Q_reg ( .D(g4255), .SI(g818), .SE(n2803), .CLK(n2907), .Q(
        g1747), .QN(n2714) );
  SDFFX1 DFF_389_Q_reg ( .D(g5543), .SI(g1747), .SE(n2803), .CLK(n2907), .Q(
        g802), .QN(n1622) );
  SDFFX1 DFF_390_Q_reg ( .D(g6915), .SI(g802), .SE(n2808), .CLK(n2905), .Q(
        g275) );
  SDFFX1 DFF_391_Q_reg ( .D(g6513), .SI(g275), .SE(n2808), .CLK(n2905), .Q(
        g1524), .QN(n1649) );
  SDFFX1 DFF_392_Q_reg ( .D(g6480), .SI(g1524), .SE(n2808), .CLK(n2905), .Q(
        g1577), .QN(n2537) );
  SDFFX1 DFF_393_Q_reg ( .D(g6733), .SI(g1577), .SE(n2807), .CLK(n2905), .Q(
        g810), .QN(n2737) );
  SDFFX1 DFF_394_Q_reg ( .D(g11264), .SI(g810), .SE(n2830), .CLK(n2894), .Q(
        g391), .QN(n2703) );
  SDFFX1 DFF_395_Q_reg ( .D(g8973), .SI(g391), .SE(n2817), .CLK(n2900), .Q(
        g658), .QN(n1615) );
  SDFFX1 DFF_396_Q_reg ( .D(g6833), .SI(g658), .SE(n2777), .CLK(n2920), .Q(
        g1386), .QN(n2668) );
  SDFFX1 DFF_397_Q_reg ( .D(g5996), .SI(g1386), .SE(n2778), .CLK(n2919), .Q(
        g253) );
  SDFFX1 DFF_398_Q_reg ( .D(n1587), .SI(g253), .SE(n2778), .CLK(n2920), .Q(
        g875) );
  SDFFX1 DFF_399_Q_reg ( .D(g4473), .SI(g875), .SE(n2776), .CLK(n2921), .Q(
        g1125), .QN(n1708) );
  SDFFX1 DFF_400_Q_reg ( .D(g5755), .SI(g1125), .SE(n2764), .CLK(n2926), .Q(
        g201), .QN(n1619) );
  SDFFX1 DFF_401_Q_reg ( .D(g7295), .SI(g201), .SE(n2821), .CLK(n2898), .Q(
        g1280), .QN(n1862) );
  SDFFX1 DFF_402_Q_reg ( .D(g6068), .SI(g1280), .SE(n2820), .CLK(n2898), .Q(
        g1083) );
  SDFFX1 DFF_403_Q_reg ( .D(g7137), .SI(g1083), .SE(n2820), .CLK(n2898), .Q(
        g650), .QN(n1709) );
  SDFFX1 DFF_404_Q_reg ( .D(g8779), .SI(g650), .SE(n2789), .CLK(n2914), .Q(
        g1636) );
  SDFFX1 DFF_405_Q_reg ( .D(g818), .SI(g1636), .SE(n2789), .CLK(n2914), .Q(
        g853), .QN(n2465) );
  SDFFX1 DFF_406_Q_reg ( .D(g11270), .SI(g853), .SE(n2829), .CLK(n2894), .Q(
        g421), .QN(n2684) );
  SDFFX1 DFF_407_Q_reg ( .D(g5529), .SI(g421), .SE(n2838), .CLK(n2889), .Q(
        g4174), .QN(n2520) );
  SDFFX1 DFF_408_Q_reg ( .D(g11306), .SI(g4174), .SE(n2807), .CLK(n2905), .Q(
        g956) );
  SDFFX1 DFF_409_Q_reg ( .D(g11291), .SI(g956), .SE(n2807), .CLK(n2905), .Q(
        g378), .QN(n2615) );
  SDFFX1 DFF_410_Q_reg ( .D(g4283), .SI(g378), .SE(n2764), .CLK(n2927), .Q(
        g1756) );
  SDFFX1 DFF_411_Q_reg ( .D(g29), .SI(g1756), .SE(n2764), .CLK(n2927), .Q(
        g2604) );
  SDFFX1 DFF_412_Q_reg ( .D(g806), .SI(g2604), .SE(n2764), .CLK(n2927), .Q(
        g841) );
  SDFFX1 DFF_413_Q_reg ( .D(g6894), .SI(g841), .SE(n2844), .CLK(n2886), .Q(
        g1027), .QN(n2746) );
  SDFFX1 DFF_414_Q_reg ( .D(g6902), .SI(g1027), .SE(n2800), .CLK(n2908), .Q(
        g1003), .QN(n2700) );
  SDFFX1 DFF_415_Q_reg ( .D(g8765), .SI(g1003), .SE(n2800), .CLK(n2908), .Q(
        g1403), .QN(n2655) );
  SDFFX1 DFF_416_Q_reg ( .D(g4498), .SI(g1403), .SE(n2800), .CLK(n2909), .Q(
        g1145), .QN(n1617) );
  SDFFX1 DFF_417_Q_reg ( .D(g5148), .SI(g1145), .SE(n2793), .CLK(n2912), .Q(
        g1107), .QN(n1614) );
  SDFFX1 DFF_418_Q_reg ( .D(g7581), .SI(g1107), .SE(n2793), .CLK(n2912), .Q(
        g1223), .QN(n2509) );
  SDFFX1 DFF_419_Q_reg ( .D(g11267), .SI(g1223), .SE(n2829), .CLK(n2894), .Q(
        g406), .QN(n2631) );
  SDFFX1 DFF_420_Q_reg ( .D(g10936), .SI(g406), .SE(n2842), .CLK(n2887), .Q(
        g1811) );
  SDFFX1 DFF_421_Q_reg ( .D(g10784), .SI(g1811), .SE(n2799), .CLK(n2909), .Q(
        n3029), .QN(n4953) );
  SDFFX1 DFF_423_Q_reg ( .D(g10765), .SI(n3029), .SE(n2792), .CLK(n2912), .Q(
        g1654) );
  SDFFX1 DFF_424_Q_reg ( .D(g6332), .SI(g1654), .SE(n2806), .CLK(n2905), .Q(
        g197), .QN(n1678) );
  SDFFX1 DFF_425_Q_reg ( .D(g6479), .SI(g197), .SE(n2782), .CLK(n2917), .Q(
        g1595) );
  SDFFX1 DFF_426_Q_reg ( .D(g6537), .SI(g1595), .SE(n2766), .CLK(n2925), .Q(
        g1537) );
  SDFFX1 DFF_427_Q_reg ( .D(g8434), .SI(g1537), .SE(n2812), .CLK(n2903), .Q(
        g727) );
  SDFFX1 DFF_428_Q_reg ( .D(g6908), .SI(g727), .SE(n2761), .CLK(n2928), .Q(
        test_so8) );
  SDFFX1 DFF_429_Q_reg ( .D(g6243), .SI(test_si9), .SE(n2781), .CLK(n2918), 
        .Q(g798), .QN(n1717) );
  SDFFX1 DFF_430_Q_reg ( .D(g11324), .SI(g798), .SE(n2781), .CLK(n2918), .Q(
        g481) );
  SDFFX1 DFF_431_Q_reg ( .D(g3462), .SI(g481), .SE(n2781), .CLK(n2918), .Q(
        g4172), .QN(n1647) );
  SDFFX1 DFF_432_Q_reg ( .D(g11609), .SI(g4172), .SE(n2837), .CLK(n2890), .Q(
        g1330) );
  SDFFX1 DFF_433_Q_reg ( .D(g810), .SI(g1330), .SE(n2807), .CLK(n2905), .Q(
        g845), .QN(n2491) );
  SDFFX1 DFF_434_Q_reg ( .D(g8244), .SI(g845), .SE(n2788), .CLK(n2915), .Q(
        g4181), .QN(n2519) );
  SDFFX1 DFF_435_Q_reg ( .D(g8194), .SI(g4181), .SE(n2787), .CLK(n2915), .Q(
        g1512) );
  SDFFX1 DFF_436_Q_reg ( .D(g113), .SI(g1512), .SE(n2787), .CLK(n2915), .Q(
        n3027), .QN(n4930) );
  SDFFX1 DFF_437_Q_reg ( .D(g8052), .SI(n3027), .SE(n2787), .CLK(n2915), .Q(
        g1490) );
  SDFFX1 DFF_438_Q_reg ( .D(g4325), .SI(g1490), .SE(n2787), .CLK(n2915), .Q(
        g1166), .QN(n2667) );
  SDFFX1 DFF_440_Q_reg ( .D(g11481), .SI(g1166), .SE(n2787), .CLK(n2915), .Q(
        g348) );
  SDFFX1 DFF_441_Q_reg ( .D(g874), .SI(g348), .SE(n2787), .CLK(n2915), .Q(
        n3026), .QN(DFF_441_n1) );
  SDFFX1 DFF_442_Q_reg ( .D(g7301), .SI(n3026), .SE(n2822), .CLK(n2897), .Q(
        g1260), .QN(n2630) );
  SDFFX1 DFF_443_Q_reg ( .D(g6035), .SI(g1260), .SE(n2822), .CLK(n2897), .Q(
        g260) );
  SDFFX1 DFF_444_Q_reg ( .D(g8059), .SI(g260), .SE(n2801), .CLK(n2908), .Q(
        g131), .QN(n2644) );
  SDFFX1 DFF_445_Q_reg ( .D(g1854), .SI(g131), .SE(n2801), .CLK(n2908), .Q(
        n3025) );
  SDFFX1 DFF_446_Q_reg ( .D(g6015), .SI(n3025), .SE(n2801), .CLK(n2908), .Q(
        g258) );
  SDFFX1 DFF_447_Q_reg ( .D(g11330), .SI(g258), .SE(n2824), .CLK(n2897), .Q(
        g521), .QN(n1698) );
  SDFFX1 DFF_448_Q_reg ( .D(g11605), .SI(g521), .SE(n2824), .CLK(n2897), .Q(
        g1318) );
  SDFFX1 DFF_449_Q_reg ( .D(g8921), .SI(g1318), .SE(n2824), .CLK(n2897), .Q(
        g1872), .QN(n1616) );
  SDFFX1 DFF_450_Q_reg ( .D(g8883), .SI(g1872), .SE(n2817), .CLK(n2900), .Q(
        g677), .QN(n1656) );
  SDFFX1 DFF_451_Q_reg ( .D(g28), .SI(g677), .SE(n2817), .CLK(n2900), .Q(g2608) );
  SDFFX1 DFF_452_Q_reg ( .D(n2748), .SI(g2608), .SE(n2844), .CLK(n2887), .Q(
        n3024), .QN(n4931) );
  SDFFX1 DFF_453_Q_reg ( .D(g6523), .SI(n3024), .SE(n2798), .CLK(n2910), .Q(
        g1549), .QN(n2535) );
  SDFFX1 DFF_454_Q_reg ( .D(g11300), .SI(g1549), .SE(n2840), .CLK(n2888), .Q(
        g947), .QN(n2459) );
  SDFFX1 DFF_455_Q_reg ( .D(g9555), .SI(g947), .SE(n2840), .CLK(n2889), .Q(
        g1834), .QN(n1655) );
  SDFFX1 DFF_456_Q_reg ( .D(g6481), .SI(g1834), .SE(n2798), .CLK(n2910), .Q(
        g1598) );
  SDFFX1 DFF_457_Q_reg ( .D(g4471), .SI(g1598), .SE(n2798), .CLK(n2910), .Q(
        g1121), .QN(n1618) );
  SDFFX1 DFF_458_Q_reg ( .D(g11606), .SI(g1121), .SE(n2792), .CLK(n2913), .Q(
        g1321), .QN(n2476) );
  SDFFX1 DFF_459_Q_reg ( .D(g11335), .SI(g1321), .SE(n2778), .CLK(n2919), .Q(
        g506) );
  SDFFX1 DFF_460_Q_reg ( .D(g10791), .SI(g506), .SE(n2778), .CLK(n2919), .Q(
        g546) );
  SDFFX1 DFF_461_Q_reg ( .D(g8939), .SI(g546), .SE(n2827), .CLK(n2895), .Q(
        g1909), .QN(n2710) );
  SDFFX1 DFF_462_Q_reg ( .D(g83), .SI(g1909), .SE(n2827), .CLK(n2895), .Q(g755) );
  SDFFX1 DFF_463_Q_reg ( .D(g6529), .SI(g755), .SE(n2769), .CLK(n2924), .Q(
        g1552), .QN(n2533) );
  SDFFX1 DFF_464_Q_reg ( .D(g101), .SI(g1552), .SE(n2769), .CLK(n2924), .Q(
        g2610) );
  SDFFX1 DFF_465_Q_reg ( .D(g10776), .SI(g2610), .SE(n2769), .CLK(n2924), .Q(
        g1687) );
  SDFFX1 DFF_466_Q_reg ( .D(g6514), .SI(g1687), .SE(n2769), .CLK(n2924), .Q(
        g1586) );
  SDFFX1 DFF_467_Q_reg ( .D(g259), .SI(g1586), .SE(n2832), .CLK(n2893), .Q(
        g324), .QN(n2660) );
  SDFFX1 DFF_468_Q_reg ( .D(g4490), .SI(g324), .SE(n2832), .CLK(n2893), .Q(
        g1141), .QN(n1660) );
  SDFFX1 DFF_470_Q_reg ( .D(g11639), .SI(g1141), .SE(n2795), .CLK(n2911), .Q(
        g1341), .QN(n2705) );
  SDFFX1 DFF_471_Q_reg ( .D(g4089), .SI(g1341), .SE(n2795), .CLK(n2911), .Q(
        g1710) );
  SDFFX1 DFF_472_Q_reg ( .D(g10785), .SI(g1710), .SE(n2795), .CLK(n2911), .Q(
        n3023), .QN(n4952) );
  SDFFX1 DFF_473_Q_reg ( .D(g6179), .SI(n3023), .SE(n2843), .CLK(n2887), .Q(
        n3022), .QN(n4944) );
  SDFFX1 DFF_474_Q_reg ( .D(g8053), .SI(n3022), .SE(n2805), .CLK(n2906), .Q(
        g135), .QN(n2646) );
  SDFFX1 DFF_475_Q_reg ( .D(g11329), .SI(g135), .SE(n2824), .CLK(n2896), .Q(
        g525), .QN(n1695) );
  SDFFX1 DFF_476_Q_reg ( .D(g104), .SI(g525), .SE(n2824), .CLK(n2896), .Q(
        g2607) );
  SDFFX1 DFF_477_Q_reg ( .D(g6515), .SI(g2607), .SE(n2782), .CLK(n2917), .Q(
        g1607), .QN(n2530) );
  SDFFX1 DFF_478_Q_reg ( .D(g258), .SI(g1607), .SE(n2801), .CLK(n2908), .Q(
        g321), .QN(n2704) );
  SDFFX1 DFF_479_Q_reg ( .D(g7204), .SI(g321), .SE(n2775), .CLK(n2921), .Q(
        g8982), .QN(n1672) );
  SDFFX1 DFF_480_Q_reg ( .D(g11443), .SI(g8982), .SE(n2762), .CLK(n2928), .Q(
        g1275), .QN(n2697) );
  SDFFX1 DFF_481_Q_reg ( .D(g11603), .SI(g1275), .SE(n2762), .CLK(n2928), .Q(
        test_so9) );
  SDFFX1 DFF_482_Q_reg ( .D(g8770), .SI(test_si10), .SE(n2777), .CLK(n2920), 
        .Q(g1615) );
  SDFFX1 DFF_483_Q_reg ( .D(g11292), .SI(g1615), .SE(n2807), .CLK(n2905), .Q(
        g382) );
  SDFFX1 DFF_484_Q_reg ( .D(g6331), .SI(g382), .SE(n2807), .CLK(n2905), .Q(
        n3020), .QN(n4947) );
  SDFFX1 DFF_485_Q_reg ( .D(g6900), .SI(n3020), .SE(n2772), .CLK(n2923), .Q(
        g266), .QN(n2554) );
  SDFFX1 DFF_486_Q_reg ( .D(g7294), .SI(g266), .SE(n2821), .CLK(n2898), .Q(
        g1284), .QN(n1864) );
  SDFFX1 DFF_487_Q_reg ( .D(g6829), .SI(g1284), .SE(n2821), .CLK(n2898), .Q(
        n3019), .QN(n4945) );
  SDFFX1 DFF_488_Q_reg ( .D(g8428), .SI(n3019), .SE(n2767), .CLK(n2925), .Q(
        g673) );
  SDFFX1 DFF_489_Q_reg ( .D(g4904), .SI(g673), .SE(n2839), .CLK(n2889), .Q(
        n3018), .QN(DFF_489_n1) );
  SDFFX1 DFF_490_Q_reg ( .D(g8054), .SI(n3018), .SE(n2808), .CLK(n2904), .Q(
        g162), .QN(n2649) );
  SDFFX1 DFF_491_Q_reg ( .D(g11268), .SI(g162), .SE(n2829), .CLK(n2894), .Q(
        g411), .QN(n2686) );
  SDFFX1 DFF_492_Q_reg ( .D(g11262), .SI(g411), .SE(n2828), .CLK(n2895), .Q(
        g431) );
  SDFFX1 DFF_493_Q_reg ( .D(g8283), .SI(g431), .SE(n2828), .CLK(n2895), .Q(
        g1905), .QN(n2613) );
  SDFFX1 DFF_494_Q_reg ( .D(g6193), .SI(g1905), .SE(n2785), .CLK(n2916), .Q(
        g1515), .QN(n1627) );
  SDFFX1 DFF_495_Q_reg ( .D(g8776), .SI(g1515), .SE(n2809), .CLK(n2904), .Q(
        g1630), .QN(n2579) );
  SDFFX1 DFF_496_Q_reg ( .D(g7143), .SI(g1630), .SE(n2775), .CLK(n2921), .Q(
        g8976), .QN(n1671) );
  SDFFX1 DFF_497_Q_reg ( .D(g6898), .SI(g8976), .SE(n2762), .CLK(n2927), .Q(
        g991), .QN(n1871) );
  SDFFX1 DFF_498_Q_reg ( .D(g7291), .SI(g991), .SE(n2822), .CLK(n2898), .Q(
        g1300), .QN(n2636) );
  SDFFX1 DFF_499_Q_reg ( .D(g11478), .SI(g1300), .SE(n2833), .CLK(n2892), .Q(
        g339) );
  SDFFX1 DFF_500_Q_reg ( .D(g6000), .SI(g339), .SE(n2780), .CLK(n2918), .Q(
        g256) );
  SDFFX1 DFF_501_Q_reg ( .D(g4264), .SI(g256), .SE(n2780), .CLK(n2918), .Q(
        g1750), .QN(n2712) );
  SDFFX1 DFF_502_Q_reg ( .D(g102), .SI(g1750), .SE(n2780), .CLK(n2918), .Q(
        g2611) );
  SDFFX1 DFF_503_Q_reg ( .D(g8768), .SI(g2611), .SE(n2780), .CLK(n2919), .Q(
        g1440), .QN(n2720) );
  SDFFX1 DFF_504_Q_reg ( .D(g10863), .SI(g1440), .SE(n2780), .CLK(n2919), .Q(
        g1666) );
  SDFFX1 DFF_505_Q_reg ( .D(g6522), .SI(g1666), .SE(n2780), .CLK(n2919), .Q(
        g1528), .QN(n1635) );
  SDFFX1 DFF_506_Q_reg ( .D(g11641), .SI(g1528), .SE(n2804), .CLK(n2906), .Q(
        g1351), .QN(n1721) );
  SDFFX1 DFF_507_Q_reg ( .D(g10780), .SI(g1351), .SE(n2799), .CLK(n2909), .Q(
        n3017), .QN(n4955) );
  SDFFX1 DFF_508_Q_reg ( .D(g8044), .SI(n3017), .SE(n2765), .CLK(n2926), .Q(
        g127), .QN(n1704) );
  SDFFX1 DFF_509_Q_reg ( .D(g11579), .SI(g127), .SE(n2842), .CLK(n2888), .Q(
        g1618) );
  SDFFX1 DFF_510_Q_reg ( .D(g7296), .SI(g1618), .SE(n2762), .CLK(n2928), .Q(
        g1235), .QN(n2657) );
  SDFFX1 DFF_511_Q_reg ( .D(g6923), .SI(g1235), .SE(n2761), .CLK(n2928), .Q(
        g299) );
  SDFFX1 DFF_512_Q_reg ( .D(g11261), .SI(g299), .SE(n2828), .CLK(n2894), .Q(
        g435), .QN(n1878) );
  SDFFX1 DFF_513_Q_reg ( .D(g6638), .SI(g435), .SE(n2775), .CLK(n2921), .Q(
        g8981), .QN(n1664) );
  SDFFX1 DFF_514_Q_reg ( .D(g6534), .SI(g8981), .SE(n2767), .CLK(n2925), .Q(
        g1555), .QN(n2528) );
  SDFFX1 DFF_515_Q_reg ( .D(g6895), .SI(g1555), .SE(n2766), .CLK(n2925), .Q(
        g995), .QN(n2698) );
  SDFFX1 DFF_516_Q_reg ( .D(g8771), .SI(g995), .SE(n2836), .CLK(n2890), .Q(
        g1621) );
  SDFFX1 DFF_517_Q_reg ( .D(g4506), .SI(g1621), .SE(n2836), .CLK(n2891), .Q(
        n3016), .QN(n4950) );
  SDFFX1 DFF_518_Q_reg ( .D(g7441), .SI(n3016), .SE(n2768), .CLK(n2925), .Q(
        g643) );
  SDFFX1 DFF_519_Q_reg ( .D(g8055), .SI(g643), .SE(n2841), .CLK(n2888), .Q(
        g1494), .QN(n2687) );
  SDFFX1 DFF_520_Q_reg ( .D(g6468), .SI(g1494), .SE(n2783), .CLK(n2917), .Q(
        g1567), .QN(n2526) );
  SDFFX1 DFF_521_Q_reg ( .D(g8430), .SI(g1567), .SE(n2811), .CLK(n2903), .Q(
        g691) );
  SDFFX1 DFF_522_Q_reg ( .D(g11327), .SI(g691), .SE(n2825), .CLK(n2896), .Q(
        g534) );
  SDFFX1 DFF_523_Q_reg ( .D(g6508), .SI(g534), .SE(n2796), .CLK(n2911), .Q(
        g1776), .QN(n1715) );
  SDFFX1 DFF_524_Q_reg ( .D(g10717), .SI(g1776), .SE(n2794), .CLK(n2911), .Q(
        g569) );
  SDFFX1 DFF_525_Q_reg ( .D(g4334), .SI(g569), .SE(n2794), .CLK(n2912), .Q(
        g1160), .QN(n4932) );
  SDFFX1 DFF_526_Q_reg ( .D(n1585), .SI(g1160), .SE(n2794), .CLK(n2912), .Q(
        g1360) );
  SDFFX1 DFF_528_Q_reg ( .D(g6679), .SI(g1360), .SE(n2826), .CLK(n2896), .Q(g1) );
  SDFFX1 DFF_529_Q_reg ( .D(g11336), .SI(g1), .SE(n2826), .CLK(n2896), .Q(g511), .QN(n1679) );
  SDFFX1 DFF_530_Q_reg ( .D(g10771), .SI(g511), .SE(n2798), .CLK(n2909), .Q(
        g1724), .QN(n2484) );
  SDFFX1 DFF_531_Q_reg ( .D(g5445), .SI(g1724), .SE(n2798), .CLK(n2909), .Q(
        g12), .QN(n2622) );
  SDFFX1 DFF_532_Q_reg ( .D(g8559), .SI(g12), .SE(n2766), .CLK(n2926), .Q(
        g1878), .QN(n2620) );
  SDFFX1 DFF_533_Q_reg ( .D(g7219), .SI(g1878), .SE(n2766), .CLK(n2926), .Q(
        test_so10), .QN(n2756) );
  SDFFX1 DFF_158_Q_reg ( .D(g5390), .SI(n3053), .SE(n2793), .CLK(n2912), .Q(
        g1101), .QN(n1654) );
  AND2X2 Tg1_Trojan1 ( .IN1(g6179), .IN2(n2748), .Q(Tg1_OUT1) );
  AND2X2 Tg1_Trojan2 ( .IN1(n18), .IN2(n1132), .Q(Tg1_OUT2) );
  AND2X2 Tg1_Trojan3 ( .IN1(n1226), .IN2(n1858), .Q(Tg1_OUT3) );
  AND2X2 Tg1_Trojan4 ( .IN1(g5556), .IN2(n898), .Q(Tg1_OUT4) );
  AND4X1 Tg1_Trojan1234 ( .IN1(Tg1_OUT1), .IN2(Tg1_OUT2), .IN3(Tg1_OUT3), 
        .IN4(Tg1_OUT4) );
  NOR2X0 Tg1_Trojan5 ( .IN1(n1391), .IN2(n931), .QN(Tg1_OUT5) );
  NOR2X0 Tg1_Trojan6 ( .IN1(n857), .IN2(n902), .QN(Tg1_OUT6) );
  NOR2X0 Tg1_Trojan7 ( .IN1(n1239), .IN2(n1239), .QN(Tg1_OUT7) );
  NOR2X0 Tg1_Trojan8 ( .IN1(n1055), .IN2(n1016), .QN(Tg1_OUT8) );
  AND4X1 Tg1_Trojan5678 ( .IN1(Tg1_OUT5), .IN2(Tg1_OUT6), .IN3(Tg1_OUT7), 
        .IN4(Tg1_OUT8) );
  AND2X2 Tg2_Trojan1 ( .IN1(n938), .IN2(n16), .Q(Tg2_OUT1) );
  AND2X2 Tg2_Trojan2 ( .IN1(n16), .IN2(n16), .Q(Tg2_OUT2) );
  AND2X2 Tg2_Trojan3 ( .IN1(n16), .IN2(n16), .Q(Tg2_OUT3) );
  AND2X2 Tg2_Trojan4 ( .IN1(n16), .IN2(n16), .Q(Tg2_OUT4) );
  AND4X1 Tg2_Trojan1234 ( .IN1(Tg2_OUT1), .IN2(Tg2_OUT2), .IN3(Tg2_OUT3), 
        .IN4(Tg2_OUT4) );
  AND2X2 Tg2_Trojan5 ( .IN1(n1161), .IN2(n1154), .Q(Tg2_OUT5) );
  AND2X2 Tg2_Trojan6 ( .IN1(n1116), .IN2(n1162), .Q(Tg2_OUT6) );
  AND2X2 Tg2_Trojan7 ( .IN1(n1155), .IN2(n1107), .Q(Tg2_OUT7) );
  AND2X2 Tg2_Trojan8 ( .IN1(n929), .IN2(n97), .Q(Tg2_OUT8) );
  AND4X1 Tg2_Trojan5678 ( .IN1(Tg2_OUT5), .IN2(Tg2_OUT6), .IN3(Tg2_OUT7), 
        .IN4(Tg2_OUT8) );
  INVX0 TrojanINVtest_se ( .INP(n2846), .ZN(test_se_NOT) );
  AND2X2 Trojan_Trigger ( .IN1(1'b1), .IN2(test_se_NOT), .Q(Trigger_select) );
  MUX21X2 Trojan_Paylaod ( .IN1(g1200), .IN2(n968), .S(Trigger_select), .Q(
        g4207) );
  INVX0 U2788 ( .INP(g109), .ZN(n2757) );
  INVX0 U2789 ( .INP(g109), .ZN(n2758) );
  INVX0 U2790 ( .INP(g109), .ZN(n2759) );
  INVX0 U2791 ( .INP(g109), .ZN(n2760) );
  NAND2X1 U2792 ( .IN1(n4373), .IN2(n4374), .QN(n1239) );
  NBUFFX2 U2793 ( .INP(n2937), .Z(n2887) );
  NBUFFX2 U2794 ( .INP(n2937), .Z(n2888) );
  NBUFFX2 U2795 ( .INP(n2937), .Z(n2886) );
  NBUFFX2 U2796 ( .INP(n2930), .Z(n2919) );
  NBUFFX2 U2797 ( .INP(n2933), .Z(n2904) );
  NBUFFX2 U2798 ( .INP(n2936), .Z(n2889) );
  NBUFFX2 U2799 ( .INP(n2930), .Z(n2923) );
  NBUFFX2 U2800 ( .INP(n2932), .Z(n2910) );
  NBUFFX2 U2801 ( .INP(n2932), .Z(n2909) );
  NBUFFX2 U2802 ( .INP(n2931), .Z(n2916) );
  NBUFFX2 U2803 ( .INP(n2929), .Z(n2926) );
  NBUFFX2 U2804 ( .INP(n2931), .Z(n2914) );
  NBUFFX2 U2805 ( .INP(n2930), .Z(n2922) );
  NBUFFX2 U2806 ( .INP(n2933), .Z(n2906) );
  NBUFFX2 U2807 ( .INP(n2933), .Z(n2905) );
  NBUFFX2 U2808 ( .INP(n2930), .Z(n2921) );
  NBUFFX2 U2809 ( .INP(n2929), .Z(n2925) );
  NBUFFX2 U2810 ( .INP(n2932), .Z(n2913) );
  NBUFFX2 U2811 ( .INP(n2935), .Z(n2897) );
  NBUFFX2 U2812 ( .INP(n2929), .Z(n2927) );
  NBUFFX2 U2813 ( .INP(n2933), .Z(n2907) );
  NBUFFX2 U2814 ( .INP(n2931), .Z(n2918) );
  NBUFFX2 U2815 ( .INP(n2935), .Z(n2896) );
  NBUFFX2 U2816 ( .INP(n2929), .Z(n2924) );
  NBUFFX2 U2817 ( .INP(n2931), .Z(n2915) );
  NBUFFX2 U2818 ( .INP(n2936), .Z(n2891) );
  NBUFFX2 U2819 ( .INP(n2933), .Z(n2908) );
  NBUFFX2 U2820 ( .INP(n2935), .Z(n2898) );
  NBUFFX2 U2821 ( .INP(n2932), .Z(n2912) );
  NBUFFX2 U2822 ( .INP(n2934), .Z(n2899) );
  NBUFFX2 U2823 ( .INP(n2932), .Z(n2911) );
  NBUFFX2 U2824 ( .INP(n2934), .Z(n2902) );
  NBUFFX2 U2825 ( .INP(n2930), .Z(n2920) );
  NBUFFX2 U2826 ( .INP(n2931), .Z(n2917) );
  NBUFFX2 U2827 ( .INP(n2934), .Z(n2903) );
  NBUFFX2 U2828 ( .INP(n2936), .Z(n2893) );
  NBUFFX2 U2829 ( .INP(n2934), .Z(n2901) );
  NBUFFX2 U2830 ( .INP(n2934), .Z(n2900) );
  NBUFFX2 U2831 ( .INP(n2936), .Z(n2890) );
  NBUFFX2 U2832 ( .INP(n2935), .Z(n2894) );
  NBUFFX2 U2833 ( .INP(n2936), .Z(n2892) );
  NBUFFX2 U2834 ( .INP(n2935), .Z(n2895) );
  NBUFFX2 U2835 ( .INP(n2929), .Z(n2928) );
  NBUFFX2 U2836 ( .INP(n2875), .Z(n2761) );
  NBUFFX2 U2837 ( .INP(n2875), .Z(n2762) );
  NBUFFX2 U2838 ( .INP(n2874), .Z(n2763) );
  NBUFFX2 U2839 ( .INP(n2874), .Z(n2764) );
  NBUFFX2 U2840 ( .INP(n2874), .Z(n2765) );
  NBUFFX2 U2841 ( .INP(n2873), .Z(n2766) );
  NBUFFX2 U2842 ( .INP(n2873), .Z(n2767) );
  NBUFFX2 U2843 ( .INP(n2873), .Z(n2768) );
  NBUFFX2 U2844 ( .INP(n2872), .Z(n2769) );
  NBUFFX2 U2845 ( .INP(n2872), .Z(n2770) );
  NBUFFX2 U2849 ( .INP(n2872), .Z(n2771) );
  NBUFFX2 U2850 ( .INP(n2871), .Z(n2772) );
  NBUFFX2 U2851 ( .INP(n2871), .Z(n2773) );
  NBUFFX2 U2852 ( .INP(n2871), .Z(n2774) );
  NBUFFX2 U2853 ( .INP(n2870), .Z(n2775) );
  NBUFFX2 U2854 ( .INP(n2870), .Z(n2776) );
  NBUFFX2 U2855 ( .INP(n2870), .Z(n2777) );
  NBUFFX2 U2856 ( .INP(n2869), .Z(n2778) );
  NBUFFX2 U2857 ( .INP(n2869), .Z(n2779) );
  NBUFFX2 U2858 ( .INP(n2869), .Z(n2780) );
  NBUFFX2 U2862 ( .INP(n2868), .Z(n2781) );
  NBUFFX2 U2863 ( .INP(n2868), .Z(n2782) );
  NBUFFX2 U2864 ( .INP(n2868), .Z(n2783) );
  NBUFFX2 U2865 ( .INP(n2867), .Z(n2784) );
  NBUFFX2 U2866 ( .INP(n2867), .Z(n2785) );
  NBUFFX2 U2868 ( .INP(n2867), .Z(n2786) );
  NBUFFX2 U2869 ( .INP(n2866), .Z(n2787) );
  NBUFFX2 U2870 ( .INP(n2866), .Z(n2788) );
  NBUFFX2 U2871 ( .INP(n2866), .Z(n2789) );
  NBUFFX2 U2872 ( .INP(n2865), .Z(n2790) );
  NBUFFX2 U2873 ( .INP(n2865), .Z(n2791) );
  NBUFFX2 U2874 ( .INP(n2865), .Z(n2792) );
  NBUFFX2 U2875 ( .INP(n2864), .Z(n2793) );
  NBUFFX2 U2876 ( .INP(n2864), .Z(n2794) );
  NBUFFX2 U2877 ( .INP(n2864), .Z(n2795) );
  NBUFFX2 U2878 ( .INP(n2863), .Z(n2796) );
  NBUFFX2 U2880 ( .INP(n2863), .Z(n2797) );
  NBUFFX2 U2903 ( .INP(n2863), .Z(n2798) );
  NBUFFX2 U2904 ( .INP(n2862), .Z(n2799) );
  NBUFFX2 U2905 ( .INP(n2862), .Z(n2800) );
  NBUFFX2 U2906 ( .INP(n2862), .Z(n2801) );
  NBUFFX2 U2907 ( .INP(n2861), .Z(n2802) );
  NBUFFX2 U2908 ( .INP(n2861), .Z(n2803) );
  NBUFFX2 U2909 ( .INP(n2861), .Z(n2804) );
  NBUFFX2 U2910 ( .INP(n2860), .Z(n2805) );
  NBUFFX2 U2911 ( .INP(n2860), .Z(n2806) );
  NBUFFX2 U2912 ( .INP(n2860), .Z(n2807) );
  NBUFFX2 U2913 ( .INP(n2859), .Z(n2808) );
  NBUFFX2 U2914 ( .INP(n2859), .Z(n2809) );
  NBUFFX2 U2915 ( .INP(n2859), .Z(n2810) );
  NBUFFX2 U2916 ( .INP(n2858), .Z(n2811) );
  NBUFFX2 U2917 ( .INP(n2858), .Z(n2812) );
  NBUFFX2 U2918 ( .INP(n2858), .Z(n2813) );
  NBUFFX2 U2919 ( .INP(n2857), .Z(n2814) );
  NBUFFX2 U2920 ( .INP(n2857), .Z(n2815) );
  NBUFFX2 U2921 ( .INP(n2857), .Z(n2816) );
  NBUFFX2 U2922 ( .INP(n2856), .Z(n2817) );
  NBUFFX2 U2923 ( .INP(n2856), .Z(n2818) );
  NBUFFX2 U2924 ( .INP(n2856), .Z(n2819) );
  NBUFFX2 U2925 ( .INP(n2855), .Z(n2820) );
  NBUFFX2 U2926 ( .INP(n2855), .Z(n2821) );
  NBUFFX2 U2927 ( .INP(n2855), .Z(n2822) );
  NBUFFX2 U2928 ( .INP(n2854), .Z(n2823) );
  NBUFFX2 U2929 ( .INP(n2854), .Z(n2824) );
  NBUFFX2 U2930 ( .INP(n2854), .Z(n2825) );
  NBUFFX2 U2931 ( .INP(n2853), .Z(n2826) );
  NBUFFX2 U2932 ( .INP(n2853), .Z(n2827) );
  NBUFFX2 U2933 ( .INP(n2853), .Z(n2828) );
  NBUFFX2 U2934 ( .INP(n2852), .Z(n2829) );
  NBUFFX2 U2935 ( .INP(n2852), .Z(n2830) );
  NBUFFX2 U2936 ( .INP(n2852), .Z(n2831) );
  NBUFFX2 U2937 ( .INP(n2851), .Z(n2832) );
  NBUFFX2 U2938 ( .INP(n2851), .Z(n2833) );
  NBUFFX2 U2939 ( .INP(n2851), .Z(n2834) );
  NBUFFX2 U2940 ( .INP(n2850), .Z(n2835) );
  NBUFFX2 U2941 ( .INP(n2850), .Z(n2836) );
  NBUFFX2 U2942 ( .INP(n2850), .Z(n2837) );
  NBUFFX2 U2943 ( .INP(n2849), .Z(n2838) );
  NBUFFX2 U2944 ( .INP(n2849), .Z(n2839) );
  NBUFFX2 U2945 ( .INP(n2849), .Z(n2840) );
  NBUFFX2 U2946 ( .INP(n2848), .Z(n2841) );
  NBUFFX2 U2947 ( .INP(n2848), .Z(n2842) );
  NBUFFX2 U2948 ( .INP(n2848), .Z(n2843) );
  NBUFFX2 U2949 ( .INP(n2847), .Z(n2844) );
  NBUFFX2 U2950 ( .INP(n2847), .Z(n2845) );
  NBUFFX2 U2951 ( .INP(n2847), .Z(n2846) );
  NBUFFX2 U2952 ( .INP(n2885), .Z(n2847) );
  NBUFFX2 U2953 ( .INP(n2885), .Z(n2848) );
  NBUFFX2 U2954 ( .INP(n2884), .Z(n2849) );
  NBUFFX2 U2955 ( .INP(n2884), .Z(n2850) );
  NBUFFX2 U2956 ( .INP(n2884), .Z(n2851) );
  NBUFFX2 U2957 ( .INP(n2883), .Z(n2852) );
  NBUFFX2 U2958 ( .INP(n2883), .Z(n2853) );
  NBUFFX2 U2959 ( .INP(n2883), .Z(n2854) );
  NBUFFX2 U2960 ( .INP(n2882), .Z(n2855) );
  NBUFFX2 U2961 ( .INP(n2882), .Z(n2856) );
  NBUFFX2 U2962 ( .INP(n2882), .Z(n2857) );
  NBUFFX2 U2963 ( .INP(n2881), .Z(n2858) );
  NBUFFX2 U2964 ( .INP(n2881), .Z(n2859) );
  NBUFFX2 U2965 ( .INP(n2881), .Z(n2860) );
  NBUFFX2 U2966 ( .INP(n2880), .Z(n2861) );
  NBUFFX2 U2967 ( .INP(n2880), .Z(n2862) );
  NBUFFX2 U2968 ( .INP(n2880), .Z(n2863) );
  NBUFFX2 U2969 ( .INP(n2879), .Z(n2864) );
  NBUFFX2 U2970 ( .INP(n2879), .Z(n2865) );
  NBUFFX2 U2971 ( .INP(n2879), .Z(n2866) );
  NBUFFX2 U2972 ( .INP(n2878), .Z(n2867) );
  NBUFFX2 U2973 ( .INP(n2878), .Z(n2868) );
  NBUFFX2 U2974 ( .INP(n2878), .Z(n2869) );
  NBUFFX2 U2975 ( .INP(n2877), .Z(n2870) );
  NBUFFX2 U2976 ( .INP(n2877), .Z(n2871) );
  NBUFFX2 U2977 ( .INP(n2877), .Z(n2872) );
  NBUFFX2 U2978 ( .INP(n2876), .Z(n2873) );
  NBUFFX2 U2979 ( .INP(n2876), .Z(n2874) );
  NBUFFX2 U2980 ( .INP(n2876), .Z(n2875) );
  NBUFFX2 U2981 ( .INP(test_se), .Z(n2876) );
  NBUFFX2 U2982 ( .INP(n2881), .Z(n2877) );
  NBUFFX2 U2983 ( .INP(n2858), .Z(n2878) );
  NBUFFX2 U2984 ( .INP(n2859), .Z(n2879) );
  NBUFFX2 U2985 ( .INP(n2860), .Z(n2880) );
  NBUFFX2 U2986 ( .INP(test_se), .Z(n2881) );
  NBUFFX2 U2987 ( .INP(test_se), .Z(n2882) );
  NBUFFX2 U2988 ( .INP(n2875), .Z(n2883) );
  NBUFFX2 U2989 ( .INP(test_se), .Z(n2884) );
  NBUFFX2 U2990 ( .INP(n2876), .Z(n2885) );
  NBUFFX2 U2991 ( .INP(CK), .Z(n2929) );
  NBUFFX2 U2992 ( .INP(CK), .Z(n2930) );
  NBUFFX2 U2993 ( .INP(CK), .Z(n2931) );
  NBUFFX2 U2994 ( .INP(CK), .Z(n2932) );
  NBUFFX2 U2995 ( .INP(CK), .Z(n2933) );
  NBUFFX2 U2996 ( .INP(CK), .Z(n2934) );
  NBUFFX2 U2997 ( .INP(CK), .Z(n2935) );
  NBUFFX2 U2998 ( .INP(CK), .Z(n2936) );
  NBUFFX2 U2999 ( .INP(CK), .Z(n2937) );
  INVX0 U3001 ( .INP(n2938), .ZN(n97) );
  NAND2X0 U3002 ( .IN1(n2939), .IN2(n2940), .QN(n962) );
  OR2X1 U3003 ( .IN1(n902), .IN2(n1696), .Q(n2940) );
  NAND2X0 U3004 ( .IN1(n2941), .IN2(n1696), .QN(n2939) );
  INVX0 U3005 ( .INP(n2942), .ZN(n2941) );
  NAND2X0 U3006 ( .IN1(n2943), .IN2(n2944), .QN(n917) );
  OR2X1 U3007 ( .IN1(n857), .IN2(n1697), .Q(n2944) );
  NAND2X0 U3008 ( .IN1(n2945), .IN2(n1697), .QN(n2943) );
  NOR2X0 U3009 ( .IN1(n2946), .IN2(n2947), .QN(n838) );
  INVX0 U3010 ( .INP(n2948), .ZN(n343) );
  INVX0 U3011 ( .INP(n2949), .ZN(n28) );
  NOR2X0 U3012 ( .IN1(n2757), .IN2(n2950), .QN(n2749) );
  NOR2X0 U3013 ( .IN1(n2951), .IN2(n3064), .QN(n2950) );
  INVX0 U3014 ( .INP(n2952), .ZN(n2748) );
  INVX0 U3015 ( .INP(n2953), .ZN(n20) );
  NAND2X0 U3016 ( .IN1(n2954), .IN2(n2955), .QN(n1588) );
  NOR2X0 U3017 ( .IN1(g47), .IN2(g42), .QN(n2955) );
  NOR2X0 U3018 ( .IN1(n2956), .IN2(n2957), .QN(n2954) );
  NAND2X0 U3019 ( .IN1(n2958), .IN2(g46), .QN(n1587) );
  NAND2X0 U3020 ( .IN1(n2959), .IN2(n2960), .QN(n1586) );
  NOR2X0 U3021 ( .IN1(n2961), .IN2(n2962), .QN(n2959) );
  NAND2X0 U3022 ( .IN1(n2963), .IN2(n2960), .QN(n1585) );
  NOR2X0 U3023 ( .IN1(g42), .IN2(n2962), .QN(n2963) );
  OR2X1 U3024 ( .IN1(n2521), .IN2(n2520), .Q(n1214) );
  NAND2X0 U3025 ( .IN1(n1193), .IN2(g4176), .QN(n1153) );
  NAND2X0 U3026 ( .IN1(n2964), .IN2(g806), .QN(n1151) );
  INVX0 U3027 ( .INP(n2965), .ZN(n11) );
  NAND2X0 U3028 ( .IN1(n1125), .IN2(g4178), .QN(n1099) );
  NAND2X0 U3029 ( .IN1(n1123), .IN2(g814), .QN(n1097) );
  NOR2X0 U3030 ( .IN1(n2966), .IN2(n2967), .QN(g9721) );
  XOR2X1 U3031 ( .IN1(g611), .IN2(n2968), .Q(n2966) );
  NOR2X0 U3032 ( .IN1(n2969), .IN2(n2970), .QN(n2968) );
  INVX0 U3033 ( .INP(n2971), .ZN(n2970) );
  NOR2X0 U3034 ( .IN1(n2972), .IN2(n2973), .QN(n2969) );
  NOR2X0 U3035 ( .IN1(n2974), .IN2(g617), .QN(n2972) );
  NOR2X0 U3036 ( .IN1(n804), .IN2(n2975), .QN(n2974) );
  NOR2X0 U3037 ( .IN1(n2967), .IN2(n2976), .QN(g9555) );
  NAND2X0 U3038 ( .IN1(n2977), .IN2(n2978), .QN(n2976) );
  OR2X1 U3039 ( .IN1(n806), .IN2(g1834), .Q(n2978) );
  NAND2X0 U3040 ( .IN1(n2979), .IN2(g1834), .QN(n2977) );
  AND2X1 U3041 ( .IN1(n808), .IN2(n926), .Q(n2979) );
  NAND2X0 U3042 ( .IN1(n2695), .IN2(n2980), .QN(n808) );
  NAND2X0 U3043 ( .IN1(n168), .IN2(n2981), .QN(n2980) );
  INVX0 U3044 ( .INP(n2982), .ZN(n168) );
  NAND2X0 U3045 ( .IN1(n2983), .IN2(n2984), .QN(g9451) );
  NOR2X0 U3046 ( .IN1(g31), .IN2(g30), .QN(n2983) );
  NOR2X0 U3047 ( .IN1(n2967), .IN2(n2985), .QN(g9272) );
  NAND2X0 U3048 ( .IN1(n2986), .IN2(n2987), .QN(n2985) );
  NAND2X0 U3049 ( .IN1(n2988), .IN2(g1828), .QN(n2987) );
  NAND2X0 U3050 ( .IN1(n2989), .IN2(n1605), .QN(n2986) );
  NOR2X0 U3051 ( .IN1(n2990), .IN2(n2988), .QN(n2989) );
  AND2X1 U3052 ( .IN1(n812), .IN2(n2991), .Q(n2988) );
  NAND2X0 U3053 ( .IN1(n2992), .IN2(n2993), .QN(n2991) );
  NOR2X0 U3054 ( .IN1(n2994), .IN2(n2995), .QN(n2992) );
  NOR2X0 U3055 ( .IN1(n1605), .IN2(n2996), .QN(n2994) );
  NAND2X0 U3056 ( .IN1(g1814), .IN2(g1822), .QN(n2996) );
  NOR2X0 U3057 ( .IN1(n2997), .IN2(n2967), .QN(g9269) );
  XOR2X1 U3058 ( .IN1(g1822), .IN2(n2998), .Q(n2997) );
  NOR2X0 U3059 ( .IN1(n2999), .IN2(n3000), .QN(n2998) );
  NOR2X0 U3060 ( .IN1(n3001), .IN2(n2981), .QN(n3000) );
  NOR2X0 U3061 ( .IN1(n3002), .IN2(n3003), .QN(n3001) );
  NOR2X0 U3062 ( .IN1(n2981), .IN2(n3004), .QN(n2999) );
  NAND2X0 U3063 ( .IN1(n1643), .IN2(n3005), .QN(n3004) );
  NOR2X0 U3064 ( .IN1(n2967), .IN2(n3006), .QN(g9266) );
  XOR2X1 U3065 ( .IN1(n1608), .IN2(n3007), .Q(n3006) );
  NOR2X0 U3066 ( .IN1(n3008), .IN2(n2981), .QN(n3007) );
  INVX0 U3067 ( .INP(n812), .ZN(n2981) );
  NOR2X0 U3068 ( .IN1(n3009), .IN2(n3010), .QN(n3008) );
  NAND2X0 U3069 ( .IN1(n2982), .IN2(n3011), .QN(n3010) );
  NOR2X0 U3070 ( .IN1(n817), .IN2(g1822), .QN(n3009) );
  NOR2X0 U3071 ( .IN1(n2967), .IN2(n3012), .QN(g9150) );
  NAND2X0 U3072 ( .IN1(n3013), .IN2(n3014), .QN(n3012) );
  NAND2X0 U3073 ( .IN1(n3015), .IN2(g605), .QN(n3014) );
  NAND2X0 U3074 ( .IN1(n3021), .IN2(n1593), .QN(n3013) );
  NOR2X0 U3075 ( .IN1(n3015), .IN2(n3028), .QN(n3021) );
  AND2X1 U3076 ( .IN1(n804), .IN2(n3032), .Q(n3015) );
  NAND2X0 U3077 ( .IN1(n3039), .IN2(n3043), .QN(n3032) );
  NOR2X0 U3078 ( .IN1(n3049), .IN2(n3052), .QN(n3039) );
  NOR2X0 U3079 ( .IN1(n1644), .IN2(n3060), .QN(n3052) );
  NOR2X0 U3080 ( .IN1(n2975), .IN2(g622), .QN(n3049) );
  NOR2X0 U3081 ( .IN1(n3063), .IN2(n2967), .QN(g9124) );
  XOR2X1 U3082 ( .IN1(g599), .IN2(n836), .Q(n3063) );
  NOR2X0 U3083 ( .IN1(n3066), .IN2(n2967), .QN(g9110) );
  XOR2X1 U3084 ( .IN1(n3067), .IN2(n1607), .Q(n3066) );
  NAND2X0 U3085 ( .IN1(n837), .IN2(n3068), .QN(n3067) );
  NAND2X0 U3086 ( .IN1(n804), .IN2(n3069), .QN(n3068) );
  NAND2X0 U3087 ( .IN1(n2975), .IN2(n3070), .QN(n3069) );
  NAND2X0 U3088 ( .IN1(n3071), .IN2(n3072), .QN(n837) );
  NOR2X0 U3089 ( .IN1(g599), .IN2(n2947), .QN(n3071) );
  NAND2X0 U3091 ( .IN1(n3073), .IN2(n3074), .QN(g8973) );
  NAND2X0 U3093 ( .IN1(n3075), .IN2(n3076), .QN(n3074) );
  XNOR2X1 U3095 ( .IN1(n1615), .IN2(n3077), .Q(n3075) );
  NOR2X0 U3097 ( .IN1(n3078), .IN2(n3079), .QN(n3077) );
  NOR2X0 U3099 ( .IN1(n3080), .IN2(g664), .QN(n3078) );
  NAND2X0 U3100 ( .IN1(n3081), .IN2(n3082), .QN(g8945) );
  NAND2X0 U3101 ( .IN1(n3083), .IN2(n3084), .QN(n3082) );
  XNOR2X1 U3102 ( .IN1(n1697), .IN2(n3085), .Q(n3083) );
  NOR2X0 U3103 ( .IN1(n3086), .IN2(n3087), .QN(n3085) );
  NAND2X0 U3104 ( .IN1(n3088), .IN2(n3089), .QN(n3087) );
  NAND2X0 U3105 ( .IN1(n2696), .IN2(n3090), .QN(n3089) );
  NAND2X0 U3106 ( .IN1(n3091), .IN2(n3092), .QN(n3088) );
  NOR2X0 U3107 ( .IN1(n2945), .IN2(n3093), .QN(n3091) );
  INVX0 U3108 ( .INP(n857), .ZN(n3093) );
  NAND2X0 U3109 ( .IN1(n3094), .IN2(n3095), .QN(n857) );
  NOR2X0 U3110 ( .IN1(n1616), .IN2(n3096), .QN(n3095) );
  NAND2X0 U3111 ( .IN1(g1882), .IN2(g1936), .QN(n3096) );
  NOR2X0 U3112 ( .IN1(n3097), .IN2(n3098), .QN(n3094) );
  OR2X1 U3113 ( .IN1(n3099), .IN2(n3100), .Q(n3098) );
  AND2X1 U3114 ( .IN1(n3101), .IN2(n3102), .Q(n2945) );
  NOR2X0 U3115 ( .IN1(n3103), .IN2(n3104), .QN(n3102) );
  NOR2X0 U3116 ( .IN1(g1936), .IN2(g1927), .QN(n3101) );
  NAND2X0 U3117 ( .IN1(n3081), .IN2(n3105), .QN(g8944) );
  NAND2X0 U3118 ( .IN1(n3106), .IN2(n3084), .QN(n3105) );
  XOR2X1 U3119 ( .IN1(g1936), .IN2(n3107), .Q(n3106) );
  NOR2X0 U3120 ( .IN1(n3108), .IN2(n3086), .QN(n3107) );
  NOR2X0 U3121 ( .IN1(n3109), .IN2(n3110), .QN(n3108) );
  NAND2X0 U3122 ( .IN1(n3111), .IN2(n3112), .QN(n3110) );
  NAND2X0 U3123 ( .IN1(n3113), .IN2(n3114), .QN(n3112) );
  NOR2X0 U3125 ( .IN1(n3099), .IN2(n3097), .QN(n3113) );
  INVX0 U3126 ( .INP(n921), .ZN(n3097) );
  NAND2X0 U3127 ( .IN1(n3115), .IN2(n3116), .QN(n3111) );
  NOR2X0 U3128 ( .IN1(n3104), .IN2(g1927), .QN(n3115) );
  NOR2X0 U3129 ( .IN1(n2626), .IN2(n3092), .QN(n3109) );
  NAND2X0 U3130 ( .IN1(n3081), .IN2(n3117), .QN(g8943) );
  NAND2X0 U3131 ( .IN1(n3118), .IN2(n3084), .QN(n3117) );
  XOR2X1 U3132 ( .IN1(n3119), .IN2(n1663), .Q(n3118) );
  NAND2X0 U3133 ( .IN1(n3120), .IN2(n3121), .QN(n3119) );
  INVX0 U3134 ( .INP(n3122), .ZN(n3121) );
  NOR2X0 U3135 ( .IN1(n3123), .IN2(n3124), .QN(n3120) );
  NOR2X0 U3136 ( .IN1(n3092), .IN2(g1887), .QN(n3124) );
  NOR2X0 U3137 ( .IN1(n3125), .IN2(n3126), .QN(n3123) );
  NAND2X0 U3138 ( .IN1(n3081), .IN2(n3127), .QN(g8941) );
  NAND2X0 U3139 ( .IN1(n3128), .IN2(n3084), .QN(n3127) );
  XOR2X1 U3140 ( .IN1(n3129), .IN2(n2627), .Q(n3128) );
  NAND2X0 U3141 ( .IN1(n3130), .IN2(n3131), .QN(n3129) );
  NAND2X0 U3142 ( .IN1(n3132), .IN2(n3133), .QN(n3131) );
  NAND2X0 U3143 ( .IN1(n3090), .IN2(g1932), .QN(n3133) );
  NOR2X0 U3144 ( .IN1(n3134), .IN2(n3135), .QN(n3132) );
  NOR2X0 U3145 ( .IN1(n3104), .IN2(n3136), .QN(n3135) );
  NAND2X0 U3146 ( .IN1(n3137), .IN2(n2710), .QN(n3104) );
  AND2X1 U3147 ( .IN1(n1675), .IN2(n2681), .Q(n3137) );
  NOR2X0 U3148 ( .IN1(n3099), .IN2(n3138), .QN(n3134) );
  NAND2X0 U3149 ( .IN1(n3139), .IN2(g1900), .QN(n3099) );
  NOR2X0 U3150 ( .IN1(n2710), .IN2(n2681), .QN(n3139) );
  NAND2X0 U3151 ( .IN1(n3081), .IN2(n3140), .QN(g8940) );
  NAND2X0 U3152 ( .IN1(n3141), .IN2(n3084), .QN(n3140) );
  XNOR2X1 U3153 ( .IN1(n2681), .IN2(n3142), .Q(n3141) );
  NOR2X0 U3154 ( .IN1(n3143), .IN2(n3086), .QN(n3142) );
  NOR2X0 U3155 ( .IN1(n3144), .IN2(n3145), .QN(n3143) );
  NAND2X0 U3156 ( .IN1(n3146), .IN2(n3147), .QN(n3145) );
  NAND2X0 U3157 ( .IN1(n3148), .IN2(g1909), .QN(n3147) );
  NAND2X0 U3158 ( .IN1(n3149), .IN2(n2710), .QN(n3146) );
  NOR2X0 U3159 ( .IN1(n1718), .IN2(n3092), .QN(n3144) );
  NAND2X0 U3160 ( .IN1(n3081), .IN2(n3150), .QN(g8939) );
  NAND2X0 U3161 ( .IN1(n3151), .IN2(n3084), .QN(n3150) );
  XOR2X1 U3162 ( .IN1(n3152), .IN2(n2710), .Q(n3151) );
  NAND2X0 U3163 ( .IN1(n3153), .IN2(n3130), .QN(n3152) );
  NAND2X0 U3164 ( .IN1(n3154), .IN2(n3155), .QN(n3153) );
  NAND2X0 U3165 ( .IN1(n3090), .IN2(g1914), .QN(n3155) );
  NOR2X0 U3166 ( .IN1(n3148), .IN2(n3149), .QN(n3154) );
  NOR2X0 U3167 ( .IN1(g1900), .IN2(n3136), .QN(n3149) );
  NOR2X0 U3168 ( .IN1(n1675), .IN2(n3138), .QN(n3148) );
  NAND2X0 U3169 ( .IN1(n3081), .IN2(n3156), .QN(g8938) );
  NAND2X0 U3170 ( .IN1(n3157), .IN2(n3084), .QN(n3156) );
  XOR2X1 U3172 ( .IN1(g1900), .IN2(n3158), .Q(n3157) );
  NOR2X0 U3173 ( .IN1(n3086), .IN2(n3159), .QN(n3158) );
  NOR2X0 U3174 ( .IN1(n3160), .IN2(n3161), .QN(n3159) );
  NAND2X0 U3175 ( .IN1(n3136), .IN2(n3138), .QN(n3161) );
  NAND2X0 U3176 ( .IN1(n3114), .IN2(g1891), .QN(n3138) );
  NOR2X0 U3177 ( .IN1(n3162), .IN2(n3126), .QN(n3114) );
  NAND2X0 U3178 ( .IN1(g1882), .IN2(n3125), .QN(n3162) );
  INVX0 U3179 ( .INP(n3116), .ZN(n3136) );
  NOR2X0 U3180 ( .IN1(n3090), .IN2(n3103), .QN(n3116) );
  NAND2X0 U3181 ( .IN1(n3163), .IN2(n3164), .QN(n3103) );
  NOR2X0 U3182 ( .IN1(n3125), .IN2(g1872), .QN(n3164) );
  NOR2X0 U3183 ( .IN1(g1891), .IN2(g1882), .QN(n3163) );
  NOR2X0 U3184 ( .IN1(n2613), .IN2(n3092), .QN(n3160) );
  INVX0 U3185 ( .INP(n3130), .ZN(n3086) );
  NAND2X0 U3186 ( .IN1(n3081), .IN2(n3165), .QN(g8937) );
  NAND2X0 U3187 ( .IN1(n3166), .IN2(n3084), .QN(n3165) );
  XOR2X1 U3188 ( .IN1(n3167), .IN2(n1657), .Q(n3166) );
  NAND2X0 U3189 ( .IN1(n3168), .IN2(n3169), .QN(n3167) );
  NOR2X0 U3190 ( .IN1(n3170), .IN2(n3171), .QN(n3169) );
  NOR2X0 U3191 ( .IN1(g1882), .IN2(n3126), .QN(n3171) );
  NAND2X0 U3192 ( .IN1(n3092), .IN2(g1872), .QN(n3126) );
  NOR2X0 U3193 ( .IN1(n1663), .IN2(n3172), .QN(n3170) );
  NAND2X0 U3194 ( .IN1(n3092), .IN2(n3100), .QN(n3172) );
  NOR2X0 U3195 ( .IN1(n3173), .IN2(n3122), .QN(n3168) );
  NAND2X0 U3196 ( .IN1(n3130), .IN2(n3174), .QN(n3122) );
  NAND2X0 U3197 ( .IN1(n3175), .IN2(n3092), .QN(n3174) );
  NOR2X0 U3198 ( .IN1(n3100), .IN2(g1872), .QN(n3175) );
  INVX0 U3199 ( .INP(n3125), .ZN(n3100) );
  NAND2X0 U3200 ( .IN1(n3176), .IN2(n3177), .QN(n3125) );
  NAND2X0 U3201 ( .IN1(n1643), .IN2(g1814), .QN(n3177) );
  NOR2X0 U3202 ( .IN1(n3002), .IN2(n2995), .QN(n3176) );
  NOR2X0 U3203 ( .IN1(g1828), .IN2(n3011), .QN(n2995) );
  NOR2X0 U3204 ( .IN1(n3092), .IN2(g1896), .QN(n3173) );
  NAND2X0 U3205 ( .IN1(n3073), .IN2(n3178), .QN(g8926) );
  NAND2X0 U3206 ( .IN1(n3179), .IN2(n3076), .QN(n3178) );
  XNOR2X1 U3207 ( .IN1(n1696), .IN2(n898), .Q(n3179) );
  AND2X1 U3208 ( .IN1(n3180), .IN2(n3181), .Q(n898) );
  NOR2X0 U3209 ( .IN1(n3182), .IN2(n3183), .QN(n3180) );
  NOR2X0 U3210 ( .IN1(n3080), .IN2(g736), .QN(n3183) );
  NOR2X0 U3211 ( .IN1(n3184), .IN2(n3185), .QN(n3182) );
  NAND2X0 U3212 ( .IN1(n2942), .IN2(n902), .QN(n3185) );
  NAND2X0 U3213 ( .IN1(n3186), .IN2(n3187), .QN(n902) );
  NOR2X0 U3214 ( .IN1(n1615), .IN2(n3188), .QN(n3187) );
  NAND2X0 U3215 ( .IN1(g668), .IN2(g722), .QN(n3188) );
  NOR2X0 U3216 ( .IN1(n3189), .IN2(n3190), .QN(n3186) );
  NAND2X0 U3217 ( .IN1(n3191), .IN2(n3192), .QN(n3190) );
  INVX0 U3218 ( .INP(n967), .ZN(n3189) );
  NAND2X0 U3219 ( .IN1(n3193), .IN2(n3194), .QN(n2942) );
  NOR2X0 U3220 ( .IN1(g722), .IN2(n3195), .QN(n3194) );
  NAND2X0 U3221 ( .IN1(n1676), .IN2(n3196), .QN(n3195) );
  NOR2X0 U3222 ( .IN1(g695), .IN2(n3197), .QN(n3193) );
  NAND2X0 U3223 ( .IN1(n3073), .IN2(n3198), .QN(g8923) );
  NAND2X0 U3224 ( .IN1(n3199), .IN2(n3076), .QN(n3198) );
  XOR2X1 U3225 ( .IN1(n3200), .IN2(n1693), .Q(n3199) );
  NAND2X0 U3226 ( .IN1(n3181), .IN2(n3201), .QN(n3200) );
  NAND2X0 U3227 ( .IN1(n3202), .IN2(n3203), .QN(n3201) );
  NAND2X0 U3228 ( .IN1(n3184), .IN2(g727), .QN(n3203) );
  NOR2X0 U3229 ( .IN1(n3204), .IN2(n3205), .QN(n3202) );
  NOR2X0 U3230 ( .IN1(n3206), .IN2(n3197), .QN(n3205) );
  NAND2X0 U3231 ( .IN1(n2682), .IN2(n2515), .QN(n3197) );
  NOR2X0 U3232 ( .IN1(n3207), .IN2(n3208), .QN(n3204) );
  NAND2X0 U3233 ( .IN1(n967), .IN2(n3191), .QN(n3208) );
  INVX0 U3234 ( .INP(n3209), .ZN(n3191) );
  NAND2X0 U3235 ( .IN1(n3073), .IN2(n3210), .QN(g8922) );
  NAND2X0 U3236 ( .IN1(n3211), .IN2(n3076), .QN(n3210) );
  XOR2X1 U3237 ( .IN1(n3212), .IN2(n1662), .Q(n3211) );
  NAND2X0 U3238 ( .IN1(n3213), .IN2(n3214), .QN(n3212) );
  INVX0 U3239 ( .INP(n3215), .ZN(n3214) );
  NOR2X0 U3240 ( .IN1(n3216), .IN2(n3217), .QN(n3213) );
  NOR2X0 U3241 ( .IN1(n3080), .IN2(g673), .QN(n3217) );
  NOR2X0 U3242 ( .IN1(n3192), .IN2(n3218), .QN(n3216) );
  NAND2X0 U3243 ( .IN1(n3081), .IN2(n3219), .QN(g8921) );
  NAND2X0 U3244 ( .IN1(n3220), .IN2(n3084), .QN(n3219) );
  XOR2X1 U3245 ( .IN1(n3221), .IN2(n1616), .Q(n3220) );
  NAND2X0 U3246 ( .IN1(n3130), .IN2(n3222), .QN(n3221) );
  NAND2X0 U3247 ( .IN1(n2620), .IN2(n3090), .QN(n3222) );
  INVX0 U3248 ( .INP(n3092), .ZN(n3090) );
  NAND2X0 U3249 ( .IN1(n3092), .IN2(n918), .QN(n3130) );
  NAND2X0 U3250 ( .IN1(n3223), .IN2(n926), .QN(n918) );
  NAND2X0 U3251 ( .IN1(n3224), .IN2(n2982), .QN(n3223) );
  NAND2X0 U3252 ( .IN1(n3225), .IN2(n2695), .QN(n2982) );
  NOR2X0 U3253 ( .IN1(n1655), .IN2(n1608), .QN(n3225) );
  NAND2X0 U3254 ( .IN1(g1857), .IN2(n3226), .QN(n3224) );
  NAND2X0 U3255 ( .IN1(n1643), .IN2(n1605), .QN(n3226) );
  NOR2X0 U3256 ( .IN1(n3227), .IN2(n929), .QN(n3092) );
  NAND2X0 U3257 ( .IN1(n3228), .IN2(n3229), .QN(n3081) );
  NOR2X0 U3258 ( .IN1(n3084), .IN2(n3002), .QN(n3229) );
  INVX0 U3259 ( .INP(n2993), .ZN(n3002) );
  NOR2X0 U3260 ( .IN1(n2990), .IN2(n812), .QN(n3084) );
  AND2X1 U3261 ( .IN1(n916), .IN2(n3230), .Q(n3228) );
  NAND2X0 U3262 ( .IN1(n3073), .IN2(n3231), .QN(g8920) );
  NAND2X0 U3263 ( .IN1(n3232), .IN2(n3076), .QN(n3231) );
  XOR2X1 U3264 ( .IN1(n2515), .IN2(n931), .Q(n3232) );
  NAND2X0 U3265 ( .IN1(n3181), .IN2(n3233), .QN(n931) );
  NAND2X0 U3266 ( .IN1(n3234), .IN2(n3235), .QN(n3233) );
  NAND2X0 U3267 ( .IN1(n3184), .IN2(g718), .QN(n3235) );
  NOR2X0 U3268 ( .IN1(n3236), .IN2(n3237), .QN(n3234) );
  AND2X1 U3269 ( .IN1(n2682), .IN2(n3238), .Q(n3237) );
  NOR2X0 U3270 ( .IN1(n3209), .IN2(n3239), .QN(n3236) );
  NAND2X0 U3271 ( .IN1(n3240), .IN2(g686), .QN(n3209) );
  NOR2X0 U3272 ( .IN1(n2711), .IN2(n2682), .QN(n3240) );
  NAND2X0 U3273 ( .IN1(n3073), .IN2(n3241), .QN(g8889) );
  NAND2X0 U3274 ( .IN1(n3242), .IN2(n3076), .QN(n3241) );
  XNOR2X1 U3275 ( .IN1(n938), .IN2(n2682), .Q(n3242) );
  AND2X1 U3276 ( .IN1(n3243), .IN2(n3181), .Q(n938) );
  NAND2X0 U3277 ( .IN1(n3244), .IN2(n3245), .QN(n3243) );
  NAND2X0 U3278 ( .IN1(n3184), .IN2(g709), .QN(n3245) );
  NOR2X0 U3279 ( .IN1(n3238), .IN2(n3246), .QN(n3244) );
  NOR2X0 U3280 ( .IN1(n3239), .IN2(n3247), .QN(n3246) );
  NAND2X0 U3281 ( .IN1(g686), .IN2(g695), .QN(n3247) );
  INVX0 U3282 ( .INP(n3248), .ZN(n3239) );
  INVX0 U3283 ( .INP(n3206), .ZN(n3238) );
  NAND2X0 U3284 ( .IN1(n3249), .IN2(n3250), .QN(n3206) );
  NOR2X0 U3285 ( .IN1(g686), .IN2(g695), .QN(n3249) );
  NAND2X0 U3286 ( .IN1(n3073), .IN2(n3251), .QN(g8887) );
  NAND2X0 U3287 ( .IN1(n3252), .IN2(n3076), .QN(n3251) );
  XOR2X1 U3288 ( .IN1(g695), .IN2(n3253), .Q(n3252) );
  NOR2X0 U3289 ( .IN1(n3079), .IN2(n3254), .QN(n3253) );
  NOR2X0 U3290 ( .IN1(n3255), .IN2(n3256), .QN(n3254) );
  NAND2X0 U3291 ( .IN1(n3257), .IN2(n3258), .QN(n3256) );
  NAND2X0 U3292 ( .IN1(n3248), .IN2(g686), .QN(n3258) );
  NAND2X0 U3293 ( .IN1(n3250), .IN2(n1676), .QN(n3257) );
  NOR2X0 U3294 ( .IN1(n2680), .IN2(n3080), .QN(n3255) );
  INVX0 U3295 ( .INP(n3181), .ZN(n3079) );
  NAND2X0 U3296 ( .IN1(n3073), .IN2(n3259), .QN(g8885) );
  NAND2X0 U3297 ( .IN1(n3260), .IN2(n3076), .QN(n3259) );
  XOR2X1 U3298 ( .IN1(n3261), .IN2(n1676), .Q(n3260) );
  NAND2X0 U3299 ( .IN1(n3262), .IN2(n3181), .QN(n3261) );
  NAND2X0 U3300 ( .IN1(n3263), .IN2(n3264), .QN(n3262) );
  NAND2X0 U3301 ( .IN1(n3184), .IN2(g691), .QN(n3264) );
  NOR2X0 U3302 ( .IN1(n3248), .IN2(n3250), .QN(n3263) );
  AND2X1 U3303 ( .IN1(n3196), .IN2(n3080), .Q(n3250) );
  AND2X1 U3304 ( .IN1(n3265), .IN2(n3266), .Q(n3196) );
  AND2X1 U3305 ( .IN1(n3267), .IN2(n1615), .Q(n3266) );
  AND2X1 U3306 ( .IN1(n1656), .IN2(n1662), .Q(n3265) );
  NOR2X0 U3307 ( .IN1(n3207), .IN2(n1656), .QN(n3248) );
  NAND2X0 U3308 ( .IN1(n3268), .IN2(n3269), .QN(n3207) );
  NOR2X0 U3309 ( .IN1(n1662), .IN2(n3267), .QN(n3268) );
  NAND2X0 U3310 ( .IN1(n3073), .IN2(n3270), .QN(g8883) );
  NAND2X0 U3311 ( .IN1(n3271), .IN2(n3076), .QN(n3270) );
  INVX0 U3312 ( .INP(n3272), .ZN(n3076) );
  XOR2X1 U3313 ( .IN1(n3273), .IN2(n1656), .Q(n3271) );
  NAND2X0 U3314 ( .IN1(n3274), .IN2(n3275), .QN(n3273) );
  NOR2X0 U3315 ( .IN1(n3276), .IN2(n3277), .QN(n3275) );
  NOR2X0 U3316 ( .IN1(g668), .IN2(n3218), .QN(n3277) );
  INVX0 U3317 ( .INP(n3269), .ZN(n3218) );
  NOR2X0 U3318 ( .IN1(n3184), .IN2(n1615), .QN(n3269) );
  NOR2X0 U3319 ( .IN1(n1662), .IN2(n3278), .QN(n3276) );
  NAND2X0 U3320 ( .IN1(n3267), .IN2(n3080), .QN(n3278) );
  NOR2X0 U3321 ( .IN1(n3279), .IN2(n3215), .QN(n3274) );
  NAND2X0 U3322 ( .IN1(n3181), .IN2(n3280), .QN(n3215) );
  NAND2X0 U3323 ( .IN1(n3281), .IN2(n1615), .QN(n3280) );
  NOR2X0 U3324 ( .IN1(n3184), .IN2(n3267), .QN(n3281) );
  INVX0 U3325 ( .INP(n3192), .ZN(n3267) );
  NAND2X0 U3326 ( .IN1(n3043), .IN2(n3282), .QN(n3192) );
  NAND2X0 U3327 ( .IN1(n1644), .IN2(g591), .QN(n3282) );
  AND2X1 U3328 ( .IN1(n3283), .IN2(n3284), .Q(n3043) );
  NAND2X0 U3329 ( .IN1(n1593), .IN2(n3285), .QN(n3284) );
  INVX0 U3330 ( .INP(n3080), .ZN(n3184) );
  NAND2X0 U3331 ( .IN1(n958), .IN2(n3080), .QN(n3181) );
  NAND2X0 U3332 ( .IN1(n3286), .IN2(n3287), .QN(n958) );
  NAND2X0 U3333 ( .IN1(n3288), .IN2(n2975), .QN(n3287) );
  NAND2X0 U3334 ( .IN1(g639), .IN2(n3289), .QN(n3288) );
  NAND2X0 U3335 ( .IN1(n1644), .IN2(n1593), .QN(n3289) );
  NOR2X0 U3336 ( .IN1(n3080), .IN2(g682), .QN(n3279) );
  NAND2X0 U3337 ( .IN1(n3286), .IN2(n3290), .QN(n3080) );
  NAND2X0 U3338 ( .IN1(n1645), .IN2(n3291), .QN(n3290) );
  NAND2X0 U3339 ( .IN1(n3292), .IN2(n3293), .QN(n3291) );
  NAND2X0 U3340 ( .IN1(n3294), .IN2(n3295), .QN(n3073) );
  AND2X1 U3341 ( .IN1(n3272), .IN2(n2975), .Q(n3295) );
  NOR2X0 U3342 ( .IN1(n3028), .IN2(n3296), .QN(n3294) );
  NAND2X0 U3343 ( .IN1(n2971), .IN2(n3297), .QN(g8820) );
  NAND2X0 U3344 ( .IN1(n3298), .IN2(g622), .QN(n3297) );
  NAND2X0 U3345 ( .IN1(n3272), .IN2(n3299), .QN(n3298) );
  NAND2X0 U3346 ( .IN1(n3300), .IN2(n2975), .QN(n3299) );
  NAND2X0 U3347 ( .IN1(n3300), .IN2(n2947), .QN(n3272) );
  NAND2X0 U3348 ( .IN1(n3301), .IN2(n1713), .QN(n2971) );
  NOR2X0 U3349 ( .IN1(n2947), .IN2(n2975), .QN(n3301) );
  NAND2X0 U3350 ( .IN1(n3302), .IN2(n1645), .QN(n2975) );
  NOR2X0 U3351 ( .IN1(n1609), .IN2(n1607), .QN(n3302) );
  INVX0 U3352 ( .INP(n804), .ZN(n2947) );
  NAND2X0 U3353 ( .IN1(n3303), .IN2(n3304), .QN(g8779) );
  NAND2X0 U3354 ( .IN1(n968), .IN2(g1636), .QN(n3304) );
  NAND2X0 U3355 ( .IN1(n3305), .IN2(n3306), .QN(n3303) );
  NAND2X0 U3356 ( .IN1(n3307), .IN2(n3308), .QN(g8777) );
  NAND2X0 U3357 ( .IN1(n968), .IN2(g1633), .QN(n3308) );
  NAND2X0 U3358 ( .IN1(n3309), .IN2(n3306), .QN(n3307) );
  NAND2X0 U3359 ( .IN1(n3310), .IN2(n3311), .QN(g8776) );
  OR2X1 U3360 ( .IN1(n3306), .IN2(n2579), .Q(n3311) );
  NAND2X0 U3361 ( .IN1(n3312), .IN2(n3306), .QN(n3310) );
  NOR2X0 U3362 ( .IN1(n2758), .IN2(n3313), .QN(g8775) );
  XOR2X1 U3363 ( .IN1(n3314), .IN2(n2719), .Q(n3313) );
  NAND2X0 U3364 ( .IN1(n3315), .IN2(n3316), .QN(g8774) );
  OR2X1 U3365 ( .IN1(n3306), .IN2(n2582), .Q(n3316) );
  NAND2X0 U3366 ( .IN1(n3314), .IN2(n3306), .QN(n3315) );
  NAND2X0 U3367 ( .IN1(n3317), .IN2(n3318), .QN(n3314) );
  NAND2X0 U3368 ( .IN1(n3319), .IN2(n2967), .QN(n3318) );
  XOR2X1 U3369 ( .IN1(n3320), .IN2(n1706), .Q(n3319) );
  NAND2X0 U3370 ( .IN1(n3321), .IN2(n3322), .QN(n3320) );
  NOR2X0 U3371 ( .IN1(n1614), .IN2(g1101), .QN(n3321) );
  NAND2X0 U3372 ( .IN1(n3323), .IN2(n3324), .QN(g8773) );
  NAND2X0 U3373 ( .IN1(n968), .IN2(g1624), .QN(n3324) );
  NAND2X0 U3374 ( .IN1(n3325), .IN2(n3306), .QN(n3323) );
  NOR2X0 U3375 ( .IN1(n2759), .IN2(n3326), .QN(g8772) );
  XOR2X1 U3376 ( .IN1(n3312), .IN2(n2720), .Q(n3326) );
  NAND2X0 U3377 ( .IN1(n3327), .IN2(n3328), .QN(n3312) );
  NAND2X0 U3378 ( .IN1(n3329), .IN2(n2967), .QN(n3328) );
  XOR2X1 U3379 ( .IN1(n3330), .IN2(n1597), .Q(n3329) );
  NAND2X0 U3380 ( .IN1(n3331), .IN2(n3322), .QN(n3330) );
  INVX0 U3381 ( .INP(n3332), .ZN(n3322) );
  NOR2X0 U3382 ( .IN1(n1654), .IN2(n1614), .QN(n3331) );
  NAND2X0 U3383 ( .IN1(n3333), .IN2(n3334), .QN(g8771) );
  NAND2X0 U3384 ( .IN1(n968), .IN2(g1621), .QN(n3334) );
  NAND2X0 U3385 ( .IN1(n3335), .IN2(n3306), .QN(n3333) );
  NAND2X0 U3386 ( .IN1(n3336), .IN2(n3337), .QN(g8770) );
  NAND2X0 U3387 ( .IN1(n968), .IN2(g1615), .QN(n3337) );
  NAND2X0 U3388 ( .IN1(n3338), .IN2(n3306), .QN(n3336) );
  NOR2X0 U3389 ( .IN1(n2760), .IN2(n3339), .QN(g8769) );
  XOR2X1 U3390 ( .IN1(n3338), .IN2(n2721), .Q(n3339) );
  NAND2X0 U3391 ( .IN1(n3340), .IN2(n3341), .QN(n3338) );
  NAND2X0 U3392 ( .IN1(n3342), .IN2(n2967), .QN(n3341) );
  XOR2X1 U3393 ( .IN1(n3343), .IN2(n1618), .Q(n3342) );
  OR2X1 U3394 ( .IN1(n3332), .IN2(n3344), .Q(n3343) );
  NOR2X0 U3395 ( .IN1(n2757), .IN2(n3345), .QN(g8768) );
  XOR2X1 U3396 ( .IN1(n3309), .IN2(n2722), .Q(n3345) );
  NAND2X0 U3397 ( .IN1(n3346), .IN2(n3347), .QN(n3309) );
  NAND2X0 U3398 ( .IN1(n3348), .IN2(n2967), .QN(n3346) );
  XNOR2X1 U3399 ( .IN1(n1660), .IN2(n3349), .Q(n3348) );
  NOR2X0 U3400 ( .IN1(n3350), .IN2(g1101), .QN(n3349) );
  NOR2X0 U3401 ( .IN1(n2758), .IN2(n3351), .QN(g8767) );
  XOR2X1 U3402 ( .IN1(n3335), .IN2(n2655), .Q(n3351) );
  NAND2X0 U3403 ( .IN1(n3352), .IN2(n3353), .QN(n3335) );
  NAND2X0 U3404 ( .IN1(n3354), .IN2(n2967), .QN(n3353) );
  XOR2X1 U3405 ( .IN1(n3355), .IN2(n1708), .Q(n3354) );
  NAND2X0 U3406 ( .IN1(n3356), .IN2(n1654), .QN(n3355) );
  NOR2X0 U3407 ( .IN1(n2759), .IN2(n3357), .QN(g8766) );
  XOR2X1 U3408 ( .IN1(n3305), .IN2(n2653), .Q(n3357) );
  NAND2X0 U3409 ( .IN1(n3358), .IN2(n3359), .QN(n3305) );
  NAND2X0 U3410 ( .IN1(n3360), .IN2(n2967), .QN(n3358) );
  XOR2X1 U3411 ( .IN1(n3361), .IN2(n1617), .Q(n3360) );
  OR2X1 U3412 ( .IN1(n3350), .IN2(n1654), .Q(n3361) );
  NAND2X0 U3413 ( .IN1(n3362), .IN2(n1658), .QN(n3350) );
  AND2X1 U3414 ( .IN1(g1110), .IN2(n1614), .Q(n3362) );
  NOR2X0 U3415 ( .IN1(n2760), .IN2(n3363), .QN(g8765) );
  XOR2X1 U3416 ( .IN1(n3325), .IN2(n2654), .Q(n3363) );
  NAND2X0 U3417 ( .IN1(n3364), .IN2(n3365), .QN(n3325) );
  NAND2X0 U3418 ( .IN1(n3366), .IN2(n2967), .QN(n3365) );
  XOR2X1 U3419 ( .IN1(n3367), .IN2(n1705), .Q(n3366) );
  NAND2X0 U3420 ( .IN1(n3356), .IN2(g1101), .QN(n3367) );
  AND2X1 U3421 ( .IN1(n3368), .IN2(n1677), .Q(n3356) );
  NOR2X0 U3422 ( .IN1(n1614), .IN2(g1104), .QN(n3368) );
  NAND2X0 U3423 ( .IN1(n3369), .IN2(n3300), .QN(g8649) );
  NOR2X0 U3424 ( .IN1(n3370), .IN2(n3371), .QN(n3369) );
  NOR2X0 U3425 ( .IN1(n2621), .IN2(n3372), .QN(n3371) );
  NOR2X0 U3426 ( .IN1(n2694), .IN2(n1016), .QN(n3370) );
  NAND2X0 U3427 ( .IN1(n3373), .IN2(n3374), .QN(g8631) );
  NAND2X0 U3428 ( .IN1(n3375), .IN2(n3300), .QN(n3374) );
  NAND2X0 U3429 ( .IN1(n3376), .IN2(n3377), .QN(n3375) );
  NAND2X0 U3430 ( .IN1(n3378), .IN2(g636), .QN(n3377) );
  NAND2X0 U3431 ( .IN1(n3379), .IN2(n3380), .QN(n3378) );
  XOR2X1 U3432 ( .IN1(n3381), .IN2(n3382), .Q(n3380) );
  NAND2X0 U3433 ( .IN1(n3383), .IN2(n3384), .QN(n3382) );
  NAND2X0 U3434 ( .IN1(n3070), .IN2(g639), .QN(n3384) );
  NAND2X0 U3435 ( .IN1(n3385), .IN2(n1692), .QN(n3383) );
  NOR2X0 U3436 ( .IN1(n3072), .IN2(g611), .QN(n3385) );
  NAND2X0 U3437 ( .IN1(g255), .IN2(g622), .QN(n3381) );
  NOR2X0 U3438 ( .IN1(n3386), .IN2(n3387), .QN(n3379) );
  NOR2X0 U3439 ( .IN1(n3388), .IN2(n3389), .QN(n3386) );
  NAND2X0 U3440 ( .IN1(n3390), .IN2(n3060), .QN(n3389) );
  OR2X1 U3441 ( .IN1(n3283), .IN2(g622), .Q(n3376) );
  NAND2X0 U3442 ( .IN1(n3028), .IN2(n3391), .QN(n3373) );
  NAND2X0 U3443 ( .IN1(n3392), .IN2(n3393), .QN(n3391) );
  NAND2X0 U3444 ( .IN1(n3394), .IN2(n3395), .QN(n3393) );
  OR2X1 U3445 ( .IN1(n2726), .IN2(n1622), .Q(n3394) );
  NOR2X0 U3446 ( .IN1(n1716), .IN2(n3396), .QN(n3392) );
  NOR2X0 U3447 ( .IN1(n3397), .IN2(n3398), .QN(n3396) );
  NOR2X0 U3448 ( .IN1(n2739), .IN2(n2740), .QN(n3398) );
  NOR2X0 U3449 ( .IN1(n2737), .IN2(n2738), .QN(n3397) );
  NAND2X0 U3450 ( .IN1(n3399), .IN2(n3400), .QN(g8566) );
  NAND2X0 U3451 ( .IN1(n1653), .IN2(g1669), .QN(n3400) );
  NAND2X0 U3452 ( .IN1(g1690), .IN2(g1687), .QN(n3399) );
  NAND2X0 U3453 ( .IN1(n3401), .IN2(n3402), .QN(g8565) );
  NAND2X0 U3454 ( .IN1(n1653), .IN2(g1666), .QN(n3402) );
  NAND2X0 U3455 ( .IN1(g1690), .IN2(g1684), .QN(n3401) );
  NAND2X0 U3456 ( .IN1(n3403), .IN2(n3404), .QN(g8564) );
  NAND2X0 U3457 ( .IN1(n1653), .IN2(g1663), .QN(n3404) );
  NAND2X0 U3458 ( .IN1(g1690), .IN2(g1681), .QN(n3403) );
  NAND2X0 U3459 ( .IN1(n3405), .IN2(n3406), .QN(g8563) );
  NAND2X0 U3460 ( .IN1(n1653), .IN2(g1660), .QN(n3406) );
  NAND2X0 U3461 ( .IN1(g1690), .IN2(g1678), .QN(n3405) );
  NAND2X0 U3462 ( .IN1(n3407), .IN2(n3408), .QN(g8562) );
  NAND2X0 U3463 ( .IN1(n1653), .IN2(g1657), .QN(n3408) );
  NAND2X0 U3464 ( .IN1(g1690), .IN2(g1675), .QN(n3407) );
  NAND2X0 U3465 ( .IN1(n3409), .IN2(n3410), .QN(g8561) );
  NAND2X0 U3466 ( .IN1(n1653), .IN2(g1654), .QN(n3410) );
  NAND2X0 U3467 ( .IN1(g1690), .IN2(g1672), .QN(n3409) );
  NAND2X0 U3468 ( .IN1(n3411), .IN2(n3412), .QN(g8559) );
  NAND2X0 U3469 ( .IN1(n3413), .IN2(g1878), .QN(n3412) );
  NOR2X0 U3470 ( .IN1(n2990), .IN2(n3414), .QN(n3411) );
  NOR2X0 U3471 ( .IN1(n3415), .IN2(n2967), .QN(g8505) );
  XOR2X1 U3472 ( .IN1(n3416), .IN2(n1645), .Q(n3415) );
  NAND2X0 U3473 ( .IN1(n3417), .IN2(n3418), .QN(n3416) );
  NAND2X0 U3474 ( .IN1(n3419), .IN2(n3420), .QN(n3418) );
  INVX0 U3475 ( .INP(n3390), .ZN(n3420) );
  NAND2X0 U3476 ( .IN1(n3292), .IN2(n1645), .QN(n3390) );
  NOR2X0 U3477 ( .IN1(n1607), .IN2(g605), .QN(n3292) );
  NOR2X0 U3478 ( .IN1(n2973), .IN2(n3388), .QN(n3419) );
  NAND2X0 U3479 ( .IN1(n3372), .IN2(g736), .QN(n3417) );
  NAND2X0 U3480 ( .IN1(n3421), .IN2(n3422), .QN(g8435) );
  NAND2X0 U3481 ( .IN1(n3423), .IN2(g736), .QN(n3422) );
  NAND2X0 U3482 ( .IN1(n3372), .IN2(g727), .QN(n3421) );
  NAND2X0 U3483 ( .IN1(n3424), .IN2(n3425), .QN(g8434) );
  NAND2X0 U3484 ( .IN1(n3423), .IN2(g727), .QN(n3425) );
  NAND2X0 U3485 ( .IN1(n3372), .IN2(g718), .QN(n3424) );
  NAND2X0 U3486 ( .IN1(n3426), .IN2(n3427), .QN(g8433) );
  NAND2X0 U3487 ( .IN1(n3423), .IN2(g718), .QN(n3427) );
  NAND2X0 U3488 ( .IN1(n3372), .IN2(g709), .QN(n3426) );
  NAND2X0 U3489 ( .IN1(n3428), .IN2(n3429), .QN(g8432) );
  NAND2X0 U3490 ( .IN1(n3423), .IN2(g709), .QN(n3429) );
  NAND2X0 U3491 ( .IN1(n3372), .IN2(g700), .QN(n3428) );
  NAND2X0 U3492 ( .IN1(n3430), .IN2(n3431), .QN(g8431) );
  NAND2X0 U3493 ( .IN1(n3423), .IN2(g700), .QN(n3431) );
  NAND2X0 U3494 ( .IN1(n3372), .IN2(g691), .QN(n3430) );
  NAND2X0 U3495 ( .IN1(n3432), .IN2(n3433), .QN(g8430) );
  NAND2X0 U3496 ( .IN1(n3423), .IN2(g691), .QN(n3433) );
  NAND2X0 U3497 ( .IN1(n3372), .IN2(g682), .QN(n3432) );
  NAND2X0 U3498 ( .IN1(n3434), .IN2(n3435), .QN(g8429) );
  NAND2X0 U3499 ( .IN1(n3423), .IN2(g682), .QN(n3435) );
  NAND2X0 U3500 ( .IN1(n3372), .IN2(g673), .QN(n3434) );
  NAND2X0 U3501 ( .IN1(n3436), .IN2(n3437), .QN(g8428) );
  NAND2X0 U3502 ( .IN1(n3423), .IN2(g673), .QN(n3437) );
  NOR2X0 U3503 ( .IN1(n3372), .IN2(n3028), .QN(n3423) );
  NAND2X0 U3504 ( .IN1(n3372), .IN2(g664), .QN(n3436) );
  INVX0 U3505 ( .INP(n1016), .ZN(n3372) );
  NAND2X0 U3506 ( .IN1(n3438), .IN2(n1609), .QN(n1016) );
  NOR2X0 U3507 ( .IN1(n1645), .IN2(n2973), .QN(n3438) );
  NOR2X0 U3508 ( .IN1(n3439), .IN2(n2967), .QN(g8384) );
  XNOR2X1 U3509 ( .IN1(n2695), .IN2(n3440), .Q(n3439) );
  NOR2X0 U3510 ( .IN1(n3414), .IN2(n929), .QN(n3440) );
  AND2X1 U3511 ( .IN1(n3441), .IN2(n1643), .Q(n929) );
  NOR2X0 U3512 ( .IN1(n346), .IN2(n3442), .QN(n3441) );
  NOR2X0 U3513 ( .IN1(n3413), .IN2(n2696), .QN(n3414) );
  NAND2X0 U3514 ( .IN1(n1665), .IN2(n3443), .QN(g8352) );
  NAND2X0 U3515 ( .IN1(n1669), .IN2(n3443), .QN(g8349) );
  NAND2X0 U3516 ( .IN1(n1671), .IN2(n3443), .QN(g8347) );
  NAND2X0 U3517 ( .IN1(n2756), .IN2(n3443), .QN(g8340) );
  NAND2X0 U3518 ( .IN1(n1666), .IN2(n3443), .QN(g8335) );
  NAND2X0 U3519 ( .IN1(n1672), .IN2(n3443), .QN(g8331) );
  NAND2X0 U3520 ( .IN1(n1664), .IN2(n3443), .QN(g8328) );
  NAND2X0 U3521 ( .IN1(n1673), .IN2(n3443), .QN(g8323) );
  NAND2X0 U3522 ( .IN1(n1667), .IN2(n3443), .QN(g8318) );
  NAND2X0 U3523 ( .IN1(n1674), .IN2(n3443), .QN(g8316) );
  NAND2X0 U3524 ( .IN1(n1668), .IN2(n3443), .QN(g8313) );
  INVX0 U3525 ( .INP(g82), .ZN(n3443) );
  NAND2X0 U3526 ( .IN1(n3444), .IN2(n3445), .QN(g8288) );
  NAND2X0 U3527 ( .IN1(n3446), .IN2(g1950), .QN(n3445) );
  NAND2X0 U3528 ( .IN1(n3447), .IN2(g1941), .QN(n3444) );
  NAND2X0 U3529 ( .IN1(n3448), .IN2(n3449), .QN(g8287) );
  NAND2X0 U3530 ( .IN1(n3446), .IN2(g1941), .QN(n3449) );
  NAND2X0 U3531 ( .IN1(n3447), .IN2(g1932), .QN(n3448) );
  NAND2X0 U3532 ( .IN1(n3450), .IN2(n3451), .QN(g8286) );
  NAND2X0 U3533 ( .IN1(n3446), .IN2(g1932), .QN(n3451) );
  NAND2X0 U3534 ( .IN1(n3447), .IN2(g1923), .QN(n3450) );
  NAND2X0 U3535 ( .IN1(n3452), .IN2(n3453), .QN(g8285) );
  NAND2X0 U3536 ( .IN1(n3446), .IN2(g1923), .QN(n3453) );
  NAND2X0 U3537 ( .IN1(n3447), .IN2(g1914), .QN(n3452) );
  NAND2X0 U3538 ( .IN1(n3454), .IN2(n3455), .QN(g8284) );
  NAND2X0 U3539 ( .IN1(n3446), .IN2(g1914), .QN(n3455) );
  NAND2X0 U3540 ( .IN1(n3447), .IN2(g1905), .QN(n3454) );
  NAND2X0 U3541 ( .IN1(n3456), .IN2(n3457), .QN(g8283) );
  NAND2X0 U3542 ( .IN1(n3446), .IN2(g1905), .QN(n3457) );
  NAND2X0 U3543 ( .IN1(n3447), .IN2(g1896), .QN(n3456) );
  NAND2X0 U3544 ( .IN1(n3458), .IN2(n3459), .QN(g8282) );
  NAND2X0 U3545 ( .IN1(n3446), .IN2(g1896), .QN(n3459) );
  NAND2X0 U3546 ( .IN1(n3447), .IN2(g1887), .QN(n3458) );
  NAND2X0 U3547 ( .IN1(n3460), .IN2(n3461), .QN(g8281) );
  NAND2X0 U3548 ( .IN1(n3446), .IN2(g1887), .QN(n3461) );
  NOR2X0 U3549 ( .IN1(n3447), .IN2(n2990), .QN(n3446) );
  NAND2X0 U3550 ( .IN1(n3447), .IN2(g1878), .QN(n3460) );
  INVX0 U3551 ( .INP(n3413), .ZN(n3447) );
  NAND2X0 U3552 ( .IN1(n3227), .IN2(n1655), .QN(n3413) );
  NOR2X0 U3553 ( .IN1(n346), .IN2(n2695), .QN(n3227) );
  NOR2X0 U3554 ( .IN1(n1712), .IN2(n3462), .QN(g8260) );
  NOR2X0 U3555 ( .IN1(n1630), .IN2(n3462), .QN(g8254) );
  NOR2X0 U3556 ( .IN1(n1591), .IN2(n3462), .QN(g8250) );
  NOR2X0 U3557 ( .IN1(n3463), .IN2(n3464), .QN(g8245) );
  XOR2X1 U3558 ( .IN1(n1716), .IN2(n3465), .Q(n3464) );
  NOR2X0 U3559 ( .IN1(n2740), .IN2(n3466), .QN(n3465) );
  INVX0 U3560 ( .INP(n1090), .ZN(n3466) );
  NOR2X0 U3561 ( .IN1(n3467), .IN2(n3468), .QN(g8244) );
  NAND2X0 U3562 ( .IN1(n3469), .IN2(n3470), .QN(n3468) );
  NAND2X0 U3563 ( .IN1(n2519), .IN2(n3471), .QN(n3469) );
  NAND2X0 U3564 ( .IN1(n1093), .IN2(g4180), .QN(n3471) );
  NAND2X0 U3565 ( .IN1(n3472), .IN2(n3473), .QN(g8194) );
  NAND2X0 U3566 ( .IN1(n968), .IN2(g1512), .QN(n3473) );
  NAND2X0 U3567 ( .IN1(n3474), .IN2(n3306), .QN(n3472) );
  XOR2X1 U3568 ( .IN1(n3016), .IN2(n3475), .Q(n3474) );
  NOR2X0 U3569 ( .IN1(n3476), .IN2(n3477), .QN(n3475) );
  NAND2X0 U3570 ( .IN1(g1104), .IN2(g1110), .QN(n3477) );
  NAND2X0 U3571 ( .IN1(n3478), .IN2(n3479), .QN(g8193) );
  NAND2X0 U3572 ( .IN1(n968), .IN2(g1639), .QN(n3479) );
  NAND2X0 U3573 ( .IN1(n3480), .IN2(n3306), .QN(n3478) );
  XOR2X1 U3574 ( .IN1(test_so4), .IN2(n3481), .Q(n3480) );
  NOR2X0 U3575 ( .IN1(n3332), .IN2(n3476), .QN(n3481) );
  NAND2X0 U3576 ( .IN1(n1654), .IN2(n1614), .QN(n3476) );
  NAND2X0 U3577 ( .IN1(n1677), .IN2(g1104), .QN(n3332) );
  NOR2X0 U3578 ( .IN1(n3482), .IN2(g1713), .QN(g8173) );
  NOR2X0 U3579 ( .IN1(n3483), .IN2(n3484), .QN(n3482) );
  NOR2X0 U3580 ( .IN1(n2734), .IN2(n3485), .QN(n3484) );
  NOR2X0 U3581 ( .IN1(n1055), .IN2(n1054), .QN(n3485) );
  NOR2X0 U3582 ( .IN1(n3486), .IN2(n3487), .QN(n3483) );
  NAND2X0 U3583 ( .IN1(n1055), .IN2(g1801), .QN(n3487) );
  NAND2X0 U3584 ( .IN1(n3488), .IN2(n1057), .QN(n1055) );
  NOR2X0 U3585 ( .IN1(n3489), .IN2(n1626), .QN(n1057) );
  NOR2X0 U3586 ( .IN1(n2734), .IN2(n2733), .QN(n3488) );
  INVX0 U3587 ( .INP(n1056), .ZN(n3486) );
  NOR2X0 U3588 ( .IN1(n1604), .IN2(n3462), .QN(g8147) );
  NAND2X0 U3589 ( .IN1(n3490), .IN2(g109), .QN(n3462) );
  NAND2X0 U3590 ( .IN1(n3491), .IN2(n4930), .QN(n3490) );
  NOR2X0 U3591 ( .IN1(g881), .IN2(n3492), .QN(n3491) );
  NOR2X0 U3592 ( .IN1(n2757), .IN2(n3493), .QN(g8060) );
  XOR2X1 U3593 ( .IN1(g6002), .IN2(n2649), .Q(n3493) );
  NOR2X0 U3594 ( .IN1(n2758), .IN2(n3494), .QN(g8059) );
  XOR2X1 U3595 ( .IN1(g6042), .IN2(n2646), .Q(n3494) );
  NOR2X0 U3596 ( .IN1(n2759), .IN2(n3495), .QN(g8055) );
  XOR2X1 U3597 ( .IN1(n3496), .IN2(g1490), .Q(n3495) );
  NOR2X0 U3598 ( .IN1(n2760), .IN2(n3497), .QN(g8054) );
  XOR2X1 U3599 ( .IN1(g6015), .IN2(n2741), .Q(n3497) );
  NOR2X0 U3600 ( .IN1(n2757), .IN2(n3498), .QN(g8053) );
  XOR2X1 U3601 ( .IN1(g6045), .IN2(n2645), .Q(n3498) );
  NOR2X0 U3602 ( .IN1(n2758), .IN2(n3499), .QN(g8052) );
  XOR2X1 U3603 ( .IN1(n3500), .IN2(n2647), .Q(n3499) );
  NOR2X0 U3604 ( .IN1(n2759), .IN2(n3501), .QN(g8051) );
  XNOR2X1 U3605 ( .IN1(n3502), .IN2(n2651), .Q(n3501) );
  NOR2X0 U3606 ( .IN1(n2760), .IN2(n3503), .QN(g8050) );
  XOR2X1 U3607 ( .IN1(g6026), .IN2(n2742), .Q(n3503) );
  NOR2X0 U3608 ( .IN1(n2757), .IN2(n3504), .QN(g8049) );
  XOR2X1 U3609 ( .IN1(g6049), .IN2(n2648), .Q(n3504) );
  NOR2X0 U3610 ( .IN1(n2758), .IN2(n3505), .QN(g8048) );
  XOR2X1 U3611 ( .IN1(g5996), .IN2(n2670), .Q(n3505) );
  NOR2X0 U3612 ( .IN1(n2759), .IN2(n3506), .QN(g8047) );
  XOR2X1 U3613 ( .IN1(g6035), .IN2(n1704), .Q(n3506) );
  NOR2X0 U3614 ( .IN1(n2760), .IN2(n3507), .QN(g8046) );
  XOR2X1 U3615 ( .IN1(n3508), .IN2(n2652), .Q(n3507) );
  NOR2X0 U3616 ( .IN1(n2757), .IN2(n3509), .QN(g8045) );
  XOR2X1 U3617 ( .IN1(n3510), .IN2(g1462), .Q(n3509) );
  NOR2X0 U3618 ( .IN1(n2758), .IN2(n3511), .QN(g8044) );
  XOR2X1 U3619 ( .IN1(g6038), .IN2(n2644), .Q(n3511) );
  NOR2X0 U3620 ( .IN1(n2759), .IN2(n3512), .QN(g8043) );
  XOR2X1 U3621 ( .IN1(n3513), .IN2(n2725), .Q(n3512) );
  NOR2X0 U3622 ( .IN1(n2760), .IN2(n3514), .QN(g8042) );
  XNOR2X1 U3623 ( .IN1(n3515), .IN2(n1703), .Q(n3514) );
  NOR2X0 U3624 ( .IN1(n2757), .IN2(n3516), .QN(g8041) );
  XOR2X1 U3625 ( .IN1(n3517), .IN2(n2687), .Q(n3516) );
  NOR2X0 U3626 ( .IN1(n2758), .IN2(n3518), .QN(g8040) );
  XOR2X1 U3627 ( .IN1(g1474), .IN2(n3519), .Q(n3518) );
  NOR2X0 U3628 ( .IN1(n2759), .IN2(n3520), .QN(g8039) );
  XOR2X1 U3629 ( .IN1(g1470), .IN2(n3521), .Q(n3520) );
  NOR2X0 U3630 ( .IN1(n3463), .IN2(n3522), .QN(g8024) );
  XOR2X1 U3631 ( .IN1(n2740), .IN2(n1090), .Q(n3522) );
  NOR2X0 U3632 ( .IN1(n3467), .IN2(n3523), .QN(g8019) );
  XOR2X1 U3633 ( .IN1(n2524), .IN2(n1093), .Q(n3523) );
  NOR2X0 U3634 ( .IN1(g1713), .IN2(n3524), .QN(g7930) );
  XOR2X1 U3635 ( .IN1(n2733), .IN2(n1056), .Q(n3524) );
  NOR2X0 U3636 ( .IN1(n2760), .IN2(n3525), .QN(g7843) );
  XOR2X1 U3637 ( .IN1(g6000), .IN2(n2650), .Q(n3525) );
  NOR2X0 U3638 ( .IN1(n3463), .IN2(n3526), .QN(g7709) );
  OR2X1 U3639 ( .IN1(n1096), .IN2(n1090), .Q(n3526) );
  NOR2X0 U3640 ( .IN1(n3467), .IN2(n3527), .QN(g7705) );
  OR2X1 U3641 ( .IN1(n1098), .IN2(n1093), .Q(n3527) );
  NAND2X0 U3642 ( .IN1(n3528), .IN2(n3529), .QN(g7660) );
  OR2X1 U3643 ( .IN1(n3530), .IN2(n2729), .Q(n3529) );
  NOR2X0 U3644 ( .IN1(n3286), .IN2(n3028), .QN(n3528) );
  INVX0 U3645 ( .INP(n3300), .ZN(n3028) );
  NOR2X0 U3646 ( .IN1(n3531), .IN2(n3532), .QN(g7632) );
  XNOR2X1 U3647 ( .IN1(n2508), .IN2(n3533), .Q(n3532) );
  NAND2X0 U3648 ( .IN1(n3534), .IN2(n3300), .QN(g7626) );
  NOR2X0 U3649 ( .IN1(n3535), .IN2(n3536), .QN(n3534) );
  NOR2X0 U3650 ( .IN1(g639), .IN2(n3537), .QN(n3536) );
  NAND2X0 U3651 ( .IN1(n3286), .IN2(n3538), .QN(n3537) );
  NAND2X0 U3652 ( .IN1(n3539), .IN2(n2946), .QN(n3538) );
  INVX0 U3653 ( .INP(n3296), .ZN(n2946) );
  NAND2X0 U3654 ( .IN1(n3283), .IN2(n3540), .QN(n3296) );
  NAND2X0 U3655 ( .IN1(n1593), .IN2(g599), .QN(n3540) );
  NAND2X0 U3656 ( .IN1(n3541), .IN2(n1644), .QN(n3283) );
  NOR2X0 U3657 ( .IN1(n1593), .IN2(g591), .QN(n3541) );
  NOR2X0 U3658 ( .IN1(n3072), .IN2(n3285), .QN(n3539) );
  INVX0 U3659 ( .INP(n3070), .ZN(n3285) );
  NAND2X0 U3660 ( .IN1(n1607), .IN2(g599), .QN(n3070) );
  INVX0 U3661 ( .INP(n3060), .ZN(n3072) );
  NAND2X0 U3662 ( .IN1(g605), .IN2(g591), .QN(n3060) );
  NOR2X0 U3663 ( .IN1(n1692), .IN2(n3286), .QN(n3535) );
  INVX0 U3664 ( .INP(n2973), .ZN(n3286) );
  NOR2X0 U3665 ( .IN1(n3542), .IN2(n3531), .QN(g7590) );
  NOR2X0 U3666 ( .IN1(n3543), .IN2(g1231), .QN(n3542) );
  NOR2X0 U3667 ( .IN1(n3544), .IN2(n3531), .QN(g7586) );
  NOR2X0 U3668 ( .IN1(n3545), .IN2(n1107), .QN(n3544) );
  AND2X1 U3669 ( .IN1(n3546), .IN2(n3547), .Q(n1107) );
  NOR2X0 U3670 ( .IN1(n2509), .IN2(n2508), .QN(n3547) );
  NOR2X0 U3671 ( .IN1(n3548), .IN2(n3533), .QN(n3546) );
  NOR2X0 U3672 ( .IN1(n2507), .IN2(n3543), .QN(n3545) );
  NOR2X0 U3673 ( .IN1(n3549), .IN2(n3533), .QN(n3543) );
  INVX0 U3674 ( .INP(n3548), .ZN(n3549) );
  NOR2X0 U3675 ( .IN1(n3531), .IN2(n3550), .QN(g7581) );
  XOR2X1 U3676 ( .IN1(n2509), .IN2(n3551), .Q(n3550) );
  NOR2X0 U3677 ( .IN1(n2508), .IN2(n3533), .QN(n3551) );
  NAND2X0 U3678 ( .IN1(n3552), .IN2(n3553), .QN(n3533) );
  NAND2X0 U3679 ( .IN1(n2743), .IN2(g109), .QN(n3531) );
  NOR2X0 U3680 ( .IN1(g1713), .IN2(n3554), .QN(g7541) );
  NAND2X0 U3681 ( .IN1(n3555), .IN2(n3556), .QN(n3554) );
  NAND2X0 U3682 ( .IN1(n1056), .IN2(g1796), .QN(n3556) );
  OR2X1 U3683 ( .IN1(g1796), .IN2(n1116), .Q(n3555) );
  NAND2X0 U3684 ( .IN1(n3557), .IN2(n3300), .QN(g7441) );
  XOR2X1 U3685 ( .IN1(g643), .IN2(n1701), .Q(n3557) );
  NAND2X0 U3686 ( .IN1(n3558), .IN2(n3559), .QN(g7303) );
  NAND2X0 U3687 ( .IN1(n3560), .IN2(test_so6), .QN(n3559) );
  NAND2X0 U3688 ( .IN1(n3552), .IN2(g1265), .QN(n3558) );
  NAND2X0 U3689 ( .IN1(n3561), .IN2(n3562), .QN(g7302) );
  NAND2X0 U3690 ( .IN1(n3560), .IN2(g1265), .QN(n3562) );
  NAND2X0 U3691 ( .IN1(n3552), .IN2(g1260), .QN(n3561) );
  NAND2X0 U3692 ( .IN1(n3563), .IN2(n3564), .QN(g7301) );
  NAND2X0 U3693 ( .IN1(n3560), .IN2(g1260), .QN(n3564) );
  NAND2X0 U3694 ( .IN1(n3552), .IN2(g1255), .QN(n3563) );
  NAND2X0 U3695 ( .IN1(n3565), .IN2(n3566), .QN(g7300) );
  NAND2X0 U3696 ( .IN1(n3560), .IN2(g1255), .QN(n3566) );
  NAND2X0 U3697 ( .IN1(n3552), .IN2(g1250), .QN(n3565) );
  NAND2X0 U3698 ( .IN1(n3567), .IN2(n3568), .QN(g7299) );
  NAND2X0 U3699 ( .IN1(n3560), .IN2(g1250), .QN(n3568) );
  NAND2X0 U3700 ( .IN1(n3552), .IN2(g1245), .QN(n3567) );
  NAND2X0 U3701 ( .IN1(n3569), .IN2(n3570), .QN(g7298) );
  NAND2X0 U3702 ( .IN1(n3560), .IN2(g1245), .QN(n3570) );
  NAND2X0 U3703 ( .IN1(n3552), .IN2(g1240), .QN(n3569) );
  NAND2X0 U3704 ( .IN1(n3571), .IN2(n3572), .QN(g7297) );
  NAND2X0 U3705 ( .IN1(n3560), .IN2(g1240), .QN(n3572) );
  NAND2X0 U3706 ( .IN1(n3552), .IN2(g1235), .QN(n3571) );
  NAND2X0 U3707 ( .IN1(n3573), .IN2(n3574), .QN(g7296) );
  NAND2X0 U3708 ( .IN1(n3560), .IN2(g1235), .QN(n3574) );
  NAND2X0 U3709 ( .IN1(n3552), .IN2(g1275), .QN(n3573) );
  NAND2X0 U3710 ( .IN1(n3575), .IN2(n3576), .QN(g7295) );
  NAND2X0 U3711 ( .IN1(n3560), .IN2(g1280), .QN(n3576) );
  NAND2X0 U3712 ( .IN1(n3552), .IN2(g1284), .QN(n3575) );
  NAND2X0 U3713 ( .IN1(n3577), .IN2(n3578), .QN(g7294) );
  NAND2X0 U3714 ( .IN1(n3560), .IN2(g1284), .QN(n3578) );
  NAND2X0 U3715 ( .IN1(n3552), .IN2(g1292), .QN(n3577) );
  NAND2X0 U3716 ( .IN1(n3579), .IN2(n3580), .QN(g7293) );
  NAND2X0 U3717 ( .IN1(n3560), .IN2(g1292), .QN(n3580) );
  NAND2X0 U3718 ( .IN1(n3552), .IN2(g1296), .QN(n3579) );
  NAND2X0 U3719 ( .IN1(n3581), .IN2(n3582), .QN(g7292) );
  NAND2X0 U3720 ( .IN1(n3560), .IN2(g1296), .QN(n3582) );
  NAND2X0 U3721 ( .IN1(n3552), .IN2(g1300), .QN(n3581) );
  NAND2X0 U3722 ( .IN1(n3583), .IN2(n3584), .QN(g7291) );
  NAND2X0 U3723 ( .IN1(n3560), .IN2(g1300), .QN(n3584) );
  NAND2X0 U3724 ( .IN1(n3552), .IN2(g1304), .QN(n3583) );
  NAND2X0 U3725 ( .IN1(n3585), .IN2(n3586), .QN(g7290) );
  NAND2X0 U3726 ( .IN1(n3560), .IN2(g1304), .QN(n3586) );
  NAND2X0 U3727 ( .IN1(n3552), .IN2(test_so6), .QN(n3585) );
  NAND2X0 U3728 ( .IN1(n3587), .IN2(n3588), .QN(g7257) );
  NAND2X0 U3729 ( .IN1(n3306), .IN2(g1077), .QN(n3588) );
  NAND2X0 U3730 ( .IN1(n968), .IN2(g1032), .QN(n3587) );
  NAND2X0 U3731 ( .IN1(n3589), .IN2(n3590), .QN(g7244) );
  NAND2X0 U3732 ( .IN1(n3306), .IN2(g1071), .QN(n3590) );
  OR2X1 U3733 ( .IN1(n3306), .IN2(n2593), .Q(n3589) );
  NAND2X0 U3734 ( .IN1(n2756), .IN2(n3591), .QN(g7219) );
  NAND2X0 U3735 ( .IN1(n1672), .IN2(n3591), .QN(g7204) );
  NOR2X0 U3736 ( .IN1(n3463), .IN2(n3592), .QN(g7202) );
  XOR2X1 U3737 ( .IN1(n2738), .IN2(n1123), .Q(n3592) );
  NOR2X0 U3738 ( .IN1(n3467), .IN2(n3593), .QN(g7191) );
  XOR2X1 U3739 ( .IN1(n2523), .IN2(n1125), .Q(n3593) );
  NAND2X0 U3740 ( .IN1(n1673), .IN2(n3591), .QN(g7189) );
  NAND2X0 U3741 ( .IN1(n1674), .IN2(n3591), .QN(g7183) );
  NAND2X0 U3742 ( .IN1(n1671), .IN2(n3591), .QN(g7143) );
  NOR2X0 U3743 ( .IN1(n3594), .IN2(n3595), .QN(g7137) );
  NOR2X0 U3744 ( .IN1(n3596), .IN2(n3530), .QN(n3594) );
  NOR2X0 U3745 ( .IN1(n1709), .IN2(n3597), .QN(n3596) );
  NOR2X0 U3746 ( .IN1(n3598), .IN2(n3595), .QN(g7134) );
  NAND2X0 U3747 ( .IN1(n3300), .IN2(n2973), .QN(n3595) );
  NAND2X0 U3748 ( .IN1(n2729), .IN2(n3530), .QN(n2973) );
  AND2X1 U3749 ( .IN1(n1709), .IN2(n3597), .Q(n3530) );
  NOR2X0 U3750 ( .IN1(n3599), .IN2(n3597), .QN(n3598) );
  AND2X1 U3751 ( .IN1(n3600), .IN2(n4940), .Q(n3597) );
  NOR2X0 U3752 ( .IN1(n4940), .IN2(n3600), .QN(n3599) );
  NOR2X0 U3753 ( .IN1(n1701), .IN2(g643), .QN(n3600) );
  NAND2X0 U3754 ( .IN1(n1610), .IN2(n3601), .QN(g7133) );
  XOR2X1 U3755 ( .IN1(g1766), .IN2(n1054), .Q(n3601) );
  NAND2X0 U3756 ( .IN1(n3602), .IN2(n3603), .QN(g7032) );
  OR2X1 U3757 ( .IN1(n2758), .IN2(n2488), .Q(n3603) );
  INVX0 U3758 ( .INP(n1132), .ZN(n3602) );
  NOR2X0 U3759 ( .IN1(n3604), .IN2(n3605), .QN(n1132) );
  NAND2X0 U3760 ( .IN1(n3606), .IN2(n3607), .QN(n3605) );
  NOR2X0 U3761 ( .IN1(n3608), .IN2(n3609), .QN(n3607) );
  NAND2X0 U3762 ( .IN1(n2649), .IN2(n2646), .QN(n3609) );
  NAND2X0 U3763 ( .IN1(n2645), .IN2(n2644), .QN(n3608) );
  NOR2X0 U3764 ( .IN1(n3610), .IN2(n3611), .QN(n3606) );
  NAND2X0 U3765 ( .IN1(n2672), .IN2(n2671), .QN(n3611) );
  NAND2X0 U3766 ( .IN1(n2670), .IN2(n2650), .QN(n3610) );
  NAND2X0 U3767 ( .IN1(n3612), .IN2(n3613), .QN(n3604) );
  NOR2X0 U3768 ( .IN1(n3614), .IN2(n3615), .QN(n3613) );
  NAND2X0 U3769 ( .IN1(g166), .IN2(g182), .QN(n3615) );
  NAND2X0 U3770 ( .IN1(g174), .IN2(g170), .QN(n3614) );
  NOR2X0 U3771 ( .IN1(n3616), .IN2(n3617), .QN(n3612) );
  NAND2X0 U3772 ( .IN1(n1704), .IN2(n1613), .QN(n3617) );
  NAND2X0 U3773 ( .IN1(g6786), .IN2(n1137), .QN(n3616) );
  NOR2X0 U3774 ( .IN1(n3618), .IN2(g1713), .QN(g6983) );
  NOR2X0 U3775 ( .IN1(n3619), .IN2(n3620), .QN(n3618) );
  NOR2X0 U3776 ( .IN1(n1702), .IN2(n1116), .QN(n3620) );
  NOR2X0 U3777 ( .IN1(n3489), .IN2(n1054), .QN(n1116) );
  NOR2X0 U3778 ( .IN1(n2938), .IN2(n3621), .QN(n3619) );
  NAND2X0 U3779 ( .IN1(n3489), .IN2(g1786), .QN(n3621) );
  NAND2X0 U3780 ( .IN1(n3622), .IN2(n3623), .QN(n3489) );
  NOR2X0 U3781 ( .IN1(n2735), .IN2(n1702), .QN(n3623) );
  NOR2X0 U3782 ( .IN1(n1659), .IN2(n3624), .QN(n3622) );
  NAND2X0 U3783 ( .IN1(n3625), .IN2(n3626), .QN(g6934) );
  OR2X1 U3784 ( .IN1(n3627), .IN2(n2565), .Q(n3626) );
  NAND2X0 U3785 ( .IN1(n3627), .IN2(g170), .QN(n3625) );
  NAND2X0 U3786 ( .IN1(n3628), .IN2(n3629), .QN(g6930) );
  NAND2X0 U3787 ( .IN1(n3306), .IN2(g1074), .QN(n3629) );
  OR2X1 U3788 ( .IN1(n3306), .IN2(n2618), .Q(n3628) );
  NAND2X0 U3789 ( .IN1(n3630), .IN2(n3631), .QN(g6929) );
  NAND2X0 U3790 ( .IN1(n3632), .IN2(g302), .QN(n3631) );
  OR2X1 U3791 ( .IN1(n3632), .IN2(n2671), .Q(n3630) );
  NAND2X0 U3792 ( .IN1(n3633), .IN2(n3634), .QN(g6928) );
  OR2X1 U3793 ( .IN1(n3627), .IN2(n2564), .Q(n3634) );
  NAND2X0 U3794 ( .IN1(n3627), .IN2(g174), .QN(n3633) );
  NAND2X0 U3795 ( .IN1(n3635), .IN2(n3636), .QN(g6924) );
  NAND2X0 U3796 ( .IN1(n3306), .IN2(g1098), .QN(n3636) );
  OR2X1 U3797 ( .IN1(n3306), .IN2(n2619), .Q(n3635) );
  NAND2X0 U3798 ( .IN1(n3637), .IN2(n3638), .QN(g6923) );
  NAND2X0 U3799 ( .IN1(n3632), .IN2(g299), .QN(n3638) );
  NAND2X0 U3800 ( .IN1(n3627), .IN2(g166), .QN(n3637) );
  NAND2X0 U3801 ( .IN1(n3639), .IN2(n3640), .QN(g6922) );
  NAND2X0 U3802 ( .IN1(n3632), .IN2(g278), .QN(n3640) );
  OR2X1 U3803 ( .IN1(n3632), .IN2(n2649), .Q(n3639) );
  NAND2X0 U3804 ( .IN1(n3641), .IN2(n3642), .QN(g6918) );
  NAND2X0 U3805 ( .IN1(n3306), .IN2(g1095), .QN(n3642) );
  NAND2X0 U3806 ( .IN1(test_so2), .IN2(n968), .QN(n3641) );
  NAND2X0 U3807 ( .IN1(n3643), .IN2(n3644), .QN(g6916) );
  NAND2X0 U3808 ( .IN1(n3632), .IN2(g296), .QN(n3644) );
  OR2X1 U3809 ( .IN1(n3632), .IN2(n2645), .Q(n3643) );
  NAND2X0 U3810 ( .IN1(n3645), .IN2(n3646), .QN(g6915) );
  NAND2X0 U3811 ( .IN1(n3632), .IN2(g275), .QN(n3646) );
  OR2X1 U3812 ( .IN1(n3632), .IN2(n2650), .Q(n3645) );
  NAND2X0 U3813 ( .IN1(n3647), .IN2(n3648), .QN(g6912) );
  NAND2X0 U3814 ( .IN1(n3306), .IN2(g1092), .QN(n3648) );
  OR2X1 U3815 ( .IN1(n3306), .IN2(n2658), .Q(n3647) );
  NAND2X0 U3816 ( .IN1(n3649), .IN2(n3650), .QN(g6911) );
  NAND2X0 U3817 ( .IN1(n3632), .IN2(g293), .QN(n3650) );
  OR2X1 U3818 ( .IN1(n3632), .IN2(n2646), .Q(n3649) );
  NAND2X0 U3819 ( .IN1(n3651), .IN2(n3652), .QN(g6910) );
  OR2X1 U3820 ( .IN1(n3627), .IN2(n2557), .Q(n3652) );
  OR2X1 U3821 ( .IN1(n3632), .IN2(n2670), .Q(n3651) );
  NAND2X0 U3822 ( .IN1(n3653), .IN2(n3654), .QN(g6909) );
  NAND2X0 U3823 ( .IN1(n3655), .IN2(g1868), .QN(n3654) );
  INVX0 U3824 ( .INP(n3656), .ZN(n3653) );
  NAND2X0 U3825 ( .IN1(n3657), .IN2(n3658), .QN(g6908) );
  NAND2X0 U3826 ( .IN1(n3306), .IN2(g1089), .QN(n3658) );
  NAND2X0 U3827 ( .IN1(test_so8), .IN2(n968), .QN(n3657) );
  NAND2X0 U3828 ( .IN1(n3659), .IN2(n3660), .QN(g6907) );
  NAND2X0 U3829 ( .IN1(n3632), .IN2(g290), .QN(n3660) );
  OR2X1 U3830 ( .IN1(n3632), .IN2(n2644), .Q(n3659) );
  NAND2X0 U3831 ( .IN1(n3661), .IN2(n3662), .QN(g6906) );
  OR2X1 U3832 ( .IN1(n3627), .IN2(n2563), .Q(n3662) );
  OR2X1 U3833 ( .IN1(n3632), .IN2(n2672), .Q(n3661) );
  NAND2X0 U3834 ( .IN1(n3663), .IN2(n3664), .QN(g6902) );
  NAND2X0 U3835 ( .IN1(n3306), .IN2(g1086), .QN(n3664) );
  NAND2X0 U3836 ( .IN1(n968), .IN2(g1003), .QN(n3663) );
  NAND2X0 U3837 ( .IN1(n3665), .IN2(n3666), .QN(g6901) );
  NAND2X0 U3838 ( .IN1(n3632), .IN2(g287), .QN(n3666) );
  OR2X1 U3839 ( .IN1(n3632), .IN2(n1704), .Q(n3665) );
  NAND2X0 U3840 ( .IN1(n3667), .IN2(n3668), .QN(g6900) );
  OR2X1 U3841 ( .IN1(n3627), .IN2(n2554), .Q(n3668) );
  NAND2X0 U3842 ( .IN1(n3627), .IN2(g178), .QN(n3667) );
  NAND2X0 U3843 ( .IN1(n3669), .IN2(n3670), .QN(g6898) );
  NAND2X0 U3844 ( .IN1(n3306), .IN2(g1083), .QN(n3670) );
  OR2X1 U3845 ( .IN1(n3306), .IN2(n1871), .Q(n3669) );
  NAND2X0 U3846 ( .IN1(n3671), .IN2(n3672), .QN(g6897) );
  NAND2X0 U3847 ( .IN1(n3632), .IN2(g263), .QN(n3672) );
  INVX0 U3848 ( .INP(n3627), .ZN(n3632) );
  NAND2X0 U3849 ( .IN1(n3627), .IN2(g182), .QN(n3671) );
  NAND2X0 U3850 ( .IN1(n3673), .IN2(g109), .QN(n3627) );
  NAND2X0 U3851 ( .IN1(n1613), .IN2(n1137), .QN(n3673) );
  NOR2X0 U3852 ( .IN1(n2967), .IN2(n4944), .QN(n1137) );
  NAND2X0 U3853 ( .IN1(n3674), .IN2(n3675), .QN(g6895) );
  NAND2X0 U3854 ( .IN1(n3306), .IN2(g1080), .QN(n3675) );
  OR2X1 U3855 ( .IN1(n3306), .IN2(n2698), .Q(n3674) );
  NAND2X0 U3856 ( .IN1(n3676), .IN2(n3677), .QN(g6894) );
  NAND2X0 U3857 ( .IN1(test_so7), .IN2(n3306), .QN(n3677) );
  NAND2X0 U3858 ( .IN1(n968), .IN2(g1027), .QN(n3676) );
  NOR2X0 U3859 ( .IN1(g1696), .IN2(g4089), .QN(g6842) );
  NOR2X0 U3860 ( .IN1(n1629), .IN2(n2757), .QN(g6841) );
  NOR2X0 U3861 ( .IN1(n1598), .IN2(n2757), .QN(g6840) );
  NOR2X0 U3862 ( .IN1(n1711), .IN2(n2758), .QN(g6839) );
  NOR2X0 U3863 ( .IN1(n4942), .IN2(n2759), .QN(g6834) );
  NOR2X0 U3864 ( .IN1(n4945), .IN2(n2760), .QN(g6830) );
  NOR2X0 U3865 ( .IN1(n4943), .IN2(n2757), .QN(g6828) );
  NOR2X0 U3866 ( .IN1(n4941), .IN2(n2758), .QN(g6820) );
  NOR2X0 U3867 ( .IN1(n3678), .IN2(n3656), .QN(g6795) );
  NOR2X0 U3868 ( .IN1(n3679), .IN2(n34), .QN(n3678) );
  INVX0 U3869 ( .INP(n3655), .ZN(n34) );
  NAND2X0 U3870 ( .IN1(n2730), .IN2(n3680), .QN(n3655) );
  NOR2X0 U3871 ( .IN1(n2730), .IN2(n3680), .QN(n3679) );
  NAND2X0 U3872 ( .IN1(n4946), .IN2(n3681), .QN(g6755) );
  NOR2X0 U3873 ( .IN1(n3022), .IN2(n3682), .QN(g6747) );
  NAND2X0 U3874 ( .IN1(n3683), .IN2(g109), .QN(n3682) );
  NAND2X0 U3875 ( .IN1(n4931), .IN2(n4948), .QN(n3683) );
  NOR2X0 U3876 ( .IN1(n3463), .IN2(n3684), .QN(g6733) );
  OR2X1 U3877 ( .IN1(n1150), .IN2(n1123), .Q(n3684) );
  NOR2X0 U3878 ( .IN1(n3467), .IN2(n3685), .QN(g6728) );
  OR2X1 U3879 ( .IN1(n1152), .IN2(n1125), .Q(n3685) );
  NAND2X0 U3880 ( .IN1(n3686), .IN2(n3687), .QN(g6679) );
  NAND2X0 U3881 ( .IN1(n1155), .IN2(n1154), .QN(n3687) );
  AND2X1 U3882 ( .IN1(n3688), .IN2(n3689), .Q(n1154) );
  NOR2X0 U3883 ( .IN1(n3690), .IN2(n3691), .QN(n3689) );
  NAND2X0 U3884 ( .IN1(g1515), .IN2(g1520), .QN(n3691) );
  NAND2X0 U3885 ( .IN1(g1448), .IN2(g1432), .QN(n3690) );
  AND2X1 U3886 ( .IN1(n3692), .IN2(g6234), .Q(n3688) );
  NOR2X0 U3887 ( .IN1(n1602), .IN2(n3693), .QN(n3692) );
  AND2X1 U3888 ( .IN1(n3694), .IN2(n3695), .Q(n1155) );
  NOR2X0 U3889 ( .IN1(n3696), .IN2(n3697), .QN(n3695) );
  NAND2X0 U3890 ( .IN1(g1436), .IN2(g1440), .QN(n3697) );
  NAND2X0 U3891 ( .IN1(g1428), .IN2(g1444), .QN(n3696) );
  NOR2X0 U3892 ( .IN1(n3698), .IN2(n3699), .QN(n3694) );
  NAND2X0 U3893 ( .IN1(n2655), .IN2(n2550), .QN(n3699) );
  NAND2X0 U3894 ( .IN1(n2532), .IN2(n2527), .QN(n3698) );
  NAND2X0 U3895 ( .IN1(g109), .IN2(g1), .QN(n3686) );
  NAND2X0 U3896 ( .IN1(n1701), .IN2(n3700), .QN(g6672) );
  NAND2X0 U3897 ( .IN1(n3701), .IN2(n3702), .QN(g6656) );
  NAND2X0 U3898 ( .IN1(n1162), .IN2(n1161), .QN(n3702) );
  AND2X1 U3899 ( .IN1(n3703), .IN2(n3704), .Q(n1161) );
  NOR2X0 U3900 ( .IN1(n3705), .IN2(n3706), .QN(n3704) );
  NAND2X0 U3901 ( .IN1(g1508), .IN2(g1494), .QN(n3706) );
  NAND2X0 U3902 ( .IN1(g1474), .IN2(g1470), .QN(n3705) );
  NOR2X0 U3903 ( .IN1(n3693), .IN2(n3707), .QN(n3703) );
  NAND2X0 U3904 ( .IN1(n2750), .IN2(g1453), .QN(n3707) );
  NOR2X0 U3905 ( .IN1(n2757), .IN2(n2529), .QN(n2750) );
  AND2X1 U3906 ( .IN1(n3708), .IN2(n3709), .Q(n1162) );
  NOR2X0 U3907 ( .IN1(n3710), .IN2(n3711), .QN(n3709) );
  NAND2X0 U3908 ( .IN1(n1703), .IN2(g1490), .QN(n3711) );
  NAND2X0 U3909 ( .IN1(g1462), .IN2(g1478), .QN(n3710) );
  NOR2X0 U3910 ( .IN1(n3712), .IN2(n3713), .QN(n3708) );
  NAND2X0 U3911 ( .IN1(n2673), .IN2(n2652), .QN(n3713) );
  NAND2X0 U3912 ( .IN1(n2651), .IN2(n2647), .QN(n3712) );
  NAND2X0 U3913 ( .IN1(g109), .IN2(g4), .QN(n3701) );
  NOR2X0 U3914 ( .IN1(n1666), .IN2(n3714), .QN(g6653) );
  NOR2X0 U3915 ( .IN1(n1664), .IN2(n3714), .QN(g6638) );
  NOR2X0 U3916 ( .IN1(n1667), .IN2(n3714), .QN(g6627) );
  NOR2X0 U3917 ( .IN1(n1668), .IN2(n3714), .QN(g6621) );
  NAND2X0 U3918 ( .IN1(n3715), .IN2(n3716), .QN(g6551) );
  NAND2X0 U3919 ( .IN1(n3717), .IN2(g1546), .QN(n3716) );
  NAND2X0 U3920 ( .IN1(n3718), .IN2(g1478), .QN(n3715) );
  NAND2X0 U3921 ( .IN1(n3719), .IN2(n3720), .QN(g6546) );
  OR2X1 U3922 ( .IN1(n3718), .IN2(n2546), .Q(n3720) );
  NAND2X0 U3923 ( .IN1(n3718), .IN2(g1453), .QN(n3719) );
  NAND2X0 U3924 ( .IN1(n3721), .IN2(n3722), .QN(g6545) );
  OR2X1 U3925 ( .IN1(n3718), .IN2(n2548), .Q(n3722) );
  OR2X1 U3926 ( .IN1(n3717), .IN2(n2652), .Q(n3721) );
  NAND2X0 U3927 ( .IN1(n3723), .IN2(n3724), .QN(g6542) );
  NAND2X0 U3928 ( .IN1(n3717), .IN2(g1561), .QN(n3724) );
  OR2X1 U3929 ( .IN1(n3717), .IN2(n1703), .Q(n3723) );
  NAND2X0 U3930 ( .IN1(n3725), .IN2(n3726), .QN(g6541) );
  NAND2X0 U3931 ( .IN1(n3717), .IN2(g1540), .QN(n3726) );
  OR2X1 U3932 ( .IN1(n3717), .IN2(n2647), .Q(n3725) );
  NAND2X0 U3933 ( .IN1(n3727), .IN2(n3728), .QN(g6538) );
  OR2X1 U3934 ( .IN1(n3718), .IN2(n2552), .Q(n3728) );
  NAND2X0 U3935 ( .IN1(n3718), .IN2(g1462), .QN(n3727) );
  NAND2X0 U3936 ( .IN1(n3729), .IN2(n3730), .QN(g6537) );
  NAND2X0 U3937 ( .IN1(n3717), .IN2(g1537), .QN(n3730) );
  NAND2X0 U3938 ( .IN1(n3718), .IN2(g1490), .QN(n3729) );
  NAND2X0 U3939 ( .IN1(n3731), .IN2(n3732), .QN(g6534) );
  OR2X1 U3940 ( .IN1(n3718), .IN2(n2528), .Q(n3732) );
  OR2X1 U3941 ( .IN1(n3717), .IN2(n2651), .Q(n3731) );
  NAND2X0 U3942 ( .IN1(n3733), .IN2(n3734), .QN(g6533) );
  OR2X1 U3943 ( .IN1(n3718), .IN2(n1632), .Q(n3734) );
  NAND2X0 U3944 ( .IN1(n3718), .IN2(g1494), .QN(n3733) );
  NOR2X0 U3945 ( .IN1(n1665), .IN2(n3714), .QN(g6531) );
  NAND2X0 U3946 ( .IN1(n3735), .IN2(n3736), .QN(g6529) );
  OR2X1 U3947 ( .IN1(n3718), .IN2(n2533), .Q(n3736) );
  NAND2X0 U3948 ( .IN1(n3718), .IN2(g1470), .QN(n3735) );
  NAND2X0 U3949 ( .IN1(n3737), .IN2(n3738), .QN(g6528) );
  OR2X1 U3950 ( .IN1(n3718), .IN2(n1652), .Q(n3738) );
  OR2X1 U3951 ( .IN1(n3717), .IN2(n2673), .Q(n3737) );
  NOR2X0 U3952 ( .IN1(n1669), .IN2(n3714), .QN(g6526) );
  NOR2X0 U3953 ( .IN1(g1713), .IN2(n3739), .QN(g6525) );
  XOR2X1 U3954 ( .IN1(g1786), .IN2(n2938), .Q(n3739) );
  NAND2X0 U3955 ( .IN1(n3740), .IN2(n3741), .QN(g6524) );
  NAND2X0 U3956 ( .IN1(n3717), .IN2(g1589), .QN(n3741) );
  NAND2X0 U3957 ( .IN1(n3718), .IN2(g1428), .QN(n3740) );
  NAND2X0 U3958 ( .IN1(n3742), .IN2(n3743), .QN(g6523) );
  OR2X1 U3959 ( .IN1(n3718), .IN2(n2535), .Q(n3743) );
  NAND2X0 U3960 ( .IN1(n3718), .IN2(g1474), .QN(n3742) );
  NAND2X0 U3961 ( .IN1(n3744), .IN2(n3745), .QN(g6522) );
  OR2X1 U3962 ( .IN1(n3718), .IN2(n1635), .Q(n3745) );
  OR2X1 U3963 ( .IN1(n3717), .IN2(n2529), .Q(n3744) );
  NOR2X0 U3964 ( .IN1(g1713), .IN2(n3746), .QN(g6516) );
  NAND2X0 U3965 ( .IN1(n3747), .IN2(n2938), .QN(n3746) );
  NAND2X0 U3966 ( .IN1(n3748), .IN2(g1781), .QN(n2938) );
  OR2X1 U3967 ( .IN1(g1781), .IN2(n3748), .Q(n3747) );
  NAND2X0 U3968 ( .IN1(n3749), .IN2(n3750), .QN(g6515) );
  OR2X1 U3969 ( .IN1(n3718), .IN2(n2530), .Q(n3750) );
  NAND2X0 U3970 ( .IN1(n3718), .IN2(g1448), .QN(n3749) );
  NAND2X0 U3971 ( .IN1(n3751), .IN2(n3752), .QN(g6514) );
  NAND2X0 U3972 ( .IN1(n3717), .IN2(g1586), .QN(n3752) );
  OR2X1 U3973 ( .IN1(n3717), .IN2(n2532), .Q(n3751) );
  NAND2X0 U3974 ( .IN1(n3753), .IN2(n3754), .QN(g6513) );
  OR2X1 U3975 ( .IN1(n3718), .IN2(n1649), .Q(n3754) );
  NAND2X0 U3976 ( .IN1(n3718), .IN2(g1508), .QN(n3753) );
  NOR2X0 U3977 ( .IN1(n3755), .IN2(g1713), .QN(g6508) );
  NOR2X0 U3978 ( .IN1(n3756), .IN2(n3757), .QN(n3755) );
  NOR2X0 U3979 ( .IN1(n1715), .IN2(n3748), .QN(n3757) );
  NOR2X0 U3980 ( .IN1(n3624), .IN2(n1054), .QN(n3748) );
  NOR2X0 U3981 ( .IN1(n3758), .IN2(n3759), .QN(n3756) );
  NAND2X0 U3982 ( .IN1(test_so5), .IN2(n3624), .QN(n3759) );
  NAND2X0 U3983 ( .IN1(n3760), .IN2(n3761), .QN(g6507) );
  NAND2X0 U3984 ( .IN1(n3717), .IN2(g1604), .QN(n3761) );
  NAND2X0 U3985 ( .IN1(n3718), .IN2(g1444), .QN(n3760) );
  NAND2X0 U3986 ( .IN1(n3762), .IN2(n3763), .QN(g6506) );
  NAND2X0 U3987 ( .IN1(n3717), .IN2(g1583), .QN(n3763) );
  NAND2X0 U3988 ( .IN1(n3718), .IN2(g1424), .QN(n3762) );
  NOR2X0 U3989 ( .IN1(n3764), .IN2(g1713), .QN(g6502) );
  XOR2X1 U3990 ( .IN1(test_so5), .IN2(n3758), .Q(n3764) );
  NAND2X0 U3991 ( .IN1(n256), .IN2(g1766), .QN(n3758) );
  NAND2X0 U3992 ( .IN1(n3765), .IN2(n3766), .QN(g6501) );
  NAND2X0 U3993 ( .IN1(n3717), .IN2(g1601), .QN(n3766) );
  NAND2X0 U3994 ( .IN1(n3718), .IN2(g1440), .QN(n3765) );
  NAND2X0 U3995 ( .IN1(n3767), .IN2(n3768), .QN(g6500) );
  NAND2X0 U3996 ( .IN1(n3717), .IN2(g1580), .QN(n3768) );
  OR2X1 U3997 ( .IN1(n3717), .IN2(n2550), .Q(n3767) );
  NAND2X0 U3998 ( .IN1(n3769), .IN2(n3770), .QN(g6481) );
  NAND2X0 U3999 ( .IN1(n3717), .IN2(g1598), .QN(n3770) );
  NAND2X0 U4000 ( .IN1(n3718), .IN2(g1436), .QN(n3769) );
  NAND2X0 U4001 ( .IN1(n3771), .IN2(n3772), .QN(g6480) );
  OR2X1 U4002 ( .IN1(n3718), .IN2(n2537), .Q(n3772) );
  NAND2X0 U4003 ( .IN1(n3718), .IN2(g1419), .QN(n3771) );
  NAND2X0 U4004 ( .IN1(n3773), .IN2(n3774), .QN(g6479) );
  NAND2X0 U4005 ( .IN1(n3717), .IN2(g1595), .QN(n3774) );
  NAND2X0 U4006 ( .IN1(n3718), .IN2(g1432), .QN(n3773) );
  NAND2X0 U4007 ( .IN1(n3775), .IN2(n3776), .QN(g6478) );
  OR2X1 U4008 ( .IN1(n3718), .IN2(n2551), .Q(n3776) );
  NAND2X0 U4009 ( .IN1(n3718), .IN2(g1515), .QN(n3775) );
  NOR2X0 U4010 ( .IN1(n3777), .IN2(n3656), .QN(g6471) );
  NOR2X0 U4011 ( .IN1(n3778), .IN2(n3680), .QN(n3777) );
  AND2X1 U4012 ( .IN1(n2732), .IN2(n3033), .Q(n3680) );
  NOR2X0 U4013 ( .IN1(n2732), .IN2(n3033), .QN(n3778) );
  NAND2X0 U4014 ( .IN1(n3779), .IN2(n3780), .QN(g6470) );
  OR2X1 U4015 ( .IN1(n3718), .IN2(n2538), .Q(n3780) );
  OR2X1 U4016 ( .IN1(n3717), .IN2(n2655), .Q(n3779) );
  NAND2X0 U4017 ( .IN1(n3781), .IN2(n3782), .QN(g6469) );
  OR2X1 U4018 ( .IN1(n3718), .IN2(n2544), .Q(n3782) );
  NAND2X0 U4019 ( .IN1(n3718), .IN2(g1520), .QN(n3781) );
  NAND2X0 U4020 ( .IN1(n3783), .IN2(n3784), .QN(g6468) );
  OR2X1 U4021 ( .IN1(n3718), .IN2(n2526), .Q(n3784) );
  OR2X1 U4022 ( .IN1(n3717), .IN2(n2527), .Q(n3783) );
  INVX0 U4023 ( .INP(n3718), .ZN(n3717) );
  NAND2X0 U4024 ( .IN1(g109), .IN2(n3693), .QN(n3718) );
  INVX0 U4025 ( .INP(n1159), .ZN(n3693) );
  NOR2X0 U4026 ( .IN1(n2758), .IN2(n3785), .QN(g6439) );
  XOR2X1 U4027 ( .IN1(n3786), .IN2(n3787), .Q(n3785) );
  XOR2X1 U4028 ( .IN1(n2672), .IN2(n2671), .Q(n3787) );
  XOR2X1 U4029 ( .IN1(g182), .IN2(n2670), .Q(n3786) );
  NOR2X0 U4030 ( .IN1(n3492), .IN2(n3788), .QN(g6392) );
  AND2X1 U4031 ( .IN1(g109), .IN2(g881), .Q(n3788) );
  NOR2X0 U4032 ( .IN1(n1603), .IN2(n2759), .QN(g6334) );
  NOR2X0 U4033 ( .IN1(n4947), .IN2(n2760), .QN(g6332) );
  NAND2X0 U4034 ( .IN1(n3789), .IN2(n3790), .QN(g6243) );
  INVX0 U4035 ( .INP(n3463), .ZN(n3790) );
  XNOR2X1 U4036 ( .IN1(n1717), .IN2(n2632), .Q(n3789) );
  NOR2X0 U4037 ( .IN1(n1710), .IN2(n2757), .QN(g6224) );
  NOR2X0 U4038 ( .IN1(n1627), .IN2(n2758), .QN(g6205) );
  NOR2X0 U4039 ( .IN1(n4948), .IN2(n2952), .QN(g6179) );
  NAND2X0 U4040 ( .IN1(g6331), .IN2(n3791), .QN(n2952) );
  NAND2X0 U4041 ( .IN1(n3792), .IN2(n3793), .QN(g6155) );
  NAND2X0 U4042 ( .IN1(g4076), .IN2(g1690), .QN(n3793) );
  NAND2X0 U4043 ( .IN1(n3794), .IN2(n1653), .QN(n3792) );
  NOR2X0 U4044 ( .IN1(n2736), .IN2(n356), .QN(n3794) );
  NOR2X0 U4045 ( .IN1(n3463), .IN2(n3795), .QN(g6126) );
  XOR2X1 U4046 ( .IN1(n2726), .IN2(n2964), .Q(n3795) );
  NOR2X0 U4047 ( .IN1(n3467), .IN2(n3796), .QN(g6123) );
  XOR2X1 U4048 ( .IN1(n2522), .IN2(n1193), .Q(n3796) );
  NAND2X0 U4049 ( .IN1(n3797), .IN2(n3798), .QN(g6099) );
  NAND2X0 U4050 ( .IN1(n3799), .IN2(g342), .QN(n3798) );
  NAND2X0 U4051 ( .IN1(n3800), .IN2(g1074), .QN(n3797) );
  NAND2X0 U4052 ( .IN1(n3801), .IN2(n3802), .QN(g6096) );
  NAND2X0 U4053 ( .IN1(n3799), .IN2(g366), .QN(n3802) );
  NAND2X0 U4054 ( .IN1(n3800), .IN2(g1098), .QN(n3801) );
  NAND2X0 U4055 ( .IN1(n3803), .IN2(n3804), .QN(g6093) );
  NAND2X0 U4056 ( .IN1(n3799), .IN2(g363), .QN(n3804) );
  NAND2X0 U4057 ( .IN1(n3800), .IN2(g1095), .QN(n3803) );
  NAND2X0 U4058 ( .IN1(n3805), .IN2(n3806), .QN(g6088) );
  NAND2X0 U4059 ( .IN1(n3799), .IN2(g360), .QN(n3806) );
  NAND2X0 U4060 ( .IN1(n3800), .IN2(g1092), .QN(n3805) );
  NAND2X0 U4061 ( .IN1(n3807), .IN2(n3808), .QN(g6080) );
  NAND2X0 U4062 ( .IN1(n3799), .IN2(g357), .QN(n3808) );
  NAND2X0 U4063 ( .IN1(n3800), .IN2(g1089), .QN(n3807) );
  NAND2X0 U4064 ( .IN1(n3809), .IN2(n3810), .QN(g6071) );
  NAND2X0 U4065 ( .IN1(n3799), .IN2(g354), .QN(n3810) );
  NAND2X0 U4066 ( .IN1(n3800), .IN2(g1086), .QN(n3809) );
  NAND2X0 U4067 ( .IN1(n3811), .IN2(n3812), .QN(g6068) );
  NAND2X0 U4068 ( .IN1(n3799), .IN2(g351), .QN(n3812) );
  NAND2X0 U4069 ( .IN1(n3800), .IN2(g1083), .QN(n3811) );
  NAND2X0 U4070 ( .IN1(n3813), .IN2(n3814), .QN(g6059) );
  NAND2X0 U4071 ( .IN1(n3799), .IN2(g348), .QN(n3814) );
  NAND2X0 U4072 ( .IN1(n3800), .IN2(g1080), .QN(n3813) );
  NAND2X0 U4073 ( .IN1(n3815), .IN2(n3816), .QN(g6054) );
  NAND2X0 U4074 ( .IN1(n3799), .IN2(g336), .QN(n3816) );
  NAND2X0 U4075 ( .IN1(test_so7), .IN2(n3800), .QN(n3815) );
  NAND2X0 U4076 ( .IN1(n3817), .IN2(n3818), .QN(g6049) );
  NAND2X0 U4077 ( .IN1(n2967), .IN2(g549), .QN(n3817) );
  NAND2X0 U4078 ( .IN1(n3819), .IN2(n3820), .QN(g6045) );
  NAND2X0 U4079 ( .IN1(n2967), .IN2(g575), .QN(n3819) );
  NAND2X0 U4080 ( .IN1(n3821), .IN2(n3822), .QN(g6042) );
  NAND2X0 U4081 ( .IN1(n2967), .IN2(g572), .QN(n3821) );
  NAND2X0 U4082 ( .IN1(n3823), .IN2(n3359), .QN(g6038) );
  NAND2X0 U4083 ( .IN1(g18), .IN2(g237), .QN(n3359) );
  NAND2X0 U4084 ( .IN1(n2967), .IN2(g569), .QN(n3823) );
  NAND2X0 U4085 ( .IN1(n3824), .IN2(n3347), .QN(g6035) );
  NAND2X0 U4086 ( .IN1(g18), .IN2(g231), .QN(n3347) );
  NAND2X0 U4087 ( .IN1(n2967), .IN2(g566), .QN(n3824) );
  NAND2X0 U4088 ( .IN1(n3327), .IN2(n3825), .QN(g6026) );
  NAND2X0 U4089 ( .IN1(n2967), .IN2(g563), .QN(n3825) );
  NAND2X0 U4090 ( .IN1(n3317), .IN2(n3826), .QN(g6015) );
  NAND2X0 U4091 ( .IN1(n2967), .IN2(g560), .QN(n3826) );
  NAND2X0 U4092 ( .IN1(n3364), .IN2(n3827), .QN(g6002) );
  NAND2X0 U4093 ( .IN1(n2967), .IN2(g557), .QN(n3827) );
  NAND2X0 U4094 ( .IN1(n3352), .IN2(n3828), .QN(g6000) );
  NAND2X0 U4095 ( .IN1(n2967), .IN2(g554), .QN(n3828) );
  NAND2X0 U4096 ( .IN1(n3340), .IN2(n3829), .QN(g5996) );
  NAND2X0 U4097 ( .IN1(n2967), .IN2(g546), .QN(n3829) );
  NAND2X0 U4098 ( .IN1(n3830), .IN2(n3831), .QN(g5918) );
  NAND2X0 U4099 ( .IN1(g109), .IN2(g119), .QN(n3831) );
  NAND2X0 U4100 ( .IN1(n3832), .IN2(n3833), .QN(g5914) );
  NAND2X0 U4101 ( .IN1(n3799), .IN2(g345), .QN(n3833) );
  NAND2X0 U4102 ( .IN1(n3800), .IN2(g1077), .QN(n3832) );
  NAND2X0 U4103 ( .IN1(n3834), .IN2(n3835), .QN(g5910) );
  NAND2X0 U4104 ( .IN1(n3799), .IN2(g339), .QN(n3835) );
  NAND2X0 U4105 ( .IN1(n3800), .IN2(g1071), .QN(n3834) );
  NAND2X0 U4106 ( .IN1(n3836), .IN2(n3837), .QN(g5770) );
  NAND2X0 U4107 ( .IN1(n3838), .IN2(n3839), .QN(n3837) );
  NOR2X0 U4108 ( .IN1(n2759), .IN2(g1453), .QN(n3838) );
  NAND2X0 U4109 ( .IN1(g6180), .IN2(n3840), .QN(n3836) );
  INVX0 U4110 ( .INP(n3839), .ZN(n3840) );
  XOR2X1 U4111 ( .IN1(g1508), .IN2(n3841), .Q(n3839) );
  XOR2X1 U4112 ( .IN1(n2687), .IN2(n2673), .Q(n3841) );
  NOR2X0 U4113 ( .IN1(n2760), .IN2(n1628), .QN(g6180) );
  NOR2X0 U4114 ( .IN1(n3842), .IN2(n3843), .QN(g5763) );
  NOR2X0 U4115 ( .IN1(n4949), .IN2(n2759), .QN(n3843) );
  NAND2X0 U4116 ( .IN1(n3844), .IN2(n3845), .QN(g5755) );
  NAND2X0 U4117 ( .IN1(g6333), .IN2(n3846), .QN(n3845) );
  XOR2X1 U4118 ( .IN1(n1619), .IN2(n3847), .Q(n3846) );
  NOR2X0 U4119 ( .IN1(n2757), .IN2(n1678), .QN(g6333) );
  NAND2X0 U4120 ( .IN1(n3848), .IN2(n1678), .QN(n3844) );
  NOR2X0 U4121 ( .IN1(n3849), .IN2(n3850), .QN(n3848) );
  NOR2X0 U4122 ( .IN1(g6331), .IN2(n3847), .QN(n3850) );
  INVX0 U4123 ( .INP(n3851), .ZN(n3847) );
  NOR2X0 U4124 ( .IN1(n2758), .IN2(n1619), .QN(g6331) );
  NOR2X0 U4125 ( .IN1(n3852), .IN2(n3851), .QN(n3849) );
  XOR2X1 U4126 ( .IN1(g1389), .IN2(n3853), .Q(n3851) );
  NOR2X0 U4127 ( .IN1(n18), .IN2(g1386), .QN(n3853) );
  AND2X1 U4128 ( .IN1(n1619), .IN2(n3791), .Q(n18) );
  AND2X1 U4129 ( .IN1(n3854), .IN2(n3855), .Q(n3791) );
  NOR2X0 U4130 ( .IN1(n3856), .IN2(n3857), .QN(n3855) );
  NAND2X0 U4131 ( .IN1(n3858), .IN2(n3859), .QN(n3857) );
  NOR2X0 U4132 ( .IN1(g207), .IN2(n3860), .QN(n3859) );
  NAND2X0 U4133 ( .IN1(n2511), .IN2(n2510), .QN(n3860) );
  NOR2X0 U4134 ( .IN1(g192), .IN2(n3861), .QN(n3858) );
  NAND2X0 U4135 ( .IN1(n2514), .IN2(n2513), .QN(n3861) );
  NAND2X0 U4136 ( .IN1(n3862), .IN2(n3863), .QN(n3856) );
  NOR2X0 U4137 ( .IN1(g1389), .IN2(n3864), .QN(n3863) );
  NAND2X0 U4138 ( .IN1(n1598), .IN2(n2674), .QN(n3864) );
  NOR2X0 U4139 ( .IN1(g1397), .IN2(n3865), .QN(n3862) );
  NAND2X0 U4140 ( .IN1(n1678), .IN2(n1629), .QN(n3865) );
  NOR2X0 U4141 ( .IN1(n3866), .IN2(n3867), .QN(n3854) );
  NAND2X0 U4142 ( .IN1(n3868), .IN2(n3869), .QN(n3867) );
  NOR2X0 U4143 ( .IN1(n3038), .IN2(n3870), .QN(n3869) );
  NAND2X0 U4144 ( .IN1(n4945), .IN2(n4947), .QN(n3870) );
  AND2X1 U4145 ( .IN1(n4942), .IN2(n4941), .Q(n3868) );
  NAND2X0 U4146 ( .IN1(n3871), .IN2(n3872), .QN(n3866) );
  NOR2X0 U4147 ( .IN1(g225), .IN2(n3873), .QN(n3872) );
  NAND2X0 U4148 ( .IN1(n2675), .IN2(n2668), .QN(n3873) );
  NOR2X0 U4149 ( .IN1(g243), .IN2(n3874), .QN(n3871) );
  NAND2X0 U4150 ( .IN1(n2678), .IN2(n2677), .QN(n3874) );
  NOR2X0 U4151 ( .IN1(n2759), .IN2(g201), .QN(n3852) );
  AND2X1 U4152 ( .IN1(n3875), .IN2(g744), .Q(g5659) );
  AND2X1 U4153 ( .IN1(g743), .IN2(g109), .Q(n3875) );
  AND2X1 U4154 ( .IN1(n3876), .IN2(g742), .Q(g5658) );
  AND2X1 U4155 ( .IN1(g741), .IN2(g109), .Q(n3876) );
  NOR2X0 U4156 ( .IN1(n3877), .IN2(n3878), .QN(g5556) );
  NAND2X0 U4157 ( .IN1(n3879), .IN2(n3880), .QN(n3878) );
  NOR2X0 U4158 ( .IN1(n1653), .IN2(n1626), .QN(n3880) );
  NOR2X0 U4159 ( .IN1(n3624), .IN2(g1781), .QN(n3879) );
  NAND2X0 U4160 ( .IN1(n3881), .IN2(test_so5), .QN(n3624) );
  NOR2X0 U4161 ( .IN1(n2728), .IN2(n1715), .QN(n3881) );
  NAND2X0 U4162 ( .IN1(n3882), .IN2(n3883), .QN(n3877) );
  NOR2X0 U4163 ( .IN1(n2734), .IN2(n3884), .QN(n3883) );
  NAND2X0 U4164 ( .IN1(g1786), .IN2(g1707), .QN(n3884) );
  NOR2X0 U4165 ( .IN1(n2733), .IN2(n1702), .QN(n3882) );
  NOR2X0 U4166 ( .IN1(n2964), .IN2(n3885), .QN(g5543) );
  NOR2X0 U4167 ( .IN1(n3886), .IN2(n3887), .QN(n3885) );
  NOR2X0 U4168 ( .IN1(n1717), .IN2(g5849), .QN(n3887) );
  OR2X1 U4169 ( .IN1(n3463), .IN2(n2632), .Q(g5849) );
  NOR2X0 U4170 ( .IN1(n1622), .IN2(n3463), .QN(n3886) );
  NAND2X0 U4171 ( .IN1(n3888), .IN2(g109), .QN(n3463) );
  NOR2X0 U4172 ( .IN1(n2731), .IN2(n2505), .QN(n3888) );
  NOR2X0 U4173 ( .IN1(n3395), .IN2(n1622), .QN(n2964) );
  OR2X1 U4174 ( .IN1(n2632), .IN2(n1717), .Q(n3395) );
  NOR2X0 U4175 ( .IN1(n3467), .IN2(n3889), .QN(g5536) );
  OR2X1 U4176 ( .IN1(n1213), .IN2(n1193), .Q(n3889) );
  NAND2X0 U4177 ( .IN1(n3890), .IN2(n3891), .QN(g5529) );
  NAND2X0 U4178 ( .IN1(g4940), .IN2(g4174), .QN(n3891) );
  NAND2X0 U4179 ( .IN1(n3892), .IN2(n2520), .QN(n3890) );
  NOR2X0 U4180 ( .IN1(n2521), .IN2(n3467), .QN(n3892) );
  INVX0 U4181 ( .INP(n3893), .ZN(n3467) );
  NAND2X0 U4182 ( .IN1(n3830), .IN2(n3894), .QN(g5445) );
  OR2X1 U4183 ( .IN1(n2759), .IN2(n2622), .Q(n3894) );
  NAND2X0 U4184 ( .IN1(n3830), .IN2(n3895), .QN(g5421) );
  OR2X1 U4185 ( .IN1(n2760), .IN2(n2623), .Q(n3895) );
  INVX0 U4186 ( .INP(n1195), .ZN(n3830) );
  NAND2X0 U4187 ( .IN1(n3896), .IN2(n3897), .QN(g5404) );
  NAND2X0 U4188 ( .IN1(n3306), .IN2(g1713), .QN(n3897) );
  NAND2X0 U4189 ( .IN1(n968), .IN2(g1718), .QN(n3896) );
  NAND2X0 U4190 ( .IN1(n3898), .IN2(n3899), .QN(g5396) );
  NAND2X0 U4191 ( .IN1(n3306), .IN2(g1710), .QN(n3899) );
  NAND2X0 U4192 ( .IN1(n968), .IN2(g1713), .QN(n3898) );
  NOR2X0 U4193 ( .IN1(n1654), .IN2(n3900), .QN(g5390) );
  NOR2X0 U4194 ( .IN1(n1677), .IN2(n3900), .QN(g5173) );
  NOR2X0 U4195 ( .IN1(n1614), .IN2(n3900), .QN(g5148) );
  NOR2X0 U4196 ( .IN1(n1658), .IN2(n3900), .QN(g5126) );
  NAND2X0 U4197 ( .IN1(g109), .IN2(DFF_126_n1), .QN(n3900) );
  NOR2X0 U4198 ( .IN1(n3306), .IN2(n3901), .QN(g5083) );
  OR2X1 U4199 ( .IN1(n3902), .IN2(g4089), .Q(n3901) );
  AND2X1 U4200 ( .IN1(n2521), .IN2(n3893), .Q(g4940) );
  NOR2X0 U4201 ( .IN1(n2760), .IN2(test_so1), .QN(n3893) );
  NOR2X0 U4202 ( .IN1(n2753), .IN2(DFF_489_n1), .QN(g4905) );
  INVX0 U4203 ( .INP(n3903), .ZN(g4904) );
  NOR2X0 U4204 ( .IN1(n2753), .IN2(DFF_330_n1), .QN(g4903) );
  NOR2X0 U4205 ( .IN1(n2753), .IN2(DFF_385_n1), .QN(g4902) );
  NOR2X0 U4206 ( .IN1(n2751), .IN2(DFF_157_n1), .QN(g4893) );
  INVX0 U4207 ( .INP(n3387), .ZN(g4892) );
  NAND2X0 U4208 ( .IN1(n3700), .IN2(n3059), .QN(n3387) );
  INVX0 U4209 ( .INP(n2751), .ZN(n3700) );
  NOR2X0 U4210 ( .IN1(n2751), .IN2(DFF_136_n1), .QN(g4891) );
  NOR2X0 U4211 ( .IN1(n2751), .IN2(DFF_336_n1), .QN(g4890) );
  NAND2X0 U4212 ( .IN1(n3300), .IN2(n3904), .QN(n2751) );
  NAND2X0 U4213 ( .IN1(n1607), .IN2(g611), .QN(n3904) );
  NAND2X0 U4214 ( .IN1(n3905), .IN2(n3293), .QN(n3300) );
  INVX0 U4215 ( .INP(n3388), .ZN(n3293) );
  NAND2X0 U4216 ( .IN1(n1609), .IN2(n1644), .QN(n3388) );
  NOR2X0 U4217 ( .IN1(g591), .IN2(g605), .QN(n3905) );
  NAND2X0 U4218 ( .IN1(n2744), .IN2(n2743), .QN(g4556) );
  NOR2X0 U4219 ( .IN1(n4950), .IN2(n2760), .QN(g4506) );
  NOR2X0 U4220 ( .IN1(n4951), .IN2(n3306), .QN(g4500) );
  NOR2X0 U4221 ( .IN1(n1617), .IN2(n2757), .QN(g4498) );
  NOR2X0 U4222 ( .IN1(n1660), .IN2(n2758), .QN(g4490) );
  NOR2X0 U4223 ( .IN1(n1597), .IN2(n2759), .QN(g4484) );
  NOR2X0 U4224 ( .IN1(n1706), .IN2(n2760), .QN(g4480) );
  NOR2X0 U4225 ( .IN1(n1705), .IN2(n2757), .QN(g4477) );
  NOR2X0 U4226 ( .IN1(n1708), .IN2(n2758), .QN(g4473) );
  NOR2X0 U4227 ( .IN1(n1618), .IN2(n2759), .QN(g4471) );
  NOR2X0 U4228 ( .IN1(n2757), .IN2(n2755), .QN(g4465) );
  NOR2X0 U4229 ( .IN1(n1685), .IN2(n2760), .QN(g4342) );
  NOR2X0 U4230 ( .IN1(n1686), .IN2(n2757), .QN(g4340) );
  NAND2X0 U4231 ( .IN1(n3906), .IN2(n3907), .QN(g4309) );
  NAND2X0 U4232 ( .IN1(n3908), .IN2(g1806), .QN(n3907) );
  OR2X1 U4233 ( .IN1(n3908), .IN2(n2715), .Q(n3906) );
  NAND2X0 U4234 ( .IN1(n3909), .IN2(n3910), .QN(g4293) );
  NAND2X0 U4235 ( .IN1(n3908), .IN2(g1801), .QN(n3910) );
  OR2X1 U4236 ( .IN1(n3908), .IN2(n2717), .Q(n3909) );
  NAND2X0 U4237 ( .IN1(n3911), .IN2(n3912), .QN(g4283) );
  NAND2X0 U4238 ( .IN1(n3908), .IN2(g1796), .QN(n3912) );
  NAND2X0 U4239 ( .IN1(n3913), .IN2(g1756), .QN(n3911) );
  NAND2X0 U4240 ( .IN1(n3914), .IN2(n3915), .QN(g4274) );
  NAND2X0 U4241 ( .IN1(n3908), .IN2(g1791), .QN(n3915) );
  OR2X1 U4242 ( .IN1(n3908), .IN2(n2716), .Q(n3914) );
  NAND2X0 U4243 ( .IN1(n3916), .IN2(n3917), .QN(g4264) );
  NAND2X0 U4244 ( .IN1(n3908), .IN2(g1786), .QN(n3917) );
  OR2X1 U4245 ( .IN1(n3908), .IN2(n2712), .Q(n3916) );
  NAND2X0 U4246 ( .IN1(n3918), .IN2(n3919), .QN(g4255) );
  NAND2X0 U4247 ( .IN1(n3908), .IN2(g1781), .QN(n3919) );
  OR2X1 U4248 ( .IN1(n3908), .IN2(n2714), .Q(n3918) );
  NAND2X0 U4249 ( .IN1(n3920), .IN2(n3921), .QN(g4239) );
  NAND2X0 U4250 ( .IN1(n3908), .IN2(g1776), .QN(n3921) );
  NAND2X0 U4251 ( .IN1(n3913), .IN2(g1744), .QN(n3920) );
  NAND2X0 U4252 ( .IN1(n3922), .IN2(n3923), .QN(g4238) );
  NAND2X0 U4253 ( .IN1(n3908), .IN2(test_so5), .QN(n3923) );
  NAND2X0 U4254 ( .IN1(n3913), .IN2(g1741), .QN(n3922) );
  NAND2X0 U4255 ( .IN1(n3924), .IN2(n3925), .QN(g4231) );
  NAND2X0 U4256 ( .IN1(n3908), .IN2(g1766), .QN(n3925) );
  OR2X1 U4257 ( .IN1(n3908), .IN2(n1640), .Q(n3924) );
  INVX0 U4258 ( .INP(n3913), .ZN(n3908) );
  NAND2X0 U4259 ( .IN1(g1700), .IN2(DFF_275_n1), .QN(g4089) );
  NOR2X0 U4260 ( .IN1(g1707), .IN2(n356), .QN(g4076) );
  INVX0 U4261 ( .INP(g1700), .ZN(n356) );
  NOR2X0 U4262 ( .IN1(n2731), .IN2(n3926), .QN(g3462) );
  NOR2X0 U4263 ( .IN1(n3927), .IN2(n3714), .QN(n3926) );
  NOR2X0 U4264 ( .IN1(n1647), .IN2(g750), .QN(n3927) );
  NOR2X0 U4265 ( .IN1(n3928), .IN2(n3929), .QN(g3381) );
  OR2X1 U4266 ( .IN1(n1591), .IN2(n1604), .Q(n3929) );
  NAND2X0 U4267 ( .IN1(g936), .IN2(g940), .QN(n3928) );
  INVX0 U4268 ( .INP(g23), .ZN(g3327) );
  NOR2X0 U4269 ( .IN1(g1610), .IN2(g1737), .QN(g2478) );
  NAND2X0 U4270 ( .IN1(n3930), .IN2(n3931), .QN(g11647) );
  NAND2X0 U4271 ( .IN1(n3591), .IN2(g336), .QN(n3931) );
  NAND2X0 U4272 ( .IN1(n3714), .IN2(n3932), .QN(n3930) );
  NAND2X0 U4273 ( .IN1(n3933), .IN2(n3934), .QN(n3932) );
  NAND2X0 U4274 ( .IN1(n3935), .IN2(n3936), .QN(n3934) );
  NAND2X0 U4275 ( .IN1(n3937), .IN2(n3938), .QN(n3933) );
  INVX0 U4276 ( .INP(n3936), .ZN(n3937) );
  NOR2X0 U4277 ( .IN1(n3939), .IN2(n3940), .QN(g11641) );
  NOR2X0 U4278 ( .IN1(n3941), .IN2(n3942), .QN(n3939) );
  NOR2X0 U4279 ( .IN1(n1721), .IN2(n1226), .QN(n3942) );
  NOR2X0 U4280 ( .IN1(n3943), .IN2(n1227), .QN(n1226) );
  NOR2X0 U4281 ( .IN1(n3944), .IN2(n3945), .QN(n3941) );
  NAND2X0 U4282 ( .IN1(n3), .IN2(n3943), .QN(n3945) );
  INVX0 U4283 ( .INP(n2752), .ZN(n3943) );
  NOR2X0 U4284 ( .IN1(n3944), .IN2(n1721), .QN(n2752) );
  INVX0 U4285 ( .INP(n1229), .ZN(n3944) );
  NOR2X0 U4286 ( .IN1(n3946), .IN2(n2705), .QN(n1229) );
  OR2X1 U4287 ( .IN1(n2707), .IN2(n2706), .Q(n3946) );
  NOR2X0 U4288 ( .IN1(n3947), .IN2(n3940), .QN(g11640) );
  NOR2X0 U4289 ( .IN1(n3948), .IN2(n3949), .QN(n3947) );
  AND2X1 U4290 ( .IN1(n1232), .IN2(n1231), .Q(n3949) );
  NOR2X0 U4291 ( .IN1(n2706), .IN2(n3950), .QN(n3948) );
  NOR2X0 U4292 ( .IN1(n1227), .IN2(n3951), .QN(n3950) );
  OR2X1 U4293 ( .IN1(n2705), .IN2(n2707), .Q(n3951) );
  NOR2X0 U4294 ( .IN1(n3940), .IN2(n3952), .QN(g11639) );
  XOR2X1 U4295 ( .IN1(n2705), .IN2(n1231), .Q(n3952) );
  NOR2X0 U4296 ( .IN1(n3940), .IN2(n3953), .QN(g11636) );
  XOR2X1 U4297 ( .IN1(n2707), .IN2(n3), .Q(n3953) );
  NAND2X0 U4298 ( .IN1(n3954), .IN2(g109), .QN(n3940) );
  NAND2X0 U4299 ( .IN1(n3955), .IN2(n4949), .QN(n3954) );
  NOR2X0 U4300 ( .IN1(n2743), .IN2(n3842), .QN(n3955) );
  INVX0 U4301 ( .INP(n3956), .ZN(n3842) );
  NAND2X0 U4302 ( .IN1(n3957), .IN2(n3958), .QN(g11625) );
  NAND2X0 U4303 ( .IN1(n3591), .IN2(g345), .QN(n3958) );
  NAND2X0 U4304 ( .IN1(n3714), .IN2(n3959), .QN(n3957) );
  XOR2X1 U4305 ( .IN1(n3935), .IN2(n3938), .Q(n3959) );
  AND2X1 U4306 ( .IN1(n3960), .IN2(n3961), .Q(n3938) );
  OR2X1 U4307 ( .IN1(n1239), .IN2(n1681), .Q(n3961) );
  NAND2X0 U4308 ( .IN1(n3962), .IN2(n1239), .QN(n3960) );
  XNOR2X1 U4309 ( .IN1(n3963), .IN2(n3964), .Q(n3962) );
  NAND2X0 U4310 ( .IN1(n1646), .IN2(n3965), .QN(n3963) );
  XOR2X1 U4311 ( .IN1(n3966), .IN2(n3967), .Q(n3935) );
  XOR2X1 U4312 ( .IN1(n3968), .IN2(n3969), .Q(n3967) );
  XOR2X1 U4313 ( .IN1(n3970), .IN2(n3971), .Q(n3969) );
  XOR2X1 U4314 ( .IN1(n3972), .IN2(n3973), .Q(n3971) );
  XOR2X1 U4315 ( .IN1(n3974), .IN2(n3975), .Q(n3970) );
  XOR2X1 U4316 ( .IN1(n3976), .IN2(n3977), .Q(n3968) );
  XOR2X1 U4317 ( .IN1(n3978), .IN2(n3979), .Q(n3977) );
  XOR2X1 U4318 ( .IN1(n3980), .IN2(n3981), .Q(n3976) );
  NAND2X0 U4319 ( .IN1(n3982), .IN2(n3983), .QN(g11610) );
  NAND2X0 U4320 ( .IN1(n3984), .IN2(g1806), .QN(n3983) );
  OR2X1 U4321 ( .IN1(n3984), .IN2(n2478), .Q(n3982) );
  NAND2X0 U4322 ( .IN1(n3985), .IN2(n3986), .QN(g11609) );
  NAND2X0 U4323 ( .IN1(n3984), .IN2(g1801), .QN(n3986) );
  NAND2X0 U4324 ( .IN1(n3987), .IN2(g1330), .QN(n3985) );
  NAND2X0 U4325 ( .IN1(n3988), .IN2(n3989), .QN(g11608) );
  NAND2X0 U4326 ( .IN1(n3984), .IN2(g1796), .QN(n3989) );
  NAND2X0 U4327 ( .IN1(n3987), .IN2(g1327), .QN(n3988) );
  NAND2X0 U4328 ( .IN1(n3990), .IN2(n3991), .QN(g11607) );
  NAND2X0 U4329 ( .IN1(n3984), .IN2(g1791), .QN(n3991) );
  OR2X1 U4330 ( .IN1(n3984), .IN2(n2472), .Q(n3990) );
  NAND2X0 U4331 ( .IN1(n3992), .IN2(n3993), .QN(g11606) );
  NAND2X0 U4332 ( .IN1(n3984), .IN2(g1786), .QN(n3993) );
  OR2X1 U4333 ( .IN1(n3984), .IN2(n2476), .Q(n3992) );
  NAND2X0 U4334 ( .IN1(n3994), .IN2(n3995), .QN(g11605) );
  NAND2X0 U4335 ( .IN1(n3984), .IN2(g1781), .QN(n3995) );
  NAND2X0 U4336 ( .IN1(n3987), .IN2(g1318), .QN(n3994) );
  NAND2X0 U4337 ( .IN1(n3996), .IN2(n3997), .QN(g11604) );
  NAND2X0 U4338 ( .IN1(n3984), .IN2(g1776), .QN(n3997) );
  NAND2X0 U4339 ( .IN1(n3987), .IN2(g1314), .QN(n3996) );
  NAND2X0 U4340 ( .IN1(n3998), .IN2(n3999), .QN(g11603) );
  NAND2X0 U4341 ( .IN1(test_so9), .IN2(n3987), .QN(n3999) );
  NAND2X0 U4342 ( .IN1(n3984), .IN2(test_so5), .QN(n3998) );
  NAND2X0 U4343 ( .IN1(n4000), .IN2(n4001), .QN(g11602) );
  NAND2X0 U4344 ( .IN1(n3984), .IN2(g1766), .QN(n4001) );
  OR2X1 U4345 ( .IN1(n3984), .IN2(n2479), .Q(n4000) );
  INVX0 U4346 ( .INP(n3987), .ZN(n3984) );
  NAND2X0 U4347 ( .IN1(n3), .IN2(g1317), .QN(n3987) );
  INVX0 U4348 ( .INP(n1227), .ZN(n3) );
  NAND2X0 U4349 ( .IN1(n4002), .IN2(n3552), .QN(n1227) );
  NOR2X0 U4350 ( .IN1(n4003), .IN2(n3553), .QN(n4002) );
  NOR2X0 U4351 ( .IN1(n4004), .IN2(n4005), .QN(n4003) );
  NAND2X0 U4352 ( .IN1(n4006), .IN2(n4007), .QN(n4005) );
  NOR2X0 U4353 ( .IN1(n4008), .IN2(n4009), .QN(n4007) );
  NAND2X0 U4354 ( .IN1(n4010), .IN2(n4011), .QN(n4009) );
  XOR2X1 U4355 ( .IN1(n2658), .IN2(g1250), .Q(n4011) );
  XOR2X1 U4356 ( .IN1(n1871), .IN2(g1235), .Q(n4010) );
  XOR2X1 U4357 ( .IN1(n2630), .IN2(n2619), .Q(n4008) );
  NOR2X0 U4358 ( .IN1(n4012), .IN2(n4013), .QN(n4006) );
  XOR2X1 U4359 ( .IN1(n2700), .IN2(n2699), .Q(n4013) );
  XOR2X1 U4360 ( .IN1(n2698), .IN2(n2697), .Q(n4012) );
  NAND2X0 U4361 ( .IN1(n4014), .IN2(n4015), .QN(n4004) );
  NOR2X0 U4362 ( .IN1(n4016), .IN2(n4017), .QN(n4015) );
  NAND2X0 U4363 ( .IN1(n4018), .IN2(n4019), .QN(n4017) );
  XOR2X1 U4364 ( .IN1(test_so2), .IN2(n2629), .Q(n4019) );
  XOR2X1 U4365 ( .IN1(n4020), .IN2(n4021), .Q(n4018) );
  XNOR2X1 U4366 ( .IN1(n2593), .IN2(test_so6), .Q(n4016) );
  NOR2X0 U4367 ( .IN1(n4022), .IN2(n4023), .QN(n4014) );
  XOR2X1 U4368 ( .IN1(n2633), .IN2(n2618), .Q(n4023) );
  XOR2X1 U4369 ( .IN1(test_so8), .IN2(g1245), .Q(n4022) );
  NAND2X0 U4370 ( .IN1(n4024), .IN2(n4025), .QN(g11579) );
  NAND2X0 U4371 ( .IN1(n968), .IN2(g1618), .QN(n4025) );
  NAND2X0 U4372 ( .IN1(n4026), .IN2(n3306), .QN(n4024) );
  XOR2X1 U4373 ( .IN1(g1610), .IN2(n4027), .Q(n4026) );
  NAND2X0 U4374 ( .IN1(n4028), .IN2(n4029), .QN(n4027) );
  NAND2X0 U4375 ( .IN1(n4030), .IN2(n4031), .QN(n4029) );
  NAND2X0 U4376 ( .IN1(n1262), .IN2(n2953), .QN(n4031) );
  NAND2X0 U4377 ( .IN1(n4032), .IN2(n4033), .QN(n2953) );
  NAND2X0 U4378 ( .IN1(n4034), .IN2(n1677), .QN(n4033) );
  NOR2X0 U4379 ( .IN1(n4035), .IN2(n4036), .QN(n4032) );
  NOR2X0 U4380 ( .IN1(n4037), .IN2(g1149), .QN(n4036) );
  NOR2X0 U4381 ( .IN1(n1685), .IN2(g1153), .QN(n4035) );
  NAND2X0 U4382 ( .IN1(n4038), .IN2(n4034), .QN(n1262) );
  NOR2X0 U4383 ( .IN1(n3344), .IN2(g1104), .QN(n4034) );
  NAND2X0 U4384 ( .IN1(n1614), .IN2(g1101), .QN(n3344) );
  NOR2X0 U4385 ( .IN1(g1110), .IN2(n4039), .QN(n4038) );
  NAND2X0 U4386 ( .IN1(n4040), .IN2(n4041), .QN(n4039) );
  NAND2X0 U4387 ( .IN1(g1149), .IN2(g1153), .QN(n4041) );
  NAND2X0 U4388 ( .IN1(n1685), .IN2(n4037), .QN(n4040) );
  AND2X1 U4389 ( .IN1(n1686), .IN2(n4042), .Q(n4037) );
  NAND2X0 U4390 ( .IN1(n4043), .IN2(n4044), .QN(n4042) );
  NOR2X0 U4391 ( .IN1(n4045), .IN2(n4046), .QN(n4044) );
  NAND2X0 U4392 ( .IN1(n4047), .IN2(n1706), .QN(n4046) );
  AND2X1 U4393 ( .IN1(n1660), .IN2(n1705), .Q(n4047) );
  NAND2X0 U4394 ( .IN1(n4048), .IN2(n4049), .QN(n4045) );
  AND2X1 U4395 ( .IN1(n2755), .IN2(n1597), .Q(n4049) );
  AND2X1 U4396 ( .IN1(n1617), .IN2(n1618), .Q(n4048) );
  NOR2X0 U4397 ( .IN1(n4050), .IN2(n4051), .QN(n4043) );
  NAND2X0 U4398 ( .IN1(n4052), .IN2(n4932), .QN(n4051) );
  NOR2X0 U4399 ( .IN1(n3016), .IN2(g1163), .QN(n4052) );
  NAND2X0 U4400 ( .IN1(n4053), .IN2(n2667), .QN(n4050) );
  NOR2X0 U4401 ( .IN1(g1125), .IN2(g1157), .QN(n4053) );
  NAND2X0 U4402 ( .IN1(n1260), .IN2(n4054), .QN(n4028) );
  NAND2X0 U4403 ( .IN1(n4055), .IN2(n4056), .QN(g11514) );
  NAND2X0 U4404 ( .IN1(n4057), .IN2(n4058), .QN(n4056) );
  INVX0 U4405 ( .INP(n4059), .ZN(n4058) );
  NOR2X0 U4406 ( .IN1(n2758), .IN2(g1419), .QN(n4057) );
  NAND2X0 U4407 ( .IN1(g6193), .IN2(n4059), .QN(n4055) );
  XOR2X1 U4408 ( .IN1(n4060), .IN2(n4061), .Q(n4059) );
  XOR2X1 U4409 ( .IN1(n2653), .IN2(n2527), .Q(n4061) );
  XOR2X1 U4410 ( .IN1(g1515), .IN2(n4054), .Q(n4060) );
  INVX0 U4411 ( .INP(n4030), .ZN(n4054) );
  NAND2X0 U4412 ( .IN1(n4062), .IN2(n4063), .QN(n4030) );
  NAND2X0 U4413 ( .IN1(g18), .IN2(g201), .QN(n4063) );
  NAND2X0 U4414 ( .IN1(n4064), .IN2(n2967), .QN(n4062) );
  NAND2X0 U4415 ( .IN1(n4065), .IN2(n4066), .QN(n4064) );
  OR2X1 U4416 ( .IN1(n4067), .IN2(g1811), .Q(n4066) );
  NAND2X0 U4417 ( .IN1(n4067), .IN2(n4068), .QN(n4065) );
  NAND2X0 U4418 ( .IN1(n4069), .IN2(n4070), .QN(n4068) );
  NAND2X0 U4419 ( .IN1(n4071), .IN2(n4072), .QN(n4067) );
  AND2X1 U4420 ( .IN1(n4955), .IN2(n4954), .Q(n4072) );
  AND2X1 U4421 ( .IN1(n4953), .IN2(n4952), .Q(n4071) );
  NOR2X0 U4422 ( .IN1(n2759), .IN2(n1602), .QN(g6193) );
  NAND2X0 U4423 ( .IN1(n4073), .IN2(n4074), .QN(g11488) );
  NAND2X0 U4424 ( .IN1(n3591), .IN2(g342), .QN(n4074) );
  NAND2X0 U4425 ( .IN1(n3714), .IN2(n3981), .QN(n4073) );
  NAND2X0 U4426 ( .IN1(n4075), .IN2(n4076), .QN(n3981) );
  OR2X1 U4427 ( .IN1(n1239), .IN2(n2458), .Q(n4076) );
  NAND2X0 U4428 ( .IN1(n4077), .IN2(n1239), .QN(n4075) );
  XOR2X1 U4429 ( .IN1(n4078), .IN2(n1620), .Q(n4077) );
  NAND2X0 U4430 ( .IN1(n4079), .IN2(n4080), .QN(n4078) );
  NOR2X0 U4431 ( .IN1(n1641), .IN2(n1606), .QN(n4080) );
  NOR2X0 U4432 ( .IN1(g461), .IN2(g466), .QN(n4079) );
  NAND2X0 U4433 ( .IN1(n4081), .IN2(n4082), .QN(g11487) );
  NAND2X0 U4434 ( .IN1(n3591), .IN2(g366), .QN(n4082) );
  NAND2X0 U4435 ( .IN1(n3714), .IN2(n3980), .QN(n4081) );
  NAND2X0 U4436 ( .IN1(n4083), .IN2(n4084), .QN(n3980) );
  OR2X1 U4437 ( .IN1(n1239), .IN2(n2685), .Q(n4084) );
  NAND2X0 U4438 ( .IN1(n4085), .IN2(n1239), .QN(n4083) );
  XOR2X1 U4439 ( .IN1(n4086), .IN2(n1679), .Q(n4085) );
  NAND2X0 U4440 ( .IN1(n4087), .IN2(n1594), .QN(n4086) );
  NAND2X0 U4441 ( .IN1(n4088), .IN2(n4089), .QN(g11486) );
  NAND2X0 U4442 ( .IN1(n3591), .IN2(g363), .QN(n4089) );
  NAND2X0 U4443 ( .IN1(n3714), .IN2(n3979), .QN(n4088) );
  NAND2X0 U4444 ( .IN1(n4090), .IN2(n4091), .QN(n3979) );
  OR2X1 U4445 ( .IN1(n1239), .IN2(n2457), .Q(n4091) );
  NAND2X0 U4446 ( .IN1(n4092), .IN2(n1239), .QN(n4090) );
  XOR2X1 U4447 ( .IN1(g506), .IN2(n4093), .Q(n4092) );
  NOR2X0 U4448 ( .IN1(g471), .IN2(n4094), .QN(n4093) );
  NAND2X0 U4449 ( .IN1(n4095), .IN2(n4096), .QN(g11485) );
  NAND2X0 U4450 ( .IN1(n3591), .IN2(g360), .QN(n4096) );
  NAND2X0 U4451 ( .IN1(n3714), .IN2(n3975), .QN(n4095) );
  NAND2X0 U4452 ( .IN1(n4097), .IN2(n4098), .QN(n3975) );
  OR2X1 U4453 ( .IN1(n1239), .IN2(n2664), .Q(n4098) );
  NAND2X0 U4454 ( .IN1(n4099), .IN2(n1239), .QN(n4097) );
  XOR2X1 U4455 ( .IN1(n4100), .IN2(n1690), .Q(n4099) );
  NAND2X0 U4456 ( .IN1(n4101), .IN2(g461), .QN(n4100) );
  NAND2X0 U4457 ( .IN1(n4102), .IN2(n4103), .QN(g11484) );
  NAND2X0 U4458 ( .IN1(n3591), .IN2(g357), .QN(n4103) );
  NAND2X0 U4459 ( .IN1(n3714), .IN2(n3974), .QN(n4102) );
  NAND2X0 U4460 ( .IN1(n4104), .IN2(n4105), .QN(n3974) );
  OR2X1 U4461 ( .IN1(n1239), .IN2(n2660), .Q(n4105) );
  NAND2X0 U4462 ( .IN1(n4106), .IN2(n1239), .QN(n4104) );
  XOR2X1 U4463 ( .IN1(n4107), .IN2(n1689), .Q(n4106) );
  NAND2X0 U4464 ( .IN1(n3965), .IN2(g466), .QN(n4107) );
  AND2X1 U4465 ( .IN1(n4108), .IN2(n1606), .Q(n3965) );
  NOR2X0 U4466 ( .IN1(n1641), .IN2(g461), .QN(n4108) );
  NAND2X0 U4467 ( .IN1(n4109), .IN2(n4110), .QN(g11483) );
  NAND2X0 U4468 ( .IN1(n3591), .IN2(g354), .QN(n4110) );
  NAND2X0 U4469 ( .IN1(n3714), .IN2(n3973), .QN(n4109) );
  NAND2X0 U4470 ( .IN1(n4111), .IN2(n4112), .QN(n3973) );
  OR2X1 U4471 ( .IN1(n1239), .IN2(n2704), .Q(n4112) );
  NAND2X0 U4472 ( .IN1(n4113), .IN2(n1239), .QN(n4111) );
  XOR2X1 U4473 ( .IN1(n4114), .IN2(n1691), .Q(n4113) );
  NAND2X0 U4474 ( .IN1(n4101), .IN2(n1594), .QN(n4114) );
  AND2X1 U4475 ( .IN1(n4115), .IN2(n1641), .Q(n4101) );
  NOR2X0 U4476 ( .IN1(n1646), .IN2(g471), .QN(n4115) );
  NAND2X0 U4477 ( .IN1(n4116), .IN2(n4117), .QN(g11482) );
  NAND2X0 U4478 ( .IN1(n3591), .IN2(g351), .QN(n4117) );
  NAND2X0 U4479 ( .IN1(n3714), .IN2(n3966), .QN(n4116) );
  NAND2X0 U4480 ( .IN1(n4118), .IN2(n4119), .QN(n3966) );
  OR2X1 U4481 ( .IN1(n1239), .IN2(n2662), .Q(n4119) );
  NAND2X0 U4482 ( .IN1(n4120), .IN2(n1239), .QN(n4118) );
  XOR2X1 U4483 ( .IN1(n4121), .IN2(n1621), .Q(n4120) );
  OR2X1 U4484 ( .IN1(n4122), .IN2(n1641), .Q(n4121) );
  NAND2X0 U4485 ( .IN1(n4123), .IN2(n4124), .QN(g11481) );
  NAND2X0 U4486 ( .IN1(n3591), .IN2(g348), .QN(n4124) );
  NAND2X0 U4487 ( .IN1(n3714), .IN2(n3972), .QN(n4123) );
  NAND2X0 U4488 ( .IN1(n4125), .IN2(n4126), .QN(n3972) );
  OR2X1 U4489 ( .IN1(n1239), .IN2(n2702), .Q(n4126) );
  NAND2X0 U4490 ( .IN1(n4127), .IN2(n1239), .QN(n4125) );
  XOR2X1 U4491 ( .IN1(g481), .IN2(n4128), .Q(n4127) );
  NOR2X0 U4492 ( .IN1(n4122), .IN2(g456), .QN(n4128) );
  NAND2X0 U4493 ( .IN1(n4129), .IN2(n1646), .QN(n4122) );
  NOR2X0 U4494 ( .IN1(n1594), .IN2(g471), .QN(n4129) );
  NAND2X0 U4495 ( .IN1(n4130), .IN2(n4131), .QN(g11478) );
  NAND2X0 U4496 ( .IN1(n3591), .IN2(g339), .QN(n4131) );
  NAND2X0 U4497 ( .IN1(n3714), .IN2(n3978), .QN(n4130) );
  NAND2X0 U4498 ( .IN1(n4132), .IN2(n4133), .QN(n3978) );
  OR2X1 U4499 ( .IN1(n1239), .IN2(n2683), .Q(n4133) );
  NAND2X0 U4500 ( .IN1(n4134), .IN2(n1239), .QN(n4132) );
  XOR2X1 U4501 ( .IN1(n4135), .IN2(n1599), .Q(n4134) );
  NAND2X0 U4502 ( .IN1(n4087), .IN2(g461), .QN(n4135) );
  AND2X1 U4503 ( .IN1(n4136), .IN2(n1641), .Q(n4087) );
  NOR2X0 U4504 ( .IN1(n1606), .IN2(g466), .QN(n4136) );
  INVX0 U4505 ( .INP(n3591), .ZN(n3714) );
  NAND2X0 U4506 ( .IN1(n1647), .IN2(g750), .QN(n3591) );
  NAND2X0 U4507 ( .IN1(n4137), .IN2(n4138), .QN(g11443) );
  NAND2X0 U4508 ( .IN1(n3560), .IN2(g1275), .QN(n4138) );
  NOR2X0 U4509 ( .IN1(n3552), .IN2(n2758), .QN(n3560) );
  NAND2X0 U4510 ( .IN1(n3552), .IN2(n4020), .QN(n4137) );
  NAND2X0 U4511 ( .IN1(n4139), .IN2(n4140), .QN(n4020) );
  OR2X1 U4512 ( .IN1(n4021), .IN2(n4141), .Q(n4140) );
  XNOR2X1 U4513 ( .IN1(n4142), .IN2(n2746), .Q(n4021) );
  NAND2X0 U4514 ( .IN1(g1032), .IN2(n3936), .QN(n4142) );
  NAND2X0 U4515 ( .IN1(n4143), .IN2(n4141), .QN(n4139) );
  INVX0 U4516 ( .INP(n3553), .ZN(n4141) );
  NAND2X0 U4517 ( .IN1(n3548), .IN2(g1231), .QN(n3553) );
  NOR2X0 U4518 ( .IN1(n4144), .IN2(n2507), .QN(n3548) );
  OR2X1 U4519 ( .IN1(n2509), .IN2(n2508), .Q(n4144) );
  NAND2X0 U4520 ( .IN1(n4145), .IN2(n4146), .QN(n4143) );
  NAND2X0 U4521 ( .IN1(n1864), .IN2(g1280), .QN(n4146) );
  NAND2X0 U4522 ( .IN1(n1862), .IN2(n4147), .QN(n4145) );
  NAND2X0 U4523 ( .IN1(n1864), .IN2(n4148), .QN(n4147) );
  NAND2X0 U4524 ( .IN1(n4149), .IN2(n4150), .QN(n4148) );
  NOR2X0 U4525 ( .IN1(n4151), .IN2(n4152), .QN(n4150) );
  NAND2X0 U4526 ( .IN1(n4153), .IN2(n2636), .QN(n4152) );
  NOR2X0 U4527 ( .IN1(g1292), .IN2(g1296), .QN(n4153) );
  NAND2X0 U4528 ( .IN1(n4154), .IN2(n4155), .QN(n4151) );
  NOR2X0 U4529 ( .IN1(test_so6), .IN2(g1255), .QN(n4155) );
  NOR2X0 U4530 ( .IN1(g1260), .IN2(g1265), .QN(n4154) );
  NOR2X0 U4531 ( .IN1(n4156), .IN2(n4157), .QN(n4149) );
  NAND2X0 U4532 ( .IN1(n4158), .IN2(n2699), .QN(n4157) );
  NOR2X0 U4533 ( .IN1(g1250), .IN2(g1275), .QN(n4158) );
  NAND2X0 U4534 ( .IN1(n4159), .IN2(n2657), .QN(n4156) );
  NOR2X0 U4535 ( .IN1(g1304), .IN2(g1245), .QN(n4159) );
  AND2X1 U4536 ( .IN1(n4160), .IN2(n1610), .Q(n3552) );
  NOR2X0 U4537 ( .IN1(n2744), .IN2(n968), .QN(n4160) );
  NOR2X0 U4538 ( .IN1(n4161), .IN2(n4162), .QN(g11393) );
  NOR2X0 U4539 ( .IN1(n4163), .IN2(n4164), .QN(n4161) );
  NOR2X0 U4540 ( .IN1(n1722), .IN2(n4165), .QN(n4164) );
  NOR2X0 U4541 ( .IN1(n2965), .IN2(n2949), .QN(n4165) );
  NOR2X0 U4542 ( .IN1(n4166), .IN2(n4167), .QN(n4163) );
  NAND2X0 U4543 ( .IN1(n2949), .IN2(g981), .QN(n4167) );
  NAND2X0 U4544 ( .IN1(n4168), .IN2(n4169), .QN(n2949) );
  NOR2X0 U4545 ( .IN1(n2709), .IN2(n2708), .QN(n4169) );
  NOR2X0 U4546 ( .IN1(n1722), .IN2(n1720), .QN(n4168) );
  NOR2X0 U4547 ( .IN1(n4162), .IN2(n4170), .QN(g11392) );
  XOR2X1 U4548 ( .IN1(g981), .IN2(n4166), .Q(n4170) );
  NAND2X0 U4549 ( .IN1(n4171), .IN2(g976), .QN(n4166) );
  NOR2X0 U4550 ( .IN1(n4162), .IN2(n4172), .QN(g11391) );
  XOR2X1 U4551 ( .IN1(n2708), .IN2(n4171), .Q(n4172) );
  NOR2X0 U4552 ( .IN1(n4173), .IN2(n4174), .QN(g11380) );
  NOR2X0 U4553 ( .IN1(n4175), .IN2(g471), .QN(n4173) );
  NOR2X0 U4554 ( .IN1(n4176), .IN2(n4174), .QN(g11376) );
  NOR2X0 U4555 ( .IN1(n4177), .IN2(n4178), .QN(n4176) );
  NOR2X0 U4556 ( .IN1(n1646), .IN2(n4175), .QN(n4178) );
  AND2X1 U4557 ( .IN1(n4179), .IN2(n4180), .Q(n4175) );
  NOR2X0 U4558 ( .IN1(n4181), .IN2(n4182), .QN(n4177) );
  NAND2X0 U4559 ( .IN1(n4094), .IN2(g461), .QN(n4182) );
  NOR2X0 U4560 ( .IN1(n4174), .IN2(n4183), .QN(g11372) );
  XOR2X1 U4561 ( .IN1(g461), .IN2(n4181), .Q(n4183) );
  NAND2X0 U4562 ( .IN1(n4179), .IN2(g456), .QN(n4181) );
  NOR2X0 U4563 ( .IN1(n4162), .IN2(n4184), .QN(g11349) );
  NAND2X0 U4564 ( .IN1(n4185), .IN2(n4186), .QN(n4184) );
  INVX0 U4565 ( .INP(n4171), .ZN(n4186) );
  NOR2X0 U4566 ( .IN1(n2965), .IN2(n2709), .QN(n4171) );
  NAND2X0 U4567 ( .IN1(n2709), .IN2(n2965), .QN(n4185) );
  NAND2X0 U4568 ( .IN1(n4187), .IN2(n1420), .QN(n2965) );
  NOR2X0 U4569 ( .IN1(n16), .IN2(n4188), .QN(n4187) );
  NOR2X0 U4570 ( .IN1(n4189), .IN2(n4190), .QN(n4188) );
  NAND2X0 U4571 ( .IN1(n4191), .IN2(n4192), .QN(n4190) );
  NOR2X0 U4572 ( .IN1(n4193), .IN2(n4194), .QN(n4192) );
  NAND2X0 U4573 ( .IN1(n4195), .IN2(n4196), .QN(n4194) );
  XOR2X1 U4574 ( .IN1(n2664), .IN2(g401), .Q(n4196) );
  XOR2X1 U4575 ( .IN1(n2660), .IN2(g396), .Q(n4195) );
  XOR2X1 U4576 ( .IN1(n2663), .IN2(n2662), .Q(n4193) );
  NOR2X0 U4577 ( .IN1(n4197), .IN2(n4198), .QN(n4191) );
  XOR2X1 U4578 ( .IN1(n2686), .IN2(n2685), .Q(n4198) );
  XOR2X1 U4579 ( .IN1(n2684), .IN2(n2683), .Q(n4197) );
  NAND2X0 U4580 ( .IN1(n4199), .IN2(n4200), .QN(n4189) );
  NOR2X0 U4581 ( .IN1(n4201), .IN2(n4202), .QN(n4200) );
  NAND2X0 U4582 ( .IN1(n4203), .IN2(n4204), .QN(n4202) );
  XOR2X1 U4583 ( .IN1(n2458), .IN2(g416), .Q(n4204) );
  XNOR2X1 U4584 ( .IN1(n1681), .IN2(n4205), .Q(n4203) );
  XOR2X1 U4585 ( .IN1(n2631), .IN2(n2457), .Q(n4201) );
  NOR2X0 U4586 ( .IN1(n4206), .IN2(n4207), .QN(n4199) );
  XOR2X1 U4587 ( .IN1(n2704), .IN2(n2703), .Q(n4207) );
  XOR2X1 U4588 ( .IN1(n2702), .IN2(n2701), .Q(n4206) );
  NAND2X0 U4589 ( .IN1(n4208), .IN2(g109), .QN(n4162) );
  NAND2X0 U4590 ( .IN1(n4209), .IN2(n4933), .QN(n4208) );
  NOR2X0 U4591 ( .IN1(n2504), .IN2(n2951), .QN(n4209) );
  NOR2X0 U4592 ( .IN1(n4174), .IN2(n4210), .QN(g11340) );
  XOR2X1 U4593 ( .IN1(n1641), .IN2(n4179), .Q(n4210) );
  AND2X1 U4594 ( .IN1(n1239), .IN2(n4211), .Q(n4179) );
  NAND2X0 U4595 ( .IN1(n4180), .IN2(g471), .QN(n4211) );
  INVX0 U4596 ( .INP(n4094), .ZN(n4180) );
  NAND2X0 U4597 ( .IN1(n4212), .IN2(g461), .QN(n4094) );
  NOR2X0 U4598 ( .IN1(n1646), .IN2(n1641), .QN(n4212) );
  NAND2X0 U4599 ( .IN1(g109), .IN2(DFF_441_n1), .QN(n4174) );
  NAND2X0 U4600 ( .IN1(n4213), .IN2(n4214), .QN(g11338) );
  NAND2X0 U4601 ( .IN1(n16), .IN2(g476), .QN(n4214) );
  NAND2X0 U4602 ( .IN1(n1239), .IN2(g516), .QN(n4213) );
  NAND2X0 U4603 ( .IN1(n4215), .IN2(n4216), .QN(g11337) );
  NAND2X0 U4604 ( .IN1(n16), .IN2(g516), .QN(n4216) );
  NAND2X0 U4605 ( .IN1(n1239), .IN2(g511), .QN(n4215) );
  NAND2X0 U4606 ( .IN1(n4217), .IN2(n4218), .QN(g11336) );
  NAND2X0 U4607 ( .IN1(n16), .IN2(g511), .QN(n4218) );
  NAND2X0 U4608 ( .IN1(n1239), .IN2(g506), .QN(n4217) );
  NAND2X0 U4609 ( .IN1(n4219), .IN2(n4220), .QN(g11335) );
  NAND2X0 U4610 ( .IN1(n16), .IN2(g506), .QN(n4220) );
  NAND2X0 U4611 ( .IN1(n1239), .IN2(g501), .QN(n4219) );
  NAND2X0 U4612 ( .IN1(n4221), .IN2(n4222), .QN(g11334) );
  NAND2X0 U4613 ( .IN1(n16), .IN2(g501), .QN(n4222) );
  NAND2X0 U4614 ( .IN1(n1239), .IN2(g496), .QN(n4221) );
  NAND2X0 U4615 ( .IN1(n4223), .IN2(n4224), .QN(g11333) );
  NAND2X0 U4616 ( .IN1(n16), .IN2(g496), .QN(n4224) );
  NAND2X0 U4617 ( .IN1(n1239), .IN2(g491), .QN(n4223) );
  NAND2X0 U4618 ( .IN1(n4225), .IN2(n4226), .QN(g11332) );
  NAND2X0 U4619 ( .IN1(n16), .IN2(g491), .QN(n4226) );
  NAND2X0 U4620 ( .IN1(n1239), .IN2(g486), .QN(n4225) );
  NAND2X0 U4621 ( .IN1(n4227), .IN2(n4228), .QN(g11331) );
  NAND2X0 U4622 ( .IN1(n16), .IN2(g486), .QN(n4228) );
  NAND2X0 U4623 ( .IN1(n1239), .IN2(g481), .QN(n4227) );
  NAND2X0 U4624 ( .IN1(n4229), .IN2(n4230), .QN(g11330) );
  NAND2X0 U4625 ( .IN1(n16), .IN2(g521), .QN(n4230) );
  NAND2X0 U4626 ( .IN1(n1239), .IN2(g525), .QN(n4229) );
  NAND2X0 U4627 ( .IN1(n4231), .IN2(n4232), .QN(g11329) );
  NAND2X0 U4628 ( .IN1(n16), .IN2(g525), .QN(n4232) );
  NAND2X0 U4629 ( .IN1(n1239), .IN2(g530), .QN(n4231) );
  NAND2X0 U4630 ( .IN1(n4233), .IN2(n4234), .QN(g11328) );
  NAND2X0 U4631 ( .IN1(n16), .IN2(g530), .QN(n4234) );
  NAND2X0 U4632 ( .IN1(n1239), .IN2(g534), .QN(n4233) );
  NAND2X0 U4633 ( .IN1(n4235), .IN2(n4236), .QN(g11327) );
  NAND2X0 U4634 ( .IN1(n16), .IN2(g534), .QN(n4236) );
  NAND2X0 U4635 ( .IN1(n1239), .IN2(g538), .QN(n4235) );
  NAND2X0 U4636 ( .IN1(n4237), .IN2(n4238), .QN(g11326) );
  NAND2X0 U4637 ( .IN1(n16), .IN2(g538), .QN(n4238) );
  NAND2X0 U4638 ( .IN1(n1239), .IN2(g542), .QN(n4237) );
  NAND2X0 U4639 ( .IN1(n4239), .IN2(n4240), .QN(g11325) );
  NAND2X0 U4640 ( .IN1(n16), .IN2(g542), .QN(n4240) );
  NAND2X0 U4641 ( .IN1(n1239), .IN2(g476), .QN(n4239) );
  NAND2X0 U4642 ( .IN1(n4241), .IN2(n4242), .QN(g11324) );
  NAND2X0 U4643 ( .IN1(n16), .IN2(g481), .QN(n4242) );
  NAND2X0 U4644 ( .IN1(n3964), .IN2(n1239), .QN(n4241) );
  NAND2X0 U4645 ( .IN1(n4243), .IN2(n4244), .QN(n3964) );
  NAND2X0 U4646 ( .IN1(n1695), .IN2(g521), .QN(n4244) );
  NAND2X0 U4647 ( .IN1(n1698), .IN2(n4245), .QN(n4243) );
  NAND2X0 U4648 ( .IN1(n1695), .IN2(n4246), .QN(n4245) );
  NAND2X0 U4649 ( .IN1(n4247), .IN2(n4248), .QN(n4246) );
  NOR2X0 U4650 ( .IN1(n4249), .IN2(n4250), .QN(n4248) );
  NAND2X0 U4651 ( .IN1(n4251), .IN2(n1689), .QN(n4250) );
  NOR2X0 U4652 ( .IN1(g511), .IN2(g481), .QN(n4251) );
  NAND2X0 U4653 ( .IN1(n4252), .IN2(n4253), .QN(n4249) );
  NOR2X0 U4654 ( .IN1(g476), .IN2(g506), .QN(n4253) );
  NOR2X0 U4655 ( .IN1(g516), .IN2(g486), .QN(n4252) );
  NOR2X0 U4656 ( .IN1(n4254), .IN2(n4255), .QN(n4247) );
  NAND2X0 U4657 ( .IN1(n4256), .IN2(n2693), .QN(n4255) );
  NOR2X0 U4658 ( .IN1(g534), .IN2(g538), .QN(n4256) );
  NAND2X0 U4659 ( .IN1(n4257), .IN2(n2690), .QN(n4254) );
  NOR2X0 U4660 ( .IN1(g501), .IN2(g491), .QN(n4257) );
  NOR2X0 U4661 ( .IN1(n4258), .IN2(n4259), .QN(g11320) );
  NAND2X0 U4662 ( .IN1(n4260), .IN2(n4261), .QN(n4259) );
  NAND2X0 U4663 ( .IN1(n2616), .IN2(n4262), .QN(n4260) );
  NAND2X0 U4664 ( .IN1(n1239), .IN2(n4263), .QN(n4262) );
  NAND2X0 U4665 ( .IN1(n4264), .IN2(n4265), .QN(g11314) );
  OR2X1 U4666 ( .IN1(n4266), .IN2(n2462), .Q(n4265) );
  NAND2X0 U4667 ( .IN1(n4266), .IN2(g968), .QN(n4264) );
  NAND2X0 U4668 ( .IN1(n4267), .IN2(n4268), .QN(g11312) );
  NAND2X0 U4669 ( .IN1(n1855), .IN2(g857), .QN(n4268) );
  NAND2X0 U4670 ( .IN1(g965), .IN2(n4266), .QN(n4267) );
  NAND2X0 U4671 ( .IN1(n4269), .IN2(n4270), .QN(g11310) );
  OR2X1 U4672 ( .IN1(n4266), .IN2(n2465), .Q(n4270) );
  NAND2X0 U4673 ( .IN1(g962), .IN2(n4266), .QN(n4269) );
  NAND2X0 U4674 ( .IN1(n4271), .IN2(n4272), .QN(g11308) );
  OR2X1 U4675 ( .IN1(n4266), .IN2(n2490), .Q(n4272) );
  NAND2X0 U4676 ( .IN1(n4266), .IN2(g959), .QN(n4271) );
  NAND2X0 U4677 ( .IN1(n4273), .IN2(n4274), .QN(g11306) );
  OR2X1 U4678 ( .IN1(n4266), .IN2(n2491), .Q(n4274) );
  NAND2X0 U4679 ( .IN1(n4266), .IN2(g956), .QN(n4273) );
  NAND2X0 U4680 ( .IN1(n4275), .IN2(n4276), .QN(g11305) );
  NAND2X0 U4681 ( .IN1(n1855), .IN2(g841), .QN(n4276) );
  OR2X1 U4682 ( .IN1(n1855), .IN2(n2468), .Q(n4275) );
  NAND2X0 U4683 ( .IN1(n4277), .IN2(n4278), .QN(g11303) );
  OR2X1 U4684 ( .IN1(n4266), .IN2(n2461), .Q(n4278) );
  OR2X1 U4685 ( .IN1(n1855), .IN2(n2470), .Q(n4277) );
  NAND2X0 U4686 ( .IN1(n4279), .IN2(n4280), .QN(g11300) );
  OR2X1 U4687 ( .IN1(n4266), .IN2(n2460), .Q(n4280) );
  INVX0 U4688 ( .INP(n1855), .ZN(n4266) );
  OR2X1 U4689 ( .IN1(n1855), .IN2(n2459), .Q(n4279) );
  NAND2X0 U4690 ( .IN1(n4281), .IN2(n4282), .QN(g11298) );
  OR2X1 U4691 ( .IN1(n1855), .IN2(n2469), .Q(n4282) );
  NAND2X0 U4692 ( .IN1(n1855), .IN2(g829), .QN(n4281) );
  NAND2X0 U4693 ( .IN1(n4283), .IN2(n4284), .QN(g11294) );
  NAND2X0 U4694 ( .IN1(n4285), .IN2(n2990), .QN(n4284) );
  NOR2X0 U4695 ( .IN1(n4286), .IN2(n4287), .QN(n4285) );
  NOR2X0 U4696 ( .IN1(g1690), .IN2(n4288), .QN(n4287) );
  NAND2X0 U4697 ( .IN1(n4289), .IN2(n4290), .QN(n4288) );
  NAND2X0 U4698 ( .IN1(n4291), .IN2(n4292), .QN(n4290) );
  NAND2X0 U4699 ( .IN1(g1796), .IN2(g1801), .QN(n4292) );
  NAND2X0 U4700 ( .IN1(g1791), .IN2(g1786), .QN(n4291) );
  NAND2X0 U4701 ( .IN1(n4293), .IN2(n4294), .QN(n4289) );
  NAND2X0 U4702 ( .IN1(g1781), .IN2(g1776), .QN(n4294) );
  NAND2X0 U4703 ( .IN1(test_so5), .IN2(g1766), .QN(n4293) );
  NOR2X0 U4704 ( .IN1(n1653), .IN2(n4295), .QN(n4286) );
  NAND2X0 U4705 ( .IN1(n4296), .IN2(n4297), .QN(n4295) );
  NAND2X0 U4706 ( .IN1(n4298), .IN2(n4299), .QN(n4297) );
  NAND2X0 U4707 ( .IN1(n53), .IN2(n36), .QN(n4299) );
  NAND2X0 U4708 ( .IN1(g10664), .IN2(n38), .QN(n4298) );
  NAND2X0 U4709 ( .IN1(n4300), .IN2(n4301), .QN(n4296) );
  NAND2X0 U4710 ( .IN1(g10719), .IN2(g10720), .QN(n4301) );
  NAND2X0 U4711 ( .IN1(g10721), .IN2(g10722), .QN(n4300) );
  NOR2X0 U4712 ( .IN1(n4302), .IN2(n4303), .QN(n4283) );
  NOR2X0 U4713 ( .IN1(g1857), .IN2(n4304), .QN(n4303) );
  NAND2X0 U4714 ( .IN1(n926), .IN2(n4305), .QN(n4304) );
  NAND2X0 U4715 ( .IN1(n4306), .IN2(n4307), .QN(n4305) );
  AND2X1 U4716 ( .IN1(n3011), .IN2(n2993), .Q(n4307) );
  NOR2X0 U4717 ( .IN1(n3003), .IN2(n3005), .QN(n4306) );
  INVX0 U4718 ( .INP(n817), .ZN(n3005) );
  NAND2X0 U4719 ( .IN1(g1814), .IN2(g1828), .QN(n817) );
  INVX0 U4720 ( .INP(n822), .ZN(n3003) );
  NOR2X0 U4721 ( .IN1(n1682), .IN2(n3656), .QN(n4302) );
  NAND2X0 U4722 ( .IN1(n3230), .IN2(n346), .QN(n3656) );
  INVX0 U4723 ( .INP(n926), .ZN(n346) );
  NAND2X0 U4724 ( .IN1(n4308), .IN2(n4309), .QN(g11293) );
  NAND2X0 U4725 ( .IN1(n4310), .IN2(n3230), .QN(n4309) );
  NAND2X0 U4726 ( .IN1(n2993), .IN2(n4311), .QN(n4310) );
  NAND2X0 U4727 ( .IN1(n4312), .IN2(g1854), .QN(n4311) );
  NAND2X0 U4728 ( .IN1(n4313), .IN2(n4314), .QN(n4312) );
  NOR2X0 U4729 ( .IN1(n4315), .IN2(n4316), .QN(n4314) );
  NOR2X0 U4730 ( .IN1(n4317), .IN2(g1857), .QN(n4316) );
  XNOR2X1 U4731 ( .IN1(n1380), .IN2(n4318), .Q(n4317) );
  NOR2X0 U4732 ( .IN1(n1682), .IN2(n4319), .QN(n4315) );
  XNOR2X1 U4733 ( .IN1(n3011), .IN2(n4318), .Q(n4319) );
  NOR2X0 U4734 ( .IN1(n4320), .IN2(n3903), .QN(n4313) );
  NAND2X0 U4735 ( .IN1(n3681), .IN2(n3044), .QN(n3903) );
  INVX0 U4736 ( .INP(n2753), .ZN(n3681) );
  NAND2X0 U4737 ( .IN1(n3230), .IN2(n4321), .QN(n2753) );
  NAND2X0 U4738 ( .IN1(n1608), .IN2(g1834), .QN(n4321) );
  NOR2X0 U4739 ( .IN1(n4322), .IN2(n4323), .QN(n4320) );
  NAND2X0 U4740 ( .IN1(n1380), .IN2(n822), .QN(n4323) );
  NAND2X0 U4741 ( .IN1(n1605), .IN2(g1822), .QN(n822) );
  NAND2X0 U4742 ( .IN1(n3442), .IN2(n3011), .QN(n4322) );
  NAND2X0 U4743 ( .IN1(n1608), .IN2(g1822), .QN(n3011) );
  NAND2X0 U4744 ( .IN1(n4324), .IN2(n4325), .QN(n3442) );
  NOR2X0 U4745 ( .IN1(n1608), .IN2(g1828), .QN(n4325) );
  AND2X1 U4746 ( .IN1(n1655), .IN2(n2695), .Q(n4324) );
  NAND2X0 U4747 ( .IN1(n4326), .IN2(n1608), .QN(n2993) );
  NOR2X0 U4748 ( .IN1(n1605), .IN2(g1822), .QN(n4326) );
  NAND2X0 U4749 ( .IN1(n4327), .IN2(n2990), .QN(n4308) );
  INVX0 U4750 ( .INP(n3230), .ZN(n2990) );
  NAND2X0 U4751 ( .IN1(n4328), .IN2(n4329), .QN(n3230) );
  NOR2X0 U4752 ( .IN1(g1828), .IN2(g1834), .QN(n4329) );
  NOR2X0 U4753 ( .IN1(g1822), .IN2(g1814), .QN(n4328) );
  NAND2X0 U4754 ( .IN1(n4330), .IN2(n4331), .QN(n4327) );
  NAND2X0 U4755 ( .IN1(n4332), .IN2(g1690), .QN(n4331) );
  NAND2X0 U4756 ( .IN1(n1653), .IN2(n2734), .QN(n4330) );
  NOR2X0 U4757 ( .IN1(n4333), .IN2(n4258), .QN(g11292) );
  NOR2X0 U4758 ( .IN1(n4334), .IN2(g382), .QN(n4333) );
  NOR2X0 U4759 ( .IN1(n4335), .IN2(n4258), .QN(g11291) );
  NOR2X0 U4760 ( .IN1(n4336), .IN2(n4337), .QN(n4335) );
  NOR2X0 U4761 ( .IN1(n2615), .IN2(n4334), .QN(n4337) );
  AND2X1 U4762 ( .IN1(n4338), .IN2(n1239), .Q(n4334) );
  NOR2X0 U4763 ( .IN1(n1420), .IN2(n1385), .QN(n4338) );
  NAND2X0 U4764 ( .IN1(n4339), .IN2(g374), .QN(n1385) );
  NOR2X0 U4765 ( .IN1(n4261), .IN2(n4340), .QN(n4336) );
  OR2X1 U4766 ( .IN1(n4339), .IN2(n2617), .Q(n4340) );
  NOR2X0 U4767 ( .IN1(n2616), .IN2(n2615), .QN(n4339) );
  NOR2X0 U4768 ( .IN1(n4258), .IN2(n4341), .QN(g11290) );
  XOR2X1 U4769 ( .IN1(g374), .IN2(n4261), .Q(n4341) );
  NAND2X0 U4770 ( .IN1(n4342), .IN2(n1239), .QN(n4261) );
  NOR2X0 U4771 ( .IN1(n2616), .IN2(n1420), .QN(n4342) );
  NAND2X0 U4772 ( .IN1(n2504), .IN2(g109), .QN(n4258) );
  NAND2X0 U4773 ( .IN1(n4343), .IN2(n4344), .QN(g11270) );
  NAND2X0 U4774 ( .IN1(n16), .IN2(g421), .QN(n4344) );
  NAND2X0 U4775 ( .IN1(n1239), .IN2(g416), .QN(n4343) );
  NAND2X0 U4776 ( .IN1(n4345), .IN2(n4346), .QN(g11269) );
  NAND2X0 U4777 ( .IN1(n16), .IN2(g416), .QN(n4346) );
  NAND2X0 U4778 ( .IN1(n1239), .IN2(g411), .QN(n4345) );
  NAND2X0 U4779 ( .IN1(n4347), .IN2(n4348), .QN(g11268) );
  NAND2X0 U4780 ( .IN1(n16), .IN2(g411), .QN(n4348) );
  NAND2X0 U4781 ( .IN1(n1239), .IN2(g406), .QN(n4347) );
  NAND2X0 U4782 ( .IN1(n4349), .IN2(n4350), .QN(g11267) );
  NAND2X0 U4783 ( .IN1(n16), .IN2(g406), .QN(n4350) );
  NAND2X0 U4784 ( .IN1(n1239), .IN2(g401), .QN(n4349) );
  NAND2X0 U4785 ( .IN1(n4351), .IN2(n4352), .QN(g11266) );
  NAND2X0 U4786 ( .IN1(n16), .IN2(g401), .QN(n4352) );
  NAND2X0 U4787 ( .IN1(n1239), .IN2(g396), .QN(n4351) );
  NAND2X0 U4788 ( .IN1(n4353), .IN2(n4354), .QN(g11265) );
  NAND2X0 U4789 ( .IN1(n16), .IN2(g396), .QN(n4354) );
  NAND2X0 U4790 ( .IN1(n1239), .IN2(g391), .QN(n4353) );
  NAND2X0 U4791 ( .IN1(n4355), .IN2(n4356), .QN(g11264) );
  NAND2X0 U4792 ( .IN1(n16), .IN2(g391), .QN(n4356) );
  NAND2X0 U4793 ( .IN1(n1239), .IN2(g386), .QN(n4355) );
  NAND2X0 U4794 ( .IN1(n4357), .IN2(n4358), .QN(g11263) );
  NAND2X0 U4795 ( .IN1(n16), .IN2(g386), .QN(n4358) );
  NAND2X0 U4796 ( .IN1(n1239), .IN2(g426), .QN(n4357) );
  NAND2X0 U4797 ( .IN1(n4359), .IN2(n4360), .QN(g11262) );
  NAND2X0 U4798 ( .IN1(n16), .IN2(g431), .QN(n4360) );
  NAND2X0 U4799 ( .IN1(n1239), .IN2(g435), .QN(n4359) );
  NAND2X0 U4800 ( .IN1(n4361), .IN2(n4362), .QN(g11261) );
  NAND2X0 U4801 ( .IN1(n16), .IN2(g435), .QN(n4362) );
  NAND2X0 U4802 ( .IN1(n1239), .IN2(g440), .QN(n4361) );
  NAND2X0 U4803 ( .IN1(n4363), .IN2(n4364), .QN(g11260) );
  NAND2X0 U4804 ( .IN1(n16), .IN2(g440), .QN(n4364) );
  NAND2X0 U4805 ( .IN1(n1239), .IN2(g444), .QN(n4363) );
  NAND2X0 U4806 ( .IN1(n4365), .IN2(n4366), .QN(g11259) );
  NAND2X0 U4807 ( .IN1(n16), .IN2(g444), .QN(n4366) );
  NAND2X0 U4808 ( .IN1(n1239), .IN2(g448), .QN(n4365) );
  NAND2X0 U4809 ( .IN1(n4367), .IN2(n4368), .QN(g11258) );
  NAND2X0 U4810 ( .IN1(n16), .IN2(g448), .QN(n4368) );
  NAND2X0 U4811 ( .IN1(n1239), .IN2(g452), .QN(n4367) );
  NAND2X0 U4812 ( .IN1(n4369), .IN2(n4370), .QN(g11257) );
  NAND2X0 U4813 ( .IN1(n16), .IN2(g452), .QN(n4370) );
  NAND2X0 U4814 ( .IN1(n1239), .IN2(g421), .QN(n4369) );
  NAND2X0 U4815 ( .IN1(n4371), .IN2(n4372), .QN(g11256) );
  NAND2X0 U4816 ( .IN1(n16), .IN2(g426), .QN(n4372) );
  OR2X1 U4817 ( .IN1(n4205), .IN2(n16), .Q(n4371) );
  INVX0 U4818 ( .INP(n1239), .ZN(n16) );
  NOR2X0 U4819 ( .IN1(n4375), .IN2(n4376), .QN(n4374) );
  NAND2X0 U4820 ( .IN1(n2462), .IN2(n2461), .QN(n4376) );
  NAND2X0 U4821 ( .IN1(n4377), .IN2(n2460), .QN(n4375) );
  NOR2X0 U4822 ( .IN1(n4378), .IN2(g829), .QN(n4377) );
  NOR2X0 U4823 ( .IN1(n4379), .IN2(n4380), .QN(n4378) );
  OR2X1 U4824 ( .IN1(n4381), .IN2(n4382), .Q(n4380) );
  NOR2X0 U4825 ( .IN1(n2760), .IN2(n4383), .QN(n4379) );
  NOR2X0 U4826 ( .IN1(n4384), .IN2(n4385), .QN(n4383) );
  NOR2X0 U4827 ( .IN1(n4386), .IN2(n4387), .QN(n4373) );
  NAND2X0 U4828 ( .IN1(n2491), .IN2(n2490), .QN(n4387) );
  NAND2X0 U4829 ( .IN1(n4388), .IN2(n2465), .QN(n4386) );
  NOR2X0 U4830 ( .IN1(g841), .IN2(g857), .QN(n4388) );
  NAND2X0 U4831 ( .IN1(n4389), .IN2(n4390), .QN(n4205) );
  NAND2X0 U4832 ( .IN1(n1681), .IN2(n4263), .QN(n4390) );
  INVX0 U4833 ( .INP(n1420), .ZN(n4263) );
  NAND2X0 U4834 ( .IN1(n4391), .IN2(n1420), .QN(n4389) );
  NAND2X0 U4835 ( .IN1(n4392), .IN2(n4393), .QN(n4391) );
  NAND2X0 U4836 ( .IN1(g431), .IN2(g435), .QN(n4393) );
  NAND2X0 U4837 ( .IN1(n4394), .IN2(n1878), .QN(n4392) );
  NOR2X0 U4838 ( .IN1(n4395), .IN2(g431), .QN(n4394) );
  NOR2X0 U4839 ( .IN1(n4396), .IN2(n4397), .QN(n4395) );
  NAND2X0 U4840 ( .IN1(n4398), .IN2(n4399), .QN(n4397) );
  NOR2X0 U4841 ( .IN1(g421), .IN2(n4400), .QN(n4399) );
  NAND2X0 U4842 ( .IN1(n2665), .IN2(n2663), .QN(n4400) );
  NOR2X0 U4843 ( .IN1(g391), .IN2(n4401), .QN(n4398) );
  NAND2X0 U4844 ( .IN1(n2701), .IN2(n2686), .QN(n4401) );
  NAND2X0 U4845 ( .IN1(n4402), .IN2(n4403), .QN(n4396) );
  NOR2X0 U4846 ( .IN1(n4404), .IN2(n4405), .QN(n4403) );
  NAND2X0 U4847 ( .IN1(n2640), .IN2(n2639), .QN(n4405) );
  NAND2X0 U4848 ( .IN1(n2631), .IN2(n2638), .QN(n4404) );
  NOR2X0 U4849 ( .IN1(g396), .IN2(n4406), .QN(n4402) );
  NAND2X0 U4850 ( .IN1(n2642), .IN2(n2641), .QN(n4406) );
  NOR2X0 U4851 ( .IN1(n4407), .IN2(n4408), .QN(g11206) );
  XOR2X1 U4852 ( .IN1(n4409), .IN2(n4407), .Q(g11163) );
  NAND2X0 U4853 ( .IN1(n4410), .IN2(n4411), .QN(n4407) );
  NAND2X0 U4854 ( .IN1(g5392), .IN2(n38), .QN(n4411) );
  NOR2X0 U4855 ( .IN1(n3913), .IN2(n2759), .QN(g5392) );
  NAND2X0 U4856 ( .IN1(g1765), .IN2(g1610), .QN(n3913) );
  NOR2X0 U4857 ( .IN1(n4412), .IN2(n4413), .QN(n4410) );
  NOR2X0 U4858 ( .IN1(n4414), .IN2(n3956), .QN(n4413) );
  NAND2X0 U4859 ( .IN1(n4415), .IN2(n4935), .QN(n3956) );
  NOR2X0 U4860 ( .IN1(n2482), .IN2(n2760), .QN(n4415) );
  NOR2X0 U4861 ( .IN1(n2757), .IN2(n4416), .QN(n4412) );
  NOR2X0 U4862 ( .IN1(n4417), .IN2(n4418), .QN(n4416) );
  NAND2X0 U4863 ( .IN1(n4419), .IN2(n4420), .QN(n4418) );
  OR2X1 U4864 ( .IN1(n4421), .IN2(n4949), .Q(n4420) );
  NAND2X0 U4865 ( .IN1(n2483), .IN2(n53), .QN(n4419) );
  NOR2X0 U4866 ( .IN1(n4936), .IN2(n4422), .QN(n4417) );
  NAND2X0 U4867 ( .IN1(n4423), .IN2(n4424), .QN(g10936) );
  NAND2X0 U4868 ( .IN1(n1054), .IN2(g1811), .QN(n4424) );
  NAND2X0 U4869 ( .IN1(n1391), .IN2(n256), .QN(n4423) );
  NAND2X0 U4870 ( .IN1(n4425), .IN2(n4426), .QN(n1391) );
  NOR2X0 U4871 ( .IN1(g10721), .IN2(n4427), .QN(n4426) );
  NOR2X0 U4872 ( .IN1(g46), .IN2(n4428), .QN(n4427) );
  NOR2X0 U4873 ( .IN1(n4385), .IN2(n4421), .QN(n4425) );
  NAND2X0 U4874 ( .IN1(n4429), .IN2(n4430), .QN(g10898) );
  OR2X1 U4875 ( .IN1(n3306), .IN2(n2483), .Q(n4430) );
  NAND2X0 U4876 ( .IN1(n4431), .IN2(n3306), .QN(n4429) );
  NAND2X0 U4877 ( .IN1(n4432), .IN2(n3936), .QN(n4431) );
  NAND2X0 U4878 ( .IN1(n4069), .IN2(n4433), .QN(n3936) );
  NAND2X0 U4879 ( .IN1(n2958), .IN2(n2956), .QN(n4069) );
  INVX0 U4880 ( .INP(n4428), .ZN(n2958) );
  NAND2X0 U4881 ( .IN1(n4434), .IN2(n2960), .QN(n4428) );
  INVX0 U4882 ( .INP(n2957), .ZN(n2960) );
  NAND2X0 U4883 ( .IN1(n4435), .IN2(n4436), .QN(n2957) );
  NOR2X0 U4884 ( .IN1(g44), .IN2(n4437), .QN(n4436) );
  NAND2X0 U4885 ( .IN1(n4438), .IN2(n4439), .QN(n4437) );
  AND2X1 U4886 ( .IN1(n4440), .IN2(n2984), .Q(n4435) );
  NOR2X0 U4887 ( .IN1(g47), .IN2(n2961), .QN(n4434) );
  XOR2X1 U4888 ( .IN1(n4441), .IN2(n4442), .Q(n4432) );
  XOR2X1 U4889 ( .IN1(n4443), .IN2(n4444), .Q(n4442) );
  XOR2X1 U4890 ( .IN1(n4445), .IN2(n4446), .Q(n4444) );
  XOR2X1 U4891 ( .IN1(n2593), .IN2(n1871), .Q(n4446) );
  XOR2X1 U4892 ( .IN1(n2658), .IN2(n2618), .Q(n4445) );
  XOR2X1 U4893 ( .IN1(n4447), .IN2(n4448), .Q(n4443) );
  XOR2X1 U4894 ( .IN1(n2700), .IN2(n2698), .Q(n4448) );
  XOR2X1 U4895 ( .IN1(test_so2), .IN2(n2746), .Q(n4447) );
  XNOR2X1 U4896 ( .IN1(n2619), .IN2(test_so8), .Q(n4441) );
  NAND2X0 U4897 ( .IN1(n4449), .IN2(n4450), .QN(g10866) );
  NAND2X0 U4898 ( .IN1(n968), .IN2(g1684), .QN(n4450) );
  NAND2X0 U4899 ( .IN1(n4451), .IN2(n4452), .QN(g10865) );
  NAND2X0 U4900 ( .IN1(n3800), .IN2(g1669), .QN(n4452) );
  NAND2X0 U4901 ( .IN1(n4453), .IN2(n3799), .QN(n4451) );
  NOR2X0 U4902 ( .IN1(n4454), .IN2(n4455), .QN(n4453) );
  NOR2X0 U4903 ( .IN1(n2758), .IN2(g10722), .QN(n4454) );
  NAND2X0 U4904 ( .IN1(n4456), .IN2(n4457), .QN(g10864) );
  NAND2X0 U4905 ( .IN1(n968), .IN2(g1681), .QN(n4457) );
  NAND2X0 U4906 ( .IN1(n4458), .IN2(n4459), .QN(g10863) );
  NAND2X0 U4907 ( .IN1(n3800), .IN2(g1666), .QN(n4459) );
  NAND2X0 U4908 ( .IN1(n4460), .IN2(n3799), .QN(n4458) );
  NOR2X0 U4909 ( .IN1(n4461), .IN2(n4462), .QN(n4460) );
  NOR2X0 U4910 ( .IN1(n4382), .IN2(g1718), .QN(n4462) );
  NAND2X0 U4911 ( .IN1(n4463), .IN2(n4464), .QN(g10862) );
  NAND2X0 U4912 ( .IN1(n968), .IN2(g1678), .QN(n4464) );
  NAND2X0 U4913 ( .IN1(n4465), .IN2(n4466), .QN(g10861) );
  NAND2X0 U4914 ( .IN1(n3800), .IN2(g1663), .QN(n4466) );
  NAND2X0 U4915 ( .IN1(n3799), .IN2(n4467), .QN(n4465) );
  NAND2X0 U4916 ( .IN1(n4468), .IN2(n4469), .QN(g10860) );
  NAND2X0 U4917 ( .IN1(n968), .IN2(g1675), .QN(n4469) );
  NAND2X0 U4918 ( .IN1(n4470), .IN2(n4471), .QN(g10859) );
  NAND2X0 U4919 ( .IN1(n3800), .IN2(g1660), .QN(n4471) );
  NAND2X0 U4920 ( .IN1(n3799), .IN2(n4472), .QN(n4470) );
  NAND2X0 U4921 ( .IN1(n4473), .IN2(n4474), .QN(g10858) );
  NAND2X0 U4922 ( .IN1(n968), .IN2(g1672), .QN(n4474) );
  NAND2X0 U4923 ( .IN1(n4475), .IN2(n4476), .QN(g10855) );
  NAND2X0 U4924 ( .IN1(n968), .IN2(g549), .QN(n4476) );
  NAND2X0 U4925 ( .IN1(n4467), .IN2(n3306), .QN(n4475) );
  NAND2X0 U4926 ( .IN1(n4477), .IN2(n1611), .QN(n4467) );
  NOR2X0 U4927 ( .IN1(n4478), .IN2(n4479), .QN(n4477) );
  NOR2X0 U4928 ( .IN1(n4480), .IN2(n3515), .QN(n4479) );
  AND2X1 U4929 ( .IN1(n4481), .IN2(n3818), .Q(n3515) );
  NAND2X0 U4930 ( .IN1(g18), .IN2(g192), .QN(n3818) );
  NAND2X0 U4931 ( .IN1(n2967), .IN2(g1512), .QN(n4481) );
  NOR2X0 U4932 ( .IN1(n4461), .IN2(n4482), .QN(n4478) );
  NAND2X0 U4933 ( .IN1(g109), .IN2(g10720), .QN(n4482) );
  NAND2X0 U4934 ( .IN1(n2754), .IN2(n4409), .QN(g10801) );
  INVX0 U4935 ( .INP(n2747), .ZN(n4409) );
  XOR2X1 U4936 ( .IN1(n4483), .IN2(n4484), .Q(n2747) );
  XOR2X1 U4937 ( .IN1(n4485), .IN2(n4486), .Q(n4484) );
  NAND2X0 U4938 ( .IN1(n4937), .IN2(n4487), .QN(n4486) );
  NAND2X0 U4939 ( .IN1(n4488), .IN2(n4384), .QN(n4485) );
  NAND2X0 U4940 ( .IN1(n4489), .IN2(n4422), .QN(n4384) );
  NOR2X0 U4941 ( .IN1(n53), .IN2(n38), .QN(n4489) );
  NOR2X0 U4942 ( .IN1(n4490), .IN2(n4491), .QN(n4488) );
  NOR2X0 U4943 ( .IN1(g10664), .IN2(n4492), .QN(n4491) );
  NAND2X0 U4944 ( .IN1(n53), .IN2(n38), .QN(n4492) );
  NOR2X0 U4945 ( .IN1(n4422), .IN2(n4493), .QN(n4490) );
  XOR2X1 U4946 ( .IN1(n53), .IN2(n4433), .Q(n4493) );
  INVX0 U4947 ( .INP(g10664), .ZN(n4422) );
  XNOR2X1 U4948 ( .IN1(n4494), .IN2(n1858), .Q(n4483) );
  XNOR2X1 U4949 ( .IN1(g10722), .IN2(g10721), .Q(n1858) );
  NAND2X0 U4950 ( .IN1(n4495), .IN2(n4385), .QN(n4494) );
  NAND2X0 U4951 ( .IN1(n4496), .IN2(n4332), .QN(n4385) );
  NOR2X0 U4952 ( .IN1(n36), .IN2(g10720), .QN(n4496) );
  NOR2X0 U4953 ( .IN1(n4497), .IN2(n4498), .QN(n4495) );
  NOR2X0 U4954 ( .IN1(g10720), .IN2(n4499), .QN(n4498) );
  NAND2X0 U4955 ( .IN1(g10719), .IN2(n36), .QN(n4499) );
  NOR2X0 U4956 ( .IN1(n4500), .IN2(n4501), .QN(n4497) );
  XOR2X1 U4957 ( .IN1(n36), .IN2(n4332), .Q(n4501) );
  NAND2X0 U4958 ( .IN1(n4502), .IN2(n4503), .QN(g10800) );
  NAND2X0 U4959 ( .IN1(n968), .IN2(g575), .QN(n4503) );
  NAND2X0 U4960 ( .IN1(n4472), .IN2(n3306), .QN(n4502) );
  NAND2X0 U4961 ( .IN1(n4504), .IN2(n1611), .QN(n4472) );
  NOR2X0 U4962 ( .IN1(n4505), .IN2(n4506), .QN(n4504) );
  NOR2X0 U4963 ( .IN1(n4480), .IN2(n3510), .QN(n4506) );
  AND2X1 U4964 ( .IN1(n4507), .IN2(n3820), .Q(n3510) );
  NAND2X0 U4965 ( .IN1(g18), .IN2(g248), .QN(n3820) );
  NAND2X0 U4966 ( .IN1(n2967), .IN2(g1636), .QN(n4507) );
  NOR2X0 U4967 ( .IN1(n4461), .IN2(n4508), .QN(n4505) );
  NOR2X0 U4968 ( .IN1(n2759), .IN2(g10719), .QN(n4508) );
  NAND2X0 U4969 ( .IN1(n4509), .IN2(n4510), .QN(g10799) );
  NAND2X0 U4970 ( .IN1(n968), .IN2(g566), .QN(n4510) );
  NAND2X0 U4971 ( .IN1(n4449), .IN2(n4511), .QN(g10798) );
  NAND2X0 U4972 ( .IN1(n968), .IN2(g563), .QN(n4511) );
  NAND2X0 U4973 ( .IN1(n4512), .IN2(n3306), .QN(n4449) );
  NAND2X0 U4974 ( .IN1(n4513), .IN2(n4514), .QN(n4512) );
  NAND2X0 U4975 ( .IN1(n4461), .IN2(n3513), .QN(n4514) );
  NAND2X0 U4976 ( .IN1(n3327), .IN2(n4515), .QN(n3513) );
  NAND2X0 U4977 ( .IN1(n2967), .IN2(g1624), .QN(n4515) );
  NAND2X0 U4978 ( .IN1(g18), .IN2(g225), .QN(n3327) );
  NAND2X0 U4979 ( .IN1(n1404), .IN2(n4318), .QN(n4513) );
  NAND2X0 U4980 ( .IN1(n4456), .IN2(n4516), .QN(g10797) );
  NAND2X0 U4981 ( .IN1(n968), .IN2(g560), .QN(n4516) );
  NAND2X0 U4982 ( .IN1(n4517), .IN2(n3306), .QN(n4456) );
  NAND2X0 U4983 ( .IN1(n4518), .IN2(n4519), .QN(n4517) );
  NAND2X0 U4984 ( .IN1(n4461), .IN2(n3508), .QN(n4519) );
  NAND2X0 U4985 ( .IN1(n3317), .IN2(n4520), .QN(n3508) );
  NAND2X0 U4986 ( .IN1(n2967), .IN2(g1621), .QN(n4520) );
  OR2X1 U4987 ( .IN1(n2967), .IN2(n2514), .Q(n3317) );
  NAND2X0 U4988 ( .IN1(n1404), .IN2(n4381), .QN(n4518) );
  NAND2X0 U4989 ( .IN1(n4463), .IN2(n4521), .QN(g10795) );
  NAND2X0 U4990 ( .IN1(n968), .IN2(g557), .QN(n4521) );
  NAND2X0 U4991 ( .IN1(n4522), .IN2(n3306), .QN(n4463) );
  NAND2X0 U4992 ( .IN1(n4523), .IN2(n4524), .QN(n4522) );
  NAND2X0 U4993 ( .IN1(n4461), .IN2(n3500), .QN(n4524) );
  NAND2X0 U4994 ( .IN1(n3364), .IN2(n4525), .QN(n3500) );
  NAND2X0 U4995 ( .IN1(n2967), .IN2(g1615), .QN(n4525) );
  OR2X1 U4996 ( .IN1(n2967), .IN2(n2513), .Q(n3364) );
  NAND2X0 U4997 ( .IN1(n1404), .IN2(n4382), .QN(n4523) );
  NAND2X0 U4998 ( .IN1(n4468), .IN2(n4526), .QN(g10793) );
  NAND2X0 U4999 ( .IN1(n968), .IN2(g554), .QN(n4526) );
  NAND2X0 U5000 ( .IN1(n4527), .IN2(n4528), .QN(n4468) );
  NAND2X0 U5001 ( .IN1(n4461), .IN2(n3496), .QN(n4528) );
  AND2X1 U5002 ( .IN1(n3352), .IN2(n4529), .Q(n3496) );
  NAND2X0 U5003 ( .IN1(n2967), .IN2(g1639), .QN(n4529) );
  NAND2X0 U5004 ( .IN1(g18), .IN2(g207), .QN(n3352) );
  NOR2X0 U5005 ( .IN1(n968), .IN2(n4530), .QN(n4527) );
  NOR2X0 U5006 ( .IN1(n4455), .IN2(n4531), .QN(n4530) );
  NAND2X0 U5007 ( .IN1(n4500), .IN2(g109), .QN(n4531) );
  NAND2X0 U5008 ( .IN1(n4473), .IN2(n4532), .QN(g10791) );
  NAND2X0 U5009 ( .IN1(n968), .IN2(g546), .QN(n4532) );
  NAND2X0 U5010 ( .IN1(n4533), .IN2(n3306), .QN(n4473) );
  NAND2X0 U5011 ( .IN1(n4534), .IN2(n4535), .QN(n4533) );
  NAND2X0 U5012 ( .IN1(n4536), .IN2(n1404), .QN(n4535) );
  NAND2X0 U5013 ( .IN1(n4461), .IN2(n3517), .QN(n4534) );
  NAND2X0 U5014 ( .IN1(n3340), .IN2(n4537), .QN(n3517) );
  NAND2X0 U5015 ( .IN1(n2967), .IN2(g1618), .QN(n4537) );
  OR2X1 U5016 ( .IN1(n2967), .IN2(n2511), .Q(n3340) );
  NOR2X0 U5017 ( .IN1(n4952), .IN2(n256), .QN(g10785) );
  NOR2X0 U5018 ( .IN1(n4953), .IN2(n256), .QN(g10784) );
  NOR2X0 U5019 ( .IN1(n4954), .IN2(n256), .QN(g10782) );
  NOR2X0 U5020 ( .IN1(n4955), .IN2(n256), .QN(g10780) );
  INVX0 U5021 ( .INP(n1054), .ZN(n256) );
  NAND2X0 U5022 ( .IN1(n2745), .IN2(g1696), .QN(n1054) );
  NAND2X0 U5023 ( .IN1(n4509), .IN2(n4538), .QN(g10776) );
  NAND2X0 U5024 ( .IN1(n968), .IN2(g1687), .QN(n4538) );
  NAND2X0 U5025 ( .IN1(n4539), .IN2(n3306), .QN(n4509) );
  NAND2X0 U5026 ( .IN1(n4540), .IN2(n4541), .QN(n4539) );
  NAND2X0 U5027 ( .IN1(n1404), .IN2(n53), .QN(n4541) );
  INVX0 U5028 ( .INP(n4070), .ZN(n53) );
  NOR2X0 U5029 ( .IN1(n1450), .IN2(n4542), .QN(n4540) );
  NOR2X0 U5030 ( .IN1(n3519), .IN2(n4480), .QN(n4542) );
  NAND2X0 U5031 ( .IN1(n4543), .IN2(n4544), .QN(n3519) );
  NAND2X0 U5032 ( .IN1(n2582), .IN2(n2967), .QN(n4544) );
  NAND2X0 U5033 ( .IN1(g18), .IN2(n2677), .QN(n4543) );
  NAND2X0 U5034 ( .IN1(n4545), .IN2(n4546), .QN(g10773) );
  NAND2X0 U5035 ( .IN1(n3902), .IN2(n4382), .QN(n4546) );
  OR2X1 U5036 ( .IN1(n3902), .IN2(n2486), .Q(n4545) );
  NAND2X0 U5037 ( .IN1(n4547), .IN2(n4548), .QN(g10771) );
  OR2X1 U5038 ( .IN1(n3902), .IN2(n2484), .Q(n4548) );
  NAND2X0 U5039 ( .IN1(n4549), .IN2(n3902), .QN(n4547) );
  NOR2X0 U5040 ( .IN1(n4500), .IN2(n2757), .QN(n4549) );
  NAND2X0 U5041 ( .IN1(n4550), .IN2(n4551), .QN(g10770) );
  OR2X1 U5042 ( .IN1(n3902), .IN2(n2487), .Q(n4551) );
  NAND2X0 U5043 ( .IN1(n4536), .IN2(n3902), .QN(n4550) );
  NOR2X0 U5044 ( .IN1(n4332), .IN2(n2758), .QN(n4536) );
  NAND2X0 U5045 ( .IN1(n4552), .IN2(n4553), .QN(g10767) );
  NAND2X0 U5046 ( .IN1(n3800), .IN2(g1657), .QN(n4553) );
  NAND2X0 U5047 ( .IN1(n3799), .IN2(n4554), .QN(n4552) );
  NAND2X0 U5048 ( .IN1(n4555), .IN2(n4556), .QN(g10765) );
  NAND2X0 U5049 ( .IN1(n3800), .IN2(g1654), .QN(n4556) );
  INVX0 U5050 ( .INP(n3799), .ZN(n3800) );
  NAND2X0 U5051 ( .IN1(n3799), .IN2(n4557), .QN(n4555) );
  NOR2X0 U5052 ( .IN1(g1696), .IN2(n2745), .QN(n3799) );
  NAND2X0 U5053 ( .IN1(n4558), .IN2(n4559), .QN(g10718) );
  NAND2X0 U5054 ( .IN1(n968), .IN2(g572), .QN(n4559) );
  NAND2X0 U5055 ( .IN1(n4554), .IN2(n3306), .QN(n4558) );
  NAND2X0 U5056 ( .IN1(n4560), .IN2(n1611), .QN(n4554) );
  NOR2X0 U5057 ( .IN1(n4561), .IN2(n4562), .QN(n4560) );
  NOR2X0 U5058 ( .IN1(n4480), .IN2(n3502), .QN(n4562) );
  AND2X1 U5059 ( .IN1(n4563), .IN2(n3822), .Q(n3502) );
  NAND2X0 U5060 ( .IN1(g18), .IN2(g243), .QN(n3822) );
  NAND2X0 U5061 ( .IN1(n2967), .IN2(g1633), .QN(n4563) );
  NOR2X0 U5062 ( .IN1(n4461), .IN2(n4564), .QN(n4561) );
  NAND2X0 U5063 ( .IN1(g109), .IN2(g10664), .QN(n4564) );
  INVX0 U5064 ( .INP(n4480), .ZN(n4461) );
  NAND2X0 U5065 ( .IN1(n4565), .IN2(n4566), .QN(g10717) );
  NAND2X0 U5066 ( .IN1(n968), .IN2(g569), .QN(n4566) );
  NAND2X0 U5067 ( .IN1(n4557), .IN2(n3306), .QN(n4565) );
  INVX0 U5068 ( .INP(n968), .ZN(n3306) );
  NAND2X0 U5069 ( .IN1(n2745), .IN2(n4567), .QN(n968) );
  NAND2X0 U5070 ( .IN1(n4568), .IN2(n4569), .QN(n4557) );
  NAND2X0 U5071 ( .IN1(n1404), .IN2(n38), .QN(n4569) );
  INVX0 U5072 ( .INP(n4455), .ZN(n1404) );
  NAND2X0 U5073 ( .IN1(n1611), .IN2(n4480), .QN(n4455) );
  NOR2X0 U5074 ( .IN1(n1450), .IN2(n4570), .QN(n4568) );
  NOR2X0 U5075 ( .IN1(n3521), .IN2(n4480), .QN(n4570) );
  NAND2X0 U5076 ( .IN1(n4951), .IN2(n1611), .QN(n4480) );
  NAND2X0 U5077 ( .IN1(n4571), .IN2(n4572), .QN(n3521) );
  NAND2X0 U5078 ( .IN1(n2579), .IN2(n2967), .QN(n4572) );
  INVX0 U5079 ( .INP(g18), .ZN(n2967) );
  NAND2X0 U5080 ( .IN1(g18), .IN2(n2678), .QN(n4571) );
  NAND2X0 U5081 ( .IN1(n4573), .IN2(n4574), .QN(g10711) );
  OR2X1 U5082 ( .IN1(n3902), .IN2(n2485), .Q(n4574) );
  NAND2X0 U5083 ( .IN1(n3902), .IN2(n4318), .QN(n4573) );
  NAND2X0 U5084 ( .IN1(g109), .IN2(n4414), .QN(n4318) );
  NAND2X0 U5085 ( .IN1(n4575), .IN2(n4576), .QN(g10707) );
  NAND2X0 U5086 ( .IN1(n3902), .IN2(n4381), .QN(n4576) );
  OR2X1 U5087 ( .IN1(n3902), .IN2(n2467), .Q(n4575) );
  NOR2X0 U5088 ( .IN1(n4567), .IN2(n2745), .QN(n3902) );
  INVX0 U5089 ( .INP(g1696), .ZN(n4567) );
  NAND2X0 U5090 ( .IN1(n4577), .IN2(n4578), .QN(g10664) );
  NOR2X0 U5091 ( .IN1(n4579), .IN2(n4580), .QN(n4578) );
  NAND2X0 U5092 ( .IN1(n4581), .IN2(n4582), .QN(n4580) );
  NAND2X0 U5093 ( .IN1(n4583), .IN2(g1741), .QN(n4582) );
  NAND2X0 U5094 ( .IN1(n3040), .IN2(n4487), .QN(n4581) );
  NAND2X0 U5095 ( .IN1(n4584), .IN2(n4585), .QN(n4579) );
  NAND2X0 U5096 ( .IN1(g919), .IN2(n4586), .QN(n4585) );
  NOR2X0 U5097 ( .IN1(n4587), .IN2(n4588), .QN(n4584) );
  NOR2X0 U5098 ( .IN1(n2459), .IN2(n4589), .QN(n4588) );
  NOR2X0 U5099 ( .IN1(n2565), .IN2(n4590), .QN(n4587) );
  NOR2X0 U5100 ( .IN1(n4591), .IN2(n4592), .QN(n4577) );
  NAND2X0 U5101 ( .IN1(n4593), .IN2(n4594), .QN(n4592) );
  NAND2X0 U5102 ( .IN1(g1191), .IN2(n4595), .QN(n4594) );
  NOR2X0 U5103 ( .IN1(n4596), .IN2(n4597), .QN(n4593) );
  AND2X1 U5104 ( .IN1(n4598), .IN2(test_so9), .Q(n4597) );
  NOR2X0 U5105 ( .IN1(n4598), .IN2(n4599), .QN(n4596) );
  NAND2X0 U5106 ( .IN1(n1478), .IN2(n4600), .QN(n4599) );
  NAND2X0 U5107 ( .IN1(n4601), .IN2(n4602), .QN(n4591) );
  NAND2X0 U5108 ( .IN1(n1485), .IN2(g1589), .QN(n4602) );
  NAND2X0 U5109 ( .IN1(n1486), .IN2(g1546), .QN(n4601) );
  INVX0 U5110 ( .INP(n4408), .ZN(g10628) );
  NAND2X0 U5111 ( .IN1(n4603), .IN2(n4604), .QN(n4408) );
  NAND2X0 U5112 ( .IN1(n4605), .IN2(g109), .QN(n4604) );
  OR2X1 U5113 ( .IN1(n4606), .IN2(n4607), .Q(n4605) );
  NAND2X0 U5114 ( .IN1(n4608), .IN2(n4609), .QN(n4607) );
  NAND2X0 U5115 ( .IN1(g877), .IN2(g10719), .QN(n4609) );
  NAND2X0 U5116 ( .IN1(g881), .IN2(g10720), .QN(n4608) );
  NAND2X0 U5117 ( .IN1(n4610), .IN2(n4611), .QN(n4606) );
  NAND2X0 U5118 ( .IN1(n2951), .IN2(n36), .QN(n4611) );
  INVX0 U5119 ( .INP(n4414), .ZN(n36) );
  AND2X1 U5120 ( .IN1(n2480), .IN2(g3007), .Q(n2951) );
  NAND2X0 U5121 ( .IN1(n4381), .IN2(n3064), .QN(n4610) );
  INVX0 U5122 ( .INP(n4421), .ZN(n4381) );
  NAND2X0 U5123 ( .IN1(g10722), .IN2(g109), .QN(n4421) );
  NAND2X0 U5124 ( .IN1(n4612), .IN2(n4613), .QN(g10722) );
  NOR2X0 U5125 ( .IN1(n4614), .IN2(n4615), .QN(n4613) );
  NAND2X0 U5126 ( .IN1(n4616), .IN2(n4617), .QN(n4615) );
  NOR2X0 U5127 ( .IN1(n4618), .IN2(n4619), .QN(n4617) );
  NAND2X0 U5128 ( .IN1(n4620), .IN2(n4621), .QN(n4619) );
  NAND2X0 U5129 ( .IN1(n4622), .IN2(g296), .QN(n4621) );
  NAND2X0 U5130 ( .IN1(n373), .IN2(g1601), .QN(n4620) );
  AND2X1 U5131 ( .IN1(g1179), .IN2(n4595), .Q(n4618) );
  NOR2X0 U5132 ( .IN1(n4623), .IN2(n4624), .QN(n4616) );
  NOR2X0 U5133 ( .IN1(n1721), .IN2(n4625), .QN(n4624) );
  NOR2X0 U5134 ( .IN1(n2716), .IN2(n4626), .QN(n4623) );
  NAND2X0 U5135 ( .IN1(n4627), .IN2(n4628), .QN(n4614) );
  NOR2X0 U5136 ( .IN1(n4629), .IN2(n4630), .QN(n4628) );
  NAND2X0 U5137 ( .IN1(n4631), .IN2(n4632), .QN(n4630) );
  NAND2X0 U5138 ( .IN1(n4633), .IN2(g8), .QN(n4631) );
  NOR2X0 U5139 ( .IN1(n4938), .IN2(n4634), .QN(n4629) );
  NOR2X0 U5140 ( .IN1(n4635), .IN2(n4636), .QN(n4627) );
  NAND2X0 U5141 ( .IN1(n4637), .IN2(n4638), .QN(n4636) );
  NAND2X0 U5142 ( .IN1(g895), .IN2(n4639), .QN(n4638) );
  NAND2X0 U5143 ( .IN1(n4640), .IN2(g940), .QN(n4637) );
  NOR2X0 U5144 ( .IN1(n2557), .IN2(n4590), .QN(n4635) );
  NOR2X0 U5145 ( .IN1(n4641), .IN2(n4642), .QN(n4612) );
  NAND2X0 U5146 ( .IN1(n4643), .IN2(n4644), .QN(n4642) );
  NOR2X0 U5147 ( .IN1(n4645), .IN2(n4646), .QN(n4644) );
  NAND2X0 U5148 ( .IN1(n4647), .IN2(n4648), .QN(n4646) );
  NAND2X0 U5149 ( .IN1(n4649), .IN2(g959), .QN(n4648) );
  NAND2X0 U5150 ( .IN1(g1203), .IN2(n1512), .QN(n4647) );
  NOR2X0 U5151 ( .IN1(n2552), .IN2(n4650), .QN(n4645) );
  NOR2X0 U5152 ( .IN1(n4651), .IN2(n4652), .QN(n4643) );
  NOR2X0 U5153 ( .IN1(n1632), .IN2(n4653), .QN(n4652) );
  NOR2X0 U5154 ( .IN1(n2537), .IN2(n4654), .QN(n4651) );
  NAND2X0 U5155 ( .IN1(n4655), .IN2(n4656), .QN(n4641) );
  NOR2X0 U5156 ( .IN1(n4657), .IN2(n4658), .QN(n4656) );
  NAND2X0 U5157 ( .IN1(n4659), .IN2(n4660), .QN(n4658) );
  OR2X1 U5158 ( .IN1(n4589), .IN2(n1722), .Q(n4660) );
  NAND2X0 U5159 ( .IN1(g907), .IN2(n4586), .QN(n4659) );
  NOR2X0 U5160 ( .IN1(n2467), .IN2(n4661), .QN(n4657) );
  NOR2X0 U5161 ( .IN1(n4662), .IN2(n4663), .QN(n4655) );
  NOR2X0 U5162 ( .IN1(n4664), .IN2(DFF_228_n1), .QN(n4663) );
  NOR2X0 U5163 ( .IN1(n2472), .IN2(n4665), .QN(n4662) );
  NAND2X0 U5164 ( .IN1(n4382), .IN2(n3492), .QN(n4603) );
  AND2X1 U5165 ( .IN1(n4666), .IN2(n4934), .Q(n3492) );
  NOR2X0 U5166 ( .IN1(n2481), .IN2(n2759), .QN(n4666) );
  NOR2X0 U5167 ( .IN1(n4667), .IN2(n2760), .QN(n4382) );
  NAND2X0 U5168 ( .IN1(n2754), .IN2(n4070), .QN(g10465) );
  NOR2X0 U5169 ( .IN1(n4668), .IN2(n4669), .QN(n4070) );
  NAND2X0 U5170 ( .IN1(n4670), .IN2(n4671), .QN(n4669) );
  NOR2X0 U5171 ( .IN1(n4672), .IN2(n4673), .QN(n4671) );
  NAND2X0 U5172 ( .IN1(n4674), .IN2(n4675), .QN(n4673) );
  NAND2X0 U5173 ( .IN1(n4487), .IN2(n1650), .QN(n4675) );
  NAND2X0 U5174 ( .IN1(n4649), .IN2(g965), .QN(n4674) );
  NOR2X0 U5175 ( .IN1(n2546), .IN2(n4650), .QN(n4672) );
  NOR2X0 U5176 ( .IN1(n4676), .IN2(n4677), .QN(n4670) );
  NAND2X0 U5177 ( .IN1(n4678), .IN2(n4679), .QN(n4677) );
  NAND2X0 U5178 ( .IN1(n1485), .IN2(g1583), .QN(n4679) );
  NAND2X0 U5179 ( .IN1(n1486), .IN2(g1540), .QN(n4678) );
  NOR2X0 U5180 ( .IN1(n2717), .IN2(n4626), .QN(n4676) );
  NAND2X0 U5181 ( .IN1(n4680), .IN2(n4681), .QN(n4668) );
  NOR2X0 U5182 ( .IN1(n4682), .IN2(n4683), .QN(n4681) );
  NAND2X0 U5183 ( .IN1(n4684), .IN2(n4685), .QN(n4683) );
  NAND2X0 U5184 ( .IN1(g913), .IN2(n4586), .QN(n4684) );
  NAND2X0 U5185 ( .IN1(n4686), .IN2(n4687), .QN(n4682) );
  NAND2X0 U5186 ( .IN1(n4688), .IN2(g278), .QN(n4687) );
  NAND2X0 U5187 ( .IN1(n4622), .IN2(g302), .QN(n4686) );
  NOR2X0 U5188 ( .IN1(n4689), .IN2(n4690), .QN(n4680) );
  NAND2X0 U5189 ( .IN1(n4691), .IN2(n4692), .QN(n4690) );
  NAND2X0 U5190 ( .IN1(g1185), .IN2(n4595), .QN(n4692) );
  NAND2X0 U5191 ( .IN1(n4693), .IN2(g1330), .QN(n4691) );
  NOR2X0 U5192 ( .IN1(n2530), .IN2(n4694), .QN(n4689) );
  NAND2X0 U5193 ( .IN1(n2754), .IN2(n4414), .QN(g10463) );
  NOR2X0 U5194 ( .IN1(n4695), .IN2(n4696), .QN(n4414) );
  NAND2X0 U5195 ( .IN1(n4697), .IN2(n4698), .QN(n4696) );
  NOR2X0 U5196 ( .IN1(n4699), .IN2(n4700), .QN(n4698) );
  NAND2X0 U5197 ( .IN1(n4701), .IN2(n4702), .QN(n4700) );
  NAND2X0 U5198 ( .IN1(n4622), .IN2(g299), .QN(n4702) );
  NAND2X0 U5199 ( .IN1(n4703), .IN2(g1756), .QN(n4701) );
  NAND2X0 U5200 ( .IN1(n4704), .IN2(n4705), .QN(n4699) );
  NAND2X0 U5201 ( .IN1(n1485), .IN2(g1580), .QN(n4705) );
  NAND2X0 U5202 ( .IN1(n1486), .IN2(g1537), .QN(n4704) );
  NOR2X0 U5203 ( .IN1(n4706), .IN2(n4707), .QN(n4697) );
  NAND2X0 U5204 ( .IN1(n4708), .IN2(n4709), .QN(n4707) );
  NAND2X0 U5205 ( .IN1(n4487), .IN2(n3034), .QN(n4709) );
  NAND2X0 U5206 ( .IN1(n4649), .IN2(g962), .QN(n4708) );
  NAND2X0 U5207 ( .IN1(n4710), .IN2(n4711), .QN(n4706) );
  NAND2X0 U5208 ( .IN1(n4712), .IN2(n3057), .QN(n4711) );
  OR2X1 U5209 ( .IN1(n4713), .IN2(n4712), .Q(n4710) );
  NAND2X0 U5210 ( .IN1(n4714), .IN2(n4715), .QN(n4695) );
  NOR2X0 U5211 ( .IN1(n4716), .IN2(n4717), .QN(n4715) );
  NAND2X0 U5212 ( .IN1(n4718), .IN2(n4719), .QN(n4717) );
  NAND2X0 U5213 ( .IN1(n4688), .IN2(g275), .QN(n4719) );
  NAND2X0 U5214 ( .IN1(g1182), .IN2(n4595), .QN(n4718) );
  NAND2X0 U5215 ( .IN1(n4720), .IN2(n4721), .QN(n4716) );
  OR2X1 U5216 ( .IN1(n4661), .IN2(n2485), .Q(n4721) );
  NAND2X0 U5217 ( .IN1(n4693), .IN2(g1327), .QN(n4720) );
  NOR2X0 U5218 ( .IN1(n4722), .IN2(n4723), .QN(n4714) );
  NAND2X0 U5219 ( .IN1(n4724), .IN2(n4725), .QN(n4723) );
  NAND2X0 U5220 ( .IN1(n373), .IN2(g1604), .QN(n4725) );
  NAND2X0 U5221 ( .IN1(n1479), .IN2(g1561), .QN(n4724) );
  NAND2X0 U5222 ( .IN1(n4726), .IN2(n4727), .QN(n4722) );
  NAND2X0 U5223 ( .IN1(n4633), .IN2(n3025), .QN(n4727) );
  NAND2X0 U5224 ( .IN1(g910), .IN2(n4586), .QN(n4726) );
  NAND2X0 U5225 ( .IN1(n2754), .IN2(n4667), .QN(g10459) );
  INVX0 U5226 ( .INP(g10721), .ZN(n4667) );
  NAND2X0 U5227 ( .IN1(n4728), .IN2(n4729), .QN(g10721) );
  NOR2X0 U5228 ( .IN1(n4730), .IN2(n4731), .QN(n4729) );
  NAND2X0 U5229 ( .IN1(n4732), .IN2(n4733), .QN(n4731) );
  NOR2X0 U5230 ( .IN1(n4734), .IN2(n4735), .QN(n4733) );
  NAND2X0 U5231 ( .IN1(n4736), .IN2(n4737), .QN(n4735) );
  NAND2X0 U5232 ( .IN1(n4622), .IN2(g293), .QN(n4737) );
  NAND2X0 U5233 ( .IN1(n373), .IN2(g1598), .QN(n4736) );
  AND2X1 U5234 ( .IN1(g1176), .IN2(n4595), .Q(n4734) );
  NOR2X0 U5235 ( .IN1(n4738), .IN2(n4739), .QN(n4732) );
  NOR2X0 U5236 ( .IN1(n2706), .IN2(n4625), .QN(n4739) );
  NOR2X0 U5237 ( .IN1(n2712), .IN2(n4626), .QN(n4738) );
  NAND2X0 U5238 ( .IN1(n4740), .IN2(n4741), .QN(n4730) );
  NOR2X0 U5239 ( .IN1(n4742), .IN2(n4743), .QN(n4741) );
  NAND2X0 U5240 ( .IN1(n4744), .IN2(n4632), .QN(n4743) );
  NAND2X0 U5241 ( .IN1(n4633), .IN2(g1), .QN(n4744) );
  NOR2X0 U5242 ( .IN1(n2623), .IN2(n4634), .QN(n4742) );
  NOR2X0 U5243 ( .IN1(n4745), .IN2(n4746), .QN(n4740) );
  NAND2X0 U5244 ( .IN1(n4747), .IN2(n4748), .QN(n4746) );
  NAND2X0 U5245 ( .IN1(g892), .IN2(n4639), .QN(n4748) );
  NAND2X0 U5246 ( .IN1(n4640), .IN2(g936), .QN(n4747) );
  INVX0 U5247 ( .INP(n4749), .ZN(n4640) );
  NOR2X0 U5248 ( .IN1(n2563), .IN2(n4590), .QN(n4745) );
  NOR2X0 U5249 ( .IN1(n4750), .IN2(n4751), .QN(n4728) );
  NAND2X0 U5250 ( .IN1(n4752), .IN2(n4753), .QN(n4751) );
  NOR2X0 U5251 ( .IN1(n4754), .IN2(n4755), .QN(n4753) );
  NAND2X0 U5252 ( .IN1(n4756), .IN2(n4757), .QN(n4755) );
  NAND2X0 U5253 ( .IN1(n4649), .IN2(g956), .QN(n4757) );
  INVX0 U5254 ( .INP(n1472), .ZN(n4649) );
  NAND2X0 U5255 ( .IN1(g1200), .IN2(n1512), .QN(n4756) );
  NOR2X0 U5256 ( .IN1(n2528), .IN2(n4650), .QN(n4754) );
  NOR2X0 U5257 ( .IN1(n4758), .IN2(n4759), .QN(n4752) );
  NOR2X0 U5258 ( .IN1(n1652), .IN2(n4653), .QN(n4759) );
  NOR2X0 U5259 ( .IN1(n2551), .IN2(n4654), .QN(n4758) );
  NAND2X0 U5260 ( .IN1(n4760), .IN2(n4761), .QN(n4750) );
  NOR2X0 U5261 ( .IN1(n4762), .IN2(n4763), .QN(n4761) );
  NAND2X0 U5262 ( .IN1(n4764), .IN2(n4765), .QN(n4763) );
  NAND2X0 U5263 ( .IN1(n4766), .IN2(g981), .QN(n4765) );
  NAND2X0 U5264 ( .IN1(g904), .IN2(n4586), .QN(n4764) );
  NOR2X0 U5265 ( .IN1(n2486), .IN2(n4661), .QN(n4762) );
  NOR2X0 U5266 ( .IN1(n4767), .IN2(n4768), .QN(n4760) );
  NOR2X0 U5267 ( .IN1(n4664), .IN2(DFF_242_n1), .QN(n4768) );
  NOR2X0 U5268 ( .IN1(n2476), .IN2(n4665), .QN(n4767) );
  NAND2X0 U5269 ( .IN1(n2754), .IN2(n4500), .QN(g10457) );
  INVX0 U5270 ( .INP(g10720), .ZN(n4500) );
  NAND2X0 U5271 ( .IN1(n4769), .IN2(n4770), .QN(g10720) );
  NOR2X0 U5272 ( .IN1(n4771), .IN2(n4772), .QN(n4770) );
  NAND2X0 U5273 ( .IN1(n4773), .IN2(n4774), .QN(n4772) );
  NOR2X0 U5274 ( .IN1(n4775), .IN2(n4776), .QN(n4774) );
  NAND2X0 U5275 ( .IN1(n4777), .IN2(n4778), .QN(n4776) );
  NAND2X0 U5276 ( .IN1(n4622), .IN2(g290), .QN(n4778) );
  NAND2X0 U5277 ( .IN1(n373), .IN2(g1595), .QN(n4777) );
  INVX0 U5278 ( .INP(n4694), .ZN(n373) );
  AND2X1 U5279 ( .IN1(g1173), .IN2(n4595), .Q(n4775) );
  NOR2X0 U5280 ( .IN1(n4779), .IN2(n4780), .QN(n4773) );
  NOR2X0 U5281 ( .IN1(n2705), .IN2(n4625), .QN(n4780) );
  NOR2X0 U5282 ( .IN1(n2714), .IN2(n4626), .QN(n4779) );
  NAND2X0 U5283 ( .IN1(n4781), .IN2(n4782), .QN(n4771) );
  NOR2X0 U5284 ( .IN1(n4783), .IN2(n4784), .QN(n4782) );
  NAND2X0 U5285 ( .IN1(n4785), .IN2(n4632), .QN(n4784) );
  NAND2X0 U5286 ( .IN1(n4633), .IN2(g4), .QN(n4785) );
  NOR2X0 U5287 ( .IN1(n2622), .IN2(n4634), .QN(n4783) );
  NOR2X0 U5288 ( .IN1(n4786), .IN2(n4787), .QN(n4781) );
  NAND2X0 U5289 ( .IN1(n4788), .IN2(n4789), .QN(n4787) );
  NAND2X0 U5290 ( .IN1(g889), .IN2(n4639), .QN(n4789) );
  OR2X1 U5291 ( .IN1(n4749), .IN2(n1591), .Q(n4788) );
  NOR2X0 U5292 ( .IN1(n2554), .IN2(n4590), .QN(n4786) );
  NOR2X0 U5293 ( .IN1(n4790), .IN2(n4791), .QN(n4769) );
  NAND2X0 U5294 ( .IN1(n4792), .IN2(n4793), .QN(n4791) );
  NOR2X0 U5295 ( .IN1(n4794), .IN2(n4795), .QN(n4793) );
  NAND2X0 U5296 ( .IN1(n4796), .IN2(n4797), .QN(n4795) );
  NAND2X0 U5297 ( .IN1(n1512), .IN2(g1197), .QN(n4797) );
  NAND2X0 U5298 ( .IN1(n1530), .IN2(g925), .QN(n4796) );
  NOR2X0 U5299 ( .IN1(n2533), .IN2(n4650), .QN(n4794) );
  NOR2X0 U5300 ( .IN1(n4798), .IN2(n4799), .QN(n4792) );
  NOR2X0 U5301 ( .IN1(n1635), .IN2(n4653), .QN(n4799) );
  NOR2X0 U5302 ( .IN1(n2544), .IN2(n4654), .QN(n4798) );
  NAND2X0 U5303 ( .IN1(n4800), .IN2(n4801), .QN(n4790) );
  NOR2X0 U5304 ( .IN1(n4802), .IN2(n4803), .QN(n4801) );
  NAND2X0 U5305 ( .IN1(n4804), .IN2(n4805), .QN(n4803) );
  NAND2X0 U5306 ( .IN1(n4766), .IN2(g976), .QN(n4805) );
  INVX0 U5307 ( .INP(n4589), .ZN(n4766) );
  NAND2X0 U5308 ( .IN1(g901), .IN2(n4586), .QN(n4804) );
  NOR2X0 U5309 ( .IN1(n2484), .IN2(n4661), .QN(n4802) );
  NOR2X0 U5310 ( .IN1(n4806), .IN2(n4807), .QN(n4800) );
  NAND2X0 U5311 ( .IN1(n4808), .IN2(n4809), .QN(n4807) );
  NAND2X0 U5312 ( .IN1(n4693), .IN2(g1318), .QN(n4809) );
  NAND2X0 U5313 ( .IN1(n4487), .IN2(n3031), .QN(n4808) );
  NOR2X0 U5314 ( .IN1(n2468), .IN2(n1472), .QN(n4806) );
  NAND2X0 U5315 ( .IN1(n2754), .IN2(n4332), .QN(g10455) );
  INVX0 U5316 ( .INP(g10719), .ZN(n4332) );
  NAND2X0 U5317 ( .IN1(n4810), .IN2(n4811), .QN(g10719) );
  NOR2X0 U5318 ( .IN1(n4812), .IN2(n4813), .QN(n4811) );
  NAND2X0 U5319 ( .IN1(n4814), .IN2(n4815), .QN(n4813) );
  NOR2X0 U5320 ( .IN1(n4816), .IN2(n4817), .QN(n4815) );
  NAND2X0 U5321 ( .IN1(n4818), .IN2(n4819), .QN(n4817) );
  NAND2X0 U5322 ( .IN1(n4688), .IN2(g263), .QN(n4819) );
  INVX0 U5323 ( .INP(n4590), .ZN(n4688) );
  NAND2X0 U5324 ( .IN1(n4622), .IN2(g287), .QN(n4818) );
  INVX0 U5325 ( .INP(n4820), .ZN(n4622) );
  NOR2X0 U5326 ( .IN1(n2538), .IN2(n4694), .QN(n4816) );
  NOR2X0 U5327 ( .IN1(n4821), .IN2(n4822), .QN(n4814) );
  NAND2X0 U5328 ( .IN1(n4823), .IN2(n4824), .QN(n4822) );
  NAND2X0 U5329 ( .IN1(g1170), .IN2(n4595), .QN(n4824) );
  NAND2X0 U5330 ( .IN1(n4703), .IN2(g1744), .QN(n4823) );
  NOR2X0 U5331 ( .IN1(n2707), .IN2(n4625), .QN(n4821) );
  NAND2X0 U5332 ( .IN1(n4825), .IN2(n4826), .QN(n4812) );
  NOR2X0 U5333 ( .IN1(n4827), .IN2(n4828), .QN(n4826) );
  NAND2X0 U5334 ( .IN1(n4632), .IN2(n4829), .QN(n4828) );
  NAND2X0 U5335 ( .IN1(n4830), .IN2(n4831), .QN(n4632) );
  NOR2X0 U5336 ( .IN1(n1512), .IN2(n4598), .QN(n4831) );
  NOR2X0 U5337 ( .IN1(n4712), .IN2(n4713), .QN(n4830) );
  NAND2X0 U5338 ( .IN1(n4832), .IN2(n4833), .QN(n4713) );
  NOR2X0 U5339 ( .IN1(n369), .IN2(n4633), .QN(n4833) );
  INVX0 U5340 ( .INP(n4834), .ZN(n4633) );
  NOR2X0 U5341 ( .IN1(n4835), .IN2(n2948), .QN(n4832) );
  NAND2X0 U5342 ( .IN1(n4836), .IN2(n4837), .QN(n2948) );
  NOR2X0 U5343 ( .IN1(n4838), .IN2(n4839), .QN(n4837) );
  NAND2X0 U5344 ( .IN1(n1472), .IN2(n4820), .QN(n4839) );
  NAND2X0 U5345 ( .IN1(n4840), .IN2(n4841), .QN(n4820) );
  NOR2X0 U5346 ( .IN1(g43), .IN2(n4842), .QN(n4840) );
  NAND2X0 U5347 ( .IN1(n4843), .IN2(n4590), .QN(n4838) );
  NOR2X0 U5348 ( .IN1(n1530), .IN2(n4586), .QN(n4843) );
  NOR2X0 U5349 ( .IN1(n4844), .IN2(n4845), .QN(n4836) );
  NAND2X0 U5350 ( .IN1(n4664), .IN2(n4846), .QN(n4845) );
  NAND2X0 U5351 ( .IN1(n4749), .IN2(n4589), .QN(n4844) );
  NOR2X0 U5352 ( .IN1(n2488), .IN2(n4834), .QN(n4827) );
  NAND2X0 U5353 ( .IN1(n4847), .IN2(g42), .QN(n4834) );
  NOR2X0 U5354 ( .IN1(n4848), .IN2(n4849), .QN(n4825) );
  NAND2X0 U5355 ( .IN1(n4850), .IN2(n4851), .QN(n4849) );
  NAND2X0 U5356 ( .IN1(n4712), .IN2(g119), .QN(n4851) );
  INVX0 U5357 ( .INP(n4634), .ZN(n4712) );
  NAND2X0 U5358 ( .IN1(n4847), .IN2(n2961), .QN(n4634) );
  AND2X1 U5359 ( .IN1(n4852), .IN2(n4853), .Q(n4847) );
  NOR2X0 U5360 ( .IN1(g45), .IN2(g44), .QN(n4853) );
  NOR2X0 U5361 ( .IN1(n4842), .IN2(n4440), .QN(n4852) );
  INVX0 U5362 ( .INP(n1548), .ZN(n4842) );
  NAND2X0 U5363 ( .IN1(g886), .IN2(n4639), .QN(n4850) );
  INVX0 U5364 ( .INP(n4846), .ZN(n4639) );
  NAND2X0 U5365 ( .IN1(n4854), .IN2(n4855), .QN(n4846) );
  NOR2X0 U5366 ( .IN1(g44), .IN2(n4440), .QN(n4854) );
  NOR2X0 U5367 ( .IN1(n1604), .IN2(n4749), .QN(n4848) );
  NAND2X0 U5368 ( .IN1(n4856), .IN2(n4855), .QN(n4749) );
  AND2X1 U5369 ( .IN1(n4857), .IN2(n366), .Q(n4855) );
  NOR2X0 U5370 ( .IN1(g43), .IN2(n4858), .QN(n4856) );
  NOR2X0 U5371 ( .IN1(n4859), .IN2(n4860), .QN(n4810) );
  NAND2X0 U5372 ( .IN1(n4861), .IN2(n4862), .QN(n4860) );
  NOR2X0 U5373 ( .IN1(n4863), .IN2(n4864), .QN(n4862) );
  NAND2X0 U5374 ( .IN1(n4865), .IN2(n4866), .QN(n4864) );
  NAND2X0 U5375 ( .IN1(g1194), .IN2(n1512), .QN(n4866) );
  NAND2X0 U5376 ( .IN1(g922), .IN2(n1530), .QN(n4865) );
  NOR2X0 U5377 ( .IN1(n2535), .IN2(n4650), .QN(n4863) );
  NOR2X0 U5378 ( .IN1(n4867), .IN2(n4868), .QN(n4861) );
  NOR2X0 U5379 ( .IN1(n1649), .IN2(n4653), .QN(n4868) );
  NOR2X0 U5380 ( .IN1(n2526), .IN2(n4654), .QN(n4867) );
  INVX0 U5381 ( .INP(n1485), .ZN(n4654) );
  NAND2X0 U5382 ( .IN1(n4869), .IN2(n4870), .QN(n4859) );
  NOR2X0 U5383 ( .IN1(n4871), .IN2(n4872), .QN(n4870) );
  NAND2X0 U5384 ( .IN1(n4873), .IN2(n4874), .QN(n4872) );
  OR2X1 U5385 ( .IN1(n4589), .IN2(n2709), .Q(n4874) );
  NAND2X0 U5386 ( .IN1(g898), .IN2(n4586), .QN(n4873) );
  NOR2X0 U5387 ( .IN1(n2487), .IN2(n4661), .QN(n4871) );
  NOR2X0 U5388 ( .IN1(n4875), .IN2(n4876), .QN(n4869) );
  NAND2X0 U5389 ( .IN1(n4877), .IN2(n4878), .QN(n4876) );
  NAND2X0 U5390 ( .IN1(n4693), .IN2(g1314), .QN(n4878) );
  NAND2X0 U5391 ( .IN1(n4487), .IN2(n3051), .QN(n4877) );
  NOR2X0 U5392 ( .IN1(n2470), .IN2(n1472), .QN(n4875) );
  NAND2X0 U5393 ( .IN1(n366), .IN2(n4879), .QN(n1472) );
  NAND2X0 U5394 ( .IN1(n2754), .IN2(n4433), .QN(g10377) );
  INVX0 U5395 ( .INP(n38), .ZN(n4433) );
  NAND2X0 U5396 ( .IN1(n4880), .IN2(n4881), .QN(n38) );
  NOR2X0 U5397 ( .IN1(n4882), .IN2(n4883), .QN(n4881) );
  NAND2X0 U5398 ( .IN1(n4884), .IN2(n4885), .QN(n4883) );
  NAND2X0 U5399 ( .IN1(g1188), .IN2(n4595), .QN(n4885) );
  NOR2X0 U5400 ( .IN1(n4886), .IN2(n4887), .QN(n4884) );
  NOR2X0 U5401 ( .IN1(n2564), .IN2(n4590), .QN(n4887) );
  NAND2X0 U5402 ( .IN1(n4888), .IN2(n1548), .QN(n4590) );
  NOR2X0 U5403 ( .IN1(g43), .IN2(n4889), .QN(n4888) );
  NOR2X0 U5404 ( .IN1(n2469), .IN2(n4589), .QN(n4886) );
  NAND2X0 U5405 ( .IN1(n366), .IN2(n4890), .QN(n4589) );
  NAND2X0 U5406 ( .IN1(n4891), .IN2(n4892), .QN(n4882) );
  NOR2X0 U5407 ( .IN1(n1564), .IN2(n4893), .QN(n4892) );
  AND2X1 U5408 ( .IN1(g916), .IN2(n4586), .Q(n4893) );
  AND2X1 U5409 ( .IN1(n366), .IN2(n4894), .Q(n4586) );
  AND2X1 U5410 ( .IN1(n4895), .IN2(g46), .Q(n366) );
  NOR2X0 U5411 ( .IN1(g47), .IN2(n4896), .QN(n4895) );
  NOR2X0 U5412 ( .IN1(n4897), .IN2(n369), .QN(n4891) );
  INVX0 U5413 ( .INP(n4829), .ZN(n369) );
  NAND2X0 U5414 ( .IN1(n4898), .IN2(n4899), .QN(n4829) );
  NOR2X0 U5415 ( .IN1(n1545), .IN2(n4896), .QN(n4899) );
  NAND2X0 U5416 ( .IN1(g43), .IN2(n4841), .QN(n1545) );
  AND2X1 U5417 ( .IN1(n4900), .IN2(g44), .Q(n4841) );
  NOR2X0 U5418 ( .IN1(g45), .IN2(g42), .QN(n4900) );
  AND2X1 U5419 ( .IN1(g47), .IN2(g46), .Q(n4898) );
  NOR2X0 U5420 ( .IN1(n1640), .IN2(n4661), .QN(n4897) );
  NOR2X0 U5421 ( .IN1(n4901), .IN2(n4902), .QN(n4880) );
  NAND2X0 U5422 ( .IN1(n4903), .IN2(n4904), .QN(n4902) );
  NOR2X0 U5423 ( .IN1(n4905), .IN2(n4906), .QN(n4904) );
  NOR2X0 U5424 ( .IN1(n4598), .IN2(n4685), .QN(n4906) );
  NAND2X0 U5425 ( .IN1(n1478), .IN2(n4907), .QN(n4685) );
  INVX0 U5426 ( .INP(n4835), .ZN(n4907) );
  NAND2X0 U5427 ( .IN1(n4908), .IN2(n4600), .QN(n4835) );
  AND2X1 U5428 ( .IN1(n4909), .IN2(n4910), .Q(n4600) );
  NOR2X0 U5429 ( .IN1(n1567), .IN2(n1566), .QN(n4910) );
  NAND2X0 U5430 ( .IN1(n4650), .IN2(n4911), .QN(n1566) );
  NAND2X0 U5431 ( .IN1(n4894), .IN2(n1548), .QN(n4911) );
  INVX0 U5432 ( .INP(n1479), .ZN(n4650) );
  NAND2X0 U5433 ( .IN1(n4694), .IN2(n4912), .QN(n1567) );
  NAND2X0 U5434 ( .IN1(n4890), .IN2(n1548), .QN(n4912) );
  NAND2X0 U5435 ( .IN1(n4879), .IN2(n1548), .QN(n4694) );
  NOR2X0 U5436 ( .IN1(n4913), .IN2(n4896), .QN(n1548) );
  OR2X1 U5437 ( .IN1(g47), .IN2(g46), .Q(n4913) );
  NOR2X0 U5438 ( .IN1(n4583), .IN2(n4595), .QN(n4909) );
  AND2X1 U5439 ( .IN1(n4894), .IN2(n362), .Q(n4595) );
  NOR2X0 U5440 ( .IN1(n4440), .IN2(n4889), .QN(n4894) );
  NAND2X0 U5441 ( .IN1(n4914), .IN2(g44), .QN(n4889) );
  NOR2X0 U5442 ( .IN1(g45), .IN2(n2961), .QN(n4914) );
  INVX0 U5443 ( .INP(g43), .ZN(n4440) );
  INVX0 U5444 ( .INP(n4661), .ZN(n4583) );
  NAND2X0 U5445 ( .IN1(n4915), .IN2(g42), .QN(n4661) );
  NOR2X0 U5446 ( .IN1(n4693), .IN2(n4703), .QN(n4908) );
  INVX0 U5447 ( .INP(n4626), .ZN(n4703) );
  INVX0 U5448 ( .INP(n4665), .ZN(n4693) );
  INVX0 U5449 ( .INP(n4625), .ZN(n4598) );
  NOR2X0 U5450 ( .IN1(n2479), .IN2(n4625), .QN(n4905) );
  NAND2X0 U5451 ( .IN1(n4890), .IN2(n362), .QN(n4625) );
  AND2X1 U5452 ( .IN1(n4857), .IN2(n4916), .Q(n4890) );
  NOR2X0 U5453 ( .IN1(n2961), .IN2(n4438), .QN(n4857) );
  NOR2X0 U5454 ( .IN1(n4917), .IN2(n4918), .QN(n4903) );
  NOR2X0 U5455 ( .IN1(n2478), .IN2(n4665), .QN(n4918) );
  NAND2X0 U5456 ( .IN1(n4879), .IN2(n362), .QN(n4665) );
  AND2X1 U5457 ( .IN1(n4919), .IN2(n4916), .Q(n4879) );
  NOR2X0 U5458 ( .IN1(g44), .IN2(g43), .QN(n4916) );
  NOR2X0 U5459 ( .IN1(g42), .IN2(n4438), .QN(n4919) );
  NOR2X0 U5460 ( .IN1(n2548), .IN2(n4653), .QN(n4917) );
  INVX0 U5461 ( .INP(n1486), .ZN(n4653) );
  NAND2X0 U5462 ( .IN1(n4920), .IN2(n4921), .QN(n4901) );
  NAND2X0 U5463 ( .IN1(n1485), .IN2(g1586), .QN(n4921) );
  NOR2X0 U5464 ( .IN1(n4922), .IN2(n4923), .QN(n4920) );
  NOR2X0 U5465 ( .IN1(n4939), .IN2(n4664), .QN(n4923) );
  NOR2X0 U5466 ( .IN1(n2715), .IN2(n4626), .QN(n4922) );
  NAND2X0 U5467 ( .IN1(n4915), .IN2(n2961), .QN(n4626) );
  INVX0 U5468 ( .INP(g42), .ZN(n2961) );
  AND2X1 U5469 ( .IN1(n4924), .IN2(n4925), .Q(n4915) );
  NOR2X0 U5470 ( .IN1(n4858), .IN2(n4438), .QN(n4925) );
  INVX0 U5471 ( .INP(g45), .ZN(n4438) );
  INVX0 U5472 ( .INP(g44), .ZN(n4858) );
  AND2X1 U5473 ( .IN1(n362), .IN2(g43), .Q(n4924) );
  NOR2X0 U5474 ( .IN1(n2962), .IN2(n4896), .QN(n362) );
  NAND2X0 U5475 ( .IN1(n2984), .IN2(g48), .QN(n4896) );
  NOR2X0 U5476 ( .IN1(g41), .IN2(n4926), .QN(n2984) );
  NAND2X0 U5477 ( .IN1(n4927), .IN2(n4928), .QN(n4926) );
  NAND2X0 U5478 ( .IN1(g30), .IN2(n4439), .QN(n4928) );
  NAND2X0 U5479 ( .IN1(g48), .IN2(n4487), .QN(n4927) );
  NAND2X0 U5480 ( .IN1(g47), .IN2(n2956), .QN(n2962) );
  INVX0 U5481 ( .INP(g46), .ZN(n2956) );
  NOR2X0 U5482 ( .IN1(n4487), .IN2(g30), .QN(n2754) );
  INVX0 U5483 ( .INP(n4664), .ZN(n4487) );
  NOR2X0 U5484 ( .IN1(n4439), .IN2(g31), .QN(n4664) );
  INVX0 U5485 ( .INP(g48), .ZN(n4439) );
  XNOR2X1 U5486 ( .IN1(test_so1), .IN2(n3470), .Q(N599) );
  NAND2X0 U5487 ( .IN1(n4929), .IN2(n1093), .QN(n3470) );
  NOR2X0 U5488 ( .IN1(n2524), .IN2(n2519), .QN(n4929) );
  OR2X1 U1550_U1 ( .IN1(g10722), .IN2(n2754), .Q(g10461) );
  OR2X1 U1551_U1 ( .IN1(g10664), .IN2(n2754), .Q(g10379) );
  INVX0 U1586_U2 ( .INP(n11), .ZN(U1586_n1) );
  NOR2X0 U1586_U1 ( .IN1(n2749), .IN2(U1586_n1), .QN(n1855) );
  INVX0 U1754_U2 ( .INP(n1548), .ZN(U1754_n1) );
  NOR2X0 U1754_U1 ( .IN1(n1545), .IN2(U1754_n1), .QN(n1479) );
  INVX0 U1798_U2 ( .INP(n1567), .ZN(U1798_n1) );
  NOR2X0 U1798_U1 ( .IN1(n373), .IN2(U1798_n1), .QN(n1485) );
  INVX0 U1839_U2 ( .INP(n1566), .ZN(U1839_n1) );
  NOR2X0 U1839_U1 ( .IN1(n1479), .IN2(U1839_n1), .QN(n1486) );
  INVX0 U1843_U2 ( .INP(n343), .ZN(U1843_n1) );
  NOR2X0 U1843_U1 ( .IN1(n369), .IN2(U1843_n1), .QN(n1478) );
  INVX0 U1877_U2 ( .INP(n1137), .ZN(U1877_n1) );
  NOR2X0 U1877_U1 ( .IN1(n2757), .IN2(U1877_n1), .QN(n1195) );
  INVX0 U1908_U2 ( .INP(n362), .ZN(U1908_n1) );
  NOR2X0 U1908_U1 ( .IN1(n1545), .IN2(U1908_n1), .QN(n1512) );
  INVX0 U1909_U2 ( .INP(n366), .ZN(U1909_n1) );
  NOR2X0 U1909_U1 ( .IN1(n1545), .IN2(U1909_n1), .QN(n1530) );
  INVX0 U1987_U2 ( .INP(n822), .ZN(U1987_n1) );
  NOR2X0 U1987_U1 ( .IN1(n168), .IN2(U1987_n1), .QN(n916) );
  INVX0 U2031_U2 ( .INP(n1057), .ZN(U2031_n1) );
  NOR2X0 U2031_U1 ( .IN1(n1054), .IN2(U2031_n1), .QN(n1056) );
  INVX0 U2035_U2 ( .INP(n1404), .ZN(U2035_n1) );
  NOR2X0 U2035_U1 ( .IN1(g109), .IN2(U2035_n1), .QN(n1450) );
  INVX0 U2418_U2 ( .INP(g968), .ZN(U2418_n1) );
  NOR2X0 U2418_U1 ( .IN1(n1472), .IN2(U2418_n1), .QN(n1564) );
  INVX0 U2468_U2 ( .INP(g1336), .ZN(U2468_n1) );
  NOR2X0 U2468_U1 ( .IN1(n1227), .IN2(U2468_n1), .QN(n1231) );
  INVX0 U2478_U2 ( .INP(g1341), .ZN(U2478_n1) );
  NOR2X0 U2478_U1 ( .IN1(n1229), .IN2(U2478_n1), .QN(n1232) );
  INVX0 U2488_U2 ( .INP(n1262), .ZN(U2488_n1) );
  NOR2X0 U2488_U1 ( .IN1(n20), .IN2(U2488_n1), .QN(n1260) );
  INVX0 U2533_U2 ( .INP(g178), .ZN(U2533_n1) );
  NOR2X0 U2533_U1 ( .IN1(n2758), .IN2(U2533_n1), .QN(g6786) );
  INVX0 U2534_U2 ( .INP(g1424), .ZN(U2534_n1) );
  NOR2X0 U2534_U1 ( .IN1(n2759), .IN2(U2534_n1), .QN(g6234) );
  INVX0 U2639_U2 ( .INP(n962), .ZN(U2639_n1) );
  NOR2X0 U2639_U1 ( .IN1(n958), .IN2(U2639_n1), .QN(n804) );
  INVX0 U2641_U2 ( .INP(n34), .ZN(U2641_n1) );
  NOR2X0 U2641_U1 ( .IN1(g1868), .IN2(U2641_n1), .QN(n926) );
  INVX0 U2654_U2 ( .INP(g746), .ZN(U2654_n1) );
  NOR2X0 U2654_U1 ( .IN1(g750), .IN2(U2654_n1), .QN(g4171) );
  INVX0 U2658_U2 ( .INP(n917), .ZN(U2658_n1) );
  NOR2X0 U2658_U1 ( .IN1(n918), .IN2(U2658_n1), .QN(n812) );
  INVX0 U2683_U2 ( .INP(g382), .ZN(U2683_n1) );
  NOR2X0 U2683_U1 ( .IN1(n1385), .IN2(U2683_n1), .QN(n1420) );
  INVX0 U2699_U2 ( .INP(n808), .ZN(U2699_n1) );
  NOR2X0 U2699_U1 ( .IN1(n346), .IN2(U2699_n1), .QN(n806) );
  INVX0 U2846_U2 ( .INP(g4175), .ZN(U2846_n1) );
  NOR2X0 U2846_U1 ( .IN1(n1214), .IN2(U2846_n1), .QN(n1193) );
  INVX0 U2847_U2 ( .INP(g4177), .ZN(U2847_n1) );
  NOR2X0 U2847_U1 ( .IN1(n1153), .IN2(U2847_n1), .QN(n1125) );
  INVX0 U2848_U2 ( .INP(g4179), .ZN(U2848_n1) );
  NOR2X0 U2848_U1 ( .IN1(n1099), .IN2(U2848_n1), .QN(n1093) );
  INVX0 U2859_U2 ( .INP(n1137), .ZN(U2859_n1) );
  NOR2X0 U2859_U1 ( .IN1(g12), .IN2(U2859_n1), .QN(n1159) );
  INVX0 U2860_U2 ( .INP(g810), .ZN(U2860_n1) );
  NOR2X0 U2860_U1 ( .IN1(n1151), .IN2(U2860_n1), .QN(n1123) );
  INVX0 U2861_U2 ( .INP(g818), .ZN(U2861_n1) );
  NOR2X0 U2861_U1 ( .IN1(n1097), .IN2(U2861_n1), .QN(n1090) );
  INVX0 U2867_U2 ( .INP(n817), .ZN(U2867_n1) );
  NOR2X0 U2867_U1 ( .IN1(g1834), .IN2(U2867_n1), .QN(n1380) );
  INVX0 U2879_U2 ( .INP(g713), .ZN(U2879_n1) );
  NOR2X0 U2879_U1 ( .IN1(n1656), .IN2(U2879_n1), .QN(n967) );
  INVX0 U2881_U2 ( .INP(g1927), .ZN(U2881_n1) );
  NOR2X0 U2881_U1 ( .IN1(n1657), .IN2(U2881_n1), .QN(n921) );
  INVX0 U2882_U2 ( .INP(g1160), .ZN(U2882_n1) );
  NOR2X0 U2882_U1 ( .IN1(n2760), .IN2(U2882_n1), .QN(g4334) );
  INVX0 U2883_U2 ( .INP(g1166), .ZN(U2883_n1) );
  NOR2X0 U2883_U1 ( .IN1(n2757), .IN2(U2883_n1), .QN(g4325) );
  INVX0 U2884_U2 ( .INP(g148), .ZN(U2884_n1) );
  NOR2X0 U2884_U1 ( .IN1(n2758), .IN2(U2884_n1), .QN(g6759) );
  INVX0 U2885_U2 ( .INP(g1157), .ZN(U2885_n1) );
  NOR2X0 U2885_U1 ( .IN1(n2759), .IN2(U2885_n1), .QN(g4338) );
  INVX0 U2886_U2 ( .INP(g1163), .ZN(U2886_n1) );
  NOR2X0 U2886_U1 ( .IN1(n2760), .IN2(U2886_n1), .QN(g4330) );
  INVX0 U2887_U2 ( .INP(g237), .ZN(U2887_n1) );
  NOR2X0 U2887_U1 ( .IN1(n2757), .IN2(U2887_n1), .QN(g6821) );
  INVX0 U2888_U2 ( .INP(g1499), .ZN(U2888_n1) );
  NOR2X0 U2888_U1 ( .IN1(n2758), .IN2(U2888_n1), .QN(g6198) );
  INVX0 U2889_U2 ( .INP(g1411), .ZN(U2889_n1) );
  NOR2X0 U2889_U1 ( .IN1(n2759), .IN2(U2889_n1), .QN(g6244) );
  INVX0 U2890_U2 ( .INP(g225), .ZN(U2890_n1) );
  NOR2X0 U2890_U1 ( .IN1(n2760), .IN2(U2890_n1), .QN(g6826) );
  INVX0 U2891_U2 ( .INP(g1407), .ZN(U2891_n1) );
  NOR2X0 U2891_U1 ( .IN1(n2757), .IN2(U2891_n1), .QN(g6216) );
  INVX0 U2892_U2 ( .INP(g213), .ZN(U2892_n1) );
  NOR2X0 U2892_U1 ( .IN1(n2758), .IN2(U2892_n1), .QN(g6829) );
  INVX0 U2893_U2 ( .INP(g186), .ZN(U2893_n1) );
  NOR2X0 U2893_U1 ( .IN1(n2759), .IN2(U2893_n1), .QN(g6833) );
  INVX0 U2894_U2 ( .INP(g219), .ZN(U2894_n1) );
  NOR2X0 U2894_U1 ( .IN1(n2760), .IN2(U2894_n1), .QN(g6827) );
  INVX0 U2895_U2 ( .INP(g143), .ZN(U2895_n1) );
  NOR2X0 U2895_U1 ( .IN1(n2757), .IN2(U2895_n1), .QN(g6757) );
  INVX0 U2896_U2 ( .INP(g207), .ZN(U2896_n1) );
  NOR2X0 U2896_U1 ( .IN1(n2758), .IN2(U2896_n1), .QN(g6831) );
  INVX0 U2897_U2 ( .INP(g231), .ZN(U2897_n1) );
  NOR2X0 U2897_U1 ( .IN1(n2759), .IN2(U2897_n1), .QN(g6822) );
  INVX0 U2898_U2 ( .INP(g192), .ZN(U2898_n1) );
  NOR2X0 U2898_U1 ( .IN1(n2760), .IN2(U2898_n1), .QN(g6838) );
  INVX0 U2899_U2 ( .INP(test_so3), .ZN(U2899_n1) );
  NOR2X0 U2899_U1 ( .IN1(n2757), .IN2(U2899_n1), .QN(g6823) );
  INVX0 U2900_U2 ( .INP(g1371), .ZN(U2900_n1) );
  NOR2X0 U2900_U1 ( .IN1(n2758), .IN2(U2900_n1), .QN(g6824) );
  INVX0 U2901_U2 ( .INP(g1383), .ZN(U2901_n1) );
  NOR2X0 U2901_U1 ( .IN1(n2759), .IN2(U2901_n1), .QN(g6832) );
  INVX0 U2902_U2 ( .INP(g243), .ZN(U2902_n1) );
  NOR2X0 U2902_U1 ( .IN1(n2760), .IN2(U2902_n1), .QN(g6819) );
  INVX0 U3090_U2 ( .INP(n1151), .ZN(U3090_n1) );
  NOR2X0 U3090_U1 ( .IN1(g810), .IN2(U3090_n1), .QN(n1150) );
  INVX0 U3092_U2 ( .INP(n1097), .ZN(U3092_n1) );
  NOR2X0 U3092_U1 ( .IN1(g818), .IN2(U3092_n1), .QN(n1096) );
  INVX0 U3094_U2 ( .INP(n1099), .ZN(U3094_n1) );
  NOR2X0 U3094_U1 ( .IN1(g4179), .IN2(U3094_n1), .QN(n1098) );
  INVX0 U3096_U2 ( .INP(n1214), .ZN(U3096_n1) );
  NOR2X0 U3096_U1 ( .IN1(g4175), .IN2(U3096_n1), .QN(n1213) );
  INVX0 U3098_U2 ( .INP(n1153), .ZN(U3098_n1) );
  NOR2X0 U3098_U1 ( .IN1(g4177), .IN2(U3098_n1), .QN(n1152) );
  INVX0 U3124_U2 ( .INP(n837), .ZN(U3124_n1) );
  NOR2X0 U3124_U1 ( .IN1(n838), .IN2(U3124_n1), .QN(n836) );
  INVX0 U3171_U2 ( .INP(g1610), .ZN(U3171_n1) );
  NOR2X0 U3171_U1 ( .IN1(n256), .IN2(U3171_n1), .QN(g5194) );
endmodule

