module add_mul_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, 
        a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, 
        a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, 
        b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, 
        b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, 
        b_28_, b_29_, b_30_, b_31_, operation, Result_0_, Result_1_, Result_2_, 
        Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, 
        Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, 
        Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, 
        Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, 
        Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, Result_32_, 
        Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, Result_38_, 
        Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, Result_44_, 
        Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, Result_50_, 
        Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, Result_56_, 
        Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, Result_62_, 
        Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803;

  INV_X4 U8483 ( .A(operation), .ZN(n8421) );
  INV_X2 U8484 ( .A(b_26_), .ZN(n10156) );
  INV_X2 U8485 ( .A(b_21_), .ZN(n8599) );
  INV_X2 U8486 ( .A(b_23_), .ZN(n8570) );
  INV_X2 U8487 ( .A(b_15_), .ZN(n8690) );
  INV_X2 U8488 ( .A(b_19_), .ZN(n8628) );
  INV_X2 U8489 ( .A(b_22_), .ZN(n8983) );
  INV_X2 U8490 ( .A(b_25_), .ZN(n8543) );
  INV_X2 U8491 ( .A(b_2_), .ZN(n8997) );
  INV_X2 U8492 ( .A(b_14_), .ZN(n8990) );
  INV_X2 U8493 ( .A(b_11_), .ZN(n8751) );
  INV_X2 U8494 ( .A(a_17_), .ZN(n8662) );
  INV_X2 U8495 ( .A(a_12_), .ZN(n8739) );
  INV_X2 U8496 ( .A(a_20_), .ZN(n8986) );
  INV_X2 U8497 ( .A(a_26_), .ZN(n9893) );
  INV_X2 U8498 ( .A(a_10_), .ZN(n8769) );
  INV_X2 U8499 ( .A(a_2_), .ZN(n8998) );
  NAND2_X2 U8500 ( .A1(a_31_), .A2(a_30_), .ZN(n8979) );
  INV_X2 U8501 ( .A(a_3_), .ZN(n8877) );
  INV_X2 U8502 ( .A(a_18_), .ZN(n8988) );
  INV_X2 U8503 ( .A(a_25_), .ZN(n8541) );
  INV_X2 U8504 ( .A(a_7_), .ZN(n8817) );
  NAND2_X2 U8505 ( .A1(a_31_), .A2(n16582), .ZN(n8456) );
  NAND2_X2 U8506 ( .A1(a_30_), .A2(n8978), .ZN(n8459) );
  INV_X2 U8507 ( .A(a_13_), .ZN(n8721) );
  INV_X2 U8508 ( .A(a_27_), .ZN(n8512) );
  INV_X2 U8509 ( .A(a_24_), .ZN(n8982) );
  INV_X2 U8510 ( .A(b_9_), .ZN(n8781) );
  INV_X2 U8511 ( .A(a_9_), .ZN(n8779) );
  INV_X2 U8512 ( .A(a_28_), .ZN(n8493) );
  INV_X2 U8513 ( .A(b_17_), .ZN(n8660) );
  INV_X2 U8514 ( .A(b_8_), .ZN(n14458) );
  INV_X2 U8515 ( .A(b_10_), .ZN(n8992) );
  INV_X2 U8516 ( .A(b_7_), .ZN(n8819) );
  INV_X2 U8517 ( .A(a_29_), .ZN(n8473) );
  INV_X2 U8518 ( .A(b_1_), .ZN(n8907) );
  INV_X2 U8519 ( .A(b_13_), .ZN(n8719) );
  INV_X2 U8520 ( .A(b_4_), .ZN(n8995) );
  INV_X2 U8521 ( .A(b_3_), .ZN(n8875) );
  INV_X2 U8522 ( .A(a_11_), .ZN(n8749) );
  INV_X2 U8523 ( .A(a_5_), .ZN(n8848) );
  INV_X2 U8524 ( .A(a_21_), .ZN(n8601) );
  INV_X2 U8525 ( .A(b_6_), .ZN(n8993) );
  INV_X2 U8526 ( .A(a_15_), .ZN(n8692) );
  INV_X2 U8527 ( .A(b_5_), .ZN(n8846) );
  NOR2_X1 U8528 ( .A1(n8420), .A2(n8421), .ZN(Result_9_) );
  XOR2_X1 U8529 ( .A(n8422), .B(n8423), .Z(n8420) );
  NAND2_X1 U8530 ( .A1(n8424), .A2(n8425), .ZN(n8422) );
  NAND2_X1 U8531 ( .A1(n8426), .A2(n8427), .ZN(n8425) );
  NAND2_X1 U8532 ( .A1(n8428), .A2(n8429), .ZN(n8426) );
  NOR2_X1 U8533 ( .A1(n8430), .A2(n8421), .ZN(Result_8_) );
  XNOR2_X1 U8534 ( .A(n8431), .B(n8432), .ZN(n8430) );
  NOR2_X1 U8535 ( .A1(n8433), .A2(n8421), .ZN(Result_7_) );
  XNOR2_X1 U8536 ( .A(n8434), .B(n8435), .ZN(n8433) );
  NAND2_X1 U8537 ( .A1(n8436), .A2(n8437), .ZN(n8434) );
  NAND2_X1 U8538 ( .A1(n8438), .A2(n8439), .ZN(n8437) );
  NAND2_X1 U8539 ( .A1(n8440), .A2(n8441), .ZN(n8438) );
  NOR2_X1 U8540 ( .A1(n8442), .A2(n8421), .ZN(Result_6_) );
  XNOR2_X1 U8541 ( .A(n8443), .B(n8444), .ZN(n8442) );
  NAND2_X1 U8542 ( .A1(n8445), .A2(n8446), .ZN(Result_63_) );
  NAND2_X1 U8543 ( .A1(n8447), .A2(n8421), .ZN(n8446) );
  XNOR2_X1 U8544 ( .A(n8448), .B(a_31_), .ZN(n8447) );
  NAND2_X1 U8545 ( .A1(n8449), .A2(operation), .ZN(n8445) );
  NAND2_X1 U8546 ( .A1(n8450), .A2(n8451), .ZN(Result_62_) );
  NAND2_X1 U8547 ( .A1(operation), .A2(n8452), .ZN(n8451) );
  NAND2_X1 U8548 ( .A1(n8453), .A2(n8454), .ZN(n8452) );
  NAND2_X1 U8549 ( .A1(b_30_), .A2(n8455), .ZN(n8454) );
  NAND2_X1 U8550 ( .A1(n8456), .A2(n8457), .ZN(n8455) );
  NAND2_X1 U8551 ( .A1(a_31_), .A2(n8448), .ZN(n8457) );
  NAND2_X1 U8552 ( .A1(b_31_), .A2(n8458), .ZN(n8453) );
  NAND2_X1 U8553 ( .A1(n8459), .A2(n8460), .ZN(n8458) );
  NAND2_X1 U8554 ( .A1(a_30_), .A2(n8461), .ZN(n8460) );
  NAND2_X1 U8555 ( .A1(n8462), .A2(n8421), .ZN(n8450) );
  XNOR2_X1 U8556 ( .A(n8449), .B(n8463), .ZN(n8462) );
  XNOR2_X1 U8557 ( .A(a_30_), .B(b_30_), .ZN(n8463) );
  NAND2_X1 U8558 ( .A1(n8464), .A2(n8465), .ZN(Result_61_) );
  NAND2_X1 U8559 ( .A1(n8466), .A2(n8421), .ZN(n8465) );
  NAND3_X1 U8560 ( .A1(n8467), .A2(n8468), .A3(n8469), .ZN(n8466) );
  NAND2_X1 U8561 ( .A1(n8470), .A2(n8471), .ZN(n8469) );
  NAND3_X1 U8562 ( .A1(n8472), .A2(n8473), .A3(b_29_), .ZN(n8468) );
  NAND2_X1 U8563 ( .A1(n8474), .A2(n8475), .ZN(n8467) );
  XNOR2_X1 U8564 ( .A(a_29_), .B(n8472), .ZN(n8474) );
  NAND2_X1 U8565 ( .A1(n8476), .A2(operation), .ZN(n8464) );
  XNOR2_X1 U8566 ( .A(n8477), .B(n8478), .ZN(n8476) );
  XOR2_X1 U8567 ( .A(n8479), .B(n8480), .Z(n8478) );
  NAND2_X1 U8568 ( .A1(n8481), .A2(n8482), .ZN(Result_60_) );
  NAND2_X1 U8569 ( .A1(n8483), .A2(n8421), .ZN(n8482) );
  XNOR2_X1 U8570 ( .A(n8484), .B(n8485), .ZN(n8483) );
  NAND2_X1 U8571 ( .A1(n8486), .A2(n8487), .ZN(n8484) );
  NAND2_X1 U8572 ( .A1(n8488), .A2(operation), .ZN(n8481) );
  XOR2_X1 U8573 ( .A(n8489), .B(n8490), .Z(n8488) );
  XOR2_X1 U8574 ( .A(n8491), .B(n8492), .Z(n8489) );
  NOR2_X1 U8575 ( .A1(n8493), .A2(n8448), .ZN(n8492) );
  NOR2_X1 U8576 ( .A1(n8494), .A2(n8421), .ZN(Result_5_) );
  XNOR2_X1 U8577 ( .A(n8495), .B(n8496), .ZN(n8494) );
  NAND2_X1 U8578 ( .A1(n8497), .A2(n8498), .ZN(n8495) );
  NAND2_X1 U8579 ( .A1(n8499), .A2(n8500), .ZN(n8498) );
  NAND2_X1 U8580 ( .A1(n8501), .A2(n8502), .ZN(n8499) );
  NAND2_X1 U8581 ( .A1(n8503), .A2(n8504), .ZN(Result_59_) );
  NAND2_X1 U8582 ( .A1(n8505), .A2(n8421), .ZN(n8504) );
  NAND3_X1 U8583 ( .A1(n8506), .A2(n8507), .A3(n8508), .ZN(n8505) );
  NAND2_X1 U8584 ( .A1(n8509), .A2(n8510), .ZN(n8508) );
  NAND3_X1 U8585 ( .A1(n8511), .A2(n8512), .A3(b_27_), .ZN(n8507) );
  NAND2_X1 U8586 ( .A1(n8513), .A2(n8514), .ZN(n8506) );
  XNOR2_X1 U8587 ( .A(a_27_), .B(n8511), .ZN(n8513) );
  NAND2_X1 U8588 ( .A1(n8515), .A2(operation), .ZN(n8503) );
  XOR2_X1 U8589 ( .A(n8516), .B(n8517), .Z(n8515) );
  XOR2_X1 U8590 ( .A(n8518), .B(n8519), .Z(n8517) );
  NAND2_X1 U8591 ( .A1(n8520), .A2(n8521), .ZN(Result_58_) );
  NAND2_X1 U8592 ( .A1(n8522), .A2(n8421), .ZN(n8521) );
  XNOR2_X1 U8593 ( .A(n8523), .B(n8524), .ZN(n8522) );
  NOR2_X1 U8594 ( .A1(n8525), .A2(n8526), .ZN(n8524) );
  NAND2_X1 U8595 ( .A1(n8527), .A2(operation), .ZN(n8520) );
  XNOR2_X1 U8596 ( .A(n8528), .B(n8529), .ZN(n8527) );
  XOR2_X1 U8597 ( .A(n8530), .B(n8531), .Z(n8529) );
  NAND2_X1 U8598 ( .A1(n8532), .A2(n8533), .ZN(Result_57_) );
  NAND2_X1 U8599 ( .A1(n8534), .A2(n8421), .ZN(n8533) );
  NAND3_X1 U8600 ( .A1(n8535), .A2(n8536), .A3(n8537), .ZN(n8534) );
  NAND2_X1 U8601 ( .A1(n8538), .A2(n8539), .ZN(n8537) );
  NAND3_X1 U8602 ( .A1(n8540), .A2(n8541), .A3(b_25_), .ZN(n8536) );
  NAND2_X1 U8603 ( .A1(n8542), .A2(n8543), .ZN(n8535) );
  XNOR2_X1 U8604 ( .A(n8540), .B(a_25_), .ZN(n8542) );
  NAND2_X1 U8605 ( .A1(n8544), .A2(operation), .ZN(n8532) );
  XNOR2_X1 U8606 ( .A(n8545), .B(n8546), .ZN(n8544) );
  XNOR2_X1 U8607 ( .A(n8547), .B(n8548), .ZN(n8545) );
  NAND2_X1 U8608 ( .A1(n8549), .A2(n8550), .ZN(Result_56_) );
  NAND2_X1 U8609 ( .A1(n8551), .A2(n8421), .ZN(n8550) );
  XNOR2_X1 U8610 ( .A(n8552), .B(n8553), .ZN(n8551) );
  NAND2_X1 U8611 ( .A1(n8554), .A2(n8555), .ZN(n8553) );
  NAND2_X1 U8612 ( .A1(n8556), .A2(operation), .ZN(n8549) );
  XNOR2_X1 U8613 ( .A(n8557), .B(n8558), .ZN(n8556) );
  XNOR2_X1 U8614 ( .A(n8559), .B(n8560), .ZN(n8558) );
  NAND2_X1 U8615 ( .A1(n8561), .A2(n8562), .ZN(Result_55_) );
  NAND2_X1 U8616 ( .A1(n8563), .A2(n8421), .ZN(n8562) );
  NAND3_X1 U8617 ( .A1(n8564), .A2(n8565), .A3(n8566), .ZN(n8563) );
  NAND2_X1 U8618 ( .A1(n8567), .A2(n8568), .ZN(n8566) );
  INV_X1 U8619 ( .A(n8569), .ZN(n8565) );
  NOR3_X1 U8620 ( .A1(n8568), .A2(a_23_), .A3(n8570), .ZN(n8569) );
  NAND2_X1 U8621 ( .A1(n8571), .A2(n8570), .ZN(n8564) );
  XNOR2_X1 U8622 ( .A(n8568), .B(n8572), .ZN(n8571) );
  NAND2_X1 U8623 ( .A1(n8573), .A2(operation), .ZN(n8561) );
  XNOR2_X1 U8624 ( .A(n8574), .B(n8575), .ZN(n8573) );
  NAND2_X1 U8625 ( .A1(n8576), .A2(n8577), .ZN(n8574) );
  NAND2_X1 U8626 ( .A1(n8578), .A2(n8579), .ZN(Result_54_) );
  NAND2_X1 U8627 ( .A1(n8580), .A2(n8421), .ZN(n8579) );
  XNOR2_X1 U8628 ( .A(n8581), .B(n8582), .ZN(n8580) );
  NAND2_X1 U8629 ( .A1(n8583), .A2(n8584), .ZN(n8582) );
  NAND2_X1 U8630 ( .A1(n8585), .A2(operation), .ZN(n8578) );
  XOR2_X1 U8631 ( .A(n8586), .B(n8587), .Z(n8585) );
  XNOR2_X1 U8632 ( .A(n8588), .B(n8589), .ZN(n8586) );
  NAND2_X1 U8633 ( .A1(n8590), .A2(n8591), .ZN(Result_53_) );
  NAND2_X1 U8634 ( .A1(n8592), .A2(n8421), .ZN(n8591) );
  NAND3_X1 U8635 ( .A1(n8593), .A2(n8594), .A3(n8595), .ZN(n8592) );
  NAND2_X1 U8636 ( .A1(n8596), .A2(n8597), .ZN(n8595) );
  INV_X1 U8637 ( .A(n8598), .ZN(n8594) );
  NOR3_X1 U8638 ( .A1(n8597), .A2(a_21_), .A3(n8599), .ZN(n8598) );
  NAND2_X1 U8639 ( .A1(n8600), .A2(n8599), .ZN(n8593) );
  XNOR2_X1 U8640 ( .A(n8597), .B(n8601), .ZN(n8600) );
  NAND2_X1 U8641 ( .A1(n8602), .A2(operation), .ZN(n8590) );
  XNOR2_X1 U8642 ( .A(n8603), .B(n8604), .ZN(n8602) );
  NAND2_X1 U8643 ( .A1(n8605), .A2(n8606), .ZN(n8603) );
  NAND2_X1 U8644 ( .A1(n8607), .A2(n8608), .ZN(Result_52_) );
  NAND2_X1 U8645 ( .A1(n8609), .A2(n8421), .ZN(n8608) );
  XNOR2_X1 U8646 ( .A(n8610), .B(n8611), .ZN(n8609) );
  NAND2_X1 U8647 ( .A1(n8612), .A2(n8613), .ZN(n8611) );
  NAND2_X1 U8648 ( .A1(n8614), .A2(operation), .ZN(n8607) );
  XNOR2_X1 U8649 ( .A(n8615), .B(n8616), .ZN(n8614) );
  XOR2_X1 U8650 ( .A(n8617), .B(n8618), .Z(n8616) );
  NAND2_X1 U8651 ( .A1(n8619), .A2(n8620), .ZN(Result_51_) );
  NAND2_X1 U8652 ( .A1(n8621), .A2(n8421), .ZN(n8620) );
  NAND3_X1 U8653 ( .A1(n8622), .A2(n8623), .A3(n8624), .ZN(n8621) );
  NAND2_X1 U8654 ( .A1(n8625), .A2(n8626), .ZN(n8624) );
  INV_X1 U8655 ( .A(n8627), .ZN(n8623) );
  NOR3_X1 U8656 ( .A1(n8626), .A2(a_19_), .A3(n8628), .ZN(n8627) );
  NAND2_X1 U8657 ( .A1(n8629), .A2(n8628), .ZN(n8622) );
  XNOR2_X1 U8658 ( .A(n8626), .B(n8630), .ZN(n8629) );
  NAND2_X1 U8659 ( .A1(n8631), .A2(operation), .ZN(n8619) );
  XNOR2_X1 U8660 ( .A(n8632), .B(n8633), .ZN(n8631) );
  NAND2_X1 U8661 ( .A1(n8634), .A2(n8635), .ZN(n8632) );
  NAND2_X1 U8662 ( .A1(n8636), .A2(n8637), .ZN(Result_50_) );
  NAND2_X1 U8663 ( .A1(n8638), .A2(n8421), .ZN(n8637) );
  XNOR2_X1 U8664 ( .A(n8639), .B(n8640), .ZN(n8638) );
  NAND2_X1 U8665 ( .A1(n8641), .A2(n8642), .ZN(n8640) );
  NAND2_X1 U8666 ( .A1(n8643), .A2(operation), .ZN(n8636) );
  XNOR2_X1 U8667 ( .A(n8644), .B(n8645), .ZN(n8643) );
  XOR2_X1 U8668 ( .A(n8646), .B(n8647), .Z(n8645) );
  NAND2_X1 U8669 ( .A1(b_31_), .A2(a_18_), .ZN(n8647) );
  NOR2_X1 U8670 ( .A1(n8648), .A2(n8421), .ZN(Result_4_) );
  XNOR2_X1 U8671 ( .A(n8649), .B(n8650), .ZN(n8648) );
  NAND2_X1 U8672 ( .A1(n8651), .A2(n8652), .ZN(Result_49_) );
  NAND2_X1 U8673 ( .A1(n8653), .A2(n8421), .ZN(n8652) );
  NAND3_X1 U8674 ( .A1(n8654), .A2(n8655), .A3(n8656), .ZN(n8653) );
  NAND2_X1 U8675 ( .A1(n8657), .A2(n8658), .ZN(n8656) );
  INV_X1 U8676 ( .A(n8659), .ZN(n8655) );
  NOR3_X1 U8677 ( .A1(n8658), .A2(a_17_), .A3(n8660), .ZN(n8659) );
  NAND2_X1 U8678 ( .A1(n8661), .A2(n8660), .ZN(n8654) );
  XNOR2_X1 U8679 ( .A(n8658), .B(n8662), .ZN(n8661) );
  NAND2_X1 U8680 ( .A1(n8663), .A2(operation), .ZN(n8651) );
  XOR2_X1 U8681 ( .A(n8664), .B(n8665), .Z(n8663) );
  XOR2_X1 U8682 ( .A(n8666), .B(n8667), .Z(n8664) );
  NOR2_X1 U8683 ( .A1(n8662), .A2(n8448), .ZN(n8667) );
  NAND2_X1 U8684 ( .A1(n8668), .A2(n8669), .ZN(Result_48_) );
  NAND2_X1 U8685 ( .A1(n8670), .A2(n8421), .ZN(n8669) );
  XNOR2_X1 U8686 ( .A(n8671), .B(n8672), .ZN(n8670) );
  NAND2_X1 U8687 ( .A1(n8673), .A2(n8674), .ZN(n8672) );
  NAND2_X1 U8688 ( .A1(n8675), .A2(operation), .ZN(n8668) );
  XNOR2_X1 U8689 ( .A(n8676), .B(n8677), .ZN(n8675) );
  XNOR2_X1 U8690 ( .A(n8678), .B(n8679), .ZN(n8676) );
  NOR2_X1 U8691 ( .A1(n8680), .A2(n8448), .ZN(n8679) );
  NAND2_X1 U8692 ( .A1(n8681), .A2(n8682), .ZN(Result_47_) );
  NAND2_X1 U8693 ( .A1(n8683), .A2(n8421), .ZN(n8682) );
  NAND3_X1 U8694 ( .A1(n8684), .A2(n8685), .A3(n8686), .ZN(n8683) );
  NAND2_X1 U8695 ( .A1(n8687), .A2(n8688), .ZN(n8686) );
  INV_X1 U8696 ( .A(n8689), .ZN(n8685) );
  NOR3_X1 U8697 ( .A1(n8688), .A2(a_15_), .A3(n8690), .ZN(n8689) );
  NAND2_X1 U8698 ( .A1(n8691), .A2(n8690), .ZN(n8684) );
  XNOR2_X1 U8699 ( .A(n8688), .B(n8692), .ZN(n8691) );
  NAND2_X1 U8700 ( .A1(n8693), .A2(operation), .ZN(n8681) );
  XOR2_X1 U8701 ( .A(n8694), .B(n8695), .Z(n8693) );
  XNOR2_X1 U8702 ( .A(n8696), .B(n8697), .ZN(n8695) );
  NAND2_X1 U8703 ( .A1(b_31_), .A2(a_15_), .ZN(n8697) );
  NAND2_X1 U8704 ( .A1(n8698), .A2(n8699), .ZN(Result_46_) );
  NAND2_X1 U8705 ( .A1(n8700), .A2(n8421), .ZN(n8699) );
  XNOR2_X1 U8706 ( .A(n8701), .B(n8702), .ZN(n8700) );
  NAND2_X1 U8707 ( .A1(n8703), .A2(n8704), .ZN(n8702) );
  NAND2_X1 U8708 ( .A1(n8705), .A2(operation), .ZN(n8698) );
  XOR2_X1 U8709 ( .A(n8706), .B(n8707), .Z(n8705) );
  XNOR2_X1 U8710 ( .A(n8708), .B(n8709), .ZN(n8707) );
  NAND2_X1 U8711 ( .A1(b_31_), .A2(a_14_), .ZN(n8709) );
  NAND2_X1 U8712 ( .A1(n8710), .A2(n8711), .ZN(Result_45_) );
  NAND2_X1 U8713 ( .A1(n8712), .A2(n8421), .ZN(n8711) );
  NAND3_X1 U8714 ( .A1(n8713), .A2(n8714), .A3(n8715), .ZN(n8712) );
  NAND2_X1 U8715 ( .A1(n8716), .A2(n8717), .ZN(n8715) );
  INV_X1 U8716 ( .A(n8718), .ZN(n8714) );
  NOR3_X1 U8717 ( .A1(n8717), .A2(a_13_), .A3(n8719), .ZN(n8718) );
  NAND2_X1 U8718 ( .A1(n8720), .A2(n8719), .ZN(n8713) );
  XNOR2_X1 U8719 ( .A(n8717), .B(n8721), .ZN(n8720) );
  NAND2_X1 U8720 ( .A1(n8722), .A2(operation), .ZN(n8710) );
  XOR2_X1 U8721 ( .A(n8723), .B(n8724), .Z(n8722) );
  XNOR2_X1 U8722 ( .A(n8725), .B(n8726), .ZN(n8724) );
  NAND2_X1 U8723 ( .A1(b_31_), .A2(a_13_), .ZN(n8726) );
  NAND2_X1 U8724 ( .A1(n8727), .A2(n8728), .ZN(Result_44_) );
  NAND2_X1 U8725 ( .A1(n8729), .A2(n8421), .ZN(n8728) );
  XNOR2_X1 U8726 ( .A(n8730), .B(n8731), .ZN(n8729) );
  NOR2_X1 U8727 ( .A1(n8732), .A2(n8733), .ZN(n8731) );
  NAND2_X1 U8728 ( .A1(n8734), .A2(operation), .ZN(n8727) );
  XOR2_X1 U8729 ( .A(n8735), .B(n8736), .Z(n8734) );
  XOR2_X1 U8730 ( .A(n8737), .B(n8738), .Z(n8735) );
  NOR2_X1 U8731 ( .A1(n8739), .A2(n8448), .ZN(n8738) );
  NAND2_X1 U8732 ( .A1(n8740), .A2(n8741), .ZN(Result_43_) );
  NAND2_X1 U8733 ( .A1(n8742), .A2(n8421), .ZN(n8741) );
  NAND3_X1 U8734 ( .A1(n8743), .A2(n8744), .A3(n8745), .ZN(n8742) );
  NAND2_X1 U8735 ( .A1(n8746), .A2(n8747), .ZN(n8745) );
  NAND3_X1 U8736 ( .A1(n8748), .A2(n8749), .A3(b_11_), .ZN(n8744) );
  NAND2_X1 U8737 ( .A1(n8750), .A2(n8751), .ZN(n8743) );
  XNOR2_X1 U8738 ( .A(n8748), .B(a_11_), .ZN(n8750) );
  NAND2_X1 U8739 ( .A1(n8752), .A2(operation), .ZN(n8740) );
  XOR2_X1 U8740 ( .A(n8753), .B(n8754), .Z(n8752) );
  XNOR2_X1 U8741 ( .A(n8755), .B(n8756), .ZN(n8754) );
  NAND2_X1 U8742 ( .A1(b_31_), .A2(a_11_), .ZN(n8756) );
  NAND2_X1 U8743 ( .A1(n8757), .A2(n8758), .ZN(Result_42_) );
  NAND2_X1 U8744 ( .A1(n8759), .A2(n8421), .ZN(n8758) );
  XNOR2_X1 U8745 ( .A(n8760), .B(n8761), .ZN(n8759) );
  NAND2_X1 U8746 ( .A1(n8762), .A2(n8763), .ZN(n8761) );
  NAND2_X1 U8747 ( .A1(n8764), .A2(operation), .ZN(n8757) );
  XNOR2_X1 U8748 ( .A(n8765), .B(n8766), .ZN(n8764) );
  XNOR2_X1 U8749 ( .A(n8767), .B(n8768), .ZN(n8765) );
  NOR2_X1 U8750 ( .A1(n8769), .A2(n8448), .ZN(n8768) );
  NAND2_X1 U8751 ( .A1(n8770), .A2(n8771), .ZN(Result_41_) );
  NAND2_X1 U8752 ( .A1(n8772), .A2(n8421), .ZN(n8771) );
  NAND3_X1 U8753 ( .A1(n8773), .A2(n8774), .A3(n8775), .ZN(n8772) );
  NAND2_X1 U8754 ( .A1(n8776), .A2(n8777), .ZN(n8775) );
  NAND3_X1 U8755 ( .A1(n8778), .A2(n8779), .A3(b_9_), .ZN(n8774) );
  NAND2_X1 U8756 ( .A1(n8780), .A2(n8781), .ZN(n8773) );
  XNOR2_X1 U8757 ( .A(n8777), .B(n8779), .ZN(n8780) );
  NAND2_X1 U8758 ( .A1(n8782), .A2(operation), .ZN(n8770) );
  XOR2_X1 U8759 ( .A(n8783), .B(n8784), .Z(n8782) );
  XNOR2_X1 U8760 ( .A(n8785), .B(n8786), .ZN(n8784) );
  NAND2_X1 U8761 ( .A1(b_31_), .A2(a_9_), .ZN(n8786) );
  NAND2_X1 U8762 ( .A1(n8787), .A2(n8788), .ZN(Result_40_) );
  NAND2_X1 U8763 ( .A1(n8789), .A2(n8421), .ZN(n8788) );
  XNOR2_X1 U8764 ( .A(n8790), .B(n8791), .ZN(n8789) );
  NOR2_X1 U8765 ( .A1(n8792), .A2(n8793), .ZN(n8791) );
  NAND2_X1 U8766 ( .A1(n8794), .A2(operation), .ZN(n8787) );
  XOR2_X1 U8767 ( .A(n8795), .B(n8796), .Z(n8794) );
  XNOR2_X1 U8768 ( .A(n8797), .B(n8798), .ZN(n8796) );
  NAND2_X1 U8769 ( .A1(b_31_), .A2(a_8_), .ZN(n8798) );
  NOR2_X1 U8770 ( .A1(n8799), .A2(n8421), .ZN(Result_3_) );
  XNOR2_X1 U8771 ( .A(n8800), .B(n8801), .ZN(n8799) );
  NAND2_X1 U8772 ( .A1(n8802), .A2(n8803), .ZN(n8800) );
  NAND2_X1 U8773 ( .A1(n8804), .A2(n8805), .ZN(n8803) );
  NAND2_X1 U8774 ( .A1(n8806), .A2(n8807), .ZN(n8804) );
  NAND2_X1 U8775 ( .A1(n8808), .A2(n8809), .ZN(Result_39_) );
  NAND2_X1 U8776 ( .A1(n8810), .A2(n8421), .ZN(n8809) );
  NAND3_X1 U8777 ( .A1(n8811), .A2(n8812), .A3(n8813), .ZN(n8810) );
  NAND2_X1 U8778 ( .A1(n8814), .A2(n8815), .ZN(n8813) );
  NAND3_X1 U8779 ( .A1(n8816), .A2(n8817), .A3(b_7_), .ZN(n8812) );
  NAND2_X1 U8780 ( .A1(n8818), .A2(n8819), .ZN(n8811) );
  XNOR2_X1 U8781 ( .A(n8816), .B(a_7_), .ZN(n8818) );
  NAND2_X1 U8782 ( .A1(n8820), .A2(operation), .ZN(n8808) );
  XOR2_X1 U8783 ( .A(n8821), .B(n8822), .Z(n8820) );
  XNOR2_X1 U8784 ( .A(n8823), .B(n8824), .ZN(n8822) );
  NAND2_X1 U8785 ( .A1(b_31_), .A2(a_7_), .ZN(n8824) );
  NAND2_X1 U8786 ( .A1(n8825), .A2(n8826), .ZN(Result_38_) );
  NAND2_X1 U8787 ( .A1(n8827), .A2(n8421), .ZN(n8826) );
  XNOR2_X1 U8788 ( .A(n8828), .B(n8829), .ZN(n8827) );
  NAND2_X1 U8789 ( .A1(n8830), .A2(n8831), .ZN(n8829) );
  NAND2_X1 U8790 ( .A1(n8832), .A2(operation), .ZN(n8825) );
  XOR2_X1 U8791 ( .A(n8833), .B(n8834), .Z(n8832) );
  XNOR2_X1 U8792 ( .A(n8835), .B(n8836), .ZN(n8834) );
  NAND2_X1 U8793 ( .A1(b_31_), .A2(a_6_), .ZN(n8836) );
  NAND2_X1 U8794 ( .A1(n8837), .A2(n8838), .ZN(Result_37_) );
  NAND2_X1 U8795 ( .A1(n8839), .A2(n8421), .ZN(n8838) );
  NAND3_X1 U8796 ( .A1(n8840), .A2(n8841), .A3(n8842), .ZN(n8839) );
  NAND2_X1 U8797 ( .A1(n8843), .A2(n8844), .ZN(n8842) );
  INV_X1 U8798 ( .A(n8845), .ZN(n8841) );
  NOR3_X1 U8799 ( .A1(n8844), .A2(a_5_), .A3(n8846), .ZN(n8845) );
  NAND2_X1 U8800 ( .A1(n8847), .A2(n8846), .ZN(n8840) );
  XNOR2_X1 U8801 ( .A(n8844), .B(n8848), .ZN(n8847) );
  NAND2_X1 U8802 ( .A1(n8849), .A2(operation), .ZN(n8837) );
  XOR2_X1 U8803 ( .A(n8850), .B(n8851), .Z(n8849) );
  XNOR2_X1 U8804 ( .A(n8852), .B(n8853), .ZN(n8851) );
  NAND2_X1 U8805 ( .A1(b_31_), .A2(a_5_), .ZN(n8853) );
  NAND2_X1 U8806 ( .A1(n8854), .A2(n8855), .ZN(Result_36_) );
  NAND2_X1 U8807 ( .A1(n8856), .A2(n8421), .ZN(n8855) );
  XNOR2_X1 U8808 ( .A(n8857), .B(n8858), .ZN(n8856) );
  NAND2_X1 U8809 ( .A1(n8859), .A2(n8860), .ZN(n8858) );
  NAND2_X1 U8810 ( .A1(n8861), .A2(operation), .ZN(n8854) );
  XOR2_X1 U8811 ( .A(n8862), .B(n8863), .Z(n8861) );
  XNOR2_X1 U8812 ( .A(n8864), .B(n8865), .ZN(n8863) );
  NAND2_X1 U8813 ( .A1(b_31_), .A2(a_4_), .ZN(n8865) );
  NAND2_X1 U8814 ( .A1(n8866), .A2(n8867), .ZN(Result_35_) );
  NAND2_X1 U8815 ( .A1(n8868), .A2(n8421), .ZN(n8867) );
  NAND3_X1 U8816 ( .A1(n8869), .A2(n8870), .A3(n8871), .ZN(n8868) );
  NAND2_X1 U8817 ( .A1(n8872), .A2(n8873), .ZN(n8871) );
  INV_X1 U8818 ( .A(n8874), .ZN(n8870) );
  NOR3_X1 U8819 ( .A1(n8873), .A2(a_3_), .A3(n8875), .ZN(n8874) );
  NAND2_X1 U8820 ( .A1(n8876), .A2(n8875), .ZN(n8869) );
  XNOR2_X1 U8821 ( .A(n8873), .B(n8877), .ZN(n8876) );
  NAND2_X1 U8822 ( .A1(n8878), .A2(operation), .ZN(n8866) );
  XNOR2_X1 U8823 ( .A(n8879), .B(n8880), .ZN(n8878) );
  XNOR2_X1 U8824 ( .A(n8881), .B(n8882), .ZN(n8879) );
  NOR2_X1 U8825 ( .A1(n8877), .A2(n8448), .ZN(n8882) );
  NAND2_X1 U8826 ( .A1(n8883), .A2(n8884), .ZN(Result_34_) );
  NAND2_X1 U8827 ( .A1(n8885), .A2(n8421), .ZN(n8884) );
  XNOR2_X1 U8828 ( .A(n8886), .B(n8887), .ZN(n8885) );
  NAND2_X1 U8829 ( .A1(n8888), .A2(n8889), .ZN(n8887) );
  NAND2_X1 U8830 ( .A1(n8890), .A2(operation), .ZN(n8883) );
  XOR2_X1 U8831 ( .A(n8891), .B(n8892), .Z(n8890) );
  XNOR2_X1 U8832 ( .A(n8893), .B(n8894), .ZN(n8892) );
  NAND2_X1 U8833 ( .A1(b_31_), .A2(a_2_), .ZN(n8894) );
  NAND2_X1 U8834 ( .A1(n8895), .A2(n8896), .ZN(Result_33_) );
  NAND2_X1 U8835 ( .A1(n8897), .A2(n8421), .ZN(n8896) );
  NAND2_X1 U8836 ( .A1(n8898), .A2(n8899), .ZN(n8897) );
  INV_X1 U8837 ( .A(n8900), .ZN(n8899) );
  NOR2_X1 U8838 ( .A1(n8901), .A2(n8902), .ZN(n8900) );
  NOR2_X1 U8839 ( .A1(n8903), .A2(n8904), .ZN(n8901) );
  NAND2_X1 U8840 ( .A1(n8905), .A2(n8902), .ZN(n8898) );
  INV_X1 U8841 ( .A(n8906), .ZN(n8902) );
  XNOR2_X1 U8842 ( .A(n8907), .B(a_1_), .ZN(n8905) );
  NAND2_X1 U8843 ( .A1(n8908), .A2(operation), .ZN(n8895) );
  XOR2_X1 U8844 ( .A(n8909), .B(n8910), .Z(n8908) );
  XNOR2_X1 U8845 ( .A(n8911), .B(n8912), .ZN(n8910) );
  NAND2_X1 U8846 ( .A1(b_31_), .A2(a_1_), .ZN(n8912) );
  NAND2_X1 U8847 ( .A1(n8913), .A2(n8914), .ZN(Result_32_) );
  NAND2_X1 U8848 ( .A1(n8915), .A2(n8421), .ZN(n8914) );
  XOR2_X1 U8849 ( .A(n8916), .B(n8917), .Z(n8915) );
  NOR2_X1 U8850 ( .A1(n8918), .A2(n8919), .ZN(n8917) );
  NOR2_X1 U8851 ( .A1(b_0_), .A2(a_0_), .ZN(n8918) );
  NOR2_X1 U8852 ( .A1(n8904), .A2(n8920), .ZN(n8916) );
  NOR2_X1 U8853 ( .A1(n8903), .A2(n8906), .ZN(n8920) );
  NAND2_X1 U8854 ( .A1(n8889), .A2(n8921), .ZN(n8906) );
  NAND2_X1 U8855 ( .A1(n8888), .A2(n8886), .ZN(n8921) );
  NAND2_X1 U8856 ( .A1(n8922), .A2(n8923), .ZN(n8886) );
  NAND2_X1 U8857 ( .A1(n8924), .A2(n8873), .ZN(n8923) );
  NAND2_X1 U8858 ( .A1(n8860), .A2(n8925), .ZN(n8873) );
  NAND2_X1 U8859 ( .A1(n8859), .A2(n8857), .ZN(n8925) );
  NAND2_X1 U8860 ( .A1(n8926), .A2(n8927), .ZN(n8857) );
  NAND2_X1 U8861 ( .A1(n8928), .A2(n8844), .ZN(n8927) );
  NAND2_X1 U8862 ( .A1(n8831), .A2(n8929), .ZN(n8844) );
  NAND2_X1 U8863 ( .A1(n8830), .A2(n8828), .ZN(n8929) );
  NAND2_X1 U8864 ( .A1(n8930), .A2(n8931), .ZN(n8828) );
  NAND2_X1 U8865 ( .A1(n8932), .A2(n8815), .ZN(n8931) );
  INV_X1 U8866 ( .A(n8816), .ZN(n8815) );
  NOR2_X1 U8867 ( .A1(n8793), .A2(n8933), .ZN(n8816) );
  NOR2_X1 U8868 ( .A1(n8792), .A2(n8790), .ZN(n8933) );
  NOR2_X1 U8869 ( .A1(n8776), .A2(n8934), .ZN(n8790) );
  NOR2_X1 U8870 ( .A1(n8935), .A2(n8778), .ZN(n8934) );
  INV_X1 U8871 ( .A(n8777), .ZN(n8778) );
  NAND2_X1 U8872 ( .A1(n8763), .A2(n8936), .ZN(n8777) );
  NAND2_X1 U8873 ( .A1(n8762), .A2(n8760), .ZN(n8936) );
  NAND2_X1 U8874 ( .A1(n8937), .A2(n8938), .ZN(n8760) );
  NAND2_X1 U8875 ( .A1(n8939), .A2(n8747), .ZN(n8938) );
  INV_X1 U8876 ( .A(n8748), .ZN(n8747) );
  NOR2_X1 U8877 ( .A1(n8733), .A2(n8940), .ZN(n8748) );
  NOR2_X1 U8878 ( .A1(n8732), .A2(n8730), .ZN(n8940) );
  NOR2_X1 U8879 ( .A1(n8716), .A2(n8941), .ZN(n8730) );
  INV_X1 U8880 ( .A(n8942), .ZN(n8941) );
  NAND2_X1 U8881 ( .A1(n8943), .A2(n8717), .ZN(n8942) );
  NAND2_X1 U8882 ( .A1(n8704), .A2(n8944), .ZN(n8717) );
  NAND2_X1 U8883 ( .A1(n8703), .A2(n8701), .ZN(n8944) );
  NAND2_X1 U8884 ( .A1(n8945), .A2(n8946), .ZN(n8701) );
  NAND2_X1 U8885 ( .A1(n8947), .A2(n8688), .ZN(n8946) );
  NAND2_X1 U8886 ( .A1(n8674), .A2(n8948), .ZN(n8688) );
  NAND2_X1 U8887 ( .A1(n8673), .A2(n8671), .ZN(n8948) );
  NAND2_X1 U8888 ( .A1(n8949), .A2(n8950), .ZN(n8671) );
  NAND2_X1 U8889 ( .A1(n8951), .A2(n8658), .ZN(n8950) );
  NAND2_X1 U8890 ( .A1(n8642), .A2(n8952), .ZN(n8658) );
  NAND2_X1 U8891 ( .A1(n8641), .A2(n8639), .ZN(n8952) );
  NAND2_X1 U8892 ( .A1(n8953), .A2(n8954), .ZN(n8639) );
  NAND2_X1 U8893 ( .A1(n8955), .A2(n8626), .ZN(n8954) );
  NAND2_X1 U8894 ( .A1(n8613), .A2(n8956), .ZN(n8626) );
  NAND2_X1 U8895 ( .A1(n8612), .A2(n8610), .ZN(n8956) );
  NAND2_X1 U8896 ( .A1(n8957), .A2(n8958), .ZN(n8610) );
  NAND2_X1 U8897 ( .A1(n8959), .A2(n8597), .ZN(n8958) );
  NAND2_X1 U8898 ( .A1(n8584), .A2(n8960), .ZN(n8597) );
  NAND2_X1 U8899 ( .A1(n8583), .A2(n8581), .ZN(n8960) );
  NAND2_X1 U8900 ( .A1(n8961), .A2(n8962), .ZN(n8581) );
  NAND2_X1 U8901 ( .A1(n8963), .A2(n8568), .ZN(n8962) );
  NAND2_X1 U8902 ( .A1(n8555), .A2(n8964), .ZN(n8568) );
  NAND2_X1 U8903 ( .A1(n8554), .A2(n8552), .ZN(n8964) );
  NAND2_X1 U8904 ( .A1(n8965), .A2(n8966), .ZN(n8552) );
  NAND2_X1 U8905 ( .A1(n8967), .A2(n8539), .ZN(n8966) );
  INV_X1 U8906 ( .A(n8540), .ZN(n8539) );
  NOR2_X1 U8907 ( .A1(n8526), .A2(n8968), .ZN(n8540) );
  NOR2_X1 U8908 ( .A1(n8525), .A2(n8523), .ZN(n8968) );
  NOR2_X1 U8909 ( .A1(n8509), .A2(n8969), .ZN(n8523) );
  NOR2_X1 U8910 ( .A1(n8970), .A2(n8511), .ZN(n8969) );
  INV_X1 U8911 ( .A(n8510), .ZN(n8511) );
  NAND2_X1 U8912 ( .A1(n8486), .A2(n8971), .ZN(n8510) );
  NAND2_X1 U8913 ( .A1(n8487), .A2(n8485), .ZN(n8971) );
  NAND2_X1 U8914 ( .A1(n8972), .A2(n8973), .ZN(n8485) );
  NAND2_X1 U8915 ( .A1(n8974), .A2(n8471), .ZN(n8973) );
  INV_X1 U8916 ( .A(n8472), .ZN(n8471) );
  NOR2_X1 U8917 ( .A1(n8975), .A2(n8976), .ZN(n8472) );
  NOR2_X1 U8918 ( .A1(n8461), .A2(n8977), .ZN(n8976) );
  NOR2_X1 U8919 ( .A1(a_30_), .A2(n8449), .ZN(n8977) );
  NOR2_X1 U8920 ( .A1(n8448), .A2(n8978), .ZN(n8449) );
  NOR2_X1 U8921 ( .A1(n8448), .A2(n8979), .ZN(n8975) );
  NAND2_X1 U8922 ( .A1(n8475), .A2(n8473), .ZN(n8974) );
  NAND2_X1 U8923 ( .A1(n8980), .A2(n8493), .ZN(n8487) );
  NOR2_X1 U8924 ( .A1(b_27_), .A2(a_27_), .ZN(n8970) );
  NOR2_X1 U8925 ( .A1(b_26_), .A2(a_26_), .ZN(n8525) );
  NAND2_X1 U8926 ( .A1(n8543), .A2(n8541), .ZN(n8967) );
  NAND2_X1 U8927 ( .A1(n8981), .A2(n8982), .ZN(n8554) );
  NAND2_X1 U8928 ( .A1(n8570), .A2(n8572), .ZN(n8963) );
  NAND2_X1 U8929 ( .A1(n8983), .A2(n8984), .ZN(n8583) );
  NAND2_X1 U8930 ( .A1(n8599), .A2(n8601), .ZN(n8959) );
  INV_X1 U8931 ( .A(n8596), .ZN(n8957) );
  NAND2_X1 U8932 ( .A1(n8985), .A2(n8986), .ZN(n8612) );
  NAND2_X1 U8933 ( .A1(n8628), .A2(n8630), .ZN(n8955) );
  NAND2_X1 U8934 ( .A1(n8987), .A2(n8988), .ZN(n8641) );
  NAND2_X1 U8935 ( .A1(n8660), .A2(n8662), .ZN(n8951) );
  NAND2_X1 U8936 ( .A1(n8989), .A2(n8680), .ZN(n8673) );
  NAND2_X1 U8937 ( .A1(n8690), .A2(n8692), .ZN(n8947) );
  NAND2_X1 U8938 ( .A1(n8990), .A2(n8991), .ZN(n8703) );
  NAND2_X1 U8939 ( .A1(n8719), .A2(n8721), .ZN(n8943) );
  NOR2_X1 U8940 ( .A1(b_12_), .A2(a_12_), .ZN(n8732) );
  NAND2_X1 U8941 ( .A1(n8751), .A2(n8749), .ZN(n8939) );
  NAND2_X1 U8942 ( .A1(n8992), .A2(n8769), .ZN(n8762) );
  NOR2_X1 U8943 ( .A1(b_9_), .A2(a_9_), .ZN(n8935) );
  NOR2_X1 U8944 ( .A1(b_8_), .A2(a_8_), .ZN(n8792) );
  NAND2_X1 U8945 ( .A1(n8819), .A2(n8817), .ZN(n8932) );
  NAND2_X1 U8946 ( .A1(n8993), .A2(n8994), .ZN(n8830) );
  NAND2_X1 U8947 ( .A1(n8846), .A2(n8848), .ZN(n8928) );
  NAND2_X1 U8948 ( .A1(n8995), .A2(n8996), .ZN(n8859) );
  NAND2_X1 U8949 ( .A1(n8875), .A2(n8877), .ZN(n8924) );
  NAND2_X1 U8950 ( .A1(n8997), .A2(n8998), .ZN(n8888) );
  NOR2_X1 U8951 ( .A1(b_1_), .A2(a_1_), .ZN(n8904) );
  NAND2_X1 U8952 ( .A1(n8999), .A2(operation), .ZN(n8913) );
  XOR2_X1 U8953 ( .A(n9000), .B(n9001), .Z(n8999) );
  XNOR2_X1 U8954 ( .A(n9002), .B(n9003), .ZN(n9001) );
  NAND2_X1 U8955 ( .A1(b_31_), .A2(a_0_), .ZN(n9003) );
  NOR2_X1 U8956 ( .A1(n8421), .A2(n9004), .ZN(Result_31_) );
  XNOR2_X1 U8957 ( .A(n9005), .B(n9006), .ZN(n9004) );
  NOR3_X1 U8958 ( .A1(n8421), .A2(n9007), .A3(n9008), .ZN(Result_30_) );
  NOR2_X1 U8959 ( .A1(n9009), .A2(n9010), .ZN(n9008) );
  XOR2_X1 U8960 ( .A(n9011), .B(n9012), .Z(n9010) );
  NOR2_X1 U8961 ( .A1(n9005), .A2(n9006), .ZN(n9009) );
  NOR2_X1 U8962 ( .A1(n8421), .A2(n9013), .ZN(Result_2_) );
  XNOR2_X1 U8963 ( .A(n9014), .B(n9015), .ZN(n9013) );
  NOR2_X1 U8964 ( .A1(n9016), .A2(n8421), .ZN(Result_29_) );
  XOR2_X1 U8965 ( .A(n9017), .B(n9007), .Z(n9016) );
  NAND2_X1 U8966 ( .A1(n9018), .A2(n9019), .ZN(n9017) );
  NOR2_X1 U8967 ( .A1(n8421), .A2(n9020), .ZN(Result_28_) );
  XOR2_X1 U8968 ( .A(n9021), .B(n9022), .Z(n9020) );
  NAND2_X1 U8969 ( .A1(n9023), .A2(n9024), .ZN(n9022) );
  NOR2_X1 U8970 ( .A1(n8421), .A2(n9025), .ZN(Result_27_) );
  XOR2_X1 U8971 ( .A(n9026), .B(n9027), .Z(n9025) );
  NAND2_X1 U8972 ( .A1(n9028), .A2(n9029), .ZN(n9027) );
  NOR2_X1 U8973 ( .A1(n8421), .A2(n9030), .ZN(Result_26_) );
  XOR2_X1 U8974 ( .A(n9031), .B(n9032), .Z(n9030) );
  NAND2_X1 U8975 ( .A1(n9033), .A2(n9034), .ZN(n9032) );
  NAND2_X1 U8976 ( .A1(n9035), .A2(n9036), .ZN(n9034) );
  INV_X1 U8977 ( .A(n9037), .ZN(n9035) );
  NOR2_X1 U8978 ( .A1(n8421), .A2(n9038), .ZN(Result_25_) );
  XOR2_X1 U8979 ( .A(n9039), .B(n9040), .Z(n9038) );
  NAND2_X1 U8980 ( .A1(n9041), .A2(n9042), .ZN(n9040) );
  NOR2_X1 U8981 ( .A1(n8421), .A2(n9043), .ZN(Result_24_) );
  XOR2_X1 U8982 ( .A(n9044), .B(n9045), .Z(n9043) );
  NAND2_X1 U8983 ( .A1(n9046), .A2(n9047), .ZN(n9045) );
  NOR2_X1 U8984 ( .A1(n8421), .A2(n9048), .ZN(Result_23_) );
  XOR2_X1 U8985 ( .A(n9049), .B(n9050), .Z(n9048) );
  NAND2_X1 U8986 ( .A1(n9051), .A2(n9052), .ZN(n9050) );
  NOR2_X1 U8987 ( .A1(n8421), .A2(n9053), .ZN(Result_22_) );
  XOR2_X1 U8988 ( .A(n9054), .B(n9055), .Z(n9053) );
  NAND2_X1 U8989 ( .A1(n9056), .A2(n9057), .ZN(n9055) );
  NOR2_X1 U8990 ( .A1(n8421), .A2(n9058), .ZN(Result_21_) );
  XOR2_X1 U8991 ( .A(n9059), .B(n9060), .Z(n9058) );
  NAND2_X1 U8992 ( .A1(n9061), .A2(n9062), .ZN(n9060) );
  NOR2_X1 U8993 ( .A1(n8421), .A2(n9063), .ZN(Result_20_) );
  XOR2_X1 U8994 ( .A(n9064), .B(n9065), .Z(n9063) );
  NAND2_X1 U8995 ( .A1(n9066), .A2(n9067), .ZN(n9065) );
  NOR2_X1 U8996 ( .A1(n9068), .A2(n8421), .ZN(Result_1_) );
  XNOR2_X1 U8997 ( .A(n9069), .B(n9070), .ZN(n9068) );
  NAND2_X1 U8998 ( .A1(n9071), .A2(n9072), .ZN(n9069) );
  NOR2_X1 U8999 ( .A1(n8421), .A2(n9073), .ZN(Result_19_) );
  XOR2_X1 U9000 ( .A(n9074), .B(n9075), .Z(n9073) );
  NAND2_X1 U9001 ( .A1(n9076), .A2(n9077), .ZN(n9075) );
  NOR2_X1 U9002 ( .A1(n8421), .A2(n9078), .ZN(Result_18_) );
  XOR2_X1 U9003 ( .A(n9079), .B(n9080), .Z(n9078) );
  NAND2_X1 U9004 ( .A1(n9081), .A2(n9082), .ZN(n9080) );
  NOR2_X1 U9005 ( .A1(n8421), .A2(n9083), .ZN(Result_17_) );
  XOR2_X1 U9006 ( .A(n9084), .B(n9085), .Z(n9083) );
  NAND2_X1 U9007 ( .A1(n9086), .A2(n9087), .ZN(n9085) );
  NAND2_X1 U9008 ( .A1(n9088), .A2(n9089), .ZN(n9087) );
  INV_X1 U9009 ( .A(n9090), .ZN(n9089) );
  NAND2_X1 U9010 ( .A1(n9091), .A2(n9092), .ZN(n9088) );
  NOR2_X1 U9011 ( .A1(n8421), .A2(n9093), .ZN(Result_16_) );
  XOR2_X1 U9012 ( .A(n9094), .B(n9095), .Z(n9093) );
  NAND2_X1 U9013 ( .A1(n9096), .A2(n9097), .ZN(n9095) );
  NOR2_X1 U9014 ( .A1(n8421), .A2(n9098), .ZN(Result_15_) );
  XOR2_X1 U9015 ( .A(n9099), .B(n9100), .Z(n9098) );
  NAND2_X1 U9016 ( .A1(n9101), .A2(n9102), .ZN(n9100) );
  NOR2_X1 U9017 ( .A1(n9103), .A2(n8421), .ZN(Result_14_) );
  XNOR2_X1 U9018 ( .A(n9104), .B(n9105), .ZN(n9103) );
  NOR2_X1 U9019 ( .A1(n9106), .A2(n8421), .ZN(Result_13_) );
  XOR2_X1 U9020 ( .A(n9107), .B(n9108), .Z(n9106) );
  NAND2_X1 U9021 ( .A1(n9109), .A2(n9110), .ZN(n9107) );
  NAND2_X1 U9022 ( .A1(n9111), .A2(n9112), .ZN(n9110) );
  NAND2_X1 U9023 ( .A1(n9113), .A2(n9114), .ZN(n9111) );
  NOR2_X1 U9024 ( .A1(n9115), .A2(n8421), .ZN(Result_12_) );
  XNOR2_X1 U9025 ( .A(n9116), .B(n9117), .ZN(n9115) );
  NOR2_X1 U9026 ( .A1(n9118), .A2(n8421), .ZN(Result_11_) );
  XOR2_X1 U9027 ( .A(n9119), .B(n9120), .Z(n9118) );
  NAND2_X1 U9028 ( .A1(n9121), .A2(n9122), .ZN(n9119) );
  NAND2_X1 U9029 ( .A1(n9123), .A2(n9124), .ZN(n9122) );
  NAND2_X1 U9030 ( .A1(n9125), .A2(n9126), .ZN(n9123) );
  NOR2_X1 U9031 ( .A1(n8421), .A2(n9127), .ZN(Result_10_) );
  XNOR2_X1 U9032 ( .A(n9128), .B(n9129), .ZN(n9127) );
  NOR2_X1 U9033 ( .A1(n9130), .A2(n8421), .ZN(Result_0_) );
  NOR3_X1 U9034 ( .A1(n9131), .A2(n9132), .A3(n9133), .ZN(n9130) );
  NOR2_X1 U9035 ( .A1(n9134), .A2(n9070), .ZN(n9133) );
  NAND2_X1 U9036 ( .A1(n9015), .A2(n9014), .ZN(n9070) );
  NAND2_X1 U9037 ( .A1(n9135), .A2(n9136), .ZN(n9014) );
  NOR2_X1 U9038 ( .A1(n9137), .A2(n9138), .ZN(n9135) );
  NOR2_X1 U9039 ( .A1(n8801), .A2(n8805), .ZN(n9138) );
  NAND2_X1 U9040 ( .A1(n8649), .A2(n8650), .ZN(n8801) );
  NAND2_X1 U9041 ( .A1(n9139), .A2(n9140), .ZN(n8650) );
  NOR2_X1 U9042 ( .A1(n9141), .A2(n9142), .ZN(n9139) );
  NOR2_X1 U9043 ( .A1(n8496), .A2(n8500), .ZN(n9142) );
  NAND2_X1 U9044 ( .A1(n8443), .A2(n8444), .ZN(n8496) );
  NAND2_X1 U9045 ( .A1(n9143), .A2(n9144), .ZN(n8444) );
  NOR2_X1 U9046 ( .A1(n9145), .A2(n9146), .ZN(n9143) );
  NOR2_X1 U9047 ( .A1(n8435), .A2(n8439), .ZN(n9146) );
  NAND2_X1 U9048 ( .A1(n8431), .A2(n8432), .ZN(n8435) );
  NAND2_X1 U9049 ( .A1(n9147), .A2(n9148), .ZN(n8432) );
  INV_X1 U9050 ( .A(n9149), .ZN(n9147) );
  NAND2_X1 U9051 ( .A1(n8424), .A2(n9150), .ZN(n9149) );
  NAND2_X1 U9052 ( .A1(n8423), .A2(n9151), .ZN(n9150) );
  NOR2_X1 U9053 ( .A1(n9129), .A2(n9128), .ZN(n8423) );
  NOR2_X1 U9054 ( .A1(n9152), .A2(n9153), .ZN(n9128) );
  NAND2_X1 U9055 ( .A1(n9121), .A2(n9154), .ZN(n9153) );
  NAND2_X1 U9056 ( .A1(n9155), .A2(n9120), .ZN(n9154) );
  NOR2_X1 U9057 ( .A1(n9116), .A2(n9117), .ZN(n9120) );
  NOR2_X1 U9058 ( .A1(n9156), .A2(n9157), .ZN(n9117) );
  NAND2_X1 U9059 ( .A1(n9109), .A2(n9158), .ZN(n9157) );
  NAND2_X1 U9060 ( .A1(n9159), .A2(n9108), .ZN(n9158) );
  NOR2_X1 U9061 ( .A1(n9104), .A2(n9105), .ZN(n9108) );
  NOR2_X1 U9062 ( .A1(n9160), .A2(n9161), .ZN(n9105) );
  NAND2_X1 U9063 ( .A1(n9101), .A2(n9162), .ZN(n9161) );
  NAND2_X1 U9064 ( .A1(n9102), .A2(n9099), .ZN(n9162) );
  NAND2_X1 U9065 ( .A1(n9096), .A2(n9163), .ZN(n9099) );
  NAND2_X1 U9066 ( .A1(n9097), .A2(n9094), .ZN(n9163) );
  NAND2_X1 U9067 ( .A1(n9086), .A2(n9164), .ZN(n9094) );
  NAND2_X1 U9068 ( .A1(n9090), .A2(n9084), .ZN(n9164) );
  NAND2_X1 U9069 ( .A1(n9165), .A2(n9082), .ZN(n9084) );
  NAND2_X1 U9070 ( .A1(n9166), .A2(n9167), .ZN(n9082) );
  NAND2_X1 U9071 ( .A1(n9079), .A2(n9081), .ZN(n9165) );
  INV_X1 U9072 ( .A(n9168), .ZN(n9081) );
  NOR2_X1 U9073 ( .A1(n9167), .A2(n9166), .ZN(n9168) );
  XOR2_X1 U9074 ( .A(n9092), .B(n9091), .Z(n9167) );
  NAND2_X1 U9075 ( .A1(n9077), .A2(n9169), .ZN(n9079) );
  NAND2_X1 U9076 ( .A1(n9074), .A2(n9076), .ZN(n9169) );
  NAND2_X1 U9077 ( .A1(n9170), .A2(n9171), .ZN(n9076) );
  NAND2_X1 U9078 ( .A1(n9172), .A2(n9173), .ZN(n9171) );
  NAND2_X1 U9079 ( .A1(n9174), .A2(n9175), .ZN(n9170) );
  NAND2_X1 U9080 ( .A1(n9067), .A2(n9176), .ZN(n9074) );
  NAND2_X1 U9081 ( .A1(n9064), .A2(n9066), .ZN(n9176) );
  NAND2_X1 U9082 ( .A1(n9177), .A2(n9178), .ZN(n9066) );
  NAND2_X1 U9083 ( .A1(n9179), .A2(n9180), .ZN(n9178) );
  XNOR2_X1 U9084 ( .A(n9175), .B(n9174), .ZN(n9177) );
  NAND2_X1 U9085 ( .A1(n9062), .A2(n9181), .ZN(n9064) );
  NAND2_X1 U9086 ( .A1(n9061), .A2(n9059), .ZN(n9181) );
  NAND2_X1 U9087 ( .A1(n9182), .A2(n9057), .ZN(n9059) );
  NAND2_X1 U9088 ( .A1(n9183), .A2(n9184), .ZN(n9057) );
  NAND2_X1 U9089 ( .A1(n9054), .A2(n9056), .ZN(n9182) );
  INV_X1 U9090 ( .A(n9185), .ZN(n9056) );
  NOR2_X1 U9091 ( .A1(n9184), .A2(n9183), .ZN(n9185) );
  XOR2_X1 U9092 ( .A(n9186), .B(n9187), .Z(n9184) );
  NAND2_X1 U9093 ( .A1(n9052), .A2(n9188), .ZN(n9054) );
  NAND2_X1 U9094 ( .A1(n9049), .A2(n9051), .ZN(n9188) );
  NAND2_X1 U9095 ( .A1(n9189), .A2(n9190), .ZN(n9051) );
  NAND2_X1 U9096 ( .A1(n9191), .A2(n9192), .ZN(n9190) );
  NAND2_X1 U9097 ( .A1(n9193), .A2(n9194), .ZN(n9189) );
  NAND2_X1 U9098 ( .A1(n9047), .A2(n9195), .ZN(n9049) );
  NAND2_X1 U9099 ( .A1(n9044), .A2(n9046), .ZN(n9195) );
  NAND2_X1 U9100 ( .A1(n9196), .A2(n9197), .ZN(n9046) );
  XNOR2_X1 U9101 ( .A(n9194), .B(n9193), .ZN(n9196) );
  NAND2_X1 U9102 ( .A1(n9042), .A2(n9198), .ZN(n9044) );
  NAND2_X1 U9103 ( .A1(n9039), .A2(n9041), .ZN(n9198) );
  NAND2_X1 U9104 ( .A1(n9199), .A2(n9200), .ZN(n9041) );
  NAND2_X1 U9105 ( .A1(n9201), .A2(n9197), .ZN(n9200) );
  NAND2_X1 U9106 ( .A1(n9202), .A2(n9203), .ZN(n9199) );
  NAND2_X1 U9107 ( .A1(n9033), .A2(n9204), .ZN(n9039) );
  NAND2_X1 U9108 ( .A1(n9037), .A2(n9031), .ZN(n9204) );
  NAND2_X1 U9109 ( .A1(n9028), .A2(n9205), .ZN(n9031) );
  NAND2_X1 U9110 ( .A1(n9026), .A2(n9029), .ZN(n9205) );
  NAND2_X1 U9111 ( .A1(n9206), .A2(n9207), .ZN(n9029) );
  NAND2_X1 U9112 ( .A1(n9208), .A2(n9036), .ZN(n9207) );
  NAND2_X1 U9113 ( .A1(n9209), .A2(n9210), .ZN(n9206) );
  NAND2_X1 U9114 ( .A1(n9023), .A2(n9211), .ZN(n9026) );
  NAND2_X1 U9115 ( .A1(n9021), .A2(n9024), .ZN(n9211) );
  NAND2_X1 U9116 ( .A1(n9212), .A2(n9213), .ZN(n9024) );
  NAND2_X1 U9117 ( .A1(n9214), .A2(n9215), .ZN(n9213) );
  XNOR2_X1 U9118 ( .A(n9210), .B(n9209), .ZN(n9212) );
  NAND2_X1 U9119 ( .A1(n9019), .A2(n9216), .ZN(n9021) );
  NAND2_X1 U9120 ( .A1(n9007), .A2(n9018), .ZN(n9216) );
  NAND2_X1 U9121 ( .A1(n9217), .A2(n9218), .ZN(n9018) );
  NAND2_X1 U9122 ( .A1(n9012), .A2(n9011), .ZN(n9218) );
  XNOR2_X1 U9123 ( .A(n9215), .B(n9214), .ZN(n9217) );
  NOR3_X1 U9124 ( .A1(n9219), .A2(n9005), .A3(n9006), .ZN(n9007) );
  XOR2_X1 U9125 ( .A(n9220), .B(n9221), .Z(n9006) );
  XOR2_X1 U9126 ( .A(n9222), .B(n9223), .Z(n9221) );
  NAND2_X1 U9127 ( .A1(b_30_), .A2(a_0_), .ZN(n9223) );
  NOR2_X1 U9128 ( .A1(n9224), .A2(n9225), .ZN(n9005) );
  INV_X1 U9129 ( .A(n9226), .ZN(n9225) );
  NAND3_X1 U9130 ( .A1(a_0_), .A2(n9227), .A3(b_31_), .ZN(n9226) );
  NAND2_X1 U9131 ( .A1(n9002), .A2(n9000), .ZN(n9227) );
  NOR2_X1 U9132 ( .A1(n9000), .A2(n9002), .ZN(n9224) );
  NOR2_X1 U9133 ( .A1(n9228), .A2(n9229), .ZN(n9002) );
  INV_X1 U9134 ( .A(n9230), .ZN(n9229) );
  NAND3_X1 U9135 ( .A1(a_1_), .A2(n9231), .A3(b_31_), .ZN(n9230) );
  NAND2_X1 U9136 ( .A1(n8911), .A2(n8909), .ZN(n9231) );
  NOR2_X1 U9137 ( .A1(n8909), .A2(n8911), .ZN(n9228) );
  NOR2_X1 U9138 ( .A1(n9232), .A2(n9233), .ZN(n8911) );
  INV_X1 U9139 ( .A(n9234), .ZN(n9233) );
  NAND3_X1 U9140 ( .A1(a_2_), .A2(n9235), .A3(b_31_), .ZN(n9234) );
  NAND2_X1 U9141 ( .A1(n8893), .A2(n8891), .ZN(n9235) );
  NOR2_X1 U9142 ( .A1(n8891), .A2(n8893), .ZN(n9232) );
  NOR2_X1 U9143 ( .A1(n9236), .A2(n9237), .ZN(n8893) );
  NOR3_X1 U9144 ( .A1(n8877), .A2(n9238), .A3(n8448), .ZN(n9237) );
  INV_X1 U9145 ( .A(n9239), .ZN(n9238) );
  NAND2_X1 U9146 ( .A1(n8881), .A2(n8880), .ZN(n9239) );
  NOR2_X1 U9147 ( .A1(n8880), .A2(n8881), .ZN(n9236) );
  NOR2_X1 U9148 ( .A1(n9240), .A2(n9241), .ZN(n8881) );
  INV_X1 U9149 ( .A(n9242), .ZN(n9241) );
  NAND3_X1 U9150 ( .A1(a_4_), .A2(n9243), .A3(b_31_), .ZN(n9242) );
  NAND2_X1 U9151 ( .A1(n8864), .A2(n8862), .ZN(n9243) );
  NOR2_X1 U9152 ( .A1(n8862), .A2(n8864), .ZN(n9240) );
  NOR2_X1 U9153 ( .A1(n9244), .A2(n9245), .ZN(n8864) );
  NOR3_X1 U9154 ( .A1(n8848), .A2(n9246), .A3(n8448), .ZN(n9245) );
  INV_X1 U9155 ( .A(n9247), .ZN(n9246) );
  NAND2_X1 U9156 ( .A1(n8852), .A2(n8850), .ZN(n9247) );
  NOR2_X1 U9157 ( .A1(n8850), .A2(n8852), .ZN(n9244) );
  NOR2_X1 U9158 ( .A1(n9248), .A2(n9249), .ZN(n8852) );
  INV_X1 U9159 ( .A(n9250), .ZN(n9249) );
  NAND3_X1 U9160 ( .A1(a_6_), .A2(n9251), .A3(b_31_), .ZN(n9250) );
  NAND2_X1 U9161 ( .A1(n8835), .A2(n8833), .ZN(n9251) );
  NOR2_X1 U9162 ( .A1(n8833), .A2(n8835), .ZN(n9248) );
  NOR2_X1 U9163 ( .A1(n9252), .A2(n9253), .ZN(n8835) );
  INV_X1 U9164 ( .A(n9254), .ZN(n9253) );
  NAND3_X1 U9165 ( .A1(a_7_), .A2(n9255), .A3(b_31_), .ZN(n9254) );
  NAND2_X1 U9166 ( .A1(n8823), .A2(n8821), .ZN(n9255) );
  NOR2_X1 U9167 ( .A1(n8821), .A2(n8823), .ZN(n9252) );
  NOR2_X1 U9168 ( .A1(n9256), .A2(n9257), .ZN(n8823) );
  INV_X1 U9169 ( .A(n9258), .ZN(n9257) );
  NAND3_X1 U9170 ( .A1(a_8_), .A2(n9259), .A3(b_31_), .ZN(n9258) );
  NAND2_X1 U9171 ( .A1(n8797), .A2(n8795), .ZN(n9259) );
  NOR2_X1 U9172 ( .A1(n8795), .A2(n8797), .ZN(n9256) );
  NOR2_X1 U9173 ( .A1(n9260), .A2(n9261), .ZN(n8797) );
  INV_X1 U9174 ( .A(n9262), .ZN(n9261) );
  NAND3_X1 U9175 ( .A1(a_9_), .A2(n9263), .A3(b_31_), .ZN(n9262) );
  NAND2_X1 U9176 ( .A1(n8785), .A2(n8783), .ZN(n9263) );
  NOR2_X1 U9177 ( .A1(n8783), .A2(n8785), .ZN(n9260) );
  NOR2_X1 U9178 ( .A1(n9264), .A2(n9265), .ZN(n8785) );
  NOR3_X1 U9179 ( .A1(n8769), .A2(n9266), .A3(n8448), .ZN(n9265) );
  INV_X1 U9180 ( .A(n9267), .ZN(n9266) );
  NAND2_X1 U9181 ( .A1(n8767), .A2(n8766), .ZN(n9267) );
  NOR2_X1 U9182 ( .A1(n8766), .A2(n8767), .ZN(n9264) );
  NOR2_X1 U9183 ( .A1(n9268), .A2(n9269), .ZN(n8767) );
  INV_X1 U9184 ( .A(n9270), .ZN(n9269) );
  NAND3_X1 U9185 ( .A1(a_11_), .A2(n9271), .A3(b_31_), .ZN(n9270) );
  NAND2_X1 U9186 ( .A1(n8755), .A2(n8753), .ZN(n9271) );
  NOR2_X1 U9187 ( .A1(n8753), .A2(n8755), .ZN(n9268) );
  NOR2_X1 U9188 ( .A1(n9272), .A2(n9273), .ZN(n8755) );
  NOR3_X1 U9189 ( .A1(n8739), .A2(n9274), .A3(n8448), .ZN(n9273) );
  NOR2_X1 U9190 ( .A1(n8737), .A2(n8736), .ZN(n9274) );
  INV_X1 U9191 ( .A(n9275), .ZN(n9272) );
  NAND2_X1 U9192 ( .A1(n8736), .A2(n8737), .ZN(n9275) );
  NAND2_X1 U9193 ( .A1(n9276), .A2(n9277), .ZN(n8737) );
  NAND3_X1 U9194 ( .A1(a_13_), .A2(n9278), .A3(b_31_), .ZN(n9277) );
  NAND2_X1 U9195 ( .A1(n8725), .A2(n8723), .ZN(n9278) );
  INV_X1 U9196 ( .A(n9279), .ZN(n9276) );
  NOR2_X1 U9197 ( .A1(n8723), .A2(n8725), .ZN(n9279) );
  NOR2_X1 U9198 ( .A1(n9280), .A2(n9281), .ZN(n8725) );
  INV_X1 U9199 ( .A(n9282), .ZN(n9281) );
  NAND3_X1 U9200 ( .A1(a_14_), .A2(n9283), .A3(b_31_), .ZN(n9282) );
  NAND2_X1 U9201 ( .A1(n8708), .A2(n8706), .ZN(n9283) );
  NOR2_X1 U9202 ( .A1(n8706), .A2(n8708), .ZN(n9280) );
  NOR2_X1 U9203 ( .A1(n9284), .A2(n9285), .ZN(n8708) );
  INV_X1 U9204 ( .A(n9286), .ZN(n9285) );
  NAND3_X1 U9205 ( .A1(a_15_), .A2(n9287), .A3(b_31_), .ZN(n9286) );
  NAND2_X1 U9206 ( .A1(n8696), .A2(n8694), .ZN(n9287) );
  NOR2_X1 U9207 ( .A1(n8694), .A2(n8696), .ZN(n9284) );
  NOR2_X1 U9208 ( .A1(n9288), .A2(n9289), .ZN(n8696) );
  NOR3_X1 U9209 ( .A1(n8680), .A2(n9290), .A3(n8448), .ZN(n9289) );
  INV_X1 U9210 ( .A(n9291), .ZN(n9290) );
  NAND2_X1 U9211 ( .A1(n8678), .A2(n8677), .ZN(n9291) );
  NOR2_X1 U9212 ( .A1(n8677), .A2(n8678), .ZN(n9288) );
  NOR2_X1 U9213 ( .A1(n9292), .A2(n9293), .ZN(n8678) );
  NOR3_X1 U9214 ( .A1(n8662), .A2(n9294), .A3(n8448), .ZN(n9293) );
  NOR2_X1 U9215 ( .A1(n8666), .A2(n8665), .ZN(n9294) );
  INV_X1 U9216 ( .A(n9295), .ZN(n9292) );
  NAND2_X1 U9217 ( .A1(n8665), .A2(n8666), .ZN(n9295) );
  NAND2_X1 U9218 ( .A1(n9296), .A2(n9297), .ZN(n8666) );
  NAND3_X1 U9219 ( .A1(a_18_), .A2(n9298), .A3(b_31_), .ZN(n9297) );
  INV_X1 U9220 ( .A(n9299), .ZN(n9298) );
  NOR2_X1 U9221 ( .A1(n8646), .A2(n8644), .ZN(n9299) );
  NAND2_X1 U9222 ( .A1(n8644), .A2(n8646), .ZN(n9296) );
  NAND2_X1 U9223 ( .A1(n8634), .A2(n9300), .ZN(n8646) );
  NAND2_X1 U9224 ( .A1(n8633), .A2(n8635), .ZN(n9300) );
  NAND2_X1 U9225 ( .A1(n9301), .A2(n9302), .ZN(n8635) );
  NAND2_X1 U9226 ( .A1(b_31_), .A2(a_19_), .ZN(n9301) );
  XNOR2_X1 U9227 ( .A(n9303), .B(n9304), .ZN(n8633) );
  NAND2_X1 U9228 ( .A1(n9305), .A2(n9306), .ZN(n9303) );
  INV_X1 U9229 ( .A(n9307), .ZN(n8634) );
  NOR2_X1 U9230 ( .A1(n9302), .A2(n8630), .ZN(n9307) );
  NAND2_X1 U9231 ( .A1(n9308), .A2(n9309), .ZN(n9302) );
  NAND2_X1 U9232 ( .A1(n9310), .A2(n8617), .ZN(n9309) );
  NAND2_X1 U9233 ( .A1(b_31_), .A2(a_20_), .ZN(n8617) );
  NAND2_X1 U9234 ( .A1(n8615), .A2(n8618), .ZN(n9310) );
  INV_X1 U9235 ( .A(n9311), .ZN(n9308) );
  NOR2_X1 U9236 ( .A1(n8618), .A2(n8615), .ZN(n9311) );
  XNOR2_X1 U9237 ( .A(n9312), .B(n9313), .ZN(n8615) );
  XOR2_X1 U9238 ( .A(n9314), .B(n9315), .Z(n9313) );
  NAND2_X1 U9239 ( .A1(b_30_), .A2(a_21_), .ZN(n9315) );
  NAND2_X1 U9240 ( .A1(n8605), .A2(n9316), .ZN(n8618) );
  NAND2_X1 U9241 ( .A1(n8604), .A2(n8606), .ZN(n9316) );
  NAND2_X1 U9242 ( .A1(n9317), .A2(n9318), .ZN(n8606) );
  NAND2_X1 U9243 ( .A1(b_31_), .A2(a_21_), .ZN(n9317) );
  XNOR2_X1 U9244 ( .A(n9319), .B(n9320), .ZN(n8604) );
  NAND2_X1 U9245 ( .A1(n9321), .A2(n9322), .ZN(n9319) );
  INV_X1 U9246 ( .A(n9323), .ZN(n8605) );
  NOR2_X1 U9247 ( .A1(n9318), .A2(n8601), .ZN(n9323) );
  NAND2_X1 U9248 ( .A1(n9324), .A2(n9325), .ZN(n9318) );
  NAND2_X1 U9249 ( .A1(n9326), .A2(n8589), .ZN(n9325) );
  NAND2_X1 U9250 ( .A1(b_31_), .A2(a_22_), .ZN(n8589) );
  NAND2_X1 U9251 ( .A1(n8587), .A2(n8588), .ZN(n9326) );
  INV_X1 U9252 ( .A(n9327), .ZN(n9324) );
  NOR2_X1 U9253 ( .A1(n8588), .A2(n8587), .ZN(n9327) );
  XNOR2_X1 U9254 ( .A(n9328), .B(n9329), .ZN(n8587) );
  NAND2_X1 U9255 ( .A1(n9330), .A2(n9331), .ZN(n9328) );
  NAND2_X1 U9256 ( .A1(n8576), .A2(n9332), .ZN(n8588) );
  NAND2_X1 U9257 ( .A1(n8575), .A2(n8577), .ZN(n9332) );
  NAND2_X1 U9258 ( .A1(n9333), .A2(n9334), .ZN(n8577) );
  INV_X1 U9259 ( .A(n9335), .ZN(n9334) );
  NAND2_X1 U9260 ( .A1(b_31_), .A2(a_23_), .ZN(n9333) );
  XNOR2_X1 U9261 ( .A(n9336), .B(n9337), .ZN(n8575) );
  XNOR2_X1 U9262 ( .A(n9338), .B(n9339), .ZN(n9336) );
  NAND2_X1 U9263 ( .A1(n9335), .A2(a_23_), .ZN(n8576) );
  NOR2_X1 U9264 ( .A1(n9340), .A2(n9341), .ZN(n9335) );
  NOR2_X1 U9265 ( .A1(n9342), .A2(n8559), .ZN(n9341) );
  NOR2_X1 U9266 ( .A1(n8448), .A2(n8982), .ZN(n8559) );
  INV_X1 U9267 ( .A(n9343), .ZN(n9342) );
  NAND2_X1 U9268 ( .A1(n8557), .A2(n8560), .ZN(n9343) );
  NOR2_X1 U9269 ( .A1(n8560), .A2(n8557), .ZN(n9340) );
  XOR2_X1 U9270 ( .A(n9344), .B(n9345), .Z(n8557) );
  XOR2_X1 U9271 ( .A(n9346), .B(n9347), .Z(n9344) );
  NAND2_X1 U9272 ( .A1(n9348), .A2(n9349), .ZN(n8560) );
  NAND2_X1 U9273 ( .A1(n8548), .A2(n9350), .ZN(n9349) );
  NAND2_X1 U9274 ( .A1(n8547), .A2(n8546), .ZN(n9350) );
  NOR2_X1 U9275 ( .A1(n8448), .A2(n8541), .ZN(n8548) );
  INV_X1 U9276 ( .A(n9351), .ZN(n9348) );
  NOR2_X1 U9277 ( .A1(n8546), .A2(n8547), .ZN(n9351) );
  NOR2_X1 U9278 ( .A1(n9352), .A2(n9353), .ZN(n8547) );
  NOR2_X1 U9279 ( .A1(n8530), .A2(n9354), .ZN(n9353) );
  NOR2_X1 U9280 ( .A1(n8531), .A2(n8528), .ZN(n9354) );
  NAND2_X1 U9281 ( .A1(b_31_), .A2(a_26_), .ZN(n8530) );
  INV_X1 U9282 ( .A(n9355), .ZN(n9352) );
  NAND2_X1 U9283 ( .A1(n8528), .A2(n8531), .ZN(n9355) );
  NAND2_X1 U9284 ( .A1(n9356), .A2(n9357), .ZN(n8531) );
  NAND2_X1 U9285 ( .A1(n8518), .A2(n9358), .ZN(n9357) );
  NAND2_X1 U9286 ( .A1(n8519), .A2(n8516), .ZN(n9358) );
  NOR2_X1 U9287 ( .A1(n8448), .A2(n8512), .ZN(n8518) );
  INV_X1 U9288 ( .A(n9359), .ZN(n9356) );
  NOR2_X1 U9289 ( .A1(n8516), .A2(n8519), .ZN(n9359) );
  NOR2_X1 U9290 ( .A1(n9360), .A2(n9361), .ZN(n8519) );
  INV_X1 U9291 ( .A(n9362), .ZN(n9361) );
  NAND3_X1 U9292 ( .A1(a_28_), .A2(n9363), .A3(b_31_), .ZN(n9362) );
  NAND2_X1 U9293 ( .A1(n8490), .A2(n8491), .ZN(n9363) );
  NOR2_X1 U9294 ( .A1(n8491), .A2(n8490), .ZN(n9360) );
  XNOR2_X1 U9295 ( .A(n9364), .B(n9365), .ZN(n8490) );
  XNOR2_X1 U9296 ( .A(n9366), .B(n9367), .ZN(n9364) );
  NAND2_X1 U9297 ( .A1(n9368), .A2(n9369), .ZN(n8491) );
  NAND2_X1 U9298 ( .A1(n9370), .A2(n8479), .ZN(n9369) );
  NAND2_X1 U9299 ( .A1(b_31_), .A2(a_29_), .ZN(n8479) );
  NAND2_X1 U9300 ( .A1(n8477), .A2(n8480), .ZN(n9370) );
  INV_X1 U9301 ( .A(n9371), .ZN(n9368) );
  NOR2_X1 U9302 ( .A1(n8480), .A2(n8477), .ZN(n9371) );
  NOR3_X1 U9303 ( .A1(n8461), .A2(n8979), .A3(n8448), .ZN(n8477) );
  INV_X1 U9304 ( .A(b_31_), .ZN(n8448) );
  NAND2_X1 U9305 ( .A1(n9372), .A2(n9373), .ZN(n8480) );
  NAND2_X1 U9306 ( .A1(b_29_), .A2(n9374), .ZN(n9373) );
  NAND2_X1 U9307 ( .A1(n8456), .A2(n9375), .ZN(n9374) );
  NAND2_X1 U9308 ( .A1(a_31_), .A2(n8461), .ZN(n9375) );
  NAND2_X1 U9309 ( .A1(b_30_), .A2(n9376), .ZN(n9372) );
  NAND2_X1 U9310 ( .A1(n8459), .A2(n9377), .ZN(n9376) );
  NAND2_X1 U9311 ( .A1(a_30_), .A2(n8475), .ZN(n9377) );
  XOR2_X1 U9312 ( .A(n9378), .B(n9379), .Z(n8516) );
  XNOR2_X1 U9313 ( .A(n9380), .B(n9381), .ZN(n9378) );
  XNOR2_X1 U9314 ( .A(n9382), .B(n9383), .ZN(n8528) );
  XNOR2_X1 U9315 ( .A(n9384), .B(n9385), .ZN(n9382) );
  NOR2_X1 U9316 ( .A1(n8512), .A2(n8461), .ZN(n9385) );
  XNOR2_X1 U9317 ( .A(n9386), .B(n9387), .ZN(n8546) );
  XNOR2_X1 U9318 ( .A(n9388), .B(n9389), .ZN(n9387) );
  XNOR2_X1 U9319 ( .A(n9390), .B(n9391), .ZN(n8644) );
  XOR2_X1 U9320 ( .A(n9392), .B(n9393), .Z(n9391) );
  NAND2_X1 U9321 ( .A1(b_30_), .A2(a_19_), .ZN(n9393) );
  XOR2_X1 U9322 ( .A(n9394), .B(n9395), .Z(n8665) );
  XNOR2_X1 U9323 ( .A(n9396), .B(n9397), .ZN(n9395) );
  XOR2_X1 U9324 ( .A(n9398), .B(n9399), .Z(n8677) );
  XOR2_X1 U9325 ( .A(n9400), .B(n9401), .Z(n9399) );
  NAND2_X1 U9326 ( .A1(b_30_), .A2(a_17_), .ZN(n9401) );
  XOR2_X1 U9327 ( .A(n9402), .B(n9403), .Z(n8694) );
  NAND2_X1 U9328 ( .A1(n9404), .A2(n9405), .ZN(n9402) );
  XNOR2_X1 U9329 ( .A(n9406), .B(n9407), .ZN(n8706) );
  XOR2_X1 U9330 ( .A(n9408), .B(n9409), .Z(n9406) );
  NOR2_X1 U9331 ( .A1(n8692), .A2(n8461), .ZN(n9409) );
  XOR2_X1 U9332 ( .A(n9410), .B(n9411), .Z(n8723) );
  NAND2_X1 U9333 ( .A1(n9412), .A2(n9413), .ZN(n9410) );
  XNOR2_X1 U9334 ( .A(n9414), .B(n9415), .ZN(n8736) );
  XOR2_X1 U9335 ( .A(n9416), .B(n9417), .Z(n9415) );
  NAND2_X1 U9336 ( .A1(b_30_), .A2(a_13_), .ZN(n9417) );
  XOR2_X1 U9337 ( .A(n9418), .B(n9419), .Z(n8753) );
  NAND2_X1 U9338 ( .A1(n9420), .A2(n9421), .ZN(n9418) );
  XNOR2_X1 U9339 ( .A(n9422), .B(n9423), .ZN(n8766) );
  XOR2_X1 U9340 ( .A(n9424), .B(n9425), .Z(n9422) );
  NOR2_X1 U9341 ( .A1(n8749), .A2(n8461), .ZN(n9425) );
  XOR2_X1 U9342 ( .A(n9426), .B(n9427), .Z(n8783) );
  NAND2_X1 U9343 ( .A1(n9428), .A2(n9429), .ZN(n9426) );
  XOR2_X1 U9344 ( .A(n9430), .B(n9431), .Z(n8795) );
  XOR2_X1 U9345 ( .A(n9432), .B(n9433), .Z(n9431) );
  NAND2_X1 U9346 ( .A1(b_30_), .A2(a_9_), .ZN(n9433) );
  XOR2_X1 U9347 ( .A(n9434), .B(n9435), .Z(n8821) );
  NAND2_X1 U9348 ( .A1(n9436), .A2(n9437), .ZN(n9434) );
  XNOR2_X1 U9349 ( .A(n9438), .B(n9439), .ZN(n8833) );
  XOR2_X1 U9350 ( .A(n9440), .B(n9441), .Z(n9438) );
  NOR2_X1 U9351 ( .A1(n8817), .A2(n8461), .ZN(n9441) );
  XOR2_X1 U9352 ( .A(n9442), .B(n9443), .Z(n8850) );
  NAND2_X1 U9353 ( .A1(n9444), .A2(n9445), .ZN(n9442) );
  XOR2_X1 U9354 ( .A(n9446), .B(n9447), .Z(n8862) );
  XOR2_X1 U9355 ( .A(n9448), .B(n9449), .Z(n9447) );
  NAND2_X1 U9356 ( .A1(b_30_), .A2(a_5_), .ZN(n9449) );
  XOR2_X1 U9357 ( .A(n9450), .B(n9451), .Z(n8880) );
  NAND2_X1 U9358 ( .A1(n9452), .A2(n9453), .ZN(n9450) );
  XOR2_X1 U9359 ( .A(n9454), .B(n9455), .Z(n8891) );
  NAND2_X1 U9360 ( .A1(n9456), .A2(n9457), .ZN(n9454) );
  XOR2_X1 U9361 ( .A(n9458), .B(n9459), .Z(n8909) );
  XOR2_X1 U9362 ( .A(n9460), .B(n9461), .Z(n9458) );
  XOR2_X1 U9363 ( .A(n9462), .B(n9463), .Z(n9000) );
  XNOR2_X1 U9364 ( .A(n9464), .B(n9465), .ZN(n9463) );
  NAND2_X1 U9365 ( .A1(b_30_), .A2(a_1_), .ZN(n9465) );
  XNOR2_X1 U9366 ( .A(n9011), .B(n9012), .ZN(n9219) );
  NAND3_X1 U9367 ( .A1(n9012), .A2(n9011), .A3(n9466), .ZN(n9019) );
  XNOR2_X1 U9368 ( .A(n9467), .B(n9215), .ZN(n9466) );
  INV_X1 U9369 ( .A(n9214), .ZN(n9467) );
  NAND2_X1 U9370 ( .A1(n9468), .A2(n9469), .ZN(n9011) );
  INV_X1 U9371 ( .A(n9470), .ZN(n9469) );
  NOR3_X1 U9372 ( .A1(n9471), .A2(n9472), .A3(n8461), .ZN(n9470) );
  NOR2_X1 U9373 ( .A1(n9222), .A2(n9220), .ZN(n9472) );
  NAND2_X1 U9374 ( .A1(n9220), .A2(n9222), .ZN(n9468) );
  NAND2_X1 U9375 ( .A1(n9473), .A2(n9474), .ZN(n9222) );
  NAND3_X1 U9376 ( .A1(a_1_), .A2(n9475), .A3(b_30_), .ZN(n9474) );
  NAND2_X1 U9377 ( .A1(n9462), .A2(n9476), .ZN(n9475) );
  INV_X1 U9378 ( .A(n9464), .ZN(n9476) );
  NAND2_X1 U9379 ( .A1(n9464), .A2(n9477), .ZN(n9473) );
  INV_X1 U9380 ( .A(n9462), .ZN(n9477) );
  XOR2_X1 U9381 ( .A(n9478), .B(n9479), .Z(n9462) );
  XNOR2_X1 U9382 ( .A(n9480), .B(n9481), .ZN(n9479) );
  NOR2_X1 U9383 ( .A1(n9482), .A2(n9483), .ZN(n9464) );
  INV_X1 U9384 ( .A(n9484), .ZN(n9483) );
  NAND2_X1 U9385 ( .A1(n9459), .A2(n9485), .ZN(n9484) );
  NAND2_X1 U9386 ( .A1(n9461), .A2(n9460), .ZN(n9485) );
  XOR2_X1 U9387 ( .A(n9486), .B(n9487), .Z(n9459) );
  NAND2_X1 U9388 ( .A1(n9488), .A2(n9489), .ZN(n9486) );
  NOR2_X1 U9389 ( .A1(n9460), .A2(n9461), .ZN(n9482) );
  NOR2_X1 U9390 ( .A1(n8461), .A2(n8998), .ZN(n9461) );
  NAND2_X1 U9391 ( .A1(n9456), .A2(n9490), .ZN(n9460) );
  NAND2_X1 U9392 ( .A1(n9455), .A2(n9457), .ZN(n9490) );
  NAND2_X1 U9393 ( .A1(n9491), .A2(n9492), .ZN(n9457) );
  NAND2_X1 U9394 ( .A1(b_30_), .A2(a_3_), .ZN(n9492) );
  INV_X1 U9395 ( .A(n9493), .ZN(n9491) );
  XNOR2_X1 U9396 ( .A(n9494), .B(n9495), .ZN(n9455) );
  NAND2_X1 U9397 ( .A1(n9496), .A2(n9497), .ZN(n9494) );
  NAND2_X1 U9398 ( .A1(a_3_), .A2(n9493), .ZN(n9456) );
  NAND2_X1 U9399 ( .A1(n9452), .A2(n9498), .ZN(n9493) );
  NAND2_X1 U9400 ( .A1(n9451), .A2(n9453), .ZN(n9498) );
  NAND2_X1 U9401 ( .A1(n9499), .A2(n9500), .ZN(n9453) );
  NAND2_X1 U9402 ( .A1(b_30_), .A2(a_4_), .ZN(n9500) );
  INV_X1 U9403 ( .A(n9501), .ZN(n9499) );
  XOR2_X1 U9404 ( .A(n9502), .B(n9503), .Z(n9451) );
  XOR2_X1 U9405 ( .A(n9504), .B(n9505), .Z(n9502) );
  NOR2_X1 U9406 ( .A1(n8848), .A2(n8475), .ZN(n9505) );
  NAND2_X1 U9407 ( .A1(a_4_), .A2(n9501), .ZN(n9452) );
  NAND2_X1 U9408 ( .A1(n9506), .A2(n9507), .ZN(n9501) );
  INV_X1 U9409 ( .A(n9508), .ZN(n9507) );
  NOR3_X1 U9410 ( .A1(n8848), .A2(n9509), .A3(n8461), .ZN(n9508) );
  NOR2_X1 U9411 ( .A1(n9448), .A2(n9446), .ZN(n9509) );
  NAND2_X1 U9412 ( .A1(n9446), .A2(n9448), .ZN(n9506) );
  NAND2_X1 U9413 ( .A1(n9444), .A2(n9510), .ZN(n9448) );
  NAND2_X1 U9414 ( .A1(n9443), .A2(n9445), .ZN(n9510) );
  NAND2_X1 U9415 ( .A1(n9511), .A2(n9512), .ZN(n9445) );
  NAND2_X1 U9416 ( .A1(b_30_), .A2(a_6_), .ZN(n9512) );
  INV_X1 U9417 ( .A(n9513), .ZN(n9511) );
  XOR2_X1 U9418 ( .A(n9514), .B(n9515), .Z(n9443) );
  XOR2_X1 U9419 ( .A(n9516), .B(n9517), .Z(n9514) );
  NOR2_X1 U9420 ( .A1(n8817), .A2(n8475), .ZN(n9517) );
  NAND2_X1 U9421 ( .A1(a_6_), .A2(n9513), .ZN(n9444) );
  NAND2_X1 U9422 ( .A1(n9518), .A2(n9519), .ZN(n9513) );
  INV_X1 U9423 ( .A(n9520), .ZN(n9519) );
  NOR3_X1 U9424 ( .A1(n8817), .A2(n9521), .A3(n8461), .ZN(n9520) );
  NOR2_X1 U9425 ( .A1(n9440), .A2(n9439), .ZN(n9521) );
  NAND2_X1 U9426 ( .A1(n9439), .A2(n9440), .ZN(n9518) );
  NAND2_X1 U9427 ( .A1(n9436), .A2(n9522), .ZN(n9440) );
  NAND2_X1 U9428 ( .A1(n9435), .A2(n9437), .ZN(n9522) );
  NAND2_X1 U9429 ( .A1(n9523), .A2(n9524), .ZN(n9437) );
  NAND2_X1 U9430 ( .A1(b_30_), .A2(a_8_), .ZN(n9524) );
  INV_X1 U9431 ( .A(n9525), .ZN(n9523) );
  XNOR2_X1 U9432 ( .A(n9526), .B(n9527), .ZN(n9435) );
  XOR2_X1 U9433 ( .A(n9528), .B(n9529), .Z(n9527) );
  NAND2_X1 U9434 ( .A1(b_29_), .A2(a_9_), .ZN(n9529) );
  NAND2_X1 U9435 ( .A1(a_8_), .A2(n9525), .ZN(n9436) );
  NAND2_X1 U9436 ( .A1(n9530), .A2(n9531), .ZN(n9525) );
  INV_X1 U9437 ( .A(n9532), .ZN(n9531) );
  NOR3_X1 U9438 ( .A1(n8779), .A2(n9533), .A3(n8461), .ZN(n9532) );
  NOR2_X1 U9439 ( .A1(n9432), .A2(n9430), .ZN(n9533) );
  NAND2_X1 U9440 ( .A1(n9430), .A2(n9432), .ZN(n9530) );
  NAND2_X1 U9441 ( .A1(n9428), .A2(n9534), .ZN(n9432) );
  NAND2_X1 U9442 ( .A1(n9427), .A2(n9429), .ZN(n9534) );
  NAND2_X1 U9443 ( .A1(n9535), .A2(n9536), .ZN(n9429) );
  NAND2_X1 U9444 ( .A1(b_30_), .A2(a_10_), .ZN(n9536) );
  XOR2_X1 U9445 ( .A(n9537), .B(n9538), .Z(n9427) );
  XOR2_X1 U9446 ( .A(n9539), .B(n9540), .Z(n9537) );
  NOR2_X1 U9447 ( .A1(n8749), .A2(n8475), .ZN(n9540) );
  INV_X1 U9448 ( .A(n9541), .ZN(n9428) );
  NOR2_X1 U9449 ( .A1(n8769), .A2(n9535), .ZN(n9541) );
  NOR2_X1 U9450 ( .A1(n9542), .A2(n9543), .ZN(n9535) );
  NOR3_X1 U9451 ( .A1(n8749), .A2(n9544), .A3(n8461), .ZN(n9543) );
  NOR2_X1 U9452 ( .A1(n9424), .A2(n9423), .ZN(n9544) );
  INV_X1 U9453 ( .A(n9545), .ZN(n9542) );
  NAND2_X1 U9454 ( .A1(n9423), .A2(n9424), .ZN(n9545) );
  NAND2_X1 U9455 ( .A1(n9420), .A2(n9546), .ZN(n9424) );
  NAND2_X1 U9456 ( .A1(n9419), .A2(n9421), .ZN(n9546) );
  NAND2_X1 U9457 ( .A1(n9547), .A2(n9548), .ZN(n9421) );
  NAND2_X1 U9458 ( .A1(b_30_), .A2(a_12_), .ZN(n9548) );
  XNOR2_X1 U9459 ( .A(n9549), .B(n9550), .ZN(n9419) );
  XOR2_X1 U9460 ( .A(n9551), .B(n9552), .Z(n9550) );
  NAND2_X1 U9461 ( .A1(b_29_), .A2(a_13_), .ZN(n9552) );
  INV_X1 U9462 ( .A(n9553), .ZN(n9420) );
  NOR2_X1 U9463 ( .A1(n8739), .A2(n9547), .ZN(n9553) );
  NOR2_X1 U9464 ( .A1(n9554), .A2(n9555), .ZN(n9547) );
  NOR3_X1 U9465 ( .A1(n8721), .A2(n9556), .A3(n8461), .ZN(n9555) );
  NOR2_X1 U9466 ( .A1(n9416), .A2(n9414), .ZN(n9556) );
  INV_X1 U9467 ( .A(n9557), .ZN(n9554) );
  NAND2_X1 U9468 ( .A1(n9414), .A2(n9416), .ZN(n9557) );
  NAND2_X1 U9469 ( .A1(n9412), .A2(n9558), .ZN(n9416) );
  NAND2_X1 U9470 ( .A1(n9411), .A2(n9413), .ZN(n9558) );
  NAND2_X1 U9471 ( .A1(n9559), .A2(n9560), .ZN(n9413) );
  NAND2_X1 U9472 ( .A1(b_30_), .A2(a_14_), .ZN(n9560) );
  INV_X1 U9473 ( .A(n9561), .ZN(n9559) );
  XOR2_X1 U9474 ( .A(n9562), .B(n9563), .Z(n9411) );
  XOR2_X1 U9475 ( .A(n9564), .B(n9565), .Z(n9562) );
  NOR2_X1 U9476 ( .A1(n8692), .A2(n8475), .ZN(n9565) );
  NAND2_X1 U9477 ( .A1(a_14_), .A2(n9561), .ZN(n9412) );
  NAND2_X1 U9478 ( .A1(n9566), .A2(n9567), .ZN(n9561) );
  INV_X1 U9479 ( .A(n9568), .ZN(n9567) );
  NOR3_X1 U9480 ( .A1(n8692), .A2(n9569), .A3(n8461), .ZN(n9568) );
  NOR2_X1 U9481 ( .A1(n9408), .A2(n9407), .ZN(n9569) );
  NAND2_X1 U9482 ( .A1(n9407), .A2(n9408), .ZN(n9566) );
  NAND2_X1 U9483 ( .A1(n9404), .A2(n9570), .ZN(n9408) );
  NAND2_X1 U9484 ( .A1(n9403), .A2(n9405), .ZN(n9570) );
  NAND2_X1 U9485 ( .A1(n9571), .A2(n9572), .ZN(n9405) );
  NAND2_X1 U9486 ( .A1(b_30_), .A2(a_16_), .ZN(n9572) );
  XNOR2_X1 U9487 ( .A(n9573), .B(n9574), .ZN(n9403) );
  XOR2_X1 U9488 ( .A(n9575), .B(n9576), .Z(n9574) );
  NAND2_X1 U9489 ( .A1(b_29_), .A2(a_17_), .ZN(n9576) );
  NAND2_X1 U9490 ( .A1(a_16_), .A2(n9577), .ZN(n9404) );
  INV_X1 U9491 ( .A(n9571), .ZN(n9577) );
  NOR2_X1 U9492 ( .A1(n9578), .A2(n9579), .ZN(n9571) );
  NOR3_X1 U9493 ( .A1(n8662), .A2(n9580), .A3(n8461), .ZN(n9579) );
  INV_X1 U9494 ( .A(n9581), .ZN(n9580) );
  NAND2_X1 U9495 ( .A1(n9398), .A2(n9400), .ZN(n9581) );
  NOR2_X1 U9496 ( .A1(n9400), .A2(n9398), .ZN(n9578) );
  XOR2_X1 U9497 ( .A(n9582), .B(n9583), .Z(n9398) );
  XOR2_X1 U9498 ( .A(n9584), .B(n9585), .Z(n9582) );
  NAND2_X1 U9499 ( .A1(n9586), .A2(n9587), .ZN(n9400) );
  NAND2_X1 U9500 ( .A1(n9394), .A2(n9588), .ZN(n9587) );
  INV_X1 U9501 ( .A(n9589), .ZN(n9588) );
  NOR2_X1 U9502 ( .A1(n9397), .A2(n9396), .ZN(n9589) );
  XNOR2_X1 U9503 ( .A(n9590), .B(n9591), .ZN(n9394) );
  XOR2_X1 U9504 ( .A(n9592), .B(n9593), .Z(n9590) );
  NOR2_X1 U9505 ( .A1(n8630), .A2(n8475), .ZN(n9593) );
  NAND2_X1 U9506 ( .A1(n9396), .A2(n9397), .ZN(n9586) );
  NAND2_X1 U9507 ( .A1(b_30_), .A2(a_18_), .ZN(n9397) );
  NOR2_X1 U9508 ( .A1(n9594), .A2(n9595), .ZN(n9396) );
  NOR3_X1 U9509 ( .A1(n8630), .A2(n9596), .A3(n8461), .ZN(n9595) );
  NOR2_X1 U9510 ( .A1(n9392), .A2(n9390), .ZN(n9596) );
  INV_X1 U9511 ( .A(n9597), .ZN(n9594) );
  NAND2_X1 U9512 ( .A1(n9390), .A2(n9392), .ZN(n9597) );
  NAND2_X1 U9513 ( .A1(n9305), .A2(n9598), .ZN(n9392) );
  NAND2_X1 U9514 ( .A1(n9304), .A2(n9306), .ZN(n9598) );
  NAND2_X1 U9515 ( .A1(n9599), .A2(n9600), .ZN(n9306) );
  NAND2_X1 U9516 ( .A1(b_30_), .A2(a_20_), .ZN(n9600) );
  XOR2_X1 U9517 ( .A(n9601), .B(n9602), .Z(n9304) );
  XOR2_X1 U9518 ( .A(n9603), .B(n9604), .Z(n9601) );
  NOR2_X1 U9519 ( .A1(n8601), .A2(n8475), .ZN(n9604) );
  INV_X1 U9520 ( .A(n9605), .ZN(n9305) );
  NOR2_X1 U9521 ( .A1(n8986), .A2(n9599), .ZN(n9605) );
  NOR2_X1 U9522 ( .A1(n9606), .A2(n9607), .ZN(n9599) );
  NOR3_X1 U9523 ( .A1(n8601), .A2(n9608), .A3(n8461), .ZN(n9607) );
  NOR2_X1 U9524 ( .A1(n9314), .A2(n9312), .ZN(n9608) );
  INV_X1 U9525 ( .A(n9609), .ZN(n9606) );
  NAND2_X1 U9526 ( .A1(n9312), .A2(n9314), .ZN(n9609) );
  NAND2_X1 U9527 ( .A1(n9321), .A2(n9610), .ZN(n9314) );
  NAND2_X1 U9528 ( .A1(n9320), .A2(n9322), .ZN(n9610) );
  NAND2_X1 U9529 ( .A1(n9611), .A2(n9612), .ZN(n9322) );
  NAND2_X1 U9530 ( .A1(b_30_), .A2(a_22_), .ZN(n9612) );
  INV_X1 U9531 ( .A(n9613), .ZN(n9611) );
  XNOR2_X1 U9532 ( .A(n9614), .B(n9615), .ZN(n9320) );
  NAND2_X1 U9533 ( .A1(n9616), .A2(n9617), .ZN(n9614) );
  NAND2_X1 U9534 ( .A1(a_22_), .A2(n9613), .ZN(n9321) );
  NAND2_X1 U9535 ( .A1(n9330), .A2(n9618), .ZN(n9613) );
  NAND2_X1 U9536 ( .A1(n9329), .A2(n9331), .ZN(n9618) );
  NAND2_X1 U9537 ( .A1(n9619), .A2(n9620), .ZN(n9331) );
  NAND2_X1 U9538 ( .A1(b_30_), .A2(a_23_), .ZN(n9620) );
  INV_X1 U9539 ( .A(n9621), .ZN(n9619) );
  XNOR2_X1 U9540 ( .A(n9622), .B(n9623), .ZN(n9329) );
  XNOR2_X1 U9541 ( .A(n9624), .B(n9625), .ZN(n9622) );
  NAND2_X1 U9542 ( .A1(a_23_), .A2(n9621), .ZN(n9330) );
  NAND2_X1 U9543 ( .A1(n9626), .A2(n9627), .ZN(n9621) );
  NAND2_X1 U9544 ( .A1(n9339), .A2(n9628), .ZN(n9627) );
  NAND2_X1 U9545 ( .A1(n9338), .A2(n9337), .ZN(n9628) );
  NOR2_X1 U9546 ( .A1(n8461), .A2(n8982), .ZN(n9339) );
  NAND2_X1 U9547 ( .A1(n9629), .A2(n9630), .ZN(n9626) );
  INV_X1 U9548 ( .A(n9338), .ZN(n9630) );
  NOR2_X1 U9549 ( .A1(n9631), .A2(n9632), .ZN(n9338) );
  INV_X1 U9550 ( .A(n9633), .ZN(n9632) );
  NAND2_X1 U9551 ( .A1(n9347), .A2(n9634), .ZN(n9633) );
  NAND2_X1 U9552 ( .A1(n9345), .A2(n9346), .ZN(n9634) );
  NOR2_X1 U9553 ( .A1(n8461), .A2(n8541), .ZN(n9347) );
  NOR2_X1 U9554 ( .A1(n9346), .A2(n9345), .ZN(n9631) );
  XNOR2_X1 U9555 ( .A(n9635), .B(n9636), .ZN(n9345) );
  XNOR2_X1 U9556 ( .A(n9637), .B(n9638), .ZN(n9636) );
  NAND2_X1 U9557 ( .A1(n9639), .A2(n9640), .ZN(n9346) );
  NAND2_X1 U9558 ( .A1(n9386), .A2(n9641), .ZN(n9640) );
  INV_X1 U9559 ( .A(n9642), .ZN(n9641) );
  NOR2_X1 U9560 ( .A1(n9389), .A2(n9388), .ZN(n9642) );
  XOR2_X1 U9561 ( .A(n9643), .B(n9644), .Z(n9386) );
  XNOR2_X1 U9562 ( .A(n9645), .B(n9646), .ZN(n9644) );
  NAND2_X1 U9563 ( .A1(b_29_), .A2(a_27_), .ZN(n9646) );
  NAND2_X1 U9564 ( .A1(n9388), .A2(n9389), .ZN(n9639) );
  NAND2_X1 U9565 ( .A1(b_30_), .A2(a_26_), .ZN(n9389) );
  NOR2_X1 U9566 ( .A1(n9647), .A2(n9648), .ZN(n9388) );
  INV_X1 U9567 ( .A(n9649), .ZN(n9648) );
  NAND3_X1 U9568 ( .A1(a_27_), .A2(n9650), .A3(b_30_), .ZN(n9649) );
  NAND2_X1 U9569 ( .A1(n9384), .A2(n9383), .ZN(n9650) );
  NOR2_X1 U9570 ( .A1(n9383), .A2(n9384), .ZN(n9647) );
  NOR2_X1 U9571 ( .A1(n9651), .A2(n9652), .ZN(n9384) );
  INV_X1 U9572 ( .A(n9653), .ZN(n9652) );
  NAND2_X1 U9573 ( .A1(n9380), .A2(n9654), .ZN(n9653) );
  NAND2_X1 U9574 ( .A1(n9381), .A2(n9379), .ZN(n9654) );
  NOR2_X1 U9575 ( .A1(n8461), .A2(n8493), .ZN(n9380) );
  NOR2_X1 U9576 ( .A1(n9379), .A2(n9381), .ZN(n9651) );
  NOR2_X1 U9577 ( .A1(n9655), .A2(n9656), .ZN(n9381) );
  INV_X1 U9578 ( .A(n9657), .ZN(n9656) );
  NAND2_X1 U9579 ( .A1(n9365), .A2(n9658), .ZN(n9657) );
  NAND2_X1 U9580 ( .A1(n9659), .A2(n9367), .ZN(n9658) );
  NOR2_X1 U9581 ( .A1(n8461), .A2(n8473), .ZN(n9365) );
  INV_X1 U9582 ( .A(b_30_), .ZN(n8461) );
  NOR2_X1 U9583 ( .A1(n9367), .A2(n9659), .ZN(n9655) );
  INV_X1 U9584 ( .A(n9366), .ZN(n9659) );
  NAND2_X1 U9585 ( .A1(n9660), .A2(n9661), .ZN(n9366) );
  NAND2_X1 U9586 ( .A1(b_28_), .A2(n9662), .ZN(n9661) );
  NAND2_X1 U9587 ( .A1(n8456), .A2(n9663), .ZN(n9662) );
  NAND2_X1 U9588 ( .A1(a_31_), .A2(n8475), .ZN(n9663) );
  NAND2_X1 U9589 ( .A1(b_29_), .A2(n9664), .ZN(n9660) );
  NAND2_X1 U9590 ( .A1(n8459), .A2(n9665), .ZN(n9664) );
  NAND2_X1 U9591 ( .A1(a_30_), .A2(n8980), .ZN(n9665) );
  NAND3_X1 U9592 ( .A1(b_29_), .A2(n9666), .A3(b_30_), .ZN(n9367) );
  XOR2_X1 U9593 ( .A(n9667), .B(n8972), .Z(n9379) );
  INV_X1 U9594 ( .A(n8470), .ZN(n8972) );
  XNOR2_X1 U9595 ( .A(n9668), .B(n9669), .ZN(n9667) );
  XNOR2_X1 U9596 ( .A(n9670), .B(n9671), .ZN(n9383) );
  XOR2_X1 U9597 ( .A(n9672), .B(n9673), .Z(n9670) );
  INV_X1 U9598 ( .A(n9337), .ZN(n9629) );
  XOR2_X1 U9599 ( .A(n9674), .B(n9675), .Z(n9337) );
  XNOR2_X1 U9600 ( .A(n9676), .B(n9677), .ZN(n9675) );
  XNOR2_X1 U9601 ( .A(n9678), .B(n9679), .ZN(n9312) );
  NAND2_X1 U9602 ( .A1(n9680), .A2(n9681), .ZN(n9678) );
  XNOR2_X1 U9603 ( .A(n9682), .B(n9683), .ZN(n9390) );
  NAND2_X1 U9604 ( .A1(n9684), .A2(n9685), .ZN(n9682) );
  XNOR2_X1 U9605 ( .A(n9686), .B(n9687), .ZN(n9407) );
  NAND2_X1 U9606 ( .A1(n9688), .A2(n9689), .ZN(n9686) );
  XNOR2_X1 U9607 ( .A(n9690), .B(n9691), .ZN(n9414) );
  NAND2_X1 U9608 ( .A1(n9692), .A2(n9693), .ZN(n9690) );
  XNOR2_X1 U9609 ( .A(n9694), .B(n9695), .ZN(n9423) );
  NAND2_X1 U9610 ( .A1(n9696), .A2(n9697), .ZN(n9694) );
  XNOR2_X1 U9611 ( .A(n9698), .B(n9699), .ZN(n9430) );
  NAND2_X1 U9612 ( .A1(n9700), .A2(n9701), .ZN(n9698) );
  XNOR2_X1 U9613 ( .A(n9702), .B(n9703), .ZN(n9439) );
  NAND2_X1 U9614 ( .A1(n9704), .A2(n9705), .ZN(n9702) );
  XNOR2_X1 U9615 ( .A(n9706), .B(n9707), .ZN(n9446) );
  NAND2_X1 U9616 ( .A1(n9708), .A2(n9709), .ZN(n9706) );
  XOR2_X1 U9617 ( .A(n9710), .B(n9711), .Z(n9220) );
  XOR2_X1 U9618 ( .A(n9712), .B(n9713), .Z(n9710) );
  XNOR2_X1 U9619 ( .A(n9714), .B(n9715), .ZN(n9012) );
  NAND2_X1 U9620 ( .A1(n9716), .A2(n9717), .ZN(n9714) );
  NAND3_X1 U9621 ( .A1(n9214), .A2(n9215), .A3(n9718), .ZN(n9023) );
  XOR2_X1 U9622 ( .A(n9209), .B(n9210), .Z(n9718) );
  NAND2_X1 U9623 ( .A1(n9716), .A2(n9719), .ZN(n9215) );
  NAND2_X1 U9624 ( .A1(n9715), .A2(n9717), .ZN(n9719) );
  NAND2_X1 U9625 ( .A1(n9720), .A2(n9721), .ZN(n9717) );
  NAND2_X1 U9626 ( .A1(b_29_), .A2(a_0_), .ZN(n9721) );
  INV_X1 U9627 ( .A(n9722), .ZN(n9720) );
  XOR2_X1 U9628 ( .A(n9723), .B(n9724), .Z(n9715) );
  XOR2_X1 U9629 ( .A(n9725), .B(n9726), .Z(n9723) );
  NAND2_X1 U9630 ( .A1(a_0_), .A2(n9722), .ZN(n9716) );
  NAND2_X1 U9631 ( .A1(n9727), .A2(n9728), .ZN(n9722) );
  NAND2_X1 U9632 ( .A1(n9713), .A2(n9729), .ZN(n9728) );
  INV_X1 U9633 ( .A(n9730), .ZN(n9729) );
  NOR2_X1 U9634 ( .A1(n9712), .A2(n9711), .ZN(n9730) );
  NOR2_X1 U9635 ( .A1(n8475), .A2(n9731), .ZN(n9713) );
  NAND2_X1 U9636 ( .A1(n9711), .A2(n9712), .ZN(n9727) );
  NAND2_X1 U9637 ( .A1(n9732), .A2(n9733), .ZN(n9712) );
  NAND2_X1 U9638 ( .A1(n9480), .A2(n9734), .ZN(n9733) );
  NAND2_X1 U9639 ( .A1(n9735), .A2(n9736), .ZN(n9734) );
  INV_X1 U9640 ( .A(n9481), .ZN(n9736) );
  INV_X1 U9641 ( .A(n9478), .ZN(n9735) );
  NAND2_X1 U9642 ( .A1(n9488), .A2(n9737), .ZN(n9480) );
  NAND2_X1 U9643 ( .A1(n9487), .A2(n9489), .ZN(n9737) );
  NAND2_X1 U9644 ( .A1(n9738), .A2(n9739), .ZN(n9489) );
  NAND2_X1 U9645 ( .A1(b_29_), .A2(a_3_), .ZN(n9739) );
  INV_X1 U9646 ( .A(n9740), .ZN(n9738) );
  XNOR2_X1 U9647 ( .A(n9741), .B(n9742), .ZN(n9487) );
  XOR2_X1 U9648 ( .A(n9743), .B(n9744), .Z(n9742) );
  NAND2_X1 U9649 ( .A1(b_28_), .A2(a_4_), .ZN(n9744) );
  NAND2_X1 U9650 ( .A1(a_3_), .A2(n9740), .ZN(n9488) );
  NAND2_X1 U9651 ( .A1(n9496), .A2(n9745), .ZN(n9740) );
  NAND2_X1 U9652 ( .A1(n9495), .A2(n9497), .ZN(n9745) );
  NAND2_X1 U9653 ( .A1(n9746), .A2(n9747), .ZN(n9497) );
  NAND2_X1 U9654 ( .A1(b_29_), .A2(a_4_), .ZN(n9747) );
  XOR2_X1 U9655 ( .A(n9748), .B(n9749), .Z(n9495) );
  XOR2_X1 U9656 ( .A(n9750), .B(n9751), .Z(n9748) );
  NOR2_X1 U9657 ( .A1(n8848), .A2(n8980), .ZN(n9751) );
  INV_X1 U9658 ( .A(n9752), .ZN(n9496) );
  NOR2_X1 U9659 ( .A1(n8996), .A2(n9746), .ZN(n9752) );
  NOR2_X1 U9660 ( .A1(n9753), .A2(n9754), .ZN(n9746) );
  NOR3_X1 U9661 ( .A1(n8848), .A2(n9755), .A3(n8475), .ZN(n9754) );
  NOR2_X1 U9662 ( .A1(n9504), .A2(n9503), .ZN(n9755) );
  INV_X1 U9663 ( .A(n9756), .ZN(n9753) );
  NAND2_X1 U9664 ( .A1(n9503), .A2(n9504), .ZN(n9756) );
  NAND2_X1 U9665 ( .A1(n9708), .A2(n9757), .ZN(n9504) );
  NAND2_X1 U9666 ( .A1(n9707), .A2(n9709), .ZN(n9757) );
  NAND2_X1 U9667 ( .A1(n9758), .A2(n9759), .ZN(n9709) );
  NAND2_X1 U9668 ( .A1(b_29_), .A2(a_6_), .ZN(n9759) );
  XNOR2_X1 U9669 ( .A(n9760), .B(n9761), .ZN(n9707) );
  XOR2_X1 U9670 ( .A(n9762), .B(n9763), .Z(n9761) );
  NAND2_X1 U9671 ( .A1(b_28_), .A2(a_7_), .ZN(n9763) );
  INV_X1 U9672 ( .A(n9764), .ZN(n9708) );
  NOR2_X1 U9673 ( .A1(n8994), .A2(n9758), .ZN(n9764) );
  NOR2_X1 U9674 ( .A1(n9765), .A2(n9766), .ZN(n9758) );
  NOR3_X1 U9675 ( .A1(n8817), .A2(n9767), .A3(n8475), .ZN(n9766) );
  NOR2_X1 U9676 ( .A1(n9516), .A2(n9515), .ZN(n9767) );
  INV_X1 U9677 ( .A(n9768), .ZN(n9765) );
  NAND2_X1 U9678 ( .A1(n9515), .A2(n9516), .ZN(n9768) );
  NAND2_X1 U9679 ( .A1(n9704), .A2(n9769), .ZN(n9516) );
  NAND2_X1 U9680 ( .A1(n9703), .A2(n9705), .ZN(n9769) );
  NAND2_X1 U9681 ( .A1(n9770), .A2(n9771), .ZN(n9705) );
  NAND2_X1 U9682 ( .A1(b_29_), .A2(a_8_), .ZN(n9771) );
  INV_X1 U9683 ( .A(n9772), .ZN(n9770) );
  XNOR2_X1 U9684 ( .A(n9773), .B(n9774), .ZN(n9703) );
  XOR2_X1 U9685 ( .A(n9775), .B(n9776), .Z(n9774) );
  NAND2_X1 U9686 ( .A1(b_28_), .A2(a_9_), .ZN(n9776) );
  NAND2_X1 U9687 ( .A1(a_8_), .A2(n9772), .ZN(n9704) );
  NAND2_X1 U9688 ( .A1(n9777), .A2(n9778), .ZN(n9772) );
  INV_X1 U9689 ( .A(n9779), .ZN(n9778) );
  NOR3_X1 U9690 ( .A1(n8779), .A2(n9780), .A3(n8475), .ZN(n9779) );
  NOR2_X1 U9691 ( .A1(n9528), .A2(n9526), .ZN(n9780) );
  NAND2_X1 U9692 ( .A1(n9526), .A2(n9528), .ZN(n9777) );
  NAND2_X1 U9693 ( .A1(n9700), .A2(n9781), .ZN(n9528) );
  NAND2_X1 U9694 ( .A1(n9699), .A2(n9701), .ZN(n9781) );
  NAND2_X1 U9695 ( .A1(n9782), .A2(n9783), .ZN(n9701) );
  NAND2_X1 U9696 ( .A1(b_29_), .A2(a_10_), .ZN(n9783) );
  INV_X1 U9697 ( .A(n9784), .ZN(n9782) );
  XOR2_X1 U9698 ( .A(n9785), .B(n9786), .Z(n9699) );
  XOR2_X1 U9699 ( .A(n9787), .B(n9788), .Z(n9785) );
  NOR2_X1 U9700 ( .A1(n8749), .A2(n8980), .ZN(n9788) );
  NAND2_X1 U9701 ( .A1(a_10_), .A2(n9784), .ZN(n9700) );
  NAND2_X1 U9702 ( .A1(n9789), .A2(n9790), .ZN(n9784) );
  INV_X1 U9703 ( .A(n9791), .ZN(n9790) );
  NOR3_X1 U9704 ( .A1(n8749), .A2(n9792), .A3(n8475), .ZN(n9791) );
  NOR2_X1 U9705 ( .A1(n9539), .A2(n9538), .ZN(n9792) );
  NAND2_X1 U9706 ( .A1(n9538), .A2(n9539), .ZN(n9789) );
  NAND2_X1 U9707 ( .A1(n9696), .A2(n9793), .ZN(n9539) );
  NAND2_X1 U9708 ( .A1(n9695), .A2(n9697), .ZN(n9793) );
  NAND2_X1 U9709 ( .A1(n9794), .A2(n9795), .ZN(n9697) );
  NAND2_X1 U9710 ( .A1(b_29_), .A2(a_12_), .ZN(n9795) );
  INV_X1 U9711 ( .A(n9796), .ZN(n9794) );
  XNOR2_X1 U9712 ( .A(n9797), .B(n9798), .ZN(n9695) );
  XOR2_X1 U9713 ( .A(n9799), .B(n9800), .Z(n9798) );
  NAND2_X1 U9714 ( .A1(b_28_), .A2(a_13_), .ZN(n9800) );
  NAND2_X1 U9715 ( .A1(a_12_), .A2(n9796), .ZN(n9696) );
  NAND2_X1 U9716 ( .A1(n9801), .A2(n9802), .ZN(n9796) );
  INV_X1 U9717 ( .A(n9803), .ZN(n9802) );
  NOR3_X1 U9718 ( .A1(n8721), .A2(n9804), .A3(n8475), .ZN(n9803) );
  NOR2_X1 U9719 ( .A1(n9551), .A2(n9549), .ZN(n9804) );
  NAND2_X1 U9720 ( .A1(n9549), .A2(n9551), .ZN(n9801) );
  NAND2_X1 U9721 ( .A1(n9692), .A2(n9805), .ZN(n9551) );
  NAND2_X1 U9722 ( .A1(n9691), .A2(n9693), .ZN(n9805) );
  NAND2_X1 U9723 ( .A1(n9806), .A2(n9807), .ZN(n9693) );
  NAND2_X1 U9724 ( .A1(b_29_), .A2(a_14_), .ZN(n9807) );
  XOR2_X1 U9725 ( .A(n9808), .B(n9809), .Z(n9691) );
  XOR2_X1 U9726 ( .A(n9810), .B(n9811), .Z(n9808) );
  NOR2_X1 U9727 ( .A1(n8692), .A2(n8980), .ZN(n9811) );
  INV_X1 U9728 ( .A(n9812), .ZN(n9692) );
  NOR2_X1 U9729 ( .A1(n8991), .A2(n9806), .ZN(n9812) );
  NOR2_X1 U9730 ( .A1(n9813), .A2(n9814), .ZN(n9806) );
  NOR3_X1 U9731 ( .A1(n8692), .A2(n9815), .A3(n8475), .ZN(n9814) );
  NOR2_X1 U9732 ( .A1(n9564), .A2(n9563), .ZN(n9815) );
  INV_X1 U9733 ( .A(n9816), .ZN(n9813) );
  NAND2_X1 U9734 ( .A1(n9563), .A2(n9564), .ZN(n9816) );
  NAND2_X1 U9735 ( .A1(n9688), .A2(n9817), .ZN(n9564) );
  NAND2_X1 U9736 ( .A1(n9687), .A2(n9689), .ZN(n9817) );
  NAND2_X1 U9737 ( .A1(n9818), .A2(n9819), .ZN(n9689) );
  NAND2_X1 U9738 ( .A1(b_29_), .A2(a_16_), .ZN(n9819) );
  INV_X1 U9739 ( .A(n9820), .ZN(n9818) );
  XNOR2_X1 U9740 ( .A(n9821), .B(n9822), .ZN(n9687) );
  XOR2_X1 U9741 ( .A(n9823), .B(n9824), .Z(n9822) );
  NAND2_X1 U9742 ( .A1(b_28_), .A2(a_17_), .ZN(n9824) );
  NAND2_X1 U9743 ( .A1(a_16_), .A2(n9820), .ZN(n9688) );
  NAND2_X1 U9744 ( .A1(n9825), .A2(n9826), .ZN(n9820) );
  NAND3_X1 U9745 ( .A1(a_17_), .A2(n9827), .A3(b_29_), .ZN(n9826) );
  NAND2_X1 U9746 ( .A1(n9573), .A2(n9575), .ZN(n9827) );
  INV_X1 U9747 ( .A(n9828), .ZN(n9825) );
  NOR2_X1 U9748 ( .A1(n9575), .A2(n9573), .ZN(n9828) );
  XNOR2_X1 U9749 ( .A(n9829), .B(n9830), .ZN(n9573) );
  XNOR2_X1 U9750 ( .A(n9831), .B(n9832), .ZN(n9830) );
  NAND2_X1 U9751 ( .A1(n9833), .A2(n9834), .ZN(n9575) );
  NAND2_X1 U9752 ( .A1(n9583), .A2(n9835), .ZN(n9834) );
  NAND2_X1 U9753 ( .A1(n9585), .A2(n9584), .ZN(n9835) );
  XNOR2_X1 U9754 ( .A(n9836), .B(n9837), .ZN(n9583) );
  XOR2_X1 U9755 ( .A(n9838), .B(n9839), .Z(n9836) );
  NOR2_X1 U9756 ( .A1(n8630), .A2(n8980), .ZN(n9839) );
  INV_X1 U9757 ( .A(n9840), .ZN(n9833) );
  NOR2_X1 U9758 ( .A1(n9584), .A2(n9585), .ZN(n9840) );
  NOR2_X1 U9759 ( .A1(n8475), .A2(n8988), .ZN(n9585) );
  NAND2_X1 U9760 ( .A1(n9841), .A2(n9842), .ZN(n9584) );
  NAND3_X1 U9761 ( .A1(a_19_), .A2(n9843), .A3(b_29_), .ZN(n9842) );
  INV_X1 U9762 ( .A(n9844), .ZN(n9843) );
  NOR2_X1 U9763 ( .A1(n9592), .A2(n9591), .ZN(n9844) );
  NAND2_X1 U9764 ( .A1(n9591), .A2(n9592), .ZN(n9841) );
  NAND2_X1 U9765 ( .A1(n9684), .A2(n9845), .ZN(n9592) );
  NAND2_X1 U9766 ( .A1(n9683), .A2(n9685), .ZN(n9845) );
  NAND2_X1 U9767 ( .A1(n9846), .A2(n9847), .ZN(n9685) );
  NAND2_X1 U9768 ( .A1(b_29_), .A2(a_20_), .ZN(n9847) );
  XNOR2_X1 U9769 ( .A(n9848), .B(n9849), .ZN(n9683) );
  XOR2_X1 U9770 ( .A(n9850), .B(n9851), .Z(n9849) );
  NAND2_X1 U9771 ( .A1(b_28_), .A2(a_21_), .ZN(n9851) );
  INV_X1 U9772 ( .A(n9852), .ZN(n9684) );
  NOR2_X1 U9773 ( .A1(n8986), .A2(n9846), .ZN(n9852) );
  NOR2_X1 U9774 ( .A1(n9853), .A2(n9854), .ZN(n9846) );
  NOR3_X1 U9775 ( .A1(n8601), .A2(n9855), .A3(n8475), .ZN(n9854) );
  NOR2_X1 U9776 ( .A1(n9603), .A2(n9602), .ZN(n9855) );
  INV_X1 U9777 ( .A(n9856), .ZN(n9853) );
  NAND2_X1 U9778 ( .A1(n9602), .A2(n9603), .ZN(n9856) );
  NAND2_X1 U9779 ( .A1(n9680), .A2(n9857), .ZN(n9603) );
  NAND2_X1 U9780 ( .A1(n9679), .A2(n9681), .ZN(n9857) );
  NAND2_X1 U9781 ( .A1(n9858), .A2(n9859), .ZN(n9681) );
  NAND2_X1 U9782 ( .A1(b_29_), .A2(a_22_), .ZN(n9859) );
  INV_X1 U9783 ( .A(n9860), .ZN(n9858) );
  XNOR2_X1 U9784 ( .A(n9861), .B(n9862), .ZN(n9679) );
  NAND2_X1 U9785 ( .A1(n9863), .A2(n9864), .ZN(n9861) );
  NAND2_X1 U9786 ( .A1(a_22_), .A2(n9860), .ZN(n9680) );
  NAND2_X1 U9787 ( .A1(n9616), .A2(n9865), .ZN(n9860) );
  NAND2_X1 U9788 ( .A1(n9615), .A2(n9617), .ZN(n9865) );
  NAND2_X1 U9789 ( .A1(n9866), .A2(n9867), .ZN(n9617) );
  NAND2_X1 U9790 ( .A1(b_29_), .A2(a_23_), .ZN(n9867) );
  XNOR2_X1 U9791 ( .A(n9868), .B(n9869), .ZN(n9615) );
  XNOR2_X1 U9792 ( .A(n9870), .B(n9871), .ZN(n9868) );
  NAND2_X1 U9793 ( .A1(a_23_), .A2(n9872), .ZN(n9616) );
  INV_X1 U9794 ( .A(n9866), .ZN(n9872) );
  NOR2_X1 U9795 ( .A1(n9873), .A2(n9874), .ZN(n9866) );
  INV_X1 U9796 ( .A(n9875), .ZN(n9874) );
  NAND2_X1 U9797 ( .A1(n9625), .A2(n9876), .ZN(n9875) );
  NAND2_X1 U9798 ( .A1(n9624), .A2(n9623), .ZN(n9876) );
  NOR2_X1 U9799 ( .A1(n8475), .A2(n8982), .ZN(n9625) );
  NOR2_X1 U9800 ( .A1(n9623), .A2(n9624), .ZN(n9873) );
  NOR2_X1 U9801 ( .A1(n9877), .A2(n9878), .ZN(n9624) );
  INV_X1 U9802 ( .A(n9879), .ZN(n9878) );
  NAND2_X1 U9803 ( .A1(n9677), .A2(n9880), .ZN(n9879) );
  NAND2_X1 U9804 ( .A1(n9674), .A2(n9676), .ZN(n9880) );
  NOR2_X1 U9805 ( .A1(n8475), .A2(n8541), .ZN(n9677) );
  NOR2_X1 U9806 ( .A1(n9676), .A2(n9674), .ZN(n9877) );
  XNOR2_X1 U9807 ( .A(n9881), .B(n9882), .ZN(n9674) );
  XNOR2_X1 U9808 ( .A(n9883), .B(n9884), .ZN(n9882) );
  NAND2_X1 U9809 ( .A1(n9885), .A2(n9886), .ZN(n9676) );
  NAND2_X1 U9810 ( .A1(n9635), .A2(n9887), .ZN(n9886) );
  NAND2_X1 U9811 ( .A1(n9638), .A2(n9637), .ZN(n9887) );
  XNOR2_X1 U9812 ( .A(n9888), .B(n9889), .ZN(n9635) );
  XOR2_X1 U9813 ( .A(n9890), .B(n9891), .Z(n9888) );
  INV_X1 U9814 ( .A(n9892), .ZN(n9885) );
  NOR2_X1 U9815 ( .A1(n9637), .A2(n9638), .ZN(n9892) );
  NOR2_X1 U9816 ( .A1(n8475), .A2(n9893), .ZN(n9638) );
  NAND2_X1 U9817 ( .A1(n9894), .A2(n9895), .ZN(n9637) );
  NAND3_X1 U9818 ( .A1(a_27_), .A2(n9896), .A3(b_29_), .ZN(n9895) );
  NAND2_X1 U9819 ( .A1(n9645), .A2(n9897), .ZN(n9896) );
  INV_X1 U9820 ( .A(n9643), .ZN(n9897) );
  NAND2_X1 U9821 ( .A1(n9643), .A2(n9898), .ZN(n9894) );
  INV_X1 U9822 ( .A(n9645), .ZN(n9898) );
  NOR2_X1 U9823 ( .A1(n9899), .A2(n9900), .ZN(n9645) );
  INV_X1 U9824 ( .A(n9901), .ZN(n9900) );
  NAND2_X1 U9825 ( .A1(n9673), .A2(n9902), .ZN(n9901) );
  NAND2_X1 U9826 ( .A1(n9671), .A2(n9672), .ZN(n9902) );
  NOR2_X1 U9827 ( .A1(n8475), .A2(n8493), .ZN(n9673) );
  NOR2_X1 U9828 ( .A1(n9672), .A2(n9671), .ZN(n9899) );
  XNOR2_X1 U9829 ( .A(n9903), .B(n9904), .ZN(n9671) );
  XNOR2_X1 U9830 ( .A(n9905), .B(n9906), .ZN(n9903) );
  NAND2_X1 U9831 ( .A1(n9907), .A2(n9908), .ZN(n9672) );
  NAND2_X1 U9832 ( .A1(n9909), .A2(n9669), .ZN(n9908) );
  NAND3_X1 U9833 ( .A1(b_28_), .A2(n9666), .A3(b_29_), .ZN(n9669) );
  NAND2_X1 U9834 ( .A1(n8470), .A2(n9668), .ZN(n9909) );
  INV_X1 U9835 ( .A(n9910), .ZN(n9907) );
  NOR2_X1 U9836 ( .A1(n9668), .A2(n8470), .ZN(n9910) );
  NOR2_X1 U9837 ( .A1(n8475), .A2(n8473), .ZN(n8470) );
  NAND2_X1 U9838 ( .A1(n9911), .A2(n9912), .ZN(n9668) );
  NAND2_X1 U9839 ( .A1(b_27_), .A2(n9913), .ZN(n9912) );
  NAND2_X1 U9840 ( .A1(n8456), .A2(n9914), .ZN(n9913) );
  NAND2_X1 U9841 ( .A1(a_31_), .A2(n8980), .ZN(n9914) );
  NAND2_X1 U9842 ( .A1(b_28_), .A2(n9915), .ZN(n9911) );
  NAND2_X1 U9843 ( .A1(n8459), .A2(n9916), .ZN(n9915) );
  NAND2_X1 U9844 ( .A1(a_30_), .A2(n8514), .ZN(n9916) );
  XNOR2_X1 U9845 ( .A(n9917), .B(n9918), .ZN(n9643) );
  XOR2_X1 U9846 ( .A(n8486), .B(n9919), .Z(n9917) );
  XOR2_X1 U9847 ( .A(n9920), .B(n9921), .Z(n9623) );
  XNOR2_X1 U9848 ( .A(n9922), .B(n9923), .ZN(n9921) );
  XNOR2_X1 U9849 ( .A(n9924), .B(n9925), .ZN(n9602) );
  NAND2_X1 U9850 ( .A1(n9926), .A2(n9927), .ZN(n9924) );
  XNOR2_X1 U9851 ( .A(n9928), .B(n9929), .ZN(n9591) );
  NAND2_X1 U9852 ( .A1(n9930), .A2(n9931), .ZN(n9928) );
  XNOR2_X1 U9853 ( .A(n9932), .B(n9933), .ZN(n9563) );
  NAND2_X1 U9854 ( .A1(n9934), .A2(n9935), .ZN(n9932) );
  XNOR2_X1 U9855 ( .A(n9936), .B(n9937), .ZN(n9549) );
  NAND2_X1 U9856 ( .A1(n9938), .A2(n9939), .ZN(n9936) );
  XNOR2_X1 U9857 ( .A(n9940), .B(n9941), .ZN(n9538) );
  NAND2_X1 U9858 ( .A1(n9942), .A2(n9943), .ZN(n9940) );
  XNOR2_X1 U9859 ( .A(n9944), .B(n9945), .ZN(n9526) );
  NAND2_X1 U9860 ( .A1(n9946), .A2(n9947), .ZN(n9944) );
  XNOR2_X1 U9861 ( .A(n9948), .B(n9949), .ZN(n9515) );
  NAND2_X1 U9862 ( .A1(n9950), .A2(n9951), .ZN(n9948) );
  XNOR2_X1 U9863 ( .A(n9952), .B(n9953), .ZN(n9503) );
  NAND2_X1 U9864 ( .A1(n9954), .A2(n9955), .ZN(n9952) );
  NAND2_X1 U9865 ( .A1(n9481), .A2(n9478), .ZN(n9732) );
  XNOR2_X1 U9866 ( .A(n9956), .B(n9957), .ZN(n9478) );
  XOR2_X1 U9867 ( .A(n9958), .B(n9959), .Z(n9957) );
  NAND2_X1 U9868 ( .A1(b_28_), .A2(a_3_), .ZN(n9959) );
  NOR2_X1 U9869 ( .A1(n8475), .A2(n8998), .ZN(n9481) );
  INV_X1 U9870 ( .A(b_29_), .ZN(n8475) );
  XOR2_X1 U9871 ( .A(n9960), .B(n9961), .Z(n9711) );
  XOR2_X1 U9872 ( .A(n9962), .B(n9963), .Z(n9961) );
  XOR2_X1 U9873 ( .A(n9964), .B(n9965), .Z(n9214) );
  XOR2_X1 U9874 ( .A(n9966), .B(n9967), .Z(n9964) );
  NOR2_X1 U9875 ( .A1(n9471), .A2(n8980), .ZN(n9967) );
  NAND4_X1 U9876 ( .A1(n9209), .A2(n9208), .A3(n9210), .A4(n9036), .ZN(n9028)
         );
  INV_X1 U9877 ( .A(n9968), .ZN(n9036) );
  NAND2_X1 U9878 ( .A1(n9969), .A2(n9970), .ZN(n9210) );
  NAND3_X1 U9879 ( .A1(a_0_), .A2(n9971), .A3(b_28_), .ZN(n9970) );
  INV_X1 U9880 ( .A(n9972), .ZN(n9971) );
  NOR2_X1 U9881 ( .A1(n9966), .A2(n9965), .ZN(n9972) );
  NAND2_X1 U9882 ( .A1(n9965), .A2(n9966), .ZN(n9969) );
  NAND2_X1 U9883 ( .A1(n9973), .A2(n9974), .ZN(n9966) );
  NAND2_X1 U9884 ( .A1(n9726), .A2(n9975), .ZN(n9974) );
  INV_X1 U9885 ( .A(n9976), .ZN(n9975) );
  NOR2_X1 U9886 ( .A1(n9725), .A2(n9724), .ZN(n9976) );
  NOR2_X1 U9887 ( .A1(n8980), .A2(n9731), .ZN(n9726) );
  NAND2_X1 U9888 ( .A1(n9724), .A2(n9725), .ZN(n9973) );
  NAND2_X1 U9889 ( .A1(n9977), .A2(n9978), .ZN(n9725) );
  NAND2_X1 U9890 ( .A1(n9962), .A2(n9979), .ZN(n9978) );
  NAND2_X1 U9891 ( .A1(n9963), .A2(n9960), .ZN(n9979) );
  NOR2_X1 U9892 ( .A1(n8980), .A2(n8998), .ZN(n9962) );
  INV_X1 U9893 ( .A(n9980), .ZN(n9977) );
  NOR2_X1 U9894 ( .A1(n9960), .A2(n9963), .ZN(n9980) );
  NOR2_X1 U9895 ( .A1(n9981), .A2(n9982), .ZN(n9963) );
  NOR3_X1 U9896 ( .A1(n8877), .A2(n9983), .A3(n8980), .ZN(n9982) );
  NOR2_X1 U9897 ( .A1(n9958), .A2(n9956), .ZN(n9983) );
  INV_X1 U9898 ( .A(n9984), .ZN(n9981) );
  NAND2_X1 U9899 ( .A1(n9956), .A2(n9958), .ZN(n9984) );
  NAND2_X1 U9900 ( .A1(n9985), .A2(n9986), .ZN(n9958) );
  INV_X1 U9901 ( .A(n9987), .ZN(n9986) );
  NOR3_X1 U9902 ( .A1(n8996), .A2(n9988), .A3(n8980), .ZN(n9987) );
  NOR2_X1 U9903 ( .A1(n9743), .A2(n9741), .ZN(n9988) );
  NAND2_X1 U9904 ( .A1(n9741), .A2(n9743), .ZN(n9985) );
  NAND2_X1 U9905 ( .A1(n9989), .A2(n9990), .ZN(n9743) );
  NAND3_X1 U9906 ( .A1(a_5_), .A2(n9991), .A3(b_28_), .ZN(n9990) );
  INV_X1 U9907 ( .A(n9992), .ZN(n9991) );
  NOR2_X1 U9908 ( .A1(n9750), .A2(n9749), .ZN(n9992) );
  NAND2_X1 U9909 ( .A1(n9749), .A2(n9750), .ZN(n9989) );
  NAND2_X1 U9910 ( .A1(n9954), .A2(n9993), .ZN(n9750) );
  NAND2_X1 U9911 ( .A1(n9953), .A2(n9955), .ZN(n9993) );
  NAND2_X1 U9912 ( .A1(n9994), .A2(n9995), .ZN(n9955) );
  NAND2_X1 U9913 ( .A1(b_28_), .A2(a_6_), .ZN(n9995) );
  INV_X1 U9914 ( .A(n9996), .ZN(n9994) );
  XOR2_X1 U9915 ( .A(n9997), .B(n9998), .Z(n9953) );
  XOR2_X1 U9916 ( .A(n9999), .B(n10000), .Z(n9997) );
  NOR2_X1 U9917 ( .A1(n8817), .A2(n8514), .ZN(n10000) );
  NAND2_X1 U9918 ( .A1(a_6_), .A2(n9996), .ZN(n9954) );
  NAND2_X1 U9919 ( .A1(n10001), .A2(n10002), .ZN(n9996) );
  INV_X1 U9920 ( .A(n10003), .ZN(n10002) );
  NOR3_X1 U9921 ( .A1(n8817), .A2(n10004), .A3(n8980), .ZN(n10003) );
  NOR2_X1 U9922 ( .A1(n9762), .A2(n9760), .ZN(n10004) );
  NAND2_X1 U9923 ( .A1(n9760), .A2(n9762), .ZN(n10001) );
  NAND2_X1 U9924 ( .A1(n9950), .A2(n10005), .ZN(n9762) );
  NAND2_X1 U9925 ( .A1(n9949), .A2(n9951), .ZN(n10005) );
  NAND2_X1 U9926 ( .A1(n10006), .A2(n10007), .ZN(n9951) );
  NAND2_X1 U9927 ( .A1(b_28_), .A2(a_8_), .ZN(n10007) );
  INV_X1 U9928 ( .A(n10008), .ZN(n10006) );
  XNOR2_X1 U9929 ( .A(n10009), .B(n10010), .ZN(n9949) );
  XOR2_X1 U9930 ( .A(n10011), .B(n10012), .Z(n10010) );
  NAND2_X1 U9931 ( .A1(b_27_), .A2(a_9_), .ZN(n10012) );
  NAND2_X1 U9932 ( .A1(a_8_), .A2(n10008), .ZN(n9950) );
  NAND2_X1 U9933 ( .A1(n10013), .A2(n10014), .ZN(n10008) );
  INV_X1 U9934 ( .A(n10015), .ZN(n10014) );
  NOR3_X1 U9935 ( .A1(n8779), .A2(n10016), .A3(n8980), .ZN(n10015) );
  NOR2_X1 U9936 ( .A1(n9775), .A2(n9773), .ZN(n10016) );
  NAND2_X1 U9937 ( .A1(n9773), .A2(n9775), .ZN(n10013) );
  NAND2_X1 U9938 ( .A1(n9946), .A2(n10017), .ZN(n9775) );
  NAND2_X1 U9939 ( .A1(n9945), .A2(n9947), .ZN(n10017) );
  NAND2_X1 U9940 ( .A1(n10018), .A2(n10019), .ZN(n9947) );
  NAND2_X1 U9941 ( .A1(b_28_), .A2(a_10_), .ZN(n10019) );
  XOR2_X1 U9942 ( .A(n10020), .B(n10021), .Z(n9945) );
  XOR2_X1 U9943 ( .A(n10022), .B(n10023), .Z(n10020) );
  NOR2_X1 U9944 ( .A1(n8749), .A2(n8514), .ZN(n10023) );
  INV_X1 U9945 ( .A(n10024), .ZN(n9946) );
  NOR2_X1 U9946 ( .A1(n8769), .A2(n10018), .ZN(n10024) );
  NOR2_X1 U9947 ( .A1(n10025), .A2(n10026), .ZN(n10018) );
  NOR3_X1 U9948 ( .A1(n8749), .A2(n10027), .A3(n8980), .ZN(n10026) );
  NOR2_X1 U9949 ( .A1(n9787), .A2(n9786), .ZN(n10027) );
  INV_X1 U9950 ( .A(n10028), .ZN(n10025) );
  NAND2_X1 U9951 ( .A1(n9786), .A2(n9787), .ZN(n10028) );
  NAND2_X1 U9952 ( .A1(n9942), .A2(n10029), .ZN(n9787) );
  NAND2_X1 U9953 ( .A1(n9941), .A2(n9943), .ZN(n10029) );
  NAND2_X1 U9954 ( .A1(n10030), .A2(n10031), .ZN(n9943) );
  NAND2_X1 U9955 ( .A1(b_28_), .A2(a_12_), .ZN(n10031) );
  INV_X1 U9956 ( .A(n10032), .ZN(n10030) );
  XNOR2_X1 U9957 ( .A(n10033), .B(n10034), .ZN(n9941) );
  XOR2_X1 U9958 ( .A(n10035), .B(n10036), .Z(n10034) );
  NAND2_X1 U9959 ( .A1(b_27_), .A2(a_13_), .ZN(n10036) );
  NAND2_X1 U9960 ( .A1(a_12_), .A2(n10032), .ZN(n9942) );
  NAND2_X1 U9961 ( .A1(n10037), .A2(n10038), .ZN(n10032) );
  INV_X1 U9962 ( .A(n10039), .ZN(n10038) );
  NOR3_X1 U9963 ( .A1(n8721), .A2(n10040), .A3(n8980), .ZN(n10039) );
  NOR2_X1 U9964 ( .A1(n9799), .A2(n9797), .ZN(n10040) );
  NAND2_X1 U9965 ( .A1(n9797), .A2(n9799), .ZN(n10037) );
  NAND2_X1 U9966 ( .A1(n9938), .A2(n10041), .ZN(n9799) );
  NAND2_X1 U9967 ( .A1(n9937), .A2(n9939), .ZN(n10041) );
  NAND2_X1 U9968 ( .A1(n10042), .A2(n10043), .ZN(n9939) );
  NAND2_X1 U9969 ( .A1(b_28_), .A2(a_14_), .ZN(n10043) );
  INV_X1 U9970 ( .A(n10044), .ZN(n10042) );
  XOR2_X1 U9971 ( .A(n10045), .B(n10046), .Z(n9937) );
  XOR2_X1 U9972 ( .A(n10047), .B(n10048), .Z(n10045) );
  NOR2_X1 U9973 ( .A1(n8692), .A2(n8514), .ZN(n10048) );
  NAND2_X1 U9974 ( .A1(a_14_), .A2(n10044), .ZN(n9938) );
  NAND2_X1 U9975 ( .A1(n10049), .A2(n10050), .ZN(n10044) );
  INV_X1 U9976 ( .A(n10051), .ZN(n10050) );
  NOR3_X1 U9977 ( .A1(n8692), .A2(n10052), .A3(n8980), .ZN(n10051) );
  NOR2_X1 U9978 ( .A1(n9810), .A2(n9809), .ZN(n10052) );
  NAND2_X1 U9979 ( .A1(n9809), .A2(n9810), .ZN(n10049) );
  NAND2_X1 U9980 ( .A1(n9934), .A2(n10053), .ZN(n9810) );
  NAND2_X1 U9981 ( .A1(n9933), .A2(n9935), .ZN(n10053) );
  NAND2_X1 U9982 ( .A1(n10054), .A2(n10055), .ZN(n9935) );
  NAND2_X1 U9983 ( .A1(b_28_), .A2(a_16_), .ZN(n10055) );
  XNOR2_X1 U9984 ( .A(n10056), .B(n10057), .ZN(n9933) );
  XOR2_X1 U9985 ( .A(n10058), .B(n10059), .Z(n10057) );
  NAND2_X1 U9986 ( .A1(b_27_), .A2(a_17_), .ZN(n10059) );
  NAND2_X1 U9987 ( .A1(a_16_), .A2(n10060), .ZN(n9934) );
  INV_X1 U9988 ( .A(n10054), .ZN(n10060) );
  NOR2_X1 U9989 ( .A1(n10061), .A2(n10062), .ZN(n10054) );
  NOR3_X1 U9990 ( .A1(n8662), .A2(n10063), .A3(n8980), .ZN(n10062) );
  INV_X1 U9991 ( .A(n10064), .ZN(n10063) );
  NAND2_X1 U9992 ( .A1(n9821), .A2(n9823), .ZN(n10064) );
  NOR2_X1 U9993 ( .A1(n9823), .A2(n9821), .ZN(n10061) );
  XOR2_X1 U9994 ( .A(n10065), .B(n10066), .Z(n9821) );
  XOR2_X1 U9995 ( .A(n10067), .B(n10068), .Z(n10065) );
  NAND2_X1 U9996 ( .A1(n10069), .A2(n10070), .ZN(n9823) );
  NAND2_X1 U9997 ( .A1(n9829), .A2(n10071), .ZN(n10070) );
  NAND2_X1 U9998 ( .A1(n9832), .A2(n9831), .ZN(n10071) );
  XOR2_X1 U9999 ( .A(n10072), .B(n10073), .Z(n9829) );
  XOR2_X1 U10000 ( .A(n10074), .B(n10075), .Z(n10073) );
  NAND2_X1 U10001 ( .A1(b_27_), .A2(a_19_), .ZN(n10075) );
  INV_X1 U10002 ( .A(n10076), .ZN(n10069) );
  NOR2_X1 U10003 ( .A1(n9831), .A2(n9832), .ZN(n10076) );
  NOR2_X1 U10004 ( .A1(n8980), .A2(n8988), .ZN(n9832) );
  NAND2_X1 U10005 ( .A1(n10077), .A2(n10078), .ZN(n9831) );
  NAND3_X1 U10006 ( .A1(a_19_), .A2(n10079), .A3(b_28_), .ZN(n10078) );
  INV_X1 U10007 ( .A(n10080), .ZN(n10079) );
  NOR2_X1 U10008 ( .A1(n9838), .A2(n9837), .ZN(n10080) );
  NAND2_X1 U10009 ( .A1(n9837), .A2(n9838), .ZN(n10077) );
  NAND2_X1 U10010 ( .A1(n9930), .A2(n10081), .ZN(n9838) );
  NAND2_X1 U10011 ( .A1(n9929), .A2(n9931), .ZN(n10081) );
  NAND2_X1 U10012 ( .A1(n10082), .A2(n10083), .ZN(n9931) );
  NAND2_X1 U10013 ( .A1(b_28_), .A2(a_20_), .ZN(n10083) );
  INV_X1 U10014 ( .A(n10084), .ZN(n10082) );
  XNOR2_X1 U10015 ( .A(n10085), .B(n10086), .ZN(n9929) );
  XOR2_X1 U10016 ( .A(n10087), .B(n10088), .Z(n10086) );
  NAND2_X1 U10017 ( .A1(b_27_), .A2(a_21_), .ZN(n10088) );
  NAND2_X1 U10018 ( .A1(a_20_), .A2(n10084), .ZN(n9930) );
  NAND2_X1 U10019 ( .A1(n10089), .A2(n10090), .ZN(n10084) );
  INV_X1 U10020 ( .A(n10091), .ZN(n10090) );
  NOR3_X1 U10021 ( .A1(n8601), .A2(n10092), .A3(n8980), .ZN(n10091) );
  NOR2_X1 U10022 ( .A1(n9850), .A2(n9848), .ZN(n10092) );
  NAND2_X1 U10023 ( .A1(n9848), .A2(n9850), .ZN(n10089) );
  NAND2_X1 U10024 ( .A1(n9926), .A2(n10093), .ZN(n9850) );
  NAND2_X1 U10025 ( .A1(n9925), .A2(n9927), .ZN(n10093) );
  NAND2_X1 U10026 ( .A1(n10094), .A2(n10095), .ZN(n9927) );
  NAND2_X1 U10027 ( .A1(b_28_), .A2(a_22_), .ZN(n10095) );
  INV_X1 U10028 ( .A(n10096), .ZN(n10094) );
  XNOR2_X1 U10029 ( .A(n10097), .B(n10098), .ZN(n9925) );
  NAND2_X1 U10030 ( .A1(n10099), .A2(n10100), .ZN(n10097) );
  NAND2_X1 U10031 ( .A1(a_22_), .A2(n10096), .ZN(n9926) );
  NAND2_X1 U10032 ( .A1(n9863), .A2(n10101), .ZN(n10096) );
  NAND2_X1 U10033 ( .A1(n9862), .A2(n9864), .ZN(n10101) );
  NAND2_X1 U10034 ( .A1(n10102), .A2(n10103), .ZN(n9864) );
  NAND2_X1 U10035 ( .A1(b_28_), .A2(a_23_), .ZN(n10103) );
  INV_X1 U10036 ( .A(n10104), .ZN(n10102) );
  XNOR2_X1 U10037 ( .A(n10105), .B(n10106), .ZN(n9862) );
  XOR2_X1 U10038 ( .A(n10107), .B(n10108), .Z(n10106) );
  NAND2_X1 U10039 ( .A1(a_23_), .A2(n10104), .ZN(n9863) );
  NAND2_X1 U10040 ( .A1(n10109), .A2(n10110), .ZN(n10104) );
  NAND2_X1 U10041 ( .A1(n9871), .A2(n10111), .ZN(n10110) );
  NAND2_X1 U10042 ( .A1(n9870), .A2(n9869), .ZN(n10111) );
  NOR2_X1 U10043 ( .A1(n8980), .A2(n8982), .ZN(n9871) );
  NAND2_X1 U10044 ( .A1(n10112), .A2(n10113), .ZN(n10109) );
  INV_X1 U10045 ( .A(n9870), .ZN(n10113) );
  NOR2_X1 U10046 ( .A1(n10114), .A2(n10115), .ZN(n9870) );
  INV_X1 U10047 ( .A(n10116), .ZN(n10115) );
  NAND2_X1 U10048 ( .A1(n9923), .A2(n10117), .ZN(n10116) );
  NAND2_X1 U10049 ( .A1(n9920), .A2(n9922), .ZN(n10117) );
  NOR2_X1 U10050 ( .A1(n8980), .A2(n8541), .ZN(n9923) );
  NOR2_X1 U10051 ( .A1(n9922), .A2(n9920), .ZN(n10114) );
  XOR2_X1 U10052 ( .A(n10118), .B(n10119), .Z(n9920) );
  NAND2_X1 U10053 ( .A1(n10120), .A2(n10121), .ZN(n10118) );
  NAND2_X1 U10054 ( .A1(n10122), .A2(n10123), .ZN(n9922) );
  NAND2_X1 U10055 ( .A1(n9881), .A2(n10124), .ZN(n10123) );
  INV_X1 U10056 ( .A(n10125), .ZN(n10124) );
  NOR2_X1 U10057 ( .A1(n9884), .A2(n9883), .ZN(n10125) );
  XOR2_X1 U10058 ( .A(n10126), .B(n10127), .Z(n9881) );
  XOR2_X1 U10059 ( .A(n10128), .B(n8509), .Z(n10126) );
  NAND2_X1 U10060 ( .A1(n9883), .A2(n9884), .ZN(n10122) );
  NAND2_X1 U10061 ( .A1(b_28_), .A2(a_26_), .ZN(n9884) );
  NOR2_X1 U10062 ( .A1(n10129), .A2(n10130), .ZN(n9883) );
  INV_X1 U10063 ( .A(n10131), .ZN(n10130) );
  NAND2_X1 U10064 ( .A1(n9891), .A2(n10132), .ZN(n10131) );
  NAND2_X1 U10065 ( .A1(n9889), .A2(n9890), .ZN(n10132) );
  NOR2_X1 U10066 ( .A1(n8980), .A2(n8512), .ZN(n9891) );
  NOR2_X1 U10067 ( .A1(n9890), .A2(n9889), .ZN(n10129) );
  XNOR2_X1 U10068 ( .A(n10133), .B(n10134), .ZN(n9889) );
  XOR2_X1 U10069 ( .A(n10135), .B(n10136), .Z(n10133) );
  NAND2_X1 U10070 ( .A1(n10137), .A2(n10138), .ZN(n9890) );
  NAND2_X1 U10071 ( .A1(n9918), .A2(n10139), .ZN(n10138) );
  INV_X1 U10072 ( .A(n10140), .ZN(n10139) );
  NOR2_X1 U10073 ( .A1(n8486), .A2(n9919), .ZN(n10140) );
  XNOR2_X1 U10074 ( .A(n10141), .B(n10142), .ZN(n9918) );
  XOR2_X1 U10075 ( .A(n10143), .B(n10144), .Z(n10141) );
  NAND2_X1 U10076 ( .A1(n9919), .A2(n8486), .ZN(n10137) );
  NAND2_X1 U10077 ( .A1(b_28_), .A2(a_28_), .ZN(n8486) );
  NOR2_X1 U10078 ( .A1(n10145), .A2(n10146), .ZN(n9919) );
  INV_X1 U10079 ( .A(n10147), .ZN(n10146) );
  NAND2_X1 U10080 ( .A1(n9904), .A2(n10148), .ZN(n10147) );
  NAND2_X1 U10081 ( .A1(n10149), .A2(n9906), .ZN(n10148) );
  NOR2_X1 U10082 ( .A1(n8980), .A2(n8473), .ZN(n9904) );
  INV_X1 U10083 ( .A(b_28_), .ZN(n8980) );
  NOR2_X1 U10084 ( .A1(n9906), .A2(n10149), .ZN(n10145) );
  INV_X1 U10085 ( .A(n9905), .ZN(n10149) );
  NAND2_X1 U10086 ( .A1(n10150), .A2(n10151), .ZN(n9905) );
  NAND2_X1 U10087 ( .A1(b_26_), .A2(n10152), .ZN(n10151) );
  NAND2_X1 U10088 ( .A1(n8456), .A2(n10153), .ZN(n10152) );
  NAND2_X1 U10089 ( .A1(a_31_), .A2(n8514), .ZN(n10153) );
  NAND2_X1 U10090 ( .A1(b_27_), .A2(n10154), .ZN(n10150) );
  NAND2_X1 U10091 ( .A1(n8459), .A2(n10155), .ZN(n10154) );
  NAND2_X1 U10092 ( .A1(a_30_), .A2(n10156), .ZN(n10155) );
  NAND3_X1 U10093 ( .A1(b_27_), .A2(n9666), .A3(b_28_), .ZN(n9906) );
  INV_X1 U10094 ( .A(n9869), .ZN(n10112) );
  XOR2_X1 U10095 ( .A(n10157), .B(n10158), .Z(n9869) );
  NAND2_X1 U10096 ( .A1(n10159), .A2(n10160), .ZN(n10157) );
  XNOR2_X1 U10097 ( .A(n10161), .B(n10162), .ZN(n9848) );
  NAND2_X1 U10098 ( .A1(n10163), .A2(n10164), .ZN(n10161) );
  XNOR2_X1 U10099 ( .A(n10165), .B(n10166), .ZN(n9837) );
  NAND2_X1 U10100 ( .A1(n10167), .A2(n10168), .ZN(n10165) );
  XNOR2_X1 U10101 ( .A(n10169), .B(n10170), .ZN(n9809) );
  NAND2_X1 U10102 ( .A1(n10171), .A2(n10172), .ZN(n10169) );
  XNOR2_X1 U10103 ( .A(n10173), .B(n10174), .ZN(n9797) );
  NAND2_X1 U10104 ( .A1(n10175), .A2(n10176), .ZN(n10173) );
  XNOR2_X1 U10105 ( .A(n10177), .B(n10178), .ZN(n9786) );
  NAND2_X1 U10106 ( .A1(n10179), .A2(n10180), .ZN(n10177) );
  XNOR2_X1 U10107 ( .A(n10181), .B(n10182), .ZN(n9773) );
  NAND2_X1 U10108 ( .A1(n10183), .A2(n10184), .ZN(n10181) );
  XNOR2_X1 U10109 ( .A(n10185), .B(n10186), .ZN(n9760) );
  NAND2_X1 U10110 ( .A1(n10187), .A2(n10188), .ZN(n10185) );
  XOR2_X1 U10111 ( .A(n10189), .B(n10190), .Z(n9749) );
  XNOR2_X1 U10112 ( .A(n10191), .B(n10192), .ZN(n10190) );
  XOR2_X1 U10113 ( .A(n10193), .B(n10194), .Z(n9741) );
  XOR2_X1 U10114 ( .A(n10195), .B(n10196), .Z(n10193) );
  XOR2_X1 U10115 ( .A(n10197), .B(n10198), .Z(n9956) );
  XOR2_X1 U10116 ( .A(n10199), .B(n10200), .Z(n10197) );
  XNOR2_X1 U10117 ( .A(n10201), .B(n10202), .ZN(n9960) );
  XOR2_X1 U10118 ( .A(n10203), .B(n10204), .Z(n10201) );
  NOR2_X1 U10119 ( .A1(n8877), .A2(n8514), .ZN(n10204) );
  XNOR2_X1 U10120 ( .A(n10205), .B(n10206), .ZN(n9724) );
  NAND2_X1 U10121 ( .A1(n10207), .A2(n10208), .ZN(n10205) );
  XOR2_X1 U10122 ( .A(n10209), .B(n10210), .Z(n9965) );
  XOR2_X1 U10123 ( .A(n10211), .B(n10212), .Z(n10209) );
  NOR2_X1 U10124 ( .A1(n9731), .A2(n8514), .ZN(n10212) );
  NAND2_X1 U10125 ( .A1(n10213), .A2(n10214), .ZN(n9208) );
  XOR2_X1 U10126 ( .A(n10215), .B(n10216), .Z(n9209) );
  XNOR2_X1 U10127 ( .A(n10217), .B(n10218), .ZN(n10216) );
  NAND2_X1 U10128 ( .A1(n9968), .A2(n9037), .ZN(n9033) );
  XOR2_X1 U10129 ( .A(n9203), .B(n9202), .Z(n9037) );
  NOR2_X1 U10130 ( .A1(n10214), .A2(n10213), .ZN(n9968) );
  XOR2_X1 U10131 ( .A(n10219), .B(n10220), .Z(n10213) );
  NAND2_X1 U10132 ( .A1(n10221), .A2(n10222), .ZN(n10219) );
  NAND2_X1 U10133 ( .A1(n10223), .A2(n10224), .ZN(n10214) );
  NAND2_X1 U10134 ( .A1(n10215), .A2(n10225), .ZN(n10224) );
  NAND2_X1 U10135 ( .A1(n10218), .A2(n10217), .ZN(n10225) );
  XOR2_X1 U10136 ( .A(n10226), .B(n10227), .Z(n10215) );
  XOR2_X1 U10137 ( .A(n10228), .B(n10229), .Z(n10226) );
  INV_X1 U10138 ( .A(n10230), .ZN(n10223) );
  NOR2_X1 U10139 ( .A1(n10217), .A2(n10218), .ZN(n10230) );
  NOR2_X1 U10140 ( .A1(n8514), .A2(n9471), .ZN(n10218) );
  NAND2_X1 U10141 ( .A1(n10231), .A2(n10232), .ZN(n10217) );
  NAND3_X1 U10142 ( .A1(a_1_), .A2(n10233), .A3(b_27_), .ZN(n10232) );
  INV_X1 U10143 ( .A(n10234), .ZN(n10233) );
  NOR2_X1 U10144 ( .A1(n10211), .A2(n10210), .ZN(n10234) );
  NAND2_X1 U10145 ( .A1(n10210), .A2(n10211), .ZN(n10231) );
  NAND2_X1 U10146 ( .A1(n10207), .A2(n10235), .ZN(n10211) );
  NAND2_X1 U10147 ( .A1(n10206), .A2(n10208), .ZN(n10235) );
  NAND2_X1 U10148 ( .A1(n10236), .A2(n10237), .ZN(n10208) );
  NAND2_X1 U10149 ( .A1(b_27_), .A2(a_2_), .ZN(n10237) );
  INV_X1 U10150 ( .A(n10238), .ZN(n10236) );
  XNOR2_X1 U10151 ( .A(n10239), .B(n10240), .ZN(n10206) );
  XNOR2_X1 U10152 ( .A(n10241), .B(n10242), .ZN(n10239) );
  NOR2_X1 U10153 ( .A1(n8877), .A2(n10156), .ZN(n10242) );
  NAND2_X1 U10154 ( .A1(a_2_), .A2(n10238), .ZN(n10207) );
  NAND2_X1 U10155 ( .A1(n10243), .A2(n10244), .ZN(n10238) );
  INV_X1 U10156 ( .A(n10245), .ZN(n10244) );
  NOR3_X1 U10157 ( .A1(n8877), .A2(n10246), .A3(n8514), .ZN(n10245) );
  NOR2_X1 U10158 ( .A1(n10203), .A2(n10202), .ZN(n10246) );
  NAND2_X1 U10159 ( .A1(n10202), .A2(n10203), .ZN(n10243) );
  NAND2_X1 U10160 ( .A1(n10247), .A2(n10248), .ZN(n10203) );
  NAND2_X1 U10161 ( .A1(n10200), .A2(n10249), .ZN(n10248) );
  INV_X1 U10162 ( .A(n10250), .ZN(n10249) );
  NOR2_X1 U10163 ( .A1(n10199), .A2(n10198), .ZN(n10250) );
  NOR2_X1 U10164 ( .A1(n8514), .A2(n8996), .ZN(n10200) );
  NAND2_X1 U10165 ( .A1(n10198), .A2(n10199), .ZN(n10247) );
  NAND2_X1 U10166 ( .A1(n10251), .A2(n10252), .ZN(n10199) );
  NAND2_X1 U10167 ( .A1(n10196), .A2(n10253), .ZN(n10252) );
  INV_X1 U10168 ( .A(n10254), .ZN(n10253) );
  NOR2_X1 U10169 ( .A1(n10195), .A2(n10194), .ZN(n10254) );
  NOR2_X1 U10170 ( .A1(n8514), .A2(n8848), .ZN(n10196) );
  NAND2_X1 U10171 ( .A1(n10194), .A2(n10195), .ZN(n10251) );
  NAND2_X1 U10172 ( .A1(n10255), .A2(n10256), .ZN(n10195) );
  NAND2_X1 U10173 ( .A1(n10191), .A2(n10257), .ZN(n10256) );
  NAND2_X1 U10174 ( .A1(n10189), .A2(n10258), .ZN(n10257) );
  INV_X1 U10175 ( .A(n10192), .ZN(n10258) );
  NAND2_X1 U10176 ( .A1(n10259), .A2(n10260), .ZN(n10191) );
  INV_X1 U10177 ( .A(n10261), .ZN(n10260) );
  NOR3_X1 U10178 ( .A1(n8817), .A2(n10262), .A3(n8514), .ZN(n10261) );
  NOR2_X1 U10179 ( .A1(n9999), .A2(n9998), .ZN(n10262) );
  NAND2_X1 U10180 ( .A1(n9998), .A2(n9999), .ZN(n10259) );
  NAND2_X1 U10181 ( .A1(n10187), .A2(n10263), .ZN(n9999) );
  NAND2_X1 U10182 ( .A1(n10186), .A2(n10188), .ZN(n10263) );
  NAND2_X1 U10183 ( .A1(n10264), .A2(n10265), .ZN(n10188) );
  NAND2_X1 U10184 ( .A1(b_27_), .A2(a_8_), .ZN(n10265) );
  INV_X1 U10185 ( .A(n10266), .ZN(n10264) );
  XOR2_X1 U10186 ( .A(n10267), .B(n10268), .Z(n10186) );
  XOR2_X1 U10187 ( .A(n10269), .B(n10270), .Z(n10267) );
  NOR2_X1 U10188 ( .A1(n8779), .A2(n10156), .ZN(n10270) );
  NAND2_X1 U10189 ( .A1(a_8_), .A2(n10266), .ZN(n10187) );
  NAND2_X1 U10190 ( .A1(n10271), .A2(n10272), .ZN(n10266) );
  INV_X1 U10191 ( .A(n10273), .ZN(n10272) );
  NOR3_X1 U10192 ( .A1(n8779), .A2(n10274), .A3(n8514), .ZN(n10273) );
  NOR2_X1 U10193 ( .A1(n10011), .A2(n10009), .ZN(n10274) );
  NAND2_X1 U10194 ( .A1(n10009), .A2(n10011), .ZN(n10271) );
  NAND2_X1 U10195 ( .A1(n10183), .A2(n10275), .ZN(n10011) );
  NAND2_X1 U10196 ( .A1(n10182), .A2(n10184), .ZN(n10275) );
  NAND2_X1 U10197 ( .A1(n10276), .A2(n10277), .ZN(n10184) );
  NAND2_X1 U10198 ( .A1(b_27_), .A2(a_10_), .ZN(n10277) );
  XNOR2_X1 U10199 ( .A(n10278), .B(n10279), .ZN(n10182) );
  XOR2_X1 U10200 ( .A(n10280), .B(n10281), .Z(n10279) );
  NAND2_X1 U10201 ( .A1(b_26_), .A2(a_11_), .ZN(n10281) );
  INV_X1 U10202 ( .A(n10282), .ZN(n10183) );
  NOR2_X1 U10203 ( .A1(n8769), .A2(n10276), .ZN(n10282) );
  NOR2_X1 U10204 ( .A1(n10283), .A2(n10284), .ZN(n10276) );
  NOR3_X1 U10205 ( .A1(n8749), .A2(n10285), .A3(n8514), .ZN(n10284) );
  NOR2_X1 U10206 ( .A1(n10022), .A2(n10021), .ZN(n10285) );
  INV_X1 U10207 ( .A(n10286), .ZN(n10283) );
  NAND2_X1 U10208 ( .A1(n10021), .A2(n10022), .ZN(n10286) );
  NAND2_X1 U10209 ( .A1(n10179), .A2(n10287), .ZN(n10022) );
  NAND2_X1 U10210 ( .A1(n10178), .A2(n10180), .ZN(n10287) );
  NAND2_X1 U10211 ( .A1(n10288), .A2(n10289), .ZN(n10180) );
  NAND2_X1 U10212 ( .A1(b_27_), .A2(a_12_), .ZN(n10289) );
  INV_X1 U10213 ( .A(n10290), .ZN(n10288) );
  XNOR2_X1 U10214 ( .A(n10291), .B(n10292), .ZN(n10178) );
  XOR2_X1 U10215 ( .A(n10293), .B(n10294), .Z(n10292) );
  NAND2_X1 U10216 ( .A1(b_26_), .A2(a_13_), .ZN(n10294) );
  NAND2_X1 U10217 ( .A1(a_12_), .A2(n10290), .ZN(n10179) );
  NAND2_X1 U10218 ( .A1(n10295), .A2(n10296), .ZN(n10290) );
  INV_X1 U10219 ( .A(n10297), .ZN(n10296) );
  NOR3_X1 U10220 ( .A1(n8721), .A2(n10298), .A3(n8514), .ZN(n10297) );
  NOR2_X1 U10221 ( .A1(n10035), .A2(n10033), .ZN(n10298) );
  NAND2_X1 U10222 ( .A1(n10033), .A2(n10035), .ZN(n10295) );
  NAND2_X1 U10223 ( .A1(n10175), .A2(n10299), .ZN(n10035) );
  NAND2_X1 U10224 ( .A1(n10174), .A2(n10176), .ZN(n10299) );
  NAND2_X1 U10225 ( .A1(n10300), .A2(n10301), .ZN(n10176) );
  NAND2_X1 U10226 ( .A1(b_27_), .A2(a_14_), .ZN(n10301) );
  XOR2_X1 U10227 ( .A(n10302), .B(n10303), .Z(n10174) );
  XOR2_X1 U10228 ( .A(n10304), .B(n10305), .Z(n10302) );
  NOR2_X1 U10229 ( .A1(n8692), .A2(n10156), .ZN(n10305) );
  INV_X1 U10230 ( .A(n10306), .ZN(n10175) );
  NOR2_X1 U10231 ( .A1(n8991), .A2(n10300), .ZN(n10306) );
  NOR2_X1 U10232 ( .A1(n10307), .A2(n10308), .ZN(n10300) );
  NOR3_X1 U10233 ( .A1(n8692), .A2(n10309), .A3(n8514), .ZN(n10308) );
  NOR2_X1 U10234 ( .A1(n10047), .A2(n10046), .ZN(n10309) );
  INV_X1 U10235 ( .A(n10310), .ZN(n10307) );
  NAND2_X1 U10236 ( .A1(n10046), .A2(n10047), .ZN(n10310) );
  NAND2_X1 U10237 ( .A1(n10171), .A2(n10311), .ZN(n10047) );
  NAND2_X1 U10238 ( .A1(n10170), .A2(n10172), .ZN(n10311) );
  NAND2_X1 U10239 ( .A1(n10312), .A2(n10313), .ZN(n10172) );
  NAND2_X1 U10240 ( .A1(b_27_), .A2(a_16_), .ZN(n10313) );
  INV_X1 U10241 ( .A(n10314), .ZN(n10312) );
  XNOR2_X1 U10242 ( .A(n10315), .B(n10316), .ZN(n10170) );
  XOR2_X1 U10243 ( .A(n10317), .B(n10318), .Z(n10316) );
  NAND2_X1 U10244 ( .A1(b_26_), .A2(a_17_), .ZN(n10318) );
  NAND2_X1 U10245 ( .A1(a_16_), .A2(n10314), .ZN(n10171) );
  NAND2_X1 U10246 ( .A1(n10319), .A2(n10320), .ZN(n10314) );
  NAND3_X1 U10247 ( .A1(a_17_), .A2(n10321), .A3(b_27_), .ZN(n10320) );
  NAND2_X1 U10248 ( .A1(n10056), .A2(n10058), .ZN(n10321) );
  INV_X1 U10249 ( .A(n10322), .ZN(n10319) );
  NOR2_X1 U10250 ( .A1(n10058), .A2(n10056), .ZN(n10322) );
  XOR2_X1 U10251 ( .A(n10323), .B(n10324), .Z(n10056) );
  XOR2_X1 U10252 ( .A(n10325), .B(n10326), .Z(n10323) );
  NAND2_X1 U10253 ( .A1(n10327), .A2(n10328), .ZN(n10058) );
  NAND2_X1 U10254 ( .A1(n10066), .A2(n10329), .ZN(n10328) );
  NAND2_X1 U10255 ( .A1(n10068), .A2(n10067), .ZN(n10329) );
  XNOR2_X1 U10256 ( .A(n10330), .B(n10331), .ZN(n10066) );
  XOR2_X1 U10257 ( .A(n10332), .B(n10333), .Z(n10330) );
  NOR2_X1 U10258 ( .A1(n8630), .A2(n10156), .ZN(n10333) );
  INV_X1 U10259 ( .A(n10334), .ZN(n10327) );
  NOR2_X1 U10260 ( .A1(n10067), .A2(n10068), .ZN(n10334) );
  NOR2_X1 U10261 ( .A1(n8514), .A2(n8988), .ZN(n10068) );
  NAND2_X1 U10262 ( .A1(n10335), .A2(n10336), .ZN(n10067) );
  NAND3_X1 U10263 ( .A1(a_19_), .A2(n10337), .A3(b_27_), .ZN(n10336) );
  INV_X1 U10264 ( .A(n10338), .ZN(n10337) );
  NOR2_X1 U10265 ( .A1(n10074), .A2(n10072), .ZN(n10338) );
  NAND2_X1 U10266 ( .A1(n10072), .A2(n10074), .ZN(n10335) );
  NAND2_X1 U10267 ( .A1(n10167), .A2(n10339), .ZN(n10074) );
  NAND2_X1 U10268 ( .A1(n10166), .A2(n10168), .ZN(n10339) );
  NAND2_X1 U10269 ( .A1(n10340), .A2(n10341), .ZN(n10168) );
  NAND2_X1 U10270 ( .A1(b_27_), .A2(a_20_), .ZN(n10341) );
  INV_X1 U10271 ( .A(n10342), .ZN(n10340) );
  XNOR2_X1 U10272 ( .A(n10343), .B(n10344), .ZN(n10166) );
  XOR2_X1 U10273 ( .A(n10345), .B(n10346), .Z(n10344) );
  NAND2_X1 U10274 ( .A1(b_26_), .A2(a_21_), .ZN(n10346) );
  NAND2_X1 U10275 ( .A1(a_20_), .A2(n10342), .ZN(n10167) );
  NAND2_X1 U10276 ( .A1(n10347), .A2(n10348), .ZN(n10342) );
  INV_X1 U10277 ( .A(n10349), .ZN(n10348) );
  NOR3_X1 U10278 ( .A1(n8601), .A2(n10350), .A3(n8514), .ZN(n10349) );
  NOR2_X1 U10279 ( .A1(n10087), .A2(n10085), .ZN(n10350) );
  NAND2_X1 U10280 ( .A1(n10085), .A2(n10087), .ZN(n10347) );
  NAND2_X1 U10281 ( .A1(n10163), .A2(n10351), .ZN(n10087) );
  NAND2_X1 U10282 ( .A1(n10162), .A2(n10164), .ZN(n10351) );
  NAND2_X1 U10283 ( .A1(n10352), .A2(n10353), .ZN(n10164) );
  NAND2_X1 U10284 ( .A1(b_27_), .A2(a_22_), .ZN(n10353) );
  INV_X1 U10285 ( .A(n10354), .ZN(n10352) );
  XNOR2_X1 U10286 ( .A(n10355), .B(n10356), .ZN(n10162) );
  NAND2_X1 U10287 ( .A1(n10357), .A2(n10358), .ZN(n10355) );
  NAND2_X1 U10288 ( .A1(a_22_), .A2(n10354), .ZN(n10163) );
  NAND2_X1 U10289 ( .A1(n10099), .A2(n10359), .ZN(n10354) );
  NAND2_X1 U10290 ( .A1(n10098), .A2(n10100), .ZN(n10359) );
  NAND2_X1 U10291 ( .A1(n10360), .A2(n10361), .ZN(n10100) );
  NAND2_X1 U10292 ( .A1(b_27_), .A2(a_23_), .ZN(n10361) );
  XOR2_X1 U10293 ( .A(n10362), .B(n10363), .Z(n10098) );
  XOR2_X1 U10294 ( .A(n10364), .B(n10365), .Z(n10362) );
  NAND2_X1 U10295 ( .A1(a_23_), .A2(n10366), .ZN(n10099) );
  INV_X1 U10296 ( .A(n10360), .ZN(n10366) );
  NOR2_X1 U10297 ( .A1(n10367), .A2(n10368), .ZN(n10360) );
  NOR2_X1 U10298 ( .A1(n10108), .A2(n10369), .ZN(n10368) );
  NOR2_X1 U10299 ( .A1(n10107), .A2(n10105), .ZN(n10369) );
  NAND2_X1 U10300 ( .A1(b_27_), .A2(a_24_), .ZN(n10108) );
  INV_X1 U10301 ( .A(n10370), .ZN(n10367) );
  NAND2_X1 U10302 ( .A1(n10105), .A2(n10107), .ZN(n10370) );
  NAND2_X1 U10303 ( .A1(n10159), .A2(n10371), .ZN(n10107) );
  NAND2_X1 U10304 ( .A1(n10158), .A2(n10160), .ZN(n10371) );
  NAND2_X1 U10305 ( .A1(n10372), .A2(n10373), .ZN(n10160) );
  NAND2_X1 U10306 ( .A1(b_27_), .A2(a_25_), .ZN(n10373) );
  INV_X1 U10307 ( .A(n10374), .ZN(n10372) );
  XOR2_X1 U10308 ( .A(n10375), .B(n10376), .Z(n10158) );
  XNOR2_X1 U10309 ( .A(n10377), .B(n8526), .ZN(n10376) );
  NAND2_X1 U10310 ( .A1(a_25_), .A2(n10374), .ZN(n10159) );
  NAND2_X1 U10311 ( .A1(n10120), .A2(n10378), .ZN(n10374) );
  NAND2_X1 U10312 ( .A1(n10119), .A2(n10121), .ZN(n10378) );
  NAND2_X1 U10313 ( .A1(n10379), .A2(n10380), .ZN(n10121) );
  NAND2_X1 U10314 ( .A1(b_27_), .A2(a_26_), .ZN(n10379) );
  XOR2_X1 U10315 ( .A(n10381), .B(n10382), .Z(n10119) );
  XOR2_X1 U10316 ( .A(n10383), .B(n10384), .Z(n10381) );
  NAND2_X1 U10317 ( .A1(n10385), .A2(a_26_), .ZN(n10120) );
  INV_X1 U10318 ( .A(n10380), .ZN(n10385) );
  NAND2_X1 U10319 ( .A1(n10386), .A2(n10387), .ZN(n10380) );
  NAND2_X1 U10320 ( .A1(n10127), .A2(n10388), .ZN(n10387) );
  NAND2_X1 U10321 ( .A1(n8509), .A2(n10128), .ZN(n10388) );
  XNOR2_X1 U10322 ( .A(n10389), .B(n10390), .ZN(n10127) );
  XOR2_X1 U10323 ( .A(n10391), .B(n10392), .Z(n10389) );
  INV_X1 U10324 ( .A(n10393), .ZN(n10386) );
  NOR2_X1 U10325 ( .A1(n10128), .A2(n8509), .ZN(n10393) );
  NOR2_X1 U10326 ( .A1(n8514), .A2(n8512), .ZN(n8509) );
  NAND2_X1 U10327 ( .A1(n10394), .A2(n10395), .ZN(n10128) );
  NAND2_X1 U10328 ( .A1(n10135), .A2(n10396), .ZN(n10395) );
  INV_X1 U10329 ( .A(n10397), .ZN(n10396) );
  NOR2_X1 U10330 ( .A1(n10136), .A2(n10134), .ZN(n10397) );
  NOR2_X1 U10331 ( .A1(n8514), .A2(n8493), .ZN(n10135) );
  NAND2_X1 U10332 ( .A1(n10134), .A2(n10136), .ZN(n10394) );
  NAND2_X1 U10333 ( .A1(n10398), .A2(n10399), .ZN(n10136) );
  NAND2_X1 U10334 ( .A1(n10142), .A2(n10400), .ZN(n10399) );
  INV_X1 U10335 ( .A(n10401), .ZN(n10400) );
  NOR2_X1 U10336 ( .A1(n10143), .A2(n10144), .ZN(n10401) );
  NOR2_X1 U10337 ( .A1(n8514), .A2(n8473), .ZN(n10142) );
  NAND2_X1 U10338 ( .A1(n10144), .A2(n10143), .ZN(n10398) );
  NAND2_X1 U10339 ( .A1(n10402), .A2(n10403), .ZN(n10143) );
  NAND2_X1 U10340 ( .A1(b_25_), .A2(n10404), .ZN(n10403) );
  NAND2_X1 U10341 ( .A1(n8456), .A2(n10405), .ZN(n10404) );
  NAND2_X1 U10342 ( .A1(a_31_), .A2(n10156), .ZN(n10405) );
  NAND2_X1 U10343 ( .A1(b_26_), .A2(n10406), .ZN(n10402) );
  NAND2_X1 U10344 ( .A1(n8459), .A2(n10407), .ZN(n10406) );
  NAND2_X1 U10345 ( .A1(a_30_), .A2(n8543), .ZN(n10407) );
  NOR3_X1 U10346 ( .A1(n10156), .A2(n8979), .A3(n8514), .ZN(n10144) );
  XOR2_X1 U10347 ( .A(n10408), .B(n10409), .Z(n10134) );
  XOR2_X1 U10348 ( .A(n10410), .B(n10411), .Z(n10408) );
  XNOR2_X1 U10349 ( .A(n10412), .B(n10413), .ZN(n10105) );
  XNOR2_X1 U10350 ( .A(n10414), .B(n10415), .ZN(n10413) );
  XNOR2_X1 U10351 ( .A(n10416), .B(n10417), .ZN(n10085) );
  NAND2_X1 U10352 ( .A1(n10418), .A2(n10419), .ZN(n10416) );
  XNOR2_X1 U10353 ( .A(n10420), .B(n10421), .ZN(n10072) );
  NAND2_X1 U10354 ( .A1(n10422), .A2(n10423), .ZN(n10420) );
  XNOR2_X1 U10355 ( .A(n10424), .B(n10425), .ZN(n10046) );
  NAND2_X1 U10356 ( .A1(n10426), .A2(n10427), .ZN(n10424) );
  XNOR2_X1 U10357 ( .A(n10428), .B(n10429), .ZN(n10033) );
  NAND2_X1 U10358 ( .A1(n10430), .A2(n10431), .ZN(n10428) );
  XNOR2_X1 U10359 ( .A(n10432), .B(n10433), .ZN(n10021) );
  NAND2_X1 U10360 ( .A1(n10434), .A2(n10435), .ZN(n10432) );
  XNOR2_X1 U10361 ( .A(n10436), .B(n10437), .ZN(n10009) );
  NAND2_X1 U10362 ( .A1(n10438), .A2(n10439), .ZN(n10436) );
  XNOR2_X1 U10363 ( .A(n10440), .B(n10441), .ZN(n9998) );
  XOR2_X1 U10364 ( .A(n10442), .B(n10443), .Z(n10441) );
  NAND2_X1 U10365 ( .A1(b_26_), .A2(a_8_), .ZN(n10443) );
  NAND2_X1 U10366 ( .A1(n10192), .A2(n10444), .ZN(n10255) );
  INV_X1 U10367 ( .A(n10189), .ZN(n10444) );
  XOR2_X1 U10368 ( .A(n10445), .B(n10446), .Z(n10189) );
  XOR2_X1 U10369 ( .A(n10447), .B(n10448), .Z(n10446) );
  NAND2_X1 U10370 ( .A1(b_26_), .A2(a_7_), .ZN(n10448) );
  NOR2_X1 U10371 ( .A1(n8514), .A2(n8994), .ZN(n10192) );
  INV_X1 U10372 ( .A(b_27_), .ZN(n8514) );
  XNOR2_X1 U10373 ( .A(n10449), .B(n10450), .ZN(n10194) );
  XNOR2_X1 U10374 ( .A(n10451), .B(n10452), .ZN(n10449) );
  XNOR2_X1 U10375 ( .A(n10453), .B(n10454), .ZN(n10198) );
  XNOR2_X1 U10376 ( .A(n10455), .B(n10456), .ZN(n10453) );
  NOR2_X1 U10377 ( .A1(n8848), .A2(n10156), .ZN(n10456) );
  XOR2_X1 U10378 ( .A(n10457), .B(n10458), .Z(n10202) );
  XNOR2_X1 U10379 ( .A(n10459), .B(n10460), .ZN(n10458) );
  NAND2_X1 U10380 ( .A1(b_26_), .A2(a_4_), .ZN(n10460) );
  XNOR2_X1 U10381 ( .A(n10461), .B(n10462), .ZN(n10210) );
  NAND2_X1 U10382 ( .A1(n10463), .A2(n10464), .ZN(n10461) );
  NAND4_X1 U10383 ( .A1(n9202), .A2(n9201), .A3(n9203), .A4(n9197), .ZN(n9042)
         );
  INV_X1 U10384 ( .A(n10465), .ZN(n9197) );
  NAND2_X1 U10385 ( .A1(n10221), .A2(n10466), .ZN(n9203) );
  NAND2_X1 U10386 ( .A1(n10220), .A2(n10222), .ZN(n10466) );
  NAND2_X1 U10387 ( .A1(n10467), .A2(n10468), .ZN(n10222) );
  NAND2_X1 U10388 ( .A1(b_26_), .A2(a_0_), .ZN(n10467) );
  XNOR2_X1 U10389 ( .A(n10469), .B(n10470), .ZN(n10220) );
  XNOR2_X1 U10390 ( .A(n10471), .B(n10472), .ZN(n10469) );
  NOR2_X1 U10391 ( .A1(n9731), .A2(n8543), .ZN(n10472) );
  INV_X1 U10392 ( .A(n10473), .ZN(n10221) );
  NOR2_X1 U10393 ( .A1(n10468), .A2(n9471), .ZN(n10473) );
  NAND2_X1 U10394 ( .A1(n10474), .A2(n10475), .ZN(n10468) );
  NAND2_X1 U10395 ( .A1(n10227), .A2(n10476), .ZN(n10475) );
  NAND2_X1 U10396 ( .A1(n10229), .A2(n10228), .ZN(n10476) );
  XOR2_X1 U10397 ( .A(n10477), .B(n10478), .Z(n10227) );
  XNOR2_X1 U10398 ( .A(n10479), .B(n10480), .ZN(n10477) );
  NOR2_X1 U10399 ( .A1(n8998), .A2(n8543), .ZN(n10480) );
  INV_X1 U10400 ( .A(n10481), .ZN(n10474) );
  NOR2_X1 U10401 ( .A1(n10228), .A2(n10229), .ZN(n10481) );
  NOR2_X1 U10402 ( .A1(n10156), .A2(n9731), .ZN(n10229) );
  NAND2_X1 U10403 ( .A1(n10463), .A2(n10482), .ZN(n10228) );
  NAND2_X1 U10404 ( .A1(n10462), .A2(n10464), .ZN(n10482) );
  NAND2_X1 U10405 ( .A1(n10483), .A2(n10484), .ZN(n10464) );
  NAND2_X1 U10406 ( .A1(b_26_), .A2(a_2_), .ZN(n10484) );
  XOR2_X1 U10407 ( .A(n10485), .B(n10486), .Z(n10462) );
  XOR2_X1 U10408 ( .A(n10487), .B(n10488), .Z(n10485) );
  NOR2_X1 U10409 ( .A1(n8877), .A2(n8543), .ZN(n10488) );
  NAND2_X1 U10410 ( .A1(a_2_), .A2(n10489), .ZN(n10463) );
  INV_X1 U10411 ( .A(n10483), .ZN(n10489) );
  NOR2_X1 U10412 ( .A1(n10490), .A2(n10491), .ZN(n10483) );
  NOR3_X1 U10413 ( .A1(n8877), .A2(n10492), .A3(n10156), .ZN(n10491) );
  INV_X1 U10414 ( .A(n10493), .ZN(n10492) );
  NAND2_X1 U10415 ( .A1(n10241), .A2(n10240), .ZN(n10493) );
  NOR2_X1 U10416 ( .A1(n10240), .A2(n10241), .ZN(n10490) );
  NOR2_X1 U10417 ( .A1(n10494), .A2(n10495), .ZN(n10241) );
  NOR3_X1 U10418 ( .A1(n8996), .A2(n10496), .A3(n10156), .ZN(n10495) );
  INV_X1 U10419 ( .A(n10497), .ZN(n10496) );
  NAND2_X1 U10420 ( .A1(n10459), .A2(n10457), .ZN(n10497) );
  NOR2_X1 U10421 ( .A1(n10457), .A2(n10459), .ZN(n10494) );
  NOR2_X1 U10422 ( .A1(n10498), .A2(n10499), .ZN(n10459) );
  INV_X1 U10423 ( .A(n10500), .ZN(n10499) );
  NAND3_X1 U10424 ( .A1(a_5_), .A2(n10501), .A3(b_26_), .ZN(n10500) );
  NAND2_X1 U10425 ( .A1(n10455), .A2(n10454), .ZN(n10501) );
  NOR2_X1 U10426 ( .A1(n10454), .A2(n10455), .ZN(n10498) );
  NOR2_X1 U10427 ( .A1(n10502), .A2(n10503), .ZN(n10455) );
  INV_X1 U10428 ( .A(n10504), .ZN(n10503) );
  NAND2_X1 U10429 ( .A1(n10451), .A2(n10505), .ZN(n10504) );
  NAND2_X1 U10430 ( .A1(n10450), .A2(n10452), .ZN(n10505) );
  NAND2_X1 U10431 ( .A1(n10506), .A2(n10507), .ZN(n10451) );
  INV_X1 U10432 ( .A(n10508), .ZN(n10507) );
  NOR3_X1 U10433 ( .A1(n8817), .A2(n10509), .A3(n10156), .ZN(n10508) );
  NOR2_X1 U10434 ( .A1(n10447), .A2(n10445), .ZN(n10509) );
  NAND2_X1 U10435 ( .A1(n10445), .A2(n10447), .ZN(n10506) );
  NAND2_X1 U10436 ( .A1(n10510), .A2(n10511), .ZN(n10447) );
  INV_X1 U10437 ( .A(n10512), .ZN(n10511) );
  NOR3_X1 U10438 ( .A1(n10513), .A2(n10514), .A3(n10156), .ZN(n10512) );
  NOR2_X1 U10439 ( .A1(n10442), .A2(n10440), .ZN(n10514) );
  NAND2_X1 U10440 ( .A1(n10440), .A2(n10442), .ZN(n10510) );
  NAND2_X1 U10441 ( .A1(n10515), .A2(n10516), .ZN(n10442) );
  NAND3_X1 U10442 ( .A1(a_9_), .A2(n10517), .A3(b_26_), .ZN(n10516) );
  INV_X1 U10443 ( .A(n10518), .ZN(n10517) );
  NOR2_X1 U10444 ( .A1(n10269), .A2(n10268), .ZN(n10518) );
  NAND2_X1 U10445 ( .A1(n10268), .A2(n10269), .ZN(n10515) );
  NAND2_X1 U10446 ( .A1(n10438), .A2(n10519), .ZN(n10269) );
  NAND2_X1 U10447 ( .A1(n10437), .A2(n10439), .ZN(n10519) );
  NAND2_X1 U10448 ( .A1(n10520), .A2(n10521), .ZN(n10439) );
  NAND2_X1 U10449 ( .A1(b_26_), .A2(a_10_), .ZN(n10521) );
  INV_X1 U10450 ( .A(n10522), .ZN(n10520) );
  XOR2_X1 U10451 ( .A(n10523), .B(n10524), .Z(n10437) );
  XOR2_X1 U10452 ( .A(n10525), .B(n10526), .Z(n10523) );
  NOR2_X1 U10453 ( .A1(n8749), .A2(n8543), .ZN(n10526) );
  NAND2_X1 U10454 ( .A1(a_10_), .A2(n10522), .ZN(n10438) );
  NAND2_X1 U10455 ( .A1(n10527), .A2(n10528), .ZN(n10522) );
  INV_X1 U10456 ( .A(n10529), .ZN(n10528) );
  NOR3_X1 U10457 ( .A1(n8749), .A2(n10530), .A3(n10156), .ZN(n10529) );
  NOR2_X1 U10458 ( .A1(n10280), .A2(n10278), .ZN(n10530) );
  NAND2_X1 U10459 ( .A1(n10278), .A2(n10280), .ZN(n10527) );
  NAND2_X1 U10460 ( .A1(n10434), .A2(n10531), .ZN(n10280) );
  NAND2_X1 U10461 ( .A1(n10433), .A2(n10435), .ZN(n10531) );
  NAND2_X1 U10462 ( .A1(n10532), .A2(n10533), .ZN(n10435) );
  NAND2_X1 U10463 ( .A1(b_26_), .A2(a_12_), .ZN(n10533) );
  INV_X1 U10464 ( .A(n10534), .ZN(n10532) );
  XOR2_X1 U10465 ( .A(n10535), .B(n10536), .Z(n10433) );
  XOR2_X1 U10466 ( .A(n10537), .B(n10538), .Z(n10535) );
  NOR2_X1 U10467 ( .A1(n8721), .A2(n8543), .ZN(n10538) );
  NAND2_X1 U10468 ( .A1(a_12_), .A2(n10534), .ZN(n10434) );
  NAND2_X1 U10469 ( .A1(n10539), .A2(n10540), .ZN(n10534) );
  INV_X1 U10470 ( .A(n10541), .ZN(n10540) );
  NOR3_X1 U10471 ( .A1(n8721), .A2(n10542), .A3(n10156), .ZN(n10541) );
  NOR2_X1 U10472 ( .A1(n10293), .A2(n10291), .ZN(n10542) );
  NAND2_X1 U10473 ( .A1(n10291), .A2(n10293), .ZN(n10539) );
  NAND2_X1 U10474 ( .A1(n10430), .A2(n10543), .ZN(n10293) );
  NAND2_X1 U10475 ( .A1(n10429), .A2(n10431), .ZN(n10543) );
  NAND2_X1 U10476 ( .A1(n10544), .A2(n10545), .ZN(n10431) );
  NAND2_X1 U10477 ( .A1(b_26_), .A2(a_14_), .ZN(n10545) );
  XOR2_X1 U10478 ( .A(n10546), .B(n10547), .Z(n10429) );
  XOR2_X1 U10479 ( .A(n10548), .B(n10549), .Z(n10546) );
  NOR2_X1 U10480 ( .A1(n8692), .A2(n8543), .ZN(n10549) );
  INV_X1 U10481 ( .A(n10550), .ZN(n10430) );
  NOR2_X1 U10482 ( .A1(n8991), .A2(n10544), .ZN(n10550) );
  NOR2_X1 U10483 ( .A1(n10551), .A2(n10552), .ZN(n10544) );
  NOR3_X1 U10484 ( .A1(n8692), .A2(n10553), .A3(n10156), .ZN(n10552) );
  NOR2_X1 U10485 ( .A1(n10304), .A2(n10303), .ZN(n10553) );
  INV_X1 U10486 ( .A(n10554), .ZN(n10551) );
  NAND2_X1 U10487 ( .A1(n10303), .A2(n10304), .ZN(n10554) );
  NAND2_X1 U10488 ( .A1(n10426), .A2(n10555), .ZN(n10304) );
  NAND2_X1 U10489 ( .A1(n10425), .A2(n10427), .ZN(n10555) );
  NAND2_X1 U10490 ( .A1(n10556), .A2(n10557), .ZN(n10427) );
  NAND2_X1 U10491 ( .A1(b_26_), .A2(a_16_), .ZN(n10557) );
  XNOR2_X1 U10492 ( .A(n10558), .B(n10559), .ZN(n10425) );
  XOR2_X1 U10493 ( .A(n10560), .B(n10561), .Z(n10559) );
  NAND2_X1 U10494 ( .A1(b_25_), .A2(a_17_), .ZN(n10561) );
  INV_X1 U10495 ( .A(n10562), .ZN(n10426) );
  NOR2_X1 U10496 ( .A1(n8680), .A2(n10556), .ZN(n10562) );
  NOR2_X1 U10497 ( .A1(n10563), .A2(n10564), .ZN(n10556) );
  NOR3_X1 U10498 ( .A1(n8662), .A2(n10565), .A3(n10156), .ZN(n10564) );
  INV_X1 U10499 ( .A(n10566), .ZN(n10565) );
  NAND2_X1 U10500 ( .A1(n10315), .A2(n10317), .ZN(n10566) );
  NOR2_X1 U10501 ( .A1(n10317), .A2(n10315), .ZN(n10563) );
  XOR2_X1 U10502 ( .A(n10567), .B(n10568), .Z(n10315) );
  XOR2_X1 U10503 ( .A(n10569), .B(n10570), .Z(n10567) );
  NAND2_X1 U10504 ( .A1(n10571), .A2(n10572), .ZN(n10317) );
  NAND2_X1 U10505 ( .A1(n10324), .A2(n10573), .ZN(n10572) );
  NAND2_X1 U10506 ( .A1(n10326), .A2(n10325), .ZN(n10573) );
  XNOR2_X1 U10507 ( .A(n10574), .B(n10575), .ZN(n10324) );
  XOR2_X1 U10508 ( .A(n10576), .B(n10577), .Z(n10574) );
  NOR2_X1 U10509 ( .A1(n8630), .A2(n8543), .ZN(n10577) );
  INV_X1 U10510 ( .A(n10578), .ZN(n10571) );
  NOR2_X1 U10511 ( .A1(n10325), .A2(n10326), .ZN(n10578) );
  NOR2_X1 U10512 ( .A1(n10156), .A2(n8988), .ZN(n10326) );
  NAND2_X1 U10513 ( .A1(n10579), .A2(n10580), .ZN(n10325) );
  NAND3_X1 U10514 ( .A1(a_19_), .A2(n10581), .A3(b_26_), .ZN(n10580) );
  INV_X1 U10515 ( .A(n10582), .ZN(n10581) );
  NOR2_X1 U10516 ( .A1(n10332), .A2(n10331), .ZN(n10582) );
  NAND2_X1 U10517 ( .A1(n10331), .A2(n10332), .ZN(n10579) );
  NAND2_X1 U10518 ( .A1(n10422), .A2(n10583), .ZN(n10332) );
  NAND2_X1 U10519 ( .A1(n10421), .A2(n10423), .ZN(n10583) );
  NAND2_X1 U10520 ( .A1(n10584), .A2(n10585), .ZN(n10423) );
  NAND2_X1 U10521 ( .A1(b_26_), .A2(a_20_), .ZN(n10585) );
  INV_X1 U10522 ( .A(n10586), .ZN(n10584) );
  XNOR2_X1 U10523 ( .A(n10587), .B(n10588), .ZN(n10421) );
  XOR2_X1 U10524 ( .A(n10589), .B(n10590), .Z(n10588) );
  NAND2_X1 U10525 ( .A1(b_25_), .A2(a_21_), .ZN(n10590) );
  NAND2_X1 U10526 ( .A1(a_20_), .A2(n10586), .ZN(n10422) );
  NAND2_X1 U10527 ( .A1(n10591), .A2(n10592), .ZN(n10586) );
  INV_X1 U10528 ( .A(n10593), .ZN(n10592) );
  NOR3_X1 U10529 ( .A1(n8601), .A2(n10594), .A3(n10156), .ZN(n10593) );
  NOR2_X1 U10530 ( .A1(n10345), .A2(n10343), .ZN(n10594) );
  NAND2_X1 U10531 ( .A1(n10343), .A2(n10345), .ZN(n10591) );
  NAND2_X1 U10532 ( .A1(n10418), .A2(n10595), .ZN(n10345) );
  NAND2_X1 U10533 ( .A1(n10417), .A2(n10419), .ZN(n10595) );
  NAND2_X1 U10534 ( .A1(n10596), .A2(n10597), .ZN(n10419) );
  NAND2_X1 U10535 ( .A1(b_26_), .A2(a_22_), .ZN(n10597) );
  INV_X1 U10536 ( .A(n10598), .ZN(n10596) );
  XNOR2_X1 U10537 ( .A(n10599), .B(n10600), .ZN(n10417) );
  NAND2_X1 U10538 ( .A1(n10601), .A2(n10602), .ZN(n10599) );
  NAND2_X1 U10539 ( .A1(a_22_), .A2(n10598), .ZN(n10418) );
  NAND2_X1 U10540 ( .A1(n10357), .A2(n10603), .ZN(n10598) );
  NAND2_X1 U10541 ( .A1(n10356), .A2(n10358), .ZN(n10603) );
  NAND2_X1 U10542 ( .A1(n10604), .A2(n10605), .ZN(n10358) );
  NAND2_X1 U10543 ( .A1(b_26_), .A2(a_23_), .ZN(n10605) );
  INV_X1 U10544 ( .A(n10606), .ZN(n10604) );
  XNOR2_X1 U10545 ( .A(n10607), .B(n10608), .ZN(n10356) );
  XNOR2_X1 U10546 ( .A(n10609), .B(n10610), .ZN(n10608) );
  NAND2_X1 U10547 ( .A1(a_23_), .A2(n10606), .ZN(n10357) );
  NAND2_X1 U10548 ( .A1(n10611), .A2(n10612), .ZN(n10606) );
  NAND2_X1 U10549 ( .A1(n10365), .A2(n10613), .ZN(n10612) );
  INV_X1 U10550 ( .A(n10614), .ZN(n10613) );
  NOR2_X1 U10551 ( .A1(n10364), .A2(n10363), .ZN(n10614) );
  NOR2_X1 U10552 ( .A1(n10156), .A2(n8982), .ZN(n10365) );
  NAND2_X1 U10553 ( .A1(n10363), .A2(n10364), .ZN(n10611) );
  NAND2_X1 U10554 ( .A1(n10615), .A2(n10616), .ZN(n10364) );
  NAND2_X1 U10555 ( .A1(n10415), .A2(n10617), .ZN(n10616) );
  NAND2_X1 U10556 ( .A1(n10412), .A2(n10414), .ZN(n10617) );
  NOR2_X1 U10557 ( .A1(n10156), .A2(n8541), .ZN(n10415) );
  INV_X1 U10558 ( .A(n10618), .ZN(n10615) );
  NOR2_X1 U10559 ( .A1(n10414), .A2(n10412), .ZN(n10618) );
  XNOR2_X1 U10560 ( .A(n10619), .B(n10620), .ZN(n10412) );
  XNOR2_X1 U10561 ( .A(n10621), .B(n10622), .ZN(n10620) );
  NAND2_X1 U10562 ( .A1(n10623), .A2(n10624), .ZN(n10414) );
  NAND2_X1 U10563 ( .A1(n10375), .A2(n10625), .ZN(n10624) );
  NAND2_X1 U10564 ( .A1(n8526), .A2(n10377), .ZN(n10625) );
  XNOR2_X1 U10565 ( .A(n10626), .B(n10627), .ZN(n10375) );
  XOR2_X1 U10566 ( .A(n10628), .B(n10629), .Z(n10626) );
  INV_X1 U10567 ( .A(n10630), .ZN(n10623) );
  NOR2_X1 U10568 ( .A1(n10377), .A2(n8526), .ZN(n10630) );
  NOR2_X1 U10569 ( .A1(n10156), .A2(n9893), .ZN(n8526) );
  NAND2_X1 U10570 ( .A1(n10631), .A2(n10632), .ZN(n10377) );
  NAND2_X1 U10571 ( .A1(n10384), .A2(n10633), .ZN(n10632) );
  INV_X1 U10572 ( .A(n10634), .ZN(n10633) );
  NOR2_X1 U10573 ( .A1(n10383), .A2(n10382), .ZN(n10634) );
  NOR2_X1 U10574 ( .A1(n10156), .A2(n8512), .ZN(n10384) );
  NAND2_X1 U10575 ( .A1(n10382), .A2(n10383), .ZN(n10631) );
  NAND2_X1 U10576 ( .A1(n10635), .A2(n10636), .ZN(n10383) );
  NAND2_X1 U10577 ( .A1(n10391), .A2(n10637), .ZN(n10636) );
  INV_X1 U10578 ( .A(n10638), .ZN(n10637) );
  NOR2_X1 U10579 ( .A1(n10392), .A2(n10390), .ZN(n10638) );
  NOR2_X1 U10580 ( .A1(n10156), .A2(n8493), .ZN(n10391) );
  NAND2_X1 U10581 ( .A1(n10390), .A2(n10392), .ZN(n10635) );
  NAND2_X1 U10582 ( .A1(n10639), .A2(n10640), .ZN(n10392) );
  NAND2_X1 U10583 ( .A1(n10409), .A2(n10641), .ZN(n10640) );
  INV_X1 U10584 ( .A(n10642), .ZN(n10641) );
  NOR2_X1 U10585 ( .A1(n10410), .A2(n10411), .ZN(n10642) );
  NOR2_X1 U10586 ( .A1(n10156), .A2(n8473), .ZN(n10409) );
  NAND2_X1 U10587 ( .A1(n10411), .A2(n10410), .ZN(n10639) );
  NAND2_X1 U10588 ( .A1(n10643), .A2(n10644), .ZN(n10410) );
  NAND2_X1 U10589 ( .A1(b_24_), .A2(n10645), .ZN(n10644) );
  NAND2_X1 U10590 ( .A1(n8456), .A2(n10646), .ZN(n10645) );
  NAND2_X1 U10591 ( .A1(a_31_), .A2(n8543), .ZN(n10646) );
  NAND2_X1 U10592 ( .A1(b_25_), .A2(n10647), .ZN(n10643) );
  NAND2_X1 U10593 ( .A1(n8459), .A2(n10648), .ZN(n10647) );
  NAND2_X1 U10594 ( .A1(a_30_), .A2(n8981), .ZN(n10648) );
  NOR3_X1 U10595 ( .A1(n8543), .A2(n8979), .A3(n10156), .ZN(n10411) );
  XOR2_X1 U10596 ( .A(n10649), .B(n10650), .Z(n10390) );
  XOR2_X1 U10597 ( .A(n10651), .B(n10652), .Z(n10649) );
  XOR2_X1 U10598 ( .A(n10653), .B(n10654), .Z(n10382) );
  XOR2_X1 U10599 ( .A(n10655), .B(n10656), .Z(n10653) );
  XNOR2_X1 U10600 ( .A(n10657), .B(n10658), .ZN(n10363) );
  XNOR2_X1 U10601 ( .A(n10659), .B(n8965), .ZN(n10658) );
  XNOR2_X1 U10602 ( .A(n10660), .B(n10661), .ZN(n10343) );
  NAND2_X1 U10603 ( .A1(n10662), .A2(n10663), .ZN(n10660) );
  XNOR2_X1 U10604 ( .A(n10664), .B(n10665), .ZN(n10331) );
  NAND2_X1 U10605 ( .A1(n10666), .A2(n10667), .ZN(n10664) );
  XNOR2_X1 U10606 ( .A(n10668), .B(n10669), .ZN(n10303) );
  NAND2_X1 U10607 ( .A1(n10670), .A2(n10671), .ZN(n10668) );
  XNOR2_X1 U10608 ( .A(n10672), .B(n10673), .ZN(n10291) );
  NAND2_X1 U10609 ( .A1(n10674), .A2(n10675), .ZN(n10672) );
  XNOR2_X1 U10610 ( .A(n10676), .B(n10677), .ZN(n10278) );
  NAND2_X1 U10611 ( .A1(n10678), .A2(n10679), .ZN(n10676) );
  XOR2_X1 U10612 ( .A(n10680), .B(n10681), .Z(n10268) );
  XNOR2_X1 U10613 ( .A(n10682), .B(n10683), .ZN(n10681) );
  XOR2_X1 U10614 ( .A(n10684), .B(n10685), .Z(n10440) );
  XOR2_X1 U10615 ( .A(n10686), .B(n10687), .Z(n10684) );
  NOR2_X1 U10616 ( .A1(n8779), .A2(n8543), .ZN(n10687) );
  XNOR2_X1 U10617 ( .A(n10688), .B(n10689), .ZN(n10445) );
  XNOR2_X1 U10618 ( .A(n10690), .B(n10691), .ZN(n10688) );
  NOR2_X1 U10619 ( .A1(n10513), .A2(n8543), .ZN(n10691) );
  NOR2_X1 U10620 ( .A1(n10452), .A2(n10450), .ZN(n10502) );
  XNOR2_X1 U10621 ( .A(n10692), .B(n10693), .ZN(n10450) );
  XNOR2_X1 U10622 ( .A(n10694), .B(n10695), .ZN(n10693) );
  NAND2_X1 U10623 ( .A1(b_25_), .A2(a_7_), .ZN(n10695) );
  NAND2_X1 U10624 ( .A1(b_26_), .A2(a_6_), .ZN(n10452) );
  XOR2_X1 U10625 ( .A(n10696), .B(n10697), .Z(n10454) );
  NAND2_X1 U10626 ( .A1(n10698), .A2(n10699), .ZN(n10696) );
  XOR2_X1 U10627 ( .A(n10700), .B(n10701), .Z(n10457) );
  XOR2_X1 U10628 ( .A(n10702), .B(n10703), .Z(n10701) );
  NAND2_X1 U10629 ( .A1(b_25_), .A2(a_5_), .ZN(n10703) );
  XOR2_X1 U10630 ( .A(n10704), .B(n10705), .Z(n10240) );
  XOR2_X1 U10631 ( .A(n10706), .B(n10707), .Z(n10705) );
  NAND2_X1 U10632 ( .A1(b_25_), .A2(a_4_), .ZN(n10707) );
  NAND2_X1 U10633 ( .A1(n10708), .A2(n10709), .ZN(n9201) );
  XOR2_X1 U10634 ( .A(n10710), .B(n10711), .Z(n9202) );
  XNOR2_X1 U10635 ( .A(n10712), .B(n10713), .ZN(n10711) );
  NAND2_X1 U10636 ( .A1(b_25_), .A2(a_0_), .ZN(n10713) );
  NAND2_X1 U10637 ( .A1(n10465), .A2(n10714), .ZN(n9047) );
  XOR2_X1 U10638 ( .A(n9194), .B(n9193), .Z(n10714) );
  NOR2_X1 U10639 ( .A1(n10709), .A2(n10708), .ZN(n10465) );
  NOR2_X1 U10640 ( .A1(n10715), .A2(n10716), .ZN(n10708) );
  NOR3_X1 U10641 ( .A1(n9471), .A2(n10717), .A3(n8543), .ZN(n10716) );
  INV_X1 U10642 ( .A(n10718), .ZN(n10717) );
  NAND2_X1 U10643 ( .A1(n10712), .A2(n10710), .ZN(n10718) );
  NOR2_X1 U10644 ( .A1(n10710), .A2(n10712), .ZN(n10715) );
  NOR2_X1 U10645 ( .A1(n10719), .A2(n10720), .ZN(n10712) );
  INV_X1 U10646 ( .A(n10721), .ZN(n10720) );
  NAND3_X1 U10647 ( .A1(a_1_), .A2(n10722), .A3(b_25_), .ZN(n10721) );
  NAND2_X1 U10648 ( .A1(n10471), .A2(n10470), .ZN(n10722) );
  NOR2_X1 U10649 ( .A1(n10470), .A2(n10471), .ZN(n10719) );
  NOR2_X1 U10650 ( .A1(n10723), .A2(n10724), .ZN(n10471) );
  INV_X1 U10651 ( .A(n10725), .ZN(n10724) );
  NAND3_X1 U10652 ( .A1(a_2_), .A2(n10726), .A3(b_25_), .ZN(n10725) );
  NAND2_X1 U10653 ( .A1(n10479), .A2(n10478), .ZN(n10726) );
  NOR2_X1 U10654 ( .A1(n10478), .A2(n10479), .ZN(n10723) );
  NOR2_X1 U10655 ( .A1(n10727), .A2(n10728), .ZN(n10479) );
  NOR3_X1 U10656 ( .A1(n8877), .A2(n10729), .A3(n8543), .ZN(n10728) );
  NOR2_X1 U10657 ( .A1(n10487), .A2(n10486), .ZN(n10729) );
  INV_X1 U10658 ( .A(n10730), .ZN(n10727) );
  NAND2_X1 U10659 ( .A1(n10486), .A2(n10487), .ZN(n10730) );
  NAND2_X1 U10660 ( .A1(n10731), .A2(n10732), .ZN(n10487) );
  NAND3_X1 U10661 ( .A1(a_4_), .A2(n10733), .A3(b_25_), .ZN(n10732) );
  INV_X1 U10662 ( .A(n10734), .ZN(n10733) );
  NOR2_X1 U10663 ( .A1(n10706), .A2(n10704), .ZN(n10734) );
  NAND2_X1 U10664 ( .A1(n10704), .A2(n10706), .ZN(n10731) );
  NAND2_X1 U10665 ( .A1(n10735), .A2(n10736), .ZN(n10706) );
  NAND3_X1 U10666 ( .A1(a_5_), .A2(n10737), .A3(b_25_), .ZN(n10736) );
  INV_X1 U10667 ( .A(n10738), .ZN(n10737) );
  NOR2_X1 U10668 ( .A1(n10702), .A2(n10700), .ZN(n10738) );
  NAND2_X1 U10669 ( .A1(n10700), .A2(n10702), .ZN(n10735) );
  NAND2_X1 U10670 ( .A1(n10698), .A2(n10739), .ZN(n10702) );
  NAND2_X1 U10671 ( .A1(n10697), .A2(n10699), .ZN(n10739) );
  NAND2_X1 U10672 ( .A1(n10740), .A2(n10741), .ZN(n10699) );
  NAND2_X1 U10673 ( .A1(b_25_), .A2(a_6_), .ZN(n10741) );
  XNOR2_X1 U10674 ( .A(n10742), .B(n10743), .ZN(n10697) );
  NAND2_X1 U10675 ( .A1(n10744), .A2(n10745), .ZN(n10742) );
  INV_X1 U10676 ( .A(n10746), .ZN(n10698) );
  NOR2_X1 U10677 ( .A1(n8994), .A2(n10740), .ZN(n10746) );
  NOR2_X1 U10678 ( .A1(n10747), .A2(n10748), .ZN(n10740) );
  INV_X1 U10679 ( .A(n10749), .ZN(n10748) );
  NAND3_X1 U10680 ( .A1(a_7_), .A2(n10750), .A3(b_25_), .ZN(n10749) );
  NAND2_X1 U10681 ( .A1(n10694), .A2(n10692), .ZN(n10750) );
  NOR2_X1 U10682 ( .A1(n10692), .A2(n10694), .ZN(n10747) );
  NOR2_X1 U10683 ( .A1(n10751), .A2(n10752), .ZN(n10694) );
  INV_X1 U10684 ( .A(n10753), .ZN(n10752) );
  NAND3_X1 U10685 ( .A1(a_8_), .A2(n10754), .A3(b_25_), .ZN(n10753) );
  NAND2_X1 U10686 ( .A1(n10690), .A2(n10689), .ZN(n10754) );
  NOR2_X1 U10687 ( .A1(n10689), .A2(n10690), .ZN(n10751) );
  NOR2_X1 U10688 ( .A1(n10755), .A2(n10756), .ZN(n10690) );
  NOR3_X1 U10689 ( .A1(n8779), .A2(n10757), .A3(n8543), .ZN(n10756) );
  NOR2_X1 U10690 ( .A1(n10686), .A2(n10685), .ZN(n10757) );
  INV_X1 U10691 ( .A(n10758), .ZN(n10755) );
  NAND2_X1 U10692 ( .A1(n10685), .A2(n10686), .ZN(n10758) );
  NAND2_X1 U10693 ( .A1(n10759), .A2(n10760), .ZN(n10686) );
  NAND2_X1 U10694 ( .A1(n10682), .A2(n10761), .ZN(n10760) );
  NAND2_X1 U10695 ( .A1(n10680), .A2(n10762), .ZN(n10761) );
  INV_X1 U10696 ( .A(n10683), .ZN(n10762) );
  NAND2_X1 U10697 ( .A1(n10763), .A2(n10764), .ZN(n10682) );
  INV_X1 U10698 ( .A(n10765), .ZN(n10764) );
  NOR3_X1 U10699 ( .A1(n8749), .A2(n10766), .A3(n8543), .ZN(n10765) );
  NOR2_X1 U10700 ( .A1(n10525), .A2(n10524), .ZN(n10766) );
  NAND2_X1 U10701 ( .A1(n10524), .A2(n10525), .ZN(n10763) );
  NAND2_X1 U10702 ( .A1(n10678), .A2(n10767), .ZN(n10525) );
  NAND2_X1 U10703 ( .A1(n10677), .A2(n10679), .ZN(n10767) );
  NAND2_X1 U10704 ( .A1(n10768), .A2(n10769), .ZN(n10679) );
  NAND2_X1 U10705 ( .A1(b_25_), .A2(a_12_), .ZN(n10769) );
  INV_X1 U10706 ( .A(n10770), .ZN(n10768) );
  XOR2_X1 U10707 ( .A(n10771), .B(n10772), .Z(n10677) );
  XOR2_X1 U10708 ( .A(n10773), .B(n10774), .Z(n10771) );
  NOR2_X1 U10709 ( .A1(n8721), .A2(n8981), .ZN(n10774) );
  NAND2_X1 U10710 ( .A1(a_12_), .A2(n10770), .ZN(n10678) );
  NAND2_X1 U10711 ( .A1(n10775), .A2(n10776), .ZN(n10770) );
  INV_X1 U10712 ( .A(n10777), .ZN(n10776) );
  NOR3_X1 U10713 ( .A1(n8721), .A2(n10778), .A3(n8543), .ZN(n10777) );
  NOR2_X1 U10714 ( .A1(n10537), .A2(n10536), .ZN(n10778) );
  NAND2_X1 U10715 ( .A1(n10536), .A2(n10537), .ZN(n10775) );
  NAND2_X1 U10716 ( .A1(n10674), .A2(n10779), .ZN(n10537) );
  NAND2_X1 U10717 ( .A1(n10673), .A2(n10675), .ZN(n10779) );
  NAND2_X1 U10718 ( .A1(n10780), .A2(n10781), .ZN(n10675) );
  NAND2_X1 U10719 ( .A1(b_25_), .A2(a_14_), .ZN(n10781) );
  INV_X1 U10720 ( .A(n10782), .ZN(n10780) );
  XOR2_X1 U10721 ( .A(n10783), .B(n10784), .Z(n10673) );
  XOR2_X1 U10722 ( .A(n10785), .B(n10786), .Z(n10783) );
  NOR2_X1 U10723 ( .A1(n8692), .A2(n8981), .ZN(n10786) );
  NAND2_X1 U10724 ( .A1(a_14_), .A2(n10782), .ZN(n10674) );
  NAND2_X1 U10725 ( .A1(n10787), .A2(n10788), .ZN(n10782) );
  INV_X1 U10726 ( .A(n10789), .ZN(n10788) );
  NOR3_X1 U10727 ( .A1(n8692), .A2(n10790), .A3(n8543), .ZN(n10789) );
  NOR2_X1 U10728 ( .A1(n10548), .A2(n10547), .ZN(n10790) );
  NAND2_X1 U10729 ( .A1(n10547), .A2(n10548), .ZN(n10787) );
  NAND2_X1 U10730 ( .A1(n10670), .A2(n10791), .ZN(n10548) );
  NAND2_X1 U10731 ( .A1(n10669), .A2(n10671), .ZN(n10791) );
  NAND2_X1 U10732 ( .A1(n10792), .A2(n10793), .ZN(n10671) );
  NAND2_X1 U10733 ( .A1(b_25_), .A2(a_16_), .ZN(n10793) );
  INV_X1 U10734 ( .A(n10794), .ZN(n10792) );
  XNOR2_X1 U10735 ( .A(n10795), .B(n10796), .ZN(n10669) );
  XNOR2_X1 U10736 ( .A(n10797), .B(n10798), .ZN(n10796) );
  NAND2_X1 U10737 ( .A1(a_16_), .A2(n10794), .ZN(n10670) );
  NAND2_X1 U10738 ( .A1(n10799), .A2(n10800), .ZN(n10794) );
  NAND3_X1 U10739 ( .A1(a_17_), .A2(n10801), .A3(b_25_), .ZN(n10800) );
  NAND2_X1 U10740 ( .A1(n10558), .A2(n10560), .ZN(n10801) );
  INV_X1 U10741 ( .A(n10802), .ZN(n10799) );
  NOR2_X1 U10742 ( .A1(n10560), .A2(n10558), .ZN(n10802) );
  XOR2_X1 U10743 ( .A(n10803), .B(n10804), .Z(n10558) );
  XOR2_X1 U10744 ( .A(n10805), .B(n10806), .Z(n10803) );
  NAND2_X1 U10745 ( .A1(n10807), .A2(n10808), .ZN(n10560) );
  NAND2_X1 U10746 ( .A1(n10568), .A2(n10809), .ZN(n10808) );
  NAND2_X1 U10747 ( .A1(n10570), .A2(n10569), .ZN(n10809) );
  XNOR2_X1 U10748 ( .A(n10810), .B(n10811), .ZN(n10568) );
  XOR2_X1 U10749 ( .A(n10812), .B(n10813), .Z(n10810) );
  NOR2_X1 U10750 ( .A1(n8630), .A2(n8981), .ZN(n10813) );
  INV_X1 U10751 ( .A(n10814), .ZN(n10807) );
  NOR2_X1 U10752 ( .A1(n10569), .A2(n10570), .ZN(n10814) );
  NOR2_X1 U10753 ( .A1(n8543), .A2(n8988), .ZN(n10570) );
  NAND2_X1 U10754 ( .A1(n10815), .A2(n10816), .ZN(n10569) );
  NAND3_X1 U10755 ( .A1(a_19_), .A2(n10817), .A3(b_25_), .ZN(n10816) );
  INV_X1 U10756 ( .A(n10818), .ZN(n10817) );
  NOR2_X1 U10757 ( .A1(n10576), .A2(n10575), .ZN(n10818) );
  NAND2_X1 U10758 ( .A1(n10575), .A2(n10576), .ZN(n10815) );
  NAND2_X1 U10759 ( .A1(n10666), .A2(n10819), .ZN(n10576) );
  NAND2_X1 U10760 ( .A1(n10665), .A2(n10667), .ZN(n10819) );
  NAND2_X1 U10761 ( .A1(n10820), .A2(n10821), .ZN(n10667) );
  NAND2_X1 U10762 ( .A1(b_25_), .A2(a_20_), .ZN(n10821) );
  INV_X1 U10763 ( .A(n10822), .ZN(n10820) );
  XOR2_X1 U10764 ( .A(n10823), .B(n10824), .Z(n10665) );
  XOR2_X1 U10765 ( .A(n10825), .B(n10826), .Z(n10823) );
  NOR2_X1 U10766 ( .A1(n8601), .A2(n8981), .ZN(n10826) );
  NAND2_X1 U10767 ( .A1(a_20_), .A2(n10822), .ZN(n10666) );
  NAND2_X1 U10768 ( .A1(n10827), .A2(n10828), .ZN(n10822) );
  INV_X1 U10769 ( .A(n10829), .ZN(n10828) );
  NOR3_X1 U10770 ( .A1(n8601), .A2(n10830), .A3(n8543), .ZN(n10829) );
  NOR2_X1 U10771 ( .A1(n10589), .A2(n10587), .ZN(n10830) );
  NAND2_X1 U10772 ( .A1(n10587), .A2(n10589), .ZN(n10827) );
  NAND2_X1 U10773 ( .A1(n10662), .A2(n10831), .ZN(n10589) );
  NAND2_X1 U10774 ( .A1(n10661), .A2(n10663), .ZN(n10831) );
  NAND2_X1 U10775 ( .A1(n10832), .A2(n10833), .ZN(n10663) );
  NAND2_X1 U10776 ( .A1(b_25_), .A2(a_22_), .ZN(n10833) );
  INV_X1 U10777 ( .A(n10834), .ZN(n10832) );
  XNOR2_X1 U10778 ( .A(n10835), .B(n10836), .ZN(n10661) );
  NAND2_X1 U10779 ( .A1(n10837), .A2(n10838), .ZN(n10835) );
  NAND2_X1 U10780 ( .A1(a_22_), .A2(n10834), .ZN(n10662) );
  NAND2_X1 U10781 ( .A1(n10601), .A2(n10839), .ZN(n10834) );
  NAND2_X1 U10782 ( .A1(n10600), .A2(n10602), .ZN(n10839) );
  NAND2_X1 U10783 ( .A1(n10840), .A2(n10841), .ZN(n10602) );
  NAND2_X1 U10784 ( .A1(b_25_), .A2(a_23_), .ZN(n10841) );
  XNOR2_X1 U10785 ( .A(n10842), .B(n10843), .ZN(n10600) );
  XOR2_X1 U10786 ( .A(n10844), .B(n8555), .Z(n10842) );
  NAND2_X1 U10787 ( .A1(a_23_), .A2(n10845), .ZN(n10601) );
  INV_X1 U10788 ( .A(n10840), .ZN(n10845) );
  NOR2_X1 U10789 ( .A1(n10846), .A2(n10847), .ZN(n10840) );
  INV_X1 U10790 ( .A(n10848), .ZN(n10847) );
  NAND2_X1 U10791 ( .A1(n10610), .A2(n10849), .ZN(n10848) );
  NAND2_X1 U10792 ( .A1(n10607), .A2(n10609), .ZN(n10849) );
  NOR2_X1 U10793 ( .A1(n8543), .A2(n8982), .ZN(n10610) );
  NOR2_X1 U10794 ( .A1(n10609), .A2(n10607), .ZN(n10846) );
  XOR2_X1 U10795 ( .A(n10850), .B(n10851), .Z(n10607) );
  XNOR2_X1 U10796 ( .A(n10852), .B(n10853), .ZN(n10851) );
  NAND2_X1 U10797 ( .A1(n10854), .A2(n10855), .ZN(n10609) );
  NAND2_X1 U10798 ( .A1(n10657), .A2(n10856), .ZN(n10855) );
  NAND2_X1 U10799 ( .A1(n10659), .A2(n8538), .ZN(n10856) );
  XNOR2_X1 U10800 ( .A(n10857), .B(n10858), .ZN(n10657) );
  XNOR2_X1 U10801 ( .A(n10859), .B(n10860), .ZN(n10858) );
  NAND2_X1 U10802 ( .A1(n8965), .A2(n10861), .ZN(n10854) );
  INV_X1 U10803 ( .A(n10659), .ZN(n10861) );
  NOR2_X1 U10804 ( .A1(n10862), .A2(n10863), .ZN(n10659) );
  INV_X1 U10805 ( .A(n10864), .ZN(n10863) );
  NAND2_X1 U10806 ( .A1(n10619), .A2(n10865), .ZN(n10864) );
  NAND2_X1 U10807 ( .A1(n10622), .A2(n10621), .ZN(n10865) );
  XNOR2_X1 U10808 ( .A(n10866), .B(n10867), .ZN(n10619) );
  XOR2_X1 U10809 ( .A(n10868), .B(n10869), .Z(n10866) );
  NOR2_X1 U10810 ( .A1(n10621), .A2(n10622), .ZN(n10862) );
  NOR2_X1 U10811 ( .A1(n8543), .A2(n9893), .ZN(n10622) );
  NAND2_X1 U10812 ( .A1(n10870), .A2(n10871), .ZN(n10621) );
  NAND2_X1 U10813 ( .A1(n10629), .A2(n10872), .ZN(n10871) );
  INV_X1 U10814 ( .A(n10873), .ZN(n10872) );
  NOR2_X1 U10815 ( .A1(n10628), .A2(n10627), .ZN(n10873) );
  NOR2_X1 U10816 ( .A1(n8543), .A2(n8512), .ZN(n10629) );
  NAND2_X1 U10817 ( .A1(n10627), .A2(n10628), .ZN(n10870) );
  NAND2_X1 U10818 ( .A1(n10874), .A2(n10875), .ZN(n10628) );
  NAND2_X1 U10819 ( .A1(n10655), .A2(n10876), .ZN(n10875) );
  INV_X1 U10820 ( .A(n10877), .ZN(n10876) );
  NOR2_X1 U10821 ( .A1(n10656), .A2(n10654), .ZN(n10877) );
  NOR2_X1 U10822 ( .A1(n8543), .A2(n8493), .ZN(n10655) );
  NAND2_X1 U10823 ( .A1(n10654), .A2(n10656), .ZN(n10874) );
  NAND2_X1 U10824 ( .A1(n10878), .A2(n10879), .ZN(n10656) );
  NAND2_X1 U10825 ( .A1(n10650), .A2(n10880), .ZN(n10879) );
  INV_X1 U10826 ( .A(n10881), .ZN(n10880) );
  NOR2_X1 U10827 ( .A1(n10651), .A2(n10652), .ZN(n10881) );
  NOR2_X1 U10828 ( .A1(n8543), .A2(n8473), .ZN(n10650) );
  NAND2_X1 U10829 ( .A1(n10652), .A2(n10651), .ZN(n10878) );
  NAND2_X1 U10830 ( .A1(n10882), .A2(n10883), .ZN(n10651) );
  NAND2_X1 U10831 ( .A1(b_23_), .A2(n10884), .ZN(n10883) );
  NAND2_X1 U10832 ( .A1(n8456), .A2(n10885), .ZN(n10884) );
  NAND2_X1 U10833 ( .A1(a_31_), .A2(n8981), .ZN(n10885) );
  NAND2_X1 U10834 ( .A1(b_24_), .A2(n10886), .ZN(n10882) );
  NAND2_X1 U10835 ( .A1(n8459), .A2(n10887), .ZN(n10886) );
  NAND2_X1 U10836 ( .A1(a_30_), .A2(n8570), .ZN(n10887) );
  NOR3_X1 U10837 ( .A1(n8981), .A2(n8979), .A3(n8543), .ZN(n10652) );
  XOR2_X1 U10838 ( .A(n10888), .B(n10889), .Z(n10654) );
  XOR2_X1 U10839 ( .A(n10890), .B(n10891), .Z(n10888) );
  XOR2_X1 U10840 ( .A(n10892), .B(n10893), .Z(n10627) );
  XOR2_X1 U10841 ( .A(n10894), .B(n10895), .Z(n10892) );
  INV_X1 U10842 ( .A(n8538), .ZN(n8965) );
  NOR2_X1 U10843 ( .A1(n8543), .A2(n8541), .ZN(n8538) );
  XNOR2_X1 U10844 ( .A(n10896), .B(n10897), .ZN(n10587) );
  NAND2_X1 U10845 ( .A1(n10898), .A2(n10899), .ZN(n10896) );
  XNOR2_X1 U10846 ( .A(n10900), .B(n10901), .ZN(n10575) );
  NAND2_X1 U10847 ( .A1(n10902), .A2(n10903), .ZN(n10900) );
  XNOR2_X1 U10848 ( .A(n10904), .B(n10905), .ZN(n10547) );
  NAND2_X1 U10849 ( .A1(n10906), .A2(n10907), .ZN(n10904) );
  XNOR2_X1 U10850 ( .A(n10908), .B(n10909), .ZN(n10536) );
  NAND2_X1 U10851 ( .A1(n10910), .A2(n10911), .ZN(n10908) );
  XOR2_X1 U10852 ( .A(n10912), .B(n10913), .Z(n10524) );
  XNOR2_X1 U10853 ( .A(n10914), .B(n10915), .ZN(n10913) );
  NAND2_X1 U10854 ( .A1(b_24_), .A2(a_12_), .ZN(n10915) );
  NAND2_X1 U10855 ( .A1(n10683), .A2(n10916), .ZN(n10759) );
  INV_X1 U10856 ( .A(n10680), .ZN(n10916) );
  XOR2_X1 U10857 ( .A(n10917), .B(n10918), .Z(n10680) );
  NAND2_X1 U10858 ( .A1(n10919), .A2(n10920), .ZN(n10917) );
  NOR2_X1 U10859 ( .A1(n8543), .A2(n8769), .ZN(n10683) );
  XNOR2_X1 U10860 ( .A(n10921), .B(n10922), .ZN(n10685) );
  NAND2_X1 U10861 ( .A1(n10923), .A2(n10924), .ZN(n10921) );
  XOR2_X1 U10862 ( .A(n10925), .B(n10926), .Z(n10689) );
  XOR2_X1 U10863 ( .A(n10927), .B(n10928), .Z(n10926) );
  NAND2_X1 U10864 ( .A1(b_24_), .A2(a_9_), .ZN(n10928) );
  XOR2_X1 U10865 ( .A(n10929), .B(n10930), .Z(n10692) );
  XOR2_X1 U10866 ( .A(n10931), .B(n10932), .Z(n10930) );
  NAND2_X1 U10867 ( .A1(b_24_), .A2(a_8_), .ZN(n10932) );
  XNOR2_X1 U10868 ( .A(n10933), .B(n10934), .ZN(n10700) );
  XNOR2_X1 U10869 ( .A(n10935), .B(n10936), .ZN(n10933) );
  XNOR2_X1 U10870 ( .A(n10937), .B(n10938), .ZN(n10704) );
  XNOR2_X1 U10871 ( .A(n10939), .B(n10940), .ZN(n10937) );
  XNOR2_X1 U10872 ( .A(n10941), .B(n10942), .ZN(n10486) );
  XNOR2_X1 U10873 ( .A(n10943), .B(n10944), .ZN(n10942) );
  NAND2_X1 U10874 ( .A1(b_24_), .A2(a_4_), .ZN(n10944) );
  XNOR2_X1 U10875 ( .A(n10945), .B(n10946), .ZN(n10478) );
  XOR2_X1 U10876 ( .A(n10947), .B(n10948), .Z(n10945) );
  XOR2_X1 U10877 ( .A(n10949), .B(n10950), .Z(n10470) );
  XOR2_X1 U10878 ( .A(n10951), .B(n10952), .Z(n10950) );
  NAND2_X1 U10879 ( .A1(b_24_), .A2(a_2_), .ZN(n10952) );
  XOR2_X1 U10880 ( .A(n10953), .B(n10954), .Z(n10710) );
  XNOR2_X1 U10881 ( .A(n10955), .B(n10956), .ZN(n10953) );
  XNOR2_X1 U10882 ( .A(n10957), .B(n10958), .ZN(n10709) );
  XNOR2_X1 U10883 ( .A(n10959), .B(n10960), .ZN(n10958) );
  NAND2_X1 U10884 ( .A1(b_24_), .A2(a_0_), .ZN(n10960) );
  NAND4_X1 U10885 ( .A1(n9193), .A2(n9191), .A3(n9194), .A4(n9192), .ZN(n9052)
         );
  INV_X1 U10886 ( .A(n9183), .ZN(n9192) );
  NOR2_X1 U10887 ( .A1(n10961), .A2(n10962), .ZN(n9183) );
  NAND2_X1 U10888 ( .A1(n10963), .A2(n10964), .ZN(n9194) );
  NAND3_X1 U10889 ( .A1(a_0_), .A2(n10965), .A3(b_24_), .ZN(n10964) );
  NAND2_X1 U10890 ( .A1(n10959), .A2(n10957), .ZN(n10965) );
  INV_X1 U10891 ( .A(n10966), .ZN(n10963) );
  NOR2_X1 U10892 ( .A1(n10957), .A2(n10959), .ZN(n10966) );
  NOR2_X1 U10893 ( .A1(n10967), .A2(n10968), .ZN(n10959) );
  INV_X1 U10894 ( .A(n10969), .ZN(n10968) );
  NAND2_X1 U10895 ( .A1(n10955), .A2(n10970), .ZN(n10969) );
  NAND2_X1 U10896 ( .A1(n10954), .A2(n10956), .ZN(n10970) );
  NAND2_X1 U10897 ( .A1(n10971), .A2(n10972), .ZN(n10955) );
  INV_X1 U10898 ( .A(n10973), .ZN(n10972) );
  NOR3_X1 U10899 ( .A1(n8998), .A2(n10974), .A3(n8981), .ZN(n10973) );
  NOR2_X1 U10900 ( .A1(n10951), .A2(n10949), .ZN(n10974) );
  NAND2_X1 U10901 ( .A1(n10949), .A2(n10951), .ZN(n10971) );
  NAND2_X1 U10902 ( .A1(n10975), .A2(n10976), .ZN(n10951) );
  NAND2_X1 U10903 ( .A1(n10947), .A2(n10977), .ZN(n10976) );
  INV_X1 U10904 ( .A(n10978), .ZN(n10977) );
  NOR2_X1 U10905 ( .A1(n10946), .A2(n10948), .ZN(n10978) );
  NAND2_X1 U10906 ( .A1(n10979), .A2(n10980), .ZN(n10947) );
  NAND3_X1 U10907 ( .A1(a_4_), .A2(n10981), .A3(b_24_), .ZN(n10980) );
  NAND2_X1 U10908 ( .A1(n10943), .A2(n10982), .ZN(n10981) );
  INV_X1 U10909 ( .A(n10941), .ZN(n10982) );
  NAND2_X1 U10910 ( .A1(n10941), .A2(n10983), .ZN(n10979) );
  INV_X1 U10911 ( .A(n10943), .ZN(n10983) );
  NOR2_X1 U10912 ( .A1(n10984), .A2(n10985), .ZN(n10943) );
  INV_X1 U10913 ( .A(n10986), .ZN(n10985) );
  NAND2_X1 U10914 ( .A1(n10940), .A2(n10987), .ZN(n10986) );
  NAND2_X1 U10915 ( .A1(n10939), .A2(n10938), .ZN(n10987) );
  NOR2_X1 U10916 ( .A1(n8981), .A2(n8848), .ZN(n10940) );
  NOR2_X1 U10917 ( .A1(n10938), .A2(n10939), .ZN(n10984) );
  NOR2_X1 U10918 ( .A1(n10988), .A2(n10989), .ZN(n10939) );
  INV_X1 U10919 ( .A(n10990), .ZN(n10989) );
  NAND2_X1 U10920 ( .A1(n10936), .A2(n10991), .ZN(n10990) );
  NAND2_X1 U10921 ( .A1(n10935), .A2(n10934), .ZN(n10991) );
  NOR2_X1 U10922 ( .A1(n8981), .A2(n8994), .ZN(n10936) );
  NOR2_X1 U10923 ( .A1(n10934), .A2(n10935), .ZN(n10988) );
  INV_X1 U10924 ( .A(n10992), .ZN(n10935) );
  NAND2_X1 U10925 ( .A1(n10744), .A2(n10993), .ZN(n10992) );
  NAND2_X1 U10926 ( .A1(n10743), .A2(n10745), .ZN(n10993) );
  NAND2_X1 U10927 ( .A1(n10994), .A2(n10995), .ZN(n10745) );
  NAND2_X1 U10928 ( .A1(b_24_), .A2(a_7_), .ZN(n10995) );
  XNOR2_X1 U10929 ( .A(n10996), .B(n10997), .ZN(n10743) );
  XOR2_X1 U10930 ( .A(n10998), .B(n10999), .Z(n10996) );
  INV_X1 U10931 ( .A(n11000), .ZN(n10744) );
  NOR2_X1 U10932 ( .A1(n8817), .A2(n10994), .ZN(n11000) );
  NOR2_X1 U10933 ( .A1(n11001), .A2(n11002), .ZN(n10994) );
  NOR3_X1 U10934 ( .A1(n10513), .A2(n11003), .A3(n8981), .ZN(n11002) );
  NOR2_X1 U10935 ( .A1(n10931), .A2(n10929), .ZN(n11003) );
  INV_X1 U10936 ( .A(n11004), .ZN(n11001) );
  NAND2_X1 U10937 ( .A1(n10929), .A2(n10931), .ZN(n11004) );
  NAND2_X1 U10938 ( .A1(n11005), .A2(n11006), .ZN(n10931) );
  INV_X1 U10939 ( .A(n11007), .ZN(n11006) );
  NOR3_X1 U10940 ( .A1(n8779), .A2(n11008), .A3(n8981), .ZN(n11007) );
  NOR2_X1 U10941 ( .A1(n10927), .A2(n10925), .ZN(n11008) );
  NAND2_X1 U10942 ( .A1(n10925), .A2(n10927), .ZN(n11005) );
  NAND2_X1 U10943 ( .A1(n10923), .A2(n11009), .ZN(n10927) );
  NAND2_X1 U10944 ( .A1(n10922), .A2(n10924), .ZN(n11009) );
  NAND2_X1 U10945 ( .A1(n11010), .A2(n11011), .ZN(n10924) );
  NAND2_X1 U10946 ( .A1(b_24_), .A2(a_10_), .ZN(n11011) );
  INV_X1 U10947 ( .A(n11012), .ZN(n11010) );
  XNOR2_X1 U10948 ( .A(n11013), .B(n11014), .ZN(n10922) );
  XOR2_X1 U10949 ( .A(n11015), .B(n11016), .Z(n11014) );
  NAND2_X1 U10950 ( .A1(b_23_), .A2(a_11_), .ZN(n11016) );
  NAND2_X1 U10951 ( .A1(a_10_), .A2(n11012), .ZN(n10923) );
  NAND2_X1 U10952 ( .A1(n10919), .A2(n11017), .ZN(n11012) );
  NAND2_X1 U10953 ( .A1(n10918), .A2(n10920), .ZN(n11017) );
  NAND2_X1 U10954 ( .A1(n11018), .A2(n11019), .ZN(n10920) );
  NAND2_X1 U10955 ( .A1(b_24_), .A2(a_11_), .ZN(n11019) );
  XOR2_X1 U10956 ( .A(n11020), .B(n11021), .Z(n10918) );
  XNOR2_X1 U10957 ( .A(n11022), .B(n11023), .ZN(n11021) );
  INV_X1 U10958 ( .A(n11024), .ZN(n10919) );
  NOR2_X1 U10959 ( .A1(n8749), .A2(n11018), .ZN(n11024) );
  NOR2_X1 U10960 ( .A1(n11025), .A2(n11026), .ZN(n11018) );
  INV_X1 U10961 ( .A(n11027), .ZN(n11026) );
  NAND3_X1 U10962 ( .A1(a_12_), .A2(n11028), .A3(b_24_), .ZN(n11027) );
  NAND2_X1 U10963 ( .A1(n10914), .A2(n10912), .ZN(n11028) );
  NOR2_X1 U10964 ( .A1(n10912), .A2(n10914), .ZN(n11025) );
  NOR2_X1 U10965 ( .A1(n11029), .A2(n11030), .ZN(n10914) );
  NOR3_X1 U10966 ( .A1(n8721), .A2(n11031), .A3(n8981), .ZN(n11030) );
  NOR2_X1 U10967 ( .A1(n10773), .A2(n10772), .ZN(n11031) );
  INV_X1 U10968 ( .A(n11032), .ZN(n11029) );
  NAND2_X1 U10969 ( .A1(n10772), .A2(n10773), .ZN(n11032) );
  NAND2_X1 U10970 ( .A1(n10910), .A2(n11033), .ZN(n10773) );
  NAND2_X1 U10971 ( .A1(n10909), .A2(n10911), .ZN(n11033) );
  NAND2_X1 U10972 ( .A1(n11034), .A2(n11035), .ZN(n10911) );
  NAND2_X1 U10973 ( .A1(b_24_), .A2(a_14_), .ZN(n11035) );
  XOR2_X1 U10974 ( .A(n11036), .B(n11037), .Z(n10909) );
  XOR2_X1 U10975 ( .A(n11038), .B(n11039), .Z(n11036) );
  NOR2_X1 U10976 ( .A1(n8692), .A2(n8570), .ZN(n11039) );
  INV_X1 U10977 ( .A(n11040), .ZN(n10910) );
  NOR2_X1 U10978 ( .A1(n8991), .A2(n11034), .ZN(n11040) );
  NOR2_X1 U10979 ( .A1(n11041), .A2(n11042), .ZN(n11034) );
  NOR3_X1 U10980 ( .A1(n8692), .A2(n11043), .A3(n8981), .ZN(n11042) );
  NOR2_X1 U10981 ( .A1(n10785), .A2(n10784), .ZN(n11043) );
  INV_X1 U10982 ( .A(n11044), .ZN(n11041) );
  NAND2_X1 U10983 ( .A1(n10784), .A2(n10785), .ZN(n11044) );
  NAND2_X1 U10984 ( .A1(n10906), .A2(n11045), .ZN(n10785) );
  NAND2_X1 U10985 ( .A1(n10905), .A2(n10907), .ZN(n11045) );
  NAND2_X1 U10986 ( .A1(n11046), .A2(n11047), .ZN(n10907) );
  NAND2_X1 U10987 ( .A1(b_24_), .A2(a_16_), .ZN(n11047) );
  INV_X1 U10988 ( .A(n11048), .ZN(n11046) );
  XNOR2_X1 U10989 ( .A(n11049), .B(n11050), .ZN(n10905) );
  XOR2_X1 U10990 ( .A(n11051), .B(n11052), .Z(n11050) );
  NAND2_X1 U10991 ( .A1(b_23_), .A2(a_17_), .ZN(n11052) );
  NAND2_X1 U10992 ( .A1(a_16_), .A2(n11048), .ZN(n10906) );
  NAND2_X1 U10993 ( .A1(n11053), .A2(n11054), .ZN(n11048) );
  NAND2_X1 U10994 ( .A1(n10798), .A2(n11055), .ZN(n11054) );
  NAND2_X1 U10995 ( .A1(n10795), .A2(n10797), .ZN(n11055) );
  NOR2_X1 U10996 ( .A1(n8981), .A2(n8662), .ZN(n10798) );
  INV_X1 U10997 ( .A(n11056), .ZN(n11053) );
  NOR2_X1 U10998 ( .A1(n10797), .A2(n10795), .ZN(n11056) );
  XNOR2_X1 U10999 ( .A(n11057), .B(n11058), .ZN(n10795) );
  XNOR2_X1 U11000 ( .A(n11059), .B(n11060), .ZN(n11058) );
  NAND2_X1 U11001 ( .A1(n11061), .A2(n11062), .ZN(n10797) );
  NAND2_X1 U11002 ( .A1(n10804), .A2(n11063), .ZN(n11062) );
  NAND2_X1 U11003 ( .A1(n10806), .A2(n10805), .ZN(n11063) );
  XNOR2_X1 U11004 ( .A(n11064), .B(n11065), .ZN(n10804) );
  XOR2_X1 U11005 ( .A(n11066), .B(n11067), .Z(n11064) );
  NOR2_X1 U11006 ( .A1(n8630), .A2(n8570), .ZN(n11067) );
  INV_X1 U11007 ( .A(n11068), .ZN(n11061) );
  NOR2_X1 U11008 ( .A1(n10805), .A2(n10806), .ZN(n11068) );
  NOR2_X1 U11009 ( .A1(n8981), .A2(n8988), .ZN(n10806) );
  NAND2_X1 U11010 ( .A1(n11069), .A2(n11070), .ZN(n10805) );
  NAND3_X1 U11011 ( .A1(a_19_), .A2(n11071), .A3(b_24_), .ZN(n11070) );
  INV_X1 U11012 ( .A(n11072), .ZN(n11071) );
  NOR2_X1 U11013 ( .A1(n10812), .A2(n10811), .ZN(n11072) );
  NAND2_X1 U11014 ( .A1(n10811), .A2(n10812), .ZN(n11069) );
  NAND2_X1 U11015 ( .A1(n10902), .A2(n11073), .ZN(n10812) );
  NAND2_X1 U11016 ( .A1(n10901), .A2(n10903), .ZN(n11073) );
  NAND2_X1 U11017 ( .A1(n11074), .A2(n11075), .ZN(n10903) );
  NAND2_X1 U11018 ( .A1(b_24_), .A2(a_20_), .ZN(n11075) );
  XNOR2_X1 U11019 ( .A(n11076), .B(n11077), .ZN(n10901) );
  XOR2_X1 U11020 ( .A(n11078), .B(n11079), .Z(n11077) );
  NAND2_X1 U11021 ( .A1(b_23_), .A2(a_21_), .ZN(n11079) );
  INV_X1 U11022 ( .A(n11080), .ZN(n10902) );
  NOR2_X1 U11023 ( .A1(n8986), .A2(n11074), .ZN(n11080) );
  NOR2_X1 U11024 ( .A1(n11081), .A2(n11082), .ZN(n11074) );
  NOR3_X1 U11025 ( .A1(n8601), .A2(n11083), .A3(n8981), .ZN(n11082) );
  NOR2_X1 U11026 ( .A1(n10825), .A2(n10824), .ZN(n11083) );
  INV_X1 U11027 ( .A(n11084), .ZN(n11081) );
  NAND2_X1 U11028 ( .A1(n10824), .A2(n10825), .ZN(n11084) );
  NAND2_X1 U11029 ( .A1(n10898), .A2(n11085), .ZN(n10825) );
  NAND2_X1 U11030 ( .A1(n10897), .A2(n10899), .ZN(n11085) );
  NAND2_X1 U11031 ( .A1(n11086), .A2(n11087), .ZN(n10899) );
  NAND2_X1 U11032 ( .A1(b_24_), .A2(a_22_), .ZN(n11087) );
  INV_X1 U11033 ( .A(n11088), .ZN(n11086) );
  XNOR2_X1 U11034 ( .A(n11089), .B(n11090), .ZN(n10897) );
  XNOR2_X1 U11035 ( .A(n11091), .B(n8961), .ZN(n11089) );
  NAND2_X1 U11036 ( .A1(a_22_), .A2(n11088), .ZN(n10898) );
  NAND2_X1 U11037 ( .A1(n10837), .A2(n11092), .ZN(n11088) );
  NAND2_X1 U11038 ( .A1(n10836), .A2(n10838), .ZN(n11092) );
  NAND2_X1 U11039 ( .A1(n11093), .A2(n11094), .ZN(n10838) );
  NAND2_X1 U11040 ( .A1(b_24_), .A2(a_23_), .ZN(n11093) );
  XOR2_X1 U11041 ( .A(n11095), .B(n11096), .Z(n10836) );
  XOR2_X1 U11042 ( .A(n11097), .B(n11098), .Z(n11095) );
  NAND2_X1 U11043 ( .A1(n11099), .A2(a_23_), .ZN(n10837) );
  INV_X1 U11044 ( .A(n11094), .ZN(n11099) );
  NAND2_X1 U11045 ( .A1(n11100), .A2(n11101), .ZN(n11094) );
  NAND2_X1 U11046 ( .A1(n10843), .A2(n11102), .ZN(n11101) );
  INV_X1 U11047 ( .A(n11103), .ZN(n11102) );
  NOR2_X1 U11048 ( .A1(n8555), .A2(n10844), .ZN(n11103) );
  XOR2_X1 U11049 ( .A(n11104), .B(n11105), .Z(n10843) );
  XNOR2_X1 U11050 ( .A(n11106), .B(n11107), .ZN(n11105) );
  NAND2_X1 U11051 ( .A1(n10844), .A2(n8555), .ZN(n11100) );
  NAND2_X1 U11052 ( .A1(b_24_), .A2(a_24_), .ZN(n8555) );
  NOR2_X1 U11053 ( .A1(n11108), .A2(n11109), .ZN(n10844) );
  INV_X1 U11054 ( .A(n11110), .ZN(n11109) );
  NAND2_X1 U11055 ( .A1(n10853), .A2(n11111), .ZN(n11110) );
  NAND2_X1 U11056 ( .A1(n10850), .A2(n10852), .ZN(n11111) );
  NOR2_X1 U11057 ( .A1(n8981), .A2(n8541), .ZN(n10853) );
  NOR2_X1 U11058 ( .A1(n10852), .A2(n10850), .ZN(n11108) );
  XNOR2_X1 U11059 ( .A(n11112), .B(n11113), .ZN(n10850) );
  XNOR2_X1 U11060 ( .A(n11114), .B(n11115), .ZN(n11113) );
  NAND2_X1 U11061 ( .A1(n11116), .A2(n11117), .ZN(n10852) );
  NAND2_X1 U11062 ( .A1(n10857), .A2(n11118), .ZN(n11117) );
  NAND2_X1 U11063 ( .A1(n10860), .A2(n10859), .ZN(n11118) );
  XNOR2_X1 U11064 ( .A(n11119), .B(n11120), .ZN(n10857) );
  XOR2_X1 U11065 ( .A(n11121), .B(n11122), .Z(n11119) );
  INV_X1 U11066 ( .A(n11123), .ZN(n11116) );
  NOR2_X1 U11067 ( .A1(n10859), .A2(n10860), .ZN(n11123) );
  NOR2_X1 U11068 ( .A1(n8981), .A2(n9893), .ZN(n10860) );
  NAND2_X1 U11069 ( .A1(n11124), .A2(n11125), .ZN(n10859) );
  NAND2_X1 U11070 ( .A1(n10869), .A2(n11126), .ZN(n11125) );
  INV_X1 U11071 ( .A(n11127), .ZN(n11126) );
  NOR2_X1 U11072 ( .A1(n10868), .A2(n10867), .ZN(n11127) );
  NOR2_X1 U11073 ( .A1(n8981), .A2(n8512), .ZN(n10869) );
  NAND2_X1 U11074 ( .A1(n10867), .A2(n10868), .ZN(n11124) );
  NAND2_X1 U11075 ( .A1(n11128), .A2(n11129), .ZN(n10868) );
  NAND2_X1 U11076 ( .A1(n10894), .A2(n11130), .ZN(n11129) );
  INV_X1 U11077 ( .A(n11131), .ZN(n11130) );
  NOR2_X1 U11078 ( .A1(n10895), .A2(n10893), .ZN(n11131) );
  NOR2_X1 U11079 ( .A1(n8981), .A2(n8493), .ZN(n10894) );
  NAND2_X1 U11080 ( .A1(n10893), .A2(n10895), .ZN(n11128) );
  NAND2_X1 U11081 ( .A1(n11132), .A2(n11133), .ZN(n10895) );
  NAND2_X1 U11082 ( .A1(n10889), .A2(n11134), .ZN(n11133) );
  INV_X1 U11083 ( .A(n11135), .ZN(n11134) );
  NOR2_X1 U11084 ( .A1(n10890), .A2(n10891), .ZN(n11135) );
  NOR2_X1 U11085 ( .A1(n8981), .A2(n8473), .ZN(n10889) );
  NAND2_X1 U11086 ( .A1(n10891), .A2(n10890), .ZN(n11132) );
  NAND2_X1 U11087 ( .A1(n11136), .A2(n11137), .ZN(n10890) );
  NAND2_X1 U11088 ( .A1(b_22_), .A2(n11138), .ZN(n11137) );
  NAND2_X1 U11089 ( .A1(n8456), .A2(n11139), .ZN(n11138) );
  NAND2_X1 U11090 ( .A1(a_31_), .A2(n8570), .ZN(n11139) );
  NAND2_X1 U11091 ( .A1(b_23_), .A2(n11140), .ZN(n11136) );
  NAND2_X1 U11092 ( .A1(n8459), .A2(n11141), .ZN(n11140) );
  NAND2_X1 U11093 ( .A1(a_30_), .A2(n8983), .ZN(n11141) );
  NOR3_X1 U11094 ( .A1(n8570), .A2(n8979), .A3(n8981), .ZN(n10891) );
  XOR2_X1 U11095 ( .A(n11142), .B(n11143), .Z(n10893) );
  XOR2_X1 U11096 ( .A(n11144), .B(n11145), .Z(n11142) );
  XOR2_X1 U11097 ( .A(n11146), .B(n11147), .Z(n10867) );
  XOR2_X1 U11098 ( .A(n11148), .B(n11149), .Z(n11146) );
  XNOR2_X1 U11099 ( .A(n11150), .B(n11151), .ZN(n10824) );
  NAND2_X1 U11100 ( .A1(n11152), .A2(n11153), .ZN(n11150) );
  XNOR2_X1 U11101 ( .A(n11154), .B(n11155), .ZN(n10811) );
  NAND2_X1 U11102 ( .A1(n11156), .A2(n11157), .ZN(n11154) );
  XOR2_X1 U11103 ( .A(n11158), .B(n11159), .Z(n10784) );
  XNOR2_X1 U11104 ( .A(n11160), .B(n11161), .ZN(n11159) );
  XNOR2_X1 U11105 ( .A(n11162), .B(n11163), .ZN(n10772) );
  NAND2_X1 U11106 ( .A1(n11164), .A2(n11165), .ZN(n11162) );
  XOR2_X1 U11107 ( .A(n11166), .B(n11167), .Z(n10912) );
  XOR2_X1 U11108 ( .A(n11168), .B(n11169), .Z(n11167) );
  NAND2_X1 U11109 ( .A1(b_23_), .A2(a_13_), .ZN(n11169) );
  XNOR2_X1 U11110 ( .A(n11170), .B(n11171), .ZN(n10925) );
  XNOR2_X1 U11111 ( .A(n11172), .B(n11173), .ZN(n11170) );
  XOR2_X1 U11112 ( .A(n11174), .B(n11175), .Z(n10929) );
  XOR2_X1 U11113 ( .A(n11176), .B(n11177), .Z(n11175) );
  XOR2_X1 U11114 ( .A(n11178), .B(n11179), .Z(n10934) );
  XOR2_X1 U11115 ( .A(n11180), .B(n11181), .Z(n11179) );
  NAND2_X1 U11116 ( .A1(b_23_), .A2(a_7_), .ZN(n11181) );
  XOR2_X1 U11117 ( .A(n11182), .B(n11183), .Z(n10938) );
  NAND2_X1 U11118 ( .A1(n11184), .A2(n11185), .ZN(n11182) );
  XOR2_X1 U11119 ( .A(n11186), .B(n11187), .Z(n10941) );
  XOR2_X1 U11120 ( .A(n11188), .B(n11189), .Z(n11186) );
  NOR2_X1 U11121 ( .A1(n8848), .A2(n8570), .ZN(n11189) );
  NAND2_X1 U11122 ( .A1(n10948), .A2(n10946), .ZN(n10975) );
  XNOR2_X1 U11123 ( .A(n11190), .B(n11191), .ZN(n10946) );
  XNOR2_X1 U11124 ( .A(n11192), .B(n11193), .ZN(n11190) );
  NOR2_X1 U11125 ( .A1(n8996), .A2(n8570), .ZN(n11193) );
  NOR2_X1 U11126 ( .A1(n8981), .A2(n8877), .ZN(n10948) );
  INV_X1 U11127 ( .A(b_24_), .ZN(n8981) );
  XOR2_X1 U11128 ( .A(n11194), .B(n11195), .Z(n10949) );
  XNOR2_X1 U11129 ( .A(n11196), .B(n11197), .ZN(n11195) );
  NAND2_X1 U11130 ( .A1(b_23_), .A2(a_3_), .ZN(n11197) );
  NOR2_X1 U11131 ( .A1(n10956), .A2(n10954), .ZN(n10967) );
  XNOR2_X1 U11132 ( .A(n11198), .B(n11199), .ZN(n10954) );
  XOR2_X1 U11133 ( .A(n11200), .B(n11201), .Z(n11198) );
  NOR2_X1 U11134 ( .A1(n8998), .A2(n8570), .ZN(n11201) );
  NAND2_X1 U11135 ( .A1(b_24_), .A2(a_1_), .ZN(n10956) );
  XOR2_X1 U11136 ( .A(n11202), .B(n11203), .Z(n10957) );
  XOR2_X1 U11137 ( .A(n11204), .B(n11205), .Z(n11203) );
  NAND2_X1 U11138 ( .A1(b_23_), .A2(a_1_), .ZN(n11205) );
  NAND2_X1 U11139 ( .A1(n10962), .A2(n10961), .ZN(n9191) );
  XOR2_X1 U11140 ( .A(n11206), .B(n11207), .Z(n10961) );
  NAND2_X1 U11141 ( .A1(n11208), .A2(n11209), .ZN(n11206) );
  NOR2_X1 U11142 ( .A1(n11210), .A2(n11211), .ZN(n10962) );
  NOR3_X1 U11143 ( .A1(n9471), .A2(n11212), .A3(n8570), .ZN(n11211) );
  NOR2_X1 U11144 ( .A1(n11213), .A2(n11214), .ZN(n11212) );
  INV_X1 U11145 ( .A(n11215), .ZN(n11210) );
  NAND2_X1 U11146 ( .A1(n11214), .A2(n11213), .ZN(n11215) );
  XNOR2_X1 U11147 ( .A(n11214), .B(n11216), .ZN(n9193) );
  XOR2_X1 U11148 ( .A(n11213), .B(n11217), .Z(n11216) );
  NAND2_X1 U11149 ( .A1(b_23_), .A2(a_0_), .ZN(n11217) );
  NAND2_X1 U11150 ( .A1(n11218), .A2(n11219), .ZN(n11213) );
  INV_X1 U11151 ( .A(n11220), .ZN(n11219) );
  NOR3_X1 U11152 ( .A1(n9731), .A2(n11221), .A3(n8570), .ZN(n11220) );
  NOR2_X1 U11153 ( .A1(n11204), .A2(n11202), .ZN(n11221) );
  NAND2_X1 U11154 ( .A1(n11202), .A2(n11204), .ZN(n11218) );
  NAND2_X1 U11155 ( .A1(n11222), .A2(n11223), .ZN(n11204) );
  NAND3_X1 U11156 ( .A1(a_2_), .A2(n11224), .A3(b_23_), .ZN(n11223) );
  INV_X1 U11157 ( .A(n11225), .ZN(n11224) );
  NOR2_X1 U11158 ( .A1(n11200), .A2(n11199), .ZN(n11225) );
  NAND2_X1 U11159 ( .A1(n11199), .A2(n11200), .ZN(n11222) );
  NAND2_X1 U11160 ( .A1(n11226), .A2(n11227), .ZN(n11200) );
  NAND3_X1 U11161 ( .A1(a_3_), .A2(n11228), .A3(b_23_), .ZN(n11227) );
  NAND2_X1 U11162 ( .A1(n11196), .A2(n11194), .ZN(n11228) );
  INV_X1 U11163 ( .A(n11229), .ZN(n11226) );
  NOR2_X1 U11164 ( .A1(n11194), .A2(n11196), .ZN(n11229) );
  NOR2_X1 U11165 ( .A1(n11230), .A2(n11231), .ZN(n11196) );
  NOR3_X1 U11166 ( .A1(n8996), .A2(n11232), .A3(n8570), .ZN(n11231) );
  INV_X1 U11167 ( .A(n11233), .ZN(n11232) );
  NAND2_X1 U11168 ( .A1(n11192), .A2(n11191), .ZN(n11233) );
  NOR2_X1 U11169 ( .A1(n11191), .A2(n11192), .ZN(n11230) );
  NOR2_X1 U11170 ( .A1(n11234), .A2(n11235), .ZN(n11192) );
  NOR3_X1 U11171 ( .A1(n8848), .A2(n11236), .A3(n8570), .ZN(n11235) );
  NOR2_X1 U11172 ( .A1(n11188), .A2(n11187), .ZN(n11236) );
  INV_X1 U11173 ( .A(n11237), .ZN(n11234) );
  NAND2_X1 U11174 ( .A1(n11187), .A2(n11188), .ZN(n11237) );
  NAND2_X1 U11175 ( .A1(n11184), .A2(n11238), .ZN(n11188) );
  NAND2_X1 U11176 ( .A1(n11183), .A2(n11185), .ZN(n11238) );
  NAND2_X1 U11177 ( .A1(n11239), .A2(n11240), .ZN(n11185) );
  NAND2_X1 U11178 ( .A1(b_23_), .A2(a_6_), .ZN(n11240) );
  XOR2_X1 U11179 ( .A(n11241), .B(n11242), .Z(n11183) );
  XOR2_X1 U11180 ( .A(n11243), .B(n11244), .Z(n11241) );
  NOR2_X1 U11181 ( .A1(n8817), .A2(n8983), .ZN(n11244) );
  NAND2_X1 U11182 ( .A1(a_6_), .A2(n11245), .ZN(n11184) );
  INV_X1 U11183 ( .A(n11239), .ZN(n11245) );
  NOR2_X1 U11184 ( .A1(n11246), .A2(n11247), .ZN(n11239) );
  NOR3_X1 U11185 ( .A1(n8817), .A2(n11248), .A3(n8570), .ZN(n11247) );
  INV_X1 U11186 ( .A(n11249), .ZN(n11248) );
  NAND2_X1 U11187 ( .A1(n11178), .A2(n11180), .ZN(n11249) );
  NOR2_X1 U11188 ( .A1(n11180), .A2(n11178), .ZN(n11246) );
  XOR2_X1 U11189 ( .A(n11250), .B(n11251), .Z(n11178) );
  XOR2_X1 U11190 ( .A(n11252), .B(n11253), .Z(n11251) );
  NAND2_X1 U11191 ( .A1(b_22_), .A2(a_8_), .ZN(n11253) );
  NAND2_X1 U11192 ( .A1(n11254), .A2(n11255), .ZN(n11180) );
  NAND2_X1 U11193 ( .A1(n10997), .A2(n11256), .ZN(n11255) );
  INV_X1 U11194 ( .A(n11257), .ZN(n11256) );
  NOR2_X1 U11195 ( .A1(n10998), .A2(n10999), .ZN(n11257) );
  XOR2_X1 U11196 ( .A(n11258), .B(n11259), .Z(n10997) );
  NAND2_X1 U11197 ( .A1(n11260), .A2(n11261), .ZN(n11258) );
  NAND2_X1 U11198 ( .A1(n10999), .A2(n10998), .ZN(n11254) );
  NAND2_X1 U11199 ( .A1(b_23_), .A2(a_8_), .ZN(n10998) );
  NOR2_X1 U11200 ( .A1(n11262), .A2(n11263), .ZN(n10999) );
  INV_X1 U11201 ( .A(n11264), .ZN(n11263) );
  NAND2_X1 U11202 ( .A1(n11177), .A2(n11265), .ZN(n11264) );
  NAND2_X1 U11203 ( .A1(n11176), .A2(n11174), .ZN(n11265) );
  NOR2_X1 U11204 ( .A1(n8570), .A2(n8779), .ZN(n11177) );
  NOR2_X1 U11205 ( .A1(n11174), .A2(n11176), .ZN(n11262) );
  NOR2_X1 U11206 ( .A1(n11266), .A2(n11267), .ZN(n11176) );
  INV_X1 U11207 ( .A(n11268), .ZN(n11267) );
  NAND2_X1 U11208 ( .A1(n11172), .A2(n11269), .ZN(n11268) );
  NAND2_X1 U11209 ( .A1(n11171), .A2(n11173), .ZN(n11269) );
  NAND2_X1 U11210 ( .A1(n11270), .A2(n11271), .ZN(n11172) );
  NAND3_X1 U11211 ( .A1(a_11_), .A2(n11272), .A3(b_23_), .ZN(n11271) );
  NAND2_X1 U11212 ( .A1(n11013), .A2(n11015), .ZN(n11272) );
  INV_X1 U11213 ( .A(n11273), .ZN(n11270) );
  NOR2_X1 U11214 ( .A1(n11015), .A2(n11013), .ZN(n11273) );
  XOR2_X1 U11215 ( .A(n11274), .B(n11275), .Z(n11013) );
  XNOR2_X1 U11216 ( .A(n11276), .B(n11277), .ZN(n11274) );
  NOR2_X1 U11217 ( .A1(n8739), .A2(n8983), .ZN(n11277) );
  NAND2_X1 U11218 ( .A1(n11278), .A2(n11279), .ZN(n11015) );
  NAND2_X1 U11219 ( .A1(n11020), .A2(n11280), .ZN(n11279) );
  INV_X1 U11220 ( .A(n11281), .ZN(n11280) );
  NOR2_X1 U11221 ( .A1(n11023), .A2(n11022), .ZN(n11281) );
  XOR2_X1 U11222 ( .A(n11282), .B(n11283), .Z(n11020) );
  XOR2_X1 U11223 ( .A(n11284), .B(n11285), .Z(n11283) );
  NAND2_X1 U11224 ( .A1(b_22_), .A2(a_13_), .ZN(n11285) );
  NAND2_X1 U11225 ( .A1(n11022), .A2(n11023), .ZN(n11278) );
  NAND2_X1 U11226 ( .A1(b_23_), .A2(a_12_), .ZN(n11023) );
  NOR2_X1 U11227 ( .A1(n11286), .A2(n11287), .ZN(n11022) );
  NOR3_X1 U11228 ( .A1(n8721), .A2(n11288), .A3(n8570), .ZN(n11287) );
  NOR2_X1 U11229 ( .A1(n11168), .A2(n11166), .ZN(n11288) );
  INV_X1 U11230 ( .A(n11289), .ZN(n11286) );
  NAND2_X1 U11231 ( .A1(n11166), .A2(n11168), .ZN(n11289) );
  NAND2_X1 U11232 ( .A1(n11164), .A2(n11290), .ZN(n11168) );
  NAND2_X1 U11233 ( .A1(n11163), .A2(n11165), .ZN(n11290) );
  NAND2_X1 U11234 ( .A1(n11291), .A2(n11292), .ZN(n11165) );
  NAND2_X1 U11235 ( .A1(b_23_), .A2(a_14_), .ZN(n11292) );
  XOR2_X1 U11236 ( .A(n11293), .B(n11294), .Z(n11163) );
  XOR2_X1 U11237 ( .A(n11295), .B(n11296), .Z(n11293) );
  NOR2_X1 U11238 ( .A1(n8692), .A2(n8983), .ZN(n11296) );
  NAND2_X1 U11239 ( .A1(a_14_), .A2(n11297), .ZN(n11164) );
  INV_X1 U11240 ( .A(n11291), .ZN(n11297) );
  NOR2_X1 U11241 ( .A1(n11298), .A2(n11299), .ZN(n11291) );
  NOR3_X1 U11242 ( .A1(n8692), .A2(n11300), .A3(n8570), .ZN(n11299) );
  INV_X1 U11243 ( .A(n11301), .ZN(n11300) );
  NAND2_X1 U11244 ( .A1(n11037), .A2(n11038), .ZN(n11301) );
  NOR2_X1 U11245 ( .A1(n11038), .A2(n11037), .ZN(n11298) );
  XOR2_X1 U11246 ( .A(n11302), .B(n11303), .Z(n11037) );
  NAND2_X1 U11247 ( .A1(n11304), .A2(n11305), .ZN(n11302) );
  NAND2_X1 U11248 ( .A1(n11306), .A2(n11307), .ZN(n11038) );
  NAND2_X1 U11249 ( .A1(n11158), .A2(n11308), .ZN(n11307) );
  INV_X1 U11250 ( .A(n11309), .ZN(n11308) );
  NOR2_X1 U11251 ( .A1(n11161), .A2(n11160), .ZN(n11309) );
  XOR2_X1 U11252 ( .A(n11310), .B(n11311), .Z(n11158) );
  XNOR2_X1 U11253 ( .A(n11312), .B(n11313), .ZN(n11310) );
  NOR2_X1 U11254 ( .A1(n8662), .A2(n8983), .ZN(n11313) );
  NAND2_X1 U11255 ( .A1(n11160), .A2(n11161), .ZN(n11306) );
  NAND2_X1 U11256 ( .A1(b_23_), .A2(a_16_), .ZN(n11161) );
  NOR2_X1 U11257 ( .A1(n11314), .A2(n11315), .ZN(n11160) );
  INV_X1 U11258 ( .A(n11316), .ZN(n11315) );
  NAND3_X1 U11259 ( .A1(a_17_), .A2(n11317), .A3(b_23_), .ZN(n11316) );
  NAND2_X1 U11260 ( .A1(n11049), .A2(n11051), .ZN(n11317) );
  NOR2_X1 U11261 ( .A1(n11051), .A2(n11049), .ZN(n11314) );
  XOR2_X1 U11262 ( .A(n11318), .B(n11319), .Z(n11049) );
  XOR2_X1 U11263 ( .A(n11320), .B(n11321), .Z(n11318) );
  NAND2_X1 U11264 ( .A1(n11322), .A2(n11323), .ZN(n11051) );
  NAND2_X1 U11265 ( .A1(n11057), .A2(n11324), .ZN(n11323) );
  INV_X1 U11266 ( .A(n11325), .ZN(n11324) );
  NOR2_X1 U11267 ( .A1(n11060), .A2(n11059), .ZN(n11325) );
  XOR2_X1 U11268 ( .A(n11326), .B(n11327), .Z(n11057) );
  XNOR2_X1 U11269 ( .A(n11328), .B(n11329), .ZN(n11327) );
  NAND2_X1 U11270 ( .A1(n11059), .A2(n11060), .ZN(n11322) );
  NAND2_X1 U11271 ( .A1(b_23_), .A2(a_18_), .ZN(n11060) );
  NOR2_X1 U11272 ( .A1(n11330), .A2(n11331), .ZN(n11059) );
  NOR3_X1 U11273 ( .A1(n8630), .A2(n11332), .A3(n8570), .ZN(n11331) );
  NOR2_X1 U11274 ( .A1(n11066), .A2(n11065), .ZN(n11332) );
  INV_X1 U11275 ( .A(n11333), .ZN(n11330) );
  NAND2_X1 U11276 ( .A1(n11065), .A2(n11066), .ZN(n11333) );
  NAND2_X1 U11277 ( .A1(n11156), .A2(n11334), .ZN(n11066) );
  NAND2_X1 U11278 ( .A1(n11155), .A2(n11157), .ZN(n11334) );
  NAND2_X1 U11279 ( .A1(n11335), .A2(n11336), .ZN(n11157) );
  NAND2_X1 U11280 ( .A1(b_23_), .A2(a_20_), .ZN(n11336) );
  INV_X1 U11281 ( .A(n11337), .ZN(n11335) );
  XOR2_X1 U11282 ( .A(n11338), .B(n11339), .Z(n11155) );
  XNOR2_X1 U11283 ( .A(n11340), .B(n11341), .ZN(n11339) );
  NAND2_X1 U11284 ( .A1(b_22_), .A2(a_21_), .ZN(n11341) );
  NAND2_X1 U11285 ( .A1(a_20_), .A2(n11337), .ZN(n11156) );
  NAND2_X1 U11286 ( .A1(n11342), .A2(n11343), .ZN(n11337) );
  INV_X1 U11287 ( .A(n11344), .ZN(n11343) );
  NOR3_X1 U11288 ( .A1(n8601), .A2(n11345), .A3(n8570), .ZN(n11344) );
  NOR2_X1 U11289 ( .A1(n11078), .A2(n11076), .ZN(n11345) );
  NAND2_X1 U11290 ( .A1(n11076), .A2(n11078), .ZN(n11342) );
  NAND2_X1 U11291 ( .A1(n11152), .A2(n11346), .ZN(n11078) );
  NAND2_X1 U11292 ( .A1(n11151), .A2(n11153), .ZN(n11346) );
  NAND2_X1 U11293 ( .A1(n11347), .A2(n11348), .ZN(n11153) );
  NAND2_X1 U11294 ( .A1(b_23_), .A2(a_22_), .ZN(n11347) );
  XNOR2_X1 U11295 ( .A(n11349), .B(n11350), .ZN(n11151) );
  NAND2_X1 U11296 ( .A1(n11351), .A2(n11352), .ZN(n11349) );
  INV_X1 U11297 ( .A(n11353), .ZN(n11152) );
  NOR2_X1 U11298 ( .A1(n11348), .A2(n8984), .ZN(n11353) );
  NAND2_X1 U11299 ( .A1(n11354), .A2(n11355), .ZN(n11348) );
  NAND2_X1 U11300 ( .A1(n11090), .A2(n11356), .ZN(n11355) );
  NAND2_X1 U11301 ( .A1(n8567), .A2(n11091), .ZN(n11356) );
  XNOR2_X1 U11302 ( .A(n11357), .B(n11358), .ZN(n11090) );
  XOR2_X1 U11303 ( .A(n11359), .B(n11360), .Z(n11357) );
  NAND2_X1 U11304 ( .A1(n11361), .A2(n8961), .ZN(n11354) );
  INV_X1 U11305 ( .A(n8567), .ZN(n8961) );
  NOR2_X1 U11306 ( .A1(n8570), .A2(n8572), .ZN(n8567) );
  INV_X1 U11307 ( .A(n11091), .ZN(n11361) );
  NAND2_X1 U11308 ( .A1(n11362), .A2(n11363), .ZN(n11091) );
  NAND2_X1 U11309 ( .A1(n11098), .A2(n11364), .ZN(n11363) );
  INV_X1 U11310 ( .A(n11365), .ZN(n11364) );
  NOR2_X1 U11311 ( .A1(n11097), .A2(n11096), .ZN(n11365) );
  NOR2_X1 U11312 ( .A1(n8570), .A2(n8982), .ZN(n11098) );
  NAND2_X1 U11313 ( .A1(n11096), .A2(n11097), .ZN(n11362) );
  NAND2_X1 U11314 ( .A1(n11366), .A2(n11367), .ZN(n11097) );
  NAND2_X1 U11315 ( .A1(n11107), .A2(n11368), .ZN(n11367) );
  NAND2_X1 U11316 ( .A1(n11104), .A2(n11106), .ZN(n11368) );
  NOR2_X1 U11317 ( .A1(n8570), .A2(n8541), .ZN(n11107) );
  INV_X1 U11318 ( .A(n11369), .ZN(n11366) );
  NOR2_X1 U11319 ( .A1(n11106), .A2(n11104), .ZN(n11369) );
  XNOR2_X1 U11320 ( .A(n11370), .B(n11371), .ZN(n11104) );
  XNOR2_X1 U11321 ( .A(n11372), .B(n11373), .ZN(n11371) );
  NAND2_X1 U11322 ( .A1(n11374), .A2(n11375), .ZN(n11106) );
  NAND2_X1 U11323 ( .A1(n11112), .A2(n11376), .ZN(n11375) );
  NAND2_X1 U11324 ( .A1(n11115), .A2(n11114), .ZN(n11376) );
  XNOR2_X1 U11325 ( .A(n11377), .B(n11378), .ZN(n11112) );
  XOR2_X1 U11326 ( .A(n11379), .B(n11380), .Z(n11377) );
  INV_X1 U11327 ( .A(n11381), .ZN(n11374) );
  NOR2_X1 U11328 ( .A1(n11114), .A2(n11115), .ZN(n11381) );
  NOR2_X1 U11329 ( .A1(n8570), .A2(n9893), .ZN(n11115) );
  NAND2_X1 U11330 ( .A1(n11382), .A2(n11383), .ZN(n11114) );
  NAND2_X1 U11331 ( .A1(n11122), .A2(n11384), .ZN(n11383) );
  INV_X1 U11332 ( .A(n11385), .ZN(n11384) );
  NOR2_X1 U11333 ( .A1(n11121), .A2(n11120), .ZN(n11385) );
  NOR2_X1 U11334 ( .A1(n8570), .A2(n8512), .ZN(n11122) );
  NAND2_X1 U11335 ( .A1(n11120), .A2(n11121), .ZN(n11382) );
  NAND2_X1 U11336 ( .A1(n11386), .A2(n11387), .ZN(n11121) );
  NAND2_X1 U11337 ( .A1(n11148), .A2(n11388), .ZN(n11387) );
  INV_X1 U11338 ( .A(n11389), .ZN(n11388) );
  NOR2_X1 U11339 ( .A1(n11149), .A2(n11147), .ZN(n11389) );
  NOR2_X1 U11340 ( .A1(n8570), .A2(n8493), .ZN(n11148) );
  NAND2_X1 U11341 ( .A1(n11147), .A2(n11149), .ZN(n11386) );
  NAND2_X1 U11342 ( .A1(n11390), .A2(n11391), .ZN(n11149) );
  NAND2_X1 U11343 ( .A1(n11143), .A2(n11392), .ZN(n11391) );
  INV_X1 U11344 ( .A(n11393), .ZN(n11392) );
  NOR2_X1 U11345 ( .A1(n11144), .A2(n11145), .ZN(n11393) );
  NOR2_X1 U11346 ( .A1(n8570), .A2(n8473), .ZN(n11143) );
  NAND2_X1 U11347 ( .A1(n11145), .A2(n11144), .ZN(n11390) );
  NAND2_X1 U11348 ( .A1(n11394), .A2(n11395), .ZN(n11144) );
  NAND2_X1 U11349 ( .A1(b_21_), .A2(n11396), .ZN(n11395) );
  NAND2_X1 U11350 ( .A1(n8456), .A2(n11397), .ZN(n11396) );
  NAND2_X1 U11351 ( .A1(a_31_), .A2(n8983), .ZN(n11397) );
  NAND2_X1 U11352 ( .A1(b_22_), .A2(n11398), .ZN(n11394) );
  NAND2_X1 U11353 ( .A1(n8459), .A2(n11399), .ZN(n11398) );
  NAND2_X1 U11354 ( .A1(a_30_), .A2(n8599), .ZN(n11399) );
  NOR3_X1 U11355 ( .A1(n8570), .A2(n8979), .A3(n8983), .ZN(n11145) );
  XOR2_X1 U11356 ( .A(n11400), .B(n11401), .Z(n11147) );
  XOR2_X1 U11357 ( .A(n11402), .B(n11403), .Z(n11400) );
  XOR2_X1 U11358 ( .A(n11404), .B(n11405), .Z(n11120) );
  XOR2_X1 U11359 ( .A(n11406), .B(n11407), .Z(n11404) );
  XNOR2_X1 U11360 ( .A(n11408), .B(n11409), .ZN(n11096) );
  XNOR2_X1 U11361 ( .A(n11410), .B(n11411), .ZN(n11409) );
  XNOR2_X1 U11362 ( .A(n11412), .B(n11413), .ZN(n11076) );
  XNOR2_X1 U11363 ( .A(n11414), .B(n11415), .ZN(n11412) );
  XOR2_X1 U11364 ( .A(n11416), .B(n11417), .Z(n11065) );
  XNOR2_X1 U11365 ( .A(n11418), .B(n11419), .ZN(n11417) );
  XNOR2_X1 U11366 ( .A(n11420), .B(n11421), .ZN(n11166) );
  NAND2_X1 U11367 ( .A1(n11422), .A2(n11423), .ZN(n11420) );
  NOR2_X1 U11368 ( .A1(n11173), .A2(n11171), .ZN(n11266) );
  XOR2_X1 U11369 ( .A(n11424), .B(n11425), .Z(n11171) );
  XNOR2_X1 U11370 ( .A(n11426), .B(n11427), .ZN(n11424) );
  NOR2_X1 U11371 ( .A1(n8749), .A2(n8983), .ZN(n11427) );
  NAND2_X1 U11372 ( .A1(b_23_), .A2(a_10_), .ZN(n11173) );
  XNOR2_X1 U11373 ( .A(n11428), .B(n11429), .ZN(n11174) );
  XNOR2_X1 U11374 ( .A(n11430), .B(n11431), .ZN(n11429) );
  XNOR2_X1 U11375 ( .A(n11432), .B(n11433), .ZN(n11187) );
  NAND2_X1 U11376 ( .A1(n11434), .A2(n11435), .ZN(n11432) );
  XNOR2_X1 U11377 ( .A(n11436), .B(n11437), .ZN(n11191) );
  XOR2_X1 U11378 ( .A(n11438), .B(n11439), .Z(n11436) );
  NOR2_X1 U11379 ( .A1(n8848), .A2(n8983), .ZN(n11439) );
  XOR2_X1 U11380 ( .A(n11440), .B(n11441), .Z(n11194) );
  NAND2_X1 U11381 ( .A1(n11442), .A2(n11443), .ZN(n11440) );
  XNOR2_X1 U11382 ( .A(n11444), .B(n11445), .ZN(n11199) );
  XOR2_X1 U11383 ( .A(n11446), .B(n11447), .Z(n11444) );
  XNOR2_X1 U11384 ( .A(n11448), .B(n11449), .ZN(n11202) );
  XNOR2_X1 U11385 ( .A(n11450), .B(n11451), .ZN(n11448) );
  XOR2_X1 U11386 ( .A(n11452), .B(n11453), .Z(n11214) );
  XOR2_X1 U11387 ( .A(n11454), .B(n11455), .Z(n11452) );
  NAND2_X1 U11388 ( .A1(n11456), .A2(n11457), .ZN(n9061) );
  NAND2_X1 U11389 ( .A1(n9186), .A2(n9187), .ZN(n11457) );
  XNOR2_X1 U11390 ( .A(n9180), .B(n9179), .ZN(n11456) );
  NAND3_X1 U11391 ( .A1(n9186), .A2(n9187), .A3(n11458), .ZN(n9062) );
  XNOR2_X1 U11392 ( .A(n9180), .B(n11459), .ZN(n11458) );
  INV_X1 U11393 ( .A(n9179), .ZN(n11459) );
  NAND2_X1 U11394 ( .A1(n11208), .A2(n11460), .ZN(n9187) );
  NAND2_X1 U11395 ( .A1(n11207), .A2(n11209), .ZN(n11460) );
  NAND2_X1 U11396 ( .A1(n11461), .A2(n11462), .ZN(n11209) );
  NAND2_X1 U11397 ( .A1(b_22_), .A2(a_0_), .ZN(n11462) );
  INV_X1 U11398 ( .A(n11463), .ZN(n11461) );
  XNOR2_X1 U11399 ( .A(n11464), .B(n11465), .ZN(n11207) );
  XOR2_X1 U11400 ( .A(n11466), .B(n11467), .Z(n11465) );
  NAND2_X1 U11401 ( .A1(b_21_), .A2(a_1_), .ZN(n11467) );
  NAND2_X1 U11402 ( .A1(a_0_), .A2(n11463), .ZN(n11208) );
  NAND2_X1 U11403 ( .A1(n11468), .A2(n11469), .ZN(n11463) );
  NAND2_X1 U11404 ( .A1(n11455), .A2(n11470), .ZN(n11469) );
  INV_X1 U11405 ( .A(n11471), .ZN(n11470) );
  NOR2_X1 U11406 ( .A1(n11454), .A2(n11453), .ZN(n11471) );
  NOR2_X1 U11407 ( .A1(n8983), .A2(n9731), .ZN(n11455) );
  NAND2_X1 U11408 ( .A1(n11453), .A2(n11454), .ZN(n11468) );
  NAND2_X1 U11409 ( .A1(n11472), .A2(n11473), .ZN(n11454) );
  NAND2_X1 U11410 ( .A1(n11451), .A2(n11474), .ZN(n11473) );
  INV_X1 U11411 ( .A(n11475), .ZN(n11474) );
  NOR2_X1 U11412 ( .A1(n11449), .A2(n11450), .ZN(n11475) );
  NOR2_X1 U11413 ( .A1(n8983), .A2(n8998), .ZN(n11451) );
  NAND2_X1 U11414 ( .A1(n11450), .A2(n11449), .ZN(n11472) );
  XNOR2_X1 U11415 ( .A(n11476), .B(n11477), .ZN(n11449) );
  XOR2_X1 U11416 ( .A(n11478), .B(n11479), .Z(n11477) );
  NAND2_X1 U11417 ( .A1(b_21_), .A2(a_3_), .ZN(n11479) );
  NOR2_X1 U11418 ( .A1(n11480), .A2(n11481), .ZN(n11450) );
  INV_X1 U11419 ( .A(n11482), .ZN(n11481) );
  NAND2_X1 U11420 ( .A1(n11445), .A2(n11483), .ZN(n11482) );
  NAND2_X1 U11421 ( .A1(n11447), .A2(n11446), .ZN(n11483) );
  XNOR2_X1 U11422 ( .A(n11484), .B(n11485), .ZN(n11445) );
  XOR2_X1 U11423 ( .A(n11486), .B(n11487), .Z(n11484) );
  NOR2_X1 U11424 ( .A1(n8996), .A2(n8599), .ZN(n11487) );
  NOR2_X1 U11425 ( .A1(n11446), .A2(n11447), .ZN(n11480) );
  NOR2_X1 U11426 ( .A1(n8983), .A2(n8877), .ZN(n11447) );
  NAND2_X1 U11427 ( .A1(n11442), .A2(n11488), .ZN(n11446) );
  NAND2_X1 U11428 ( .A1(n11441), .A2(n11443), .ZN(n11488) );
  NAND2_X1 U11429 ( .A1(n11489), .A2(n11490), .ZN(n11443) );
  NAND2_X1 U11430 ( .A1(b_22_), .A2(a_4_), .ZN(n11490) );
  INV_X1 U11431 ( .A(n11491), .ZN(n11489) );
  XNOR2_X1 U11432 ( .A(n11492), .B(n11493), .ZN(n11441) );
  XOR2_X1 U11433 ( .A(n11494), .B(n11495), .Z(n11493) );
  NAND2_X1 U11434 ( .A1(b_21_), .A2(a_5_), .ZN(n11495) );
  NAND2_X1 U11435 ( .A1(a_4_), .A2(n11491), .ZN(n11442) );
  NAND2_X1 U11436 ( .A1(n11496), .A2(n11497), .ZN(n11491) );
  INV_X1 U11437 ( .A(n11498), .ZN(n11497) );
  NOR3_X1 U11438 ( .A1(n8848), .A2(n11499), .A3(n8983), .ZN(n11498) );
  NOR2_X1 U11439 ( .A1(n11437), .A2(n11438), .ZN(n11499) );
  NAND2_X1 U11440 ( .A1(n11437), .A2(n11438), .ZN(n11496) );
  NAND2_X1 U11441 ( .A1(n11434), .A2(n11500), .ZN(n11438) );
  NAND2_X1 U11442 ( .A1(n11433), .A2(n11435), .ZN(n11500) );
  NAND2_X1 U11443 ( .A1(n11501), .A2(n11502), .ZN(n11435) );
  NAND2_X1 U11444 ( .A1(b_22_), .A2(a_6_), .ZN(n11502) );
  INV_X1 U11445 ( .A(n11503), .ZN(n11501) );
  XOR2_X1 U11446 ( .A(n11504), .B(n11505), .Z(n11433) );
  XOR2_X1 U11447 ( .A(n11506), .B(n11507), .Z(n11504) );
  NOR2_X1 U11448 ( .A1(n8817), .A2(n8599), .ZN(n11507) );
  NAND2_X1 U11449 ( .A1(a_6_), .A2(n11503), .ZN(n11434) );
  NAND2_X1 U11450 ( .A1(n11508), .A2(n11509), .ZN(n11503) );
  INV_X1 U11451 ( .A(n11510), .ZN(n11509) );
  NOR3_X1 U11452 ( .A1(n8817), .A2(n11511), .A3(n8983), .ZN(n11510) );
  NOR2_X1 U11453 ( .A1(n11242), .A2(n11243), .ZN(n11511) );
  NAND2_X1 U11454 ( .A1(n11242), .A2(n11243), .ZN(n11508) );
  NAND2_X1 U11455 ( .A1(n11512), .A2(n11513), .ZN(n11243) );
  NAND3_X1 U11456 ( .A1(a_8_), .A2(n11514), .A3(b_22_), .ZN(n11513) );
  INV_X1 U11457 ( .A(n11515), .ZN(n11514) );
  NOR2_X1 U11458 ( .A1(n11250), .A2(n11252), .ZN(n11515) );
  NAND2_X1 U11459 ( .A1(n11250), .A2(n11252), .ZN(n11512) );
  NAND2_X1 U11460 ( .A1(n11260), .A2(n11516), .ZN(n11252) );
  NAND2_X1 U11461 ( .A1(n11259), .A2(n11261), .ZN(n11516) );
  NAND2_X1 U11462 ( .A1(n11517), .A2(n11518), .ZN(n11261) );
  NAND2_X1 U11463 ( .A1(b_22_), .A2(a_9_), .ZN(n11517) );
  XNOR2_X1 U11464 ( .A(n11519), .B(n11520), .ZN(n11259) );
  XNOR2_X1 U11465 ( .A(n11521), .B(n11522), .ZN(n11519) );
  NAND2_X1 U11466 ( .A1(n11523), .A2(a_9_), .ZN(n11260) );
  INV_X1 U11467 ( .A(n11518), .ZN(n11523) );
  NAND2_X1 U11468 ( .A1(n11524), .A2(n11525), .ZN(n11518) );
  NAND2_X1 U11469 ( .A1(n11428), .A2(n11526), .ZN(n11525) );
  NAND2_X1 U11470 ( .A1(n11431), .A2(n11430), .ZN(n11526) );
  XOR2_X1 U11471 ( .A(n11527), .B(n11528), .Z(n11428) );
  XNOR2_X1 U11472 ( .A(n11529), .B(n11530), .ZN(n11528) );
  INV_X1 U11473 ( .A(n11531), .ZN(n11524) );
  NOR2_X1 U11474 ( .A1(n11430), .A2(n11431), .ZN(n11531) );
  NOR2_X1 U11475 ( .A1(n8983), .A2(n8769), .ZN(n11431) );
  NAND2_X1 U11476 ( .A1(n11532), .A2(n11533), .ZN(n11430) );
  NAND3_X1 U11477 ( .A1(a_11_), .A2(n11534), .A3(b_22_), .ZN(n11533) );
  NAND2_X1 U11478 ( .A1(n11425), .A2(n11426), .ZN(n11534) );
  INV_X1 U11479 ( .A(n11535), .ZN(n11532) );
  NOR2_X1 U11480 ( .A1(n11425), .A2(n11426), .ZN(n11535) );
  NOR2_X1 U11481 ( .A1(n11536), .A2(n11537), .ZN(n11426) );
  INV_X1 U11482 ( .A(n11538), .ZN(n11537) );
  NAND3_X1 U11483 ( .A1(a_12_), .A2(n11539), .A3(b_22_), .ZN(n11538) );
  NAND2_X1 U11484 ( .A1(n11276), .A2(n11275), .ZN(n11539) );
  NOR2_X1 U11485 ( .A1(n11275), .A2(n11276), .ZN(n11536) );
  NOR2_X1 U11486 ( .A1(n11540), .A2(n11541), .ZN(n11276) );
  NOR3_X1 U11487 ( .A1(n8721), .A2(n11542), .A3(n8983), .ZN(n11541) );
  NOR2_X1 U11488 ( .A1(n11284), .A2(n11282), .ZN(n11542) );
  INV_X1 U11489 ( .A(n11543), .ZN(n11540) );
  NAND2_X1 U11490 ( .A1(n11282), .A2(n11284), .ZN(n11543) );
  NAND2_X1 U11491 ( .A1(n11422), .A2(n11544), .ZN(n11284) );
  NAND2_X1 U11492 ( .A1(n11421), .A2(n11423), .ZN(n11544) );
  NAND2_X1 U11493 ( .A1(n11545), .A2(n11546), .ZN(n11423) );
  NAND2_X1 U11494 ( .A1(b_22_), .A2(a_14_), .ZN(n11546) );
  INV_X1 U11495 ( .A(n11547), .ZN(n11545) );
  XOR2_X1 U11496 ( .A(n11548), .B(n11549), .Z(n11421) );
  XOR2_X1 U11497 ( .A(n11550), .B(n11551), .Z(n11548) );
  NOR2_X1 U11498 ( .A1(n8692), .A2(n8599), .ZN(n11551) );
  NAND2_X1 U11499 ( .A1(a_14_), .A2(n11547), .ZN(n11422) );
  NAND2_X1 U11500 ( .A1(n11552), .A2(n11553), .ZN(n11547) );
  INV_X1 U11501 ( .A(n11554), .ZN(n11553) );
  NOR3_X1 U11502 ( .A1(n8692), .A2(n11555), .A3(n8983), .ZN(n11554) );
  NOR2_X1 U11503 ( .A1(n11295), .A2(n11294), .ZN(n11555) );
  NAND2_X1 U11504 ( .A1(n11294), .A2(n11295), .ZN(n11552) );
  NAND2_X1 U11505 ( .A1(n11304), .A2(n11556), .ZN(n11295) );
  NAND2_X1 U11506 ( .A1(n11303), .A2(n11305), .ZN(n11556) );
  NAND2_X1 U11507 ( .A1(n11557), .A2(n11558), .ZN(n11305) );
  NAND2_X1 U11508 ( .A1(b_22_), .A2(a_16_), .ZN(n11558) );
  INV_X1 U11509 ( .A(n11559), .ZN(n11557) );
  XNOR2_X1 U11510 ( .A(n11560), .B(n11561), .ZN(n11303) );
  XOR2_X1 U11511 ( .A(n11562), .B(n11563), .Z(n11561) );
  NAND2_X1 U11512 ( .A1(b_21_), .A2(a_17_), .ZN(n11563) );
  NAND2_X1 U11513 ( .A1(a_16_), .A2(n11559), .ZN(n11304) );
  NAND2_X1 U11514 ( .A1(n11564), .A2(n11565), .ZN(n11559) );
  INV_X1 U11515 ( .A(n11566), .ZN(n11565) );
  NOR3_X1 U11516 ( .A1(n8662), .A2(n11567), .A3(n8983), .ZN(n11566) );
  NOR2_X1 U11517 ( .A1(n11311), .A2(n11312), .ZN(n11567) );
  NAND2_X1 U11518 ( .A1(n11312), .A2(n11311), .ZN(n11564) );
  XOR2_X1 U11519 ( .A(n11568), .B(n11569), .Z(n11311) );
  XNOR2_X1 U11520 ( .A(n11570), .B(n11571), .ZN(n11569) );
  NOR2_X1 U11521 ( .A1(n11572), .A2(n11573), .ZN(n11312) );
  INV_X1 U11522 ( .A(n11574), .ZN(n11573) );
  NAND2_X1 U11523 ( .A1(n11319), .A2(n11575), .ZN(n11574) );
  NAND2_X1 U11524 ( .A1(n11321), .A2(n11320), .ZN(n11575) );
  XOR2_X1 U11525 ( .A(n11576), .B(n11577), .Z(n11319) );
  XOR2_X1 U11526 ( .A(n11578), .B(n11579), .Z(n11577) );
  NAND2_X1 U11527 ( .A1(b_21_), .A2(a_19_), .ZN(n11579) );
  NOR2_X1 U11528 ( .A1(n11320), .A2(n11321), .ZN(n11572) );
  NOR2_X1 U11529 ( .A1(n8983), .A2(n8988), .ZN(n11321) );
  NAND2_X1 U11530 ( .A1(n11580), .A2(n11581), .ZN(n11320) );
  NAND2_X1 U11531 ( .A1(n11329), .A2(n11582), .ZN(n11581) );
  NAND2_X1 U11532 ( .A1(n11326), .A2(n11328), .ZN(n11582) );
  NOR2_X1 U11533 ( .A1(n8983), .A2(n8630), .ZN(n11329) );
  INV_X1 U11534 ( .A(n11583), .ZN(n11580) );
  NOR2_X1 U11535 ( .A1(n11328), .A2(n11326), .ZN(n11583) );
  XOR2_X1 U11536 ( .A(n11584), .B(n11585), .Z(n11326) );
  NAND2_X1 U11537 ( .A1(n11586), .A2(n11587), .ZN(n11584) );
  NAND2_X1 U11538 ( .A1(n11588), .A2(n11589), .ZN(n11328) );
  NAND2_X1 U11539 ( .A1(n11416), .A2(n11590), .ZN(n11589) );
  NAND2_X1 U11540 ( .A1(n11419), .A2(n11418), .ZN(n11590) );
  XOR2_X1 U11541 ( .A(n11591), .B(n11592), .Z(n11416) );
  XNOR2_X1 U11542 ( .A(n8596), .B(n11593), .ZN(n11592) );
  INV_X1 U11543 ( .A(n11594), .ZN(n11588) );
  NOR2_X1 U11544 ( .A1(n11418), .A2(n11419), .ZN(n11594) );
  NOR2_X1 U11545 ( .A1(n8983), .A2(n8986), .ZN(n11419) );
  NAND2_X1 U11546 ( .A1(n11595), .A2(n11596), .ZN(n11418) );
  NAND3_X1 U11547 ( .A1(a_21_), .A2(n11597), .A3(b_22_), .ZN(n11596) );
  NAND2_X1 U11548 ( .A1(n11340), .A2(n11338), .ZN(n11597) );
  INV_X1 U11549 ( .A(n11598), .ZN(n11595) );
  NOR2_X1 U11550 ( .A1(n11338), .A2(n11340), .ZN(n11598) );
  NOR2_X1 U11551 ( .A1(n11599), .A2(n11600), .ZN(n11340) );
  NOR2_X1 U11552 ( .A1(n11413), .A2(n11601), .ZN(n11600) );
  NOR2_X1 U11553 ( .A1(n11602), .A2(n11415), .ZN(n11601) );
  INV_X1 U11554 ( .A(n8584), .ZN(n11415) );
  XOR2_X1 U11555 ( .A(n11603), .B(n11604), .Z(n11413) );
  NAND2_X1 U11556 ( .A1(n11605), .A2(n11606), .ZN(n11603) );
  NOR2_X1 U11557 ( .A1(n8584), .A2(n11414), .ZN(n11599) );
  INV_X1 U11558 ( .A(n11602), .ZN(n11414) );
  NAND2_X1 U11559 ( .A1(n11351), .A2(n11607), .ZN(n11602) );
  NAND2_X1 U11560 ( .A1(n11350), .A2(n11352), .ZN(n11607) );
  NAND2_X1 U11561 ( .A1(n11608), .A2(n11609), .ZN(n11352) );
  NAND2_X1 U11562 ( .A1(b_22_), .A2(a_23_), .ZN(n11609) );
  INV_X1 U11563 ( .A(n11610), .ZN(n11608) );
  XOR2_X1 U11564 ( .A(n11611), .B(n11612), .Z(n11350) );
  XOR2_X1 U11565 ( .A(n11613), .B(n11614), .Z(n11611) );
  NAND2_X1 U11566 ( .A1(a_23_), .A2(n11610), .ZN(n11351) );
  NAND2_X1 U11567 ( .A1(n11615), .A2(n11616), .ZN(n11610) );
  NAND2_X1 U11568 ( .A1(n11360), .A2(n11617), .ZN(n11616) );
  INV_X1 U11569 ( .A(n11618), .ZN(n11617) );
  NOR2_X1 U11570 ( .A1(n11359), .A2(n11358), .ZN(n11618) );
  NOR2_X1 U11571 ( .A1(n8983), .A2(n8982), .ZN(n11360) );
  NAND2_X1 U11572 ( .A1(n11358), .A2(n11359), .ZN(n11615) );
  NAND2_X1 U11573 ( .A1(n11619), .A2(n11620), .ZN(n11359) );
  NAND2_X1 U11574 ( .A1(n11411), .A2(n11621), .ZN(n11620) );
  NAND2_X1 U11575 ( .A1(n11408), .A2(n11410), .ZN(n11621) );
  NOR2_X1 U11576 ( .A1(n8983), .A2(n8541), .ZN(n11411) );
  INV_X1 U11577 ( .A(n11622), .ZN(n11619) );
  NOR2_X1 U11578 ( .A1(n11410), .A2(n11408), .ZN(n11622) );
  XNOR2_X1 U11579 ( .A(n11623), .B(n11624), .ZN(n11408) );
  XNOR2_X1 U11580 ( .A(n11625), .B(n11626), .ZN(n11624) );
  NAND2_X1 U11581 ( .A1(n11627), .A2(n11628), .ZN(n11410) );
  NAND2_X1 U11582 ( .A1(n11370), .A2(n11629), .ZN(n11628) );
  NAND2_X1 U11583 ( .A1(n11373), .A2(n11372), .ZN(n11629) );
  XNOR2_X1 U11584 ( .A(n11630), .B(n11631), .ZN(n11370) );
  XOR2_X1 U11585 ( .A(n11632), .B(n11633), .Z(n11630) );
  INV_X1 U11586 ( .A(n11634), .ZN(n11627) );
  NOR2_X1 U11587 ( .A1(n11372), .A2(n11373), .ZN(n11634) );
  NOR2_X1 U11588 ( .A1(n8983), .A2(n9893), .ZN(n11373) );
  NAND2_X1 U11589 ( .A1(n11635), .A2(n11636), .ZN(n11372) );
  NAND2_X1 U11590 ( .A1(n11380), .A2(n11637), .ZN(n11636) );
  INV_X1 U11591 ( .A(n11638), .ZN(n11637) );
  NOR2_X1 U11592 ( .A1(n11379), .A2(n11378), .ZN(n11638) );
  NOR2_X1 U11593 ( .A1(n8983), .A2(n8512), .ZN(n11380) );
  NAND2_X1 U11594 ( .A1(n11378), .A2(n11379), .ZN(n11635) );
  NAND2_X1 U11595 ( .A1(n11639), .A2(n11640), .ZN(n11379) );
  NAND2_X1 U11596 ( .A1(n11406), .A2(n11641), .ZN(n11640) );
  INV_X1 U11597 ( .A(n11642), .ZN(n11641) );
  NOR2_X1 U11598 ( .A1(n11407), .A2(n11405), .ZN(n11642) );
  NOR2_X1 U11599 ( .A1(n8983), .A2(n8493), .ZN(n11406) );
  NAND2_X1 U11600 ( .A1(n11405), .A2(n11407), .ZN(n11639) );
  NAND2_X1 U11601 ( .A1(n11643), .A2(n11644), .ZN(n11407) );
  NAND2_X1 U11602 ( .A1(n11401), .A2(n11645), .ZN(n11644) );
  INV_X1 U11603 ( .A(n11646), .ZN(n11645) );
  NOR2_X1 U11604 ( .A1(n11402), .A2(n11403), .ZN(n11646) );
  NOR2_X1 U11605 ( .A1(n8983), .A2(n8473), .ZN(n11401) );
  NAND2_X1 U11606 ( .A1(n11403), .A2(n11402), .ZN(n11643) );
  NAND2_X1 U11607 ( .A1(n11647), .A2(n11648), .ZN(n11402) );
  NAND2_X1 U11608 ( .A1(b_20_), .A2(n11649), .ZN(n11648) );
  NAND2_X1 U11609 ( .A1(n8456), .A2(n11650), .ZN(n11649) );
  NAND2_X1 U11610 ( .A1(a_31_), .A2(n8599), .ZN(n11650) );
  NAND2_X1 U11611 ( .A1(b_21_), .A2(n11651), .ZN(n11647) );
  NAND2_X1 U11612 ( .A1(n8459), .A2(n11652), .ZN(n11651) );
  NAND2_X1 U11613 ( .A1(a_30_), .A2(n8985), .ZN(n11652) );
  NOR3_X1 U11614 ( .A1(n8599), .A2(n8979), .A3(n8983), .ZN(n11403) );
  XOR2_X1 U11615 ( .A(n11653), .B(n11654), .Z(n11405) );
  XOR2_X1 U11616 ( .A(n11655), .B(n11656), .Z(n11653) );
  XOR2_X1 U11617 ( .A(n11657), .B(n11658), .Z(n11378) );
  XOR2_X1 U11618 ( .A(n11659), .B(n11660), .Z(n11657) );
  XNOR2_X1 U11619 ( .A(n11661), .B(n11662), .ZN(n11358) );
  XNOR2_X1 U11620 ( .A(n11663), .B(n11664), .ZN(n11662) );
  NAND2_X1 U11621 ( .A1(b_22_), .A2(a_22_), .ZN(n8584) );
  XOR2_X1 U11622 ( .A(n11665), .B(n11666), .Z(n11338) );
  NAND2_X1 U11623 ( .A1(n11667), .A2(n11668), .ZN(n11665) );
  XNOR2_X1 U11624 ( .A(n11669), .B(n11670), .ZN(n11294) );
  NAND2_X1 U11625 ( .A1(n11671), .A2(n11672), .ZN(n11669) );
  XNOR2_X1 U11626 ( .A(n11673), .B(n11674), .ZN(n11282) );
  XOR2_X1 U11627 ( .A(n11675), .B(n11676), .Z(n11674) );
  NAND2_X1 U11628 ( .A1(b_21_), .A2(a_14_), .ZN(n11676) );
  XOR2_X1 U11629 ( .A(n11677), .B(n11678), .Z(n11275) );
  NAND2_X1 U11630 ( .A1(n11679), .A2(n11680), .ZN(n11677) );
  XOR2_X1 U11631 ( .A(n11681), .B(n11682), .Z(n11425) );
  XOR2_X1 U11632 ( .A(n11683), .B(n11684), .Z(n11681) );
  XNOR2_X1 U11633 ( .A(n11685), .B(n11686), .ZN(n11250) );
  XNOR2_X1 U11634 ( .A(n11687), .B(n11688), .ZN(n11685) );
  XOR2_X1 U11635 ( .A(n11689), .B(n11690), .Z(n11242) );
  XNOR2_X1 U11636 ( .A(n11691), .B(n11692), .ZN(n11690) );
  NAND2_X1 U11637 ( .A1(b_21_), .A2(a_8_), .ZN(n11692) );
  XNOR2_X1 U11638 ( .A(n11693), .B(n11694), .ZN(n11437) );
  XOR2_X1 U11639 ( .A(n11695), .B(n11696), .Z(n11694) );
  NAND2_X1 U11640 ( .A1(b_21_), .A2(a_6_), .ZN(n11696) );
  XNOR2_X1 U11641 ( .A(n11697), .B(n11698), .ZN(n11453) );
  XOR2_X1 U11642 ( .A(n11699), .B(n11700), .Z(n11698) );
  NAND2_X1 U11643 ( .A1(b_21_), .A2(a_2_), .ZN(n11700) );
  XOR2_X1 U11644 ( .A(n11701), .B(n11702), .Z(n9186) );
  XOR2_X1 U11645 ( .A(n11703), .B(n11704), .Z(n11701) );
  NOR2_X1 U11646 ( .A1(n9471), .A2(n8599), .ZN(n11704) );
  NAND3_X1 U11647 ( .A1(n9179), .A2(n9180), .A3(n11705), .ZN(n9067) );
  XOR2_X1 U11648 ( .A(n9175), .B(n9174), .Z(n11705) );
  NAND2_X1 U11649 ( .A1(n11706), .A2(n11707), .ZN(n9180) );
  INV_X1 U11650 ( .A(n11708), .ZN(n11707) );
  NOR3_X1 U11651 ( .A1(n9471), .A2(n11709), .A3(n8599), .ZN(n11708) );
  NOR2_X1 U11652 ( .A1(n11703), .A2(n11702), .ZN(n11709) );
  NAND2_X1 U11653 ( .A1(n11702), .A2(n11703), .ZN(n11706) );
  NAND2_X1 U11654 ( .A1(n11710), .A2(n11711), .ZN(n11703) );
  NAND3_X1 U11655 ( .A1(a_1_), .A2(n11712), .A3(b_21_), .ZN(n11711) );
  INV_X1 U11656 ( .A(n11713), .ZN(n11712) );
  NOR2_X1 U11657 ( .A1(n11466), .A2(n11464), .ZN(n11713) );
  NAND2_X1 U11658 ( .A1(n11464), .A2(n11466), .ZN(n11710) );
  NAND2_X1 U11659 ( .A1(n11714), .A2(n11715), .ZN(n11466) );
  NAND3_X1 U11660 ( .A1(a_2_), .A2(n11716), .A3(b_21_), .ZN(n11715) );
  INV_X1 U11661 ( .A(n11717), .ZN(n11716) );
  NOR2_X1 U11662 ( .A1(n11699), .A2(n11697), .ZN(n11717) );
  NAND2_X1 U11663 ( .A1(n11697), .A2(n11699), .ZN(n11714) );
  NAND2_X1 U11664 ( .A1(n11718), .A2(n11719), .ZN(n11699) );
  NAND3_X1 U11665 ( .A1(a_3_), .A2(n11720), .A3(b_21_), .ZN(n11719) );
  INV_X1 U11666 ( .A(n11721), .ZN(n11720) );
  NOR2_X1 U11667 ( .A1(n11478), .A2(n11476), .ZN(n11721) );
  NAND2_X1 U11668 ( .A1(n11476), .A2(n11478), .ZN(n11718) );
  NAND2_X1 U11669 ( .A1(n11722), .A2(n11723), .ZN(n11478) );
  NAND3_X1 U11670 ( .A1(a_4_), .A2(n11724), .A3(b_21_), .ZN(n11723) );
  INV_X1 U11671 ( .A(n11725), .ZN(n11724) );
  NOR2_X1 U11672 ( .A1(n11486), .A2(n11485), .ZN(n11725) );
  NAND2_X1 U11673 ( .A1(n11485), .A2(n11486), .ZN(n11722) );
  NAND2_X1 U11674 ( .A1(n11726), .A2(n11727), .ZN(n11486) );
  NAND3_X1 U11675 ( .A1(a_5_), .A2(n11728), .A3(b_21_), .ZN(n11727) );
  INV_X1 U11676 ( .A(n11729), .ZN(n11728) );
  NOR2_X1 U11677 ( .A1(n11494), .A2(n11492), .ZN(n11729) );
  NAND2_X1 U11678 ( .A1(n11492), .A2(n11494), .ZN(n11726) );
  NAND2_X1 U11679 ( .A1(n11730), .A2(n11731), .ZN(n11494) );
  INV_X1 U11680 ( .A(n11732), .ZN(n11731) );
  NOR3_X1 U11681 ( .A1(n8994), .A2(n11733), .A3(n8599), .ZN(n11732) );
  NOR2_X1 U11682 ( .A1(n11695), .A2(n11693), .ZN(n11733) );
  NAND2_X1 U11683 ( .A1(n11693), .A2(n11695), .ZN(n11730) );
  NAND2_X1 U11684 ( .A1(n11734), .A2(n11735), .ZN(n11695) );
  NAND3_X1 U11685 ( .A1(a_7_), .A2(n11736), .A3(b_21_), .ZN(n11735) );
  INV_X1 U11686 ( .A(n11737), .ZN(n11736) );
  NOR2_X1 U11687 ( .A1(n11506), .A2(n11505), .ZN(n11737) );
  NAND2_X1 U11688 ( .A1(n11505), .A2(n11506), .ZN(n11734) );
  NAND2_X1 U11689 ( .A1(n11738), .A2(n11739), .ZN(n11506) );
  NAND3_X1 U11690 ( .A1(a_8_), .A2(n11740), .A3(b_21_), .ZN(n11739) );
  NAND2_X1 U11691 ( .A1(n11691), .A2(n11689), .ZN(n11740) );
  NAND2_X1 U11692 ( .A1(n11741), .A2(n11742), .ZN(n11738) );
  INV_X1 U11693 ( .A(n11691), .ZN(n11742) );
  NOR2_X1 U11694 ( .A1(n11743), .A2(n11744), .ZN(n11691) );
  INV_X1 U11695 ( .A(n11745), .ZN(n11744) );
  NAND2_X1 U11696 ( .A1(n11688), .A2(n11746), .ZN(n11745) );
  NAND2_X1 U11697 ( .A1(n11687), .A2(n11686), .ZN(n11746) );
  NOR2_X1 U11698 ( .A1(n8599), .A2(n8779), .ZN(n11688) );
  NOR2_X1 U11699 ( .A1(n11686), .A2(n11687), .ZN(n11743) );
  NOR2_X1 U11700 ( .A1(n11747), .A2(n11748), .ZN(n11687) );
  INV_X1 U11701 ( .A(n11749), .ZN(n11748) );
  NAND2_X1 U11702 ( .A1(n11522), .A2(n11750), .ZN(n11749) );
  NAND2_X1 U11703 ( .A1(n11521), .A2(n11520), .ZN(n11750) );
  NOR2_X1 U11704 ( .A1(n8599), .A2(n8769), .ZN(n11522) );
  NOR2_X1 U11705 ( .A1(n11520), .A2(n11521), .ZN(n11747) );
  NOR2_X1 U11706 ( .A1(n11751), .A2(n11752), .ZN(n11521) );
  INV_X1 U11707 ( .A(n11753), .ZN(n11752) );
  NAND2_X1 U11708 ( .A1(n11530), .A2(n11754), .ZN(n11753) );
  NAND2_X1 U11709 ( .A1(n11527), .A2(n11529), .ZN(n11754) );
  NOR2_X1 U11710 ( .A1(n8599), .A2(n8749), .ZN(n11530) );
  NOR2_X1 U11711 ( .A1(n11529), .A2(n11527), .ZN(n11751) );
  XOR2_X1 U11712 ( .A(n11755), .B(n11756), .Z(n11527) );
  XOR2_X1 U11713 ( .A(n11757), .B(n11758), .Z(n11755) );
  NAND2_X1 U11714 ( .A1(n11759), .A2(n11760), .ZN(n11529) );
  NAND2_X1 U11715 ( .A1(n11682), .A2(n11761), .ZN(n11760) );
  NAND2_X1 U11716 ( .A1(n11684), .A2(n11683), .ZN(n11761) );
  XOR2_X1 U11717 ( .A(n11762), .B(n11763), .Z(n11682) );
  NAND2_X1 U11718 ( .A1(n11764), .A2(n11765), .ZN(n11762) );
  INV_X1 U11719 ( .A(n11766), .ZN(n11759) );
  NOR2_X1 U11720 ( .A1(n11683), .A2(n11684), .ZN(n11766) );
  NOR2_X1 U11721 ( .A1(n8599), .A2(n8739), .ZN(n11684) );
  NAND2_X1 U11722 ( .A1(n11679), .A2(n11767), .ZN(n11683) );
  NAND2_X1 U11723 ( .A1(n11678), .A2(n11680), .ZN(n11767) );
  NAND2_X1 U11724 ( .A1(n11768), .A2(n11769), .ZN(n11680) );
  NAND2_X1 U11725 ( .A1(b_21_), .A2(a_13_), .ZN(n11769) );
  XOR2_X1 U11726 ( .A(n11770), .B(n11771), .Z(n11678) );
  XNOR2_X1 U11727 ( .A(n11772), .B(n11773), .ZN(n11771) );
  INV_X1 U11728 ( .A(n11774), .ZN(n11679) );
  NOR2_X1 U11729 ( .A1(n8721), .A2(n11768), .ZN(n11774) );
  NOR2_X1 U11730 ( .A1(n11775), .A2(n11776), .ZN(n11768) );
  NOR3_X1 U11731 ( .A1(n8991), .A2(n11777), .A3(n8599), .ZN(n11776) );
  NOR2_X1 U11732 ( .A1(n11675), .A2(n11673), .ZN(n11777) );
  INV_X1 U11733 ( .A(n11778), .ZN(n11775) );
  NAND2_X1 U11734 ( .A1(n11673), .A2(n11675), .ZN(n11778) );
  NAND2_X1 U11735 ( .A1(n11779), .A2(n11780), .ZN(n11675) );
  NAND3_X1 U11736 ( .A1(a_15_), .A2(n11781), .A3(b_21_), .ZN(n11780) );
  INV_X1 U11737 ( .A(n11782), .ZN(n11781) );
  NOR2_X1 U11738 ( .A1(n11550), .A2(n11549), .ZN(n11782) );
  NAND2_X1 U11739 ( .A1(n11549), .A2(n11550), .ZN(n11779) );
  NAND2_X1 U11740 ( .A1(n11671), .A2(n11783), .ZN(n11550) );
  NAND2_X1 U11741 ( .A1(n11670), .A2(n11672), .ZN(n11783) );
  NAND2_X1 U11742 ( .A1(n11784), .A2(n11785), .ZN(n11672) );
  NAND2_X1 U11743 ( .A1(b_21_), .A2(a_16_), .ZN(n11785) );
  XNOR2_X1 U11744 ( .A(n11786), .B(n11787), .ZN(n11670) );
  XOR2_X1 U11745 ( .A(n11788), .B(n11789), .Z(n11787) );
  NAND2_X1 U11746 ( .A1(b_20_), .A2(a_17_), .ZN(n11789) );
  NAND2_X1 U11747 ( .A1(a_16_), .A2(n11790), .ZN(n11671) );
  INV_X1 U11748 ( .A(n11784), .ZN(n11790) );
  NOR2_X1 U11749 ( .A1(n11791), .A2(n11792), .ZN(n11784) );
  NOR3_X1 U11750 ( .A1(n8662), .A2(n11793), .A3(n8599), .ZN(n11792) );
  INV_X1 U11751 ( .A(n11794), .ZN(n11793) );
  NAND2_X1 U11752 ( .A1(n11560), .A2(n11562), .ZN(n11794) );
  NOR2_X1 U11753 ( .A1(n11562), .A2(n11560), .ZN(n11791) );
  XNOR2_X1 U11754 ( .A(n11795), .B(n11796), .ZN(n11560) );
  XNOR2_X1 U11755 ( .A(n11797), .B(n11798), .ZN(n11796) );
  NAND2_X1 U11756 ( .A1(n11799), .A2(n11800), .ZN(n11562) );
  NAND2_X1 U11757 ( .A1(n11568), .A2(n11801), .ZN(n11800) );
  NAND2_X1 U11758 ( .A1(n11571), .A2(n11570), .ZN(n11801) );
  XOR2_X1 U11759 ( .A(n11802), .B(n11803), .Z(n11568) );
  XOR2_X1 U11760 ( .A(n11804), .B(n11805), .Z(n11803) );
  NAND2_X1 U11761 ( .A1(b_20_), .A2(a_19_), .ZN(n11805) );
  INV_X1 U11762 ( .A(n11806), .ZN(n11799) );
  NOR2_X1 U11763 ( .A1(n11570), .A2(n11571), .ZN(n11806) );
  NOR2_X1 U11764 ( .A1(n8599), .A2(n8988), .ZN(n11571) );
  NAND2_X1 U11765 ( .A1(n11807), .A2(n11808), .ZN(n11570) );
  NAND3_X1 U11766 ( .A1(a_19_), .A2(n11809), .A3(b_21_), .ZN(n11808) );
  INV_X1 U11767 ( .A(n11810), .ZN(n11809) );
  NOR2_X1 U11768 ( .A1(n11578), .A2(n11576), .ZN(n11810) );
  NAND2_X1 U11769 ( .A1(n11576), .A2(n11578), .ZN(n11807) );
  NAND2_X1 U11770 ( .A1(n11586), .A2(n11811), .ZN(n11578) );
  NAND2_X1 U11771 ( .A1(n11585), .A2(n11587), .ZN(n11811) );
  NAND2_X1 U11772 ( .A1(n11812), .A2(n11813), .ZN(n11587) );
  NAND2_X1 U11773 ( .A1(b_21_), .A2(a_20_), .ZN(n11813) );
  INV_X1 U11774 ( .A(n11814), .ZN(n11812) );
  XNOR2_X1 U11775 ( .A(n11815), .B(n11816), .ZN(n11585) );
  XOR2_X1 U11776 ( .A(n11817), .B(n11818), .Z(n11816) );
  NAND2_X1 U11777 ( .A1(b_20_), .A2(a_21_), .ZN(n11818) );
  NAND2_X1 U11778 ( .A1(a_20_), .A2(n11814), .ZN(n11586) );
  NAND2_X1 U11779 ( .A1(n11819), .A2(n11820), .ZN(n11814) );
  NAND2_X1 U11780 ( .A1(n11591), .A2(n11821), .ZN(n11820) );
  INV_X1 U11781 ( .A(n11822), .ZN(n11821) );
  NOR2_X1 U11782 ( .A1(n11593), .A2(n8596), .ZN(n11822) );
  XNOR2_X1 U11783 ( .A(n11823), .B(n11824), .ZN(n11591) );
  NAND2_X1 U11784 ( .A1(n11825), .A2(n11826), .ZN(n11823) );
  NAND2_X1 U11785 ( .A1(n8596), .A2(n11593), .ZN(n11819) );
  NAND2_X1 U11786 ( .A1(n11667), .A2(n11827), .ZN(n11593) );
  NAND2_X1 U11787 ( .A1(n11666), .A2(n11668), .ZN(n11827) );
  NAND2_X1 U11788 ( .A1(n11828), .A2(n11829), .ZN(n11668) );
  NAND2_X1 U11789 ( .A1(b_21_), .A2(a_22_), .ZN(n11829) );
  INV_X1 U11790 ( .A(n11830), .ZN(n11828) );
  XNOR2_X1 U11791 ( .A(n11831), .B(n11832), .ZN(n11666) );
  NAND2_X1 U11792 ( .A1(n11833), .A2(n11834), .ZN(n11831) );
  NAND2_X1 U11793 ( .A1(a_22_), .A2(n11830), .ZN(n11667) );
  NAND2_X1 U11794 ( .A1(n11605), .A2(n11835), .ZN(n11830) );
  NAND2_X1 U11795 ( .A1(n11604), .A2(n11606), .ZN(n11835) );
  NAND2_X1 U11796 ( .A1(n11836), .A2(n11837), .ZN(n11606) );
  NAND2_X1 U11797 ( .A1(b_21_), .A2(a_23_), .ZN(n11837) );
  INV_X1 U11798 ( .A(n11838), .ZN(n11836) );
  XOR2_X1 U11799 ( .A(n11839), .B(n11840), .Z(n11604) );
  XOR2_X1 U11800 ( .A(n11841), .B(n11842), .Z(n11839) );
  NAND2_X1 U11801 ( .A1(a_23_), .A2(n11838), .ZN(n11605) );
  NAND2_X1 U11802 ( .A1(n11843), .A2(n11844), .ZN(n11838) );
  NAND2_X1 U11803 ( .A1(n11614), .A2(n11845), .ZN(n11844) );
  INV_X1 U11804 ( .A(n11846), .ZN(n11845) );
  NOR2_X1 U11805 ( .A1(n11613), .A2(n11612), .ZN(n11846) );
  NOR2_X1 U11806 ( .A1(n8599), .A2(n8982), .ZN(n11614) );
  NAND2_X1 U11807 ( .A1(n11612), .A2(n11613), .ZN(n11843) );
  NAND2_X1 U11808 ( .A1(n11847), .A2(n11848), .ZN(n11613) );
  NAND2_X1 U11809 ( .A1(n11664), .A2(n11849), .ZN(n11848) );
  NAND2_X1 U11810 ( .A1(n11661), .A2(n11663), .ZN(n11849) );
  NOR2_X1 U11811 ( .A1(n8599), .A2(n8541), .ZN(n11664) );
  INV_X1 U11812 ( .A(n11850), .ZN(n11847) );
  NOR2_X1 U11813 ( .A1(n11663), .A2(n11661), .ZN(n11850) );
  XNOR2_X1 U11814 ( .A(n11851), .B(n11852), .ZN(n11661) );
  XNOR2_X1 U11815 ( .A(n11853), .B(n11854), .ZN(n11852) );
  NAND2_X1 U11816 ( .A1(n11855), .A2(n11856), .ZN(n11663) );
  NAND2_X1 U11817 ( .A1(n11623), .A2(n11857), .ZN(n11856) );
  NAND2_X1 U11818 ( .A1(n11626), .A2(n11625), .ZN(n11857) );
  XNOR2_X1 U11819 ( .A(n11858), .B(n11859), .ZN(n11623) );
  XOR2_X1 U11820 ( .A(n11860), .B(n11861), .Z(n11858) );
  INV_X1 U11821 ( .A(n11862), .ZN(n11855) );
  NOR2_X1 U11822 ( .A1(n11625), .A2(n11626), .ZN(n11862) );
  NOR2_X1 U11823 ( .A1(n8599), .A2(n9893), .ZN(n11626) );
  NAND2_X1 U11824 ( .A1(n11863), .A2(n11864), .ZN(n11625) );
  NAND2_X1 U11825 ( .A1(n11633), .A2(n11865), .ZN(n11864) );
  INV_X1 U11826 ( .A(n11866), .ZN(n11865) );
  NOR2_X1 U11827 ( .A1(n11632), .A2(n11631), .ZN(n11866) );
  NOR2_X1 U11828 ( .A1(n8599), .A2(n8512), .ZN(n11633) );
  NAND2_X1 U11829 ( .A1(n11631), .A2(n11632), .ZN(n11863) );
  NAND2_X1 U11830 ( .A1(n11867), .A2(n11868), .ZN(n11632) );
  NAND2_X1 U11831 ( .A1(n11659), .A2(n11869), .ZN(n11868) );
  INV_X1 U11832 ( .A(n11870), .ZN(n11869) );
  NOR2_X1 U11833 ( .A1(n11660), .A2(n11658), .ZN(n11870) );
  NOR2_X1 U11834 ( .A1(n8599), .A2(n8493), .ZN(n11659) );
  NAND2_X1 U11835 ( .A1(n11658), .A2(n11660), .ZN(n11867) );
  NAND2_X1 U11836 ( .A1(n11871), .A2(n11872), .ZN(n11660) );
  NAND2_X1 U11837 ( .A1(n11654), .A2(n11873), .ZN(n11872) );
  INV_X1 U11838 ( .A(n11874), .ZN(n11873) );
  NOR2_X1 U11839 ( .A1(n11655), .A2(n11656), .ZN(n11874) );
  NOR2_X1 U11840 ( .A1(n8599), .A2(n8473), .ZN(n11654) );
  NAND2_X1 U11841 ( .A1(n11656), .A2(n11655), .ZN(n11871) );
  NAND2_X1 U11842 ( .A1(n11875), .A2(n11876), .ZN(n11655) );
  NAND2_X1 U11843 ( .A1(b_19_), .A2(n11877), .ZN(n11876) );
  NAND2_X1 U11844 ( .A1(n8456), .A2(n11878), .ZN(n11877) );
  NAND2_X1 U11845 ( .A1(a_31_), .A2(n8985), .ZN(n11878) );
  NAND2_X1 U11846 ( .A1(b_20_), .A2(n11879), .ZN(n11875) );
  NAND2_X1 U11847 ( .A1(n8459), .A2(n11880), .ZN(n11879) );
  NAND2_X1 U11848 ( .A1(a_30_), .A2(n8628), .ZN(n11880) );
  NOR3_X1 U11849 ( .A1(n8985), .A2(n8979), .A3(n8599), .ZN(n11656) );
  XOR2_X1 U11850 ( .A(n11881), .B(n11882), .Z(n11658) );
  XOR2_X1 U11851 ( .A(n11883), .B(n11884), .Z(n11881) );
  XOR2_X1 U11852 ( .A(n11885), .B(n11886), .Z(n11631) );
  XOR2_X1 U11853 ( .A(n11887), .B(n11888), .Z(n11885) );
  XNOR2_X1 U11854 ( .A(n11889), .B(n11890), .ZN(n11612) );
  XNOR2_X1 U11855 ( .A(n11891), .B(n11892), .ZN(n11890) );
  NOR2_X1 U11856 ( .A1(n8599), .A2(n8601), .ZN(n8596) );
  XOR2_X1 U11857 ( .A(n11893), .B(n11894), .Z(n11576) );
  XOR2_X1 U11858 ( .A(n11895), .B(n8613), .Z(n11893) );
  XNOR2_X1 U11859 ( .A(n11896), .B(n11897), .ZN(n11549) );
  XNOR2_X1 U11860 ( .A(n11898), .B(n11899), .ZN(n11896) );
  NOR2_X1 U11861 ( .A1(n8680), .A2(n8985), .ZN(n11899) );
  XNOR2_X1 U11862 ( .A(n11900), .B(n11901), .ZN(n11673) );
  XNOR2_X1 U11863 ( .A(n11902), .B(n11903), .ZN(n11900) );
  NOR2_X1 U11864 ( .A1(n8692), .A2(n8985), .ZN(n11903) );
  XOR2_X1 U11865 ( .A(n11904), .B(n11905), .Z(n11520) );
  XNOR2_X1 U11866 ( .A(n11906), .B(n11907), .ZN(n11905) );
  NAND2_X1 U11867 ( .A1(b_20_), .A2(a_11_), .ZN(n11907) );
  XNOR2_X1 U11868 ( .A(n11908), .B(n11909), .ZN(n11686) );
  XNOR2_X1 U11869 ( .A(n11910), .B(n11911), .ZN(n11909) );
  INV_X1 U11870 ( .A(n11689), .ZN(n11741) );
  XNOR2_X1 U11871 ( .A(n11912), .B(n11913), .ZN(n11689) );
  XOR2_X1 U11872 ( .A(n11914), .B(n11915), .Z(n11912) );
  XNOR2_X1 U11873 ( .A(n11916), .B(n11917), .ZN(n11505) );
  XNOR2_X1 U11874 ( .A(n11918), .B(n11919), .ZN(n11916) );
  XNOR2_X1 U11875 ( .A(n11920), .B(n11921), .ZN(n11693) );
  XNOR2_X1 U11876 ( .A(n11922), .B(n11923), .ZN(n11921) );
  NAND2_X1 U11877 ( .A1(b_20_), .A2(a_7_), .ZN(n11923) );
  XNOR2_X1 U11878 ( .A(n11924), .B(n11925), .ZN(n11492) );
  NAND2_X1 U11879 ( .A1(n11926), .A2(n11927), .ZN(n11924) );
  XNOR2_X1 U11880 ( .A(n11928), .B(n11929), .ZN(n11485) );
  XOR2_X1 U11881 ( .A(n11930), .B(n11931), .Z(n11928) );
  XOR2_X1 U11882 ( .A(n11932), .B(n11933), .Z(n11476) );
  XOR2_X1 U11883 ( .A(n11934), .B(n11935), .Z(n11932) );
  XNOR2_X1 U11884 ( .A(n11936), .B(n11937), .ZN(n11697) );
  XNOR2_X1 U11885 ( .A(n11938), .B(n11939), .ZN(n11936) );
  XNOR2_X1 U11886 ( .A(n11940), .B(n11941), .ZN(n11464) );
  XNOR2_X1 U11887 ( .A(n11942), .B(n11943), .ZN(n11941) );
  XOR2_X1 U11888 ( .A(n11944), .B(n11945), .Z(n11702) );
  XOR2_X1 U11889 ( .A(n11946), .B(n11947), .Z(n11944) );
  XNOR2_X1 U11890 ( .A(n11948), .B(n11949), .ZN(n9179) );
  NAND2_X1 U11891 ( .A1(n11950), .A2(n11951), .ZN(n11948) );
  NAND4_X1 U11892 ( .A1(n9174), .A2(n9172), .A3(n9175), .A4(n9173), .ZN(n9077)
         );
  INV_X1 U11893 ( .A(n9166), .ZN(n9173) );
  NOR2_X1 U11894 ( .A1(n11952), .A2(n11953), .ZN(n9166) );
  NAND2_X1 U11895 ( .A1(n11950), .A2(n11954), .ZN(n9175) );
  NAND2_X1 U11896 ( .A1(n11949), .A2(n11951), .ZN(n11954) );
  NAND2_X1 U11897 ( .A1(n11955), .A2(n11956), .ZN(n11951) );
  NAND2_X1 U11898 ( .A1(b_20_), .A2(a_0_), .ZN(n11956) );
  INV_X1 U11899 ( .A(n11957), .ZN(n11955) );
  XOR2_X1 U11900 ( .A(n11958), .B(n11959), .Z(n11949) );
  XNOR2_X1 U11901 ( .A(n11960), .B(n11961), .ZN(n11959) );
  NAND2_X1 U11902 ( .A1(b_19_), .A2(a_1_), .ZN(n11961) );
  NAND2_X1 U11903 ( .A1(a_0_), .A2(n11957), .ZN(n11950) );
  NAND2_X1 U11904 ( .A1(n11962), .A2(n11963), .ZN(n11957) );
  NAND2_X1 U11905 ( .A1(n11947), .A2(n11964), .ZN(n11963) );
  INV_X1 U11906 ( .A(n11965), .ZN(n11964) );
  NOR2_X1 U11907 ( .A1(n11946), .A2(n11945), .ZN(n11965) );
  NOR2_X1 U11908 ( .A1(n8985), .A2(n9731), .ZN(n11947) );
  NAND2_X1 U11909 ( .A1(n11945), .A2(n11946), .ZN(n11962) );
  NAND2_X1 U11910 ( .A1(n11966), .A2(n11967), .ZN(n11946) );
  NAND2_X1 U11911 ( .A1(n11943), .A2(n11968), .ZN(n11967) );
  INV_X1 U11912 ( .A(n11969), .ZN(n11968) );
  NOR2_X1 U11913 ( .A1(n11942), .A2(n11940), .ZN(n11969) );
  NOR2_X1 U11914 ( .A1(n8985), .A2(n8998), .ZN(n11943) );
  NAND2_X1 U11915 ( .A1(n11940), .A2(n11942), .ZN(n11966) );
  NAND2_X1 U11916 ( .A1(n11970), .A2(n11971), .ZN(n11942) );
  NAND2_X1 U11917 ( .A1(n11939), .A2(n11972), .ZN(n11971) );
  NAND2_X1 U11918 ( .A1(n11938), .A2(n11937), .ZN(n11972) );
  NOR2_X1 U11919 ( .A1(n8985), .A2(n8877), .ZN(n11939) );
  INV_X1 U11920 ( .A(n11973), .ZN(n11970) );
  NOR2_X1 U11921 ( .A1(n11937), .A2(n11938), .ZN(n11973) );
  NOR2_X1 U11922 ( .A1(n11974), .A2(n11975), .ZN(n11938) );
  INV_X1 U11923 ( .A(n11976), .ZN(n11975) );
  NAND2_X1 U11924 ( .A1(n11935), .A2(n11977), .ZN(n11976) );
  NAND2_X1 U11925 ( .A1(n11933), .A2(n11934), .ZN(n11977) );
  NOR2_X1 U11926 ( .A1(n8985), .A2(n8996), .ZN(n11935) );
  NOR2_X1 U11927 ( .A1(n11934), .A2(n11933), .ZN(n11974) );
  XOR2_X1 U11928 ( .A(n11978), .B(n11979), .Z(n11933) );
  XOR2_X1 U11929 ( .A(n11980), .B(n11981), .Z(n11979) );
  NAND2_X1 U11930 ( .A1(b_19_), .A2(a_5_), .ZN(n11981) );
  NAND2_X1 U11931 ( .A1(n11982), .A2(n11983), .ZN(n11934) );
  NAND2_X1 U11932 ( .A1(n11929), .A2(n11984), .ZN(n11983) );
  NAND2_X1 U11933 ( .A1(n11931), .A2(n11930), .ZN(n11984) );
  XNOR2_X1 U11934 ( .A(n11985), .B(n11986), .ZN(n11929) );
  XOR2_X1 U11935 ( .A(n11987), .B(n11988), .Z(n11985) );
  NOR2_X1 U11936 ( .A1(n8994), .A2(n8628), .ZN(n11988) );
  INV_X1 U11937 ( .A(n11989), .ZN(n11982) );
  NOR2_X1 U11938 ( .A1(n11930), .A2(n11931), .ZN(n11989) );
  NOR2_X1 U11939 ( .A1(n8985), .A2(n8848), .ZN(n11931) );
  NAND2_X1 U11940 ( .A1(n11926), .A2(n11990), .ZN(n11930) );
  NAND2_X1 U11941 ( .A1(n11925), .A2(n11927), .ZN(n11990) );
  NAND2_X1 U11942 ( .A1(n11991), .A2(n11992), .ZN(n11927) );
  NAND2_X1 U11943 ( .A1(b_20_), .A2(a_6_), .ZN(n11992) );
  INV_X1 U11944 ( .A(n11993), .ZN(n11991) );
  XOR2_X1 U11945 ( .A(n11994), .B(n11995), .Z(n11925) );
  XNOR2_X1 U11946 ( .A(n11996), .B(n11997), .ZN(n11995) );
  NAND2_X1 U11947 ( .A1(b_19_), .A2(a_7_), .ZN(n11997) );
  NAND2_X1 U11948 ( .A1(a_6_), .A2(n11993), .ZN(n11926) );
  NAND2_X1 U11949 ( .A1(n11998), .A2(n11999), .ZN(n11993) );
  NAND3_X1 U11950 ( .A1(a_7_), .A2(n12000), .A3(b_20_), .ZN(n11999) );
  NAND2_X1 U11951 ( .A1(n11922), .A2(n12001), .ZN(n12000) );
  INV_X1 U11952 ( .A(n11920), .ZN(n12001) );
  NAND2_X1 U11953 ( .A1(n11920), .A2(n12002), .ZN(n11998) );
  INV_X1 U11954 ( .A(n11922), .ZN(n12002) );
  NOR2_X1 U11955 ( .A1(n12003), .A2(n12004), .ZN(n11922) );
  INV_X1 U11956 ( .A(n12005), .ZN(n12004) );
  NAND2_X1 U11957 ( .A1(n11919), .A2(n12006), .ZN(n12005) );
  NAND2_X1 U11958 ( .A1(n11918), .A2(n11917), .ZN(n12006) );
  NOR2_X1 U11959 ( .A1(n8985), .A2(n10513), .ZN(n11919) );
  NOR2_X1 U11960 ( .A1(n11917), .A2(n11918), .ZN(n12003) );
  NOR2_X1 U11961 ( .A1(n12007), .A2(n12008), .ZN(n11918) );
  INV_X1 U11962 ( .A(n12009), .ZN(n12008) );
  NAND2_X1 U11963 ( .A1(n11915), .A2(n12010), .ZN(n12009) );
  NAND2_X1 U11964 ( .A1(n11913), .A2(n11914), .ZN(n12010) );
  NOR2_X1 U11965 ( .A1(n8985), .A2(n8779), .ZN(n11915) );
  NOR2_X1 U11966 ( .A1(n11914), .A2(n11913), .ZN(n12007) );
  XOR2_X1 U11967 ( .A(n12011), .B(n12012), .Z(n11913) );
  XOR2_X1 U11968 ( .A(n12013), .B(n12014), .Z(n12012) );
  NAND2_X1 U11969 ( .A1(b_19_), .A2(a_10_), .ZN(n12014) );
  NAND2_X1 U11970 ( .A1(n12015), .A2(n12016), .ZN(n11914) );
  NAND2_X1 U11971 ( .A1(n11908), .A2(n12017), .ZN(n12016) );
  NAND2_X1 U11972 ( .A1(n11911), .A2(n11910), .ZN(n12017) );
  XOR2_X1 U11973 ( .A(n12018), .B(n12019), .Z(n11908) );
  XNOR2_X1 U11974 ( .A(n12020), .B(n12021), .ZN(n12019) );
  INV_X1 U11975 ( .A(n12022), .ZN(n12015) );
  NOR2_X1 U11976 ( .A1(n11910), .A2(n11911), .ZN(n12022) );
  NOR2_X1 U11977 ( .A1(n8985), .A2(n8769), .ZN(n11911) );
  NAND2_X1 U11978 ( .A1(n12023), .A2(n12024), .ZN(n11910) );
  NAND3_X1 U11979 ( .A1(a_11_), .A2(n12025), .A3(b_20_), .ZN(n12024) );
  NAND2_X1 U11980 ( .A1(n11904), .A2(n12026), .ZN(n12025) );
  INV_X1 U11981 ( .A(n11906), .ZN(n12026) );
  NAND2_X1 U11982 ( .A1(n11906), .A2(n12027), .ZN(n12023) );
  INV_X1 U11983 ( .A(n11904), .ZN(n12027) );
  XNOR2_X1 U11984 ( .A(n12028), .B(n12029), .ZN(n11904) );
  XNOR2_X1 U11985 ( .A(n12030), .B(n12031), .ZN(n12029) );
  NOR2_X1 U11986 ( .A1(n12032), .A2(n12033), .ZN(n11906) );
  INV_X1 U11987 ( .A(n12034), .ZN(n12033) );
  NAND2_X1 U11988 ( .A1(n11756), .A2(n12035), .ZN(n12034) );
  NAND2_X1 U11989 ( .A1(n11758), .A2(n11757), .ZN(n12035) );
  XNOR2_X1 U11990 ( .A(n12036), .B(n12037), .ZN(n11756) );
  XNOR2_X1 U11991 ( .A(n12038), .B(n12039), .ZN(n12037) );
  NAND2_X1 U11992 ( .A1(b_19_), .A2(a_13_), .ZN(n12039) );
  NOR2_X1 U11993 ( .A1(n11757), .A2(n11758), .ZN(n12032) );
  NOR2_X1 U11994 ( .A1(n8985), .A2(n8739), .ZN(n11758) );
  NAND2_X1 U11995 ( .A1(n11764), .A2(n12040), .ZN(n11757) );
  NAND2_X1 U11996 ( .A1(n11763), .A2(n11765), .ZN(n12040) );
  NAND2_X1 U11997 ( .A1(n12041), .A2(n12042), .ZN(n11765) );
  NAND2_X1 U11998 ( .A1(b_20_), .A2(a_13_), .ZN(n12041) );
  XNOR2_X1 U11999 ( .A(n12043), .B(n12044), .ZN(n11763) );
  XNOR2_X1 U12000 ( .A(n12045), .B(n12046), .ZN(n12043) );
  NOR2_X1 U12001 ( .A1(n8991), .A2(n8628), .ZN(n12046) );
  INV_X1 U12002 ( .A(n12047), .ZN(n11764) );
  NOR2_X1 U12003 ( .A1(n12042), .A2(n8721), .ZN(n12047) );
  NAND2_X1 U12004 ( .A1(n12048), .A2(n12049), .ZN(n12042) );
  NAND2_X1 U12005 ( .A1(n11770), .A2(n12050), .ZN(n12049) );
  INV_X1 U12006 ( .A(n12051), .ZN(n12050) );
  NOR2_X1 U12007 ( .A1(n11773), .A2(n11772), .ZN(n12051) );
  XNOR2_X1 U12008 ( .A(n12052), .B(n12053), .ZN(n11770) );
  XOR2_X1 U12009 ( .A(n12054), .B(n12055), .Z(n12052) );
  NOR2_X1 U12010 ( .A1(n8692), .A2(n8628), .ZN(n12055) );
  NAND2_X1 U12011 ( .A1(n11772), .A2(n11773), .ZN(n12048) );
  NAND2_X1 U12012 ( .A1(b_20_), .A2(a_14_), .ZN(n11773) );
  NOR2_X1 U12013 ( .A1(n12056), .A2(n12057), .ZN(n11772) );
  INV_X1 U12014 ( .A(n12058), .ZN(n12057) );
  NAND3_X1 U12015 ( .A1(a_15_), .A2(n12059), .A3(b_20_), .ZN(n12058) );
  NAND2_X1 U12016 ( .A1(n11902), .A2(n11901), .ZN(n12059) );
  NOR2_X1 U12017 ( .A1(n11901), .A2(n11902), .ZN(n12056) );
  NOR2_X1 U12018 ( .A1(n12060), .A2(n12061), .ZN(n11902) );
  INV_X1 U12019 ( .A(n12062), .ZN(n12061) );
  NAND3_X1 U12020 ( .A1(a_16_), .A2(n12063), .A3(b_20_), .ZN(n12062) );
  NAND2_X1 U12021 ( .A1(n11898), .A2(n11897), .ZN(n12063) );
  NOR2_X1 U12022 ( .A1(n11897), .A2(n11898), .ZN(n12060) );
  NOR2_X1 U12023 ( .A1(n12064), .A2(n12065), .ZN(n11898) );
  INV_X1 U12024 ( .A(n12066), .ZN(n12065) );
  NAND3_X1 U12025 ( .A1(a_17_), .A2(n12067), .A3(b_20_), .ZN(n12066) );
  NAND2_X1 U12026 ( .A1(n11786), .A2(n11788), .ZN(n12067) );
  NOR2_X1 U12027 ( .A1(n11788), .A2(n11786), .ZN(n12064) );
  XNOR2_X1 U12028 ( .A(n12068), .B(n12069), .ZN(n11786) );
  XOR2_X1 U12029 ( .A(n12070), .B(n12071), .Z(n12068) );
  NAND2_X1 U12030 ( .A1(n12072), .A2(n12073), .ZN(n11788) );
  NAND2_X1 U12031 ( .A1(n11795), .A2(n12074), .ZN(n12073) );
  NAND2_X1 U12032 ( .A1(n11798), .A2(n11797), .ZN(n12074) );
  XOR2_X1 U12033 ( .A(n12075), .B(n12076), .Z(n11795) );
  XNOR2_X1 U12034 ( .A(n12077), .B(n8953), .ZN(n12076) );
  INV_X1 U12035 ( .A(n12078), .ZN(n12072) );
  NOR2_X1 U12036 ( .A1(n11797), .A2(n11798), .ZN(n12078) );
  NOR2_X1 U12037 ( .A1(n8985), .A2(n8988), .ZN(n11798) );
  NAND2_X1 U12038 ( .A1(n12079), .A2(n12080), .ZN(n11797) );
  NAND3_X1 U12039 ( .A1(a_19_), .A2(n12081), .A3(b_20_), .ZN(n12080) );
  INV_X1 U12040 ( .A(n12082), .ZN(n12081) );
  NOR2_X1 U12041 ( .A1(n11804), .A2(n11802), .ZN(n12082) );
  NAND2_X1 U12042 ( .A1(n11802), .A2(n11804), .ZN(n12079) );
  NAND2_X1 U12043 ( .A1(n12083), .A2(n12084), .ZN(n11804) );
  NAND2_X1 U12044 ( .A1(n11894), .A2(n12085), .ZN(n12084) );
  NAND2_X1 U12045 ( .A1(n11895), .A2(n8613), .ZN(n12085) );
  XNOR2_X1 U12046 ( .A(n12086), .B(n12087), .ZN(n11894) );
  XOR2_X1 U12047 ( .A(n12088), .B(n12089), .Z(n12087) );
  NAND2_X1 U12048 ( .A1(b_19_), .A2(a_21_), .ZN(n12089) );
  INV_X1 U12049 ( .A(n12090), .ZN(n12083) );
  NOR2_X1 U12050 ( .A1(n8613), .A2(n11895), .ZN(n12090) );
  NOR2_X1 U12051 ( .A1(n12091), .A2(n12092), .ZN(n11895) );
  NOR3_X1 U12052 ( .A1(n8601), .A2(n12093), .A3(n8985), .ZN(n12092) );
  NOR2_X1 U12053 ( .A1(n11817), .A2(n11815), .ZN(n12093) );
  INV_X1 U12054 ( .A(n12094), .ZN(n12091) );
  NAND2_X1 U12055 ( .A1(n11815), .A2(n11817), .ZN(n12094) );
  NAND2_X1 U12056 ( .A1(n11825), .A2(n12095), .ZN(n11817) );
  NAND2_X1 U12057 ( .A1(n11824), .A2(n11826), .ZN(n12095) );
  NAND2_X1 U12058 ( .A1(n12096), .A2(n12097), .ZN(n11826) );
  NAND2_X1 U12059 ( .A1(b_20_), .A2(a_22_), .ZN(n12097) );
  INV_X1 U12060 ( .A(n12098), .ZN(n12096) );
  XNOR2_X1 U12061 ( .A(n12099), .B(n12100), .ZN(n11824) );
  NAND2_X1 U12062 ( .A1(n12101), .A2(n12102), .ZN(n12099) );
  NAND2_X1 U12063 ( .A1(a_22_), .A2(n12098), .ZN(n11825) );
  NAND2_X1 U12064 ( .A1(n11833), .A2(n12103), .ZN(n12098) );
  NAND2_X1 U12065 ( .A1(n11832), .A2(n11834), .ZN(n12103) );
  NAND2_X1 U12066 ( .A1(n12104), .A2(n12105), .ZN(n11834) );
  NAND2_X1 U12067 ( .A1(b_20_), .A2(a_23_), .ZN(n12105) );
  INV_X1 U12068 ( .A(n12106), .ZN(n12104) );
  XOR2_X1 U12069 ( .A(n12107), .B(n12108), .Z(n11832) );
  XOR2_X1 U12070 ( .A(n12109), .B(n12110), .Z(n12107) );
  NAND2_X1 U12071 ( .A1(a_23_), .A2(n12106), .ZN(n11833) );
  NAND2_X1 U12072 ( .A1(n12111), .A2(n12112), .ZN(n12106) );
  NAND2_X1 U12073 ( .A1(n11842), .A2(n12113), .ZN(n12112) );
  INV_X1 U12074 ( .A(n12114), .ZN(n12113) );
  NOR2_X1 U12075 ( .A1(n11841), .A2(n11840), .ZN(n12114) );
  NOR2_X1 U12076 ( .A1(n8985), .A2(n8982), .ZN(n11842) );
  NAND2_X1 U12077 ( .A1(n11840), .A2(n11841), .ZN(n12111) );
  NAND2_X1 U12078 ( .A1(n12115), .A2(n12116), .ZN(n11841) );
  NAND2_X1 U12079 ( .A1(n11892), .A2(n12117), .ZN(n12116) );
  NAND2_X1 U12080 ( .A1(n11889), .A2(n11891), .ZN(n12117) );
  NOR2_X1 U12081 ( .A1(n8985), .A2(n8541), .ZN(n11892) );
  INV_X1 U12082 ( .A(n12118), .ZN(n12115) );
  NOR2_X1 U12083 ( .A1(n11891), .A2(n11889), .ZN(n12118) );
  XNOR2_X1 U12084 ( .A(n12119), .B(n12120), .ZN(n11889) );
  XNOR2_X1 U12085 ( .A(n12121), .B(n12122), .ZN(n12120) );
  NAND2_X1 U12086 ( .A1(n12123), .A2(n12124), .ZN(n11891) );
  NAND2_X1 U12087 ( .A1(n11851), .A2(n12125), .ZN(n12124) );
  NAND2_X1 U12088 ( .A1(n11854), .A2(n11853), .ZN(n12125) );
  XNOR2_X1 U12089 ( .A(n12126), .B(n12127), .ZN(n11851) );
  XOR2_X1 U12090 ( .A(n12128), .B(n12129), .Z(n12126) );
  INV_X1 U12091 ( .A(n12130), .ZN(n12123) );
  NOR2_X1 U12092 ( .A1(n11853), .A2(n11854), .ZN(n12130) );
  NOR2_X1 U12093 ( .A1(n8985), .A2(n9893), .ZN(n11854) );
  NAND2_X1 U12094 ( .A1(n12131), .A2(n12132), .ZN(n11853) );
  NAND2_X1 U12095 ( .A1(n11861), .A2(n12133), .ZN(n12132) );
  INV_X1 U12096 ( .A(n12134), .ZN(n12133) );
  NOR2_X1 U12097 ( .A1(n11860), .A2(n11859), .ZN(n12134) );
  NOR2_X1 U12098 ( .A1(n8985), .A2(n8512), .ZN(n11861) );
  NAND2_X1 U12099 ( .A1(n11859), .A2(n11860), .ZN(n12131) );
  NAND2_X1 U12100 ( .A1(n12135), .A2(n12136), .ZN(n11860) );
  NAND2_X1 U12101 ( .A1(n11887), .A2(n12137), .ZN(n12136) );
  INV_X1 U12102 ( .A(n12138), .ZN(n12137) );
  NOR2_X1 U12103 ( .A1(n11888), .A2(n11886), .ZN(n12138) );
  NOR2_X1 U12104 ( .A1(n8985), .A2(n8493), .ZN(n11887) );
  NAND2_X1 U12105 ( .A1(n11886), .A2(n11888), .ZN(n12135) );
  NAND2_X1 U12106 ( .A1(n12139), .A2(n12140), .ZN(n11888) );
  NAND2_X1 U12107 ( .A1(n11882), .A2(n12141), .ZN(n12140) );
  INV_X1 U12108 ( .A(n12142), .ZN(n12141) );
  NOR2_X1 U12109 ( .A1(n11883), .A2(n11884), .ZN(n12142) );
  NOR2_X1 U12110 ( .A1(n8985), .A2(n8473), .ZN(n11882) );
  NAND2_X1 U12111 ( .A1(n11884), .A2(n11883), .ZN(n12139) );
  NAND2_X1 U12112 ( .A1(n12143), .A2(n12144), .ZN(n11883) );
  NAND2_X1 U12113 ( .A1(b_18_), .A2(n12145), .ZN(n12144) );
  NAND2_X1 U12114 ( .A1(n8456), .A2(n12146), .ZN(n12145) );
  NAND2_X1 U12115 ( .A1(a_31_), .A2(n8628), .ZN(n12146) );
  NAND2_X1 U12116 ( .A1(b_19_), .A2(n12147), .ZN(n12143) );
  NAND2_X1 U12117 ( .A1(n8459), .A2(n12148), .ZN(n12147) );
  NAND2_X1 U12118 ( .A1(a_30_), .A2(n8987), .ZN(n12148) );
  NOR3_X1 U12119 ( .A1(n8628), .A2(n8979), .A3(n8985), .ZN(n11884) );
  INV_X1 U12120 ( .A(b_20_), .ZN(n8985) );
  XOR2_X1 U12121 ( .A(n12149), .B(n12150), .Z(n11886) );
  XOR2_X1 U12122 ( .A(n12151), .B(n12152), .Z(n12149) );
  XOR2_X1 U12123 ( .A(n12153), .B(n12154), .Z(n11859) );
  XOR2_X1 U12124 ( .A(n12155), .B(n12156), .Z(n12153) );
  XNOR2_X1 U12125 ( .A(n12157), .B(n12158), .ZN(n11840) );
  XNOR2_X1 U12126 ( .A(n12159), .B(n12160), .ZN(n12158) );
  XNOR2_X1 U12127 ( .A(n12161), .B(n12162), .ZN(n11815) );
  NAND2_X1 U12128 ( .A1(n12163), .A2(n12164), .ZN(n12161) );
  NAND2_X1 U12129 ( .A1(b_20_), .A2(a_20_), .ZN(n8613) );
  XNOR2_X1 U12130 ( .A(n12165), .B(n12166), .ZN(n11802) );
  XOR2_X1 U12131 ( .A(n12167), .B(n12168), .Z(n12165) );
  XOR2_X1 U12132 ( .A(n12169), .B(n12170), .Z(n11897) );
  NAND2_X1 U12133 ( .A1(n12171), .A2(n12172), .ZN(n12169) );
  XOR2_X1 U12134 ( .A(n12173), .B(n12174), .Z(n11901) );
  NAND2_X1 U12135 ( .A1(n12175), .A2(n12176), .ZN(n12173) );
  XOR2_X1 U12136 ( .A(n12177), .B(n12178), .Z(n11917) );
  XOR2_X1 U12137 ( .A(n12179), .B(n12180), .Z(n12178) );
  NAND2_X1 U12138 ( .A1(b_19_), .A2(a_9_), .ZN(n12180) );
  XOR2_X1 U12139 ( .A(n12181), .B(n12182), .Z(n11920) );
  XNOR2_X1 U12140 ( .A(n12183), .B(n12184), .ZN(n12182) );
  NAND2_X1 U12141 ( .A1(b_19_), .A2(a_8_), .ZN(n12184) );
  XNOR2_X1 U12142 ( .A(n12185), .B(n12186), .ZN(n11937) );
  XOR2_X1 U12143 ( .A(n12187), .B(n12188), .Z(n12185) );
  NOR2_X1 U12144 ( .A1(n8996), .A2(n8628), .ZN(n12188) );
  XNOR2_X1 U12145 ( .A(n12189), .B(n12190), .ZN(n11940) );
  XOR2_X1 U12146 ( .A(n12191), .B(n12192), .Z(n12190) );
  NAND2_X1 U12147 ( .A1(b_19_), .A2(a_3_), .ZN(n12192) );
  XOR2_X1 U12148 ( .A(n12193), .B(n12194), .Z(n11945) );
  XOR2_X1 U12149 ( .A(n12195), .B(n12196), .Z(n12193) );
  NOR2_X1 U12150 ( .A1(n8998), .A2(n8628), .ZN(n12196) );
  NAND2_X1 U12151 ( .A1(n11953), .A2(n11952), .ZN(n9172) );
  XOR2_X1 U12152 ( .A(n12197), .B(n12198), .Z(n11952) );
  NAND2_X1 U12153 ( .A1(n12199), .A2(n12200), .ZN(n12197) );
  NOR2_X1 U12154 ( .A1(n12201), .A2(n12202), .ZN(n11953) );
  INV_X1 U12155 ( .A(n12203), .ZN(n12202) );
  NAND3_X1 U12156 ( .A1(a_0_), .A2(n12204), .A3(b_19_), .ZN(n12203) );
  NAND2_X1 U12157 ( .A1(n12205), .A2(n12206), .ZN(n12204) );
  NOR2_X1 U12158 ( .A1(n12206), .A2(n12205), .ZN(n12201) );
  XOR2_X1 U12159 ( .A(n12206), .B(n12207), .Z(n9174) );
  XNOR2_X1 U12160 ( .A(n12205), .B(n12208), .ZN(n12207) );
  NAND2_X1 U12161 ( .A1(b_19_), .A2(a_0_), .ZN(n12208) );
  NOR2_X1 U12162 ( .A1(n12209), .A2(n12210), .ZN(n12205) );
  NOR3_X1 U12163 ( .A1(n9731), .A2(n12211), .A3(n8628), .ZN(n12210) );
  INV_X1 U12164 ( .A(n12212), .ZN(n12211) );
  NAND2_X1 U12165 ( .A1(n11960), .A2(n11958), .ZN(n12212) );
  NOR2_X1 U12166 ( .A1(n11958), .A2(n11960), .ZN(n12209) );
  NOR2_X1 U12167 ( .A1(n12213), .A2(n12214), .ZN(n11960) );
  NOR3_X1 U12168 ( .A1(n8998), .A2(n12215), .A3(n8628), .ZN(n12214) );
  NOR2_X1 U12169 ( .A1(n12195), .A2(n12194), .ZN(n12215) );
  INV_X1 U12170 ( .A(n12216), .ZN(n12213) );
  NAND2_X1 U12171 ( .A1(n12194), .A2(n12195), .ZN(n12216) );
  NAND2_X1 U12172 ( .A1(n12217), .A2(n12218), .ZN(n12195) );
  NAND3_X1 U12173 ( .A1(a_3_), .A2(n12219), .A3(b_19_), .ZN(n12218) );
  INV_X1 U12174 ( .A(n12220), .ZN(n12219) );
  NOR2_X1 U12175 ( .A1(n12191), .A2(n12189), .ZN(n12220) );
  NAND2_X1 U12176 ( .A1(n12189), .A2(n12191), .ZN(n12217) );
  NAND2_X1 U12177 ( .A1(n12221), .A2(n12222), .ZN(n12191) );
  NAND3_X1 U12178 ( .A1(a_4_), .A2(n12223), .A3(b_19_), .ZN(n12222) );
  INV_X1 U12179 ( .A(n12224), .ZN(n12223) );
  NOR2_X1 U12180 ( .A1(n12187), .A2(n12186), .ZN(n12224) );
  NAND2_X1 U12181 ( .A1(n12186), .A2(n12187), .ZN(n12221) );
  NAND2_X1 U12182 ( .A1(n12225), .A2(n12226), .ZN(n12187) );
  INV_X1 U12183 ( .A(n12227), .ZN(n12226) );
  NOR3_X1 U12184 ( .A1(n8848), .A2(n12228), .A3(n8628), .ZN(n12227) );
  NOR2_X1 U12185 ( .A1(n11980), .A2(n11978), .ZN(n12228) );
  NAND2_X1 U12186 ( .A1(n11978), .A2(n11980), .ZN(n12225) );
  NAND2_X1 U12187 ( .A1(n12229), .A2(n12230), .ZN(n11980) );
  NAND3_X1 U12188 ( .A1(a_6_), .A2(n12231), .A3(b_19_), .ZN(n12230) );
  INV_X1 U12189 ( .A(n12232), .ZN(n12231) );
  NOR2_X1 U12190 ( .A1(n11987), .A2(n11986), .ZN(n12232) );
  NAND2_X1 U12191 ( .A1(n11986), .A2(n11987), .ZN(n12229) );
  NAND2_X1 U12192 ( .A1(n12233), .A2(n12234), .ZN(n11987) );
  NAND3_X1 U12193 ( .A1(a_7_), .A2(n12235), .A3(b_19_), .ZN(n12234) );
  NAND2_X1 U12194 ( .A1(n11996), .A2(n11994), .ZN(n12235) );
  INV_X1 U12195 ( .A(n12236), .ZN(n12233) );
  NOR2_X1 U12196 ( .A1(n11994), .A2(n11996), .ZN(n12236) );
  NOR2_X1 U12197 ( .A1(n12237), .A2(n12238), .ZN(n11996) );
  INV_X1 U12198 ( .A(n12239), .ZN(n12238) );
  NAND3_X1 U12199 ( .A1(a_8_), .A2(n12240), .A3(b_19_), .ZN(n12239) );
  NAND2_X1 U12200 ( .A1(n12183), .A2(n12181), .ZN(n12240) );
  NOR2_X1 U12201 ( .A1(n12181), .A2(n12183), .ZN(n12237) );
  NOR2_X1 U12202 ( .A1(n12241), .A2(n12242), .ZN(n12183) );
  NOR3_X1 U12203 ( .A1(n8779), .A2(n12243), .A3(n8628), .ZN(n12242) );
  NOR2_X1 U12204 ( .A1(n12179), .A2(n12177), .ZN(n12243) );
  INV_X1 U12205 ( .A(n12244), .ZN(n12241) );
  NAND2_X1 U12206 ( .A1(n12177), .A2(n12179), .ZN(n12244) );
  NAND2_X1 U12207 ( .A1(n12245), .A2(n12246), .ZN(n12179) );
  NAND3_X1 U12208 ( .A1(a_10_), .A2(n12247), .A3(b_19_), .ZN(n12246) );
  INV_X1 U12209 ( .A(n12248), .ZN(n12247) );
  NOR2_X1 U12210 ( .A1(n12013), .A2(n12011), .ZN(n12248) );
  NAND2_X1 U12211 ( .A1(n12011), .A2(n12013), .ZN(n12245) );
  NAND2_X1 U12212 ( .A1(n12249), .A2(n12250), .ZN(n12013) );
  NAND2_X1 U12213 ( .A1(n12021), .A2(n12251), .ZN(n12250) );
  NAND2_X1 U12214 ( .A1(n12018), .A2(n12020), .ZN(n12251) );
  NOR2_X1 U12215 ( .A1(n8628), .A2(n8749), .ZN(n12021) );
  INV_X1 U12216 ( .A(n12252), .ZN(n12249) );
  NOR2_X1 U12217 ( .A1(n12020), .A2(n12018), .ZN(n12252) );
  XOR2_X1 U12218 ( .A(n12253), .B(n12254), .Z(n12018) );
  XNOR2_X1 U12219 ( .A(n12255), .B(n12256), .ZN(n12253) );
  NOR2_X1 U12220 ( .A1(n8739), .A2(n8987), .ZN(n12256) );
  NAND2_X1 U12221 ( .A1(n12257), .A2(n12258), .ZN(n12020) );
  NAND2_X1 U12222 ( .A1(n12028), .A2(n12259), .ZN(n12258) );
  NAND2_X1 U12223 ( .A1(n12031), .A2(n12030), .ZN(n12259) );
  XOR2_X1 U12224 ( .A(n12260), .B(n12261), .Z(n12028) );
  XNOR2_X1 U12225 ( .A(n12262), .B(n12263), .ZN(n12260) );
  NOR2_X1 U12226 ( .A1(n8721), .A2(n8987), .ZN(n12263) );
  INV_X1 U12227 ( .A(n12264), .ZN(n12257) );
  NOR2_X1 U12228 ( .A1(n12030), .A2(n12031), .ZN(n12264) );
  NOR2_X1 U12229 ( .A1(n8628), .A2(n8739), .ZN(n12031) );
  NAND2_X1 U12230 ( .A1(n12265), .A2(n12266), .ZN(n12030) );
  NAND3_X1 U12231 ( .A1(a_13_), .A2(n12267), .A3(b_19_), .ZN(n12266) );
  NAND2_X1 U12232 ( .A1(n12038), .A2(n12036), .ZN(n12267) );
  INV_X1 U12233 ( .A(n12268), .ZN(n12265) );
  NOR2_X1 U12234 ( .A1(n12036), .A2(n12038), .ZN(n12268) );
  NOR2_X1 U12235 ( .A1(n12269), .A2(n12270), .ZN(n12038) );
  INV_X1 U12236 ( .A(n12271), .ZN(n12270) );
  NAND3_X1 U12237 ( .A1(a_14_), .A2(n12272), .A3(b_19_), .ZN(n12271) );
  NAND2_X1 U12238 ( .A1(n12045), .A2(n12044), .ZN(n12272) );
  NOR2_X1 U12239 ( .A1(n12044), .A2(n12045), .ZN(n12269) );
  NOR2_X1 U12240 ( .A1(n12273), .A2(n12274), .ZN(n12045) );
  NOR3_X1 U12241 ( .A1(n8692), .A2(n12275), .A3(n8628), .ZN(n12274) );
  NOR2_X1 U12242 ( .A1(n12054), .A2(n12053), .ZN(n12275) );
  INV_X1 U12243 ( .A(n12276), .ZN(n12273) );
  NAND2_X1 U12244 ( .A1(n12053), .A2(n12054), .ZN(n12276) );
  NAND2_X1 U12245 ( .A1(n12175), .A2(n12277), .ZN(n12054) );
  NAND2_X1 U12246 ( .A1(n12174), .A2(n12176), .ZN(n12277) );
  NAND2_X1 U12247 ( .A1(n12278), .A2(n12279), .ZN(n12176) );
  NAND2_X1 U12248 ( .A1(b_19_), .A2(a_16_), .ZN(n12279) );
  INV_X1 U12249 ( .A(n12280), .ZN(n12278) );
  XNOR2_X1 U12250 ( .A(n12281), .B(n12282), .ZN(n12174) );
  NAND2_X1 U12251 ( .A1(n12283), .A2(n12284), .ZN(n12281) );
  NAND2_X1 U12252 ( .A1(a_16_), .A2(n12280), .ZN(n12175) );
  NAND2_X1 U12253 ( .A1(n12171), .A2(n12285), .ZN(n12280) );
  NAND2_X1 U12254 ( .A1(n12170), .A2(n12172), .ZN(n12285) );
  NAND2_X1 U12255 ( .A1(n12286), .A2(n12287), .ZN(n12172) );
  NAND2_X1 U12256 ( .A1(b_19_), .A2(a_17_), .ZN(n12287) );
  XOR2_X1 U12257 ( .A(n12288), .B(n12289), .Z(n12170) );
  XOR2_X1 U12258 ( .A(n12290), .B(n8642), .Z(n12288) );
  NAND2_X1 U12259 ( .A1(a_17_), .A2(n12291), .ZN(n12171) );
  INV_X1 U12260 ( .A(n12286), .ZN(n12291) );
  NOR2_X1 U12261 ( .A1(n12292), .A2(n12293), .ZN(n12286) );
  INV_X1 U12262 ( .A(n12294), .ZN(n12293) );
  NAND2_X1 U12263 ( .A1(n12071), .A2(n12295), .ZN(n12294) );
  NAND2_X1 U12264 ( .A1(n12069), .A2(n12070), .ZN(n12295) );
  NOR2_X1 U12265 ( .A1(n8628), .A2(n8988), .ZN(n12071) );
  NOR2_X1 U12266 ( .A1(n12070), .A2(n12069), .ZN(n12292) );
  XNOR2_X1 U12267 ( .A(n12296), .B(n12297), .ZN(n12069) );
  XNOR2_X1 U12268 ( .A(n12298), .B(n12299), .ZN(n12297) );
  NAND2_X1 U12269 ( .A1(b_18_), .A2(a_19_), .ZN(n12299) );
  NAND2_X1 U12270 ( .A1(n12300), .A2(n12301), .ZN(n12070) );
  NAND2_X1 U12271 ( .A1(n12075), .A2(n12302), .ZN(n12301) );
  NAND2_X1 U12272 ( .A1(n12077), .A2(n8625), .ZN(n12302) );
  XNOR2_X1 U12273 ( .A(n12303), .B(n12304), .ZN(n12075) );
  XOR2_X1 U12274 ( .A(n12305), .B(n12306), .Z(n12303) );
  NOR2_X1 U12275 ( .A1(n8986), .A2(n8987), .ZN(n12306) );
  NAND2_X1 U12276 ( .A1(n8953), .A2(n12307), .ZN(n12300) );
  INV_X1 U12277 ( .A(n12077), .ZN(n12307) );
  NOR2_X1 U12278 ( .A1(n12308), .A2(n12309), .ZN(n12077) );
  INV_X1 U12279 ( .A(n12310), .ZN(n12309) );
  NAND2_X1 U12280 ( .A1(n12166), .A2(n12311), .ZN(n12310) );
  NAND2_X1 U12281 ( .A1(n12168), .A2(n12167), .ZN(n12311) );
  XNOR2_X1 U12282 ( .A(n12312), .B(n12313), .ZN(n12166) );
  XOR2_X1 U12283 ( .A(n12314), .B(n12315), .Z(n12312) );
  NOR2_X1 U12284 ( .A1(n8601), .A2(n8987), .ZN(n12315) );
  NOR2_X1 U12285 ( .A1(n12167), .A2(n12168), .ZN(n12308) );
  NOR2_X1 U12286 ( .A1(n8628), .A2(n8986), .ZN(n12168) );
  NAND2_X1 U12287 ( .A1(n12316), .A2(n12317), .ZN(n12167) );
  NAND3_X1 U12288 ( .A1(a_21_), .A2(n12318), .A3(b_19_), .ZN(n12317) );
  INV_X1 U12289 ( .A(n12319), .ZN(n12318) );
  NOR2_X1 U12290 ( .A1(n12088), .A2(n12086), .ZN(n12319) );
  NAND2_X1 U12291 ( .A1(n12086), .A2(n12088), .ZN(n12316) );
  NAND2_X1 U12292 ( .A1(n12163), .A2(n12320), .ZN(n12088) );
  NAND2_X1 U12293 ( .A1(n12162), .A2(n12164), .ZN(n12320) );
  NAND2_X1 U12294 ( .A1(n12321), .A2(n12322), .ZN(n12164) );
  NAND2_X1 U12295 ( .A1(b_19_), .A2(a_22_), .ZN(n12322) );
  INV_X1 U12296 ( .A(n12323), .ZN(n12321) );
  XNOR2_X1 U12297 ( .A(n12324), .B(n12325), .ZN(n12162) );
  NAND2_X1 U12298 ( .A1(n12326), .A2(n12327), .ZN(n12324) );
  NAND2_X1 U12299 ( .A1(a_22_), .A2(n12323), .ZN(n12163) );
  NAND2_X1 U12300 ( .A1(n12101), .A2(n12328), .ZN(n12323) );
  NAND2_X1 U12301 ( .A1(n12100), .A2(n12102), .ZN(n12328) );
  NAND2_X1 U12302 ( .A1(n12329), .A2(n12330), .ZN(n12102) );
  NAND2_X1 U12303 ( .A1(b_19_), .A2(a_23_), .ZN(n12330) );
  INV_X1 U12304 ( .A(n12331), .ZN(n12329) );
  XOR2_X1 U12305 ( .A(n12332), .B(n12333), .Z(n12100) );
  XOR2_X1 U12306 ( .A(n12334), .B(n12335), .Z(n12332) );
  NAND2_X1 U12307 ( .A1(a_23_), .A2(n12331), .ZN(n12101) );
  NAND2_X1 U12308 ( .A1(n12336), .A2(n12337), .ZN(n12331) );
  NAND2_X1 U12309 ( .A1(n12110), .A2(n12338), .ZN(n12337) );
  INV_X1 U12310 ( .A(n12339), .ZN(n12338) );
  NOR2_X1 U12311 ( .A1(n12109), .A2(n12108), .ZN(n12339) );
  NOR2_X1 U12312 ( .A1(n8628), .A2(n8982), .ZN(n12110) );
  NAND2_X1 U12313 ( .A1(n12108), .A2(n12109), .ZN(n12336) );
  NAND2_X1 U12314 ( .A1(n12340), .A2(n12341), .ZN(n12109) );
  NAND2_X1 U12315 ( .A1(n12160), .A2(n12342), .ZN(n12341) );
  NAND2_X1 U12316 ( .A1(n12157), .A2(n12159), .ZN(n12342) );
  NOR2_X1 U12317 ( .A1(n8628), .A2(n8541), .ZN(n12160) );
  INV_X1 U12318 ( .A(n12343), .ZN(n12340) );
  NOR2_X1 U12319 ( .A1(n12159), .A2(n12157), .ZN(n12343) );
  XNOR2_X1 U12320 ( .A(n12344), .B(n12345), .ZN(n12157) );
  XNOR2_X1 U12321 ( .A(n12346), .B(n12347), .ZN(n12345) );
  NAND2_X1 U12322 ( .A1(n12348), .A2(n12349), .ZN(n12159) );
  NAND2_X1 U12323 ( .A1(n12119), .A2(n12350), .ZN(n12349) );
  NAND2_X1 U12324 ( .A1(n12122), .A2(n12121), .ZN(n12350) );
  XNOR2_X1 U12325 ( .A(n12351), .B(n12352), .ZN(n12119) );
  XOR2_X1 U12326 ( .A(n12353), .B(n12354), .Z(n12351) );
  INV_X1 U12327 ( .A(n12355), .ZN(n12348) );
  NOR2_X1 U12328 ( .A1(n12121), .A2(n12122), .ZN(n12355) );
  NOR2_X1 U12329 ( .A1(n8628), .A2(n9893), .ZN(n12122) );
  NAND2_X1 U12330 ( .A1(n12356), .A2(n12357), .ZN(n12121) );
  NAND2_X1 U12331 ( .A1(n12129), .A2(n12358), .ZN(n12357) );
  INV_X1 U12332 ( .A(n12359), .ZN(n12358) );
  NOR2_X1 U12333 ( .A1(n12128), .A2(n12127), .ZN(n12359) );
  NOR2_X1 U12334 ( .A1(n8628), .A2(n8512), .ZN(n12129) );
  NAND2_X1 U12335 ( .A1(n12127), .A2(n12128), .ZN(n12356) );
  NAND2_X1 U12336 ( .A1(n12360), .A2(n12361), .ZN(n12128) );
  NAND2_X1 U12337 ( .A1(n12155), .A2(n12362), .ZN(n12361) );
  INV_X1 U12338 ( .A(n12363), .ZN(n12362) );
  NOR2_X1 U12339 ( .A1(n12156), .A2(n12154), .ZN(n12363) );
  NOR2_X1 U12340 ( .A1(n8628), .A2(n8493), .ZN(n12155) );
  NAND2_X1 U12341 ( .A1(n12154), .A2(n12156), .ZN(n12360) );
  NAND2_X1 U12342 ( .A1(n12364), .A2(n12365), .ZN(n12156) );
  NAND2_X1 U12343 ( .A1(n12150), .A2(n12366), .ZN(n12365) );
  INV_X1 U12344 ( .A(n12367), .ZN(n12366) );
  NOR2_X1 U12345 ( .A1(n12151), .A2(n12152), .ZN(n12367) );
  NOR2_X1 U12346 ( .A1(n8628), .A2(n8473), .ZN(n12150) );
  NAND2_X1 U12347 ( .A1(n12152), .A2(n12151), .ZN(n12364) );
  NAND2_X1 U12348 ( .A1(n12368), .A2(n12369), .ZN(n12151) );
  NAND2_X1 U12349 ( .A1(b_17_), .A2(n12370), .ZN(n12369) );
  NAND2_X1 U12350 ( .A1(n8456), .A2(n12371), .ZN(n12370) );
  NAND2_X1 U12351 ( .A1(a_31_), .A2(n8987), .ZN(n12371) );
  NAND2_X1 U12352 ( .A1(b_18_), .A2(n12372), .ZN(n12368) );
  NAND2_X1 U12353 ( .A1(n8459), .A2(n12373), .ZN(n12372) );
  NAND2_X1 U12354 ( .A1(a_30_), .A2(n8660), .ZN(n12373) );
  NOR3_X1 U12355 ( .A1(n8628), .A2(n8979), .A3(n8987), .ZN(n12152) );
  XOR2_X1 U12356 ( .A(n12374), .B(n12375), .Z(n12154) );
  XOR2_X1 U12357 ( .A(n12376), .B(n12377), .Z(n12374) );
  XOR2_X1 U12358 ( .A(n12378), .B(n12379), .Z(n12127) );
  XOR2_X1 U12359 ( .A(n12380), .B(n12381), .Z(n12378) );
  XNOR2_X1 U12360 ( .A(n12382), .B(n12383), .ZN(n12108) );
  XNOR2_X1 U12361 ( .A(n12384), .B(n12385), .ZN(n12383) );
  XNOR2_X1 U12362 ( .A(n12386), .B(n12387), .ZN(n12086) );
  NAND2_X1 U12363 ( .A1(n12388), .A2(n12389), .ZN(n12386) );
  INV_X1 U12364 ( .A(n8625), .ZN(n8953) );
  NOR2_X1 U12365 ( .A1(n8628), .A2(n8630), .ZN(n8625) );
  XOR2_X1 U12366 ( .A(n12390), .B(n12391), .Z(n12053) );
  XOR2_X1 U12367 ( .A(n12392), .B(n12393), .Z(n12390) );
  NOR2_X1 U12368 ( .A1(n8680), .A2(n8987), .ZN(n12393) );
  XOR2_X1 U12369 ( .A(n12394), .B(n12395), .Z(n12044) );
  XOR2_X1 U12370 ( .A(n12396), .B(n12397), .Z(n12395) );
  NAND2_X1 U12371 ( .A1(b_18_), .A2(a_15_), .ZN(n12397) );
  XNOR2_X1 U12372 ( .A(n12398), .B(n12399), .ZN(n12036) );
  XNOR2_X1 U12373 ( .A(n12400), .B(n12401), .ZN(n12399) );
  XOR2_X1 U12374 ( .A(n12402), .B(n12403), .Z(n12011) );
  XOR2_X1 U12375 ( .A(n12404), .B(n12405), .Z(n12403) );
  XOR2_X1 U12376 ( .A(n12406), .B(n12407), .Z(n12177) );
  XNOR2_X1 U12377 ( .A(n12408), .B(n12409), .ZN(n12407) );
  XNOR2_X1 U12378 ( .A(n12410), .B(n12411), .ZN(n12181) );
  XNOR2_X1 U12379 ( .A(n12412), .B(n12413), .ZN(n12411) );
  NAND2_X1 U12380 ( .A1(b_18_), .A2(a_9_), .ZN(n12413) );
  XOR2_X1 U12381 ( .A(n12414), .B(n12415), .Z(n11994) );
  NAND2_X1 U12382 ( .A1(n12416), .A2(n12417), .ZN(n12414) );
  XNOR2_X1 U12383 ( .A(n12418), .B(n12419), .ZN(n11986) );
  NAND2_X1 U12384 ( .A1(n12420), .A2(n12421), .ZN(n12418) );
  XNOR2_X1 U12385 ( .A(n12422), .B(n12423), .ZN(n11978) );
  NAND2_X1 U12386 ( .A1(n12424), .A2(n12425), .ZN(n12422) );
  XOR2_X1 U12387 ( .A(n12426), .B(n12427), .Z(n12186) );
  XNOR2_X1 U12388 ( .A(n12428), .B(n12429), .ZN(n12427) );
  XNOR2_X1 U12389 ( .A(n12430), .B(n12431), .ZN(n12189) );
  XNOR2_X1 U12390 ( .A(n12432), .B(n12433), .ZN(n12431) );
  XNOR2_X1 U12391 ( .A(n12434), .B(n12435), .ZN(n12194) );
  XOR2_X1 U12392 ( .A(n12436), .B(n12437), .Z(n12435) );
  XOR2_X1 U12393 ( .A(n12438), .B(n12439), .Z(n11958) );
  XNOR2_X1 U12394 ( .A(n12440), .B(n12441), .ZN(n12438) );
  NOR2_X1 U12395 ( .A1(n8998), .A2(n8987), .ZN(n12441) );
  XOR2_X1 U12396 ( .A(n12442), .B(n12443), .Z(n12206) );
  NAND2_X1 U12397 ( .A1(n12444), .A2(n12445), .ZN(n12442) );
  NAND3_X1 U12398 ( .A1(n9091), .A2(n9092), .A3(n9090), .ZN(n9086) );
  NOR2_X1 U12399 ( .A1(n12446), .A2(n12447), .ZN(n9090) );
  INV_X1 U12400 ( .A(n12448), .ZN(n12447) );
  NAND2_X1 U12401 ( .A1(n12449), .A2(n12450), .ZN(n12448) );
  NAND2_X1 U12402 ( .A1(n12199), .A2(n12451), .ZN(n9092) );
  NAND2_X1 U12403 ( .A1(n12198), .A2(n12200), .ZN(n12451) );
  NAND2_X1 U12404 ( .A1(n12452), .A2(n12453), .ZN(n12200) );
  NAND2_X1 U12405 ( .A1(b_18_), .A2(a_0_), .ZN(n12453) );
  INV_X1 U12406 ( .A(n12454), .ZN(n12452) );
  XNOR2_X1 U12407 ( .A(n12455), .B(n12456), .ZN(n12198) );
  XNOR2_X1 U12408 ( .A(n12457), .B(n12458), .ZN(n12455) );
  NOR2_X1 U12409 ( .A1(n9731), .A2(n8660), .ZN(n12458) );
  NAND2_X1 U12410 ( .A1(a_0_), .A2(n12454), .ZN(n12199) );
  NAND2_X1 U12411 ( .A1(n12444), .A2(n12459), .ZN(n12454) );
  NAND2_X1 U12412 ( .A1(n12443), .A2(n12445), .ZN(n12459) );
  NAND2_X1 U12413 ( .A1(n12460), .A2(n12461), .ZN(n12445) );
  NAND2_X1 U12414 ( .A1(b_18_), .A2(a_1_), .ZN(n12461) );
  XOR2_X1 U12415 ( .A(n12462), .B(n12463), .Z(n12443) );
  XNOR2_X1 U12416 ( .A(n12464), .B(n12465), .ZN(n12463) );
  NAND2_X1 U12417 ( .A1(b_17_), .A2(a_2_), .ZN(n12465) );
  NAND2_X1 U12418 ( .A1(a_1_), .A2(n12466), .ZN(n12444) );
  INV_X1 U12419 ( .A(n12460), .ZN(n12466) );
  NOR2_X1 U12420 ( .A1(n12467), .A2(n12468), .ZN(n12460) );
  NOR3_X1 U12421 ( .A1(n8998), .A2(n12469), .A3(n8987), .ZN(n12468) );
  INV_X1 U12422 ( .A(n12470), .ZN(n12469) );
  NAND2_X1 U12423 ( .A1(n12439), .A2(n12440), .ZN(n12470) );
  NOR2_X1 U12424 ( .A1(n12439), .A2(n12440), .ZN(n12467) );
  NOR2_X1 U12425 ( .A1(n12471), .A2(n12472), .ZN(n12440) );
  NOR2_X1 U12426 ( .A1(n12437), .A2(n12473), .ZN(n12472) );
  NOR2_X1 U12427 ( .A1(n12434), .A2(n12436), .ZN(n12473) );
  NAND2_X1 U12428 ( .A1(b_18_), .A2(a_3_), .ZN(n12437) );
  INV_X1 U12429 ( .A(n12474), .ZN(n12471) );
  NAND2_X1 U12430 ( .A1(n12434), .A2(n12436), .ZN(n12474) );
  NAND2_X1 U12431 ( .A1(n12475), .A2(n12476), .ZN(n12436) );
  NAND2_X1 U12432 ( .A1(n12433), .A2(n12477), .ZN(n12476) );
  NAND2_X1 U12433 ( .A1(n12430), .A2(n12432), .ZN(n12477) );
  NOR2_X1 U12434 ( .A1(n8987), .A2(n8996), .ZN(n12433) );
  INV_X1 U12435 ( .A(n12478), .ZN(n12475) );
  NOR2_X1 U12436 ( .A1(n12432), .A2(n12430), .ZN(n12478) );
  XOR2_X1 U12437 ( .A(n12479), .B(n12480), .Z(n12430) );
  XOR2_X1 U12438 ( .A(n12481), .B(n12482), .Z(n12480) );
  NAND2_X1 U12439 ( .A1(b_17_), .A2(a_5_), .ZN(n12482) );
  NAND2_X1 U12440 ( .A1(n12483), .A2(n12484), .ZN(n12432) );
  NAND2_X1 U12441 ( .A1(n12426), .A2(n12485), .ZN(n12484) );
  NAND2_X1 U12442 ( .A1(n12429), .A2(n12428), .ZN(n12485) );
  XOR2_X1 U12443 ( .A(n12486), .B(n12487), .Z(n12426) );
  XOR2_X1 U12444 ( .A(n12488), .B(n12489), .Z(n12487) );
  NAND2_X1 U12445 ( .A1(b_17_), .A2(a_6_), .ZN(n12489) );
  INV_X1 U12446 ( .A(n12490), .ZN(n12483) );
  NOR2_X1 U12447 ( .A1(n12428), .A2(n12429), .ZN(n12490) );
  NOR2_X1 U12448 ( .A1(n8987), .A2(n8848), .ZN(n12429) );
  NAND2_X1 U12449 ( .A1(n12424), .A2(n12491), .ZN(n12428) );
  NAND2_X1 U12450 ( .A1(n12423), .A2(n12425), .ZN(n12491) );
  NAND2_X1 U12451 ( .A1(n12492), .A2(n12493), .ZN(n12425) );
  NAND2_X1 U12452 ( .A1(b_18_), .A2(a_6_), .ZN(n12493) );
  INV_X1 U12453 ( .A(n12494), .ZN(n12492) );
  XOR2_X1 U12454 ( .A(n12495), .B(n12496), .Z(n12423) );
  XNOR2_X1 U12455 ( .A(n12497), .B(n12498), .ZN(n12496) );
  NAND2_X1 U12456 ( .A1(b_17_), .A2(a_7_), .ZN(n12498) );
  NAND2_X1 U12457 ( .A1(a_6_), .A2(n12494), .ZN(n12424) );
  NAND2_X1 U12458 ( .A1(n12420), .A2(n12499), .ZN(n12494) );
  NAND2_X1 U12459 ( .A1(n12419), .A2(n12421), .ZN(n12499) );
  NAND2_X1 U12460 ( .A1(n12500), .A2(n12501), .ZN(n12421) );
  NAND2_X1 U12461 ( .A1(b_18_), .A2(a_7_), .ZN(n12501) );
  INV_X1 U12462 ( .A(n12502), .ZN(n12500) );
  XNOR2_X1 U12463 ( .A(n12503), .B(n12504), .ZN(n12419) );
  XNOR2_X1 U12464 ( .A(n12505), .B(n12506), .ZN(n12503) );
  NOR2_X1 U12465 ( .A1(n10513), .A2(n8660), .ZN(n12506) );
  NAND2_X1 U12466 ( .A1(a_7_), .A2(n12502), .ZN(n12420) );
  NAND2_X1 U12467 ( .A1(n12416), .A2(n12507), .ZN(n12502) );
  NAND2_X1 U12468 ( .A1(n12415), .A2(n12417), .ZN(n12507) );
  NAND2_X1 U12469 ( .A1(n12508), .A2(n12509), .ZN(n12417) );
  NAND2_X1 U12470 ( .A1(b_18_), .A2(a_8_), .ZN(n12509) );
  XNOR2_X1 U12471 ( .A(n12510), .B(n12511), .ZN(n12415) );
  XNOR2_X1 U12472 ( .A(n12512), .B(n12513), .ZN(n12510) );
  NOR2_X1 U12473 ( .A1(n8779), .A2(n8660), .ZN(n12513) );
  INV_X1 U12474 ( .A(n12514), .ZN(n12416) );
  NOR2_X1 U12475 ( .A1(n10513), .A2(n12508), .ZN(n12514) );
  NOR2_X1 U12476 ( .A1(n12515), .A2(n12516), .ZN(n12508) );
  INV_X1 U12477 ( .A(n12517), .ZN(n12516) );
  NAND3_X1 U12478 ( .A1(a_9_), .A2(n12518), .A3(b_18_), .ZN(n12517) );
  NAND2_X1 U12479 ( .A1(n12410), .A2(n12412), .ZN(n12518) );
  NOR2_X1 U12480 ( .A1(n12410), .A2(n12412), .ZN(n12515) );
  NOR2_X1 U12481 ( .A1(n12519), .A2(n12520), .ZN(n12412) );
  NOR2_X1 U12482 ( .A1(n12409), .A2(n12521), .ZN(n12520) );
  NOR2_X1 U12483 ( .A1(n12522), .A2(n12523), .ZN(n12521) );
  INV_X1 U12484 ( .A(n12406), .ZN(n12523) );
  INV_X1 U12485 ( .A(n12408), .ZN(n12522) );
  NAND2_X1 U12486 ( .A1(b_18_), .A2(a_10_), .ZN(n12409) );
  NOR2_X1 U12487 ( .A1(n12406), .A2(n12408), .ZN(n12519) );
  NOR2_X1 U12488 ( .A1(n12524), .A2(n12525), .ZN(n12408) );
  INV_X1 U12489 ( .A(n12526), .ZN(n12525) );
  NAND2_X1 U12490 ( .A1(n12405), .A2(n12527), .ZN(n12526) );
  NAND2_X1 U12491 ( .A1(n12404), .A2(n12402), .ZN(n12527) );
  NOR2_X1 U12492 ( .A1(n8987), .A2(n8749), .ZN(n12405) );
  NOR2_X1 U12493 ( .A1(n12402), .A2(n12404), .ZN(n12524) );
  NOR2_X1 U12494 ( .A1(n12528), .A2(n12529), .ZN(n12404) );
  INV_X1 U12495 ( .A(n12530), .ZN(n12529) );
  NAND3_X1 U12496 ( .A1(a_12_), .A2(n12531), .A3(b_18_), .ZN(n12530) );
  NAND2_X1 U12497 ( .A1(n12255), .A2(n12254), .ZN(n12531) );
  NOR2_X1 U12498 ( .A1(n12254), .A2(n12255), .ZN(n12528) );
  NOR2_X1 U12499 ( .A1(n12532), .A2(n12533), .ZN(n12255) );
  NOR3_X1 U12500 ( .A1(n8721), .A2(n12534), .A3(n8987), .ZN(n12533) );
  NOR2_X1 U12501 ( .A1(n12261), .A2(n12262), .ZN(n12534) );
  INV_X1 U12502 ( .A(n12535), .ZN(n12532) );
  NAND2_X1 U12503 ( .A1(n12262), .A2(n12261), .ZN(n12535) );
  XOR2_X1 U12504 ( .A(n12536), .B(n12537), .Z(n12261) );
  XOR2_X1 U12505 ( .A(n12538), .B(n12539), .Z(n12537) );
  NOR2_X1 U12506 ( .A1(n12540), .A2(n12541), .ZN(n12262) );
  INV_X1 U12507 ( .A(n12542), .ZN(n12541) );
  NAND2_X1 U12508 ( .A1(n12398), .A2(n12543), .ZN(n12542) );
  NAND2_X1 U12509 ( .A1(n12401), .A2(n12400), .ZN(n12543) );
  XOR2_X1 U12510 ( .A(n12544), .B(n12545), .Z(n12398) );
  XOR2_X1 U12511 ( .A(n12546), .B(n12547), .Z(n12545) );
  NAND2_X1 U12512 ( .A1(b_17_), .A2(a_15_), .ZN(n12547) );
  NOR2_X1 U12513 ( .A1(n12400), .A2(n12401), .ZN(n12540) );
  NOR2_X1 U12514 ( .A1(n8987), .A2(n8991), .ZN(n12401) );
  NAND2_X1 U12515 ( .A1(n12548), .A2(n12549), .ZN(n12400) );
  INV_X1 U12516 ( .A(n12550), .ZN(n12549) );
  NOR3_X1 U12517 ( .A1(n8692), .A2(n12551), .A3(n8987), .ZN(n12550) );
  NOR2_X1 U12518 ( .A1(n12396), .A2(n12394), .ZN(n12551) );
  NAND2_X1 U12519 ( .A1(n12394), .A2(n12396), .ZN(n12548) );
  NAND2_X1 U12520 ( .A1(n12552), .A2(n12553), .ZN(n12396) );
  NAND3_X1 U12521 ( .A1(a_16_), .A2(n12554), .A3(b_18_), .ZN(n12553) );
  INV_X1 U12522 ( .A(n12555), .ZN(n12554) );
  NOR2_X1 U12523 ( .A1(n12391), .A2(n12392), .ZN(n12555) );
  NAND2_X1 U12524 ( .A1(n12391), .A2(n12392), .ZN(n12552) );
  NAND2_X1 U12525 ( .A1(n12283), .A2(n12556), .ZN(n12392) );
  NAND2_X1 U12526 ( .A1(n12282), .A2(n12284), .ZN(n12556) );
  NAND2_X1 U12527 ( .A1(n12557), .A2(n12558), .ZN(n12284) );
  NAND2_X1 U12528 ( .A1(b_18_), .A2(a_17_), .ZN(n12558) );
  INV_X1 U12529 ( .A(n12559), .ZN(n12557) );
  XOR2_X1 U12530 ( .A(n12560), .B(n12561), .Z(n12282) );
  XOR2_X1 U12531 ( .A(n12562), .B(n12563), .Z(n12560) );
  NOR2_X1 U12532 ( .A1(n8988), .A2(n8660), .ZN(n12563) );
  NAND2_X1 U12533 ( .A1(a_17_), .A2(n12559), .ZN(n12283) );
  NAND2_X1 U12534 ( .A1(n12564), .A2(n12565), .ZN(n12559) );
  NAND2_X1 U12535 ( .A1(n12289), .A2(n12566), .ZN(n12565) );
  NAND2_X1 U12536 ( .A1(n12290), .A2(n8642), .ZN(n12566) );
  XNOR2_X1 U12537 ( .A(n12567), .B(n12568), .ZN(n12289) );
  XNOR2_X1 U12538 ( .A(n12569), .B(n12570), .ZN(n12568) );
  INV_X1 U12539 ( .A(n12571), .ZN(n12564) );
  NOR2_X1 U12540 ( .A1(n8642), .A2(n12290), .ZN(n12571) );
  NOR2_X1 U12541 ( .A1(n12572), .A2(n12573), .ZN(n12290) );
  INV_X1 U12542 ( .A(n12574), .ZN(n12573) );
  NAND3_X1 U12543 ( .A1(a_19_), .A2(n12575), .A3(b_18_), .ZN(n12574) );
  NAND2_X1 U12544 ( .A1(n12298), .A2(n12296), .ZN(n12575) );
  NOR2_X1 U12545 ( .A1(n12296), .A2(n12298), .ZN(n12572) );
  NOR2_X1 U12546 ( .A1(n12576), .A2(n12577), .ZN(n12298) );
  NOR3_X1 U12547 ( .A1(n8986), .A2(n12578), .A3(n8987), .ZN(n12577) );
  NOR2_X1 U12548 ( .A1(n12304), .A2(n12305), .ZN(n12578) );
  INV_X1 U12549 ( .A(n12579), .ZN(n12576) );
  NAND2_X1 U12550 ( .A1(n12304), .A2(n12305), .ZN(n12579) );
  NAND2_X1 U12551 ( .A1(n12580), .A2(n12581), .ZN(n12305) );
  NAND3_X1 U12552 ( .A1(a_21_), .A2(n12582), .A3(b_18_), .ZN(n12581) );
  INV_X1 U12553 ( .A(n12583), .ZN(n12582) );
  NOR2_X1 U12554 ( .A1(n12313), .A2(n12314), .ZN(n12583) );
  NAND2_X1 U12555 ( .A1(n12313), .A2(n12314), .ZN(n12580) );
  NAND2_X1 U12556 ( .A1(n12388), .A2(n12584), .ZN(n12314) );
  NAND2_X1 U12557 ( .A1(n12387), .A2(n12389), .ZN(n12584) );
  NAND2_X1 U12558 ( .A1(n12585), .A2(n12586), .ZN(n12389) );
  NAND2_X1 U12559 ( .A1(b_18_), .A2(a_22_), .ZN(n12586) );
  INV_X1 U12560 ( .A(n12587), .ZN(n12585) );
  XOR2_X1 U12561 ( .A(n12588), .B(n12589), .Z(n12387) );
  XOR2_X1 U12562 ( .A(n12590), .B(n12591), .Z(n12588) );
  NAND2_X1 U12563 ( .A1(a_22_), .A2(n12587), .ZN(n12388) );
  NAND2_X1 U12564 ( .A1(n12326), .A2(n12592), .ZN(n12587) );
  NAND2_X1 U12565 ( .A1(n12325), .A2(n12327), .ZN(n12592) );
  NAND2_X1 U12566 ( .A1(n12593), .A2(n12594), .ZN(n12327) );
  NAND2_X1 U12567 ( .A1(b_18_), .A2(a_23_), .ZN(n12594) );
  INV_X1 U12568 ( .A(n12595), .ZN(n12593) );
  XOR2_X1 U12569 ( .A(n12596), .B(n12597), .Z(n12325) );
  XOR2_X1 U12570 ( .A(n12598), .B(n12599), .Z(n12596) );
  NAND2_X1 U12571 ( .A1(a_23_), .A2(n12595), .ZN(n12326) );
  NAND2_X1 U12572 ( .A1(n12600), .A2(n12601), .ZN(n12595) );
  NAND2_X1 U12573 ( .A1(n12335), .A2(n12602), .ZN(n12601) );
  INV_X1 U12574 ( .A(n12603), .ZN(n12602) );
  NOR2_X1 U12575 ( .A1(n12333), .A2(n12334), .ZN(n12603) );
  NOR2_X1 U12576 ( .A1(n8987), .A2(n8982), .ZN(n12335) );
  NAND2_X1 U12577 ( .A1(n12333), .A2(n12334), .ZN(n12600) );
  NAND2_X1 U12578 ( .A1(n12604), .A2(n12605), .ZN(n12334) );
  NAND2_X1 U12579 ( .A1(n12385), .A2(n12606), .ZN(n12605) );
  NAND2_X1 U12580 ( .A1(n12382), .A2(n12384), .ZN(n12606) );
  NOR2_X1 U12581 ( .A1(n8987), .A2(n8541), .ZN(n12385) );
  INV_X1 U12582 ( .A(n12607), .ZN(n12604) );
  NOR2_X1 U12583 ( .A1(n12384), .A2(n12382), .ZN(n12607) );
  XNOR2_X1 U12584 ( .A(n12608), .B(n12609), .ZN(n12382) );
  XNOR2_X1 U12585 ( .A(n12610), .B(n12611), .ZN(n12609) );
  NAND2_X1 U12586 ( .A1(n12612), .A2(n12613), .ZN(n12384) );
  NAND2_X1 U12587 ( .A1(n12344), .A2(n12614), .ZN(n12613) );
  NAND2_X1 U12588 ( .A1(n12347), .A2(n12346), .ZN(n12614) );
  XNOR2_X1 U12589 ( .A(n12615), .B(n12616), .ZN(n12344) );
  XOR2_X1 U12590 ( .A(n12617), .B(n12618), .Z(n12615) );
  INV_X1 U12591 ( .A(n12619), .ZN(n12612) );
  NOR2_X1 U12592 ( .A1(n12346), .A2(n12347), .ZN(n12619) );
  NOR2_X1 U12593 ( .A1(n8987), .A2(n9893), .ZN(n12347) );
  NAND2_X1 U12594 ( .A1(n12620), .A2(n12621), .ZN(n12346) );
  NAND2_X1 U12595 ( .A1(n12354), .A2(n12622), .ZN(n12621) );
  INV_X1 U12596 ( .A(n12623), .ZN(n12622) );
  NOR2_X1 U12597 ( .A1(n12352), .A2(n12353), .ZN(n12623) );
  NOR2_X1 U12598 ( .A1(n8987), .A2(n8512), .ZN(n12354) );
  NAND2_X1 U12599 ( .A1(n12352), .A2(n12353), .ZN(n12620) );
  NAND2_X1 U12600 ( .A1(n12624), .A2(n12625), .ZN(n12353) );
  NAND2_X1 U12601 ( .A1(n12380), .A2(n12626), .ZN(n12625) );
  INV_X1 U12602 ( .A(n12627), .ZN(n12626) );
  NOR2_X1 U12603 ( .A1(n12381), .A2(n12379), .ZN(n12627) );
  NOR2_X1 U12604 ( .A1(n8987), .A2(n8493), .ZN(n12380) );
  NAND2_X1 U12605 ( .A1(n12379), .A2(n12381), .ZN(n12624) );
  NAND2_X1 U12606 ( .A1(n12628), .A2(n12629), .ZN(n12381) );
  NAND2_X1 U12607 ( .A1(n12375), .A2(n12630), .ZN(n12629) );
  INV_X1 U12608 ( .A(n12631), .ZN(n12630) );
  NOR2_X1 U12609 ( .A1(n12376), .A2(n12377), .ZN(n12631) );
  NOR2_X1 U12610 ( .A1(n8987), .A2(n8473), .ZN(n12375) );
  NAND2_X1 U12611 ( .A1(n12377), .A2(n12376), .ZN(n12628) );
  NAND2_X1 U12612 ( .A1(n12632), .A2(n12633), .ZN(n12376) );
  NAND2_X1 U12613 ( .A1(b_16_), .A2(n12634), .ZN(n12633) );
  NAND2_X1 U12614 ( .A1(n8456), .A2(n12635), .ZN(n12634) );
  NAND2_X1 U12615 ( .A1(a_31_), .A2(n8660), .ZN(n12635) );
  NAND2_X1 U12616 ( .A1(b_17_), .A2(n12636), .ZN(n12632) );
  NAND2_X1 U12617 ( .A1(n8459), .A2(n12637), .ZN(n12636) );
  NAND2_X1 U12618 ( .A1(a_30_), .A2(n8989), .ZN(n12637) );
  NOR3_X1 U12619 ( .A1(n8987), .A2(n8979), .A3(n8660), .ZN(n12377) );
  INV_X1 U12620 ( .A(b_18_), .ZN(n8987) );
  XOR2_X1 U12621 ( .A(n12638), .B(n12639), .Z(n12379) );
  XOR2_X1 U12622 ( .A(n12640), .B(n12641), .Z(n12638) );
  XOR2_X1 U12623 ( .A(n12642), .B(n12643), .Z(n12352) );
  XOR2_X1 U12624 ( .A(n12644), .B(n12645), .Z(n12642) );
  XNOR2_X1 U12625 ( .A(n12646), .B(n12647), .ZN(n12333) );
  XNOR2_X1 U12626 ( .A(n12648), .B(n12649), .ZN(n12647) );
  XNOR2_X1 U12627 ( .A(n12650), .B(n12651), .ZN(n12313) );
  XNOR2_X1 U12628 ( .A(n12652), .B(n12653), .ZN(n12651) );
  XNOR2_X1 U12629 ( .A(n12654), .B(n12655), .ZN(n12304) );
  NAND2_X1 U12630 ( .A1(n12656), .A2(n12657), .ZN(n12654) );
  XOR2_X1 U12631 ( .A(n12658), .B(n12659), .Z(n12296) );
  XOR2_X1 U12632 ( .A(n12660), .B(n12661), .Z(n12658) );
  NAND2_X1 U12633 ( .A1(b_18_), .A2(a_18_), .ZN(n8642) );
  XOR2_X1 U12634 ( .A(n12662), .B(n12663), .Z(n12391) );
  XNOR2_X1 U12635 ( .A(n12664), .B(n8657), .ZN(n12663) );
  XNOR2_X1 U12636 ( .A(n12665), .B(n12666), .ZN(n12394) );
  NAND2_X1 U12637 ( .A1(n12667), .A2(n12668), .ZN(n12665) );
  XNOR2_X1 U12638 ( .A(n12669), .B(n12670), .ZN(n12254) );
  XNOR2_X1 U12639 ( .A(n12671), .B(n12672), .ZN(n12669) );
  XOR2_X1 U12640 ( .A(n12673), .B(n12674), .Z(n12402) );
  XNOR2_X1 U12641 ( .A(n12675), .B(n12676), .ZN(n12673) );
  NOR2_X1 U12642 ( .A1(n8739), .A2(n8660), .ZN(n12676) );
  XNOR2_X1 U12643 ( .A(n12677), .B(n12678), .ZN(n12406) );
  XNOR2_X1 U12644 ( .A(n12679), .B(n12680), .ZN(n12678) );
  NAND2_X1 U12645 ( .A1(b_17_), .A2(a_11_), .ZN(n12680) );
  XOR2_X1 U12646 ( .A(n12681), .B(n12682), .Z(n12410) );
  XNOR2_X1 U12647 ( .A(n12683), .B(n12684), .ZN(n12681) );
  NOR2_X1 U12648 ( .A1(n8769), .A2(n8660), .ZN(n12684) );
  XOR2_X1 U12649 ( .A(n12685), .B(n12686), .Z(n12434) );
  XNOR2_X1 U12650 ( .A(n12687), .B(n12688), .ZN(n12686) );
  NAND2_X1 U12651 ( .A1(b_17_), .A2(a_4_), .ZN(n12688) );
  XOR2_X1 U12652 ( .A(n12689), .B(n12690), .Z(n12439) );
  XNOR2_X1 U12653 ( .A(n12691), .B(n12692), .ZN(n12689) );
  NOR2_X1 U12654 ( .A1(n8877), .A2(n8660), .ZN(n12692) );
  XOR2_X1 U12655 ( .A(n12693), .B(n12694), .Z(n9091) );
  XNOR2_X1 U12656 ( .A(n12695), .B(n12696), .ZN(n12694) );
  INV_X1 U12657 ( .A(n12697), .ZN(n9097) );
  NOR2_X1 U12658 ( .A1(n12698), .A2(n12446), .ZN(n12697) );
  NAND2_X1 U12659 ( .A1(n12446), .A2(n12698), .ZN(n9096) );
  XOR2_X1 U12660 ( .A(n12699), .B(n12700), .Z(n12698) );
  NOR2_X1 U12661 ( .A1(n12450), .A2(n12449), .ZN(n12446) );
  XOR2_X1 U12662 ( .A(n12701), .B(n12702), .Z(n12449) );
  NAND2_X1 U12663 ( .A1(n12703), .A2(n12704), .ZN(n12701) );
  NAND2_X1 U12664 ( .A1(n12705), .A2(n12706), .ZN(n12450) );
  NAND2_X1 U12665 ( .A1(n12693), .A2(n12707), .ZN(n12706) );
  INV_X1 U12666 ( .A(n12708), .ZN(n12707) );
  NOR2_X1 U12667 ( .A1(n12696), .A2(n12695), .ZN(n12708) );
  XOR2_X1 U12668 ( .A(n12709), .B(n12710), .Z(n12693) );
  NAND2_X1 U12669 ( .A1(n12711), .A2(n12712), .ZN(n12709) );
  NAND2_X1 U12670 ( .A1(n12695), .A2(n12696), .ZN(n12705) );
  NAND2_X1 U12671 ( .A1(b_17_), .A2(a_0_), .ZN(n12696) );
  NOR2_X1 U12672 ( .A1(n12713), .A2(n12714), .ZN(n12695) );
  INV_X1 U12673 ( .A(n12715), .ZN(n12714) );
  NAND3_X1 U12674 ( .A1(a_1_), .A2(n12716), .A3(b_17_), .ZN(n12715) );
  NAND2_X1 U12675 ( .A1(n12457), .A2(n12456), .ZN(n12716) );
  NOR2_X1 U12676 ( .A1(n12456), .A2(n12457), .ZN(n12713) );
  NOR2_X1 U12677 ( .A1(n12717), .A2(n12718), .ZN(n12457) );
  NOR3_X1 U12678 ( .A1(n8998), .A2(n12719), .A3(n8660), .ZN(n12718) );
  INV_X1 U12679 ( .A(n12720), .ZN(n12719) );
  NAND2_X1 U12680 ( .A1(n12464), .A2(n12462), .ZN(n12720) );
  NOR2_X1 U12681 ( .A1(n12462), .A2(n12464), .ZN(n12717) );
  NOR2_X1 U12682 ( .A1(n12721), .A2(n12722), .ZN(n12464) );
  INV_X1 U12683 ( .A(n12723), .ZN(n12722) );
  NAND3_X1 U12684 ( .A1(a_3_), .A2(n12724), .A3(b_17_), .ZN(n12723) );
  NAND2_X1 U12685 ( .A1(n12691), .A2(n12690), .ZN(n12724) );
  NOR2_X1 U12686 ( .A1(n12690), .A2(n12691), .ZN(n12721) );
  NOR2_X1 U12687 ( .A1(n12725), .A2(n12726), .ZN(n12691) );
  INV_X1 U12688 ( .A(n12727), .ZN(n12726) );
  NAND3_X1 U12689 ( .A1(a_4_), .A2(n12728), .A3(b_17_), .ZN(n12727) );
  NAND2_X1 U12690 ( .A1(n12687), .A2(n12685), .ZN(n12728) );
  NOR2_X1 U12691 ( .A1(n12685), .A2(n12687), .ZN(n12725) );
  NOR2_X1 U12692 ( .A1(n12729), .A2(n12730), .ZN(n12687) );
  NOR3_X1 U12693 ( .A1(n8848), .A2(n12731), .A3(n8660), .ZN(n12730) );
  NOR2_X1 U12694 ( .A1(n12481), .A2(n12479), .ZN(n12731) );
  INV_X1 U12695 ( .A(n12732), .ZN(n12729) );
  NAND2_X1 U12696 ( .A1(n12479), .A2(n12481), .ZN(n12732) );
  NAND2_X1 U12697 ( .A1(n12733), .A2(n12734), .ZN(n12481) );
  INV_X1 U12698 ( .A(n12735), .ZN(n12734) );
  NOR3_X1 U12699 ( .A1(n8994), .A2(n12736), .A3(n8660), .ZN(n12735) );
  NOR2_X1 U12700 ( .A1(n12486), .A2(n12488), .ZN(n12736) );
  NAND2_X1 U12701 ( .A1(n12486), .A2(n12488), .ZN(n12733) );
  NAND2_X1 U12702 ( .A1(n12737), .A2(n12738), .ZN(n12488) );
  NAND3_X1 U12703 ( .A1(a_7_), .A2(n12739), .A3(b_17_), .ZN(n12738) );
  NAND2_X1 U12704 ( .A1(n12497), .A2(n12495), .ZN(n12739) );
  INV_X1 U12705 ( .A(n12740), .ZN(n12737) );
  NOR2_X1 U12706 ( .A1(n12495), .A2(n12497), .ZN(n12740) );
  NOR2_X1 U12707 ( .A1(n12741), .A2(n12742), .ZN(n12497) );
  INV_X1 U12708 ( .A(n12743), .ZN(n12742) );
  NAND3_X1 U12709 ( .A1(a_8_), .A2(n12744), .A3(b_17_), .ZN(n12743) );
  NAND2_X1 U12710 ( .A1(n12505), .A2(n12504), .ZN(n12744) );
  NOR2_X1 U12711 ( .A1(n12504), .A2(n12505), .ZN(n12741) );
  NOR2_X1 U12712 ( .A1(n12745), .A2(n12746), .ZN(n12505) );
  NOR3_X1 U12713 ( .A1(n8779), .A2(n12747), .A3(n8660), .ZN(n12746) );
  INV_X1 U12714 ( .A(n12748), .ZN(n12747) );
  NAND2_X1 U12715 ( .A1(n12511), .A2(n12512), .ZN(n12748) );
  NOR2_X1 U12716 ( .A1(n12511), .A2(n12512), .ZN(n12745) );
  NOR2_X1 U12717 ( .A1(n12749), .A2(n12750), .ZN(n12512) );
  INV_X1 U12718 ( .A(n12751), .ZN(n12750) );
  NAND3_X1 U12719 ( .A1(a_10_), .A2(n12752), .A3(b_17_), .ZN(n12751) );
  NAND2_X1 U12720 ( .A1(n12683), .A2(n12682), .ZN(n12752) );
  NOR2_X1 U12721 ( .A1(n12682), .A2(n12683), .ZN(n12749) );
  NOR2_X1 U12722 ( .A1(n12753), .A2(n12754), .ZN(n12683) );
  NOR3_X1 U12723 ( .A1(n8749), .A2(n12755), .A3(n8660), .ZN(n12754) );
  INV_X1 U12724 ( .A(n12756), .ZN(n12755) );
  NAND2_X1 U12725 ( .A1(n12677), .A2(n12679), .ZN(n12756) );
  NOR2_X1 U12726 ( .A1(n12677), .A2(n12679), .ZN(n12753) );
  NOR2_X1 U12727 ( .A1(n12757), .A2(n12758), .ZN(n12679) );
  INV_X1 U12728 ( .A(n12759), .ZN(n12758) );
  NAND3_X1 U12729 ( .A1(a_12_), .A2(n12760), .A3(b_17_), .ZN(n12759) );
  NAND2_X1 U12730 ( .A1(n12674), .A2(n12675), .ZN(n12760) );
  NOR2_X1 U12731 ( .A1(n12674), .A2(n12675), .ZN(n12757) );
  NOR2_X1 U12732 ( .A1(n12761), .A2(n12762), .ZN(n12675) );
  NOR2_X1 U12733 ( .A1(n12671), .A2(n12763), .ZN(n12762) );
  NOR2_X1 U12734 ( .A1(n12670), .A2(n12672), .ZN(n12763) );
  NAND2_X1 U12735 ( .A1(b_17_), .A2(a_13_), .ZN(n12671) );
  INV_X1 U12736 ( .A(n12764), .ZN(n12761) );
  NAND2_X1 U12737 ( .A1(n12670), .A2(n12672), .ZN(n12764) );
  NAND2_X1 U12738 ( .A1(n12765), .A2(n12766), .ZN(n12672) );
  NAND2_X1 U12739 ( .A1(n12539), .A2(n12767), .ZN(n12766) );
  NAND2_X1 U12740 ( .A1(n12538), .A2(n12536), .ZN(n12767) );
  NOR2_X1 U12741 ( .A1(n8660), .A2(n8991), .ZN(n12539) );
  INV_X1 U12742 ( .A(n12768), .ZN(n12765) );
  NOR2_X1 U12743 ( .A1(n12536), .A2(n12538), .ZN(n12768) );
  NOR2_X1 U12744 ( .A1(n12769), .A2(n12770), .ZN(n12538) );
  NOR3_X1 U12745 ( .A1(n8692), .A2(n12771), .A3(n8660), .ZN(n12770) );
  NOR2_X1 U12746 ( .A1(n12546), .A2(n12544), .ZN(n12771) );
  INV_X1 U12747 ( .A(n12772), .ZN(n12769) );
  NAND2_X1 U12748 ( .A1(n12544), .A2(n12546), .ZN(n12772) );
  NAND2_X1 U12749 ( .A1(n12667), .A2(n12773), .ZN(n12546) );
  NAND2_X1 U12750 ( .A1(n12666), .A2(n12668), .ZN(n12773) );
  NAND2_X1 U12751 ( .A1(n12774), .A2(n12775), .ZN(n12668) );
  NAND2_X1 U12752 ( .A1(b_17_), .A2(a_16_), .ZN(n12774) );
  XOR2_X1 U12753 ( .A(n12776), .B(n12777), .Z(n12666) );
  XOR2_X1 U12754 ( .A(n12778), .B(n12779), .Z(n12776) );
  NOR2_X1 U12755 ( .A1(n8662), .A2(n8989), .ZN(n12779) );
  INV_X1 U12756 ( .A(n12780), .ZN(n12667) );
  NOR2_X1 U12757 ( .A1(n12775), .A2(n8680), .ZN(n12780) );
  NAND2_X1 U12758 ( .A1(n12781), .A2(n12782), .ZN(n12775) );
  NAND2_X1 U12759 ( .A1(n12662), .A2(n12783), .ZN(n12782) );
  NAND2_X1 U12760 ( .A1(n8657), .A2(n12664), .ZN(n12783) );
  XNOR2_X1 U12761 ( .A(n12784), .B(n12785), .ZN(n12662) );
  XNOR2_X1 U12762 ( .A(n12786), .B(n12787), .ZN(n12785) );
  NAND2_X1 U12763 ( .A1(n12788), .A2(n8949), .ZN(n12781) );
  INV_X1 U12764 ( .A(n8657), .ZN(n8949) );
  NOR2_X1 U12765 ( .A1(n8660), .A2(n8662), .ZN(n8657) );
  INV_X1 U12766 ( .A(n12664), .ZN(n12788) );
  NAND2_X1 U12767 ( .A1(n12789), .A2(n12790), .ZN(n12664) );
  NAND3_X1 U12768 ( .A1(a_18_), .A2(n12791), .A3(b_17_), .ZN(n12790) );
  INV_X1 U12769 ( .A(n12792), .ZN(n12791) );
  NOR2_X1 U12770 ( .A1(n12561), .A2(n12562), .ZN(n12792) );
  NAND2_X1 U12771 ( .A1(n12561), .A2(n12562), .ZN(n12789) );
  NAND2_X1 U12772 ( .A1(n12793), .A2(n12794), .ZN(n12562) );
  NAND2_X1 U12773 ( .A1(n12570), .A2(n12795), .ZN(n12794) );
  NAND2_X1 U12774 ( .A1(n12567), .A2(n12569), .ZN(n12795) );
  NOR2_X1 U12775 ( .A1(n8660), .A2(n8630), .ZN(n12570) );
  INV_X1 U12776 ( .A(n12796), .ZN(n12793) );
  NOR2_X1 U12777 ( .A1(n12569), .A2(n12567), .ZN(n12796) );
  XOR2_X1 U12778 ( .A(n12797), .B(n12798), .Z(n12567) );
  XNOR2_X1 U12779 ( .A(n12799), .B(n12800), .ZN(n12798) );
  NAND2_X1 U12780 ( .A1(n12801), .A2(n12802), .ZN(n12569) );
  NAND2_X1 U12781 ( .A1(n12659), .A2(n12803), .ZN(n12802) );
  NAND2_X1 U12782 ( .A1(n12661), .A2(n12660), .ZN(n12803) );
  XOR2_X1 U12783 ( .A(n12804), .B(n12805), .Z(n12659) );
  XOR2_X1 U12784 ( .A(n12806), .B(n12807), .Z(n12804) );
  INV_X1 U12785 ( .A(n12808), .ZN(n12801) );
  NOR2_X1 U12786 ( .A1(n12660), .A2(n12661), .ZN(n12808) );
  NOR2_X1 U12787 ( .A1(n8660), .A2(n8986), .ZN(n12661) );
  NAND2_X1 U12788 ( .A1(n12656), .A2(n12809), .ZN(n12660) );
  NAND2_X1 U12789 ( .A1(n12655), .A2(n12657), .ZN(n12809) );
  NAND2_X1 U12790 ( .A1(n12810), .A2(n12811), .ZN(n12657) );
  NAND2_X1 U12791 ( .A1(b_17_), .A2(a_21_), .ZN(n12811) );
  INV_X1 U12792 ( .A(n12812), .ZN(n12810) );
  XNOR2_X1 U12793 ( .A(n12813), .B(n12814), .ZN(n12655) );
  NAND2_X1 U12794 ( .A1(n12815), .A2(n12816), .ZN(n12813) );
  NAND2_X1 U12795 ( .A1(a_21_), .A2(n12812), .ZN(n12656) );
  NAND2_X1 U12796 ( .A1(n12817), .A2(n12818), .ZN(n12812) );
  NAND2_X1 U12797 ( .A1(n12653), .A2(n12819), .ZN(n12818) );
  INV_X1 U12798 ( .A(n12820), .ZN(n12819) );
  NOR2_X1 U12799 ( .A1(n12652), .A2(n12650), .ZN(n12820) );
  NOR2_X1 U12800 ( .A1(n8660), .A2(n8984), .ZN(n12653) );
  NAND2_X1 U12801 ( .A1(n12650), .A2(n12652), .ZN(n12817) );
  NAND2_X1 U12802 ( .A1(n12821), .A2(n12822), .ZN(n12652) );
  NAND2_X1 U12803 ( .A1(n12591), .A2(n12823), .ZN(n12822) );
  INV_X1 U12804 ( .A(n12824), .ZN(n12823) );
  NOR2_X1 U12805 ( .A1(n12590), .A2(n12589), .ZN(n12824) );
  NOR2_X1 U12806 ( .A1(n8660), .A2(n8572), .ZN(n12591) );
  NAND2_X1 U12807 ( .A1(n12589), .A2(n12590), .ZN(n12821) );
  NAND2_X1 U12808 ( .A1(n12825), .A2(n12826), .ZN(n12590) );
  NAND2_X1 U12809 ( .A1(n12599), .A2(n12827), .ZN(n12826) );
  INV_X1 U12810 ( .A(n12828), .ZN(n12827) );
  NOR2_X1 U12811 ( .A1(n12597), .A2(n12598), .ZN(n12828) );
  NOR2_X1 U12812 ( .A1(n8660), .A2(n8982), .ZN(n12599) );
  NAND2_X1 U12813 ( .A1(n12597), .A2(n12598), .ZN(n12825) );
  NAND2_X1 U12814 ( .A1(n12829), .A2(n12830), .ZN(n12598) );
  NAND2_X1 U12815 ( .A1(n12649), .A2(n12831), .ZN(n12830) );
  NAND2_X1 U12816 ( .A1(n12646), .A2(n12648), .ZN(n12831) );
  NOR2_X1 U12817 ( .A1(n8660), .A2(n8541), .ZN(n12649) );
  INV_X1 U12818 ( .A(n12832), .ZN(n12829) );
  NOR2_X1 U12819 ( .A1(n12648), .A2(n12646), .ZN(n12832) );
  XNOR2_X1 U12820 ( .A(n12833), .B(n12834), .ZN(n12646) );
  XNOR2_X1 U12821 ( .A(n12835), .B(n12836), .ZN(n12834) );
  NAND2_X1 U12822 ( .A1(n12837), .A2(n12838), .ZN(n12648) );
  NAND2_X1 U12823 ( .A1(n12608), .A2(n12839), .ZN(n12838) );
  NAND2_X1 U12824 ( .A1(n12611), .A2(n12610), .ZN(n12839) );
  XNOR2_X1 U12825 ( .A(n12840), .B(n12841), .ZN(n12608) );
  XOR2_X1 U12826 ( .A(n12842), .B(n12843), .Z(n12840) );
  INV_X1 U12827 ( .A(n12844), .ZN(n12837) );
  NOR2_X1 U12828 ( .A1(n12610), .A2(n12611), .ZN(n12844) );
  NOR2_X1 U12829 ( .A1(n8660), .A2(n9893), .ZN(n12611) );
  NAND2_X1 U12830 ( .A1(n12845), .A2(n12846), .ZN(n12610) );
  NAND2_X1 U12831 ( .A1(n12618), .A2(n12847), .ZN(n12846) );
  INV_X1 U12832 ( .A(n12848), .ZN(n12847) );
  NOR2_X1 U12833 ( .A1(n12616), .A2(n12617), .ZN(n12848) );
  NOR2_X1 U12834 ( .A1(n8660), .A2(n8512), .ZN(n12618) );
  NAND2_X1 U12835 ( .A1(n12616), .A2(n12617), .ZN(n12845) );
  NAND2_X1 U12836 ( .A1(n12849), .A2(n12850), .ZN(n12617) );
  NAND2_X1 U12837 ( .A1(n12644), .A2(n12851), .ZN(n12850) );
  INV_X1 U12838 ( .A(n12852), .ZN(n12851) );
  NOR2_X1 U12839 ( .A1(n12645), .A2(n12643), .ZN(n12852) );
  NOR2_X1 U12840 ( .A1(n8660), .A2(n8493), .ZN(n12644) );
  NAND2_X1 U12841 ( .A1(n12643), .A2(n12645), .ZN(n12849) );
  NAND2_X1 U12842 ( .A1(n12853), .A2(n12854), .ZN(n12645) );
  NAND2_X1 U12843 ( .A1(n12639), .A2(n12855), .ZN(n12854) );
  INV_X1 U12844 ( .A(n12856), .ZN(n12855) );
  NOR2_X1 U12845 ( .A1(n12640), .A2(n12641), .ZN(n12856) );
  NOR2_X1 U12846 ( .A1(n8660), .A2(n8473), .ZN(n12639) );
  NAND2_X1 U12847 ( .A1(n12641), .A2(n12640), .ZN(n12853) );
  NAND2_X1 U12848 ( .A1(n12857), .A2(n12858), .ZN(n12640) );
  NAND2_X1 U12849 ( .A1(b_15_), .A2(n12859), .ZN(n12858) );
  NAND2_X1 U12850 ( .A1(n8456), .A2(n12860), .ZN(n12859) );
  NAND2_X1 U12851 ( .A1(a_31_), .A2(n8989), .ZN(n12860) );
  NAND2_X1 U12852 ( .A1(b_16_), .A2(n12861), .ZN(n12857) );
  NAND2_X1 U12853 ( .A1(n8459), .A2(n12862), .ZN(n12861) );
  NAND2_X1 U12854 ( .A1(a_30_), .A2(n8690), .ZN(n12862) );
  NOR3_X1 U12855 ( .A1(n8660), .A2(n8979), .A3(n8989), .ZN(n12641) );
  XOR2_X1 U12856 ( .A(n12863), .B(n12864), .Z(n12643) );
  XOR2_X1 U12857 ( .A(n12865), .B(n12866), .Z(n12863) );
  XOR2_X1 U12858 ( .A(n12867), .B(n12868), .Z(n12616) );
  XOR2_X1 U12859 ( .A(n12869), .B(n12870), .Z(n12867) );
  XNOR2_X1 U12860 ( .A(n12871), .B(n12872), .ZN(n12597) );
  XNOR2_X1 U12861 ( .A(n12873), .B(n12874), .ZN(n12872) );
  XOR2_X1 U12862 ( .A(n12875), .B(n12876), .Z(n12589) );
  XOR2_X1 U12863 ( .A(n12877), .B(n12878), .Z(n12875) );
  XNOR2_X1 U12864 ( .A(n12879), .B(n12880), .ZN(n12650) );
  NAND2_X1 U12865 ( .A1(n12881), .A2(n12882), .ZN(n12879) );
  XOR2_X1 U12866 ( .A(n12883), .B(n12884), .Z(n12561) );
  XNOR2_X1 U12867 ( .A(n12885), .B(n12886), .ZN(n12884) );
  NAND2_X1 U12868 ( .A1(b_16_), .A2(a_19_), .ZN(n12886) );
  XNOR2_X1 U12869 ( .A(n12887), .B(n12888), .ZN(n12544) );
  XOR2_X1 U12870 ( .A(n12889), .B(n8674), .Z(n12887) );
  XOR2_X1 U12871 ( .A(n12890), .B(n12891), .Z(n12536) );
  XOR2_X1 U12872 ( .A(n12892), .B(n12893), .Z(n12891) );
  NAND2_X1 U12873 ( .A1(b_16_), .A2(a_15_), .ZN(n12893) );
  XOR2_X1 U12874 ( .A(n12894), .B(n12895), .Z(n12670) );
  XNOR2_X1 U12875 ( .A(n12896), .B(n12897), .ZN(n12895) );
  NAND2_X1 U12876 ( .A1(b_16_), .A2(a_14_), .ZN(n12897) );
  XOR2_X1 U12877 ( .A(n12898), .B(n12899), .Z(n12674) );
  XNOR2_X1 U12878 ( .A(n12900), .B(n12901), .ZN(n12898) );
  XOR2_X1 U12879 ( .A(n12902), .B(n12903), .Z(n12677) );
  XNOR2_X1 U12880 ( .A(n12904), .B(n12905), .ZN(n12902) );
  XNOR2_X1 U12881 ( .A(n12906), .B(n12907), .ZN(n12682) );
  XNOR2_X1 U12882 ( .A(n12908), .B(n12909), .ZN(n12906) );
  NOR2_X1 U12883 ( .A1(n8749), .A2(n8989), .ZN(n12909) );
  XOR2_X1 U12884 ( .A(n12910), .B(n12911), .Z(n12511) );
  NAND2_X1 U12885 ( .A1(n12912), .A2(n12913), .ZN(n12910) );
  XNOR2_X1 U12886 ( .A(n12914), .B(n12915), .ZN(n12504) );
  XOR2_X1 U12887 ( .A(n12916), .B(n12917), .Z(n12914) );
  NOR2_X1 U12888 ( .A1(n8779), .A2(n8989), .ZN(n12917) );
  XOR2_X1 U12889 ( .A(n12918), .B(n12919), .Z(n12495) );
  NAND2_X1 U12890 ( .A1(n12920), .A2(n12921), .ZN(n12918) );
  XNOR2_X1 U12891 ( .A(n12922), .B(n12923), .ZN(n12486) );
  NAND2_X1 U12892 ( .A1(n12924), .A2(n12925), .ZN(n12922) );
  XNOR2_X1 U12893 ( .A(n12926), .B(n12927), .ZN(n12479) );
  NAND2_X1 U12894 ( .A1(n12928), .A2(n12929), .ZN(n12926) );
  XNOR2_X1 U12895 ( .A(n12930), .B(n12931), .ZN(n12685) );
  XOR2_X1 U12896 ( .A(n12932), .B(n12933), .Z(n12930) );
  XNOR2_X1 U12897 ( .A(n12934), .B(n12935), .ZN(n12690) );
  XOR2_X1 U12898 ( .A(n12936), .B(n12937), .Z(n12934) );
  NOR2_X1 U12899 ( .A1(n8996), .A2(n8989), .ZN(n12937) );
  XOR2_X1 U12900 ( .A(n12938), .B(n12939), .Z(n12462) );
  NAND2_X1 U12901 ( .A1(n12940), .A2(n12941), .ZN(n12938) );
  XOR2_X1 U12902 ( .A(n12942), .B(n12943), .Z(n12456) );
  NAND2_X1 U12903 ( .A1(n12944), .A2(n12945), .ZN(n12942) );
  NAND2_X1 U12904 ( .A1(n12946), .A2(n12947), .ZN(n9102) );
  NAND2_X1 U12905 ( .A1(n12948), .A2(n12949), .ZN(n12947) );
  NAND2_X1 U12906 ( .A1(n12699), .A2(n12700), .ZN(n12946) );
  NAND4_X1 U12907 ( .A1(n12699), .A2(n12948), .A3(n12700), .A4(n12949), .ZN(
        n9101) );
  NAND2_X1 U12908 ( .A1(n12703), .A2(n12950), .ZN(n12700) );
  NAND2_X1 U12909 ( .A1(n12702), .A2(n12704), .ZN(n12950) );
  NAND2_X1 U12910 ( .A1(n12951), .A2(n12952), .ZN(n12704) );
  NAND2_X1 U12911 ( .A1(b_16_), .A2(a_0_), .ZN(n12952) );
  INV_X1 U12912 ( .A(n12953), .ZN(n12951) );
  XOR2_X1 U12913 ( .A(n12954), .B(n12955), .Z(n12702) );
  XNOR2_X1 U12914 ( .A(n12956), .B(n12957), .ZN(n12955) );
  NAND2_X1 U12915 ( .A1(a_0_), .A2(n12953), .ZN(n12703) );
  NAND2_X1 U12916 ( .A1(n12711), .A2(n12958), .ZN(n12953) );
  NAND2_X1 U12917 ( .A1(n12710), .A2(n12712), .ZN(n12958) );
  NAND2_X1 U12918 ( .A1(n12959), .A2(n12960), .ZN(n12712) );
  NAND2_X1 U12919 ( .A1(b_16_), .A2(a_1_), .ZN(n12960) );
  INV_X1 U12920 ( .A(n12961), .ZN(n12959) );
  XOR2_X1 U12921 ( .A(n12962), .B(n12963), .Z(n12710) );
  XOR2_X1 U12922 ( .A(n12964), .B(n12965), .Z(n12962) );
  NOR2_X1 U12923 ( .A1(n8998), .A2(n8690), .ZN(n12965) );
  NAND2_X1 U12924 ( .A1(a_1_), .A2(n12961), .ZN(n12711) );
  NAND2_X1 U12925 ( .A1(n12944), .A2(n12966), .ZN(n12961) );
  NAND2_X1 U12926 ( .A1(n12943), .A2(n12945), .ZN(n12966) );
  NAND2_X1 U12927 ( .A1(n12967), .A2(n12968), .ZN(n12945) );
  NAND2_X1 U12928 ( .A1(b_16_), .A2(a_2_), .ZN(n12968) );
  INV_X1 U12929 ( .A(n12969), .ZN(n12967) );
  XNOR2_X1 U12930 ( .A(n12970), .B(n12971), .ZN(n12943) );
  XOR2_X1 U12931 ( .A(n12972), .B(n12973), .Z(n12971) );
  NAND2_X1 U12932 ( .A1(b_15_), .A2(a_3_), .ZN(n12973) );
  NAND2_X1 U12933 ( .A1(a_2_), .A2(n12969), .ZN(n12944) );
  NAND2_X1 U12934 ( .A1(n12940), .A2(n12974), .ZN(n12969) );
  NAND2_X1 U12935 ( .A1(n12939), .A2(n12941), .ZN(n12974) );
  NAND2_X1 U12936 ( .A1(n12975), .A2(n12976), .ZN(n12941) );
  NAND2_X1 U12937 ( .A1(b_16_), .A2(a_3_), .ZN(n12976) );
  INV_X1 U12938 ( .A(n12977), .ZN(n12975) );
  XOR2_X1 U12939 ( .A(n12978), .B(n12979), .Z(n12939) );
  XNOR2_X1 U12940 ( .A(n12980), .B(n12981), .ZN(n12979) );
  NAND2_X1 U12941 ( .A1(b_15_), .A2(a_4_), .ZN(n12981) );
  NAND2_X1 U12942 ( .A1(a_3_), .A2(n12977), .ZN(n12940) );
  NAND2_X1 U12943 ( .A1(n12982), .A2(n12983), .ZN(n12977) );
  INV_X1 U12944 ( .A(n12984), .ZN(n12983) );
  NOR3_X1 U12945 ( .A1(n8996), .A2(n12985), .A3(n8989), .ZN(n12984) );
  NOR2_X1 U12946 ( .A1(n12935), .A2(n12936), .ZN(n12985) );
  NAND2_X1 U12947 ( .A1(n12935), .A2(n12936), .ZN(n12982) );
  NAND2_X1 U12948 ( .A1(n12986), .A2(n12987), .ZN(n12936) );
  NAND2_X1 U12949 ( .A1(n12933), .A2(n12988), .ZN(n12987) );
  INV_X1 U12950 ( .A(n12989), .ZN(n12988) );
  NOR2_X1 U12951 ( .A1(n12931), .A2(n12932), .ZN(n12989) );
  NOR2_X1 U12952 ( .A1(n8989), .A2(n8848), .ZN(n12933) );
  NAND2_X1 U12953 ( .A1(n12931), .A2(n12932), .ZN(n12986) );
  NAND2_X1 U12954 ( .A1(n12928), .A2(n12990), .ZN(n12932) );
  NAND2_X1 U12955 ( .A1(n12927), .A2(n12929), .ZN(n12990) );
  NAND2_X1 U12956 ( .A1(n12991), .A2(n12992), .ZN(n12929) );
  NAND2_X1 U12957 ( .A1(b_16_), .A2(a_6_), .ZN(n12992) );
  INV_X1 U12958 ( .A(n12993), .ZN(n12991) );
  XOR2_X1 U12959 ( .A(n12994), .B(n12995), .Z(n12927) );
  XOR2_X1 U12960 ( .A(n12996), .B(n12997), .Z(n12994) );
  NOR2_X1 U12961 ( .A1(n8817), .A2(n8690), .ZN(n12997) );
  NAND2_X1 U12962 ( .A1(a_6_), .A2(n12993), .ZN(n12928) );
  NAND2_X1 U12963 ( .A1(n12924), .A2(n12998), .ZN(n12993) );
  NAND2_X1 U12964 ( .A1(n12923), .A2(n12925), .ZN(n12998) );
  NAND2_X1 U12965 ( .A1(n12999), .A2(n13000), .ZN(n12925) );
  NAND2_X1 U12966 ( .A1(b_16_), .A2(a_7_), .ZN(n13000) );
  INV_X1 U12967 ( .A(n13001), .ZN(n12999) );
  XNOR2_X1 U12968 ( .A(n13002), .B(n13003), .ZN(n12923) );
  XOR2_X1 U12969 ( .A(n13004), .B(n13005), .Z(n13003) );
  NAND2_X1 U12970 ( .A1(b_15_), .A2(a_8_), .ZN(n13005) );
  NAND2_X1 U12971 ( .A1(a_7_), .A2(n13001), .ZN(n12924) );
  NAND2_X1 U12972 ( .A1(n12920), .A2(n13006), .ZN(n13001) );
  NAND2_X1 U12973 ( .A1(n12919), .A2(n12921), .ZN(n13006) );
  NAND2_X1 U12974 ( .A1(n13007), .A2(n13008), .ZN(n12921) );
  NAND2_X1 U12975 ( .A1(b_16_), .A2(a_8_), .ZN(n13008) );
  INV_X1 U12976 ( .A(n13009), .ZN(n13007) );
  XOR2_X1 U12977 ( .A(n13010), .B(n13011), .Z(n12919) );
  XOR2_X1 U12978 ( .A(n13012), .B(n13013), .Z(n13010) );
  NOR2_X1 U12979 ( .A1(n8779), .A2(n8690), .ZN(n13013) );
  NAND2_X1 U12980 ( .A1(a_8_), .A2(n13009), .ZN(n12920) );
  NAND2_X1 U12981 ( .A1(n13014), .A2(n13015), .ZN(n13009) );
  INV_X1 U12982 ( .A(n13016), .ZN(n13015) );
  NOR3_X1 U12983 ( .A1(n8779), .A2(n13017), .A3(n8989), .ZN(n13016) );
  NOR2_X1 U12984 ( .A1(n12915), .A2(n12916), .ZN(n13017) );
  NAND2_X1 U12985 ( .A1(n12915), .A2(n12916), .ZN(n13014) );
  NAND2_X1 U12986 ( .A1(n12912), .A2(n13018), .ZN(n12916) );
  NAND2_X1 U12987 ( .A1(n12911), .A2(n12913), .ZN(n13018) );
  NAND2_X1 U12988 ( .A1(n13019), .A2(n13020), .ZN(n12913) );
  NAND2_X1 U12989 ( .A1(b_16_), .A2(a_10_), .ZN(n13020) );
  XNOR2_X1 U12990 ( .A(n13021), .B(n13022), .ZN(n12911) );
  XNOR2_X1 U12991 ( .A(n13023), .B(n13024), .ZN(n13021) );
  NOR2_X1 U12992 ( .A1(n8749), .A2(n8690), .ZN(n13024) );
  INV_X1 U12993 ( .A(n13025), .ZN(n12912) );
  NOR2_X1 U12994 ( .A1(n8769), .A2(n13019), .ZN(n13025) );
  NOR2_X1 U12995 ( .A1(n13026), .A2(n13027), .ZN(n13019) );
  NOR3_X1 U12996 ( .A1(n8749), .A2(n13028), .A3(n8989), .ZN(n13027) );
  NOR2_X1 U12997 ( .A1(n12907), .A2(n13029), .ZN(n13028) );
  INV_X1 U12998 ( .A(n12908), .ZN(n13029) );
  NOR2_X1 U12999 ( .A1(n13030), .A2(n12908), .ZN(n13026) );
  NOR2_X1 U13000 ( .A1(n13031), .A2(n13032), .ZN(n12908) );
  INV_X1 U13001 ( .A(n13033), .ZN(n13032) );
  NAND2_X1 U13002 ( .A1(n12905), .A2(n13034), .ZN(n13033) );
  NAND2_X1 U13003 ( .A1(n12904), .A2(n12903), .ZN(n13034) );
  NOR2_X1 U13004 ( .A1(n8989), .A2(n8739), .ZN(n12905) );
  NOR2_X1 U13005 ( .A1(n12903), .A2(n12904), .ZN(n13031) );
  NOR2_X1 U13006 ( .A1(n13035), .A2(n13036), .ZN(n12904) );
  INV_X1 U13007 ( .A(n13037), .ZN(n13036) );
  NAND2_X1 U13008 ( .A1(n12901), .A2(n13038), .ZN(n13037) );
  NAND2_X1 U13009 ( .A1(n12900), .A2(n12899), .ZN(n13038) );
  NOR2_X1 U13010 ( .A1(n8989), .A2(n8721), .ZN(n12901) );
  NOR2_X1 U13011 ( .A1(n12899), .A2(n12900), .ZN(n13035) );
  NOR2_X1 U13012 ( .A1(n13039), .A2(n13040), .ZN(n12900) );
  NOR3_X1 U13013 ( .A1(n8991), .A2(n13041), .A3(n8989), .ZN(n13040) );
  INV_X1 U13014 ( .A(n13042), .ZN(n13041) );
  NAND2_X1 U13015 ( .A1(n12896), .A2(n12894), .ZN(n13042) );
  NOR2_X1 U13016 ( .A1(n12894), .A2(n12896), .ZN(n13039) );
  NOR2_X1 U13017 ( .A1(n13043), .A2(n13044), .ZN(n12896) );
  INV_X1 U13018 ( .A(n13045), .ZN(n13044) );
  NAND3_X1 U13019 ( .A1(a_15_), .A2(n13046), .A3(b_16_), .ZN(n13045) );
  NAND2_X1 U13020 ( .A1(n12890), .A2(n12892), .ZN(n13046) );
  NOR2_X1 U13021 ( .A1(n12890), .A2(n12892), .ZN(n13043) );
  NAND2_X1 U13022 ( .A1(n13047), .A2(n13048), .ZN(n12892) );
  NAND2_X1 U13023 ( .A1(n12888), .A2(n13049), .ZN(n13048) );
  INV_X1 U13024 ( .A(n13050), .ZN(n13049) );
  NOR2_X1 U13025 ( .A1(n8674), .A2(n12889), .ZN(n13050) );
  XNOR2_X1 U13026 ( .A(n13051), .B(n13052), .ZN(n12888) );
  XNOR2_X1 U13027 ( .A(n13053), .B(n13054), .ZN(n13052) );
  NAND2_X1 U13028 ( .A1(b_15_), .A2(a_17_), .ZN(n13054) );
  NAND2_X1 U13029 ( .A1(n12889), .A2(n8674), .ZN(n13047) );
  NAND2_X1 U13030 ( .A1(b_16_), .A2(a_16_), .ZN(n8674) );
  NOR2_X1 U13031 ( .A1(n13055), .A2(n13056), .ZN(n12889) );
  INV_X1 U13032 ( .A(n13057), .ZN(n13056) );
  NAND3_X1 U13033 ( .A1(a_17_), .A2(n13058), .A3(b_16_), .ZN(n13057) );
  NAND2_X1 U13034 ( .A1(n12777), .A2(n12778), .ZN(n13058) );
  NOR2_X1 U13035 ( .A1(n12777), .A2(n12778), .ZN(n13055) );
  NAND2_X1 U13036 ( .A1(n13059), .A2(n13060), .ZN(n12778) );
  NAND2_X1 U13037 ( .A1(n12784), .A2(n13061), .ZN(n13060) );
  NAND2_X1 U13038 ( .A1(n12787), .A2(n12786), .ZN(n13061) );
  XNOR2_X1 U13039 ( .A(n13062), .B(n13063), .ZN(n12784) );
  XNOR2_X1 U13040 ( .A(n13064), .B(n13065), .ZN(n13063) );
  NAND2_X1 U13041 ( .A1(b_15_), .A2(a_19_), .ZN(n13065) );
  INV_X1 U13042 ( .A(n13066), .ZN(n13059) );
  NOR2_X1 U13043 ( .A1(n12786), .A2(n12787), .ZN(n13066) );
  NOR2_X1 U13044 ( .A1(n8989), .A2(n8988), .ZN(n12787) );
  NAND2_X1 U13045 ( .A1(n13067), .A2(n13068), .ZN(n12786) );
  NAND3_X1 U13046 ( .A1(a_19_), .A2(n13069), .A3(b_16_), .ZN(n13068) );
  NAND2_X1 U13047 ( .A1(n12885), .A2(n12883), .ZN(n13069) );
  INV_X1 U13048 ( .A(n13070), .ZN(n13067) );
  NOR2_X1 U13049 ( .A1(n12883), .A2(n12885), .ZN(n13070) );
  NOR2_X1 U13050 ( .A1(n13071), .A2(n13072), .ZN(n12885) );
  INV_X1 U13051 ( .A(n13073), .ZN(n13072) );
  NAND2_X1 U13052 ( .A1(n12800), .A2(n13074), .ZN(n13073) );
  NAND2_X1 U13053 ( .A1(n12797), .A2(n12799), .ZN(n13074) );
  NOR2_X1 U13054 ( .A1(n8989), .A2(n8986), .ZN(n12800) );
  NOR2_X1 U13055 ( .A1(n12799), .A2(n12797), .ZN(n13071) );
  XOR2_X1 U13056 ( .A(n13075), .B(n13076), .Z(n12797) );
  XNOR2_X1 U13057 ( .A(n13077), .B(n13078), .ZN(n13075) );
  NOR2_X1 U13058 ( .A1(n8601), .A2(n8690), .ZN(n13078) );
  NAND2_X1 U13059 ( .A1(n13079), .A2(n13080), .ZN(n12799) );
  NAND2_X1 U13060 ( .A1(n12805), .A2(n13081), .ZN(n13080) );
  NAND2_X1 U13061 ( .A1(n12807), .A2(n12806), .ZN(n13081) );
  XNOR2_X1 U13062 ( .A(n13082), .B(n13083), .ZN(n12805) );
  XNOR2_X1 U13063 ( .A(n13084), .B(n13085), .ZN(n13083) );
  INV_X1 U13064 ( .A(n13086), .ZN(n13079) );
  NOR2_X1 U13065 ( .A1(n12806), .A2(n12807), .ZN(n13086) );
  NOR2_X1 U13066 ( .A1(n8989), .A2(n8601), .ZN(n12807) );
  NAND2_X1 U13067 ( .A1(n12815), .A2(n13087), .ZN(n12806) );
  NAND2_X1 U13068 ( .A1(n12814), .A2(n12816), .ZN(n13087) );
  NAND2_X1 U13069 ( .A1(n13088), .A2(n13089), .ZN(n12816) );
  NAND2_X1 U13070 ( .A1(b_16_), .A2(a_22_), .ZN(n13089) );
  INV_X1 U13071 ( .A(n13090), .ZN(n13088) );
  XOR2_X1 U13072 ( .A(n13091), .B(n13092), .Z(n12814) );
  XOR2_X1 U13073 ( .A(n13093), .B(n13094), .Z(n13091) );
  NAND2_X1 U13074 ( .A1(a_22_), .A2(n13090), .ZN(n12815) );
  NAND2_X1 U13075 ( .A1(n12881), .A2(n13095), .ZN(n13090) );
  NAND2_X1 U13076 ( .A1(n12880), .A2(n12882), .ZN(n13095) );
  NAND2_X1 U13077 ( .A1(n13096), .A2(n13097), .ZN(n12882) );
  NAND2_X1 U13078 ( .A1(b_16_), .A2(a_23_), .ZN(n13097) );
  INV_X1 U13079 ( .A(n13098), .ZN(n13096) );
  XOR2_X1 U13080 ( .A(n13099), .B(n13100), .Z(n12880) );
  XOR2_X1 U13081 ( .A(n13101), .B(n13102), .Z(n13099) );
  NAND2_X1 U13082 ( .A1(a_23_), .A2(n13098), .ZN(n12881) );
  NAND2_X1 U13083 ( .A1(n13103), .A2(n13104), .ZN(n13098) );
  NAND2_X1 U13084 ( .A1(n12878), .A2(n13105), .ZN(n13104) );
  INV_X1 U13085 ( .A(n13106), .ZN(n13105) );
  NOR2_X1 U13086 ( .A1(n12876), .A2(n12877), .ZN(n13106) );
  NOR2_X1 U13087 ( .A1(n8989), .A2(n8982), .ZN(n12878) );
  NAND2_X1 U13088 ( .A1(n12876), .A2(n12877), .ZN(n13103) );
  NAND2_X1 U13089 ( .A1(n13107), .A2(n13108), .ZN(n12877) );
  NAND2_X1 U13090 ( .A1(n12874), .A2(n13109), .ZN(n13108) );
  NAND2_X1 U13091 ( .A1(n12871), .A2(n12873), .ZN(n13109) );
  NOR2_X1 U13092 ( .A1(n8989), .A2(n8541), .ZN(n12874) );
  INV_X1 U13093 ( .A(n13110), .ZN(n13107) );
  NOR2_X1 U13094 ( .A1(n12873), .A2(n12871), .ZN(n13110) );
  XNOR2_X1 U13095 ( .A(n13111), .B(n13112), .ZN(n12871) );
  XNOR2_X1 U13096 ( .A(n13113), .B(n13114), .ZN(n13112) );
  NAND2_X1 U13097 ( .A1(n13115), .A2(n13116), .ZN(n12873) );
  NAND2_X1 U13098 ( .A1(n12833), .A2(n13117), .ZN(n13116) );
  NAND2_X1 U13099 ( .A1(n12836), .A2(n12835), .ZN(n13117) );
  XNOR2_X1 U13100 ( .A(n13118), .B(n13119), .ZN(n12833) );
  XOR2_X1 U13101 ( .A(n13120), .B(n13121), .Z(n13118) );
  INV_X1 U13102 ( .A(n13122), .ZN(n13115) );
  NOR2_X1 U13103 ( .A1(n12835), .A2(n12836), .ZN(n13122) );
  NOR2_X1 U13104 ( .A1(n8989), .A2(n9893), .ZN(n12836) );
  NAND2_X1 U13105 ( .A1(n13123), .A2(n13124), .ZN(n12835) );
  NAND2_X1 U13106 ( .A1(n12843), .A2(n13125), .ZN(n13124) );
  INV_X1 U13107 ( .A(n13126), .ZN(n13125) );
  NOR2_X1 U13108 ( .A1(n12841), .A2(n12842), .ZN(n13126) );
  NOR2_X1 U13109 ( .A1(n8989), .A2(n8512), .ZN(n12843) );
  NAND2_X1 U13110 ( .A1(n12841), .A2(n12842), .ZN(n13123) );
  NAND2_X1 U13111 ( .A1(n13127), .A2(n13128), .ZN(n12842) );
  NAND2_X1 U13112 ( .A1(n12869), .A2(n13129), .ZN(n13128) );
  INV_X1 U13113 ( .A(n13130), .ZN(n13129) );
  NOR2_X1 U13114 ( .A1(n12870), .A2(n12868), .ZN(n13130) );
  NOR2_X1 U13115 ( .A1(n8989), .A2(n8493), .ZN(n12869) );
  NAND2_X1 U13116 ( .A1(n12868), .A2(n12870), .ZN(n13127) );
  NAND2_X1 U13117 ( .A1(n13131), .A2(n13132), .ZN(n12870) );
  NAND2_X1 U13118 ( .A1(n12864), .A2(n13133), .ZN(n13132) );
  INV_X1 U13119 ( .A(n13134), .ZN(n13133) );
  NOR2_X1 U13120 ( .A1(n12865), .A2(n12866), .ZN(n13134) );
  NOR2_X1 U13121 ( .A1(n8989), .A2(n8473), .ZN(n12864) );
  NAND2_X1 U13122 ( .A1(n12866), .A2(n12865), .ZN(n13131) );
  NAND2_X1 U13123 ( .A1(n13135), .A2(n13136), .ZN(n12865) );
  NAND2_X1 U13124 ( .A1(b_14_), .A2(n13137), .ZN(n13136) );
  NAND2_X1 U13125 ( .A1(n8456), .A2(n13138), .ZN(n13137) );
  NAND2_X1 U13126 ( .A1(a_31_), .A2(n8690), .ZN(n13138) );
  NAND2_X1 U13127 ( .A1(b_15_), .A2(n13139), .ZN(n13135) );
  NAND2_X1 U13128 ( .A1(n8459), .A2(n13140), .ZN(n13139) );
  NAND2_X1 U13129 ( .A1(a_30_), .A2(n8990), .ZN(n13140) );
  NOR3_X1 U13130 ( .A1(n8690), .A2(n8979), .A3(n8989), .ZN(n12866) );
  INV_X1 U13131 ( .A(b_16_), .ZN(n8989) );
  XOR2_X1 U13132 ( .A(n13141), .B(n13142), .Z(n12868) );
  XOR2_X1 U13133 ( .A(n13143), .B(n13144), .Z(n13141) );
  XOR2_X1 U13134 ( .A(n13145), .B(n13146), .Z(n12841) );
  XOR2_X1 U13135 ( .A(n13147), .B(n13148), .Z(n13145) );
  XNOR2_X1 U13136 ( .A(n13149), .B(n13150), .ZN(n12876) );
  XNOR2_X1 U13137 ( .A(n13151), .B(n13152), .ZN(n13150) );
  XOR2_X1 U13138 ( .A(n13153), .B(n13154), .Z(n12883) );
  XNOR2_X1 U13139 ( .A(n13155), .B(n13156), .ZN(n13153) );
  NOR2_X1 U13140 ( .A1(n8986), .A2(n8690), .ZN(n13156) );
  XOR2_X1 U13141 ( .A(n13157), .B(n13158), .Z(n12777) );
  XOR2_X1 U13142 ( .A(n13159), .B(n13160), .Z(n13158) );
  NAND2_X1 U13143 ( .A1(b_15_), .A2(a_18_), .ZN(n13160) );
  XOR2_X1 U13144 ( .A(n13161), .B(n13162), .Z(n12890) );
  XOR2_X1 U13145 ( .A(n13163), .B(n13164), .Z(n13162) );
  XOR2_X1 U13146 ( .A(n13165), .B(n13166), .Z(n12894) );
  XNOR2_X1 U13147 ( .A(n13167), .B(n8687), .ZN(n13165) );
  XOR2_X1 U13148 ( .A(n13168), .B(n13169), .Z(n12899) );
  NAND2_X1 U13149 ( .A1(n13170), .A2(n13171), .ZN(n13168) );
  XOR2_X1 U13150 ( .A(n13172), .B(n13173), .Z(n12903) );
  XOR2_X1 U13151 ( .A(n13174), .B(n13175), .Z(n13173) );
  NAND2_X1 U13152 ( .A1(b_15_), .A2(a_13_), .ZN(n13175) );
  INV_X1 U13153 ( .A(n12907), .ZN(n13030) );
  XNOR2_X1 U13154 ( .A(n13176), .B(n13177), .ZN(n12907) );
  XOR2_X1 U13155 ( .A(n13178), .B(n13179), .Z(n13177) );
  NAND2_X1 U13156 ( .A1(b_15_), .A2(a_12_), .ZN(n13179) );
  XNOR2_X1 U13157 ( .A(n13180), .B(n13181), .ZN(n12915) );
  XOR2_X1 U13158 ( .A(n13182), .B(n13183), .Z(n13181) );
  NAND2_X1 U13159 ( .A1(b_15_), .A2(a_10_), .ZN(n13183) );
  XNOR2_X1 U13160 ( .A(n13184), .B(n13185), .ZN(n12931) );
  XOR2_X1 U13161 ( .A(n13186), .B(n13187), .Z(n13185) );
  NAND2_X1 U13162 ( .A1(b_15_), .A2(a_6_), .ZN(n13187) );
  XNOR2_X1 U13163 ( .A(n13188), .B(n13189), .ZN(n12935) );
  XOR2_X1 U13164 ( .A(n13190), .B(n13191), .Z(n13188) );
  NAND2_X1 U13165 ( .A1(b_15_), .A2(a_5_), .ZN(n13190) );
  INV_X1 U13166 ( .A(n13192), .ZN(n12948) );
  NOR2_X1 U13167 ( .A1(n13193), .A2(n13194), .ZN(n13192) );
  XOR2_X1 U13168 ( .A(n13195), .B(n13196), .Z(n12699) );
  XOR2_X1 U13169 ( .A(n13197), .B(n13198), .Z(n13195) );
  NOR2_X1 U13170 ( .A1(n9471), .A2(n8690), .ZN(n13198) );
  INV_X1 U13171 ( .A(n12949), .ZN(n9160) );
  NAND2_X1 U13172 ( .A1(n13194), .A2(n13193), .ZN(n12949) );
  NAND2_X1 U13173 ( .A1(n13199), .A2(n13200), .ZN(n13193) );
  NAND3_X1 U13174 ( .A1(a_0_), .A2(n13201), .A3(b_15_), .ZN(n13200) );
  NAND2_X1 U13175 ( .A1(n13196), .A2(n13197), .ZN(n13201) );
  INV_X1 U13176 ( .A(n13202), .ZN(n13199) );
  NOR2_X1 U13177 ( .A1(n13197), .A2(n13196), .ZN(n13202) );
  XOR2_X1 U13178 ( .A(n13203), .B(n13204), .Z(n13196) );
  NAND2_X1 U13179 ( .A1(n13205), .A2(n13206), .ZN(n13203) );
  NAND2_X1 U13180 ( .A1(n13207), .A2(n13208), .ZN(n13197) );
  NAND2_X1 U13181 ( .A1(n12954), .A2(n13209), .ZN(n13208) );
  INV_X1 U13182 ( .A(n13210), .ZN(n13209) );
  NOR2_X1 U13183 ( .A1(n12957), .A2(n12956), .ZN(n13210) );
  XOR2_X1 U13184 ( .A(n13211), .B(n13212), .Z(n12954) );
  NAND2_X1 U13185 ( .A1(n13213), .A2(n13214), .ZN(n13211) );
  NAND2_X1 U13186 ( .A1(n12956), .A2(n12957), .ZN(n13207) );
  NAND2_X1 U13187 ( .A1(b_15_), .A2(a_1_), .ZN(n12957) );
  NOR2_X1 U13188 ( .A1(n13215), .A2(n13216), .ZN(n12956) );
  NOR3_X1 U13189 ( .A1(n8998), .A2(n13217), .A3(n8690), .ZN(n13216) );
  NOR2_X1 U13190 ( .A1(n12964), .A2(n12963), .ZN(n13217) );
  INV_X1 U13191 ( .A(n13218), .ZN(n13215) );
  NAND2_X1 U13192 ( .A1(n12963), .A2(n12964), .ZN(n13218) );
  NAND2_X1 U13193 ( .A1(n13219), .A2(n13220), .ZN(n12964) );
  INV_X1 U13194 ( .A(n13221), .ZN(n13220) );
  NOR3_X1 U13195 ( .A1(n8877), .A2(n13222), .A3(n8690), .ZN(n13221) );
  NOR2_X1 U13196 ( .A1(n12972), .A2(n12970), .ZN(n13222) );
  NAND2_X1 U13197 ( .A1(n12970), .A2(n12972), .ZN(n13219) );
  NAND2_X1 U13198 ( .A1(n13223), .A2(n13224), .ZN(n12972) );
  NAND3_X1 U13199 ( .A1(a_4_), .A2(n13225), .A3(b_15_), .ZN(n13224) );
  NAND2_X1 U13200 ( .A1(n12980), .A2(n12978), .ZN(n13225) );
  INV_X1 U13201 ( .A(n13226), .ZN(n13223) );
  NOR2_X1 U13202 ( .A1(n12978), .A2(n12980), .ZN(n13226) );
  NOR2_X1 U13203 ( .A1(n13227), .A2(n13228), .ZN(n12980) );
  INV_X1 U13204 ( .A(n13229), .ZN(n13228) );
  NAND3_X1 U13205 ( .A1(a_5_), .A2(n13230), .A3(b_15_), .ZN(n13229) );
  NAND2_X1 U13206 ( .A1(n13191), .A2(n13189), .ZN(n13230) );
  NOR2_X1 U13207 ( .A1(n13189), .A2(n13191), .ZN(n13227) );
  NOR2_X1 U13208 ( .A1(n13231), .A2(n13232), .ZN(n13191) );
  NOR3_X1 U13209 ( .A1(n8994), .A2(n13233), .A3(n8690), .ZN(n13232) );
  NOR2_X1 U13210 ( .A1(n13186), .A2(n13184), .ZN(n13233) );
  INV_X1 U13211 ( .A(n13234), .ZN(n13231) );
  NAND2_X1 U13212 ( .A1(n13184), .A2(n13186), .ZN(n13234) );
  NAND2_X1 U13213 ( .A1(n13235), .A2(n13236), .ZN(n13186) );
  INV_X1 U13214 ( .A(n13237), .ZN(n13236) );
  NOR3_X1 U13215 ( .A1(n8817), .A2(n13238), .A3(n8690), .ZN(n13237) );
  NOR2_X1 U13216 ( .A1(n12996), .A2(n12995), .ZN(n13238) );
  NAND2_X1 U13217 ( .A1(n12995), .A2(n12996), .ZN(n13235) );
  NAND2_X1 U13218 ( .A1(n13239), .A2(n13240), .ZN(n12996) );
  NAND3_X1 U13219 ( .A1(a_8_), .A2(n13241), .A3(b_15_), .ZN(n13240) );
  INV_X1 U13220 ( .A(n13242), .ZN(n13241) );
  NOR2_X1 U13221 ( .A1(n13004), .A2(n13002), .ZN(n13242) );
  NAND2_X1 U13222 ( .A1(n13002), .A2(n13004), .ZN(n13239) );
  NAND2_X1 U13223 ( .A1(n13243), .A2(n13244), .ZN(n13004) );
  NAND3_X1 U13224 ( .A1(a_9_), .A2(n13245), .A3(b_15_), .ZN(n13244) );
  INV_X1 U13225 ( .A(n13246), .ZN(n13245) );
  NOR2_X1 U13226 ( .A1(n13012), .A2(n13011), .ZN(n13246) );
  NAND2_X1 U13227 ( .A1(n13011), .A2(n13012), .ZN(n13243) );
  NAND2_X1 U13228 ( .A1(n13247), .A2(n13248), .ZN(n13012) );
  NAND3_X1 U13229 ( .A1(a_10_), .A2(n13249), .A3(b_15_), .ZN(n13248) );
  INV_X1 U13230 ( .A(n13250), .ZN(n13249) );
  NOR2_X1 U13231 ( .A1(n13182), .A2(n13180), .ZN(n13250) );
  NAND2_X1 U13232 ( .A1(n13180), .A2(n13182), .ZN(n13247) );
  NAND2_X1 U13233 ( .A1(n13251), .A2(n13252), .ZN(n13182) );
  NAND3_X1 U13234 ( .A1(a_11_), .A2(n13253), .A3(b_15_), .ZN(n13252) );
  NAND2_X1 U13235 ( .A1(n13023), .A2(n13022), .ZN(n13253) );
  INV_X1 U13236 ( .A(n13254), .ZN(n13251) );
  NOR2_X1 U13237 ( .A1(n13022), .A2(n13023), .ZN(n13254) );
  NOR2_X1 U13238 ( .A1(n13255), .A2(n13256), .ZN(n13023) );
  NOR3_X1 U13239 ( .A1(n8739), .A2(n13257), .A3(n8690), .ZN(n13256) );
  NOR2_X1 U13240 ( .A1(n13178), .A2(n13176), .ZN(n13257) );
  INV_X1 U13241 ( .A(n13258), .ZN(n13255) );
  NAND2_X1 U13242 ( .A1(n13176), .A2(n13178), .ZN(n13258) );
  NAND2_X1 U13243 ( .A1(n13259), .A2(n13260), .ZN(n13178) );
  INV_X1 U13244 ( .A(n13261), .ZN(n13260) );
  NOR3_X1 U13245 ( .A1(n8721), .A2(n13262), .A3(n8690), .ZN(n13261) );
  NOR2_X1 U13246 ( .A1(n13174), .A2(n13172), .ZN(n13262) );
  NAND2_X1 U13247 ( .A1(n13172), .A2(n13174), .ZN(n13259) );
  NAND2_X1 U13248 ( .A1(n13170), .A2(n13263), .ZN(n13174) );
  NAND2_X1 U13249 ( .A1(n13169), .A2(n13171), .ZN(n13263) );
  NAND2_X1 U13250 ( .A1(n13264), .A2(n13265), .ZN(n13171) );
  NAND2_X1 U13251 ( .A1(b_15_), .A2(a_14_), .ZN(n13264) );
  XOR2_X1 U13252 ( .A(n13266), .B(n13267), .Z(n13169) );
  XOR2_X1 U13253 ( .A(n13268), .B(n13269), .Z(n13267) );
  INV_X1 U13254 ( .A(n13270), .ZN(n13170) );
  NOR2_X1 U13255 ( .A1(n13265), .A2(n8991), .ZN(n13270) );
  NAND2_X1 U13256 ( .A1(n13271), .A2(n13272), .ZN(n13265) );
  NAND2_X1 U13257 ( .A1(n13166), .A2(n13273), .ZN(n13272) );
  NAND2_X1 U13258 ( .A1(n8687), .A2(n13274), .ZN(n13273) );
  INV_X1 U13259 ( .A(n13167), .ZN(n13274) );
  XOR2_X1 U13260 ( .A(n13275), .B(n13276), .Z(n13166) );
  XNOR2_X1 U13261 ( .A(n13277), .B(n13278), .ZN(n13275) );
  NOR2_X1 U13262 ( .A1(n8680), .A2(n8990), .ZN(n13278) );
  NAND2_X1 U13263 ( .A1(n13167), .A2(n8945), .ZN(n13271) );
  INV_X1 U13264 ( .A(n8687), .ZN(n8945) );
  NOR2_X1 U13265 ( .A1(n8690), .A2(n8692), .ZN(n8687) );
  NOR2_X1 U13266 ( .A1(n13279), .A2(n13280), .ZN(n13167) );
  NOR2_X1 U13267 ( .A1(n13164), .A2(n13281), .ZN(n13280) );
  NOR2_X1 U13268 ( .A1(n13163), .A2(n13161), .ZN(n13281) );
  NAND2_X1 U13269 ( .A1(b_15_), .A2(a_16_), .ZN(n13164) );
  INV_X1 U13270 ( .A(n13282), .ZN(n13279) );
  NAND2_X1 U13271 ( .A1(n13161), .A2(n13163), .ZN(n13282) );
  NAND2_X1 U13272 ( .A1(n13283), .A2(n13284), .ZN(n13163) );
  NAND3_X1 U13273 ( .A1(a_17_), .A2(n13285), .A3(b_15_), .ZN(n13284) );
  NAND2_X1 U13274 ( .A1(n13053), .A2(n13051), .ZN(n13285) );
  INV_X1 U13275 ( .A(n13286), .ZN(n13283) );
  NOR2_X1 U13276 ( .A1(n13051), .A2(n13053), .ZN(n13286) );
  NOR2_X1 U13277 ( .A1(n13287), .A2(n13288), .ZN(n13053) );
  NOR3_X1 U13278 ( .A1(n8988), .A2(n13289), .A3(n8690), .ZN(n13288) );
  NOR2_X1 U13279 ( .A1(n13159), .A2(n13157), .ZN(n13289) );
  INV_X1 U13280 ( .A(n13290), .ZN(n13287) );
  NAND2_X1 U13281 ( .A1(n13157), .A2(n13159), .ZN(n13290) );
  NAND2_X1 U13282 ( .A1(n13291), .A2(n13292), .ZN(n13159) );
  NAND3_X1 U13283 ( .A1(a_19_), .A2(n13293), .A3(b_15_), .ZN(n13292) );
  NAND2_X1 U13284 ( .A1(n13064), .A2(n13062), .ZN(n13293) );
  INV_X1 U13285 ( .A(n13294), .ZN(n13291) );
  NOR2_X1 U13286 ( .A1(n13062), .A2(n13064), .ZN(n13294) );
  NOR2_X1 U13287 ( .A1(n13295), .A2(n13296), .ZN(n13064) );
  INV_X1 U13288 ( .A(n13297), .ZN(n13296) );
  NAND3_X1 U13289 ( .A1(a_20_), .A2(n13298), .A3(b_15_), .ZN(n13297) );
  NAND2_X1 U13290 ( .A1(n13155), .A2(n13154), .ZN(n13298) );
  NOR2_X1 U13291 ( .A1(n13154), .A2(n13155), .ZN(n13295) );
  NOR2_X1 U13292 ( .A1(n13299), .A2(n13300), .ZN(n13155) );
  INV_X1 U13293 ( .A(n13301), .ZN(n13300) );
  NAND3_X1 U13294 ( .A1(a_21_), .A2(n13302), .A3(b_15_), .ZN(n13301) );
  NAND2_X1 U13295 ( .A1(n13077), .A2(n13076), .ZN(n13302) );
  NOR2_X1 U13296 ( .A1(n13076), .A2(n13077), .ZN(n13299) );
  NOR2_X1 U13297 ( .A1(n13303), .A2(n13304), .ZN(n13077) );
  INV_X1 U13298 ( .A(n13305), .ZN(n13304) );
  NAND2_X1 U13299 ( .A1(n13085), .A2(n13306), .ZN(n13305) );
  NAND2_X1 U13300 ( .A1(n13307), .A2(n13082), .ZN(n13306) );
  NOR2_X1 U13301 ( .A1(n8690), .A2(n8984), .ZN(n13085) );
  NOR2_X1 U13302 ( .A1(n13082), .A2(n13307), .ZN(n13303) );
  INV_X1 U13303 ( .A(n13084), .ZN(n13307) );
  NAND2_X1 U13304 ( .A1(n13308), .A2(n13309), .ZN(n13084) );
  NAND2_X1 U13305 ( .A1(n13094), .A2(n13310), .ZN(n13309) );
  INV_X1 U13306 ( .A(n13311), .ZN(n13310) );
  NOR2_X1 U13307 ( .A1(n13093), .A2(n13092), .ZN(n13311) );
  NOR2_X1 U13308 ( .A1(n8690), .A2(n8572), .ZN(n13094) );
  NAND2_X1 U13309 ( .A1(n13092), .A2(n13093), .ZN(n13308) );
  NAND2_X1 U13310 ( .A1(n13312), .A2(n13313), .ZN(n13093) );
  NAND2_X1 U13311 ( .A1(n13102), .A2(n13314), .ZN(n13313) );
  INV_X1 U13312 ( .A(n13315), .ZN(n13314) );
  NOR2_X1 U13313 ( .A1(n13101), .A2(n13100), .ZN(n13315) );
  NOR2_X1 U13314 ( .A1(n8690), .A2(n8982), .ZN(n13102) );
  NAND2_X1 U13315 ( .A1(n13100), .A2(n13101), .ZN(n13312) );
  NAND2_X1 U13316 ( .A1(n13316), .A2(n13317), .ZN(n13101) );
  NAND2_X1 U13317 ( .A1(n13152), .A2(n13318), .ZN(n13317) );
  NAND2_X1 U13318 ( .A1(n13149), .A2(n13151), .ZN(n13318) );
  NOR2_X1 U13319 ( .A1(n8690), .A2(n8541), .ZN(n13152) );
  INV_X1 U13320 ( .A(n13319), .ZN(n13316) );
  NOR2_X1 U13321 ( .A1(n13151), .A2(n13149), .ZN(n13319) );
  XNOR2_X1 U13322 ( .A(n13320), .B(n13321), .ZN(n13149) );
  XNOR2_X1 U13323 ( .A(n13322), .B(n13323), .ZN(n13321) );
  NAND2_X1 U13324 ( .A1(n13324), .A2(n13325), .ZN(n13151) );
  NAND2_X1 U13325 ( .A1(n13111), .A2(n13326), .ZN(n13325) );
  NAND2_X1 U13326 ( .A1(n13114), .A2(n13113), .ZN(n13326) );
  XNOR2_X1 U13327 ( .A(n13327), .B(n13328), .ZN(n13111) );
  XOR2_X1 U13328 ( .A(n13329), .B(n13330), .Z(n13327) );
  INV_X1 U13329 ( .A(n13331), .ZN(n13324) );
  NOR2_X1 U13330 ( .A1(n13113), .A2(n13114), .ZN(n13331) );
  NOR2_X1 U13331 ( .A1(n8690), .A2(n9893), .ZN(n13114) );
  NAND2_X1 U13332 ( .A1(n13332), .A2(n13333), .ZN(n13113) );
  NAND2_X1 U13333 ( .A1(n13121), .A2(n13334), .ZN(n13333) );
  INV_X1 U13334 ( .A(n13335), .ZN(n13334) );
  NOR2_X1 U13335 ( .A1(n13120), .A2(n13119), .ZN(n13335) );
  NOR2_X1 U13336 ( .A1(n8690), .A2(n8512), .ZN(n13121) );
  NAND2_X1 U13337 ( .A1(n13119), .A2(n13120), .ZN(n13332) );
  NAND2_X1 U13338 ( .A1(n13336), .A2(n13337), .ZN(n13120) );
  NAND2_X1 U13339 ( .A1(n13147), .A2(n13338), .ZN(n13337) );
  INV_X1 U13340 ( .A(n13339), .ZN(n13338) );
  NOR2_X1 U13341 ( .A1(n13148), .A2(n13146), .ZN(n13339) );
  NOR2_X1 U13342 ( .A1(n8690), .A2(n8493), .ZN(n13147) );
  NAND2_X1 U13343 ( .A1(n13146), .A2(n13148), .ZN(n13336) );
  NAND2_X1 U13344 ( .A1(n13340), .A2(n13341), .ZN(n13148) );
  NAND2_X1 U13345 ( .A1(n13142), .A2(n13342), .ZN(n13341) );
  INV_X1 U13346 ( .A(n13343), .ZN(n13342) );
  NOR2_X1 U13347 ( .A1(n13143), .A2(n13144), .ZN(n13343) );
  NOR2_X1 U13348 ( .A1(n8690), .A2(n8473), .ZN(n13142) );
  NAND2_X1 U13349 ( .A1(n13144), .A2(n13143), .ZN(n13340) );
  NAND2_X1 U13350 ( .A1(n13344), .A2(n13345), .ZN(n13143) );
  NAND2_X1 U13351 ( .A1(b_13_), .A2(n13346), .ZN(n13345) );
  NAND2_X1 U13352 ( .A1(n8456), .A2(n13347), .ZN(n13346) );
  NAND2_X1 U13353 ( .A1(a_31_), .A2(n8990), .ZN(n13347) );
  NAND2_X1 U13354 ( .A1(b_14_), .A2(n13348), .ZN(n13344) );
  NAND2_X1 U13355 ( .A1(n8459), .A2(n13349), .ZN(n13348) );
  NAND2_X1 U13356 ( .A1(a_30_), .A2(n8719), .ZN(n13349) );
  NOR3_X1 U13357 ( .A1(n8690), .A2(n8979), .A3(n8990), .ZN(n13144) );
  XOR2_X1 U13358 ( .A(n13350), .B(n13351), .Z(n13146) );
  XOR2_X1 U13359 ( .A(n13352), .B(n13353), .Z(n13350) );
  XOR2_X1 U13360 ( .A(n13354), .B(n13355), .Z(n13119) );
  XOR2_X1 U13361 ( .A(n13356), .B(n13357), .Z(n13354) );
  XNOR2_X1 U13362 ( .A(n13358), .B(n13359), .ZN(n13100) );
  XNOR2_X1 U13363 ( .A(n13360), .B(n13361), .ZN(n13359) );
  XOR2_X1 U13364 ( .A(n13362), .B(n13363), .Z(n13092) );
  XOR2_X1 U13365 ( .A(n13364), .B(n13365), .Z(n13362) );
  XNOR2_X1 U13366 ( .A(n13366), .B(n13367), .ZN(n13082) );
  XOR2_X1 U13367 ( .A(n13368), .B(n13369), .Z(n13366) );
  XOR2_X1 U13368 ( .A(n13370), .B(n13371), .Z(n13076) );
  XNOR2_X1 U13369 ( .A(n13372), .B(n13373), .ZN(n13371) );
  XNOR2_X1 U13370 ( .A(n13374), .B(n13375), .ZN(n13154) );
  XOR2_X1 U13371 ( .A(n13376), .B(n13377), .Z(n13374) );
  NOR2_X1 U13372 ( .A1(n8601), .A2(n8990), .ZN(n13377) );
  XOR2_X1 U13373 ( .A(n13378), .B(n13379), .Z(n13062) );
  XNOR2_X1 U13374 ( .A(n13380), .B(n13381), .ZN(n13378) );
  NOR2_X1 U13375 ( .A1(n8986), .A2(n8990), .ZN(n13381) );
  XOR2_X1 U13376 ( .A(n13382), .B(n13383), .Z(n13157) );
  XNOR2_X1 U13377 ( .A(n13384), .B(n13385), .ZN(n13383) );
  NAND2_X1 U13378 ( .A1(b_14_), .A2(a_19_), .ZN(n13385) );
  XOR2_X1 U13379 ( .A(n13386), .B(n13387), .Z(n13051) );
  XOR2_X1 U13380 ( .A(n13388), .B(n13389), .Z(n13387) );
  NAND2_X1 U13381 ( .A1(b_14_), .A2(a_18_), .ZN(n13389) );
  XNOR2_X1 U13382 ( .A(n13390), .B(n13391), .ZN(n13161) );
  XOR2_X1 U13383 ( .A(n13392), .B(n13393), .Z(n13391) );
  NAND2_X1 U13384 ( .A1(b_14_), .A2(a_17_), .ZN(n13393) );
  XNOR2_X1 U13385 ( .A(n13394), .B(n13395), .ZN(n13172) );
  XOR2_X1 U13386 ( .A(n13396), .B(n8704), .Z(n13394) );
  XNOR2_X1 U13387 ( .A(n13397), .B(n13398), .ZN(n13176) );
  XNOR2_X1 U13388 ( .A(n13399), .B(n13400), .ZN(n13398) );
  XOR2_X1 U13389 ( .A(n13401), .B(n13402), .Z(n13022) );
  XOR2_X1 U13390 ( .A(n13403), .B(n13404), .Z(n13401) );
  XOR2_X1 U13391 ( .A(n13405), .B(n13406), .Z(n13180) );
  XOR2_X1 U13392 ( .A(n13407), .B(n13408), .Z(n13406) );
  XNOR2_X1 U13393 ( .A(n13409), .B(n13410), .ZN(n13011) );
  XOR2_X1 U13394 ( .A(n13411), .B(n13412), .Z(n13409) );
  XOR2_X1 U13395 ( .A(n13413), .B(n13414), .Z(n13002) );
  XOR2_X1 U13396 ( .A(n13415), .B(n13416), .Z(n13413) );
  XNOR2_X1 U13397 ( .A(n13417), .B(n13418), .ZN(n12995) );
  XOR2_X1 U13398 ( .A(n13419), .B(n13420), .Z(n13417) );
  XOR2_X1 U13399 ( .A(n13421), .B(n13422), .Z(n13184) );
  XOR2_X1 U13400 ( .A(n13423), .B(n13424), .Z(n13421) );
  NOR2_X1 U13401 ( .A1(n8817), .A2(n8990), .ZN(n13424) );
  XOR2_X1 U13402 ( .A(n13425), .B(n13426), .Z(n13189) );
  NAND2_X1 U13403 ( .A1(n13427), .A2(n13428), .ZN(n13425) );
  XOR2_X1 U13404 ( .A(n13429), .B(n13430), .Z(n12978) );
  XOR2_X1 U13405 ( .A(n13431), .B(n13432), .Z(n13430) );
  NAND2_X1 U13406 ( .A1(b_14_), .A2(a_5_), .ZN(n13432) );
  XNOR2_X1 U13407 ( .A(n13433), .B(n13434), .ZN(n12970) );
  NAND2_X1 U13408 ( .A1(n13435), .A2(n13436), .ZN(n13433) );
  XNOR2_X1 U13409 ( .A(n13437), .B(n13438), .ZN(n12963) );
  NAND2_X1 U13410 ( .A1(n13439), .A2(n13440), .ZN(n13437) );
  XNOR2_X1 U13411 ( .A(n13441), .B(n13442), .ZN(n13194) );
  NAND2_X1 U13412 ( .A1(n13443), .A2(n13444), .ZN(n13441) );
  XNOR2_X1 U13413 ( .A(n9113), .B(n9114), .ZN(n9104) );
  NAND3_X1 U13414 ( .A1(n9113), .A2(n9114), .A3(n9159), .ZN(n9109) );
  INV_X1 U13415 ( .A(n9112), .ZN(n9159) );
  NAND2_X1 U13416 ( .A1(n13445), .A2(n13446), .ZN(n9112) );
  INV_X1 U13417 ( .A(n9156), .ZN(n13446) );
  NAND2_X1 U13418 ( .A1(n13447), .A2(n13448), .ZN(n13445) );
  NAND2_X1 U13419 ( .A1(n13443), .A2(n13449), .ZN(n9114) );
  NAND2_X1 U13420 ( .A1(n13442), .A2(n13444), .ZN(n13449) );
  NAND2_X1 U13421 ( .A1(n13450), .A2(n13451), .ZN(n13444) );
  NAND2_X1 U13422 ( .A1(b_14_), .A2(a_0_), .ZN(n13451) );
  INV_X1 U13423 ( .A(n13452), .ZN(n13450) );
  XNOR2_X1 U13424 ( .A(n13453), .B(n13454), .ZN(n13442) );
  XOR2_X1 U13425 ( .A(n13455), .B(n13456), .Z(n13454) );
  NAND2_X1 U13426 ( .A1(b_13_), .A2(a_1_), .ZN(n13456) );
  NAND2_X1 U13427 ( .A1(a_0_), .A2(n13452), .ZN(n13443) );
  NAND2_X1 U13428 ( .A1(n13205), .A2(n13457), .ZN(n13452) );
  NAND2_X1 U13429 ( .A1(n13204), .A2(n13206), .ZN(n13457) );
  NAND2_X1 U13430 ( .A1(n13458), .A2(n13459), .ZN(n13206) );
  NAND2_X1 U13431 ( .A1(b_14_), .A2(a_1_), .ZN(n13459) );
  INV_X1 U13432 ( .A(n13460), .ZN(n13458) );
  XOR2_X1 U13433 ( .A(n13461), .B(n13462), .Z(n13204) );
  XOR2_X1 U13434 ( .A(n13463), .B(n13464), .Z(n13461) );
  NOR2_X1 U13435 ( .A1(n8998), .A2(n8719), .ZN(n13464) );
  NAND2_X1 U13436 ( .A1(a_1_), .A2(n13460), .ZN(n13205) );
  NAND2_X1 U13437 ( .A1(n13213), .A2(n13465), .ZN(n13460) );
  NAND2_X1 U13438 ( .A1(n13212), .A2(n13214), .ZN(n13465) );
  NAND2_X1 U13439 ( .A1(n13466), .A2(n13467), .ZN(n13214) );
  NAND2_X1 U13440 ( .A1(b_14_), .A2(a_2_), .ZN(n13467) );
  INV_X1 U13441 ( .A(n13468), .ZN(n13466) );
  XOR2_X1 U13442 ( .A(n13469), .B(n13470), .Z(n13212) );
  XNOR2_X1 U13443 ( .A(n13471), .B(n13472), .ZN(n13470) );
  NAND2_X1 U13444 ( .A1(b_13_), .A2(a_3_), .ZN(n13472) );
  NAND2_X1 U13445 ( .A1(a_2_), .A2(n13468), .ZN(n13213) );
  NAND2_X1 U13446 ( .A1(n13439), .A2(n13473), .ZN(n13468) );
  NAND2_X1 U13447 ( .A1(n13438), .A2(n13440), .ZN(n13473) );
  NAND2_X1 U13448 ( .A1(n13474), .A2(n13475), .ZN(n13440) );
  NAND2_X1 U13449 ( .A1(b_14_), .A2(a_3_), .ZN(n13475) );
  INV_X1 U13450 ( .A(n13476), .ZN(n13474) );
  XNOR2_X1 U13451 ( .A(n13477), .B(n13478), .ZN(n13438) );
  XNOR2_X1 U13452 ( .A(n13479), .B(n13480), .ZN(n13477) );
  NOR2_X1 U13453 ( .A1(n8996), .A2(n8719), .ZN(n13480) );
  NAND2_X1 U13454 ( .A1(a_3_), .A2(n13476), .ZN(n13439) );
  NAND2_X1 U13455 ( .A1(n13435), .A2(n13481), .ZN(n13476) );
  NAND2_X1 U13456 ( .A1(n13434), .A2(n13436), .ZN(n13481) );
  NAND2_X1 U13457 ( .A1(n13482), .A2(n13483), .ZN(n13436) );
  NAND2_X1 U13458 ( .A1(b_14_), .A2(a_4_), .ZN(n13483) );
  XOR2_X1 U13459 ( .A(n13484), .B(n13485), .Z(n13434) );
  XOR2_X1 U13460 ( .A(n13486), .B(n13487), .Z(n13484) );
  NOR2_X1 U13461 ( .A1(n8848), .A2(n8719), .ZN(n13487) );
  INV_X1 U13462 ( .A(n13488), .ZN(n13435) );
  NOR2_X1 U13463 ( .A1(n8996), .A2(n13482), .ZN(n13488) );
  NOR2_X1 U13464 ( .A1(n13489), .A2(n13490), .ZN(n13482) );
  NOR3_X1 U13465 ( .A1(n8848), .A2(n13491), .A3(n8990), .ZN(n13490) );
  NOR2_X1 U13466 ( .A1(n13431), .A2(n13429), .ZN(n13491) );
  INV_X1 U13467 ( .A(n13492), .ZN(n13489) );
  NAND2_X1 U13468 ( .A1(n13429), .A2(n13431), .ZN(n13492) );
  NAND2_X1 U13469 ( .A1(n13427), .A2(n13493), .ZN(n13431) );
  NAND2_X1 U13470 ( .A1(n13426), .A2(n13428), .ZN(n13493) );
  NAND2_X1 U13471 ( .A1(n13494), .A2(n13495), .ZN(n13428) );
  NAND2_X1 U13472 ( .A1(b_14_), .A2(a_6_), .ZN(n13495) );
  XOR2_X1 U13473 ( .A(n13496), .B(n13497), .Z(n13426) );
  XOR2_X1 U13474 ( .A(n13498), .B(n13499), .Z(n13496) );
  NOR2_X1 U13475 ( .A1(n8817), .A2(n8719), .ZN(n13499) );
  NAND2_X1 U13476 ( .A1(a_6_), .A2(n13500), .ZN(n13427) );
  INV_X1 U13477 ( .A(n13494), .ZN(n13500) );
  NOR2_X1 U13478 ( .A1(n13501), .A2(n13502), .ZN(n13494) );
  NOR3_X1 U13479 ( .A1(n8817), .A2(n13503), .A3(n8990), .ZN(n13502) );
  INV_X1 U13480 ( .A(n13504), .ZN(n13503) );
  NAND2_X1 U13481 ( .A1(n13422), .A2(n13423), .ZN(n13504) );
  NOR2_X1 U13482 ( .A1(n13422), .A2(n13423), .ZN(n13501) );
  NAND2_X1 U13483 ( .A1(n13505), .A2(n13506), .ZN(n13423) );
  NAND2_X1 U13484 ( .A1(n13418), .A2(n13507), .ZN(n13506) );
  NAND2_X1 U13485 ( .A1(n13420), .A2(n13419), .ZN(n13507) );
  XNOR2_X1 U13486 ( .A(n13508), .B(n13509), .ZN(n13418) );
  XOR2_X1 U13487 ( .A(n13510), .B(n13511), .Z(n13508) );
  NOR2_X1 U13488 ( .A1(n8779), .A2(n8719), .ZN(n13511) );
  INV_X1 U13489 ( .A(n13512), .ZN(n13505) );
  NOR2_X1 U13490 ( .A1(n13419), .A2(n13420), .ZN(n13512) );
  NOR2_X1 U13491 ( .A1(n8990), .A2(n10513), .ZN(n13420) );
  NAND2_X1 U13492 ( .A1(n13513), .A2(n13514), .ZN(n13419) );
  NAND2_X1 U13493 ( .A1(n13416), .A2(n13515), .ZN(n13514) );
  NAND2_X1 U13494 ( .A1(n13414), .A2(n13415), .ZN(n13515) );
  NOR2_X1 U13495 ( .A1(n8990), .A2(n8779), .ZN(n13416) );
  INV_X1 U13496 ( .A(n13516), .ZN(n13513) );
  NOR2_X1 U13497 ( .A1(n13414), .A2(n13415), .ZN(n13516) );
  NAND2_X1 U13498 ( .A1(n13517), .A2(n13518), .ZN(n13415) );
  NAND2_X1 U13499 ( .A1(n13410), .A2(n13519), .ZN(n13518) );
  NAND2_X1 U13500 ( .A1(n13412), .A2(n13411), .ZN(n13519) );
  XOR2_X1 U13501 ( .A(n13520), .B(n13521), .Z(n13410) );
  XNOR2_X1 U13502 ( .A(n13522), .B(n13523), .ZN(n13520) );
  NOR2_X1 U13503 ( .A1(n8749), .A2(n8719), .ZN(n13523) );
  INV_X1 U13504 ( .A(n13524), .ZN(n13517) );
  NOR2_X1 U13505 ( .A1(n13411), .A2(n13412), .ZN(n13524) );
  NOR2_X1 U13506 ( .A1(n8990), .A2(n8769), .ZN(n13412) );
  NAND2_X1 U13507 ( .A1(n13525), .A2(n13526), .ZN(n13411) );
  NAND2_X1 U13508 ( .A1(n13408), .A2(n13527), .ZN(n13526) );
  INV_X1 U13509 ( .A(n13528), .ZN(n13527) );
  NOR2_X1 U13510 ( .A1(n13405), .A2(n13407), .ZN(n13528) );
  NOR2_X1 U13511 ( .A1(n8990), .A2(n8749), .ZN(n13408) );
  NAND2_X1 U13512 ( .A1(n13405), .A2(n13407), .ZN(n13525) );
  NOR2_X1 U13513 ( .A1(n13529), .A2(n13530), .ZN(n13407) );
  INV_X1 U13514 ( .A(n13531), .ZN(n13530) );
  NAND2_X1 U13515 ( .A1(n13402), .A2(n13532), .ZN(n13531) );
  NAND2_X1 U13516 ( .A1(n13404), .A2(n13403), .ZN(n13532) );
  XOR2_X1 U13517 ( .A(n13533), .B(n13534), .Z(n13402) );
  XNOR2_X1 U13518 ( .A(n13535), .B(n8716), .ZN(n13533) );
  NOR2_X1 U13519 ( .A1(n13403), .A2(n13404), .ZN(n13529) );
  NOR2_X1 U13520 ( .A1(n8990), .A2(n8739), .ZN(n13404) );
  NAND2_X1 U13521 ( .A1(n13536), .A2(n13537), .ZN(n13403) );
  NAND2_X1 U13522 ( .A1(n13400), .A2(n13538), .ZN(n13537) );
  NAND2_X1 U13523 ( .A1(n13397), .A2(n13399), .ZN(n13538) );
  NOR2_X1 U13524 ( .A1(n8990), .A2(n8721), .ZN(n13400) );
  INV_X1 U13525 ( .A(n13539), .ZN(n13536) );
  NOR2_X1 U13526 ( .A1(n13397), .A2(n13399), .ZN(n13539) );
  NAND2_X1 U13527 ( .A1(n13540), .A2(n13541), .ZN(n13399) );
  NAND2_X1 U13528 ( .A1(n13395), .A2(n13542), .ZN(n13541) );
  INV_X1 U13529 ( .A(n13543), .ZN(n13542) );
  NOR2_X1 U13530 ( .A1(n8704), .A2(n13396), .ZN(n13543) );
  XNOR2_X1 U13531 ( .A(n13544), .B(n13545), .ZN(n13395) );
  XNOR2_X1 U13532 ( .A(n13546), .B(n13547), .ZN(n13545) );
  NAND2_X1 U13533 ( .A1(b_13_), .A2(a_15_), .ZN(n13547) );
  NAND2_X1 U13534 ( .A1(n13396), .A2(n8704), .ZN(n13540) );
  NAND2_X1 U13535 ( .A1(b_14_), .A2(a_14_), .ZN(n8704) );
  NOR2_X1 U13536 ( .A1(n13548), .A2(n13549), .ZN(n13396) );
  INV_X1 U13537 ( .A(n13550), .ZN(n13549) );
  NAND2_X1 U13538 ( .A1(n13269), .A2(n13551), .ZN(n13550) );
  NAND2_X1 U13539 ( .A1(n13266), .A2(n13268), .ZN(n13551) );
  NOR2_X1 U13540 ( .A1(n8990), .A2(n8692), .ZN(n13269) );
  NOR2_X1 U13541 ( .A1(n13266), .A2(n13268), .ZN(n13548) );
  NOR2_X1 U13542 ( .A1(n13552), .A2(n13553), .ZN(n13268) );
  NOR3_X1 U13543 ( .A1(n8680), .A2(n13554), .A3(n8990), .ZN(n13553) );
  INV_X1 U13544 ( .A(n13555), .ZN(n13554) );
  NAND2_X1 U13545 ( .A1(n13277), .A2(n13276), .ZN(n13555) );
  NOR2_X1 U13546 ( .A1(n13276), .A2(n13277), .ZN(n13552) );
  NOR2_X1 U13547 ( .A1(n13556), .A2(n13557), .ZN(n13277) );
  NOR3_X1 U13548 ( .A1(n8662), .A2(n13558), .A3(n8990), .ZN(n13557) );
  NOR2_X1 U13549 ( .A1(n13392), .A2(n13390), .ZN(n13558) );
  INV_X1 U13550 ( .A(n13559), .ZN(n13556) );
  NAND2_X1 U13551 ( .A1(n13390), .A2(n13392), .ZN(n13559) );
  NAND2_X1 U13552 ( .A1(n13560), .A2(n13561), .ZN(n13392) );
  INV_X1 U13553 ( .A(n13562), .ZN(n13561) );
  NOR3_X1 U13554 ( .A1(n8988), .A2(n13563), .A3(n8990), .ZN(n13562) );
  NOR2_X1 U13555 ( .A1(n13386), .A2(n13388), .ZN(n13563) );
  NAND2_X1 U13556 ( .A1(n13386), .A2(n13388), .ZN(n13560) );
  NAND2_X1 U13557 ( .A1(n13564), .A2(n13565), .ZN(n13388) );
  NAND3_X1 U13558 ( .A1(a_19_), .A2(n13566), .A3(b_14_), .ZN(n13565) );
  NAND2_X1 U13559 ( .A1(n13384), .A2(n13382), .ZN(n13566) );
  INV_X1 U13560 ( .A(n13567), .ZN(n13564) );
  NOR2_X1 U13561 ( .A1(n13382), .A2(n13384), .ZN(n13567) );
  NOR2_X1 U13562 ( .A1(n13568), .A2(n13569), .ZN(n13384) );
  INV_X1 U13563 ( .A(n13570), .ZN(n13569) );
  NAND3_X1 U13564 ( .A1(a_20_), .A2(n13571), .A3(b_14_), .ZN(n13570) );
  NAND2_X1 U13565 ( .A1(n13379), .A2(n13380), .ZN(n13571) );
  NOR2_X1 U13566 ( .A1(n13379), .A2(n13380), .ZN(n13568) );
  NOR2_X1 U13567 ( .A1(n13572), .A2(n13573), .ZN(n13380) );
  NOR3_X1 U13568 ( .A1(n8601), .A2(n13574), .A3(n8990), .ZN(n13573) );
  NOR2_X1 U13569 ( .A1(n13376), .A2(n13375), .ZN(n13574) );
  INV_X1 U13570 ( .A(n13575), .ZN(n13572) );
  NAND2_X1 U13571 ( .A1(n13375), .A2(n13376), .ZN(n13575) );
  NAND2_X1 U13572 ( .A1(n13576), .A2(n13577), .ZN(n13376) );
  NAND2_X1 U13573 ( .A1(n13373), .A2(n13578), .ZN(n13577) );
  INV_X1 U13574 ( .A(n13579), .ZN(n13578) );
  NOR2_X1 U13575 ( .A1(n13370), .A2(n13372), .ZN(n13579) );
  NOR2_X1 U13576 ( .A1(n8990), .A2(n8984), .ZN(n13373) );
  NAND2_X1 U13577 ( .A1(n13370), .A2(n13372), .ZN(n13576) );
  NAND2_X1 U13578 ( .A1(n13580), .A2(n13581), .ZN(n13372) );
  NAND2_X1 U13579 ( .A1(n13369), .A2(n13582), .ZN(n13581) );
  INV_X1 U13580 ( .A(n13583), .ZN(n13582) );
  NOR2_X1 U13581 ( .A1(n13368), .A2(n13367), .ZN(n13583) );
  NOR2_X1 U13582 ( .A1(n8990), .A2(n8572), .ZN(n13369) );
  NAND2_X1 U13583 ( .A1(n13367), .A2(n13368), .ZN(n13580) );
  NAND2_X1 U13584 ( .A1(n13584), .A2(n13585), .ZN(n13368) );
  NAND2_X1 U13585 ( .A1(n13365), .A2(n13586), .ZN(n13585) );
  INV_X1 U13586 ( .A(n13587), .ZN(n13586) );
  NOR2_X1 U13587 ( .A1(n13363), .A2(n13364), .ZN(n13587) );
  NOR2_X1 U13588 ( .A1(n8990), .A2(n8982), .ZN(n13365) );
  NAND2_X1 U13589 ( .A1(n13363), .A2(n13364), .ZN(n13584) );
  NAND2_X1 U13590 ( .A1(n13588), .A2(n13589), .ZN(n13364) );
  NAND2_X1 U13591 ( .A1(n13361), .A2(n13590), .ZN(n13589) );
  NAND2_X1 U13592 ( .A1(n13358), .A2(n13360), .ZN(n13590) );
  NOR2_X1 U13593 ( .A1(n8990), .A2(n8541), .ZN(n13361) );
  INV_X1 U13594 ( .A(n13591), .ZN(n13588) );
  NOR2_X1 U13595 ( .A1(n13360), .A2(n13358), .ZN(n13591) );
  XNOR2_X1 U13596 ( .A(n13592), .B(n13593), .ZN(n13358) );
  XNOR2_X1 U13597 ( .A(n13594), .B(n13595), .ZN(n13593) );
  NAND2_X1 U13598 ( .A1(n13596), .A2(n13597), .ZN(n13360) );
  NAND2_X1 U13599 ( .A1(n13320), .A2(n13598), .ZN(n13597) );
  NAND2_X1 U13600 ( .A1(n13323), .A2(n13322), .ZN(n13598) );
  XNOR2_X1 U13601 ( .A(n13599), .B(n13600), .ZN(n13320) );
  XOR2_X1 U13602 ( .A(n13601), .B(n13602), .Z(n13599) );
  INV_X1 U13603 ( .A(n13603), .ZN(n13596) );
  NOR2_X1 U13604 ( .A1(n13322), .A2(n13323), .ZN(n13603) );
  NOR2_X1 U13605 ( .A1(n8990), .A2(n9893), .ZN(n13323) );
  NAND2_X1 U13606 ( .A1(n13604), .A2(n13605), .ZN(n13322) );
  NAND2_X1 U13607 ( .A1(n13330), .A2(n13606), .ZN(n13605) );
  INV_X1 U13608 ( .A(n13607), .ZN(n13606) );
  NOR2_X1 U13609 ( .A1(n13328), .A2(n13329), .ZN(n13607) );
  NOR2_X1 U13610 ( .A1(n8990), .A2(n8512), .ZN(n13330) );
  NAND2_X1 U13611 ( .A1(n13328), .A2(n13329), .ZN(n13604) );
  NAND2_X1 U13612 ( .A1(n13608), .A2(n13609), .ZN(n13329) );
  NAND2_X1 U13613 ( .A1(n13356), .A2(n13610), .ZN(n13609) );
  INV_X1 U13614 ( .A(n13611), .ZN(n13610) );
  NOR2_X1 U13615 ( .A1(n13357), .A2(n13355), .ZN(n13611) );
  NOR2_X1 U13616 ( .A1(n8990), .A2(n8493), .ZN(n13356) );
  NAND2_X1 U13617 ( .A1(n13355), .A2(n13357), .ZN(n13608) );
  NAND2_X1 U13618 ( .A1(n13612), .A2(n13613), .ZN(n13357) );
  NAND2_X1 U13619 ( .A1(n13351), .A2(n13614), .ZN(n13613) );
  INV_X1 U13620 ( .A(n13615), .ZN(n13614) );
  NOR2_X1 U13621 ( .A1(n13352), .A2(n13353), .ZN(n13615) );
  NOR2_X1 U13622 ( .A1(n8990), .A2(n8473), .ZN(n13351) );
  NAND2_X1 U13623 ( .A1(n13353), .A2(n13352), .ZN(n13612) );
  NAND2_X1 U13624 ( .A1(n13616), .A2(n13617), .ZN(n13352) );
  NAND2_X1 U13625 ( .A1(b_12_), .A2(n13618), .ZN(n13617) );
  NAND2_X1 U13626 ( .A1(n8456), .A2(n13619), .ZN(n13618) );
  NAND2_X1 U13627 ( .A1(a_31_), .A2(n8719), .ZN(n13619) );
  NAND2_X1 U13628 ( .A1(b_13_), .A2(n13620), .ZN(n13616) );
  NAND2_X1 U13629 ( .A1(n8459), .A2(n13621), .ZN(n13620) );
  NAND2_X1 U13630 ( .A1(a_30_), .A2(n13622), .ZN(n13621) );
  NOR3_X1 U13631 ( .A1(n8719), .A2(n8979), .A3(n8990), .ZN(n13353) );
  XOR2_X1 U13632 ( .A(n13623), .B(n13624), .Z(n13355) );
  XOR2_X1 U13633 ( .A(n13625), .B(n13626), .Z(n13623) );
  XOR2_X1 U13634 ( .A(n13627), .B(n13628), .Z(n13328) );
  XOR2_X1 U13635 ( .A(n13629), .B(n13630), .Z(n13627) );
  XNOR2_X1 U13636 ( .A(n13631), .B(n13632), .ZN(n13363) );
  XNOR2_X1 U13637 ( .A(n13633), .B(n13634), .ZN(n13632) );
  XOR2_X1 U13638 ( .A(n13635), .B(n13636), .Z(n13367) );
  XOR2_X1 U13639 ( .A(n13637), .B(n13638), .Z(n13635) );
  XOR2_X1 U13640 ( .A(n13639), .B(n13640), .Z(n13370) );
  XOR2_X1 U13641 ( .A(n13641), .B(n13642), .Z(n13639) );
  XNOR2_X1 U13642 ( .A(n13643), .B(n13644), .ZN(n13375) );
  XNOR2_X1 U13643 ( .A(n13645), .B(n13646), .ZN(n13644) );
  XNOR2_X1 U13644 ( .A(n13647), .B(n13648), .ZN(n13379) );
  XOR2_X1 U13645 ( .A(n13649), .B(n13650), .Z(n13647) );
  NOR2_X1 U13646 ( .A1(n8601), .A2(n8719), .ZN(n13650) );
  XOR2_X1 U13647 ( .A(n13651), .B(n13652), .Z(n13382) );
  XNOR2_X1 U13648 ( .A(n13653), .B(n13654), .ZN(n13651) );
  NOR2_X1 U13649 ( .A1(n8986), .A2(n8719), .ZN(n13654) );
  XOR2_X1 U13650 ( .A(n13655), .B(n13656), .Z(n13386) );
  XNOR2_X1 U13651 ( .A(n13657), .B(n13658), .ZN(n13656) );
  NAND2_X1 U13652 ( .A1(b_13_), .A2(a_19_), .ZN(n13658) );
  XNOR2_X1 U13653 ( .A(n13659), .B(n13660), .ZN(n13390) );
  XOR2_X1 U13654 ( .A(n13661), .B(n13662), .Z(n13660) );
  XNOR2_X1 U13655 ( .A(n13663), .B(n13664), .ZN(n13276) );
  XNOR2_X1 U13656 ( .A(n13665), .B(n13666), .ZN(n13663) );
  XNOR2_X1 U13657 ( .A(n13667), .B(n13668), .ZN(n13266) );
  XOR2_X1 U13658 ( .A(n13669), .B(n13670), .Z(n13667) );
  NOR2_X1 U13659 ( .A1(n8680), .A2(n8719), .ZN(n13670) );
  XOR2_X1 U13660 ( .A(n13671), .B(n13672), .Z(n13397) );
  XOR2_X1 U13661 ( .A(n13673), .B(n13674), .Z(n13672) );
  NAND2_X1 U13662 ( .A1(b_13_), .A2(a_14_), .ZN(n13674) );
  XNOR2_X1 U13663 ( .A(n13675), .B(n13676), .ZN(n13405) );
  XOR2_X1 U13664 ( .A(n13677), .B(n13678), .Z(n13676) );
  NAND2_X1 U13665 ( .A1(b_13_), .A2(a_12_), .ZN(n13678) );
  XNOR2_X1 U13666 ( .A(n13679), .B(n13680), .ZN(n13414) );
  XNOR2_X1 U13667 ( .A(n13681), .B(n13682), .ZN(n13680) );
  NAND2_X1 U13668 ( .A1(b_13_), .A2(a_10_), .ZN(n13682) );
  XOR2_X1 U13669 ( .A(n13683), .B(n13684), .Z(n13422) );
  XOR2_X1 U13670 ( .A(n13685), .B(n13686), .Z(n13684) );
  NAND2_X1 U13671 ( .A1(b_13_), .A2(a_8_), .ZN(n13686) );
  XNOR2_X1 U13672 ( .A(n13687), .B(n13688), .ZN(n13429) );
  XOR2_X1 U13673 ( .A(n13689), .B(n13690), .Z(n13688) );
  NAND2_X1 U13674 ( .A1(b_13_), .A2(a_6_), .ZN(n13690) );
  XOR2_X1 U13675 ( .A(n13691), .B(n13692), .Z(n9113) );
  XOR2_X1 U13676 ( .A(n13693), .B(n13694), .Z(n13691) );
  NOR2_X1 U13677 ( .A1(n9471), .A2(n8719), .ZN(n13694) );
  NOR2_X1 U13678 ( .A1(n13448), .A2(n13447), .ZN(n9156) );
  NOR2_X1 U13679 ( .A1(n13695), .A2(n13696), .ZN(n13447) );
  NOR3_X1 U13680 ( .A1(n9471), .A2(n13697), .A3(n8719), .ZN(n13696) );
  NOR2_X1 U13681 ( .A1(n13693), .A2(n13692), .ZN(n13697) );
  INV_X1 U13682 ( .A(n13698), .ZN(n13695) );
  NAND2_X1 U13683 ( .A1(n13692), .A2(n13693), .ZN(n13698) );
  NAND2_X1 U13684 ( .A1(n13699), .A2(n13700), .ZN(n13693) );
  NAND3_X1 U13685 ( .A1(a_1_), .A2(n13701), .A3(b_13_), .ZN(n13700) );
  INV_X1 U13686 ( .A(n13702), .ZN(n13701) );
  NOR2_X1 U13687 ( .A1(n13455), .A2(n13453), .ZN(n13702) );
  NAND2_X1 U13688 ( .A1(n13453), .A2(n13455), .ZN(n13699) );
  NAND2_X1 U13689 ( .A1(n13703), .A2(n13704), .ZN(n13455) );
  NAND3_X1 U13690 ( .A1(a_2_), .A2(n13705), .A3(b_13_), .ZN(n13704) );
  INV_X1 U13691 ( .A(n13706), .ZN(n13705) );
  NOR2_X1 U13692 ( .A1(n13463), .A2(n13462), .ZN(n13706) );
  NAND2_X1 U13693 ( .A1(n13462), .A2(n13463), .ZN(n13703) );
  NAND2_X1 U13694 ( .A1(n13707), .A2(n13708), .ZN(n13463) );
  NAND3_X1 U13695 ( .A1(a_3_), .A2(n13709), .A3(b_13_), .ZN(n13708) );
  NAND2_X1 U13696 ( .A1(n13471), .A2(n13469), .ZN(n13709) );
  INV_X1 U13697 ( .A(n13710), .ZN(n13707) );
  NOR2_X1 U13698 ( .A1(n13469), .A2(n13471), .ZN(n13710) );
  NOR2_X1 U13699 ( .A1(n13711), .A2(n13712), .ZN(n13471) );
  INV_X1 U13700 ( .A(n13713), .ZN(n13712) );
  NAND3_X1 U13701 ( .A1(a_4_), .A2(n13714), .A3(b_13_), .ZN(n13713) );
  NAND2_X1 U13702 ( .A1(n13479), .A2(n13478), .ZN(n13714) );
  NOR2_X1 U13703 ( .A1(n13478), .A2(n13479), .ZN(n13711) );
  NOR2_X1 U13704 ( .A1(n13715), .A2(n13716), .ZN(n13479) );
  NOR3_X1 U13705 ( .A1(n8848), .A2(n13717), .A3(n8719), .ZN(n13716) );
  NOR2_X1 U13706 ( .A1(n13486), .A2(n13485), .ZN(n13717) );
  INV_X1 U13707 ( .A(n13718), .ZN(n13715) );
  NAND2_X1 U13708 ( .A1(n13485), .A2(n13486), .ZN(n13718) );
  NAND2_X1 U13709 ( .A1(n13719), .A2(n13720), .ZN(n13486) );
  NAND3_X1 U13710 ( .A1(a_6_), .A2(n13721), .A3(b_13_), .ZN(n13720) );
  INV_X1 U13711 ( .A(n13722), .ZN(n13721) );
  NOR2_X1 U13712 ( .A1(n13689), .A2(n13687), .ZN(n13722) );
  NAND2_X1 U13713 ( .A1(n13687), .A2(n13689), .ZN(n13719) );
  NAND2_X1 U13714 ( .A1(n13723), .A2(n13724), .ZN(n13689) );
  NAND3_X1 U13715 ( .A1(a_7_), .A2(n13725), .A3(b_13_), .ZN(n13724) );
  INV_X1 U13716 ( .A(n13726), .ZN(n13725) );
  NOR2_X1 U13717 ( .A1(n13498), .A2(n13497), .ZN(n13726) );
  NAND2_X1 U13718 ( .A1(n13497), .A2(n13498), .ZN(n13723) );
  NAND2_X1 U13719 ( .A1(n13727), .A2(n13728), .ZN(n13498) );
  INV_X1 U13720 ( .A(n13729), .ZN(n13728) );
  NOR3_X1 U13721 ( .A1(n10513), .A2(n13730), .A3(n8719), .ZN(n13729) );
  NOR2_X1 U13722 ( .A1(n13685), .A2(n13683), .ZN(n13730) );
  NAND2_X1 U13723 ( .A1(n13683), .A2(n13685), .ZN(n13727) );
  NAND2_X1 U13724 ( .A1(n13731), .A2(n13732), .ZN(n13685) );
  NAND3_X1 U13725 ( .A1(a_9_), .A2(n13733), .A3(b_13_), .ZN(n13732) );
  INV_X1 U13726 ( .A(n13734), .ZN(n13733) );
  NOR2_X1 U13727 ( .A1(n13510), .A2(n13509), .ZN(n13734) );
  NAND2_X1 U13728 ( .A1(n13509), .A2(n13510), .ZN(n13731) );
  NAND2_X1 U13729 ( .A1(n13735), .A2(n13736), .ZN(n13510) );
  NAND3_X1 U13730 ( .A1(a_10_), .A2(n13737), .A3(b_13_), .ZN(n13736) );
  NAND2_X1 U13731 ( .A1(n13681), .A2(n13679), .ZN(n13737) );
  INV_X1 U13732 ( .A(n13738), .ZN(n13735) );
  NOR2_X1 U13733 ( .A1(n13679), .A2(n13681), .ZN(n13738) );
  NOR2_X1 U13734 ( .A1(n13739), .A2(n13740), .ZN(n13681) );
  INV_X1 U13735 ( .A(n13741), .ZN(n13740) );
  NAND3_X1 U13736 ( .A1(a_11_), .A2(n13742), .A3(b_13_), .ZN(n13741) );
  NAND2_X1 U13737 ( .A1(n13522), .A2(n13521), .ZN(n13742) );
  NOR2_X1 U13738 ( .A1(n13521), .A2(n13522), .ZN(n13739) );
  NOR2_X1 U13739 ( .A1(n13743), .A2(n13744), .ZN(n13522) );
  INV_X1 U13740 ( .A(n13745), .ZN(n13744) );
  NAND3_X1 U13741 ( .A1(a_12_), .A2(n13746), .A3(b_13_), .ZN(n13745) );
  NAND2_X1 U13742 ( .A1(n13675), .A2(n13677), .ZN(n13746) );
  NOR2_X1 U13743 ( .A1(n13677), .A2(n13675), .ZN(n13743) );
  XOR2_X1 U13744 ( .A(n13747), .B(n13748), .Z(n13675) );
  NAND2_X1 U13745 ( .A1(n13749), .A2(n13750), .ZN(n13747) );
  NAND2_X1 U13746 ( .A1(n13751), .A2(n13752), .ZN(n13677) );
  NAND2_X1 U13747 ( .A1(n13534), .A2(n13753), .ZN(n13752) );
  NAND2_X1 U13748 ( .A1(n8716), .A2(n13754), .ZN(n13753) );
  XOR2_X1 U13749 ( .A(n13755), .B(n13756), .Z(n13534) );
  NAND2_X1 U13750 ( .A1(n13757), .A2(n13758), .ZN(n13755) );
  INV_X1 U13751 ( .A(n13759), .ZN(n13751) );
  NOR2_X1 U13752 ( .A1(n13754), .A2(n8716), .ZN(n13759) );
  NOR2_X1 U13753 ( .A1(n8719), .A2(n8721), .ZN(n8716) );
  INV_X1 U13754 ( .A(n13535), .ZN(n13754) );
  NOR2_X1 U13755 ( .A1(n13760), .A2(n13761), .ZN(n13535) );
  NOR3_X1 U13756 ( .A1(n8991), .A2(n13762), .A3(n8719), .ZN(n13761) );
  NOR2_X1 U13757 ( .A1(n13673), .A2(n13671), .ZN(n13762) );
  INV_X1 U13758 ( .A(n13763), .ZN(n13760) );
  NAND2_X1 U13759 ( .A1(n13671), .A2(n13673), .ZN(n13763) );
  NAND2_X1 U13760 ( .A1(n13764), .A2(n13765), .ZN(n13673) );
  NAND3_X1 U13761 ( .A1(a_15_), .A2(n13766), .A3(b_13_), .ZN(n13765) );
  NAND2_X1 U13762 ( .A1(n13546), .A2(n13544), .ZN(n13766) );
  INV_X1 U13763 ( .A(n13767), .ZN(n13764) );
  NOR2_X1 U13764 ( .A1(n13544), .A2(n13546), .ZN(n13767) );
  NOR2_X1 U13765 ( .A1(n13768), .A2(n13769), .ZN(n13546) );
  NOR3_X1 U13766 ( .A1(n8680), .A2(n13770), .A3(n8719), .ZN(n13769) );
  NOR2_X1 U13767 ( .A1(n13669), .A2(n13668), .ZN(n13770) );
  INV_X1 U13768 ( .A(n13771), .ZN(n13768) );
  NAND2_X1 U13769 ( .A1(n13668), .A2(n13669), .ZN(n13771) );
  NAND2_X1 U13770 ( .A1(n13772), .A2(n13773), .ZN(n13669) );
  NAND2_X1 U13771 ( .A1(n13666), .A2(n13774), .ZN(n13773) );
  NAND2_X1 U13772 ( .A1(n13665), .A2(n13775), .ZN(n13774) );
  INV_X1 U13773 ( .A(n13664), .ZN(n13775) );
  NOR2_X1 U13774 ( .A1(n8719), .A2(n8662), .ZN(n13666) );
  NAND2_X1 U13775 ( .A1(n13664), .A2(n13776), .ZN(n13772) );
  INV_X1 U13776 ( .A(n13665), .ZN(n13776) );
  NOR2_X1 U13777 ( .A1(n13777), .A2(n13778), .ZN(n13665) );
  NOR2_X1 U13778 ( .A1(n13662), .A2(n13779), .ZN(n13778) );
  NOR2_X1 U13779 ( .A1(n13661), .A2(n13659), .ZN(n13779) );
  NAND2_X1 U13780 ( .A1(b_13_), .A2(a_18_), .ZN(n13662) );
  INV_X1 U13781 ( .A(n13780), .ZN(n13777) );
  NAND2_X1 U13782 ( .A1(n13659), .A2(n13661), .ZN(n13780) );
  NAND2_X1 U13783 ( .A1(n13781), .A2(n13782), .ZN(n13661) );
  NAND3_X1 U13784 ( .A1(a_19_), .A2(n13783), .A3(b_13_), .ZN(n13782) );
  NAND2_X1 U13785 ( .A1(n13657), .A2(n13655), .ZN(n13783) );
  INV_X1 U13786 ( .A(n13784), .ZN(n13781) );
  NOR2_X1 U13787 ( .A1(n13655), .A2(n13657), .ZN(n13784) );
  NOR2_X1 U13788 ( .A1(n13785), .A2(n13786), .ZN(n13657) );
  INV_X1 U13789 ( .A(n13787), .ZN(n13786) );
  NAND3_X1 U13790 ( .A1(a_20_), .A2(n13788), .A3(b_13_), .ZN(n13787) );
  NAND2_X1 U13791 ( .A1(n13653), .A2(n13652), .ZN(n13788) );
  NOR2_X1 U13792 ( .A1(n13652), .A2(n13653), .ZN(n13785) );
  NOR2_X1 U13793 ( .A1(n13789), .A2(n13790), .ZN(n13653) );
  NOR3_X1 U13794 ( .A1(n8601), .A2(n13791), .A3(n8719), .ZN(n13790) );
  NOR2_X1 U13795 ( .A1(n13649), .A2(n13648), .ZN(n13791) );
  INV_X1 U13796 ( .A(n13792), .ZN(n13789) );
  NAND2_X1 U13797 ( .A1(n13648), .A2(n13649), .ZN(n13792) );
  NAND2_X1 U13798 ( .A1(n13793), .A2(n13794), .ZN(n13649) );
  NAND2_X1 U13799 ( .A1(n13646), .A2(n13795), .ZN(n13794) );
  INV_X1 U13800 ( .A(n13796), .ZN(n13795) );
  NOR2_X1 U13801 ( .A1(n13645), .A2(n13643), .ZN(n13796) );
  NOR2_X1 U13802 ( .A1(n8719), .A2(n8984), .ZN(n13646) );
  NAND2_X1 U13803 ( .A1(n13643), .A2(n13645), .ZN(n13793) );
  NAND2_X1 U13804 ( .A1(n13797), .A2(n13798), .ZN(n13645) );
  NAND2_X1 U13805 ( .A1(n13642), .A2(n13799), .ZN(n13798) );
  INV_X1 U13806 ( .A(n13800), .ZN(n13799) );
  NOR2_X1 U13807 ( .A1(n13641), .A2(n13640), .ZN(n13800) );
  NOR2_X1 U13808 ( .A1(n8719), .A2(n8572), .ZN(n13642) );
  NAND2_X1 U13809 ( .A1(n13640), .A2(n13641), .ZN(n13797) );
  NAND2_X1 U13810 ( .A1(n13801), .A2(n13802), .ZN(n13641) );
  NAND2_X1 U13811 ( .A1(n13638), .A2(n13803), .ZN(n13802) );
  INV_X1 U13812 ( .A(n13804), .ZN(n13803) );
  NOR2_X1 U13813 ( .A1(n13637), .A2(n13636), .ZN(n13804) );
  NOR2_X1 U13814 ( .A1(n8719), .A2(n8982), .ZN(n13638) );
  NAND2_X1 U13815 ( .A1(n13636), .A2(n13637), .ZN(n13801) );
  NAND2_X1 U13816 ( .A1(n13805), .A2(n13806), .ZN(n13637) );
  NAND2_X1 U13817 ( .A1(n13634), .A2(n13807), .ZN(n13806) );
  NAND2_X1 U13818 ( .A1(n13631), .A2(n13633), .ZN(n13807) );
  NOR2_X1 U13819 ( .A1(n8719), .A2(n8541), .ZN(n13634) );
  INV_X1 U13820 ( .A(n13808), .ZN(n13805) );
  NOR2_X1 U13821 ( .A1(n13633), .A2(n13631), .ZN(n13808) );
  XNOR2_X1 U13822 ( .A(n13809), .B(n13810), .ZN(n13631) );
  XNOR2_X1 U13823 ( .A(n13811), .B(n13812), .ZN(n13810) );
  NAND2_X1 U13824 ( .A1(n13813), .A2(n13814), .ZN(n13633) );
  NAND2_X1 U13825 ( .A1(n13592), .A2(n13815), .ZN(n13814) );
  NAND2_X1 U13826 ( .A1(n13595), .A2(n13594), .ZN(n13815) );
  XNOR2_X1 U13827 ( .A(n13816), .B(n13817), .ZN(n13592) );
  XOR2_X1 U13828 ( .A(n13818), .B(n13819), .Z(n13816) );
  INV_X1 U13829 ( .A(n13820), .ZN(n13813) );
  NOR2_X1 U13830 ( .A1(n13594), .A2(n13595), .ZN(n13820) );
  NOR2_X1 U13831 ( .A1(n8719), .A2(n9893), .ZN(n13595) );
  NAND2_X1 U13832 ( .A1(n13821), .A2(n13822), .ZN(n13594) );
  NAND2_X1 U13833 ( .A1(n13602), .A2(n13823), .ZN(n13822) );
  INV_X1 U13834 ( .A(n13824), .ZN(n13823) );
  NOR2_X1 U13835 ( .A1(n13601), .A2(n13600), .ZN(n13824) );
  NOR2_X1 U13836 ( .A1(n8719), .A2(n8512), .ZN(n13602) );
  NAND2_X1 U13837 ( .A1(n13600), .A2(n13601), .ZN(n13821) );
  NAND2_X1 U13838 ( .A1(n13825), .A2(n13826), .ZN(n13601) );
  NAND2_X1 U13839 ( .A1(n13629), .A2(n13827), .ZN(n13826) );
  INV_X1 U13840 ( .A(n13828), .ZN(n13827) );
  NOR2_X1 U13841 ( .A1(n13630), .A2(n13628), .ZN(n13828) );
  NOR2_X1 U13842 ( .A1(n8719), .A2(n8493), .ZN(n13629) );
  NAND2_X1 U13843 ( .A1(n13628), .A2(n13630), .ZN(n13825) );
  NAND2_X1 U13844 ( .A1(n13829), .A2(n13830), .ZN(n13630) );
  NAND2_X1 U13845 ( .A1(n13624), .A2(n13831), .ZN(n13830) );
  INV_X1 U13846 ( .A(n13832), .ZN(n13831) );
  NOR2_X1 U13847 ( .A1(n13625), .A2(n13626), .ZN(n13832) );
  NOR2_X1 U13848 ( .A1(n8719), .A2(n8473), .ZN(n13624) );
  NAND2_X1 U13849 ( .A1(n13626), .A2(n13625), .ZN(n13829) );
  NAND2_X1 U13850 ( .A1(n13833), .A2(n13834), .ZN(n13625) );
  NAND2_X1 U13851 ( .A1(b_11_), .A2(n13835), .ZN(n13834) );
  NAND2_X1 U13852 ( .A1(n8456), .A2(n13836), .ZN(n13835) );
  NAND2_X1 U13853 ( .A1(a_31_), .A2(n13622), .ZN(n13836) );
  NAND2_X1 U13854 ( .A1(b_12_), .A2(n13837), .ZN(n13833) );
  NAND2_X1 U13855 ( .A1(n8459), .A2(n13838), .ZN(n13837) );
  NAND2_X1 U13856 ( .A1(a_30_), .A2(n8751), .ZN(n13838) );
  NOR3_X1 U13857 ( .A1(n8719), .A2(n8979), .A3(n13622), .ZN(n13626) );
  XOR2_X1 U13858 ( .A(n13839), .B(n13840), .Z(n13628) );
  XOR2_X1 U13859 ( .A(n13841), .B(n13842), .Z(n13839) );
  XOR2_X1 U13860 ( .A(n13843), .B(n13844), .Z(n13600) );
  XOR2_X1 U13861 ( .A(n13845), .B(n13846), .Z(n13843) );
  XNOR2_X1 U13862 ( .A(n13847), .B(n13848), .ZN(n13636) );
  XNOR2_X1 U13863 ( .A(n13849), .B(n13850), .ZN(n13848) );
  XOR2_X1 U13864 ( .A(n13851), .B(n13852), .Z(n13640) );
  XOR2_X1 U13865 ( .A(n13853), .B(n13854), .Z(n13851) );
  XOR2_X1 U13866 ( .A(n13855), .B(n13856), .Z(n13643) );
  XOR2_X1 U13867 ( .A(n13857), .B(n13858), .Z(n13855) );
  XNOR2_X1 U13868 ( .A(n13859), .B(n13860), .ZN(n13648) );
  XNOR2_X1 U13869 ( .A(n13861), .B(n13862), .ZN(n13860) );
  XNOR2_X1 U13870 ( .A(n13863), .B(n13864), .ZN(n13652) );
  XOR2_X1 U13871 ( .A(n13865), .B(n13866), .Z(n13863) );
  NOR2_X1 U13872 ( .A1(n8601), .A2(n13622), .ZN(n13866) );
  XOR2_X1 U13873 ( .A(n13867), .B(n13868), .Z(n13655) );
  XNOR2_X1 U13874 ( .A(n13869), .B(n13870), .ZN(n13867) );
  NOR2_X1 U13875 ( .A1(n8986), .A2(n13622), .ZN(n13870) );
  XOR2_X1 U13876 ( .A(n13871), .B(n13872), .Z(n13659) );
  XNOR2_X1 U13877 ( .A(n13873), .B(n13874), .ZN(n13872) );
  NAND2_X1 U13878 ( .A1(b_12_), .A2(a_19_), .ZN(n13874) );
  XOR2_X1 U13879 ( .A(n13875), .B(n13876), .Z(n13664) );
  XNOR2_X1 U13880 ( .A(n13877), .B(n13878), .ZN(n13876) );
  NAND2_X1 U13881 ( .A1(b_12_), .A2(a_18_), .ZN(n13878) );
  XNOR2_X1 U13882 ( .A(n13879), .B(n13880), .ZN(n13668) );
  XNOR2_X1 U13883 ( .A(n13881), .B(n13882), .ZN(n13879) );
  XNOR2_X1 U13884 ( .A(n13883), .B(n13884), .ZN(n13544) );
  XOR2_X1 U13885 ( .A(n13885), .B(n13886), .Z(n13883) );
  XNOR2_X1 U13886 ( .A(n13887), .B(n13888), .ZN(n13671) );
  XOR2_X1 U13887 ( .A(n13889), .B(n13890), .Z(n13888) );
  NAND2_X1 U13888 ( .A1(b_12_), .A2(a_15_), .ZN(n13890) );
  XOR2_X1 U13889 ( .A(n13891), .B(n13892), .Z(n13521) );
  XNOR2_X1 U13890 ( .A(n8733), .B(n13893), .ZN(n13892) );
  XNOR2_X1 U13891 ( .A(n13894), .B(n13895), .ZN(n13679) );
  XNOR2_X1 U13892 ( .A(n13896), .B(n13897), .ZN(n13895) );
  XOR2_X1 U13893 ( .A(n13898), .B(n13899), .Z(n13509) );
  NOR2_X1 U13894 ( .A1(n13900), .A2(n13901), .ZN(n13899) );
  NOR2_X1 U13895 ( .A1(n13902), .A2(n13903), .ZN(n13900) );
  NOR2_X1 U13896 ( .A1(n8769), .A2(n13622), .ZN(n13903) );
  XNOR2_X1 U13897 ( .A(n13904), .B(n13905), .ZN(n13683) );
  NAND2_X1 U13898 ( .A1(n13906), .A2(n13907), .ZN(n13904) );
  XOR2_X1 U13899 ( .A(n13908), .B(n13909), .Z(n13497) );
  NOR2_X1 U13900 ( .A1(n13910), .A2(n13911), .ZN(n13909) );
  NOR2_X1 U13901 ( .A1(n13912), .A2(n13913), .ZN(n13910) );
  NOR2_X1 U13902 ( .A1(n10513), .A2(n13622), .ZN(n13912) );
  XNOR2_X1 U13903 ( .A(n13914), .B(n13915), .ZN(n13687) );
  NAND2_X1 U13904 ( .A1(n13916), .A2(n13917), .ZN(n13914) );
  XNOR2_X1 U13905 ( .A(n13918), .B(n13919), .ZN(n13485) );
  NAND2_X1 U13906 ( .A1(n13920), .A2(n13921), .ZN(n13918) );
  XOR2_X1 U13907 ( .A(n13922), .B(n13923), .Z(n13478) );
  NAND2_X1 U13908 ( .A1(n13924), .A2(n13925), .ZN(n13922) );
  XOR2_X1 U13909 ( .A(n13926), .B(n13927), .Z(n13469) );
  NAND2_X1 U13910 ( .A1(n13928), .A2(n13929), .ZN(n13926) );
  XNOR2_X1 U13911 ( .A(n13930), .B(n13931), .ZN(n13462) );
  NAND2_X1 U13912 ( .A1(n13932), .A2(n13933), .ZN(n13930) );
  XNOR2_X1 U13913 ( .A(n13934), .B(n13935), .ZN(n13453) );
  NAND2_X1 U13914 ( .A1(n13936), .A2(n13937), .ZN(n13934) );
  XNOR2_X1 U13915 ( .A(n13938), .B(n13939), .ZN(n13692) );
  XOR2_X1 U13916 ( .A(n13940), .B(n13941), .Z(n13939) );
  XNOR2_X1 U13917 ( .A(n13942), .B(n13943), .ZN(n13448) );
  XOR2_X1 U13918 ( .A(n13944), .B(n13945), .Z(n13942) );
  NOR2_X1 U13919 ( .A1(n9471), .A2(n13622), .ZN(n13945) );
  XNOR2_X1 U13920 ( .A(n9126), .B(n9125), .ZN(n9116) );
  NAND3_X1 U13921 ( .A1(n9125), .A2(n9126), .A3(n9155), .ZN(n9121) );
  INV_X1 U13922 ( .A(n9124), .ZN(n9155) );
  NAND2_X1 U13923 ( .A1(n13946), .A2(n13947), .ZN(n9124) );
  INV_X1 U13924 ( .A(n9152), .ZN(n13947) );
  NAND2_X1 U13925 ( .A1(n13948), .A2(n13949), .ZN(n13946) );
  NAND2_X1 U13926 ( .A1(n13950), .A2(n13951), .ZN(n9126) );
  INV_X1 U13927 ( .A(n13952), .ZN(n13951) );
  NOR3_X1 U13928 ( .A1(n9471), .A2(n13953), .A3(n13622), .ZN(n13952) );
  NOR2_X1 U13929 ( .A1(n13943), .A2(n13944), .ZN(n13953) );
  NAND2_X1 U13930 ( .A1(n13943), .A2(n13944), .ZN(n13950) );
  NAND2_X1 U13931 ( .A1(n13954), .A2(n13955), .ZN(n13944) );
  INV_X1 U13932 ( .A(n13956), .ZN(n13955) );
  NOR2_X1 U13933 ( .A1(n13941), .A2(n13957), .ZN(n13956) );
  NOR2_X1 U13934 ( .A1(n13938), .A2(n13940), .ZN(n13957) );
  NAND2_X1 U13935 ( .A1(b_12_), .A2(a_1_), .ZN(n13941) );
  NAND2_X1 U13936 ( .A1(n13938), .A2(n13940), .ZN(n13954) );
  NAND2_X1 U13937 ( .A1(n13936), .A2(n13958), .ZN(n13940) );
  NAND2_X1 U13938 ( .A1(n13935), .A2(n13937), .ZN(n13958) );
  NAND2_X1 U13939 ( .A1(n13959), .A2(n13960), .ZN(n13937) );
  NAND2_X1 U13940 ( .A1(b_12_), .A2(a_2_), .ZN(n13960) );
  INV_X1 U13941 ( .A(n13961), .ZN(n13959) );
  XNOR2_X1 U13942 ( .A(n13962), .B(n13963), .ZN(n13935) );
  XOR2_X1 U13943 ( .A(n13964), .B(n13965), .Z(n13963) );
  NAND2_X1 U13944 ( .A1(a_3_), .A2(b_11_), .ZN(n13965) );
  NAND2_X1 U13945 ( .A1(a_2_), .A2(n13961), .ZN(n13936) );
  NAND2_X1 U13946 ( .A1(n13932), .A2(n13966), .ZN(n13961) );
  NAND2_X1 U13947 ( .A1(n13931), .A2(n13933), .ZN(n13966) );
  NAND2_X1 U13948 ( .A1(n13967), .A2(n13968), .ZN(n13933) );
  NAND2_X1 U13949 ( .A1(b_12_), .A2(a_3_), .ZN(n13968) );
  INV_X1 U13950 ( .A(n13969), .ZN(n13967) );
  XOR2_X1 U13951 ( .A(n13970), .B(n13971), .Z(n13931) );
  XNOR2_X1 U13952 ( .A(n13972), .B(n13973), .ZN(n13971) );
  NAND2_X1 U13953 ( .A1(a_4_), .A2(b_11_), .ZN(n13973) );
  NAND2_X1 U13954 ( .A1(a_3_), .A2(n13969), .ZN(n13932) );
  NAND2_X1 U13955 ( .A1(n13928), .A2(n13974), .ZN(n13969) );
  NAND2_X1 U13956 ( .A1(n13927), .A2(n13929), .ZN(n13974) );
  NAND2_X1 U13957 ( .A1(n13975), .A2(n13976), .ZN(n13929) );
  NAND2_X1 U13958 ( .A1(b_12_), .A2(a_4_), .ZN(n13976) );
  INV_X1 U13959 ( .A(n13977), .ZN(n13975) );
  XOR2_X1 U13960 ( .A(n13978), .B(n13979), .Z(n13927) );
  XOR2_X1 U13961 ( .A(n13980), .B(n13981), .Z(n13978) );
  NOR2_X1 U13962 ( .A1(n8751), .A2(n8848), .ZN(n13981) );
  NAND2_X1 U13963 ( .A1(a_4_), .A2(n13977), .ZN(n13928) );
  NAND2_X1 U13964 ( .A1(n13924), .A2(n13982), .ZN(n13977) );
  NAND2_X1 U13965 ( .A1(n13923), .A2(n13925), .ZN(n13982) );
  NAND2_X1 U13966 ( .A1(n13983), .A2(n13984), .ZN(n13925) );
  NAND2_X1 U13967 ( .A1(b_12_), .A2(a_5_), .ZN(n13984) );
  INV_X1 U13968 ( .A(n13985), .ZN(n13983) );
  XNOR2_X1 U13969 ( .A(n13986), .B(n13987), .ZN(n13923) );
  XOR2_X1 U13970 ( .A(n13988), .B(n13989), .Z(n13987) );
  NAND2_X1 U13971 ( .A1(a_6_), .A2(b_11_), .ZN(n13989) );
  NAND2_X1 U13972 ( .A1(a_5_), .A2(n13985), .ZN(n13924) );
  NAND2_X1 U13973 ( .A1(n13920), .A2(n13990), .ZN(n13985) );
  NAND2_X1 U13974 ( .A1(n13919), .A2(n13921), .ZN(n13990) );
  NAND2_X1 U13975 ( .A1(n13991), .A2(n13992), .ZN(n13921) );
  NAND2_X1 U13976 ( .A1(b_12_), .A2(a_6_), .ZN(n13992) );
  INV_X1 U13977 ( .A(n13993), .ZN(n13991) );
  XOR2_X1 U13978 ( .A(n13994), .B(n13995), .Z(n13919) );
  XOR2_X1 U13979 ( .A(n13996), .B(n13997), .Z(n13994) );
  NOR2_X1 U13980 ( .A1(n8751), .A2(n8817), .ZN(n13997) );
  NAND2_X1 U13981 ( .A1(a_6_), .A2(n13993), .ZN(n13920) );
  NAND2_X1 U13982 ( .A1(n13916), .A2(n13998), .ZN(n13993) );
  NAND2_X1 U13983 ( .A1(n13915), .A2(n13917), .ZN(n13998) );
  NAND2_X1 U13984 ( .A1(n13999), .A2(n14000), .ZN(n13917) );
  NAND2_X1 U13985 ( .A1(b_12_), .A2(a_7_), .ZN(n14000) );
  INV_X1 U13986 ( .A(n14001), .ZN(n13999) );
  XOR2_X1 U13987 ( .A(n14002), .B(n14003), .Z(n13915) );
  XNOR2_X1 U13988 ( .A(n14004), .B(n14005), .ZN(n14003) );
  NAND2_X1 U13989 ( .A1(a_8_), .A2(b_11_), .ZN(n14005) );
  NAND2_X1 U13990 ( .A1(a_7_), .A2(n14001), .ZN(n13916) );
  NAND2_X1 U13991 ( .A1(n14006), .A2(n14007), .ZN(n14001) );
  NAND2_X1 U13992 ( .A1(n13908), .A2(n14008), .ZN(n14007) );
  NAND2_X1 U13993 ( .A1(n14009), .A2(n14010), .ZN(n14008) );
  NAND2_X1 U13994 ( .A1(b_12_), .A2(a_8_), .ZN(n14010) );
  XNOR2_X1 U13995 ( .A(n14011), .B(n14012), .ZN(n13908) );
  XNOR2_X1 U13996 ( .A(n14013), .B(n14014), .ZN(n14011) );
  NOR2_X1 U13997 ( .A1(n8751), .A2(n8779), .ZN(n14014) );
  INV_X1 U13998 ( .A(n13911), .ZN(n14006) );
  NOR2_X1 U13999 ( .A1(n10513), .A2(n14009), .ZN(n13911) );
  INV_X1 U14000 ( .A(n13913), .ZN(n14009) );
  NAND2_X1 U14001 ( .A1(n13906), .A2(n14015), .ZN(n13913) );
  NAND2_X1 U14002 ( .A1(n13905), .A2(n13907), .ZN(n14015) );
  NAND2_X1 U14003 ( .A1(n14016), .A2(n14017), .ZN(n13907) );
  NAND2_X1 U14004 ( .A1(b_12_), .A2(a_9_), .ZN(n14017) );
  INV_X1 U14005 ( .A(n14018), .ZN(n14016) );
  XOR2_X1 U14006 ( .A(n14019), .B(n14020), .Z(n13905) );
  XOR2_X1 U14007 ( .A(n14021), .B(n14022), .Z(n14019) );
  NOR2_X1 U14008 ( .A1(n8751), .A2(n8769), .ZN(n14022) );
  NAND2_X1 U14009 ( .A1(a_9_), .A2(n14018), .ZN(n13906) );
  NAND2_X1 U14010 ( .A1(n14023), .A2(n14024), .ZN(n14018) );
  NAND2_X1 U14011 ( .A1(n13898), .A2(n14025), .ZN(n14024) );
  NAND2_X1 U14012 ( .A1(n14026), .A2(n14027), .ZN(n14025) );
  NAND2_X1 U14013 ( .A1(b_12_), .A2(a_10_), .ZN(n14027) );
  XNOR2_X1 U14014 ( .A(n14028), .B(n14029), .ZN(n13898) );
  XNOR2_X1 U14015 ( .A(n14030), .B(n8746), .ZN(n14028) );
  INV_X1 U14016 ( .A(n13901), .ZN(n14023) );
  NOR2_X1 U14017 ( .A1(n14026), .A2(n8769), .ZN(n13901) );
  INV_X1 U14018 ( .A(n13902), .ZN(n14026) );
  NOR2_X1 U14019 ( .A1(n14031), .A2(n14032), .ZN(n13902) );
  INV_X1 U14020 ( .A(n14033), .ZN(n14032) );
  NAND2_X1 U14021 ( .A1(n13894), .A2(n14034), .ZN(n14033) );
  NAND2_X1 U14022 ( .A1(n13897), .A2(n13896), .ZN(n14034) );
  XNOR2_X1 U14023 ( .A(n14035), .B(n14036), .ZN(n13894) );
  XOR2_X1 U14024 ( .A(n14037), .B(n14038), .Z(n14035) );
  NOR2_X1 U14025 ( .A1(n8751), .A2(n8739), .ZN(n14038) );
  NOR2_X1 U14026 ( .A1(n13896), .A2(n13897), .ZN(n14031) );
  NOR2_X1 U14027 ( .A1(n13622), .A2(n8749), .ZN(n13897) );
  NAND2_X1 U14028 ( .A1(n14039), .A2(n14040), .ZN(n13896) );
  NAND2_X1 U14029 ( .A1(n13891), .A2(n14041), .ZN(n14040) );
  INV_X1 U14030 ( .A(n14042), .ZN(n14041) );
  NOR2_X1 U14031 ( .A1(n13893), .A2(n8733), .ZN(n14042) );
  XNOR2_X1 U14032 ( .A(n14043), .B(n14044), .ZN(n13891) );
  XOR2_X1 U14033 ( .A(n14045), .B(n14046), .Z(n14044) );
  NAND2_X1 U14034 ( .A1(a_13_), .A2(b_11_), .ZN(n14046) );
  NAND2_X1 U14035 ( .A1(n8733), .A2(n13893), .ZN(n14039) );
  NAND2_X1 U14036 ( .A1(n13749), .A2(n14047), .ZN(n13893) );
  NAND2_X1 U14037 ( .A1(n13748), .A2(n13750), .ZN(n14047) );
  NAND2_X1 U14038 ( .A1(n14048), .A2(n14049), .ZN(n13750) );
  NAND2_X1 U14039 ( .A1(b_12_), .A2(a_13_), .ZN(n14049) );
  INV_X1 U14040 ( .A(n14050), .ZN(n14048) );
  XNOR2_X1 U14041 ( .A(n14051), .B(n14052), .ZN(n13748) );
  XOR2_X1 U14042 ( .A(n14053), .B(n14054), .Z(n14052) );
  NAND2_X1 U14043 ( .A1(a_14_), .A2(b_11_), .ZN(n14054) );
  NAND2_X1 U14044 ( .A1(a_13_), .A2(n14050), .ZN(n13749) );
  NAND2_X1 U14045 ( .A1(n13757), .A2(n14055), .ZN(n14050) );
  NAND2_X1 U14046 ( .A1(n13756), .A2(n13758), .ZN(n14055) );
  NAND2_X1 U14047 ( .A1(n14056), .A2(n14057), .ZN(n13758) );
  NAND2_X1 U14048 ( .A1(b_12_), .A2(a_14_), .ZN(n14057) );
  INV_X1 U14049 ( .A(n14058), .ZN(n14056) );
  XOR2_X1 U14050 ( .A(n14059), .B(n14060), .Z(n13756) );
  XOR2_X1 U14051 ( .A(n14061), .B(n14062), .Z(n14059) );
  NOR2_X1 U14052 ( .A1(n8751), .A2(n8692), .ZN(n14062) );
  NAND2_X1 U14053 ( .A1(a_14_), .A2(n14058), .ZN(n13757) );
  NAND2_X1 U14054 ( .A1(n14063), .A2(n14064), .ZN(n14058) );
  INV_X1 U14055 ( .A(n14065), .ZN(n14064) );
  NOR3_X1 U14056 ( .A1(n8692), .A2(n14066), .A3(n13622), .ZN(n14065) );
  NOR2_X1 U14057 ( .A1(n13889), .A2(n13887), .ZN(n14066) );
  NAND2_X1 U14058 ( .A1(n13887), .A2(n13889), .ZN(n14063) );
  NAND2_X1 U14059 ( .A1(n14067), .A2(n14068), .ZN(n13889) );
  NAND2_X1 U14060 ( .A1(n13886), .A2(n14069), .ZN(n14068) );
  INV_X1 U14061 ( .A(n14070), .ZN(n14069) );
  NOR2_X1 U14062 ( .A1(n13885), .A2(n13884), .ZN(n14070) );
  NOR2_X1 U14063 ( .A1(n13622), .A2(n8680), .ZN(n13886) );
  NAND2_X1 U14064 ( .A1(n13884), .A2(n13885), .ZN(n14067) );
  NAND2_X1 U14065 ( .A1(n14071), .A2(n14072), .ZN(n13885) );
  NAND2_X1 U14066 ( .A1(n13882), .A2(n14073), .ZN(n14072) );
  NAND2_X1 U14067 ( .A1(n13880), .A2(n13881), .ZN(n14073) );
  NOR2_X1 U14068 ( .A1(n13622), .A2(n8662), .ZN(n13882) );
  INV_X1 U14069 ( .A(n14074), .ZN(n14071) );
  NOR2_X1 U14070 ( .A1(n13880), .A2(n13881), .ZN(n14074) );
  NOR2_X1 U14071 ( .A1(n14075), .A2(n14076), .ZN(n13881) );
  INV_X1 U14072 ( .A(n14077), .ZN(n14076) );
  NAND3_X1 U14073 ( .A1(a_18_), .A2(n14078), .A3(b_12_), .ZN(n14077) );
  NAND2_X1 U14074 ( .A1(n13877), .A2(n13875), .ZN(n14078) );
  NOR2_X1 U14075 ( .A1(n13875), .A2(n13877), .ZN(n14075) );
  NOR2_X1 U14076 ( .A1(n14079), .A2(n14080), .ZN(n13877) );
  NOR3_X1 U14077 ( .A1(n8630), .A2(n14081), .A3(n13622), .ZN(n14080) );
  INV_X1 U14078 ( .A(n14082), .ZN(n14081) );
  NAND2_X1 U14079 ( .A1(n13873), .A2(n13871), .ZN(n14082) );
  NOR2_X1 U14080 ( .A1(n13871), .A2(n13873), .ZN(n14079) );
  NOR2_X1 U14081 ( .A1(n14083), .A2(n14084), .ZN(n13873) );
  INV_X1 U14082 ( .A(n14085), .ZN(n14084) );
  NAND3_X1 U14083 ( .A1(a_20_), .A2(n14086), .A3(b_12_), .ZN(n14085) );
  NAND2_X1 U14084 ( .A1(n13868), .A2(n13869), .ZN(n14086) );
  NOR2_X1 U14085 ( .A1(n13868), .A2(n13869), .ZN(n14083) );
  NOR2_X1 U14086 ( .A1(n14087), .A2(n14088), .ZN(n13869) );
  NOR3_X1 U14087 ( .A1(n8601), .A2(n14089), .A3(n13622), .ZN(n14088) );
  NOR2_X1 U14088 ( .A1(n13865), .A2(n13864), .ZN(n14089) );
  INV_X1 U14089 ( .A(n14090), .ZN(n14087) );
  NAND2_X1 U14090 ( .A1(n13864), .A2(n13865), .ZN(n14090) );
  NAND2_X1 U14091 ( .A1(n14091), .A2(n14092), .ZN(n13865) );
  NAND2_X1 U14092 ( .A1(n13862), .A2(n14093), .ZN(n14092) );
  INV_X1 U14093 ( .A(n14094), .ZN(n14093) );
  NOR2_X1 U14094 ( .A1(n13859), .A2(n13861), .ZN(n14094) );
  NOR2_X1 U14095 ( .A1(n13622), .A2(n8984), .ZN(n13862) );
  NAND2_X1 U14096 ( .A1(n13859), .A2(n13861), .ZN(n14091) );
  NAND2_X1 U14097 ( .A1(n14095), .A2(n14096), .ZN(n13861) );
  NAND2_X1 U14098 ( .A1(n13858), .A2(n14097), .ZN(n14096) );
  INV_X1 U14099 ( .A(n14098), .ZN(n14097) );
  NOR2_X1 U14100 ( .A1(n13857), .A2(n13856), .ZN(n14098) );
  NOR2_X1 U14101 ( .A1(n13622), .A2(n8572), .ZN(n13858) );
  NAND2_X1 U14102 ( .A1(n13856), .A2(n13857), .ZN(n14095) );
  NAND2_X1 U14103 ( .A1(n14099), .A2(n14100), .ZN(n13857) );
  NAND2_X1 U14104 ( .A1(n13854), .A2(n14101), .ZN(n14100) );
  INV_X1 U14105 ( .A(n14102), .ZN(n14101) );
  NOR2_X1 U14106 ( .A1(n13852), .A2(n13853), .ZN(n14102) );
  NOR2_X1 U14107 ( .A1(n13622), .A2(n8982), .ZN(n13854) );
  NAND2_X1 U14108 ( .A1(n13852), .A2(n13853), .ZN(n14099) );
  NAND2_X1 U14109 ( .A1(n14103), .A2(n14104), .ZN(n13853) );
  NAND2_X1 U14110 ( .A1(n13850), .A2(n14105), .ZN(n14104) );
  NAND2_X1 U14111 ( .A1(n13847), .A2(n13849), .ZN(n14105) );
  NOR2_X1 U14112 ( .A1(n13622), .A2(n8541), .ZN(n13850) );
  INV_X1 U14113 ( .A(n14106), .ZN(n14103) );
  NOR2_X1 U14114 ( .A1(n13849), .A2(n13847), .ZN(n14106) );
  XNOR2_X1 U14115 ( .A(n14107), .B(n14108), .ZN(n13847) );
  XNOR2_X1 U14116 ( .A(n14109), .B(n14110), .ZN(n14108) );
  NAND2_X1 U14117 ( .A1(n14111), .A2(n14112), .ZN(n13849) );
  NAND2_X1 U14118 ( .A1(n13809), .A2(n14113), .ZN(n14112) );
  NAND2_X1 U14119 ( .A1(n13812), .A2(n13811), .ZN(n14113) );
  XNOR2_X1 U14120 ( .A(n14114), .B(n14115), .ZN(n13809) );
  XOR2_X1 U14121 ( .A(n14116), .B(n14117), .Z(n14114) );
  INV_X1 U14122 ( .A(n14118), .ZN(n14111) );
  NOR2_X1 U14123 ( .A1(n13811), .A2(n13812), .ZN(n14118) );
  NOR2_X1 U14124 ( .A1(n13622), .A2(n9893), .ZN(n13812) );
  NAND2_X1 U14125 ( .A1(n14119), .A2(n14120), .ZN(n13811) );
  NAND2_X1 U14126 ( .A1(n13819), .A2(n14121), .ZN(n14120) );
  INV_X1 U14127 ( .A(n14122), .ZN(n14121) );
  NOR2_X1 U14128 ( .A1(n13817), .A2(n13818), .ZN(n14122) );
  NOR2_X1 U14129 ( .A1(n13622), .A2(n8512), .ZN(n13819) );
  NAND2_X1 U14130 ( .A1(n13817), .A2(n13818), .ZN(n14119) );
  NAND2_X1 U14131 ( .A1(n14123), .A2(n14124), .ZN(n13818) );
  NAND2_X1 U14132 ( .A1(n13845), .A2(n14125), .ZN(n14124) );
  INV_X1 U14133 ( .A(n14126), .ZN(n14125) );
  NOR2_X1 U14134 ( .A1(n13846), .A2(n13844), .ZN(n14126) );
  NOR2_X1 U14135 ( .A1(n13622), .A2(n8493), .ZN(n13845) );
  NAND2_X1 U14136 ( .A1(n13844), .A2(n13846), .ZN(n14123) );
  NAND2_X1 U14137 ( .A1(n14127), .A2(n14128), .ZN(n13846) );
  NAND2_X1 U14138 ( .A1(n13840), .A2(n14129), .ZN(n14128) );
  INV_X1 U14139 ( .A(n14130), .ZN(n14129) );
  NOR2_X1 U14140 ( .A1(n13841), .A2(n13842), .ZN(n14130) );
  NOR2_X1 U14141 ( .A1(n13622), .A2(n8473), .ZN(n13840) );
  NAND2_X1 U14142 ( .A1(n13842), .A2(n13841), .ZN(n14127) );
  NAND2_X1 U14143 ( .A1(n14131), .A2(n14132), .ZN(n13841) );
  NAND2_X1 U14144 ( .A1(b_10_), .A2(n14133), .ZN(n14132) );
  NAND2_X1 U14145 ( .A1(n8456), .A2(n14134), .ZN(n14133) );
  NAND2_X1 U14146 ( .A1(a_31_), .A2(n8751), .ZN(n14134) );
  NAND2_X1 U14147 ( .A1(b_11_), .A2(n14135), .ZN(n14131) );
  NAND2_X1 U14148 ( .A1(n8459), .A2(n14136), .ZN(n14135) );
  NAND2_X1 U14149 ( .A1(a_30_), .A2(n8992), .ZN(n14136) );
  NOR3_X1 U14150 ( .A1(n8979), .A2(n8751), .A3(n13622), .ZN(n13842) );
  XOR2_X1 U14151 ( .A(n14137), .B(n14138), .Z(n13844) );
  XOR2_X1 U14152 ( .A(n14139), .B(n14140), .Z(n14137) );
  XOR2_X1 U14153 ( .A(n14141), .B(n14142), .Z(n13817) );
  XOR2_X1 U14154 ( .A(n14143), .B(n14144), .Z(n14141) );
  XNOR2_X1 U14155 ( .A(n14145), .B(n14146), .ZN(n13852) );
  XNOR2_X1 U14156 ( .A(n14147), .B(n14148), .ZN(n14146) );
  XOR2_X1 U14157 ( .A(n14149), .B(n14150), .Z(n13856) );
  XOR2_X1 U14158 ( .A(n14151), .B(n14152), .Z(n14149) );
  XOR2_X1 U14159 ( .A(n14153), .B(n14154), .Z(n13859) );
  XOR2_X1 U14160 ( .A(n14155), .B(n14156), .Z(n14153) );
  XNOR2_X1 U14161 ( .A(n14157), .B(n14158), .ZN(n13864) );
  XNOR2_X1 U14162 ( .A(n14159), .B(n14160), .ZN(n14158) );
  XNOR2_X1 U14163 ( .A(n14161), .B(n14162), .ZN(n13868) );
  XOR2_X1 U14164 ( .A(n14163), .B(n14164), .Z(n14161) );
  XNOR2_X1 U14165 ( .A(n14165), .B(n14166), .ZN(n13871) );
  XOR2_X1 U14166 ( .A(n14167), .B(n14168), .Z(n14165) );
  XOR2_X1 U14167 ( .A(n14169), .B(n14170), .Z(n13875) );
  XOR2_X1 U14168 ( .A(n14171), .B(n14172), .Z(n14170) );
  XOR2_X1 U14169 ( .A(n14173), .B(n14174), .Z(n13880) );
  NAND2_X1 U14170 ( .A1(n14175), .A2(n14176), .ZN(n14173) );
  XOR2_X1 U14171 ( .A(n14177), .B(n14178), .Z(n13884) );
  XOR2_X1 U14172 ( .A(n14179), .B(n14180), .Z(n14177) );
  NOR2_X1 U14173 ( .A1(n8751), .A2(n8662), .ZN(n14180) );
  XNOR2_X1 U14174 ( .A(n14181), .B(n14182), .ZN(n13887) );
  XOR2_X1 U14175 ( .A(n14183), .B(n14184), .Z(n14182) );
  NAND2_X1 U14176 ( .A1(a_16_), .A2(b_11_), .ZN(n14184) );
  NOR2_X1 U14177 ( .A1(n13622), .A2(n8739), .ZN(n8733) );
  INV_X1 U14178 ( .A(b_12_), .ZN(n13622) );
  XNOR2_X1 U14179 ( .A(n14185), .B(n14186), .ZN(n13938) );
  XOR2_X1 U14180 ( .A(n14187), .B(n14188), .Z(n14186) );
  NAND2_X1 U14181 ( .A1(a_2_), .A2(b_11_), .ZN(n14188) );
  XOR2_X1 U14182 ( .A(n14189), .B(n14190), .Z(n13943) );
  XNOR2_X1 U14183 ( .A(n14191), .B(n14192), .ZN(n14190) );
  NAND2_X1 U14184 ( .A1(a_1_), .A2(b_11_), .ZN(n14192) );
  XNOR2_X1 U14185 ( .A(n14193), .B(n14194), .ZN(n9125) );
  XNOR2_X1 U14186 ( .A(n14195), .B(n14196), .ZN(n14193) );
  NOR2_X1 U14187 ( .A1(n8751), .A2(n9471), .ZN(n14196) );
  NOR2_X1 U14188 ( .A1(n13949), .A2(n13948), .ZN(n9152) );
  NOR2_X1 U14189 ( .A1(n14197), .A2(n14198), .ZN(n13948) );
  INV_X1 U14190 ( .A(n14199), .ZN(n14198) );
  NAND3_X1 U14191 ( .A1(b_11_), .A2(n14200), .A3(a_0_), .ZN(n14199) );
  NAND2_X1 U14192 ( .A1(n14195), .A2(n14194), .ZN(n14200) );
  NOR2_X1 U14193 ( .A1(n14194), .A2(n14195), .ZN(n14197) );
  NOR2_X1 U14194 ( .A1(n14201), .A2(n14202), .ZN(n14195) );
  INV_X1 U14195 ( .A(n14203), .ZN(n14202) );
  NAND3_X1 U14196 ( .A1(b_11_), .A2(n14204), .A3(a_1_), .ZN(n14203) );
  NAND2_X1 U14197 ( .A1(n14191), .A2(n14189), .ZN(n14204) );
  NOR2_X1 U14198 ( .A1(n14189), .A2(n14191), .ZN(n14201) );
  NOR2_X1 U14199 ( .A1(n14205), .A2(n14206), .ZN(n14191) );
  NOR3_X1 U14200 ( .A1(n8751), .A2(n14207), .A3(n8998), .ZN(n14206) );
  NOR2_X1 U14201 ( .A1(n14187), .A2(n14185), .ZN(n14207) );
  INV_X1 U14202 ( .A(n14208), .ZN(n14205) );
  NAND2_X1 U14203 ( .A1(n14185), .A2(n14187), .ZN(n14208) );
  NAND2_X1 U14204 ( .A1(n14209), .A2(n14210), .ZN(n14187) );
  INV_X1 U14205 ( .A(n14211), .ZN(n14210) );
  NOR3_X1 U14206 ( .A1(n8751), .A2(n14212), .A3(n8877), .ZN(n14211) );
  NOR2_X1 U14207 ( .A1(n13964), .A2(n13962), .ZN(n14212) );
  NAND2_X1 U14208 ( .A1(n13962), .A2(n13964), .ZN(n14209) );
  NAND2_X1 U14209 ( .A1(n14213), .A2(n14214), .ZN(n13964) );
  NAND3_X1 U14210 ( .A1(b_11_), .A2(n14215), .A3(a_4_), .ZN(n14214) );
  NAND2_X1 U14211 ( .A1(n13972), .A2(n13970), .ZN(n14215) );
  INV_X1 U14212 ( .A(n14216), .ZN(n14213) );
  NOR2_X1 U14213 ( .A1(n13970), .A2(n13972), .ZN(n14216) );
  NOR2_X1 U14214 ( .A1(n14217), .A2(n14218), .ZN(n13972) );
  NOR3_X1 U14215 ( .A1(n8751), .A2(n14219), .A3(n8848), .ZN(n14218) );
  NOR2_X1 U14216 ( .A1(n13980), .A2(n13979), .ZN(n14219) );
  INV_X1 U14217 ( .A(n14220), .ZN(n14217) );
  NAND2_X1 U14218 ( .A1(n13979), .A2(n13980), .ZN(n14220) );
  NAND2_X1 U14219 ( .A1(n14221), .A2(n14222), .ZN(n13980) );
  NAND3_X1 U14220 ( .A1(b_11_), .A2(n14223), .A3(a_6_), .ZN(n14222) );
  INV_X1 U14221 ( .A(n14224), .ZN(n14223) );
  NOR2_X1 U14222 ( .A1(n13988), .A2(n13986), .ZN(n14224) );
  NAND2_X1 U14223 ( .A1(n13986), .A2(n13988), .ZN(n14221) );
  NAND2_X1 U14224 ( .A1(n14225), .A2(n14226), .ZN(n13988) );
  NAND3_X1 U14225 ( .A1(b_11_), .A2(n14227), .A3(a_7_), .ZN(n14226) );
  INV_X1 U14226 ( .A(n14228), .ZN(n14227) );
  NOR2_X1 U14227 ( .A1(n13996), .A2(n13995), .ZN(n14228) );
  NAND2_X1 U14228 ( .A1(n13995), .A2(n13996), .ZN(n14225) );
  NAND2_X1 U14229 ( .A1(n14229), .A2(n14230), .ZN(n13996) );
  NAND3_X1 U14230 ( .A1(b_11_), .A2(n14231), .A3(a_8_), .ZN(n14230) );
  NAND2_X1 U14231 ( .A1(n14004), .A2(n14002), .ZN(n14231) );
  INV_X1 U14232 ( .A(n14232), .ZN(n14229) );
  NOR2_X1 U14233 ( .A1(n14002), .A2(n14004), .ZN(n14232) );
  NOR2_X1 U14234 ( .A1(n14233), .A2(n14234), .ZN(n14004) );
  INV_X1 U14235 ( .A(n14235), .ZN(n14234) );
  NAND3_X1 U14236 ( .A1(b_11_), .A2(n14236), .A3(a_9_), .ZN(n14235) );
  NAND2_X1 U14237 ( .A1(n14013), .A2(n14012), .ZN(n14236) );
  NOR2_X1 U14238 ( .A1(n14012), .A2(n14013), .ZN(n14233) );
  NOR2_X1 U14239 ( .A1(n14237), .A2(n14238), .ZN(n14013) );
  INV_X1 U14240 ( .A(n14239), .ZN(n14238) );
  NAND3_X1 U14241 ( .A1(b_11_), .A2(n14240), .A3(a_10_), .ZN(n14239) );
  NAND2_X1 U14242 ( .A1(n14020), .A2(n14021), .ZN(n14240) );
  NOR2_X1 U14243 ( .A1(n14021), .A2(n14020), .ZN(n14237) );
  XOR2_X1 U14244 ( .A(n14241), .B(n14242), .Z(n14020) );
  NAND2_X1 U14245 ( .A1(n14243), .A2(n14244), .ZN(n14241) );
  NAND2_X1 U14246 ( .A1(n14245), .A2(n14246), .ZN(n14021) );
  NAND2_X1 U14247 ( .A1(n14029), .A2(n14247), .ZN(n14246) );
  NAND2_X1 U14248 ( .A1(n8746), .A2(n14248), .ZN(n14247) );
  XNOR2_X1 U14249 ( .A(n14249), .B(n14250), .ZN(n14029) );
  XOR2_X1 U14250 ( .A(n14251), .B(n14252), .Z(n14249) );
  NOR2_X1 U14251 ( .A1(n8992), .A2(n8739), .ZN(n14252) );
  NAND2_X1 U14252 ( .A1(n14030), .A2(n8937), .ZN(n14245) );
  INV_X1 U14253 ( .A(n8746), .ZN(n8937) );
  NOR2_X1 U14254 ( .A1(n8749), .A2(n8751), .ZN(n8746) );
  INV_X1 U14255 ( .A(n14248), .ZN(n14030) );
  NAND2_X1 U14256 ( .A1(n14253), .A2(n14254), .ZN(n14248) );
  NAND3_X1 U14257 ( .A1(b_11_), .A2(n14255), .A3(a_12_), .ZN(n14254) );
  INV_X1 U14258 ( .A(n14256), .ZN(n14255) );
  NOR2_X1 U14259 ( .A1(n14037), .A2(n14036), .ZN(n14256) );
  NAND2_X1 U14260 ( .A1(n14036), .A2(n14037), .ZN(n14253) );
  NAND2_X1 U14261 ( .A1(n14257), .A2(n14258), .ZN(n14037) );
  NAND3_X1 U14262 ( .A1(b_11_), .A2(n14259), .A3(a_13_), .ZN(n14258) );
  INV_X1 U14263 ( .A(n14260), .ZN(n14259) );
  NOR2_X1 U14264 ( .A1(n14045), .A2(n14043), .ZN(n14260) );
  NAND2_X1 U14265 ( .A1(n14043), .A2(n14045), .ZN(n14257) );
  NAND2_X1 U14266 ( .A1(n14261), .A2(n14262), .ZN(n14045) );
  INV_X1 U14267 ( .A(n14263), .ZN(n14262) );
  NOR3_X1 U14268 ( .A1(n8751), .A2(n14264), .A3(n8991), .ZN(n14263) );
  NOR2_X1 U14269 ( .A1(n14053), .A2(n14051), .ZN(n14264) );
  NAND2_X1 U14270 ( .A1(n14051), .A2(n14053), .ZN(n14261) );
  NAND2_X1 U14271 ( .A1(n14265), .A2(n14266), .ZN(n14053) );
  NAND3_X1 U14272 ( .A1(b_11_), .A2(n14267), .A3(a_15_), .ZN(n14266) );
  INV_X1 U14273 ( .A(n14268), .ZN(n14267) );
  NOR2_X1 U14274 ( .A1(n14061), .A2(n14060), .ZN(n14268) );
  NAND2_X1 U14275 ( .A1(n14060), .A2(n14061), .ZN(n14265) );
  NAND2_X1 U14276 ( .A1(n14269), .A2(n14270), .ZN(n14061) );
  INV_X1 U14277 ( .A(n14271), .ZN(n14270) );
  NOR3_X1 U14278 ( .A1(n8751), .A2(n14272), .A3(n8680), .ZN(n14271) );
  NOR2_X1 U14279 ( .A1(n14183), .A2(n14181), .ZN(n14272) );
  NAND2_X1 U14280 ( .A1(n14181), .A2(n14183), .ZN(n14269) );
  NAND2_X1 U14281 ( .A1(n14273), .A2(n14274), .ZN(n14183) );
  NAND3_X1 U14282 ( .A1(b_11_), .A2(n14275), .A3(a_17_), .ZN(n14274) );
  INV_X1 U14283 ( .A(n14276), .ZN(n14275) );
  NOR2_X1 U14284 ( .A1(n14179), .A2(n14178), .ZN(n14276) );
  NAND2_X1 U14285 ( .A1(n14178), .A2(n14179), .ZN(n14273) );
  NAND2_X1 U14286 ( .A1(n14175), .A2(n14277), .ZN(n14179) );
  NAND2_X1 U14287 ( .A1(n14174), .A2(n14176), .ZN(n14277) );
  NAND2_X1 U14288 ( .A1(n14278), .A2(n14279), .ZN(n14176) );
  NAND2_X1 U14289 ( .A1(a_18_), .A2(b_11_), .ZN(n14279) );
  XOR2_X1 U14290 ( .A(n14280), .B(n14281), .Z(n14174) );
  XOR2_X1 U14291 ( .A(n14282), .B(n14283), .Z(n14281) );
  NAND2_X1 U14292 ( .A1(a_18_), .A2(n14284), .ZN(n14175) );
  INV_X1 U14293 ( .A(n14278), .ZN(n14284) );
  NOR2_X1 U14294 ( .A1(n14285), .A2(n14286), .ZN(n14278) );
  NOR2_X1 U14295 ( .A1(n14172), .A2(n14287), .ZN(n14286) );
  NOR2_X1 U14296 ( .A1(n14171), .A2(n14169), .ZN(n14287) );
  NAND2_X1 U14297 ( .A1(b_11_), .A2(a_19_), .ZN(n14172) );
  INV_X1 U14298 ( .A(n14288), .ZN(n14285) );
  NAND2_X1 U14299 ( .A1(n14169), .A2(n14171), .ZN(n14288) );
  NAND2_X1 U14300 ( .A1(n14289), .A2(n14290), .ZN(n14171) );
  NAND2_X1 U14301 ( .A1(n14168), .A2(n14291), .ZN(n14290) );
  INV_X1 U14302 ( .A(n14292), .ZN(n14291) );
  NOR2_X1 U14303 ( .A1(n14167), .A2(n14166), .ZN(n14292) );
  NOR2_X1 U14304 ( .A1(n8986), .A2(n8751), .ZN(n14168) );
  NAND2_X1 U14305 ( .A1(n14166), .A2(n14167), .ZN(n14289) );
  NAND2_X1 U14306 ( .A1(n14293), .A2(n14294), .ZN(n14167) );
  NAND2_X1 U14307 ( .A1(n14164), .A2(n14295), .ZN(n14294) );
  INV_X1 U14308 ( .A(n14296), .ZN(n14295) );
  NOR2_X1 U14309 ( .A1(n14163), .A2(n14162), .ZN(n14296) );
  NOR2_X1 U14310 ( .A1(n8601), .A2(n8751), .ZN(n14164) );
  NAND2_X1 U14311 ( .A1(n14162), .A2(n14163), .ZN(n14293) );
  NAND2_X1 U14312 ( .A1(n14297), .A2(n14298), .ZN(n14163) );
  NAND2_X1 U14313 ( .A1(n14160), .A2(n14299), .ZN(n14298) );
  INV_X1 U14314 ( .A(n14300), .ZN(n14299) );
  NOR2_X1 U14315 ( .A1(n14159), .A2(n14157), .ZN(n14300) );
  NOR2_X1 U14316 ( .A1(n8984), .A2(n8751), .ZN(n14160) );
  NAND2_X1 U14317 ( .A1(n14157), .A2(n14159), .ZN(n14297) );
  NAND2_X1 U14318 ( .A1(n14301), .A2(n14302), .ZN(n14159) );
  NAND2_X1 U14319 ( .A1(n14156), .A2(n14303), .ZN(n14302) );
  INV_X1 U14320 ( .A(n14304), .ZN(n14303) );
  NOR2_X1 U14321 ( .A1(n14155), .A2(n14154), .ZN(n14304) );
  NOR2_X1 U14322 ( .A1(n8572), .A2(n8751), .ZN(n14156) );
  NAND2_X1 U14323 ( .A1(n14154), .A2(n14155), .ZN(n14301) );
  NAND2_X1 U14324 ( .A1(n14305), .A2(n14306), .ZN(n14155) );
  NAND2_X1 U14325 ( .A1(n14152), .A2(n14307), .ZN(n14306) );
  INV_X1 U14326 ( .A(n14308), .ZN(n14307) );
  NOR2_X1 U14327 ( .A1(n14151), .A2(n14150), .ZN(n14308) );
  NOR2_X1 U14328 ( .A1(n8982), .A2(n8751), .ZN(n14152) );
  NAND2_X1 U14329 ( .A1(n14150), .A2(n14151), .ZN(n14305) );
  NAND2_X1 U14330 ( .A1(n14309), .A2(n14310), .ZN(n14151) );
  NAND2_X1 U14331 ( .A1(n14148), .A2(n14311), .ZN(n14310) );
  NAND2_X1 U14332 ( .A1(n14145), .A2(n14147), .ZN(n14311) );
  NOR2_X1 U14333 ( .A1(n8541), .A2(n8751), .ZN(n14148) );
  INV_X1 U14334 ( .A(n14312), .ZN(n14309) );
  NOR2_X1 U14335 ( .A1(n14147), .A2(n14145), .ZN(n14312) );
  XNOR2_X1 U14336 ( .A(n14313), .B(n14314), .ZN(n14145) );
  XNOR2_X1 U14337 ( .A(n14315), .B(n14316), .ZN(n14314) );
  NAND2_X1 U14338 ( .A1(n14317), .A2(n14318), .ZN(n14147) );
  NAND2_X1 U14339 ( .A1(n14107), .A2(n14319), .ZN(n14318) );
  NAND2_X1 U14340 ( .A1(n14110), .A2(n14109), .ZN(n14319) );
  XNOR2_X1 U14341 ( .A(n14320), .B(n14321), .ZN(n14107) );
  XOR2_X1 U14342 ( .A(n14322), .B(n14323), .Z(n14320) );
  INV_X1 U14343 ( .A(n14324), .ZN(n14317) );
  NOR2_X1 U14344 ( .A1(n14109), .A2(n14110), .ZN(n14324) );
  NOR2_X1 U14345 ( .A1(n9893), .A2(n8751), .ZN(n14110) );
  NAND2_X1 U14346 ( .A1(n14325), .A2(n14326), .ZN(n14109) );
  NAND2_X1 U14347 ( .A1(n14117), .A2(n14327), .ZN(n14326) );
  INV_X1 U14348 ( .A(n14328), .ZN(n14327) );
  NOR2_X1 U14349 ( .A1(n14116), .A2(n14115), .ZN(n14328) );
  NOR2_X1 U14350 ( .A1(n8512), .A2(n8751), .ZN(n14117) );
  NAND2_X1 U14351 ( .A1(n14115), .A2(n14116), .ZN(n14325) );
  NAND2_X1 U14352 ( .A1(n14329), .A2(n14330), .ZN(n14116) );
  NAND2_X1 U14353 ( .A1(n14143), .A2(n14331), .ZN(n14330) );
  INV_X1 U14354 ( .A(n14332), .ZN(n14331) );
  NOR2_X1 U14355 ( .A1(n14144), .A2(n14142), .ZN(n14332) );
  NOR2_X1 U14356 ( .A1(n8493), .A2(n8751), .ZN(n14143) );
  NAND2_X1 U14357 ( .A1(n14142), .A2(n14144), .ZN(n14329) );
  NAND2_X1 U14358 ( .A1(n14333), .A2(n14334), .ZN(n14144) );
  NAND2_X1 U14359 ( .A1(n14138), .A2(n14335), .ZN(n14334) );
  INV_X1 U14360 ( .A(n14336), .ZN(n14335) );
  NOR2_X1 U14361 ( .A1(n14139), .A2(n14140), .ZN(n14336) );
  NOR2_X1 U14362 ( .A1(n8473), .A2(n8751), .ZN(n14138) );
  NAND2_X1 U14363 ( .A1(n14140), .A2(n14139), .ZN(n14333) );
  NAND2_X1 U14364 ( .A1(n14337), .A2(n14338), .ZN(n14139) );
  NAND2_X1 U14365 ( .A1(b_10_), .A2(n14339), .ZN(n14338) );
  NAND2_X1 U14366 ( .A1(n8459), .A2(n14340), .ZN(n14339) );
  NAND2_X1 U14367 ( .A1(a_30_), .A2(n8781), .ZN(n14340) );
  NAND2_X1 U14368 ( .A1(b_9_), .A2(n14341), .ZN(n14337) );
  NAND2_X1 U14369 ( .A1(n8456), .A2(n14342), .ZN(n14341) );
  NAND2_X1 U14370 ( .A1(a_31_), .A2(n8992), .ZN(n14342) );
  NOR3_X1 U14371 ( .A1(n8979), .A2(n8751), .A3(n8992), .ZN(n14140) );
  XOR2_X1 U14372 ( .A(n14343), .B(n14344), .Z(n14142) );
  XOR2_X1 U14373 ( .A(n14345), .B(n14346), .Z(n14343) );
  XOR2_X1 U14374 ( .A(n14347), .B(n14348), .Z(n14115) );
  XOR2_X1 U14375 ( .A(n14349), .B(n14350), .Z(n14347) );
  XNOR2_X1 U14376 ( .A(n14351), .B(n14352), .ZN(n14150) );
  XNOR2_X1 U14377 ( .A(n14353), .B(n14354), .ZN(n14352) );
  XOR2_X1 U14378 ( .A(n14355), .B(n14356), .Z(n14154) );
  XOR2_X1 U14379 ( .A(n14357), .B(n14358), .Z(n14355) );
  XOR2_X1 U14380 ( .A(n14359), .B(n14360), .Z(n14157) );
  XOR2_X1 U14381 ( .A(n14361), .B(n14362), .Z(n14359) );
  XNOR2_X1 U14382 ( .A(n14363), .B(n14364), .ZN(n14162) );
  XNOR2_X1 U14383 ( .A(n14365), .B(n14366), .ZN(n14364) );
  XOR2_X1 U14384 ( .A(n14367), .B(n14368), .Z(n14166) );
  XOR2_X1 U14385 ( .A(n14369), .B(n14370), .Z(n14367) );
  NOR2_X1 U14386 ( .A1(n8601), .A2(n8992), .ZN(n14370) );
  XNOR2_X1 U14387 ( .A(n14371), .B(n14372), .ZN(n14169) );
  XNOR2_X1 U14388 ( .A(n14373), .B(n14374), .ZN(n14371) );
  NOR2_X1 U14389 ( .A1(n8986), .A2(n8992), .ZN(n14374) );
  XOR2_X1 U14390 ( .A(n14375), .B(n14376), .Z(n14178) );
  XOR2_X1 U14391 ( .A(n14377), .B(n14378), .Z(n14375) );
  NOR2_X1 U14392 ( .A1(n8992), .A2(n8988), .ZN(n14378) );
  XNOR2_X1 U14393 ( .A(n14379), .B(n14380), .ZN(n14181) );
  NAND2_X1 U14394 ( .A1(n14381), .A2(n14382), .ZN(n14379) );
  XNOR2_X1 U14395 ( .A(n14383), .B(n14384), .ZN(n14060) );
  NAND2_X1 U14396 ( .A1(n14385), .A2(n14386), .ZN(n14383) );
  XNOR2_X1 U14397 ( .A(n14387), .B(n14388), .ZN(n14051) );
  NAND2_X1 U14398 ( .A1(n14389), .A2(n14390), .ZN(n14387) );
  XNOR2_X1 U14399 ( .A(n14391), .B(n14392), .ZN(n14043) );
  XOR2_X1 U14400 ( .A(n14393), .B(n14394), .Z(n14392) );
  NAND2_X1 U14401 ( .A1(a_14_), .A2(b_10_), .ZN(n14394) );
  XNOR2_X1 U14402 ( .A(n14395), .B(n14396), .ZN(n14036) );
  NAND2_X1 U14403 ( .A1(n14397), .A2(n14398), .ZN(n14395) );
  XNOR2_X1 U14404 ( .A(n14399), .B(n14400), .ZN(n14012) );
  XOR2_X1 U14405 ( .A(n14401), .B(n8763), .Z(n14399) );
  XOR2_X1 U14406 ( .A(n14402), .B(n14403), .Z(n14002) );
  NAND2_X1 U14407 ( .A1(n14404), .A2(n14405), .ZN(n14402) );
  XNOR2_X1 U14408 ( .A(n14406), .B(n14407), .ZN(n13995) );
  XOR2_X1 U14409 ( .A(n14408), .B(n14409), .Z(n14406) );
  XNOR2_X1 U14410 ( .A(n14410), .B(n14411), .ZN(n13986) );
  XNOR2_X1 U14411 ( .A(n14412), .B(n14413), .ZN(n14411) );
  XOR2_X1 U14412 ( .A(n14414), .B(n14415), .Z(n13979) );
  XOR2_X1 U14413 ( .A(n14416), .B(n14417), .Z(n14414) );
  XNOR2_X1 U14414 ( .A(n14418), .B(n14419), .ZN(n13970) );
  XOR2_X1 U14415 ( .A(n14420), .B(n14421), .Z(n14418) );
  XOR2_X1 U14416 ( .A(n14422), .B(n14423), .Z(n13962) );
  XOR2_X1 U14417 ( .A(n14424), .B(n14425), .Z(n14422) );
  XOR2_X1 U14418 ( .A(n14426), .B(n14427), .Z(n14185) );
  XOR2_X1 U14419 ( .A(n14428), .B(n14429), .Z(n14426) );
  XNOR2_X1 U14420 ( .A(n14430), .B(n14431), .ZN(n14189) );
  XOR2_X1 U14421 ( .A(n14432), .B(n14433), .Z(n14430) );
  XNOR2_X1 U14422 ( .A(n14434), .B(n14435), .ZN(n14194) );
  XOR2_X1 U14423 ( .A(n14436), .B(n14437), .Z(n14434) );
  NOR2_X1 U14424 ( .A1(n8992), .A2(n9731), .ZN(n14437) );
  XOR2_X1 U14425 ( .A(n14438), .B(n14439), .Z(n13949) );
  XNOR2_X1 U14426 ( .A(n14440), .B(n14441), .ZN(n14439) );
  NOR2_X1 U14427 ( .A1(n8992), .A2(n9471), .ZN(n14441) );
  XNOR2_X1 U14428 ( .A(n8429), .B(n8428), .ZN(n9129) );
  NAND3_X1 U14429 ( .A1(n8428), .A2(n8429), .A3(n9151), .ZN(n8424) );
  INV_X1 U14430 ( .A(n8427), .ZN(n9151) );
  NAND2_X1 U14431 ( .A1(n9148), .A2(n14442), .ZN(n8427) );
  NAND2_X1 U14432 ( .A1(n14443), .A2(n14444), .ZN(n14442) );
  XNOR2_X1 U14433 ( .A(n14445), .B(n14446), .ZN(n14444) );
  NAND2_X1 U14434 ( .A1(n14447), .A2(n14448), .ZN(n9148) );
  INV_X1 U14435 ( .A(n14443), .ZN(n14448) );
  NOR2_X1 U14436 ( .A1(n14449), .A2(n14450), .ZN(n14443) );
  INV_X1 U14437 ( .A(n14451), .ZN(n14450) );
  NAND2_X1 U14438 ( .A1(n14452), .A2(n14453), .ZN(n14451) );
  NAND2_X1 U14439 ( .A1(n14454), .A2(n14455), .ZN(n14453) );
  NOR2_X1 U14440 ( .A1(n14454), .A2(n14455), .ZN(n14449) );
  XOR2_X1 U14441 ( .A(n14445), .B(n14446), .Z(n14447) );
  XOR2_X1 U14442 ( .A(n14456), .B(n14457), .Z(n14445) );
  NOR2_X1 U14443 ( .A1(n14458), .A2(n9471), .ZN(n14457) );
  NAND2_X1 U14444 ( .A1(n14459), .A2(n14460), .ZN(n8429) );
  NAND3_X1 U14445 ( .A1(b_10_), .A2(n14461), .A3(a_0_), .ZN(n14460) );
  INV_X1 U14446 ( .A(n14462), .ZN(n14461) );
  NOR2_X1 U14447 ( .A1(n14438), .A2(n14440), .ZN(n14462) );
  NAND2_X1 U14448 ( .A1(n14438), .A2(n14440), .ZN(n14459) );
  NAND2_X1 U14449 ( .A1(n14463), .A2(n14464), .ZN(n14440) );
  NAND3_X1 U14450 ( .A1(b_10_), .A2(n14465), .A3(a_1_), .ZN(n14464) );
  INV_X1 U14451 ( .A(n14466), .ZN(n14465) );
  NOR2_X1 U14452 ( .A1(n14435), .A2(n14436), .ZN(n14466) );
  NAND2_X1 U14453 ( .A1(n14435), .A2(n14436), .ZN(n14463) );
  NAND2_X1 U14454 ( .A1(n14467), .A2(n14468), .ZN(n14436) );
  NAND2_X1 U14455 ( .A1(n14433), .A2(n14469), .ZN(n14468) );
  INV_X1 U14456 ( .A(n14470), .ZN(n14469) );
  NOR2_X1 U14457 ( .A1(n14431), .A2(n14432), .ZN(n14470) );
  NOR2_X1 U14458 ( .A1(n8998), .A2(n8992), .ZN(n14433) );
  NAND2_X1 U14459 ( .A1(n14431), .A2(n14432), .ZN(n14467) );
  NAND2_X1 U14460 ( .A1(n14471), .A2(n14472), .ZN(n14432) );
  NAND2_X1 U14461 ( .A1(n14429), .A2(n14473), .ZN(n14472) );
  INV_X1 U14462 ( .A(n14474), .ZN(n14473) );
  NOR2_X1 U14463 ( .A1(n14427), .A2(n14428), .ZN(n14474) );
  NOR2_X1 U14464 ( .A1(n8877), .A2(n8992), .ZN(n14429) );
  NAND2_X1 U14465 ( .A1(n14427), .A2(n14428), .ZN(n14471) );
  NAND2_X1 U14466 ( .A1(n14475), .A2(n14476), .ZN(n14428) );
  NAND2_X1 U14467 ( .A1(n14425), .A2(n14477), .ZN(n14476) );
  INV_X1 U14468 ( .A(n14478), .ZN(n14477) );
  NOR2_X1 U14469 ( .A1(n14423), .A2(n14424), .ZN(n14478) );
  NOR2_X1 U14470 ( .A1(n8996), .A2(n8992), .ZN(n14425) );
  NAND2_X1 U14471 ( .A1(n14423), .A2(n14424), .ZN(n14475) );
  NAND2_X1 U14472 ( .A1(n14479), .A2(n14480), .ZN(n14424) );
  NAND2_X1 U14473 ( .A1(n14421), .A2(n14481), .ZN(n14480) );
  INV_X1 U14474 ( .A(n14482), .ZN(n14481) );
  NOR2_X1 U14475 ( .A1(n14419), .A2(n14420), .ZN(n14482) );
  NOR2_X1 U14476 ( .A1(n8848), .A2(n8992), .ZN(n14421) );
  NAND2_X1 U14477 ( .A1(n14419), .A2(n14420), .ZN(n14479) );
  NAND2_X1 U14478 ( .A1(n14483), .A2(n14484), .ZN(n14420) );
  NAND2_X1 U14479 ( .A1(n14417), .A2(n14485), .ZN(n14484) );
  INV_X1 U14480 ( .A(n14486), .ZN(n14485) );
  NOR2_X1 U14481 ( .A1(n14415), .A2(n14416), .ZN(n14486) );
  NOR2_X1 U14482 ( .A1(n8994), .A2(n8992), .ZN(n14417) );
  NAND2_X1 U14483 ( .A1(n14415), .A2(n14416), .ZN(n14483) );
  NAND2_X1 U14484 ( .A1(n14487), .A2(n14488), .ZN(n14416) );
  NAND2_X1 U14485 ( .A1(n14413), .A2(n14489), .ZN(n14488) );
  NAND2_X1 U14486 ( .A1(n14410), .A2(n14412), .ZN(n14489) );
  NOR2_X1 U14487 ( .A1(n8817), .A2(n8992), .ZN(n14413) );
  INV_X1 U14488 ( .A(n14490), .ZN(n14487) );
  NOR2_X1 U14489 ( .A1(n14412), .A2(n14410), .ZN(n14490) );
  XOR2_X1 U14490 ( .A(n14491), .B(n14492), .Z(n14410) );
  XOR2_X1 U14491 ( .A(n14493), .B(n14494), .Z(n14492) );
  NAND2_X1 U14492 ( .A1(a_8_), .A2(b_9_), .ZN(n14494) );
  NAND2_X1 U14493 ( .A1(n14495), .A2(n14496), .ZN(n14412) );
  NAND2_X1 U14494 ( .A1(n14407), .A2(n14497), .ZN(n14496) );
  NAND2_X1 U14495 ( .A1(n14409), .A2(n14408), .ZN(n14497) );
  XNOR2_X1 U14496 ( .A(n14498), .B(n14499), .ZN(n14407) );
  XNOR2_X1 U14497 ( .A(n14500), .B(n8776), .ZN(n14499) );
  INV_X1 U14498 ( .A(n14501), .ZN(n14495) );
  NOR2_X1 U14499 ( .A1(n14408), .A2(n14409), .ZN(n14501) );
  NOR2_X1 U14500 ( .A1(n10513), .A2(n8992), .ZN(n14409) );
  NAND2_X1 U14501 ( .A1(n14404), .A2(n14502), .ZN(n14408) );
  NAND2_X1 U14502 ( .A1(n14403), .A2(n14405), .ZN(n14502) );
  NAND2_X1 U14503 ( .A1(n14503), .A2(n14504), .ZN(n14405) );
  NAND2_X1 U14504 ( .A1(a_9_), .A2(b_10_), .ZN(n14504) );
  INV_X1 U14505 ( .A(n14505), .ZN(n14503) );
  XNOR2_X1 U14506 ( .A(n14506), .B(n14507), .ZN(n14403) );
  XOR2_X1 U14507 ( .A(n14508), .B(n14509), .Z(n14507) );
  NAND2_X1 U14508 ( .A1(a_10_), .A2(b_9_), .ZN(n14509) );
  NAND2_X1 U14509 ( .A1(a_9_), .A2(n14505), .ZN(n14404) );
  NAND2_X1 U14510 ( .A1(n14510), .A2(n14511), .ZN(n14505) );
  NAND2_X1 U14511 ( .A1(n14400), .A2(n14512), .ZN(n14511) );
  NAND2_X1 U14512 ( .A1(n14401), .A2(n8763), .ZN(n14512) );
  INV_X1 U14513 ( .A(n14513), .ZN(n14401) );
  XOR2_X1 U14514 ( .A(n14514), .B(n14515), .Z(n14400) );
  XNOR2_X1 U14515 ( .A(n14516), .B(n14517), .ZN(n14515) );
  NAND2_X1 U14516 ( .A1(a_11_), .A2(b_9_), .ZN(n14517) );
  NAND2_X1 U14517 ( .A1(n14518), .A2(n14513), .ZN(n14510) );
  NAND2_X1 U14518 ( .A1(n14243), .A2(n14519), .ZN(n14513) );
  NAND2_X1 U14519 ( .A1(n14242), .A2(n14244), .ZN(n14519) );
  NAND2_X1 U14520 ( .A1(n14520), .A2(n14521), .ZN(n14244) );
  NAND2_X1 U14521 ( .A1(a_11_), .A2(b_10_), .ZN(n14521) );
  XNOR2_X1 U14522 ( .A(n14522), .B(n14523), .ZN(n14242) );
  XNOR2_X1 U14523 ( .A(n14524), .B(n14525), .ZN(n14522) );
  NOR2_X1 U14524 ( .A1(n8781), .A2(n8739), .ZN(n14525) );
  NAND2_X1 U14525 ( .A1(a_11_), .A2(n14526), .ZN(n14243) );
  INV_X1 U14526 ( .A(n14520), .ZN(n14526) );
  NOR2_X1 U14527 ( .A1(n14527), .A2(n14528), .ZN(n14520) );
  NOR3_X1 U14528 ( .A1(n8992), .A2(n14529), .A3(n8739), .ZN(n14528) );
  NOR2_X1 U14529 ( .A1(n14250), .A2(n14251), .ZN(n14529) );
  INV_X1 U14530 ( .A(n14530), .ZN(n14527) );
  NAND2_X1 U14531 ( .A1(n14250), .A2(n14251), .ZN(n14530) );
  NAND2_X1 U14532 ( .A1(n14397), .A2(n14531), .ZN(n14251) );
  NAND2_X1 U14533 ( .A1(n14396), .A2(n14398), .ZN(n14531) );
  NAND2_X1 U14534 ( .A1(n14532), .A2(n14533), .ZN(n14398) );
  NAND2_X1 U14535 ( .A1(a_13_), .A2(b_10_), .ZN(n14533) );
  XNOR2_X1 U14536 ( .A(n14534), .B(n14535), .ZN(n14396) );
  XNOR2_X1 U14537 ( .A(n14536), .B(n14537), .ZN(n14534) );
  NOR2_X1 U14538 ( .A1(n8781), .A2(n8991), .ZN(n14537) );
  INV_X1 U14539 ( .A(n14538), .ZN(n14397) );
  NOR2_X1 U14540 ( .A1(n8721), .A2(n14532), .ZN(n14538) );
  NOR2_X1 U14541 ( .A1(n14539), .A2(n14540), .ZN(n14532) );
  NOR3_X1 U14542 ( .A1(n8992), .A2(n14541), .A3(n8991), .ZN(n14540) );
  NOR2_X1 U14543 ( .A1(n14393), .A2(n14391), .ZN(n14541) );
  INV_X1 U14544 ( .A(n14542), .ZN(n14539) );
  NAND2_X1 U14545 ( .A1(n14391), .A2(n14393), .ZN(n14542) );
  NAND2_X1 U14546 ( .A1(n14389), .A2(n14543), .ZN(n14393) );
  NAND2_X1 U14547 ( .A1(n14388), .A2(n14390), .ZN(n14543) );
  NAND2_X1 U14548 ( .A1(n14544), .A2(n14545), .ZN(n14390) );
  NAND2_X1 U14549 ( .A1(a_15_), .A2(b_10_), .ZN(n14545) );
  INV_X1 U14550 ( .A(n14546), .ZN(n14544) );
  XOR2_X1 U14551 ( .A(n14547), .B(n14548), .Z(n14388) );
  XNOR2_X1 U14552 ( .A(n14549), .B(n14550), .ZN(n14548) );
  NAND2_X1 U14553 ( .A1(a_16_), .A2(b_9_), .ZN(n14550) );
  NAND2_X1 U14554 ( .A1(a_15_), .A2(n14546), .ZN(n14389) );
  NAND2_X1 U14555 ( .A1(n14385), .A2(n14551), .ZN(n14546) );
  NAND2_X1 U14556 ( .A1(n14384), .A2(n14386), .ZN(n14551) );
  NAND2_X1 U14557 ( .A1(n14552), .A2(n14553), .ZN(n14386) );
  NAND2_X1 U14558 ( .A1(a_16_), .A2(b_10_), .ZN(n14553) );
  INV_X1 U14559 ( .A(n14554), .ZN(n14552) );
  XNOR2_X1 U14560 ( .A(n14555), .B(n14556), .ZN(n14384) );
  XNOR2_X1 U14561 ( .A(n14557), .B(n14558), .ZN(n14555) );
  NOR2_X1 U14562 ( .A1(n8781), .A2(n8662), .ZN(n14558) );
  NAND2_X1 U14563 ( .A1(a_16_), .A2(n14554), .ZN(n14385) );
  NAND2_X1 U14564 ( .A1(n14381), .A2(n14559), .ZN(n14554) );
  NAND2_X1 U14565 ( .A1(n14380), .A2(n14382), .ZN(n14559) );
  NAND2_X1 U14566 ( .A1(n14560), .A2(n14561), .ZN(n14382) );
  NAND2_X1 U14567 ( .A1(a_17_), .A2(b_10_), .ZN(n14561) );
  XNOR2_X1 U14568 ( .A(n14562), .B(n14563), .ZN(n14380) );
  XOR2_X1 U14569 ( .A(n14564), .B(n14565), .Z(n14563) );
  NAND2_X1 U14570 ( .A1(a_18_), .A2(b_9_), .ZN(n14565) );
  INV_X1 U14571 ( .A(n14566), .ZN(n14381) );
  NOR2_X1 U14572 ( .A1(n8662), .A2(n14560), .ZN(n14566) );
  NOR2_X1 U14573 ( .A1(n14567), .A2(n14568), .ZN(n14560) );
  NOR3_X1 U14574 ( .A1(n8992), .A2(n14569), .A3(n8988), .ZN(n14568) );
  NOR2_X1 U14575 ( .A1(n14377), .A2(n14376), .ZN(n14569) );
  INV_X1 U14576 ( .A(n14570), .ZN(n14567) );
  NAND2_X1 U14577 ( .A1(n14376), .A2(n14377), .ZN(n14570) );
  NAND2_X1 U14578 ( .A1(n14571), .A2(n14572), .ZN(n14377) );
  NAND2_X1 U14579 ( .A1(n14283), .A2(n14573), .ZN(n14572) );
  NAND2_X1 U14580 ( .A1(n14282), .A2(n14280), .ZN(n14573) );
  NOR2_X1 U14581 ( .A1(n8992), .A2(n8630), .ZN(n14283) );
  INV_X1 U14582 ( .A(n14574), .ZN(n14571) );
  NOR2_X1 U14583 ( .A1(n14280), .A2(n14282), .ZN(n14574) );
  NOR2_X1 U14584 ( .A1(n14575), .A2(n14576), .ZN(n14282) );
  NOR3_X1 U14585 ( .A1(n8986), .A2(n14577), .A3(n8992), .ZN(n14576) );
  INV_X1 U14586 ( .A(n14578), .ZN(n14577) );
  NAND2_X1 U14587 ( .A1(n14373), .A2(n14372), .ZN(n14578) );
  NOR2_X1 U14588 ( .A1(n14372), .A2(n14373), .ZN(n14575) );
  NOR2_X1 U14589 ( .A1(n14579), .A2(n14580), .ZN(n14373) );
  NOR3_X1 U14590 ( .A1(n8601), .A2(n14581), .A3(n8992), .ZN(n14580) );
  NOR2_X1 U14591 ( .A1(n14369), .A2(n14368), .ZN(n14581) );
  INV_X1 U14592 ( .A(n14582), .ZN(n14579) );
  NAND2_X1 U14593 ( .A1(n14368), .A2(n14369), .ZN(n14582) );
  NAND2_X1 U14594 ( .A1(n14583), .A2(n14584), .ZN(n14369) );
  NAND2_X1 U14595 ( .A1(n14366), .A2(n14585), .ZN(n14584) );
  INV_X1 U14596 ( .A(n14586), .ZN(n14585) );
  NOR2_X1 U14597 ( .A1(n14363), .A2(n14365), .ZN(n14586) );
  NOR2_X1 U14598 ( .A1(n8992), .A2(n8984), .ZN(n14366) );
  NAND2_X1 U14599 ( .A1(n14363), .A2(n14365), .ZN(n14583) );
  NAND2_X1 U14600 ( .A1(n14587), .A2(n14588), .ZN(n14365) );
  NAND2_X1 U14601 ( .A1(n14362), .A2(n14589), .ZN(n14588) );
  INV_X1 U14602 ( .A(n14590), .ZN(n14589) );
  NOR2_X1 U14603 ( .A1(n14361), .A2(n14360), .ZN(n14590) );
  NOR2_X1 U14604 ( .A1(n8992), .A2(n8572), .ZN(n14362) );
  NAND2_X1 U14605 ( .A1(n14360), .A2(n14361), .ZN(n14587) );
  NAND2_X1 U14606 ( .A1(n14591), .A2(n14592), .ZN(n14361) );
  NAND2_X1 U14607 ( .A1(n14358), .A2(n14593), .ZN(n14592) );
  INV_X1 U14608 ( .A(n14594), .ZN(n14593) );
  NOR2_X1 U14609 ( .A1(n14356), .A2(n14357), .ZN(n14594) );
  NOR2_X1 U14610 ( .A1(n8992), .A2(n8982), .ZN(n14358) );
  NAND2_X1 U14611 ( .A1(n14356), .A2(n14357), .ZN(n14591) );
  NAND2_X1 U14612 ( .A1(n14595), .A2(n14596), .ZN(n14357) );
  NAND2_X1 U14613 ( .A1(n14354), .A2(n14597), .ZN(n14596) );
  NAND2_X1 U14614 ( .A1(n14351), .A2(n14353), .ZN(n14597) );
  NOR2_X1 U14615 ( .A1(n8992), .A2(n8541), .ZN(n14354) );
  INV_X1 U14616 ( .A(n14598), .ZN(n14595) );
  NOR2_X1 U14617 ( .A1(n14353), .A2(n14351), .ZN(n14598) );
  XNOR2_X1 U14618 ( .A(n14599), .B(n14600), .ZN(n14351) );
  XNOR2_X1 U14619 ( .A(n14601), .B(n14602), .ZN(n14600) );
  NAND2_X1 U14620 ( .A1(n14603), .A2(n14604), .ZN(n14353) );
  NAND2_X1 U14621 ( .A1(n14313), .A2(n14605), .ZN(n14604) );
  NAND2_X1 U14622 ( .A1(n14316), .A2(n14315), .ZN(n14605) );
  XNOR2_X1 U14623 ( .A(n14606), .B(n14607), .ZN(n14313) );
  XOR2_X1 U14624 ( .A(n14608), .B(n14609), .Z(n14606) );
  INV_X1 U14625 ( .A(n14610), .ZN(n14603) );
  NOR2_X1 U14626 ( .A1(n14315), .A2(n14316), .ZN(n14610) );
  NOR2_X1 U14627 ( .A1(n9893), .A2(n8992), .ZN(n14316) );
  NAND2_X1 U14628 ( .A1(n14611), .A2(n14612), .ZN(n14315) );
  NAND2_X1 U14629 ( .A1(n14323), .A2(n14613), .ZN(n14612) );
  INV_X1 U14630 ( .A(n14614), .ZN(n14613) );
  NOR2_X1 U14631 ( .A1(n14321), .A2(n14322), .ZN(n14614) );
  NOR2_X1 U14632 ( .A1(n8992), .A2(n8512), .ZN(n14323) );
  NAND2_X1 U14633 ( .A1(n14321), .A2(n14322), .ZN(n14611) );
  NAND2_X1 U14634 ( .A1(n14615), .A2(n14616), .ZN(n14322) );
  NAND2_X1 U14635 ( .A1(n14349), .A2(n14617), .ZN(n14616) );
  INV_X1 U14636 ( .A(n14618), .ZN(n14617) );
  NOR2_X1 U14637 ( .A1(n14350), .A2(n14348), .ZN(n14618) );
  NOR2_X1 U14638 ( .A1(n8992), .A2(n8493), .ZN(n14349) );
  NAND2_X1 U14639 ( .A1(n14348), .A2(n14350), .ZN(n14615) );
  NAND2_X1 U14640 ( .A1(n14619), .A2(n14620), .ZN(n14350) );
  NAND2_X1 U14641 ( .A1(n14344), .A2(n14621), .ZN(n14620) );
  INV_X1 U14642 ( .A(n14622), .ZN(n14621) );
  NOR2_X1 U14643 ( .A1(n14345), .A2(n14346), .ZN(n14622) );
  NOR2_X1 U14644 ( .A1(n8992), .A2(n8473), .ZN(n14344) );
  NAND2_X1 U14645 ( .A1(n14346), .A2(n14345), .ZN(n14619) );
  NAND2_X1 U14646 ( .A1(n14623), .A2(n14624), .ZN(n14345) );
  NAND2_X1 U14647 ( .A1(b_8_), .A2(n14625), .ZN(n14624) );
  NAND2_X1 U14648 ( .A1(n8456), .A2(n14626), .ZN(n14625) );
  NAND2_X1 U14649 ( .A1(a_31_), .A2(n8781), .ZN(n14626) );
  NAND2_X1 U14650 ( .A1(b_9_), .A2(n14627), .ZN(n14623) );
  NAND2_X1 U14651 ( .A1(n8459), .A2(n14628), .ZN(n14627) );
  NAND2_X1 U14652 ( .A1(a_30_), .A2(n14458), .ZN(n14628) );
  NOR3_X1 U14653 ( .A1(n8992), .A2(n8979), .A3(n8781), .ZN(n14346) );
  XOR2_X1 U14654 ( .A(n14629), .B(n14630), .Z(n14348) );
  XOR2_X1 U14655 ( .A(n14631), .B(n14632), .Z(n14629) );
  XOR2_X1 U14656 ( .A(n14633), .B(n14634), .Z(n14321) );
  XOR2_X1 U14657 ( .A(n14635), .B(n14636), .Z(n14633) );
  XNOR2_X1 U14658 ( .A(n14637), .B(n14638), .ZN(n14356) );
  XNOR2_X1 U14659 ( .A(n14639), .B(n14640), .ZN(n14638) );
  XOR2_X1 U14660 ( .A(n14641), .B(n14642), .Z(n14360) );
  XOR2_X1 U14661 ( .A(n14643), .B(n14644), .Z(n14641) );
  XOR2_X1 U14662 ( .A(n14645), .B(n14646), .Z(n14363) );
  XOR2_X1 U14663 ( .A(n14647), .B(n14648), .Z(n14645) );
  XNOR2_X1 U14664 ( .A(n14649), .B(n14650), .ZN(n14368) );
  XNOR2_X1 U14665 ( .A(n14651), .B(n14652), .ZN(n14650) );
  XNOR2_X1 U14666 ( .A(n14653), .B(n14654), .ZN(n14372) );
  XOR2_X1 U14667 ( .A(n14655), .B(n14656), .Z(n14653) );
  XOR2_X1 U14668 ( .A(n14657), .B(n14658), .Z(n14280) );
  NAND2_X1 U14669 ( .A1(n14659), .A2(n14660), .ZN(n14657) );
  XOR2_X1 U14670 ( .A(n14661), .B(n14662), .Z(n14376) );
  XOR2_X1 U14671 ( .A(n14663), .B(n14664), .Z(n14661) );
  NOR2_X1 U14672 ( .A1(n8630), .A2(n8781), .ZN(n14664) );
  XOR2_X1 U14673 ( .A(n14665), .B(n14666), .Z(n14391) );
  XOR2_X1 U14674 ( .A(n14667), .B(n14668), .Z(n14665) );
  NOR2_X1 U14675 ( .A1(n8781), .A2(n8692), .ZN(n14668) );
  XOR2_X1 U14676 ( .A(n14669), .B(n14670), .Z(n14250) );
  XNOR2_X1 U14677 ( .A(n14671), .B(n14672), .ZN(n14670) );
  NAND2_X1 U14678 ( .A1(a_13_), .A2(b_9_), .ZN(n14672) );
  INV_X1 U14679 ( .A(n8763), .ZN(n14518) );
  NAND2_X1 U14680 ( .A1(a_10_), .A2(b_10_), .ZN(n8763) );
  XOR2_X1 U14681 ( .A(n14673), .B(n14674), .Z(n14415) );
  XNOR2_X1 U14682 ( .A(n14675), .B(n14676), .ZN(n14674) );
  NAND2_X1 U14683 ( .A1(a_7_), .A2(b_9_), .ZN(n14676) );
  XNOR2_X1 U14684 ( .A(n14677), .B(n14678), .ZN(n14419) );
  XNOR2_X1 U14685 ( .A(n14679), .B(n14680), .ZN(n14677) );
  NOR2_X1 U14686 ( .A1(n8781), .A2(n8994), .ZN(n14680) );
  XNOR2_X1 U14687 ( .A(n14681), .B(n14682), .ZN(n14423) );
  XNOR2_X1 U14688 ( .A(n14683), .B(n14684), .ZN(n14681) );
  NOR2_X1 U14689 ( .A1(n8781), .A2(n8848), .ZN(n14684) );
  XNOR2_X1 U14690 ( .A(n14685), .B(n14686), .ZN(n14427) );
  XNOR2_X1 U14691 ( .A(n14687), .B(n14688), .ZN(n14685) );
  NOR2_X1 U14692 ( .A1(n8781), .A2(n8996), .ZN(n14688) );
  XNOR2_X1 U14693 ( .A(n14689), .B(n14690), .ZN(n14431) );
  XNOR2_X1 U14694 ( .A(n14691), .B(n14692), .ZN(n14689) );
  NOR2_X1 U14695 ( .A1(n8781), .A2(n8877), .ZN(n14692) );
  XNOR2_X1 U14696 ( .A(n14693), .B(n14694), .ZN(n14435) );
  XNOR2_X1 U14697 ( .A(n14695), .B(n14696), .ZN(n14693) );
  NOR2_X1 U14698 ( .A1(n8781), .A2(n8998), .ZN(n14696) );
  XOR2_X1 U14699 ( .A(n14697), .B(n14698), .Z(n14438) );
  XNOR2_X1 U14700 ( .A(n14699), .B(n14700), .ZN(n14698) );
  NAND2_X1 U14701 ( .A1(a_1_), .A2(b_9_), .ZN(n14700) );
  XNOR2_X1 U14702 ( .A(n14701), .B(n14454), .ZN(n8428) );
  XNOR2_X1 U14703 ( .A(n14702), .B(n14703), .ZN(n14454) );
  XOR2_X1 U14704 ( .A(n14704), .B(n14705), .Z(n14702) );
  NOR2_X1 U14705 ( .A1(n14458), .A2(n9731), .ZN(n14705) );
  XNOR2_X1 U14706 ( .A(n14455), .B(n14452), .ZN(n14701) );
  NOR2_X1 U14707 ( .A1(n9471), .A2(n8781), .ZN(n14452) );
  NOR2_X1 U14708 ( .A1(n14706), .A2(n14707), .ZN(n14455) );
  NOR3_X1 U14709 ( .A1(n8781), .A2(n14708), .A3(n9731), .ZN(n14707) );
  INV_X1 U14710 ( .A(n14709), .ZN(n14708) );
  NAND2_X1 U14711 ( .A1(n14699), .A2(n14697), .ZN(n14709) );
  NOR2_X1 U14712 ( .A1(n14697), .A2(n14699), .ZN(n14706) );
  NOR2_X1 U14713 ( .A1(n14710), .A2(n14711), .ZN(n14699) );
  INV_X1 U14714 ( .A(n14712), .ZN(n14711) );
  NAND3_X1 U14715 ( .A1(b_9_), .A2(n14713), .A3(a_2_), .ZN(n14712) );
  NAND2_X1 U14716 ( .A1(n14695), .A2(n14694), .ZN(n14713) );
  NOR2_X1 U14717 ( .A1(n14694), .A2(n14695), .ZN(n14710) );
  NOR2_X1 U14718 ( .A1(n14714), .A2(n14715), .ZN(n14695) );
  INV_X1 U14719 ( .A(n14716), .ZN(n14715) );
  NAND3_X1 U14720 ( .A1(b_9_), .A2(n14717), .A3(a_3_), .ZN(n14716) );
  NAND2_X1 U14721 ( .A1(n14691), .A2(n14690), .ZN(n14717) );
  NOR2_X1 U14722 ( .A1(n14690), .A2(n14691), .ZN(n14714) );
  NOR2_X1 U14723 ( .A1(n14718), .A2(n14719), .ZN(n14691) );
  INV_X1 U14724 ( .A(n14720), .ZN(n14719) );
  NAND3_X1 U14725 ( .A1(b_9_), .A2(n14721), .A3(a_4_), .ZN(n14720) );
  NAND2_X1 U14726 ( .A1(n14687), .A2(n14686), .ZN(n14721) );
  NOR2_X1 U14727 ( .A1(n14686), .A2(n14687), .ZN(n14718) );
  NOR2_X1 U14728 ( .A1(n14722), .A2(n14723), .ZN(n14687) );
  INV_X1 U14729 ( .A(n14724), .ZN(n14723) );
  NAND3_X1 U14730 ( .A1(b_9_), .A2(n14725), .A3(a_5_), .ZN(n14724) );
  NAND2_X1 U14731 ( .A1(n14683), .A2(n14682), .ZN(n14725) );
  NOR2_X1 U14732 ( .A1(n14682), .A2(n14683), .ZN(n14722) );
  NOR2_X1 U14733 ( .A1(n14726), .A2(n14727), .ZN(n14683) );
  INV_X1 U14734 ( .A(n14728), .ZN(n14727) );
  NAND3_X1 U14735 ( .A1(b_9_), .A2(n14729), .A3(a_6_), .ZN(n14728) );
  NAND2_X1 U14736 ( .A1(n14679), .A2(n14678), .ZN(n14729) );
  NOR2_X1 U14737 ( .A1(n14678), .A2(n14679), .ZN(n14726) );
  NOR2_X1 U14738 ( .A1(n14730), .A2(n14731), .ZN(n14679) );
  NOR3_X1 U14739 ( .A1(n8781), .A2(n14732), .A3(n8817), .ZN(n14731) );
  INV_X1 U14740 ( .A(n14733), .ZN(n14732) );
  NAND2_X1 U14741 ( .A1(n14675), .A2(n14673), .ZN(n14733) );
  NOR2_X1 U14742 ( .A1(n14673), .A2(n14675), .ZN(n14730) );
  NOR2_X1 U14743 ( .A1(n14734), .A2(n14735), .ZN(n14675) );
  INV_X1 U14744 ( .A(n14736), .ZN(n14735) );
  NAND3_X1 U14745 ( .A1(b_9_), .A2(n14737), .A3(a_8_), .ZN(n14736) );
  NAND2_X1 U14746 ( .A1(n14491), .A2(n14493), .ZN(n14737) );
  NOR2_X1 U14747 ( .A1(n14493), .A2(n14491), .ZN(n14734) );
  XNOR2_X1 U14748 ( .A(n14738), .B(n14739), .ZN(n14491) );
  XOR2_X1 U14749 ( .A(n14740), .B(n14741), .Z(n14739) );
  NAND2_X1 U14750 ( .A1(n14742), .A2(n14743), .ZN(n14493) );
  NAND2_X1 U14751 ( .A1(n14498), .A2(n14744), .ZN(n14743) );
  NAND2_X1 U14752 ( .A1(n8776), .A2(n14500), .ZN(n14744) );
  XOR2_X1 U14753 ( .A(n14745), .B(n14746), .Z(n14498) );
  XNOR2_X1 U14754 ( .A(n14747), .B(n14748), .ZN(n14745) );
  INV_X1 U14755 ( .A(n14749), .ZN(n14742) );
  NOR2_X1 U14756 ( .A1(n14500), .A2(n8776), .ZN(n14749) );
  NOR2_X1 U14757 ( .A1(n8779), .A2(n8781), .ZN(n8776) );
  NAND2_X1 U14758 ( .A1(n14750), .A2(n14751), .ZN(n14500) );
  NAND3_X1 U14759 ( .A1(b_9_), .A2(n14752), .A3(a_10_), .ZN(n14751) );
  INV_X1 U14760 ( .A(n14753), .ZN(n14752) );
  NOR2_X1 U14761 ( .A1(n14506), .A2(n14508), .ZN(n14753) );
  NAND2_X1 U14762 ( .A1(n14506), .A2(n14508), .ZN(n14750) );
  NAND2_X1 U14763 ( .A1(n14754), .A2(n14755), .ZN(n14508) );
  NAND3_X1 U14764 ( .A1(b_9_), .A2(n14756), .A3(a_11_), .ZN(n14755) );
  NAND2_X1 U14765 ( .A1(n14516), .A2(n14514), .ZN(n14756) );
  INV_X1 U14766 ( .A(n14757), .ZN(n14754) );
  NOR2_X1 U14767 ( .A1(n14514), .A2(n14516), .ZN(n14757) );
  NOR2_X1 U14768 ( .A1(n14758), .A2(n14759), .ZN(n14516) );
  INV_X1 U14769 ( .A(n14760), .ZN(n14759) );
  NAND3_X1 U14770 ( .A1(b_9_), .A2(n14761), .A3(a_12_), .ZN(n14760) );
  NAND2_X1 U14771 ( .A1(n14524), .A2(n14523), .ZN(n14761) );
  NOR2_X1 U14772 ( .A1(n14523), .A2(n14524), .ZN(n14758) );
  NOR2_X1 U14773 ( .A1(n14762), .A2(n14763), .ZN(n14524) );
  NOR3_X1 U14774 ( .A1(n8781), .A2(n14764), .A3(n8721), .ZN(n14763) );
  INV_X1 U14775 ( .A(n14765), .ZN(n14764) );
  NAND2_X1 U14776 ( .A1(n14671), .A2(n14669), .ZN(n14765) );
  NOR2_X1 U14777 ( .A1(n14669), .A2(n14671), .ZN(n14762) );
  NOR2_X1 U14778 ( .A1(n14766), .A2(n14767), .ZN(n14671) );
  INV_X1 U14779 ( .A(n14768), .ZN(n14767) );
  NAND3_X1 U14780 ( .A1(b_9_), .A2(n14769), .A3(a_14_), .ZN(n14768) );
  NAND2_X1 U14781 ( .A1(n14536), .A2(n14535), .ZN(n14769) );
  NOR2_X1 U14782 ( .A1(n14535), .A2(n14536), .ZN(n14766) );
  NOR2_X1 U14783 ( .A1(n14770), .A2(n14771), .ZN(n14536) );
  NOR3_X1 U14784 ( .A1(n8781), .A2(n14772), .A3(n8692), .ZN(n14771) );
  NOR2_X1 U14785 ( .A1(n14666), .A2(n14667), .ZN(n14772) );
  INV_X1 U14786 ( .A(n14773), .ZN(n14770) );
  NAND2_X1 U14787 ( .A1(n14666), .A2(n14667), .ZN(n14773) );
  NAND2_X1 U14788 ( .A1(n14774), .A2(n14775), .ZN(n14667) );
  NAND3_X1 U14789 ( .A1(b_9_), .A2(n14776), .A3(a_16_), .ZN(n14775) );
  NAND2_X1 U14790 ( .A1(n14549), .A2(n14547), .ZN(n14776) );
  INV_X1 U14791 ( .A(n14777), .ZN(n14774) );
  NOR2_X1 U14792 ( .A1(n14547), .A2(n14549), .ZN(n14777) );
  NOR2_X1 U14793 ( .A1(n14778), .A2(n14779), .ZN(n14549) );
  INV_X1 U14794 ( .A(n14780), .ZN(n14779) );
  NAND3_X1 U14795 ( .A1(b_9_), .A2(n14781), .A3(a_17_), .ZN(n14780) );
  NAND2_X1 U14796 ( .A1(n14557), .A2(n14556), .ZN(n14781) );
  NOR2_X1 U14797 ( .A1(n14556), .A2(n14557), .ZN(n14778) );
  NOR2_X1 U14798 ( .A1(n14782), .A2(n14783), .ZN(n14557) );
  NOR3_X1 U14799 ( .A1(n8781), .A2(n14784), .A3(n8988), .ZN(n14783) );
  NOR2_X1 U14800 ( .A1(n14564), .A2(n14562), .ZN(n14784) );
  INV_X1 U14801 ( .A(n14785), .ZN(n14782) );
  NAND2_X1 U14802 ( .A1(n14562), .A2(n14564), .ZN(n14785) );
  NAND2_X1 U14803 ( .A1(n14786), .A2(n14787), .ZN(n14564) );
  NAND3_X1 U14804 ( .A1(a_19_), .A2(n14788), .A3(b_9_), .ZN(n14787) );
  INV_X1 U14805 ( .A(n14789), .ZN(n14788) );
  NOR2_X1 U14806 ( .A1(n14662), .A2(n14663), .ZN(n14789) );
  NAND2_X1 U14807 ( .A1(n14662), .A2(n14663), .ZN(n14786) );
  NAND2_X1 U14808 ( .A1(n14659), .A2(n14790), .ZN(n14663) );
  NAND2_X1 U14809 ( .A1(n14658), .A2(n14660), .ZN(n14790) );
  NAND2_X1 U14810 ( .A1(n14791), .A2(n14792), .ZN(n14660) );
  NAND2_X1 U14811 ( .A1(b_9_), .A2(a_20_), .ZN(n14792) );
  INV_X1 U14812 ( .A(n14793), .ZN(n14791) );
  XNOR2_X1 U14813 ( .A(n14794), .B(n14795), .ZN(n14658) );
  XOR2_X1 U14814 ( .A(n14796), .B(n14797), .Z(n14795) );
  NAND2_X1 U14815 ( .A1(a_20_), .A2(n14793), .ZN(n14659) );
  NAND2_X1 U14816 ( .A1(n14798), .A2(n14799), .ZN(n14793) );
  NAND2_X1 U14817 ( .A1(n14656), .A2(n14800), .ZN(n14799) );
  INV_X1 U14818 ( .A(n14801), .ZN(n14800) );
  NOR2_X1 U14819 ( .A1(n14654), .A2(n14655), .ZN(n14801) );
  NOR2_X1 U14820 ( .A1(n8781), .A2(n8601), .ZN(n14656) );
  NAND2_X1 U14821 ( .A1(n14654), .A2(n14655), .ZN(n14798) );
  NAND2_X1 U14822 ( .A1(n14802), .A2(n14803), .ZN(n14655) );
  NAND2_X1 U14823 ( .A1(n14652), .A2(n14804), .ZN(n14803) );
  INV_X1 U14824 ( .A(n14805), .ZN(n14804) );
  NOR2_X1 U14825 ( .A1(n14649), .A2(n14651), .ZN(n14805) );
  NOR2_X1 U14826 ( .A1(n8781), .A2(n8984), .ZN(n14652) );
  NAND2_X1 U14827 ( .A1(n14649), .A2(n14651), .ZN(n14802) );
  NAND2_X1 U14828 ( .A1(n14806), .A2(n14807), .ZN(n14651) );
  NAND2_X1 U14829 ( .A1(n14648), .A2(n14808), .ZN(n14807) );
  INV_X1 U14830 ( .A(n14809), .ZN(n14808) );
  NOR2_X1 U14831 ( .A1(n14647), .A2(n14646), .ZN(n14809) );
  NOR2_X1 U14832 ( .A1(n8781), .A2(n8572), .ZN(n14648) );
  NAND2_X1 U14833 ( .A1(n14646), .A2(n14647), .ZN(n14806) );
  NAND2_X1 U14834 ( .A1(n14810), .A2(n14811), .ZN(n14647) );
  NAND2_X1 U14835 ( .A1(n14644), .A2(n14812), .ZN(n14811) );
  INV_X1 U14836 ( .A(n14813), .ZN(n14812) );
  NOR2_X1 U14837 ( .A1(n14642), .A2(n14643), .ZN(n14813) );
  NOR2_X1 U14838 ( .A1(n8781), .A2(n8982), .ZN(n14644) );
  NAND2_X1 U14839 ( .A1(n14642), .A2(n14643), .ZN(n14810) );
  NAND2_X1 U14840 ( .A1(n14814), .A2(n14815), .ZN(n14643) );
  NAND2_X1 U14841 ( .A1(n14640), .A2(n14816), .ZN(n14815) );
  NAND2_X1 U14842 ( .A1(n14637), .A2(n14639), .ZN(n14816) );
  NOR2_X1 U14843 ( .A1(n8781), .A2(n8541), .ZN(n14640) );
  INV_X1 U14844 ( .A(n14817), .ZN(n14814) );
  NOR2_X1 U14845 ( .A1(n14639), .A2(n14637), .ZN(n14817) );
  XNOR2_X1 U14846 ( .A(n14818), .B(n14819), .ZN(n14637) );
  XNOR2_X1 U14847 ( .A(n14820), .B(n14821), .ZN(n14819) );
  NAND2_X1 U14848 ( .A1(n14822), .A2(n14823), .ZN(n14639) );
  NAND2_X1 U14849 ( .A1(n14599), .A2(n14824), .ZN(n14823) );
  NAND2_X1 U14850 ( .A1(n14602), .A2(n14601), .ZN(n14824) );
  XNOR2_X1 U14851 ( .A(n14825), .B(n14826), .ZN(n14599) );
  XOR2_X1 U14852 ( .A(n14827), .B(n14828), .Z(n14825) );
  INV_X1 U14853 ( .A(n14829), .ZN(n14822) );
  NOR2_X1 U14854 ( .A1(n14601), .A2(n14602), .ZN(n14829) );
  NOR2_X1 U14855 ( .A1(n9893), .A2(n8781), .ZN(n14602) );
  NAND2_X1 U14856 ( .A1(n14830), .A2(n14831), .ZN(n14601) );
  NAND2_X1 U14857 ( .A1(n14609), .A2(n14832), .ZN(n14831) );
  INV_X1 U14858 ( .A(n14833), .ZN(n14832) );
  NOR2_X1 U14859 ( .A1(n14607), .A2(n14608), .ZN(n14833) );
  NOR2_X1 U14860 ( .A1(n8781), .A2(n8512), .ZN(n14609) );
  NAND2_X1 U14861 ( .A1(n14607), .A2(n14608), .ZN(n14830) );
  NAND2_X1 U14862 ( .A1(n14834), .A2(n14835), .ZN(n14608) );
  NAND2_X1 U14863 ( .A1(n14635), .A2(n14836), .ZN(n14835) );
  INV_X1 U14864 ( .A(n14837), .ZN(n14836) );
  NOR2_X1 U14865 ( .A1(n14636), .A2(n14634), .ZN(n14837) );
  NOR2_X1 U14866 ( .A1(n8781), .A2(n8493), .ZN(n14635) );
  NAND2_X1 U14867 ( .A1(n14634), .A2(n14636), .ZN(n14834) );
  NAND2_X1 U14868 ( .A1(n14838), .A2(n14839), .ZN(n14636) );
  NAND2_X1 U14869 ( .A1(n14630), .A2(n14840), .ZN(n14839) );
  INV_X1 U14870 ( .A(n14841), .ZN(n14840) );
  NOR2_X1 U14871 ( .A1(n14631), .A2(n14632), .ZN(n14841) );
  NOR2_X1 U14872 ( .A1(n8781), .A2(n8473), .ZN(n14630) );
  NAND2_X1 U14873 ( .A1(n14632), .A2(n14631), .ZN(n14838) );
  NAND2_X1 U14874 ( .A1(n14842), .A2(n14843), .ZN(n14631) );
  NAND2_X1 U14875 ( .A1(b_7_), .A2(n14844), .ZN(n14843) );
  NAND2_X1 U14876 ( .A1(n8456), .A2(n14845), .ZN(n14844) );
  NAND2_X1 U14877 ( .A1(a_31_), .A2(n14458), .ZN(n14845) );
  NAND2_X1 U14878 ( .A1(b_8_), .A2(n14846), .ZN(n14842) );
  NAND2_X1 U14879 ( .A1(n8459), .A2(n14847), .ZN(n14846) );
  NAND2_X1 U14880 ( .A1(a_30_), .A2(n8819), .ZN(n14847) );
  NOR3_X1 U14881 ( .A1(n8781), .A2(n8979), .A3(n14458), .ZN(n14632) );
  XOR2_X1 U14882 ( .A(n14848), .B(n14849), .Z(n14634) );
  XOR2_X1 U14883 ( .A(n14850), .B(n14851), .Z(n14848) );
  XOR2_X1 U14884 ( .A(n14852), .B(n14853), .Z(n14607) );
  XOR2_X1 U14885 ( .A(n14854), .B(n14855), .Z(n14852) );
  XNOR2_X1 U14886 ( .A(n14856), .B(n14857), .ZN(n14642) );
  XNOR2_X1 U14887 ( .A(n14858), .B(n14859), .ZN(n14857) );
  XOR2_X1 U14888 ( .A(n14860), .B(n14861), .Z(n14646) );
  XOR2_X1 U14889 ( .A(n14862), .B(n14863), .Z(n14860) );
  XOR2_X1 U14890 ( .A(n14864), .B(n14865), .Z(n14649) );
  XOR2_X1 U14891 ( .A(n14866), .B(n14867), .Z(n14864) );
  XNOR2_X1 U14892 ( .A(n14868), .B(n14869), .ZN(n14654) );
  XNOR2_X1 U14893 ( .A(n14870), .B(n14871), .ZN(n14869) );
  XNOR2_X1 U14894 ( .A(n14872), .B(n14873), .ZN(n14662) );
  XNOR2_X1 U14895 ( .A(n14874), .B(n14875), .ZN(n14872) );
  XOR2_X1 U14896 ( .A(n14876), .B(n14877), .Z(n14562) );
  XOR2_X1 U14897 ( .A(n14878), .B(n14879), .Z(n14877) );
  XOR2_X1 U14898 ( .A(n14880), .B(n14881), .Z(n14556) );
  XOR2_X1 U14899 ( .A(n14882), .B(n14883), .Z(n14880) );
  XOR2_X1 U14900 ( .A(n14884), .B(n14885), .Z(n14547) );
  XNOR2_X1 U14901 ( .A(n14886), .B(n14887), .ZN(n14885) );
  XOR2_X1 U14902 ( .A(n14888), .B(n14889), .Z(n14666) );
  XNOR2_X1 U14903 ( .A(n14890), .B(n14891), .ZN(n14889) );
  XNOR2_X1 U14904 ( .A(n14892), .B(n14893), .ZN(n14535) );
  XOR2_X1 U14905 ( .A(n14894), .B(n14895), .Z(n14893) );
  XNOR2_X1 U14906 ( .A(n14896), .B(n14897), .ZN(n14669) );
  XNOR2_X1 U14907 ( .A(n14898), .B(n14899), .ZN(n14897) );
  XNOR2_X1 U14908 ( .A(n14900), .B(n14901), .ZN(n14523) );
  XOR2_X1 U14909 ( .A(n14902), .B(n14903), .Z(n14901) );
  XNOR2_X1 U14910 ( .A(n14904), .B(n14905), .ZN(n14514) );
  XOR2_X1 U14911 ( .A(n14906), .B(n14907), .Z(n14904) );
  XNOR2_X1 U14912 ( .A(n14908), .B(n14909), .ZN(n14506) );
  XNOR2_X1 U14913 ( .A(n14910), .B(n14911), .ZN(n14908) );
  XNOR2_X1 U14914 ( .A(n14912), .B(n14913), .ZN(n14673) );
  XNOR2_X1 U14915 ( .A(n14914), .B(n8793), .ZN(n14913) );
  XNOR2_X1 U14916 ( .A(n14915), .B(n14916), .ZN(n14678) );
  XOR2_X1 U14917 ( .A(n14917), .B(n14918), .Z(n14916) );
  XOR2_X1 U14918 ( .A(n14919), .B(n14920), .Z(n14682) );
  XOR2_X1 U14919 ( .A(n14921), .B(n14922), .Z(n14920) );
  XOR2_X1 U14920 ( .A(n14923), .B(n14924), .Z(n14686) );
  XNOR2_X1 U14921 ( .A(n14925), .B(n14926), .ZN(n14923) );
  XNOR2_X1 U14922 ( .A(n14927), .B(n14928), .ZN(n14690) );
  XNOR2_X1 U14923 ( .A(n14929), .B(n14930), .ZN(n14927) );
  XOR2_X1 U14924 ( .A(n14931), .B(n14932), .Z(n14694) );
  XNOR2_X1 U14925 ( .A(n14933), .B(n14934), .ZN(n14931) );
  XNOR2_X1 U14926 ( .A(n14935), .B(n14936), .ZN(n14697) );
  XOR2_X1 U14927 ( .A(n14937), .B(n14938), .Z(n14935) );
  XOR2_X1 U14928 ( .A(n8441), .B(n8440), .Z(n8431) );
  INV_X1 U14929 ( .A(n8436), .ZN(n9145) );
  NAND3_X1 U14930 ( .A1(n8440), .A2(n8441), .A3(n14939), .ZN(n8436) );
  INV_X1 U14931 ( .A(n8439), .ZN(n14939) );
  NAND2_X1 U14932 ( .A1(n9144), .A2(n14940), .ZN(n8439) );
  NAND2_X1 U14933 ( .A1(n14941), .A2(n14942), .ZN(n14940) );
  INV_X1 U14934 ( .A(n14943), .ZN(n9144) );
  NOR2_X1 U14935 ( .A1(n14941), .A2(n14942), .ZN(n14943) );
  NOR2_X1 U14936 ( .A1(n14944), .A2(n14945), .ZN(n14942) );
  INV_X1 U14937 ( .A(n14946), .ZN(n14945) );
  NAND2_X1 U14938 ( .A1(n14947), .A2(n14948), .ZN(n14946) );
  NAND2_X1 U14939 ( .A1(n14949), .A2(n14950), .ZN(n14948) );
  NOR2_X1 U14940 ( .A1(n14950), .A2(n14949), .ZN(n14944) );
  XOR2_X1 U14941 ( .A(n14951), .B(n14952), .Z(n14941) );
  XNOR2_X1 U14942 ( .A(n14953), .B(n14954), .ZN(n14951) );
  NOR2_X1 U14943 ( .A1(n8993), .A2(n9471), .ZN(n14954) );
  NAND2_X1 U14944 ( .A1(n14955), .A2(n14956), .ZN(n8441) );
  NAND3_X1 U14945 ( .A1(b_8_), .A2(n14957), .A3(a_0_), .ZN(n14956) );
  NAND2_X1 U14946 ( .A1(n14446), .A2(n14456), .ZN(n14957) );
  INV_X1 U14947 ( .A(n14958), .ZN(n14955) );
  NOR2_X1 U14948 ( .A1(n14446), .A2(n14456), .ZN(n14958) );
  NOR2_X1 U14949 ( .A1(n14959), .A2(n14960), .ZN(n14456) );
  NOR3_X1 U14950 ( .A1(n14458), .A2(n14961), .A3(n9731), .ZN(n14960) );
  NOR2_X1 U14951 ( .A1(n14704), .A2(n14703), .ZN(n14961) );
  INV_X1 U14952 ( .A(n14962), .ZN(n14959) );
  NAND2_X1 U14953 ( .A1(n14703), .A2(n14704), .ZN(n14962) );
  NAND2_X1 U14954 ( .A1(n14963), .A2(n14964), .ZN(n14704) );
  NAND2_X1 U14955 ( .A1(n14938), .A2(n14965), .ZN(n14964) );
  INV_X1 U14956 ( .A(n14966), .ZN(n14965) );
  NOR2_X1 U14957 ( .A1(n14936), .A2(n14937), .ZN(n14966) );
  NOR2_X1 U14958 ( .A1(n8998), .A2(n14458), .ZN(n14938) );
  NAND2_X1 U14959 ( .A1(n14936), .A2(n14937), .ZN(n14963) );
  NAND2_X1 U14960 ( .A1(n14967), .A2(n14968), .ZN(n14937) );
  NAND2_X1 U14961 ( .A1(n14934), .A2(n14969), .ZN(n14968) );
  NAND2_X1 U14962 ( .A1(n14932), .A2(n14933), .ZN(n14969) );
  NOR2_X1 U14963 ( .A1(n8877), .A2(n14458), .ZN(n14934) );
  INV_X1 U14964 ( .A(n14970), .ZN(n14967) );
  NOR2_X1 U14965 ( .A1(n14932), .A2(n14933), .ZN(n14970) );
  NOR2_X1 U14966 ( .A1(n14971), .A2(n14972), .ZN(n14933) );
  NOR2_X1 U14967 ( .A1(n14929), .A2(n14973), .ZN(n14972) );
  NOR2_X1 U14968 ( .A1(n14928), .A2(n14930), .ZN(n14973) );
  NAND2_X1 U14969 ( .A1(a_4_), .A2(b_8_), .ZN(n14929) );
  INV_X1 U14970 ( .A(n14974), .ZN(n14971) );
  NAND2_X1 U14971 ( .A1(n14928), .A2(n14930), .ZN(n14974) );
  NAND2_X1 U14972 ( .A1(n14975), .A2(n14976), .ZN(n14930) );
  NAND2_X1 U14973 ( .A1(n14926), .A2(n14977), .ZN(n14976) );
  NAND2_X1 U14974 ( .A1(n14924), .A2(n14925), .ZN(n14977) );
  NOR2_X1 U14975 ( .A1(n8848), .A2(n14458), .ZN(n14926) );
  INV_X1 U14976 ( .A(n14978), .ZN(n14975) );
  NOR2_X1 U14977 ( .A1(n14924), .A2(n14925), .ZN(n14978) );
  NOR2_X1 U14978 ( .A1(n14979), .A2(n14980), .ZN(n14925) );
  NOR2_X1 U14979 ( .A1(n14922), .A2(n14981), .ZN(n14980) );
  NOR2_X1 U14980 ( .A1(n14919), .A2(n14921), .ZN(n14981) );
  NAND2_X1 U14981 ( .A1(a_6_), .A2(b_8_), .ZN(n14922) );
  INV_X1 U14982 ( .A(n14982), .ZN(n14979) );
  NAND2_X1 U14983 ( .A1(n14919), .A2(n14921), .ZN(n14982) );
  NAND2_X1 U14984 ( .A1(n14983), .A2(n14984), .ZN(n14921) );
  NAND2_X1 U14985 ( .A1(n14918), .A2(n14985), .ZN(n14984) );
  INV_X1 U14986 ( .A(n14986), .ZN(n14985) );
  NOR2_X1 U14987 ( .A1(n14915), .A2(n14917), .ZN(n14986) );
  NOR2_X1 U14988 ( .A1(n8817), .A2(n14458), .ZN(n14918) );
  NAND2_X1 U14989 ( .A1(n14915), .A2(n14917), .ZN(n14983) );
  NOR2_X1 U14990 ( .A1(n14987), .A2(n14988), .ZN(n14917) );
  INV_X1 U14991 ( .A(n14989), .ZN(n14988) );
  NAND2_X1 U14992 ( .A1(n14912), .A2(n14990), .ZN(n14989) );
  NAND2_X1 U14993 ( .A1(n8793), .A2(n14914), .ZN(n14990) );
  XOR2_X1 U14994 ( .A(n14991), .B(n14992), .Z(n14912) );
  XNOR2_X1 U14995 ( .A(n14993), .B(n14994), .ZN(n14991) );
  NOR2_X1 U14996 ( .A1(n8819), .A2(n8779), .ZN(n14994) );
  NOR2_X1 U14997 ( .A1(n14914), .A2(n8793), .ZN(n14987) );
  NOR2_X1 U14998 ( .A1(n10513), .A2(n14458), .ZN(n8793) );
  NAND2_X1 U14999 ( .A1(n14995), .A2(n14996), .ZN(n14914) );
  NAND2_X1 U15000 ( .A1(n14741), .A2(n14997), .ZN(n14996) );
  NAND2_X1 U15001 ( .A1(n14740), .A2(n14738), .ZN(n14997) );
  NOR2_X1 U15002 ( .A1(n8779), .A2(n14458), .ZN(n14741) );
  INV_X1 U15003 ( .A(n14998), .ZN(n14995) );
  NOR2_X1 U15004 ( .A1(n14738), .A2(n14740), .ZN(n14998) );
  NOR2_X1 U15005 ( .A1(n14999), .A2(n15000), .ZN(n14740) );
  INV_X1 U15006 ( .A(n15001), .ZN(n15000) );
  NAND2_X1 U15007 ( .A1(n14748), .A2(n15002), .ZN(n15001) );
  NAND2_X1 U15008 ( .A1(n14747), .A2(n14746), .ZN(n15002) );
  NOR2_X1 U15009 ( .A1(n8769), .A2(n14458), .ZN(n14748) );
  NOR2_X1 U15010 ( .A1(n14746), .A2(n14747), .ZN(n14999) );
  NOR2_X1 U15011 ( .A1(n15003), .A2(n15004), .ZN(n14747) );
  INV_X1 U15012 ( .A(n15005), .ZN(n15004) );
  NAND2_X1 U15013 ( .A1(n14911), .A2(n15006), .ZN(n15005) );
  NAND2_X1 U15014 ( .A1(n14910), .A2(n14909), .ZN(n15006) );
  NOR2_X1 U15015 ( .A1(n8749), .A2(n14458), .ZN(n14911) );
  NOR2_X1 U15016 ( .A1(n14909), .A2(n14910), .ZN(n15003) );
  INV_X1 U15017 ( .A(n15007), .ZN(n14910) );
  NAND2_X1 U15018 ( .A1(n15008), .A2(n15009), .ZN(n15007) );
  NAND2_X1 U15019 ( .A1(n14907), .A2(n15010), .ZN(n15009) );
  INV_X1 U15020 ( .A(n15011), .ZN(n15010) );
  NOR2_X1 U15021 ( .A1(n14905), .A2(n14906), .ZN(n15011) );
  NOR2_X1 U15022 ( .A1(n8739), .A2(n14458), .ZN(n14907) );
  NAND2_X1 U15023 ( .A1(n14905), .A2(n14906), .ZN(n15008) );
  NAND2_X1 U15024 ( .A1(n15012), .A2(n15013), .ZN(n14906) );
  NAND2_X1 U15025 ( .A1(n14903), .A2(n15014), .ZN(n15013) );
  INV_X1 U15026 ( .A(n15015), .ZN(n15014) );
  NOR2_X1 U15027 ( .A1(n14900), .A2(n14902), .ZN(n15015) );
  NOR2_X1 U15028 ( .A1(n8721), .A2(n14458), .ZN(n14903) );
  NAND2_X1 U15029 ( .A1(n14900), .A2(n14902), .ZN(n15012) );
  NOR2_X1 U15030 ( .A1(n15016), .A2(n15017), .ZN(n14902) );
  INV_X1 U15031 ( .A(n15018), .ZN(n15017) );
  NAND2_X1 U15032 ( .A1(n14896), .A2(n15019), .ZN(n15018) );
  NAND2_X1 U15033 ( .A1(n14899), .A2(n14898), .ZN(n15019) );
  XOR2_X1 U15034 ( .A(n15020), .B(n15021), .Z(n14896) );
  XOR2_X1 U15035 ( .A(n15022), .B(n15023), .Z(n15021) );
  NAND2_X1 U15036 ( .A1(a_15_), .A2(b_7_), .ZN(n15023) );
  NOR2_X1 U15037 ( .A1(n14898), .A2(n14899), .ZN(n15016) );
  NOR2_X1 U15038 ( .A1(n8991), .A2(n14458), .ZN(n14899) );
  NAND2_X1 U15039 ( .A1(n15024), .A2(n15025), .ZN(n14898) );
  NAND2_X1 U15040 ( .A1(n14895), .A2(n15026), .ZN(n15025) );
  INV_X1 U15041 ( .A(n15027), .ZN(n15026) );
  NOR2_X1 U15042 ( .A1(n14892), .A2(n14894), .ZN(n15027) );
  NOR2_X1 U15043 ( .A1(n8692), .A2(n14458), .ZN(n14895) );
  NAND2_X1 U15044 ( .A1(n14892), .A2(n14894), .ZN(n15024) );
  NOR2_X1 U15045 ( .A1(n15028), .A2(n15029), .ZN(n14894) );
  INV_X1 U15046 ( .A(n15030), .ZN(n15029) );
  NAND2_X1 U15047 ( .A1(n14888), .A2(n15031), .ZN(n15030) );
  NAND2_X1 U15048 ( .A1(n14891), .A2(n14890), .ZN(n15031) );
  XNOR2_X1 U15049 ( .A(n15032), .B(n15033), .ZN(n14888) );
  XNOR2_X1 U15050 ( .A(n15034), .B(n15035), .ZN(n15033) );
  NAND2_X1 U15051 ( .A1(a_17_), .A2(b_7_), .ZN(n15035) );
  NOR2_X1 U15052 ( .A1(n14890), .A2(n14891), .ZN(n15028) );
  NOR2_X1 U15053 ( .A1(n8680), .A2(n14458), .ZN(n14891) );
  NAND2_X1 U15054 ( .A1(n15036), .A2(n15037), .ZN(n14890) );
  NAND2_X1 U15055 ( .A1(n14887), .A2(n15038), .ZN(n15037) );
  NAND2_X1 U15056 ( .A1(n14884), .A2(n14886), .ZN(n15038) );
  NOR2_X1 U15057 ( .A1(n8662), .A2(n14458), .ZN(n14887) );
  INV_X1 U15058 ( .A(n15039), .ZN(n15036) );
  NOR2_X1 U15059 ( .A1(n14884), .A2(n14886), .ZN(n15039) );
  NAND2_X1 U15060 ( .A1(n15040), .A2(n15041), .ZN(n14886) );
  NAND2_X1 U15061 ( .A1(n14881), .A2(n15042), .ZN(n15041) );
  NAND2_X1 U15062 ( .A1(n14883), .A2(n14882), .ZN(n15042) );
  XOR2_X1 U15063 ( .A(n15043), .B(n15044), .Z(n14881) );
  XOR2_X1 U15064 ( .A(n15045), .B(n15046), .Z(n15044) );
  NAND2_X1 U15065 ( .A1(b_7_), .A2(a_19_), .ZN(n15046) );
  INV_X1 U15066 ( .A(n15047), .ZN(n15040) );
  NOR2_X1 U15067 ( .A1(n14882), .A2(n14883), .ZN(n15047) );
  NOR2_X1 U15068 ( .A1(n8988), .A2(n14458), .ZN(n14883) );
  NAND2_X1 U15069 ( .A1(n15048), .A2(n15049), .ZN(n14882) );
  NAND2_X1 U15070 ( .A1(n14879), .A2(n15050), .ZN(n15049) );
  NAND2_X1 U15071 ( .A1(n14876), .A2(n14878), .ZN(n15050) );
  NOR2_X1 U15072 ( .A1(n14458), .A2(n8630), .ZN(n14879) );
  INV_X1 U15073 ( .A(n15051), .ZN(n15048) );
  NOR2_X1 U15074 ( .A1(n14876), .A2(n14878), .ZN(n15051) );
  NOR2_X1 U15075 ( .A1(n15052), .A2(n15053), .ZN(n14878) );
  INV_X1 U15076 ( .A(n15054), .ZN(n15053) );
  NAND2_X1 U15077 ( .A1(n14875), .A2(n15055), .ZN(n15054) );
  NAND2_X1 U15078 ( .A1(n14874), .A2(n14873), .ZN(n15055) );
  NOR2_X1 U15079 ( .A1(n14458), .A2(n8986), .ZN(n14875) );
  NOR2_X1 U15080 ( .A1(n14873), .A2(n14874), .ZN(n15052) );
  NOR2_X1 U15081 ( .A1(n15056), .A2(n15057), .ZN(n14874) );
  NOR2_X1 U15082 ( .A1(n14797), .A2(n15058), .ZN(n15057) );
  NOR2_X1 U15083 ( .A1(n14794), .A2(n14796), .ZN(n15058) );
  NAND2_X1 U15084 ( .A1(b_8_), .A2(a_21_), .ZN(n14797) );
  INV_X1 U15085 ( .A(n15059), .ZN(n15056) );
  NAND2_X1 U15086 ( .A1(n14794), .A2(n14796), .ZN(n15059) );
  NAND2_X1 U15087 ( .A1(n15060), .A2(n15061), .ZN(n14796) );
  NAND2_X1 U15088 ( .A1(n14871), .A2(n15062), .ZN(n15061) );
  INV_X1 U15089 ( .A(n15063), .ZN(n15062) );
  NOR2_X1 U15090 ( .A1(n14870), .A2(n14868), .ZN(n15063) );
  NOR2_X1 U15091 ( .A1(n14458), .A2(n8984), .ZN(n14871) );
  NAND2_X1 U15092 ( .A1(n14868), .A2(n14870), .ZN(n15060) );
  NAND2_X1 U15093 ( .A1(n15064), .A2(n15065), .ZN(n14870) );
  NAND2_X1 U15094 ( .A1(n14867), .A2(n15066), .ZN(n15065) );
  INV_X1 U15095 ( .A(n15067), .ZN(n15066) );
  NOR2_X1 U15096 ( .A1(n14866), .A2(n14865), .ZN(n15067) );
  NOR2_X1 U15097 ( .A1(n14458), .A2(n8572), .ZN(n14867) );
  NAND2_X1 U15098 ( .A1(n14865), .A2(n14866), .ZN(n15064) );
  NAND2_X1 U15099 ( .A1(n15068), .A2(n15069), .ZN(n14866) );
  NAND2_X1 U15100 ( .A1(n14863), .A2(n15070), .ZN(n15069) );
  INV_X1 U15101 ( .A(n15071), .ZN(n15070) );
  NOR2_X1 U15102 ( .A1(n14861), .A2(n14862), .ZN(n15071) );
  NOR2_X1 U15103 ( .A1(n14458), .A2(n8982), .ZN(n14863) );
  NAND2_X1 U15104 ( .A1(n14861), .A2(n14862), .ZN(n15068) );
  NAND2_X1 U15105 ( .A1(n15072), .A2(n15073), .ZN(n14862) );
  NAND2_X1 U15106 ( .A1(n14859), .A2(n15074), .ZN(n15073) );
  NAND2_X1 U15107 ( .A1(n14856), .A2(n14858), .ZN(n15074) );
  NOR2_X1 U15108 ( .A1(n14458), .A2(n8541), .ZN(n14859) );
  INV_X1 U15109 ( .A(n15075), .ZN(n15072) );
  NOR2_X1 U15110 ( .A1(n14858), .A2(n14856), .ZN(n15075) );
  XNOR2_X1 U15111 ( .A(n15076), .B(n15077), .ZN(n14856) );
  XNOR2_X1 U15112 ( .A(n15078), .B(n15079), .ZN(n15077) );
  NAND2_X1 U15113 ( .A1(n15080), .A2(n15081), .ZN(n14858) );
  NAND2_X1 U15114 ( .A1(n14818), .A2(n15082), .ZN(n15081) );
  NAND2_X1 U15115 ( .A1(n14821), .A2(n14820), .ZN(n15082) );
  XNOR2_X1 U15116 ( .A(n15083), .B(n15084), .ZN(n14818) );
  XOR2_X1 U15117 ( .A(n15085), .B(n15086), .Z(n15083) );
  INV_X1 U15118 ( .A(n15087), .ZN(n15080) );
  NOR2_X1 U15119 ( .A1(n14820), .A2(n14821), .ZN(n15087) );
  NOR2_X1 U15120 ( .A1(n9893), .A2(n14458), .ZN(n14821) );
  NAND2_X1 U15121 ( .A1(n15088), .A2(n15089), .ZN(n14820) );
  NAND2_X1 U15122 ( .A1(n14828), .A2(n15090), .ZN(n15089) );
  INV_X1 U15123 ( .A(n15091), .ZN(n15090) );
  NOR2_X1 U15124 ( .A1(n14826), .A2(n14827), .ZN(n15091) );
  NOR2_X1 U15125 ( .A1(n14458), .A2(n8512), .ZN(n14828) );
  NAND2_X1 U15126 ( .A1(n14826), .A2(n14827), .ZN(n15088) );
  NAND2_X1 U15127 ( .A1(n15092), .A2(n15093), .ZN(n14827) );
  NAND2_X1 U15128 ( .A1(n14854), .A2(n15094), .ZN(n15093) );
  INV_X1 U15129 ( .A(n15095), .ZN(n15094) );
  NOR2_X1 U15130 ( .A1(n14855), .A2(n14853), .ZN(n15095) );
  NOR2_X1 U15131 ( .A1(n14458), .A2(n8493), .ZN(n14854) );
  NAND2_X1 U15132 ( .A1(n14853), .A2(n14855), .ZN(n15092) );
  NAND2_X1 U15133 ( .A1(n15096), .A2(n15097), .ZN(n14855) );
  NAND2_X1 U15134 ( .A1(n14849), .A2(n15098), .ZN(n15097) );
  INV_X1 U15135 ( .A(n15099), .ZN(n15098) );
  NOR2_X1 U15136 ( .A1(n14850), .A2(n14851), .ZN(n15099) );
  NOR2_X1 U15137 ( .A1(n14458), .A2(n8473), .ZN(n14849) );
  NAND2_X1 U15138 ( .A1(n14851), .A2(n14850), .ZN(n15096) );
  NAND2_X1 U15139 ( .A1(n15100), .A2(n15101), .ZN(n14850) );
  NAND2_X1 U15140 ( .A1(b_6_), .A2(n15102), .ZN(n15101) );
  NAND2_X1 U15141 ( .A1(n8456), .A2(n15103), .ZN(n15102) );
  NAND2_X1 U15142 ( .A1(a_31_), .A2(n8819), .ZN(n15103) );
  NAND2_X1 U15143 ( .A1(b_7_), .A2(n15104), .ZN(n15100) );
  NAND2_X1 U15144 ( .A1(n8459), .A2(n15105), .ZN(n15104) );
  NAND2_X1 U15145 ( .A1(a_30_), .A2(n8993), .ZN(n15105) );
  NOR3_X1 U15146 ( .A1(n14458), .A2(n8979), .A3(n8819), .ZN(n14851) );
  XOR2_X1 U15147 ( .A(n15106), .B(n15107), .Z(n14853) );
  XOR2_X1 U15148 ( .A(n15108), .B(n15109), .Z(n15106) );
  XOR2_X1 U15149 ( .A(n15110), .B(n15111), .Z(n14826) );
  XOR2_X1 U15150 ( .A(n15112), .B(n15113), .Z(n15110) );
  XNOR2_X1 U15151 ( .A(n15114), .B(n15115), .ZN(n14861) );
  XNOR2_X1 U15152 ( .A(n15116), .B(n15117), .ZN(n15115) );
  XOR2_X1 U15153 ( .A(n15118), .B(n15119), .Z(n14865) );
  XOR2_X1 U15154 ( .A(n15120), .B(n15121), .Z(n15118) );
  XOR2_X1 U15155 ( .A(n15122), .B(n15123), .Z(n14868) );
  XOR2_X1 U15156 ( .A(n15124), .B(n15125), .Z(n15122) );
  XNOR2_X1 U15157 ( .A(n15126), .B(n15127), .ZN(n14794) );
  NAND2_X1 U15158 ( .A1(n15128), .A2(n15129), .ZN(n15126) );
  XOR2_X1 U15159 ( .A(n15130), .B(n15131), .Z(n14873) );
  XOR2_X1 U15160 ( .A(n15132), .B(n15133), .Z(n15130) );
  XNOR2_X1 U15161 ( .A(n15134), .B(n15135), .ZN(n14876) );
  XNOR2_X1 U15162 ( .A(n15136), .B(n15137), .ZN(n15135) );
  NAND2_X1 U15163 ( .A1(b_7_), .A2(a_20_), .ZN(n15137) );
  XOR2_X1 U15164 ( .A(n15138), .B(n15139), .Z(n14884) );
  XNOR2_X1 U15165 ( .A(n15140), .B(n15141), .ZN(n15138) );
  NOR2_X1 U15166 ( .A1(n8819), .A2(n8988), .ZN(n15141) );
  XOR2_X1 U15167 ( .A(n15142), .B(n15143), .Z(n14892) );
  XOR2_X1 U15168 ( .A(n15144), .B(n15145), .Z(n15142) );
  NOR2_X1 U15169 ( .A1(n8819), .A2(n8680), .ZN(n15145) );
  XNOR2_X1 U15170 ( .A(n15146), .B(n15147), .ZN(n14900) );
  XOR2_X1 U15171 ( .A(n15148), .B(n15149), .Z(n15147) );
  NAND2_X1 U15172 ( .A1(a_14_), .A2(b_7_), .ZN(n15149) );
  XNOR2_X1 U15173 ( .A(n15150), .B(n15151), .ZN(n14905) );
  XNOR2_X1 U15174 ( .A(n15152), .B(n15153), .ZN(n15150) );
  NOR2_X1 U15175 ( .A1(n8819), .A2(n8721), .ZN(n15153) );
  XOR2_X1 U15176 ( .A(n15154), .B(n15155), .Z(n14909) );
  XNOR2_X1 U15177 ( .A(n15156), .B(n15157), .ZN(n15154) );
  NOR2_X1 U15178 ( .A1(n8819), .A2(n8739), .ZN(n15157) );
  XOR2_X1 U15179 ( .A(n15158), .B(n15159), .Z(n14746) );
  XNOR2_X1 U15180 ( .A(n15160), .B(n15161), .ZN(n15158) );
  NOR2_X1 U15181 ( .A1(n8819), .A2(n8749), .ZN(n15161) );
  XOR2_X1 U15182 ( .A(n15162), .B(n15163), .Z(n14738) );
  XNOR2_X1 U15183 ( .A(n15164), .B(n15165), .ZN(n15162) );
  NOR2_X1 U15184 ( .A1(n8819), .A2(n8769), .ZN(n15165) );
  XOR2_X1 U15185 ( .A(n15166), .B(n15167), .Z(n14915) );
  XNOR2_X1 U15186 ( .A(n15168), .B(n15169), .ZN(n15167) );
  NAND2_X1 U15187 ( .A1(a_8_), .A2(b_7_), .ZN(n15169) );
  XNOR2_X1 U15188 ( .A(n15170), .B(n15171), .ZN(n14919) );
  XOR2_X1 U15189 ( .A(n15172), .B(n8814), .Z(n15170) );
  XOR2_X1 U15190 ( .A(n15173), .B(n15174), .Z(n14924) );
  XNOR2_X1 U15191 ( .A(n15175), .B(n15176), .ZN(n15174) );
  XNOR2_X1 U15192 ( .A(n15177), .B(n15178), .ZN(n14928) );
  XNOR2_X1 U15193 ( .A(n15179), .B(n15180), .ZN(n15177) );
  XNOR2_X1 U15194 ( .A(n15181), .B(n15182), .ZN(n14932) );
  XOR2_X1 U15195 ( .A(n15183), .B(n15184), .Z(n15182) );
  XNOR2_X1 U15196 ( .A(n15185), .B(n15186), .ZN(n14936) );
  XNOR2_X1 U15197 ( .A(n15187), .B(n15188), .ZN(n15185) );
  XNOR2_X1 U15198 ( .A(n15189), .B(n15190), .ZN(n14703) );
  XNOR2_X1 U15199 ( .A(n15191), .B(n15192), .ZN(n15189) );
  XNOR2_X1 U15200 ( .A(n15193), .B(n15194), .ZN(n14446) );
  XOR2_X1 U15201 ( .A(n15195), .B(n15196), .Z(n15194) );
  XNOR2_X1 U15202 ( .A(n15197), .B(n14950), .ZN(n8440) );
  XOR2_X1 U15203 ( .A(n15198), .B(n15199), .Z(n14950) );
  XOR2_X1 U15204 ( .A(n15200), .B(n15201), .Z(n15199) );
  NAND2_X1 U15205 ( .A1(a_1_), .A2(b_6_), .ZN(n15201) );
  XNOR2_X1 U15206 ( .A(n14949), .B(n14947), .ZN(n15197) );
  NOR2_X1 U15207 ( .A1(n9471), .A2(n8819), .ZN(n14947) );
  NOR2_X1 U15208 ( .A1(n15202), .A2(n15203), .ZN(n14949) );
  INV_X1 U15209 ( .A(n15204), .ZN(n15203) );
  NAND2_X1 U15210 ( .A1(n15196), .A2(n15205), .ZN(n15204) );
  NAND2_X1 U15211 ( .A1(n15195), .A2(n15193), .ZN(n15205) );
  NOR2_X1 U15212 ( .A1(n9731), .A2(n8819), .ZN(n15196) );
  NOR2_X1 U15213 ( .A1(n15193), .A2(n15195), .ZN(n15202) );
  NOR2_X1 U15214 ( .A1(n15206), .A2(n15207), .ZN(n15195) );
  INV_X1 U15215 ( .A(n15208), .ZN(n15207) );
  NAND2_X1 U15216 ( .A1(n15192), .A2(n15209), .ZN(n15208) );
  NAND2_X1 U15217 ( .A1(n15190), .A2(n15191), .ZN(n15209) );
  NOR2_X1 U15218 ( .A1(n8998), .A2(n8819), .ZN(n15192) );
  NOR2_X1 U15219 ( .A1(n15190), .A2(n15191), .ZN(n15206) );
  NOR2_X1 U15220 ( .A1(n15210), .A2(n15211), .ZN(n15191) );
  INV_X1 U15221 ( .A(n15212), .ZN(n15211) );
  NAND2_X1 U15222 ( .A1(n15188), .A2(n15213), .ZN(n15212) );
  NAND2_X1 U15223 ( .A1(n15187), .A2(n15186), .ZN(n15213) );
  NOR2_X1 U15224 ( .A1(n8877), .A2(n8819), .ZN(n15188) );
  NOR2_X1 U15225 ( .A1(n15186), .A2(n15187), .ZN(n15210) );
  NOR2_X1 U15226 ( .A1(n15214), .A2(n15215), .ZN(n15187) );
  INV_X1 U15227 ( .A(n15216), .ZN(n15215) );
  NAND2_X1 U15228 ( .A1(n15184), .A2(n15217), .ZN(n15216) );
  NAND2_X1 U15229 ( .A1(n15183), .A2(n15181), .ZN(n15217) );
  NOR2_X1 U15230 ( .A1(n8996), .A2(n8819), .ZN(n15184) );
  NOR2_X1 U15231 ( .A1(n15181), .A2(n15183), .ZN(n15214) );
  NOR2_X1 U15232 ( .A1(n15218), .A2(n15219), .ZN(n15183) );
  INV_X1 U15233 ( .A(n15220), .ZN(n15219) );
  NAND2_X1 U15234 ( .A1(n15180), .A2(n15221), .ZN(n15220) );
  NAND2_X1 U15235 ( .A1(n15179), .A2(n15178), .ZN(n15221) );
  NOR2_X1 U15236 ( .A1(n8848), .A2(n8819), .ZN(n15180) );
  NOR2_X1 U15237 ( .A1(n15178), .A2(n15179), .ZN(n15218) );
  NOR2_X1 U15238 ( .A1(n15222), .A2(n15223), .ZN(n15179) );
  INV_X1 U15239 ( .A(n15224), .ZN(n15223) );
  NAND2_X1 U15240 ( .A1(n15176), .A2(n15225), .ZN(n15224) );
  NAND2_X1 U15241 ( .A1(n15173), .A2(n15175), .ZN(n15225) );
  NOR2_X1 U15242 ( .A1(n8994), .A2(n8819), .ZN(n15176) );
  NOR2_X1 U15243 ( .A1(n15175), .A2(n15173), .ZN(n15222) );
  XNOR2_X1 U15244 ( .A(n15226), .B(n15227), .ZN(n15173) );
  XOR2_X1 U15245 ( .A(n15228), .B(n15229), .Z(n15227) );
  NAND2_X1 U15246 ( .A1(n15230), .A2(n15231), .ZN(n15175) );
  NAND2_X1 U15247 ( .A1(n15171), .A2(n15232), .ZN(n15231) );
  NAND2_X1 U15248 ( .A1(n8814), .A2(n15172), .ZN(n15232) );
  INV_X1 U15249 ( .A(n15233), .ZN(n15172) );
  INV_X1 U15250 ( .A(n8930), .ZN(n8814) );
  XOR2_X1 U15251 ( .A(n15234), .B(n15235), .Z(n15171) );
  XNOR2_X1 U15252 ( .A(n15236), .B(n15237), .ZN(n15234) );
  NAND2_X1 U15253 ( .A1(n15233), .A2(n8930), .ZN(n15230) );
  NAND2_X1 U15254 ( .A1(a_7_), .A2(b_7_), .ZN(n8930) );
  NOR2_X1 U15255 ( .A1(n15238), .A2(n15239), .ZN(n15233) );
  INV_X1 U15256 ( .A(n15240), .ZN(n15239) );
  NAND3_X1 U15257 ( .A1(b_7_), .A2(n15241), .A3(a_8_), .ZN(n15240) );
  NAND2_X1 U15258 ( .A1(n15166), .A2(n15168), .ZN(n15241) );
  NOR2_X1 U15259 ( .A1(n15166), .A2(n15168), .ZN(n15238) );
  NOR2_X1 U15260 ( .A1(n15242), .A2(n15243), .ZN(n15168) );
  INV_X1 U15261 ( .A(n15244), .ZN(n15243) );
  NAND3_X1 U15262 ( .A1(b_7_), .A2(n15245), .A3(a_9_), .ZN(n15244) );
  NAND2_X1 U15263 ( .A1(n14993), .A2(n14992), .ZN(n15245) );
  NOR2_X1 U15264 ( .A1(n14992), .A2(n14993), .ZN(n15242) );
  NOR2_X1 U15265 ( .A1(n15246), .A2(n15247), .ZN(n14993) );
  NOR3_X1 U15266 ( .A1(n8819), .A2(n15248), .A3(n8769), .ZN(n15247) );
  INV_X1 U15267 ( .A(n15249), .ZN(n15248) );
  NAND2_X1 U15268 ( .A1(n15163), .A2(n15164), .ZN(n15249) );
  NOR2_X1 U15269 ( .A1(n15163), .A2(n15164), .ZN(n15246) );
  NOR2_X1 U15270 ( .A1(n15250), .A2(n15251), .ZN(n15164) );
  INV_X1 U15271 ( .A(n15252), .ZN(n15251) );
  NAND3_X1 U15272 ( .A1(b_7_), .A2(n15253), .A3(a_11_), .ZN(n15252) );
  NAND2_X1 U15273 ( .A1(n15159), .A2(n15160), .ZN(n15253) );
  NOR2_X1 U15274 ( .A1(n15159), .A2(n15160), .ZN(n15250) );
  NOR2_X1 U15275 ( .A1(n15254), .A2(n15255), .ZN(n15160) );
  INV_X1 U15276 ( .A(n15256), .ZN(n15255) );
  NAND3_X1 U15277 ( .A1(b_7_), .A2(n15257), .A3(a_12_), .ZN(n15256) );
  NAND2_X1 U15278 ( .A1(n15155), .A2(n15156), .ZN(n15257) );
  NOR2_X1 U15279 ( .A1(n15155), .A2(n15156), .ZN(n15254) );
  NOR2_X1 U15280 ( .A1(n15258), .A2(n15259), .ZN(n15156) );
  INV_X1 U15281 ( .A(n15260), .ZN(n15259) );
  NAND3_X1 U15282 ( .A1(b_7_), .A2(n15261), .A3(a_13_), .ZN(n15260) );
  NAND2_X1 U15283 ( .A1(n15152), .A2(n15151), .ZN(n15261) );
  NOR2_X1 U15284 ( .A1(n15151), .A2(n15152), .ZN(n15258) );
  NOR2_X1 U15285 ( .A1(n15262), .A2(n15263), .ZN(n15152) );
  NOR3_X1 U15286 ( .A1(n8819), .A2(n15264), .A3(n8991), .ZN(n15263) );
  NOR2_X1 U15287 ( .A1(n15146), .A2(n15148), .ZN(n15264) );
  INV_X1 U15288 ( .A(n15265), .ZN(n15262) );
  NAND2_X1 U15289 ( .A1(n15146), .A2(n15148), .ZN(n15265) );
  NAND2_X1 U15290 ( .A1(n15266), .A2(n15267), .ZN(n15148) );
  INV_X1 U15291 ( .A(n15268), .ZN(n15267) );
  NOR3_X1 U15292 ( .A1(n8819), .A2(n15269), .A3(n8692), .ZN(n15268) );
  NOR2_X1 U15293 ( .A1(n15022), .A2(n15020), .ZN(n15269) );
  NAND2_X1 U15294 ( .A1(n15020), .A2(n15022), .ZN(n15266) );
  NAND2_X1 U15295 ( .A1(n15270), .A2(n15271), .ZN(n15022) );
  NAND3_X1 U15296 ( .A1(b_7_), .A2(n15272), .A3(a_16_), .ZN(n15271) );
  INV_X1 U15297 ( .A(n15273), .ZN(n15272) );
  NOR2_X1 U15298 ( .A1(n15143), .A2(n15144), .ZN(n15273) );
  NAND2_X1 U15299 ( .A1(n15143), .A2(n15144), .ZN(n15270) );
  NAND2_X1 U15300 ( .A1(n15274), .A2(n15275), .ZN(n15144) );
  NAND3_X1 U15301 ( .A1(b_7_), .A2(n15276), .A3(a_17_), .ZN(n15275) );
  NAND2_X1 U15302 ( .A1(n15032), .A2(n15034), .ZN(n15276) );
  INV_X1 U15303 ( .A(n15277), .ZN(n15274) );
  NOR2_X1 U15304 ( .A1(n15032), .A2(n15034), .ZN(n15277) );
  NOR2_X1 U15305 ( .A1(n15278), .A2(n15279), .ZN(n15034) );
  INV_X1 U15306 ( .A(n15280), .ZN(n15279) );
  NAND3_X1 U15307 ( .A1(b_7_), .A2(n15281), .A3(a_18_), .ZN(n15280) );
  NAND2_X1 U15308 ( .A1(n15139), .A2(n15140), .ZN(n15281) );
  NOR2_X1 U15309 ( .A1(n15139), .A2(n15140), .ZN(n15278) );
  NOR2_X1 U15310 ( .A1(n15282), .A2(n15283), .ZN(n15140) );
  NOR3_X1 U15311 ( .A1(n8630), .A2(n15284), .A3(n8819), .ZN(n15283) );
  NOR2_X1 U15312 ( .A1(n15045), .A2(n15043), .ZN(n15284) );
  INV_X1 U15313 ( .A(n15285), .ZN(n15282) );
  NAND2_X1 U15314 ( .A1(n15043), .A2(n15045), .ZN(n15285) );
  NAND2_X1 U15315 ( .A1(n15286), .A2(n15287), .ZN(n15045) );
  NAND3_X1 U15316 ( .A1(a_20_), .A2(n15288), .A3(b_7_), .ZN(n15287) );
  NAND2_X1 U15317 ( .A1(n15289), .A2(n15290), .ZN(n15288) );
  INV_X1 U15318 ( .A(n15136), .ZN(n15290) );
  INV_X1 U15319 ( .A(n15134), .ZN(n15289) );
  NAND2_X1 U15320 ( .A1(n15136), .A2(n15134), .ZN(n15286) );
  XOR2_X1 U15321 ( .A(n15291), .B(n15292), .Z(n15134) );
  XOR2_X1 U15322 ( .A(n15293), .B(n15294), .Z(n15291) );
  NOR2_X1 U15323 ( .A1(n8601), .A2(n8993), .ZN(n15294) );
  NOR2_X1 U15324 ( .A1(n15295), .A2(n15296), .ZN(n15136) );
  INV_X1 U15325 ( .A(n15297), .ZN(n15296) );
  NAND2_X1 U15326 ( .A1(n15131), .A2(n15298), .ZN(n15297) );
  NAND2_X1 U15327 ( .A1(n15133), .A2(n15132), .ZN(n15298) );
  XOR2_X1 U15328 ( .A(n15299), .B(n15300), .Z(n15131) );
  NAND2_X1 U15329 ( .A1(n15301), .A2(n15302), .ZN(n15299) );
  NOR2_X1 U15330 ( .A1(n15132), .A2(n15133), .ZN(n15295) );
  NOR2_X1 U15331 ( .A1(n8819), .A2(n8601), .ZN(n15133) );
  NAND2_X1 U15332 ( .A1(n15128), .A2(n15303), .ZN(n15132) );
  NAND2_X1 U15333 ( .A1(n15127), .A2(n15129), .ZN(n15303) );
  NAND2_X1 U15334 ( .A1(n15304), .A2(n15305), .ZN(n15129) );
  NAND2_X1 U15335 ( .A1(b_7_), .A2(a_22_), .ZN(n15305) );
  INV_X1 U15336 ( .A(n15306), .ZN(n15304) );
  XNOR2_X1 U15337 ( .A(n15307), .B(n15308), .ZN(n15127) );
  XNOR2_X1 U15338 ( .A(n15309), .B(n15310), .ZN(n15307) );
  NOR2_X1 U15339 ( .A1(n8572), .A2(n8993), .ZN(n15310) );
  NAND2_X1 U15340 ( .A1(a_22_), .A2(n15306), .ZN(n15128) );
  NAND2_X1 U15341 ( .A1(n15311), .A2(n15312), .ZN(n15306) );
  NAND2_X1 U15342 ( .A1(n15125), .A2(n15313), .ZN(n15312) );
  INV_X1 U15343 ( .A(n15314), .ZN(n15313) );
  NOR2_X1 U15344 ( .A1(n15123), .A2(n15124), .ZN(n15314) );
  NOR2_X1 U15345 ( .A1(n8819), .A2(n8572), .ZN(n15125) );
  NAND2_X1 U15346 ( .A1(n15123), .A2(n15124), .ZN(n15311) );
  NAND2_X1 U15347 ( .A1(n15315), .A2(n15316), .ZN(n15124) );
  NAND2_X1 U15348 ( .A1(n15121), .A2(n15317), .ZN(n15316) );
  INV_X1 U15349 ( .A(n15318), .ZN(n15317) );
  NOR2_X1 U15350 ( .A1(n15119), .A2(n15120), .ZN(n15318) );
  NOR2_X1 U15351 ( .A1(n8819), .A2(n8982), .ZN(n15121) );
  NAND2_X1 U15352 ( .A1(n15119), .A2(n15120), .ZN(n15315) );
  NAND2_X1 U15353 ( .A1(n15319), .A2(n15320), .ZN(n15120) );
  NAND2_X1 U15354 ( .A1(n15117), .A2(n15321), .ZN(n15320) );
  NAND2_X1 U15355 ( .A1(n15114), .A2(n15116), .ZN(n15321) );
  NOR2_X1 U15356 ( .A1(n8819), .A2(n8541), .ZN(n15117) );
  INV_X1 U15357 ( .A(n15322), .ZN(n15319) );
  NOR2_X1 U15358 ( .A1(n15116), .A2(n15114), .ZN(n15322) );
  XNOR2_X1 U15359 ( .A(n15323), .B(n15324), .ZN(n15114) );
  XNOR2_X1 U15360 ( .A(n15325), .B(n15326), .ZN(n15324) );
  NAND2_X1 U15361 ( .A1(n15327), .A2(n15328), .ZN(n15116) );
  NAND2_X1 U15362 ( .A1(n15076), .A2(n15329), .ZN(n15328) );
  NAND2_X1 U15363 ( .A1(n15079), .A2(n15078), .ZN(n15329) );
  XNOR2_X1 U15364 ( .A(n15330), .B(n15331), .ZN(n15076) );
  XOR2_X1 U15365 ( .A(n15332), .B(n15333), .Z(n15330) );
  INV_X1 U15366 ( .A(n15334), .ZN(n15327) );
  NOR2_X1 U15367 ( .A1(n15078), .A2(n15079), .ZN(n15334) );
  NOR2_X1 U15368 ( .A1(n9893), .A2(n8819), .ZN(n15079) );
  NAND2_X1 U15369 ( .A1(n15335), .A2(n15336), .ZN(n15078) );
  NAND2_X1 U15370 ( .A1(n15086), .A2(n15337), .ZN(n15336) );
  INV_X1 U15371 ( .A(n15338), .ZN(n15337) );
  NOR2_X1 U15372 ( .A1(n15084), .A2(n15085), .ZN(n15338) );
  NOR2_X1 U15373 ( .A1(n8819), .A2(n8512), .ZN(n15086) );
  NAND2_X1 U15374 ( .A1(n15084), .A2(n15085), .ZN(n15335) );
  NAND2_X1 U15375 ( .A1(n15339), .A2(n15340), .ZN(n15085) );
  NAND2_X1 U15376 ( .A1(n15112), .A2(n15341), .ZN(n15340) );
  INV_X1 U15377 ( .A(n15342), .ZN(n15341) );
  NOR2_X1 U15378 ( .A1(n15113), .A2(n15111), .ZN(n15342) );
  NOR2_X1 U15379 ( .A1(n8819), .A2(n8493), .ZN(n15112) );
  NAND2_X1 U15380 ( .A1(n15111), .A2(n15113), .ZN(n15339) );
  NAND2_X1 U15381 ( .A1(n15343), .A2(n15344), .ZN(n15113) );
  NAND2_X1 U15382 ( .A1(n15107), .A2(n15345), .ZN(n15344) );
  INV_X1 U15383 ( .A(n15346), .ZN(n15345) );
  NOR2_X1 U15384 ( .A1(n15108), .A2(n15109), .ZN(n15346) );
  NOR2_X1 U15385 ( .A1(n8819), .A2(n8473), .ZN(n15107) );
  NAND2_X1 U15386 ( .A1(n15109), .A2(n15108), .ZN(n15343) );
  NAND2_X1 U15387 ( .A1(n15347), .A2(n15348), .ZN(n15108) );
  NAND2_X1 U15388 ( .A1(b_5_), .A2(n15349), .ZN(n15348) );
  NAND2_X1 U15389 ( .A1(n8456), .A2(n15350), .ZN(n15349) );
  NAND2_X1 U15390 ( .A1(a_31_), .A2(n8993), .ZN(n15350) );
  NAND2_X1 U15391 ( .A1(b_6_), .A2(n15351), .ZN(n15347) );
  NAND2_X1 U15392 ( .A1(n8459), .A2(n15352), .ZN(n15351) );
  NAND2_X1 U15393 ( .A1(a_30_), .A2(n8846), .ZN(n15352) );
  NOR3_X1 U15394 ( .A1(n8819), .A2(n8979), .A3(n8993), .ZN(n15109) );
  XOR2_X1 U15395 ( .A(n15353), .B(n15354), .Z(n15111) );
  XOR2_X1 U15396 ( .A(n15355), .B(n15356), .Z(n15353) );
  XOR2_X1 U15397 ( .A(n15357), .B(n15358), .Z(n15084) );
  XOR2_X1 U15398 ( .A(n15359), .B(n15360), .Z(n15357) );
  XNOR2_X1 U15399 ( .A(n15361), .B(n15362), .ZN(n15119) );
  XNOR2_X1 U15400 ( .A(n15363), .B(n15364), .ZN(n15362) );
  XNOR2_X1 U15401 ( .A(n15365), .B(n15366), .ZN(n15123) );
  XNOR2_X1 U15402 ( .A(n15367), .B(n15368), .ZN(n15365) );
  NOR2_X1 U15403 ( .A1(n8982), .A2(n8993), .ZN(n15368) );
  XNOR2_X1 U15404 ( .A(n15369), .B(n15370), .ZN(n15043) );
  NAND2_X1 U15405 ( .A1(n15371), .A2(n15372), .ZN(n15369) );
  XOR2_X1 U15406 ( .A(n15373), .B(n15374), .Z(n15139) );
  XOR2_X1 U15407 ( .A(n15375), .B(n15376), .Z(n15373) );
  XOR2_X1 U15408 ( .A(n15377), .B(n15378), .Z(n15032) );
  XNOR2_X1 U15409 ( .A(n15379), .B(n15380), .ZN(n15377) );
  XNOR2_X1 U15410 ( .A(n15381), .B(n15382), .ZN(n15143) );
  XNOR2_X1 U15411 ( .A(n15383), .B(n15384), .ZN(n15382) );
  XNOR2_X1 U15412 ( .A(n15385), .B(n15386), .ZN(n15020) );
  XNOR2_X1 U15413 ( .A(n15387), .B(n15388), .ZN(n15386) );
  XOR2_X1 U15414 ( .A(n15389), .B(n15390), .Z(n15146) );
  XOR2_X1 U15415 ( .A(n15391), .B(n15392), .Z(n15389) );
  XOR2_X1 U15416 ( .A(n15393), .B(n15394), .Z(n15151) );
  XNOR2_X1 U15417 ( .A(n15395), .B(n15396), .ZN(n15393) );
  XOR2_X1 U15418 ( .A(n15397), .B(n15398), .Z(n15155) );
  XNOR2_X1 U15419 ( .A(n15399), .B(n15400), .ZN(n15397) );
  XOR2_X1 U15420 ( .A(n15401), .B(n15402), .Z(n15159) );
  XNOR2_X1 U15421 ( .A(n15403), .B(n15404), .ZN(n15401) );
  XNOR2_X1 U15422 ( .A(n15405), .B(n15406), .ZN(n15163) );
  XOR2_X1 U15423 ( .A(n15407), .B(n15408), .Z(n15406) );
  XNOR2_X1 U15424 ( .A(n15409), .B(n15410), .ZN(n14992) );
  XOR2_X1 U15425 ( .A(n15411), .B(n15412), .Z(n15409) );
  XNOR2_X1 U15426 ( .A(n15413), .B(n15414), .ZN(n15166) );
  XOR2_X1 U15427 ( .A(n15415), .B(n15416), .Z(n15413) );
  XOR2_X1 U15428 ( .A(n15417), .B(n15418), .Z(n15178) );
  XNOR2_X1 U15429 ( .A(n15419), .B(n15420), .ZN(n15417) );
  XOR2_X1 U15430 ( .A(n15421), .B(n15422), .Z(n15181) );
  XNOR2_X1 U15431 ( .A(n15423), .B(n15424), .ZN(n15422) );
  XOR2_X1 U15432 ( .A(n15425), .B(n15426), .Z(n15186) );
  XNOR2_X1 U15433 ( .A(n15427), .B(n15428), .ZN(n15426) );
  XNOR2_X1 U15434 ( .A(n15429), .B(n15430), .ZN(n15190) );
  XOR2_X1 U15435 ( .A(n15431), .B(n15432), .Z(n15429) );
  XNOR2_X1 U15436 ( .A(n15433), .B(n15434), .ZN(n15193) );
  XOR2_X1 U15437 ( .A(n15435), .B(n15436), .Z(n15433) );
  XOR2_X1 U15438 ( .A(n8502), .B(n8501), .Z(n8443) );
  INV_X1 U15439 ( .A(n8497), .ZN(n9141) );
  NAND3_X1 U15440 ( .A1(n8501), .A2(n8502), .A3(n15437), .ZN(n8497) );
  INV_X1 U15441 ( .A(n8500), .ZN(n15437) );
  NAND2_X1 U15442 ( .A1(n9140), .A2(n15438), .ZN(n8500) );
  NAND2_X1 U15443 ( .A1(n15439), .A2(n15440), .ZN(n15438) );
  INV_X1 U15444 ( .A(n15441), .ZN(n9140) );
  NOR2_X1 U15445 ( .A1(n15440), .A2(n15439), .ZN(n15441) );
  NOR2_X1 U15446 ( .A1(n15442), .A2(n15443), .ZN(n15439) );
  INV_X1 U15447 ( .A(n15444), .ZN(n15443) );
  NAND2_X1 U15448 ( .A1(n15445), .A2(n15446), .ZN(n15444) );
  NAND2_X1 U15449 ( .A1(n15447), .A2(n15448), .ZN(n15446) );
  NOR2_X1 U15450 ( .A1(n15448), .A2(n15447), .ZN(n15442) );
  XNOR2_X1 U15451 ( .A(n15449), .B(n15450), .ZN(n15440) );
  XOR2_X1 U15452 ( .A(n15451), .B(n15452), .Z(n15449) );
  NOR2_X1 U15453 ( .A1(n8995), .A2(n9471), .ZN(n15452) );
  NAND2_X1 U15454 ( .A1(n15453), .A2(n15454), .ZN(n8502) );
  NAND3_X1 U15455 ( .A1(b_6_), .A2(n15455), .A3(a_0_), .ZN(n15454) );
  NAND2_X1 U15456 ( .A1(n14953), .A2(n14952), .ZN(n15455) );
  INV_X1 U15457 ( .A(n15456), .ZN(n15453) );
  NOR2_X1 U15458 ( .A1(n14952), .A2(n14953), .ZN(n15456) );
  NOR2_X1 U15459 ( .A1(n15457), .A2(n15458), .ZN(n14953) );
  NOR3_X1 U15460 ( .A1(n8993), .A2(n15459), .A3(n9731), .ZN(n15458) );
  NOR2_X1 U15461 ( .A1(n15198), .A2(n15200), .ZN(n15459) );
  INV_X1 U15462 ( .A(n15460), .ZN(n15457) );
  NAND2_X1 U15463 ( .A1(n15198), .A2(n15200), .ZN(n15460) );
  NAND2_X1 U15464 ( .A1(n15461), .A2(n15462), .ZN(n15200) );
  NAND2_X1 U15465 ( .A1(n15436), .A2(n15463), .ZN(n15462) );
  INV_X1 U15466 ( .A(n15464), .ZN(n15463) );
  NOR2_X1 U15467 ( .A1(n15434), .A2(n15435), .ZN(n15464) );
  NOR2_X1 U15468 ( .A1(n8998), .A2(n8993), .ZN(n15436) );
  NAND2_X1 U15469 ( .A1(n15434), .A2(n15435), .ZN(n15461) );
  NAND2_X1 U15470 ( .A1(n15465), .A2(n15466), .ZN(n15435) );
  NAND2_X1 U15471 ( .A1(n15432), .A2(n15467), .ZN(n15466) );
  INV_X1 U15472 ( .A(n15468), .ZN(n15467) );
  NOR2_X1 U15473 ( .A1(n15431), .A2(n15430), .ZN(n15468) );
  NOR2_X1 U15474 ( .A1(n8877), .A2(n8993), .ZN(n15432) );
  NAND2_X1 U15475 ( .A1(n15430), .A2(n15431), .ZN(n15465) );
  NAND2_X1 U15476 ( .A1(n15469), .A2(n15470), .ZN(n15431) );
  NAND2_X1 U15477 ( .A1(n15428), .A2(n15471), .ZN(n15470) );
  INV_X1 U15478 ( .A(n15472), .ZN(n15471) );
  NOR2_X1 U15479 ( .A1(n15425), .A2(n15427), .ZN(n15472) );
  NOR2_X1 U15480 ( .A1(n8996), .A2(n8993), .ZN(n15428) );
  NAND2_X1 U15481 ( .A1(n15425), .A2(n15427), .ZN(n15469) );
  NAND2_X1 U15482 ( .A1(n15473), .A2(n15474), .ZN(n15427) );
  NAND2_X1 U15483 ( .A1(n15424), .A2(n15475), .ZN(n15474) );
  NAND2_X1 U15484 ( .A1(n15421), .A2(n15423), .ZN(n15475) );
  NOR2_X1 U15485 ( .A1(n8848), .A2(n8993), .ZN(n15424) );
  INV_X1 U15486 ( .A(n15476), .ZN(n15473) );
  NOR2_X1 U15487 ( .A1(n15421), .A2(n15423), .ZN(n15476) );
  NAND2_X1 U15488 ( .A1(n15477), .A2(n15478), .ZN(n15423) );
  NAND2_X1 U15489 ( .A1(n15418), .A2(n15479), .ZN(n15478) );
  NAND2_X1 U15490 ( .A1(n15420), .A2(n15480), .ZN(n15479) );
  INV_X1 U15491 ( .A(n15419), .ZN(n15480) );
  XOR2_X1 U15492 ( .A(n15481), .B(n15482), .Z(n15418) );
  XNOR2_X1 U15493 ( .A(n15483), .B(n15484), .ZN(n15481) );
  NOR2_X1 U15494 ( .A1(n8846), .A2(n8817), .ZN(n15484) );
  NAND2_X1 U15495 ( .A1(n15419), .A2(n8831), .ZN(n15477) );
  INV_X1 U15496 ( .A(n15420), .ZN(n8831) );
  NOR2_X1 U15497 ( .A1(n8994), .A2(n8993), .ZN(n15420) );
  NOR2_X1 U15498 ( .A1(n15485), .A2(n15486), .ZN(n15419) );
  INV_X1 U15499 ( .A(n15487), .ZN(n15486) );
  NAND2_X1 U15500 ( .A1(n15229), .A2(n15488), .ZN(n15487) );
  NAND2_X1 U15501 ( .A1(n15228), .A2(n15226), .ZN(n15488) );
  NOR2_X1 U15502 ( .A1(n8817), .A2(n8993), .ZN(n15229) );
  NOR2_X1 U15503 ( .A1(n15226), .A2(n15228), .ZN(n15485) );
  NOR2_X1 U15504 ( .A1(n15489), .A2(n15490), .ZN(n15228) );
  INV_X1 U15505 ( .A(n15491), .ZN(n15490) );
  NAND2_X1 U15506 ( .A1(n15237), .A2(n15492), .ZN(n15491) );
  NAND2_X1 U15507 ( .A1(n15235), .A2(n15236), .ZN(n15492) );
  NOR2_X1 U15508 ( .A1(n10513), .A2(n8993), .ZN(n15237) );
  NOR2_X1 U15509 ( .A1(n15235), .A2(n15236), .ZN(n15489) );
  INV_X1 U15510 ( .A(n15493), .ZN(n15236) );
  NAND2_X1 U15511 ( .A1(n15494), .A2(n15495), .ZN(n15493) );
  NAND2_X1 U15512 ( .A1(n15416), .A2(n15496), .ZN(n15495) );
  INV_X1 U15513 ( .A(n15497), .ZN(n15496) );
  NOR2_X1 U15514 ( .A1(n15415), .A2(n15414), .ZN(n15497) );
  NOR2_X1 U15515 ( .A1(n8779), .A2(n8993), .ZN(n15416) );
  NAND2_X1 U15516 ( .A1(n15414), .A2(n15415), .ZN(n15494) );
  NAND2_X1 U15517 ( .A1(n15498), .A2(n15499), .ZN(n15415) );
  NAND2_X1 U15518 ( .A1(n15412), .A2(n15500), .ZN(n15499) );
  INV_X1 U15519 ( .A(n15501), .ZN(n15500) );
  NOR2_X1 U15520 ( .A1(n15410), .A2(n15411), .ZN(n15501) );
  NOR2_X1 U15521 ( .A1(n8769), .A2(n8993), .ZN(n15412) );
  NAND2_X1 U15522 ( .A1(n15410), .A2(n15411), .ZN(n15498) );
  NAND2_X1 U15523 ( .A1(n15502), .A2(n15503), .ZN(n15411) );
  NAND2_X1 U15524 ( .A1(n15408), .A2(n15504), .ZN(n15503) );
  NAND2_X1 U15525 ( .A1(n15407), .A2(n15405), .ZN(n15504) );
  NOR2_X1 U15526 ( .A1(n8749), .A2(n8993), .ZN(n15408) );
  INV_X1 U15527 ( .A(n15505), .ZN(n15502) );
  NOR2_X1 U15528 ( .A1(n15405), .A2(n15407), .ZN(n15505) );
  NOR2_X1 U15529 ( .A1(n15506), .A2(n15507), .ZN(n15407) );
  INV_X1 U15530 ( .A(n15508), .ZN(n15507) );
  NAND2_X1 U15531 ( .A1(n15404), .A2(n15509), .ZN(n15508) );
  NAND2_X1 U15532 ( .A1(n15403), .A2(n15402), .ZN(n15509) );
  NOR2_X1 U15533 ( .A1(n8739), .A2(n8993), .ZN(n15404) );
  NOR2_X1 U15534 ( .A1(n15402), .A2(n15403), .ZN(n15506) );
  NOR2_X1 U15535 ( .A1(n15510), .A2(n15511), .ZN(n15403) );
  INV_X1 U15536 ( .A(n15512), .ZN(n15511) );
  NAND2_X1 U15537 ( .A1(n15400), .A2(n15513), .ZN(n15512) );
  NAND2_X1 U15538 ( .A1(n15399), .A2(n15398), .ZN(n15513) );
  NOR2_X1 U15539 ( .A1(n8721), .A2(n8993), .ZN(n15400) );
  NOR2_X1 U15540 ( .A1(n15398), .A2(n15399), .ZN(n15510) );
  NOR2_X1 U15541 ( .A1(n15514), .A2(n15515), .ZN(n15399) );
  INV_X1 U15542 ( .A(n15516), .ZN(n15515) );
  NAND2_X1 U15543 ( .A1(n15396), .A2(n15517), .ZN(n15516) );
  NAND2_X1 U15544 ( .A1(n15394), .A2(n15395), .ZN(n15517) );
  NOR2_X1 U15545 ( .A1(n8991), .A2(n8993), .ZN(n15396) );
  NOR2_X1 U15546 ( .A1(n15394), .A2(n15395), .ZN(n15514) );
  INV_X1 U15547 ( .A(n15518), .ZN(n15395) );
  NAND2_X1 U15548 ( .A1(n15519), .A2(n15520), .ZN(n15518) );
  NAND2_X1 U15549 ( .A1(n15392), .A2(n15521), .ZN(n15520) );
  INV_X1 U15550 ( .A(n15522), .ZN(n15521) );
  NOR2_X1 U15551 ( .A1(n15391), .A2(n15390), .ZN(n15522) );
  NOR2_X1 U15552 ( .A1(n8692), .A2(n8993), .ZN(n15392) );
  NAND2_X1 U15553 ( .A1(n15390), .A2(n15391), .ZN(n15519) );
  NAND2_X1 U15554 ( .A1(n15523), .A2(n15524), .ZN(n15391) );
  NAND2_X1 U15555 ( .A1(n15388), .A2(n15525), .ZN(n15524) );
  INV_X1 U15556 ( .A(n15526), .ZN(n15525) );
  NOR2_X1 U15557 ( .A1(n15385), .A2(n15387), .ZN(n15526) );
  NOR2_X1 U15558 ( .A1(n8680), .A2(n8993), .ZN(n15388) );
  NAND2_X1 U15559 ( .A1(n15385), .A2(n15387), .ZN(n15523) );
  NAND2_X1 U15560 ( .A1(n15527), .A2(n15528), .ZN(n15387) );
  NAND2_X1 U15561 ( .A1(n15384), .A2(n15529), .ZN(n15528) );
  INV_X1 U15562 ( .A(n15530), .ZN(n15529) );
  NOR2_X1 U15563 ( .A1(n15383), .A2(n15381), .ZN(n15530) );
  NOR2_X1 U15564 ( .A1(n8662), .A2(n8993), .ZN(n15384) );
  NAND2_X1 U15565 ( .A1(n15381), .A2(n15383), .ZN(n15527) );
  NAND2_X1 U15566 ( .A1(n15531), .A2(n15532), .ZN(n15383) );
  NAND2_X1 U15567 ( .A1(n15380), .A2(n15533), .ZN(n15532) );
  INV_X1 U15568 ( .A(n15534), .ZN(n15533) );
  NOR2_X1 U15569 ( .A1(n15378), .A2(n15379), .ZN(n15534) );
  NOR2_X1 U15570 ( .A1(n8988), .A2(n8993), .ZN(n15380) );
  NAND2_X1 U15571 ( .A1(n15379), .A2(n15378), .ZN(n15531) );
  XNOR2_X1 U15572 ( .A(n15535), .B(n15536), .ZN(n15378) );
  XNOR2_X1 U15573 ( .A(n15537), .B(n15538), .ZN(n15535) );
  NOR2_X1 U15574 ( .A1(n8630), .A2(n8846), .ZN(n15538) );
  NOR2_X1 U15575 ( .A1(n15539), .A2(n15540), .ZN(n15379) );
  INV_X1 U15576 ( .A(n15541), .ZN(n15540) );
  NAND2_X1 U15577 ( .A1(n15374), .A2(n15542), .ZN(n15541) );
  NAND2_X1 U15578 ( .A1(n15376), .A2(n15375), .ZN(n15542) );
  XNOR2_X1 U15579 ( .A(n15543), .B(n15544), .ZN(n15374) );
  XOR2_X1 U15580 ( .A(n15545), .B(n15546), .Z(n15543) );
  NOR2_X1 U15581 ( .A1(n8986), .A2(n8846), .ZN(n15546) );
  NOR2_X1 U15582 ( .A1(n15375), .A2(n15376), .ZN(n15539) );
  NOR2_X1 U15583 ( .A1(n8993), .A2(n8630), .ZN(n15376) );
  NAND2_X1 U15584 ( .A1(n15371), .A2(n15547), .ZN(n15375) );
  NAND2_X1 U15585 ( .A1(n15370), .A2(n15372), .ZN(n15547) );
  NAND2_X1 U15586 ( .A1(n15548), .A2(n15549), .ZN(n15372) );
  NAND2_X1 U15587 ( .A1(b_6_), .A2(a_20_), .ZN(n15549) );
  XOR2_X1 U15588 ( .A(n15550), .B(n15551), .Z(n15370) );
  XNOR2_X1 U15589 ( .A(n15552), .B(n15553), .ZN(n15551) );
  NAND2_X1 U15590 ( .A1(b_5_), .A2(a_21_), .ZN(n15553) );
  INV_X1 U15591 ( .A(n15554), .ZN(n15371) );
  NOR2_X1 U15592 ( .A1(n8986), .A2(n15548), .ZN(n15554) );
  NOR2_X1 U15593 ( .A1(n15555), .A2(n15556), .ZN(n15548) );
  NOR3_X1 U15594 ( .A1(n8601), .A2(n15557), .A3(n8993), .ZN(n15556) );
  NOR2_X1 U15595 ( .A1(n15293), .A2(n15292), .ZN(n15557) );
  INV_X1 U15596 ( .A(n15558), .ZN(n15555) );
  NAND2_X1 U15597 ( .A1(n15292), .A2(n15293), .ZN(n15558) );
  NAND2_X1 U15598 ( .A1(n15301), .A2(n15559), .ZN(n15293) );
  NAND2_X1 U15599 ( .A1(n15300), .A2(n15302), .ZN(n15559) );
  NAND2_X1 U15600 ( .A1(n15560), .A2(n15561), .ZN(n15302) );
  NAND2_X1 U15601 ( .A1(b_6_), .A2(a_22_), .ZN(n15561) );
  XNOR2_X1 U15602 ( .A(n15562), .B(n15563), .ZN(n15300) );
  XOR2_X1 U15603 ( .A(n15564), .B(n15565), .Z(n15562) );
  NAND2_X1 U15604 ( .A1(a_22_), .A2(n15566), .ZN(n15301) );
  INV_X1 U15605 ( .A(n15560), .ZN(n15566) );
  NOR2_X1 U15606 ( .A1(n15567), .A2(n15568), .ZN(n15560) );
  NOR3_X1 U15607 ( .A1(n8572), .A2(n15569), .A3(n8993), .ZN(n15568) );
  INV_X1 U15608 ( .A(n15570), .ZN(n15569) );
  NAND2_X1 U15609 ( .A1(n15309), .A2(n15308), .ZN(n15570) );
  NOR2_X1 U15610 ( .A1(n15308), .A2(n15309), .ZN(n15567) );
  NOR2_X1 U15611 ( .A1(n15571), .A2(n15572), .ZN(n15309) );
  INV_X1 U15612 ( .A(n15573), .ZN(n15572) );
  NAND3_X1 U15613 ( .A1(a_24_), .A2(n15574), .A3(b_6_), .ZN(n15573) );
  NAND2_X1 U15614 ( .A1(n15367), .A2(n15366), .ZN(n15574) );
  NOR2_X1 U15615 ( .A1(n15366), .A2(n15367), .ZN(n15571) );
  NOR2_X1 U15616 ( .A1(n15575), .A2(n15576), .ZN(n15367) );
  INV_X1 U15617 ( .A(n15577), .ZN(n15576) );
  NAND2_X1 U15618 ( .A1(n15364), .A2(n15578), .ZN(n15577) );
  NAND2_X1 U15619 ( .A1(n15361), .A2(n15363), .ZN(n15578) );
  NOR2_X1 U15620 ( .A1(n8993), .A2(n8541), .ZN(n15364) );
  NOR2_X1 U15621 ( .A1(n15363), .A2(n15361), .ZN(n15575) );
  XNOR2_X1 U15622 ( .A(n15579), .B(n15580), .ZN(n15361) );
  XNOR2_X1 U15623 ( .A(n15581), .B(n15582), .ZN(n15580) );
  NAND2_X1 U15624 ( .A1(n15583), .A2(n15584), .ZN(n15363) );
  NAND2_X1 U15625 ( .A1(n15323), .A2(n15585), .ZN(n15584) );
  NAND2_X1 U15626 ( .A1(n15326), .A2(n15325), .ZN(n15585) );
  XNOR2_X1 U15627 ( .A(n15586), .B(n15587), .ZN(n15323) );
  XOR2_X1 U15628 ( .A(n15588), .B(n15589), .Z(n15586) );
  INV_X1 U15629 ( .A(n15590), .ZN(n15583) );
  NOR2_X1 U15630 ( .A1(n15325), .A2(n15326), .ZN(n15590) );
  NOR2_X1 U15631 ( .A1(n8993), .A2(n9893), .ZN(n15326) );
  NAND2_X1 U15632 ( .A1(n15591), .A2(n15592), .ZN(n15325) );
  NAND2_X1 U15633 ( .A1(n15333), .A2(n15593), .ZN(n15592) );
  INV_X1 U15634 ( .A(n15594), .ZN(n15593) );
  NOR2_X1 U15635 ( .A1(n15331), .A2(n15332), .ZN(n15594) );
  NOR2_X1 U15636 ( .A1(n8993), .A2(n8512), .ZN(n15333) );
  NAND2_X1 U15637 ( .A1(n15331), .A2(n15332), .ZN(n15591) );
  NAND2_X1 U15638 ( .A1(n15595), .A2(n15596), .ZN(n15332) );
  NAND2_X1 U15639 ( .A1(n15359), .A2(n15597), .ZN(n15596) );
  INV_X1 U15640 ( .A(n15598), .ZN(n15597) );
  NOR2_X1 U15641 ( .A1(n15360), .A2(n15358), .ZN(n15598) );
  NOR2_X1 U15642 ( .A1(n8993), .A2(n8493), .ZN(n15359) );
  NAND2_X1 U15643 ( .A1(n15358), .A2(n15360), .ZN(n15595) );
  NAND2_X1 U15644 ( .A1(n15599), .A2(n15600), .ZN(n15360) );
  NAND2_X1 U15645 ( .A1(n15354), .A2(n15601), .ZN(n15600) );
  INV_X1 U15646 ( .A(n15602), .ZN(n15601) );
  NOR2_X1 U15647 ( .A1(n15355), .A2(n15356), .ZN(n15602) );
  NOR2_X1 U15648 ( .A1(n8993), .A2(n8473), .ZN(n15354) );
  NAND2_X1 U15649 ( .A1(n15356), .A2(n15355), .ZN(n15599) );
  NAND2_X1 U15650 ( .A1(n15603), .A2(n15604), .ZN(n15355) );
  NAND2_X1 U15651 ( .A1(b_4_), .A2(n15605), .ZN(n15604) );
  NAND2_X1 U15652 ( .A1(n8456), .A2(n15606), .ZN(n15605) );
  NAND2_X1 U15653 ( .A1(a_31_), .A2(n8846), .ZN(n15606) );
  NAND2_X1 U15654 ( .A1(b_5_), .A2(n15607), .ZN(n15603) );
  NAND2_X1 U15655 ( .A1(n8459), .A2(n15608), .ZN(n15607) );
  NAND2_X1 U15656 ( .A1(a_30_), .A2(n8995), .ZN(n15608) );
  NOR3_X1 U15657 ( .A1(n8993), .A2(n8979), .A3(n8846), .ZN(n15356) );
  XOR2_X1 U15658 ( .A(n15609), .B(n15610), .Z(n15358) );
  XOR2_X1 U15659 ( .A(n15611), .B(n15612), .Z(n15609) );
  XOR2_X1 U15660 ( .A(n15613), .B(n15614), .Z(n15331) );
  XOR2_X1 U15661 ( .A(n15615), .B(n15616), .Z(n15613) );
  XNOR2_X1 U15662 ( .A(n15617), .B(n15618), .ZN(n15366) );
  XOR2_X1 U15663 ( .A(n15619), .B(n15620), .Z(n15617) );
  XOR2_X1 U15664 ( .A(n15621), .B(n15622), .Z(n15308) );
  XNOR2_X1 U15665 ( .A(n15623), .B(n15624), .ZN(n15621) );
  NOR2_X1 U15666 ( .A1(n8982), .A2(n8846), .ZN(n15624) );
  XOR2_X1 U15667 ( .A(n15625), .B(n15626), .Z(n15292) );
  XOR2_X1 U15668 ( .A(n15627), .B(n15628), .Z(n15625) );
  NOR2_X1 U15669 ( .A1(n8984), .A2(n8846), .ZN(n15628) );
  XNOR2_X1 U15670 ( .A(n15629), .B(n15630), .ZN(n15381) );
  XNOR2_X1 U15671 ( .A(n15631), .B(n15632), .ZN(n15629) );
  NOR2_X1 U15672 ( .A1(n8846), .A2(n8988), .ZN(n15632) );
  XNOR2_X1 U15673 ( .A(n15633), .B(n15634), .ZN(n15385) );
  XNOR2_X1 U15674 ( .A(n15635), .B(n15636), .ZN(n15633) );
  NOR2_X1 U15675 ( .A1(n8846), .A2(n8662), .ZN(n15636) );
  XNOR2_X1 U15676 ( .A(n15637), .B(n15638), .ZN(n15390) );
  XNOR2_X1 U15677 ( .A(n15639), .B(n15640), .ZN(n15637) );
  NOR2_X1 U15678 ( .A1(n8846), .A2(n8680), .ZN(n15640) );
  XOR2_X1 U15679 ( .A(n15641), .B(n15642), .Z(n15394) );
  XNOR2_X1 U15680 ( .A(n15643), .B(n15644), .ZN(n15641) );
  NOR2_X1 U15681 ( .A1(n8846), .A2(n8692), .ZN(n15644) );
  XOR2_X1 U15682 ( .A(n15645), .B(n15646), .Z(n15398) );
  XNOR2_X1 U15683 ( .A(n15647), .B(n15648), .ZN(n15645) );
  NOR2_X1 U15684 ( .A1(n8846), .A2(n8991), .ZN(n15648) );
  XOR2_X1 U15685 ( .A(n15649), .B(n15650), .Z(n15402) );
  XNOR2_X1 U15686 ( .A(n15651), .B(n15652), .ZN(n15649) );
  NOR2_X1 U15687 ( .A1(n8846), .A2(n8721), .ZN(n15652) );
  XOR2_X1 U15688 ( .A(n15653), .B(n15654), .Z(n15405) );
  XNOR2_X1 U15689 ( .A(n15655), .B(n15656), .ZN(n15653) );
  NOR2_X1 U15690 ( .A1(n8846), .A2(n8739), .ZN(n15656) );
  XNOR2_X1 U15691 ( .A(n15657), .B(n15658), .ZN(n15410) );
  XNOR2_X1 U15692 ( .A(n15659), .B(n15660), .ZN(n15657) );
  NOR2_X1 U15693 ( .A1(n8846), .A2(n8749), .ZN(n15660) );
  XNOR2_X1 U15694 ( .A(n15661), .B(n15662), .ZN(n15414) );
  XNOR2_X1 U15695 ( .A(n15663), .B(n15664), .ZN(n15661) );
  NOR2_X1 U15696 ( .A1(n8846), .A2(n8769), .ZN(n15664) );
  XOR2_X1 U15697 ( .A(n15665), .B(n15666), .Z(n15235) );
  XNOR2_X1 U15698 ( .A(n15667), .B(n15668), .ZN(n15665) );
  NOR2_X1 U15699 ( .A1(n8846), .A2(n8779), .ZN(n15668) );
  XOR2_X1 U15700 ( .A(n15669), .B(n15670), .Z(n15226) );
  XNOR2_X1 U15701 ( .A(n15671), .B(n15672), .ZN(n15669) );
  NOR2_X1 U15702 ( .A1(n8846), .A2(n10513), .ZN(n15672) );
  XOR2_X1 U15703 ( .A(n15673), .B(n15674), .Z(n15421) );
  XNOR2_X1 U15704 ( .A(n15675), .B(n15676), .ZN(n15673) );
  NOR2_X1 U15705 ( .A1(n8846), .A2(n8994), .ZN(n15676) );
  XNOR2_X1 U15706 ( .A(n15677), .B(n15678), .ZN(n15425) );
  XNOR2_X1 U15707 ( .A(n8926), .B(n15679), .ZN(n15678) );
  XNOR2_X1 U15708 ( .A(n15680), .B(n15681), .ZN(n15430) );
  XNOR2_X1 U15709 ( .A(n15682), .B(n15683), .ZN(n15680) );
  NOR2_X1 U15710 ( .A1(n8846), .A2(n8996), .ZN(n15683) );
  XNOR2_X1 U15711 ( .A(n15684), .B(n15685), .ZN(n15434) );
  XNOR2_X1 U15712 ( .A(n15686), .B(n15687), .ZN(n15684) );
  NOR2_X1 U15713 ( .A1(n8846), .A2(n8877), .ZN(n15687) );
  XNOR2_X1 U15714 ( .A(n15688), .B(n15689), .ZN(n15198) );
  XNOR2_X1 U15715 ( .A(n15690), .B(n15691), .ZN(n15688) );
  NOR2_X1 U15716 ( .A1(n8846), .A2(n8998), .ZN(n15691) );
  XOR2_X1 U15717 ( .A(n15692), .B(n15693), .Z(n14952) );
  XNOR2_X1 U15718 ( .A(n15694), .B(n15695), .ZN(n15692) );
  NOR2_X1 U15719 ( .A1(n8846), .A2(n9731), .ZN(n15695) );
  XNOR2_X1 U15720 ( .A(n15696), .B(n15448), .ZN(n8501) );
  XOR2_X1 U15721 ( .A(n15697), .B(n15698), .Z(n15448) );
  XNOR2_X1 U15722 ( .A(n15699), .B(n15700), .ZN(n15697) );
  NOR2_X1 U15723 ( .A1(n8995), .A2(n9731), .ZN(n15700) );
  XNOR2_X1 U15724 ( .A(n15447), .B(n15445), .ZN(n15696) );
  NOR2_X1 U15725 ( .A1(n9471), .A2(n8846), .ZN(n15445) );
  NOR2_X1 U15726 ( .A1(n15701), .A2(n15702), .ZN(n15447) );
  INV_X1 U15727 ( .A(n15703), .ZN(n15702) );
  NAND3_X1 U15728 ( .A1(b_5_), .A2(n15704), .A3(a_1_), .ZN(n15703) );
  NAND2_X1 U15729 ( .A1(n15693), .A2(n15694), .ZN(n15704) );
  NOR2_X1 U15730 ( .A1(n15693), .A2(n15694), .ZN(n15701) );
  NOR2_X1 U15731 ( .A1(n15705), .A2(n15706), .ZN(n15694) );
  INV_X1 U15732 ( .A(n15707), .ZN(n15706) );
  NAND3_X1 U15733 ( .A1(b_5_), .A2(n15708), .A3(a_2_), .ZN(n15707) );
  NAND2_X1 U15734 ( .A1(n15690), .A2(n15689), .ZN(n15708) );
  NOR2_X1 U15735 ( .A1(n15689), .A2(n15690), .ZN(n15705) );
  NOR2_X1 U15736 ( .A1(n15709), .A2(n15710), .ZN(n15690) );
  INV_X1 U15737 ( .A(n15711), .ZN(n15710) );
  NAND3_X1 U15738 ( .A1(b_5_), .A2(n15712), .A3(a_3_), .ZN(n15711) );
  NAND2_X1 U15739 ( .A1(n15686), .A2(n15685), .ZN(n15712) );
  NOR2_X1 U15740 ( .A1(n15685), .A2(n15686), .ZN(n15709) );
  NOR2_X1 U15741 ( .A1(n15713), .A2(n15714), .ZN(n15686) );
  INV_X1 U15742 ( .A(n15715), .ZN(n15714) );
  NAND3_X1 U15743 ( .A1(b_5_), .A2(n15716), .A3(a_4_), .ZN(n15715) );
  NAND2_X1 U15744 ( .A1(n15681), .A2(n15682), .ZN(n15716) );
  NOR2_X1 U15745 ( .A1(n15681), .A2(n15682), .ZN(n15713) );
  NOR2_X1 U15746 ( .A1(n15717), .A2(n15718), .ZN(n15682) );
  INV_X1 U15747 ( .A(n15719), .ZN(n15718) );
  NAND2_X1 U15748 ( .A1(n15677), .A2(n15720), .ZN(n15719) );
  NAND2_X1 U15749 ( .A1(n15679), .A2(n8926), .ZN(n15720) );
  XNOR2_X1 U15750 ( .A(n15721), .B(n15722), .ZN(n15677) );
  XNOR2_X1 U15751 ( .A(n15723), .B(n15724), .ZN(n15722) );
  NOR2_X1 U15752 ( .A1(n8926), .A2(n15679), .ZN(n15717) );
  NOR2_X1 U15753 ( .A1(n15725), .A2(n15726), .ZN(n15679) );
  INV_X1 U15754 ( .A(n15727), .ZN(n15726) );
  NAND3_X1 U15755 ( .A1(b_5_), .A2(n15728), .A3(a_6_), .ZN(n15727) );
  NAND2_X1 U15756 ( .A1(n15674), .A2(n15675), .ZN(n15728) );
  NOR2_X1 U15757 ( .A1(n15674), .A2(n15675), .ZN(n15725) );
  NOR2_X1 U15758 ( .A1(n15729), .A2(n15730), .ZN(n15675) );
  INV_X1 U15759 ( .A(n15731), .ZN(n15730) );
  NAND3_X1 U15760 ( .A1(b_5_), .A2(n15732), .A3(a_7_), .ZN(n15731) );
  NAND2_X1 U15761 ( .A1(n15483), .A2(n15482), .ZN(n15732) );
  NOR2_X1 U15762 ( .A1(n15482), .A2(n15483), .ZN(n15729) );
  NOR2_X1 U15763 ( .A1(n15733), .A2(n15734), .ZN(n15483) );
  NOR3_X1 U15764 ( .A1(n8846), .A2(n15735), .A3(n10513), .ZN(n15734) );
  INV_X1 U15765 ( .A(n15736), .ZN(n15735) );
  NAND2_X1 U15766 ( .A1(n15670), .A2(n15671), .ZN(n15736) );
  NOR2_X1 U15767 ( .A1(n15670), .A2(n15671), .ZN(n15733) );
  NOR2_X1 U15768 ( .A1(n15737), .A2(n15738), .ZN(n15671) );
  INV_X1 U15769 ( .A(n15739), .ZN(n15738) );
  NAND3_X1 U15770 ( .A1(b_5_), .A2(n15740), .A3(a_9_), .ZN(n15739) );
  NAND2_X1 U15771 ( .A1(n15667), .A2(n15666), .ZN(n15740) );
  NOR2_X1 U15772 ( .A1(n15666), .A2(n15667), .ZN(n15737) );
  NOR2_X1 U15773 ( .A1(n15741), .A2(n15742), .ZN(n15667) );
  NOR3_X1 U15774 ( .A1(n8846), .A2(n15743), .A3(n8769), .ZN(n15742) );
  INV_X1 U15775 ( .A(n15744), .ZN(n15743) );
  NAND2_X1 U15776 ( .A1(n15662), .A2(n15663), .ZN(n15744) );
  NOR2_X1 U15777 ( .A1(n15662), .A2(n15663), .ZN(n15741) );
  NOR2_X1 U15778 ( .A1(n15745), .A2(n15746), .ZN(n15663) );
  INV_X1 U15779 ( .A(n15747), .ZN(n15746) );
  NAND3_X1 U15780 ( .A1(b_5_), .A2(n15748), .A3(a_11_), .ZN(n15747) );
  NAND2_X1 U15781 ( .A1(n15659), .A2(n15658), .ZN(n15748) );
  NOR2_X1 U15782 ( .A1(n15658), .A2(n15659), .ZN(n15745) );
  NOR2_X1 U15783 ( .A1(n15749), .A2(n15750), .ZN(n15659) );
  NOR3_X1 U15784 ( .A1(n8846), .A2(n15751), .A3(n8739), .ZN(n15750) );
  INV_X1 U15785 ( .A(n15752), .ZN(n15751) );
  NAND2_X1 U15786 ( .A1(n15654), .A2(n15655), .ZN(n15752) );
  NOR2_X1 U15787 ( .A1(n15654), .A2(n15655), .ZN(n15749) );
  NOR2_X1 U15788 ( .A1(n15753), .A2(n15754), .ZN(n15655) );
  INV_X1 U15789 ( .A(n15755), .ZN(n15754) );
  NAND3_X1 U15790 ( .A1(b_5_), .A2(n15756), .A3(a_13_), .ZN(n15755) );
  NAND2_X1 U15791 ( .A1(n15650), .A2(n15651), .ZN(n15756) );
  NOR2_X1 U15792 ( .A1(n15650), .A2(n15651), .ZN(n15753) );
  NOR2_X1 U15793 ( .A1(n15757), .A2(n15758), .ZN(n15651) );
  INV_X1 U15794 ( .A(n15759), .ZN(n15758) );
  NAND3_X1 U15795 ( .A1(b_5_), .A2(n15760), .A3(a_14_), .ZN(n15759) );
  NAND2_X1 U15796 ( .A1(n15646), .A2(n15647), .ZN(n15760) );
  NOR2_X1 U15797 ( .A1(n15646), .A2(n15647), .ZN(n15757) );
  NOR2_X1 U15798 ( .A1(n15761), .A2(n15762), .ZN(n15647) );
  INV_X1 U15799 ( .A(n15763), .ZN(n15762) );
  NAND3_X1 U15800 ( .A1(b_5_), .A2(n15764), .A3(a_15_), .ZN(n15763) );
  NAND2_X1 U15801 ( .A1(n15643), .A2(n15642), .ZN(n15764) );
  NOR2_X1 U15802 ( .A1(n15642), .A2(n15643), .ZN(n15761) );
  NOR2_X1 U15803 ( .A1(n15765), .A2(n15766), .ZN(n15643) );
  NOR3_X1 U15804 ( .A1(n8846), .A2(n15767), .A3(n8680), .ZN(n15766) );
  INV_X1 U15805 ( .A(n15768), .ZN(n15767) );
  NAND2_X1 U15806 ( .A1(n15638), .A2(n15639), .ZN(n15768) );
  NOR2_X1 U15807 ( .A1(n15638), .A2(n15639), .ZN(n15765) );
  NOR2_X1 U15808 ( .A1(n15769), .A2(n15770), .ZN(n15639) );
  INV_X1 U15809 ( .A(n15771), .ZN(n15770) );
  NAND3_X1 U15810 ( .A1(b_5_), .A2(n15772), .A3(a_17_), .ZN(n15771) );
  NAND2_X1 U15811 ( .A1(n15635), .A2(n15634), .ZN(n15772) );
  NOR2_X1 U15812 ( .A1(n15634), .A2(n15635), .ZN(n15769) );
  NOR2_X1 U15813 ( .A1(n15773), .A2(n15774), .ZN(n15635) );
  NOR3_X1 U15814 ( .A1(n8846), .A2(n15775), .A3(n8988), .ZN(n15774) );
  INV_X1 U15815 ( .A(n15776), .ZN(n15775) );
  NAND2_X1 U15816 ( .A1(n15630), .A2(n15631), .ZN(n15776) );
  NOR2_X1 U15817 ( .A1(n15630), .A2(n15631), .ZN(n15773) );
  NOR2_X1 U15818 ( .A1(n15777), .A2(n15778), .ZN(n15631) );
  INV_X1 U15819 ( .A(n15779), .ZN(n15778) );
  NAND3_X1 U15820 ( .A1(a_19_), .A2(n15780), .A3(b_5_), .ZN(n15779) );
  NAND2_X1 U15821 ( .A1(n15537), .A2(n15536), .ZN(n15780) );
  NOR2_X1 U15822 ( .A1(n15536), .A2(n15537), .ZN(n15777) );
  NOR2_X1 U15823 ( .A1(n15781), .A2(n15782), .ZN(n15537) );
  NOR3_X1 U15824 ( .A1(n8986), .A2(n15783), .A3(n8846), .ZN(n15782) );
  NOR2_X1 U15825 ( .A1(n15544), .A2(n15545), .ZN(n15783) );
  INV_X1 U15826 ( .A(n15784), .ZN(n15781) );
  NAND2_X1 U15827 ( .A1(n15544), .A2(n15545), .ZN(n15784) );
  NAND2_X1 U15828 ( .A1(n15785), .A2(n15786), .ZN(n15545) );
  NAND3_X1 U15829 ( .A1(a_21_), .A2(n15787), .A3(b_5_), .ZN(n15786) );
  NAND2_X1 U15830 ( .A1(n15550), .A2(n15552), .ZN(n15787) );
  INV_X1 U15831 ( .A(n15788), .ZN(n15785) );
  NOR2_X1 U15832 ( .A1(n15550), .A2(n15552), .ZN(n15788) );
  NOR2_X1 U15833 ( .A1(n15789), .A2(n15790), .ZN(n15552) );
  INV_X1 U15834 ( .A(n15791), .ZN(n15790) );
  NAND3_X1 U15835 ( .A1(a_22_), .A2(n15792), .A3(b_5_), .ZN(n15791) );
  NAND2_X1 U15836 ( .A1(n15626), .A2(n15627), .ZN(n15792) );
  NOR2_X1 U15837 ( .A1(n15626), .A2(n15627), .ZN(n15789) );
  NAND2_X1 U15838 ( .A1(n15793), .A2(n15794), .ZN(n15627) );
  NAND2_X1 U15839 ( .A1(n15563), .A2(n15795), .ZN(n15794) );
  NAND2_X1 U15840 ( .A1(n15565), .A2(n15564), .ZN(n15795) );
  XOR2_X1 U15841 ( .A(n15796), .B(n15797), .Z(n15563) );
  XNOR2_X1 U15842 ( .A(n15798), .B(n15799), .ZN(n15796) );
  INV_X1 U15843 ( .A(n15800), .ZN(n15793) );
  NOR2_X1 U15844 ( .A1(n15564), .A2(n15565), .ZN(n15800) );
  NOR2_X1 U15845 ( .A1(n8846), .A2(n8572), .ZN(n15565) );
  NAND2_X1 U15846 ( .A1(n15801), .A2(n15802), .ZN(n15564) );
  NAND3_X1 U15847 ( .A1(a_24_), .A2(n15803), .A3(b_5_), .ZN(n15802) );
  NAND2_X1 U15848 ( .A1(n15622), .A2(n15623), .ZN(n15803) );
  INV_X1 U15849 ( .A(n15804), .ZN(n15801) );
  NOR2_X1 U15850 ( .A1(n15622), .A2(n15623), .ZN(n15804) );
  NOR2_X1 U15851 ( .A1(n15805), .A2(n15806), .ZN(n15623) );
  INV_X1 U15852 ( .A(n15807), .ZN(n15806) );
  NAND2_X1 U15853 ( .A1(n15620), .A2(n15808), .ZN(n15807) );
  NAND2_X1 U15854 ( .A1(n15618), .A2(n15619), .ZN(n15808) );
  NOR2_X1 U15855 ( .A1(n8846), .A2(n8541), .ZN(n15620) );
  NOR2_X1 U15856 ( .A1(n15618), .A2(n15619), .ZN(n15805) );
  NAND2_X1 U15857 ( .A1(n15809), .A2(n15810), .ZN(n15619) );
  NAND2_X1 U15858 ( .A1(n15579), .A2(n15811), .ZN(n15810) );
  NAND2_X1 U15859 ( .A1(n15582), .A2(n15581), .ZN(n15811) );
  XNOR2_X1 U15860 ( .A(n15812), .B(n15813), .ZN(n15579) );
  XOR2_X1 U15861 ( .A(n15814), .B(n15815), .Z(n15812) );
  NOR2_X1 U15862 ( .A1(n8512), .A2(n8995), .ZN(n15815) );
  INV_X1 U15863 ( .A(n15816), .ZN(n15809) );
  NOR2_X1 U15864 ( .A1(n15581), .A2(n15582), .ZN(n15816) );
  NOR2_X1 U15865 ( .A1(n8846), .A2(n9893), .ZN(n15582) );
  NAND2_X1 U15866 ( .A1(n15817), .A2(n15818), .ZN(n15581) );
  NAND2_X1 U15867 ( .A1(n15589), .A2(n15819), .ZN(n15818) );
  INV_X1 U15868 ( .A(n15820), .ZN(n15819) );
  NOR2_X1 U15869 ( .A1(n15587), .A2(n15588), .ZN(n15820) );
  NOR2_X1 U15870 ( .A1(n8846), .A2(n8512), .ZN(n15589) );
  NAND2_X1 U15871 ( .A1(n15587), .A2(n15588), .ZN(n15817) );
  NAND2_X1 U15872 ( .A1(n15821), .A2(n15822), .ZN(n15588) );
  NAND2_X1 U15873 ( .A1(n15615), .A2(n15823), .ZN(n15822) );
  INV_X1 U15874 ( .A(n15824), .ZN(n15823) );
  NOR2_X1 U15875 ( .A1(n15616), .A2(n15614), .ZN(n15824) );
  NOR2_X1 U15876 ( .A1(n8846), .A2(n8493), .ZN(n15615) );
  NAND2_X1 U15877 ( .A1(n15614), .A2(n15616), .ZN(n15821) );
  NAND2_X1 U15878 ( .A1(n15825), .A2(n15826), .ZN(n15616) );
  NAND2_X1 U15879 ( .A1(n15610), .A2(n15827), .ZN(n15826) );
  INV_X1 U15880 ( .A(n15828), .ZN(n15827) );
  NOR2_X1 U15881 ( .A1(n15611), .A2(n15612), .ZN(n15828) );
  NOR2_X1 U15882 ( .A1(n8846), .A2(n8473), .ZN(n15610) );
  NAND2_X1 U15883 ( .A1(n15612), .A2(n15611), .ZN(n15825) );
  NAND2_X1 U15884 ( .A1(n15829), .A2(n15830), .ZN(n15611) );
  NAND2_X1 U15885 ( .A1(b_3_), .A2(n15831), .ZN(n15830) );
  NAND2_X1 U15886 ( .A1(n8456), .A2(n15832), .ZN(n15831) );
  NAND2_X1 U15887 ( .A1(a_31_), .A2(n8995), .ZN(n15832) );
  NAND2_X1 U15888 ( .A1(b_4_), .A2(n15833), .ZN(n15829) );
  NAND2_X1 U15889 ( .A1(n8459), .A2(n15834), .ZN(n15833) );
  NAND2_X1 U15890 ( .A1(a_30_), .A2(n8875), .ZN(n15834) );
  NOR3_X1 U15891 ( .A1(n8846), .A2(n8979), .A3(n8995), .ZN(n15612) );
  XOR2_X1 U15892 ( .A(n15835), .B(n15836), .Z(n15614) );
  XOR2_X1 U15893 ( .A(n15837), .B(n15838), .Z(n15835) );
  XOR2_X1 U15894 ( .A(n15839), .B(n15840), .Z(n15587) );
  XOR2_X1 U15895 ( .A(n15841), .B(n15842), .Z(n15839) );
  XNOR2_X1 U15896 ( .A(n15843), .B(n15844), .ZN(n15618) );
  XNOR2_X1 U15897 ( .A(n15845), .B(n15846), .ZN(n15844) );
  XOR2_X1 U15898 ( .A(n15847), .B(n15848), .Z(n15622) );
  XNOR2_X1 U15899 ( .A(n15849), .B(n15850), .ZN(n15848) );
  XNOR2_X1 U15900 ( .A(n15851), .B(n15852), .ZN(n15626) );
  XOR2_X1 U15901 ( .A(n15853), .B(n15854), .Z(n15851) );
  XOR2_X1 U15902 ( .A(n15855), .B(n15856), .Z(n15550) );
  XOR2_X1 U15903 ( .A(n15857), .B(n15858), .Z(n15856) );
  XNOR2_X1 U15904 ( .A(n15859), .B(n15860), .ZN(n15544) );
  XNOR2_X1 U15905 ( .A(n15861), .B(n15862), .ZN(n15859) );
  XNOR2_X1 U15906 ( .A(n15863), .B(n15864), .ZN(n15536) );
  XOR2_X1 U15907 ( .A(n15865), .B(n15866), .Z(n15864) );
  XOR2_X1 U15908 ( .A(n15867), .B(n15868), .Z(n15630) );
  XNOR2_X1 U15909 ( .A(n15869), .B(n15870), .ZN(n15867) );
  XOR2_X1 U15910 ( .A(n15871), .B(n15872), .Z(n15634) );
  XOR2_X1 U15911 ( .A(n15873), .B(n15874), .Z(n15872) );
  XNOR2_X1 U15912 ( .A(n15875), .B(n15876), .ZN(n15638) );
  XOR2_X1 U15913 ( .A(n15877), .B(n15878), .Z(n15875) );
  XOR2_X1 U15914 ( .A(n15879), .B(n15880), .Z(n15642) );
  XNOR2_X1 U15915 ( .A(n15881), .B(n15882), .ZN(n15880) );
  XNOR2_X1 U15916 ( .A(n15883), .B(n15884), .ZN(n15646) );
  XOR2_X1 U15917 ( .A(n15885), .B(n15886), .Z(n15883) );
  XOR2_X1 U15918 ( .A(n15887), .B(n15888), .Z(n15650) );
  XNOR2_X1 U15919 ( .A(n15889), .B(n15890), .ZN(n15888) );
  XNOR2_X1 U15920 ( .A(n15891), .B(n15892), .ZN(n15654) );
  XOR2_X1 U15921 ( .A(n15893), .B(n15894), .Z(n15891) );
  XOR2_X1 U15922 ( .A(n15895), .B(n15896), .Z(n15658) );
  XNOR2_X1 U15923 ( .A(n15897), .B(n15898), .ZN(n15896) );
  XNOR2_X1 U15924 ( .A(n15899), .B(n15900), .ZN(n15662) );
  XOR2_X1 U15925 ( .A(n15901), .B(n15902), .Z(n15899) );
  XOR2_X1 U15926 ( .A(n15903), .B(n15904), .Z(n15666) );
  XNOR2_X1 U15927 ( .A(n15905), .B(n15906), .ZN(n15904) );
  XNOR2_X1 U15928 ( .A(n15907), .B(n15908), .ZN(n15670) );
  XOR2_X1 U15929 ( .A(n15909), .B(n15910), .Z(n15907) );
  XOR2_X1 U15930 ( .A(n15911), .B(n15912), .Z(n15482) );
  XNOR2_X1 U15931 ( .A(n15913), .B(n15914), .ZN(n15912) );
  XNOR2_X1 U15932 ( .A(n15915), .B(n15916), .ZN(n15674) );
  XOR2_X1 U15933 ( .A(n15917), .B(n15918), .Z(n15915) );
  INV_X1 U15934 ( .A(n8843), .ZN(n8926) );
  NOR2_X1 U15935 ( .A1(n8848), .A2(n8846), .ZN(n8843) );
  XNOR2_X1 U15936 ( .A(n15919), .B(n15920), .ZN(n15681) );
  XOR2_X1 U15937 ( .A(n15921), .B(n15922), .Z(n15919) );
  XNOR2_X1 U15938 ( .A(n15923), .B(n15924), .ZN(n15685) );
  XNOR2_X1 U15939 ( .A(n15925), .B(n15926), .ZN(n15924) );
  XOR2_X1 U15940 ( .A(n15927), .B(n15928), .Z(n15689) );
  XNOR2_X1 U15941 ( .A(n15929), .B(n15930), .ZN(n15928) );
  XNOR2_X1 U15942 ( .A(n15931), .B(n15932), .ZN(n15693) );
  XOR2_X1 U15943 ( .A(n15933), .B(n15934), .Z(n15932) );
  XOR2_X1 U15944 ( .A(n8807), .B(n8806), .Z(n8649) );
  INV_X1 U15945 ( .A(n8802), .ZN(n9137) );
  NAND3_X1 U15946 ( .A1(n8806), .A2(n8807), .A3(n15935), .ZN(n8802) );
  INV_X1 U15947 ( .A(n8805), .ZN(n15935) );
  NAND2_X1 U15948 ( .A1(n9136), .A2(n15936), .ZN(n8805) );
  NAND2_X1 U15949 ( .A1(n15937), .A2(n15938), .ZN(n15936) );
  INV_X1 U15950 ( .A(n15939), .ZN(n9136) );
  NOR2_X1 U15951 ( .A1(n15938), .A2(n15937), .ZN(n15939) );
  NOR2_X1 U15952 ( .A1(n15940), .A2(n15941), .ZN(n15937) );
  INV_X1 U15953 ( .A(n15942), .ZN(n15941) );
  NAND2_X1 U15954 ( .A1(n15943), .A2(n15944), .ZN(n15942) );
  NAND2_X1 U15955 ( .A1(n15945), .A2(n15946), .ZN(n15944) );
  NOR2_X1 U15956 ( .A1(n15946), .A2(n15945), .ZN(n15940) );
  XOR2_X1 U15957 ( .A(n15947), .B(n15948), .Z(n15938) );
  NAND2_X1 U15958 ( .A1(n15949), .A2(n15950), .ZN(n15947) );
  NAND2_X1 U15959 ( .A1(n15951), .A2(n15952), .ZN(n8807) );
  NAND3_X1 U15960 ( .A1(b_4_), .A2(n15953), .A3(a_0_), .ZN(n15952) );
  NAND2_X1 U15961 ( .A1(n15450), .A2(n15451), .ZN(n15953) );
  INV_X1 U15962 ( .A(n15954), .ZN(n15951) );
  NOR2_X1 U15963 ( .A1(n15450), .A2(n15451), .ZN(n15954) );
  NOR2_X1 U15964 ( .A1(n15955), .A2(n15956), .ZN(n15451) );
  INV_X1 U15965 ( .A(n15957), .ZN(n15956) );
  NAND3_X1 U15966 ( .A1(b_4_), .A2(n15958), .A3(a_1_), .ZN(n15957) );
  NAND2_X1 U15967 ( .A1(n15698), .A2(n15699), .ZN(n15958) );
  NOR2_X1 U15968 ( .A1(n15698), .A2(n15699), .ZN(n15955) );
  NOR2_X1 U15969 ( .A1(n15959), .A2(n15960), .ZN(n15699) );
  INV_X1 U15970 ( .A(n15961), .ZN(n15960) );
  NAND2_X1 U15971 ( .A1(n15934), .A2(n15962), .ZN(n15961) );
  NAND2_X1 U15972 ( .A1(n15933), .A2(n15931), .ZN(n15962) );
  NOR2_X1 U15973 ( .A1(n8998), .A2(n8995), .ZN(n15934) );
  NOR2_X1 U15974 ( .A1(n15931), .A2(n15933), .ZN(n15959) );
  NOR2_X1 U15975 ( .A1(n15963), .A2(n15964), .ZN(n15933) );
  INV_X1 U15976 ( .A(n15965), .ZN(n15964) );
  NAND2_X1 U15977 ( .A1(n15930), .A2(n15966), .ZN(n15965) );
  NAND2_X1 U15978 ( .A1(n15927), .A2(n15929), .ZN(n15966) );
  NOR2_X1 U15979 ( .A1(n8877), .A2(n8995), .ZN(n15930) );
  NOR2_X1 U15980 ( .A1(n15927), .A2(n15929), .ZN(n15963) );
  NAND2_X1 U15981 ( .A1(n15967), .A2(n15968), .ZN(n15929) );
  NAND2_X1 U15982 ( .A1(n15923), .A2(n15969), .ZN(n15968) );
  NAND2_X1 U15983 ( .A1(n15926), .A2(n15925), .ZN(n15969) );
  XOR2_X1 U15984 ( .A(n15970), .B(n15971), .Z(n15923) );
  NAND2_X1 U15985 ( .A1(n15972), .A2(n15973), .ZN(n15970) );
  INV_X1 U15986 ( .A(n15974), .ZN(n15967) );
  NOR2_X1 U15987 ( .A1(n15925), .A2(n15926), .ZN(n15974) );
  INV_X1 U15988 ( .A(n8860), .ZN(n15926) );
  NAND2_X1 U15989 ( .A1(a_4_), .A2(b_4_), .ZN(n8860) );
  NAND2_X1 U15990 ( .A1(n15975), .A2(n15976), .ZN(n15925) );
  NAND2_X1 U15991 ( .A1(n15922), .A2(n15977), .ZN(n15976) );
  INV_X1 U15992 ( .A(n15978), .ZN(n15977) );
  NOR2_X1 U15993 ( .A1(n15921), .A2(n15920), .ZN(n15978) );
  NOR2_X1 U15994 ( .A1(n8848), .A2(n8995), .ZN(n15922) );
  NAND2_X1 U15995 ( .A1(n15920), .A2(n15921), .ZN(n15975) );
  NAND2_X1 U15996 ( .A1(n15979), .A2(n15980), .ZN(n15921) );
  NAND2_X1 U15997 ( .A1(n15724), .A2(n15981), .ZN(n15980) );
  INV_X1 U15998 ( .A(n15982), .ZN(n15981) );
  NOR2_X1 U15999 ( .A1(n15721), .A2(n15723), .ZN(n15982) );
  NOR2_X1 U16000 ( .A1(n8994), .A2(n8995), .ZN(n15724) );
  NAND2_X1 U16001 ( .A1(n15721), .A2(n15723), .ZN(n15979) );
  NAND2_X1 U16002 ( .A1(n15983), .A2(n15984), .ZN(n15723) );
  NAND2_X1 U16003 ( .A1(n15918), .A2(n15985), .ZN(n15984) );
  INV_X1 U16004 ( .A(n15986), .ZN(n15985) );
  NOR2_X1 U16005 ( .A1(n15917), .A2(n15916), .ZN(n15986) );
  NOR2_X1 U16006 ( .A1(n8817), .A2(n8995), .ZN(n15918) );
  NAND2_X1 U16007 ( .A1(n15916), .A2(n15917), .ZN(n15983) );
  NAND2_X1 U16008 ( .A1(n15987), .A2(n15988), .ZN(n15917) );
  NAND2_X1 U16009 ( .A1(n15914), .A2(n15989), .ZN(n15988) );
  INV_X1 U16010 ( .A(n15990), .ZN(n15989) );
  NOR2_X1 U16011 ( .A1(n15911), .A2(n15913), .ZN(n15990) );
  NOR2_X1 U16012 ( .A1(n10513), .A2(n8995), .ZN(n15914) );
  NAND2_X1 U16013 ( .A1(n15911), .A2(n15913), .ZN(n15987) );
  NAND2_X1 U16014 ( .A1(n15991), .A2(n15992), .ZN(n15913) );
  NAND2_X1 U16015 ( .A1(n15910), .A2(n15993), .ZN(n15992) );
  INV_X1 U16016 ( .A(n15994), .ZN(n15993) );
  NOR2_X1 U16017 ( .A1(n15909), .A2(n15908), .ZN(n15994) );
  NOR2_X1 U16018 ( .A1(n8779), .A2(n8995), .ZN(n15910) );
  NAND2_X1 U16019 ( .A1(n15908), .A2(n15909), .ZN(n15991) );
  NAND2_X1 U16020 ( .A1(n15995), .A2(n15996), .ZN(n15909) );
  NAND2_X1 U16021 ( .A1(n15906), .A2(n15997), .ZN(n15996) );
  INV_X1 U16022 ( .A(n15998), .ZN(n15997) );
  NOR2_X1 U16023 ( .A1(n15903), .A2(n15905), .ZN(n15998) );
  NOR2_X1 U16024 ( .A1(n8769), .A2(n8995), .ZN(n15906) );
  NAND2_X1 U16025 ( .A1(n15903), .A2(n15905), .ZN(n15995) );
  NAND2_X1 U16026 ( .A1(n15999), .A2(n16000), .ZN(n15905) );
  NAND2_X1 U16027 ( .A1(n15902), .A2(n16001), .ZN(n16000) );
  INV_X1 U16028 ( .A(n16002), .ZN(n16001) );
  NOR2_X1 U16029 ( .A1(n15901), .A2(n15900), .ZN(n16002) );
  NOR2_X1 U16030 ( .A1(n8749), .A2(n8995), .ZN(n15902) );
  NAND2_X1 U16031 ( .A1(n15900), .A2(n15901), .ZN(n15999) );
  NAND2_X1 U16032 ( .A1(n16003), .A2(n16004), .ZN(n15901) );
  NAND2_X1 U16033 ( .A1(n15898), .A2(n16005), .ZN(n16004) );
  INV_X1 U16034 ( .A(n16006), .ZN(n16005) );
  NOR2_X1 U16035 ( .A1(n15895), .A2(n15897), .ZN(n16006) );
  NOR2_X1 U16036 ( .A1(n8739), .A2(n8995), .ZN(n15898) );
  NAND2_X1 U16037 ( .A1(n15895), .A2(n15897), .ZN(n16003) );
  NAND2_X1 U16038 ( .A1(n16007), .A2(n16008), .ZN(n15897) );
  NAND2_X1 U16039 ( .A1(n15893), .A2(n16009), .ZN(n16008) );
  INV_X1 U16040 ( .A(n16010), .ZN(n16009) );
  NOR2_X1 U16041 ( .A1(n15894), .A2(n15892), .ZN(n16010) );
  NOR2_X1 U16042 ( .A1(n8721), .A2(n8995), .ZN(n15893) );
  NAND2_X1 U16043 ( .A1(n15892), .A2(n15894), .ZN(n16007) );
  NAND2_X1 U16044 ( .A1(n16011), .A2(n16012), .ZN(n15894) );
  NAND2_X1 U16045 ( .A1(n15890), .A2(n16013), .ZN(n16012) );
  INV_X1 U16046 ( .A(n16014), .ZN(n16013) );
  NOR2_X1 U16047 ( .A1(n15889), .A2(n15887), .ZN(n16014) );
  NOR2_X1 U16048 ( .A1(n8991), .A2(n8995), .ZN(n15890) );
  NAND2_X1 U16049 ( .A1(n15887), .A2(n15889), .ZN(n16011) );
  NAND2_X1 U16050 ( .A1(n16015), .A2(n16016), .ZN(n15889) );
  NAND2_X1 U16051 ( .A1(n15886), .A2(n16017), .ZN(n16016) );
  INV_X1 U16052 ( .A(n16018), .ZN(n16017) );
  NOR2_X1 U16053 ( .A1(n15885), .A2(n15884), .ZN(n16018) );
  NOR2_X1 U16054 ( .A1(n8692), .A2(n8995), .ZN(n15886) );
  NAND2_X1 U16055 ( .A1(n15884), .A2(n15885), .ZN(n16015) );
  NAND2_X1 U16056 ( .A1(n16019), .A2(n16020), .ZN(n15885) );
  NAND2_X1 U16057 ( .A1(n15882), .A2(n16021), .ZN(n16020) );
  INV_X1 U16058 ( .A(n16022), .ZN(n16021) );
  NOR2_X1 U16059 ( .A1(n15879), .A2(n15881), .ZN(n16022) );
  NOR2_X1 U16060 ( .A1(n8680), .A2(n8995), .ZN(n15882) );
  NAND2_X1 U16061 ( .A1(n15879), .A2(n15881), .ZN(n16019) );
  NAND2_X1 U16062 ( .A1(n16023), .A2(n16024), .ZN(n15881) );
  NAND2_X1 U16063 ( .A1(n15878), .A2(n16025), .ZN(n16024) );
  INV_X1 U16064 ( .A(n16026), .ZN(n16025) );
  NOR2_X1 U16065 ( .A1(n15877), .A2(n15876), .ZN(n16026) );
  NOR2_X1 U16066 ( .A1(n8662), .A2(n8995), .ZN(n15878) );
  NAND2_X1 U16067 ( .A1(n15876), .A2(n15877), .ZN(n16023) );
  NAND2_X1 U16068 ( .A1(n16027), .A2(n16028), .ZN(n15877) );
  NAND2_X1 U16069 ( .A1(n15874), .A2(n16029), .ZN(n16028) );
  NAND2_X1 U16070 ( .A1(n16030), .A2(n15873), .ZN(n16029) );
  INV_X1 U16071 ( .A(n15871), .ZN(n16030) );
  NOR2_X1 U16072 ( .A1(n8988), .A2(n8995), .ZN(n15874) );
  NAND2_X1 U16073 ( .A1(n15871), .A2(n16031), .ZN(n16027) );
  INV_X1 U16074 ( .A(n15873), .ZN(n16031) );
  NOR2_X1 U16075 ( .A1(n16032), .A2(n16033), .ZN(n15873) );
  INV_X1 U16076 ( .A(n16034), .ZN(n16033) );
  NAND2_X1 U16077 ( .A1(n15870), .A2(n16035), .ZN(n16034) );
  NAND2_X1 U16078 ( .A1(n15869), .A2(n15868), .ZN(n16035) );
  NOR2_X1 U16079 ( .A1(n8995), .A2(n8630), .ZN(n15870) );
  NOR2_X1 U16080 ( .A1(n15868), .A2(n15869), .ZN(n16032) );
  NOR2_X1 U16081 ( .A1(n16036), .A2(n16037), .ZN(n15869) );
  INV_X1 U16082 ( .A(n16038), .ZN(n16037) );
  NAND2_X1 U16083 ( .A1(n15866), .A2(n16039), .ZN(n16038) );
  NAND2_X1 U16084 ( .A1(n15863), .A2(n15865), .ZN(n16039) );
  NOR2_X1 U16085 ( .A1(n8995), .A2(n8986), .ZN(n15866) );
  NOR2_X1 U16086 ( .A1(n15863), .A2(n15865), .ZN(n16036) );
  NOR2_X1 U16087 ( .A1(n16040), .A2(n16041), .ZN(n15865) );
  INV_X1 U16088 ( .A(n16042), .ZN(n16041) );
  NAND2_X1 U16089 ( .A1(n15861), .A2(n16043), .ZN(n16042) );
  NAND2_X1 U16090 ( .A1(n15862), .A2(n15860), .ZN(n16043) );
  NOR2_X1 U16091 ( .A1(n8995), .A2(n8601), .ZN(n15861) );
  NOR2_X1 U16092 ( .A1(n15860), .A2(n15862), .ZN(n16040) );
  NOR2_X1 U16093 ( .A1(n16044), .A2(n16045), .ZN(n15862) );
  NOR2_X1 U16094 ( .A1(n15858), .A2(n16046), .ZN(n16045) );
  NOR2_X1 U16095 ( .A1(n15857), .A2(n15855), .ZN(n16046) );
  NAND2_X1 U16096 ( .A1(b_4_), .A2(a_22_), .ZN(n15858) );
  INV_X1 U16097 ( .A(n16047), .ZN(n16044) );
  NAND2_X1 U16098 ( .A1(n15855), .A2(n15857), .ZN(n16047) );
  NAND2_X1 U16099 ( .A1(n16048), .A2(n16049), .ZN(n15857) );
  NAND2_X1 U16100 ( .A1(n15854), .A2(n16050), .ZN(n16049) );
  INV_X1 U16101 ( .A(n16051), .ZN(n16050) );
  NOR2_X1 U16102 ( .A1(n15852), .A2(n15853), .ZN(n16051) );
  NOR2_X1 U16103 ( .A1(n8995), .A2(n8572), .ZN(n15854) );
  NAND2_X1 U16104 ( .A1(n15852), .A2(n15853), .ZN(n16048) );
  NAND2_X1 U16105 ( .A1(n16052), .A2(n16053), .ZN(n15853) );
  NAND2_X1 U16106 ( .A1(n15799), .A2(n16054), .ZN(n16053) );
  NAND2_X1 U16107 ( .A1(n15797), .A2(n15798), .ZN(n16054) );
  NOR2_X1 U16108 ( .A1(n8995), .A2(n8982), .ZN(n15799) );
  INV_X1 U16109 ( .A(n16055), .ZN(n16052) );
  NOR2_X1 U16110 ( .A1(n15797), .A2(n15798), .ZN(n16055) );
  NOR2_X1 U16111 ( .A1(n16056), .A2(n16057), .ZN(n15798) );
  INV_X1 U16112 ( .A(n16058), .ZN(n16057) );
  NAND2_X1 U16113 ( .A1(n15850), .A2(n16059), .ZN(n16058) );
  NAND2_X1 U16114 ( .A1(n15847), .A2(n15849), .ZN(n16059) );
  NOR2_X1 U16115 ( .A1(n8995), .A2(n8541), .ZN(n15850) );
  NOR2_X1 U16116 ( .A1(n15849), .A2(n15847), .ZN(n16056) );
  XOR2_X1 U16117 ( .A(n16060), .B(n16061), .Z(n15847) );
  XNOR2_X1 U16118 ( .A(n16062), .B(n16063), .ZN(n16061) );
  NAND2_X1 U16119 ( .A1(n16064), .A2(n16065), .ZN(n15849) );
  NAND2_X1 U16120 ( .A1(n15843), .A2(n16066), .ZN(n16065) );
  INV_X1 U16121 ( .A(n16067), .ZN(n16066) );
  NOR2_X1 U16122 ( .A1(n15846), .A2(n15845), .ZN(n16067) );
  XOR2_X1 U16123 ( .A(n16068), .B(n16069), .Z(n15843) );
  XNOR2_X1 U16124 ( .A(n16070), .B(n16071), .ZN(n16068) );
  NAND2_X1 U16125 ( .A1(n15845), .A2(n15846), .ZN(n16064) );
  NAND2_X1 U16126 ( .A1(b_4_), .A2(a_26_), .ZN(n15846) );
  NOR2_X1 U16127 ( .A1(n16072), .A2(n16073), .ZN(n15845) );
  NOR3_X1 U16128 ( .A1(n8512), .A2(n16074), .A3(n8995), .ZN(n16073) );
  NOR2_X1 U16129 ( .A1(n15813), .A2(n15814), .ZN(n16074) );
  INV_X1 U16130 ( .A(n16075), .ZN(n16072) );
  NAND2_X1 U16131 ( .A1(n15813), .A2(n15814), .ZN(n16075) );
  NAND2_X1 U16132 ( .A1(n16076), .A2(n16077), .ZN(n15814) );
  NAND2_X1 U16133 ( .A1(n15841), .A2(n16078), .ZN(n16077) );
  INV_X1 U16134 ( .A(n16079), .ZN(n16078) );
  NOR2_X1 U16135 ( .A1(n15842), .A2(n15840), .ZN(n16079) );
  NOR2_X1 U16136 ( .A1(n8995), .A2(n8493), .ZN(n15841) );
  NAND2_X1 U16137 ( .A1(n15840), .A2(n15842), .ZN(n16076) );
  NAND2_X1 U16138 ( .A1(n16080), .A2(n16081), .ZN(n15842) );
  NAND2_X1 U16139 ( .A1(n15836), .A2(n16082), .ZN(n16081) );
  INV_X1 U16140 ( .A(n16083), .ZN(n16082) );
  NOR2_X1 U16141 ( .A1(n15837), .A2(n15838), .ZN(n16083) );
  NOR2_X1 U16142 ( .A1(n8995), .A2(n8473), .ZN(n15836) );
  NAND2_X1 U16143 ( .A1(n15838), .A2(n15837), .ZN(n16080) );
  NAND2_X1 U16144 ( .A1(n16084), .A2(n16085), .ZN(n15837) );
  NAND2_X1 U16145 ( .A1(b_2_), .A2(n16086), .ZN(n16085) );
  NAND2_X1 U16146 ( .A1(n8456), .A2(n16087), .ZN(n16086) );
  NAND2_X1 U16147 ( .A1(a_31_), .A2(n8875), .ZN(n16087) );
  NAND2_X1 U16148 ( .A1(b_3_), .A2(n16088), .ZN(n16084) );
  NAND2_X1 U16149 ( .A1(n8459), .A2(n16089), .ZN(n16088) );
  NAND2_X1 U16150 ( .A1(a_30_), .A2(n8997), .ZN(n16089) );
  NOR3_X1 U16151 ( .A1(n8995), .A2(n8979), .A3(n8875), .ZN(n15838) );
  XOR2_X1 U16152 ( .A(n16090), .B(n16091), .Z(n15840) );
  XNOR2_X1 U16153 ( .A(n16092), .B(n16093), .ZN(n16090) );
  XNOR2_X1 U16154 ( .A(n16094), .B(n16095), .ZN(n15813) );
  XNOR2_X1 U16155 ( .A(n16096), .B(n16097), .ZN(n16094) );
  XOR2_X1 U16156 ( .A(n16098), .B(n16099), .Z(n15797) );
  NAND2_X1 U16157 ( .A1(n16100), .A2(n16101), .ZN(n16098) );
  XOR2_X1 U16158 ( .A(n16102), .B(n16103), .Z(n15852) );
  XOR2_X1 U16159 ( .A(n16104), .B(n16105), .Z(n16102) );
  NOR2_X1 U16160 ( .A1(n8982), .A2(n8875), .ZN(n16105) );
  XNOR2_X1 U16161 ( .A(n16106), .B(n16107), .ZN(n15855) );
  NAND2_X1 U16162 ( .A1(n16108), .A2(n16109), .ZN(n16106) );
  XNOR2_X1 U16163 ( .A(n16110), .B(n16111), .ZN(n15860) );
  XOR2_X1 U16164 ( .A(n16112), .B(n16113), .Z(n16110) );
  NOR2_X1 U16165 ( .A1(n8984), .A2(n8875), .ZN(n16113) );
  XOR2_X1 U16166 ( .A(n16114), .B(n16115), .Z(n15863) );
  NAND2_X1 U16167 ( .A1(n16116), .A2(n16117), .ZN(n16114) );
  XNOR2_X1 U16168 ( .A(n16118), .B(n16119), .ZN(n15868) );
  XOR2_X1 U16169 ( .A(n16120), .B(n16121), .Z(n16118) );
  NOR2_X1 U16170 ( .A1(n8986), .A2(n8875), .ZN(n16121) );
  XNOR2_X1 U16171 ( .A(n16122), .B(n16123), .ZN(n15871) );
  NAND2_X1 U16172 ( .A1(n16124), .A2(n16125), .ZN(n16122) );
  XOR2_X1 U16173 ( .A(n16126), .B(n16127), .Z(n15876) );
  XOR2_X1 U16174 ( .A(n16128), .B(n16129), .Z(n16126) );
  NOR2_X1 U16175 ( .A1(n8875), .A2(n8988), .ZN(n16129) );
  XNOR2_X1 U16176 ( .A(n16130), .B(n16131), .ZN(n15879) );
  NAND2_X1 U16177 ( .A1(n16132), .A2(n16133), .ZN(n16130) );
  XOR2_X1 U16178 ( .A(n16134), .B(n16135), .Z(n15884) );
  XOR2_X1 U16179 ( .A(n16136), .B(n16137), .Z(n16134) );
  NOR2_X1 U16180 ( .A1(n8875), .A2(n8680), .ZN(n16137) );
  XNOR2_X1 U16181 ( .A(n16138), .B(n16139), .ZN(n15887) );
  NAND2_X1 U16182 ( .A1(n16140), .A2(n16141), .ZN(n16138) );
  XOR2_X1 U16183 ( .A(n16142), .B(n16143), .Z(n15892) );
  XOR2_X1 U16184 ( .A(n16144), .B(n16145), .Z(n16142) );
  NOR2_X1 U16185 ( .A1(n8875), .A2(n8991), .ZN(n16145) );
  XNOR2_X1 U16186 ( .A(n16146), .B(n16147), .ZN(n15895) );
  NAND2_X1 U16187 ( .A1(n16148), .A2(n16149), .ZN(n16146) );
  XOR2_X1 U16188 ( .A(n16150), .B(n16151), .Z(n15900) );
  XOR2_X1 U16189 ( .A(n16152), .B(n16153), .Z(n16150) );
  NOR2_X1 U16190 ( .A1(n8875), .A2(n8739), .ZN(n16153) );
  XNOR2_X1 U16191 ( .A(n16154), .B(n16155), .ZN(n15903) );
  NAND2_X1 U16192 ( .A1(n16156), .A2(n16157), .ZN(n16154) );
  XOR2_X1 U16193 ( .A(n16158), .B(n16159), .Z(n15908) );
  XOR2_X1 U16194 ( .A(n16160), .B(n16161), .Z(n16158) );
  NOR2_X1 U16195 ( .A1(n8875), .A2(n8769), .ZN(n16161) );
  XNOR2_X1 U16196 ( .A(n16162), .B(n16163), .ZN(n15911) );
  NAND2_X1 U16197 ( .A1(n16164), .A2(n16165), .ZN(n16162) );
  XOR2_X1 U16198 ( .A(n16166), .B(n16167), .Z(n15916) );
  XOR2_X1 U16199 ( .A(n16168), .B(n16169), .Z(n16166) );
  NOR2_X1 U16200 ( .A1(n8875), .A2(n10513), .ZN(n16169) );
  XNOR2_X1 U16201 ( .A(n16170), .B(n16171), .ZN(n15721) );
  NAND2_X1 U16202 ( .A1(n16172), .A2(n16173), .ZN(n16170) );
  XOR2_X1 U16203 ( .A(n16174), .B(n16175), .Z(n15920) );
  XOR2_X1 U16204 ( .A(n16176), .B(n16177), .Z(n16174) );
  NOR2_X1 U16205 ( .A1(n8875), .A2(n8994), .ZN(n16177) );
  XNOR2_X1 U16206 ( .A(n16178), .B(n16179), .ZN(n15927) );
  XOR2_X1 U16207 ( .A(n16180), .B(n16181), .Z(n16178) );
  NOR2_X1 U16208 ( .A1(n8875), .A2(n8996), .ZN(n16181) );
  XOR2_X1 U16209 ( .A(n16182), .B(n16183), .Z(n15931) );
  XNOR2_X1 U16210 ( .A(n16184), .B(n8872), .ZN(n16182) );
  XOR2_X1 U16211 ( .A(n16185), .B(n16186), .Z(n15698) );
  XOR2_X1 U16212 ( .A(n16187), .B(n16188), .Z(n16186) );
  NAND2_X1 U16213 ( .A1(a_2_), .A2(b_3_), .ZN(n16188) );
  XOR2_X1 U16214 ( .A(n16189), .B(n16190), .Z(n15450) );
  NAND2_X1 U16215 ( .A1(n16191), .A2(n16192), .ZN(n16189) );
  XNOR2_X1 U16216 ( .A(n16193), .B(n15946), .ZN(n8806) );
  XOR2_X1 U16217 ( .A(n16194), .B(n16195), .Z(n15946) );
  XNOR2_X1 U16218 ( .A(n16196), .B(n16197), .ZN(n16195) );
  NOR2_X1 U16219 ( .A1(n8997), .A2(n9731), .ZN(n16197) );
  XNOR2_X1 U16220 ( .A(n15945), .B(n15943), .ZN(n16193) );
  NOR2_X1 U16221 ( .A1(n9471), .A2(n8875), .ZN(n15943) );
  INV_X1 U16222 ( .A(n16198), .ZN(n15945) );
  NAND2_X1 U16223 ( .A1(n16191), .A2(n16199), .ZN(n16198) );
  NAND2_X1 U16224 ( .A1(n16190), .A2(n16192), .ZN(n16199) );
  NAND2_X1 U16225 ( .A1(n16200), .A2(n16201), .ZN(n16192) );
  NAND2_X1 U16226 ( .A1(a_1_), .A2(b_3_), .ZN(n16201) );
  XNOR2_X1 U16227 ( .A(n16202), .B(n16203), .ZN(n16190) );
  XOR2_X1 U16228 ( .A(n16204), .B(n8889), .Z(n16202) );
  INV_X1 U16229 ( .A(n16205), .ZN(n16191) );
  NOR2_X1 U16230 ( .A1(n9731), .A2(n16200), .ZN(n16205) );
  NOR2_X1 U16231 ( .A1(n16206), .A2(n16207), .ZN(n16200) );
  NOR3_X1 U16232 ( .A1(n8875), .A2(n16208), .A3(n8998), .ZN(n16207) );
  INV_X1 U16233 ( .A(n16209), .ZN(n16208) );
  NAND2_X1 U16234 ( .A1(n16185), .A2(n16187), .ZN(n16209) );
  NOR2_X1 U16235 ( .A1(n16187), .A2(n16185), .ZN(n16206) );
  XOR2_X1 U16236 ( .A(n16210), .B(n16211), .Z(n16185) );
  XNOR2_X1 U16237 ( .A(n16212), .B(n16213), .ZN(n16210) );
  NAND2_X1 U16238 ( .A1(n16214), .A2(n16215), .ZN(n16187) );
  NAND2_X1 U16239 ( .A1(n16183), .A2(n16216), .ZN(n16215) );
  NAND2_X1 U16240 ( .A1(n8872), .A2(n16217), .ZN(n16216) );
  XOR2_X1 U16241 ( .A(n16218), .B(n16219), .Z(n16183) );
  XNOR2_X1 U16242 ( .A(n16220), .B(n16221), .ZN(n16218) );
  NAND2_X1 U16243 ( .A1(n16184), .A2(n8922), .ZN(n16214) );
  INV_X1 U16244 ( .A(n8872), .ZN(n8922) );
  NOR2_X1 U16245 ( .A1(n8877), .A2(n8875), .ZN(n8872) );
  INV_X1 U16246 ( .A(n16217), .ZN(n16184) );
  NAND2_X1 U16247 ( .A1(n16222), .A2(n16223), .ZN(n16217) );
  NAND3_X1 U16248 ( .A1(b_3_), .A2(n16224), .A3(a_4_), .ZN(n16223) );
  INV_X1 U16249 ( .A(n16225), .ZN(n16224) );
  NOR2_X1 U16250 ( .A1(n16179), .A2(n16180), .ZN(n16225) );
  NAND2_X1 U16251 ( .A1(n16179), .A2(n16180), .ZN(n16222) );
  NAND2_X1 U16252 ( .A1(n15972), .A2(n16226), .ZN(n16180) );
  NAND2_X1 U16253 ( .A1(n15971), .A2(n15973), .ZN(n16226) );
  NAND2_X1 U16254 ( .A1(n16227), .A2(n16228), .ZN(n15973) );
  NAND2_X1 U16255 ( .A1(a_5_), .A2(b_3_), .ZN(n16228) );
  XNOR2_X1 U16256 ( .A(n16229), .B(n16230), .ZN(n15971) );
  XNOR2_X1 U16257 ( .A(n16231), .B(n16232), .ZN(n16229) );
  NAND2_X1 U16258 ( .A1(a_5_), .A2(n16233), .ZN(n15972) );
  INV_X1 U16259 ( .A(n16227), .ZN(n16233) );
  NOR2_X1 U16260 ( .A1(n16234), .A2(n16235), .ZN(n16227) );
  NOR3_X1 U16261 ( .A1(n8875), .A2(n16236), .A3(n8994), .ZN(n16235) );
  NOR2_X1 U16262 ( .A1(n16175), .A2(n16176), .ZN(n16236) );
  INV_X1 U16263 ( .A(n16237), .ZN(n16234) );
  NAND2_X1 U16264 ( .A1(n16175), .A2(n16176), .ZN(n16237) );
  NAND2_X1 U16265 ( .A1(n16172), .A2(n16238), .ZN(n16176) );
  NAND2_X1 U16266 ( .A1(n16171), .A2(n16173), .ZN(n16238) );
  NAND2_X1 U16267 ( .A1(n16239), .A2(n16240), .ZN(n16173) );
  NAND2_X1 U16268 ( .A1(a_7_), .A2(b_3_), .ZN(n16240) );
  XNOR2_X1 U16269 ( .A(n16241), .B(n16242), .ZN(n16171) );
  XNOR2_X1 U16270 ( .A(n16243), .B(n16244), .ZN(n16241) );
  NAND2_X1 U16271 ( .A1(a_7_), .A2(n16245), .ZN(n16172) );
  INV_X1 U16272 ( .A(n16239), .ZN(n16245) );
  NOR2_X1 U16273 ( .A1(n16246), .A2(n16247), .ZN(n16239) );
  NOR3_X1 U16274 ( .A1(n8875), .A2(n16248), .A3(n10513), .ZN(n16247) );
  NOR2_X1 U16275 ( .A1(n16167), .A2(n16168), .ZN(n16248) );
  INV_X1 U16276 ( .A(n16249), .ZN(n16246) );
  NAND2_X1 U16277 ( .A1(n16167), .A2(n16168), .ZN(n16249) );
  NAND2_X1 U16278 ( .A1(n16164), .A2(n16250), .ZN(n16168) );
  NAND2_X1 U16279 ( .A1(n16163), .A2(n16165), .ZN(n16250) );
  NAND2_X1 U16280 ( .A1(n16251), .A2(n16252), .ZN(n16165) );
  NAND2_X1 U16281 ( .A1(a_9_), .A2(b_3_), .ZN(n16252) );
  INV_X1 U16282 ( .A(n16253), .ZN(n16251) );
  XNOR2_X1 U16283 ( .A(n16254), .B(n16255), .ZN(n16163) );
  XNOR2_X1 U16284 ( .A(n16256), .B(n16257), .ZN(n16254) );
  NAND2_X1 U16285 ( .A1(a_9_), .A2(n16253), .ZN(n16164) );
  NAND2_X1 U16286 ( .A1(n16258), .A2(n16259), .ZN(n16253) );
  INV_X1 U16287 ( .A(n16260), .ZN(n16259) );
  NOR3_X1 U16288 ( .A1(n8875), .A2(n16261), .A3(n8769), .ZN(n16260) );
  NOR2_X1 U16289 ( .A1(n16159), .A2(n16160), .ZN(n16261) );
  NAND2_X1 U16290 ( .A1(n16159), .A2(n16160), .ZN(n16258) );
  NAND2_X1 U16291 ( .A1(n16156), .A2(n16262), .ZN(n16160) );
  NAND2_X1 U16292 ( .A1(n16155), .A2(n16157), .ZN(n16262) );
  NAND2_X1 U16293 ( .A1(n16263), .A2(n16264), .ZN(n16157) );
  NAND2_X1 U16294 ( .A1(a_11_), .A2(b_3_), .ZN(n16264) );
  INV_X1 U16295 ( .A(n16265), .ZN(n16263) );
  XNOR2_X1 U16296 ( .A(n16266), .B(n16267), .ZN(n16155) );
  XNOR2_X1 U16297 ( .A(n16268), .B(n16269), .ZN(n16266) );
  NAND2_X1 U16298 ( .A1(a_11_), .A2(n16265), .ZN(n16156) );
  NAND2_X1 U16299 ( .A1(n16270), .A2(n16271), .ZN(n16265) );
  INV_X1 U16300 ( .A(n16272), .ZN(n16271) );
  NOR3_X1 U16301 ( .A1(n8875), .A2(n16273), .A3(n8739), .ZN(n16272) );
  NOR2_X1 U16302 ( .A1(n16151), .A2(n16152), .ZN(n16273) );
  NAND2_X1 U16303 ( .A1(n16151), .A2(n16152), .ZN(n16270) );
  NAND2_X1 U16304 ( .A1(n16148), .A2(n16274), .ZN(n16152) );
  NAND2_X1 U16305 ( .A1(n16147), .A2(n16149), .ZN(n16274) );
  NAND2_X1 U16306 ( .A1(n16275), .A2(n16276), .ZN(n16149) );
  NAND2_X1 U16307 ( .A1(a_13_), .A2(b_3_), .ZN(n16276) );
  INV_X1 U16308 ( .A(n16277), .ZN(n16275) );
  XNOR2_X1 U16309 ( .A(n16278), .B(n16279), .ZN(n16147) );
  XNOR2_X1 U16310 ( .A(n16280), .B(n16281), .ZN(n16278) );
  NAND2_X1 U16311 ( .A1(a_13_), .A2(n16277), .ZN(n16148) );
  NAND2_X1 U16312 ( .A1(n16282), .A2(n16283), .ZN(n16277) );
  INV_X1 U16313 ( .A(n16284), .ZN(n16283) );
  NOR3_X1 U16314 ( .A1(n8875), .A2(n16285), .A3(n8991), .ZN(n16284) );
  NOR2_X1 U16315 ( .A1(n16143), .A2(n16144), .ZN(n16285) );
  NAND2_X1 U16316 ( .A1(n16143), .A2(n16144), .ZN(n16282) );
  NAND2_X1 U16317 ( .A1(n16140), .A2(n16286), .ZN(n16144) );
  NAND2_X1 U16318 ( .A1(n16139), .A2(n16141), .ZN(n16286) );
  NAND2_X1 U16319 ( .A1(n16287), .A2(n16288), .ZN(n16141) );
  NAND2_X1 U16320 ( .A1(a_15_), .A2(b_3_), .ZN(n16288) );
  INV_X1 U16321 ( .A(n16289), .ZN(n16287) );
  XNOR2_X1 U16322 ( .A(n16290), .B(n16291), .ZN(n16139) );
  XNOR2_X1 U16323 ( .A(n16292), .B(n16293), .ZN(n16291) );
  NAND2_X1 U16324 ( .A1(a_15_), .A2(n16289), .ZN(n16140) );
  NAND2_X1 U16325 ( .A1(n16294), .A2(n16295), .ZN(n16289) );
  INV_X1 U16326 ( .A(n16296), .ZN(n16295) );
  NOR3_X1 U16327 ( .A1(n8875), .A2(n16297), .A3(n8680), .ZN(n16296) );
  NOR2_X1 U16328 ( .A1(n16135), .A2(n16136), .ZN(n16297) );
  NAND2_X1 U16329 ( .A1(n16135), .A2(n16136), .ZN(n16294) );
  NAND2_X1 U16330 ( .A1(n16132), .A2(n16298), .ZN(n16136) );
  NAND2_X1 U16331 ( .A1(n16131), .A2(n16133), .ZN(n16298) );
  NAND2_X1 U16332 ( .A1(n16299), .A2(n16300), .ZN(n16133) );
  NAND2_X1 U16333 ( .A1(a_17_), .A2(b_3_), .ZN(n16300) );
  INV_X1 U16334 ( .A(n16301), .ZN(n16299) );
  XNOR2_X1 U16335 ( .A(n16302), .B(n16303), .ZN(n16131) );
  XNOR2_X1 U16336 ( .A(n16304), .B(n16305), .ZN(n16303) );
  NAND2_X1 U16337 ( .A1(a_17_), .A2(n16301), .ZN(n16132) );
  NAND2_X1 U16338 ( .A1(n16306), .A2(n16307), .ZN(n16301) );
  INV_X1 U16339 ( .A(n16308), .ZN(n16307) );
  NOR3_X1 U16340 ( .A1(n8875), .A2(n16309), .A3(n8988), .ZN(n16308) );
  NOR2_X1 U16341 ( .A1(n16127), .A2(n16128), .ZN(n16309) );
  NAND2_X1 U16342 ( .A1(n16127), .A2(n16128), .ZN(n16306) );
  NAND2_X1 U16343 ( .A1(n16124), .A2(n16310), .ZN(n16128) );
  NAND2_X1 U16344 ( .A1(n16123), .A2(n16125), .ZN(n16310) );
  NAND2_X1 U16345 ( .A1(n16311), .A2(n16312), .ZN(n16125) );
  NAND2_X1 U16346 ( .A1(b_3_), .A2(a_19_), .ZN(n16312) );
  INV_X1 U16347 ( .A(n16313), .ZN(n16311) );
  XNOR2_X1 U16348 ( .A(n16314), .B(n16315), .ZN(n16123) );
  XNOR2_X1 U16349 ( .A(n16316), .B(n16317), .ZN(n16315) );
  NAND2_X1 U16350 ( .A1(a_19_), .A2(n16313), .ZN(n16124) );
  NAND2_X1 U16351 ( .A1(n16318), .A2(n16319), .ZN(n16313) );
  INV_X1 U16352 ( .A(n16320), .ZN(n16319) );
  NOR3_X1 U16353 ( .A1(n8986), .A2(n16321), .A3(n8875), .ZN(n16320) );
  NOR2_X1 U16354 ( .A1(n16119), .A2(n16120), .ZN(n16321) );
  NAND2_X1 U16355 ( .A1(n16119), .A2(n16120), .ZN(n16318) );
  NAND2_X1 U16356 ( .A1(n16116), .A2(n16322), .ZN(n16120) );
  NAND2_X1 U16357 ( .A1(n16115), .A2(n16117), .ZN(n16322) );
  NAND2_X1 U16358 ( .A1(n16323), .A2(n16324), .ZN(n16117) );
  NAND2_X1 U16359 ( .A1(b_3_), .A2(a_21_), .ZN(n16324) );
  INV_X1 U16360 ( .A(n16325), .ZN(n16323) );
  XNOR2_X1 U16361 ( .A(n16326), .B(n16327), .ZN(n16115) );
  XOR2_X1 U16362 ( .A(n16328), .B(n16329), .Z(n16327) );
  NAND2_X1 U16363 ( .A1(a_21_), .A2(n16325), .ZN(n16116) );
  NAND2_X1 U16364 ( .A1(n16330), .A2(n16331), .ZN(n16325) );
  INV_X1 U16365 ( .A(n16332), .ZN(n16331) );
  NOR3_X1 U16366 ( .A1(n8984), .A2(n16333), .A3(n8875), .ZN(n16332) );
  NOR2_X1 U16367 ( .A1(n16111), .A2(n16112), .ZN(n16333) );
  NAND2_X1 U16368 ( .A1(n16111), .A2(n16112), .ZN(n16330) );
  NAND2_X1 U16369 ( .A1(n16108), .A2(n16334), .ZN(n16112) );
  NAND2_X1 U16370 ( .A1(n16107), .A2(n16109), .ZN(n16334) );
  NAND2_X1 U16371 ( .A1(n16335), .A2(n16336), .ZN(n16109) );
  NAND2_X1 U16372 ( .A1(b_3_), .A2(a_23_), .ZN(n16336) );
  XNOR2_X1 U16373 ( .A(n16337), .B(n16338), .ZN(n16107) );
  NAND2_X1 U16374 ( .A1(n16339), .A2(n16340), .ZN(n16337) );
  INV_X1 U16375 ( .A(n16341), .ZN(n16108) );
  NOR2_X1 U16376 ( .A1(n8572), .A2(n16335), .ZN(n16341) );
  NOR2_X1 U16377 ( .A1(n16342), .A2(n16343), .ZN(n16335) );
  NOR3_X1 U16378 ( .A1(n8982), .A2(n16344), .A3(n8875), .ZN(n16343) );
  NOR2_X1 U16379 ( .A1(n16104), .A2(n16103), .ZN(n16344) );
  INV_X1 U16380 ( .A(n16345), .ZN(n16342) );
  NAND2_X1 U16381 ( .A1(n16103), .A2(n16104), .ZN(n16345) );
  NAND2_X1 U16382 ( .A1(n16100), .A2(n16346), .ZN(n16104) );
  NAND2_X1 U16383 ( .A1(n16099), .A2(n16101), .ZN(n16346) );
  NAND2_X1 U16384 ( .A1(n16347), .A2(n16348), .ZN(n16101) );
  NAND2_X1 U16385 ( .A1(b_3_), .A2(a_25_), .ZN(n16348) );
  INV_X1 U16386 ( .A(n16349), .ZN(n16347) );
  XNOR2_X1 U16387 ( .A(n16350), .B(n16351), .ZN(n16099) );
  XNOR2_X1 U16388 ( .A(n16352), .B(n16353), .ZN(n16351) );
  NOR2_X1 U16389 ( .A1(n9893), .A2(n8997), .ZN(n16353) );
  NAND2_X1 U16390 ( .A1(a_25_), .A2(n16349), .ZN(n16100) );
  NAND2_X1 U16391 ( .A1(n16354), .A2(n16355), .ZN(n16349) );
  NAND2_X1 U16392 ( .A1(n16063), .A2(n16356), .ZN(n16355) );
  INV_X1 U16393 ( .A(n16357), .ZN(n16356) );
  NOR2_X1 U16394 ( .A1(n16062), .A2(n16060), .ZN(n16357) );
  NOR2_X1 U16395 ( .A1(n8875), .A2(n9893), .ZN(n16063) );
  NAND2_X1 U16396 ( .A1(n16060), .A2(n16062), .ZN(n16354) );
  NAND2_X1 U16397 ( .A1(n16358), .A2(n16359), .ZN(n16062) );
  NAND2_X1 U16398 ( .A1(n16071), .A2(n16360), .ZN(n16359) );
  NAND2_X1 U16399 ( .A1(n16070), .A2(n16069), .ZN(n16360) );
  NOR2_X1 U16400 ( .A1(n8875), .A2(n8512), .ZN(n16071) );
  INV_X1 U16401 ( .A(n16361), .ZN(n16358) );
  NOR2_X1 U16402 ( .A1(n16069), .A2(n16070), .ZN(n16361) );
  NOR2_X1 U16403 ( .A1(n16362), .A2(n16363), .ZN(n16070) );
  INV_X1 U16404 ( .A(n16364), .ZN(n16363) );
  NAND2_X1 U16405 ( .A1(n16096), .A2(n16365), .ZN(n16364) );
  NAND2_X1 U16406 ( .A1(n16097), .A2(n16095), .ZN(n16365) );
  NOR2_X1 U16407 ( .A1(n8875), .A2(n8493), .ZN(n16096) );
  NOR2_X1 U16408 ( .A1(n16095), .A2(n16097), .ZN(n16362) );
  NOR2_X1 U16409 ( .A1(n16366), .A2(n16367), .ZN(n16097) );
  INV_X1 U16410 ( .A(n16368), .ZN(n16367) );
  NAND2_X1 U16411 ( .A1(n16091), .A2(n16369), .ZN(n16368) );
  NAND2_X1 U16412 ( .A1(n16370), .A2(n16093), .ZN(n16369) );
  NOR2_X1 U16413 ( .A1(n8875), .A2(n8473), .ZN(n16091) );
  NOR2_X1 U16414 ( .A1(n16093), .A2(n16370), .ZN(n16366) );
  INV_X1 U16415 ( .A(n16092), .ZN(n16370) );
  NAND2_X1 U16416 ( .A1(n16371), .A2(n16372), .ZN(n16092) );
  NAND2_X1 U16417 ( .A1(b_1_), .A2(n16373), .ZN(n16372) );
  NAND2_X1 U16418 ( .A1(n8456), .A2(n16374), .ZN(n16373) );
  NAND2_X1 U16419 ( .A1(a_31_), .A2(n8997), .ZN(n16374) );
  NAND2_X1 U16420 ( .A1(b_2_), .A2(n16375), .ZN(n16371) );
  NAND2_X1 U16421 ( .A1(n8459), .A2(n16376), .ZN(n16375) );
  NAND2_X1 U16422 ( .A1(a_30_), .A2(n8907), .ZN(n16376) );
  NAND3_X1 U16423 ( .A1(b_3_), .A2(n9666), .A3(b_2_), .ZN(n16093) );
  XNOR2_X1 U16424 ( .A(n16377), .B(n16378), .ZN(n16095) );
  XOR2_X1 U16425 ( .A(n16379), .B(n16380), .Z(n16377) );
  XNOR2_X1 U16426 ( .A(n16381), .B(n16382), .ZN(n16069) );
  XNOR2_X1 U16427 ( .A(n16383), .B(n16384), .ZN(n16381) );
  NAND2_X1 U16428 ( .A1(b_2_), .A2(a_28_), .ZN(n16383) );
  XNOR2_X1 U16429 ( .A(n16385), .B(n16386), .ZN(n16060) );
  NAND2_X1 U16430 ( .A1(n16387), .A2(n16388), .ZN(n16385) );
  XNOR2_X1 U16431 ( .A(n16389), .B(n16390), .ZN(n16103) );
  NAND2_X1 U16432 ( .A1(n16391), .A2(n16392), .ZN(n16389) );
  XNOR2_X1 U16433 ( .A(n16393), .B(n16394), .ZN(n16111) );
  XNOR2_X1 U16434 ( .A(n16395), .B(n16396), .ZN(n16394) );
  XNOR2_X1 U16435 ( .A(n16397), .B(n16398), .ZN(n16119) );
  XNOR2_X1 U16436 ( .A(n16399), .B(n16400), .ZN(n16397) );
  XOR2_X1 U16437 ( .A(n16401), .B(n16402), .Z(n16127) );
  XOR2_X1 U16438 ( .A(n16403), .B(n16404), .Z(n16401) );
  XOR2_X1 U16439 ( .A(n16405), .B(n16406), .Z(n16135) );
  XOR2_X1 U16440 ( .A(n16407), .B(n16408), .Z(n16405) );
  XNOR2_X1 U16441 ( .A(n16409), .B(n16410), .ZN(n16143) );
  XNOR2_X1 U16442 ( .A(n16411), .B(n16412), .ZN(n16409) );
  XNOR2_X1 U16443 ( .A(n16413), .B(n16414), .ZN(n16151) );
  XNOR2_X1 U16444 ( .A(n16415), .B(n16416), .ZN(n16413) );
  XNOR2_X1 U16445 ( .A(n16417), .B(n16418), .ZN(n16159) );
  XNOR2_X1 U16446 ( .A(n16419), .B(n16420), .ZN(n16417) );
  XNOR2_X1 U16447 ( .A(n16421), .B(n16422), .ZN(n16167) );
  XNOR2_X1 U16448 ( .A(n16423), .B(n16424), .ZN(n16421) );
  XNOR2_X1 U16449 ( .A(n16425), .B(n16426), .ZN(n16175) );
  XNOR2_X1 U16450 ( .A(n16427), .B(n16428), .ZN(n16425) );
  XNOR2_X1 U16451 ( .A(n16429), .B(n16430), .ZN(n16179) );
  XNOR2_X1 U16452 ( .A(n16431), .B(n16432), .ZN(n16429) );
  XOR2_X1 U16453 ( .A(n16433), .B(n16434), .Z(n9015) );
  INV_X1 U16454 ( .A(n9071), .ZN(n9134) );
  NAND2_X1 U16455 ( .A1(n16435), .A2(n16436), .ZN(n9071) );
  NAND2_X1 U16456 ( .A1(n16434), .A2(n16433), .ZN(n16436) );
  XOR2_X1 U16457 ( .A(n8919), .B(n16437), .Z(n16435) );
  INV_X1 U16458 ( .A(n9072), .ZN(n9132) );
  NAND4_X1 U16459 ( .A1(n8919), .A2(n16437), .A3(n16434), .A4(n16433), .ZN(
        n9072) );
  NAND2_X1 U16460 ( .A1(n15949), .A2(n16438), .ZN(n16433) );
  NAND2_X1 U16461 ( .A1(n15948), .A2(n15950), .ZN(n16438) );
  NAND2_X1 U16462 ( .A1(n16439), .A2(n16440), .ZN(n15950) );
  NAND2_X1 U16463 ( .A1(a_0_), .A2(b_2_), .ZN(n16440) );
  XOR2_X1 U16464 ( .A(n16441), .B(n16442), .Z(n15948) );
  XOR2_X1 U16465 ( .A(n16443), .B(n8903), .Z(n16441) );
  NAND2_X1 U16466 ( .A1(a_0_), .A2(n16444), .ZN(n15949) );
  INV_X1 U16467 ( .A(n16439), .ZN(n16444) );
  NOR2_X1 U16468 ( .A1(n16445), .A2(n16446), .ZN(n16439) );
  NOR3_X1 U16469 ( .A1(n8997), .A2(n16447), .A3(n9731), .ZN(n16446) );
  INV_X1 U16470 ( .A(n16448), .ZN(n16447) );
  NAND2_X1 U16471 ( .A1(n16194), .A2(n16196), .ZN(n16448) );
  NOR2_X1 U16472 ( .A1(n16194), .A2(n16196), .ZN(n16445) );
  NAND2_X1 U16473 ( .A1(n16449), .A2(n16450), .ZN(n16196) );
  NAND2_X1 U16474 ( .A1(n16203), .A2(n16451), .ZN(n16450) );
  INV_X1 U16475 ( .A(n16452), .ZN(n16451) );
  NOR2_X1 U16476 ( .A1(n8889), .A2(n16204), .ZN(n16452) );
  XNOR2_X1 U16477 ( .A(n16453), .B(n16454), .ZN(n16203) );
  XOR2_X1 U16478 ( .A(n16455), .B(n16456), .Z(n16453) );
  NAND2_X1 U16479 ( .A1(n16204), .A2(n8889), .ZN(n16449) );
  NAND2_X1 U16480 ( .A1(a_2_), .A2(b_2_), .ZN(n8889) );
  NOR2_X1 U16481 ( .A1(n16457), .A2(n16458), .ZN(n16204) );
  INV_X1 U16482 ( .A(n16459), .ZN(n16458) );
  NAND2_X1 U16483 ( .A1(n16213), .A2(n16460), .ZN(n16459) );
  NAND2_X1 U16484 ( .A1(n16212), .A2(n16211), .ZN(n16460) );
  NOR2_X1 U16485 ( .A1(n8877), .A2(n8997), .ZN(n16213) );
  NOR2_X1 U16486 ( .A1(n16211), .A2(n16212), .ZN(n16457) );
  NOR2_X1 U16487 ( .A1(n16461), .A2(n16462), .ZN(n16212) );
  INV_X1 U16488 ( .A(n16463), .ZN(n16462) );
  NAND2_X1 U16489 ( .A1(n16221), .A2(n16464), .ZN(n16463) );
  NAND2_X1 U16490 ( .A1(n16220), .A2(n16219), .ZN(n16464) );
  NOR2_X1 U16491 ( .A1(n8996), .A2(n8997), .ZN(n16221) );
  NOR2_X1 U16492 ( .A1(n16219), .A2(n16220), .ZN(n16461) );
  NOR2_X1 U16493 ( .A1(n16465), .A2(n16466), .ZN(n16220) );
  INV_X1 U16494 ( .A(n16467), .ZN(n16466) );
  NAND2_X1 U16495 ( .A1(n16432), .A2(n16468), .ZN(n16467) );
  NAND2_X1 U16496 ( .A1(n16431), .A2(n16430), .ZN(n16468) );
  NOR2_X1 U16497 ( .A1(n8848), .A2(n8997), .ZN(n16432) );
  NOR2_X1 U16498 ( .A1(n16430), .A2(n16431), .ZN(n16465) );
  NOR2_X1 U16499 ( .A1(n16469), .A2(n16470), .ZN(n16431) );
  INV_X1 U16500 ( .A(n16471), .ZN(n16470) );
  NAND2_X1 U16501 ( .A1(n16232), .A2(n16472), .ZN(n16471) );
  NAND2_X1 U16502 ( .A1(n16231), .A2(n16230), .ZN(n16472) );
  NOR2_X1 U16503 ( .A1(n8994), .A2(n8997), .ZN(n16232) );
  NOR2_X1 U16504 ( .A1(n16230), .A2(n16231), .ZN(n16469) );
  NOR2_X1 U16505 ( .A1(n16473), .A2(n16474), .ZN(n16231) );
  INV_X1 U16506 ( .A(n16475), .ZN(n16474) );
  NAND2_X1 U16507 ( .A1(n16428), .A2(n16476), .ZN(n16475) );
  NAND2_X1 U16508 ( .A1(n16427), .A2(n16426), .ZN(n16476) );
  NOR2_X1 U16509 ( .A1(n8817), .A2(n8997), .ZN(n16428) );
  NOR2_X1 U16510 ( .A1(n16426), .A2(n16427), .ZN(n16473) );
  NOR2_X1 U16511 ( .A1(n16477), .A2(n16478), .ZN(n16427) );
  INV_X1 U16512 ( .A(n16479), .ZN(n16478) );
  NAND2_X1 U16513 ( .A1(n16244), .A2(n16480), .ZN(n16479) );
  NAND2_X1 U16514 ( .A1(n16243), .A2(n16242), .ZN(n16480) );
  NOR2_X1 U16515 ( .A1(n10513), .A2(n8997), .ZN(n16244) );
  NOR2_X1 U16516 ( .A1(n16242), .A2(n16243), .ZN(n16477) );
  NOR2_X1 U16517 ( .A1(n16481), .A2(n16482), .ZN(n16243) );
  INV_X1 U16518 ( .A(n16483), .ZN(n16482) );
  NAND2_X1 U16519 ( .A1(n16424), .A2(n16484), .ZN(n16483) );
  NAND2_X1 U16520 ( .A1(n16423), .A2(n16422), .ZN(n16484) );
  NOR2_X1 U16521 ( .A1(n8779), .A2(n8997), .ZN(n16424) );
  NOR2_X1 U16522 ( .A1(n16422), .A2(n16423), .ZN(n16481) );
  NOR2_X1 U16523 ( .A1(n16485), .A2(n16486), .ZN(n16423) );
  INV_X1 U16524 ( .A(n16487), .ZN(n16486) );
  NAND2_X1 U16525 ( .A1(n16257), .A2(n16488), .ZN(n16487) );
  NAND2_X1 U16526 ( .A1(n16256), .A2(n16255), .ZN(n16488) );
  NOR2_X1 U16527 ( .A1(n8769), .A2(n8997), .ZN(n16257) );
  NOR2_X1 U16528 ( .A1(n16255), .A2(n16256), .ZN(n16485) );
  NOR2_X1 U16529 ( .A1(n16489), .A2(n16490), .ZN(n16256) );
  INV_X1 U16530 ( .A(n16491), .ZN(n16490) );
  NAND2_X1 U16531 ( .A1(n16420), .A2(n16492), .ZN(n16491) );
  NAND2_X1 U16532 ( .A1(n16419), .A2(n16418), .ZN(n16492) );
  NOR2_X1 U16533 ( .A1(n8749), .A2(n8997), .ZN(n16420) );
  NOR2_X1 U16534 ( .A1(n16418), .A2(n16419), .ZN(n16489) );
  NOR2_X1 U16535 ( .A1(n16493), .A2(n16494), .ZN(n16419) );
  INV_X1 U16536 ( .A(n16495), .ZN(n16494) );
  NAND2_X1 U16537 ( .A1(n16269), .A2(n16496), .ZN(n16495) );
  NAND2_X1 U16538 ( .A1(n16268), .A2(n16267), .ZN(n16496) );
  NOR2_X1 U16539 ( .A1(n8739), .A2(n8997), .ZN(n16269) );
  NOR2_X1 U16540 ( .A1(n16267), .A2(n16268), .ZN(n16493) );
  NOR2_X1 U16541 ( .A1(n16497), .A2(n16498), .ZN(n16268) );
  INV_X1 U16542 ( .A(n16499), .ZN(n16498) );
  NAND2_X1 U16543 ( .A1(n16416), .A2(n16500), .ZN(n16499) );
  NAND2_X1 U16544 ( .A1(n16415), .A2(n16414), .ZN(n16500) );
  NOR2_X1 U16545 ( .A1(n8721), .A2(n8997), .ZN(n16416) );
  NOR2_X1 U16546 ( .A1(n16414), .A2(n16415), .ZN(n16497) );
  NOR2_X1 U16547 ( .A1(n16501), .A2(n16502), .ZN(n16415) );
  INV_X1 U16548 ( .A(n16503), .ZN(n16502) );
  NAND2_X1 U16549 ( .A1(n16281), .A2(n16504), .ZN(n16503) );
  NAND2_X1 U16550 ( .A1(n16280), .A2(n16279), .ZN(n16504) );
  NOR2_X1 U16551 ( .A1(n8991), .A2(n8997), .ZN(n16281) );
  NOR2_X1 U16552 ( .A1(n16279), .A2(n16280), .ZN(n16501) );
  NOR2_X1 U16553 ( .A1(n16505), .A2(n16506), .ZN(n16280) );
  INV_X1 U16554 ( .A(n16507), .ZN(n16506) );
  NAND2_X1 U16555 ( .A1(n16412), .A2(n16508), .ZN(n16507) );
  NAND2_X1 U16556 ( .A1(n16411), .A2(n16410), .ZN(n16508) );
  NOR2_X1 U16557 ( .A1(n8692), .A2(n8997), .ZN(n16412) );
  NOR2_X1 U16558 ( .A1(n16410), .A2(n16411), .ZN(n16505) );
  INV_X1 U16559 ( .A(n16509), .ZN(n16411) );
  NAND2_X1 U16560 ( .A1(n16510), .A2(n16511), .ZN(n16509) );
  NAND2_X1 U16561 ( .A1(n16293), .A2(n16512), .ZN(n16511) );
  INV_X1 U16562 ( .A(n16513), .ZN(n16512) );
  NOR2_X1 U16563 ( .A1(n16290), .A2(n16292), .ZN(n16513) );
  NOR2_X1 U16564 ( .A1(n8680), .A2(n8997), .ZN(n16293) );
  INV_X1 U16565 ( .A(a_16_), .ZN(n8680) );
  NAND2_X1 U16566 ( .A1(n16290), .A2(n16292), .ZN(n16510) );
  NAND2_X1 U16567 ( .A1(n16514), .A2(n16515), .ZN(n16292) );
  NAND2_X1 U16568 ( .A1(n16407), .A2(n16516), .ZN(n16515) );
  INV_X1 U16569 ( .A(n16517), .ZN(n16516) );
  NOR2_X1 U16570 ( .A1(n16408), .A2(n16406), .ZN(n16517) );
  NOR2_X1 U16571 ( .A1(n8662), .A2(n8997), .ZN(n16407) );
  NAND2_X1 U16572 ( .A1(n16406), .A2(n16408), .ZN(n16514) );
  NAND2_X1 U16573 ( .A1(n16518), .A2(n16519), .ZN(n16408) );
  NAND2_X1 U16574 ( .A1(n16305), .A2(n16520), .ZN(n16519) );
  INV_X1 U16575 ( .A(n16521), .ZN(n16520) );
  NOR2_X1 U16576 ( .A1(n16304), .A2(n16302), .ZN(n16521) );
  NOR2_X1 U16577 ( .A1(n8988), .A2(n8997), .ZN(n16305) );
  NAND2_X1 U16578 ( .A1(n16302), .A2(n16304), .ZN(n16518) );
  NAND2_X1 U16579 ( .A1(n16522), .A2(n16523), .ZN(n16304) );
  NAND2_X1 U16580 ( .A1(n16403), .A2(n16524), .ZN(n16523) );
  INV_X1 U16581 ( .A(n16525), .ZN(n16524) );
  NOR2_X1 U16582 ( .A1(n16404), .A2(n16402), .ZN(n16525) );
  NOR2_X1 U16583 ( .A1(n8997), .A2(n8630), .ZN(n16403) );
  NAND2_X1 U16584 ( .A1(n16402), .A2(n16404), .ZN(n16522) );
  NAND2_X1 U16585 ( .A1(n16526), .A2(n16527), .ZN(n16404) );
  NAND2_X1 U16586 ( .A1(n16317), .A2(n16528), .ZN(n16527) );
  INV_X1 U16587 ( .A(n16529), .ZN(n16528) );
  NOR2_X1 U16588 ( .A1(n16316), .A2(n16314), .ZN(n16529) );
  NOR2_X1 U16589 ( .A1(n8997), .A2(n8986), .ZN(n16317) );
  NAND2_X1 U16590 ( .A1(n16314), .A2(n16316), .ZN(n16526) );
  NAND2_X1 U16591 ( .A1(n16530), .A2(n16531), .ZN(n16316) );
  NAND2_X1 U16592 ( .A1(n16399), .A2(n16532), .ZN(n16531) );
  NAND2_X1 U16593 ( .A1(n16400), .A2(n16398), .ZN(n16532) );
  NOR2_X1 U16594 ( .A1(n8997), .A2(n8601), .ZN(n16399) );
  INV_X1 U16595 ( .A(n16533), .ZN(n16530) );
  NOR2_X1 U16596 ( .A1(n16398), .A2(n16400), .ZN(n16533) );
  NOR2_X1 U16597 ( .A1(n16534), .A2(n16535), .ZN(n16400) );
  NOR2_X1 U16598 ( .A1(n16329), .A2(n16536), .ZN(n16535) );
  NOR2_X1 U16599 ( .A1(n16328), .A2(n16326), .ZN(n16536) );
  NAND2_X1 U16600 ( .A1(b_2_), .A2(a_22_), .ZN(n16329) );
  INV_X1 U16601 ( .A(n16537), .ZN(n16534) );
  NAND2_X1 U16602 ( .A1(n16326), .A2(n16328), .ZN(n16537) );
  NAND2_X1 U16603 ( .A1(n16538), .A2(n16539), .ZN(n16328) );
  NAND2_X1 U16604 ( .A1(n16396), .A2(n16540), .ZN(n16539) );
  INV_X1 U16605 ( .A(n16541), .ZN(n16540) );
  NOR2_X1 U16606 ( .A1(n16395), .A2(n16393), .ZN(n16541) );
  NOR2_X1 U16607 ( .A1(n8997), .A2(n8572), .ZN(n16396) );
  NAND2_X1 U16608 ( .A1(n16393), .A2(n16395), .ZN(n16538) );
  NAND2_X1 U16609 ( .A1(n16339), .A2(n16542), .ZN(n16395) );
  NAND2_X1 U16610 ( .A1(n16338), .A2(n16340), .ZN(n16542) );
  NAND2_X1 U16611 ( .A1(n16543), .A2(n16544), .ZN(n16340) );
  NAND2_X1 U16612 ( .A1(b_2_), .A2(a_24_), .ZN(n16544) );
  INV_X1 U16613 ( .A(n16545), .ZN(n16543) );
  XOR2_X1 U16614 ( .A(n16546), .B(n16547), .Z(n16338) );
  XNOR2_X1 U16615 ( .A(n16548), .B(n16549), .ZN(n16547) );
  NAND2_X1 U16616 ( .A1(b_1_), .A2(a_25_), .ZN(n16546) );
  NAND2_X1 U16617 ( .A1(a_24_), .A2(n16545), .ZN(n16339) );
  NAND2_X1 U16618 ( .A1(n16391), .A2(n16550), .ZN(n16545) );
  NAND2_X1 U16619 ( .A1(n16390), .A2(n16392), .ZN(n16550) );
  NAND2_X1 U16620 ( .A1(n16551), .A2(n16552), .ZN(n16392) );
  NAND2_X1 U16621 ( .A1(b_2_), .A2(a_25_), .ZN(n16552) );
  XOR2_X1 U16622 ( .A(n16553), .B(n16554), .Z(n16390) );
  NOR2_X1 U16623 ( .A1(n9893), .A2(n8907), .ZN(n16554) );
  XOR2_X1 U16624 ( .A(n16555), .B(n16556), .Z(n16553) );
  NAND2_X1 U16625 ( .A1(a_25_), .A2(n16557), .ZN(n16391) );
  INV_X1 U16626 ( .A(n16551), .ZN(n16557) );
  NOR2_X1 U16627 ( .A1(n16558), .A2(n16559), .ZN(n16551) );
  NOR3_X1 U16628 ( .A1(n9893), .A2(n16560), .A3(n8997), .ZN(n16559) );
  NOR2_X1 U16629 ( .A1(n16352), .A2(n16350), .ZN(n16560) );
  INV_X1 U16630 ( .A(n16561), .ZN(n16558) );
  NAND2_X1 U16631 ( .A1(n16350), .A2(n16352), .ZN(n16561) );
  NAND2_X1 U16632 ( .A1(n16387), .A2(n16562), .ZN(n16352) );
  NAND2_X1 U16633 ( .A1(n16386), .A2(n16388), .ZN(n16562) );
  NAND2_X1 U16634 ( .A1(n16563), .A2(n16564), .ZN(n16388) );
  NAND2_X1 U16635 ( .A1(b_2_), .A2(a_27_), .ZN(n16564) );
  INV_X1 U16636 ( .A(n16565), .ZN(n16563) );
  XOR2_X1 U16637 ( .A(n16566), .B(n16567), .Z(n16386) );
  XNOR2_X1 U16638 ( .A(n16568), .B(n16569), .ZN(n16567) );
  NAND2_X1 U16639 ( .A1(b_1_), .A2(a_28_), .ZN(n16566) );
  NAND2_X1 U16640 ( .A1(a_27_), .A2(n16565), .ZN(n16387) );
  NAND2_X1 U16641 ( .A1(n16570), .A2(n16571), .ZN(n16565) );
  INV_X1 U16642 ( .A(n16572), .ZN(n16571) );
  NOR3_X1 U16643 ( .A1(n8493), .A2(n16573), .A3(n8997), .ZN(n16572) );
  NOR2_X1 U16644 ( .A1(n16382), .A2(n16384), .ZN(n16573) );
  NAND2_X1 U16645 ( .A1(n16382), .A2(n16384), .ZN(n16570) );
  NAND2_X1 U16646 ( .A1(n16574), .A2(n16575), .ZN(n16384) );
  NAND2_X1 U16647 ( .A1(n16378), .A2(n16576), .ZN(n16575) );
  INV_X1 U16648 ( .A(n16577), .ZN(n16576) );
  NOR2_X1 U16649 ( .A1(n16379), .A2(n16380), .ZN(n16577) );
  NOR2_X1 U16650 ( .A1(n8997), .A2(n8473), .ZN(n16378) );
  NAND2_X1 U16651 ( .A1(n16380), .A2(n16379), .ZN(n16574) );
  NAND2_X1 U16652 ( .A1(n16578), .A2(n16579), .ZN(n16379) );
  NAND2_X1 U16653 ( .A1(b_0_), .A2(n16580), .ZN(n16579) );
  NAND2_X1 U16654 ( .A1(n8456), .A2(n16581), .ZN(n16580) );
  NAND2_X1 U16655 ( .A1(a_31_), .A2(n8907), .ZN(n16581) );
  INV_X1 U16656 ( .A(a_30_), .ZN(n16582) );
  NAND2_X1 U16657 ( .A1(b_1_), .A2(n16583), .ZN(n16578) );
  NAND2_X1 U16658 ( .A1(n8459), .A2(n16584), .ZN(n16583) );
  NAND2_X1 U16659 ( .A1(a_30_), .A2(n16585), .ZN(n16584) );
  INV_X1 U16660 ( .A(a_31_), .ZN(n8978) );
  NOR3_X1 U16661 ( .A1(n8997), .A2(n8979), .A3(n8907), .ZN(n16380) );
  XNOR2_X1 U16662 ( .A(n16586), .B(n16587), .ZN(n16382) );
  XNOR2_X1 U16663 ( .A(n16588), .B(n16589), .ZN(n16587) );
  NAND2_X1 U16664 ( .A1(b_0_), .A2(a_30_), .ZN(n16586) );
  XOR2_X1 U16665 ( .A(n16590), .B(n16591), .Z(n16350) );
  XNOR2_X1 U16666 ( .A(n16592), .B(n16593), .ZN(n16591) );
  NAND2_X1 U16667 ( .A1(b_1_), .A2(a_27_), .ZN(n16590) );
  XOR2_X1 U16668 ( .A(n16594), .B(n16595), .Z(n16393) );
  NOR2_X1 U16669 ( .A1(n8982), .A2(n8907), .ZN(n16595) );
  XOR2_X1 U16670 ( .A(n16596), .B(n16597), .Z(n16594) );
  XOR2_X1 U16671 ( .A(n16598), .B(n16599), .Z(n16326) );
  XNOR2_X1 U16672 ( .A(n16600), .B(n16601), .ZN(n16599) );
  NAND2_X1 U16673 ( .A1(b_1_), .A2(a_23_), .ZN(n16598) );
  XNOR2_X1 U16674 ( .A(n16602), .B(n16603), .ZN(n16398) );
  NOR2_X1 U16675 ( .A1(n8984), .A2(n8907), .ZN(n16603) );
  XNOR2_X1 U16676 ( .A(n16604), .B(n16605), .ZN(n16602) );
  XOR2_X1 U16677 ( .A(n16606), .B(n16607), .Z(n16314) );
  XNOR2_X1 U16678 ( .A(n16608), .B(n16609), .ZN(n16607) );
  NAND2_X1 U16679 ( .A1(b_1_), .A2(a_21_), .ZN(n16606) );
  XOR2_X1 U16680 ( .A(n16610), .B(n16611), .Z(n16402) );
  NOR2_X1 U16681 ( .A1(n8986), .A2(n8907), .ZN(n16611) );
  XOR2_X1 U16682 ( .A(n16612), .B(n16613), .Z(n16610) );
  XOR2_X1 U16683 ( .A(n16614), .B(n16615), .Z(n16302) );
  XNOR2_X1 U16684 ( .A(n16616), .B(n16617), .ZN(n16615) );
  NAND2_X1 U16685 ( .A1(b_1_), .A2(a_19_), .ZN(n16614) );
  XOR2_X1 U16686 ( .A(n16618), .B(n16619), .Z(n16406) );
  XNOR2_X1 U16687 ( .A(n16620), .B(n16621), .ZN(n16618) );
  XNOR2_X1 U16688 ( .A(n16622), .B(n16623), .ZN(n16290) );
  XNOR2_X1 U16689 ( .A(n16624), .B(n16625), .ZN(n16622) );
  XNOR2_X1 U16690 ( .A(n16626), .B(n16627), .ZN(n16410) );
  XNOR2_X1 U16691 ( .A(n16628), .B(n16629), .ZN(n16627) );
  XNOR2_X1 U16692 ( .A(n16630), .B(n16631), .ZN(n16279) );
  XOR2_X1 U16693 ( .A(n16632), .B(n16633), .Z(n16630) );
  XOR2_X1 U16694 ( .A(n16634), .B(n16635), .Z(n16414) );
  XNOR2_X1 U16695 ( .A(n16636), .B(n16637), .ZN(n16635) );
  XNOR2_X1 U16696 ( .A(n16638), .B(n16639), .ZN(n16267) );
  XOR2_X1 U16697 ( .A(n16640), .B(n16641), .Z(n16638) );
  XOR2_X1 U16698 ( .A(n16642), .B(n16643), .Z(n16418) );
  XNOR2_X1 U16699 ( .A(n16644), .B(n16645), .ZN(n16643) );
  XOR2_X1 U16700 ( .A(n16646), .B(n16647), .Z(n16255) );
  XNOR2_X1 U16701 ( .A(n16648), .B(n16649), .ZN(n16647) );
  XNOR2_X1 U16702 ( .A(n16650), .B(n16651), .ZN(n16422) );
  XOR2_X1 U16703 ( .A(n16652), .B(n16653), .Z(n16650) );
  XNOR2_X1 U16704 ( .A(n16654), .B(n16655), .ZN(n16242) );
  XOR2_X1 U16705 ( .A(n16656), .B(n16657), .Z(n16654) );
  XNOR2_X1 U16706 ( .A(n16658), .B(n16659), .ZN(n16426) );
  XOR2_X1 U16707 ( .A(n16660), .B(n16661), .Z(n16658) );
  XNOR2_X1 U16708 ( .A(n16662), .B(n16663), .ZN(n16230) );
  XOR2_X1 U16709 ( .A(n16664), .B(n16665), .Z(n16662) );
  XNOR2_X1 U16710 ( .A(n16666), .B(n16667), .ZN(n16430) );
  XOR2_X1 U16711 ( .A(n16668), .B(n16669), .Z(n16666) );
  XNOR2_X1 U16712 ( .A(n16670), .B(n16671), .ZN(n16219) );
  XOR2_X1 U16713 ( .A(n16672), .B(n16673), .Z(n16670) );
  XNOR2_X1 U16714 ( .A(n16674), .B(n16675), .ZN(n16211) );
  XOR2_X1 U16715 ( .A(n16676), .B(n16677), .Z(n16674) );
  XNOR2_X1 U16716 ( .A(n16678), .B(n16679), .ZN(n16194) );
  XOR2_X1 U16717 ( .A(n16680), .B(n16681), .Z(n16678) );
  XOR2_X1 U16718 ( .A(n16682), .B(n16683), .Z(n16434) );
  NOR2_X1 U16719 ( .A1(n16585), .A2(n9731), .ZN(n16683) );
  XOR2_X1 U16720 ( .A(n16684), .B(n16685), .Z(n16682) );
  NOR2_X1 U16721 ( .A1(n9471), .A2(n16585), .ZN(n8919) );
  NOR2_X1 U16722 ( .A1(n16437), .A2(n9471), .ZN(n9131) );
  NOR2_X1 U16723 ( .A1(n16686), .A2(n16687), .ZN(n16437) );
  NOR3_X1 U16724 ( .A1(n16585), .A2(n16688), .A3(n9731), .ZN(n16687) );
  NOR2_X1 U16725 ( .A1(n16684), .A2(n16685), .ZN(n16688) );
  INV_X1 U16726 ( .A(n16689), .ZN(n16686) );
  NAND2_X1 U16727 ( .A1(n16685), .A2(n16684), .ZN(n16689) );
  NAND2_X1 U16728 ( .A1(n16690), .A2(n16691), .ZN(n16684) );
  NAND2_X1 U16729 ( .A1(n16442), .A2(n16692), .ZN(n16691) );
  INV_X1 U16730 ( .A(n16693), .ZN(n16692) );
  NOR2_X1 U16731 ( .A1(n16443), .A2(n8903), .ZN(n16693) );
  NOR2_X1 U16732 ( .A1(n8998), .A2(n16585), .ZN(n16442) );
  NAND2_X1 U16733 ( .A1(n8903), .A2(n16443), .ZN(n16690) );
  NAND2_X1 U16734 ( .A1(n16694), .A2(n16695), .ZN(n16443) );
  NAND2_X1 U16735 ( .A1(n16679), .A2(n16696), .ZN(n16695) );
  INV_X1 U16736 ( .A(n16697), .ZN(n16696) );
  NOR2_X1 U16737 ( .A1(n16680), .A2(n16681), .ZN(n16697) );
  NOR2_X1 U16738 ( .A1(n8998), .A2(n8907), .ZN(n16679) );
  NAND2_X1 U16739 ( .A1(n16681), .A2(n16680), .ZN(n16694) );
  NAND2_X1 U16740 ( .A1(n16698), .A2(n16699), .ZN(n16680) );
  NAND2_X1 U16741 ( .A1(n16454), .A2(n16700), .ZN(n16699) );
  INV_X1 U16742 ( .A(n16701), .ZN(n16700) );
  NOR2_X1 U16743 ( .A1(n16455), .A2(n16456), .ZN(n16701) );
  NOR2_X1 U16744 ( .A1(n8877), .A2(n8907), .ZN(n16454) );
  NAND2_X1 U16745 ( .A1(n16456), .A2(n16455), .ZN(n16698) );
  NAND2_X1 U16746 ( .A1(n16702), .A2(n16703), .ZN(n16455) );
  NAND2_X1 U16747 ( .A1(n16675), .A2(n16704), .ZN(n16703) );
  INV_X1 U16748 ( .A(n16705), .ZN(n16704) );
  NOR2_X1 U16749 ( .A1(n16676), .A2(n16677), .ZN(n16705) );
  NOR2_X1 U16750 ( .A1(n8996), .A2(n8907), .ZN(n16675) );
  NAND2_X1 U16751 ( .A1(n16677), .A2(n16676), .ZN(n16702) );
  NAND2_X1 U16752 ( .A1(n16706), .A2(n16707), .ZN(n16676) );
  NAND2_X1 U16753 ( .A1(n16671), .A2(n16708), .ZN(n16707) );
  INV_X1 U16754 ( .A(n16709), .ZN(n16708) );
  NOR2_X1 U16755 ( .A1(n16672), .A2(n16673), .ZN(n16709) );
  NOR2_X1 U16756 ( .A1(n8848), .A2(n8907), .ZN(n16671) );
  NAND2_X1 U16757 ( .A1(n16673), .A2(n16672), .ZN(n16706) );
  NAND2_X1 U16758 ( .A1(n16710), .A2(n16711), .ZN(n16672) );
  NAND2_X1 U16759 ( .A1(n16667), .A2(n16712), .ZN(n16711) );
  INV_X1 U16760 ( .A(n16713), .ZN(n16712) );
  NOR2_X1 U16761 ( .A1(n16668), .A2(n16669), .ZN(n16713) );
  NOR2_X1 U16762 ( .A1(n8994), .A2(n8907), .ZN(n16667) );
  NAND2_X1 U16763 ( .A1(n16669), .A2(n16668), .ZN(n16710) );
  NAND2_X1 U16764 ( .A1(n16714), .A2(n16715), .ZN(n16668) );
  NAND2_X1 U16765 ( .A1(n16663), .A2(n16716), .ZN(n16715) );
  INV_X1 U16766 ( .A(n16717), .ZN(n16716) );
  NOR2_X1 U16767 ( .A1(n16664), .A2(n16665), .ZN(n16717) );
  NOR2_X1 U16768 ( .A1(n8817), .A2(n8907), .ZN(n16663) );
  NAND2_X1 U16769 ( .A1(n16665), .A2(n16664), .ZN(n16714) );
  NAND2_X1 U16770 ( .A1(n16718), .A2(n16719), .ZN(n16664) );
  NAND2_X1 U16771 ( .A1(n16659), .A2(n16720), .ZN(n16719) );
  INV_X1 U16772 ( .A(n16721), .ZN(n16720) );
  NOR2_X1 U16773 ( .A1(n16660), .A2(n16661), .ZN(n16721) );
  NOR2_X1 U16774 ( .A1(n10513), .A2(n8907), .ZN(n16659) );
  NAND2_X1 U16775 ( .A1(n16661), .A2(n16660), .ZN(n16718) );
  NAND2_X1 U16776 ( .A1(n16722), .A2(n16723), .ZN(n16660) );
  NAND2_X1 U16777 ( .A1(n16655), .A2(n16724), .ZN(n16723) );
  INV_X1 U16778 ( .A(n16725), .ZN(n16724) );
  NOR2_X1 U16779 ( .A1(n16656), .A2(n16657), .ZN(n16725) );
  NOR2_X1 U16780 ( .A1(n8779), .A2(n8907), .ZN(n16655) );
  NAND2_X1 U16781 ( .A1(n16657), .A2(n16656), .ZN(n16722) );
  NAND2_X1 U16782 ( .A1(n16726), .A2(n16727), .ZN(n16656) );
  NAND2_X1 U16783 ( .A1(n16651), .A2(n16728), .ZN(n16727) );
  INV_X1 U16784 ( .A(n16729), .ZN(n16728) );
  NOR2_X1 U16785 ( .A1(n16652), .A2(n16653), .ZN(n16729) );
  NOR2_X1 U16786 ( .A1(n8769), .A2(n8907), .ZN(n16651) );
  NAND2_X1 U16787 ( .A1(n16653), .A2(n16652), .ZN(n16726) );
  NAND2_X1 U16788 ( .A1(n16730), .A2(n16731), .ZN(n16652) );
  NAND2_X1 U16789 ( .A1(n16646), .A2(n16732), .ZN(n16731) );
  NAND2_X1 U16790 ( .A1(n16648), .A2(n16649), .ZN(n16732) );
  NOR2_X1 U16791 ( .A1(n8749), .A2(n8907), .ZN(n16646) );
  INV_X1 U16792 ( .A(n16733), .ZN(n16730) );
  NOR2_X1 U16793 ( .A1(n16649), .A2(n16648), .ZN(n16733) );
  NOR2_X1 U16794 ( .A1(n16734), .A2(n16735), .ZN(n16648) );
  INV_X1 U16795 ( .A(n16736), .ZN(n16735) );
  NAND2_X1 U16796 ( .A1(n16642), .A2(n16737), .ZN(n16736) );
  NAND2_X1 U16797 ( .A1(n16644), .A2(n16645), .ZN(n16737) );
  NOR2_X1 U16798 ( .A1(n8739), .A2(n8907), .ZN(n16642) );
  NOR2_X1 U16799 ( .A1(n16645), .A2(n16644), .ZN(n16734) );
  NOR2_X1 U16800 ( .A1(n16738), .A2(n16739), .ZN(n16644) );
  INV_X1 U16801 ( .A(n16740), .ZN(n16739) );
  NAND2_X1 U16802 ( .A1(n16639), .A2(n16741), .ZN(n16740) );
  NAND2_X1 U16803 ( .A1(n16641), .A2(n16640), .ZN(n16741) );
  NOR2_X1 U16804 ( .A1(n8721), .A2(n8907), .ZN(n16639) );
  NOR2_X1 U16805 ( .A1(n16640), .A2(n16641), .ZN(n16738) );
  NOR2_X1 U16806 ( .A1(n16742), .A2(n16743), .ZN(n16641) );
  INV_X1 U16807 ( .A(n16744), .ZN(n16743) );
  NAND2_X1 U16808 ( .A1(n16634), .A2(n16745), .ZN(n16744) );
  NAND2_X1 U16809 ( .A1(n16636), .A2(n16637), .ZN(n16745) );
  NOR2_X1 U16810 ( .A1(n8991), .A2(n8907), .ZN(n16634) );
  INV_X1 U16811 ( .A(a_14_), .ZN(n8991) );
  NOR2_X1 U16812 ( .A1(n16637), .A2(n16636), .ZN(n16742) );
  NOR2_X1 U16813 ( .A1(n16746), .A2(n16747), .ZN(n16636) );
  INV_X1 U16814 ( .A(n16748), .ZN(n16747) );
  NAND2_X1 U16815 ( .A1(n16631), .A2(n16749), .ZN(n16748) );
  NAND2_X1 U16816 ( .A1(n16633), .A2(n16632), .ZN(n16749) );
  NOR2_X1 U16817 ( .A1(n8692), .A2(n8907), .ZN(n16631) );
  NOR2_X1 U16818 ( .A1(n16632), .A2(n16633), .ZN(n16746) );
  NOR2_X1 U16819 ( .A1(n16750), .A2(n16751), .ZN(n16633) );
  NOR2_X1 U16820 ( .A1(n16626), .A2(n16752), .ZN(n16751) );
  NOR2_X1 U16821 ( .A1(n16628), .A2(n16629), .ZN(n16752) );
  NAND2_X1 U16822 ( .A1(a_16_), .A2(b_1_), .ZN(n16626) );
  INV_X1 U16823 ( .A(n16753), .ZN(n16750) );
  NAND2_X1 U16824 ( .A1(n16629), .A2(n16628), .ZN(n16753) );
  NAND2_X1 U16825 ( .A1(n16754), .A2(n16755), .ZN(n16628) );
  NAND2_X1 U16826 ( .A1(n16623), .A2(n16756), .ZN(n16755) );
  INV_X1 U16827 ( .A(n16757), .ZN(n16756) );
  NOR2_X1 U16828 ( .A1(n16624), .A2(n16625), .ZN(n16757) );
  NOR2_X1 U16829 ( .A1(n8662), .A2(n8907), .ZN(n16623) );
  NAND2_X1 U16830 ( .A1(n16624), .A2(n16625), .ZN(n16754) );
  NOR2_X1 U16831 ( .A1(n8988), .A2(n16585), .ZN(n16625) );
  NOR2_X1 U16832 ( .A1(n16758), .A2(n16759), .ZN(n16624) );
  INV_X1 U16833 ( .A(n16760), .ZN(n16759) );
  NAND2_X1 U16834 ( .A1(n16761), .A2(n16620), .ZN(n16760) );
  NAND2_X1 U16835 ( .A1(b_0_), .A2(a_19_), .ZN(n16620) );
  NAND2_X1 U16836 ( .A1(n16619), .A2(n16621), .ZN(n16761) );
  NOR2_X1 U16837 ( .A1(n16621), .A2(n16619), .ZN(n16758) );
  NOR2_X1 U16838 ( .A1(n8988), .A2(n8907), .ZN(n16619) );
  NAND2_X1 U16839 ( .A1(n16762), .A2(n16763), .ZN(n16621) );
  INV_X1 U16840 ( .A(n16764), .ZN(n16763) );
  NOR3_X1 U16841 ( .A1(n8630), .A2(n16765), .A3(n8907), .ZN(n16764) );
  NOR2_X1 U16842 ( .A1(n16617), .A2(n16616), .ZN(n16765) );
  INV_X1 U16843 ( .A(a_19_), .ZN(n8630) );
  NAND2_X1 U16844 ( .A1(n16616), .A2(n16617), .ZN(n16762) );
  NAND2_X1 U16845 ( .A1(n16766), .A2(n16767), .ZN(n16617) );
  NAND3_X1 U16846 ( .A1(a_20_), .A2(n16768), .A3(b_1_), .ZN(n16767) );
  NAND2_X1 U16847 ( .A1(n16613), .A2(n16612), .ZN(n16768) );
  INV_X1 U16848 ( .A(n16769), .ZN(n16766) );
  NOR2_X1 U16849 ( .A1(n16612), .A2(n16613), .ZN(n16769) );
  NOR2_X1 U16850 ( .A1(n16770), .A2(n16771), .ZN(n16613) );
  NOR3_X1 U16851 ( .A1(n8601), .A2(n16772), .A3(n8907), .ZN(n16771) );
  NOR2_X1 U16852 ( .A1(n16609), .A2(n16608), .ZN(n16772) );
  INV_X1 U16853 ( .A(n16773), .ZN(n16770) );
  NAND2_X1 U16854 ( .A1(n16608), .A2(n16609), .ZN(n16773) );
  NAND2_X1 U16855 ( .A1(n16774), .A2(n16775), .ZN(n16609) );
  NAND3_X1 U16856 ( .A1(a_22_), .A2(n16776), .A3(b_1_), .ZN(n16775) );
  NAND2_X1 U16857 ( .A1(n16605), .A2(n16777), .ZN(n16776) );
  INV_X1 U16858 ( .A(n16778), .ZN(n16774) );
  NOR2_X1 U16859 ( .A1(n16777), .A2(n16605), .ZN(n16778) );
  NOR2_X1 U16860 ( .A1(n16779), .A2(n16780), .ZN(n16605) );
  NOR3_X1 U16861 ( .A1(n8572), .A2(n16781), .A3(n8907), .ZN(n16780) );
  NOR2_X1 U16862 ( .A1(n16601), .A2(n16600), .ZN(n16781) );
  INV_X1 U16863 ( .A(n16782), .ZN(n16779) );
  NAND2_X1 U16864 ( .A1(n16600), .A2(n16601), .ZN(n16782) );
  NAND2_X1 U16865 ( .A1(n16783), .A2(n16784), .ZN(n16601) );
  NAND3_X1 U16866 ( .A1(a_24_), .A2(n16785), .A3(b_1_), .ZN(n16784) );
  NAND2_X1 U16867 ( .A1(n16597), .A2(n16596), .ZN(n16785) );
  INV_X1 U16868 ( .A(n16786), .ZN(n16783) );
  NOR2_X1 U16869 ( .A1(n16596), .A2(n16597), .ZN(n16786) );
  NOR2_X1 U16870 ( .A1(n16787), .A2(n16788), .ZN(n16597) );
  NOR3_X1 U16871 ( .A1(n8541), .A2(n16789), .A3(n8907), .ZN(n16788) );
  NOR2_X1 U16872 ( .A1(n16549), .A2(n16548), .ZN(n16789) );
  INV_X1 U16873 ( .A(n16790), .ZN(n16787) );
  NAND2_X1 U16874 ( .A1(n16548), .A2(n16549), .ZN(n16790) );
  NAND2_X1 U16875 ( .A1(n16791), .A2(n16792), .ZN(n16549) );
  NAND3_X1 U16876 ( .A1(a_26_), .A2(n16793), .A3(b_1_), .ZN(n16792) );
  NAND2_X1 U16877 ( .A1(n16556), .A2(n16555), .ZN(n16793) );
  INV_X1 U16878 ( .A(n16794), .ZN(n16791) );
  NOR2_X1 U16879 ( .A1(n16555), .A2(n16556), .ZN(n16794) );
  NOR2_X1 U16880 ( .A1(n16795), .A2(n16796), .ZN(n16556) );
  NOR3_X1 U16881 ( .A1(n8512), .A2(n16797), .A3(n8907), .ZN(n16796) );
  NOR2_X1 U16882 ( .A1(n16593), .A2(n16592), .ZN(n16797) );
  INV_X1 U16883 ( .A(n16798), .ZN(n16795) );
  NAND2_X1 U16884 ( .A1(n16592), .A2(n16593), .ZN(n16798) );
  NAND2_X1 U16885 ( .A1(n16799), .A2(n16800), .ZN(n16593) );
  INV_X1 U16886 ( .A(n16801), .ZN(n16800) );
  NOR3_X1 U16887 ( .A1(n8493), .A2(n16802), .A3(n8907), .ZN(n16801) );
  NOR2_X1 U16888 ( .A1(n16569), .A2(n16568), .ZN(n16802) );
  NAND2_X1 U16889 ( .A1(n16568), .A2(n16569), .ZN(n16799) );
  NAND2_X1 U16890 ( .A1(n16589), .A2(n16803), .ZN(n16569) );
  NAND3_X1 U16891 ( .A1(b_0_), .A2(a_30_), .A3(n16588), .ZN(n16803) );
  NOR2_X1 U16892 ( .A1(n8907), .A2(n8473), .ZN(n16588) );
  NAND3_X1 U16893 ( .A1(b_1_), .A2(n9666), .A3(b_0_), .ZN(n16589) );
  INV_X1 U16894 ( .A(n8979), .ZN(n9666) );
  NOR2_X1 U16895 ( .A1(n16585), .A2(n8473), .ZN(n16568) );
  NOR2_X1 U16896 ( .A1(n16585), .A2(n8493), .ZN(n16592) );
  NAND2_X1 U16897 ( .A1(b_0_), .A2(a_27_), .ZN(n16555) );
  NOR2_X1 U16898 ( .A1(n16585), .A2(n9893), .ZN(n16548) );
  NAND2_X1 U16899 ( .A1(b_0_), .A2(a_25_), .ZN(n16596) );
  NOR2_X1 U16900 ( .A1(n16585), .A2(n8982), .ZN(n16600) );
  INV_X1 U16901 ( .A(n16604), .ZN(n16777) );
  NOR2_X1 U16902 ( .A1(n16585), .A2(n8572), .ZN(n16604) );
  INV_X1 U16903 ( .A(a_23_), .ZN(n8572) );
  NOR2_X1 U16904 ( .A1(n16585), .A2(n8984), .ZN(n16608) );
  INV_X1 U16905 ( .A(a_22_), .ZN(n8984) );
  NAND2_X1 U16906 ( .A1(b_0_), .A2(a_21_), .ZN(n16612) );
  NOR2_X1 U16907 ( .A1(n16585), .A2(n8986), .ZN(n16616) );
  NOR2_X1 U16908 ( .A1(n8662), .A2(n16585), .ZN(n16629) );
  NAND2_X1 U16909 ( .A1(a_16_), .A2(b_0_), .ZN(n16632) );
  NAND2_X1 U16910 ( .A1(a_15_), .A2(b_0_), .ZN(n16637) );
  NAND2_X1 U16911 ( .A1(a_14_), .A2(b_0_), .ZN(n16640) );
  NAND2_X1 U16912 ( .A1(a_13_), .A2(b_0_), .ZN(n16645) );
  NAND2_X1 U16913 ( .A1(a_12_), .A2(b_0_), .ZN(n16649) );
  NOR2_X1 U16914 ( .A1(n8749), .A2(n16585), .ZN(n16653) );
  NOR2_X1 U16915 ( .A1(n8769), .A2(n16585), .ZN(n16657) );
  NOR2_X1 U16916 ( .A1(n8779), .A2(n16585), .ZN(n16661) );
  NOR2_X1 U16917 ( .A1(n10513), .A2(n16585), .ZN(n16665) );
  INV_X1 U16918 ( .A(a_8_), .ZN(n10513) );
  NOR2_X1 U16919 ( .A1(n8817), .A2(n16585), .ZN(n16669) );
  NOR2_X1 U16920 ( .A1(n8994), .A2(n16585), .ZN(n16673) );
  INV_X1 U16921 ( .A(a_6_), .ZN(n8994) );
  NOR2_X1 U16922 ( .A1(n8848), .A2(n16585), .ZN(n16677) );
  NOR2_X1 U16923 ( .A1(n8996), .A2(n16585), .ZN(n16456) );
  INV_X1 U16924 ( .A(a_4_), .ZN(n8996) );
  NOR2_X1 U16925 ( .A1(n8877), .A2(n16585), .ZN(n16681) );
  INV_X1 U16926 ( .A(b_0_), .ZN(n16585) );
  NOR2_X1 U16927 ( .A1(n9731), .A2(n8907), .ZN(n8903) );
  INV_X1 U16928 ( .A(a_1_), .ZN(n9731) );
  NOR2_X1 U16929 ( .A1(n9471), .A2(n8907), .ZN(n16685) );
  INV_X1 U16930 ( .A(a_0_), .ZN(n9471) );
endmodule

