module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n155_, new_n384_, new_n410_, new_n445_, new_n236_, new_n238_, new_n479_, new_n92_, new_n79_, new_n543_, new_n250_, new_n113_, new_n501_, new_n288_, new_n371_, new_n509_, new_n97_, new_n454_, new_n421_, new_n202_, new_n296_, new_n308_, new_n368_, new_n232_, new_n258_, new_n76_, new_n439_, new_n176_, new_n283_, new_n223_, new_n390_, new_n156_, new_n306_, new_n366_, new_n494_, new_n291_, new_n241_, new_n261_, new_n309_, new_n566_, new_n186_, new_n365_, new_n339_, new_n197_, new_n529_, new_n386_, new_n82_, new_n401_, new_n389_, new_n323_, new_n259_, new_n362_, new_n514_, new_n227_, new_n416_, new_n222_, new_n456_, new_n170_, new_n246_, new_n571_, new_n400_, new_n328_, new_n460_, new_n367_, new_n548_, new_n173_, new_n220_, new_n130_, new_n505_, new_n419_, new_n471_, new_n268_, new_n374_, new_n534_, new_n376_, new_n380_, new_n214_, new_n451_, new_n489_, new_n424_, new_n138_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n240_, new_n413_, new_n526_, new_n352_, new_n442_, new_n485_, new_n525_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n562_, new_n126_, new_n462_, new_n564_, new_n177_, new_n493_, new_n264_, new_n379_, new_n500_, new_n273_, new_n224_, new_n270_, new_n570_, new_n317_, new_n102_, new_n344_, new_n143_, new_n520_, new_n287_, new_n125_, new_n145_, new_n253_, new_n504_, new_n475_, new_n90_, new_n237_, new_n427_, new_n234_, new_n532_, new_n149_, new_n472_, new_n557_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n106_, new_n411_, new_n215_, new_n507_, new_n152_, new_n157_, new_n107_, new_n93_, new_n182_, new_n153_, new_n407_, new_n81_, new_n480_, new_n133_, new_n257_, new_n481_, new_n212_, new_n151_, new_n513_, new_n364_, new_n449_, new_n558_, new_n484_, new_n219_, new_n231_, new_n313_, new_n78_, new_n239_, new_n272_, new_n282_, new_n382_, new_n522_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n146_, new_n88_, new_n487_, new_n360_, new_n98_, new_n546_, new_n110_, new_n315_, new_n302_, new_n191_, new_n124_, new_n326_, new_n554_, new_n95_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n87_, new_n387_, new_n544_, new_n103_, new_n476_, new_n112_, new_n248_, new_n350_, new_n117_, new_n121_, new_n415_, new_n167_, new_n537_, new_n221_, new_n385_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n478_, new_n461_, new_n459_, new_n569_, new_n555_, new_n174_, new_n297_, new_n361_, new_n565_, new_n468_, new_n150_, new_n354_, new_n392_, new_n444_, new_n518_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n105_, new_n340_, new_n147_, new_n510_, new_n285_, new_n502_, new_n80_, new_n351_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n517_, new_n325_, new_n417_, new_n180_, new_n515_, new_n530_, new_n332_, new_n318_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n531_, new_n111_, new_n158_, new_n252_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n160_, new_n312_, new_n271_, new_n535_, new_n274_, new_n372_, new_n100_, new_n242_, new_n503_, new_n527_, new_n218_, new_n497_, new_n115_, new_n307_, new_n190_, new_n305_, new_n420_, new_n568_, new_n408_, new_n470_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n213_, new_n134_, new_n433_, new_n435_, new_n206_, new_n109_, new_n254_, new_n429_, new_n355_, new_n353_, new_n85_, new_n432_, new_n265_, new_n506_, new_n370_, new_n256_, new_n452_, new_n278_, new_n304_, new_n381_, new_n523_, new_n388_, new_n550_, new_n217_, new_n101_, new_n269_, new_n508_, new_n512_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n129_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n412_, new_n165_, new_n441_, new_n477_, new_n327_, new_n216_, new_n561_, new_n495_, new_n431_, new_n77_, new_n196_, new_n280_, new_n426_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n338_, new_n207_, new_n267_, new_n473_, new_n140_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n86_, new_n465_, new_n84_, new_n195_, new_n567_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n245_, new_n402_, new_n474_, new_n89_, new_n467_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n490_, new_n560_, new_n91_, new_n346_, new_n396_, new_n198_, new_n438_, new_n128_, new_n358_, new_n208_, new_n348_, new_n159_, new_n83_, new_n322_, new_n228_, new_n545_, new_n289_, new_n528_, new_n179_, new_n572_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n104_, new_n185_, new_n399_, new_n373_, new_n171_, new_n559_, new_n540_, new_n434_, new_n200_, new_n422_, new_n99_, new_n329_, new_n249_, new_n233_, new_n136_, new_n469_, new_n284_, new_n119_, new_n391_, new_n293_, new_n96_, new_n178_, new_n437_, new_n551_, new_n168_, new_n279_, new_n455_, new_n295_, new_n359_, new_n132_, new_n120_, new_n521_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n406_, new_n356_, new_n333_, new_n229_, new_n536_, new_n290_, new_n464_, new_n94_, new_n204_, new_n369_, new_n181_, new_n135_, new_n448_, new_n573_, new_n276_, new_n405_;

not g000 ( new_n76_, N56 );
or g001 ( new_n77_, new_n76_, N50 );
not g002 ( new_n78_, N69 );
or g003 ( new_n79_, new_n78_, N63 );
and g004 ( new_n80_, new_n77_, new_n79_ );
not g005 ( new_n81_, N82 );
or g006 ( new_n82_, new_n81_, N76 );
not g007 ( new_n83_, N95 );
or g008 ( new_n84_, new_n83_, N89 );
and g009 ( new_n85_, new_n82_, new_n84_ );
and g010 ( new_n86_, new_n80_, new_n85_ );
not g011 ( new_n87_, N4 );
or g012 ( new_n88_, new_n87_, N1 );
not g013 ( new_n89_, N17 );
or g014 ( new_n90_, new_n89_, N11 );
and g015 ( new_n91_, new_n88_, new_n90_ );
not g016 ( new_n92_, N30 );
or g017 ( new_n93_, new_n92_, N24 );
not g018 ( new_n94_, N43 );
or g019 ( new_n95_, new_n94_, N37 );
and g020 ( new_n96_, new_n93_, new_n95_ );
and g021 ( new_n97_, new_n91_, new_n96_ );
and g022 ( new_n98_, new_n86_, new_n97_ );
not g023 ( new_n99_, keyIn_0_4 );
not g024 ( new_n100_, N102 );
and g025 ( new_n101_, new_n100_, N108 );
and g026 ( new_n102_, new_n101_, new_n99_ );
not g027 ( new_n103_, new_n102_ );
or g028 ( new_n104_, new_n101_, new_n99_ );
and g029 ( new_n105_, new_n103_, new_n104_ );
not g030 ( new_n106_, new_n105_ );
and g031 ( new_n107_, new_n98_, new_n106_ );
not g032 ( N223, new_n107_ );
not g033 ( new_n109_, N89 );
and g034 ( new_n110_, new_n109_, N95 );
or g035 ( new_n111_, new_n107_, new_n110_ );
not g036 ( new_n112_, N99 );
and g037 ( new_n113_, new_n83_, keyIn_0_2 );
not g038 ( new_n114_, new_n113_ );
or g039 ( new_n115_, new_n83_, keyIn_0_2 );
and g040 ( new_n116_, new_n114_, new_n115_ );
not g041 ( new_n117_, new_n116_ );
and g042 ( new_n118_, new_n117_, new_n112_ );
and g043 ( new_n119_, new_n111_, new_n118_ );
and g044 ( new_n120_, new_n119_, keyIn_0_17 );
not g045 ( new_n121_, new_n120_ );
or g046 ( new_n122_, new_n119_, keyIn_0_17 );
and g047 ( new_n123_, new_n121_, new_n122_ );
not g048 ( new_n124_, new_n123_ );
and g049 ( new_n125_, N223, new_n77_ );
not g050 ( new_n126_, N50 );
and g051 ( new_n127_, new_n126_, N56 );
and g052 ( new_n128_, new_n107_, new_n127_ );
or g053 ( new_n129_, new_n125_, new_n128_ );
not g054 ( new_n130_, N60 );
and g055 ( new_n131_, new_n130_, N56 );
not g056 ( new_n132_, new_n131_ );
or g057 ( new_n133_, new_n129_, new_n132_ );
not g058 ( new_n134_, N1 );
and g059 ( new_n135_, new_n134_, N4 );
and g060 ( new_n136_, N223, new_n135_ );
and g061 ( new_n137_, new_n107_, new_n88_ );
or g062 ( new_n138_, new_n136_, new_n137_ );
not g063 ( new_n139_, new_n138_ );
and g064 ( new_n140_, new_n87_, keyIn_0_0 );
not g065 ( new_n141_, new_n140_ );
or g066 ( new_n142_, new_n87_, keyIn_0_0 );
and g067 ( new_n143_, new_n141_, new_n142_ );
or g068 ( new_n144_, new_n143_, N8 );
or g069 ( new_n145_, new_n139_, new_n144_ );
and g070 ( new_n146_, N223, new_n82_ );
not g071 ( new_n147_, N86 );
and g072 ( new_n148_, new_n147_, N82 );
not g073 ( new_n149_, new_n148_ );
or g074 ( new_n150_, new_n146_, new_n149_ );
and g075 ( new_n151_, new_n145_, new_n150_ );
and g076 ( new_n152_, new_n151_, new_n133_ );
and g077 ( new_n153_, new_n152_, new_n124_ );
not g078 ( new_n154_, keyIn_0_12 );
and g079 ( new_n155_, N223, new_n95_ );
not g080 ( new_n156_, N37 );
and g081 ( new_n157_, new_n156_, N43 );
and g082 ( new_n158_, new_n107_, new_n157_ );
or g083 ( new_n159_, new_n155_, new_n158_ );
or g084 ( new_n160_, new_n159_, new_n154_ );
or g085 ( new_n161_, new_n107_, new_n157_ );
not g086 ( new_n162_, new_n158_ );
and g087 ( new_n163_, new_n162_, new_n161_ );
or g088 ( new_n164_, new_n163_, keyIn_0_12 );
and g089 ( new_n165_, new_n160_, new_n164_ );
not g090 ( new_n166_, keyIn_0_6 );
not g091 ( new_n167_, N47 );
and g092 ( new_n168_, new_n167_, N43 );
and g093 ( new_n169_, new_n168_, new_n166_ );
not g094 ( new_n170_, new_n169_ );
or g095 ( new_n171_, new_n168_, new_n166_ );
and g096 ( new_n172_, new_n170_, new_n171_ );
not g097 ( new_n173_, new_n172_ );
or g098 ( new_n174_, new_n165_, new_n173_ );
not g099 ( new_n175_, keyIn_0_10 );
and g100 ( new_n176_, N223, new_n90_ );
not g101 ( new_n177_, N11 );
and g102 ( new_n178_, new_n177_, N17 );
and g103 ( new_n179_, new_n107_, new_n178_ );
or g104 ( new_n180_, new_n176_, new_n179_ );
or g105 ( new_n181_, new_n180_, new_n175_ );
or g106 ( new_n182_, new_n107_, new_n178_ );
not g107 ( new_n183_, new_n179_ );
and g108 ( new_n184_, new_n183_, new_n182_ );
or g109 ( new_n185_, new_n184_, keyIn_0_10 );
and g110 ( new_n186_, new_n181_, new_n185_ );
not g111 ( new_n187_, N21 );
and g112 ( new_n188_, new_n89_, keyIn_0_1 );
not g113 ( new_n189_, new_n188_ );
or g114 ( new_n190_, new_n89_, keyIn_0_1 );
and g115 ( new_n191_, new_n189_, new_n190_ );
and g116 ( new_n192_, new_n191_, new_n187_ );
not g117 ( new_n193_, new_n192_ );
or g118 ( new_n194_, new_n186_, new_n193_ );
and g119 ( new_n195_, new_n174_, new_n194_ );
and g120 ( new_n196_, N223, new_n79_ );
not g121 ( new_n197_, N63 );
and g122 ( new_n198_, new_n197_, N69 );
and g123 ( new_n199_, new_n107_, new_n198_ );
or g124 ( new_n200_, new_n196_, new_n199_ );
or g125 ( new_n201_, new_n200_, keyIn_0_13 );
not g126 ( new_n202_, keyIn_0_13 );
or g127 ( new_n203_, new_n107_, new_n198_ );
not g128 ( new_n204_, new_n199_ );
and g129 ( new_n205_, new_n204_, new_n203_ );
or g130 ( new_n206_, new_n205_, new_n202_ );
and g131 ( new_n207_, new_n201_, new_n206_ );
not g132 ( new_n208_, N73 );
and g133 ( new_n209_, new_n208_, N69 );
not g134 ( new_n210_, new_n209_ );
or g135 ( new_n211_, new_n207_, new_n210_ );
not g136 ( new_n212_, keyIn_0_18 );
or g137 ( new_n213_, new_n127_, new_n198_ );
not g138 ( new_n214_, N76 );
and g139 ( new_n215_, new_n214_, N82 );
or g140 ( new_n216_, new_n215_, new_n110_ );
or g141 ( new_n217_, new_n213_, new_n216_ );
or g142 ( new_n218_, new_n135_, new_n178_ );
not g143 ( new_n219_, N24 );
and g144 ( new_n220_, new_n219_, N30 );
or g145 ( new_n221_, new_n220_, new_n157_ );
or g146 ( new_n222_, new_n218_, new_n221_ );
or g147 ( new_n223_, new_n217_, new_n222_ );
and g148 ( new_n224_, new_n223_, new_n106_ );
or g149 ( new_n225_, new_n224_, keyIn_0_14 );
not g150 ( new_n226_, keyIn_0_14 );
or g151 ( new_n227_, new_n98_, new_n105_ );
or g152 ( new_n228_, new_n227_, new_n226_ );
and g153 ( new_n229_, new_n225_, new_n228_ );
not g154 ( new_n230_, N112 );
and g155 ( new_n231_, keyIn_0_3, N108 );
not g156 ( new_n232_, new_n231_ );
or g157 ( new_n233_, keyIn_0_3, N108 );
and g158 ( new_n234_, new_n232_, new_n233_ );
not g159 ( new_n235_, new_n234_ );
and g160 ( new_n236_, new_n235_, new_n230_ );
not g161 ( new_n237_, new_n236_ );
or g162 ( new_n238_, new_n229_, new_n237_ );
and g163 ( new_n239_, new_n238_, new_n212_ );
and g164 ( new_n240_, new_n227_, new_n226_ );
and g165 ( new_n241_, new_n224_, keyIn_0_14 );
or g166 ( new_n242_, new_n241_, new_n240_ );
and g167 ( new_n243_, new_n242_, new_n236_ );
and g168 ( new_n244_, new_n243_, keyIn_0_18 );
or g169 ( new_n245_, new_n239_, new_n244_ );
and g170 ( new_n246_, new_n211_, new_n245_ );
and g171 ( new_n247_, new_n195_, new_n246_ );
and g172 ( new_n248_, new_n247_, new_n153_ );
not g173 ( new_n249_, keyIn_0_16 );
not g174 ( new_n250_, keyIn_0_11 );
and g175 ( new_n251_, N223, new_n93_ );
and g176 ( new_n252_, new_n107_, new_n220_ );
or g177 ( new_n253_, new_n251_, new_n252_ );
not g178 ( new_n254_, new_n253_ );
and g179 ( new_n255_, new_n254_, new_n250_ );
and g180 ( new_n256_, new_n253_, keyIn_0_11 );
or g181 ( new_n257_, new_n255_, new_n256_ );
not g182 ( new_n258_, N34 );
and g183 ( new_n259_, new_n258_, N30 );
and g184 ( new_n260_, new_n257_, new_n259_ );
not g185 ( new_n261_, new_n260_ );
and g186 ( new_n262_, new_n261_, new_n249_ );
and g187 ( new_n263_, new_n260_, keyIn_0_16 );
or g188 ( new_n264_, new_n262_, new_n263_ );
and g189 ( new_n265_, new_n248_, new_n264_ );
not g190 ( N329, new_n265_ );
and g191 ( new_n267_, new_n184_, keyIn_0_10 );
and g192 ( new_n268_, new_n180_, new_n175_ );
or g193 ( new_n269_, new_n268_, new_n267_ );
and g194 ( new_n270_, new_n269_, new_n192_ );
and g195 ( new_n271_, new_n265_, new_n270_ );
not g196 ( new_n272_, new_n271_ );
or g197 ( new_n273_, new_n265_, new_n270_ );
not g198 ( new_n274_, N27 );
and g199 ( new_n275_, new_n191_, new_n274_ );
and g200 ( new_n276_, new_n269_, new_n275_ );
and g201 ( new_n277_, new_n273_, new_n276_ );
and g202 ( new_n278_, new_n277_, new_n272_ );
or g203 ( new_n279_, new_n278_, keyIn_0_26 );
not g204 ( new_n280_, new_n279_ );
and g205 ( new_n281_, new_n278_, keyIn_0_26 );
and g206 ( new_n282_, new_n205_, new_n202_ );
and g207 ( new_n283_, new_n200_, keyIn_0_13 );
or g208 ( new_n284_, new_n283_, new_n282_ );
and g209 ( new_n285_, new_n284_, new_n209_ );
or g210 ( new_n286_, new_n265_, new_n285_ );
not g211 ( new_n287_, N79 );
and g212 ( new_n288_, new_n287_, N69 );
and g213 ( new_n289_, new_n284_, new_n288_ );
and g214 ( new_n290_, new_n286_, new_n289_ );
not g215 ( new_n291_, new_n150_ );
or g216 ( new_n292_, new_n265_, new_n291_ );
not g217 ( new_n293_, new_n146_ );
not g218 ( new_n294_, N92 );
and g219 ( new_n295_, new_n294_, N82 );
and g220 ( new_n296_, new_n293_, new_n295_ );
and g221 ( new_n297_, new_n292_, new_n296_ );
or g222 ( new_n298_, new_n290_, new_n297_ );
or g223 ( new_n299_, new_n265_, new_n123_ );
not g224 ( new_n300_, keyIn_0_8 );
not g225 ( new_n301_, N105 );
and g226 ( new_n302_, new_n117_, new_n301_ );
and g227 ( new_n303_, new_n302_, new_n300_ );
not g228 ( new_n304_, new_n303_ );
or g229 ( new_n305_, new_n302_, new_n300_ );
and g230 ( new_n306_, new_n304_, new_n305_ );
and g231 ( new_n307_, new_n306_, new_n111_ );
and g232 ( new_n308_, new_n299_, new_n307_ );
or g233 ( new_n309_, new_n243_, keyIn_0_18 );
or g234 ( new_n310_, new_n238_, new_n212_ );
and g235 ( new_n311_, new_n310_, new_n309_ );
or g236 ( new_n312_, new_n265_, new_n311_ );
not g237 ( new_n313_, keyIn_0_19 );
not g238 ( new_n314_, N115 );
and g239 ( new_n315_, new_n235_, new_n314_ );
and g240 ( new_n316_, new_n242_, new_n315_ );
and g241 ( new_n317_, new_n316_, new_n313_ );
not g242 ( new_n318_, new_n317_ );
or g243 ( new_n319_, new_n316_, new_n313_ );
and g244 ( new_n320_, new_n318_, new_n319_ );
and g245 ( new_n321_, new_n312_, new_n320_ );
or g246 ( new_n322_, new_n308_, new_n321_ );
or g247 ( new_n323_, new_n298_, new_n322_ );
or g248 ( new_n324_, new_n323_, new_n281_ );
or g249 ( new_n325_, new_n324_, new_n280_ );
not g250 ( new_n326_, keyIn_0_22 );
not g251 ( new_n327_, new_n145_ );
and g252 ( new_n328_, new_n265_, new_n327_ );
not g253 ( new_n329_, new_n328_ );
or g254 ( new_n330_, new_n265_, new_n327_ );
and g255 ( new_n331_, new_n329_, new_n330_ );
and g256 ( new_n332_, new_n331_, new_n326_ );
not g257 ( new_n333_, new_n332_ );
or g258 ( new_n334_, new_n331_, new_n326_ );
or g259 ( new_n335_, new_n143_, N14 );
or g260 ( new_n336_, new_n139_, new_n335_ );
not g261 ( new_n337_, new_n336_ );
and g262 ( new_n338_, new_n334_, new_n337_ );
and g263 ( new_n339_, new_n338_, new_n333_ );
not g264 ( new_n340_, new_n133_ );
and g265 ( new_n341_, new_n265_, new_n340_ );
not g266 ( new_n342_, new_n341_ );
or g267 ( new_n343_, new_n265_, new_n340_ );
not g268 ( new_n344_, keyIn_0_21 );
not g269 ( new_n345_, new_n129_ );
not g270 ( new_n346_, N66 );
and g271 ( new_n347_, new_n346_, N56 );
and g272 ( new_n348_, new_n345_, new_n347_ );
not g273 ( new_n349_, new_n348_ );
and g274 ( new_n350_, new_n349_, new_n344_ );
and g275 ( new_n351_, new_n348_, keyIn_0_21 );
or g276 ( new_n352_, new_n350_, new_n351_ );
and g277 ( new_n353_, new_n343_, new_n352_ );
and g278 ( new_n354_, new_n353_, new_n342_ );
not g279 ( new_n355_, keyIn_0_23 );
not g280 ( new_n356_, new_n153_ );
and g281 ( new_n357_, new_n163_, keyIn_0_12 );
and g282 ( new_n358_, new_n159_, new_n154_ );
or g283 ( new_n359_, new_n358_, new_n357_ );
and g284 ( new_n360_, new_n359_, new_n172_ );
or g285 ( new_n361_, new_n360_, new_n270_ );
or g286 ( new_n362_, new_n311_, new_n285_ );
or g287 ( new_n363_, new_n361_, new_n362_ );
or g288 ( new_n364_, new_n363_, new_n356_ );
and g289 ( new_n365_, new_n364_, new_n264_ );
and g290 ( new_n366_, new_n365_, new_n355_ );
not g291 ( new_n367_, new_n366_ );
or g292 ( new_n368_, new_n365_, new_n355_ );
not g293 ( new_n369_, keyIn_0_20 );
not g294 ( new_n370_, new_n255_ );
not g295 ( new_n371_, new_n256_ );
and g296 ( new_n372_, new_n370_, new_n371_ );
not g297 ( new_n373_, keyIn_0_5 );
not g298 ( new_n374_, N40 );
and g299 ( new_n375_, new_n374_, N30 );
and g300 ( new_n376_, new_n375_, new_n373_ );
not g301 ( new_n377_, new_n376_ );
or g302 ( new_n378_, new_n375_, new_n373_ );
and g303 ( new_n379_, new_n377_, new_n378_ );
or g304 ( new_n380_, new_n372_, new_n379_ );
and g305 ( new_n381_, new_n380_, new_n369_ );
not g306 ( new_n382_, new_n381_ );
or g307 ( new_n383_, new_n380_, new_n369_ );
and g308 ( new_n384_, new_n382_, new_n383_ );
and g309 ( new_n385_, new_n368_, new_n384_ );
and g310 ( new_n386_, new_n385_, new_n367_ );
and g311 ( new_n387_, new_n265_, new_n360_ );
not g312 ( new_n388_, new_n387_ );
or g313 ( new_n389_, new_n265_, new_n360_ );
not g314 ( new_n390_, keyIn_0_7 );
not g315 ( new_n391_, N53 );
and g316 ( new_n392_, new_n391_, N43 );
not g317 ( new_n393_, new_n392_ );
and g318 ( new_n394_, new_n393_, new_n390_ );
and g319 ( new_n395_, new_n392_, keyIn_0_7 );
or g320 ( new_n396_, new_n394_, new_n395_ );
and g321 ( new_n397_, new_n359_, new_n396_ );
and g322 ( new_n398_, new_n389_, new_n397_ );
and g323 ( new_n399_, new_n398_, new_n388_ );
or g324 ( new_n400_, new_n386_, new_n399_ );
or g325 ( new_n401_, new_n400_, new_n354_ );
or g326 ( new_n402_, new_n401_, new_n339_ );
or g327 ( N370, new_n402_, new_n325_ );
not g328 ( new_n404_, keyIn_0_29 );
and g329 ( new_n405_, N370, N79 );
or g330 ( new_n406_, new_n405_, keyIn_0_27 );
not g331 ( new_n407_, keyIn_0_27 );
not g332 ( new_n408_, new_n281_ );
not g333 ( new_n409_, new_n290_ );
not g334 ( new_n410_, new_n297_ );
and g335 ( new_n411_, new_n409_, new_n410_ );
not g336 ( new_n412_, new_n308_ );
not g337 ( new_n413_, new_n321_ );
and g338 ( new_n414_, new_n412_, new_n413_ );
and g339 ( new_n415_, new_n411_, new_n414_ );
and g340 ( new_n416_, new_n415_, new_n408_ );
and g341 ( new_n417_, new_n416_, new_n279_ );
and g342 ( new_n418_, N329, new_n145_ );
or g343 ( new_n419_, new_n418_, new_n328_ );
and g344 ( new_n420_, new_n419_, keyIn_0_22 );
or g345 ( new_n421_, new_n420_, new_n336_ );
or g346 ( new_n422_, new_n421_, new_n332_ );
not g347 ( new_n423_, new_n354_ );
or g348 ( new_n424_, new_n260_, keyIn_0_16 );
not g349 ( new_n425_, new_n263_ );
and g350 ( new_n426_, new_n425_, new_n424_ );
or g351 ( new_n427_, new_n248_, new_n426_ );
and g352 ( new_n428_, new_n427_, keyIn_0_23 );
not g353 ( new_n429_, new_n384_ );
or g354 ( new_n430_, new_n428_, new_n429_ );
or g355 ( new_n431_, new_n430_, new_n366_ );
not g356 ( new_n432_, new_n399_ );
and g357 ( new_n433_, new_n432_, new_n431_ );
and g358 ( new_n434_, new_n433_, new_n423_ );
and g359 ( new_n435_, new_n422_, new_n434_ );
and g360 ( new_n436_, new_n435_, new_n417_ );
or g361 ( new_n437_, new_n436_, new_n287_ );
or g362 ( new_n438_, new_n437_, new_n407_ );
and g363 ( new_n439_, new_n406_, new_n438_ );
not g364 ( new_n440_, keyIn_0_24 );
and g365 ( new_n441_, N329, N73 );
and g366 ( new_n442_, new_n441_, new_n440_ );
not g367 ( new_n443_, new_n442_ );
or g368 ( new_n444_, new_n441_, new_n440_ );
and g369 ( new_n445_, new_n107_, keyIn_0_9 );
not g370 ( new_n446_, new_n445_ );
or g371 ( new_n447_, new_n107_, keyIn_0_9 );
and g372 ( new_n448_, new_n446_, new_n447_ );
not g373 ( new_n449_, new_n448_ );
and g374 ( new_n450_, new_n449_, N63 );
or g375 ( new_n451_, new_n450_, new_n78_ );
not g376 ( new_n452_, new_n451_ );
and g377 ( new_n453_, new_n444_, new_n452_ );
and g378 ( new_n454_, new_n453_, new_n443_ );
not g379 ( new_n455_, new_n454_ );
or g380 ( new_n456_, new_n439_, new_n455_ );
or g381 ( new_n457_, new_n456_, new_n404_ );
and g382 ( new_n458_, new_n437_, new_n407_ );
and g383 ( new_n459_, new_n405_, keyIn_0_27 );
or g384 ( new_n460_, new_n459_, new_n458_ );
and g385 ( new_n461_, new_n460_, new_n454_ );
or g386 ( new_n462_, new_n461_, keyIn_0_29 );
and g387 ( new_n463_, new_n457_, new_n462_ );
not g388 ( new_n464_, keyIn_0_28 );
and g389 ( new_n465_, N370, N40 );
and g390 ( new_n466_, N329, N34 );
and g391 ( new_n467_, new_n449_, N24 );
or g392 ( new_n468_, new_n467_, new_n92_ );
or g393 ( new_n469_, new_n466_, new_n468_ );
or g394 ( new_n470_, new_n465_, new_n469_ );
not g395 ( new_n471_, new_n470_ );
and g396 ( new_n472_, new_n471_, new_n464_ );
and g397 ( new_n473_, new_n470_, keyIn_0_28 );
or g398 ( new_n474_, new_n472_, new_n473_ );
and g399 ( new_n475_, N370, N27 );
and g400 ( new_n476_, N329, N21 );
and g401 ( new_n477_, new_n449_, N11 );
or g402 ( new_n478_, new_n477_, new_n89_ );
or g403 ( new_n479_, new_n476_, new_n478_ );
or g404 ( new_n480_, new_n475_, new_n479_ );
not g405 ( new_n481_, new_n480_ );
or g406 ( new_n482_, new_n474_, new_n481_ );
or g407 ( new_n483_, new_n436_, new_n391_ );
and g408 ( new_n484_, N329, N47 );
and g409 ( new_n485_, new_n449_, N37 );
or g410 ( new_n486_, new_n485_, new_n94_ );
or g411 ( new_n487_, new_n484_, new_n486_ );
not g412 ( new_n488_, new_n487_ );
and g413 ( new_n489_, new_n483_, new_n488_ );
or g414 ( new_n490_, new_n436_, new_n346_ );
and g415 ( new_n491_, N329, N60 );
and g416 ( new_n492_, new_n449_, N50 );
or g417 ( new_n493_, new_n492_, new_n76_ );
or g418 ( new_n494_, new_n491_, new_n493_ );
not g419 ( new_n495_, new_n494_ );
and g420 ( new_n496_, new_n490_, new_n495_ );
or g421 ( new_n497_, new_n489_, new_n496_ );
or g422 ( new_n498_, new_n482_, new_n497_ );
or g423 ( new_n499_, new_n436_, new_n314_ );
or g424 ( new_n500_, new_n265_, new_n230_ );
or g425 ( new_n501_, new_n448_, new_n100_ );
and g426 ( new_n502_, new_n501_, N108 );
and g427 ( new_n503_, new_n500_, new_n502_ );
and g428 ( new_n504_, new_n499_, new_n503_ );
and g429 ( new_n505_, N370, N92 );
and g430 ( new_n506_, N329, N86 );
not g431 ( new_n507_, new_n506_ );
not g432 ( new_n508_, keyIn_0_15 );
and g433 ( new_n509_, new_n449_, N76 );
and g434 ( new_n510_, new_n509_, new_n508_ );
not g435 ( new_n511_, new_n510_ );
or g436 ( new_n512_, new_n509_, new_n508_ );
and g437 ( new_n513_, new_n512_, N82 );
and g438 ( new_n514_, new_n513_, new_n511_ );
and g439 ( new_n515_, new_n507_, new_n514_ );
not g440 ( new_n516_, new_n515_ );
or g441 ( new_n517_, new_n505_, new_n516_ );
not g442 ( new_n518_, new_n517_ );
and g443 ( new_n519_, N370, N105 );
not g444 ( new_n520_, new_n519_ );
and g445 ( new_n521_, N329, N99 );
not g446 ( new_n522_, new_n521_ );
and g447 ( new_n523_, new_n522_, keyIn_0_25 );
not g448 ( new_n524_, new_n523_ );
or g449 ( new_n525_, new_n522_, keyIn_0_25 );
and g450 ( new_n526_, new_n449_, N89 );
or g451 ( new_n527_, new_n526_, new_n83_ );
not g452 ( new_n528_, new_n527_ );
and g453 ( new_n529_, new_n525_, new_n528_ );
and g454 ( new_n530_, new_n529_, new_n524_ );
and g455 ( new_n531_, new_n520_, new_n530_ );
or g456 ( new_n532_, new_n518_, new_n531_ );
or g457 ( new_n533_, new_n532_, new_n504_ );
or g458 ( new_n534_, new_n498_, new_n533_ );
or g459 ( new_n535_, new_n534_, new_n463_ );
and g460 ( new_n536_, N370, N14 );
and g461 ( new_n537_, N329, N8 );
and g462 ( new_n538_, new_n449_, N1 );
or g463 ( new_n539_, new_n538_, new_n87_ );
or g464 ( new_n540_, new_n537_, new_n539_ );
or g465 ( new_n541_, new_n536_, new_n540_ );
and g466 ( N421, new_n535_, new_n541_ );
not g467 ( new_n543_, keyIn_0_30 );
not g468 ( new_n544_, new_n498_ );
and g469 ( new_n545_, new_n544_, new_n543_ );
and g470 ( new_n546_, new_n498_, keyIn_0_30 );
or g471 ( N430, new_n545_, new_n546_ );
not g472 ( new_n548_, new_n472_ );
not g473 ( new_n549_, new_n473_ );
and g474 ( new_n550_, new_n548_, new_n549_ );
not g475 ( new_n551_, new_n497_ );
and g476 ( new_n552_, new_n550_, new_n551_ );
and g477 ( new_n553_, new_n463_, new_n552_ );
and g478 ( new_n554_, new_n551_, new_n518_ );
or g479 ( new_n555_, new_n482_, new_n554_ );
or g480 ( N431, new_n553_, new_n555_ );
and g481 ( new_n557_, new_n461_, keyIn_0_29 );
and g482 ( new_n558_, new_n456_, new_n404_ );
or g483 ( new_n559_, new_n558_, new_n557_ );
or g484 ( new_n560_, new_n474_, new_n497_ );
or g485 ( new_n561_, new_n559_, new_n560_ );
and g486 ( new_n562_, new_n531_, new_n517_ );
or g487 ( new_n563_, new_n562_, new_n489_ );
not g488 ( new_n564_, new_n563_ );
or g489 ( new_n565_, new_n564_, new_n474_ );
and g490 ( new_n566_, new_n565_, new_n480_ );
and g491 ( new_n567_, new_n561_, new_n566_ );
and g492 ( new_n568_, new_n567_, keyIn_0_31 );
not g493 ( new_n569_, keyIn_0_31 );
and g494 ( new_n570_, new_n550_, new_n563_ );
or g495 ( new_n571_, new_n570_, new_n481_ );
or g496 ( new_n572_, new_n553_, new_n571_ );
and g497 ( new_n573_, new_n572_, new_n569_ );
or g498 ( N432, new_n568_, new_n573_ );
endmodule