module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n691_, new_n456_, new_n170_, new_n246_, new_n682_, new_n911_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n903_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n912_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n882_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n867_, new_n276_, new_n155_, new_n384_, new_n900_, new_n410_, new_n851_, new_n878_, new_n543_, new_n113_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n897_, new_n379_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n904_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n881_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, N65 );
nor g001 ( new_n107_, new_n106_, N69 );
not g002 ( new_n108_, N69 );
nor g003 ( new_n109_, new_n108_, N65 );
nor g004 ( new_n110_, new_n107_, new_n109_ );
not g005 ( new_n111_, new_n110_ );
nor g006 ( new_n112_, N73, N77 );
nand g007 ( new_n113_, N73, N77 );
not g008 ( new_n114_, new_n113_ );
nor g009 ( new_n115_, new_n114_, new_n112_ );
not g010 ( new_n116_, new_n115_ );
nor g011 ( new_n117_, new_n111_, new_n116_ );
nor g012 ( new_n118_, new_n110_, new_n115_ );
nor g013 ( new_n119_, new_n117_, new_n118_ );
not g014 ( new_n120_, new_n119_ );
not g015 ( new_n121_, N81 );
nor g016 ( new_n122_, new_n121_, N85 );
not g017 ( new_n123_, N85 );
nor g018 ( new_n124_, new_n123_, N81 );
nor g019 ( new_n125_, new_n122_, new_n124_ );
not g020 ( new_n126_, new_n125_ );
nor g021 ( new_n127_, N89, N93 );
nand g022 ( new_n128_, N89, N93 );
not g023 ( new_n129_, new_n128_ );
nor g024 ( new_n130_, new_n129_, new_n127_ );
not g025 ( new_n131_, new_n130_ );
nor g026 ( new_n132_, new_n126_, new_n131_ );
nor g027 ( new_n133_, new_n125_, new_n130_ );
nor g028 ( new_n134_, new_n132_, new_n133_ );
nand g029 ( new_n135_, new_n120_, new_n134_ );
not g030 ( new_n136_, new_n134_ );
nand g031 ( new_n137_, new_n136_, new_n119_ );
nand g032 ( new_n138_, new_n135_, new_n137_ );
nand g033 ( new_n139_, N129, N137 );
nand g034 ( new_n140_, new_n138_, new_n139_ );
nor g035 ( new_n141_, new_n138_, new_n139_ );
not g036 ( new_n142_, new_n141_ );
nand g037 ( new_n143_, new_n142_, new_n140_ );
not g038 ( new_n144_, keyIn_0_9 );
not g039 ( new_n145_, N33 );
nor g040 ( new_n146_, new_n145_, N49 );
not g041 ( new_n147_, N49 );
nor g042 ( new_n148_, new_n147_, N33 );
nor g043 ( new_n149_, new_n146_, new_n148_ );
not g044 ( new_n150_, new_n149_ );
nor g045 ( new_n151_, N1, N17 );
nand g046 ( new_n152_, N1, N17 );
not g047 ( new_n153_, new_n152_ );
nor g048 ( new_n154_, new_n153_, new_n151_ );
not g049 ( new_n155_, new_n154_ );
nor g050 ( new_n156_, new_n150_, new_n155_ );
nor g051 ( new_n157_, new_n149_, new_n154_ );
nor g052 ( new_n158_, new_n156_, new_n157_ );
nor g053 ( new_n159_, new_n158_, new_n144_ );
nand g054 ( new_n160_, new_n158_, new_n144_ );
not g055 ( new_n161_, new_n160_ );
nor g056 ( new_n162_, new_n161_, new_n159_ );
nand g057 ( new_n163_, new_n143_, new_n162_ );
not g058 ( new_n164_, new_n140_ );
nor g059 ( new_n165_, new_n164_, new_n141_ );
not g060 ( new_n166_, new_n162_ );
nand g061 ( new_n167_, new_n165_, new_n166_ );
nand g062 ( new_n168_, new_n167_, new_n163_ );
not g063 ( new_n169_, keyIn_0_19 );
not g064 ( new_n170_, keyIn_0_3 );
nor g065 ( new_n171_, N105, N109 );
nand g066 ( new_n172_, N105, N109 );
not g067 ( new_n173_, new_n172_ );
nor g068 ( new_n174_, new_n173_, new_n171_ );
nor g069 ( new_n175_, new_n174_, new_n170_ );
nand g070 ( new_n176_, new_n174_, new_n170_ );
not g071 ( new_n177_, new_n176_ );
nor g072 ( new_n178_, new_n177_, new_n175_ );
not g073 ( new_n179_, N97 );
nor g074 ( new_n180_, new_n179_, N101 );
not g075 ( new_n181_, N101 );
nor g076 ( new_n182_, new_n181_, N97 );
nor g077 ( new_n183_, new_n180_, new_n182_ );
nor g078 ( new_n184_, new_n178_, new_n183_ );
nand g079 ( new_n185_, new_n178_, new_n183_ );
not g080 ( new_n186_, new_n185_ );
nor g081 ( new_n187_, new_n186_, new_n184_ );
nor g082 ( new_n188_, new_n187_, new_n120_ );
nand g083 ( new_n189_, new_n187_, new_n120_ );
not g084 ( new_n190_, new_n189_ );
nor g085 ( new_n191_, new_n190_, new_n188_ );
nand g086 ( new_n192_, N131, N137 );
not g087 ( new_n193_, new_n192_ );
nand g088 ( new_n194_, new_n191_, new_n193_ );
not g089 ( new_n195_, new_n188_ );
nand g090 ( new_n196_, new_n195_, new_n189_ );
nand g091 ( new_n197_, new_n196_, new_n192_ );
nand g092 ( new_n198_, new_n194_, new_n197_ );
not g093 ( new_n199_, keyIn_0_6 );
nor g094 ( new_n200_, N41, N57 );
nand g095 ( new_n201_, N41, N57 );
not g096 ( new_n202_, new_n201_ );
nor g097 ( new_n203_, new_n202_, new_n200_ );
nor g098 ( new_n204_, new_n203_, new_n199_ );
nand g099 ( new_n205_, new_n203_, new_n199_ );
not g100 ( new_n206_, new_n205_ );
nor g101 ( new_n207_, new_n206_, new_n204_ );
nor g102 ( new_n208_, N9, N25 );
nand g103 ( new_n209_, N9, N25 );
not g104 ( new_n210_, new_n209_ );
nor g105 ( new_n211_, new_n210_, new_n208_ );
nor g106 ( new_n212_, new_n207_, new_n211_ );
nand g107 ( new_n213_, new_n207_, new_n211_ );
not g108 ( new_n214_, new_n213_ );
nor g109 ( new_n215_, new_n214_, new_n212_ );
not g110 ( new_n216_, new_n215_ );
nor g111 ( new_n217_, new_n198_, new_n216_ );
nand g112 ( new_n218_, new_n198_, new_n216_ );
not g113 ( new_n219_, new_n218_ );
nor g114 ( new_n220_, new_n219_, new_n217_ );
not g115 ( new_n221_, keyIn_0_4 );
nor g116 ( new_n222_, N113, N117 );
nand g117 ( new_n223_, N113, N117 );
not g118 ( new_n224_, new_n223_ );
nor g119 ( new_n225_, new_n224_, new_n222_ );
nor g120 ( new_n226_, new_n225_, new_n221_ );
nand g121 ( new_n227_, new_n225_, new_n221_ );
not g122 ( new_n228_, new_n227_ );
nor g123 ( new_n229_, new_n228_, new_n226_ );
not g124 ( new_n230_, new_n229_ );
nor g125 ( new_n231_, N121, N125 );
nand g126 ( new_n232_, N121, N125 );
not g127 ( new_n233_, new_n232_ );
nor g128 ( new_n234_, new_n233_, new_n231_ );
not g129 ( new_n235_, new_n234_ );
nand g130 ( new_n236_, new_n230_, new_n235_ );
not g131 ( new_n237_, new_n236_ );
nor g132 ( new_n238_, new_n230_, new_n235_ );
nor g133 ( new_n239_, new_n237_, new_n238_ );
nand g134 ( new_n240_, new_n239_, new_n136_ );
not g135 ( new_n241_, new_n238_ );
nand g136 ( new_n242_, new_n241_, new_n236_ );
nand g137 ( new_n243_, new_n242_, new_n134_ );
nand g138 ( new_n244_, new_n240_, new_n243_ );
nand g139 ( new_n245_, N132, N137 );
nand g140 ( new_n246_, new_n244_, new_n245_ );
not g141 ( new_n247_, new_n244_ );
not g142 ( new_n248_, new_n245_ );
nand g143 ( new_n249_, new_n247_, new_n248_ );
nand g144 ( new_n250_, new_n249_, new_n246_ );
not g145 ( new_n251_, new_n250_ );
nor g146 ( new_n252_, N45, N61 );
nand g147 ( new_n253_, N45, N61 );
not g148 ( new_n254_, new_n253_ );
nor g149 ( new_n255_, new_n254_, new_n252_ );
not g150 ( new_n256_, new_n255_ );
nor g151 ( new_n257_, N13, N29 );
nand g152 ( new_n258_, N13, N29 );
not g153 ( new_n259_, new_n258_ );
nor g154 ( new_n260_, new_n259_, new_n257_ );
not g155 ( new_n261_, new_n260_ );
nor g156 ( new_n262_, new_n256_, new_n261_ );
nor g157 ( new_n263_, new_n255_, new_n260_ );
nor g158 ( new_n264_, new_n262_, new_n263_ );
nand g159 ( new_n265_, new_n251_, new_n264_ );
not g160 ( new_n266_, new_n264_ );
nand g161 ( new_n267_, new_n250_, new_n266_ );
nand g162 ( new_n268_, new_n265_, new_n267_ );
nand g163 ( new_n269_, new_n268_, new_n220_ );
not g164 ( new_n270_, new_n187_ );
nand g165 ( new_n271_, new_n239_, new_n270_ );
nand g166 ( new_n272_, new_n242_, new_n187_ );
nand g167 ( new_n273_, new_n271_, new_n272_ );
nand g168 ( new_n274_, N130, N137 );
nand g169 ( new_n275_, new_n273_, new_n274_ );
nor g170 ( new_n276_, new_n273_, new_n274_ );
not g171 ( new_n277_, new_n276_ );
nand g172 ( new_n278_, new_n277_, new_n275_ );
nor g173 ( new_n279_, N37, N53 );
nand g174 ( new_n280_, N37, N53 );
not g175 ( new_n281_, new_n280_ );
nor g176 ( new_n282_, new_n281_, new_n279_ );
not g177 ( new_n283_, new_n282_ );
nor g178 ( new_n284_, N5, N21 );
nand g179 ( new_n285_, N5, N21 );
not g180 ( new_n286_, new_n285_ );
nor g181 ( new_n287_, new_n286_, new_n284_ );
not g182 ( new_n288_, new_n287_ );
nor g183 ( new_n289_, new_n283_, new_n288_ );
nor g184 ( new_n290_, new_n282_, new_n287_ );
nor g185 ( new_n291_, new_n289_, new_n290_ );
nand g186 ( new_n292_, new_n278_, new_n291_ );
not g187 ( new_n293_, new_n275_ );
nor g188 ( new_n294_, new_n293_, new_n276_ );
not g189 ( new_n295_, new_n291_ );
nand g190 ( new_n296_, new_n294_, new_n295_ );
nand g191 ( new_n297_, new_n296_, new_n292_ );
not g192 ( new_n298_, keyIn_0_11 );
nor g193 ( new_n299_, new_n168_, new_n298_ );
not g194 ( new_n300_, new_n299_ );
nand g195 ( new_n301_, new_n168_, new_n298_ );
nand g196 ( new_n302_, new_n300_, new_n301_ );
nand g197 ( new_n303_, new_n302_, new_n297_ );
nor g198 ( new_n304_, new_n303_, new_n269_ );
nor g199 ( new_n305_, new_n304_, new_n169_ );
not g200 ( new_n306_, new_n305_ );
not g201 ( new_n307_, new_n198_ );
nand g202 ( new_n308_, new_n307_, new_n215_ );
nand g203 ( new_n309_, new_n308_, new_n218_ );
nor g204 ( new_n310_, new_n250_, new_n266_ );
not g205 ( new_n311_, new_n267_ );
nor g206 ( new_n312_, new_n311_, new_n310_ );
nor g207 ( new_n313_, new_n312_, new_n309_ );
not g208 ( new_n314_, new_n297_ );
not g209 ( new_n315_, new_n301_ );
nor g210 ( new_n316_, new_n315_, new_n299_ );
nor g211 ( new_n317_, new_n314_, new_n316_ );
nand g212 ( new_n318_, new_n317_, new_n313_ );
nor g213 ( new_n319_, new_n318_, keyIn_0_19 );
not g214 ( new_n320_, new_n319_ );
nand g215 ( new_n321_, new_n320_, new_n306_ );
nand g216 ( new_n322_, new_n309_, keyIn_0_12 );
nand g217 ( new_n323_, new_n322_, new_n297_ );
nor g218 ( new_n324_, new_n322_, new_n297_ );
not g219 ( new_n325_, new_n168_ );
nand g220 ( new_n326_, new_n312_, new_n325_ );
nor g221 ( new_n327_, new_n324_, new_n326_ );
nand g222 ( new_n328_, new_n327_, new_n323_ );
nand g223 ( new_n329_, new_n220_, new_n168_ );
nor g224 ( new_n330_, new_n329_, new_n268_ );
nand g225 ( new_n331_, new_n297_, keyIn_0_13 );
not g226 ( new_n332_, new_n331_ );
nor g227 ( new_n333_, new_n297_, keyIn_0_13 );
nor g228 ( new_n334_, new_n332_, new_n333_ );
nand g229 ( new_n335_, new_n334_, new_n330_ );
nand g230 ( new_n336_, new_n328_, new_n335_ );
not g231 ( new_n337_, new_n336_ );
nand g232 ( new_n338_, new_n337_, new_n321_ );
not g233 ( new_n339_, keyIn_0_15 );
not g234 ( new_n340_, keyIn_0_10 );
nor g235 ( new_n341_, N49, N53 );
nand g236 ( new_n342_, N49, N53 );
not g237 ( new_n343_, new_n342_ );
nor g238 ( new_n344_, new_n343_, new_n341_ );
nor g239 ( new_n345_, N57, N61 );
nand g240 ( new_n346_, N57, N61 );
not g241 ( new_n347_, new_n346_ );
nor g242 ( new_n348_, new_n347_, new_n345_ );
nor g243 ( new_n349_, new_n344_, new_n348_ );
nand g244 ( new_n350_, new_n344_, new_n348_ );
not g245 ( new_n351_, new_n350_ );
nor g246 ( new_n352_, new_n351_, new_n349_ );
not g247 ( new_n353_, keyIn_0_0 );
not g248 ( new_n354_, N17 );
not g249 ( new_n355_, N21 );
nand g250 ( new_n356_, new_n354_, new_n355_ );
nand g251 ( new_n357_, N17, N21 );
nand g252 ( new_n358_, new_n356_, new_n357_ );
nand g253 ( new_n359_, new_n358_, new_n353_ );
nor g254 ( new_n360_, N17, N21 );
not g255 ( new_n361_, new_n357_ );
nor g256 ( new_n362_, new_n361_, new_n360_ );
nand g257 ( new_n363_, new_n362_, keyIn_0_0 );
nand g258 ( new_n364_, new_n363_, new_n359_ );
nor g259 ( new_n365_, N25, N29 );
nand g260 ( new_n366_, N25, N29 );
not g261 ( new_n367_, new_n366_ );
nor g262 ( new_n368_, new_n367_, new_n365_ );
nand g263 ( new_n369_, new_n364_, new_n368_ );
nor g264 ( new_n370_, new_n362_, keyIn_0_0 );
nor g265 ( new_n371_, new_n358_, new_n353_ );
nor g266 ( new_n372_, new_n370_, new_n371_ );
not g267 ( new_n373_, new_n368_ );
nand g268 ( new_n374_, new_n372_, new_n373_ );
nand g269 ( new_n375_, new_n374_, new_n369_ );
nand g270 ( new_n376_, new_n375_, new_n352_ );
not g271 ( new_n377_, new_n352_ );
not g272 ( new_n378_, new_n369_ );
nor g273 ( new_n379_, new_n364_, new_n368_ );
nor g274 ( new_n380_, new_n378_, new_n379_ );
nand g275 ( new_n381_, new_n380_, new_n377_ );
nand g276 ( new_n382_, new_n381_, new_n376_ );
nand g277 ( new_n383_, N136, N137 );
nand g278 ( new_n384_, new_n382_, new_n383_ );
not g279 ( new_n385_, new_n376_ );
nor g280 ( new_n386_, new_n375_, new_n352_ );
nor g281 ( new_n387_, new_n385_, new_n386_ );
not g282 ( new_n388_, new_n383_ );
nand g283 ( new_n389_, new_n387_, new_n388_ );
nand g284 ( new_n390_, new_n389_, new_n384_ );
nand g285 ( new_n391_, new_n390_, new_n340_ );
not g286 ( new_n392_, new_n384_ );
nor g287 ( new_n393_, new_n382_, new_n383_ );
nor g288 ( new_n394_, new_n392_, new_n393_ );
nand g289 ( new_n395_, new_n394_, keyIn_0_10 );
nand g290 ( new_n396_, new_n395_, new_n391_ );
nor g291 ( new_n397_, N109, N125 );
nand g292 ( new_n398_, N109, N125 );
not g293 ( new_n399_, new_n398_ );
nor g294 ( new_n400_, new_n399_, new_n397_ );
not g295 ( new_n401_, new_n400_ );
nor g296 ( new_n402_, N77, N93 );
nand g297 ( new_n403_, N77, N93 );
not g298 ( new_n404_, new_n403_ );
nor g299 ( new_n405_, new_n404_, new_n402_ );
not g300 ( new_n406_, new_n405_ );
nor g301 ( new_n407_, new_n401_, new_n406_ );
nor g302 ( new_n408_, new_n400_, new_n405_ );
nor g303 ( new_n409_, new_n407_, new_n408_ );
nand g304 ( new_n410_, new_n396_, new_n409_ );
not g305 ( new_n411_, new_n391_ );
nor g306 ( new_n412_, new_n390_, new_n340_ );
nor g307 ( new_n413_, new_n411_, new_n412_ );
not g308 ( new_n414_, new_n409_ );
nand g309 ( new_n415_, new_n413_, new_n414_ );
nand g310 ( new_n416_, new_n415_, new_n410_ );
nand g311 ( new_n417_, new_n416_, new_n339_ );
not g312 ( new_n418_, new_n417_ );
nor g313 ( new_n419_, new_n416_, new_n339_ );
nor g314 ( new_n420_, new_n418_, new_n419_ );
not g315 ( new_n421_, new_n420_ );
not g316 ( new_n422_, keyIn_0_8 );
not g317 ( new_n423_, N37 );
nand g318 ( new_n424_, new_n423_, N33 );
nand g319 ( new_n425_, new_n145_, N37 );
nand g320 ( new_n426_, new_n424_, new_n425_ );
nand g321 ( new_n427_, new_n426_, keyIn_0_1 );
not g322 ( new_n428_, keyIn_0_1 );
not g323 ( new_n429_, new_n426_ );
nand g324 ( new_n430_, new_n429_, new_n428_ );
nand g325 ( new_n431_, new_n430_, new_n427_ );
not g326 ( new_n432_, N41 );
not g327 ( new_n433_, N45 );
nand g328 ( new_n434_, new_n432_, new_n433_ );
nand g329 ( new_n435_, N41, N45 );
nand g330 ( new_n436_, new_n434_, new_n435_ );
nand g331 ( new_n437_, new_n436_, keyIn_0_2 );
not g332 ( new_n438_, keyIn_0_2 );
nor g333 ( new_n439_, N41, N45 );
not g334 ( new_n440_, new_n435_ );
nor g335 ( new_n441_, new_n440_, new_n439_ );
nand g336 ( new_n442_, new_n441_, new_n438_ );
nand g337 ( new_n443_, new_n442_, new_n437_ );
nor g338 ( new_n444_, new_n431_, new_n443_ );
not g339 ( new_n445_, new_n427_ );
nor g340 ( new_n446_, new_n426_, keyIn_0_1 );
nor g341 ( new_n447_, new_n445_, new_n446_ );
nor g342 ( new_n448_, new_n441_, new_n438_ );
nor g343 ( new_n449_, new_n436_, keyIn_0_2 );
nor g344 ( new_n450_, new_n448_, new_n449_ );
nor g345 ( new_n451_, new_n447_, new_n450_ );
nor g346 ( new_n452_, new_n451_, new_n444_ );
nand g347 ( new_n453_, new_n452_, new_n422_ );
nand g348 ( new_n454_, new_n447_, new_n450_ );
nand g349 ( new_n455_, new_n431_, new_n443_ );
nand g350 ( new_n456_, new_n454_, new_n455_ );
nand g351 ( new_n457_, new_n456_, keyIn_0_8 );
nand g352 ( new_n458_, new_n453_, new_n457_ );
nand g353 ( new_n459_, new_n458_, new_n377_ );
nor g354 ( new_n460_, new_n456_, keyIn_0_8 );
nor g355 ( new_n461_, new_n452_, new_n422_ );
nor g356 ( new_n462_, new_n461_, new_n460_ );
nand g357 ( new_n463_, new_n462_, new_n352_ );
nand g358 ( new_n464_, new_n463_, new_n459_ );
nand g359 ( new_n465_, N134, N137 );
not g360 ( new_n466_, new_n465_ );
nand g361 ( new_n467_, new_n464_, new_n466_ );
not g362 ( new_n468_, new_n459_ );
nor g363 ( new_n469_, new_n458_, new_n377_ );
nor g364 ( new_n470_, new_n468_, new_n469_ );
nand g365 ( new_n471_, new_n470_, new_n465_ );
nand g366 ( new_n472_, new_n471_, new_n467_ );
nor g367 ( new_n473_, N101, N117 );
nand g368 ( new_n474_, N101, N117 );
not g369 ( new_n475_, new_n474_ );
nor g370 ( new_n476_, new_n475_, new_n473_ );
not g371 ( new_n477_, new_n476_ );
nor g372 ( new_n478_, N69, N85 );
nand g373 ( new_n479_, N69, N85 );
not g374 ( new_n480_, new_n479_ );
nor g375 ( new_n481_, new_n480_, new_n478_ );
not g376 ( new_n482_, new_n481_ );
nor g377 ( new_n483_, new_n477_, new_n482_ );
nor g378 ( new_n484_, new_n476_, new_n481_ );
nor g379 ( new_n485_, new_n483_, new_n484_ );
nand g380 ( new_n486_, new_n472_, new_n485_ );
not g381 ( new_n487_, new_n467_ );
nor g382 ( new_n488_, new_n464_, new_n466_ );
nor g383 ( new_n489_, new_n487_, new_n488_ );
not g384 ( new_n490_, new_n485_ );
nand g385 ( new_n491_, new_n489_, new_n490_ );
nand g386 ( new_n492_, new_n491_, new_n486_ );
nand g387 ( new_n493_, new_n492_, keyIn_0_14 );
nor g388 ( new_n494_, new_n492_, keyIn_0_14 );
nor g389 ( new_n495_, N9, N13 );
nand g390 ( new_n496_, N9, N13 );
not g391 ( new_n497_, new_n496_ );
nor g392 ( new_n498_, new_n497_, new_n495_ );
not g393 ( new_n499_, new_n498_ );
nor g394 ( new_n500_, N1, N5 );
nand g395 ( new_n501_, N1, N5 );
not g396 ( new_n502_, new_n501_ );
nor g397 ( new_n503_, new_n502_, new_n500_ );
not g398 ( new_n504_, new_n503_ );
nor g399 ( new_n505_, new_n499_, new_n504_ );
nor g400 ( new_n506_, new_n498_, new_n503_ );
nor g401 ( new_n507_, new_n505_, new_n506_ );
not g402 ( new_n508_, new_n507_ );
nor g403 ( new_n509_, new_n462_, new_n508_ );
nor g404 ( new_n510_, new_n458_, new_n507_ );
nor g405 ( new_n511_, new_n509_, new_n510_ );
nand g406 ( new_n512_, N135, N137 );
nor g407 ( new_n513_, new_n512_, keyIn_0_5 );
nand g408 ( new_n514_, new_n512_, keyIn_0_5 );
not g409 ( new_n515_, new_n514_ );
nor g410 ( new_n516_, new_n515_, new_n513_ );
nor g411 ( new_n517_, new_n511_, new_n516_ );
nand g412 ( new_n518_, new_n458_, new_n507_ );
nand g413 ( new_n519_, new_n462_, new_n508_ );
nand g414 ( new_n520_, new_n519_, new_n518_ );
not g415 ( new_n521_, new_n516_ );
nor g416 ( new_n522_, new_n520_, new_n521_ );
nor g417 ( new_n523_, new_n517_, new_n522_ );
not g418 ( new_n524_, keyIn_0_7 );
nor g419 ( new_n525_, N105, N121 );
nand g420 ( new_n526_, N105, N121 );
not g421 ( new_n527_, new_n526_ );
nor g422 ( new_n528_, new_n527_, new_n525_ );
nor g423 ( new_n529_, new_n528_, new_n524_ );
nand g424 ( new_n530_, new_n528_, new_n524_ );
not g425 ( new_n531_, new_n530_ );
nor g426 ( new_n532_, new_n531_, new_n529_ );
nor g427 ( new_n533_, N73, N89 );
nand g428 ( new_n534_, N73, N89 );
not g429 ( new_n535_, new_n534_ );
nor g430 ( new_n536_, new_n535_, new_n533_ );
nor g431 ( new_n537_, new_n532_, new_n536_ );
nand g432 ( new_n538_, new_n532_, new_n536_ );
not g433 ( new_n539_, new_n538_ );
nor g434 ( new_n540_, new_n539_, new_n537_ );
not g435 ( new_n541_, new_n540_ );
nand g436 ( new_n542_, new_n523_, new_n541_ );
nand g437 ( new_n543_, new_n520_, new_n521_ );
nand g438 ( new_n544_, new_n511_, new_n516_ );
nand g439 ( new_n545_, new_n544_, new_n543_ );
nand g440 ( new_n546_, new_n545_, new_n540_ );
nand g441 ( new_n547_, new_n542_, new_n546_ );
nand g442 ( new_n548_, new_n375_, new_n507_ );
not g443 ( new_n549_, new_n548_ );
nor g444 ( new_n550_, new_n375_, new_n507_ );
nor g445 ( new_n551_, new_n549_, new_n550_ );
not g446 ( new_n552_, new_n551_ );
nand g447 ( new_n553_, N133, N137 );
nand g448 ( new_n554_, new_n552_, new_n553_ );
not g449 ( new_n555_, new_n553_ );
nand g450 ( new_n556_, new_n551_, new_n555_ );
nand g451 ( new_n557_, new_n554_, new_n556_ );
nor g452 ( new_n558_, new_n179_, N113 );
not g453 ( new_n559_, N113 );
nor g454 ( new_n560_, new_n559_, N97 );
nor g455 ( new_n561_, new_n558_, new_n560_ );
not g456 ( new_n562_, new_n561_ );
nor g457 ( new_n563_, N65, N81 );
nand g458 ( new_n564_, N65, N81 );
not g459 ( new_n565_, new_n564_ );
nor g460 ( new_n566_, new_n565_, new_n563_ );
not g461 ( new_n567_, new_n566_ );
nor g462 ( new_n568_, new_n562_, new_n567_ );
nor g463 ( new_n569_, new_n561_, new_n566_ );
nor g464 ( new_n570_, new_n568_, new_n569_ );
not g465 ( new_n571_, new_n570_ );
nor g466 ( new_n572_, new_n557_, new_n571_ );
nand g467 ( new_n573_, new_n557_, new_n571_ );
not g468 ( new_n574_, new_n573_ );
nor g469 ( new_n575_, new_n574_, new_n572_ );
not g470 ( new_n576_, new_n575_ );
nor g471 ( new_n577_, new_n547_, new_n576_ );
not g472 ( new_n578_, new_n577_ );
nor g473 ( new_n579_, new_n578_, new_n494_ );
nand g474 ( new_n580_, new_n579_, new_n493_ );
nor g475 ( new_n581_, new_n580_, new_n421_ );
nand g476 ( new_n582_, new_n338_, new_n581_ );
nand g477 ( new_n583_, new_n582_, keyIn_0_24 );
not g478 ( new_n584_, keyIn_0_24 );
nor g479 ( new_n585_, new_n319_, new_n305_ );
nor g480 ( new_n586_, new_n585_, new_n336_ );
not g481 ( new_n587_, new_n581_ );
nor g482 ( new_n588_, new_n587_, new_n586_ );
nand g483 ( new_n589_, new_n588_, new_n584_ );
nand g484 ( new_n590_, new_n589_, new_n583_ );
nand g485 ( new_n591_, new_n590_, new_n168_ );
nand g486 ( new_n592_, new_n591_, N1 );
not g487 ( new_n593_, N1 );
not g488 ( new_n594_, new_n591_ );
nand g489 ( new_n595_, new_n594_, new_n593_ );
nand g490 ( N724, new_n595_, new_n592_ );
nand g491 ( new_n597_, new_n590_, new_n314_ );
nand g492 ( new_n598_, new_n597_, N5 );
not g493 ( new_n599_, N5 );
not g494 ( new_n600_, new_n597_ );
nand g495 ( new_n601_, new_n600_, new_n599_ );
nand g496 ( N725, new_n601_, new_n598_ );
not g497 ( new_n603_, keyIn_0_30 );
nand g498 ( new_n604_, new_n590_, new_n309_ );
nand g499 ( new_n605_, new_n604_, N9 );
not g500 ( new_n606_, new_n605_ );
nor g501 ( new_n607_, new_n604_, N9 );
nor g502 ( new_n608_, new_n606_, new_n607_ );
nand g503 ( new_n609_, new_n608_, new_n603_ );
not g504 ( new_n610_, new_n608_ );
nand g505 ( new_n611_, new_n610_, keyIn_0_30 );
nand g506 ( N726, new_n611_, new_n609_ );
not g507 ( new_n613_, keyIn_0_31 );
nor g508 ( new_n614_, new_n420_, new_n584_ );
nor g509 ( new_n615_, new_n590_, new_n614_ );
nor g510 ( new_n616_, new_n615_, new_n312_ );
nand g511 ( new_n617_, new_n616_, N13 );
not g512 ( new_n618_, N13 );
not g513 ( new_n619_, new_n590_ );
not g514 ( new_n620_, new_n614_ );
nand g515 ( new_n621_, new_n619_, new_n620_ );
nand g516 ( new_n622_, new_n621_, new_n268_ );
nand g517 ( new_n623_, new_n622_, new_n618_ );
nand g518 ( new_n624_, new_n623_, new_n617_ );
nand g519 ( new_n625_, new_n624_, new_n613_ );
nor g520 ( new_n626_, new_n622_, new_n618_ );
nor g521 ( new_n627_, new_n616_, N13 );
nor g522 ( new_n628_, new_n626_, new_n627_ );
nand g523 ( new_n629_, new_n628_, keyIn_0_31 );
nand g524 ( N727, new_n629_, new_n625_ );
nor g525 ( new_n631_, new_n413_, new_n414_ );
nor g526 ( new_n632_, new_n396_, new_n409_ );
nor g527 ( new_n633_, new_n631_, new_n632_ );
nand g528 ( new_n634_, new_n633_, new_n547_ );
nor g529 ( new_n635_, new_n492_, new_n576_ );
not g530 ( new_n636_, new_n635_ );
nor g531 ( new_n637_, new_n636_, new_n634_ );
nand g532 ( new_n638_, new_n338_, new_n637_ );
nor g533 ( new_n639_, new_n638_, new_n325_ );
not g534 ( new_n640_, new_n639_ );
nand g535 ( new_n641_, new_n640_, N17 );
nand g536 ( new_n642_, new_n639_, new_n354_ );
nand g537 ( N728, new_n641_, new_n642_ );
nor g538 ( new_n644_, new_n638_, new_n297_ );
not g539 ( new_n645_, new_n644_ );
nand g540 ( new_n646_, new_n645_, N21 );
nand g541 ( new_n647_, new_n644_, new_n355_ );
nand g542 ( N729, new_n646_, new_n647_ );
not g543 ( new_n649_, keyIn_0_25 );
nor g544 ( new_n650_, new_n638_, new_n220_ );
not g545 ( new_n651_, new_n650_ );
nor g546 ( new_n652_, new_n651_, new_n649_ );
nor g547 ( new_n653_, new_n650_, keyIn_0_25 );
nor g548 ( new_n654_, new_n652_, new_n653_ );
not g549 ( new_n655_, new_n654_ );
nand g550 ( new_n656_, new_n655_, N25 );
not g551 ( new_n657_, N25 );
nand g552 ( new_n658_, new_n654_, new_n657_ );
nand g553 ( N730, new_n656_, new_n658_ );
not g554 ( new_n660_, N29 );
not g555 ( new_n661_, keyIn_0_26 );
nor g556 ( new_n662_, new_n638_, new_n312_ );
not g557 ( new_n663_, new_n662_ );
nor g558 ( new_n664_, new_n663_, new_n661_ );
nor g559 ( new_n665_, new_n662_, keyIn_0_26 );
nor g560 ( new_n666_, new_n664_, new_n665_ );
not g561 ( new_n667_, new_n666_ );
nand g562 ( new_n668_, new_n667_, new_n660_ );
nand g563 ( new_n669_, new_n666_, N29 );
nand g564 ( N731, new_n668_, new_n669_ );
nor g565 ( new_n671_, new_n489_, new_n490_ );
nor g566 ( new_n672_, new_n472_, new_n485_ );
nor g567 ( new_n673_, new_n671_, new_n672_ );
nor g568 ( new_n674_, new_n586_, new_n673_ );
not g569 ( new_n675_, new_n674_ );
nor g570 ( new_n676_, new_n633_, new_n547_ );
nor g571 ( new_n677_, new_n575_, keyIn_0_16 );
nand g572 ( new_n678_, new_n575_, keyIn_0_16 );
not g573 ( new_n679_, new_n678_ );
nor g574 ( new_n680_, new_n679_, new_n677_ );
nand g575 ( new_n681_, new_n680_, new_n676_ );
nor g576 ( new_n682_, new_n675_, new_n681_ );
not g577 ( new_n683_, new_n682_ );
nor g578 ( new_n684_, new_n683_, new_n325_ );
not g579 ( new_n685_, new_n684_ );
nand g580 ( new_n686_, new_n685_, N33 );
nand g581 ( new_n687_, new_n684_, new_n145_ );
nand g582 ( N732, new_n686_, new_n687_ );
nor g583 ( new_n689_, new_n683_, new_n297_ );
not g584 ( new_n690_, new_n689_ );
nand g585 ( new_n691_, new_n690_, N37 );
nand g586 ( new_n692_, new_n689_, new_n423_ );
nand g587 ( N733, new_n691_, new_n692_ );
nor g588 ( new_n694_, new_n683_, new_n220_ );
not g589 ( new_n695_, new_n694_ );
nand g590 ( new_n696_, new_n695_, N41 );
nand g591 ( new_n697_, new_n694_, new_n432_ );
nand g592 ( N734, new_n696_, new_n697_ );
nor g593 ( new_n699_, new_n683_, new_n312_ );
not g594 ( new_n700_, new_n699_ );
nand g595 ( new_n701_, new_n700_, N45 );
nand g596 ( new_n702_, new_n699_, new_n433_ );
nand g597 ( N735, new_n701_, new_n702_ );
nor g598 ( new_n704_, new_n575_, keyIn_0_17 );
nand g599 ( new_n705_, new_n575_, keyIn_0_17 );
not g600 ( new_n706_, new_n705_ );
nor g601 ( new_n707_, new_n706_, new_n704_ );
nor g602 ( new_n708_, new_n707_, new_n634_ );
nand g603 ( new_n709_, new_n674_, new_n708_ );
nor g604 ( new_n710_, new_n709_, new_n325_ );
not g605 ( new_n711_, new_n710_ );
nand g606 ( new_n712_, new_n711_, N49 );
nand g607 ( new_n713_, new_n710_, new_n147_ );
nand g608 ( N736, new_n712_, new_n713_ );
nor g609 ( new_n715_, new_n709_, new_n297_ );
not g610 ( new_n716_, new_n715_ );
nand g611 ( new_n717_, new_n716_, N53 );
not g612 ( new_n718_, N53 );
nand g613 ( new_n719_, new_n715_, new_n718_ );
nand g614 ( N737, new_n717_, new_n719_ );
nor g615 ( new_n721_, new_n709_, new_n220_ );
not g616 ( new_n722_, new_n721_ );
nand g617 ( new_n723_, new_n722_, N57 );
not g618 ( new_n724_, N57 );
nand g619 ( new_n725_, new_n721_, new_n724_ );
nand g620 ( N738, new_n723_, new_n725_ );
nor g621 ( new_n727_, new_n709_, new_n312_ );
not g622 ( new_n728_, new_n727_ );
nand g623 ( new_n729_, new_n728_, N61 );
not g624 ( new_n730_, N61 );
nand g625 ( new_n731_, new_n727_, new_n730_ );
nand g626 ( N739, new_n729_, new_n731_ );
nand g627 ( new_n733_, new_n673_, new_n576_ );
nor g628 ( new_n734_, new_n733_, new_n634_ );
nor g629 ( new_n735_, new_n734_, keyIn_0_20 );
nand g630 ( new_n736_, new_n547_, keyIn_0_18 );
nor g631 ( new_n737_, new_n547_, keyIn_0_18 );
not g632 ( new_n738_, new_n737_ );
nand g633 ( new_n739_, new_n738_, new_n736_ );
nand g634 ( new_n740_, new_n635_, new_n416_ );
not g635 ( new_n741_, new_n740_ );
nand g636 ( new_n742_, new_n741_, new_n739_ );
nand g637 ( new_n743_, new_n734_, keyIn_0_20 );
nand g638 ( new_n744_, new_n742_, new_n743_ );
nor g639 ( new_n745_, new_n744_, new_n735_ );
not g640 ( new_n746_, keyIn_0_21 );
nor g641 ( new_n747_, new_n545_, new_n540_ );
nor g642 ( new_n748_, new_n523_, new_n541_ );
nor g643 ( new_n749_, new_n748_, new_n747_ );
nand g644 ( new_n750_, new_n749_, new_n416_ );
nor g645 ( new_n751_, new_n733_, new_n750_ );
nand g646 ( new_n752_, new_n751_, new_n746_ );
nor g647 ( new_n753_, new_n492_, new_n575_ );
nand g648 ( new_n754_, new_n676_, new_n753_ );
nand g649 ( new_n755_, new_n754_, keyIn_0_21 );
nand g650 ( new_n756_, new_n752_, new_n755_ );
nand g651 ( new_n757_, new_n492_, new_n576_ );
not g652 ( new_n758_, new_n757_ );
nor g653 ( new_n759_, new_n749_, new_n633_ );
nand g654 ( new_n760_, new_n758_, new_n759_ );
nand g655 ( new_n761_, new_n760_, keyIn_0_22 );
not g656 ( new_n762_, keyIn_0_22 );
nand g657 ( new_n763_, new_n547_, new_n416_ );
nor g658 ( new_n764_, new_n757_, new_n763_ );
nand g659 ( new_n765_, new_n764_, new_n762_ );
nand g660 ( new_n766_, new_n761_, new_n765_ );
nand g661 ( new_n767_, new_n756_, new_n766_ );
not g662 ( new_n768_, new_n767_ );
nand g663 ( new_n769_, new_n768_, new_n745_ );
nand g664 ( new_n770_, new_n769_, keyIn_0_23 );
not g665 ( new_n771_, keyIn_0_23 );
not g666 ( new_n772_, new_n735_ );
not g667 ( new_n773_, keyIn_0_18 );
nor g668 ( new_n774_, new_n749_, new_n773_ );
nor g669 ( new_n775_, new_n774_, new_n737_ );
nor g670 ( new_n776_, new_n775_, new_n740_ );
not g671 ( new_n777_, keyIn_0_20 );
nor g672 ( new_n778_, new_n749_, new_n416_ );
nand g673 ( new_n779_, new_n778_, new_n753_ );
nor g674 ( new_n780_, new_n779_, new_n777_ );
nor g675 ( new_n781_, new_n776_, new_n780_ );
nand g676 ( new_n782_, new_n781_, new_n772_ );
nor g677 ( new_n783_, new_n782_, new_n767_ );
nand g678 ( new_n784_, new_n783_, new_n771_ );
nand g679 ( new_n785_, new_n770_, new_n784_ );
nand g680 ( new_n786_, new_n312_, new_n309_ );
nor g681 ( new_n787_, new_n314_, new_n325_ );
not g682 ( new_n788_, new_n787_ );
nor g683 ( new_n789_, new_n788_, new_n786_ );
nand g684 ( new_n790_, new_n785_, new_n789_ );
nor g685 ( new_n791_, new_n790_, new_n576_ );
not g686 ( new_n792_, new_n791_ );
nand g687 ( new_n793_, new_n792_, N65 );
nand g688 ( new_n794_, new_n791_, new_n106_ );
nand g689 ( N740, new_n793_, new_n794_ );
nor g690 ( new_n796_, new_n790_, new_n673_ );
not g691 ( new_n797_, new_n796_ );
nand g692 ( new_n798_, new_n797_, N69 );
nand g693 ( new_n799_, new_n796_, new_n108_ );
nand g694 ( N741, new_n798_, new_n799_ );
nor g695 ( new_n801_, new_n790_, new_n547_ );
not g696 ( new_n802_, new_n801_ );
nand g697 ( new_n803_, new_n802_, N73 );
not g698 ( new_n804_, N73 );
nand g699 ( new_n805_, new_n801_, new_n804_ );
nand g700 ( N742, new_n803_, new_n805_ );
nor g701 ( new_n807_, new_n790_, new_n416_ );
not g702 ( new_n808_, new_n807_ );
nand g703 ( new_n809_, new_n808_, N77 );
not g704 ( new_n810_, N77 );
nand g705 ( new_n811_, new_n807_, new_n810_ );
nand g706 ( N743, new_n809_, new_n811_ );
nor g707 ( new_n813_, new_n788_, new_n269_ );
nand g708 ( new_n814_, new_n785_, new_n813_ );
nor g709 ( new_n815_, new_n814_, new_n576_ );
not g710 ( new_n816_, new_n815_ );
nand g711 ( new_n817_, new_n816_, N81 );
nand g712 ( new_n818_, new_n815_, new_n121_ );
nand g713 ( N744, new_n817_, new_n818_ );
not g714 ( new_n820_, keyIn_0_27 );
nand g715 ( new_n821_, new_n785_, new_n492_ );
not g716 ( new_n822_, new_n821_ );
nand g717 ( new_n823_, new_n822_, new_n813_ );
nand g718 ( new_n824_, new_n823_, new_n820_ );
not g719 ( new_n825_, new_n813_ );
nor g720 ( new_n826_, new_n821_, new_n825_ );
nand g721 ( new_n827_, new_n826_, keyIn_0_27 );
nand g722 ( new_n828_, new_n824_, new_n827_ );
nand g723 ( new_n829_, new_n828_, new_n123_ );
nor g724 ( new_n830_, new_n826_, keyIn_0_27 );
nor g725 ( new_n831_, new_n823_, new_n820_ );
nor g726 ( new_n832_, new_n831_, new_n830_ );
nand g727 ( new_n833_, new_n832_, N85 );
nand g728 ( N745, new_n833_, new_n829_ );
nor g729 ( new_n835_, new_n814_, new_n547_ );
not g730 ( new_n836_, new_n835_ );
nand g731 ( new_n837_, new_n836_, N89 );
not g732 ( new_n838_, N89 );
nand g733 ( new_n839_, new_n835_, new_n838_ );
nand g734 ( N746, new_n837_, new_n839_ );
nor g735 ( new_n841_, new_n814_, new_n416_ );
not g736 ( new_n842_, new_n841_ );
nand g737 ( new_n843_, new_n842_, N93 );
not g738 ( new_n844_, N93 );
nand g739 ( new_n845_, new_n841_, new_n844_ );
nand g740 ( N747, new_n843_, new_n845_ );
nor g741 ( new_n847_, new_n297_, new_n168_ );
not g742 ( new_n848_, new_n847_ );
nor g743 ( new_n849_, new_n848_, new_n786_ );
nand g744 ( new_n850_, new_n785_, new_n849_ );
nor g745 ( new_n851_, new_n850_, new_n576_ );
not g746 ( new_n852_, new_n851_ );
nand g747 ( new_n853_, new_n852_, N97 );
nand g748 ( new_n854_, new_n851_, new_n179_ );
nand g749 ( N748, new_n853_, new_n854_ );
nor g750 ( new_n856_, new_n850_, new_n673_ );
not g751 ( new_n857_, new_n856_ );
nand g752 ( new_n858_, new_n857_, N101 );
nand g753 ( new_n859_, new_n856_, new_n181_ );
nand g754 ( N749, new_n858_, new_n859_ );
nor g755 ( new_n861_, new_n850_, new_n547_ );
not g756 ( new_n862_, new_n861_ );
nand g757 ( new_n863_, new_n862_, N105 );
not g758 ( new_n864_, N105 );
nand g759 ( new_n865_, new_n861_, new_n864_ );
nand g760 ( N750, new_n863_, new_n865_ );
not g761 ( new_n867_, N109 );
not g762 ( new_n868_, new_n850_ );
nand g763 ( new_n869_, new_n868_, new_n633_ );
nand g764 ( new_n870_, new_n869_, keyIn_0_28 );
not g765 ( new_n871_, keyIn_0_28 );
nor g766 ( new_n872_, new_n850_, new_n416_ );
nand g767 ( new_n873_, new_n872_, new_n871_ );
nand g768 ( new_n874_, new_n870_, new_n873_ );
nand g769 ( new_n875_, new_n874_, new_n867_ );
nor g770 ( new_n876_, new_n872_, new_n871_ );
nor g771 ( new_n877_, new_n869_, keyIn_0_28 );
nor g772 ( new_n878_, new_n877_, new_n876_ );
nand g773 ( new_n879_, new_n878_, N109 );
nand g774 ( N751, new_n879_, new_n875_ );
nor g775 ( new_n881_, new_n848_, new_n269_ );
nand g776 ( new_n882_, new_n785_, new_n881_ );
nor g777 ( new_n883_, new_n882_, new_n576_ );
not g778 ( new_n884_, new_n883_ );
nand g779 ( new_n885_, new_n884_, N113 );
nand g780 ( new_n886_, new_n883_, new_n559_ );
nand g781 ( N752, new_n885_, new_n886_ );
nand g782 ( new_n888_, new_n822_, new_n881_ );
nand g783 ( new_n889_, new_n888_, keyIn_0_29 );
not g784 ( new_n890_, keyIn_0_29 );
not g785 ( new_n891_, new_n881_ );
nor g786 ( new_n892_, new_n821_, new_n891_ );
nand g787 ( new_n893_, new_n892_, new_n890_ );
nand g788 ( new_n894_, new_n889_, new_n893_ );
nand g789 ( new_n895_, new_n894_, N117 );
not g790 ( new_n896_, N117 );
nor g791 ( new_n897_, new_n892_, new_n890_ );
nor g792 ( new_n898_, new_n888_, keyIn_0_29 );
nor g793 ( new_n899_, new_n898_, new_n897_ );
nand g794 ( new_n900_, new_n899_, new_n896_ );
nand g795 ( N753, new_n900_, new_n895_ );
nor g796 ( new_n902_, new_n882_, new_n547_ );
not g797 ( new_n903_, new_n902_ );
nand g798 ( new_n904_, new_n903_, N121 );
not g799 ( new_n905_, N121 );
nand g800 ( new_n906_, new_n902_, new_n905_ );
nand g801 ( N754, new_n904_, new_n906_ );
nor g802 ( new_n908_, new_n882_, new_n416_ );
not g803 ( new_n909_, new_n908_ );
nand g804 ( new_n910_, new_n909_, N125 );
not g805 ( new_n911_, N125 );
nand g806 ( new_n912_, new_n908_, new_n911_ );
nand g807 ( N755, new_n910_, new_n912_ );
endmodule