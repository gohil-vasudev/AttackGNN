module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n1359_, new_n595_, new_n1233_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n608_, new_n501_, new_n1157_, new_n1345_, new_n421_, new_n777_, new_n1048_, new_n885_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n1327_, new_n566_, new_n641_, new_n339_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n1351_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n728_, new_n1071_, new_n1294_, new_n894_, new_n853_, new_n695_, new_n660_, new_n1311_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n1213_, new_n752_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n721_, new_n504_, new_n742_, new_n892_, new_n472_, new_n873_, new_n1167_, new_n1300_, new_n774_, new_n792_, new_n953_, new_n257_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n983_, new_n822_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n655_, new_n1054_, new_n630_, new_n385_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n297_, new_n565_, new_n1196_, new_n1366_, new_n511_, new_n303_, new_n325_, new_n1285_, new_n1031_, new_n1216_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n324_, new_n960_, new_n491_, new_n549_, new_n676_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n1362_, new_n497_, new_n816_, new_n1355_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1062_, new_n506_, new_n680_, new_n872_, new_n981_, new_n1275_, new_n1277_, new_n1198_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n1333_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n267_, new_n473_, new_n1147_, new_n1229_, new_n969_, new_n334_, new_n331_, new_n835_, new_n1234_, new_n1360_, new_n378_, new_n621_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1321_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n1315_, new_n1003_, new_n696_, new_n1039_, new_n1365_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n729_, new_n1111_, new_n1218_, new_n1346_, new_n559_, new_n1201_, new_n1282_, new_n762_, new_n1349_, new_n1193_, new_n1187_, new_n1205_, new_n1154_, new_n1253_, new_n295_, new_n1256_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n1032_, new_n867_, new_n954_, new_n901_, new_n1171_, new_n276_, new_n688_, new_n1255_, new_n410_, new_n985_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n296_, new_n661_, new_n797_, new_n232_, new_n1358_, new_n724_, new_n1070_, new_n1109_, new_n261_, new_n672_, new_n1269_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n604_, new_n1104_, new_n571_, new_n758_, new_n328_, new_n460_, new_n1267_, new_n1299_, new_n380_, new_n1079_, new_n861_, new_n1252_, new_n352_, new_n931_, new_n575_, new_n562_, new_n944_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n963_, new_n586_, new_n1325_, new_n993_, new_n1191_, new_n1357_, new_n824_, new_n717_, new_n403_, new_n475_, new_n868_, new_n1242_, new_n858_, new_n1343_, new_n936_, new_n411_, new_n1016_, new_n673_, new_n1144_, new_n407_, new_n666_, new_n1290_, new_n736_, new_n879_, new_n513_, new_n558_, new_n219_, new_n313_, new_n382_, new_n239_, new_n718_, new_n1310_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n1040_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n345_, new_n499_, new_n255_, new_n533_, new_n1130_, new_n795_, new_n459_, new_n1122_, new_n1185_, new_n1240_, new_n354_, new_n1174_, new_n968_, new_n613_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n591_, new_n837_, new_n801_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1334_, new_n531_, new_n593_, new_n974_, new_n252_, new_n1248_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n470_, new_n769_, new_n433_, new_n871_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1367_, new_n278_, new_n304_, new_n1052_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1220_, new_n989_, new_n1117_, new_n644_, new_n836_, new_n1116_, new_n904_, new_n1276_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n818_, new_n881_, new_n1268_, new_n640_, new_n684_, new_n1274_, new_n754_, new_n653_, new_n377_, new_n905_, new_n1258_, new_n375_, new_n962_, new_n760_, new_n627_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1353_, new_n1153_, new_n357_, new_n1339_, new_n320_, new_n780_, new_n984_, new_n1183_, new_n643_, new_n1316_, new_n1338_, new_n1230_, new_n1027_, new_n610_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1165_, new_n1259_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n770_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n889_, new_n536_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n1249_, new_n1354_, new_n955_, new_n847_, new_n250_, new_n888_, new_n288_, new_n1340_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1361_, new_n738_, new_n941_, new_n827_, new_n1356_, new_n1363_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n1211_, new_n1207_, new_n1176_, new_n601_, new_n842_, new_n1057_, new_n682_, new_n1075_, new_n812_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n1342_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n413_, new_n442_, new_n677_, new_n642_, new_n462_, new_n603_, new_n564_, new_n761_, new_n840_, new_n735_, new_n1283_, new_n898_, new_n799_, new_n1304_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n862_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n1264_, new_n215_, new_n1319_, new_n626_, new_n959_, new_n990_, new_n716_, new_n701_, new_n1238_, new_n1058_, new_n1162_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n414_, new_n1101_, new_n1250_, new_n315_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n281_, new_n430_, new_n844_, new_n482_, new_n1302_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n1297_, new_n1257_, new_n1306_, new_n988_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n906_, new_n361_, new_n764_, new_n683_, new_n463_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n1292_, new_n517_, new_n609_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1051_, new_n899_, new_n1053_, new_n492_, new_n1200_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1219_, new_n920_, new_n1121_, new_n1341_, new_n820_, new_n771_, new_n979_, new_n508_, new_n714_, new_n1280_, new_n1007_, new_n1241_, new_n882_, new_n1145_, new_n929_, new_n986_, new_n314_, new_n1159_, new_n1337_, new_n216_, new_n1348_, new_n917_, new_n1322_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n541_, new_n447_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n1247_, new_n465_, new_n739_, new_n783_, new_n263_, new_n341_, new_n996_, new_n1318_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n848_, new_n277_, new_n1245_, new_n663_, new_n579_, new_n286_, new_n1254_, new_n438_, new_n1344_, new_n939_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n397_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n948_, new_n1231_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n457_, new_n1301_, new_n1128_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1161_, new_n1329_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n1000_, new_n633_, new_n784_, new_n1273_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n1166_, new_n259_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n693_, new_n1272_, new_n1287_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1289_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n578_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n1178_, new_n270_, new_n570_, new_n598_, new_n893_, new_n520_, new_n1001_, new_n1347_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n1286_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n1326_, new_n592_, new_n726_, new_n1263_, new_n231_, new_n583_, new_n617_, new_n1080_, new_n1279_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n1155_, new_n1186_, new_n1261_, new_n225_, new_n1246_, new_n922_, new_n387_, new_n476_, new_n987_, new_n949_, new_n221_, new_n243_, new_n450_, new_n1179_, new_n298_, new_n1088_, new_n1148_, new_n1146_, new_n569_, new_n555_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n623_, new_n446_, new_n316_, new_n590_, new_n826_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n1350_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n307_, new_n1181_, new_n597_, new_n1093_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1296_, new_n435_, new_n1309_, new_n1010_, new_n776_, new_n687_, new_n370_, new_n1029_, new_n638_, new_n523_, new_n909_, new_n788_, new_n841_, new_n1204_, new_n1112_, new_n711_, new_n1156_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n645_, new_n1096_, new_n1087_, new_n723_, new_n756_, new_n823_, new_n574_, new_n928_, new_n319_, new_n1008_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n1291_, new_n247_, new_n539_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n294_, new_n1295_, new_n1173_, new_n704_, new_n1189_, new_n1197_, new_n1312_, new_n474_, new_n1223_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1243_, new_n1077_, new_n490_, new_n1100_, new_n865_, new_n358_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n947_, new_n994_, new_n982_, new_n964_, new_n1078_, new_n551_, new_n279_, new_n455_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n464_, new_n573_, new_n765_, new_n1314_, new_n1103_;

not g0000 ( new_n215_, N75 );
nand g0001 ( new_n216_, N29, N42 );
nor g0002 ( N388, new_n216_, new_n215_ );
not g0003 ( new_n218_, N80 );
nand g0004 ( new_n219_, N29, N36 );
nor g0005 ( N389, new_n219_, new_n218_ );
not g0006 ( new_n221_, N42 );
nor g0007 ( N390, new_n219_, new_n221_ );
nand g0008 ( new_n223_, N85, N86 );
not g0009 ( N391, new_n223_ );
not g0010 ( new_n225_, N17 );
nand g0011 ( new_n226_, N1, N8 );
not g0012 ( new_n227_, new_n226_ );
nand g0013 ( new_n228_, new_n227_, N13 );
nor g0014 ( N418, new_n228_, new_n225_ );
not g0015 ( new_n230_, N390 );
nand g0016 ( new_n231_, N1, N26 );
nand g0017 ( new_n232_, N13, N17 );
nor g0018 ( new_n233_, new_n231_, new_n232_ );
nand g0019 ( N419, new_n230_, new_n233_ );
nand g0020 ( new_n235_, N59, N75 );
not g0021 ( new_n236_, new_n235_ );
nand g0022 ( N420, new_n236_, N80 );
nand g0023 ( new_n238_, N36, N59 );
not g0024 ( new_n239_, new_n238_ );
nand g0025 ( N421, new_n239_, N80 );
nand g0026 ( N422, new_n239_, N42 );
not g0027 ( new_n242_, N90 );
nor g0028 ( new_n243_, N87, N88 );
nor g0029 ( N423, new_n243_, new_n242_ );
nand g0030 ( N446, new_n233_, N390 );
not g0031 ( new_n246_, new_n231_ );
nand g0032 ( new_n247_, new_n246_, N51 );
nand g0033 ( new_n248_, new_n247_, keyIn_0_0 );
not g0034 ( new_n249_, keyIn_0_0 );
not g0035 ( new_n250_, N51 );
nor g0036 ( new_n251_, new_n231_, new_n250_ );
nand g0037 ( new_n252_, new_n251_, new_n249_ );
nand g0038 ( N447, new_n248_, new_n252_ );
not g0039 ( new_n254_, N55 );
nor g0040 ( new_n255_, new_n228_, new_n254_ );
not g0041 ( new_n256_, new_n255_ );
nand g0042 ( new_n257_, N29, N68 );
nor g0043 ( N448, new_n256_, new_n257_ );
nand g0044 ( new_n259_, N59, N68 );
nor g0045 ( new_n260_, new_n256_, new_n259_ );
nand g0046 ( new_n261_, new_n260_, N74 );
nand g0047 ( new_n262_, new_n261_, keyIn_0_10 );
not g0048 ( new_n263_, keyIn_0_10 );
not g0049 ( new_n264_, new_n261_ );
nand g0050 ( new_n265_, new_n264_, new_n263_ );
nand g0051 ( N449, new_n265_, new_n262_ );
not g0052 ( new_n267_, N89 );
nor g0053 ( N450, new_n243_, new_n267_ );
not g0054 ( new_n269_, N111 );
nor g0055 ( new_n270_, new_n269_, N116 );
not g0056 ( new_n271_, N116 );
nor g0057 ( new_n272_, new_n271_, N111 );
nor g0058 ( new_n273_, new_n270_, new_n272_ );
nand g0059 ( new_n274_, N121, N126 );
not g0060 ( new_n275_, new_n274_ );
nor g0061 ( new_n276_, N121, N126 );
nor g0062 ( new_n277_, new_n275_, new_n276_ );
nor g0063 ( new_n278_, new_n273_, new_n277_ );
nand g0064 ( new_n279_, new_n273_, new_n277_ );
not g0065 ( new_n280_, new_n279_ );
nor g0066 ( new_n281_, new_n280_, new_n278_ );
nor g0067 ( new_n282_, new_n281_, N135 );
nand g0068 ( new_n283_, new_n281_, N135 );
not g0069 ( new_n284_, new_n283_ );
nor g0070 ( new_n285_, new_n284_, new_n282_ );
not g0071 ( new_n286_, new_n285_ );
not g0072 ( new_n287_, N130 );
not g0073 ( new_n288_, N101 );
nor g0074 ( new_n289_, new_n288_, N106 );
not g0075 ( new_n290_, N106 );
nor g0076 ( new_n291_, new_n290_, N101 );
nor g0077 ( new_n292_, new_n289_, new_n291_ );
nor g0078 ( new_n293_, N91, N96 );
nand g0079 ( new_n294_, N91, N96 );
nand g0080 ( new_n295_, new_n294_, keyIn_0_15 );
nor g0081 ( new_n296_, new_n295_, new_n293_ );
nor g0082 ( new_n297_, new_n292_, new_n296_ );
nand g0083 ( new_n298_, new_n292_, new_n296_ );
not g0084 ( new_n299_, new_n298_ );
nor g0085 ( new_n300_, new_n299_, new_n297_ );
nor g0086 ( new_n301_, new_n300_, new_n287_ );
nand g0087 ( new_n302_, new_n300_, new_n287_ );
not g0088 ( new_n303_, new_n302_ );
nor g0089 ( new_n304_, new_n303_, new_n301_ );
not g0090 ( new_n305_, new_n304_ );
nand g0091 ( new_n306_, new_n305_, new_n286_ );
nand g0092 ( new_n307_, new_n304_, new_n285_ );
nand g0093 ( N767, new_n306_, new_n307_ );
not g0094 ( new_n309_, N207 );
not g0095 ( new_n310_, N183 );
nor g0096 ( new_n311_, new_n310_, N189 );
not g0097 ( new_n312_, N189 );
nor g0098 ( new_n313_, new_n312_, N183 );
nor g0099 ( new_n314_, new_n311_, new_n313_ );
nand g0100 ( new_n315_, N195, N201 );
not g0101 ( new_n316_, new_n315_ );
nor g0102 ( new_n317_, N195, N201 );
nor g0103 ( new_n318_, new_n316_, new_n317_ );
nor g0104 ( new_n319_, new_n314_, new_n318_ );
nand g0105 ( new_n320_, new_n314_, new_n318_ );
not g0106 ( new_n321_, new_n320_ );
nor g0107 ( new_n322_, new_n321_, new_n319_ );
nor g0108 ( new_n323_, new_n322_, new_n309_ );
nand g0109 ( new_n324_, new_n322_, new_n309_ );
not g0110 ( new_n325_, new_n324_ );
nor g0111 ( new_n326_, new_n325_, new_n323_ );
not g0112 ( new_n327_, new_n326_ );
nand g0113 ( new_n328_, N159, N165 );
not g0114 ( new_n329_, new_n328_ );
nor g0115 ( new_n330_, N159, N165 );
nor g0116 ( new_n331_, new_n329_, new_n330_ );
nand g0117 ( new_n332_, N171, N177 );
not g0118 ( new_n333_, new_n332_ );
nor g0119 ( new_n334_, N171, N177 );
nor g0120 ( new_n335_, new_n333_, new_n334_ );
nor g0121 ( new_n336_, new_n331_, new_n335_ );
nand g0122 ( new_n337_, new_n331_, new_n335_ );
not g0123 ( new_n338_, new_n337_ );
nor g0124 ( new_n339_, new_n338_, new_n336_ );
not g0125 ( new_n340_, new_n339_ );
nand g0126 ( new_n341_, new_n340_, N130 );
not g0127 ( new_n342_, new_n341_ );
nor g0128 ( new_n343_, new_n340_, N130 );
nor g0129 ( new_n344_, new_n342_, new_n343_ );
not g0130 ( new_n345_, new_n344_ );
nand g0131 ( new_n346_, new_n345_, new_n327_ );
nand g0132 ( new_n347_, new_n344_, new_n326_ );
nand g0133 ( N768, new_n346_, new_n347_ );
not g0134 ( new_n349_, N261 );
not g0135 ( new_n350_, keyIn_0_38 );
not g0136 ( new_n351_, keyIn_0_21 );
nand g0137 ( new_n352_, N447, keyIn_0_8 );
not g0138 ( new_n353_, keyIn_0_8 );
nor g0139 ( new_n354_, new_n251_, new_n249_ );
nor g0140 ( new_n355_, new_n247_, keyIn_0_0 );
nor g0141 ( new_n356_, new_n355_, new_n354_ );
nand g0142 ( new_n357_, new_n356_, new_n353_ );
nand g0143 ( new_n358_, new_n357_, new_n352_ );
nand g0144 ( new_n359_, new_n358_, keyIn_0_14 );
not g0145 ( new_n360_, keyIn_0_14 );
nor g0146 ( new_n361_, new_n356_, new_n353_ );
nor g0147 ( new_n362_, N447, keyIn_0_8 );
nor g0148 ( new_n363_, new_n361_, new_n362_ );
nand g0149 ( new_n364_, new_n363_, new_n360_ );
nand g0150 ( new_n365_, new_n364_, new_n359_ );
nand g0151 ( new_n366_, N59, N156 );
nand g0152 ( new_n367_, new_n366_, keyIn_0_5 );
not g0153 ( new_n368_, new_n367_ );
nor g0154 ( new_n369_, new_n366_, keyIn_0_5 );
nor g0155 ( new_n370_, new_n368_, new_n369_ );
nor g0156 ( new_n371_, new_n370_, new_n225_ );
nand g0157 ( new_n372_, new_n365_, new_n371_ );
nor g0158 ( new_n373_, new_n372_, new_n351_ );
not g0159 ( new_n374_, new_n373_ );
nand g0160 ( new_n375_, new_n372_, new_n351_ );
nand g0161 ( new_n376_, new_n375_, N1 );
not g0162 ( new_n377_, new_n376_ );
nand g0163 ( new_n378_, new_n377_, new_n374_ );
nand g0164 ( new_n379_, new_n378_, keyIn_0_25 );
not g0165 ( new_n380_, keyIn_0_25 );
nor g0166 ( new_n381_, new_n376_, new_n373_ );
nand g0167 ( new_n382_, new_n381_, new_n380_ );
nand g0168 ( new_n383_, new_n379_, new_n382_ );
nand g0169 ( new_n384_, new_n383_, N153 );
nand g0170 ( new_n385_, new_n384_, new_n350_ );
not g0171 ( new_n386_, new_n384_ );
nand g0172 ( new_n387_, new_n386_, keyIn_0_38 );
nand g0173 ( new_n388_, new_n387_, new_n385_ );
nand g0174 ( new_n389_, N17, N42 );
nand g0175 ( new_n390_, new_n389_, keyIn_0_7 );
not g0176 ( new_n391_, new_n390_ );
not g0177 ( new_n392_, keyIn_0_6 );
nor g0178 ( new_n393_, N17, N42 );
nor g0179 ( new_n394_, new_n393_, new_n392_ );
nor g0180 ( new_n395_, new_n391_, new_n394_ );
nor g0181 ( new_n396_, new_n389_, keyIn_0_7 );
nand g0182 ( new_n397_, new_n393_, new_n392_ );
not g0183 ( new_n398_, new_n397_ );
nor g0184 ( new_n399_, new_n398_, new_n396_ );
nand g0185 ( new_n400_, new_n399_, new_n395_ );
nor g0186 ( new_n401_, new_n400_, keyIn_0_13 );
not g0187 ( new_n402_, new_n366_ );
nand g0188 ( new_n403_, new_n400_, keyIn_0_13 );
nand g0189 ( new_n404_, new_n403_, new_n402_ );
nor g0190 ( new_n405_, new_n404_, new_n401_ );
nand g0191 ( new_n406_, new_n365_, new_n405_ );
nor g0192 ( new_n407_, new_n406_, keyIn_0_20 );
nand g0193 ( new_n408_, new_n406_, keyIn_0_20 );
not g0194 ( new_n409_, keyIn_0_16 );
not g0195 ( new_n410_, keyIn_0_3 );
nand g0196 ( new_n411_, N42, N59 );
nor g0197 ( new_n412_, new_n411_, new_n215_ );
nor g0198 ( new_n413_, new_n412_, new_n410_ );
not g0199 ( new_n414_, new_n413_ );
nand g0200 ( new_n415_, new_n412_, new_n410_ );
nand g0201 ( new_n416_, new_n414_, new_n415_ );
nand g0202 ( new_n417_, new_n416_, keyIn_0_11 );
nor g0203 ( new_n418_, new_n416_, keyIn_0_11 );
not g0204 ( new_n419_, new_n418_ );
nand g0205 ( new_n420_, new_n419_, new_n417_ );
not g0206 ( new_n421_, keyIn_0_1 );
nand g0207 ( new_n422_, N17, N51 );
nor g0208 ( new_n423_, new_n226_, new_n422_ );
nor g0209 ( new_n424_, new_n423_, new_n421_ );
not g0210 ( new_n425_, new_n424_ );
nand g0211 ( new_n426_, new_n423_, new_n421_ );
nand g0212 ( new_n427_, new_n425_, new_n426_ );
nand g0213 ( new_n428_, new_n427_, keyIn_0_9 );
not g0214 ( new_n429_, keyIn_0_9 );
not g0215 ( new_n430_, new_n426_ );
nor g0216 ( new_n431_, new_n430_, new_n424_ );
nand g0217 ( new_n432_, new_n431_, new_n429_ );
nand g0218 ( new_n433_, new_n432_, new_n428_ );
not g0219 ( new_n434_, new_n433_ );
nand g0220 ( new_n435_, new_n434_, new_n420_ );
nand g0221 ( new_n436_, new_n435_, new_n409_ );
not g0222 ( new_n437_, new_n417_ );
nor g0223 ( new_n438_, new_n437_, new_n418_ );
nor g0224 ( new_n439_, new_n438_, new_n433_ );
nand g0225 ( new_n440_, new_n439_, keyIn_0_16 );
nand g0226 ( new_n441_, new_n440_, new_n436_ );
nand g0227 ( new_n442_, new_n408_, new_n441_ );
nor g0228 ( new_n443_, new_n442_, new_n407_ );
nor g0229 ( new_n444_, new_n443_, keyIn_0_22 );
not g0230 ( new_n445_, keyIn_0_22 );
not g0231 ( new_n446_, new_n407_ );
not g0232 ( new_n447_, new_n442_ );
nand g0233 ( new_n448_, new_n447_, new_n446_ );
nor g0234 ( new_n449_, new_n448_, new_n445_ );
nor g0235 ( new_n450_, new_n449_, new_n444_ );
nand g0236 ( new_n451_, new_n450_, N126 );
nand g0237 ( new_n452_, new_n451_, keyIn_0_39 );
not g0238 ( new_n453_, keyIn_0_39 );
not g0239 ( new_n454_, N126 );
nand g0240 ( new_n455_, new_n448_, new_n445_ );
nand g0241 ( new_n456_, new_n443_, keyIn_0_22 );
nand g0242 ( new_n457_, new_n455_, new_n456_ );
nor g0243 ( new_n458_, new_n457_, new_n454_ );
nand g0244 ( new_n459_, new_n458_, new_n453_ );
nand g0245 ( new_n460_, new_n452_, new_n459_ );
nand g0246 ( new_n461_, new_n388_, new_n460_ );
nand g0247 ( new_n462_, new_n461_, keyIn_0_45 );
not g0248 ( new_n463_, keyIn_0_45 );
not g0249 ( new_n464_, new_n385_ );
nor g0250 ( new_n465_, new_n384_, new_n350_ );
nor g0251 ( new_n466_, new_n464_, new_n465_ );
nor g0252 ( new_n467_, new_n458_, new_n453_ );
nor g0253 ( new_n468_, new_n451_, keyIn_0_39 );
nor g0254 ( new_n469_, new_n468_, new_n467_ );
nor g0255 ( new_n470_, new_n466_, new_n469_ );
nand g0256 ( new_n471_, new_n470_, new_n463_ );
nand g0257 ( new_n472_, new_n471_, new_n462_ );
not g0258 ( new_n473_, keyIn_0_19 );
not g0259 ( new_n474_, new_n365_ );
nand g0260 ( new_n475_, N29, N75 );
nor g0261 ( new_n476_, new_n475_, new_n218_ );
nor g0262 ( new_n477_, new_n476_, keyIn_0_2 );
nand g0263 ( new_n478_, new_n476_, keyIn_0_2 );
not g0264 ( new_n479_, new_n478_ );
nor g0265 ( new_n480_, new_n479_, new_n477_ );
nor g0266 ( new_n481_, new_n474_, new_n480_ );
not g0267 ( new_n482_, new_n481_ );
nor g0268 ( new_n483_, new_n482_, new_n254_ );
nor g0269 ( new_n484_, new_n483_, new_n473_ );
nand g0270 ( new_n485_, new_n483_, new_n473_ );
not g0271 ( new_n486_, new_n485_ );
nor g0272 ( new_n487_, new_n486_, new_n484_ );
not g0273 ( new_n488_, keyIn_0_4 );
nor g0274 ( new_n489_, new_n488_, N268 );
nand g0275 ( new_n490_, new_n488_, N268 );
not g0276 ( new_n491_, new_n490_ );
nor g0277 ( new_n492_, new_n491_, new_n489_ );
not g0278 ( new_n493_, new_n492_ );
nand g0279 ( new_n494_, new_n493_, keyIn_0_12 );
not g0280 ( new_n495_, new_n494_ );
nor g0281 ( new_n496_, new_n493_, keyIn_0_12 );
nor g0282 ( new_n497_, new_n495_, new_n496_ );
nor g0283 ( new_n498_, new_n487_, new_n497_ );
not g0284 ( new_n499_, new_n498_ );
nand g0285 ( new_n500_, new_n499_, keyIn_0_29 );
not g0286 ( new_n501_, new_n500_ );
nor g0287 ( new_n502_, new_n499_, keyIn_0_29 );
nor g0288 ( new_n503_, new_n501_, new_n502_ );
not g0289 ( new_n504_, new_n503_ );
nand g0290 ( new_n505_, new_n472_, new_n504_ );
nand g0291 ( new_n506_, new_n505_, keyIn_0_50 );
not g0292 ( new_n507_, keyIn_0_50 );
not g0293 ( new_n508_, new_n462_ );
nor g0294 ( new_n509_, new_n461_, keyIn_0_45 );
nor g0295 ( new_n510_, new_n508_, new_n509_ );
nor g0296 ( new_n511_, new_n510_, new_n503_ );
nand g0297 ( new_n512_, new_n511_, new_n507_ );
nand g0298 ( new_n513_, new_n512_, new_n506_ );
nand g0299 ( new_n514_, new_n513_, N201 );
nand g0300 ( new_n515_, new_n514_, keyIn_0_60 );
not g0301 ( new_n516_, keyIn_0_60 );
not g0302 ( new_n517_, new_n514_ );
nand g0303 ( new_n518_, new_n517_, new_n516_ );
nand g0304 ( new_n519_, new_n518_, new_n515_ );
not g0305 ( new_n520_, N201 );
not g0306 ( new_n521_, new_n506_ );
nor g0307 ( new_n522_, new_n505_, keyIn_0_50 );
nor g0308 ( new_n523_, new_n521_, new_n522_ );
nand g0309 ( new_n524_, new_n523_, new_n520_ );
nand g0310 ( new_n525_, new_n524_, keyIn_0_61 );
not g0311 ( new_n526_, keyIn_0_61 );
nor g0312 ( new_n527_, new_n513_, N201 );
nand g0313 ( new_n528_, new_n527_, new_n526_ );
nand g0314 ( new_n529_, new_n525_, new_n528_ );
nand g0315 ( new_n530_, new_n519_, new_n529_ );
nand g0316 ( new_n531_, new_n530_, new_n349_ );
not g0317 ( new_n532_, N219 );
nor g0318 ( new_n533_, new_n530_, new_n349_ );
nor g0319 ( new_n534_, new_n533_, new_n532_ );
nand g0320 ( new_n535_, new_n534_, new_n531_ );
not g0321 ( new_n536_, keyIn_0_67 );
nand g0322 ( new_n537_, new_n519_, new_n536_ );
not g0323 ( new_n538_, new_n515_ );
nor g0324 ( new_n539_, new_n514_, keyIn_0_60 );
nor g0325 ( new_n540_, new_n538_, new_n539_ );
nand g0326 ( new_n541_, new_n540_, keyIn_0_67 );
nand g0327 ( new_n542_, new_n541_, new_n537_ );
nand g0328 ( new_n543_, new_n542_, N237 );
not g0329 ( new_n544_, N228 );
nor g0330 ( new_n545_, new_n530_, new_n544_ );
nand g0331 ( new_n546_, new_n513_, N246 );
not g0332 ( new_n547_, N73 );
nand g0333 ( new_n548_, N42, N72 );
nor g0334 ( new_n549_, new_n548_, new_n547_ );
nand g0335 ( new_n550_, new_n260_, new_n549_ );
nor g0336 ( new_n551_, new_n550_, new_n520_ );
nand g0337 ( new_n552_, N255, N267 );
nand g0338 ( new_n553_, N121, N210 );
nand g0339 ( new_n554_, new_n552_, new_n553_ );
nor g0340 ( new_n555_, new_n551_, new_n554_ );
nand g0341 ( new_n556_, new_n546_, new_n555_ );
nor g0342 ( new_n557_, new_n545_, new_n556_ );
nand g0343 ( new_n558_, new_n557_, new_n543_ );
not g0344 ( new_n559_, new_n558_ );
nand g0345 ( N850, new_n559_, new_n535_ );
not g0346 ( new_n561_, keyIn_0_112 );
not g0347 ( new_n562_, keyIn_0_106 );
not g0348 ( new_n563_, keyIn_0_100 );
not g0349 ( new_n564_, keyIn_0_92 );
not g0350 ( new_n565_, keyIn_0_83 );
not g0351 ( new_n566_, keyIn_0_76 );
not g0352 ( new_n567_, keyIn_0_32 );
not g0353 ( new_n568_, N143 );
nor g0354 ( new_n569_, new_n381_, new_n380_ );
not g0355 ( new_n570_, new_n382_ );
nor g0356 ( new_n571_, new_n570_, new_n569_ );
nor g0357 ( new_n572_, new_n571_, new_n568_ );
not g0358 ( new_n573_, new_n572_ );
nor g0359 ( new_n574_, new_n573_, new_n567_ );
not g0360 ( new_n575_, keyIn_0_33 );
nor g0361 ( new_n576_, new_n457_, new_n269_ );
nor g0362 ( new_n577_, new_n576_, new_n575_ );
nor g0363 ( new_n578_, new_n574_, new_n577_ );
not g0364 ( new_n579_, new_n578_ );
nand g0365 ( new_n580_, new_n576_, new_n575_ );
nand g0366 ( new_n581_, new_n573_, new_n567_ );
nand g0367 ( new_n582_, new_n581_, new_n580_ );
nor g0368 ( new_n583_, new_n579_, new_n582_ );
not g0369 ( new_n584_, new_n583_ );
nand g0370 ( new_n585_, new_n584_, keyIn_0_42 );
not g0371 ( new_n586_, keyIn_0_42 );
nand g0372 ( new_n587_, new_n583_, new_n586_ );
nand g0373 ( new_n588_, new_n585_, new_n587_ );
not g0374 ( new_n589_, keyIn_0_26 );
nand g0375 ( new_n590_, new_n499_, new_n589_ );
nand g0376 ( new_n591_, new_n498_, keyIn_0_26 );
nand g0377 ( new_n592_, new_n590_, new_n591_ );
nand g0378 ( new_n593_, new_n588_, new_n592_ );
nand g0379 ( new_n594_, new_n593_, keyIn_0_47 );
not g0380 ( new_n595_, new_n594_ );
nor g0381 ( new_n596_, new_n593_, keyIn_0_47 );
nor g0382 ( new_n597_, new_n595_, new_n596_ );
not g0383 ( new_n598_, new_n597_ );
nor g0384 ( new_n599_, new_n598_, new_n310_ );
not g0385 ( new_n600_, new_n599_ );
nor g0386 ( new_n601_, new_n600_, keyIn_0_54 );
nand g0387 ( new_n602_, new_n600_, keyIn_0_54 );
not g0388 ( new_n603_, new_n602_ );
nor g0389 ( new_n604_, new_n603_, new_n601_ );
not g0390 ( new_n605_, keyIn_0_55 );
nor g0391 ( new_n606_, new_n597_, N183 );
nor g0392 ( new_n607_, new_n606_, new_n605_ );
nand g0393 ( new_n608_, new_n606_, new_n605_ );
not g0394 ( new_n609_, new_n608_ );
nor g0395 ( new_n610_, new_n609_, new_n607_ );
not g0396 ( new_n611_, new_n610_ );
nor g0397 ( new_n612_, new_n604_, new_n611_ );
not g0398 ( new_n613_, new_n612_ );
not g0399 ( new_n614_, keyIn_0_75 );
nand g0400 ( new_n615_, new_n383_, N146 );
nand g0401 ( new_n616_, new_n615_, keyIn_0_34 );
not g0402 ( new_n617_, new_n616_ );
not g0403 ( new_n618_, keyIn_0_35 );
nor g0404 ( new_n619_, new_n457_, new_n271_ );
nor g0405 ( new_n620_, new_n619_, new_n618_ );
nor g0406 ( new_n621_, new_n617_, new_n620_ );
nand g0407 ( new_n622_, new_n450_, N116 );
nor g0408 ( new_n623_, new_n622_, keyIn_0_35 );
nor g0409 ( new_n624_, new_n615_, keyIn_0_34 );
nor g0410 ( new_n625_, new_n623_, new_n624_ );
nand g0411 ( new_n626_, new_n621_, new_n625_ );
nor g0412 ( new_n627_, new_n626_, keyIn_0_43 );
not g0413 ( new_n628_, new_n627_ );
nand g0414 ( new_n629_, new_n499_, keyIn_0_27 );
not g0415 ( new_n630_, new_n629_ );
nor g0416 ( new_n631_, new_n499_, keyIn_0_27 );
nor g0417 ( new_n632_, new_n630_, new_n631_ );
not g0418 ( new_n633_, keyIn_0_43 );
nand g0419 ( new_n634_, new_n622_, keyIn_0_35 );
nand g0420 ( new_n635_, new_n634_, new_n616_ );
nand g0421 ( new_n636_, new_n619_, new_n618_ );
not g0422 ( new_n637_, keyIn_0_34 );
not g0423 ( new_n638_, new_n615_ );
nand g0424 ( new_n639_, new_n638_, new_n637_ );
nand g0425 ( new_n640_, new_n639_, new_n636_ );
nor g0426 ( new_n641_, new_n640_, new_n635_ );
nor g0427 ( new_n642_, new_n641_, new_n633_ );
nor g0428 ( new_n643_, new_n642_, new_n632_ );
nand g0429 ( new_n644_, new_n643_, new_n628_ );
nand g0430 ( new_n645_, new_n644_, keyIn_0_48 );
not g0431 ( new_n646_, keyIn_0_48 );
not g0432 ( new_n647_, new_n632_ );
nand g0433 ( new_n648_, new_n626_, keyIn_0_43 );
nand g0434 ( new_n649_, new_n648_, new_n647_ );
nor g0435 ( new_n650_, new_n649_, new_n627_ );
nand g0436 ( new_n651_, new_n650_, new_n646_ );
nand g0437 ( new_n652_, new_n645_, new_n651_ );
not g0438 ( new_n653_, new_n652_ );
nand g0439 ( new_n654_, new_n653_, new_n312_ );
nand g0440 ( new_n655_, new_n654_, keyIn_0_57 );
not g0441 ( new_n656_, keyIn_0_57 );
nor g0442 ( new_n657_, new_n652_, N189 );
nand g0443 ( new_n658_, new_n657_, new_n656_ );
nand g0444 ( new_n659_, new_n655_, new_n658_ );
not g0445 ( new_n660_, keyIn_0_66 );
not g0446 ( new_n661_, N195 );
not g0447 ( new_n662_, keyIn_0_49 );
not g0448 ( new_n663_, keyIn_0_44 );
nand g0449 ( new_n664_, new_n383_, N149 );
nand g0450 ( new_n665_, new_n664_, keyIn_0_36 );
not g0451 ( new_n666_, keyIn_0_36 );
not g0452 ( new_n667_, new_n664_ );
nand g0453 ( new_n668_, new_n667_, new_n666_ );
nand g0454 ( new_n669_, new_n668_, new_n665_ );
nand g0455 ( new_n670_, new_n450_, N121 );
nand g0456 ( new_n671_, new_n670_, keyIn_0_37 );
not g0457 ( new_n672_, keyIn_0_37 );
not g0458 ( new_n673_, N121 );
nor g0459 ( new_n674_, new_n457_, new_n673_ );
nand g0460 ( new_n675_, new_n674_, new_n672_ );
nand g0461 ( new_n676_, new_n671_, new_n675_ );
nand g0462 ( new_n677_, new_n669_, new_n676_ );
nor g0463 ( new_n678_, new_n677_, new_n663_ );
not g0464 ( new_n679_, new_n678_ );
not g0465 ( new_n680_, keyIn_0_28 );
nand g0466 ( new_n681_, new_n499_, new_n680_ );
nand g0467 ( new_n682_, new_n498_, keyIn_0_28 );
nand g0468 ( new_n683_, new_n681_, new_n682_ );
nand g0469 ( new_n684_, new_n677_, new_n663_ );
nand g0470 ( new_n685_, new_n684_, new_n683_ );
not g0471 ( new_n686_, new_n685_ );
nand g0472 ( new_n687_, new_n686_, new_n679_ );
nand g0473 ( new_n688_, new_n687_, new_n662_ );
nor g0474 ( new_n689_, new_n685_, new_n678_ );
nand g0475 ( new_n690_, new_n689_, keyIn_0_49 );
nand g0476 ( new_n691_, new_n688_, new_n690_ );
nor g0477 ( new_n692_, new_n691_, new_n661_ );
nor g0478 ( new_n693_, new_n692_, keyIn_0_58 );
nand g0479 ( new_n694_, new_n692_, keyIn_0_58 );
not g0480 ( new_n695_, new_n694_ );
nor g0481 ( new_n696_, new_n695_, new_n693_ );
not g0482 ( new_n697_, new_n696_ );
nand g0483 ( new_n698_, new_n697_, new_n660_ );
nand g0484 ( new_n699_, new_n696_, keyIn_0_66 );
nand g0485 ( new_n700_, new_n698_, new_n699_ );
nand g0486 ( new_n701_, new_n700_, new_n659_ );
nand g0487 ( new_n702_, new_n701_, keyIn_0_72 );
nor g0488 ( new_n703_, new_n701_, keyIn_0_72 );
not g0489 ( new_n704_, new_n703_ );
nand g0490 ( new_n705_, new_n704_, new_n702_ );
not g0491 ( new_n706_, keyIn_0_71 );
not g0492 ( new_n707_, keyIn_0_65 );
not g0493 ( new_n708_, keyIn_0_56 );
nand g0494 ( new_n709_, new_n652_, N189 );
nand g0495 ( new_n710_, new_n709_, new_n708_ );
not g0496 ( new_n711_, new_n709_ );
nand g0497 ( new_n712_, new_n711_, keyIn_0_56 );
nand g0498 ( new_n713_, new_n712_, new_n710_ );
nand g0499 ( new_n714_, new_n713_, new_n707_ );
not g0500 ( new_n715_, new_n710_ );
nor g0501 ( new_n716_, new_n709_, new_n708_ );
nor g0502 ( new_n717_, new_n715_, new_n716_ );
nand g0503 ( new_n718_, new_n717_, keyIn_0_65 );
nand g0504 ( new_n719_, new_n718_, new_n714_ );
nand g0505 ( new_n720_, new_n719_, new_n706_ );
not g0506 ( new_n721_, new_n720_ );
not g0507 ( new_n722_, keyIn_0_68 );
nand g0508 ( new_n723_, new_n529_, N261 );
not g0509 ( new_n724_, keyIn_0_59 );
nand g0510 ( new_n725_, new_n691_, new_n661_ );
nand g0511 ( new_n726_, new_n725_, new_n724_ );
not g0512 ( new_n727_, new_n726_ );
nor g0513 ( new_n728_, new_n725_, new_n724_ );
nor g0514 ( new_n729_, new_n727_, new_n728_ );
nand g0515 ( new_n730_, new_n729_, new_n659_ );
nor g0516 ( new_n731_, new_n730_, new_n723_ );
nor g0517 ( new_n732_, new_n731_, new_n722_ );
nor g0518 ( new_n733_, new_n721_, new_n732_ );
nor g0519 ( new_n734_, new_n719_, new_n706_ );
not g0520 ( new_n735_, new_n723_ );
nor g0521 ( new_n736_, new_n657_, new_n656_ );
not g0522 ( new_n737_, new_n658_ );
nor g0523 ( new_n738_, new_n737_, new_n736_ );
not g0524 ( new_n739_, new_n728_ );
nand g0525 ( new_n740_, new_n739_, new_n726_ );
nor g0526 ( new_n741_, new_n738_, new_n740_ );
nand g0527 ( new_n742_, new_n735_, new_n741_ );
nor g0528 ( new_n743_, new_n742_, keyIn_0_68 );
nor g0529 ( new_n744_, new_n743_, new_n734_ );
nand g0530 ( new_n745_, new_n744_, new_n733_ );
not g0531 ( new_n746_, keyIn_0_73 );
nand g0532 ( new_n747_, new_n542_, new_n741_ );
nand g0533 ( new_n748_, new_n747_, new_n746_ );
not g0534 ( new_n749_, new_n747_ );
nand g0535 ( new_n750_, new_n749_, keyIn_0_73 );
nand g0536 ( new_n751_, new_n750_, new_n748_ );
nor g0537 ( new_n752_, new_n751_, new_n745_ );
nand g0538 ( new_n753_, new_n752_, new_n705_ );
nand g0539 ( new_n754_, new_n753_, new_n614_ );
not g0540 ( new_n755_, new_n702_ );
nor g0541 ( new_n756_, new_n755_, new_n703_ );
nand g0542 ( new_n757_, new_n742_, keyIn_0_68 );
nand g0543 ( new_n758_, new_n757_, new_n720_ );
nor g0544 ( new_n759_, new_n717_, keyIn_0_65 );
nor g0545 ( new_n760_, new_n713_, new_n707_ );
nor g0546 ( new_n761_, new_n759_, new_n760_ );
nand g0547 ( new_n762_, new_n761_, keyIn_0_71 );
nand g0548 ( new_n763_, new_n731_, new_n722_ );
nand g0549 ( new_n764_, new_n762_, new_n763_ );
nor g0550 ( new_n765_, new_n758_, new_n764_ );
not g0551 ( new_n766_, new_n748_ );
nor g0552 ( new_n767_, new_n747_, new_n746_ );
nor g0553 ( new_n768_, new_n766_, new_n767_ );
nand g0554 ( new_n769_, new_n768_, new_n765_ );
nor g0555 ( new_n770_, new_n769_, new_n756_ );
nand g0556 ( new_n771_, new_n770_, keyIn_0_75 );
nand g0557 ( new_n772_, new_n771_, new_n754_ );
nand g0558 ( new_n773_, new_n772_, new_n613_ );
nor g0559 ( new_n774_, new_n773_, new_n566_ );
nor g0560 ( new_n775_, new_n772_, new_n613_ );
nor g0561 ( new_n776_, new_n775_, keyIn_0_77 );
nor g0562 ( new_n777_, new_n776_, new_n774_ );
not g0563 ( new_n778_, new_n777_ );
nand g0564 ( new_n779_, new_n775_, keyIn_0_77 );
nand g0565 ( new_n780_, new_n773_, new_n566_ );
nand g0566 ( new_n781_, new_n779_, new_n780_ );
nor g0567 ( new_n782_, new_n778_, new_n781_ );
not g0568 ( new_n783_, new_n782_ );
nor g0569 ( new_n784_, new_n783_, keyIn_0_80 );
nand g0570 ( new_n785_, new_n783_, keyIn_0_80 );
nand g0571 ( new_n786_, new_n785_, N219 );
nor g0572 ( new_n787_, new_n786_, new_n784_ );
nor g0573 ( new_n788_, new_n787_, new_n565_ );
nand g0574 ( new_n789_, new_n787_, new_n565_ );
not g0575 ( new_n790_, new_n789_ );
nor g0576 ( new_n791_, new_n790_, new_n788_ );
nand g0577 ( new_n792_, N106, N210 );
not g0578 ( new_n793_, new_n792_ );
nor g0579 ( new_n794_, new_n791_, new_n793_ );
not g0580 ( new_n795_, new_n794_ );
nand g0581 ( new_n796_, new_n795_, new_n564_ );
not g0582 ( new_n797_, new_n796_ );
nor g0583 ( new_n798_, new_n795_, new_n564_ );
nor g0584 ( new_n799_, new_n797_, new_n798_ );
not g0585 ( new_n800_, N237 );
not g0586 ( new_n801_, new_n604_ );
nand g0587 ( new_n802_, new_n801_, keyIn_0_64 );
not g0588 ( new_n803_, new_n802_ );
nor g0589 ( new_n804_, new_n801_, keyIn_0_64 );
nor g0590 ( new_n805_, new_n803_, new_n804_ );
nor g0591 ( new_n806_, new_n805_, new_n800_ );
nor g0592 ( new_n807_, new_n613_, new_n544_ );
not g0593 ( new_n808_, N246 );
nor g0594 ( new_n809_, new_n598_, new_n808_ );
nor g0595 ( new_n810_, new_n550_, new_n310_ );
nor g0596 ( new_n811_, new_n809_, new_n810_ );
not g0597 ( new_n812_, new_n811_ );
nor g0598 ( new_n813_, new_n807_, new_n812_ );
not g0599 ( new_n814_, new_n813_ );
nor g0600 ( new_n815_, new_n814_, new_n806_ );
not g0601 ( new_n816_, new_n815_ );
nor g0602 ( new_n817_, new_n799_, new_n816_ );
nor g0603 ( new_n818_, new_n817_, new_n563_ );
nand g0604 ( new_n819_, new_n817_, new_n563_ );
not g0605 ( new_n820_, new_n819_ );
nor g0606 ( new_n821_, new_n820_, new_n818_ );
nor g0607 ( new_n822_, new_n821_, new_n562_ );
nand g0608 ( new_n823_, new_n821_, new_n562_ );
not g0609 ( new_n824_, new_n823_ );
nor g0610 ( new_n825_, new_n824_, new_n822_ );
not g0611 ( new_n826_, new_n825_ );
nand g0612 ( new_n827_, new_n826_, new_n561_ );
nand g0613 ( new_n828_, new_n825_, keyIn_0_112 );
nand g0614 ( N863, new_n827_, new_n828_ );
nor g0615 ( new_n830_, new_n738_, new_n717_ );
not g0616 ( new_n831_, new_n830_ );
nor g0617 ( new_n832_, new_n542_, new_n735_ );
nor g0618 ( new_n833_, new_n832_, new_n740_ );
nor g0619 ( new_n834_, new_n833_, new_n700_ );
nand g0620 ( new_n835_, new_n834_, new_n831_ );
nor g0621 ( new_n836_, new_n834_, new_n831_ );
nor g0622 ( new_n837_, new_n836_, new_n532_ );
nand g0623 ( new_n838_, new_n837_, new_n835_ );
nor g0624 ( new_n839_, new_n761_, new_n800_ );
nand g0625 ( new_n840_, new_n830_, N228 );
nand g0626 ( new_n841_, new_n652_, N246 );
nor g0627 ( new_n842_, new_n550_, new_n312_ );
nand g0628 ( new_n843_, N255, N259 );
nand g0629 ( new_n844_, N111, N210 );
nand g0630 ( new_n845_, new_n843_, new_n844_ );
nor g0631 ( new_n846_, new_n842_, new_n845_ );
nand g0632 ( new_n847_, new_n841_, new_n846_ );
not g0633 ( new_n848_, new_n847_ );
nand g0634 ( new_n849_, new_n840_, new_n848_ );
nor g0635 ( new_n850_, new_n839_, new_n849_ );
nand g0636 ( N864, new_n838_, new_n850_ );
not g0637 ( new_n852_, new_n832_ );
nor g0638 ( new_n853_, new_n697_, new_n740_ );
nor g0639 ( new_n854_, new_n852_, new_n853_ );
nand g0640 ( new_n855_, new_n852_, new_n853_ );
nand g0641 ( new_n856_, new_n855_, N219 );
nor g0642 ( new_n857_, new_n856_, new_n854_ );
not g0643 ( new_n858_, new_n857_ );
nand g0644 ( new_n859_, new_n858_, keyIn_0_84 );
not g0645 ( new_n860_, keyIn_0_84 );
nand g0646 ( new_n861_, new_n857_, new_n860_ );
nand g0647 ( new_n862_, new_n859_, new_n861_ );
not g0648 ( new_n863_, new_n700_ );
nor g0649 ( new_n864_, new_n863_, new_n800_ );
nand g0650 ( new_n865_, new_n853_, N228 );
nor g0651 ( new_n866_, new_n691_, new_n808_ );
not g0652 ( new_n867_, new_n550_ );
nand g0653 ( new_n868_, new_n867_, N195 );
nand g0654 ( new_n869_, N255, N260 );
nand g0655 ( new_n870_, N116, N210 );
nand g0656 ( new_n871_, new_n869_, new_n870_ );
not g0657 ( new_n872_, new_n871_ );
nand g0658 ( new_n873_, new_n868_, new_n872_ );
nor g0659 ( new_n874_, new_n866_, new_n873_ );
nand g0660 ( new_n875_, new_n865_, new_n874_ );
nor g0661 ( new_n876_, new_n864_, new_n875_ );
nand g0662 ( N865, new_n862_, new_n876_ );
not g0663 ( new_n878_, keyIn_0_113 );
not g0664 ( new_n879_, keyIn_0_107 );
not g0665 ( new_n880_, keyIn_0_40 );
nand g0666 ( new_n881_, new_n450_, N91 );
nand g0667 ( new_n882_, N8, N138 );
nand g0668 ( new_n883_, new_n881_, new_n882_ );
nor g0669 ( new_n884_, new_n883_, new_n880_ );
nand g0670 ( new_n885_, new_n883_, new_n880_ );
not g0671 ( new_n886_, keyIn_0_18 );
nor g0672 ( new_n887_, new_n482_, new_n225_ );
not g0673 ( new_n888_, new_n887_ );
nor g0674 ( new_n889_, new_n888_, new_n886_ );
nor g0675 ( new_n890_, new_n887_, keyIn_0_18 );
nor g0676 ( new_n891_, new_n890_, new_n492_ );
not g0677 ( new_n892_, new_n891_ );
nor g0678 ( new_n893_, new_n892_, new_n889_ );
not g0679 ( new_n894_, keyIn_0_17 );
nor g0680 ( new_n895_, new_n370_, new_n254_ );
nand g0681 ( new_n896_, new_n365_, new_n895_ );
nand g0682 ( new_n897_, new_n896_, new_n894_ );
not g0683 ( new_n898_, new_n897_ );
nor g0684 ( new_n899_, new_n896_, new_n894_ );
nor g0685 ( new_n900_, new_n898_, new_n899_ );
nor g0686 ( new_n901_, new_n900_, new_n568_ );
nor g0687 ( new_n902_, new_n893_, new_n901_ );
nand g0688 ( new_n903_, new_n885_, new_n902_ );
nor g0689 ( new_n904_, new_n903_, new_n884_ );
not g0690 ( new_n905_, new_n904_ );
nor g0691 ( new_n906_, new_n905_, N159 );
nand g0692 ( new_n907_, new_n450_, N96 );
not g0693 ( new_n908_, new_n907_ );
not g0694 ( new_n909_, new_n893_ );
nand g0695 ( new_n910_, N51, N138 );
not g0696 ( new_n911_, new_n910_ );
not g0697 ( new_n912_, N146 );
nor g0698 ( new_n913_, new_n900_, new_n912_ );
nor g0699 ( new_n914_, new_n913_, new_n911_ );
nand g0700 ( new_n915_, new_n909_, new_n914_ );
nor g0701 ( new_n916_, new_n915_, new_n908_ );
not g0702 ( new_n917_, new_n916_ );
nor g0703 ( new_n918_, new_n917_, N165 );
nor g0704 ( new_n919_, new_n457_, new_n288_ );
nand g0705 ( new_n920_, N17, N138 );
not g0706 ( new_n921_, new_n920_ );
not g0707 ( new_n922_, N149 );
nor g0708 ( new_n923_, new_n900_, new_n922_ );
nor g0709 ( new_n924_, new_n923_, new_n921_ );
nand g0710 ( new_n925_, new_n909_, new_n924_ );
nor g0711 ( new_n926_, new_n925_, new_n919_ );
not g0712 ( new_n927_, new_n926_ );
nor g0713 ( new_n928_, new_n927_, N171 );
nor g0714 ( new_n929_, new_n918_, new_n928_ );
not g0715 ( new_n930_, keyIn_0_79 );
not g0716 ( new_n931_, keyIn_0_78 );
nor g0717 ( new_n932_, new_n770_, keyIn_0_75 );
nor g0718 ( new_n933_, new_n753_, new_n614_ );
nor g0719 ( new_n934_, new_n932_, new_n933_ );
nand g0720 ( new_n935_, new_n934_, new_n610_ );
nand g0721 ( new_n936_, new_n935_, new_n931_ );
nor g0722 ( new_n937_, new_n772_, new_n611_ );
nand g0723 ( new_n938_, new_n937_, keyIn_0_78 );
nand g0724 ( new_n939_, new_n936_, new_n938_ );
not g0725 ( new_n940_, keyIn_0_70 );
nor g0726 ( new_n941_, new_n805_, new_n940_ );
not g0727 ( new_n942_, new_n941_ );
nand g0728 ( new_n943_, new_n805_, new_n940_ );
nand g0729 ( new_n944_, new_n942_, new_n943_ );
nand g0730 ( new_n945_, new_n939_, new_n944_ );
nand g0731 ( new_n946_, new_n945_, new_n930_ );
nor g0732 ( new_n947_, new_n945_, new_n930_ );
not g0733 ( new_n948_, new_n947_ );
nand g0734 ( new_n949_, new_n948_, new_n946_ );
not g0735 ( new_n950_, keyIn_0_41 );
not g0736 ( new_n951_, keyIn_0_30 );
nor g0737 ( new_n952_, new_n457_, new_n290_ );
not g0738 ( new_n953_, new_n952_ );
nor g0739 ( new_n954_, new_n953_, new_n951_ );
nand g0740 ( new_n955_, N138, N152 );
not g0741 ( new_n956_, new_n955_ );
nor g0742 ( new_n957_, new_n952_, keyIn_0_30 );
nor g0743 ( new_n958_, new_n957_, new_n956_ );
not g0744 ( new_n959_, new_n958_ );
nor g0745 ( new_n960_, new_n959_, new_n954_ );
not g0746 ( new_n961_, new_n960_ );
nand g0747 ( new_n962_, new_n961_, new_n950_ );
nand g0748 ( new_n963_, new_n960_, keyIn_0_41 );
nand g0749 ( new_n964_, new_n962_, new_n963_ );
not g0750 ( new_n965_, keyIn_0_31 );
nor g0751 ( new_n966_, new_n893_, keyIn_0_24 );
nand g0752 ( new_n967_, new_n893_, keyIn_0_24 );
not g0753 ( new_n968_, new_n967_ );
not g0754 ( new_n969_, keyIn_0_23 );
not g0755 ( new_n970_, N153 );
nor g0756 ( new_n971_, new_n900_, new_n970_ );
nor g0757 ( new_n972_, new_n971_, new_n969_ );
nand g0758 ( new_n973_, new_n971_, new_n969_ );
not g0759 ( new_n974_, new_n973_ );
nor g0760 ( new_n975_, new_n974_, new_n972_ );
nor g0761 ( new_n976_, new_n968_, new_n975_ );
not g0762 ( new_n977_, new_n976_ );
nor g0763 ( new_n978_, new_n977_, new_n966_ );
not g0764 ( new_n979_, new_n978_ );
nand g0765 ( new_n980_, new_n979_, new_n965_ );
nand g0766 ( new_n981_, new_n978_, keyIn_0_31 );
nand g0767 ( new_n982_, new_n980_, new_n981_ );
nand g0768 ( new_n983_, new_n982_, new_n964_ );
nand g0769 ( new_n984_, new_n983_, keyIn_0_46 );
not g0770 ( new_n985_, new_n984_ );
nor g0771 ( new_n986_, new_n983_, keyIn_0_46 );
nor g0772 ( new_n987_, new_n985_, new_n986_ );
not g0773 ( new_n988_, new_n987_ );
nor g0774 ( new_n989_, new_n988_, N177 );
not g0775 ( new_n990_, new_n989_ );
nor g0776 ( new_n991_, new_n990_, keyIn_0_53 );
nand g0777 ( new_n992_, new_n990_, keyIn_0_53 );
not g0778 ( new_n993_, new_n992_ );
nor g0779 ( new_n994_, new_n993_, new_n991_ );
not g0780 ( new_n995_, new_n994_ );
nor g0781 ( new_n996_, new_n949_, new_n995_ );
nand g0782 ( new_n997_, new_n996_, new_n929_ );
nand g0783 ( new_n998_, new_n997_, keyIn_0_87 );
not g0784 ( new_n999_, new_n946_ );
nor g0785 ( new_n1000_, new_n999_, new_n947_ );
nand g0786 ( new_n1001_, new_n1000_, new_n994_ );
not g0787 ( new_n1002_, new_n929_ );
nor g0788 ( new_n1003_, new_n1002_, keyIn_0_87 );
not g0789 ( new_n1004_, new_n1003_ );
nor g0790 ( new_n1005_, new_n1001_, new_n1004_ );
not g0791 ( new_n1006_, keyIn_0_74 );
not g0792 ( new_n1007_, keyIn_0_63 );
not g0793 ( new_n1008_, keyIn_0_52 );
nand g0794 ( new_n1009_, new_n988_, N177 );
not g0795 ( new_n1010_, new_n1009_ );
nor g0796 ( new_n1011_, new_n1010_, new_n1008_ );
nor g0797 ( new_n1012_, new_n1009_, keyIn_0_52 );
nor g0798 ( new_n1013_, new_n1011_, new_n1012_ );
nor g0799 ( new_n1014_, new_n1013_, new_n1007_ );
not g0800 ( new_n1015_, new_n1013_ );
nor g0801 ( new_n1016_, new_n1015_, keyIn_0_63 );
nor g0802 ( new_n1017_, new_n1016_, new_n1014_ );
nor g0803 ( new_n1018_, new_n1017_, new_n1002_ );
not g0804 ( new_n1019_, new_n1018_ );
nor g0805 ( new_n1020_, new_n1019_, new_n1006_ );
nand g0806 ( new_n1021_, new_n1019_, new_n1006_ );
not g0807 ( new_n1022_, N165 );
nor g0808 ( new_n1023_, new_n916_, new_n1022_ );
not g0809 ( new_n1024_, N171 );
nor g0810 ( new_n1025_, new_n926_, new_n1024_ );
not g0811 ( new_n1026_, new_n1025_ );
nor g0812 ( new_n1027_, new_n918_, new_n1026_ );
nor g0813 ( new_n1028_, new_n1027_, new_n1023_ );
nand g0814 ( new_n1029_, new_n1021_, new_n1028_ );
nor g0815 ( new_n1030_, new_n1029_, new_n1020_ );
not g0816 ( new_n1031_, new_n1030_ );
nor g0817 ( new_n1032_, new_n1005_, new_n1031_ );
nand g0818 ( new_n1033_, new_n1032_, new_n998_ );
nand g0819 ( new_n1034_, new_n1033_, keyIn_0_88 );
not g0820 ( new_n1035_, keyIn_0_88 );
not g0821 ( new_n1036_, keyIn_0_87 );
nor g0822 ( new_n1037_, new_n1001_, new_n1002_ );
nor g0823 ( new_n1038_, new_n1037_, new_n1036_ );
nand g0824 ( new_n1039_, new_n996_, new_n1003_ );
nand g0825 ( new_n1040_, new_n1039_, new_n1030_ );
nor g0826 ( new_n1041_, new_n1038_, new_n1040_ );
nand g0827 ( new_n1042_, new_n1041_, new_n1035_ );
nand g0828 ( new_n1043_, new_n1042_, new_n1034_ );
nor g0829 ( new_n1044_, new_n1043_, new_n906_ );
nor g0830 ( new_n1045_, new_n1044_, keyIn_0_101 );
not g0831 ( new_n1046_, N159 );
nor g0832 ( new_n1047_, new_n904_, new_n1046_ );
nor g0833 ( new_n1048_, new_n1047_, keyIn_0_51 );
nand g0834 ( new_n1049_, new_n1047_, keyIn_0_51 );
not g0835 ( new_n1050_, new_n1049_ );
nor g0836 ( new_n1051_, new_n1050_, new_n1048_ );
not g0837 ( new_n1052_, new_n1051_ );
nand g0838 ( new_n1053_, new_n1044_, keyIn_0_101 );
nand g0839 ( new_n1054_, new_n1053_, new_n1052_ );
nor g0840 ( new_n1055_, new_n1054_, new_n1045_ );
nor g0841 ( new_n1056_, new_n1055_, new_n879_ );
nand g0842 ( new_n1057_, new_n1055_, new_n879_ );
not g0843 ( new_n1058_, new_n1057_ );
nor g0844 ( new_n1059_, new_n1058_, new_n1056_ );
not g0845 ( new_n1060_, new_n1059_ );
nand g0846 ( new_n1061_, new_n1060_, new_n878_ );
nand g0847 ( new_n1062_, new_n1059_, keyIn_0_113 );
nand g0848 ( N866, new_n1061_, new_n1062_ );
not g0849 ( new_n1064_, keyIn_0_111 );
not g0850 ( new_n1065_, keyIn_0_105 );
not g0851 ( new_n1066_, keyIn_0_91 );
nor g0852 ( new_n1067_, new_n995_, new_n1013_ );
not g0853 ( new_n1068_, new_n1067_ );
nor g0854 ( new_n1069_, new_n949_, new_n1068_ );
nand g0855 ( new_n1070_, new_n1069_, keyIn_0_82 );
not g0856 ( new_n1071_, keyIn_0_82 );
not g0857 ( new_n1072_, new_n1069_ );
nand g0858 ( new_n1073_, new_n1072_, new_n1071_ );
nand g0859 ( new_n1074_, new_n1073_, new_n1070_ );
nor g0860 ( new_n1075_, new_n1000_, new_n1067_ );
not g0861 ( new_n1076_, new_n1075_ );
nand g0862 ( new_n1077_, new_n1076_, keyIn_0_81 );
not g0863 ( new_n1078_, keyIn_0_81 );
nand g0864 ( new_n1079_, new_n1075_, new_n1078_ );
nand g0865 ( new_n1080_, new_n1077_, new_n1079_ );
nand g0866 ( new_n1081_, new_n1080_, new_n1074_ );
nand g0867 ( new_n1082_, new_n1081_, new_n1066_ );
nor g0868 ( new_n1083_, new_n1081_, new_n1066_ );
nor g0869 ( new_n1084_, new_n1083_, new_n532_ );
nand g0870 ( new_n1085_, new_n1084_, new_n1082_ );
not g0871 ( new_n1086_, new_n1085_ );
nor g0872 ( new_n1087_, new_n1086_, keyIn_0_99 );
nand g0873 ( new_n1088_, N101, N210 );
nand g0874 ( new_n1089_, new_n1086_, keyIn_0_99 );
nand g0875 ( new_n1090_, new_n1089_, new_n1088_ );
nor g0876 ( new_n1091_, new_n1090_, new_n1087_ );
nor g0877 ( new_n1092_, new_n1091_, new_n1065_ );
nand g0878 ( new_n1093_, new_n1091_, new_n1065_ );
not g0879 ( new_n1094_, new_n1093_ );
nor g0880 ( new_n1095_, new_n1094_, new_n1092_ );
nor g0881 ( new_n1096_, new_n1017_, new_n800_ );
not g0882 ( new_n1097_, new_n1096_ );
nor g0883 ( new_n1098_, new_n1097_, keyIn_0_69 );
nand g0884 ( new_n1099_, new_n1097_, keyIn_0_69 );
nor g0885 ( new_n1100_, new_n1068_, new_n544_ );
nand g0886 ( new_n1101_, new_n988_, N246 );
nand g0887 ( new_n1102_, new_n867_, N177 );
nand g0888 ( new_n1103_, new_n1101_, new_n1102_ );
nor g0889 ( new_n1104_, new_n1100_, new_n1103_ );
nand g0890 ( new_n1105_, new_n1099_, new_n1104_ );
nor g0891 ( new_n1106_, new_n1105_, new_n1098_ );
not g0892 ( new_n1107_, new_n1106_ );
nor g0893 ( new_n1108_, new_n1095_, new_n1107_ );
not g0894 ( new_n1109_, new_n1108_ );
nand g0895 ( new_n1110_, new_n1109_, new_n1064_ );
not g0896 ( new_n1111_, new_n1110_ );
nor g0897 ( new_n1112_, new_n1109_, new_n1064_ );
nor g0898 ( new_n1113_, new_n1111_, new_n1112_ );
not g0899 ( new_n1114_, new_n1113_ );
nor g0900 ( new_n1115_, new_n1114_, keyIn_0_117 );
nand g0901 ( new_n1116_, new_n1114_, keyIn_0_117 );
not g0902 ( new_n1117_, new_n1116_ );
nor g0903 ( new_n1118_, new_n1117_, new_n1115_ );
not g0904 ( new_n1119_, new_n1118_ );
nand g0905 ( new_n1120_, new_n1119_, keyIn_0_121 );
not g0906 ( new_n1121_, keyIn_0_121 );
nand g0907 ( new_n1122_, new_n1118_, new_n1121_ );
nand g0908 ( N874, new_n1120_, new_n1122_ );
not g0909 ( new_n1124_, keyIn_0_125 );
not g0910 ( new_n1125_, keyIn_0_122 );
not g0911 ( new_n1126_, keyIn_0_108 );
not g0912 ( new_n1127_, keyIn_0_102 );
not g0913 ( new_n1128_, keyIn_0_62 );
not g0914 ( new_n1129_, new_n906_ );
nand g0915 ( new_n1130_, new_n1052_, new_n1129_ );
nand g0916 ( new_n1131_, new_n1130_, new_n1128_ );
not g0917 ( new_n1132_, new_n1131_ );
nor g0918 ( new_n1133_, new_n1130_, new_n1128_ );
nor g0919 ( new_n1134_, new_n1132_, new_n1133_ );
nand g0920 ( new_n1135_, new_n1043_, new_n1134_ );
nand g0921 ( new_n1136_, new_n1135_, keyIn_0_93 );
not g0922 ( new_n1137_, keyIn_0_93 );
not g0923 ( new_n1138_, new_n1135_ );
nand g0924 ( new_n1139_, new_n1138_, new_n1137_ );
nand g0925 ( new_n1140_, new_n1139_, new_n1136_ );
nor g0926 ( new_n1141_, new_n1041_, new_n1035_ );
nor g0927 ( new_n1142_, new_n1033_, keyIn_0_88 );
nor g0928 ( new_n1143_, new_n1141_, new_n1142_ );
not g0929 ( new_n1144_, new_n1134_ );
nand g0930 ( new_n1145_, new_n1143_, new_n1144_ );
nand g0931 ( new_n1146_, new_n1145_, keyIn_0_94 );
not g0932 ( new_n1147_, keyIn_0_94 );
nor g0933 ( new_n1148_, new_n1043_, new_n1134_ );
nand g0934 ( new_n1149_, new_n1148_, new_n1147_ );
nand g0935 ( new_n1150_, new_n1146_, new_n1149_ );
nand g0936 ( new_n1151_, new_n1140_, new_n1150_ );
nand g0937 ( new_n1152_, new_n1151_, new_n1127_ );
nor g0938 ( new_n1153_, new_n1151_, new_n1127_ );
nor g0939 ( new_n1154_, new_n1153_, new_n532_ );
nand g0940 ( new_n1155_, new_n1154_, new_n1152_ );
nor g0941 ( new_n1156_, new_n1155_, new_n1126_ );
not g0942 ( new_n1157_, new_n1156_ );
nand g0943 ( new_n1158_, new_n497_, N210 );
nand g0944 ( new_n1159_, new_n1155_, new_n1126_ );
nand g0945 ( new_n1160_, new_n1159_, new_n1158_ );
not g0946 ( new_n1161_, new_n1160_ );
nand g0947 ( new_n1162_, new_n1161_, new_n1157_ );
nand g0948 ( new_n1163_, new_n1162_, keyIn_0_114 );
not g0949 ( new_n1164_, keyIn_0_114 );
nor g0950 ( new_n1165_, new_n1160_, new_n1156_ );
nand g0951 ( new_n1166_, new_n1165_, new_n1164_ );
nand g0952 ( new_n1167_, new_n1163_, new_n1166_ );
nor g0953 ( new_n1168_, new_n1134_, new_n544_ );
nor g0954 ( new_n1169_, new_n1052_, new_n800_ );
nor g0955 ( new_n1170_, new_n904_, new_n808_ );
nor g0956 ( new_n1171_, new_n550_, new_n1046_ );
nor g0957 ( new_n1172_, new_n1170_, new_n1171_ );
not g0958 ( new_n1173_, new_n1172_ );
nor g0959 ( new_n1174_, new_n1169_, new_n1173_ );
not g0960 ( new_n1175_, new_n1174_ );
nor g0961 ( new_n1176_, new_n1168_, new_n1175_ );
nand g0962 ( new_n1177_, new_n1167_, new_n1176_ );
nand g0963 ( new_n1178_, new_n1177_, keyIn_0_118 );
not g0964 ( new_n1179_, new_n1178_ );
nor g0965 ( new_n1180_, new_n1177_, keyIn_0_118 );
nor g0966 ( new_n1181_, new_n1179_, new_n1180_ );
nor g0967 ( new_n1182_, new_n1181_, new_n1125_ );
not g0968 ( new_n1183_, keyIn_0_118 );
not g0969 ( new_n1184_, new_n1177_ );
nand g0970 ( new_n1185_, new_n1184_, new_n1183_ );
nand g0971 ( new_n1186_, new_n1185_, new_n1178_ );
nor g0972 ( new_n1187_, new_n1186_, keyIn_0_122 );
nor g0973 ( new_n1188_, new_n1182_, new_n1187_ );
nor g0974 ( new_n1189_, new_n1188_, new_n1124_ );
nand g0975 ( new_n1190_, new_n1186_, keyIn_0_122 );
nand g0976 ( new_n1191_, new_n1181_, new_n1125_ );
nand g0977 ( new_n1192_, new_n1191_, new_n1190_ );
nor g0978 ( new_n1193_, new_n1192_, keyIn_0_125 );
nor g0979 ( N878, new_n1189_, new_n1193_ );
not g0980 ( new_n1195_, keyIn_0_126 );
not g0981 ( new_n1196_, keyIn_0_123 );
not g0982 ( new_n1197_, keyIn_0_119 );
not g0983 ( new_n1198_, keyIn_0_115 );
not g0984 ( new_n1199_, keyIn_0_109 );
not g0985 ( new_n1200_, keyIn_0_103 );
not g0986 ( new_n1201_, keyIn_0_95 );
nor g0987 ( new_n1202_, new_n918_, new_n1023_ );
not g0988 ( new_n1203_, new_n1202_ );
not g0989 ( new_n1204_, keyIn_0_89 );
not g0990 ( new_n1205_, new_n928_ );
nand g0991 ( new_n1206_, new_n996_, new_n1205_ );
nor g0992 ( new_n1207_, new_n1206_, keyIn_0_86 );
not g0993 ( new_n1208_, new_n1207_ );
not g0994 ( new_n1209_, keyIn_0_86 );
nor g0995 ( new_n1210_, new_n1001_, new_n928_ );
nor g0996 ( new_n1211_, new_n1210_, new_n1209_ );
not g0997 ( new_n1212_, new_n1017_ );
nand g0998 ( new_n1213_, new_n1212_, new_n1205_ );
nand g0999 ( new_n1214_, new_n1213_, new_n1026_ );
nor g1000 ( new_n1215_, new_n1211_, new_n1214_ );
nand g1001 ( new_n1216_, new_n1215_, new_n1208_ );
nand g1002 ( new_n1217_, new_n1216_, new_n1204_ );
nand g1003 ( new_n1218_, new_n1206_, keyIn_0_86 );
not g1004 ( new_n1219_, new_n1214_ );
nand g1005 ( new_n1220_, new_n1218_, new_n1219_ );
nor g1006 ( new_n1221_, new_n1220_, new_n1207_ );
nand g1007 ( new_n1222_, new_n1221_, keyIn_0_89 );
nand g1008 ( new_n1223_, new_n1217_, new_n1222_ );
nand g1009 ( new_n1224_, new_n1223_, new_n1203_ );
nand g1010 ( new_n1225_, new_n1224_, new_n1201_ );
not g1011 ( new_n1226_, new_n1225_ );
not g1012 ( new_n1227_, keyIn_0_96 );
nor g1013 ( new_n1228_, new_n1223_, new_n1203_ );
nor g1014 ( new_n1229_, new_n1228_, new_n1227_ );
nor g1015 ( new_n1230_, new_n1226_, new_n1229_ );
nor g1016 ( new_n1231_, new_n1221_, keyIn_0_89 );
nor g1017 ( new_n1232_, new_n1216_, new_n1204_ );
nor g1018 ( new_n1233_, new_n1232_, new_n1231_ );
nand g1019 ( new_n1234_, new_n1233_, new_n1202_ );
nor g1020 ( new_n1235_, new_n1234_, keyIn_0_96 );
nor g1021 ( new_n1236_, new_n1224_, new_n1201_ );
nor g1022 ( new_n1237_, new_n1235_, new_n1236_ );
nand g1023 ( new_n1238_, new_n1230_, new_n1237_ );
nand g1024 ( new_n1239_, new_n1238_, new_n1200_ );
nand g1025 ( new_n1240_, new_n1234_, keyIn_0_96 );
nand g1026 ( new_n1241_, new_n1240_, new_n1225_ );
nand g1027 ( new_n1242_, new_n1228_, new_n1227_ );
nor g1028 ( new_n1243_, new_n1233_, new_n1202_ );
nand g1029 ( new_n1244_, new_n1243_, keyIn_0_95 );
nand g1030 ( new_n1245_, new_n1244_, new_n1242_ );
nor g1031 ( new_n1246_, new_n1245_, new_n1241_ );
nand g1032 ( new_n1247_, new_n1246_, keyIn_0_103 );
nand g1033 ( new_n1248_, new_n1239_, new_n1247_ );
nand g1034 ( new_n1249_, new_n1248_, N219 );
nor g1035 ( new_n1250_, new_n1249_, new_n1199_ );
nand g1036 ( new_n1251_, N91, N210 );
nand g1037 ( new_n1252_, new_n1249_, new_n1199_ );
nand g1038 ( new_n1253_, new_n1252_, new_n1251_ );
nor g1039 ( new_n1254_, new_n1253_, new_n1250_ );
nand g1040 ( new_n1255_, new_n1254_, new_n1198_ );
nor g1041 ( new_n1256_, new_n1254_, new_n1198_ );
nor g1042 ( new_n1257_, new_n1203_, new_n544_ );
nand g1043 ( new_n1258_, new_n1023_, N237 );
nor g1044 ( new_n1259_, new_n916_, new_n808_ );
nor g1045 ( new_n1260_, new_n550_, new_n1022_ );
nor g1046 ( new_n1261_, new_n1259_, new_n1260_ );
nand g1047 ( new_n1262_, new_n1261_, new_n1258_ );
nor g1048 ( new_n1263_, new_n1257_, new_n1262_ );
not g1049 ( new_n1264_, new_n1263_ );
nor g1050 ( new_n1265_, new_n1256_, new_n1264_ );
nand g1051 ( new_n1266_, new_n1265_, new_n1255_ );
nand g1052 ( new_n1267_, new_n1266_, new_n1197_ );
not g1053 ( new_n1268_, new_n1255_ );
not g1054 ( new_n1269_, new_n1250_ );
not g1055 ( new_n1270_, new_n1253_ );
nand g1056 ( new_n1271_, new_n1270_, new_n1269_ );
nand g1057 ( new_n1272_, new_n1271_, keyIn_0_115 );
nand g1058 ( new_n1273_, new_n1272_, new_n1263_ );
nor g1059 ( new_n1274_, new_n1273_, new_n1268_ );
nand g1060 ( new_n1275_, new_n1274_, keyIn_0_119 );
nand g1061 ( new_n1276_, new_n1275_, new_n1267_ );
nand g1062 ( new_n1277_, new_n1276_, new_n1196_ );
nor g1063 ( new_n1278_, new_n1274_, keyIn_0_119 );
nor g1064 ( new_n1279_, new_n1266_, new_n1197_ );
nor g1065 ( new_n1280_, new_n1278_, new_n1279_ );
nand g1066 ( new_n1281_, new_n1280_, keyIn_0_123 );
nand g1067 ( new_n1282_, new_n1281_, new_n1277_ );
nand g1068 ( new_n1283_, new_n1282_, new_n1195_ );
nor g1069 ( new_n1284_, new_n1280_, keyIn_0_123 );
nor g1070 ( new_n1285_, new_n1276_, new_n1196_ );
nor g1071 ( new_n1286_, new_n1284_, new_n1285_ );
nand g1072 ( new_n1287_, new_n1286_, keyIn_0_126 );
nand g1073 ( N879, new_n1287_, new_n1283_ );
not g1074 ( new_n1289_, keyIn_0_127 );
not g1075 ( new_n1290_, keyIn_0_85 );
nor g1076 ( new_n1291_, new_n1001_, new_n1290_ );
nand g1077 ( new_n1292_, new_n1001_, new_n1290_ );
nand g1078 ( new_n1293_, new_n1292_, new_n1017_ );
nor g1079 ( new_n1294_, new_n1293_, new_n1291_ );
nor g1080 ( new_n1295_, new_n1294_, keyIn_0_90 );
not g1081 ( new_n1296_, new_n1295_ );
nand g1082 ( new_n1297_, new_n1294_, keyIn_0_90 );
nand g1083 ( new_n1298_, new_n1296_, new_n1297_ );
nor g1084 ( new_n1299_, new_n928_, new_n1025_ );
nand g1085 ( new_n1300_, new_n1298_, new_n1299_ );
nand g1086 ( new_n1301_, new_n1300_, keyIn_0_98 );
not g1087 ( new_n1302_, new_n1297_ );
nor g1088 ( new_n1303_, new_n1302_, new_n1295_ );
not g1089 ( new_n1304_, new_n1299_ );
nand g1090 ( new_n1305_, new_n1303_, new_n1304_ );
nand g1091 ( new_n1306_, new_n1305_, keyIn_0_97 );
nand g1092 ( new_n1307_, new_n1306_, new_n1301_ );
not g1093 ( new_n1308_, new_n1307_ );
nor g1094 ( new_n1309_, new_n1305_, keyIn_0_97 );
nor g1095 ( new_n1310_, new_n1300_, keyIn_0_98 );
nor g1096 ( new_n1311_, new_n1309_, new_n1310_ );
nand g1097 ( new_n1312_, new_n1308_, new_n1311_ );
nor g1098 ( new_n1313_, new_n1312_, keyIn_0_104 );
not g1099 ( new_n1314_, new_n1313_ );
not g1100 ( new_n1315_, keyIn_0_104 );
not g1101 ( new_n1316_, keyIn_0_97 );
nor g1102 ( new_n1317_, new_n1298_, new_n1299_ );
nand g1103 ( new_n1318_, new_n1317_, new_n1316_ );
not g1104 ( new_n1319_, keyIn_0_98 );
not g1105 ( new_n1320_, new_n1300_ );
nand g1106 ( new_n1321_, new_n1320_, new_n1319_ );
nand g1107 ( new_n1322_, new_n1321_, new_n1318_ );
nor g1108 ( new_n1323_, new_n1322_, new_n1307_ );
nor g1109 ( new_n1324_, new_n1323_, new_n1315_ );
nor g1110 ( new_n1325_, new_n1324_, new_n532_ );
nand g1111 ( new_n1326_, new_n1325_, new_n1314_ );
nor g1112 ( new_n1327_, new_n1326_, keyIn_0_110 );
not g1113 ( new_n1328_, new_n1327_ );
nand g1114 ( new_n1329_, N96, N210 );
not g1115 ( new_n1330_, new_n1329_ );
not g1116 ( new_n1331_, keyIn_0_110 );
nand g1117 ( new_n1332_, new_n1312_, keyIn_0_104 );
nand g1118 ( new_n1333_, new_n1332_, N219 );
nor g1119 ( new_n1334_, new_n1333_, new_n1313_ );
nor g1120 ( new_n1335_, new_n1334_, new_n1331_ );
nor g1121 ( new_n1336_, new_n1335_, new_n1330_ );
nand g1122 ( new_n1337_, new_n1336_, new_n1328_ );
nand g1123 ( new_n1338_, new_n1337_, keyIn_0_116 );
not g1124 ( new_n1339_, keyIn_0_116 );
nand g1125 ( new_n1340_, new_n1326_, keyIn_0_110 );
nand g1126 ( new_n1341_, new_n1340_, new_n1329_ );
nor g1127 ( new_n1342_, new_n1341_, new_n1327_ );
nand g1128 ( new_n1343_, new_n1342_, new_n1339_ );
nand g1129 ( new_n1344_, new_n1343_, new_n1338_ );
nor g1130 ( new_n1345_, new_n1304_, new_n544_ );
nand g1131 ( new_n1346_, new_n1025_, N237 );
nor g1132 ( new_n1347_, new_n926_, new_n808_ );
nor g1133 ( new_n1348_, new_n550_, new_n1024_ );
nor g1134 ( new_n1349_, new_n1347_, new_n1348_ );
nand g1135 ( new_n1350_, new_n1349_, new_n1346_ );
nor g1136 ( new_n1351_, new_n1345_, new_n1350_ );
nand g1137 ( new_n1352_, new_n1344_, new_n1351_ );
nand g1138 ( new_n1353_, new_n1352_, keyIn_0_120 );
nor g1139 ( new_n1354_, new_n1352_, keyIn_0_120 );
not g1140 ( new_n1355_, new_n1354_ );
nand g1141 ( new_n1356_, new_n1355_, new_n1353_ );
nand g1142 ( new_n1357_, new_n1356_, keyIn_0_124 );
not g1143 ( new_n1358_, keyIn_0_124 );
not g1144 ( new_n1359_, new_n1353_ );
nor g1145 ( new_n1360_, new_n1359_, new_n1354_ );
nand g1146 ( new_n1361_, new_n1360_, new_n1358_ );
nand g1147 ( new_n1362_, new_n1361_, new_n1357_ );
nand g1148 ( new_n1363_, new_n1362_, new_n1289_ );
nor g1149 ( new_n1364_, new_n1360_, new_n1358_ );
nor g1150 ( new_n1365_, new_n1356_, keyIn_0_124 );
nor g1151 ( new_n1366_, new_n1364_, new_n1365_ );
nand g1152 ( new_n1367_, new_n1366_, keyIn_0_127 );
nand g1153 ( N880, new_n1367_, new_n1363_ );
endmodule