module add_mul_combine_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, Result_mul_0_, Result_mul_1_, 
        Result_mul_2_, Result_mul_3_, Result_mul_4_, Result_mul_5_, 
        Result_mul_6_, Result_mul_7_, Result_mul_8_, Result_mul_9_, 
        Result_mul_10_, Result_mul_11_, Result_mul_12_, Result_mul_13_, 
        Result_mul_14_, Result_mul_15_, Result_mul_16_, Result_mul_17_, 
        Result_mul_18_, Result_mul_19_, Result_mul_20_, Result_mul_21_, 
        Result_mul_22_, Result_mul_23_, Result_mul_24_, Result_mul_25_, 
        Result_mul_26_, Result_mul_27_, Result_mul_28_, Result_mul_29_, 
        Result_mul_30_, Result_mul_31_, Result_mul_32_, Result_mul_33_, 
        Result_mul_34_, Result_mul_35_, Result_mul_36_, Result_mul_37_, 
        Result_mul_38_, Result_mul_39_, Result_mul_40_, Result_mul_41_, 
        Result_mul_42_, Result_mul_43_, Result_mul_44_, Result_mul_45_, 
        Result_mul_46_, Result_mul_47_, Result_mul_48_, Result_mul_49_, 
        Result_mul_50_, Result_mul_51_, Result_mul_52_, Result_mul_53_, 
        Result_mul_54_, Result_mul_55_, Result_mul_56_, Result_mul_57_, 
        Result_mul_58_, Result_mul_59_, Result_mul_60_, Result_mul_61_, 
        Result_mul_62_, Result_mul_63_, Result_add_0_, Result_add_1_, 
        Result_add_2_, Result_add_3_, Result_add_4_, Result_add_5_, 
        Result_add_6_, Result_add_7_, Result_add_8_, Result_add_9_, 
        Result_add_10_, Result_add_11_, Result_add_12_, Result_add_13_, 
        Result_add_14_, Result_add_15_, Result_add_16_, Result_add_17_, 
        Result_add_18_, Result_add_19_, Result_add_20_, Result_add_21_, 
        Result_add_22_, Result_add_23_, Result_add_24_, Result_add_25_, 
        Result_add_26_, Result_add_27_, Result_add_28_, Result_add_29_, 
        Result_add_30_, Result_add_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_mul_16_, Result_mul_17_, Result_mul_18_, Result_mul_19_,
         Result_mul_20_, Result_mul_21_, Result_mul_22_, Result_mul_23_,
         Result_mul_24_, Result_mul_25_, Result_mul_26_, Result_mul_27_,
         Result_mul_28_, Result_mul_29_, Result_mul_30_, Result_mul_31_,
         Result_mul_32_, Result_mul_33_, Result_mul_34_, Result_mul_35_,
         Result_mul_36_, Result_mul_37_, Result_mul_38_, Result_mul_39_,
         Result_mul_40_, Result_mul_41_, Result_mul_42_, Result_mul_43_,
         Result_mul_44_, Result_mul_45_, Result_mul_46_, Result_mul_47_,
         Result_mul_48_, Result_mul_49_, Result_mul_50_, Result_mul_51_,
         Result_mul_52_, Result_mul_53_, Result_mul_54_, Result_mul_55_,
         Result_mul_56_, Result_mul_57_, Result_mul_58_, Result_mul_59_,
         Result_mul_60_, Result_mul_61_, Result_mul_62_, Result_mul_63_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_,
         Result_add_8_, Result_add_9_, Result_add_10_, Result_add_11_,
         Result_add_12_, Result_add_13_, Result_add_14_, Result_add_15_,
         Result_add_16_, Result_add_17_, Result_add_18_, Result_add_19_,
         Result_add_20_, Result_add_21_, Result_add_22_, Result_add_23_,
         Result_add_24_, Result_add_25_, Result_add_26_, Result_add_27_,
         Result_add_28_, Result_add_29_, Result_add_30_, Result_add_31_;
  wire   n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498;

  INV_X2 U8367 ( .A(b_24_), .ZN(n10120) );
  INV_X2 U8368 ( .A(b_18_), .ZN(n11623) );
  INV_X2 U8369 ( .A(b_16_), .ZN(n12110) );
  INV_X2 U8370 ( .A(b_8_), .ZN(n14123) );
  INV_X2 U8371 ( .A(b_19_), .ZN(n11356) );
  INV_X2 U8372 ( .A(b_11_), .ZN(n13332) );
  INV_X2 U8373 ( .A(b_28_), .ZN(n9105) );
  INV_X2 U8374 ( .A(b_2_), .ZN(n15595) );
  INV_X2 U8375 ( .A(b_21_), .ZN(n10876) );
  INV_X2 U8376 ( .A(b_10_), .ZN(n13629) );
  INV_X2 U8377 ( .A(b_25_), .ZN(n9864) );
  INV_X2 U8378 ( .A(b_17_), .ZN(n11859) );
  INV_X2 U8379 ( .A(a_7_), .ZN(n8425) );
  INV_X2 U8380 ( .A(a_17_), .ZN(n8371) );
  INV_X2 U8381 ( .A(a_20_), .ZN(n9047) );
  INV_X2 U8382 ( .A(a_13_), .ZN(n8996) );
  INV_X2 U8383 ( .A(a_18_), .ZN(n9291) );
  INV_X2 U8384 ( .A(a_10_), .ZN(n8402) );
  INV_X2 U8385 ( .A(a_4_), .ZN(n8439) );
  INV_X2 U8386 ( .A(a_26_), .ZN(n9344) );
  INV_X2 U8387 ( .A(a_1_), .ZN(n8569) );
  INV_X2 U8388 ( .A(a_25_), .ZN(n8788) );
  NAND2_X2 U8389 ( .A1(a_30_), .A2(n16108), .ZN(n8303) );
  NAND2_X2 U8390 ( .A1(a_31_), .A2(n16105), .ZN(n8299) );
  INV_X2 U8391 ( .A(a_24_), .ZN(n8779) );
  INV_X2 U8392 ( .A(a_2_), .ZN(n8448) );
  INV_X2 U8393 ( .A(a_5_), .ZN(n8938) );
  INV_X2 U8394 ( .A(a_15_), .ZN(n8850) );
  INV_X2 U8395 ( .A(a_27_), .ZN(n8797) );
  INV_X2 U8396 ( .A(a_12_), .ZN(n8393) );
  INV_X2 U8397 ( .A(b_7_), .ZN(n14345) );
  INV_X2 U8398 ( .A(a_9_), .ZN(n8971) );
  INV_X2 U8399 ( .A(a_3_), .ZN(n8900) );
  INV_X2 U8400 ( .A(b_1_), .ZN(n15890) );
  INV_X2 U8401 ( .A(a_28_), .ZN(n8314) );
  INV_X2 U8402 ( .A(b_15_), .ZN(n12340) );
  INV_X2 U8403 ( .A(b_4_), .ZN(n15110) );
  INV_X2 U8404 ( .A(b_13_), .ZN(n12835) );
  INV_X2 U8405 ( .A(a_29_), .ZN(n9098) );
  INV_X2 U8406 ( .A(b_9_), .ZN(n13840) );
  INV_X2 U8407 ( .A(b_6_), .ZN(n14621) );
  INV_X2 U8408 ( .A(a_11_), .ZN(n8867) );
  INV_X2 U8409 ( .A(b_14_), .ZN(n12609) );
  INV_X2 U8410 ( .A(a_21_), .ZN(n8759) );
  INV_X2 U8411 ( .A(b_3_), .ZN(n15343) );
  INV_X2 U8412 ( .A(b_5_), .ZN(n14859) );
  XOR2_X1 U8413 ( .A(n8272), .B(n8273), .Z(Result_mul_9_) );
  NOR2_X1 U8414 ( .A1(n8274), .A2(n8275), .ZN(n8273) );
  NOR2_X1 U8415 ( .A1(n8276), .A2(n8277), .ZN(n8275) );
  INV_X1 U8416 ( .A(n8278), .ZN(n8276) );
  NAND2_X1 U8417 ( .A1(n8279), .A2(n8280), .ZN(n8278) );
  INV_X1 U8418 ( .A(n8281), .ZN(n8274) );
  XOR2_X1 U8419 ( .A(n8282), .B(n8283), .Z(Result_mul_8_) );
  XOR2_X1 U8420 ( .A(n8284), .B(n8285), .Z(Result_mul_7_) );
  NOR2_X1 U8421 ( .A1(n8286), .A2(n8287), .ZN(n8285) );
  NOR2_X1 U8422 ( .A1(n8288), .A2(n8289), .ZN(n8287) );
  INV_X1 U8423 ( .A(n8290), .ZN(n8288) );
  NAND2_X1 U8424 ( .A1(n8291), .A2(n8292), .ZN(n8290) );
  INV_X1 U8425 ( .A(n8293), .ZN(n8286) );
  XOR2_X1 U8426 ( .A(n8294), .B(n8295), .Z(Result_mul_6_) );
  NAND2_X1 U8427 ( .A1(n8296), .A2(n8297), .ZN(Result_mul_62_) );
  NAND2_X1 U8428 ( .A1(b_30_), .A2(n8298), .ZN(n8297) );
  NAND2_X1 U8429 ( .A1(n8299), .A2(n8300), .ZN(n8298) );
  NAND2_X1 U8430 ( .A1(a_31_), .A2(n8301), .ZN(n8300) );
  NAND2_X1 U8431 ( .A1(b_31_), .A2(n8302), .ZN(n8296) );
  NAND2_X1 U8432 ( .A1(n8303), .A2(n8304), .ZN(n8302) );
  NAND2_X1 U8433 ( .A1(a_30_), .A2(n8305), .ZN(n8304) );
  XNOR2_X1 U8434 ( .A(n8306), .B(n8307), .ZN(Result_mul_61_) );
  XOR2_X1 U8435 ( .A(n8308), .B(n8309), .Z(n8307) );
  XOR2_X1 U8436 ( .A(n8310), .B(n8311), .Z(Result_mul_60_) );
  XOR2_X1 U8437 ( .A(n8312), .B(n8313), .Z(n8310) );
  NOR2_X1 U8438 ( .A1(n8314), .A2(n8301), .ZN(n8313) );
  XOR2_X1 U8439 ( .A(n8315), .B(n8316), .Z(Result_mul_5_) );
  NOR2_X1 U8440 ( .A1(n8317), .A2(n8318), .ZN(n8316) );
  NOR2_X1 U8441 ( .A1(n8319), .A2(n8320), .ZN(n8318) );
  INV_X1 U8442 ( .A(n8321), .ZN(n8319) );
  NAND2_X1 U8443 ( .A1(n8322), .A2(n8323), .ZN(n8321) );
  INV_X1 U8444 ( .A(n8324), .ZN(n8317) );
  XNOR2_X1 U8445 ( .A(n8325), .B(n8326), .ZN(Result_mul_59_) );
  XNOR2_X1 U8446 ( .A(n8327), .B(n8328), .ZN(n8325) );
  XNOR2_X1 U8447 ( .A(n8329), .B(n8330), .ZN(Result_mul_58_) );
  XOR2_X1 U8448 ( .A(n8331), .B(n8332), .Z(n8330) );
  XNOR2_X1 U8449 ( .A(n8333), .B(n8334), .ZN(Result_mul_57_) );
  XNOR2_X1 U8450 ( .A(n8335), .B(n8336), .ZN(n8333) );
  XNOR2_X1 U8451 ( .A(n8337), .B(n8338), .ZN(Result_mul_56_) );
  XNOR2_X1 U8452 ( .A(n8339), .B(n8340), .ZN(n8338) );
  XNOR2_X1 U8453 ( .A(n8341), .B(n8342), .ZN(Result_mul_55_) );
  NAND2_X1 U8454 ( .A1(n8343), .A2(n8344), .ZN(n8341) );
  XOR2_X1 U8455 ( .A(n8345), .B(n8346), .Z(Result_mul_54_) );
  XNOR2_X1 U8456 ( .A(n8347), .B(n8348), .ZN(n8345) );
  XNOR2_X1 U8457 ( .A(n8349), .B(n8350), .ZN(Result_mul_53_) );
  NAND2_X1 U8458 ( .A1(n8351), .A2(n8352), .ZN(n8349) );
  XNOR2_X1 U8459 ( .A(n8353), .B(n8354), .ZN(Result_mul_52_) );
  XOR2_X1 U8460 ( .A(n8355), .B(n8356), .Z(n8354) );
  XNOR2_X1 U8461 ( .A(n8357), .B(n8358), .ZN(Result_mul_51_) );
  NAND2_X1 U8462 ( .A1(n8359), .A2(n8360), .ZN(n8357) );
  XNOR2_X1 U8463 ( .A(n8361), .B(n8362), .ZN(Result_mul_50_) );
  XOR2_X1 U8464 ( .A(n8363), .B(n8364), .Z(n8362) );
  NAND2_X1 U8465 ( .A1(b_31_), .A2(a_18_), .ZN(n8364) );
  XOR2_X1 U8466 ( .A(n8365), .B(n8366), .Z(Result_mul_4_) );
  XOR2_X1 U8467 ( .A(n8367), .B(n8368), .Z(Result_mul_49_) );
  XOR2_X1 U8468 ( .A(n8369), .B(n8370), .Z(n8367) );
  NOR2_X1 U8469 ( .A1(n8371), .A2(n8301), .ZN(n8370) );
  XNOR2_X1 U8470 ( .A(n8372), .B(n8373), .ZN(Result_mul_48_) );
  XNOR2_X1 U8471 ( .A(n8374), .B(n8375), .ZN(n8372) );
  NOR2_X1 U8472 ( .A1(n8376), .A2(n8301), .ZN(n8375) );
  XOR2_X1 U8473 ( .A(n8377), .B(n8378), .Z(Result_mul_47_) );
  XNOR2_X1 U8474 ( .A(n8379), .B(n8380), .ZN(n8378) );
  NAND2_X1 U8475 ( .A1(b_31_), .A2(a_15_), .ZN(n8380) );
  XOR2_X1 U8476 ( .A(n8381), .B(n8382), .Z(Result_mul_46_) );
  XNOR2_X1 U8477 ( .A(n8383), .B(n8384), .ZN(n8382) );
  NAND2_X1 U8478 ( .A1(b_31_), .A2(a_14_), .ZN(n8384) );
  XOR2_X1 U8479 ( .A(n8385), .B(n8386), .Z(Result_mul_45_) );
  XNOR2_X1 U8480 ( .A(n8387), .B(n8388), .ZN(n8386) );
  NAND2_X1 U8481 ( .A1(b_31_), .A2(a_13_), .ZN(n8388) );
  XOR2_X1 U8482 ( .A(n8389), .B(n8390), .Z(Result_mul_44_) );
  XOR2_X1 U8483 ( .A(n8391), .B(n8392), .Z(n8389) );
  NOR2_X1 U8484 ( .A1(n8393), .A2(n8301), .ZN(n8392) );
  XOR2_X1 U8485 ( .A(n8394), .B(n8395), .Z(Result_mul_43_) );
  XNOR2_X1 U8486 ( .A(n8396), .B(n8397), .ZN(n8395) );
  NAND2_X1 U8487 ( .A1(b_31_), .A2(a_11_), .ZN(n8397) );
  XNOR2_X1 U8488 ( .A(n8398), .B(n8399), .ZN(Result_mul_42_) );
  XNOR2_X1 U8489 ( .A(n8400), .B(n8401), .ZN(n8398) );
  NOR2_X1 U8490 ( .A1(n8402), .A2(n8301), .ZN(n8401) );
  XOR2_X1 U8491 ( .A(n8403), .B(n8404), .Z(Result_mul_41_) );
  XNOR2_X1 U8492 ( .A(n8405), .B(n8406), .ZN(n8404) );
  NAND2_X1 U8493 ( .A1(b_31_), .A2(a_9_), .ZN(n8406) );
  XOR2_X1 U8494 ( .A(n8407), .B(n8408), .Z(Result_mul_40_) );
  XNOR2_X1 U8495 ( .A(n8409), .B(n8410), .ZN(n8408) );
  NAND2_X1 U8496 ( .A1(b_31_), .A2(a_8_), .ZN(n8410) );
  XOR2_X1 U8497 ( .A(n8411), .B(n8412), .Z(Result_mul_3_) );
  NOR2_X1 U8498 ( .A1(n8413), .A2(n8414), .ZN(n8412) );
  NOR2_X1 U8499 ( .A1(n8415), .A2(n8416), .ZN(n8414) );
  INV_X1 U8500 ( .A(n8417), .ZN(n8415) );
  NAND2_X1 U8501 ( .A1(n8418), .A2(n8419), .ZN(n8417) );
  INV_X1 U8502 ( .A(n8420), .ZN(n8413) );
  XOR2_X1 U8503 ( .A(n8421), .B(n8422), .Z(Result_mul_39_) );
  XOR2_X1 U8504 ( .A(n8423), .B(n8424), .Z(n8421) );
  NOR2_X1 U8505 ( .A1(n8425), .A2(n8301), .ZN(n8424) );
  XOR2_X1 U8506 ( .A(n8426), .B(n8427), .Z(Result_mul_38_) );
  XOR2_X1 U8507 ( .A(n8428), .B(n8429), .Z(n8426) );
  NOR2_X1 U8508 ( .A1(n8430), .A2(n8301), .ZN(n8429) );
  XOR2_X1 U8509 ( .A(n8431), .B(n8432), .Z(Result_mul_37_) );
  XNOR2_X1 U8510 ( .A(n8433), .B(n8434), .ZN(n8432) );
  NAND2_X1 U8511 ( .A1(b_31_), .A2(a_5_), .ZN(n8434) );
  XNOR2_X1 U8512 ( .A(n8435), .B(n8436), .ZN(Result_mul_36_) );
  XNOR2_X1 U8513 ( .A(n8437), .B(n8438), .ZN(n8435) );
  NOR2_X1 U8514 ( .A1(n8439), .A2(n8301), .ZN(n8438) );
  XOR2_X1 U8515 ( .A(n8440), .B(n8441), .Z(Result_mul_35_) );
  XNOR2_X1 U8516 ( .A(n8442), .B(n8443), .ZN(n8441) );
  NAND2_X1 U8517 ( .A1(b_31_), .A2(a_3_), .ZN(n8443) );
  XOR2_X1 U8518 ( .A(n8444), .B(n8445), .Z(Result_mul_34_) );
  XOR2_X1 U8519 ( .A(n8446), .B(n8447), .Z(n8444) );
  NOR2_X1 U8520 ( .A1(n8448), .A2(n8301), .ZN(n8447) );
  XOR2_X1 U8521 ( .A(n8449), .B(n8450), .Z(Result_mul_33_) );
  XNOR2_X1 U8522 ( .A(n8451), .B(n8452), .ZN(n8450) );
  NAND2_X1 U8523 ( .A1(b_31_), .A2(a_1_), .ZN(n8452) );
  XNOR2_X1 U8524 ( .A(n8453), .B(n8454), .ZN(Result_mul_32_) );
  XNOR2_X1 U8525 ( .A(n8455), .B(n8456), .ZN(n8453) );
  NOR2_X1 U8526 ( .A1(n8457), .A2(n8301), .ZN(n8456) );
  XOR2_X1 U8527 ( .A(n8458), .B(n8459), .Z(Result_mul_31_) );
  NOR2_X1 U8528 ( .A1(n8460), .A2(n8461), .ZN(Result_mul_30_) );
  NOR2_X1 U8529 ( .A1(n8462), .A2(n8463), .ZN(n8461) );
  INV_X1 U8530 ( .A(n8464), .ZN(n8463) );
  NOR2_X1 U8531 ( .A1(n8459), .A2(n8458), .ZN(n8462) );
  XOR2_X1 U8532 ( .A(n8465), .B(n8466), .Z(Result_mul_2_) );
  XNOR2_X1 U8533 ( .A(n8460), .B(n8467), .ZN(Result_mul_29_) );
  NAND2_X1 U8534 ( .A1(n8468), .A2(n8469), .ZN(n8467) );
  XNOR2_X1 U8535 ( .A(n8470), .B(n8471), .ZN(Result_mul_28_) );
  NAND2_X1 U8536 ( .A1(n8472), .A2(n8473), .ZN(n8471) );
  XNOR2_X1 U8537 ( .A(n8474), .B(n8475), .ZN(Result_mul_27_) );
  NAND2_X1 U8538 ( .A1(n8476), .A2(n8477), .ZN(n8475) );
  XNOR2_X1 U8539 ( .A(n8478), .B(n8479), .ZN(Result_mul_26_) );
  NAND2_X1 U8540 ( .A1(n8480), .A2(n8481), .ZN(n8479) );
  XNOR2_X1 U8541 ( .A(n8482), .B(n8483), .ZN(Result_mul_25_) );
  NAND2_X1 U8542 ( .A1(n8484), .A2(n8485), .ZN(n8483) );
  XNOR2_X1 U8543 ( .A(n8486), .B(n8487), .ZN(Result_mul_24_) );
  NAND2_X1 U8544 ( .A1(n8488), .A2(n8489), .ZN(n8487) );
  XNOR2_X1 U8545 ( .A(n8490), .B(n8491), .ZN(Result_mul_23_) );
  NAND2_X1 U8546 ( .A1(n8492), .A2(n8493), .ZN(n8491) );
  XNOR2_X1 U8547 ( .A(n8494), .B(n8495), .ZN(Result_mul_22_) );
  NAND2_X1 U8548 ( .A1(n8496), .A2(n8497), .ZN(n8495) );
  XNOR2_X1 U8549 ( .A(n8498), .B(n8499), .ZN(Result_mul_21_) );
  NAND2_X1 U8550 ( .A1(n8500), .A2(n8501), .ZN(n8499) );
  XNOR2_X1 U8551 ( .A(n8502), .B(n8503), .ZN(Result_mul_20_) );
  NAND2_X1 U8552 ( .A1(n8504), .A2(n8505), .ZN(n8503) );
  XNOR2_X1 U8553 ( .A(n8506), .B(n8507), .ZN(Result_mul_1_) );
  NAND2_X1 U8554 ( .A1(n8508), .A2(n8509), .ZN(n8507) );
  XOR2_X1 U8555 ( .A(n8510), .B(n8511), .Z(Result_mul_19_) );
  NOR2_X1 U8556 ( .A1(n8512), .A2(n8513), .ZN(n8511) );
  XNOR2_X1 U8557 ( .A(n8514), .B(n8515), .ZN(Result_mul_18_) );
  NAND2_X1 U8558 ( .A1(n8516), .A2(n8517), .ZN(n8515) );
  XOR2_X1 U8559 ( .A(n8518), .B(n8519), .Z(Result_mul_17_) );
  NOR2_X1 U8560 ( .A1(n8520), .A2(n8521), .ZN(n8519) );
  INV_X1 U8561 ( .A(n8522), .ZN(n8521) );
  NOR2_X1 U8562 ( .A1(n8523), .A2(n8524), .ZN(n8520) );
  INV_X1 U8563 ( .A(n8525), .ZN(n8524) );
  NAND2_X1 U8564 ( .A1(n8526), .A2(n8527), .ZN(n8525) );
  XNOR2_X1 U8565 ( .A(n8528), .B(n8529), .ZN(Result_mul_16_) );
  NAND2_X1 U8566 ( .A1(n8530), .A2(n8531), .ZN(n8529) );
  XNOR2_X1 U8567 ( .A(n8532), .B(n8533), .ZN(Result_mul_15_) );
  NAND2_X1 U8568 ( .A1(n8534), .A2(n8535), .ZN(n8533) );
  XOR2_X1 U8569 ( .A(n8536), .B(n8537), .Z(Result_mul_14_) );
  XOR2_X1 U8570 ( .A(n8538), .B(n8539), .Z(Result_mul_13_) );
  NOR2_X1 U8571 ( .A1(n8540), .A2(n8541), .ZN(n8539) );
  INV_X1 U8572 ( .A(n8542), .ZN(n8541) );
  NOR2_X1 U8573 ( .A1(n8543), .A2(n8544), .ZN(n8540) );
  XOR2_X1 U8574 ( .A(n8545), .B(n8546), .Z(Result_mul_12_) );
  XOR2_X1 U8575 ( .A(n8547), .B(n8548), .Z(Result_mul_11_) );
  NOR2_X1 U8576 ( .A1(n8549), .A2(n8550), .ZN(n8548) );
  INV_X1 U8577 ( .A(n8551), .ZN(n8550) );
  NOR2_X1 U8578 ( .A1(n8552), .A2(n8553), .ZN(n8549) );
  XOR2_X1 U8579 ( .A(n8554), .B(n8555), .Z(Result_mul_10_) );
  NAND3_X1 U8580 ( .A1(n8556), .A2(n8509), .A3(n8557), .ZN(Result_mul_0_) );
  INV_X1 U8581 ( .A(n8558), .ZN(n8557) );
  NOR2_X1 U8582 ( .A1(n8457), .A2(n8559), .ZN(n8558) );
  NAND4_X1 U8583 ( .A1(n8559), .A2(n8560), .A3(n8561), .A4(n8562), .ZN(n8509)
         );
  NAND2_X1 U8584 ( .A1(n8506), .A2(n8508), .ZN(n8556) );
  NAND2_X1 U8585 ( .A1(n8563), .A2(n8564), .ZN(n8508) );
  NAND2_X1 U8586 ( .A1(n8561), .A2(n8562), .ZN(n8564) );
  XOR2_X1 U8587 ( .A(n8560), .B(n8559), .Z(n8563) );
  NOR2_X1 U8588 ( .A1(n8565), .A2(n8566), .ZN(n8559) );
  NOR3_X1 U8589 ( .A1(n8567), .A2(n8568), .A3(n8569), .ZN(n8566) );
  NOR2_X1 U8590 ( .A1(n8570), .A2(n8571), .ZN(n8568) );
  INV_X1 U8591 ( .A(n8572), .ZN(n8565) );
  NAND2_X1 U8592 ( .A1(n8571), .A2(n8570), .ZN(n8572) );
  NOR2_X1 U8593 ( .A1(n8465), .A2(n8466), .ZN(n8506) );
  NOR2_X1 U8594 ( .A1(n8573), .A2(n8574), .ZN(n8466) );
  NAND2_X1 U8595 ( .A1(n8420), .A2(n8575), .ZN(n8573) );
  NAND2_X1 U8596 ( .A1(n8411), .A2(n8416), .ZN(n8575) );
  NOR2_X1 U8597 ( .A1(n8366), .A2(n8365), .ZN(n8411) );
  NOR2_X1 U8598 ( .A1(n8576), .A2(n8577), .ZN(n8365) );
  NAND2_X1 U8599 ( .A1(n8324), .A2(n8578), .ZN(n8576) );
  NAND2_X1 U8600 ( .A1(n8315), .A2(n8320), .ZN(n8578) );
  NOR2_X1 U8601 ( .A1(n8295), .A2(n8294), .ZN(n8315) );
  NOR2_X1 U8602 ( .A1(n8579), .A2(n8580), .ZN(n8294) );
  NAND2_X1 U8603 ( .A1(n8293), .A2(n8581), .ZN(n8579) );
  NAND2_X1 U8604 ( .A1(n8284), .A2(n8289), .ZN(n8581) );
  NOR2_X1 U8605 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  NOR2_X1 U8606 ( .A1(n8582), .A2(n8583), .ZN(n8282) );
  NAND2_X1 U8607 ( .A1(n8281), .A2(n8584), .ZN(n8582) );
  NAND2_X1 U8608 ( .A1(n8272), .A2(n8277), .ZN(n8584) );
  NOR2_X1 U8609 ( .A1(n8554), .A2(n8555), .ZN(n8272) );
  NOR2_X1 U8610 ( .A1(n8585), .A2(n8586), .ZN(n8555) );
  NAND2_X1 U8611 ( .A1(n8551), .A2(n8587), .ZN(n8586) );
  NAND2_X1 U8612 ( .A1(n8552), .A2(n8547), .ZN(n8587) );
  NOR2_X1 U8613 ( .A1(n8546), .A2(n8545), .ZN(n8547) );
  NOR2_X1 U8614 ( .A1(n8588), .A2(n8589), .ZN(n8545) );
  NAND2_X1 U8615 ( .A1(n8542), .A2(n8590), .ZN(n8589) );
  NAND2_X1 U8616 ( .A1(n8543), .A2(n8538), .ZN(n8590) );
  NOR2_X1 U8617 ( .A1(n8536), .A2(n8537), .ZN(n8538) );
  NOR2_X1 U8618 ( .A1(n8591), .A2(n8592), .ZN(n8537) );
  NAND2_X1 U8619 ( .A1(n8535), .A2(n8593), .ZN(n8592) );
  NAND2_X1 U8620 ( .A1(n8534), .A2(n8532), .ZN(n8593) );
  NAND2_X1 U8621 ( .A1(n8594), .A2(n8530), .ZN(n8532) );
  NAND2_X1 U8622 ( .A1(n8595), .A2(n8596), .ZN(n8530) );
  NAND2_X1 U8623 ( .A1(n8531), .A2(n8528), .ZN(n8594) );
  NAND2_X1 U8624 ( .A1(n8522), .A2(n8597), .ZN(n8528) );
  NAND2_X1 U8625 ( .A1(n8523), .A2(n8518), .ZN(n8597) );
  NAND2_X1 U8626 ( .A1(n8598), .A2(n8516), .ZN(n8518) );
  NAND2_X1 U8627 ( .A1(n8599), .A2(n8600), .ZN(n8516) );
  NAND2_X1 U8628 ( .A1(n8514), .A2(n8517), .ZN(n8598) );
  INV_X1 U8629 ( .A(n8601), .ZN(n8517) );
  NOR2_X1 U8630 ( .A1(n8599), .A2(n8600), .ZN(n8601) );
  XOR2_X1 U8631 ( .A(n8526), .B(n8527), .Z(n8599) );
  NAND2_X1 U8632 ( .A1(n8602), .A2(n8603), .ZN(n8514) );
  NAND2_X1 U8633 ( .A1(n8510), .A2(n8604), .ZN(n8603) );
  INV_X1 U8634 ( .A(n8513), .ZN(n8604) );
  NOR2_X1 U8635 ( .A1(n8605), .A2(n8606), .ZN(n8513) );
  NOR2_X1 U8636 ( .A1(n8607), .A2(n8600), .ZN(n8606) );
  NOR2_X1 U8637 ( .A1(n8608), .A2(n8609), .ZN(n8605) );
  NAND2_X1 U8638 ( .A1(n8504), .A2(n8610), .ZN(n8510) );
  NAND2_X1 U8639 ( .A1(n8502), .A2(n8505), .ZN(n8610) );
  NAND2_X1 U8640 ( .A1(n8611), .A2(n8612), .ZN(n8505) );
  NAND2_X1 U8641 ( .A1(n8613), .A2(n8614), .ZN(n8612) );
  XNOR2_X1 U8642 ( .A(n8609), .B(n8608), .ZN(n8611) );
  NAND2_X1 U8643 ( .A1(n8500), .A2(n8615), .ZN(n8502) );
  NAND2_X1 U8644 ( .A1(n8501), .A2(n8498), .ZN(n8615) );
  NAND2_X1 U8645 ( .A1(n8616), .A2(n8496), .ZN(n8498) );
  NAND2_X1 U8646 ( .A1(n8617), .A2(n8618), .ZN(n8496) );
  INV_X1 U8647 ( .A(n8619), .ZN(n8617) );
  NAND2_X1 U8648 ( .A1(n8494), .A2(n8497), .ZN(n8616) );
  NAND2_X1 U8649 ( .A1(n8619), .A2(n8620), .ZN(n8497) );
  XNOR2_X1 U8650 ( .A(n8621), .B(n8622), .ZN(n8619) );
  NAND2_X1 U8651 ( .A1(n8492), .A2(n8623), .ZN(n8494) );
  NAND2_X1 U8652 ( .A1(n8490), .A2(n8493), .ZN(n8623) );
  NAND2_X1 U8653 ( .A1(n8624), .A2(n8625), .ZN(n8493) );
  NAND2_X1 U8654 ( .A1(n8626), .A2(n8627), .ZN(n8625) );
  NAND2_X1 U8655 ( .A1(n8488), .A2(n8628), .ZN(n8490) );
  NAND2_X1 U8656 ( .A1(n8486), .A2(n8489), .ZN(n8628) );
  NAND2_X1 U8657 ( .A1(n8629), .A2(n8630), .ZN(n8489) );
  NAND2_X1 U8658 ( .A1(n8484), .A2(n8631), .ZN(n8486) );
  NAND2_X1 U8659 ( .A1(n8485), .A2(n8482), .ZN(n8631) );
  NAND2_X1 U8660 ( .A1(n8632), .A2(n8480), .ZN(n8482) );
  NAND2_X1 U8661 ( .A1(n8633), .A2(n8634), .ZN(n8480) );
  INV_X1 U8662 ( .A(n8635), .ZN(n8633) );
  NAND2_X1 U8663 ( .A1(n8478), .A2(n8481), .ZN(n8632) );
  NAND2_X1 U8664 ( .A1(n8635), .A2(n8636), .ZN(n8481) );
  XNOR2_X1 U8665 ( .A(n8637), .B(n8638), .ZN(n8635) );
  NAND2_X1 U8666 ( .A1(n8476), .A2(n8639), .ZN(n8478) );
  NAND2_X1 U8667 ( .A1(n8474), .A2(n8477), .ZN(n8639) );
  NAND2_X1 U8668 ( .A1(n8640), .A2(n8641), .ZN(n8477) );
  NAND2_X1 U8669 ( .A1(n8472), .A2(n8642), .ZN(n8474) );
  NAND2_X1 U8670 ( .A1(n8470), .A2(n8473), .ZN(n8642) );
  NAND2_X1 U8671 ( .A1(n8643), .A2(n8644), .ZN(n8473) );
  NAND2_X1 U8672 ( .A1(n8645), .A2(n8646), .ZN(n8644) );
  XNOR2_X1 U8673 ( .A(n8647), .B(n8648), .ZN(n8643) );
  NAND2_X1 U8674 ( .A1(n8469), .A2(n8649), .ZN(n8470) );
  NAND2_X1 U8675 ( .A1(n8460), .A2(n8468), .ZN(n8649) );
  NAND2_X1 U8676 ( .A1(n8650), .A2(n8651), .ZN(n8468) );
  NAND2_X1 U8677 ( .A1(n8652), .A2(n8653), .ZN(n8651) );
  XNOR2_X1 U8678 ( .A(n8646), .B(n8645), .ZN(n8650) );
  NOR3_X1 U8679 ( .A1(n8464), .A2(n8459), .A3(n8458), .ZN(n8460) );
  XOR2_X1 U8680 ( .A(n8654), .B(n8655), .Z(n8458) );
  XOR2_X1 U8681 ( .A(n8656), .B(n8657), .Z(n8655) );
  NAND2_X1 U8682 ( .A1(b_30_), .A2(a_0_), .ZN(n8657) );
  NOR2_X1 U8683 ( .A1(n8658), .A2(n8659), .ZN(n8459) );
  NOR3_X1 U8684 ( .A1(n8457), .A2(n8660), .A3(n8301), .ZN(n8659) );
  INV_X1 U8685 ( .A(n8661), .ZN(n8660) );
  NAND2_X1 U8686 ( .A1(n8455), .A2(n8454), .ZN(n8661) );
  NOR2_X1 U8687 ( .A1(n8454), .A2(n8455), .ZN(n8658) );
  NOR2_X1 U8688 ( .A1(n8662), .A2(n8663), .ZN(n8455) );
  INV_X1 U8689 ( .A(n8664), .ZN(n8663) );
  NAND3_X1 U8690 ( .A1(a_1_), .A2(n8665), .A3(b_31_), .ZN(n8664) );
  NAND2_X1 U8691 ( .A1(n8451), .A2(n8449), .ZN(n8665) );
  NOR2_X1 U8692 ( .A1(n8449), .A2(n8451), .ZN(n8662) );
  NOR2_X1 U8693 ( .A1(n8666), .A2(n8667), .ZN(n8451) );
  NOR3_X1 U8694 ( .A1(n8448), .A2(n8668), .A3(n8301), .ZN(n8667) );
  NOR2_X1 U8695 ( .A1(n8446), .A2(n8445), .ZN(n8668) );
  INV_X1 U8696 ( .A(n8669), .ZN(n8666) );
  NAND2_X1 U8697 ( .A1(n8445), .A2(n8446), .ZN(n8669) );
  NAND2_X1 U8698 ( .A1(n8670), .A2(n8671), .ZN(n8446) );
  NAND3_X1 U8699 ( .A1(a_3_), .A2(n8672), .A3(b_31_), .ZN(n8671) );
  NAND2_X1 U8700 ( .A1(n8442), .A2(n8440), .ZN(n8672) );
  INV_X1 U8701 ( .A(n8673), .ZN(n8670) );
  NOR2_X1 U8702 ( .A1(n8440), .A2(n8442), .ZN(n8673) );
  NOR2_X1 U8703 ( .A1(n8674), .A2(n8675), .ZN(n8442) );
  INV_X1 U8704 ( .A(n8676), .ZN(n8675) );
  NAND3_X1 U8705 ( .A1(a_4_), .A2(n8677), .A3(b_31_), .ZN(n8676) );
  NAND2_X1 U8706 ( .A1(n8437), .A2(n8436), .ZN(n8677) );
  NOR2_X1 U8707 ( .A1(n8436), .A2(n8437), .ZN(n8674) );
  NOR2_X1 U8708 ( .A1(n8678), .A2(n8679), .ZN(n8437) );
  INV_X1 U8709 ( .A(n8680), .ZN(n8679) );
  NAND3_X1 U8710 ( .A1(a_5_), .A2(n8681), .A3(b_31_), .ZN(n8680) );
  NAND2_X1 U8711 ( .A1(n8433), .A2(n8431), .ZN(n8681) );
  NOR2_X1 U8712 ( .A1(n8431), .A2(n8433), .ZN(n8678) );
  NOR2_X1 U8713 ( .A1(n8682), .A2(n8683), .ZN(n8433) );
  NOR3_X1 U8714 ( .A1(n8430), .A2(n8684), .A3(n8301), .ZN(n8683) );
  NOR2_X1 U8715 ( .A1(n8428), .A2(n8427), .ZN(n8684) );
  INV_X1 U8716 ( .A(n8685), .ZN(n8682) );
  NAND2_X1 U8717 ( .A1(n8427), .A2(n8428), .ZN(n8685) );
  NAND2_X1 U8718 ( .A1(n8686), .A2(n8687), .ZN(n8428) );
  NAND3_X1 U8719 ( .A1(a_7_), .A2(n8688), .A3(b_31_), .ZN(n8687) );
  INV_X1 U8720 ( .A(n8689), .ZN(n8688) );
  NOR2_X1 U8721 ( .A1(n8423), .A2(n8422), .ZN(n8689) );
  NAND2_X1 U8722 ( .A1(n8422), .A2(n8423), .ZN(n8686) );
  NAND2_X1 U8723 ( .A1(n8690), .A2(n8691), .ZN(n8423) );
  NAND3_X1 U8724 ( .A1(a_8_), .A2(n8692), .A3(b_31_), .ZN(n8691) );
  NAND2_X1 U8725 ( .A1(n8409), .A2(n8407), .ZN(n8692) );
  INV_X1 U8726 ( .A(n8693), .ZN(n8690) );
  NOR2_X1 U8727 ( .A1(n8407), .A2(n8409), .ZN(n8693) );
  NOR2_X1 U8728 ( .A1(n8694), .A2(n8695), .ZN(n8409) );
  INV_X1 U8729 ( .A(n8696), .ZN(n8695) );
  NAND3_X1 U8730 ( .A1(a_9_), .A2(n8697), .A3(b_31_), .ZN(n8696) );
  NAND2_X1 U8731 ( .A1(n8405), .A2(n8403), .ZN(n8697) );
  NOR2_X1 U8732 ( .A1(n8403), .A2(n8405), .ZN(n8694) );
  NOR2_X1 U8733 ( .A1(n8698), .A2(n8699), .ZN(n8405) );
  NOR3_X1 U8734 ( .A1(n8402), .A2(n8700), .A3(n8301), .ZN(n8699) );
  INV_X1 U8735 ( .A(n8701), .ZN(n8700) );
  NAND2_X1 U8736 ( .A1(n8400), .A2(n8399), .ZN(n8701) );
  NOR2_X1 U8737 ( .A1(n8399), .A2(n8400), .ZN(n8698) );
  NOR2_X1 U8738 ( .A1(n8702), .A2(n8703), .ZN(n8400) );
  INV_X1 U8739 ( .A(n8704), .ZN(n8703) );
  NAND3_X1 U8740 ( .A1(a_11_), .A2(n8705), .A3(b_31_), .ZN(n8704) );
  NAND2_X1 U8741 ( .A1(n8396), .A2(n8394), .ZN(n8705) );
  NOR2_X1 U8742 ( .A1(n8394), .A2(n8396), .ZN(n8702) );
  NOR2_X1 U8743 ( .A1(n8706), .A2(n8707), .ZN(n8396) );
  NOR3_X1 U8744 ( .A1(n8393), .A2(n8708), .A3(n8301), .ZN(n8707) );
  NOR2_X1 U8745 ( .A1(n8391), .A2(n8390), .ZN(n8708) );
  INV_X1 U8746 ( .A(n8709), .ZN(n8706) );
  NAND2_X1 U8747 ( .A1(n8390), .A2(n8391), .ZN(n8709) );
  NAND2_X1 U8748 ( .A1(n8710), .A2(n8711), .ZN(n8391) );
  NAND3_X1 U8749 ( .A1(a_13_), .A2(n8712), .A3(b_31_), .ZN(n8711) );
  NAND2_X1 U8750 ( .A1(n8387), .A2(n8385), .ZN(n8712) );
  INV_X1 U8751 ( .A(n8713), .ZN(n8710) );
  NOR2_X1 U8752 ( .A1(n8385), .A2(n8387), .ZN(n8713) );
  NOR2_X1 U8753 ( .A1(n8714), .A2(n8715), .ZN(n8387) );
  INV_X1 U8754 ( .A(n8716), .ZN(n8715) );
  NAND3_X1 U8755 ( .A1(a_14_), .A2(n8717), .A3(b_31_), .ZN(n8716) );
  NAND2_X1 U8756 ( .A1(n8383), .A2(n8381), .ZN(n8717) );
  NOR2_X1 U8757 ( .A1(n8381), .A2(n8383), .ZN(n8714) );
  NOR2_X1 U8758 ( .A1(n8718), .A2(n8719), .ZN(n8383) );
  INV_X1 U8759 ( .A(n8720), .ZN(n8719) );
  NAND3_X1 U8760 ( .A1(a_15_), .A2(n8721), .A3(b_31_), .ZN(n8720) );
  NAND2_X1 U8761 ( .A1(n8379), .A2(n8377), .ZN(n8721) );
  NOR2_X1 U8762 ( .A1(n8377), .A2(n8379), .ZN(n8718) );
  NOR2_X1 U8763 ( .A1(n8722), .A2(n8723), .ZN(n8379) );
  NOR3_X1 U8764 ( .A1(n8376), .A2(n8724), .A3(n8301), .ZN(n8723) );
  INV_X1 U8765 ( .A(n8725), .ZN(n8724) );
  NAND2_X1 U8766 ( .A1(n8374), .A2(n8373), .ZN(n8725) );
  NOR2_X1 U8767 ( .A1(n8373), .A2(n8374), .ZN(n8722) );
  NOR2_X1 U8768 ( .A1(n8726), .A2(n8727), .ZN(n8374) );
  NOR3_X1 U8769 ( .A1(n8371), .A2(n8728), .A3(n8301), .ZN(n8727) );
  NOR2_X1 U8770 ( .A1(n8369), .A2(n8368), .ZN(n8728) );
  INV_X1 U8771 ( .A(n8729), .ZN(n8726) );
  NAND2_X1 U8772 ( .A1(n8368), .A2(n8369), .ZN(n8729) );
  NAND2_X1 U8773 ( .A1(n8730), .A2(n8731), .ZN(n8369) );
  NAND3_X1 U8774 ( .A1(a_18_), .A2(n8732), .A3(b_31_), .ZN(n8731) );
  INV_X1 U8775 ( .A(n8733), .ZN(n8732) );
  NOR2_X1 U8776 ( .A1(n8363), .A2(n8361), .ZN(n8733) );
  NAND2_X1 U8777 ( .A1(n8361), .A2(n8363), .ZN(n8730) );
  NAND2_X1 U8778 ( .A1(n8359), .A2(n8734), .ZN(n8363) );
  NAND2_X1 U8779 ( .A1(n8358), .A2(n8360), .ZN(n8734) );
  NAND2_X1 U8780 ( .A1(n8735), .A2(n8736), .ZN(n8360) );
  NAND2_X1 U8781 ( .A1(b_31_), .A2(a_19_), .ZN(n8735) );
  XNOR2_X1 U8782 ( .A(n8737), .B(n8738), .ZN(n8358) );
  NAND2_X1 U8783 ( .A1(n8739), .A2(n8740), .ZN(n8737) );
  INV_X1 U8784 ( .A(n8741), .ZN(n8359) );
  NOR2_X1 U8785 ( .A1(n8736), .A2(n8742), .ZN(n8741) );
  NAND2_X1 U8786 ( .A1(n8743), .A2(n8744), .ZN(n8736) );
  NAND2_X1 U8787 ( .A1(n8745), .A2(n8355), .ZN(n8744) );
  NAND2_X1 U8788 ( .A1(b_31_), .A2(a_20_), .ZN(n8355) );
  NAND2_X1 U8789 ( .A1(n8353), .A2(n8356), .ZN(n8745) );
  INV_X1 U8790 ( .A(n8746), .ZN(n8743) );
  NOR2_X1 U8791 ( .A1(n8356), .A2(n8353), .ZN(n8746) );
  XNOR2_X1 U8792 ( .A(n8747), .B(n8748), .ZN(n8353) );
  XOR2_X1 U8793 ( .A(n8749), .B(n8750), .Z(n8748) );
  NAND2_X1 U8794 ( .A1(b_30_), .A2(a_21_), .ZN(n8750) );
  NAND2_X1 U8795 ( .A1(n8351), .A2(n8751), .ZN(n8356) );
  NAND2_X1 U8796 ( .A1(n8350), .A2(n8352), .ZN(n8751) );
  NAND2_X1 U8797 ( .A1(n8752), .A2(n8753), .ZN(n8352) );
  NAND2_X1 U8798 ( .A1(b_31_), .A2(a_21_), .ZN(n8752) );
  XNOR2_X1 U8799 ( .A(n8754), .B(n8755), .ZN(n8350) );
  NAND2_X1 U8800 ( .A1(n8756), .A2(n8757), .ZN(n8754) );
  INV_X1 U8801 ( .A(n8758), .ZN(n8351) );
  NOR2_X1 U8802 ( .A1(n8753), .A2(n8759), .ZN(n8758) );
  NAND2_X1 U8803 ( .A1(n8760), .A2(n8761), .ZN(n8753) );
  NAND2_X1 U8804 ( .A1(n8762), .A2(n8348), .ZN(n8761) );
  NAND2_X1 U8805 ( .A1(b_31_), .A2(a_22_), .ZN(n8348) );
  NAND2_X1 U8806 ( .A1(n8346), .A2(n8347), .ZN(n8762) );
  INV_X1 U8807 ( .A(n8763), .ZN(n8760) );
  NOR2_X1 U8808 ( .A1(n8347), .A2(n8346), .ZN(n8763) );
  XNOR2_X1 U8809 ( .A(n8764), .B(n8765), .ZN(n8346) );
  NAND2_X1 U8810 ( .A1(n8766), .A2(n8767), .ZN(n8764) );
  NAND2_X1 U8811 ( .A1(n8343), .A2(n8768), .ZN(n8347) );
  NAND2_X1 U8812 ( .A1(n8342), .A2(n8344), .ZN(n8768) );
  NAND2_X1 U8813 ( .A1(n8769), .A2(n8770), .ZN(n8344) );
  INV_X1 U8814 ( .A(n8771), .ZN(n8770) );
  NAND2_X1 U8815 ( .A1(b_31_), .A2(a_23_), .ZN(n8769) );
  XNOR2_X1 U8816 ( .A(n8772), .B(n8773), .ZN(n8342) );
  XNOR2_X1 U8817 ( .A(n8774), .B(n8775), .ZN(n8772) );
  NAND2_X1 U8818 ( .A1(n8771), .A2(a_23_), .ZN(n8343) );
  NOR2_X1 U8819 ( .A1(n8776), .A2(n8777), .ZN(n8771) );
  NOR2_X1 U8820 ( .A1(n8778), .A2(n8339), .ZN(n8777) );
  NOR2_X1 U8821 ( .A1(n8301), .A2(n8779), .ZN(n8339) );
  INV_X1 U8822 ( .A(n8780), .ZN(n8778) );
  NAND2_X1 U8823 ( .A1(n8337), .A2(n8340), .ZN(n8780) );
  NOR2_X1 U8824 ( .A1(n8340), .A2(n8337), .ZN(n8776) );
  XOR2_X1 U8825 ( .A(n8781), .B(n8782), .Z(n8337) );
  XOR2_X1 U8826 ( .A(n8783), .B(n8784), .Z(n8781) );
  NAND2_X1 U8827 ( .A1(n8785), .A2(n8786), .ZN(n8340) );
  NAND2_X1 U8828 ( .A1(n8336), .A2(n8787), .ZN(n8786) );
  NAND2_X1 U8829 ( .A1(n8335), .A2(n8334), .ZN(n8787) );
  NOR2_X1 U8830 ( .A1(n8301), .A2(n8788), .ZN(n8336) );
  INV_X1 U8831 ( .A(n8789), .ZN(n8785) );
  NOR2_X1 U8832 ( .A1(n8334), .A2(n8335), .ZN(n8789) );
  NOR2_X1 U8833 ( .A1(n8790), .A2(n8791), .ZN(n8335) );
  NOR2_X1 U8834 ( .A1(n8331), .A2(n8792), .ZN(n8791) );
  NOR2_X1 U8835 ( .A1(n8332), .A2(n8329), .ZN(n8792) );
  NAND2_X1 U8836 ( .A1(b_31_), .A2(a_26_), .ZN(n8331) );
  INV_X1 U8837 ( .A(n8793), .ZN(n8790) );
  NAND2_X1 U8838 ( .A1(n8329), .A2(n8332), .ZN(n8793) );
  NAND2_X1 U8839 ( .A1(n8794), .A2(n8795), .ZN(n8332) );
  NAND2_X1 U8840 ( .A1(n8328), .A2(n8796), .ZN(n8795) );
  NAND2_X1 U8841 ( .A1(n8327), .A2(n8326), .ZN(n8796) );
  NOR2_X1 U8842 ( .A1(n8301), .A2(n8797), .ZN(n8328) );
  INV_X1 U8843 ( .A(n8798), .ZN(n8794) );
  NOR2_X1 U8844 ( .A1(n8326), .A2(n8327), .ZN(n8798) );
  NOR2_X1 U8845 ( .A1(n8799), .A2(n8800), .ZN(n8327) );
  NOR3_X1 U8846 ( .A1(n8314), .A2(n8801), .A3(n8301), .ZN(n8800) );
  INV_X1 U8847 ( .A(n8802), .ZN(n8801) );
  NAND2_X1 U8848 ( .A1(n8311), .A2(n8312), .ZN(n8802) );
  NOR2_X1 U8849 ( .A1(n8312), .A2(n8311), .ZN(n8799) );
  XNOR2_X1 U8850 ( .A(n8803), .B(n8804), .ZN(n8311) );
  XNOR2_X1 U8851 ( .A(n8805), .B(n8806), .ZN(n8803) );
  NAND2_X1 U8852 ( .A1(n8807), .A2(n8808), .ZN(n8312) );
  NAND2_X1 U8853 ( .A1(n8809), .A2(n8308), .ZN(n8808) );
  NAND2_X1 U8854 ( .A1(b_31_), .A2(a_29_), .ZN(n8308) );
  NAND2_X1 U8855 ( .A1(n8306), .A2(n8309), .ZN(n8809) );
  INV_X1 U8856 ( .A(n8810), .ZN(n8807) );
  NOR2_X1 U8857 ( .A1(n8309), .A2(n8306), .ZN(n8810) );
  NAND2_X1 U8858 ( .A1(n8811), .A2(n8812), .ZN(n8309) );
  NAND2_X1 U8859 ( .A1(b_29_), .A2(n8813), .ZN(n8812) );
  NAND2_X1 U8860 ( .A1(n8299), .A2(n8814), .ZN(n8813) );
  NAND2_X1 U8861 ( .A1(a_31_), .A2(n8305), .ZN(n8814) );
  NAND2_X1 U8862 ( .A1(b_30_), .A2(n8815), .ZN(n8811) );
  NAND2_X1 U8863 ( .A1(n8303), .A2(n8816), .ZN(n8815) );
  NAND2_X1 U8864 ( .A1(a_30_), .A2(n8817), .ZN(n8816) );
  XOR2_X1 U8865 ( .A(n8818), .B(n8819), .Z(n8326) );
  XNOR2_X1 U8866 ( .A(n8820), .B(n8821), .ZN(n8818) );
  XNOR2_X1 U8867 ( .A(n8822), .B(n8823), .ZN(n8329) );
  XNOR2_X1 U8868 ( .A(n8824), .B(n8825), .ZN(n8822) );
  NOR2_X1 U8869 ( .A1(n8797), .A2(n8305), .ZN(n8825) );
  XNOR2_X1 U8870 ( .A(n8826), .B(n8827), .ZN(n8334) );
  XNOR2_X1 U8871 ( .A(n8828), .B(n8829), .ZN(n8827) );
  XNOR2_X1 U8872 ( .A(n8830), .B(n8831), .ZN(n8361) );
  XOR2_X1 U8873 ( .A(n8832), .B(n8833), .Z(n8831) );
  NAND2_X1 U8874 ( .A1(b_30_), .A2(a_19_), .ZN(n8833) );
  XOR2_X1 U8875 ( .A(n8834), .B(n8835), .Z(n8368) );
  XNOR2_X1 U8876 ( .A(n8836), .B(n8837), .ZN(n8835) );
  XOR2_X1 U8877 ( .A(n8838), .B(n8839), .Z(n8373) );
  XOR2_X1 U8878 ( .A(n8840), .B(n8841), .Z(n8839) );
  NAND2_X1 U8879 ( .A1(b_30_), .A2(a_17_), .ZN(n8841) );
  XOR2_X1 U8880 ( .A(n8842), .B(n8843), .Z(n8377) );
  NAND2_X1 U8881 ( .A1(n8844), .A2(n8845), .ZN(n8842) );
  XNOR2_X1 U8882 ( .A(n8846), .B(n8847), .ZN(n8381) );
  XOR2_X1 U8883 ( .A(n8848), .B(n8849), .Z(n8846) );
  NOR2_X1 U8884 ( .A1(n8850), .A2(n8305), .ZN(n8849) );
  XOR2_X1 U8885 ( .A(n8851), .B(n8852), .Z(n8385) );
  NAND2_X1 U8886 ( .A1(n8853), .A2(n8854), .ZN(n8851) );
  XNOR2_X1 U8887 ( .A(n8855), .B(n8856), .ZN(n8390) );
  XOR2_X1 U8888 ( .A(n8857), .B(n8858), .Z(n8856) );
  NAND2_X1 U8889 ( .A1(b_30_), .A2(a_13_), .ZN(n8858) );
  XOR2_X1 U8890 ( .A(n8859), .B(n8860), .Z(n8394) );
  NAND2_X1 U8891 ( .A1(n8861), .A2(n8862), .ZN(n8859) );
  XNOR2_X1 U8892 ( .A(n8863), .B(n8864), .ZN(n8399) );
  XOR2_X1 U8893 ( .A(n8865), .B(n8866), .Z(n8863) );
  NOR2_X1 U8894 ( .A1(n8867), .A2(n8305), .ZN(n8866) );
  XOR2_X1 U8895 ( .A(n8868), .B(n8869), .Z(n8403) );
  NAND2_X1 U8896 ( .A1(n8870), .A2(n8871), .ZN(n8868) );
  XOR2_X1 U8897 ( .A(n8872), .B(n8873), .Z(n8407) );
  XOR2_X1 U8898 ( .A(n8874), .B(n8875), .Z(n8873) );
  NAND2_X1 U8899 ( .A1(b_30_), .A2(a_9_), .ZN(n8875) );
  XNOR2_X1 U8900 ( .A(n8876), .B(n8877), .ZN(n8422) );
  NAND2_X1 U8901 ( .A1(n8878), .A2(n8879), .ZN(n8876) );
  XOR2_X1 U8902 ( .A(n8880), .B(n8881), .Z(n8427) );
  XOR2_X1 U8903 ( .A(n8882), .B(n8883), .Z(n8880) );
  NOR2_X1 U8904 ( .A1(n8425), .A2(n8305), .ZN(n8883) );
  XNOR2_X1 U8905 ( .A(n8884), .B(n8885), .ZN(n8431) );
  XNOR2_X1 U8906 ( .A(n8886), .B(n8887), .ZN(n8885) );
  XOR2_X1 U8907 ( .A(n8888), .B(n8889), .Z(n8436) );
  XOR2_X1 U8908 ( .A(n8890), .B(n8891), .Z(n8889) );
  NAND2_X1 U8909 ( .A1(b_30_), .A2(a_5_), .ZN(n8891) );
  XOR2_X1 U8910 ( .A(n8892), .B(n8893), .Z(n8440) );
  NAND2_X1 U8911 ( .A1(n8894), .A2(n8895), .ZN(n8892) );
  XOR2_X1 U8912 ( .A(n8896), .B(n8897), .Z(n8445) );
  XOR2_X1 U8913 ( .A(n8898), .B(n8899), .Z(n8896) );
  NOR2_X1 U8914 ( .A1(n8900), .A2(n8305), .ZN(n8899) );
  XOR2_X1 U8915 ( .A(n8901), .B(n8902), .Z(n8449) );
  NAND2_X1 U8916 ( .A1(n8903), .A2(n8904), .ZN(n8901) );
  XNOR2_X1 U8917 ( .A(n8905), .B(n8906), .ZN(n8454) );
  XOR2_X1 U8918 ( .A(n8907), .B(n8908), .Z(n8905) );
  NOR2_X1 U8919 ( .A1(n8569), .A2(n8305), .ZN(n8908) );
  XNOR2_X1 U8920 ( .A(n8653), .B(n8652), .ZN(n8464) );
  NAND3_X1 U8921 ( .A1(n8652), .A2(n8653), .A3(n8909), .ZN(n8469) );
  XNOR2_X1 U8922 ( .A(n8646), .B(n8910), .ZN(n8909) );
  INV_X1 U8923 ( .A(n8645), .ZN(n8910) );
  NAND2_X1 U8924 ( .A1(n8911), .A2(n8912), .ZN(n8653) );
  NAND3_X1 U8925 ( .A1(a_0_), .A2(n8913), .A3(b_30_), .ZN(n8912) );
  INV_X1 U8926 ( .A(n8914), .ZN(n8913) );
  NOR2_X1 U8927 ( .A1(n8656), .A2(n8654), .ZN(n8914) );
  NAND2_X1 U8928 ( .A1(n8654), .A2(n8656), .ZN(n8911) );
  NAND2_X1 U8929 ( .A1(n8915), .A2(n8916), .ZN(n8656) );
  INV_X1 U8930 ( .A(n8917), .ZN(n8916) );
  NOR3_X1 U8931 ( .A1(n8569), .A2(n8918), .A3(n8305), .ZN(n8917) );
  NOR2_X1 U8932 ( .A1(n8907), .A2(n8906), .ZN(n8918) );
  NAND2_X1 U8933 ( .A1(n8906), .A2(n8907), .ZN(n8915) );
  NAND2_X1 U8934 ( .A1(n8903), .A2(n8919), .ZN(n8907) );
  NAND2_X1 U8935 ( .A1(n8902), .A2(n8904), .ZN(n8919) );
  NAND2_X1 U8936 ( .A1(n8920), .A2(n8921), .ZN(n8904) );
  NAND2_X1 U8937 ( .A1(b_30_), .A2(a_2_), .ZN(n8921) );
  XNOR2_X1 U8938 ( .A(n8922), .B(n8923), .ZN(n8902) );
  XOR2_X1 U8939 ( .A(n8924), .B(n8925), .Z(n8923) );
  NAND2_X1 U8940 ( .A1(b_29_), .A2(a_3_), .ZN(n8925) );
  INV_X1 U8941 ( .A(n8926), .ZN(n8903) );
  NOR2_X1 U8942 ( .A1(n8448), .A2(n8920), .ZN(n8926) );
  NOR2_X1 U8943 ( .A1(n8927), .A2(n8928), .ZN(n8920) );
  NOR3_X1 U8944 ( .A1(n8900), .A2(n8929), .A3(n8305), .ZN(n8928) );
  NOR2_X1 U8945 ( .A1(n8898), .A2(n8897), .ZN(n8929) );
  INV_X1 U8946 ( .A(n8930), .ZN(n8927) );
  NAND2_X1 U8947 ( .A1(n8897), .A2(n8898), .ZN(n8930) );
  NAND2_X1 U8948 ( .A1(n8894), .A2(n8931), .ZN(n8898) );
  NAND2_X1 U8949 ( .A1(n8893), .A2(n8895), .ZN(n8931) );
  NAND2_X1 U8950 ( .A1(n8932), .A2(n8933), .ZN(n8895) );
  NAND2_X1 U8951 ( .A1(b_30_), .A2(a_4_), .ZN(n8933) );
  XNOR2_X1 U8952 ( .A(n8934), .B(n8935), .ZN(n8893) );
  XNOR2_X1 U8953 ( .A(n8936), .B(n8937), .ZN(n8935) );
  NOR2_X1 U8954 ( .A1(n8938), .A2(n8817), .ZN(n8937) );
  NAND2_X1 U8955 ( .A1(a_4_), .A2(n8939), .ZN(n8894) );
  INV_X1 U8956 ( .A(n8932), .ZN(n8939) );
  NOR2_X1 U8957 ( .A1(n8940), .A2(n8941), .ZN(n8932) );
  NOR3_X1 U8958 ( .A1(n8938), .A2(n8942), .A3(n8305), .ZN(n8941) );
  INV_X1 U8959 ( .A(n8943), .ZN(n8942) );
  NAND2_X1 U8960 ( .A1(n8888), .A2(n8890), .ZN(n8943) );
  NOR2_X1 U8961 ( .A1(n8890), .A2(n8888), .ZN(n8940) );
  XOR2_X1 U8962 ( .A(n8944), .B(n8945), .Z(n8888) );
  NAND2_X1 U8963 ( .A1(n8946), .A2(n8947), .ZN(n8944) );
  NAND2_X1 U8964 ( .A1(n8948), .A2(n8949), .ZN(n8890) );
  NAND2_X1 U8965 ( .A1(n8884), .A2(n8950), .ZN(n8949) );
  INV_X1 U8966 ( .A(n8951), .ZN(n8950) );
  NOR2_X1 U8967 ( .A1(n8887), .A2(n8886), .ZN(n8951) );
  XNOR2_X1 U8968 ( .A(n8952), .B(n8953), .ZN(n8884) );
  XNOR2_X1 U8969 ( .A(n8954), .B(n8955), .ZN(n8953) );
  NAND2_X1 U8970 ( .A1(b_29_), .A2(a_7_), .ZN(n8955) );
  NAND2_X1 U8971 ( .A1(n8886), .A2(n8887), .ZN(n8948) );
  NAND2_X1 U8972 ( .A1(b_30_), .A2(a_6_), .ZN(n8887) );
  NOR2_X1 U8973 ( .A1(n8956), .A2(n8957), .ZN(n8886) );
  NOR3_X1 U8974 ( .A1(n8425), .A2(n8958), .A3(n8305), .ZN(n8957) );
  NOR2_X1 U8975 ( .A1(n8882), .A2(n8881), .ZN(n8958) );
  INV_X1 U8976 ( .A(n8959), .ZN(n8956) );
  NAND2_X1 U8977 ( .A1(n8881), .A2(n8882), .ZN(n8959) );
  NAND2_X1 U8978 ( .A1(n8878), .A2(n8960), .ZN(n8882) );
  NAND2_X1 U8979 ( .A1(n8877), .A2(n8879), .ZN(n8960) );
  NAND2_X1 U8980 ( .A1(n8961), .A2(n8962), .ZN(n8879) );
  NAND2_X1 U8981 ( .A1(b_30_), .A2(a_8_), .ZN(n8962) );
  XNOR2_X1 U8982 ( .A(n8963), .B(n8964), .ZN(n8877) );
  XOR2_X1 U8983 ( .A(n8965), .B(n8966), .Z(n8964) );
  NAND2_X1 U8984 ( .A1(b_29_), .A2(a_9_), .ZN(n8966) );
  INV_X1 U8985 ( .A(n8967), .ZN(n8878) );
  NOR2_X1 U8986 ( .A1(n8968), .A2(n8961), .ZN(n8967) );
  NOR2_X1 U8987 ( .A1(n8969), .A2(n8970), .ZN(n8961) );
  NOR3_X1 U8988 ( .A1(n8971), .A2(n8972), .A3(n8305), .ZN(n8970) );
  NOR2_X1 U8989 ( .A1(n8874), .A2(n8872), .ZN(n8972) );
  INV_X1 U8990 ( .A(n8973), .ZN(n8969) );
  NAND2_X1 U8991 ( .A1(n8872), .A2(n8874), .ZN(n8973) );
  NAND2_X1 U8992 ( .A1(n8870), .A2(n8974), .ZN(n8874) );
  NAND2_X1 U8993 ( .A1(n8869), .A2(n8871), .ZN(n8974) );
  NAND2_X1 U8994 ( .A1(n8975), .A2(n8976), .ZN(n8871) );
  NAND2_X1 U8995 ( .A1(b_30_), .A2(a_10_), .ZN(n8976) );
  XOR2_X1 U8996 ( .A(n8977), .B(n8978), .Z(n8869) );
  XOR2_X1 U8997 ( .A(n8979), .B(n8980), .Z(n8977) );
  NOR2_X1 U8998 ( .A1(n8867), .A2(n8817), .ZN(n8980) );
  INV_X1 U8999 ( .A(n8981), .ZN(n8870) );
  NOR2_X1 U9000 ( .A1(n8402), .A2(n8975), .ZN(n8981) );
  NOR2_X1 U9001 ( .A1(n8982), .A2(n8983), .ZN(n8975) );
  NOR3_X1 U9002 ( .A1(n8867), .A2(n8984), .A3(n8305), .ZN(n8983) );
  NOR2_X1 U9003 ( .A1(n8865), .A2(n8864), .ZN(n8984) );
  INV_X1 U9004 ( .A(n8985), .ZN(n8982) );
  NAND2_X1 U9005 ( .A1(n8864), .A2(n8865), .ZN(n8985) );
  NAND2_X1 U9006 ( .A1(n8861), .A2(n8986), .ZN(n8865) );
  NAND2_X1 U9007 ( .A1(n8860), .A2(n8862), .ZN(n8986) );
  NAND2_X1 U9008 ( .A1(n8987), .A2(n8988), .ZN(n8862) );
  NAND2_X1 U9009 ( .A1(b_30_), .A2(a_12_), .ZN(n8988) );
  XNOR2_X1 U9010 ( .A(n8989), .B(n8990), .ZN(n8860) );
  XOR2_X1 U9011 ( .A(n8991), .B(n8992), .Z(n8990) );
  NAND2_X1 U9012 ( .A1(b_29_), .A2(a_13_), .ZN(n8992) );
  INV_X1 U9013 ( .A(n8993), .ZN(n8861) );
  NOR2_X1 U9014 ( .A1(n8393), .A2(n8987), .ZN(n8993) );
  NOR2_X1 U9015 ( .A1(n8994), .A2(n8995), .ZN(n8987) );
  NOR3_X1 U9016 ( .A1(n8996), .A2(n8997), .A3(n8305), .ZN(n8995) );
  NOR2_X1 U9017 ( .A1(n8857), .A2(n8855), .ZN(n8997) );
  INV_X1 U9018 ( .A(n8998), .ZN(n8994) );
  NAND2_X1 U9019 ( .A1(n8855), .A2(n8857), .ZN(n8998) );
  NAND2_X1 U9020 ( .A1(n8853), .A2(n8999), .ZN(n8857) );
  NAND2_X1 U9021 ( .A1(n8852), .A2(n8854), .ZN(n8999) );
  NAND2_X1 U9022 ( .A1(n9000), .A2(n9001), .ZN(n8854) );
  NAND2_X1 U9023 ( .A1(b_30_), .A2(a_14_), .ZN(n9001) );
  INV_X1 U9024 ( .A(n9002), .ZN(n9000) );
  XOR2_X1 U9025 ( .A(n9003), .B(n9004), .Z(n8852) );
  XOR2_X1 U9026 ( .A(n9005), .B(n9006), .Z(n9003) );
  NOR2_X1 U9027 ( .A1(n8850), .A2(n8817), .ZN(n9006) );
  NAND2_X1 U9028 ( .A1(a_14_), .A2(n9002), .ZN(n8853) );
  NAND2_X1 U9029 ( .A1(n9007), .A2(n9008), .ZN(n9002) );
  INV_X1 U9030 ( .A(n9009), .ZN(n9008) );
  NOR3_X1 U9031 ( .A1(n8850), .A2(n9010), .A3(n8305), .ZN(n9009) );
  NOR2_X1 U9032 ( .A1(n8847), .A2(n8848), .ZN(n9010) );
  NAND2_X1 U9033 ( .A1(n8847), .A2(n8848), .ZN(n9007) );
  NAND2_X1 U9034 ( .A1(n8844), .A2(n9011), .ZN(n8848) );
  NAND2_X1 U9035 ( .A1(n8843), .A2(n8845), .ZN(n9011) );
  NAND2_X1 U9036 ( .A1(n9012), .A2(n9013), .ZN(n8845) );
  NAND2_X1 U9037 ( .A1(b_30_), .A2(a_16_), .ZN(n9013) );
  XNOR2_X1 U9038 ( .A(n9014), .B(n9015), .ZN(n8843) );
  XOR2_X1 U9039 ( .A(n9016), .B(n9017), .Z(n9015) );
  NAND2_X1 U9040 ( .A1(b_29_), .A2(a_17_), .ZN(n9017) );
  NAND2_X1 U9041 ( .A1(a_16_), .A2(n9018), .ZN(n8844) );
  INV_X1 U9042 ( .A(n9012), .ZN(n9018) );
  NOR2_X1 U9043 ( .A1(n9019), .A2(n9020), .ZN(n9012) );
  NOR3_X1 U9044 ( .A1(n8371), .A2(n9021), .A3(n8305), .ZN(n9020) );
  INV_X1 U9045 ( .A(n9022), .ZN(n9021) );
  NAND2_X1 U9046 ( .A1(n8838), .A2(n8840), .ZN(n9022) );
  NOR2_X1 U9047 ( .A1(n8840), .A2(n8838), .ZN(n9019) );
  XOR2_X1 U9048 ( .A(n9023), .B(n9024), .Z(n8838) );
  XOR2_X1 U9049 ( .A(n9025), .B(n9026), .Z(n9023) );
  NAND2_X1 U9050 ( .A1(n9027), .A2(n9028), .ZN(n8840) );
  NAND2_X1 U9051 ( .A1(n8834), .A2(n9029), .ZN(n9028) );
  INV_X1 U9052 ( .A(n9030), .ZN(n9029) );
  NOR2_X1 U9053 ( .A1(n8837), .A2(n8836), .ZN(n9030) );
  XNOR2_X1 U9054 ( .A(n9031), .B(n9032), .ZN(n8834) );
  XOR2_X1 U9055 ( .A(n9033), .B(n9034), .Z(n9031) );
  NOR2_X1 U9056 ( .A1(n8742), .A2(n8817), .ZN(n9034) );
  NAND2_X1 U9057 ( .A1(n8836), .A2(n8837), .ZN(n9027) );
  NAND2_X1 U9058 ( .A1(b_30_), .A2(a_18_), .ZN(n8837) );
  NOR2_X1 U9059 ( .A1(n9035), .A2(n9036), .ZN(n8836) );
  NOR3_X1 U9060 ( .A1(n8742), .A2(n9037), .A3(n8305), .ZN(n9036) );
  NOR2_X1 U9061 ( .A1(n8832), .A2(n8830), .ZN(n9037) );
  INV_X1 U9062 ( .A(n9038), .ZN(n9035) );
  NAND2_X1 U9063 ( .A1(n8830), .A2(n8832), .ZN(n9038) );
  NAND2_X1 U9064 ( .A1(n8739), .A2(n9039), .ZN(n8832) );
  NAND2_X1 U9065 ( .A1(n8738), .A2(n8740), .ZN(n9039) );
  NAND2_X1 U9066 ( .A1(n9040), .A2(n9041), .ZN(n8740) );
  NAND2_X1 U9067 ( .A1(b_30_), .A2(a_20_), .ZN(n9041) );
  XOR2_X1 U9068 ( .A(n9042), .B(n9043), .Z(n8738) );
  XOR2_X1 U9069 ( .A(n9044), .B(n9045), .Z(n9042) );
  NOR2_X1 U9070 ( .A1(n8759), .A2(n8817), .ZN(n9045) );
  INV_X1 U9071 ( .A(n9046), .ZN(n8739) );
  NOR2_X1 U9072 ( .A1(n9047), .A2(n9040), .ZN(n9046) );
  NOR2_X1 U9073 ( .A1(n9048), .A2(n9049), .ZN(n9040) );
  NOR3_X1 U9074 ( .A1(n8759), .A2(n9050), .A3(n8305), .ZN(n9049) );
  NOR2_X1 U9075 ( .A1(n8749), .A2(n8747), .ZN(n9050) );
  INV_X1 U9076 ( .A(n9051), .ZN(n9048) );
  NAND2_X1 U9077 ( .A1(n8747), .A2(n8749), .ZN(n9051) );
  NAND2_X1 U9078 ( .A1(n8756), .A2(n9052), .ZN(n8749) );
  NAND2_X1 U9079 ( .A1(n8755), .A2(n8757), .ZN(n9052) );
  NAND2_X1 U9080 ( .A1(n9053), .A2(n9054), .ZN(n8757) );
  NAND2_X1 U9081 ( .A1(b_30_), .A2(a_22_), .ZN(n9054) );
  INV_X1 U9082 ( .A(n9055), .ZN(n9053) );
  XNOR2_X1 U9083 ( .A(n9056), .B(n9057), .ZN(n8755) );
  NAND2_X1 U9084 ( .A1(n9058), .A2(n9059), .ZN(n9056) );
  NAND2_X1 U9085 ( .A1(a_22_), .A2(n9055), .ZN(n8756) );
  NAND2_X1 U9086 ( .A1(n8766), .A2(n9060), .ZN(n9055) );
  NAND2_X1 U9087 ( .A1(n8765), .A2(n8767), .ZN(n9060) );
  NAND2_X1 U9088 ( .A1(n9061), .A2(n9062), .ZN(n8767) );
  NAND2_X1 U9089 ( .A1(b_30_), .A2(a_23_), .ZN(n9062) );
  INV_X1 U9090 ( .A(n9063), .ZN(n9061) );
  XNOR2_X1 U9091 ( .A(n9064), .B(n9065), .ZN(n8765) );
  XNOR2_X1 U9092 ( .A(n9066), .B(n9067), .ZN(n9064) );
  NAND2_X1 U9093 ( .A1(a_23_), .A2(n9063), .ZN(n8766) );
  NAND2_X1 U9094 ( .A1(n9068), .A2(n9069), .ZN(n9063) );
  NAND2_X1 U9095 ( .A1(n8775), .A2(n9070), .ZN(n9069) );
  NAND2_X1 U9096 ( .A1(n8773), .A2(n8774), .ZN(n9070) );
  NOR2_X1 U9097 ( .A1(n8305), .A2(n8779), .ZN(n8775) );
  NAND2_X1 U9098 ( .A1(n9071), .A2(n9072), .ZN(n9068) );
  INV_X1 U9099 ( .A(n8774), .ZN(n9072) );
  NOR2_X1 U9100 ( .A1(n9073), .A2(n9074), .ZN(n8774) );
  INV_X1 U9101 ( .A(n9075), .ZN(n9074) );
  NAND2_X1 U9102 ( .A1(n8784), .A2(n9076), .ZN(n9075) );
  NAND2_X1 U9103 ( .A1(n8782), .A2(n8783), .ZN(n9076) );
  NOR2_X1 U9104 ( .A1(n8305), .A2(n8788), .ZN(n8784) );
  NOR2_X1 U9105 ( .A1(n8782), .A2(n8783), .ZN(n9073) );
  NAND2_X1 U9106 ( .A1(n9077), .A2(n9078), .ZN(n8783) );
  NAND2_X1 U9107 ( .A1(n8826), .A2(n9079), .ZN(n9078) );
  INV_X1 U9108 ( .A(n9080), .ZN(n9079) );
  NOR2_X1 U9109 ( .A1(n8829), .A2(n8828), .ZN(n9080) );
  XOR2_X1 U9110 ( .A(n9081), .B(n9082), .Z(n8826) );
  XOR2_X1 U9111 ( .A(n9083), .B(n9084), .Z(n9082) );
  NAND2_X1 U9112 ( .A1(b_29_), .A2(a_27_), .ZN(n9084) );
  NAND2_X1 U9113 ( .A1(n8828), .A2(n8829), .ZN(n9077) );
  NAND2_X1 U9114 ( .A1(b_30_), .A2(a_26_), .ZN(n8829) );
  NOR2_X1 U9115 ( .A1(n9085), .A2(n9086), .ZN(n8828) );
  INV_X1 U9116 ( .A(n9087), .ZN(n9086) );
  NAND3_X1 U9117 ( .A1(a_27_), .A2(n9088), .A3(b_30_), .ZN(n9087) );
  NAND2_X1 U9118 ( .A1(n8824), .A2(n8823), .ZN(n9088) );
  NOR2_X1 U9119 ( .A1(n8823), .A2(n8824), .ZN(n9085) );
  NOR2_X1 U9120 ( .A1(n9089), .A2(n9090), .ZN(n8824) );
  INV_X1 U9121 ( .A(n9091), .ZN(n9090) );
  NAND2_X1 U9122 ( .A1(n8820), .A2(n9092), .ZN(n9091) );
  NAND2_X1 U9123 ( .A1(n8821), .A2(n8819), .ZN(n9092) );
  NOR2_X1 U9124 ( .A1(n8305), .A2(n8314), .ZN(n8820) );
  NOR2_X1 U9125 ( .A1(n8819), .A2(n8821), .ZN(n9089) );
  NOR2_X1 U9126 ( .A1(n9093), .A2(n9094), .ZN(n8821) );
  INV_X1 U9127 ( .A(n9095), .ZN(n9094) );
  NAND2_X1 U9128 ( .A1(n8804), .A2(n9096), .ZN(n9095) );
  NAND2_X1 U9129 ( .A1(n9097), .A2(n8806), .ZN(n9096) );
  NOR2_X1 U9130 ( .A1(n8305), .A2(n9098), .ZN(n8804) );
  NOR2_X1 U9131 ( .A1(n8806), .A2(n9097), .ZN(n9093) );
  INV_X1 U9132 ( .A(n8805), .ZN(n9097) );
  NAND2_X1 U9133 ( .A1(n9099), .A2(n9100), .ZN(n8805) );
  NAND2_X1 U9134 ( .A1(b_28_), .A2(n9101), .ZN(n9100) );
  NAND2_X1 U9135 ( .A1(n8299), .A2(n9102), .ZN(n9101) );
  NAND2_X1 U9136 ( .A1(a_31_), .A2(n8817), .ZN(n9102) );
  NAND2_X1 U9137 ( .A1(b_29_), .A2(n9103), .ZN(n9099) );
  NAND2_X1 U9138 ( .A1(n8303), .A2(n9104), .ZN(n9103) );
  NAND2_X1 U9139 ( .A1(a_30_), .A2(n9105), .ZN(n9104) );
  NAND3_X1 U9140 ( .A1(b_29_), .A2(n9106), .A3(b_30_), .ZN(n8806) );
  XNOR2_X1 U9141 ( .A(n9107), .B(n9108), .ZN(n8819) );
  XNOR2_X1 U9142 ( .A(n9109), .B(n9110), .ZN(n9107) );
  XNOR2_X1 U9143 ( .A(n9111), .B(n9112), .ZN(n8823) );
  XOR2_X1 U9144 ( .A(n9113), .B(n9114), .Z(n9111) );
  XNOR2_X1 U9145 ( .A(n9115), .B(n9116), .ZN(n8782) );
  XNOR2_X1 U9146 ( .A(n9117), .B(n9118), .ZN(n9116) );
  INV_X1 U9147 ( .A(n8773), .ZN(n9071) );
  XOR2_X1 U9148 ( .A(n9119), .B(n9120), .Z(n8773) );
  XNOR2_X1 U9149 ( .A(n9121), .B(n9122), .ZN(n9120) );
  XNOR2_X1 U9150 ( .A(n9123), .B(n9124), .ZN(n8747) );
  NAND2_X1 U9151 ( .A1(n9125), .A2(n9126), .ZN(n9123) );
  XNOR2_X1 U9152 ( .A(n9127), .B(n9128), .ZN(n8830) );
  NAND2_X1 U9153 ( .A1(n9129), .A2(n9130), .ZN(n9127) );
  XNOR2_X1 U9154 ( .A(n9131), .B(n9132), .ZN(n8847) );
  NAND2_X1 U9155 ( .A1(n9133), .A2(n9134), .ZN(n9131) );
  XNOR2_X1 U9156 ( .A(n9135), .B(n9136), .ZN(n8855) );
  NAND2_X1 U9157 ( .A1(n9137), .A2(n9138), .ZN(n9135) );
  XNOR2_X1 U9158 ( .A(n9139), .B(n9140), .ZN(n8864) );
  NAND2_X1 U9159 ( .A1(n9141), .A2(n9142), .ZN(n9139) );
  XNOR2_X1 U9160 ( .A(n9143), .B(n9144), .ZN(n8872) );
  NAND2_X1 U9161 ( .A1(n9145), .A2(n9146), .ZN(n9143) );
  XNOR2_X1 U9162 ( .A(n9147), .B(n9148), .ZN(n8881) );
  XOR2_X1 U9163 ( .A(n9149), .B(n9150), .Z(n9147) );
  XNOR2_X1 U9164 ( .A(n9151), .B(n9152), .ZN(n8897) );
  NAND2_X1 U9165 ( .A1(n9153), .A2(n9154), .ZN(n9151) );
  XNOR2_X1 U9166 ( .A(n9155), .B(n9156), .ZN(n8906) );
  XNOR2_X1 U9167 ( .A(n9157), .B(n9158), .ZN(n9156) );
  XOR2_X1 U9168 ( .A(n9159), .B(n9160), .Z(n8654) );
  XOR2_X1 U9169 ( .A(n9161), .B(n9162), .Z(n9159) );
  XNOR2_X1 U9170 ( .A(n9163), .B(n9164), .ZN(n8652) );
  NAND2_X1 U9171 ( .A1(n9165), .A2(n9166), .ZN(n9163) );
  NAND4_X1 U9172 ( .A1(n8645), .A2(n9167), .A3(n8646), .A4(n8641), .ZN(n8472)
         );
  NAND2_X1 U9173 ( .A1(n9165), .A2(n9168), .ZN(n8646) );
  NAND2_X1 U9174 ( .A1(n9164), .A2(n9166), .ZN(n9168) );
  NAND2_X1 U9175 ( .A1(n9169), .A2(n9170), .ZN(n9166) );
  NAND2_X1 U9176 ( .A1(b_29_), .A2(a_0_), .ZN(n9170) );
  INV_X1 U9177 ( .A(n9171), .ZN(n9169) );
  XOR2_X1 U9178 ( .A(n9172), .B(n9173), .Z(n9164) );
  XOR2_X1 U9179 ( .A(n9174), .B(n9175), .Z(n9172) );
  NAND2_X1 U9180 ( .A1(a_0_), .A2(n9171), .ZN(n9165) );
  NAND2_X1 U9181 ( .A1(n9176), .A2(n9177), .ZN(n9171) );
  NAND2_X1 U9182 ( .A1(n9162), .A2(n9178), .ZN(n9177) );
  INV_X1 U9183 ( .A(n9179), .ZN(n9178) );
  NOR2_X1 U9184 ( .A1(n9161), .A2(n9160), .ZN(n9179) );
  NOR2_X1 U9185 ( .A1(n8817), .A2(n8569), .ZN(n9162) );
  NAND2_X1 U9186 ( .A1(n9160), .A2(n9161), .ZN(n9176) );
  NAND2_X1 U9187 ( .A1(n9180), .A2(n9181), .ZN(n9161) );
  NAND2_X1 U9188 ( .A1(n9157), .A2(n9182), .ZN(n9181) );
  NAND2_X1 U9189 ( .A1(n9183), .A2(n9184), .ZN(n9182) );
  INV_X1 U9190 ( .A(n9158), .ZN(n9184) );
  INV_X1 U9191 ( .A(n9155), .ZN(n9183) );
  NAND2_X1 U9192 ( .A1(n9185), .A2(n9186), .ZN(n9157) );
  INV_X1 U9193 ( .A(n9187), .ZN(n9186) );
  NOR3_X1 U9194 ( .A1(n8900), .A2(n9188), .A3(n8817), .ZN(n9187) );
  NOR2_X1 U9195 ( .A1(n8924), .A2(n8922), .ZN(n9188) );
  NAND2_X1 U9196 ( .A1(n8922), .A2(n8924), .ZN(n9185) );
  NAND2_X1 U9197 ( .A1(n9153), .A2(n9189), .ZN(n8924) );
  NAND2_X1 U9198 ( .A1(n9152), .A2(n9154), .ZN(n9189) );
  NAND2_X1 U9199 ( .A1(n9190), .A2(n9191), .ZN(n9154) );
  NAND2_X1 U9200 ( .A1(b_29_), .A2(a_4_), .ZN(n9191) );
  XOR2_X1 U9201 ( .A(n9192), .B(n9193), .Z(n9152) );
  XOR2_X1 U9202 ( .A(n9194), .B(n9195), .Z(n9192) );
  NOR2_X1 U9203 ( .A1(n8938), .A2(n9105), .ZN(n9195) );
  NAND2_X1 U9204 ( .A1(a_4_), .A2(n9196), .ZN(n9153) );
  INV_X1 U9205 ( .A(n9190), .ZN(n9196) );
  NOR2_X1 U9206 ( .A1(n9197), .A2(n9198), .ZN(n9190) );
  NOR3_X1 U9207 ( .A1(n8938), .A2(n9199), .A3(n8817), .ZN(n9198) );
  NOR2_X1 U9208 ( .A1(n8936), .A2(n8934), .ZN(n9199) );
  INV_X1 U9209 ( .A(n9200), .ZN(n9197) );
  NAND2_X1 U9210 ( .A1(n8934), .A2(n8936), .ZN(n9200) );
  NAND2_X1 U9211 ( .A1(n8946), .A2(n9201), .ZN(n8936) );
  NAND2_X1 U9212 ( .A1(n8945), .A2(n8947), .ZN(n9201) );
  NAND2_X1 U9213 ( .A1(n9202), .A2(n9203), .ZN(n8947) );
  NAND2_X1 U9214 ( .A1(b_29_), .A2(a_6_), .ZN(n9203) );
  INV_X1 U9215 ( .A(n9204), .ZN(n9202) );
  XNOR2_X1 U9216 ( .A(n9205), .B(n9206), .ZN(n8945) );
  XNOR2_X1 U9217 ( .A(n9207), .B(n9208), .ZN(n9205) );
  NOR2_X1 U9218 ( .A1(n8425), .A2(n9105), .ZN(n9208) );
  NAND2_X1 U9219 ( .A1(a_6_), .A2(n9204), .ZN(n8946) );
  NAND2_X1 U9220 ( .A1(n9209), .A2(n9210), .ZN(n9204) );
  NAND3_X1 U9221 ( .A1(a_7_), .A2(n9211), .A3(b_29_), .ZN(n9210) );
  NAND2_X1 U9222 ( .A1(n9212), .A2(n9213), .ZN(n9211) );
  INV_X1 U9223 ( .A(n8954), .ZN(n9213) );
  INV_X1 U9224 ( .A(n8952), .ZN(n9212) );
  NAND2_X1 U9225 ( .A1(n8954), .A2(n8952), .ZN(n9209) );
  XNOR2_X1 U9226 ( .A(n9214), .B(n9215), .ZN(n8952) );
  XOR2_X1 U9227 ( .A(n9216), .B(n9217), .Z(n9214) );
  NOR2_X1 U9228 ( .A1(n9218), .A2(n9219), .ZN(n8954) );
  INV_X1 U9229 ( .A(n9220), .ZN(n9219) );
  NAND2_X1 U9230 ( .A1(n9148), .A2(n9221), .ZN(n9220) );
  NAND2_X1 U9231 ( .A1(n9150), .A2(n9149), .ZN(n9221) );
  XOR2_X1 U9232 ( .A(n9222), .B(n9223), .Z(n9148) );
  NAND2_X1 U9233 ( .A1(n9224), .A2(n9225), .ZN(n9222) );
  NOR2_X1 U9234 ( .A1(n9149), .A2(n9150), .ZN(n9218) );
  NOR2_X1 U9235 ( .A1(n8817), .A2(n8968), .ZN(n9150) );
  NAND2_X1 U9236 ( .A1(n9226), .A2(n9227), .ZN(n9149) );
  NAND3_X1 U9237 ( .A1(a_9_), .A2(n9228), .A3(b_29_), .ZN(n9227) );
  INV_X1 U9238 ( .A(n9229), .ZN(n9228) );
  NOR2_X1 U9239 ( .A1(n8965), .A2(n8963), .ZN(n9229) );
  NAND2_X1 U9240 ( .A1(n8963), .A2(n8965), .ZN(n9226) );
  NAND2_X1 U9241 ( .A1(n9145), .A2(n9230), .ZN(n8965) );
  NAND2_X1 U9242 ( .A1(n9144), .A2(n9146), .ZN(n9230) );
  NAND2_X1 U9243 ( .A1(n9231), .A2(n9232), .ZN(n9146) );
  NAND2_X1 U9244 ( .A1(b_29_), .A2(a_10_), .ZN(n9232) );
  INV_X1 U9245 ( .A(n9233), .ZN(n9231) );
  XOR2_X1 U9246 ( .A(n9234), .B(n9235), .Z(n9144) );
  XOR2_X1 U9247 ( .A(n9236), .B(n9237), .Z(n9234) );
  NOR2_X1 U9248 ( .A1(n8867), .A2(n9105), .ZN(n9237) );
  NAND2_X1 U9249 ( .A1(a_10_), .A2(n9233), .ZN(n9145) );
  NAND2_X1 U9250 ( .A1(n9238), .A2(n9239), .ZN(n9233) );
  INV_X1 U9251 ( .A(n9240), .ZN(n9239) );
  NOR3_X1 U9252 ( .A1(n8867), .A2(n9241), .A3(n8817), .ZN(n9240) );
  NOR2_X1 U9253 ( .A1(n8979), .A2(n8978), .ZN(n9241) );
  NAND2_X1 U9254 ( .A1(n8978), .A2(n8979), .ZN(n9238) );
  NAND2_X1 U9255 ( .A1(n9141), .A2(n9242), .ZN(n8979) );
  NAND2_X1 U9256 ( .A1(n9140), .A2(n9142), .ZN(n9242) );
  NAND2_X1 U9257 ( .A1(n9243), .A2(n9244), .ZN(n9142) );
  NAND2_X1 U9258 ( .A1(b_29_), .A2(a_12_), .ZN(n9244) );
  INV_X1 U9259 ( .A(n9245), .ZN(n9243) );
  XNOR2_X1 U9260 ( .A(n9246), .B(n9247), .ZN(n9140) );
  XOR2_X1 U9261 ( .A(n9248), .B(n9249), .Z(n9247) );
  NAND2_X1 U9262 ( .A1(b_28_), .A2(a_13_), .ZN(n9249) );
  NAND2_X1 U9263 ( .A1(a_12_), .A2(n9245), .ZN(n9141) );
  NAND2_X1 U9264 ( .A1(n9250), .A2(n9251), .ZN(n9245) );
  INV_X1 U9265 ( .A(n9252), .ZN(n9251) );
  NOR3_X1 U9266 ( .A1(n8996), .A2(n9253), .A3(n8817), .ZN(n9252) );
  NOR2_X1 U9267 ( .A1(n8991), .A2(n8989), .ZN(n9253) );
  NAND2_X1 U9268 ( .A1(n8989), .A2(n8991), .ZN(n9250) );
  NAND2_X1 U9269 ( .A1(n9137), .A2(n9254), .ZN(n8991) );
  NAND2_X1 U9270 ( .A1(n9136), .A2(n9138), .ZN(n9254) );
  NAND2_X1 U9271 ( .A1(n9255), .A2(n9256), .ZN(n9138) );
  NAND2_X1 U9272 ( .A1(b_29_), .A2(a_14_), .ZN(n9256) );
  XOR2_X1 U9273 ( .A(n9257), .B(n9258), .Z(n9136) );
  XOR2_X1 U9274 ( .A(n9259), .B(n9260), .Z(n9257) );
  NOR2_X1 U9275 ( .A1(n8850), .A2(n9105), .ZN(n9260) );
  INV_X1 U9276 ( .A(n9261), .ZN(n9137) );
  NOR2_X1 U9277 ( .A1(n9262), .A2(n9255), .ZN(n9261) );
  NOR2_X1 U9278 ( .A1(n9263), .A2(n9264), .ZN(n9255) );
  NOR3_X1 U9279 ( .A1(n8850), .A2(n9265), .A3(n8817), .ZN(n9264) );
  NOR2_X1 U9280 ( .A1(n9005), .A2(n9004), .ZN(n9265) );
  INV_X1 U9281 ( .A(n9266), .ZN(n9263) );
  NAND2_X1 U9282 ( .A1(n9004), .A2(n9005), .ZN(n9266) );
  NAND2_X1 U9283 ( .A1(n9133), .A2(n9267), .ZN(n9005) );
  NAND2_X1 U9284 ( .A1(n9132), .A2(n9134), .ZN(n9267) );
  NAND2_X1 U9285 ( .A1(n9268), .A2(n9269), .ZN(n9134) );
  NAND2_X1 U9286 ( .A1(b_29_), .A2(a_16_), .ZN(n9269) );
  INV_X1 U9287 ( .A(n9270), .ZN(n9268) );
  XNOR2_X1 U9288 ( .A(n9271), .B(n9272), .ZN(n9132) );
  XOR2_X1 U9289 ( .A(n9273), .B(n9274), .Z(n9272) );
  NAND2_X1 U9290 ( .A1(b_28_), .A2(a_17_), .ZN(n9274) );
  NAND2_X1 U9291 ( .A1(a_16_), .A2(n9270), .ZN(n9133) );
  NAND2_X1 U9292 ( .A1(n9275), .A2(n9276), .ZN(n9270) );
  NAND3_X1 U9293 ( .A1(a_17_), .A2(n9277), .A3(b_29_), .ZN(n9276) );
  NAND2_X1 U9294 ( .A1(n9014), .A2(n9016), .ZN(n9277) );
  INV_X1 U9295 ( .A(n9278), .ZN(n9275) );
  NOR2_X1 U9296 ( .A1(n9016), .A2(n9014), .ZN(n9278) );
  XNOR2_X1 U9297 ( .A(n9279), .B(n9280), .ZN(n9014) );
  XNOR2_X1 U9298 ( .A(n9281), .B(n9282), .ZN(n9280) );
  NAND2_X1 U9299 ( .A1(n9283), .A2(n9284), .ZN(n9016) );
  NAND2_X1 U9300 ( .A1(n9024), .A2(n9285), .ZN(n9284) );
  NAND2_X1 U9301 ( .A1(n9026), .A2(n9025), .ZN(n9285) );
  XNOR2_X1 U9302 ( .A(n9286), .B(n9287), .ZN(n9024) );
  XOR2_X1 U9303 ( .A(n9288), .B(n9289), .Z(n9286) );
  NOR2_X1 U9304 ( .A1(n8742), .A2(n9105), .ZN(n9289) );
  INV_X1 U9305 ( .A(n9290), .ZN(n9283) );
  NOR2_X1 U9306 ( .A1(n9025), .A2(n9026), .ZN(n9290) );
  NOR2_X1 U9307 ( .A1(n8817), .A2(n9291), .ZN(n9026) );
  NAND2_X1 U9308 ( .A1(n9292), .A2(n9293), .ZN(n9025) );
  NAND3_X1 U9309 ( .A1(a_19_), .A2(n9294), .A3(b_29_), .ZN(n9293) );
  INV_X1 U9310 ( .A(n9295), .ZN(n9294) );
  NOR2_X1 U9311 ( .A1(n9033), .A2(n9032), .ZN(n9295) );
  NAND2_X1 U9312 ( .A1(n9032), .A2(n9033), .ZN(n9292) );
  NAND2_X1 U9313 ( .A1(n9129), .A2(n9296), .ZN(n9033) );
  NAND2_X1 U9314 ( .A1(n9128), .A2(n9130), .ZN(n9296) );
  NAND2_X1 U9315 ( .A1(n9297), .A2(n9298), .ZN(n9130) );
  NAND2_X1 U9316 ( .A1(b_29_), .A2(a_20_), .ZN(n9298) );
  XNOR2_X1 U9317 ( .A(n9299), .B(n9300), .ZN(n9128) );
  XOR2_X1 U9318 ( .A(n9301), .B(n9302), .Z(n9300) );
  NAND2_X1 U9319 ( .A1(b_28_), .A2(a_21_), .ZN(n9302) );
  INV_X1 U9320 ( .A(n9303), .ZN(n9129) );
  NOR2_X1 U9321 ( .A1(n9047), .A2(n9297), .ZN(n9303) );
  NOR2_X1 U9322 ( .A1(n9304), .A2(n9305), .ZN(n9297) );
  NOR3_X1 U9323 ( .A1(n8759), .A2(n9306), .A3(n8817), .ZN(n9305) );
  NOR2_X1 U9324 ( .A1(n9044), .A2(n9043), .ZN(n9306) );
  INV_X1 U9325 ( .A(n9307), .ZN(n9304) );
  NAND2_X1 U9326 ( .A1(n9043), .A2(n9044), .ZN(n9307) );
  NAND2_X1 U9327 ( .A1(n9125), .A2(n9308), .ZN(n9044) );
  NAND2_X1 U9328 ( .A1(n9124), .A2(n9126), .ZN(n9308) );
  NAND2_X1 U9329 ( .A1(n9309), .A2(n9310), .ZN(n9126) );
  NAND2_X1 U9330 ( .A1(b_29_), .A2(a_22_), .ZN(n9310) );
  INV_X1 U9331 ( .A(n9311), .ZN(n9309) );
  XNOR2_X1 U9332 ( .A(n9312), .B(n9313), .ZN(n9124) );
  NAND2_X1 U9333 ( .A1(n9314), .A2(n9315), .ZN(n9312) );
  NAND2_X1 U9334 ( .A1(a_22_), .A2(n9311), .ZN(n9125) );
  NAND2_X1 U9335 ( .A1(n9058), .A2(n9316), .ZN(n9311) );
  NAND2_X1 U9336 ( .A1(n9057), .A2(n9059), .ZN(n9316) );
  NAND2_X1 U9337 ( .A1(n9317), .A2(n9318), .ZN(n9059) );
  NAND2_X1 U9338 ( .A1(b_29_), .A2(a_23_), .ZN(n9318) );
  XOR2_X1 U9339 ( .A(n9319), .B(n9320), .Z(n9057) );
  XOR2_X1 U9340 ( .A(n9321), .B(n9322), .Z(n9319) );
  NAND2_X1 U9341 ( .A1(a_23_), .A2(n9323), .ZN(n9058) );
  INV_X1 U9342 ( .A(n9317), .ZN(n9323) );
  NOR2_X1 U9343 ( .A1(n9324), .A2(n9325), .ZN(n9317) );
  INV_X1 U9344 ( .A(n9326), .ZN(n9325) );
  NAND2_X1 U9345 ( .A1(n9067), .A2(n9327), .ZN(n9326) );
  NAND2_X1 U9346 ( .A1(n9066), .A2(n9065), .ZN(n9327) );
  NOR2_X1 U9347 ( .A1(n8817), .A2(n8779), .ZN(n9067) );
  NOR2_X1 U9348 ( .A1(n9065), .A2(n9066), .ZN(n9324) );
  NOR2_X1 U9349 ( .A1(n9328), .A2(n9329), .ZN(n9066) );
  INV_X1 U9350 ( .A(n9330), .ZN(n9329) );
  NAND2_X1 U9351 ( .A1(n9122), .A2(n9331), .ZN(n9330) );
  NAND2_X1 U9352 ( .A1(n9119), .A2(n9121), .ZN(n9331) );
  NOR2_X1 U9353 ( .A1(n8817), .A2(n8788), .ZN(n9122) );
  NOR2_X1 U9354 ( .A1(n9121), .A2(n9119), .ZN(n9328) );
  XNOR2_X1 U9355 ( .A(n9332), .B(n9333), .ZN(n9119) );
  XNOR2_X1 U9356 ( .A(n9334), .B(n9335), .ZN(n9333) );
  NAND2_X1 U9357 ( .A1(n9336), .A2(n9337), .ZN(n9121) );
  NAND2_X1 U9358 ( .A1(n9115), .A2(n9338), .ZN(n9337) );
  NAND2_X1 U9359 ( .A1(n9118), .A2(n9117), .ZN(n9338) );
  XOR2_X1 U9360 ( .A(n9339), .B(n9340), .Z(n9115) );
  XNOR2_X1 U9361 ( .A(n9341), .B(n9342), .ZN(n9339) );
  INV_X1 U9362 ( .A(n9343), .ZN(n9336) );
  NOR2_X1 U9363 ( .A1(n9117), .A2(n9118), .ZN(n9343) );
  NOR2_X1 U9364 ( .A1(n8817), .A2(n9344), .ZN(n9118) );
  NAND2_X1 U9365 ( .A1(n9345), .A2(n9346), .ZN(n9117) );
  NAND3_X1 U9366 ( .A1(a_27_), .A2(n9347), .A3(b_29_), .ZN(n9346) );
  INV_X1 U9367 ( .A(n9348), .ZN(n9347) );
  NOR2_X1 U9368 ( .A1(n9083), .A2(n9081), .ZN(n9348) );
  NAND2_X1 U9369 ( .A1(n9081), .A2(n9083), .ZN(n9345) );
  NAND2_X1 U9370 ( .A1(n9349), .A2(n9350), .ZN(n9083) );
  NAND2_X1 U9371 ( .A1(n9114), .A2(n9351), .ZN(n9350) );
  NAND2_X1 U9372 ( .A1(n9112), .A2(n9113), .ZN(n9351) );
  NOR2_X1 U9373 ( .A1(n8817), .A2(n8314), .ZN(n9114) );
  INV_X1 U9374 ( .A(n9352), .ZN(n9349) );
  NOR2_X1 U9375 ( .A1(n9113), .A2(n9112), .ZN(n9352) );
  XNOR2_X1 U9376 ( .A(n9353), .B(n9354), .ZN(n9112) );
  XOR2_X1 U9377 ( .A(n9355), .B(n9356), .Z(n9353) );
  NAND2_X1 U9378 ( .A1(n9357), .A2(n9358), .ZN(n9113) );
  NAND2_X1 U9379 ( .A1(n9359), .A2(n9110), .ZN(n9358) );
  NAND3_X1 U9380 ( .A1(b_28_), .A2(n9106), .A3(b_29_), .ZN(n9110) );
  NAND2_X1 U9381 ( .A1(n9108), .A2(n9109), .ZN(n9359) );
  INV_X1 U9382 ( .A(n9360), .ZN(n9357) );
  NOR2_X1 U9383 ( .A1(n9109), .A2(n9108), .ZN(n9360) );
  NAND2_X1 U9384 ( .A1(n9361), .A2(n9362), .ZN(n9109) );
  NAND2_X1 U9385 ( .A1(b_27_), .A2(n9363), .ZN(n9362) );
  NAND2_X1 U9386 ( .A1(n8299), .A2(n9364), .ZN(n9363) );
  NAND2_X1 U9387 ( .A1(a_31_), .A2(n9105), .ZN(n9364) );
  NAND2_X1 U9388 ( .A1(b_28_), .A2(n9365), .ZN(n9361) );
  NAND2_X1 U9389 ( .A1(n8303), .A2(n9366), .ZN(n9365) );
  NAND2_X1 U9390 ( .A1(a_30_), .A2(n9367), .ZN(n9366) );
  XOR2_X1 U9391 ( .A(n9368), .B(n9369), .Z(n9081) );
  XOR2_X1 U9392 ( .A(n9370), .B(n9371), .Z(n9368) );
  XNOR2_X1 U9393 ( .A(n9372), .B(n9373), .ZN(n9065) );
  XOR2_X1 U9394 ( .A(n9374), .B(n9375), .Z(n9373) );
  XNOR2_X1 U9395 ( .A(n9376), .B(n9377), .ZN(n9043) );
  NAND2_X1 U9396 ( .A1(n9378), .A2(n9379), .ZN(n9376) );
  XNOR2_X1 U9397 ( .A(n9380), .B(n9381), .ZN(n9032) );
  NAND2_X1 U9398 ( .A1(n9382), .A2(n9383), .ZN(n9380) );
  XNOR2_X1 U9399 ( .A(n9384), .B(n9385), .ZN(n9004) );
  NAND2_X1 U9400 ( .A1(n9386), .A2(n9387), .ZN(n9384) );
  XNOR2_X1 U9401 ( .A(n9388), .B(n9389), .ZN(n8989) );
  NAND2_X1 U9402 ( .A1(n9390), .A2(n9391), .ZN(n9388) );
  XNOR2_X1 U9403 ( .A(n9392), .B(n9393), .ZN(n8978) );
  NAND2_X1 U9404 ( .A1(n9394), .A2(n9395), .ZN(n9392) );
  XNOR2_X1 U9405 ( .A(n9396), .B(n9397), .ZN(n8963) );
  NAND2_X1 U9406 ( .A1(n9398), .A2(n9399), .ZN(n9396) );
  XNOR2_X1 U9407 ( .A(n9400), .B(n9401), .ZN(n8934) );
  NAND2_X1 U9408 ( .A1(n9402), .A2(n9403), .ZN(n9400) );
  XNOR2_X1 U9409 ( .A(n9404), .B(n9405), .ZN(n8922) );
  XOR2_X1 U9410 ( .A(n9406), .B(n9407), .Z(n9405) );
  NAND2_X1 U9411 ( .A1(b_28_), .A2(a_4_), .ZN(n9407) );
  NAND2_X1 U9412 ( .A1(n9158), .A2(n9155), .ZN(n9180) );
  XOR2_X1 U9413 ( .A(n9408), .B(n9409), .Z(n9155) );
  XNOR2_X1 U9414 ( .A(n9410), .B(n9411), .ZN(n9409) );
  NAND2_X1 U9415 ( .A1(b_28_), .A2(a_3_), .ZN(n9411) );
  NOR2_X1 U9416 ( .A1(n8817), .A2(n8448), .ZN(n9158) );
  XOR2_X1 U9417 ( .A(n9412), .B(n9413), .Z(n9160) );
  XOR2_X1 U9418 ( .A(n9414), .B(n9415), .Z(n9413) );
  NAND2_X1 U9419 ( .A1(n8647), .A2(n8648), .ZN(n9167) );
  XOR2_X1 U9420 ( .A(n9416), .B(n9417), .Z(n8645) );
  XNOR2_X1 U9421 ( .A(n9418), .B(n9419), .ZN(n9416) );
  NAND2_X1 U9422 ( .A1(b_28_), .A2(a_0_), .ZN(n9418) );
  INV_X1 U9423 ( .A(n9420), .ZN(n8476) );
  NOR2_X1 U9424 ( .A1(n8641), .A2(n8640), .ZN(n9420) );
  NAND2_X1 U9425 ( .A1(n8636), .A2(n9421), .ZN(n8640) );
  NAND2_X1 U9426 ( .A1(n9422), .A2(n9423), .ZN(n9421) );
  INV_X1 U9427 ( .A(n8634), .ZN(n8636) );
  NOR2_X1 U9428 ( .A1(n9422), .A2(n9423), .ZN(n8634) );
  NAND2_X1 U9429 ( .A1(n9424), .A2(n9425), .ZN(n9423) );
  NAND2_X1 U9430 ( .A1(n9426), .A2(n9427), .ZN(n9425) );
  INV_X1 U9431 ( .A(n9428), .ZN(n9427) );
  NOR2_X1 U9432 ( .A1(n9429), .A2(n9430), .ZN(n9428) );
  NAND2_X1 U9433 ( .A1(n9430), .A2(n9429), .ZN(n9424) );
  XOR2_X1 U9434 ( .A(n9431), .B(n9432), .Z(n9422) );
  NAND2_X1 U9435 ( .A1(n9433), .A2(n9434), .ZN(n9431) );
  INV_X1 U9436 ( .A(n9435), .ZN(n8641) );
  NOR2_X1 U9437 ( .A1(n8648), .A2(n8647), .ZN(n9435) );
  NOR2_X1 U9438 ( .A1(n9436), .A2(n9437), .ZN(n8647) );
  NOR3_X1 U9439 ( .A1(n8457), .A2(n9438), .A3(n9105), .ZN(n9437) );
  NOR2_X1 U9440 ( .A1(n9419), .A2(n9417), .ZN(n9438) );
  INV_X1 U9441 ( .A(n9439), .ZN(n9436) );
  NAND2_X1 U9442 ( .A1(n9417), .A2(n9419), .ZN(n9439) );
  NAND2_X1 U9443 ( .A1(n9440), .A2(n9441), .ZN(n9419) );
  NAND2_X1 U9444 ( .A1(n9175), .A2(n9442), .ZN(n9441) );
  INV_X1 U9445 ( .A(n9443), .ZN(n9442) );
  NOR2_X1 U9446 ( .A1(n9174), .A2(n9173), .ZN(n9443) );
  NOR2_X1 U9447 ( .A1(n9105), .A2(n8569), .ZN(n9175) );
  NAND2_X1 U9448 ( .A1(n9173), .A2(n9174), .ZN(n9440) );
  NAND2_X1 U9449 ( .A1(n9444), .A2(n9445), .ZN(n9174) );
  NAND2_X1 U9450 ( .A1(n9414), .A2(n9446), .ZN(n9445) );
  NAND2_X1 U9451 ( .A1(n9415), .A2(n9412), .ZN(n9446) );
  NOR2_X1 U9452 ( .A1(n9105), .A2(n8448), .ZN(n9414) );
  INV_X1 U9453 ( .A(n9447), .ZN(n9444) );
  NOR2_X1 U9454 ( .A1(n9412), .A2(n9415), .ZN(n9447) );
  NOR2_X1 U9455 ( .A1(n9448), .A2(n9449), .ZN(n9415) );
  NOR3_X1 U9456 ( .A1(n8900), .A2(n9450), .A3(n9105), .ZN(n9449) );
  INV_X1 U9457 ( .A(n9451), .ZN(n9450) );
  NAND2_X1 U9458 ( .A1(n9410), .A2(n9408), .ZN(n9451) );
  NOR2_X1 U9459 ( .A1(n9408), .A2(n9410), .ZN(n9448) );
  NOR2_X1 U9460 ( .A1(n9452), .A2(n9453), .ZN(n9410) );
  NOR3_X1 U9461 ( .A1(n8439), .A2(n9454), .A3(n9105), .ZN(n9453) );
  NOR2_X1 U9462 ( .A1(n9406), .A2(n9404), .ZN(n9454) );
  INV_X1 U9463 ( .A(n9455), .ZN(n9452) );
  NAND2_X1 U9464 ( .A1(n9404), .A2(n9406), .ZN(n9455) );
  NAND2_X1 U9465 ( .A1(n9456), .A2(n9457), .ZN(n9406) );
  INV_X1 U9466 ( .A(n9458), .ZN(n9457) );
  NOR3_X1 U9467 ( .A1(n8938), .A2(n9459), .A3(n9105), .ZN(n9458) );
  NOR2_X1 U9468 ( .A1(n9194), .A2(n9193), .ZN(n9459) );
  NAND2_X1 U9469 ( .A1(n9193), .A2(n9194), .ZN(n9456) );
  NAND2_X1 U9470 ( .A1(n9402), .A2(n9460), .ZN(n9194) );
  NAND2_X1 U9471 ( .A1(n9401), .A2(n9403), .ZN(n9460) );
  NAND2_X1 U9472 ( .A1(n9461), .A2(n9462), .ZN(n9403) );
  NAND2_X1 U9473 ( .A1(b_28_), .A2(a_6_), .ZN(n9462) );
  INV_X1 U9474 ( .A(n9463), .ZN(n9461) );
  XOR2_X1 U9475 ( .A(n9464), .B(n9465), .Z(n9401) );
  XOR2_X1 U9476 ( .A(n9466), .B(n9467), .Z(n9464) );
  NOR2_X1 U9477 ( .A1(n8425), .A2(n9367), .ZN(n9467) );
  NAND2_X1 U9478 ( .A1(a_6_), .A2(n9463), .ZN(n9402) );
  NAND2_X1 U9479 ( .A1(n9468), .A2(n9469), .ZN(n9463) );
  INV_X1 U9480 ( .A(n9470), .ZN(n9469) );
  NOR3_X1 U9481 ( .A1(n8425), .A2(n9471), .A3(n9105), .ZN(n9470) );
  NOR2_X1 U9482 ( .A1(n9206), .A2(n9207), .ZN(n9471) );
  NAND2_X1 U9483 ( .A1(n9207), .A2(n9206), .ZN(n9468) );
  XNOR2_X1 U9484 ( .A(n9472), .B(n9473), .ZN(n9206) );
  NAND2_X1 U9485 ( .A1(n9474), .A2(n9475), .ZN(n9472) );
  NOR2_X1 U9486 ( .A1(n9476), .A2(n9477), .ZN(n9207) );
  INV_X1 U9487 ( .A(n9478), .ZN(n9477) );
  NAND2_X1 U9488 ( .A1(n9215), .A2(n9479), .ZN(n9478) );
  NAND2_X1 U9489 ( .A1(n9217), .A2(n9216), .ZN(n9479) );
  XOR2_X1 U9490 ( .A(n9480), .B(n9481), .Z(n9215) );
  XNOR2_X1 U9491 ( .A(n9482), .B(n9483), .ZN(n9481) );
  NOR2_X1 U9492 ( .A1(n8971), .A2(n9367), .ZN(n9483) );
  NOR2_X1 U9493 ( .A1(n9216), .A2(n9217), .ZN(n9476) );
  NOR2_X1 U9494 ( .A1(n9105), .A2(n8968), .ZN(n9217) );
  NAND2_X1 U9495 ( .A1(n9224), .A2(n9484), .ZN(n9216) );
  NAND2_X1 U9496 ( .A1(n9223), .A2(n9225), .ZN(n9484) );
  NAND2_X1 U9497 ( .A1(n9485), .A2(n9486), .ZN(n9225) );
  NAND2_X1 U9498 ( .A1(b_28_), .A2(a_9_), .ZN(n9486) );
  INV_X1 U9499 ( .A(n9487), .ZN(n9485) );
  XNOR2_X1 U9500 ( .A(n9488), .B(n9489), .ZN(n9223) );
  NAND2_X1 U9501 ( .A1(n9490), .A2(n9491), .ZN(n9488) );
  NAND2_X1 U9502 ( .A1(a_9_), .A2(n9487), .ZN(n9224) );
  NAND2_X1 U9503 ( .A1(n9398), .A2(n9492), .ZN(n9487) );
  NAND2_X1 U9504 ( .A1(n9397), .A2(n9399), .ZN(n9492) );
  NAND2_X1 U9505 ( .A1(n9493), .A2(n9494), .ZN(n9399) );
  NAND2_X1 U9506 ( .A1(b_28_), .A2(a_10_), .ZN(n9494) );
  INV_X1 U9507 ( .A(n9495), .ZN(n9493) );
  XNOR2_X1 U9508 ( .A(n9496), .B(n9497), .ZN(n9397) );
  XOR2_X1 U9509 ( .A(n9498), .B(n9499), .Z(n9497) );
  NAND2_X1 U9510 ( .A1(b_27_), .A2(a_11_), .ZN(n9499) );
  NAND2_X1 U9511 ( .A1(a_10_), .A2(n9495), .ZN(n9398) );
  NAND2_X1 U9512 ( .A1(n9500), .A2(n9501), .ZN(n9495) );
  INV_X1 U9513 ( .A(n9502), .ZN(n9501) );
  NOR3_X1 U9514 ( .A1(n8867), .A2(n9503), .A3(n9105), .ZN(n9502) );
  NOR2_X1 U9515 ( .A1(n9236), .A2(n9235), .ZN(n9503) );
  NAND2_X1 U9516 ( .A1(n9235), .A2(n9236), .ZN(n9500) );
  NAND2_X1 U9517 ( .A1(n9394), .A2(n9504), .ZN(n9236) );
  NAND2_X1 U9518 ( .A1(n9393), .A2(n9395), .ZN(n9504) );
  NAND2_X1 U9519 ( .A1(n9505), .A2(n9506), .ZN(n9395) );
  NAND2_X1 U9520 ( .A1(b_28_), .A2(a_12_), .ZN(n9506) );
  INV_X1 U9521 ( .A(n9507), .ZN(n9505) );
  XNOR2_X1 U9522 ( .A(n9508), .B(n9509), .ZN(n9393) );
  XOR2_X1 U9523 ( .A(n9510), .B(n9511), .Z(n9509) );
  NAND2_X1 U9524 ( .A1(b_27_), .A2(a_13_), .ZN(n9511) );
  NAND2_X1 U9525 ( .A1(a_12_), .A2(n9507), .ZN(n9394) );
  NAND2_X1 U9526 ( .A1(n9512), .A2(n9513), .ZN(n9507) );
  INV_X1 U9527 ( .A(n9514), .ZN(n9513) );
  NOR3_X1 U9528 ( .A1(n8996), .A2(n9515), .A3(n9105), .ZN(n9514) );
  NOR2_X1 U9529 ( .A1(n9248), .A2(n9246), .ZN(n9515) );
  NAND2_X1 U9530 ( .A1(n9246), .A2(n9248), .ZN(n9512) );
  NAND2_X1 U9531 ( .A1(n9390), .A2(n9516), .ZN(n9248) );
  NAND2_X1 U9532 ( .A1(n9389), .A2(n9391), .ZN(n9516) );
  NAND2_X1 U9533 ( .A1(n9517), .A2(n9518), .ZN(n9391) );
  NAND2_X1 U9534 ( .A1(b_28_), .A2(a_14_), .ZN(n9518) );
  INV_X1 U9535 ( .A(n9519), .ZN(n9517) );
  XOR2_X1 U9536 ( .A(n9520), .B(n9521), .Z(n9389) );
  XOR2_X1 U9537 ( .A(n9522), .B(n9523), .Z(n9520) );
  NOR2_X1 U9538 ( .A1(n8850), .A2(n9367), .ZN(n9523) );
  NAND2_X1 U9539 ( .A1(a_14_), .A2(n9519), .ZN(n9390) );
  NAND2_X1 U9540 ( .A1(n9524), .A2(n9525), .ZN(n9519) );
  INV_X1 U9541 ( .A(n9526), .ZN(n9525) );
  NOR3_X1 U9542 ( .A1(n8850), .A2(n9527), .A3(n9105), .ZN(n9526) );
  NOR2_X1 U9543 ( .A1(n9259), .A2(n9258), .ZN(n9527) );
  NAND2_X1 U9544 ( .A1(n9258), .A2(n9259), .ZN(n9524) );
  NAND2_X1 U9545 ( .A1(n9386), .A2(n9528), .ZN(n9259) );
  NAND2_X1 U9546 ( .A1(n9385), .A2(n9387), .ZN(n9528) );
  NAND2_X1 U9547 ( .A1(n9529), .A2(n9530), .ZN(n9387) );
  NAND2_X1 U9548 ( .A1(b_28_), .A2(a_16_), .ZN(n9530) );
  XNOR2_X1 U9549 ( .A(n9531), .B(n9532), .ZN(n9385) );
  XOR2_X1 U9550 ( .A(n9533), .B(n9534), .Z(n9532) );
  NAND2_X1 U9551 ( .A1(b_27_), .A2(a_17_), .ZN(n9534) );
  NAND2_X1 U9552 ( .A1(a_16_), .A2(n9535), .ZN(n9386) );
  INV_X1 U9553 ( .A(n9529), .ZN(n9535) );
  NOR2_X1 U9554 ( .A1(n9536), .A2(n9537), .ZN(n9529) );
  NOR3_X1 U9555 ( .A1(n8371), .A2(n9538), .A3(n9105), .ZN(n9537) );
  INV_X1 U9556 ( .A(n9539), .ZN(n9538) );
  NAND2_X1 U9557 ( .A1(n9271), .A2(n9273), .ZN(n9539) );
  NOR2_X1 U9558 ( .A1(n9273), .A2(n9271), .ZN(n9536) );
  XOR2_X1 U9559 ( .A(n9540), .B(n9541), .Z(n9271) );
  XOR2_X1 U9560 ( .A(n9542), .B(n9543), .Z(n9540) );
  NAND2_X1 U9561 ( .A1(n9544), .A2(n9545), .ZN(n9273) );
  NAND2_X1 U9562 ( .A1(n9279), .A2(n9546), .ZN(n9545) );
  NAND2_X1 U9563 ( .A1(n9282), .A2(n9281), .ZN(n9546) );
  XOR2_X1 U9564 ( .A(n9547), .B(n9548), .Z(n9279) );
  XOR2_X1 U9565 ( .A(n9549), .B(n9550), .Z(n9548) );
  NAND2_X1 U9566 ( .A1(b_27_), .A2(a_19_), .ZN(n9550) );
  INV_X1 U9567 ( .A(n9551), .ZN(n9544) );
  NOR2_X1 U9568 ( .A1(n9281), .A2(n9282), .ZN(n9551) );
  NOR2_X1 U9569 ( .A1(n9105), .A2(n9291), .ZN(n9282) );
  NAND2_X1 U9570 ( .A1(n9552), .A2(n9553), .ZN(n9281) );
  NAND3_X1 U9571 ( .A1(a_19_), .A2(n9554), .A3(b_28_), .ZN(n9553) );
  INV_X1 U9572 ( .A(n9555), .ZN(n9554) );
  NOR2_X1 U9573 ( .A1(n9288), .A2(n9287), .ZN(n9555) );
  NAND2_X1 U9574 ( .A1(n9287), .A2(n9288), .ZN(n9552) );
  NAND2_X1 U9575 ( .A1(n9382), .A2(n9556), .ZN(n9288) );
  NAND2_X1 U9576 ( .A1(n9381), .A2(n9383), .ZN(n9556) );
  NAND2_X1 U9577 ( .A1(n9557), .A2(n9558), .ZN(n9383) );
  NAND2_X1 U9578 ( .A1(b_28_), .A2(a_20_), .ZN(n9558) );
  INV_X1 U9579 ( .A(n9559), .ZN(n9557) );
  XNOR2_X1 U9580 ( .A(n9560), .B(n9561), .ZN(n9381) );
  XOR2_X1 U9581 ( .A(n9562), .B(n9563), .Z(n9561) );
  NAND2_X1 U9582 ( .A1(b_27_), .A2(a_21_), .ZN(n9563) );
  NAND2_X1 U9583 ( .A1(a_20_), .A2(n9559), .ZN(n9382) );
  NAND2_X1 U9584 ( .A1(n9564), .A2(n9565), .ZN(n9559) );
  INV_X1 U9585 ( .A(n9566), .ZN(n9565) );
  NOR3_X1 U9586 ( .A1(n8759), .A2(n9567), .A3(n9105), .ZN(n9566) );
  NOR2_X1 U9587 ( .A1(n9301), .A2(n9299), .ZN(n9567) );
  NAND2_X1 U9588 ( .A1(n9299), .A2(n9301), .ZN(n9564) );
  NAND2_X1 U9589 ( .A1(n9378), .A2(n9568), .ZN(n9301) );
  NAND2_X1 U9590 ( .A1(n9377), .A2(n9379), .ZN(n9568) );
  NAND2_X1 U9591 ( .A1(n9569), .A2(n9570), .ZN(n9379) );
  NAND2_X1 U9592 ( .A1(b_28_), .A2(a_22_), .ZN(n9570) );
  INV_X1 U9593 ( .A(n9571), .ZN(n9569) );
  XNOR2_X1 U9594 ( .A(n9572), .B(n9573), .ZN(n9377) );
  NAND2_X1 U9595 ( .A1(n9574), .A2(n9575), .ZN(n9572) );
  NAND2_X1 U9596 ( .A1(a_22_), .A2(n9571), .ZN(n9378) );
  NAND2_X1 U9597 ( .A1(n9314), .A2(n9576), .ZN(n9571) );
  NAND2_X1 U9598 ( .A1(n9313), .A2(n9315), .ZN(n9576) );
  NAND2_X1 U9599 ( .A1(n9577), .A2(n9578), .ZN(n9315) );
  NAND2_X1 U9600 ( .A1(b_28_), .A2(a_23_), .ZN(n9578) );
  INV_X1 U9601 ( .A(n9579), .ZN(n9577) );
  XNOR2_X1 U9602 ( .A(n9580), .B(n9581), .ZN(n9313) );
  XOR2_X1 U9603 ( .A(n9582), .B(n9583), .Z(n9581) );
  NAND2_X1 U9604 ( .A1(a_23_), .A2(n9579), .ZN(n9314) );
  NAND2_X1 U9605 ( .A1(n9584), .A2(n9585), .ZN(n9579) );
  NAND2_X1 U9606 ( .A1(n9322), .A2(n9586), .ZN(n9585) );
  INV_X1 U9607 ( .A(n9587), .ZN(n9586) );
  NOR2_X1 U9608 ( .A1(n9321), .A2(n9320), .ZN(n9587) );
  NOR2_X1 U9609 ( .A1(n9105), .A2(n8779), .ZN(n9322) );
  NAND2_X1 U9610 ( .A1(n9320), .A2(n9321), .ZN(n9584) );
  NAND2_X1 U9611 ( .A1(n9588), .A2(n9589), .ZN(n9321) );
  NAND2_X1 U9612 ( .A1(n9375), .A2(n9590), .ZN(n9589) );
  INV_X1 U9613 ( .A(n9591), .ZN(n9590) );
  NOR2_X1 U9614 ( .A1(n9372), .A2(n9374), .ZN(n9591) );
  NOR2_X1 U9615 ( .A1(n9105), .A2(n8788), .ZN(n9375) );
  NAND2_X1 U9616 ( .A1(n9374), .A2(n9372), .ZN(n9588) );
  XNOR2_X1 U9617 ( .A(n9592), .B(n9593), .ZN(n9372) );
  NAND2_X1 U9618 ( .A1(n9594), .A2(n9595), .ZN(n9592) );
  NOR2_X1 U9619 ( .A1(n9596), .A2(n9597), .ZN(n9374) );
  INV_X1 U9620 ( .A(n9598), .ZN(n9597) );
  NAND2_X1 U9621 ( .A1(n9332), .A2(n9599), .ZN(n9598) );
  NAND2_X1 U9622 ( .A1(n9335), .A2(n9334), .ZN(n9599) );
  XOR2_X1 U9623 ( .A(n9600), .B(n9601), .Z(n9332) );
  XNOR2_X1 U9624 ( .A(n9602), .B(n9603), .ZN(n9600) );
  NOR2_X1 U9625 ( .A1(n9334), .A2(n9335), .ZN(n9596) );
  NOR2_X1 U9626 ( .A1(n9105), .A2(n9344), .ZN(n9335) );
  NAND2_X1 U9627 ( .A1(n9604), .A2(n9605), .ZN(n9334) );
  NAND2_X1 U9628 ( .A1(n9342), .A2(n9606), .ZN(n9605) );
  INV_X1 U9629 ( .A(n9607), .ZN(n9606) );
  NOR2_X1 U9630 ( .A1(n9340), .A2(n9341), .ZN(n9607) );
  NOR2_X1 U9631 ( .A1(n9105), .A2(n8797), .ZN(n9342) );
  NAND2_X1 U9632 ( .A1(n9341), .A2(n9340), .ZN(n9604) );
  XOR2_X1 U9633 ( .A(n9608), .B(n9609), .Z(n9340) );
  XOR2_X1 U9634 ( .A(n9610), .B(n9611), .Z(n9608) );
  NOR2_X1 U9635 ( .A1(n9612), .A2(n9613), .ZN(n9341) );
  NOR2_X1 U9636 ( .A1(n9614), .A2(n9370), .ZN(n9613) );
  INV_X1 U9637 ( .A(n9615), .ZN(n9614) );
  NAND2_X1 U9638 ( .A1(n9369), .A2(n9371), .ZN(n9615) );
  NOR2_X1 U9639 ( .A1(n9371), .A2(n9369), .ZN(n9612) );
  XOR2_X1 U9640 ( .A(n9616), .B(n9617), .Z(n9369) );
  XOR2_X1 U9641 ( .A(n9618), .B(n9619), .Z(n9616) );
  NAND2_X1 U9642 ( .A1(n9620), .A2(n9621), .ZN(n9371) );
  NAND2_X1 U9643 ( .A1(n9354), .A2(n9622), .ZN(n9621) );
  INV_X1 U9644 ( .A(n9623), .ZN(n9622) );
  NOR2_X1 U9645 ( .A1(n9355), .A2(n9356), .ZN(n9623) );
  NOR2_X1 U9646 ( .A1(n9105), .A2(n9098), .ZN(n9354) );
  NAND2_X1 U9647 ( .A1(n9356), .A2(n9355), .ZN(n9620) );
  NAND2_X1 U9648 ( .A1(n9624), .A2(n9625), .ZN(n9355) );
  NAND2_X1 U9649 ( .A1(b_26_), .A2(n9626), .ZN(n9625) );
  NAND2_X1 U9650 ( .A1(n8299), .A2(n9627), .ZN(n9626) );
  NAND2_X1 U9651 ( .A1(a_31_), .A2(n9367), .ZN(n9627) );
  NAND2_X1 U9652 ( .A1(b_27_), .A2(n9628), .ZN(n9624) );
  NAND2_X1 U9653 ( .A1(n8303), .A2(n9629), .ZN(n9628) );
  NAND2_X1 U9654 ( .A1(a_30_), .A2(n9630), .ZN(n9629) );
  NOR3_X1 U9655 ( .A1(n9367), .A2(n9631), .A3(n9105), .ZN(n9356) );
  XNOR2_X1 U9656 ( .A(n9632), .B(n9633), .ZN(n9320) );
  NAND2_X1 U9657 ( .A1(n9634), .A2(n9635), .ZN(n9632) );
  XNOR2_X1 U9658 ( .A(n9636), .B(n9637), .ZN(n9299) );
  NAND2_X1 U9659 ( .A1(n9638), .A2(n9639), .ZN(n9636) );
  XNOR2_X1 U9660 ( .A(n9640), .B(n9641), .ZN(n9287) );
  NAND2_X1 U9661 ( .A1(n9642), .A2(n9643), .ZN(n9640) );
  XNOR2_X1 U9662 ( .A(n9644), .B(n9645), .ZN(n9258) );
  NAND2_X1 U9663 ( .A1(n9646), .A2(n9647), .ZN(n9644) );
  XNOR2_X1 U9664 ( .A(n9648), .B(n9649), .ZN(n9246) );
  NAND2_X1 U9665 ( .A1(n9650), .A2(n9651), .ZN(n9648) );
  XNOR2_X1 U9666 ( .A(n9652), .B(n9653), .ZN(n9235) );
  XOR2_X1 U9667 ( .A(n9654), .B(n9655), .Z(n9652) );
  XOR2_X1 U9668 ( .A(n9656), .B(n9657), .Z(n9193) );
  XNOR2_X1 U9669 ( .A(n9658), .B(n9659), .ZN(n9657) );
  XOR2_X1 U9670 ( .A(n9660), .B(n9661), .Z(n9404) );
  XOR2_X1 U9671 ( .A(n9662), .B(n9663), .Z(n9660) );
  XNOR2_X1 U9672 ( .A(n9664), .B(n9665), .ZN(n9408) );
  XOR2_X1 U9673 ( .A(n9666), .B(n9667), .Z(n9664) );
  XNOR2_X1 U9674 ( .A(n9668), .B(n9669), .ZN(n9412) );
  XOR2_X1 U9675 ( .A(n9670), .B(n9671), .Z(n9668) );
  NOR2_X1 U9676 ( .A1(n8900), .A2(n9367), .ZN(n9671) );
  XNOR2_X1 U9677 ( .A(n9672), .B(n9673), .ZN(n9173) );
  NAND2_X1 U9678 ( .A1(n9674), .A2(n9675), .ZN(n9672) );
  XOR2_X1 U9679 ( .A(n9676), .B(n9677), .Z(n9417) );
  XOR2_X1 U9680 ( .A(n9678), .B(n9679), .Z(n9676) );
  NOR2_X1 U9681 ( .A1(n8569), .A2(n9367), .ZN(n9679) );
  XNOR2_X1 U9682 ( .A(n9426), .B(n9680), .ZN(n8648) );
  XNOR2_X1 U9683 ( .A(n9430), .B(n9429), .ZN(n9680) );
  NAND2_X1 U9684 ( .A1(b_27_), .A2(a_0_), .ZN(n9429) );
  NOR2_X1 U9685 ( .A1(n9681), .A2(n9682), .ZN(n9430) );
  NOR3_X1 U9686 ( .A1(n8569), .A2(n9683), .A3(n9367), .ZN(n9682) );
  NOR2_X1 U9687 ( .A1(n9678), .A2(n9677), .ZN(n9683) );
  INV_X1 U9688 ( .A(n9684), .ZN(n9681) );
  NAND2_X1 U9689 ( .A1(n9677), .A2(n9678), .ZN(n9684) );
  NAND2_X1 U9690 ( .A1(n9674), .A2(n9685), .ZN(n9678) );
  NAND2_X1 U9691 ( .A1(n9673), .A2(n9675), .ZN(n9685) );
  NAND2_X1 U9692 ( .A1(n9686), .A2(n9687), .ZN(n9675) );
  NAND2_X1 U9693 ( .A1(b_27_), .A2(a_2_), .ZN(n9687) );
  INV_X1 U9694 ( .A(n9688), .ZN(n9686) );
  XOR2_X1 U9695 ( .A(n9689), .B(n9690), .Z(n9673) );
  XNOR2_X1 U9696 ( .A(n9691), .B(n9692), .ZN(n9690) );
  NAND2_X1 U9697 ( .A1(b_26_), .A2(a_3_), .ZN(n9692) );
  NAND2_X1 U9698 ( .A1(a_2_), .A2(n9688), .ZN(n9674) );
  NAND2_X1 U9699 ( .A1(n9693), .A2(n9694), .ZN(n9688) );
  INV_X1 U9700 ( .A(n9695), .ZN(n9694) );
  NOR3_X1 U9701 ( .A1(n8900), .A2(n9696), .A3(n9367), .ZN(n9695) );
  NOR2_X1 U9702 ( .A1(n9670), .A2(n9669), .ZN(n9696) );
  NAND2_X1 U9703 ( .A1(n9669), .A2(n9670), .ZN(n9693) );
  NAND2_X1 U9704 ( .A1(n9697), .A2(n9698), .ZN(n9670) );
  NAND2_X1 U9705 ( .A1(n9667), .A2(n9699), .ZN(n9698) );
  INV_X1 U9706 ( .A(n9700), .ZN(n9699) );
  NOR2_X1 U9707 ( .A1(n9666), .A2(n9665), .ZN(n9700) );
  NOR2_X1 U9708 ( .A1(n9367), .A2(n8439), .ZN(n9667) );
  NAND2_X1 U9709 ( .A1(n9665), .A2(n9666), .ZN(n9697) );
  NAND2_X1 U9710 ( .A1(n9701), .A2(n9702), .ZN(n9666) );
  NAND2_X1 U9711 ( .A1(n9663), .A2(n9703), .ZN(n9702) );
  INV_X1 U9712 ( .A(n9704), .ZN(n9703) );
  NOR2_X1 U9713 ( .A1(n9662), .A2(n9661), .ZN(n9704) );
  NOR2_X1 U9714 ( .A1(n9367), .A2(n8938), .ZN(n9663) );
  NAND2_X1 U9715 ( .A1(n9661), .A2(n9662), .ZN(n9701) );
  NAND2_X1 U9716 ( .A1(n9705), .A2(n9706), .ZN(n9662) );
  NAND2_X1 U9717 ( .A1(n9658), .A2(n9707), .ZN(n9706) );
  NAND2_X1 U9718 ( .A1(n9656), .A2(n9708), .ZN(n9707) );
  INV_X1 U9719 ( .A(n9659), .ZN(n9708) );
  NAND2_X1 U9720 ( .A1(n9709), .A2(n9710), .ZN(n9658) );
  INV_X1 U9721 ( .A(n9711), .ZN(n9710) );
  NOR3_X1 U9722 ( .A1(n8425), .A2(n9712), .A3(n9367), .ZN(n9711) );
  NOR2_X1 U9723 ( .A1(n9466), .A2(n9465), .ZN(n9712) );
  NAND2_X1 U9724 ( .A1(n9465), .A2(n9466), .ZN(n9709) );
  NAND2_X1 U9725 ( .A1(n9474), .A2(n9713), .ZN(n9466) );
  NAND2_X1 U9726 ( .A1(n9473), .A2(n9475), .ZN(n9713) );
  NAND2_X1 U9727 ( .A1(n9714), .A2(n9715), .ZN(n9475) );
  NAND2_X1 U9728 ( .A1(b_27_), .A2(a_8_), .ZN(n9715) );
  INV_X1 U9729 ( .A(n9716), .ZN(n9714) );
  XOR2_X1 U9730 ( .A(n9717), .B(n9718), .Z(n9473) );
  XOR2_X1 U9731 ( .A(n9719), .B(n9720), .Z(n9717) );
  NOR2_X1 U9732 ( .A1(n8971), .A2(n9630), .ZN(n9720) );
  NAND2_X1 U9733 ( .A1(a_8_), .A2(n9716), .ZN(n9474) );
  NAND2_X1 U9734 ( .A1(n9721), .A2(n9722), .ZN(n9716) );
  NAND3_X1 U9735 ( .A1(a_9_), .A2(n9723), .A3(b_27_), .ZN(n9722) );
  INV_X1 U9736 ( .A(n9724), .ZN(n9723) );
  NOR2_X1 U9737 ( .A1(n9482), .A2(n9480), .ZN(n9724) );
  NAND2_X1 U9738 ( .A1(n9480), .A2(n9482), .ZN(n9721) );
  NAND2_X1 U9739 ( .A1(n9490), .A2(n9725), .ZN(n9482) );
  NAND2_X1 U9740 ( .A1(n9489), .A2(n9491), .ZN(n9725) );
  NAND2_X1 U9741 ( .A1(n9726), .A2(n9727), .ZN(n9491) );
  NAND2_X1 U9742 ( .A1(b_27_), .A2(a_10_), .ZN(n9727) );
  XNOR2_X1 U9743 ( .A(n9728), .B(n9729), .ZN(n9489) );
  XNOR2_X1 U9744 ( .A(n9730), .B(n9731), .ZN(n9728) );
  NOR2_X1 U9745 ( .A1(n8867), .A2(n9630), .ZN(n9731) );
  NAND2_X1 U9746 ( .A1(a_10_), .A2(n9732), .ZN(n9490) );
  INV_X1 U9747 ( .A(n9726), .ZN(n9732) );
  NOR2_X1 U9748 ( .A1(n9733), .A2(n9734), .ZN(n9726) );
  INV_X1 U9749 ( .A(n9735), .ZN(n9734) );
  NAND3_X1 U9750 ( .A1(a_11_), .A2(n9736), .A3(b_27_), .ZN(n9735) );
  NAND2_X1 U9751 ( .A1(n9496), .A2(n9498), .ZN(n9736) );
  NOR2_X1 U9752 ( .A1(n9498), .A2(n9496), .ZN(n9733) );
  XOR2_X1 U9753 ( .A(n9737), .B(n9738), .Z(n9496) );
  XOR2_X1 U9754 ( .A(n9739), .B(n9740), .Z(n9737) );
  NAND2_X1 U9755 ( .A1(n9741), .A2(n9742), .ZN(n9498) );
  NAND2_X1 U9756 ( .A1(n9653), .A2(n9743), .ZN(n9742) );
  NAND2_X1 U9757 ( .A1(n9655), .A2(n9654), .ZN(n9743) );
  XOR2_X1 U9758 ( .A(n9744), .B(n9745), .Z(n9653) );
  NAND2_X1 U9759 ( .A1(n9746), .A2(n9747), .ZN(n9744) );
  INV_X1 U9760 ( .A(n9748), .ZN(n9741) );
  NOR2_X1 U9761 ( .A1(n9654), .A2(n9655), .ZN(n9748) );
  NOR2_X1 U9762 ( .A1(n9367), .A2(n8393), .ZN(n9655) );
  NAND2_X1 U9763 ( .A1(n9749), .A2(n9750), .ZN(n9654) );
  NAND3_X1 U9764 ( .A1(a_13_), .A2(n9751), .A3(b_27_), .ZN(n9750) );
  INV_X1 U9765 ( .A(n9752), .ZN(n9751) );
  NOR2_X1 U9766 ( .A1(n9510), .A2(n9508), .ZN(n9752) );
  NAND2_X1 U9767 ( .A1(n9508), .A2(n9510), .ZN(n9749) );
  NAND2_X1 U9768 ( .A1(n9650), .A2(n9753), .ZN(n9510) );
  NAND2_X1 U9769 ( .A1(n9649), .A2(n9651), .ZN(n9753) );
  NAND2_X1 U9770 ( .A1(n9754), .A2(n9755), .ZN(n9651) );
  NAND2_X1 U9771 ( .A1(b_27_), .A2(a_14_), .ZN(n9755) );
  XOR2_X1 U9772 ( .A(n9756), .B(n9757), .Z(n9649) );
  XOR2_X1 U9773 ( .A(n9758), .B(n9759), .Z(n9756) );
  NOR2_X1 U9774 ( .A1(n8850), .A2(n9630), .ZN(n9759) );
  INV_X1 U9775 ( .A(n9760), .ZN(n9650) );
  NOR2_X1 U9776 ( .A1(n9262), .A2(n9754), .ZN(n9760) );
  NOR2_X1 U9777 ( .A1(n9761), .A2(n9762), .ZN(n9754) );
  NOR3_X1 U9778 ( .A1(n8850), .A2(n9763), .A3(n9367), .ZN(n9762) );
  NOR2_X1 U9779 ( .A1(n9522), .A2(n9521), .ZN(n9763) );
  INV_X1 U9780 ( .A(n9764), .ZN(n9761) );
  NAND2_X1 U9781 ( .A1(n9521), .A2(n9522), .ZN(n9764) );
  NAND2_X1 U9782 ( .A1(n9646), .A2(n9765), .ZN(n9522) );
  NAND2_X1 U9783 ( .A1(n9645), .A2(n9647), .ZN(n9765) );
  NAND2_X1 U9784 ( .A1(n9766), .A2(n9767), .ZN(n9647) );
  NAND2_X1 U9785 ( .A1(b_27_), .A2(a_16_), .ZN(n9767) );
  INV_X1 U9786 ( .A(n9768), .ZN(n9766) );
  XNOR2_X1 U9787 ( .A(n9769), .B(n9770), .ZN(n9645) );
  XOR2_X1 U9788 ( .A(n9771), .B(n9772), .Z(n9770) );
  NAND2_X1 U9789 ( .A1(b_26_), .A2(a_17_), .ZN(n9772) );
  NAND2_X1 U9790 ( .A1(a_16_), .A2(n9768), .ZN(n9646) );
  NAND2_X1 U9791 ( .A1(n9773), .A2(n9774), .ZN(n9768) );
  NAND3_X1 U9792 ( .A1(a_17_), .A2(n9775), .A3(b_27_), .ZN(n9774) );
  NAND2_X1 U9793 ( .A1(n9531), .A2(n9533), .ZN(n9775) );
  INV_X1 U9794 ( .A(n9776), .ZN(n9773) );
  NOR2_X1 U9795 ( .A1(n9533), .A2(n9531), .ZN(n9776) );
  XOR2_X1 U9796 ( .A(n9777), .B(n9778), .Z(n9531) );
  XOR2_X1 U9797 ( .A(n9779), .B(n9780), .Z(n9777) );
  NAND2_X1 U9798 ( .A1(n9781), .A2(n9782), .ZN(n9533) );
  NAND2_X1 U9799 ( .A1(n9541), .A2(n9783), .ZN(n9782) );
  NAND2_X1 U9800 ( .A1(n9543), .A2(n9542), .ZN(n9783) );
  XNOR2_X1 U9801 ( .A(n9784), .B(n9785), .ZN(n9541) );
  XOR2_X1 U9802 ( .A(n9786), .B(n9787), .Z(n9784) );
  NOR2_X1 U9803 ( .A1(n8742), .A2(n9630), .ZN(n9787) );
  INV_X1 U9804 ( .A(n9788), .ZN(n9781) );
  NOR2_X1 U9805 ( .A1(n9542), .A2(n9543), .ZN(n9788) );
  NOR2_X1 U9806 ( .A1(n9367), .A2(n9291), .ZN(n9543) );
  NAND2_X1 U9807 ( .A1(n9789), .A2(n9790), .ZN(n9542) );
  NAND3_X1 U9808 ( .A1(a_19_), .A2(n9791), .A3(b_27_), .ZN(n9790) );
  INV_X1 U9809 ( .A(n9792), .ZN(n9791) );
  NOR2_X1 U9810 ( .A1(n9549), .A2(n9547), .ZN(n9792) );
  NAND2_X1 U9811 ( .A1(n9547), .A2(n9549), .ZN(n9789) );
  NAND2_X1 U9812 ( .A1(n9642), .A2(n9793), .ZN(n9549) );
  NAND2_X1 U9813 ( .A1(n9641), .A2(n9643), .ZN(n9793) );
  NAND2_X1 U9814 ( .A1(n9794), .A2(n9795), .ZN(n9643) );
  NAND2_X1 U9815 ( .A1(b_27_), .A2(a_20_), .ZN(n9795) );
  INV_X1 U9816 ( .A(n9796), .ZN(n9794) );
  XNOR2_X1 U9817 ( .A(n9797), .B(n9798), .ZN(n9641) );
  XOR2_X1 U9818 ( .A(n9799), .B(n9800), .Z(n9798) );
  NAND2_X1 U9819 ( .A1(b_26_), .A2(a_21_), .ZN(n9800) );
  NAND2_X1 U9820 ( .A1(a_20_), .A2(n9796), .ZN(n9642) );
  NAND2_X1 U9821 ( .A1(n9801), .A2(n9802), .ZN(n9796) );
  INV_X1 U9822 ( .A(n9803), .ZN(n9802) );
  NOR3_X1 U9823 ( .A1(n8759), .A2(n9804), .A3(n9367), .ZN(n9803) );
  NOR2_X1 U9824 ( .A1(n9562), .A2(n9560), .ZN(n9804) );
  NAND2_X1 U9825 ( .A1(n9560), .A2(n9562), .ZN(n9801) );
  NAND2_X1 U9826 ( .A1(n9638), .A2(n9805), .ZN(n9562) );
  NAND2_X1 U9827 ( .A1(n9637), .A2(n9639), .ZN(n9805) );
  NAND2_X1 U9828 ( .A1(n9806), .A2(n9807), .ZN(n9639) );
  NAND2_X1 U9829 ( .A1(b_27_), .A2(a_22_), .ZN(n9807) );
  INV_X1 U9830 ( .A(n9808), .ZN(n9806) );
  XNOR2_X1 U9831 ( .A(n9809), .B(n9810), .ZN(n9637) );
  NAND2_X1 U9832 ( .A1(n9811), .A2(n9812), .ZN(n9809) );
  NAND2_X1 U9833 ( .A1(a_22_), .A2(n9808), .ZN(n9638) );
  NAND2_X1 U9834 ( .A1(n9574), .A2(n9813), .ZN(n9808) );
  NAND2_X1 U9835 ( .A1(n9573), .A2(n9575), .ZN(n9813) );
  NAND2_X1 U9836 ( .A1(n9814), .A2(n9815), .ZN(n9575) );
  NAND2_X1 U9837 ( .A1(b_27_), .A2(a_23_), .ZN(n9815) );
  XOR2_X1 U9838 ( .A(n9816), .B(n9817), .Z(n9573) );
  XOR2_X1 U9839 ( .A(n9818), .B(n9819), .Z(n9816) );
  NAND2_X1 U9840 ( .A1(a_23_), .A2(n9820), .ZN(n9574) );
  INV_X1 U9841 ( .A(n9814), .ZN(n9820) );
  NOR2_X1 U9842 ( .A1(n9821), .A2(n9822), .ZN(n9814) );
  NOR2_X1 U9843 ( .A1(n9583), .A2(n9823), .ZN(n9822) );
  NOR2_X1 U9844 ( .A1(n9582), .A2(n9580), .ZN(n9823) );
  NAND2_X1 U9845 ( .A1(b_27_), .A2(a_24_), .ZN(n9583) );
  INV_X1 U9846 ( .A(n9824), .ZN(n9821) );
  NAND2_X1 U9847 ( .A1(n9580), .A2(n9582), .ZN(n9824) );
  NAND2_X1 U9848 ( .A1(n9634), .A2(n9825), .ZN(n9582) );
  NAND2_X1 U9849 ( .A1(n9633), .A2(n9635), .ZN(n9825) );
  NAND2_X1 U9850 ( .A1(n9826), .A2(n9827), .ZN(n9635) );
  NAND2_X1 U9851 ( .A1(b_27_), .A2(a_25_), .ZN(n9827) );
  INV_X1 U9852 ( .A(n9828), .ZN(n9826) );
  XNOR2_X1 U9853 ( .A(n9829), .B(n9830), .ZN(n9633) );
  XOR2_X1 U9854 ( .A(n9831), .B(n9832), .Z(n9830) );
  NAND2_X1 U9855 ( .A1(a_25_), .A2(n9828), .ZN(n9634) );
  NAND2_X1 U9856 ( .A1(n9594), .A2(n9833), .ZN(n9828) );
  NAND2_X1 U9857 ( .A1(n9593), .A2(n9595), .ZN(n9833) );
  NAND2_X1 U9858 ( .A1(n9834), .A2(n9835), .ZN(n9595) );
  NAND2_X1 U9859 ( .A1(b_27_), .A2(a_26_), .ZN(n9834) );
  XOR2_X1 U9860 ( .A(n9836), .B(n9837), .Z(n9593) );
  XOR2_X1 U9861 ( .A(n9838), .B(n9839), .Z(n9836) );
  INV_X1 U9862 ( .A(n9840), .ZN(n9594) );
  NOR2_X1 U9863 ( .A1(n9835), .A2(n9344), .ZN(n9840) );
  NAND2_X1 U9864 ( .A1(n9841), .A2(n9842), .ZN(n9835) );
  NAND2_X1 U9865 ( .A1(n9601), .A2(n9843), .ZN(n9842) );
  NAND2_X1 U9866 ( .A1(n9844), .A2(n9602), .ZN(n9843) );
  XNOR2_X1 U9867 ( .A(n9845), .B(n9846), .ZN(n9601) );
  XOR2_X1 U9868 ( .A(n9847), .B(n9848), .Z(n9845) );
  INV_X1 U9869 ( .A(n9849), .ZN(n9841) );
  NOR2_X1 U9870 ( .A1(n9602), .A2(n9844), .ZN(n9849) );
  NAND2_X1 U9871 ( .A1(n9850), .A2(n9851), .ZN(n9602) );
  NAND2_X1 U9872 ( .A1(n9610), .A2(n9852), .ZN(n9851) );
  INV_X1 U9873 ( .A(n9853), .ZN(n9852) );
  NOR2_X1 U9874 ( .A1(n9611), .A2(n9609), .ZN(n9853) );
  NOR2_X1 U9875 ( .A1(n9367), .A2(n8314), .ZN(n9610) );
  NAND2_X1 U9876 ( .A1(n9609), .A2(n9611), .ZN(n9850) );
  NAND2_X1 U9877 ( .A1(n9854), .A2(n9855), .ZN(n9611) );
  NAND2_X1 U9878 ( .A1(n9617), .A2(n9856), .ZN(n9855) );
  INV_X1 U9879 ( .A(n9857), .ZN(n9856) );
  NOR2_X1 U9880 ( .A1(n9618), .A2(n9619), .ZN(n9857) );
  NOR2_X1 U9881 ( .A1(n9367), .A2(n9098), .ZN(n9617) );
  NAND2_X1 U9882 ( .A1(n9619), .A2(n9618), .ZN(n9854) );
  NAND2_X1 U9883 ( .A1(n9858), .A2(n9859), .ZN(n9618) );
  NAND2_X1 U9884 ( .A1(b_25_), .A2(n9860), .ZN(n9859) );
  NAND2_X1 U9885 ( .A1(n8299), .A2(n9861), .ZN(n9860) );
  NAND2_X1 U9886 ( .A1(a_31_), .A2(n9630), .ZN(n9861) );
  NAND2_X1 U9887 ( .A1(b_26_), .A2(n9862), .ZN(n9858) );
  NAND2_X1 U9888 ( .A1(n8303), .A2(n9863), .ZN(n9862) );
  NAND2_X1 U9889 ( .A1(a_30_), .A2(n9864), .ZN(n9863) );
  NOR3_X1 U9890 ( .A1(n9367), .A2(n9631), .A3(n9630), .ZN(n9619) );
  XOR2_X1 U9891 ( .A(n9865), .B(n9866), .Z(n9609) );
  XOR2_X1 U9892 ( .A(n9867), .B(n9868), .Z(n9865) );
  XOR2_X1 U9893 ( .A(n9869), .B(n9870), .Z(n9580) );
  XNOR2_X1 U9894 ( .A(n9871), .B(n9872), .ZN(n9870) );
  XNOR2_X1 U9895 ( .A(n9873), .B(n9874), .ZN(n9560) );
  NAND2_X1 U9896 ( .A1(n9875), .A2(n9876), .ZN(n9873) );
  XNOR2_X1 U9897 ( .A(n9877), .B(n9878), .ZN(n9547) );
  NAND2_X1 U9898 ( .A1(n9879), .A2(n9880), .ZN(n9877) );
  XNOR2_X1 U9899 ( .A(n9881), .B(n9882), .ZN(n9521) );
  NAND2_X1 U9900 ( .A1(n9883), .A2(n9884), .ZN(n9881) );
  XNOR2_X1 U9901 ( .A(n9885), .B(n9886), .ZN(n9508) );
  NAND2_X1 U9902 ( .A1(n9887), .A2(n9888), .ZN(n9885) );
  XNOR2_X1 U9903 ( .A(n9889), .B(n9890), .ZN(n9480) );
  NAND2_X1 U9904 ( .A1(n9891), .A2(n9892), .ZN(n9889) );
  XNOR2_X1 U9905 ( .A(n9893), .B(n9894), .ZN(n9465) );
  XOR2_X1 U9906 ( .A(n9895), .B(n9896), .Z(n9894) );
  NAND2_X1 U9907 ( .A1(b_26_), .A2(a_8_), .ZN(n9896) );
  NAND2_X1 U9908 ( .A1(n9659), .A2(n9897), .ZN(n9705) );
  INV_X1 U9909 ( .A(n9656), .ZN(n9897) );
  XOR2_X1 U9910 ( .A(n9898), .B(n9899), .Z(n9656) );
  XOR2_X1 U9911 ( .A(n9900), .B(n9901), .Z(n9899) );
  NAND2_X1 U9912 ( .A1(b_26_), .A2(a_7_), .ZN(n9901) );
  NOR2_X1 U9913 ( .A1(n9367), .A2(n8430), .ZN(n9659) );
  XNOR2_X1 U9914 ( .A(n9902), .B(n9903), .ZN(n9661) );
  XNOR2_X1 U9915 ( .A(n9904), .B(n9905), .ZN(n9902) );
  XNOR2_X1 U9916 ( .A(n9906), .B(n9907), .ZN(n9665) );
  XNOR2_X1 U9917 ( .A(n9908), .B(n9909), .ZN(n9906) );
  NOR2_X1 U9918 ( .A1(n8938), .A2(n9630), .ZN(n9909) );
  XNOR2_X1 U9919 ( .A(n9910), .B(n9911), .ZN(n9669) );
  XNOR2_X1 U9920 ( .A(n9912), .B(n9913), .ZN(n9910) );
  NOR2_X1 U9921 ( .A1(n8439), .A2(n9630), .ZN(n9913) );
  XNOR2_X1 U9922 ( .A(n9914), .B(n9915), .ZN(n9677) );
  NAND2_X1 U9923 ( .A1(n9916), .A2(n9917), .ZN(n9914) );
  XNOR2_X1 U9924 ( .A(n9918), .B(n9919), .ZN(n9426) );
  XNOR2_X1 U9925 ( .A(n9920), .B(n9921), .ZN(n9919) );
  NAND2_X1 U9926 ( .A1(n9922), .A2(n9923), .ZN(n8485) );
  NAND2_X1 U9927 ( .A1(n8638), .A2(n8637), .ZN(n9923) );
  INV_X1 U9928 ( .A(n9924), .ZN(n9922) );
  NAND3_X1 U9929 ( .A1(n8638), .A2(n8637), .A3(n9924), .ZN(n8484) );
  NOR2_X1 U9930 ( .A1(n9925), .A2(n9926), .ZN(n9924) );
  NOR2_X1 U9931 ( .A1(n9927), .A2(n9928), .ZN(n9926) );
  INV_X1 U9932 ( .A(n8630), .ZN(n9925) );
  NAND2_X1 U9933 ( .A1(n9433), .A2(n9929), .ZN(n8637) );
  NAND2_X1 U9934 ( .A1(n9432), .A2(n9434), .ZN(n9929) );
  NAND2_X1 U9935 ( .A1(n9930), .A2(n9931), .ZN(n9434) );
  INV_X1 U9936 ( .A(n9932), .ZN(n9931) );
  NAND2_X1 U9937 ( .A1(b_26_), .A2(a_0_), .ZN(n9930) );
  XNOR2_X1 U9938 ( .A(n9933), .B(n9934), .ZN(n9432) );
  XNOR2_X1 U9939 ( .A(n9935), .B(n9936), .ZN(n9933) );
  NOR2_X1 U9940 ( .A1(n8569), .A2(n9864), .ZN(n9936) );
  NAND2_X1 U9941 ( .A1(n9932), .A2(a_0_), .ZN(n9433) );
  NOR2_X1 U9942 ( .A1(n9937), .A2(n9938), .ZN(n9932) );
  INV_X1 U9943 ( .A(n9939), .ZN(n9938) );
  NAND2_X1 U9944 ( .A1(n9918), .A2(n9940), .ZN(n9939) );
  NAND2_X1 U9945 ( .A1(n9921), .A2(n9920), .ZN(n9940) );
  XOR2_X1 U9946 ( .A(n9941), .B(n9942), .Z(n9918) );
  XNOR2_X1 U9947 ( .A(n9943), .B(n9944), .ZN(n9941) );
  NOR2_X1 U9948 ( .A1(n8448), .A2(n9864), .ZN(n9944) );
  NOR2_X1 U9949 ( .A1(n9920), .A2(n9921), .ZN(n9937) );
  NOR2_X1 U9950 ( .A1(n9630), .A2(n8569), .ZN(n9921) );
  NAND2_X1 U9951 ( .A1(n9916), .A2(n9945), .ZN(n9920) );
  NAND2_X1 U9952 ( .A1(n9915), .A2(n9917), .ZN(n9945) );
  NAND2_X1 U9953 ( .A1(n9946), .A2(n9947), .ZN(n9917) );
  NAND2_X1 U9954 ( .A1(b_26_), .A2(a_2_), .ZN(n9947) );
  XOR2_X1 U9955 ( .A(n9948), .B(n9949), .Z(n9915) );
  XOR2_X1 U9956 ( .A(n9950), .B(n9951), .Z(n9948) );
  NOR2_X1 U9957 ( .A1(n8900), .A2(n9864), .ZN(n9951) );
  INV_X1 U9958 ( .A(n9952), .ZN(n9916) );
  NOR2_X1 U9959 ( .A1(n8448), .A2(n9946), .ZN(n9952) );
  NOR2_X1 U9960 ( .A1(n9953), .A2(n9954), .ZN(n9946) );
  INV_X1 U9961 ( .A(n9955), .ZN(n9954) );
  NAND3_X1 U9962 ( .A1(a_3_), .A2(n9956), .A3(b_26_), .ZN(n9955) );
  NAND2_X1 U9963 ( .A1(n9691), .A2(n9689), .ZN(n9956) );
  NOR2_X1 U9964 ( .A1(n9689), .A2(n9691), .ZN(n9953) );
  NOR2_X1 U9965 ( .A1(n9957), .A2(n9958), .ZN(n9691) );
  INV_X1 U9966 ( .A(n9959), .ZN(n9958) );
  NAND3_X1 U9967 ( .A1(a_4_), .A2(n9960), .A3(b_26_), .ZN(n9959) );
  NAND2_X1 U9968 ( .A1(n9912), .A2(n9911), .ZN(n9960) );
  NOR2_X1 U9969 ( .A1(n9911), .A2(n9912), .ZN(n9957) );
  NOR2_X1 U9970 ( .A1(n9961), .A2(n9962), .ZN(n9912) );
  INV_X1 U9971 ( .A(n9963), .ZN(n9962) );
  NAND3_X1 U9972 ( .A1(a_5_), .A2(n9964), .A3(b_26_), .ZN(n9963) );
  NAND2_X1 U9973 ( .A1(n9908), .A2(n9907), .ZN(n9964) );
  NOR2_X1 U9974 ( .A1(n9907), .A2(n9908), .ZN(n9961) );
  NOR2_X1 U9975 ( .A1(n9965), .A2(n9966), .ZN(n9908) );
  INV_X1 U9976 ( .A(n9967), .ZN(n9966) );
  NAND2_X1 U9977 ( .A1(n9904), .A2(n9968), .ZN(n9967) );
  NAND2_X1 U9978 ( .A1(n9903), .A2(n9905), .ZN(n9968) );
  NAND2_X1 U9979 ( .A1(n9969), .A2(n9970), .ZN(n9904) );
  INV_X1 U9980 ( .A(n9971), .ZN(n9970) );
  NOR3_X1 U9981 ( .A1(n8425), .A2(n9972), .A3(n9630), .ZN(n9971) );
  NOR2_X1 U9982 ( .A1(n9898), .A2(n9900), .ZN(n9972) );
  NAND2_X1 U9983 ( .A1(n9898), .A2(n9900), .ZN(n9969) );
  NAND2_X1 U9984 ( .A1(n9973), .A2(n9974), .ZN(n9900) );
  NAND3_X1 U9985 ( .A1(a_8_), .A2(n9975), .A3(b_26_), .ZN(n9974) );
  INV_X1 U9986 ( .A(n9976), .ZN(n9975) );
  NOR2_X1 U9987 ( .A1(n9895), .A2(n9893), .ZN(n9976) );
  NAND2_X1 U9988 ( .A1(n9893), .A2(n9895), .ZN(n9973) );
  NAND2_X1 U9989 ( .A1(n9977), .A2(n9978), .ZN(n9895) );
  NAND3_X1 U9990 ( .A1(a_9_), .A2(n9979), .A3(b_26_), .ZN(n9978) );
  INV_X1 U9991 ( .A(n9980), .ZN(n9979) );
  NOR2_X1 U9992 ( .A1(n9719), .A2(n9718), .ZN(n9980) );
  NAND2_X1 U9993 ( .A1(n9718), .A2(n9719), .ZN(n9977) );
  NAND2_X1 U9994 ( .A1(n9891), .A2(n9981), .ZN(n9719) );
  NAND2_X1 U9995 ( .A1(n9890), .A2(n9892), .ZN(n9981) );
  NAND2_X1 U9996 ( .A1(n9982), .A2(n9983), .ZN(n9892) );
  NAND2_X1 U9997 ( .A1(b_26_), .A2(a_10_), .ZN(n9983) );
  INV_X1 U9998 ( .A(n9984), .ZN(n9982) );
  XOR2_X1 U9999 ( .A(n9985), .B(n9986), .Z(n9890) );
  XOR2_X1 U10000 ( .A(n9987), .B(n9988), .Z(n9985) );
  NOR2_X1 U10001 ( .A1(n8867), .A2(n9864), .ZN(n9988) );
  NAND2_X1 U10002 ( .A1(a_10_), .A2(n9984), .ZN(n9891) );
  NAND2_X1 U10003 ( .A1(n9989), .A2(n9990), .ZN(n9984) );
  INV_X1 U10004 ( .A(n9991), .ZN(n9990) );
  NOR3_X1 U10005 ( .A1(n8867), .A2(n9992), .A3(n9630), .ZN(n9991) );
  NOR2_X1 U10006 ( .A1(n9729), .A2(n9730), .ZN(n9992) );
  NAND2_X1 U10007 ( .A1(n9730), .A2(n9729), .ZN(n9989) );
  XNOR2_X1 U10008 ( .A(n9993), .B(n9994), .ZN(n9729) );
  NAND2_X1 U10009 ( .A1(n9995), .A2(n9996), .ZN(n9993) );
  NOR2_X1 U10010 ( .A1(n9997), .A2(n9998), .ZN(n9730) );
  INV_X1 U10011 ( .A(n9999), .ZN(n9998) );
  NAND2_X1 U10012 ( .A1(n9738), .A2(n10000), .ZN(n9999) );
  NAND2_X1 U10013 ( .A1(n9740), .A2(n9739), .ZN(n10000) );
  XNOR2_X1 U10014 ( .A(n10001), .B(n10002), .ZN(n9738) );
  XOR2_X1 U10015 ( .A(n10003), .B(n10004), .Z(n10001) );
  NOR2_X1 U10016 ( .A1(n8996), .A2(n9864), .ZN(n10004) );
  NOR2_X1 U10017 ( .A1(n9739), .A2(n9740), .ZN(n9997) );
  NOR2_X1 U10018 ( .A1(n9630), .A2(n8393), .ZN(n9740) );
  NAND2_X1 U10019 ( .A1(n9746), .A2(n10005), .ZN(n9739) );
  NAND2_X1 U10020 ( .A1(n9745), .A2(n9747), .ZN(n10005) );
  NAND2_X1 U10021 ( .A1(n10006), .A2(n10007), .ZN(n9747) );
  NAND2_X1 U10022 ( .A1(b_26_), .A2(a_13_), .ZN(n10007) );
  INV_X1 U10023 ( .A(n10008), .ZN(n10006) );
  XNOR2_X1 U10024 ( .A(n10009), .B(n10010), .ZN(n9745) );
  NAND2_X1 U10025 ( .A1(n10011), .A2(n10012), .ZN(n10009) );
  NAND2_X1 U10026 ( .A1(a_13_), .A2(n10008), .ZN(n9746) );
  NAND2_X1 U10027 ( .A1(n9887), .A2(n10013), .ZN(n10008) );
  NAND2_X1 U10028 ( .A1(n9886), .A2(n9888), .ZN(n10013) );
  NAND2_X1 U10029 ( .A1(n10014), .A2(n10015), .ZN(n9888) );
  NAND2_X1 U10030 ( .A1(b_26_), .A2(a_14_), .ZN(n10015) );
  XNOR2_X1 U10031 ( .A(n10016), .B(n10017), .ZN(n9886) );
  XOR2_X1 U10032 ( .A(n10018), .B(n10019), .Z(n10017) );
  NAND2_X1 U10033 ( .A1(b_25_), .A2(a_15_), .ZN(n10019) );
  INV_X1 U10034 ( .A(n10020), .ZN(n9887) );
  NOR2_X1 U10035 ( .A1(n9262), .A2(n10014), .ZN(n10020) );
  NOR2_X1 U10036 ( .A1(n10021), .A2(n10022), .ZN(n10014) );
  NOR3_X1 U10037 ( .A1(n8850), .A2(n10023), .A3(n9630), .ZN(n10022) );
  NOR2_X1 U10038 ( .A1(n9758), .A2(n9757), .ZN(n10023) );
  INV_X1 U10039 ( .A(n10024), .ZN(n10021) );
  NAND2_X1 U10040 ( .A1(n9757), .A2(n9758), .ZN(n10024) );
  NAND2_X1 U10041 ( .A1(n9883), .A2(n10025), .ZN(n9758) );
  NAND2_X1 U10042 ( .A1(n9882), .A2(n9884), .ZN(n10025) );
  NAND2_X1 U10043 ( .A1(n10026), .A2(n10027), .ZN(n9884) );
  NAND2_X1 U10044 ( .A1(b_26_), .A2(a_16_), .ZN(n10027) );
  XNOR2_X1 U10045 ( .A(n10028), .B(n10029), .ZN(n9882) );
  XNOR2_X1 U10046 ( .A(n10030), .B(n10031), .ZN(n10029) );
  INV_X1 U10047 ( .A(n10032), .ZN(n9883) );
  NOR2_X1 U10048 ( .A1(n8376), .A2(n10026), .ZN(n10032) );
  NOR2_X1 U10049 ( .A1(n10033), .A2(n10034), .ZN(n10026) );
  NOR3_X1 U10050 ( .A1(n8371), .A2(n10035), .A3(n9630), .ZN(n10034) );
  INV_X1 U10051 ( .A(n10036), .ZN(n10035) );
  NAND2_X1 U10052 ( .A1(n9769), .A2(n9771), .ZN(n10036) );
  NOR2_X1 U10053 ( .A1(n9771), .A2(n9769), .ZN(n10033) );
  XOR2_X1 U10054 ( .A(n10037), .B(n10038), .Z(n9769) );
  XOR2_X1 U10055 ( .A(n10039), .B(n10040), .Z(n10037) );
  NAND2_X1 U10056 ( .A1(n10041), .A2(n10042), .ZN(n9771) );
  NAND2_X1 U10057 ( .A1(n9778), .A2(n10043), .ZN(n10042) );
  NAND2_X1 U10058 ( .A1(n9780), .A2(n9779), .ZN(n10043) );
  XNOR2_X1 U10059 ( .A(n10044), .B(n10045), .ZN(n9778) );
  XOR2_X1 U10060 ( .A(n10046), .B(n10047), .Z(n10044) );
  NOR2_X1 U10061 ( .A1(n8742), .A2(n9864), .ZN(n10047) );
  INV_X1 U10062 ( .A(n10048), .ZN(n10041) );
  NOR2_X1 U10063 ( .A1(n9779), .A2(n9780), .ZN(n10048) );
  NOR2_X1 U10064 ( .A1(n9630), .A2(n9291), .ZN(n9780) );
  NAND2_X1 U10065 ( .A1(n10049), .A2(n10050), .ZN(n9779) );
  NAND3_X1 U10066 ( .A1(a_19_), .A2(n10051), .A3(b_26_), .ZN(n10050) );
  INV_X1 U10067 ( .A(n10052), .ZN(n10051) );
  NOR2_X1 U10068 ( .A1(n9786), .A2(n9785), .ZN(n10052) );
  NAND2_X1 U10069 ( .A1(n9785), .A2(n9786), .ZN(n10049) );
  NAND2_X1 U10070 ( .A1(n9879), .A2(n10053), .ZN(n9786) );
  NAND2_X1 U10071 ( .A1(n9878), .A2(n9880), .ZN(n10053) );
  NAND2_X1 U10072 ( .A1(n10054), .A2(n10055), .ZN(n9880) );
  NAND2_X1 U10073 ( .A1(b_26_), .A2(a_20_), .ZN(n10055) );
  INV_X1 U10074 ( .A(n10056), .ZN(n10054) );
  XNOR2_X1 U10075 ( .A(n10057), .B(n10058), .ZN(n9878) );
  XOR2_X1 U10076 ( .A(n10059), .B(n10060), .Z(n10058) );
  NAND2_X1 U10077 ( .A1(b_25_), .A2(a_21_), .ZN(n10060) );
  NAND2_X1 U10078 ( .A1(a_20_), .A2(n10056), .ZN(n9879) );
  NAND2_X1 U10079 ( .A1(n10061), .A2(n10062), .ZN(n10056) );
  INV_X1 U10080 ( .A(n10063), .ZN(n10062) );
  NOR3_X1 U10081 ( .A1(n8759), .A2(n10064), .A3(n9630), .ZN(n10063) );
  NOR2_X1 U10082 ( .A1(n9799), .A2(n9797), .ZN(n10064) );
  NAND2_X1 U10083 ( .A1(n9797), .A2(n9799), .ZN(n10061) );
  NAND2_X1 U10084 ( .A1(n9875), .A2(n10065), .ZN(n9799) );
  NAND2_X1 U10085 ( .A1(n9874), .A2(n9876), .ZN(n10065) );
  NAND2_X1 U10086 ( .A1(n10066), .A2(n10067), .ZN(n9876) );
  NAND2_X1 U10087 ( .A1(b_26_), .A2(a_22_), .ZN(n10067) );
  INV_X1 U10088 ( .A(n10068), .ZN(n10066) );
  XNOR2_X1 U10089 ( .A(n10069), .B(n10070), .ZN(n9874) );
  NAND2_X1 U10090 ( .A1(n10071), .A2(n10072), .ZN(n10069) );
  NAND2_X1 U10091 ( .A1(a_22_), .A2(n10068), .ZN(n9875) );
  NAND2_X1 U10092 ( .A1(n9811), .A2(n10073), .ZN(n10068) );
  NAND2_X1 U10093 ( .A1(n9810), .A2(n9812), .ZN(n10073) );
  NAND2_X1 U10094 ( .A1(n10074), .A2(n10075), .ZN(n9812) );
  NAND2_X1 U10095 ( .A1(b_26_), .A2(a_23_), .ZN(n10075) );
  INV_X1 U10096 ( .A(n10076), .ZN(n10074) );
  XNOR2_X1 U10097 ( .A(n10077), .B(n10078), .ZN(n9810) );
  XNOR2_X1 U10098 ( .A(n10079), .B(n10080), .ZN(n10078) );
  NAND2_X1 U10099 ( .A1(a_23_), .A2(n10076), .ZN(n9811) );
  NAND2_X1 U10100 ( .A1(n10081), .A2(n10082), .ZN(n10076) );
  NAND2_X1 U10101 ( .A1(n9819), .A2(n10083), .ZN(n10082) );
  INV_X1 U10102 ( .A(n10084), .ZN(n10083) );
  NOR2_X1 U10103 ( .A1(n9818), .A2(n9817), .ZN(n10084) );
  NOR2_X1 U10104 ( .A1(n9630), .A2(n8779), .ZN(n9819) );
  NAND2_X1 U10105 ( .A1(n9817), .A2(n9818), .ZN(n10081) );
  NAND2_X1 U10106 ( .A1(n10085), .A2(n10086), .ZN(n9818) );
  NAND2_X1 U10107 ( .A1(n9872), .A2(n10087), .ZN(n10086) );
  NAND2_X1 U10108 ( .A1(n10088), .A2(n9871), .ZN(n10087) );
  INV_X1 U10109 ( .A(n9869), .ZN(n10088) );
  NOR2_X1 U10110 ( .A1(n9630), .A2(n8788), .ZN(n9872) );
  NAND2_X1 U10111 ( .A1(n10089), .A2(n9869), .ZN(n10085) );
  XOR2_X1 U10112 ( .A(n10090), .B(n10091), .Z(n9869) );
  XNOR2_X1 U10113 ( .A(n10092), .B(n10093), .ZN(n10091) );
  INV_X1 U10114 ( .A(n9871), .ZN(n10089) );
  NAND2_X1 U10115 ( .A1(n10094), .A2(n10095), .ZN(n9871) );
  NAND2_X1 U10116 ( .A1(n10096), .A2(n9831), .ZN(n10095) );
  NAND2_X1 U10117 ( .A1(n9829), .A2(n9832), .ZN(n10096) );
  INV_X1 U10118 ( .A(n10097), .ZN(n10094) );
  NOR2_X1 U10119 ( .A1(n9832), .A2(n9829), .ZN(n10097) );
  XOR2_X1 U10120 ( .A(n10098), .B(n10099), .Z(n9829) );
  XOR2_X1 U10121 ( .A(n10100), .B(n10101), .Z(n10098) );
  NAND2_X1 U10122 ( .A1(n10102), .A2(n10103), .ZN(n9832) );
  NAND2_X1 U10123 ( .A1(n9839), .A2(n10104), .ZN(n10103) );
  INV_X1 U10124 ( .A(n10105), .ZN(n10104) );
  NOR2_X1 U10125 ( .A1(n9838), .A2(n9837), .ZN(n10105) );
  NOR2_X1 U10126 ( .A1(n9630), .A2(n8797), .ZN(n9839) );
  NAND2_X1 U10127 ( .A1(n9837), .A2(n9838), .ZN(n10102) );
  NAND2_X1 U10128 ( .A1(n10106), .A2(n10107), .ZN(n9838) );
  NAND2_X1 U10129 ( .A1(n9847), .A2(n10108), .ZN(n10107) );
  INV_X1 U10130 ( .A(n10109), .ZN(n10108) );
  NOR2_X1 U10131 ( .A1(n9848), .A2(n9846), .ZN(n10109) );
  NOR2_X1 U10132 ( .A1(n9630), .A2(n8314), .ZN(n9847) );
  NAND2_X1 U10133 ( .A1(n9846), .A2(n9848), .ZN(n10106) );
  NAND2_X1 U10134 ( .A1(n10110), .A2(n10111), .ZN(n9848) );
  NAND2_X1 U10135 ( .A1(n9866), .A2(n10112), .ZN(n10111) );
  INV_X1 U10136 ( .A(n10113), .ZN(n10112) );
  NOR2_X1 U10137 ( .A1(n9867), .A2(n9868), .ZN(n10113) );
  NOR2_X1 U10138 ( .A1(n9630), .A2(n9098), .ZN(n9866) );
  NAND2_X1 U10139 ( .A1(n9868), .A2(n9867), .ZN(n10110) );
  NAND2_X1 U10140 ( .A1(n10114), .A2(n10115), .ZN(n9867) );
  NAND2_X1 U10141 ( .A1(b_24_), .A2(n10116), .ZN(n10115) );
  NAND2_X1 U10142 ( .A1(n8299), .A2(n10117), .ZN(n10116) );
  NAND2_X1 U10143 ( .A1(a_31_), .A2(n9864), .ZN(n10117) );
  NAND2_X1 U10144 ( .A1(b_25_), .A2(n10118), .ZN(n10114) );
  NAND2_X1 U10145 ( .A1(n8303), .A2(n10119), .ZN(n10118) );
  NAND2_X1 U10146 ( .A1(a_30_), .A2(n10120), .ZN(n10119) );
  NOR3_X1 U10147 ( .A1(n9864), .A2(n9631), .A3(n9630), .ZN(n9868) );
  XOR2_X1 U10148 ( .A(n10121), .B(n10122), .Z(n9846) );
  XOR2_X1 U10149 ( .A(n10123), .B(n10124), .Z(n10121) );
  XOR2_X1 U10150 ( .A(n10125), .B(n10126), .Z(n9837) );
  XOR2_X1 U10151 ( .A(n10127), .B(n10128), .Z(n10125) );
  XNOR2_X1 U10152 ( .A(n10129), .B(n10130), .ZN(n9817) );
  XNOR2_X1 U10153 ( .A(n10131), .B(n10132), .ZN(n10130) );
  XNOR2_X1 U10154 ( .A(n10133), .B(n10134), .ZN(n9797) );
  NAND2_X1 U10155 ( .A1(n10135), .A2(n10136), .ZN(n10133) );
  XNOR2_X1 U10156 ( .A(n10137), .B(n10138), .ZN(n9785) );
  NAND2_X1 U10157 ( .A1(n10139), .A2(n10140), .ZN(n10137) );
  XNOR2_X1 U10158 ( .A(n10141), .B(n10142), .ZN(n9757) );
  XOR2_X1 U10159 ( .A(n10143), .B(n10144), .Z(n10141) );
  XNOR2_X1 U10160 ( .A(n10145), .B(n10146), .ZN(n9718) );
  XNOR2_X1 U10161 ( .A(n10147), .B(n10148), .ZN(n10146) );
  XOR2_X1 U10162 ( .A(n10149), .B(n10150), .Z(n9893) );
  XOR2_X1 U10163 ( .A(n10151), .B(n10152), .Z(n10149) );
  NOR2_X1 U10164 ( .A1(n8971), .A2(n9864), .ZN(n10152) );
  XNOR2_X1 U10165 ( .A(n10153), .B(n10154), .ZN(n9898) );
  XNOR2_X1 U10166 ( .A(n10155), .B(n10156), .ZN(n10153) );
  NOR2_X1 U10167 ( .A1(n8968), .A2(n9864), .ZN(n10156) );
  NOR2_X1 U10168 ( .A1(n9903), .A2(n9905), .ZN(n9965) );
  NAND2_X1 U10169 ( .A1(b_26_), .A2(a_6_), .ZN(n9905) );
  XNOR2_X1 U10170 ( .A(n10157), .B(n10158), .ZN(n9903) );
  XNOR2_X1 U10171 ( .A(n10159), .B(n10160), .ZN(n10158) );
  NAND2_X1 U10172 ( .A1(b_25_), .A2(a_7_), .ZN(n10160) );
  XOR2_X1 U10173 ( .A(n10161), .B(n10162), .Z(n9907) );
  NAND2_X1 U10174 ( .A1(n10163), .A2(n10164), .ZN(n10161) );
  XOR2_X1 U10175 ( .A(n10165), .B(n10166), .Z(n9911) );
  XOR2_X1 U10176 ( .A(n10167), .B(n10168), .Z(n10166) );
  NAND2_X1 U10177 ( .A1(b_25_), .A2(a_5_), .ZN(n10168) );
  XOR2_X1 U10178 ( .A(n10169), .B(n10170), .Z(n9689) );
  XOR2_X1 U10179 ( .A(n10171), .B(n10172), .Z(n10170) );
  NAND2_X1 U10180 ( .A1(b_25_), .A2(a_4_), .ZN(n10172) );
  XOR2_X1 U10181 ( .A(n10173), .B(n10174), .Z(n8638) );
  XNOR2_X1 U10182 ( .A(n10175), .B(n10176), .ZN(n10174) );
  NAND2_X1 U10183 ( .A1(b_25_), .A2(a_0_), .ZN(n10176) );
  INV_X1 U10184 ( .A(n10177), .ZN(n8488) );
  NOR2_X1 U10185 ( .A1(n8630), .A2(n8629), .ZN(n10177) );
  XNOR2_X1 U10186 ( .A(n8627), .B(n8626), .ZN(n8629) );
  NAND2_X1 U10187 ( .A1(n9928), .A2(n9927), .ZN(n8630) );
  NAND2_X1 U10188 ( .A1(n10178), .A2(n10179), .ZN(n9927) );
  NAND3_X1 U10189 ( .A1(a_0_), .A2(n10180), .A3(b_25_), .ZN(n10179) );
  NAND2_X1 U10190 ( .A1(n10175), .A2(n10173), .ZN(n10180) );
  INV_X1 U10191 ( .A(n10181), .ZN(n10178) );
  NOR2_X1 U10192 ( .A1(n10173), .A2(n10175), .ZN(n10181) );
  NOR2_X1 U10193 ( .A1(n10182), .A2(n10183), .ZN(n10175) );
  INV_X1 U10194 ( .A(n10184), .ZN(n10183) );
  NAND3_X1 U10195 ( .A1(a_1_), .A2(n10185), .A3(b_25_), .ZN(n10184) );
  NAND2_X1 U10196 ( .A1(n9935), .A2(n9934), .ZN(n10185) );
  NOR2_X1 U10197 ( .A1(n9934), .A2(n9935), .ZN(n10182) );
  NOR2_X1 U10198 ( .A1(n10186), .A2(n10187), .ZN(n9935) );
  INV_X1 U10199 ( .A(n10188), .ZN(n10187) );
  NAND3_X1 U10200 ( .A1(a_2_), .A2(n10189), .A3(b_25_), .ZN(n10188) );
  NAND2_X1 U10201 ( .A1(n9943), .A2(n9942), .ZN(n10189) );
  NOR2_X1 U10202 ( .A1(n9942), .A2(n9943), .ZN(n10186) );
  NOR2_X1 U10203 ( .A1(n10190), .A2(n10191), .ZN(n9943) );
  NOR3_X1 U10204 ( .A1(n8900), .A2(n10192), .A3(n9864), .ZN(n10191) );
  NOR2_X1 U10205 ( .A1(n9950), .A2(n9949), .ZN(n10192) );
  INV_X1 U10206 ( .A(n10193), .ZN(n10190) );
  NAND2_X1 U10207 ( .A1(n9949), .A2(n9950), .ZN(n10193) );
  NAND2_X1 U10208 ( .A1(n10194), .A2(n10195), .ZN(n9950) );
  NAND3_X1 U10209 ( .A1(a_4_), .A2(n10196), .A3(b_25_), .ZN(n10195) );
  INV_X1 U10210 ( .A(n10197), .ZN(n10196) );
  NOR2_X1 U10211 ( .A1(n10171), .A2(n10169), .ZN(n10197) );
  NAND2_X1 U10212 ( .A1(n10169), .A2(n10171), .ZN(n10194) );
  NAND2_X1 U10213 ( .A1(n10198), .A2(n10199), .ZN(n10171) );
  NAND3_X1 U10214 ( .A1(a_5_), .A2(n10200), .A3(b_25_), .ZN(n10199) );
  INV_X1 U10215 ( .A(n10201), .ZN(n10200) );
  NOR2_X1 U10216 ( .A1(n10167), .A2(n10165), .ZN(n10201) );
  NAND2_X1 U10217 ( .A1(n10165), .A2(n10167), .ZN(n10198) );
  NAND2_X1 U10218 ( .A1(n10163), .A2(n10202), .ZN(n10167) );
  NAND2_X1 U10219 ( .A1(n10162), .A2(n10164), .ZN(n10202) );
  NAND2_X1 U10220 ( .A1(n10203), .A2(n10204), .ZN(n10164) );
  NAND2_X1 U10221 ( .A1(b_25_), .A2(a_6_), .ZN(n10204) );
  XNOR2_X1 U10222 ( .A(n10205), .B(n10206), .ZN(n10162) );
  NAND2_X1 U10223 ( .A1(n10207), .A2(n10208), .ZN(n10205) );
  INV_X1 U10224 ( .A(n10209), .ZN(n10163) );
  NOR2_X1 U10225 ( .A1(n8430), .A2(n10203), .ZN(n10209) );
  NOR2_X1 U10226 ( .A1(n10210), .A2(n10211), .ZN(n10203) );
  INV_X1 U10227 ( .A(n10212), .ZN(n10211) );
  NAND3_X1 U10228 ( .A1(a_7_), .A2(n10213), .A3(b_25_), .ZN(n10212) );
  NAND2_X1 U10229 ( .A1(n10159), .A2(n10157), .ZN(n10213) );
  NOR2_X1 U10230 ( .A1(n10157), .A2(n10159), .ZN(n10210) );
  NOR2_X1 U10231 ( .A1(n10214), .A2(n10215), .ZN(n10159) );
  INV_X1 U10232 ( .A(n10216), .ZN(n10215) );
  NAND3_X1 U10233 ( .A1(a_8_), .A2(n10217), .A3(b_25_), .ZN(n10216) );
  NAND2_X1 U10234 ( .A1(n10155), .A2(n10154), .ZN(n10217) );
  NOR2_X1 U10235 ( .A1(n10154), .A2(n10155), .ZN(n10214) );
  NOR2_X1 U10236 ( .A1(n10218), .A2(n10219), .ZN(n10155) );
  NOR3_X1 U10237 ( .A1(n8971), .A2(n10220), .A3(n9864), .ZN(n10219) );
  NOR2_X1 U10238 ( .A1(n10151), .A2(n10150), .ZN(n10220) );
  INV_X1 U10239 ( .A(n10221), .ZN(n10218) );
  NAND2_X1 U10240 ( .A1(n10150), .A2(n10151), .ZN(n10221) );
  NAND2_X1 U10241 ( .A1(n10222), .A2(n10223), .ZN(n10151) );
  NAND2_X1 U10242 ( .A1(n10147), .A2(n10224), .ZN(n10223) );
  NAND2_X1 U10243 ( .A1(n10225), .A2(n10226), .ZN(n10224) );
  INV_X1 U10244 ( .A(n10148), .ZN(n10226) );
  INV_X1 U10245 ( .A(n10145), .ZN(n10225) );
  NAND2_X1 U10246 ( .A1(n10227), .A2(n10228), .ZN(n10147) );
  INV_X1 U10247 ( .A(n10229), .ZN(n10228) );
  NOR3_X1 U10248 ( .A1(n8867), .A2(n10230), .A3(n9864), .ZN(n10229) );
  NOR2_X1 U10249 ( .A1(n9987), .A2(n9986), .ZN(n10230) );
  NAND2_X1 U10250 ( .A1(n9986), .A2(n9987), .ZN(n10227) );
  NAND2_X1 U10251 ( .A1(n9995), .A2(n10231), .ZN(n9987) );
  NAND2_X1 U10252 ( .A1(n9994), .A2(n9996), .ZN(n10231) );
  NAND2_X1 U10253 ( .A1(n10232), .A2(n10233), .ZN(n9996) );
  NAND2_X1 U10254 ( .A1(b_25_), .A2(a_12_), .ZN(n10233) );
  XOR2_X1 U10255 ( .A(n10234), .B(n10235), .Z(n9994) );
  XOR2_X1 U10256 ( .A(n10236), .B(n10237), .Z(n10234) );
  NOR2_X1 U10257 ( .A1(n8996), .A2(n10120), .ZN(n10237) );
  INV_X1 U10258 ( .A(n10238), .ZN(n9995) );
  NOR2_X1 U10259 ( .A1(n8393), .A2(n10232), .ZN(n10238) );
  NOR2_X1 U10260 ( .A1(n10239), .A2(n10240), .ZN(n10232) );
  NOR3_X1 U10261 ( .A1(n8996), .A2(n10241), .A3(n9864), .ZN(n10240) );
  NOR2_X1 U10262 ( .A1(n10003), .A2(n10002), .ZN(n10241) );
  INV_X1 U10263 ( .A(n10242), .ZN(n10239) );
  NAND2_X1 U10264 ( .A1(n10002), .A2(n10003), .ZN(n10242) );
  NAND2_X1 U10265 ( .A1(n10011), .A2(n10243), .ZN(n10003) );
  NAND2_X1 U10266 ( .A1(n10010), .A2(n10012), .ZN(n10243) );
  NAND2_X1 U10267 ( .A1(n10244), .A2(n10245), .ZN(n10012) );
  NAND2_X1 U10268 ( .A1(b_25_), .A2(a_14_), .ZN(n10245) );
  INV_X1 U10269 ( .A(n10246), .ZN(n10244) );
  XNOR2_X1 U10270 ( .A(n10247), .B(n10248), .ZN(n10010) );
  XOR2_X1 U10271 ( .A(n10249), .B(n10250), .Z(n10248) );
  NAND2_X1 U10272 ( .A1(b_24_), .A2(a_15_), .ZN(n10250) );
  NAND2_X1 U10273 ( .A1(a_14_), .A2(n10246), .ZN(n10011) );
  NAND2_X1 U10274 ( .A1(n10251), .A2(n10252), .ZN(n10246) );
  NAND3_X1 U10275 ( .A1(a_15_), .A2(n10253), .A3(b_25_), .ZN(n10252) );
  NAND2_X1 U10276 ( .A1(n10016), .A2(n10018), .ZN(n10253) );
  INV_X1 U10277 ( .A(n10254), .ZN(n10251) );
  NOR2_X1 U10278 ( .A1(n10018), .A2(n10016), .ZN(n10254) );
  XNOR2_X1 U10279 ( .A(n10255), .B(n10256), .ZN(n10016) );
  XNOR2_X1 U10280 ( .A(n10257), .B(n10258), .ZN(n10256) );
  NAND2_X1 U10281 ( .A1(n10259), .A2(n10260), .ZN(n10018) );
  NAND2_X1 U10282 ( .A1(n10142), .A2(n10261), .ZN(n10260) );
  NAND2_X1 U10283 ( .A1(n10144), .A2(n10143), .ZN(n10261) );
  XOR2_X1 U10284 ( .A(n10262), .B(n10263), .Z(n10142) );
  NAND2_X1 U10285 ( .A1(n10264), .A2(n10265), .ZN(n10262) );
  INV_X1 U10286 ( .A(n10266), .ZN(n10259) );
  NOR2_X1 U10287 ( .A1(n10143), .A2(n10144), .ZN(n10266) );
  NOR2_X1 U10288 ( .A1(n9864), .A2(n8376), .ZN(n10144) );
  NAND2_X1 U10289 ( .A1(n10267), .A2(n10268), .ZN(n10143) );
  NAND2_X1 U10290 ( .A1(n10031), .A2(n10269), .ZN(n10268) );
  NAND2_X1 U10291 ( .A1(n10028), .A2(n10030), .ZN(n10269) );
  NOR2_X1 U10292 ( .A1(n9864), .A2(n8371), .ZN(n10031) );
  INV_X1 U10293 ( .A(n10270), .ZN(n10267) );
  NOR2_X1 U10294 ( .A1(n10030), .A2(n10028), .ZN(n10270) );
  XNOR2_X1 U10295 ( .A(n10271), .B(n10272), .ZN(n10028) );
  XNOR2_X1 U10296 ( .A(n10273), .B(n10274), .ZN(n10272) );
  NAND2_X1 U10297 ( .A1(n10275), .A2(n10276), .ZN(n10030) );
  NAND2_X1 U10298 ( .A1(n10038), .A2(n10277), .ZN(n10276) );
  NAND2_X1 U10299 ( .A1(n10040), .A2(n10039), .ZN(n10277) );
  XNOR2_X1 U10300 ( .A(n10278), .B(n10279), .ZN(n10038) );
  XOR2_X1 U10301 ( .A(n10280), .B(n10281), .Z(n10278) );
  NOR2_X1 U10302 ( .A1(n8742), .A2(n10120), .ZN(n10281) );
  INV_X1 U10303 ( .A(n10282), .ZN(n10275) );
  NOR2_X1 U10304 ( .A1(n10039), .A2(n10040), .ZN(n10282) );
  NOR2_X1 U10305 ( .A1(n9864), .A2(n9291), .ZN(n10040) );
  NAND2_X1 U10306 ( .A1(n10283), .A2(n10284), .ZN(n10039) );
  NAND3_X1 U10307 ( .A1(a_19_), .A2(n10285), .A3(b_25_), .ZN(n10284) );
  INV_X1 U10308 ( .A(n10286), .ZN(n10285) );
  NOR2_X1 U10309 ( .A1(n10046), .A2(n10045), .ZN(n10286) );
  NAND2_X1 U10310 ( .A1(n10045), .A2(n10046), .ZN(n10283) );
  NAND2_X1 U10311 ( .A1(n10139), .A2(n10287), .ZN(n10046) );
  NAND2_X1 U10312 ( .A1(n10138), .A2(n10140), .ZN(n10287) );
  NAND2_X1 U10313 ( .A1(n10288), .A2(n10289), .ZN(n10140) );
  NAND2_X1 U10314 ( .A1(b_25_), .A2(a_20_), .ZN(n10289) );
  INV_X1 U10315 ( .A(n10290), .ZN(n10288) );
  XOR2_X1 U10316 ( .A(n10291), .B(n10292), .Z(n10138) );
  XOR2_X1 U10317 ( .A(n10293), .B(n10294), .Z(n10291) );
  NOR2_X1 U10318 ( .A1(n8759), .A2(n10120), .ZN(n10294) );
  NAND2_X1 U10319 ( .A1(a_20_), .A2(n10290), .ZN(n10139) );
  NAND2_X1 U10320 ( .A1(n10295), .A2(n10296), .ZN(n10290) );
  INV_X1 U10321 ( .A(n10297), .ZN(n10296) );
  NOR3_X1 U10322 ( .A1(n8759), .A2(n10298), .A3(n9864), .ZN(n10297) );
  NOR2_X1 U10323 ( .A1(n10059), .A2(n10057), .ZN(n10298) );
  NAND2_X1 U10324 ( .A1(n10057), .A2(n10059), .ZN(n10295) );
  NAND2_X1 U10325 ( .A1(n10135), .A2(n10299), .ZN(n10059) );
  NAND2_X1 U10326 ( .A1(n10134), .A2(n10136), .ZN(n10299) );
  NAND2_X1 U10327 ( .A1(n10300), .A2(n10301), .ZN(n10136) );
  NAND2_X1 U10328 ( .A1(b_25_), .A2(a_22_), .ZN(n10301) );
  INV_X1 U10329 ( .A(n10302), .ZN(n10300) );
  XNOR2_X1 U10330 ( .A(n10303), .B(n10304), .ZN(n10134) );
  NAND2_X1 U10331 ( .A1(n10305), .A2(n10306), .ZN(n10303) );
  NAND2_X1 U10332 ( .A1(a_22_), .A2(n10302), .ZN(n10135) );
  NAND2_X1 U10333 ( .A1(n10071), .A2(n10307), .ZN(n10302) );
  NAND2_X1 U10334 ( .A1(n10070), .A2(n10072), .ZN(n10307) );
  NAND2_X1 U10335 ( .A1(n10308), .A2(n10309), .ZN(n10072) );
  NAND2_X1 U10336 ( .A1(b_25_), .A2(a_23_), .ZN(n10309) );
  XOR2_X1 U10337 ( .A(n10310), .B(n10311), .Z(n10070) );
  XNOR2_X1 U10338 ( .A(n10312), .B(n10313), .ZN(n10310) );
  NAND2_X1 U10339 ( .A1(a_23_), .A2(n10314), .ZN(n10071) );
  INV_X1 U10340 ( .A(n10308), .ZN(n10314) );
  NOR2_X1 U10341 ( .A1(n10315), .A2(n10316), .ZN(n10308) );
  INV_X1 U10342 ( .A(n10317), .ZN(n10316) );
  NAND2_X1 U10343 ( .A1(n10080), .A2(n10318), .ZN(n10317) );
  NAND2_X1 U10344 ( .A1(n10077), .A2(n10079), .ZN(n10318) );
  NOR2_X1 U10345 ( .A1(n9864), .A2(n8779), .ZN(n10080) );
  NOR2_X1 U10346 ( .A1(n10079), .A2(n10077), .ZN(n10315) );
  XOR2_X1 U10347 ( .A(n10319), .B(n10320), .Z(n10077) );
  XNOR2_X1 U10348 ( .A(n10321), .B(n10322), .ZN(n10320) );
  NAND2_X1 U10349 ( .A1(n10323), .A2(n10324), .ZN(n10079) );
  NAND2_X1 U10350 ( .A1(n10129), .A2(n10325), .ZN(n10324) );
  NAND2_X1 U10351 ( .A1(n10131), .A2(n10326), .ZN(n10325) );
  XNOR2_X1 U10352 ( .A(n10327), .B(n10328), .ZN(n10129) );
  XNOR2_X1 U10353 ( .A(n10329), .B(n10330), .ZN(n10328) );
  NAND2_X1 U10354 ( .A1(n10132), .A2(n10331), .ZN(n10323) );
  INV_X1 U10355 ( .A(n10131), .ZN(n10331) );
  NOR2_X1 U10356 ( .A1(n10332), .A2(n10333), .ZN(n10131) );
  INV_X1 U10357 ( .A(n10334), .ZN(n10333) );
  NAND2_X1 U10358 ( .A1(n10090), .A2(n10335), .ZN(n10334) );
  NAND2_X1 U10359 ( .A1(n10093), .A2(n10092), .ZN(n10335) );
  XNOR2_X1 U10360 ( .A(n10336), .B(n10337), .ZN(n10090) );
  XOR2_X1 U10361 ( .A(n10338), .B(n10339), .Z(n10336) );
  NOR2_X1 U10362 ( .A1(n10092), .A2(n10093), .ZN(n10332) );
  NOR2_X1 U10363 ( .A1(n9864), .A2(n9344), .ZN(n10093) );
  NAND2_X1 U10364 ( .A1(n10340), .A2(n10341), .ZN(n10092) );
  NAND2_X1 U10365 ( .A1(n10101), .A2(n10342), .ZN(n10341) );
  INV_X1 U10366 ( .A(n10343), .ZN(n10342) );
  NOR2_X1 U10367 ( .A1(n10100), .A2(n10099), .ZN(n10343) );
  NOR2_X1 U10368 ( .A1(n9864), .A2(n8797), .ZN(n10101) );
  NAND2_X1 U10369 ( .A1(n10099), .A2(n10100), .ZN(n10340) );
  NAND2_X1 U10370 ( .A1(n10344), .A2(n10345), .ZN(n10100) );
  NAND2_X1 U10371 ( .A1(n10127), .A2(n10346), .ZN(n10345) );
  INV_X1 U10372 ( .A(n10347), .ZN(n10346) );
  NOR2_X1 U10373 ( .A1(n10128), .A2(n10126), .ZN(n10347) );
  NOR2_X1 U10374 ( .A1(n9864), .A2(n8314), .ZN(n10127) );
  NAND2_X1 U10375 ( .A1(n10126), .A2(n10128), .ZN(n10344) );
  NAND2_X1 U10376 ( .A1(n10348), .A2(n10349), .ZN(n10128) );
  NAND2_X1 U10377 ( .A1(n10122), .A2(n10350), .ZN(n10349) );
  INV_X1 U10378 ( .A(n10351), .ZN(n10350) );
  NOR2_X1 U10379 ( .A1(n10123), .A2(n10124), .ZN(n10351) );
  NOR2_X1 U10380 ( .A1(n9864), .A2(n9098), .ZN(n10122) );
  NAND2_X1 U10381 ( .A1(n10124), .A2(n10123), .ZN(n10348) );
  NAND2_X1 U10382 ( .A1(n10352), .A2(n10353), .ZN(n10123) );
  NAND2_X1 U10383 ( .A1(b_23_), .A2(n10354), .ZN(n10353) );
  NAND2_X1 U10384 ( .A1(n8299), .A2(n10355), .ZN(n10354) );
  NAND2_X1 U10385 ( .A1(a_31_), .A2(n10120), .ZN(n10355) );
  NAND2_X1 U10386 ( .A1(b_24_), .A2(n10356), .ZN(n10352) );
  NAND2_X1 U10387 ( .A1(n8303), .A2(n10357), .ZN(n10356) );
  NAND2_X1 U10388 ( .A1(a_30_), .A2(n10358), .ZN(n10357) );
  NOR3_X1 U10389 ( .A1(n10120), .A2(n9631), .A3(n9864), .ZN(n10124) );
  XOR2_X1 U10390 ( .A(n10359), .B(n10360), .Z(n10126) );
  XOR2_X1 U10391 ( .A(n10361), .B(n10362), .Z(n10359) );
  XOR2_X1 U10392 ( .A(n10363), .B(n10364), .Z(n10099) );
  XOR2_X1 U10393 ( .A(n10365), .B(n10366), .Z(n10363) );
  XNOR2_X1 U10394 ( .A(n10367), .B(n10368), .ZN(n10057) );
  NAND2_X1 U10395 ( .A1(n10369), .A2(n10370), .ZN(n10367) );
  XNOR2_X1 U10396 ( .A(n10371), .B(n10372), .ZN(n10045) );
  NAND2_X1 U10397 ( .A1(n10373), .A2(n10374), .ZN(n10371) );
  XNOR2_X1 U10398 ( .A(n10375), .B(n10376), .ZN(n10002) );
  NAND2_X1 U10399 ( .A1(n10377), .A2(n10378), .ZN(n10375) );
  XOR2_X1 U10400 ( .A(n10379), .B(n10380), .Z(n9986) );
  XNOR2_X1 U10401 ( .A(n10381), .B(n10382), .ZN(n10380) );
  NAND2_X1 U10402 ( .A1(b_24_), .A2(a_12_), .ZN(n10382) );
  NAND2_X1 U10403 ( .A1(n10148), .A2(n10145), .ZN(n10222) );
  XNOR2_X1 U10404 ( .A(n10383), .B(n10384), .ZN(n10145) );
  NAND2_X1 U10405 ( .A1(n10385), .A2(n10386), .ZN(n10383) );
  NOR2_X1 U10406 ( .A1(n9864), .A2(n8402), .ZN(n10148) );
  XNOR2_X1 U10407 ( .A(n10387), .B(n10388), .ZN(n10150) );
  NAND2_X1 U10408 ( .A1(n10389), .A2(n10390), .ZN(n10387) );
  XNOR2_X1 U10409 ( .A(n10391), .B(n10392), .ZN(n10154) );
  XOR2_X1 U10410 ( .A(n10393), .B(n10394), .Z(n10391) );
  NOR2_X1 U10411 ( .A1(n8971), .A2(n10120), .ZN(n10394) );
  XNOR2_X1 U10412 ( .A(n10395), .B(n10396), .ZN(n10157) );
  XNOR2_X1 U10413 ( .A(n10397), .B(n10398), .ZN(n10396) );
  NAND2_X1 U10414 ( .A1(b_24_), .A2(a_8_), .ZN(n10398) );
  XNOR2_X1 U10415 ( .A(n10399), .B(n10400), .ZN(n10165) );
  XNOR2_X1 U10416 ( .A(n10401), .B(n10402), .ZN(n10399) );
  XNOR2_X1 U10417 ( .A(n10403), .B(n10404), .ZN(n10169) );
  XNOR2_X1 U10418 ( .A(n10405), .B(n10406), .ZN(n10403) );
  XOR2_X1 U10419 ( .A(n10407), .B(n10408), .Z(n9949) );
  XOR2_X1 U10420 ( .A(n10409), .B(n10410), .Z(n10407) );
  NOR2_X1 U10421 ( .A1(n8439), .A2(n10120), .ZN(n10410) );
  XNOR2_X1 U10422 ( .A(n10411), .B(n10412), .ZN(n9942) );
  XOR2_X1 U10423 ( .A(n10413), .B(n10414), .Z(n10411) );
  XNOR2_X1 U10424 ( .A(n10415), .B(n10416), .ZN(n9934) );
  XOR2_X1 U10425 ( .A(n10417), .B(n10418), .Z(n10415) );
  NOR2_X1 U10426 ( .A1(n8448), .A2(n10120), .ZN(n10418) );
  XNOR2_X1 U10427 ( .A(n10419), .B(n10420), .ZN(n10173) );
  XOR2_X1 U10428 ( .A(n10421), .B(n10422), .Z(n10420) );
  XNOR2_X1 U10429 ( .A(n10423), .B(n10424), .ZN(n9928) );
  XNOR2_X1 U10430 ( .A(n10425), .B(n10426), .ZN(n10424) );
  NAND3_X1 U10431 ( .A1(n8626), .A2(n8627), .A3(n10427), .ZN(n8492) );
  INV_X1 U10432 ( .A(n8624), .ZN(n10427) );
  NAND2_X1 U10433 ( .A1(n8620), .A2(n10428), .ZN(n8624) );
  NAND2_X1 U10434 ( .A1(n10429), .A2(n10430), .ZN(n10428) );
  INV_X1 U10435 ( .A(n8618), .ZN(n8620) );
  NOR2_X1 U10436 ( .A1(n10430), .A2(n10429), .ZN(n8618) );
  NOR2_X1 U10437 ( .A1(n10431), .A2(n10432), .ZN(n10429) );
  INV_X1 U10438 ( .A(n10433), .ZN(n10432) );
  NAND3_X1 U10439 ( .A1(a_0_), .A2(n10434), .A3(b_23_), .ZN(n10433) );
  NAND2_X1 U10440 ( .A1(n10435), .A2(n10436), .ZN(n10434) );
  NOR2_X1 U10441 ( .A1(n10436), .A2(n10435), .ZN(n10431) );
  XOR2_X1 U10442 ( .A(n10437), .B(n10438), .Z(n10430) );
  NAND2_X1 U10443 ( .A1(n10439), .A2(n10440), .ZN(n10437) );
  NAND2_X1 U10444 ( .A1(n10441), .A2(n10442), .ZN(n8627) );
  INV_X1 U10445 ( .A(n10443), .ZN(n10442) );
  NOR2_X1 U10446 ( .A1(n10444), .A2(n10445), .ZN(n10443) );
  NOR2_X1 U10447 ( .A1(n10425), .A2(n10423), .ZN(n10445) );
  INV_X1 U10448 ( .A(n10426), .ZN(n10444) );
  NOR2_X1 U10449 ( .A1(n10120), .A2(n8457), .ZN(n10426) );
  NAND2_X1 U10450 ( .A1(n10423), .A2(n10425), .ZN(n10441) );
  NAND2_X1 U10451 ( .A1(n10446), .A2(n10447), .ZN(n10425) );
  NAND2_X1 U10452 ( .A1(n10421), .A2(n10448), .ZN(n10447) );
  NAND2_X1 U10453 ( .A1(n10419), .A2(n10422), .ZN(n10448) );
  NAND2_X1 U10454 ( .A1(n10449), .A2(n10450), .ZN(n10421) );
  INV_X1 U10455 ( .A(n10451), .ZN(n10450) );
  NOR3_X1 U10456 ( .A1(n8448), .A2(n10452), .A3(n10120), .ZN(n10451) );
  NOR2_X1 U10457 ( .A1(n10417), .A2(n10416), .ZN(n10452) );
  NAND2_X1 U10458 ( .A1(n10416), .A2(n10417), .ZN(n10449) );
  NAND2_X1 U10459 ( .A1(n10453), .A2(n10454), .ZN(n10417) );
  NAND2_X1 U10460 ( .A1(n10413), .A2(n10455), .ZN(n10454) );
  INV_X1 U10461 ( .A(n10456), .ZN(n10455) );
  NOR2_X1 U10462 ( .A1(n10412), .A2(n10414), .ZN(n10456) );
  NAND2_X1 U10463 ( .A1(n10457), .A2(n10458), .ZN(n10413) );
  INV_X1 U10464 ( .A(n10459), .ZN(n10458) );
  NOR3_X1 U10465 ( .A1(n8439), .A2(n10460), .A3(n10120), .ZN(n10459) );
  NOR2_X1 U10466 ( .A1(n10409), .A2(n10408), .ZN(n10460) );
  NAND2_X1 U10467 ( .A1(n10408), .A2(n10409), .ZN(n10457) );
  NAND2_X1 U10468 ( .A1(n10461), .A2(n10462), .ZN(n10409) );
  NAND2_X1 U10469 ( .A1(n10406), .A2(n10463), .ZN(n10462) );
  NAND2_X1 U10470 ( .A1(n10405), .A2(n10404), .ZN(n10463) );
  NOR2_X1 U10471 ( .A1(n10120), .A2(n8938), .ZN(n10406) );
  INV_X1 U10472 ( .A(n10464), .ZN(n10461) );
  NOR2_X1 U10473 ( .A1(n10404), .A2(n10405), .ZN(n10464) );
  NOR2_X1 U10474 ( .A1(n10465), .A2(n10466), .ZN(n10405) );
  INV_X1 U10475 ( .A(n10467), .ZN(n10466) );
  NAND2_X1 U10476 ( .A1(n10402), .A2(n10468), .ZN(n10467) );
  NAND2_X1 U10477 ( .A1(n10401), .A2(n10400), .ZN(n10468) );
  NOR2_X1 U10478 ( .A1(n10120), .A2(n8430), .ZN(n10402) );
  NOR2_X1 U10479 ( .A1(n10400), .A2(n10401), .ZN(n10465) );
  INV_X1 U10480 ( .A(n10469), .ZN(n10401) );
  NAND2_X1 U10481 ( .A1(n10207), .A2(n10470), .ZN(n10469) );
  NAND2_X1 U10482 ( .A1(n10206), .A2(n10208), .ZN(n10470) );
  NAND2_X1 U10483 ( .A1(n10471), .A2(n10472), .ZN(n10208) );
  NAND2_X1 U10484 ( .A1(b_24_), .A2(a_7_), .ZN(n10472) );
  INV_X1 U10485 ( .A(n10473), .ZN(n10471) );
  XOR2_X1 U10486 ( .A(n10474), .B(n10475), .Z(n10206) );
  XNOR2_X1 U10487 ( .A(n10476), .B(n10477), .ZN(n10475) );
  NAND2_X1 U10488 ( .A1(a_7_), .A2(n10473), .ZN(n10207) );
  NAND2_X1 U10489 ( .A1(n10478), .A2(n10479), .ZN(n10473) );
  NAND3_X1 U10490 ( .A1(a_8_), .A2(n10480), .A3(b_24_), .ZN(n10479) );
  NAND2_X1 U10491 ( .A1(n10397), .A2(n10395), .ZN(n10480) );
  INV_X1 U10492 ( .A(n10481), .ZN(n10478) );
  NOR2_X1 U10493 ( .A1(n10395), .A2(n10397), .ZN(n10481) );
  NOR2_X1 U10494 ( .A1(n10482), .A2(n10483), .ZN(n10397) );
  NOR3_X1 U10495 ( .A1(n8971), .A2(n10484), .A3(n10120), .ZN(n10483) );
  NOR2_X1 U10496 ( .A1(n10393), .A2(n10392), .ZN(n10484) );
  INV_X1 U10497 ( .A(n10485), .ZN(n10482) );
  NAND2_X1 U10498 ( .A1(n10392), .A2(n10393), .ZN(n10485) );
  NAND2_X1 U10499 ( .A1(n10389), .A2(n10486), .ZN(n10393) );
  NAND2_X1 U10500 ( .A1(n10388), .A2(n10390), .ZN(n10486) );
  NAND2_X1 U10501 ( .A1(n10487), .A2(n10488), .ZN(n10390) );
  NAND2_X1 U10502 ( .A1(b_24_), .A2(a_10_), .ZN(n10488) );
  INV_X1 U10503 ( .A(n10489), .ZN(n10487) );
  XNOR2_X1 U10504 ( .A(n10490), .B(n10491), .ZN(n10388) );
  XOR2_X1 U10505 ( .A(n10492), .B(n10493), .Z(n10491) );
  NAND2_X1 U10506 ( .A1(b_23_), .A2(a_11_), .ZN(n10493) );
  NAND2_X1 U10507 ( .A1(a_10_), .A2(n10489), .ZN(n10389) );
  NAND2_X1 U10508 ( .A1(n10385), .A2(n10494), .ZN(n10489) );
  NAND2_X1 U10509 ( .A1(n10384), .A2(n10386), .ZN(n10494) );
  NAND2_X1 U10510 ( .A1(n10495), .A2(n10496), .ZN(n10386) );
  NAND2_X1 U10511 ( .A1(b_24_), .A2(a_11_), .ZN(n10496) );
  XOR2_X1 U10512 ( .A(n10497), .B(n10498), .Z(n10384) );
  XNOR2_X1 U10513 ( .A(n10499), .B(n10500), .ZN(n10498) );
  INV_X1 U10514 ( .A(n10501), .ZN(n10385) );
  NOR2_X1 U10515 ( .A1(n8867), .A2(n10495), .ZN(n10501) );
  NOR2_X1 U10516 ( .A1(n10502), .A2(n10503), .ZN(n10495) );
  INV_X1 U10517 ( .A(n10504), .ZN(n10503) );
  NAND3_X1 U10518 ( .A1(a_12_), .A2(n10505), .A3(b_24_), .ZN(n10504) );
  NAND2_X1 U10519 ( .A1(n10381), .A2(n10379), .ZN(n10505) );
  NOR2_X1 U10520 ( .A1(n10379), .A2(n10381), .ZN(n10502) );
  NOR2_X1 U10521 ( .A1(n10506), .A2(n10507), .ZN(n10381) );
  NOR3_X1 U10522 ( .A1(n8996), .A2(n10508), .A3(n10120), .ZN(n10507) );
  NOR2_X1 U10523 ( .A1(n10236), .A2(n10235), .ZN(n10508) );
  INV_X1 U10524 ( .A(n10509), .ZN(n10506) );
  NAND2_X1 U10525 ( .A1(n10235), .A2(n10236), .ZN(n10509) );
  NAND2_X1 U10526 ( .A1(n10377), .A2(n10510), .ZN(n10236) );
  NAND2_X1 U10527 ( .A1(n10376), .A2(n10378), .ZN(n10510) );
  NAND2_X1 U10528 ( .A1(n10511), .A2(n10512), .ZN(n10378) );
  NAND2_X1 U10529 ( .A1(b_24_), .A2(a_14_), .ZN(n10512) );
  INV_X1 U10530 ( .A(n10513), .ZN(n10511) );
  XOR2_X1 U10531 ( .A(n10514), .B(n10515), .Z(n10376) );
  XOR2_X1 U10532 ( .A(n10516), .B(n10517), .Z(n10514) );
  NOR2_X1 U10533 ( .A1(n8850), .A2(n10358), .ZN(n10517) );
  NAND2_X1 U10534 ( .A1(a_14_), .A2(n10513), .ZN(n10377) );
  NAND2_X1 U10535 ( .A1(n10518), .A2(n10519), .ZN(n10513) );
  NAND3_X1 U10536 ( .A1(a_15_), .A2(n10520), .A3(b_24_), .ZN(n10519) );
  NAND2_X1 U10537 ( .A1(n10247), .A2(n10249), .ZN(n10520) );
  INV_X1 U10538 ( .A(n10521), .ZN(n10518) );
  NOR2_X1 U10539 ( .A1(n10249), .A2(n10247), .ZN(n10521) );
  XNOR2_X1 U10540 ( .A(n10522), .B(n10523), .ZN(n10247) );
  XNOR2_X1 U10541 ( .A(n10524), .B(n10525), .ZN(n10523) );
  NAND2_X1 U10542 ( .A1(n10526), .A2(n10527), .ZN(n10249) );
  NAND2_X1 U10543 ( .A1(n10255), .A2(n10528), .ZN(n10527) );
  NAND2_X1 U10544 ( .A1(n10258), .A2(n10257), .ZN(n10528) );
  XNOR2_X1 U10545 ( .A(n10529), .B(n10530), .ZN(n10255) );
  XNOR2_X1 U10546 ( .A(n10531), .B(n10532), .ZN(n10530) );
  NAND2_X1 U10547 ( .A1(b_23_), .A2(a_17_), .ZN(n10532) );
  INV_X1 U10548 ( .A(n10533), .ZN(n10526) );
  NOR2_X1 U10549 ( .A1(n10257), .A2(n10258), .ZN(n10533) );
  NOR2_X1 U10550 ( .A1(n10120), .A2(n8376), .ZN(n10258) );
  NAND2_X1 U10551 ( .A1(n10264), .A2(n10534), .ZN(n10257) );
  NAND2_X1 U10552 ( .A1(n10263), .A2(n10265), .ZN(n10534) );
  NAND2_X1 U10553 ( .A1(n10535), .A2(n10536), .ZN(n10265) );
  NAND2_X1 U10554 ( .A1(b_24_), .A2(a_17_), .ZN(n10535) );
  XNOR2_X1 U10555 ( .A(n10537), .B(n10538), .ZN(n10263) );
  XOR2_X1 U10556 ( .A(n10539), .B(n10540), .Z(n10537) );
  INV_X1 U10557 ( .A(n10541), .ZN(n10264) );
  NOR2_X1 U10558 ( .A1(n10536), .A2(n8371), .ZN(n10541) );
  NAND2_X1 U10559 ( .A1(n10542), .A2(n10543), .ZN(n10536) );
  NAND2_X1 U10560 ( .A1(n10271), .A2(n10544), .ZN(n10543) );
  NAND2_X1 U10561 ( .A1(n10274), .A2(n10273), .ZN(n10544) );
  XOR2_X1 U10562 ( .A(n10545), .B(n10546), .Z(n10271) );
  XNOR2_X1 U10563 ( .A(n10547), .B(n10548), .ZN(n10546) );
  INV_X1 U10564 ( .A(n10549), .ZN(n10542) );
  NOR2_X1 U10565 ( .A1(n10273), .A2(n10274), .ZN(n10549) );
  NOR2_X1 U10566 ( .A1(n10120), .A2(n9291), .ZN(n10274) );
  NAND2_X1 U10567 ( .A1(n10550), .A2(n10551), .ZN(n10273) );
  NAND3_X1 U10568 ( .A1(a_19_), .A2(n10552), .A3(b_24_), .ZN(n10551) );
  INV_X1 U10569 ( .A(n10553), .ZN(n10552) );
  NOR2_X1 U10570 ( .A1(n10280), .A2(n10279), .ZN(n10553) );
  NAND2_X1 U10571 ( .A1(n10279), .A2(n10280), .ZN(n10550) );
  NAND2_X1 U10572 ( .A1(n10373), .A2(n10554), .ZN(n10280) );
  NAND2_X1 U10573 ( .A1(n10372), .A2(n10374), .ZN(n10554) );
  NAND2_X1 U10574 ( .A1(n10555), .A2(n10556), .ZN(n10374) );
  NAND2_X1 U10575 ( .A1(b_24_), .A2(a_20_), .ZN(n10556) );
  XNOR2_X1 U10576 ( .A(n10557), .B(n10558), .ZN(n10372) );
  XOR2_X1 U10577 ( .A(n10559), .B(n10560), .Z(n10558) );
  NAND2_X1 U10578 ( .A1(b_23_), .A2(a_21_), .ZN(n10560) );
  INV_X1 U10579 ( .A(n10561), .ZN(n10373) );
  NOR2_X1 U10580 ( .A1(n9047), .A2(n10555), .ZN(n10561) );
  NOR2_X1 U10581 ( .A1(n10562), .A2(n10563), .ZN(n10555) );
  NOR3_X1 U10582 ( .A1(n8759), .A2(n10564), .A3(n10120), .ZN(n10563) );
  NOR2_X1 U10583 ( .A1(n10293), .A2(n10292), .ZN(n10564) );
  INV_X1 U10584 ( .A(n10565), .ZN(n10562) );
  NAND2_X1 U10585 ( .A1(n10292), .A2(n10293), .ZN(n10565) );
  NAND2_X1 U10586 ( .A1(n10369), .A2(n10566), .ZN(n10293) );
  NAND2_X1 U10587 ( .A1(n10368), .A2(n10370), .ZN(n10566) );
  NAND2_X1 U10588 ( .A1(n10567), .A2(n10568), .ZN(n10370) );
  NAND2_X1 U10589 ( .A1(b_24_), .A2(a_22_), .ZN(n10568) );
  INV_X1 U10590 ( .A(n10569), .ZN(n10567) );
  XNOR2_X1 U10591 ( .A(n10570), .B(n10571), .ZN(n10368) );
  XOR2_X1 U10592 ( .A(n10572), .B(n10573), .Z(n10570) );
  NAND2_X1 U10593 ( .A1(a_22_), .A2(n10569), .ZN(n10369) );
  NAND2_X1 U10594 ( .A1(n10305), .A2(n10574), .ZN(n10569) );
  NAND2_X1 U10595 ( .A1(n10304), .A2(n10306), .ZN(n10574) );
  NAND2_X1 U10596 ( .A1(n10575), .A2(n10576), .ZN(n10306) );
  INV_X1 U10597 ( .A(n10577), .ZN(n10576) );
  NAND2_X1 U10598 ( .A1(b_24_), .A2(a_23_), .ZN(n10575) );
  XOR2_X1 U10599 ( .A(n10578), .B(n10579), .Z(n10304) );
  XOR2_X1 U10600 ( .A(n10580), .B(n10581), .Z(n10578) );
  NAND2_X1 U10601 ( .A1(n10577), .A2(a_23_), .ZN(n10305) );
  NOR2_X1 U10602 ( .A1(n10582), .A2(n10583), .ZN(n10577) );
  INV_X1 U10603 ( .A(n10584), .ZN(n10583) );
  NAND2_X1 U10604 ( .A1(n10585), .A2(n10313), .ZN(n10584) );
  NAND2_X1 U10605 ( .A1(n10311), .A2(n10312), .ZN(n10585) );
  NOR2_X1 U10606 ( .A1(n10312), .A2(n10311), .ZN(n10582) );
  XNOR2_X1 U10607 ( .A(n10586), .B(n10587), .ZN(n10311) );
  XNOR2_X1 U10608 ( .A(n10588), .B(n10589), .ZN(n10587) );
  NAND2_X1 U10609 ( .A1(n10590), .A2(n10591), .ZN(n10312) );
  NAND2_X1 U10610 ( .A1(n10322), .A2(n10592), .ZN(n10591) );
  NAND2_X1 U10611 ( .A1(n10319), .A2(n10321), .ZN(n10592) );
  NOR2_X1 U10612 ( .A1(n10120), .A2(n8788), .ZN(n10322) );
  INV_X1 U10613 ( .A(n10593), .ZN(n10590) );
  NOR2_X1 U10614 ( .A1(n10321), .A2(n10319), .ZN(n10593) );
  XNOR2_X1 U10615 ( .A(n10594), .B(n10595), .ZN(n10319) );
  XNOR2_X1 U10616 ( .A(n10596), .B(n10597), .ZN(n10595) );
  NAND2_X1 U10617 ( .A1(n10598), .A2(n10599), .ZN(n10321) );
  NAND2_X1 U10618 ( .A1(n10327), .A2(n10600), .ZN(n10599) );
  NAND2_X1 U10619 ( .A1(n10330), .A2(n10329), .ZN(n10600) );
  XNOR2_X1 U10620 ( .A(n10601), .B(n10602), .ZN(n10327) );
  XOR2_X1 U10621 ( .A(n10603), .B(n10604), .Z(n10601) );
  INV_X1 U10622 ( .A(n10605), .ZN(n10598) );
  NOR2_X1 U10623 ( .A1(n10329), .A2(n10330), .ZN(n10605) );
  NOR2_X1 U10624 ( .A1(n10120), .A2(n9344), .ZN(n10330) );
  NAND2_X1 U10625 ( .A1(n10606), .A2(n10607), .ZN(n10329) );
  NAND2_X1 U10626 ( .A1(n10339), .A2(n10608), .ZN(n10607) );
  INV_X1 U10627 ( .A(n10609), .ZN(n10608) );
  NOR2_X1 U10628 ( .A1(n10338), .A2(n10337), .ZN(n10609) );
  NOR2_X1 U10629 ( .A1(n10120), .A2(n8797), .ZN(n10339) );
  NAND2_X1 U10630 ( .A1(n10337), .A2(n10338), .ZN(n10606) );
  NAND2_X1 U10631 ( .A1(n10610), .A2(n10611), .ZN(n10338) );
  NAND2_X1 U10632 ( .A1(n10365), .A2(n10612), .ZN(n10611) );
  INV_X1 U10633 ( .A(n10613), .ZN(n10612) );
  NOR2_X1 U10634 ( .A1(n10366), .A2(n10364), .ZN(n10613) );
  NOR2_X1 U10635 ( .A1(n10120), .A2(n8314), .ZN(n10365) );
  NAND2_X1 U10636 ( .A1(n10364), .A2(n10366), .ZN(n10610) );
  NAND2_X1 U10637 ( .A1(n10614), .A2(n10615), .ZN(n10366) );
  NAND2_X1 U10638 ( .A1(n10360), .A2(n10616), .ZN(n10615) );
  INV_X1 U10639 ( .A(n10617), .ZN(n10616) );
  NOR2_X1 U10640 ( .A1(n10361), .A2(n10362), .ZN(n10617) );
  NOR2_X1 U10641 ( .A1(n10120), .A2(n9098), .ZN(n10360) );
  NAND2_X1 U10642 ( .A1(n10362), .A2(n10361), .ZN(n10614) );
  NAND2_X1 U10643 ( .A1(n10618), .A2(n10619), .ZN(n10361) );
  NAND2_X1 U10644 ( .A1(b_22_), .A2(n10620), .ZN(n10619) );
  NAND2_X1 U10645 ( .A1(n8299), .A2(n10621), .ZN(n10620) );
  NAND2_X1 U10646 ( .A1(a_31_), .A2(n10358), .ZN(n10621) );
  NAND2_X1 U10647 ( .A1(b_23_), .A2(n10622), .ZN(n10618) );
  NAND2_X1 U10648 ( .A1(n8303), .A2(n10623), .ZN(n10622) );
  NAND2_X1 U10649 ( .A1(a_30_), .A2(n10624), .ZN(n10623) );
  NOR3_X1 U10650 ( .A1(n10358), .A2(n9631), .A3(n10120), .ZN(n10362) );
  XOR2_X1 U10651 ( .A(n10625), .B(n10626), .Z(n10364) );
  XOR2_X1 U10652 ( .A(n10627), .B(n10628), .Z(n10625) );
  XOR2_X1 U10653 ( .A(n10629), .B(n10630), .Z(n10337) );
  XOR2_X1 U10654 ( .A(n10631), .B(n10632), .Z(n10629) );
  XNOR2_X1 U10655 ( .A(n10633), .B(n10634), .ZN(n10292) );
  NAND2_X1 U10656 ( .A1(n10635), .A2(n10636), .ZN(n10633) );
  XOR2_X1 U10657 ( .A(n10637), .B(n10638), .Z(n10279) );
  XNOR2_X1 U10658 ( .A(n10639), .B(n10640), .ZN(n10638) );
  XNOR2_X1 U10659 ( .A(n10641), .B(n10642), .ZN(n10235) );
  NAND2_X1 U10660 ( .A1(n10643), .A2(n10644), .ZN(n10641) );
  XOR2_X1 U10661 ( .A(n10645), .B(n10646), .Z(n10379) );
  XOR2_X1 U10662 ( .A(n10647), .B(n10648), .Z(n10646) );
  NAND2_X1 U10663 ( .A1(b_23_), .A2(a_13_), .ZN(n10648) );
  XNOR2_X1 U10664 ( .A(n10649), .B(n10650), .ZN(n10392) );
  XNOR2_X1 U10665 ( .A(n10651), .B(n10652), .ZN(n10649) );
  XOR2_X1 U10666 ( .A(n10653), .B(n10654), .Z(n10395) );
  XNOR2_X1 U10667 ( .A(n10655), .B(n10656), .ZN(n10653) );
  XOR2_X1 U10668 ( .A(n10657), .B(n10658), .Z(n10400) );
  XNOR2_X1 U10669 ( .A(n10659), .B(n10660), .ZN(n10658) );
  NAND2_X1 U10670 ( .A1(b_23_), .A2(a_7_), .ZN(n10660) );
  XOR2_X1 U10671 ( .A(n10661), .B(n10662), .Z(n10404) );
  NAND2_X1 U10672 ( .A1(n10663), .A2(n10664), .ZN(n10661) );
  XNOR2_X1 U10673 ( .A(n10665), .B(n10666), .ZN(n10408) );
  XOR2_X1 U10674 ( .A(n10667), .B(n10668), .Z(n10666) );
  NAND2_X1 U10675 ( .A1(b_23_), .A2(a_5_), .ZN(n10668) );
  NAND2_X1 U10676 ( .A1(n10414), .A2(n10412), .ZN(n10453) );
  XNOR2_X1 U10677 ( .A(n10669), .B(n10670), .ZN(n10412) );
  XOR2_X1 U10678 ( .A(n10671), .B(n10672), .Z(n10670) );
  NAND2_X1 U10679 ( .A1(b_23_), .A2(a_4_), .ZN(n10672) );
  NOR2_X1 U10680 ( .A1(n10120), .A2(n8900), .ZN(n10414) );
  XOR2_X1 U10681 ( .A(n10673), .B(n10674), .Z(n10416) );
  XOR2_X1 U10682 ( .A(n10675), .B(n10676), .Z(n10673) );
  NOR2_X1 U10683 ( .A1(n8900), .A2(n10358), .ZN(n10676) );
  INV_X1 U10684 ( .A(n10677), .ZN(n10446) );
  NOR2_X1 U10685 ( .A1(n10422), .A2(n10419), .ZN(n10677) );
  XNOR2_X1 U10686 ( .A(n10678), .B(n10679), .ZN(n10419) );
  XOR2_X1 U10687 ( .A(n10680), .B(n10681), .Z(n10678) );
  NOR2_X1 U10688 ( .A1(n8448), .A2(n10358), .ZN(n10681) );
  NAND2_X1 U10689 ( .A1(b_24_), .A2(a_1_), .ZN(n10422) );
  XOR2_X1 U10690 ( .A(n10682), .B(n10683), .Z(n10423) );
  XNOR2_X1 U10691 ( .A(n10684), .B(n10685), .ZN(n10683) );
  NAND2_X1 U10692 ( .A1(b_23_), .A2(a_1_), .ZN(n10685) );
  XOR2_X1 U10693 ( .A(n10436), .B(n10686), .Z(n8626) );
  XNOR2_X1 U10694 ( .A(n10435), .B(n10687), .ZN(n10686) );
  NAND2_X1 U10695 ( .A1(b_23_), .A2(a_0_), .ZN(n10687) );
  NOR2_X1 U10696 ( .A1(n10688), .A2(n10689), .ZN(n10435) );
  NOR3_X1 U10697 ( .A1(n8569), .A2(n10690), .A3(n10358), .ZN(n10689) );
  INV_X1 U10698 ( .A(n10691), .ZN(n10690) );
  NAND2_X1 U10699 ( .A1(n10684), .A2(n10682), .ZN(n10691) );
  NOR2_X1 U10700 ( .A1(n10682), .A2(n10684), .ZN(n10688) );
  NOR2_X1 U10701 ( .A1(n10692), .A2(n10693), .ZN(n10684) );
  NOR3_X1 U10702 ( .A1(n8448), .A2(n10694), .A3(n10358), .ZN(n10693) );
  NOR2_X1 U10703 ( .A1(n10680), .A2(n10679), .ZN(n10694) );
  INV_X1 U10704 ( .A(n10695), .ZN(n10692) );
  NAND2_X1 U10705 ( .A1(n10679), .A2(n10680), .ZN(n10695) );
  NAND2_X1 U10706 ( .A1(n10696), .A2(n10697), .ZN(n10680) );
  NAND3_X1 U10707 ( .A1(a_3_), .A2(n10698), .A3(b_23_), .ZN(n10697) );
  INV_X1 U10708 ( .A(n10699), .ZN(n10698) );
  NOR2_X1 U10709 ( .A1(n10675), .A2(n10674), .ZN(n10699) );
  NAND2_X1 U10710 ( .A1(n10674), .A2(n10675), .ZN(n10696) );
  NAND2_X1 U10711 ( .A1(n10700), .A2(n10701), .ZN(n10675) );
  NAND3_X1 U10712 ( .A1(a_4_), .A2(n10702), .A3(b_23_), .ZN(n10701) );
  INV_X1 U10713 ( .A(n10703), .ZN(n10702) );
  NOR2_X1 U10714 ( .A1(n10671), .A2(n10669), .ZN(n10703) );
  NAND2_X1 U10715 ( .A1(n10669), .A2(n10671), .ZN(n10700) );
  NAND2_X1 U10716 ( .A1(n10704), .A2(n10705), .ZN(n10671) );
  NAND3_X1 U10717 ( .A1(a_5_), .A2(n10706), .A3(b_23_), .ZN(n10705) );
  INV_X1 U10718 ( .A(n10707), .ZN(n10706) );
  NOR2_X1 U10719 ( .A1(n10667), .A2(n10665), .ZN(n10707) );
  NAND2_X1 U10720 ( .A1(n10665), .A2(n10667), .ZN(n10704) );
  NAND2_X1 U10721 ( .A1(n10663), .A2(n10708), .ZN(n10667) );
  NAND2_X1 U10722 ( .A1(n10662), .A2(n10664), .ZN(n10708) );
  NAND2_X1 U10723 ( .A1(n10709), .A2(n10710), .ZN(n10664) );
  NAND2_X1 U10724 ( .A1(b_23_), .A2(a_6_), .ZN(n10710) );
  INV_X1 U10725 ( .A(n10711), .ZN(n10709) );
  XNOR2_X1 U10726 ( .A(n10712), .B(n10713), .ZN(n10662) );
  XOR2_X1 U10727 ( .A(n10714), .B(n10715), .Z(n10713) );
  NAND2_X1 U10728 ( .A1(b_22_), .A2(a_7_), .ZN(n10715) );
  NAND2_X1 U10729 ( .A1(a_6_), .A2(n10711), .ZN(n10663) );
  NAND2_X1 U10730 ( .A1(n10716), .A2(n10717), .ZN(n10711) );
  NAND3_X1 U10731 ( .A1(a_7_), .A2(n10718), .A3(b_23_), .ZN(n10717) );
  NAND2_X1 U10732 ( .A1(n10657), .A2(n10719), .ZN(n10718) );
  INV_X1 U10733 ( .A(n10659), .ZN(n10719) );
  NAND2_X1 U10734 ( .A1(n10659), .A2(n10720), .ZN(n10716) );
  INV_X1 U10735 ( .A(n10657), .ZN(n10720) );
  XOR2_X1 U10736 ( .A(n10721), .B(n10722), .Z(n10657) );
  XOR2_X1 U10737 ( .A(n10723), .B(n10724), .Z(n10722) );
  NAND2_X1 U10738 ( .A1(b_22_), .A2(a_8_), .ZN(n10724) );
  NOR2_X1 U10739 ( .A1(n10725), .A2(n10726), .ZN(n10659) );
  INV_X1 U10740 ( .A(n10727), .ZN(n10726) );
  NAND2_X1 U10741 ( .A1(n10474), .A2(n10728), .ZN(n10727) );
  NAND2_X1 U10742 ( .A1(n10477), .A2(n10476), .ZN(n10728) );
  XOR2_X1 U10743 ( .A(n10729), .B(n10730), .Z(n10474) );
  NAND2_X1 U10744 ( .A1(n10731), .A2(n10732), .ZN(n10729) );
  NOR2_X1 U10745 ( .A1(n10476), .A2(n10477), .ZN(n10725) );
  NOR2_X1 U10746 ( .A1(n10358), .A2(n8968), .ZN(n10477) );
  NAND2_X1 U10747 ( .A1(n10733), .A2(n10734), .ZN(n10476) );
  NAND2_X1 U10748 ( .A1(n10656), .A2(n10735), .ZN(n10734) );
  NAND2_X1 U10749 ( .A1(n10655), .A2(n10654), .ZN(n10735) );
  NOR2_X1 U10750 ( .A1(n10358), .A2(n8971), .ZN(n10656) );
  INV_X1 U10751 ( .A(n10736), .ZN(n10733) );
  NOR2_X1 U10752 ( .A1(n10654), .A2(n10655), .ZN(n10736) );
  NOR2_X1 U10753 ( .A1(n10737), .A2(n10738), .ZN(n10655) );
  INV_X1 U10754 ( .A(n10739), .ZN(n10738) );
  NAND2_X1 U10755 ( .A1(n10651), .A2(n10740), .ZN(n10739) );
  NAND2_X1 U10756 ( .A1(n10650), .A2(n10652), .ZN(n10740) );
  NAND2_X1 U10757 ( .A1(n10741), .A2(n10742), .ZN(n10651) );
  NAND3_X1 U10758 ( .A1(a_11_), .A2(n10743), .A3(b_23_), .ZN(n10742) );
  NAND2_X1 U10759 ( .A1(n10490), .A2(n10492), .ZN(n10743) );
  INV_X1 U10760 ( .A(n10744), .ZN(n10741) );
  NOR2_X1 U10761 ( .A1(n10492), .A2(n10490), .ZN(n10744) );
  XNOR2_X1 U10762 ( .A(n10745), .B(n10746), .ZN(n10490) );
  XNOR2_X1 U10763 ( .A(n10747), .B(n10748), .ZN(n10746) );
  NAND2_X1 U10764 ( .A1(b_22_), .A2(a_12_), .ZN(n10748) );
  NAND2_X1 U10765 ( .A1(n10749), .A2(n10750), .ZN(n10492) );
  NAND2_X1 U10766 ( .A1(n10497), .A2(n10751), .ZN(n10750) );
  INV_X1 U10767 ( .A(n10752), .ZN(n10751) );
  NOR2_X1 U10768 ( .A1(n10500), .A2(n10499), .ZN(n10752) );
  XOR2_X1 U10769 ( .A(n10753), .B(n10754), .Z(n10497) );
  XOR2_X1 U10770 ( .A(n10755), .B(n10756), .Z(n10754) );
  NAND2_X1 U10771 ( .A1(b_22_), .A2(a_13_), .ZN(n10756) );
  NAND2_X1 U10772 ( .A1(n10499), .A2(n10500), .ZN(n10749) );
  NAND2_X1 U10773 ( .A1(b_23_), .A2(a_12_), .ZN(n10500) );
  NOR2_X1 U10774 ( .A1(n10757), .A2(n10758), .ZN(n10499) );
  NOR3_X1 U10775 ( .A1(n8996), .A2(n10759), .A3(n10358), .ZN(n10758) );
  NOR2_X1 U10776 ( .A1(n10647), .A2(n10645), .ZN(n10759) );
  INV_X1 U10777 ( .A(n10760), .ZN(n10757) );
  NAND2_X1 U10778 ( .A1(n10645), .A2(n10647), .ZN(n10760) );
  NAND2_X1 U10779 ( .A1(n10643), .A2(n10761), .ZN(n10647) );
  NAND2_X1 U10780 ( .A1(n10642), .A2(n10644), .ZN(n10761) );
  NAND2_X1 U10781 ( .A1(n10762), .A2(n10763), .ZN(n10644) );
  NAND2_X1 U10782 ( .A1(b_23_), .A2(a_14_), .ZN(n10763) );
  XOR2_X1 U10783 ( .A(n10764), .B(n10765), .Z(n10642) );
  XOR2_X1 U10784 ( .A(n10766), .B(n10767), .Z(n10764) );
  NOR2_X1 U10785 ( .A1(n8850), .A2(n10624), .ZN(n10767) );
  NAND2_X1 U10786 ( .A1(a_14_), .A2(n10768), .ZN(n10643) );
  INV_X1 U10787 ( .A(n10762), .ZN(n10768) );
  NOR2_X1 U10788 ( .A1(n10769), .A2(n10770), .ZN(n10762) );
  NOR3_X1 U10789 ( .A1(n8850), .A2(n10771), .A3(n10358), .ZN(n10770) );
  INV_X1 U10790 ( .A(n10772), .ZN(n10771) );
  NAND2_X1 U10791 ( .A1(n10515), .A2(n10516), .ZN(n10772) );
  NOR2_X1 U10792 ( .A1(n10516), .A2(n10515), .ZN(n10769) );
  XOR2_X1 U10793 ( .A(n10773), .B(n10774), .Z(n10515) );
  NAND2_X1 U10794 ( .A1(n10775), .A2(n10776), .ZN(n10773) );
  NAND2_X1 U10795 ( .A1(n10777), .A2(n10778), .ZN(n10516) );
  NAND2_X1 U10796 ( .A1(n10522), .A2(n10779), .ZN(n10778) );
  NAND2_X1 U10797 ( .A1(n10525), .A2(n10524), .ZN(n10779) );
  XOR2_X1 U10798 ( .A(n10780), .B(n10781), .Z(n10522) );
  XNOR2_X1 U10799 ( .A(n10782), .B(n10783), .ZN(n10780) );
  NOR2_X1 U10800 ( .A1(n8371), .A2(n10624), .ZN(n10783) );
  INV_X1 U10801 ( .A(n10784), .ZN(n10777) );
  NOR2_X1 U10802 ( .A1(n10524), .A2(n10525), .ZN(n10784) );
  NOR2_X1 U10803 ( .A1(n10358), .A2(n8376), .ZN(n10525) );
  NAND2_X1 U10804 ( .A1(n10785), .A2(n10786), .ZN(n10524) );
  NAND3_X1 U10805 ( .A1(a_17_), .A2(n10787), .A3(b_23_), .ZN(n10786) );
  NAND2_X1 U10806 ( .A1(n10788), .A2(n10789), .ZN(n10787) );
  INV_X1 U10807 ( .A(n10531), .ZN(n10789) );
  INV_X1 U10808 ( .A(n10529), .ZN(n10788) );
  NAND2_X1 U10809 ( .A1(n10531), .A2(n10529), .ZN(n10785) );
  XNOR2_X1 U10810 ( .A(n10790), .B(n10791), .ZN(n10529) );
  XOR2_X1 U10811 ( .A(n10792), .B(n10793), .Z(n10790) );
  NOR2_X1 U10812 ( .A1(n10794), .A2(n10795), .ZN(n10531) );
  INV_X1 U10813 ( .A(n10796), .ZN(n10795) );
  NAND2_X1 U10814 ( .A1(n10538), .A2(n10797), .ZN(n10796) );
  NAND2_X1 U10815 ( .A1(n10540), .A2(n10539), .ZN(n10797) );
  XNOR2_X1 U10816 ( .A(n10798), .B(n10799), .ZN(n10538) );
  XOR2_X1 U10817 ( .A(n10800), .B(n10801), .Z(n10798) );
  NOR2_X1 U10818 ( .A1(n8742), .A2(n10624), .ZN(n10801) );
  NOR2_X1 U10819 ( .A1(n10539), .A2(n10540), .ZN(n10794) );
  NOR2_X1 U10820 ( .A1(n10358), .A2(n9291), .ZN(n10540) );
  NAND2_X1 U10821 ( .A1(n10802), .A2(n10803), .ZN(n10539) );
  NAND2_X1 U10822 ( .A1(n10548), .A2(n10804), .ZN(n10803) );
  NAND2_X1 U10823 ( .A1(n10545), .A2(n10547), .ZN(n10804) );
  NOR2_X1 U10824 ( .A1(n10358), .A2(n8742), .ZN(n10548) );
  INV_X1 U10825 ( .A(n10805), .ZN(n10802) );
  NOR2_X1 U10826 ( .A1(n10547), .A2(n10545), .ZN(n10805) );
  XOR2_X1 U10827 ( .A(n10806), .B(n10807), .Z(n10545) );
  NAND2_X1 U10828 ( .A1(n10808), .A2(n10809), .ZN(n10806) );
  NAND2_X1 U10829 ( .A1(n10810), .A2(n10811), .ZN(n10547) );
  NAND2_X1 U10830 ( .A1(n10637), .A2(n10812), .ZN(n10811) );
  NAND2_X1 U10831 ( .A1(n10640), .A2(n10639), .ZN(n10812) );
  XOR2_X1 U10832 ( .A(n10813), .B(n10814), .Z(n10637) );
  NAND2_X1 U10833 ( .A1(n10815), .A2(n10816), .ZN(n10813) );
  INV_X1 U10834 ( .A(n10817), .ZN(n10810) );
  NOR2_X1 U10835 ( .A1(n10639), .A2(n10640), .ZN(n10817) );
  NOR2_X1 U10836 ( .A1(n10358), .A2(n9047), .ZN(n10640) );
  NAND2_X1 U10837 ( .A1(n10818), .A2(n10819), .ZN(n10639) );
  NAND3_X1 U10838 ( .A1(a_21_), .A2(n10820), .A3(b_23_), .ZN(n10819) );
  INV_X1 U10839 ( .A(n10821), .ZN(n10820) );
  NOR2_X1 U10840 ( .A1(n10559), .A2(n10557), .ZN(n10821) );
  NAND2_X1 U10841 ( .A1(n10557), .A2(n10559), .ZN(n10818) );
  NAND2_X1 U10842 ( .A1(n10635), .A2(n10822), .ZN(n10559) );
  NAND2_X1 U10843 ( .A1(n10634), .A2(n10636), .ZN(n10822) );
  NAND2_X1 U10844 ( .A1(n10823), .A2(n10824), .ZN(n10636) );
  NAND2_X1 U10845 ( .A1(b_23_), .A2(a_22_), .ZN(n10823) );
  XNOR2_X1 U10846 ( .A(n10825), .B(n10826), .ZN(n10634) );
  NAND2_X1 U10847 ( .A1(n10827), .A2(n10828), .ZN(n10825) );
  NAND2_X1 U10848 ( .A1(n10829), .A2(a_22_), .ZN(n10635) );
  INV_X1 U10849 ( .A(n10824), .ZN(n10829) );
  NAND2_X1 U10850 ( .A1(n10830), .A2(n10831), .ZN(n10824) );
  NAND2_X1 U10851 ( .A1(n10571), .A2(n10832), .ZN(n10831) );
  NAND2_X1 U10852 ( .A1(n10573), .A2(n10572), .ZN(n10832) );
  XNOR2_X1 U10853 ( .A(n10833), .B(n10834), .ZN(n10571) );
  XOR2_X1 U10854 ( .A(n10835), .B(n10836), .Z(n10833) );
  INV_X1 U10855 ( .A(n10837), .ZN(n10830) );
  NOR2_X1 U10856 ( .A1(n10572), .A2(n10573), .ZN(n10837) );
  NAND2_X1 U10857 ( .A1(n10838), .A2(n10839), .ZN(n10572) );
  NAND2_X1 U10858 ( .A1(n10581), .A2(n10840), .ZN(n10839) );
  INV_X1 U10859 ( .A(n10841), .ZN(n10840) );
  NOR2_X1 U10860 ( .A1(n10580), .A2(n10579), .ZN(n10841) );
  NOR2_X1 U10861 ( .A1(n10358), .A2(n8779), .ZN(n10581) );
  NAND2_X1 U10862 ( .A1(n10579), .A2(n10580), .ZN(n10838) );
  NAND2_X1 U10863 ( .A1(n10842), .A2(n10843), .ZN(n10580) );
  NAND2_X1 U10864 ( .A1(n10589), .A2(n10844), .ZN(n10843) );
  NAND2_X1 U10865 ( .A1(n10586), .A2(n10588), .ZN(n10844) );
  NOR2_X1 U10866 ( .A1(n10358), .A2(n8788), .ZN(n10589) );
  INV_X1 U10867 ( .A(n10845), .ZN(n10842) );
  NOR2_X1 U10868 ( .A1(n10588), .A2(n10586), .ZN(n10845) );
  XNOR2_X1 U10869 ( .A(n10846), .B(n10847), .ZN(n10586) );
  XNOR2_X1 U10870 ( .A(n10848), .B(n10849), .ZN(n10847) );
  NAND2_X1 U10871 ( .A1(n10850), .A2(n10851), .ZN(n10588) );
  NAND2_X1 U10872 ( .A1(n10594), .A2(n10852), .ZN(n10851) );
  NAND2_X1 U10873 ( .A1(n10597), .A2(n10596), .ZN(n10852) );
  XNOR2_X1 U10874 ( .A(n10853), .B(n10854), .ZN(n10594) );
  XOR2_X1 U10875 ( .A(n10855), .B(n10856), .Z(n10853) );
  INV_X1 U10876 ( .A(n10857), .ZN(n10850) );
  NOR2_X1 U10877 ( .A1(n10596), .A2(n10597), .ZN(n10857) );
  NOR2_X1 U10878 ( .A1(n10358), .A2(n9344), .ZN(n10597) );
  NAND2_X1 U10879 ( .A1(n10858), .A2(n10859), .ZN(n10596) );
  NAND2_X1 U10880 ( .A1(n10604), .A2(n10860), .ZN(n10859) );
  INV_X1 U10881 ( .A(n10861), .ZN(n10860) );
  NOR2_X1 U10882 ( .A1(n10603), .A2(n10602), .ZN(n10861) );
  NOR2_X1 U10883 ( .A1(n10358), .A2(n8797), .ZN(n10604) );
  NAND2_X1 U10884 ( .A1(n10602), .A2(n10603), .ZN(n10858) );
  NAND2_X1 U10885 ( .A1(n10862), .A2(n10863), .ZN(n10603) );
  NAND2_X1 U10886 ( .A1(n10631), .A2(n10864), .ZN(n10863) );
  INV_X1 U10887 ( .A(n10865), .ZN(n10864) );
  NOR2_X1 U10888 ( .A1(n10632), .A2(n10630), .ZN(n10865) );
  NOR2_X1 U10889 ( .A1(n10358), .A2(n8314), .ZN(n10631) );
  NAND2_X1 U10890 ( .A1(n10630), .A2(n10632), .ZN(n10862) );
  NAND2_X1 U10891 ( .A1(n10866), .A2(n10867), .ZN(n10632) );
  NAND2_X1 U10892 ( .A1(n10626), .A2(n10868), .ZN(n10867) );
  INV_X1 U10893 ( .A(n10869), .ZN(n10868) );
  NOR2_X1 U10894 ( .A1(n10627), .A2(n10628), .ZN(n10869) );
  NOR2_X1 U10895 ( .A1(n10358), .A2(n9098), .ZN(n10626) );
  NAND2_X1 U10896 ( .A1(n10628), .A2(n10627), .ZN(n10866) );
  NAND2_X1 U10897 ( .A1(n10870), .A2(n10871), .ZN(n10627) );
  NAND2_X1 U10898 ( .A1(b_21_), .A2(n10872), .ZN(n10871) );
  NAND2_X1 U10899 ( .A1(n8299), .A2(n10873), .ZN(n10872) );
  NAND2_X1 U10900 ( .A1(a_31_), .A2(n10624), .ZN(n10873) );
  NAND2_X1 U10901 ( .A1(b_22_), .A2(n10874), .ZN(n10870) );
  NAND2_X1 U10902 ( .A1(n8303), .A2(n10875), .ZN(n10874) );
  NAND2_X1 U10903 ( .A1(a_30_), .A2(n10876), .ZN(n10875) );
  NOR3_X1 U10904 ( .A1(n10358), .A2(n9631), .A3(n10624), .ZN(n10628) );
  XOR2_X1 U10905 ( .A(n10877), .B(n10878), .Z(n10630) );
  XOR2_X1 U10906 ( .A(n10879), .B(n10880), .Z(n10877) );
  XOR2_X1 U10907 ( .A(n10881), .B(n10882), .Z(n10602) );
  XOR2_X1 U10908 ( .A(n10883), .B(n10884), .Z(n10881) );
  XNOR2_X1 U10909 ( .A(n10885), .B(n10886), .ZN(n10579) );
  XNOR2_X1 U10910 ( .A(n10887), .B(n10888), .ZN(n10886) );
  XOR2_X1 U10911 ( .A(n10889), .B(n10890), .Z(n10557) );
  XOR2_X1 U10912 ( .A(n10891), .B(n10892), .Z(n10889) );
  XNOR2_X1 U10913 ( .A(n10893), .B(n10894), .ZN(n10645) );
  NAND2_X1 U10914 ( .A1(n10895), .A2(n10896), .ZN(n10893) );
  NOR2_X1 U10915 ( .A1(n10652), .A2(n10650), .ZN(n10737) );
  XOR2_X1 U10916 ( .A(n10897), .B(n10898), .Z(n10650) );
  XOR2_X1 U10917 ( .A(n10899), .B(n10900), .Z(n10898) );
  NAND2_X1 U10918 ( .A1(b_22_), .A2(a_11_), .ZN(n10900) );
  NAND2_X1 U10919 ( .A1(b_23_), .A2(a_10_), .ZN(n10652) );
  XOR2_X1 U10920 ( .A(n10901), .B(n10902), .Z(n10654) );
  XOR2_X1 U10921 ( .A(n10903), .B(n10904), .Z(n10901) );
  XNOR2_X1 U10922 ( .A(n10905), .B(n10906), .ZN(n10665) );
  NAND2_X1 U10923 ( .A1(n10907), .A2(n10908), .ZN(n10905) );
  XNOR2_X1 U10924 ( .A(n10909), .B(n10910), .ZN(n10669) );
  XOR2_X1 U10925 ( .A(n10911), .B(n10912), .Z(n10910) );
  NAND2_X1 U10926 ( .A1(b_22_), .A2(a_5_), .ZN(n10912) );
  XNOR2_X1 U10927 ( .A(n10913), .B(n10914), .ZN(n10674) );
  NAND2_X1 U10928 ( .A1(n10915), .A2(n10916), .ZN(n10913) );
  XNOR2_X1 U10929 ( .A(n10917), .B(n10918), .ZN(n10679) );
  XOR2_X1 U10930 ( .A(n10919), .B(n10920), .Z(n10917) );
  XNOR2_X1 U10931 ( .A(n10921), .B(n10922), .ZN(n10682) );
  XOR2_X1 U10932 ( .A(n10923), .B(n10924), .Z(n10921) );
  XOR2_X1 U10933 ( .A(n10925), .B(n10926), .Z(n10436) );
  XNOR2_X1 U10934 ( .A(n10927), .B(n10928), .ZN(n10925) );
  NAND2_X1 U10935 ( .A1(n10929), .A2(n10930), .ZN(n8501) );
  NAND2_X1 U10936 ( .A1(n8621), .A2(n8622), .ZN(n10930) );
  XNOR2_X1 U10937 ( .A(n8614), .B(n8613), .ZN(n10929) );
  NAND3_X1 U10938 ( .A1(n8621), .A2(n8622), .A3(n10931), .ZN(n8500) );
  XNOR2_X1 U10939 ( .A(n8614), .B(n10932), .ZN(n10931) );
  INV_X1 U10940 ( .A(n8613), .ZN(n10932) );
  NAND2_X1 U10941 ( .A1(n10439), .A2(n10933), .ZN(n8622) );
  NAND2_X1 U10942 ( .A1(n10438), .A2(n10440), .ZN(n10933) );
  NAND2_X1 U10943 ( .A1(n10934), .A2(n10935), .ZN(n10440) );
  NAND2_X1 U10944 ( .A1(b_22_), .A2(a_0_), .ZN(n10935) );
  XNOR2_X1 U10945 ( .A(n10936), .B(n10937), .ZN(n10438) );
  XOR2_X1 U10946 ( .A(n10938), .B(n10939), .Z(n10937) );
  NAND2_X1 U10947 ( .A1(b_21_), .A2(a_1_), .ZN(n10939) );
  NAND2_X1 U10948 ( .A1(a_0_), .A2(n10940), .ZN(n10439) );
  INV_X1 U10949 ( .A(n10934), .ZN(n10940) );
  NOR2_X1 U10950 ( .A1(n10941), .A2(n10942), .ZN(n10934) );
  INV_X1 U10951 ( .A(n10943), .ZN(n10942) );
  NAND2_X1 U10952 ( .A1(n10928), .A2(n10944), .ZN(n10943) );
  NAND2_X1 U10953 ( .A1(n10927), .A2(n10926), .ZN(n10944) );
  NOR2_X1 U10954 ( .A1(n10624), .A2(n8569), .ZN(n10928) );
  NOR2_X1 U10955 ( .A1(n10926), .A2(n10927), .ZN(n10941) );
  NOR2_X1 U10956 ( .A1(n10945), .A2(n10946), .ZN(n10927) );
  INV_X1 U10957 ( .A(n10947), .ZN(n10946) );
  NAND2_X1 U10958 ( .A1(n10924), .A2(n10948), .ZN(n10947) );
  NAND2_X1 U10959 ( .A1(n10922), .A2(n10923), .ZN(n10948) );
  NOR2_X1 U10960 ( .A1(n10624), .A2(n8448), .ZN(n10924) );
  NOR2_X1 U10961 ( .A1(n10922), .A2(n10923), .ZN(n10945) );
  NAND2_X1 U10962 ( .A1(n10949), .A2(n10950), .ZN(n10923) );
  NAND2_X1 U10963 ( .A1(n10918), .A2(n10951), .ZN(n10950) );
  NAND2_X1 U10964 ( .A1(n10920), .A2(n10919), .ZN(n10951) );
  XNOR2_X1 U10965 ( .A(n10952), .B(n10953), .ZN(n10918) );
  XOR2_X1 U10966 ( .A(n10954), .B(n10955), .Z(n10952) );
  NOR2_X1 U10967 ( .A1(n8439), .A2(n10876), .ZN(n10955) );
  INV_X1 U10968 ( .A(n10956), .ZN(n10949) );
  NOR2_X1 U10969 ( .A1(n10919), .A2(n10920), .ZN(n10956) );
  NOR2_X1 U10970 ( .A1(n10624), .A2(n8900), .ZN(n10920) );
  NAND2_X1 U10971 ( .A1(n10915), .A2(n10957), .ZN(n10919) );
  NAND2_X1 U10972 ( .A1(n10914), .A2(n10916), .ZN(n10957) );
  NAND2_X1 U10973 ( .A1(n10958), .A2(n10959), .ZN(n10916) );
  NAND2_X1 U10974 ( .A1(b_22_), .A2(a_4_), .ZN(n10959) );
  INV_X1 U10975 ( .A(n10960), .ZN(n10958) );
  XNOR2_X1 U10976 ( .A(n10961), .B(n10962), .ZN(n10914) );
  XOR2_X1 U10977 ( .A(n10963), .B(n10964), .Z(n10962) );
  NAND2_X1 U10978 ( .A1(b_21_), .A2(a_5_), .ZN(n10964) );
  NAND2_X1 U10979 ( .A1(a_4_), .A2(n10960), .ZN(n10915) );
  NAND2_X1 U10980 ( .A1(n10965), .A2(n10966), .ZN(n10960) );
  INV_X1 U10981 ( .A(n10967), .ZN(n10966) );
  NOR3_X1 U10982 ( .A1(n8938), .A2(n10968), .A3(n10624), .ZN(n10967) );
  NOR2_X1 U10983 ( .A1(n10909), .A2(n10911), .ZN(n10968) );
  NAND2_X1 U10984 ( .A1(n10909), .A2(n10911), .ZN(n10965) );
  NAND2_X1 U10985 ( .A1(n10907), .A2(n10969), .ZN(n10911) );
  NAND2_X1 U10986 ( .A1(n10906), .A2(n10908), .ZN(n10969) );
  NAND2_X1 U10987 ( .A1(n10970), .A2(n10971), .ZN(n10908) );
  NAND2_X1 U10988 ( .A1(b_22_), .A2(a_6_), .ZN(n10971) );
  XOR2_X1 U10989 ( .A(n10972), .B(n10973), .Z(n10906) );
  XOR2_X1 U10990 ( .A(n10974), .B(n10975), .Z(n10972) );
  NOR2_X1 U10991 ( .A1(n8425), .A2(n10876), .ZN(n10975) );
  INV_X1 U10992 ( .A(n10976), .ZN(n10907) );
  NOR2_X1 U10993 ( .A1(n8430), .A2(n10970), .ZN(n10976) );
  NOR2_X1 U10994 ( .A1(n10977), .A2(n10978), .ZN(n10970) );
  NOR3_X1 U10995 ( .A1(n8425), .A2(n10979), .A3(n10624), .ZN(n10978) );
  NOR2_X1 U10996 ( .A1(n10712), .A2(n10714), .ZN(n10979) );
  INV_X1 U10997 ( .A(n10980), .ZN(n10977) );
  NAND2_X1 U10998 ( .A1(n10712), .A2(n10714), .ZN(n10980) );
  NAND2_X1 U10999 ( .A1(n10981), .A2(n10982), .ZN(n10714) );
  NAND3_X1 U11000 ( .A1(a_8_), .A2(n10983), .A3(b_22_), .ZN(n10982) );
  INV_X1 U11001 ( .A(n10984), .ZN(n10983) );
  NOR2_X1 U11002 ( .A1(n10721), .A2(n10723), .ZN(n10984) );
  NAND2_X1 U11003 ( .A1(n10721), .A2(n10723), .ZN(n10981) );
  NAND2_X1 U11004 ( .A1(n10731), .A2(n10985), .ZN(n10723) );
  NAND2_X1 U11005 ( .A1(n10730), .A2(n10732), .ZN(n10985) );
  NAND2_X1 U11006 ( .A1(n10986), .A2(n10987), .ZN(n10732) );
  NAND2_X1 U11007 ( .A1(b_22_), .A2(a_9_), .ZN(n10986) );
  XNOR2_X1 U11008 ( .A(n10988), .B(n10989), .ZN(n10730) );
  XNOR2_X1 U11009 ( .A(n10990), .B(n10991), .ZN(n10988) );
  INV_X1 U11010 ( .A(n10992), .ZN(n10731) );
  NOR2_X1 U11011 ( .A1(n10987), .A2(n8971), .ZN(n10992) );
  NAND2_X1 U11012 ( .A1(n10993), .A2(n10994), .ZN(n10987) );
  NAND2_X1 U11013 ( .A1(n10902), .A2(n10995), .ZN(n10994) );
  NAND2_X1 U11014 ( .A1(n10904), .A2(n10903), .ZN(n10995) );
  XOR2_X1 U11015 ( .A(n10996), .B(n10997), .Z(n10902) );
  XNOR2_X1 U11016 ( .A(n10998), .B(n10999), .ZN(n10997) );
  INV_X1 U11017 ( .A(n11000), .ZN(n10993) );
  NOR2_X1 U11018 ( .A1(n10903), .A2(n10904), .ZN(n11000) );
  NOR2_X1 U11019 ( .A1(n10624), .A2(n8402), .ZN(n10904) );
  NAND2_X1 U11020 ( .A1(n11001), .A2(n11002), .ZN(n10903) );
  NAND3_X1 U11021 ( .A1(a_11_), .A2(n11003), .A3(b_22_), .ZN(n11002) );
  INV_X1 U11022 ( .A(n11004), .ZN(n11003) );
  NOR2_X1 U11023 ( .A1(n10897), .A2(n10899), .ZN(n11004) );
  NAND2_X1 U11024 ( .A1(n10897), .A2(n10899), .ZN(n11001) );
  NAND2_X1 U11025 ( .A1(n11005), .A2(n11006), .ZN(n10899) );
  NAND3_X1 U11026 ( .A1(a_12_), .A2(n11007), .A3(b_22_), .ZN(n11006) );
  NAND2_X1 U11027 ( .A1(n10747), .A2(n10745), .ZN(n11007) );
  INV_X1 U11028 ( .A(n11008), .ZN(n11005) );
  NOR2_X1 U11029 ( .A1(n10745), .A2(n10747), .ZN(n11008) );
  NOR2_X1 U11030 ( .A1(n11009), .A2(n11010), .ZN(n10747) );
  NOR3_X1 U11031 ( .A1(n8996), .A2(n11011), .A3(n10624), .ZN(n11010) );
  NOR2_X1 U11032 ( .A1(n10755), .A2(n10753), .ZN(n11011) );
  INV_X1 U11033 ( .A(n11012), .ZN(n11009) );
  NAND2_X1 U11034 ( .A1(n10753), .A2(n10755), .ZN(n11012) );
  NAND2_X1 U11035 ( .A1(n10895), .A2(n11013), .ZN(n10755) );
  NAND2_X1 U11036 ( .A1(n10894), .A2(n10896), .ZN(n11013) );
  NAND2_X1 U11037 ( .A1(n11014), .A2(n11015), .ZN(n10896) );
  NAND2_X1 U11038 ( .A1(b_22_), .A2(a_14_), .ZN(n11015) );
  INV_X1 U11039 ( .A(n11016), .ZN(n11014) );
  XOR2_X1 U11040 ( .A(n11017), .B(n11018), .Z(n10894) );
  XOR2_X1 U11041 ( .A(n11019), .B(n11020), .Z(n11017) );
  NOR2_X1 U11042 ( .A1(n8850), .A2(n10876), .ZN(n11020) );
  NAND2_X1 U11043 ( .A1(a_14_), .A2(n11016), .ZN(n10895) );
  NAND2_X1 U11044 ( .A1(n11021), .A2(n11022), .ZN(n11016) );
  INV_X1 U11045 ( .A(n11023), .ZN(n11022) );
  NOR3_X1 U11046 ( .A1(n8850), .A2(n11024), .A3(n10624), .ZN(n11023) );
  NOR2_X1 U11047 ( .A1(n10766), .A2(n10765), .ZN(n11024) );
  NAND2_X1 U11048 ( .A1(n10765), .A2(n10766), .ZN(n11021) );
  NAND2_X1 U11049 ( .A1(n10775), .A2(n11025), .ZN(n10766) );
  NAND2_X1 U11050 ( .A1(n10774), .A2(n10776), .ZN(n11025) );
  NAND2_X1 U11051 ( .A1(n11026), .A2(n11027), .ZN(n10776) );
  NAND2_X1 U11052 ( .A1(b_22_), .A2(a_16_), .ZN(n11027) );
  INV_X1 U11053 ( .A(n11028), .ZN(n11026) );
  XNOR2_X1 U11054 ( .A(n11029), .B(n11030), .ZN(n10774) );
  XOR2_X1 U11055 ( .A(n11031), .B(n11032), .Z(n11030) );
  NAND2_X1 U11056 ( .A1(b_21_), .A2(a_17_), .ZN(n11032) );
  NAND2_X1 U11057 ( .A1(a_16_), .A2(n11028), .ZN(n10775) );
  NAND2_X1 U11058 ( .A1(n11033), .A2(n11034), .ZN(n11028) );
  INV_X1 U11059 ( .A(n11035), .ZN(n11034) );
  NOR3_X1 U11060 ( .A1(n8371), .A2(n11036), .A3(n10624), .ZN(n11035) );
  NOR2_X1 U11061 ( .A1(n10781), .A2(n10782), .ZN(n11036) );
  NAND2_X1 U11062 ( .A1(n10782), .A2(n10781), .ZN(n11033) );
  XOR2_X1 U11063 ( .A(n11037), .B(n11038), .Z(n10781) );
  XNOR2_X1 U11064 ( .A(n11039), .B(n11040), .ZN(n11038) );
  NOR2_X1 U11065 ( .A1(n11041), .A2(n11042), .ZN(n10782) );
  INV_X1 U11066 ( .A(n11043), .ZN(n11042) );
  NAND2_X1 U11067 ( .A1(n10791), .A2(n11044), .ZN(n11043) );
  NAND2_X1 U11068 ( .A1(n10793), .A2(n10792), .ZN(n11044) );
  XOR2_X1 U11069 ( .A(n11045), .B(n11046), .Z(n10791) );
  XOR2_X1 U11070 ( .A(n11047), .B(n11048), .Z(n11046) );
  NAND2_X1 U11071 ( .A1(b_21_), .A2(a_19_), .ZN(n11048) );
  NOR2_X1 U11072 ( .A1(n10792), .A2(n10793), .ZN(n11041) );
  NOR2_X1 U11073 ( .A1(n10624), .A2(n9291), .ZN(n10793) );
  NAND2_X1 U11074 ( .A1(n11049), .A2(n11050), .ZN(n10792) );
  NAND3_X1 U11075 ( .A1(a_19_), .A2(n11051), .A3(b_22_), .ZN(n11050) );
  INV_X1 U11076 ( .A(n11052), .ZN(n11051) );
  NOR2_X1 U11077 ( .A1(n10800), .A2(n10799), .ZN(n11052) );
  NAND2_X1 U11078 ( .A1(n10799), .A2(n10800), .ZN(n11049) );
  NAND2_X1 U11079 ( .A1(n10808), .A2(n11053), .ZN(n10800) );
  NAND2_X1 U11080 ( .A1(n10807), .A2(n10809), .ZN(n11053) );
  NAND2_X1 U11081 ( .A1(n11054), .A2(n11055), .ZN(n10809) );
  NAND2_X1 U11082 ( .A1(b_22_), .A2(a_20_), .ZN(n11055) );
  INV_X1 U11083 ( .A(n11056), .ZN(n11054) );
  XNOR2_X1 U11084 ( .A(n11057), .B(n11058), .ZN(n10807) );
  XNOR2_X1 U11085 ( .A(n11059), .B(n11060), .ZN(n11058) );
  NAND2_X1 U11086 ( .A1(a_20_), .A2(n11056), .ZN(n10808) );
  NAND2_X1 U11087 ( .A1(n10815), .A2(n11061), .ZN(n11056) );
  NAND2_X1 U11088 ( .A1(n10814), .A2(n10816), .ZN(n11061) );
  NAND2_X1 U11089 ( .A1(n11062), .A2(n11063), .ZN(n10816) );
  NAND2_X1 U11090 ( .A1(b_22_), .A2(a_21_), .ZN(n11063) );
  INV_X1 U11091 ( .A(n11064), .ZN(n11062) );
  XNOR2_X1 U11092 ( .A(n11065), .B(n11066), .ZN(n10814) );
  NAND2_X1 U11093 ( .A1(n11067), .A2(n11068), .ZN(n11065) );
  NAND2_X1 U11094 ( .A1(a_21_), .A2(n11064), .ZN(n10815) );
  NAND2_X1 U11095 ( .A1(n11069), .A2(n11070), .ZN(n11064) );
  NAND2_X1 U11096 ( .A1(n10892), .A2(n11071), .ZN(n11070) );
  INV_X1 U11097 ( .A(n11072), .ZN(n11071) );
  NOR2_X1 U11098 ( .A1(n10891), .A2(n10890), .ZN(n11072) );
  NAND2_X1 U11099 ( .A1(n10890), .A2(n10891), .ZN(n11069) );
  NAND2_X1 U11100 ( .A1(n10827), .A2(n11073), .ZN(n10891) );
  NAND2_X1 U11101 ( .A1(n10826), .A2(n10828), .ZN(n11073) );
  NAND2_X1 U11102 ( .A1(n11074), .A2(n11075), .ZN(n10828) );
  NAND2_X1 U11103 ( .A1(b_22_), .A2(a_23_), .ZN(n11075) );
  INV_X1 U11104 ( .A(n11076), .ZN(n11074) );
  XOR2_X1 U11105 ( .A(n11077), .B(n11078), .Z(n10826) );
  XOR2_X1 U11106 ( .A(n11079), .B(n11080), .Z(n11077) );
  NAND2_X1 U11107 ( .A1(a_23_), .A2(n11076), .ZN(n10827) );
  NAND2_X1 U11108 ( .A1(n11081), .A2(n11082), .ZN(n11076) );
  NAND2_X1 U11109 ( .A1(n10836), .A2(n11083), .ZN(n11082) );
  INV_X1 U11110 ( .A(n11084), .ZN(n11083) );
  NOR2_X1 U11111 ( .A1(n10835), .A2(n10834), .ZN(n11084) );
  NOR2_X1 U11112 ( .A1(n10624), .A2(n8779), .ZN(n10836) );
  NAND2_X1 U11113 ( .A1(n10834), .A2(n10835), .ZN(n11081) );
  NAND2_X1 U11114 ( .A1(n11085), .A2(n11086), .ZN(n10835) );
  NAND2_X1 U11115 ( .A1(n10888), .A2(n11087), .ZN(n11086) );
  NAND2_X1 U11116 ( .A1(n10885), .A2(n10887), .ZN(n11087) );
  NOR2_X1 U11117 ( .A1(n10624), .A2(n8788), .ZN(n10888) );
  INV_X1 U11118 ( .A(n11088), .ZN(n11085) );
  NOR2_X1 U11119 ( .A1(n10887), .A2(n10885), .ZN(n11088) );
  XNOR2_X1 U11120 ( .A(n11089), .B(n11090), .ZN(n10885) );
  XNOR2_X1 U11121 ( .A(n11091), .B(n11092), .ZN(n11090) );
  NAND2_X1 U11122 ( .A1(n11093), .A2(n11094), .ZN(n10887) );
  NAND2_X1 U11123 ( .A1(n10846), .A2(n11095), .ZN(n11094) );
  NAND2_X1 U11124 ( .A1(n10849), .A2(n10848), .ZN(n11095) );
  XNOR2_X1 U11125 ( .A(n11096), .B(n11097), .ZN(n10846) );
  XOR2_X1 U11126 ( .A(n11098), .B(n11099), .Z(n11096) );
  INV_X1 U11127 ( .A(n11100), .ZN(n11093) );
  NOR2_X1 U11128 ( .A1(n10848), .A2(n10849), .ZN(n11100) );
  NOR2_X1 U11129 ( .A1(n10624), .A2(n9344), .ZN(n10849) );
  NAND2_X1 U11130 ( .A1(n11101), .A2(n11102), .ZN(n10848) );
  NAND2_X1 U11131 ( .A1(n10856), .A2(n11103), .ZN(n11102) );
  INV_X1 U11132 ( .A(n11104), .ZN(n11103) );
  NOR2_X1 U11133 ( .A1(n10855), .A2(n10854), .ZN(n11104) );
  NOR2_X1 U11134 ( .A1(n10624), .A2(n8797), .ZN(n10856) );
  NAND2_X1 U11135 ( .A1(n10854), .A2(n10855), .ZN(n11101) );
  NAND2_X1 U11136 ( .A1(n11105), .A2(n11106), .ZN(n10855) );
  NAND2_X1 U11137 ( .A1(n10883), .A2(n11107), .ZN(n11106) );
  INV_X1 U11138 ( .A(n11108), .ZN(n11107) );
  NOR2_X1 U11139 ( .A1(n10884), .A2(n10882), .ZN(n11108) );
  NOR2_X1 U11140 ( .A1(n10624), .A2(n8314), .ZN(n10883) );
  NAND2_X1 U11141 ( .A1(n10882), .A2(n10884), .ZN(n11105) );
  NAND2_X1 U11142 ( .A1(n11109), .A2(n11110), .ZN(n10884) );
  NAND2_X1 U11143 ( .A1(n10878), .A2(n11111), .ZN(n11110) );
  INV_X1 U11144 ( .A(n11112), .ZN(n11111) );
  NOR2_X1 U11145 ( .A1(n10879), .A2(n10880), .ZN(n11112) );
  NOR2_X1 U11146 ( .A1(n10624), .A2(n9098), .ZN(n10878) );
  NAND2_X1 U11147 ( .A1(n10880), .A2(n10879), .ZN(n11109) );
  NAND2_X1 U11148 ( .A1(n11113), .A2(n11114), .ZN(n10879) );
  NAND2_X1 U11149 ( .A1(b_20_), .A2(n11115), .ZN(n11114) );
  NAND2_X1 U11150 ( .A1(n8299), .A2(n11116), .ZN(n11115) );
  NAND2_X1 U11151 ( .A1(a_31_), .A2(n10876), .ZN(n11116) );
  NAND2_X1 U11152 ( .A1(b_21_), .A2(n11117), .ZN(n11113) );
  NAND2_X1 U11153 ( .A1(n8303), .A2(n11118), .ZN(n11117) );
  NAND2_X1 U11154 ( .A1(a_30_), .A2(n11119), .ZN(n11118) );
  NOR3_X1 U11155 ( .A1(n10876), .A2(n9631), .A3(n10624), .ZN(n10880) );
  XOR2_X1 U11156 ( .A(n11120), .B(n11121), .Z(n10882) );
  XOR2_X1 U11157 ( .A(n11122), .B(n11123), .Z(n11120) );
  XOR2_X1 U11158 ( .A(n11124), .B(n11125), .Z(n10854) );
  XOR2_X1 U11159 ( .A(n11126), .B(n11127), .Z(n11124) );
  XNOR2_X1 U11160 ( .A(n11128), .B(n11129), .ZN(n10834) );
  XNOR2_X1 U11161 ( .A(n11130), .B(n11131), .ZN(n11129) );
  XNOR2_X1 U11162 ( .A(n11132), .B(n11133), .ZN(n10890) );
  NAND2_X1 U11163 ( .A1(n11134), .A2(n11135), .ZN(n11132) );
  XNOR2_X1 U11164 ( .A(n11136), .B(n11137), .ZN(n10799) );
  NAND2_X1 U11165 ( .A1(n11138), .A2(n11139), .ZN(n11136) );
  XNOR2_X1 U11166 ( .A(n11140), .B(n11141), .ZN(n10765) );
  NAND2_X1 U11167 ( .A1(n11142), .A2(n11143), .ZN(n11140) );
  XNOR2_X1 U11168 ( .A(n11144), .B(n11145), .ZN(n10753) );
  XOR2_X1 U11169 ( .A(n11146), .B(n11147), .Z(n11145) );
  NAND2_X1 U11170 ( .A1(b_21_), .A2(a_14_), .ZN(n11147) );
  XNOR2_X1 U11171 ( .A(n11148), .B(n11149), .ZN(n10745) );
  XOR2_X1 U11172 ( .A(n11150), .B(n11151), .Z(n11148) );
  NOR2_X1 U11173 ( .A1(n8996), .A2(n10876), .ZN(n11151) );
  XOR2_X1 U11174 ( .A(n11152), .B(n11153), .Z(n10897) );
  XNOR2_X1 U11175 ( .A(n11154), .B(n11155), .ZN(n11153) );
  XNOR2_X1 U11176 ( .A(n11156), .B(n11157), .ZN(n10721) );
  XNOR2_X1 U11177 ( .A(n11158), .B(n11159), .ZN(n11157) );
  XNOR2_X1 U11178 ( .A(n11160), .B(n11161), .ZN(n10712) );
  NAND2_X1 U11179 ( .A1(n11162), .A2(n11163), .ZN(n11160) );
  XNOR2_X1 U11180 ( .A(n11164), .B(n11165), .ZN(n10909) );
  XOR2_X1 U11181 ( .A(n11166), .B(n11167), .Z(n11165) );
  NAND2_X1 U11182 ( .A1(b_21_), .A2(a_6_), .ZN(n11167) );
  XNOR2_X1 U11183 ( .A(n11168), .B(n11169), .ZN(n10922) );
  XNOR2_X1 U11184 ( .A(n11170), .B(n11171), .ZN(n11169) );
  NAND2_X1 U11185 ( .A1(b_21_), .A2(a_3_), .ZN(n11171) );
  XNOR2_X1 U11186 ( .A(n11172), .B(n11173), .ZN(n10926) );
  XOR2_X1 U11187 ( .A(n11174), .B(n11175), .Z(n11172) );
  NOR2_X1 U11188 ( .A1(n8448), .A2(n10876), .ZN(n11175) );
  XOR2_X1 U11189 ( .A(n11176), .B(n11177), .Z(n8621) );
  XOR2_X1 U11190 ( .A(n11178), .B(n11179), .Z(n11176) );
  NOR2_X1 U11191 ( .A1(n8457), .A2(n10876), .ZN(n11179) );
  NAND3_X1 U11192 ( .A1(n8613), .A2(n8614), .A3(n11180), .ZN(n8504) );
  XNOR2_X1 U11193 ( .A(n8608), .B(n11181), .ZN(n11180) );
  NAND2_X1 U11194 ( .A1(n11182), .A2(n11183), .ZN(n8614) );
  INV_X1 U11195 ( .A(n11184), .ZN(n11183) );
  NOR3_X1 U11196 ( .A1(n8457), .A2(n11185), .A3(n10876), .ZN(n11184) );
  NOR2_X1 U11197 ( .A1(n11178), .A2(n11177), .ZN(n11185) );
  NAND2_X1 U11198 ( .A1(n11177), .A2(n11178), .ZN(n11182) );
  NAND2_X1 U11199 ( .A1(n11186), .A2(n11187), .ZN(n11178) );
  NAND3_X1 U11200 ( .A1(a_1_), .A2(n11188), .A3(b_21_), .ZN(n11187) );
  INV_X1 U11201 ( .A(n11189), .ZN(n11188) );
  NOR2_X1 U11202 ( .A1(n10938), .A2(n10936), .ZN(n11189) );
  NAND2_X1 U11203 ( .A1(n10936), .A2(n10938), .ZN(n11186) );
  NAND2_X1 U11204 ( .A1(n11190), .A2(n11191), .ZN(n10938) );
  NAND3_X1 U11205 ( .A1(a_2_), .A2(n11192), .A3(b_21_), .ZN(n11191) );
  INV_X1 U11206 ( .A(n11193), .ZN(n11192) );
  NOR2_X1 U11207 ( .A1(n11174), .A2(n11173), .ZN(n11193) );
  NAND2_X1 U11208 ( .A1(n11173), .A2(n11174), .ZN(n11190) );
  NAND2_X1 U11209 ( .A1(n11194), .A2(n11195), .ZN(n11174) );
  NAND3_X1 U11210 ( .A1(a_3_), .A2(n11196), .A3(b_21_), .ZN(n11195) );
  NAND2_X1 U11211 ( .A1(n11170), .A2(n11168), .ZN(n11196) );
  INV_X1 U11212 ( .A(n11197), .ZN(n11194) );
  NOR2_X1 U11213 ( .A1(n11168), .A2(n11170), .ZN(n11197) );
  NOR2_X1 U11214 ( .A1(n11198), .A2(n11199), .ZN(n11170) );
  NOR3_X1 U11215 ( .A1(n8439), .A2(n11200), .A3(n10876), .ZN(n11199) );
  NOR2_X1 U11216 ( .A1(n10954), .A2(n10953), .ZN(n11200) );
  INV_X1 U11217 ( .A(n11201), .ZN(n11198) );
  NAND2_X1 U11218 ( .A1(n10953), .A2(n10954), .ZN(n11201) );
  NAND2_X1 U11219 ( .A1(n11202), .A2(n11203), .ZN(n10954) );
  NAND3_X1 U11220 ( .A1(a_5_), .A2(n11204), .A3(b_21_), .ZN(n11203) );
  INV_X1 U11221 ( .A(n11205), .ZN(n11204) );
  NOR2_X1 U11222 ( .A1(n10963), .A2(n10961), .ZN(n11205) );
  NAND2_X1 U11223 ( .A1(n10961), .A2(n10963), .ZN(n11202) );
  NAND2_X1 U11224 ( .A1(n11206), .A2(n11207), .ZN(n10963) );
  INV_X1 U11225 ( .A(n11208), .ZN(n11207) );
  NOR3_X1 U11226 ( .A1(n8430), .A2(n11209), .A3(n10876), .ZN(n11208) );
  NOR2_X1 U11227 ( .A1(n11166), .A2(n11164), .ZN(n11209) );
  NAND2_X1 U11228 ( .A1(n11164), .A2(n11166), .ZN(n11206) );
  NAND2_X1 U11229 ( .A1(n11210), .A2(n11211), .ZN(n11166) );
  NAND3_X1 U11230 ( .A1(a_7_), .A2(n11212), .A3(b_21_), .ZN(n11211) );
  INV_X1 U11231 ( .A(n11213), .ZN(n11212) );
  NOR2_X1 U11232 ( .A1(n10974), .A2(n10973), .ZN(n11213) );
  NAND2_X1 U11233 ( .A1(n10973), .A2(n10974), .ZN(n11210) );
  NAND2_X1 U11234 ( .A1(n11162), .A2(n11214), .ZN(n10974) );
  NAND2_X1 U11235 ( .A1(n11161), .A2(n11163), .ZN(n11214) );
  NAND2_X1 U11236 ( .A1(n11215), .A2(n11216), .ZN(n11163) );
  NAND2_X1 U11237 ( .A1(b_21_), .A2(a_8_), .ZN(n11216) );
  INV_X1 U11238 ( .A(n11217), .ZN(n11215) );
  XNOR2_X1 U11239 ( .A(n11218), .B(n11219), .ZN(n11161) );
  XNOR2_X1 U11240 ( .A(n11220), .B(n11221), .ZN(n11219) );
  NAND2_X1 U11241 ( .A1(a_8_), .A2(n11217), .ZN(n11162) );
  NAND2_X1 U11242 ( .A1(n11222), .A2(n11223), .ZN(n11217) );
  NAND2_X1 U11243 ( .A1(n11159), .A2(n11224), .ZN(n11223) );
  INV_X1 U11244 ( .A(n11225), .ZN(n11224) );
  NOR2_X1 U11245 ( .A1(n11158), .A2(n11156), .ZN(n11225) );
  NOR2_X1 U11246 ( .A1(n10876), .A2(n8971), .ZN(n11159) );
  NAND2_X1 U11247 ( .A1(n11156), .A2(n11158), .ZN(n11222) );
  NAND2_X1 U11248 ( .A1(n11226), .A2(n11227), .ZN(n11158) );
  NAND2_X1 U11249 ( .A1(n10991), .A2(n11228), .ZN(n11227) );
  NAND2_X1 U11250 ( .A1(n10990), .A2(n10989), .ZN(n11228) );
  NOR2_X1 U11251 ( .A1(n10876), .A2(n8402), .ZN(n10991) );
  INV_X1 U11252 ( .A(n11229), .ZN(n11226) );
  NOR2_X1 U11253 ( .A1(n10989), .A2(n10990), .ZN(n11229) );
  NOR2_X1 U11254 ( .A1(n11230), .A2(n11231), .ZN(n10990) );
  INV_X1 U11255 ( .A(n11232), .ZN(n11231) );
  NAND2_X1 U11256 ( .A1(n10999), .A2(n11233), .ZN(n11232) );
  NAND2_X1 U11257 ( .A1(n10996), .A2(n10998), .ZN(n11233) );
  NOR2_X1 U11258 ( .A1(n10876), .A2(n8867), .ZN(n10999) );
  NOR2_X1 U11259 ( .A1(n10998), .A2(n10996), .ZN(n11230) );
  XOR2_X1 U11260 ( .A(n11234), .B(n11235), .Z(n10996) );
  XOR2_X1 U11261 ( .A(n11236), .B(n11237), .Z(n11234) );
  NAND2_X1 U11262 ( .A1(n11238), .A2(n11239), .ZN(n10998) );
  NAND2_X1 U11263 ( .A1(n11152), .A2(n11240), .ZN(n11239) );
  NAND2_X1 U11264 ( .A1(n11155), .A2(n11154), .ZN(n11240) );
  XOR2_X1 U11265 ( .A(n11241), .B(n11242), .Z(n11152) );
  NAND2_X1 U11266 ( .A1(n11243), .A2(n11244), .ZN(n11241) );
  INV_X1 U11267 ( .A(n11245), .ZN(n11238) );
  NOR2_X1 U11268 ( .A1(n11154), .A2(n11155), .ZN(n11245) );
  NOR2_X1 U11269 ( .A1(n10876), .A2(n8393), .ZN(n11155) );
  NAND2_X1 U11270 ( .A1(n11246), .A2(n11247), .ZN(n11154) );
  NAND3_X1 U11271 ( .A1(a_13_), .A2(n11248), .A3(b_21_), .ZN(n11247) );
  INV_X1 U11272 ( .A(n11249), .ZN(n11248) );
  NOR2_X1 U11273 ( .A1(n11150), .A2(n11149), .ZN(n11249) );
  NAND2_X1 U11274 ( .A1(n11149), .A2(n11150), .ZN(n11246) );
  NAND2_X1 U11275 ( .A1(n11250), .A2(n11251), .ZN(n11150) );
  INV_X1 U11276 ( .A(n11252), .ZN(n11251) );
  NOR3_X1 U11277 ( .A1(n9262), .A2(n11253), .A3(n10876), .ZN(n11252) );
  NOR2_X1 U11278 ( .A1(n11146), .A2(n11144), .ZN(n11253) );
  NAND2_X1 U11279 ( .A1(n11144), .A2(n11146), .ZN(n11250) );
  NAND2_X1 U11280 ( .A1(n11254), .A2(n11255), .ZN(n11146) );
  NAND3_X1 U11281 ( .A1(a_15_), .A2(n11256), .A3(b_21_), .ZN(n11255) );
  INV_X1 U11282 ( .A(n11257), .ZN(n11256) );
  NOR2_X1 U11283 ( .A1(n11019), .A2(n11018), .ZN(n11257) );
  NAND2_X1 U11284 ( .A1(n11018), .A2(n11019), .ZN(n11254) );
  NAND2_X1 U11285 ( .A1(n11142), .A2(n11258), .ZN(n11019) );
  NAND2_X1 U11286 ( .A1(n11141), .A2(n11143), .ZN(n11258) );
  NAND2_X1 U11287 ( .A1(n11259), .A2(n11260), .ZN(n11143) );
  NAND2_X1 U11288 ( .A1(b_21_), .A2(a_16_), .ZN(n11260) );
  XNOR2_X1 U11289 ( .A(n11261), .B(n11262), .ZN(n11141) );
  XOR2_X1 U11290 ( .A(n11263), .B(n11264), .Z(n11262) );
  NAND2_X1 U11291 ( .A1(b_20_), .A2(a_17_), .ZN(n11264) );
  NAND2_X1 U11292 ( .A1(a_16_), .A2(n11265), .ZN(n11142) );
  INV_X1 U11293 ( .A(n11259), .ZN(n11265) );
  NOR2_X1 U11294 ( .A1(n11266), .A2(n11267), .ZN(n11259) );
  NOR3_X1 U11295 ( .A1(n8371), .A2(n11268), .A3(n10876), .ZN(n11267) );
  INV_X1 U11296 ( .A(n11269), .ZN(n11268) );
  NAND2_X1 U11297 ( .A1(n11029), .A2(n11031), .ZN(n11269) );
  NOR2_X1 U11298 ( .A1(n11031), .A2(n11029), .ZN(n11266) );
  XNOR2_X1 U11299 ( .A(n11270), .B(n11271), .ZN(n11029) );
  XNOR2_X1 U11300 ( .A(n11272), .B(n11273), .ZN(n11271) );
  NAND2_X1 U11301 ( .A1(n11274), .A2(n11275), .ZN(n11031) );
  NAND2_X1 U11302 ( .A1(n11037), .A2(n11276), .ZN(n11275) );
  NAND2_X1 U11303 ( .A1(n11040), .A2(n11039), .ZN(n11276) );
  XOR2_X1 U11304 ( .A(n11277), .B(n11278), .Z(n11037) );
  XNOR2_X1 U11305 ( .A(n11279), .B(n11280), .ZN(n11277) );
  NOR2_X1 U11306 ( .A1(n8742), .A2(n11119), .ZN(n11280) );
  INV_X1 U11307 ( .A(n11281), .ZN(n11274) );
  NOR2_X1 U11308 ( .A1(n11039), .A2(n11040), .ZN(n11281) );
  NOR2_X1 U11309 ( .A1(n10876), .A2(n9291), .ZN(n11040) );
  NAND2_X1 U11310 ( .A1(n11282), .A2(n11283), .ZN(n11039) );
  NAND3_X1 U11311 ( .A1(a_19_), .A2(n11284), .A3(b_21_), .ZN(n11283) );
  INV_X1 U11312 ( .A(n11285), .ZN(n11284) );
  NOR2_X1 U11313 ( .A1(n11047), .A2(n11045), .ZN(n11285) );
  NAND2_X1 U11314 ( .A1(n11045), .A2(n11047), .ZN(n11282) );
  NAND2_X1 U11315 ( .A1(n11138), .A2(n11286), .ZN(n11047) );
  NAND2_X1 U11316 ( .A1(n11137), .A2(n11139), .ZN(n11286) );
  NAND2_X1 U11317 ( .A1(n11287), .A2(n11288), .ZN(n11139) );
  NAND2_X1 U11318 ( .A1(b_21_), .A2(a_20_), .ZN(n11288) );
  INV_X1 U11319 ( .A(n11289), .ZN(n11287) );
  XNOR2_X1 U11320 ( .A(n11290), .B(n11291), .ZN(n11137) );
  XOR2_X1 U11321 ( .A(n11292), .B(n11293), .Z(n11291) );
  NAND2_X1 U11322 ( .A1(b_20_), .A2(a_21_), .ZN(n11293) );
  NAND2_X1 U11323 ( .A1(a_20_), .A2(n11289), .ZN(n11138) );
  NAND2_X1 U11324 ( .A1(n11294), .A2(n11295), .ZN(n11289) );
  NAND2_X1 U11325 ( .A1(n11057), .A2(n11296), .ZN(n11295) );
  INV_X1 U11326 ( .A(n11297), .ZN(n11296) );
  NOR2_X1 U11327 ( .A1(n11060), .A2(n11059), .ZN(n11297) );
  XNOR2_X1 U11328 ( .A(n11298), .B(n11299), .ZN(n11057) );
  NAND2_X1 U11329 ( .A1(n11300), .A2(n11301), .ZN(n11298) );
  NAND2_X1 U11330 ( .A1(n11059), .A2(n11060), .ZN(n11294) );
  NAND2_X1 U11331 ( .A1(n11067), .A2(n11302), .ZN(n11060) );
  NAND2_X1 U11332 ( .A1(n11066), .A2(n11068), .ZN(n11302) );
  NAND2_X1 U11333 ( .A1(n11303), .A2(n11304), .ZN(n11068) );
  NAND2_X1 U11334 ( .A1(b_21_), .A2(a_22_), .ZN(n11304) );
  INV_X1 U11335 ( .A(n11305), .ZN(n11303) );
  XNOR2_X1 U11336 ( .A(n11306), .B(n11307), .ZN(n11066) );
  NAND2_X1 U11337 ( .A1(n11308), .A2(n11309), .ZN(n11306) );
  NAND2_X1 U11338 ( .A1(a_22_), .A2(n11305), .ZN(n11067) );
  NAND2_X1 U11339 ( .A1(n11134), .A2(n11310), .ZN(n11305) );
  NAND2_X1 U11340 ( .A1(n11133), .A2(n11135), .ZN(n11310) );
  NAND2_X1 U11341 ( .A1(n11311), .A2(n11312), .ZN(n11135) );
  NAND2_X1 U11342 ( .A1(b_21_), .A2(a_23_), .ZN(n11312) );
  INV_X1 U11343 ( .A(n11313), .ZN(n11311) );
  XOR2_X1 U11344 ( .A(n11314), .B(n11315), .Z(n11133) );
  XOR2_X1 U11345 ( .A(n11316), .B(n11317), .Z(n11314) );
  NAND2_X1 U11346 ( .A1(a_23_), .A2(n11313), .ZN(n11134) );
  NAND2_X1 U11347 ( .A1(n11318), .A2(n11319), .ZN(n11313) );
  NAND2_X1 U11348 ( .A1(n11080), .A2(n11320), .ZN(n11319) );
  INV_X1 U11349 ( .A(n11321), .ZN(n11320) );
  NOR2_X1 U11350 ( .A1(n11079), .A2(n11078), .ZN(n11321) );
  NOR2_X1 U11351 ( .A1(n10876), .A2(n8779), .ZN(n11080) );
  NAND2_X1 U11352 ( .A1(n11078), .A2(n11079), .ZN(n11318) );
  NAND2_X1 U11353 ( .A1(n11322), .A2(n11323), .ZN(n11079) );
  NAND2_X1 U11354 ( .A1(n11131), .A2(n11324), .ZN(n11323) );
  NAND2_X1 U11355 ( .A1(n11128), .A2(n11130), .ZN(n11324) );
  NOR2_X1 U11356 ( .A1(n10876), .A2(n8788), .ZN(n11131) );
  INV_X1 U11357 ( .A(n11325), .ZN(n11322) );
  NOR2_X1 U11358 ( .A1(n11130), .A2(n11128), .ZN(n11325) );
  XNOR2_X1 U11359 ( .A(n11326), .B(n11327), .ZN(n11128) );
  XNOR2_X1 U11360 ( .A(n11328), .B(n11329), .ZN(n11327) );
  NAND2_X1 U11361 ( .A1(n11330), .A2(n11331), .ZN(n11130) );
  NAND2_X1 U11362 ( .A1(n11089), .A2(n11332), .ZN(n11331) );
  NAND2_X1 U11363 ( .A1(n11092), .A2(n11091), .ZN(n11332) );
  XNOR2_X1 U11364 ( .A(n11333), .B(n11334), .ZN(n11089) );
  XOR2_X1 U11365 ( .A(n11335), .B(n11336), .Z(n11333) );
  INV_X1 U11366 ( .A(n11337), .ZN(n11330) );
  NOR2_X1 U11367 ( .A1(n11091), .A2(n11092), .ZN(n11337) );
  NOR2_X1 U11368 ( .A1(n10876), .A2(n9344), .ZN(n11092) );
  NAND2_X1 U11369 ( .A1(n11338), .A2(n11339), .ZN(n11091) );
  NAND2_X1 U11370 ( .A1(n11099), .A2(n11340), .ZN(n11339) );
  INV_X1 U11371 ( .A(n11341), .ZN(n11340) );
  NOR2_X1 U11372 ( .A1(n11098), .A2(n11097), .ZN(n11341) );
  NOR2_X1 U11373 ( .A1(n10876), .A2(n8797), .ZN(n11099) );
  NAND2_X1 U11374 ( .A1(n11097), .A2(n11098), .ZN(n11338) );
  NAND2_X1 U11375 ( .A1(n11342), .A2(n11343), .ZN(n11098) );
  NAND2_X1 U11376 ( .A1(n11126), .A2(n11344), .ZN(n11343) );
  INV_X1 U11377 ( .A(n11345), .ZN(n11344) );
  NOR2_X1 U11378 ( .A1(n11127), .A2(n11125), .ZN(n11345) );
  NOR2_X1 U11379 ( .A1(n10876), .A2(n8314), .ZN(n11126) );
  NAND2_X1 U11380 ( .A1(n11125), .A2(n11127), .ZN(n11342) );
  NAND2_X1 U11381 ( .A1(n11346), .A2(n11347), .ZN(n11127) );
  NAND2_X1 U11382 ( .A1(n11121), .A2(n11348), .ZN(n11347) );
  INV_X1 U11383 ( .A(n11349), .ZN(n11348) );
  NOR2_X1 U11384 ( .A1(n11122), .A2(n11123), .ZN(n11349) );
  NOR2_X1 U11385 ( .A1(n10876), .A2(n9098), .ZN(n11121) );
  NAND2_X1 U11386 ( .A1(n11123), .A2(n11122), .ZN(n11346) );
  NAND2_X1 U11387 ( .A1(n11350), .A2(n11351), .ZN(n11122) );
  NAND2_X1 U11388 ( .A1(b_19_), .A2(n11352), .ZN(n11351) );
  NAND2_X1 U11389 ( .A1(n8299), .A2(n11353), .ZN(n11352) );
  NAND2_X1 U11390 ( .A1(a_31_), .A2(n11119), .ZN(n11353) );
  NAND2_X1 U11391 ( .A1(b_20_), .A2(n11354), .ZN(n11350) );
  NAND2_X1 U11392 ( .A1(n8303), .A2(n11355), .ZN(n11354) );
  NAND2_X1 U11393 ( .A1(a_30_), .A2(n11356), .ZN(n11355) );
  NOR3_X1 U11394 ( .A1(n11119), .A2(n9631), .A3(n10876), .ZN(n11123) );
  XOR2_X1 U11395 ( .A(n11357), .B(n11358), .Z(n11125) );
  XOR2_X1 U11396 ( .A(n11359), .B(n11360), .Z(n11357) );
  XOR2_X1 U11397 ( .A(n11361), .B(n11362), .Z(n11097) );
  XOR2_X1 U11398 ( .A(n11363), .B(n11364), .Z(n11361) );
  XNOR2_X1 U11399 ( .A(n11365), .B(n11366), .ZN(n11078) );
  XNOR2_X1 U11400 ( .A(n11367), .B(n11368), .ZN(n11366) );
  XNOR2_X1 U11401 ( .A(n11369), .B(n11370), .ZN(n11045) );
  XNOR2_X1 U11402 ( .A(n11371), .B(n11372), .ZN(n11369) );
  XOR2_X1 U11403 ( .A(n11373), .B(n11374), .Z(n11018) );
  XNOR2_X1 U11404 ( .A(n11375), .B(n11376), .ZN(n11374) );
  NAND2_X1 U11405 ( .A1(b_20_), .A2(a_16_), .ZN(n11376) );
  XNOR2_X1 U11406 ( .A(n11377), .B(n11378), .ZN(n11144) );
  XOR2_X1 U11407 ( .A(n11379), .B(n11380), .Z(n11378) );
  NAND2_X1 U11408 ( .A1(b_20_), .A2(a_15_), .ZN(n11380) );
  XNOR2_X1 U11409 ( .A(n11381), .B(n11382), .ZN(n11149) );
  XOR2_X1 U11410 ( .A(n11383), .B(n11384), .Z(n11381) );
  XNOR2_X1 U11411 ( .A(n11385), .B(n11386), .ZN(n10989) );
  XOR2_X1 U11412 ( .A(n11387), .B(n11388), .Z(n11385) );
  NOR2_X1 U11413 ( .A1(n8867), .A2(n11119), .ZN(n11388) );
  XNOR2_X1 U11414 ( .A(n11389), .B(n11390), .ZN(n11156) );
  XOR2_X1 U11415 ( .A(n11391), .B(n11392), .Z(n11389) );
  XNOR2_X1 U11416 ( .A(n11393), .B(n11394), .ZN(n10973) );
  XNOR2_X1 U11417 ( .A(n11395), .B(n11396), .ZN(n11393) );
  XNOR2_X1 U11418 ( .A(n11397), .B(n11398), .ZN(n11164) );
  XNOR2_X1 U11419 ( .A(n11399), .B(n11400), .ZN(n11398) );
  NAND2_X1 U11420 ( .A1(b_20_), .A2(a_7_), .ZN(n11400) );
  XNOR2_X1 U11421 ( .A(n11401), .B(n11402), .ZN(n10961) );
  NAND2_X1 U11422 ( .A1(n11403), .A2(n11404), .ZN(n11401) );
  XNOR2_X1 U11423 ( .A(n11405), .B(n11406), .ZN(n10953) );
  XOR2_X1 U11424 ( .A(n11407), .B(n11408), .Z(n11405) );
  XOR2_X1 U11425 ( .A(n11409), .B(n11410), .Z(n11168) );
  XNOR2_X1 U11426 ( .A(n11411), .B(n11412), .ZN(n11409) );
  XOR2_X1 U11427 ( .A(n11413), .B(n11414), .Z(n11173) );
  XOR2_X1 U11428 ( .A(n11415), .B(n11416), .Z(n11413) );
  XNOR2_X1 U11429 ( .A(n11417), .B(n11418), .ZN(n10936) );
  XNOR2_X1 U11430 ( .A(n11419), .B(n11420), .ZN(n11418) );
  XOR2_X1 U11431 ( .A(n11421), .B(n11422), .Z(n11177) );
  XOR2_X1 U11432 ( .A(n11423), .B(n11424), .Z(n11421) );
  XNOR2_X1 U11433 ( .A(n11425), .B(n11426), .ZN(n8613) );
  NAND2_X1 U11434 ( .A1(n11427), .A2(n11428), .ZN(n11425) );
  INV_X1 U11435 ( .A(n8512), .ZN(n8602) );
  NOR4_X1 U11436 ( .A1(n8608), .A2(n8607), .A3(n8609), .A4(n8600), .ZN(n8512)
         );
  INV_X1 U11437 ( .A(n11429), .ZN(n8600) );
  NAND2_X1 U11438 ( .A1(n11430), .A2(n11431), .ZN(n11429) );
  INV_X1 U11439 ( .A(n11181), .ZN(n8609) );
  NAND2_X1 U11440 ( .A1(n11427), .A2(n11432), .ZN(n11181) );
  NAND2_X1 U11441 ( .A1(n11426), .A2(n11428), .ZN(n11432) );
  NAND2_X1 U11442 ( .A1(n11433), .A2(n11434), .ZN(n11428) );
  NAND2_X1 U11443 ( .A1(b_20_), .A2(a_0_), .ZN(n11434) );
  INV_X1 U11444 ( .A(n11435), .ZN(n11433) );
  XNOR2_X1 U11445 ( .A(n11436), .B(n11437), .ZN(n11426) );
  XOR2_X1 U11446 ( .A(n11438), .B(n11439), .Z(n11437) );
  NAND2_X1 U11447 ( .A1(b_19_), .A2(a_1_), .ZN(n11439) );
  NAND2_X1 U11448 ( .A1(a_0_), .A2(n11435), .ZN(n11427) );
  NAND2_X1 U11449 ( .A1(n11440), .A2(n11441), .ZN(n11435) );
  NAND2_X1 U11450 ( .A1(n11424), .A2(n11442), .ZN(n11441) );
  INV_X1 U11451 ( .A(n11443), .ZN(n11442) );
  NOR2_X1 U11452 ( .A1(n11423), .A2(n11422), .ZN(n11443) );
  NOR2_X1 U11453 ( .A1(n11119), .A2(n8569), .ZN(n11424) );
  NAND2_X1 U11454 ( .A1(n11422), .A2(n11423), .ZN(n11440) );
  NAND2_X1 U11455 ( .A1(n11444), .A2(n11445), .ZN(n11423) );
  NAND2_X1 U11456 ( .A1(n11420), .A2(n11446), .ZN(n11445) );
  INV_X1 U11457 ( .A(n11447), .ZN(n11446) );
  NOR2_X1 U11458 ( .A1(n11419), .A2(n11417), .ZN(n11447) );
  NOR2_X1 U11459 ( .A1(n11119), .A2(n8448), .ZN(n11420) );
  NAND2_X1 U11460 ( .A1(n11417), .A2(n11419), .ZN(n11444) );
  NAND2_X1 U11461 ( .A1(n11448), .A2(n11449), .ZN(n11419) );
  NAND2_X1 U11462 ( .A1(n11416), .A2(n11450), .ZN(n11449) );
  INV_X1 U11463 ( .A(n11451), .ZN(n11450) );
  NOR2_X1 U11464 ( .A1(n11415), .A2(n11414), .ZN(n11451) );
  NOR2_X1 U11465 ( .A1(n11119), .A2(n8900), .ZN(n11416) );
  NAND2_X1 U11466 ( .A1(n11414), .A2(n11415), .ZN(n11448) );
  NAND2_X1 U11467 ( .A1(n11452), .A2(n11453), .ZN(n11415) );
  NAND2_X1 U11468 ( .A1(n11412), .A2(n11454), .ZN(n11453) );
  INV_X1 U11469 ( .A(n11455), .ZN(n11454) );
  NOR2_X1 U11470 ( .A1(n11410), .A2(n11411), .ZN(n11455) );
  NOR2_X1 U11471 ( .A1(n11119), .A2(n8439), .ZN(n11412) );
  NAND2_X1 U11472 ( .A1(n11411), .A2(n11410), .ZN(n11452) );
  XNOR2_X1 U11473 ( .A(n11456), .B(n11457), .ZN(n11410) );
  XOR2_X1 U11474 ( .A(n11458), .B(n11459), .Z(n11457) );
  NAND2_X1 U11475 ( .A1(b_19_), .A2(a_5_), .ZN(n11459) );
  NOR2_X1 U11476 ( .A1(n11460), .A2(n11461), .ZN(n11411) );
  INV_X1 U11477 ( .A(n11462), .ZN(n11461) );
  NAND2_X1 U11478 ( .A1(n11406), .A2(n11463), .ZN(n11462) );
  NAND2_X1 U11479 ( .A1(n11408), .A2(n11407), .ZN(n11463) );
  XNOR2_X1 U11480 ( .A(n11464), .B(n11465), .ZN(n11406) );
  XOR2_X1 U11481 ( .A(n11466), .B(n11467), .Z(n11464) );
  NOR2_X1 U11482 ( .A1(n8430), .A2(n11356), .ZN(n11467) );
  NOR2_X1 U11483 ( .A1(n11407), .A2(n11408), .ZN(n11460) );
  NOR2_X1 U11484 ( .A1(n11119), .A2(n8938), .ZN(n11408) );
  NAND2_X1 U11485 ( .A1(n11403), .A2(n11468), .ZN(n11407) );
  NAND2_X1 U11486 ( .A1(n11402), .A2(n11404), .ZN(n11468) );
  NAND2_X1 U11487 ( .A1(n11469), .A2(n11470), .ZN(n11404) );
  NAND2_X1 U11488 ( .A1(b_20_), .A2(a_6_), .ZN(n11470) );
  INV_X1 U11489 ( .A(n11471), .ZN(n11469) );
  XNOR2_X1 U11490 ( .A(n11472), .B(n11473), .ZN(n11402) );
  XOR2_X1 U11491 ( .A(n11474), .B(n11475), .Z(n11473) );
  NAND2_X1 U11492 ( .A1(b_19_), .A2(a_7_), .ZN(n11475) );
  NAND2_X1 U11493 ( .A1(a_6_), .A2(n11471), .ZN(n11403) );
  NAND2_X1 U11494 ( .A1(n11476), .A2(n11477), .ZN(n11471) );
  NAND3_X1 U11495 ( .A1(a_7_), .A2(n11478), .A3(b_20_), .ZN(n11477) );
  NAND2_X1 U11496 ( .A1(n11399), .A2(n11479), .ZN(n11478) );
  INV_X1 U11497 ( .A(n11397), .ZN(n11479) );
  NAND2_X1 U11498 ( .A1(n11397), .A2(n11480), .ZN(n11476) );
  INV_X1 U11499 ( .A(n11399), .ZN(n11480) );
  NOR2_X1 U11500 ( .A1(n11481), .A2(n11482), .ZN(n11399) );
  INV_X1 U11501 ( .A(n11483), .ZN(n11482) );
  NAND2_X1 U11502 ( .A1(n11396), .A2(n11484), .ZN(n11483) );
  NAND2_X1 U11503 ( .A1(n11395), .A2(n11394), .ZN(n11484) );
  NOR2_X1 U11504 ( .A1(n11119), .A2(n8968), .ZN(n11396) );
  NOR2_X1 U11505 ( .A1(n11394), .A2(n11395), .ZN(n11481) );
  NOR2_X1 U11506 ( .A1(n11485), .A2(n11486), .ZN(n11395) );
  INV_X1 U11507 ( .A(n11487), .ZN(n11486) );
  NAND2_X1 U11508 ( .A1(n11221), .A2(n11488), .ZN(n11487) );
  NAND2_X1 U11509 ( .A1(n11218), .A2(n11220), .ZN(n11488) );
  NOR2_X1 U11510 ( .A1(n11119), .A2(n8971), .ZN(n11221) );
  NOR2_X1 U11511 ( .A1(n11220), .A2(n11218), .ZN(n11485) );
  XNOR2_X1 U11512 ( .A(n11489), .B(n11490), .ZN(n11218) );
  XNOR2_X1 U11513 ( .A(n11491), .B(n11492), .ZN(n11490) );
  NAND2_X1 U11514 ( .A1(b_19_), .A2(a_10_), .ZN(n11492) );
  NAND2_X1 U11515 ( .A1(n11493), .A2(n11494), .ZN(n11220) );
  NAND2_X1 U11516 ( .A1(n11390), .A2(n11495), .ZN(n11494) );
  NAND2_X1 U11517 ( .A1(n11392), .A2(n11391), .ZN(n11495) );
  XOR2_X1 U11518 ( .A(n11496), .B(n11497), .Z(n11390) );
  XNOR2_X1 U11519 ( .A(n11498), .B(n11499), .ZN(n11497) );
  INV_X1 U11520 ( .A(n11500), .ZN(n11493) );
  NOR2_X1 U11521 ( .A1(n11391), .A2(n11392), .ZN(n11500) );
  NOR2_X1 U11522 ( .A1(n11119), .A2(n8402), .ZN(n11392) );
  NAND2_X1 U11523 ( .A1(n11501), .A2(n11502), .ZN(n11391) );
  NAND3_X1 U11524 ( .A1(a_11_), .A2(n11503), .A3(b_20_), .ZN(n11502) );
  NAND2_X1 U11525 ( .A1(n11386), .A2(n11387), .ZN(n11503) );
  INV_X1 U11526 ( .A(n11504), .ZN(n11501) );
  NOR2_X1 U11527 ( .A1(n11387), .A2(n11386), .ZN(n11504) );
  XNOR2_X1 U11528 ( .A(n11505), .B(n11506), .ZN(n11386) );
  XNOR2_X1 U11529 ( .A(n11507), .B(n11508), .ZN(n11506) );
  NAND2_X1 U11530 ( .A1(n11509), .A2(n11510), .ZN(n11387) );
  NAND2_X1 U11531 ( .A1(n11235), .A2(n11511), .ZN(n11510) );
  NAND2_X1 U11532 ( .A1(n11237), .A2(n11236), .ZN(n11511) );
  XNOR2_X1 U11533 ( .A(n11512), .B(n11513), .ZN(n11235) );
  XNOR2_X1 U11534 ( .A(n11514), .B(n11515), .ZN(n11513) );
  NAND2_X1 U11535 ( .A1(b_19_), .A2(a_13_), .ZN(n11515) );
  INV_X1 U11536 ( .A(n11516), .ZN(n11509) );
  NOR2_X1 U11537 ( .A1(n11236), .A2(n11237), .ZN(n11516) );
  NOR2_X1 U11538 ( .A1(n11119), .A2(n8393), .ZN(n11237) );
  NAND2_X1 U11539 ( .A1(n11243), .A2(n11517), .ZN(n11236) );
  NAND2_X1 U11540 ( .A1(n11242), .A2(n11244), .ZN(n11517) );
  NAND2_X1 U11541 ( .A1(n11518), .A2(n11519), .ZN(n11244) );
  NAND2_X1 U11542 ( .A1(b_20_), .A2(a_13_), .ZN(n11518) );
  XOR2_X1 U11543 ( .A(n11520), .B(n11521), .Z(n11242) );
  XOR2_X1 U11544 ( .A(n11522), .B(n11523), .Z(n11520) );
  NOR2_X1 U11545 ( .A1(n9262), .A2(n11356), .ZN(n11523) );
  INV_X1 U11546 ( .A(n11524), .ZN(n11243) );
  NOR2_X1 U11547 ( .A1(n11519), .A2(n8996), .ZN(n11524) );
  NAND2_X1 U11548 ( .A1(n11525), .A2(n11526), .ZN(n11519) );
  NAND2_X1 U11549 ( .A1(n11382), .A2(n11527), .ZN(n11526) );
  NAND2_X1 U11550 ( .A1(n11384), .A2(n11383), .ZN(n11527) );
  XNOR2_X1 U11551 ( .A(n11528), .B(n11529), .ZN(n11382) );
  XNOR2_X1 U11552 ( .A(n11530), .B(n11531), .ZN(n11529) );
  NAND2_X1 U11553 ( .A1(b_19_), .A2(a_15_), .ZN(n11531) );
  INV_X1 U11554 ( .A(n11532), .ZN(n11525) );
  NOR2_X1 U11555 ( .A1(n11383), .A2(n11384), .ZN(n11532) );
  NOR2_X1 U11556 ( .A1(n11119), .A2(n9262), .ZN(n11384) );
  NAND2_X1 U11557 ( .A1(n11533), .A2(n11534), .ZN(n11383) );
  NAND3_X1 U11558 ( .A1(a_15_), .A2(n11535), .A3(b_20_), .ZN(n11534) );
  INV_X1 U11559 ( .A(n11536), .ZN(n11535) );
  NOR2_X1 U11560 ( .A1(n11379), .A2(n11377), .ZN(n11536) );
  NAND2_X1 U11561 ( .A1(n11377), .A2(n11379), .ZN(n11533) );
  NAND2_X1 U11562 ( .A1(n11537), .A2(n11538), .ZN(n11379) );
  NAND3_X1 U11563 ( .A1(a_16_), .A2(n11539), .A3(b_20_), .ZN(n11538) );
  NAND2_X1 U11564 ( .A1(n11375), .A2(n11373), .ZN(n11539) );
  INV_X1 U11565 ( .A(n11540), .ZN(n11537) );
  NOR2_X1 U11566 ( .A1(n11373), .A2(n11375), .ZN(n11540) );
  NOR2_X1 U11567 ( .A1(n11541), .A2(n11542), .ZN(n11375) );
  INV_X1 U11568 ( .A(n11543), .ZN(n11542) );
  NAND3_X1 U11569 ( .A1(a_17_), .A2(n11544), .A3(b_20_), .ZN(n11543) );
  NAND2_X1 U11570 ( .A1(n11261), .A2(n11263), .ZN(n11544) );
  NOR2_X1 U11571 ( .A1(n11263), .A2(n11261), .ZN(n11541) );
  XOR2_X1 U11572 ( .A(n11545), .B(n11546), .Z(n11261) );
  XNOR2_X1 U11573 ( .A(n11547), .B(n11548), .ZN(n11546) );
  NAND2_X1 U11574 ( .A1(n11549), .A2(n11550), .ZN(n11263) );
  NAND2_X1 U11575 ( .A1(n11270), .A2(n11551), .ZN(n11550) );
  INV_X1 U11576 ( .A(n11552), .ZN(n11551) );
  NOR2_X1 U11577 ( .A1(n11273), .A2(n11272), .ZN(n11552) );
  XOR2_X1 U11578 ( .A(n11553), .B(n11554), .Z(n11270) );
  XNOR2_X1 U11579 ( .A(n11555), .B(n11556), .ZN(n11554) );
  NAND2_X1 U11580 ( .A1(n11272), .A2(n11273), .ZN(n11549) );
  NAND2_X1 U11581 ( .A1(b_20_), .A2(a_18_), .ZN(n11273) );
  NOR2_X1 U11582 ( .A1(n11557), .A2(n11558), .ZN(n11272) );
  INV_X1 U11583 ( .A(n11559), .ZN(n11558) );
  NAND3_X1 U11584 ( .A1(a_19_), .A2(n11560), .A3(b_20_), .ZN(n11559) );
  NAND2_X1 U11585 ( .A1(n11279), .A2(n11278), .ZN(n11560) );
  NOR2_X1 U11586 ( .A1(n11278), .A2(n11279), .ZN(n11557) );
  NOR2_X1 U11587 ( .A1(n11561), .A2(n11562), .ZN(n11279) );
  INV_X1 U11588 ( .A(n11563), .ZN(n11562) );
  NAND2_X1 U11589 ( .A1(n11372), .A2(n11564), .ZN(n11563) );
  NAND2_X1 U11590 ( .A1(n11371), .A2(n11370), .ZN(n11564) );
  NOR2_X1 U11591 ( .A1(n11370), .A2(n11371), .ZN(n11561) );
  NOR2_X1 U11592 ( .A1(n11565), .A2(n11566), .ZN(n11371) );
  NOR3_X1 U11593 ( .A1(n8759), .A2(n11567), .A3(n11119), .ZN(n11566) );
  NOR2_X1 U11594 ( .A1(n11292), .A2(n11290), .ZN(n11567) );
  INV_X1 U11595 ( .A(n11568), .ZN(n11565) );
  NAND2_X1 U11596 ( .A1(n11290), .A2(n11292), .ZN(n11568) );
  NAND2_X1 U11597 ( .A1(n11300), .A2(n11569), .ZN(n11292) );
  NAND2_X1 U11598 ( .A1(n11299), .A2(n11301), .ZN(n11569) );
  NAND2_X1 U11599 ( .A1(n11570), .A2(n11571), .ZN(n11301) );
  NAND2_X1 U11600 ( .A1(b_20_), .A2(a_22_), .ZN(n11571) );
  INV_X1 U11601 ( .A(n11572), .ZN(n11570) );
  XNOR2_X1 U11602 ( .A(n11573), .B(n11574), .ZN(n11299) );
  NAND2_X1 U11603 ( .A1(n11575), .A2(n11576), .ZN(n11573) );
  NAND2_X1 U11604 ( .A1(a_22_), .A2(n11572), .ZN(n11300) );
  NAND2_X1 U11605 ( .A1(n11308), .A2(n11577), .ZN(n11572) );
  NAND2_X1 U11606 ( .A1(n11307), .A2(n11309), .ZN(n11577) );
  NAND2_X1 U11607 ( .A1(n11578), .A2(n11579), .ZN(n11309) );
  NAND2_X1 U11608 ( .A1(b_20_), .A2(a_23_), .ZN(n11579) );
  INV_X1 U11609 ( .A(n11580), .ZN(n11578) );
  XOR2_X1 U11610 ( .A(n11581), .B(n11582), .Z(n11307) );
  XOR2_X1 U11611 ( .A(n11583), .B(n11584), .Z(n11581) );
  NAND2_X1 U11612 ( .A1(a_23_), .A2(n11580), .ZN(n11308) );
  NAND2_X1 U11613 ( .A1(n11585), .A2(n11586), .ZN(n11580) );
  NAND2_X1 U11614 ( .A1(n11317), .A2(n11587), .ZN(n11586) );
  INV_X1 U11615 ( .A(n11588), .ZN(n11587) );
  NOR2_X1 U11616 ( .A1(n11316), .A2(n11315), .ZN(n11588) );
  NOR2_X1 U11617 ( .A1(n11119), .A2(n8779), .ZN(n11317) );
  NAND2_X1 U11618 ( .A1(n11315), .A2(n11316), .ZN(n11585) );
  NAND2_X1 U11619 ( .A1(n11589), .A2(n11590), .ZN(n11316) );
  NAND2_X1 U11620 ( .A1(n11368), .A2(n11591), .ZN(n11590) );
  NAND2_X1 U11621 ( .A1(n11365), .A2(n11367), .ZN(n11591) );
  NOR2_X1 U11622 ( .A1(n11119), .A2(n8788), .ZN(n11368) );
  INV_X1 U11623 ( .A(n11592), .ZN(n11589) );
  NOR2_X1 U11624 ( .A1(n11367), .A2(n11365), .ZN(n11592) );
  XNOR2_X1 U11625 ( .A(n11593), .B(n11594), .ZN(n11365) );
  XNOR2_X1 U11626 ( .A(n11595), .B(n11596), .ZN(n11594) );
  NAND2_X1 U11627 ( .A1(n11597), .A2(n11598), .ZN(n11367) );
  NAND2_X1 U11628 ( .A1(n11326), .A2(n11599), .ZN(n11598) );
  NAND2_X1 U11629 ( .A1(n11329), .A2(n11328), .ZN(n11599) );
  XNOR2_X1 U11630 ( .A(n11600), .B(n11601), .ZN(n11326) );
  XOR2_X1 U11631 ( .A(n11602), .B(n11603), .Z(n11600) );
  INV_X1 U11632 ( .A(n11604), .ZN(n11597) );
  NOR2_X1 U11633 ( .A1(n11328), .A2(n11329), .ZN(n11604) );
  NOR2_X1 U11634 ( .A1(n11119), .A2(n9344), .ZN(n11329) );
  NAND2_X1 U11635 ( .A1(n11605), .A2(n11606), .ZN(n11328) );
  NAND2_X1 U11636 ( .A1(n11336), .A2(n11607), .ZN(n11606) );
  INV_X1 U11637 ( .A(n11608), .ZN(n11607) );
  NOR2_X1 U11638 ( .A1(n11335), .A2(n11334), .ZN(n11608) );
  NOR2_X1 U11639 ( .A1(n11119), .A2(n8797), .ZN(n11336) );
  NAND2_X1 U11640 ( .A1(n11334), .A2(n11335), .ZN(n11605) );
  NAND2_X1 U11641 ( .A1(n11609), .A2(n11610), .ZN(n11335) );
  NAND2_X1 U11642 ( .A1(n11363), .A2(n11611), .ZN(n11610) );
  INV_X1 U11643 ( .A(n11612), .ZN(n11611) );
  NOR2_X1 U11644 ( .A1(n11364), .A2(n11362), .ZN(n11612) );
  NOR2_X1 U11645 ( .A1(n11119), .A2(n8314), .ZN(n11363) );
  NAND2_X1 U11646 ( .A1(n11362), .A2(n11364), .ZN(n11609) );
  NAND2_X1 U11647 ( .A1(n11613), .A2(n11614), .ZN(n11364) );
  NAND2_X1 U11648 ( .A1(n11358), .A2(n11615), .ZN(n11614) );
  INV_X1 U11649 ( .A(n11616), .ZN(n11615) );
  NOR2_X1 U11650 ( .A1(n11359), .A2(n11360), .ZN(n11616) );
  NOR2_X1 U11651 ( .A1(n11119), .A2(n9098), .ZN(n11358) );
  NAND2_X1 U11652 ( .A1(n11360), .A2(n11359), .ZN(n11613) );
  NAND2_X1 U11653 ( .A1(n11617), .A2(n11618), .ZN(n11359) );
  NAND2_X1 U11654 ( .A1(b_18_), .A2(n11619), .ZN(n11618) );
  NAND2_X1 U11655 ( .A1(n8299), .A2(n11620), .ZN(n11619) );
  NAND2_X1 U11656 ( .A1(a_31_), .A2(n11356), .ZN(n11620) );
  NAND2_X1 U11657 ( .A1(b_19_), .A2(n11621), .ZN(n11617) );
  NAND2_X1 U11658 ( .A1(n8303), .A2(n11622), .ZN(n11621) );
  NAND2_X1 U11659 ( .A1(a_30_), .A2(n11623), .ZN(n11622) );
  NOR3_X1 U11660 ( .A1(n11356), .A2(n9631), .A3(n11119), .ZN(n11360) );
  XOR2_X1 U11661 ( .A(n11624), .B(n11625), .Z(n11362) );
  XOR2_X1 U11662 ( .A(n11626), .B(n11627), .Z(n11624) );
  XOR2_X1 U11663 ( .A(n11628), .B(n11629), .Z(n11334) );
  XOR2_X1 U11664 ( .A(n11630), .B(n11631), .Z(n11628) );
  XNOR2_X1 U11665 ( .A(n11632), .B(n11633), .ZN(n11315) );
  XNOR2_X1 U11666 ( .A(n11634), .B(n11635), .ZN(n11633) );
  XNOR2_X1 U11667 ( .A(n11636), .B(n11637), .ZN(n11290) );
  NAND2_X1 U11668 ( .A1(n11638), .A2(n11639), .ZN(n11636) );
  XOR2_X1 U11669 ( .A(n11640), .B(n11641), .Z(n11370) );
  XOR2_X1 U11670 ( .A(n11642), .B(n11643), .Z(n11641) );
  NAND2_X1 U11671 ( .A1(b_19_), .A2(a_21_), .ZN(n11643) );
  XOR2_X1 U11672 ( .A(n11644), .B(n11645), .Z(n11278) );
  XOR2_X1 U11673 ( .A(n11646), .B(n11647), .Z(n11644) );
  XOR2_X1 U11674 ( .A(n11648), .B(n11649), .Z(n11373) );
  XNOR2_X1 U11675 ( .A(n11650), .B(n11651), .ZN(n11648) );
  XOR2_X1 U11676 ( .A(n11652), .B(n11653), .Z(n11377) );
  XNOR2_X1 U11677 ( .A(n11654), .B(n11655), .ZN(n11653) );
  XNOR2_X1 U11678 ( .A(n11656), .B(n11657), .ZN(n11394) );
  XNOR2_X1 U11679 ( .A(n11658), .B(n11659), .ZN(n11657) );
  NAND2_X1 U11680 ( .A1(b_19_), .A2(a_9_), .ZN(n11659) );
  XOR2_X1 U11681 ( .A(n11660), .B(n11661), .Z(n11397) );
  XNOR2_X1 U11682 ( .A(n11662), .B(n11663), .ZN(n11661) );
  NAND2_X1 U11683 ( .A1(b_19_), .A2(a_8_), .ZN(n11663) );
  XOR2_X1 U11684 ( .A(n11664), .B(n11665), .Z(n11414) );
  XOR2_X1 U11685 ( .A(n11666), .B(n11667), .Z(n11664) );
  NOR2_X1 U11686 ( .A1(n8439), .A2(n11356), .ZN(n11667) );
  XNOR2_X1 U11687 ( .A(n11668), .B(n11669), .ZN(n11417) );
  XOR2_X1 U11688 ( .A(n11670), .B(n11671), .Z(n11669) );
  NAND2_X1 U11689 ( .A1(b_19_), .A2(a_3_), .ZN(n11671) );
  XNOR2_X1 U11690 ( .A(n11672), .B(n11673), .ZN(n11422) );
  XOR2_X1 U11691 ( .A(n11674), .B(n11675), .Z(n11673) );
  NAND2_X1 U11692 ( .A1(b_19_), .A2(a_2_), .ZN(n11675) );
  NOR2_X1 U11693 ( .A1(n11431), .A2(n11430), .ZN(n8607) );
  XNOR2_X1 U11694 ( .A(n11676), .B(n11677), .ZN(n11430) );
  NAND2_X1 U11695 ( .A1(n11678), .A2(n11679), .ZN(n11676) );
  NAND2_X1 U11696 ( .A1(n11680), .A2(n11681), .ZN(n11431) );
  NAND3_X1 U11697 ( .A1(a_0_), .A2(n11682), .A3(b_19_), .ZN(n11681) );
  INV_X1 U11698 ( .A(n11683), .ZN(n11682) );
  NOR2_X1 U11699 ( .A1(n11684), .A2(n11685), .ZN(n11683) );
  NAND2_X1 U11700 ( .A1(n11685), .A2(n11684), .ZN(n11680) );
  XNOR2_X1 U11701 ( .A(n11686), .B(n11685), .ZN(n8608) );
  XNOR2_X1 U11702 ( .A(n11687), .B(n11688), .ZN(n11685) );
  NAND2_X1 U11703 ( .A1(n11689), .A2(n11690), .ZN(n11687) );
  XOR2_X1 U11704 ( .A(n11684), .B(n11691), .Z(n11686) );
  NOR2_X1 U11705 ( .A1(n8457), .A2(n11356), .ZN(n11691) );
  NAND2_X1 U11706 ( .A1(n11692), .A2(n11693), .ZN(n11684) );
  INV_X1 U11707 ( .A(n11694), .ZN(n11693) );
  NOR3_X1 U11708 ( .A1(n8569), .A2(n11695), .A3(n11356), .ZN(n11694) );
  NOR2_X1 U11709 ( .A1(n11438), .A2(n11436), .ZN(n11695) );
  NAND2_X1 U11710 ( .A1(n11436), .A2(n11438), .ZN(n11692) );
  NAND2_X1 U11711 ( .A1(n11696), .A2(n11697), .ZN(n11438) );
  NAND3_X1 U11712 ( .A1(a_2_), .A2(n11698), .A3(b_19_), .ZN(n11697) );
  INV_X1 U11713 ( .A(n11699), .ZN(n11698) );
  NOR2_X1 U11714 ( .A1(n11674), .A2(n11672), .ZN(n11699) );
  NAND2_X1 U11715 ( .A1(n11672), .A2(n11674), .ZN(n11696) );
  NAND2_X1 U11716 ( .A1(n11700), .A2(n11701), .ZN(n11674) );
  INV_X1 U11717 ( .A(n11702), .ZN(n11701) );
  NOR3_X1 U11718 ( .A1(n8900), .A2(n11703), .A3(n11356), .ZN(n11702) );
  NOR2_X1 U11719 ( .A1(n11670), .A2(n11668), .ZN(n11703) );
  NAND2_X1 U11720 ( .A1(n11668), .A2(n11670), .ZN(n11700) );
  NAND2_X1 U11721 ( .A1(n11704), .A2(n11705), .ZN(n11670) );
  NAND3_X1 U11722 ( .A1(a_4_), .A2(n11706), .A3(b_19_), .ZN(n11705) );
  INV_X1 U11723 ( .A(n11707), .ZN(n11706) );
  NOR2_X1 U11724 ( .A1(n11666), .A2(n11665), .ZN(n11707) );
  NAND2_X1 U11725 ( .A1(n11665), .A2(n11666), .ZN(n11704) );
  NAND2_X1 U11726 ( .A1(n11708), .A2(n11709), .ZN(n11666) );
  INV_X1 U11727 ( .A(n11710), .ZN(n11709) );
  NOR3_X1 U11728 ( .A1(n8938), .A2(n11711), .A3(n11356), .ZN(n11710) );
  NOR2_X1 U11729 ( .A1(n11458), .A2(n11456), .ZN(n11711) );
  NAND2_X1 U11730 ( .A1(n11456), .A2(n11458), .ZN(n11708) );
  NAND2_X1 U11731 ( .A1(n11712), .A2(n11713), .ZN(n11458) );
  NAND3_X1 U11732 ( .A1(a_6_), .A2(n11714), .A3(b_19_), .ZN(n11713) );
  INV_X1 U11733 ( .A(n11715), .ZN(n11714) );
  NOR2_X1 U11734 ( .A1(n11466), .A2(n11465), .ZN(n11715) );
  NAND2_X1 U11735 ( .A1(n11465), .A2(n11466), .ZN(n11712) );
  NAND2_X1 U11736 ( .A1(n11716), .A2(n11717), .ZN(n11466) );
  INV_X1 U11737 ( .A(n11718), .ZN(n11717) );
  NOR3_X1 U11738 ( .A1(n8425), .A2(n11719), .A3(n11356), .ZN(n11718) );
  NOR2_X1 U11739 ( .A1(n11474), .A2(n11472), .ZN(n11719) );
  NAND2_X1 U11740 ( .A1(n11472), .A2(n11474), .ZN(n11716) );
  NAND2_X1 U11741 ( .A1(n11720), .A2(n11721), .ZN(n11474) );
  NAND3_X1 U11742 ( .A1(a_8_), .A2(n11722), .A3(b_19_), .ZN(n11721) );
  NAND2_X1 U11743 ( .A1(n11662), .A2(n11660), .ZN(n11722) );
  INV_X1 U11744 ( .A(n11723), .ZN(n11720) );
  NOR2_X1 U11745 ( .A1(n11660), .A2(n11662), .ZN(n11723) );
  NOR2_X1 U11746 ( .A1(n11724), .A2(n11725), .ZN(n11662) );
  INV_X1 U11747 ( .A(n11726), .ZN(n11725) );
  NAND3_X1 U11748 ( .A1(a_9_), .A2(n11727), .A3(b_19_), .ZN(n11726) );
  NAND2_X1 U11749 ( .A1(n11658), .A2(n11656), .ZN(n11727) );
  NOR2_X1 U11750 ( .A1(n11656), .A2(n11658), .ZN(n11724) );
  NOR2_X1 U11751 ( .A1(n11728), .A2(n11729), .ZN(n11658) );
  INV_X1 U11752 ( .A(n11730), .ZN(n11729) );
  NAND3_X1 U11753 ( .A1(a_10_), .A2(n11731), .A3(b_19_), .ZN(n11730) );
  NAND2_X1 U11754 ( .A1(n11491), .A2(n11489), .ZN(n11731) );
  NOR2_X1 U11755 ( .A1(n11489), .A2(n11491), .ZN(n11728) );
  NOR2_X1 U11756 ( .A1(n11732), .A2(n11733), .ZN(n11491) );
  INV_X1 U11757 ( .A(n11734), .ZN(n11733) );
  NAND2_X1 U11758 ( .A1(n11499), .A2(n11735), .ZN(n11734) );
  NAND2_X1 U11759 ( .A1(n11496), .A2(n11498), .ZN(n11735) );
  NOR2_X1 U11760 ( .A1(n11356), .A2(n8867), .ZN(n11499) );
  NOR2_X1 U11761 ( .A1(n11498), .A2(n11496), .ZN(n11732) );
  XOR2_X1 U11762 ( .A(n11736), .B(n11737), .Z(n11496) );
  XNOR2_X1 U11763 ( .A(n11738), .B(n11739), .ZN(n11736) );
  NOR2_X1 U11764 ( .A1(n8393), .A2(n11623), .ZN(n11739) );
  NAND2_X1 U11765 ( .A1(n11740), .A2(n11741), .ZN(n11498) );
  NAND2_X1 U11766 ( .A1(n11505), .A2(n11742), .ZN(n11741) );
  NAND2_X1 U11767 ( .A1(n11508), .A2(n11507), .ZN(n11742) );
  XOR2_X1 U11768 ( .A(n11743), .B(n11744), .Z(n11505) );
  XNOR2_X1 U11769 ( .A(n11745), .B(n11746), .ZN(n11743) );
  NOR2_X1 U11770 ( .A1(n8996), .A2(n11623), .ZN(n11746) );
  INV_X1 U11771 ( .A(n11747), .ZN(n11740) );
  NOR2_X1 U11772 ( .A1(n11507), .A2(n11508), .ZN(n11747) );
  NOR2_X1 U11773 ( .A1(n11356), .A2(n8393), .ZN(n11508) );
  NAND2_X1 U11774 ( .A1(n11748), .A2(n11749), .ZN(n11507) );
  NAND3_X1 U11775 ( .A1(a_13_), .A2(n11750), .A3(b_19_), .ZN(n11749) );
  NAND2_X1 U11776 ( .A1(n11514), .A2(n11512), .ZN(n11750) );
  INV_X1 U11777 ( .A(n11751), .ZN(n11748) );
  NOR2_X1 U11778 ( .A1(n11512), .A2(n11514), .ZN(n11751) );
  NOR2_X1 U11779 ( .A1(n11752), .A2(n11753), .ZN(n11514) );
  NOR3_X1 U11780 ( .A1(n9262), .A2(n11754), .A3(n11356), .ZN(n11753) );
  NOR2_X1 U11781 ( .A1(n11522), .A2(n11521), .ZN(n11754) );
  INV_X1 U11782 ( .A(n11755), .ZN(n11752) );
  NAND2_X1 U11783 ( .A1(n11521), .A2(n11522), .ZN(n11755) );
  NAND2_X1 U11784 ( .A1(n11756), .A2(n11757), .ZN(n11522) );
  NAND3_X1 U11785 ( .A1(a_15_), .A2(n11758), .A3(b_19_), .ZN(n11757) );
  INV_X1 U11786 ( .A(n11759), .ZN(n11758) );
  NOR2_X1 U11787 ( .A1(n11528), .A2(n11530), .ZN(n11759) );
  NAND2_X1 U11788 ( .A1(n11530), .A2(n11528), .ZN(n11756) );
  XNOR2_X1 U11789 ( .A(n11760), .B(n11761), .ZN(n11528) );
  XOR2_X1 U11790 ( .A(n11762), .B(n11763), .Z(n11761) );
  NAND2_X1 U11791 ( .A1(b_18_), .A2(a_16_), .ZN(n11763) );
  NOR2_X1 U11792 ( .A1(n11764), .A2(n11765), .ZN(n11530) );
  INV_X1 U11793 ( .A(n11766), .ZN(n11765) );
  NAND2_X1 U11794 ( .A1(n11652), .A2(n11767), .ZN(n11766) );
  NAND2_X1 U11795 ( .A1(n11655), .A2(n11654), .ZN(n11767) );
  XOR2_X1 U11796 ( .A(n11768), .B(n11769), .Z(n11652) );
  NAND2_X1 U11797 ( .A1(n11770), .A2(n11771), .ZN(n11768) );
  NOR2_X1 U11798 ( .A1(n11654), .A2(n11655), .ZN(n11764) );
  NOR2_X1 U11799 ( .A1(n11356), .A2(n8376), .ZN(n11655) );
  NAND2_X1 U11800 ( .A1(n11772), .A2(n11773), .ZN(n11654) );
  NAND2_X1 U11801 ( .A1(n11651), .A2(n11774), .ZN(n11773) );
  NAND2_X1 U11802 ( .A1(n11650), .A2(n11649), .ZN(n11774) );
  NOR2_X1 U11803 ( .A1(n11356), .A2(n8371), .ZN(n11651) );
  INV_X1 U11804 ( .A(n11775), .ZN(n11772) );
  NOR2_X1 U11805 ( .A1(n11649), .A2(n11650), .ZN(n11775) );
  NOR2_X1 U11806 ( .A1(n11776), .A2(n11777), .ZN(n11650) );
  INV_X1 U11807 ( .A(n11778), .ZN(n11777) );
  NAND2_X1 U11808 ( .A1(n11548), .A2(n11779), .ZN(n11778) );
  NAND2_X1 U11809 ( .A1(n11545), .A2(n11547), .ZN(n11779) );
  NOR2_X1 U11810 ( .A1(n11356), .A2(n9291), .ZN(n11548) );
  NOR2_X1 U11811 ( .A1(n11547), .A2(n11545), .ZN(n11776) );
  XNOR2_X1 U11812 ( .A(n11780), .B(n11781), .ZN(n11545) );
  XNOR2_X1 U11813 ( .A(n11782), .B(n11783), .ZN(n11781) );
  NAND2_X1 U11814 ( .A1(b_18_), .A2(a_19_), .ZN(n11783) );
  NAND2_X1 U11815 ( .A1(n11784), .A2(n11785), .ZN(n11547) );
  NAND2_X1 U11816 ( .A1(n11553), .A2(n11786), .ZN(n11785) );
  NAND2_X1 U11817 ( .A1(n11555), .A2(n11787), .ZN(n11786) );
  XOR2_X1 U11818 ( .A(n11788), .B(n11789), .Z(n11553) );
  XNOR2_X1 U11819 ( .A(n11790), .B(n11791), .ZN(n11788) );
  NOR2_X1 U11820 ( .A1(n9047), .A2(n11623), .ZN(n11791) );
  NAND2_X1 U11821 ( .A1(n11556), .A2(n11792), .ZN(n11784) );
  INV_X1 U11822 ( .A(n11555), .ZN(n11792) );
  NOR2_X1 U11823 ( .A1(n11793), .A2(n11794), .ZN(n11555) );
  INV_X1 U11824 ( .A(n11795), .ZN(n11794) );
  NAND2_X1 U11825 ( .A1(n11645), .A2(n11796), .ZN(n11795) );
  NAND2_X1 U11826 ( .A1(n11647), .A2(n11646), .ZN(n11796) );
  XNOR2_X1 U11827 ( .A(n11797), .B(n11798), .ZN(n11645) );
  XOR2_X1 U11828 ( .A(n11799), .B(n11800), .Z(n11797) );
  NOR2_X1 U11829 ( .A1(n8759), .A2(n11623), .ZN(n11800) );
  NOR2_X1 U11830 ( .A1(n11646), .A2(n11647), .ZN(n11793) );
  NOR2_X1 U11831 ( .A1(n11356), .A2(n9047), .ZN(n11647) );
  NAND2_X1 U11832 ( .A1(n11801), .A2(n11802), .ZN(n11646) );
  NAND3_X1 U11833 ( .A1(a_21_), .A2(n11803), .A3(b_19_), .ZN(n11802) );
  INV_X1 U11834 ( .A(n11804), .ZN(n11803) );
  NOR2_X1 U11835 ( .A1(n11642), .A2(n11640), .ZN(n11804) );
  NAND2_X1 U11836 ( .A1(n11640), .A2(n11642), .ZN(n11801) );
  NAND2_X1 U11837 ( .A1(n11638), .A2(n11805), .ZN(n11642) );
  NAND2_X1 U11838 ( .A1(n11637), .A2(n11639), .ZN(n11805) );
  NAND2_X1 U11839 ( .A1(n11806), .A2(n11807), .ZN(n11639) );
  NAND2_X1 U11840 ( .A1(b_19_), .A2(a_22_), .ZN(n11807) );
  INV_X1 U11841 ( .A(n11808), .ZN(n11806) );
  XNOR2_X1 U11842 ( .A(n11809), .B(n11810), .ZN(n11637) );
  NAND2_X1 U11843 ( .A1(n11811), .A2(n11812), .ZN(n11809) );
  NAND2_X1 U11844 ( .A1(a_22_), .A2(n11808), .ZN(n11638) );
  NAND2_X1 U11845 ( .A1(n11575), .A2(n11813), .ZN(n11808) );
  NAND2_X1 U11846 ( .A1(n11574), .A2(n11576), .ZN(n11813) );
  NAND2_X1 U11847 ( .A1(n11814), .A2(n11815), .ZN(n11576) );
  NAND2_X1 U11848 ( .A1(b_19_), .A2(a_23_), .ZN(n11815) );
  INV_X1 U11849 ( .A(n11816), .ZN(n11814) );
  XOR2_X1 U11850 ( .A(n11817), .B(n11818), .Z(n11574) );
  XOR2_X1 U11851 ( .A(n11819), .B(n11820), .Z(n11817) );
  NAND2_X1 U11852 ( .A1(a_23_), .A2(n11816), .ZN(n11575) );
  NAND2_X1 U11853 ( .A1(n11821), .A2(n11822), .ZN(n11816) );
  NAND2_X1 U11854 ( .A1(n11584), .A2(n11823), .ZN(n11822) );
  INV_X1 U11855 ( .A(n11824), .ZN(n11823) );
  NOR2_X1 U11856 ( .A1(n11583), .A2(n11582), .ZN(n11824) );
  NOR2_X1 U11857 ( .A1(n11356), .A2(n8779), .ZN(n11584) );
  NAND2_X1 U11858 ( .A1(n11582), .A2(n11583), .ZN(n11821) );
  NAND2_X1 U11859 ( .A1(n11825), .A2(n11826), .ZN(n11583) );
  NAND2_X1 U11860 ( .A1(n11635), .A2(n11827), .ZN(n11826) );
  NAND2_X1 U11861 ( .A1(n11632), .A2(n11634), .ZN(n11827) );
  NOR2_X1 U11862 ( .A1(n11356), .A2(n8788), .ZN(n11635) );
  INV_X1 U11863 ( .A(n11828), .ZN(n11825) );
  NOR2_X1 U11864 ( .A1(n11634), .A2(n11632), .ZN(n11828) );
  XNOR2_X1 U11865 ( .A(n11829), .B(n11830), .ZN(n11632) );
  XNOR2_X1 U11866 ( .A(n11831), .B(n11832), .ZN(n11830) );
  NAND2_X1 U11867 ( .A1(n11833), .A2(n11834), .ZN(n11634) );
  NAND2_X1 U11868 ( .A1(n11593), .A2(n11835), .ZN(n11834) );
  NAND2_X1 U11869 ( .A1(n11596), .A2(n11595), .ZN(n11835) );
  XNOR2_X1 U11870 ( .A(n11836), .B(n11837), .ZN(n11593) );
  XOR2_X1 U11871 ( .A(n11838), .B(n11839), .Z(n11836) );
  INV_X1 U11872 ( .A(n11840), .ZN(n11833) );
  NOR2_X1 U11873 ( .A1(n11595), .A2(n11596), .ZN(n11840) );
  NOR2_X1 U11874 ( .A1(n11356), .A2(n9344), .ZN(n11596) );
  NAND2_X1 U11875 ( .A1(n11841), .A2(n11842), .ZN(n11595) );
  NAND2_X1 U11876 ( .A1(n11603), .A2(n11843), .ZN(n11842) );
  INV_X1 U11877 ( .A(n11844), .ZN(n11843) );
  NOR2_X1 U11878 ( .A1(n11602), .A2(n11601), .ZN(n11844) );
  NOR2_X1 U11879 ( .A1(n11356), .A2(n8797), .ZN(n11603) );
  NAND2_X1 U11880 ( .A1(n11601), .A2(n11602), .ZN(n11841) );
  NAND2_X1 U11881 ( .A1(n11845), .A2(n11846), .ZN(n11602) );
  NAND2_X1 U11882 ( .A1(n11630), .A2(n11847), .ZN(n11846) );
  INV_X1 U11883 ( .A(n11848), .ZN(n11847) );
  NOR2_X1 U11884 ( .A1(n11631), .A2(n11629), .ZN(n11848) );
  NOR2_X1 U11885 ( .A1(n11356), .A2(n8314), .ZN(n11630) );
  NAND2_X1 U11886 ( .A1(n11629), .A2(n11631), .ZN(n11845) );
  NAND2_X1 U11887 ( .A1(n11849), .A2(n11850), .ZN(n11631) );
  NAND2_X1 U11888 ( .A1(n11625), .A2(n11851), .ZN(n11850) );
  INV_X1 U11889 ( .A(n11852), .ZN(n11851) );
  NOR2_X1 U11890 ( .A1(n11626), .A2(n11627), .ZN(n11852) );
  NOR2_X1 U11891 ( .A1(n11356), .A2(n9098), .ZN(n11625) );
  NAND2_X1 U11892 ( .A1(n11627), .A2(n11626), .ZN(n11849) );
  NAND2_X1 U11893 ( .A1(n11853), .A2(n11854), .ZN(n11626) );
  NAND2_X1 U11894 ( .A1(b_17_), .A2(n11855), .ZN(n11854) );
  NAND2_X1 U11895 ( .A1(n8299), .A2(n11856), .ZN(n11855) );
  NAND2_X1 U11896 ( .A1(a_31_), .A2(n11623), .ZN(n11856) );
  NAND2_X1 U11897 ( .A1(b_18_), .A2(n11857), .ZN(n11853) );
  NAND2_X1 U11898 ( .A1(n8303), .A2(n11858), .ZN(n11857) );
  NAND2_X1 U11899 ( .A1(a_30_), .A2(n11859), .ZN(n11858) );
  NOR3_X1 U11900 ( .A1(n11356), .A2(n9631), .A3(n11623), .ZN(n11627) );
  XOR2_X1 U11901 ( .A(n11860), .B(n11861), .Z(n11629) );
  XOR2_X1 U11902 ( .A(n11862), .B(n11863), .Z(n11860) );
  XOR2_X1 U11903 ( .A(n11864), .B(n11865), .Z(n11601) );
  XOR2_X1 U11904 ( .A(n11866), .B(n11867), .Z(n11864) );
  XNOR2_X1 U11905 ( .A(n11868), .B(n11869), .ZN(n11582) );
  XNOR2_X1 U11906 ( .A(n11870), .B(n11871), .ZN(n11869) );
  XNOR2_X1 U11907 ( .A(n11872), .B(n11873), .ZN(n11640) );
  NAND2_X1 U11908 ( .A1(n11874), .A2(n11875), .ZN(n11872) );
  XOR2_X1 U11909 ( .A(n11876), .B(n11877), .Z(n11649) );
  XNOR2_X1 U11910 ( .A(n11878), .B(n11879), .ZN(n11876) );
  XNOR2_X1 U11911 ( .A(n11880), .B(n11881), .ZN(n11521) );
  XOR2_X1 U11912 ( .A(n11882), .B(n11883), .Z(n11881) );
  NAND2_X1 U11913 ( .A1(b_18_), .A2(a_15_), .ZN(n11883) );
  XOR2_X1 U11914 ( .A(n11884), .B(n11885), .Z(n11512) );
  XOR2_X1 U11915 ( .A(n11886), .B(n11887), .Z(n11884) );
  XNOR2_X1 U11916 ( .A(n11888), .B(n11889), .ZN(n11489) );
  XOR2_X1 U11917 ( .A(n11890), .B(n11891), .Z(n11889) );
  XNOR2_X1 U11918 ( .A(n11892), .B(n11893), .ZN(n11656) );
  XOR2_X1 U11919 ( .A(n11894), .B(n11895), .Z(n11892) );
  XNOR2_X1 U11920 ( .A(n11896), .B(n11897), .ZN(n11660) );
  XOR2_X1 U11921 ( .A(n11898), .B(n11899), .Z(n11896) );
  NOR2_X1 U11922 ( .A1(n8971), .A2(n11623), .ZN(n11899) );
  XNOR2_X1 U11923 ( .A(n11900), .B(n11901), .ZN(n11472) );
  NAND2_X1 U11924 ( .A1(n11902), .A2(n11903), .ZN(n11900) );
  XNOR2_X1 U11925 ( .A(n11904), .B(n11905), .ZN(n11465) );
  NAND2_X1 U11926 ( .A1(n11906), .A2(n11907), .ZN(n11904) );
  XNOR2_X1 U11927 ( .A(n11908), .B(n11909), .ZN(n11456) );
  NAND2_X1 U11928 ( .A1(n11910), .A2(n11911), .ZN(n11908) );
  XOR2_X1 U11929 ( .A(n11912), .B(n11913), .Z(n11665) );
  XNOR2_X1 U11930 ( .A(n11914), .B(n11915), .ZN(n11913) );
  XOR2_X1 U11931 ( .A(n11916), .B(n11917), .Z(n11668) );
  XOR2_X1 U11932 ( .A(n11918), .B(n11919), .Z(n11916) );
  XNOR2_X1 U11933 ( .A(n11920), .B(n11921), .ZN(n11672) );
  XNOR2_X1 U11934 ( .A(n11922), .B(n11923), .ZN(n11920) );
  XNOR2_X1 U11935 ( .A(n11924), .B(n11925), .ZN(n11436) );
  XNOR2_X1 U11936 ( .A(n11926), .B(n11927), .ZN(n11924) );
  NOR2_X1 U11937 ( .A1(n8448), .A2(n11623), .ZN(n11927) );
  NAND3_X1 U11938 ( .A1(n8527), .A2(n8526), .A3(n8523), .ZN(n8522) );
  NOR2_X1 U11939 ( .A1(n8596), .A2(n11928), .ZN(n8523) );
  INV_X1 U11940 ( .A(n11929), .ZN(n11928) );
  NAND2_X1 U11941 ( .A1(n11930), .A2(n11931), .ZN(n11929) );
  NAND2_X1 U11942 ( .A1(n11678), .A2(n11932), .ZN(n8526) );
  NAND2_X1 U11943 ( .A1(n11677), .A2(n11679), .ZN(n11932) );
  NAND2_X1 U11944 ( .A1(n11933), .A2(n11934), .ZN(n11679) );
  NAND2_X1 U11945 ( .A1(b_18_), .A2(a_0_), .ZN(n11934) );
  INV_X1 U11946 ( .A(n11935), .ZN(n11933) );
  XNOR2_X1 U11947 ( .A(n11936), .B(n11937), .ZN(n11677) );
  XOR2_X1 U11948 ( .A(n11938), .B(n11939), .Z(n11936) );
  NAND2_X1 U11949 ( .A1(a_0_), .A2(n11935), .ZN(n11678) );
  NAND2_X1 U11950 ( .A1(n11689), .A2(n11940), .ZN(n11935) );
  NAND2_X1 U11951 ( .A1(n11688), .A2(n11690), .ZN(n11940) );
  NAND2_X1 U11952 ( .A1(n11941), .A2(n11942), .ZN(n11690) );
  NAND2_X1 U11953 ( .A1(b_18_), .A2(a_1_), .ZN(n11942) );
  XNOR2_X1 U11954 ( .A(n11943), .B(n11944), .ZN(n11688) );
  XOR2_X1 U11955 ( .A(n11945), .B(n11946), .Z(n11944) );
  NAND2_X1 U11956 ( .A1(b_17_), .A2(a_2_), .ZN(n11946) );
  NAND2_X1 U11957 ( .A1(a_1_), .A2(n11947), .ZN(n11689) );
  INV_X1 U11958 ( .A(n11941), .ZN(n11947) );
  NOR2_X1 U11959 ( .A1(n11948), .A2(n11949), .ZN(n11941) );
  NOR3_X1 U11960 ( .A1(n8448), .A2(n11950), .A3(n11623), .ZN(n11949) );
  INV_X1 U11961 ( .A(n11951), .ZN(n11950) );
  NAND2_X1 U11962 ( .A1(n11925), .A2(n11926), .ZN(n11951) );
  NOR2_X1 U11963 ( .A1(n11925), .A2(n11926), .ZN(n11948) );
  NOR2_X1 U11964 ( .A1(n11952), .A2(n11953), .ZN(n11926) );
  INV_X1 U11965 ( .A(n11954), .ZN(n11953) );
  NAND2_X1 U11966 ( .A1(n11923), .A2(n11955), .ZN(n11954) );
  NAND2_X1 U11967 ( .A1(n11922), .A2(n11921), .ZN(n11955) );
  NOR2_X1 U11968 ( .A1(n11623), .A2(n8900), .ZN(n11923) );
  NOR2_X1 U11969 ( .A1(n11921), .A2(n11922), .ZN(n11952) );
  NOR2_X1 U11970 ( .A1(n11956), .A2(n11957), .ZN(n11922) );
  INV_X1 U11971 ( .A(n11958), .ZN(n11957) );
  NAND2_X1 U11972 ( .A1(n11919), .A2(n11959), .ZN(n11958) );
  NAND2_X1 U11973 ( .A1(n11917), .A2(n11918), .ZN(n11959) );
  NOR2_X1 U11974 ( .A1(n11623), .A2(n8439), .ZN(n11919) );
  NOR2_X1 U11975 ( .A1(n11917), .A2(n11918), .ZN(n11956) );
  NAND2_X1 U11976 ( .A1(n11960), .A2(n11961), .ZN(n11918) );
  NAND2_X1 U11977 ( .A1(n11912), .A2(n11962), .ZN(n11961) );
  NAND2_X1 U11978 ( .A1(n11915), .A2(n11914), .ZN(n11962) );
  XNOR2_X1 U11979 ( .A(n11963), .B(n11964), .ZN(n11912) );
  XOR2_X1 U11980 ( .A(n11965), .B(n11966), .Z(n11963) );
  NOR2_X1 U11981 ( .A1(n8430), .A2(n11859), .ZN(n11966) );
  INV_X1 U11982 ( .A(n11967), .ZN(n11960) );
  NOR2_X1 U11983 ( .A1(n11914), .A2(n11915), .ZN(n11967) );
  NOR2_X1 U11984 ( .A1(n11623), .A2(n8938), .ZN(n11915) );
  NAND2_X1 U11985 ( .A1(n11910), .A2(n11968), .ZN(n11914) );
  NAND2_X1 U11986 ( .A1(n11909), .A2(n11911), .ZN(n11968) );
  NAND2_X1 U11987 ( .A1(n11969), .A2(n11970), .ZN(n11911) );
  NAND2_X1 U11988 ( .A1(b_18_), .A2(a_6_), .ZN(n11970) );
  INV_X1 U11989 ( .A(n11971), .ZN(n11969) );
  XOR2_X1 U11990 ( .A(n11972), .B(n11973), .Z(n11909) );
  XNOR2_X1 U11991 ( .A(n11974), .B(n11975), .ZN(n11973) );
  NAND2_X1 U11992 ( .A1(b_17_), .A2(a_7_), .ZN(n11975) );
  NAND2_X1 U11993 ( .A1(a_6_), .A2(n11971), .ZN(n11910) );
  NAND2_X1 U11994 ( .A1(n11906), .A2(n11976), .ZN(n11971) );
  NAND2_X1 U11995 ( .A1(n11905), .A2(n11907), .ZN(n11976) );
  NAND2_X1 U11996 ( .A1(n11977), .A2(n11978), .ZN(n11907) );
  NAND2_X1 U11997 ( .A1(b_18_), .A2(a_7_), .ZN(n11978) );
  INV_X1 U11998 ( .A(n11979), .ZN(n11977) );
  XNOR2_X1 U11999 ( .A(n11980), .B(n11981), .ZN(n11905) );
  XNOR2_X1 U12000 ( .A(n11982), .B(n11983), .ZN(n11980) );
  NOR2_X1 U12001 ( .A1(n8968), .A2(n11859), .ZN(n11983) );
  NAND2_X1 U12002 ( .A1(a_7_), .A2(n11979), .ZN(n11906) );
  NAND2_X1 U12003 ( .A1(n11902), .A2(n11984), .ZN(n11979) );
  NAND2_X1 U12004 ( .A1(n11901), .A2(n11903), .ZN(n11984) );
  NAND2_X1 U12005 ( .A1(n11985), .A2(n11986), .ZN(n11903) );
  NAND2_X1 U12006 ( .A1(b_18_), .A2(a_8_), .ZN(n11986) );
  INV_X1 U12007 ( .A(n11987), .ZN(n11985) );
  XNOR2_X1 U12008 ( .A(n11988), .B(n11989), .ZN(n11901) );
  XNOR2_X1 U12009 ( .A(n11990), .B(n11991), .ZN(n11988) );
  NOR2_X1 U12010 ( .A1(n8971), .A2(n11859), .ZN(n11991) );
  NAND2_X1 U12011 ( .A1(a_8_), .A2(n11987), .ZN(n11902) );
  NAND2_X1 U12012 ( .A1(n11992), .A2(n11993), .ZN(n11987) );
  INV_X1 U12013 ( .A(n11994), .ZN(n11993) );
  NOR3_X1 U12014 ( .A1(n8971), .A2(n11995), .A3(n11623), .ZN(n11994) );
  NOR2_X1 U12015 ( .A1(n11897), .A2(n11898), .ZN(n11995) );
  NAND2_X1 U12016 ( .A1(n11897), .A2(n11898), .ZN(n11992) );
  NAND2_X1 U12017 ( .A1(n11996), .A2(n11997), .ZN(n11898) );
  NAND2_X1 U12018 ( .A1(n11895), .A2(n11998), .ZN(n11997) );
  INV_X1 U12019 ( .A(n11999), .ZN(n11998) );
  NOR2_X1 U12020 ( .A1(n11894), .A2(n11893), .ZN(n11999) );
  NOR2_X1 U12021 ( .A1(n11623), .A2(n8402), .ZN(n11895) );
  NAND2_X1 U12022 ( .A1(n11893), .A2(n11894), .ZN(n11996) );
  NAND2_X1 U12023 ( .A1(n12000), .A2(n12001), .ZN(n11894) );
  NAND2_X1 U12024 ( .A1(n11891), .A2(n12002), .ZN(n12001) );
  NAND2_X1 U12025 ( .A1(n11888), .A2(n11890), .ZN(n12002) );
  NOR2_X1 U12026 ( .A1(n11623), .A2(n8867), .ZN(n11891) );
  INV_X1 U12027 ( .A(n12003), .ZN(n12000) );
  NOR2_X1 U12028 ( .A1(n11888), .A2(n11890), .ZN(n12003) );
  NOR2_X1 U12029 ( .A1(n12004), .A2(n12005), .ZN(n11890) );
  INV_X1 U12030 ( .A(n12006), .ZN(n12005) );
  NAND3_X1 U12031 ( .A1(a_12_), .A2(n12007), .A3(b_18_), .ZN(n12006) );
  NAND2_X1 U12032 ( .A1(n11738), .A2(n11737), .ZN(n12007) );
  NOR2_X1 U12033 ( .A1(n11737), .A2(n11738), .ZN(n12004) );
  NOR2_X1 U12034 ( .A1(n12008), .A2(n12009), .ZN(n11738) );
  NOR3_X1 U12035 ( .A1(n8996), .A2(n12010), .A3(n11623), .ZN(n12009) );
  NOR2_X1 U12036 ( .A1(n11744), .A2(n11745), .ZN(n12010) );
  INV_X1 U12037 ( .A(n12011), .ZN(n12008) );
  NAND2_X1 U12038 ( .A1(n11745), .A2(n11744), .ZN(n12011) );
  XNOR2_X1 U12039 ( .A(n12012), .B(n12013), .ZN(n11744) );
  XNOR2_X1 U12040 ( .A(n12014), .B(n12015), .ZN(n12013) );
  NOR2_X1 U12041 ( .A1(n12016), .A2(n12017), .ZN(n11745) );
  INV_X1 U12042 ( .A(n12018), .ZN(n12017) );
  NAND2_X1 U12043 ( .A1(n11885), .A2(n12019), .ZN(n12018) );
  NAND2_X1 U12044 ( .A1(n11887), .A2(n11886), .ZN(n12019) );
  XOR2_X1 U12045 ( .A(n12020), .B(n12021), .Z(n11885) );
  XOR2_X1 U12046 ( .A(n12022), .B(n12023), .Z(n12021) );
  NAND2_X1 U12047 ( .A1(b_17_), .A2(a_15_), .ZN(n12023) );
  NOR2_X1 U12048 ( .A1(n11886), .A2(n11887), .ZN(n12016) );
  NOR2_X1 U12049 ( .A1(n11623), .A2(n9262), .ZN(n11887) );
  NAND2_X1 U12050 ( .A1(n12024), .A2(n12025), .ZN(n11886) );
  INV_X1 U12051 ( .A(n12026), .ZN(n12025) );
  NOR3_X1 U12052 ( .A1(n8850), .A2(n12027), .A3(n11623), .ZN(n12026) );
  NOR2_X1 U12053 ( .A1(n11882), .A2(n11880), .ZN(n12027) );
  NAND2_X1 U12054 ( .A1(n11880), .A2(n11882), .ZN(n12024) );
  NAND2_X1 U12055 ( .A1(n12028), .A2(n12029), .ZN(n11882) );
  NAND3_X1 U12056 ( .A1(a_16_), .A2(n12030), .A3(b_18_), .ZN(n12029) );
  INV_X1 U12057 ( .A(n12031), .ZN(n12030) );
  NOR2_X1 U12058 ( .A1(n11760), .A2(n11762), .ZN(n12031) );
  NAND2_X1 U12059 ( .A1(n11760), .A2(n11762), .ZN(n12028) );
  NAND2_X1 U12060 ( .A1(n11770), .A2(n12032), .ZN(n11762) );
  NAND2_X1 U12061 ( .A1(n11769), .A2(n11771), .ZN(n12032) );
  NAND2_X1 U12062 ( .A1(n12033), .A2(n12034), .ZN(n11771) );
  NAND2_X1 U12063 ( .A1(b_18_), .A2(a_17_), .ZN(n12034) );
  XNOR2_X1 U12064 ( .A(n12035), .B(n12036), .ZN(n11769) );
  XOR2_X1 U12065 ( .A(n12037), .B(n12038), .Z(n12036) );
  NAND2_X1 U12066 ( .A1(b_17_), .A2(a_18_), .ZN(n12038) );
  NAND2_X1 U12067 ( .A1(a_17_), .A2(n12039), .ZN(n11770) );
  INV_X1 U12068 ( .A(n12033), .ZN(n12039) );
  NOR2_X1 U12069 ( .A1(n12040), .A2(n12041), .ZN(n12033) );
  INV_X1 U12070 ( .A(n12042), .ZN(n12041) );
  NAND2_X1 U12071 ( .A1(n11879), .A2(n12043), .ZN(n12042) );
  NAND2_X1 U12072 ( .A1(n11878), .A2(n11877), .ZN(n12043) );
  NOR2_X1 U12073 ( .A1(n11877), .A2(n11878), .ZN(n12040) );
  NOR2_X1 U12074 ( .A1(n12044), .A2(n12045), .ZN(n11878) );
  NOR3_X1 U12075 ( .A1(n8742), .A2(n12046), .A3(n11623), .ZN(n12045) );
  INV_X1 U12076 ( .A(n12047), .ZN(n12046) );
  NAND2_X1 U12077 ( .A1(n11782), .A2(n11780), .ZN(n12047) );
  NOR2_X1 U12078 ( .A1(n11780), .A2(n11782), .ZN(n12044) );
  NOR2_X1 U12079 ( .A1(n12048), .A2(n12049), .ZN(n11782) );
  INV_X1 U12080 ( .A(n12050), .ZN(n12049) );
  NAND3_X1 U12081 ( .A1(a_20_), .A2(n12051), .A3(b_18_), .ZN(n12050) );
  NAND2_X1 U12082 ( .A1(n11790), .A2(n11789), .ZN(n12051) );
  NOR2_X1 U12083 ( .A1(n11789), .A2(n11790), .ZN(n12048) );
  NOR2_X1 U12084 ( .A1(n12052), .A2(n12053), .ZN(n11790) );
  NOR3_X1 U12085 ( .A1(n8759), .A2(n12054), .A3(n11623), .ZN(n12053) );
  NOR2_X1 U12086 ( .A1(n11798), .A2(n11799), .ZN(n12054) );
  INV_X1 U12087 ( .A(n12055), .ZN(n12052) );
  NAND2_X1 U12088 ( .A1(n11798), .A2(n11799), .ZN(n12055) );
  NAND2_X1 U12089 ( .A1(n11874), .A2(n12056), .ZN(n11799) );
  NAND2_X1 U12090 ( .A1(n11873), .A2(n11875), .ZN(n12056) );
  NAND2_X1 U12091 ( .A1(n12057), .A2(n12058), .ZN(n11875) );
  NAND2_X1 U12092 ( .A1(b_18_), .A2(a_22_), .ZN(n12058) );
  INV_X1 U12093 ( .A(n12059), .ZN(n12057) );
  XOR2_X1 U12094 ( .A(n12060), .B(n12061), .Z(n11873) );
  XOR2_X1 U12095 ( .A(n12062), .B(n12063), .Z(n12060) );
  NAND2_X1 U12096 ( .A1(a_22_), .A2(n12059), .ZN(n11874) );
  NAND2_X1 U12097 ( .A1(n11811), .A2(n12064), .ZN(n12059) );
  NAND2_X1 U12098 ( .A1(n11810), .A2(n11812), .ZN(n12064) );
  NAND2_X1 U12099 ( .A1(n12065), .A2(n12066), .ZN(n11812) );
  NAND2_X1 U12100 ( .A1(b_18_), .A2(a_23_), .ZN(n12066) );
  INV_X1 U12101 ( .A(n12067), .ZN(n12065) );
  XOR2_X1 U12102 ( .A(n12068), .B(n12069), .Z(n11810) );
  XOR2_X1 U12103 ( .A(n12070), .B(n12071), .Z(n12068) );
  NAND2_X1 U12104 ( .A1(a_23_), .A2(n12067), .ZN(n11811) );
  NAND2_X1 U12105 ( .A1(n12072), .A2(n12073), .ZN(n12067) );
  NAND2_X1 U12106 ( .A1(n11820), .A2(n12074), .ZN(n12073) );
  INV_X1 U12107 ( .A(n12075), .ZN(n12074) );
  NOR2_X1 U12108 ( .A1(n11818), .A2(n11819), .ZN(n12075) );
  NOR2_X1 U12109 ( .A1(n11623), .A2(n8779), .ZN(n11820) );
  NAND2_X1 U12110 ( .A1(n11818), .A2(n11819), .ZN(n12072) );
  NAND2_X1 U12111 ( .A1(n12076), .A2(n12077), .ZN(n11819) );
  NAND2_X1 U12112 ( .A1(n11871), .A2(n12078), .ZN(n12077) );
  NAND2_X1 U12113 ( .A1(n11868), .A2(n11870), .ZN(n12078) );
  NOR2_X1 U12114 ( .A1(n11623), .A2(n8788), .ZN(n11871) );
  INV_X1 U12115 ( .A(n12079), .ZN(n12076) );
  NOR2_X1 U12116 ( .A1(n11870), .A2(n11868), .ZN(n12079) );
  XNOR2_X1 U12117 ( .A(n12080), .B(n12081), .ZN(n11868) );
  XNOR2_X1 U12118 ( .A(n12082), .B(n12083), .ZN(n12081) );
  NAND2_X1 U12119 ( .A1(n12084), .A2(n12085), .ZN(n11870) );
  NAND2_X1 U12120 ( .A1(n11829), .A2(n12086), .ZN(n12085) );
  NAND2_X1 U12121 ( .A1(n11832), .A2(n11831), .ZN(n12086) );
  XNOR2_X1 U12122 ( .A(n12087), .B(n12088), .ZN(n11829) );
  XOR2_X1 U12123 ( .A(n12089), .B(n12090), .Z(n12087) );
  INV_X1 U12124 ( .A(n12091), .ZN(n12084) );
  NOR2_X1 U12125 ( .A1(n11831), .A2(n11832), .ZN(n12091) );
  NOR2_X1 U12126 ( .A1(n11623), .A2(n9344), .ZN(n11832) );
  NAND2_X1 U12127 ( .A1(n12092), .A2(n12093), .ZN(n11831) );
  NAND2_X1 U12128 ( .A1(n11839), .A2(n12094), .ZN(n12093) );
  INV_X1 U12129 ( .A(n12095), .ZN(n12094) );
  NOR2_X1 U12130 ( .A1(n11837), .A2(n11838), .ZN(n12095) );
  NOR2_X1 U12131 ( .A1(n11623), .A2(n8797), .ZN(n11839) );
  NAND2_X1 U12132 ( .A1(n11837), .A2(n11838), .ZN(n12092) );
  NAND2_X1 U12133 ( .A1(n12096), .A2(n12097), .ZN(n11838) );
  NAND2_X1 U12134 ( .A1(n11866), .A2(n12098), .ZN(n12097) );
  INV_X1 U12135 ( .A(n12099), .ZN(n12098) );
  NOR2_X1 U12136 ( .A1(n11867), .A2(n11865), .ZN(n12099) );
  NOR2_X1 U12137 ( .A1(n11623), .A2(n8314), .ZN(n11866) );
  NAND2_X1 U12138 ( .A1(n11865), .A2(n11867), .ZN(n12096) );
  NAND2_X1 U12139 ( .A1(n12100), .A2(n12101), .ZN(n11867) );
  NAND2_X1 U12140 ( .A1(n11861), .A2(n12102), .ZN(n12101) );
  INV_X1 U12141 ( .A(n12103), .ZN(n12102) );
  NOR2_X1 U12142 ( .A1(n11862), .A2(n11863), .ZN(n12103) );
  NOR2_X1 U12143 ( .A1(n11623), .A2(n9098), .ZN(n11861) );
  NAND2_X1 U12144 ( .A1(n11863), .A2(n11862), .ZN(n12100) );
  NAND2_X1 U12145 ( .A1(n12104), .A2(n12105), .ZN(n11862) );
  NAND2_X1 U12146 ( .A1(b_16_), .A2(n12106), .ZN(n12105) );
  NAND2_X1 U12147 ( .A1(n8299), .A2(n12107), .ZN(n12106) );
  NAND2_X1 U12148 ( .A1(a_31_), .A2(n11859), .ZN(n12107) );
  NAND2_X1 U12149 ( .A1(b_17_), .A2(n12108), .ZN(n12104) );
  NAND2_X1 U12150 ( .A1(n8303), .A2(n12109), .ZN(n12108) );
  NAND2_X1 U12151 ( .A1(a_30_), .A2(n12110), .ZN(n12109) );
  NOR3_X1 U12152 ( .A1(n11859), .A2(n9631), .A3(n11623), .ZN(n11863) );
  XOR2_X1 U12153 ( .A(n12111), .B(n12112), .Z(n11865) );
  XOR2_X1 U12154 ( .A(n12113), .B(n12114), .Z(n12111) );
  XOR2_X1 U12155 ( .A(n12115), .B(n12116), .Z(n11837) );
  XOR2_X1 U12156 ( .A(n12117), .B(n12118), .Z(n12115) );
  XNOR2_X1 U12157 ( .A(n12119), .B(n12120), .ZN(n11818) );
  XNOR2_X1 U12158 ( .A(n12121), .B(n12122), .ZN(n12120) );
  XNOR2_X1 U12159 ( .A(n12123), .B(n12124), .ZN(n11798) );
  XNOR2_X1 U12160 ( .A(n12125), .B(n12126), .ZN(n12124) );
  XOR2_X1 U12161 ( .A(n12127), .B(n12128), .Z(n11789) );
  XOR2_X1 U12162 ( .A(n12129), .B(n12130), .Z(n12128) );
  XOR2_X1 U12163 ( .A(n12131), .B(n12132), .Z(n11780) );
  XOR2_X1 U12164 ( .A(n12133), .B(n12134), .Z(n12131) );
  XOR2_X1 U12165 ( .A(n12135), .B(n12136), .Z(n11877) );
  XOR2_X1 U12166 ( .A(n12137), .B(n12138), .Z(n12136) );
  NAND2_X1 U12167 ( .A1(b_17_), .A2(a_19_), .ZN(n12138) );
  XNOR2_X1 U12168 ( .A(n12139), .B(n12140), .ZN(n11760) );
  XOR2_X1 U12169 ( .A(n12141), .B(n12142), .Z(n12139) );
  XNOR2_X1 U12170 ( .A(n12143), .B(n12144), .ZN(n11880) );
  NAND2_X1 U12171 ( .A1(n12145), .A2(n12146), .ZN(n12143) );
  XNOR2_X1 U12172 ( .A(n12147), .B(n12148), .ZN(n11737) );
  XOR2_X1 U12173 ( .A(n12149), .B(n12150), .Z(n12147) );
  XNOR2_X1 U12174 ( .A(n12151), .B(n12152), .ZN(n11888) );
  XOR2_X1 U12175 ( .A(n12153), .B(n12154), .Z(n12151) );
  NOR2_X1 U12176 ( .A1(n8393), .A2(n11859), .ZN(n12154) );
  XOR2_X1 U12177 ( .A(n12155), .B(n12156), .Z(n11893) );
  XNOR2_X1 U12178 ( .A(n12157), .B(n12158), .ZN(n12156) );
  NAND2_X1 U12179 ( .A1(b_17_), .A2(a_11_), .ZN(n12158) );
  XOR2_X1 U12180 ( .A(n12159), .B(n12160), .Z(n11897) );
  XNOR2_X1 U12181 ( .A(n12161), .B(n12162), .ZN(n12160) );
  NAND2_X1 U12182 ( .A1(b_17_), .A2(a_10_), .ZN(n12162) );
  XOR2_X1 U12183 ( .A(n12163), .B(n12164), .Z(n11917) );
  XOR2_X1 U12184 ( .A(n12165), .B(n12166), .Z(n12164) );
  NAND2_X1 U12185 ( .A1(b_17_), .A2(a_5_), .ZN(n12166) );
  XNOR2_X1 U12186 ( .A(n12167), .B(n12168), .ZN(n11921) );
  XOR2_X1 U12187 ( .A(n12169), .B(n12170), .Z(n12167) );
  NOR2_X1 U12188 ( .A1(n8439), .A2(n11859), .ZN(n12170) );
  XOR2_X1 U12189 ( .A(n12171), .B(n12172), .Z(n11925) );
  XOR2_X1 U12190 ( .A(n12173), .B(n12174), .Z(n12172) );
  NAND2_X1 U12191 ( .A1(b_17_), .A2(a_3_), .ZN(n12174) );
  XNOR2_X1 U12192 ( .A(n12175), .B(n12176), .ZN(n8527) );
  XNOR2_X1 U12193 ( .A(n12177), .B(n12178), .ZN(n12176) );
  INV_X1 U12194 ( .A(n12179), .ZN(n8531) );
  NOR2_X1 U12195 ( .A1(n8595), .A2(n8596), .ZN(n12179) );
  NOR2_X1 U12196 ( .A1(n11931), .A2(n11930), .ZN(n8596) );
  NOR2_X1 U12197 ( .A1(n12180), .A2(n12181), .ZN(n11930) );
  INV_X1 U12198 ( .A(n12182), .ZN(n12181) );
  NAND2_X1 U12199 ( .A1(n12178), .A2(n12183), .ZN(n12182) );
  NAND2_X1 U12200 ( .A1(n12175), .A2(n12177), .ZN(n12183) );
  NOR2_X1 U12201 ( .A1(n11859), .A2(n8457), .ZN(n12178) );
  NOR2_X1 U12202 ( .A1(n12177), .A2(n12175), .ZN(n12180) );
  XNOR2_X1 U12203 ( .A(n12184), .B(n12185), .ZN(n12175) );
  XOR2_X1 U12204 ( .A(n12186), .B(n12187), .Z(n12184) );
  NOR2_X1 U12205 ( .A1(n8569), .A2(n12110), .ZN(n12187) );
  NAND2_X1 U12206 ( .A1(n12188), .A2(n12189), .ZN(n12177) );
  NAND2_X1 U12207 ( .A1(n11937), .A2(n12190), .ZN(n12189) );
  NAND2_X1 U12208 ( .A1(n11939), .A2(n11938), .ZN(n12190) );
  XNOR2_X1 U12209 ( .A(n12191), .B(n12192), .ZN(n11937) );
  XNOR2_X1 U12210 ( .A(n12193), .B(n12194), .ZN(n12192) );
  INV_X1 U12211 ( .A(n12195), .ZN(n12188) );
  NOR2_X1 U12212 ( .A1(n11938), .A2(n11939), .ZN(n12195) );
  NOR2_X1 U12213 ( .A1(n11859), .A2(n8569), .ZN(n11939) );
  NAND2_X1 U12214 ( .A1(n12196), .A2(n12197), .ZN(n11938) );
  NAND3_X1 U12215 ( .A1(a_2_), .A2(n12198), .A3(b_17_), .ZN(n12197) );
  INV_X1 U12216 ( .A(n12199), .ZN(n12198) );
  NOR2_X1 U12217 ( .A1(n11945), .A2(n11943), .ZN(n12199) );
  NAND2_X1 U12218 ( .A1(n11943), .A2(n11945), .ZN(n12196) );
  NAND2_X1 U12219 ( .A1(n12200), .A2(n12201), .ZN(n11945) );
  INV_X1 U12220 ( .A(n12202), .ZN(n12201) );
  NOR3_X1 U12221 ( .A1(n8900), .A2(n12203), .A3(n11859), .ZN(n12202) );
  NOR2_X1 U12222 ( .A1(n12173), .A2(n12171), .ZN(n12203) );
  NAND2_X1 U12223 ( .A1(n12171), .A2(n12173), .ZN(n12200) );
  NAND2_X1 U12224 ( .A1(n12204), .A2(n12205), .ZN(n12173) );
  NAND3_X1 U12225 ( .A1(a_4_), .A2(n12206), .A3(b_17_), .ZN(n12205) );
  INV_X1 U12226 ( .A(n12207), .ZN(n12206) );
  NOR2_X1 U12227 ( .A1(n12169), .A2(n12168), .ZN(n12207) );
  NAND2_X1 U12228 ( .A1(n12168), .A2(n12169), .ZN(n12204) );
  NAND2_X1 U12229 ( .A1(n12208), .A2(n12209), .ZN(n12169) );
  INV_X1 U12230 ( .A(n12210), .ZN(n12209) );
  NOR3_X1 U12231 ( .A1(n8938), .A2(n12211), .A3(n11859), .ZN(n12210) );
  NOR2_X1 U12232 ( .A1(n12165), .A2(n12163), .ZN(n12211) );
  NAND2_X1 U12233 ( .A1(n12163), .A2(n12165), .ZN(n12208) );
  NAND2_X1 U12234 ( .A1(n12212), .A2(n12213), .ZN(n12165) );
  NAND3_X1 U12235 ( .A1(a_6_), .A2(n12214), .A3(b_17_), .ZN(n12213) );
  INV_X1 U12236 ( .A(n12215), .ZN(n12214) );
  NOR2_X1 U12237 ( .A1(n11965), .A2(n11964), .ZN(n12215) );
  NAND2_X1 U12238 ( .A1(n11964), .A2(n11965), .ZN(n12212) );
  NAND2_X1 U12239 ( .A1(n12216), .A2(n12217), .ZN(n11965) );
  NAND3_X1 U12240 ( .A1(a_7_), .A2(n12218), .A3(b_17_), .ZN(n12217) );
  NAND2_X1 U12241 ( .A1(n11974), .A2(n11972), .ZN(n12218) );
  INV_X1 U12242 ( .A(n12219), .ZN(n12216) );
  NOR2_X1 U12243 ( .A1(n11972), .A2(n11974), .ZN(n12219) );
  NOR2_X1 U12244 ( .A1(n12220), .A2(n12221), .ZN(n11974) );
  INV_X1 U12245 ( .A(n12222), .ZN(n12221) );
  NAND3_X1 U12246 ( .A1(a_8_), .A2(n12223), .A3(b_17_), .ZN(n12222) );
  NAND2_X1 U12247 ( .A1(n11982), .A2(n11981), .ZN(n12223) );
  NOR2_X1 U12248 ( .A1(n11981), .A2(n11982), .ZN(n12220) );
  NOR2_X1 U12249 ( .A1(n12224), .A2(n12225), .ZN(n11982) );
  INV_X1 U12250 ( .A(n12226), .ZN(n12225) );
  NAND3_X1 U12251 ( .A1(a_9_), .A2(n12227), .A3(b_17_), .ZN(n12226) );
  NAND2_X1 U12252 ( .A1(n11990), .A2(n11989), .ZN(n12227) );
  NOR2_X1 U12253 ( .A1(n11989), .A2(n11990), .ZN(n12224) );
  NOR2_X1 U12254 ( .A1(n12228), .A2(n12229), .ZN(n11990) );
  NOR3_X1 U12255 ( .A1(n8402), .A2(n12230), .A3(n11859), .ZN(n12229) );
  INV_X1 U12256 ( .A(n12231), .ZN(n12230) );
  NAND2_X1 U12257 ( .A1(n12161), .A2(n12159), .ZN(n12231) );
  NOR2_X1 U12258 ( .A1(n12159), .A2(n12161), .ZN(n12228) );
  NOR2_X1 U12259 ( .A1(n12232), .A2(n12233), .ZN(n12161) );
  INV_X1 U12260 ( .A(n12234), .ZN(n12233) );
  NAND3_X1 U12261 ( .A1(a_11_), .A2(n12235), .A3(b_17_), .ZN(n12234) );
  NAND2_X1 U12262 ( .A1(n12157), .A2(n12155), .ZN(n12235) );
  NOR2_X1 U12263 ( .A1(n12155), .A2(n12157), .ZN(n12232) );
  NOR2_X1 U12264 ( .A1(n12236), .A2(n12237), .ZN(n12157) );
  NOR3_X1 U12265 ( .A1(n8393), .A2(n12238), .A3(n11859), .ZN(n12237) );
  NOR2_X1 U12266 ( .A1(n12153), .A2(n12152), .ZN(n12238) );
  INV_X1 U12267 ( .A(n12239), .ZN(n12236) );
  NAND2_X1 U12268 ( .A1(n12152), .A2(n12153), .ZN(n12239) );
  NAND2_X1 U12269 ( .A1(n12240), .A2(n12241), .ZN(n12153) );
  NAND2_X1 U12270 ( .A1(n12150), .A2(n12242), .ZN(n12241) );
  INV_X1 U12271 ( .A(n12243), .ZN(n12242) );
  NOR2_X1 U12272 ( .A1(n12149), .A2(n12148), .ZN(n12243) );
  NOR2_X1 U12273 ( .A1(n11859), .A2(n8996), .ZN(n12150) );
  NAND2_X1 U12274 ( .A1(n12148), .A2(n12149), .ZN(n12240) );
  NAND2_X1 U12275 ( .A1(n12244), .A2(n12245), .ZN(n12149) );
  NAND2_X1 U12276 ( .A1(n12015), .A2(n12246), .ZN(n12245) );
  INV_X1 U12277 ( .A(n12247), .ZN(n12246) );
  NOR2_X1 U12278 ( .A1(n12014), .A2(n12012), .ZN(n12247) );
  NOR2_X1 U12279 ( .A1(n11859), .A2(n9262), .ZN(n12015) );
  NAND2_X1 U12280 ( .A1(n12012), .A2(n12014), .ZN(n12244) );
  NAND2_X1 U12281 ( .A1(n12248), .A2(n12249), .ZN(n12014) );
  INV_X1 U12282 ( .A(n12250), .ZN(n12249) );
  NOR3_X1 U12283 ( .A1(n8850), .A2(n12251), .A3(n11859), .ZN(n12250) );
  NOR2_X1 U12284 ( .A1(n12022), .A2(n12020), .ZN(n12251) );
  NAND2_X1 U12285 ( .A1(n12020), .A2(n12022), .ZN(n12248) );
  NAND2_X1 U12286 ( .A1(n12145), .A2(n12252), .ZN(n12022) );
  NAND2_X1 U12287 ( .A1(n12144), .A2(n12146), .ZN(n12252) );
  NAND2_X1 U12288 ( .A1(n12253), .A2(n12254), .ZN(n12146) );
  NAND2_X1 U12289 ( .A1(b_17_), .A2(a_16_), .ZN(n12253) );
  XOR2_X1 U12290 ( .A(n12255), .B(n12256), .Z(n12144) );
  XOR2_X1 U12291 ( .A(n12257), .B(n12258), .Z(n12255) );
  NOR2_X1 U12292 ( .A1(n8371), .A2(n12110), .ZN(n12258) );
  NAND2_X1 U12293 ( .A1(n12259), .A2(a_16_), .ZN(n12145) );
  INV_X1 U12294 ( .A(n12254), .ZN(n12259) );
  NAND2_X1 U12295 ( .A1(n12260), .A2(n12261), .ZN(n12254) );
  NAND2_X1 U12296 ( .A1(n12140), .A2(n12262), .ZN(n12261) );
  INV_X1 U12297 ( .A(n12263), .ZN(n12262) );
  NOR2_X1 U12298 ( .A1(n12142), .A2(n12141), .ZN(n12263) );
  XNOR2_X1 U12299 ( .A(n12264), .B(n12265), .ZN(n12140) );
  XNOR2_X1 U12300 ( .A(n12266), .B(n12267), .ZN(n12265) );
  NAND2_X1 U12301 ( .A1(n12141), .A2(n12142), .ZN(n12260) );
  NOR2_X1 U12302 ( .A1(n12268), .A2(n12269), .ZN(n12141) );
  NOR3_X1 U12303 ( .A1(n9291), .A2(n12270), .A3(n11859), .ZN(n12269) );
  NOR2_X1 U12304 ( .A1(n12037), .A2(n12035), .ZN(n12270) );
  INV_X1 U12305 ( .A(n12271), .ZN(n12268) );
  NAND2_X1 U12306 ( .A1(n12035), .A2(n12037), .ZN(n12271) );
  NAND2_X1 U12307 ( .A1(n12272), .A2(n12273), .ZN(n12037) );
  NAND3_X1 U12308 ( .A1(a_19_), .A2(n12274), .A3(b_17_), .ZN(n12273) );
  NAND2_X1 U12309 ( .A1(n12135), .A2(n12137), .ZN(n12274) );
  INV_X1 U12310 ( .A(n12275), .ZN(n12272) );
  NOR2_X1 U12311 ( .A1(n12137), .A2(n12135), .ZN(n12275) );
  XOR2_X1 U12312 ( .A(n12276), .B(n12277), .Z(n12135) );
  XNOR2_X1 U12313 ( .A(n12278), .B(n12279), .ZN(n12276) );
  NOR2_X1 U12314 ( .A1(n9047), .A2(n12110), .ZN(n12279) );
  NAND2_X1 U12315 ( .A1(n12280), .A2(n12281), .ZN(n12137) );
  NAND2_X1 U12316 ( .A1(n12132), .A2(n12282), .ZN(n12281) );
  NAND2_X1 U12317 ( .A1(n12134), .A2(n12133), .ZN(n12282) );
  XNOR2_X1 U12318 ( .A(n12283), .B(n12284), .ZN(n12132) );
  XOR2_X1 U12319 ( .A(n12285), .B(n12286), .Z(n12283) );
  NOR2_X1 U12320 ( .A1(n8759), .A2(n12110), .ZN(n12286) );
  INV_X1 U12321 ( .A(n12287), .ZN(n12280) );
  NOR2_X1 U12322 ( .A1(n12133), .A2(n12134), .ZN(n12287) );
  NOR2_X1 U12323 ( .A1(n11859), .A2(n9047), .ZN(n12134) );
  NAND2_X1 U12324 ( .A1(n12288), .A2(n12289), .ZN(n12133) );
  INV_X1 U12325 ( .A(n12290), .ZN(n12289) );
  NOR2_X1 U12326 ( .A1(n12130), .A2(n12291), .ZN(n12290) );
  NOR2_X1 U12327 ( .A1(n12129), .A2(n12127), .ZN(n12291) );
  NAND2_X1 U12328 ( .A1(b_17_), .A2(a_21_), .ZN(n12130) );
  NAND2_X1 U12329 ( .A1(n12127), .A2(n12129), .ZN(n12288) );
  NAND2_X1 U12330 ( .A1(n12292), .A2(n12293), .ZN(n12129) );
  NAND2_X1 U12331 ( .A1(n12126), .A2(n12294), .ZN(n12293) );
  INV_X1 U12332 ( .A(n12295), .ZN(n12294) );
  NOR2_X1 U12333 ( .A1(n12125), .A2(n12123), .ZN(n12295) );
  NOR2_X1 U12334 ( .A1(n11859), .A2(n12296), .ZN(n12126) );
  NAND2_X1 U12335 ( .A1(n12123), .A2(n12125), .ZN(n12292) );
  NAND2_X1 U12336 ( .A1(n12297), .A2(n12298), .ZN(n12125) );
  NAND2_X1 U12337 ( .A1(n12063), .A2(n12299), .ZN(n12298) );
  INV_X1 U12338 ( .A(n12300), .ZN(n12299) );
  NOR2_X1 U12339 ( .A1(n12062), .A2(n12061), .ZN(n12300) );
  NOR2_X1 U12340 ( .A1(n11859), .A2(n12301), .ZN(n12063) );
  NAND2_X1 U12341 ( .A1(n12061), .A2(n12062), .ZN(n12297) );
  NAND2_X1 U12342 ( .A1(n12302), .A2(n12303), .ZN(n12062) );
  NAND2_X1 U12343 ( .A1(n12071), .A2(n12304), .ZN(n12303) );
  INV_X1 U12344 ( .A(n12305), .ZN(n12304) );
  NOR2_X1 U12345 ( .A1(n12070), .A2(n12069), .ZN(n12305) );
  NOR2_X1 U12346 ( .A1(n11859), .A2(n8779), .ZN(n12071) );
  NAND2_X1 U12347 ( .A1(n12069), .A2(n12070), .ZN(n12302) );
  NAND2_X1 U12348 ( .A1(n12306), .A2(n12307), .ZN(n12070) );
  NAND2_X1 U12349 ( .A1(n12122), .A2(n12308), .ZN(n12307) );
  NAND2_X1 U12350 ( .A1(n12119), .A2(n12121), .ZN(n12308) );
  NOR2_X1 U12351 ( .A1(n11859), .A2(n8788), .ZN(n12122) );
  INV_X1 U12352 ( .A(n12309), .ZN(n12306) );
  NOR2_X1 U12353 ( .A1(n12121), .A2(n12119), .ZN(n12309) );
  XNOR2_X1 U12354 ( .A(n12310), .B(n12311), .ZN(n12119) );
  XNOR2_X1 U12355 ( .A(n12312), .B(n12313), .ZN(n12311) );
  NAND2_X1 U12356 ( .A1(n12314), .A2(n12315), .ZN(n12121) );
  NAND2_X1 U12357 ( .A1(n12080), .A2(n12316), .ZN(n12315) );
  NAND2_X1 U12358 ( .A1(n12083), .A2(n12082), .ZN(n12316) );
  XNOR2_X1 U12359 ( .A(n12317), .B(n12318), .ZN(n12080) );
  XOR2_X1 U12360 ( .A(n12319), .B(n12320), .Z(n12317) );
  INV_X1 U12361 ( .A(n12321), .ZN(n12314) );
  NOR2_X1 U12362 ( .A1(n12082), .A2(n12083), .ZN(n12321) );
  NOR2_X1 U12363 ( .A1(n11859), .A2(n9344), .ZN(n12083) );
  NAND2_X1 U12364 ( .A1(n12322), .A2(n12323), .ZN(n12082) );
  NAND2_X1 U12365 ( .A1(n12090), .A2(n12324), .ZN(n12323) );
  INV_X1 U12366 ( .A(n12325), .ZN(n12324) );
  NOR2_X1 U12367 ( .A1(n12089), .A2(n12088), .ZN(n12325) );
  NOR2_X1 U12368 ( .A1(n11859), .A2(n8797), .ZN(n12090) );
  NAND2_X1 U12369 ( .A1(n12088), .A2(n12089), .ZN(n12322) );
  NAND2_X1 U12370 ( .A1(n12326), .A2(n12327), .ZN(n12089) );
  NAND2_X1 U12371 ( .A1(n12117), .A2(n12328), .ZN(n12327) );
  INV_X1 U12372 ( .A(n12329), .ZN(n12328) );
  NOR2_X1 U12373 ( .A1(n12118), .A2(n12116), .ZN(n12329) );
  NOR2_X1 U12374 ( .A1(n11859), .A2(n8314), .ZN(n12117) );
  NAND2_X1 U12375 ( .A1(n12116), .A2(n12118), .ZN(n12326) );
  NAND2_X1 U12376 ( .A1(n12330), .A2(n12331), .ZN(n12118) );
  NAND2_X1 U12377 ( .A1(n12112), .A2(n12332), .ZN(n12331) );
  INV_X1 U12378 ( .A(n12333), .ZN(n12332) );
  NOR2_X1 U12379 ( .A1(n12113), .A2(n12114), .ZN(n12333) );
  NOR2_X1 U12380 ( .A1(n11859), .A2(n9098), .ZN(n12112) );
  NAND2_X1 U12381 ( .A1(n12114), .A2(n12113), .ZN(n12330) );
  NAND2_X1 U12382 ( .A1(n12334), .A2(n12335), .ZN(n12113) );
  NAND2_X1 U12383 ( .A1(b_15_), .A2(n12336), .ZN(n12335) );
  NAND2_X1 U12384 ( .A1(n8299), .A2(n12337), .ZN(n12336) );
  NAND2_X1 U12385 ( .A1(a_31_), .A2(n12110), .ZN(n12337) );
  NAND2_X1 U12386 ( .A1(b_16_), .A2(n12338), .ZN(n12334) );
  NAND2_X1 U12387 ( .A1(n8303), .A2(n12339), .ZN(n12338) );
  NAND2_X1 U12388 ( .A1(a_30_), .A2(n12340), .ZN(n12339) );
  NOR3_X1 U12389 ( .A1(n11859), .A2(n9631), .A3(n12110), .ZN(n12114) );
  XOR2_X1 U12390 ( .A(n12341), .B(n12342), .Z(n12116) );
  XOR2_X1 U12391 ( .A(n12343), .B(n12344), .Z(n12341) );
  XOR2_X1 U12392 ( .A(n12345), .B(n12346), .Z(n12088) );
  XOR2_X1 U12393 ( .A(n12347), .B(n12348), .Z(n12345) );
  XNOR2_X1 U12394 ( .A(n12349), .B(n12350), .ZN(n12069) );
  XNOR2_X1 U12395 ( .A(n12351), .B(n12352), .ZN(n12350) );
  XOR2_X1 U12396 ( .A(n12353), .B(n12354), .Z(n12061) );
  XOR2_X1 U12397 ( .A(n12355), .B(n12356), .Z(n12353) );
  XNOR2_X1 U12398 ( .A(n12357), .B(n12358), .ZN(n12123) );
  NAND2_X1 U12399 ( .A1(n12359), .A2(n12360), .ZN(n12357) );
  XNOR2_X1 U12400 ( .A(n12361), .B(n12362), .ZN(n12127) );
  NAND2_X1 U12401 ( .A1(n12363), .A2(n12364), .ZN(n12361) );
  XOR2_X1 U12402 ( .A(n12365), .B(n12366), .Z(n12035) );
  XNOR2_X1 U12403 ( .A(n12367), .B(n12368), .ZN(n12366) );
  NAND2_X1 U12404 ( .A1(b_16_), .A2(a_19_), .ZN(n12368) );
  XOR2_X1 U12405 ( .A(n12369), .B(n12370), .Z(n12020) );
  XNOR2_X1 U12406 ( .A(n12371), .B(n12372), .ZN(n12369) );
  XOR2_X1 U12407 ( .A(n12373), .B(n12374), .Z(n12012) );
  XNOR2_X1 U12408 ( .A(n12375), .B(n12376), .ZN(n12374) );
  NAND2_X1 U12409 ( .A1(b_16_), .A2(a_15_), .ZN(n12376) );
  XNOR2_X1 U12410 ( .A(n12377), .B(n12378), .ZN(n12148) );
  XOR2_X1 U12411 ( .A(n12379), .B(n12380), .Z(n12378) );
  NAND2_X1 U12412 ( .A1(b_16_), .A2(a_14_), .ZN(n12380) );
  XNOR2_X1 U12413 ( .A(n12381), .B(n12382), .ZN(n12152) );
  XNOR2_X1 U12414 ( .A(n12383), .B(n12384), .ZN(n12381) );
  XNOR2_X1 U12415 ( .A(n12385), .B(n12386), .ZN(n12155) );
  XOR2_X1 U12416 ( .A(n12387), .B(n12388), .Z(n12385) );
  XNOR2_X1 U12417 ( .A(n12389), .B(n12390), .ZN(n12159) );
  XOR2_X1 U12418 ( .A(n12391), .B(n12392), .Z(n12389) );
  NOR2_X1 U12419 ( .A1(n8867), .A2(n12110), .ZN(n12392) );
  XOR2_X1 U12420 ( .A(n12393), .B(n12394), .Z(n11989) );
  NAND2_X1 U12421 ( .A1(n12395), .A2(n12396), .ZN(n12393) );
  XNOR2_X1 U12422 ( .A(n12397), .B(n12398), .ZN(n11981) );
  XOR2_X1 U12423 ( .A(n12399), .B(n12400), .Z(n12397) );
  NOR2_X1 U12424 ( .A1(n8971), .A2(n12110), .ZN(n12400) );
  XOR2_X1 U12425 ( .A(n12401), .B(n12402), .Z(n11972) );
  NAND2_X1 U12426 ( .A1(n12403), .A2(n12404), .ZN(n12401) );
  XNOR2_X1 U12427 ( .A(n12405), .B(n12406), .ZN(n11964) );
  NAND2_X1 U12428 ( .A1(n12407), .A2(n12408), .ZN(n12405) );
  XNOR2_X1 U12429 ( .A(n12409), .B(n12410), .ZN(n12163) );
  NAND2_X1 U12430 ( .A1(n12411), .A2(n12412), .ZN(n12409) );
  XOR2_X1 U12431 ( .A(n12413), .B(n12414), .Z(n12168) );
  XOR2_X1 U12432 ( .A(n12415), .B(n12416), .Z(n12413) );
  XOR2_X1 U12433 ( .A(n12417), .B(n12418), .Z(n12171) );
  XOR2_X1 U12434 ( .A(n12419), .B(n12420), .Z(n12417) );
  NOR2_X1 U12435 ( .A1(n8439), .A2(n12110), .ZN(n12420) );
  XNOR2_X1 U12436 ( .A(n12421), .B(n12422), .ZN(n11943) );
  NAND2_X1 U12437 ( .A1(n12423), .A2(n12424), .ZN(n12421) );
  XOR2_X1 U12438 ( .A(n12425), .B(n12426), .Z(n11931) );
  NAND2_X1 U12439 ( .A1(n12427), .A2(n12428), .ZN(n12425) );
  XOR2_X1 U12440 ( .A(n12429), .B(n12430), .Z(n8595) );
  NAND2_X1 U12441 ( .A1(n12431), .A2(n12432), .ZN(n8534) );
  NAND2_X1 U12442 ( .A1(n12433), .A2(n12434), .ZN(n12432) );
  NAND2_X1 U12443 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  NAND4_X1 U12444 ( .A1(n12430), .A2(n12433), .A3(n12429), .A4(n12434), .ZN(
        n8535) );
  INV_X1 U12445 ( .A(n8591), .ZN(n12434) );
  NAND2_X1 U12446 ( .A1(n12427), .A2(n12435), .ZN(n12429) );
  NAND2_X1 U12447 ( .A1(n12426), .A2(n12428), .ZN(n12435) );
  NAND2_X1 U12448 ( .A1(n12436), .A2(n12437), .ZN(n12428) );
  NAND2_X1 U12449 ( .A1(b_16_), .A2(a_0_), .ZN(n12437) );
  XNOR2_X1 U12450 ( .A(n12438), .B(n12439), .ZN(n12426) );
  XOR2_X1 U12451 ( .A(n12440), .B(n12441), .Z(n12438) );
  NAND2_X1 U12452 ( .A1(a_0_), .A2(n12442), .ZN(n12427) );
  INV_X1 U12453 ( .A(n12436), .ZN(n12442) );
  NOR2_X1 U12454 ( .A1(n12443), .A2(n12444), .ZN(n12436) );
  NOR3_X1 U12455 ( .A1(n8569), .A2(n12445), .A3(n12110), .ZN(n12444) );
  INV_X1 U12456 ( .A(n12446), .ZN(n12445) );
  NAND2_X1 U12457 ( .A1(n12185), .A2(n12186), .ZN(n12446) );
  NOR2_X1 U12458 ( .A1(n12185), .A2(n12186), .ZN(n12443) );
  NAND2_X1 U12459 ( .A1(n12447), .A2(n12448), .ZN(n12186) );
  NAND2_X1 U12460 ( .A1(n12191), .A2(n12449), .ZN(n12448) );
  NAND2_X1 U12461 ( .A1(n12194), .A2(n12193), .ZN(n12449) );
  XOR2_X1 U12462 ( .A(n12450), .B(n12451), .Z(n12191) );
  XNOR2_X1 U12463 ( .A(n12452), .B(n12453), .ZN(n12450) );
  NOR2_X1 U12464 ( .A1(n8900), .A2(n12340), .ZN(n12453) );
  INV_X1 U12465 ( .A(n12454), .ZN(n12447) );
  NOR2_X1 U12466 ( .A1(n12193), .A2(n12194), .ZN(n12454) );
  NOR2_X1 U12467 ( .A1(n12110), .A2(n8448), .ZN(n12194) );
  NAND2_X1 U12468 ( .A1(n12423), .A2(n12455), .ZN(n12193) );
  NAND2_X1 U12469 ( .A1(n12422), .A2(n12424), .ZN(n12455) );
  NAND2_X1 U12470 ( .A1(n12456), .A2(n12457), .ZN(n12424) );
  NAND2_X1 U12471 ( .A1(b_16_), .A2(a_3_), .ZN(n12457) );
  INV_X1 U12472 ( .A(n12458), .ZN(n12456) );
  XOR2_X1 U12473 ( .A(n12459), .B(n12460), .Z(n12422) );
  XNOR2_X1 U12474 ( .A(n12461), .B(n12462), .ZN(n12460) );
  NAND2_X1 U12475 ( .A1(b_15_), .A2(a_4_), .ZN(n12462) );
  NAND2_X1 U12476 ( .A1(a_3_), .A2(n12458), .ZN(n12423) );
  NAND2_X1 U12477 ( .A1(n12463), .A2(n12464), .ZN(n12458) );
  INV_X1 U12478 ( .A(n12465), .ZN(n12464) );
  NOR3_X1 U12479 ( .A1(n8439), .A2(n12466), .A3(n12110), .ZN(n12465) );
  NOR2_X1 U12480 ( .A1(n12418), .A2(n12419), .ZN(n12466) );
  NAND2_X1 U12481 ( .A1(n12418), .A2(n12419), .ZN(n12463) );
  NAND2_X1 U12482 ( .A1(n12467), .A2(n12468), .ZN(n12419) );
  NAND2_X1 U12483 ( .A1(n12416), .A2(n12469), .ZN(n12468) );
  INV_X1 U12484 ( .A(n12470), .ZN(n12469) );
  NOR2_X1 U12485 ( .A1(n12415), .A2(n12414), .ZN(n12470) );
  NOR2_X1 U12486 ( .A1(n12110), .A2(n8938), .ZN(n12416) );
  NAND2_X1 U12487 ( .A1(n12414), .A2(n12415), .ZN(n12467) );
  NAND2_X1 U12488 ( .A1(n12411), .A2(n12471), .ZN(n12415) );
  NAND2_X1 U12489 ( .A1(n12410), .A2(n12412), .ZN(n12471) );
  NAND2_X1 U12490 ( .A1(n12472), .A2(n12473), .ZN(n12412) );
  NAND2_X1 U12491 ( .A1(b_16_), .A2(a_6_), .ZN(n12473) );
  INV_X1 U12492 ( .A(n12474), .ZN(n12472) );
  XNOR2_X1 U12493 ( .A(n12475), .B(n12476), .ZN(n12410) );
  XNOR2_X1 U12494 ( .A(n12477), .B(n12478), .ZN(n12475) );
  NOR2_X1 U12495 ( .A1(n8425), .A2(n12340), .ZN(n12478) );
  NAND2_X1 U12496 ( .A1(a_6_), .A2(n12474), .ZN(n12411) );
  NAND2_X1 U12497 ( .A1(n12407), .A2(n12479), .ZN(n12474) );
  NAND2_X1 U12498 ( .A1(n12406), .A2(n12408), .ZN(n12479) );
  NAND2_X1 U12499 ( .A1(n12480), .A2(n12481), .ZN(n12408) );
  NAND2_X1 U12500 ( .A1(b_16_), .A2(a_7_), .ZN(n12481) );
  INV_X1 U12501 ( .A(n12482), .ZN(n12480) );
  XOR2_X1 U12502 ( .A(n12483), .B(n12484), .Z(n12406) );
  XNOR2_X1 U12503 ( .A(n12485), .B(n12486), .ZN(n12484) );
  NAND2_X1 U12504 ( .A1(b_15_), .A2(a_8_), .ZN(n12486) );
  NAND2_X1 U12505 ( .A1(a_7_), .A2(n12482), .ZN(n12407) );
  NAND2_X1 U12506 ( .A1(n12403), .A2(n12487), .ZN(n12482) );
  NAND2_X1 U12507 ( .A1(n12402), .A2(n12404), .ZN(n12487) );
  NAND2_X1 U12508 ( .A1(n12488), .A2(n12489), .ZN(n12404) );
  NAND2_X1 U12509 ( .A1(b_16_), .A2(a_8_), .ZN(n12489) );
  INV_X1 U12510 ( .A(n12490), .ZN(n12488) );
  XNOR2_X1 U12511 ( .A(n12491), .B(n12492), .ZN(n12402) );
  XNOR2_X1 U12512 ( .A(n12493), .B(n12494), .ZN(n12491) );
  NOR2_X1 U12513 ( .A1(n8971), .A2(n12340), .ZN(n12494) );
  NAND2_X1 U12514 ( .A1(a_8_), .A2(n12490), .ZN(n12403) );
  NAND2_X1 U12515 ( .A1(n12495), .A2(n12496), .ZN(n12490) );
  INV_X1 U12516 ( .A(n12497), .ZN(n12496) );
  NOR3_X1 U12517 ( .A1(n8971), .A2(n12498), .A3(n12110), .ZN(n12497) );
  NOR2_X1 U12518 ( .A1(n12398), .A2(n12399), .ZN(n12498) );
  NAND2_X1 U12519 ( .A1(n12398), .A2(n12399), .ZN(n12495) );
  NAND2_X1 U12520 ( .A1(n12395), .A2(n12499), .ZN(n12399) );
  NAND2_X1 U12521 ( .A1(n12394), .A2(n12396), .ZN(n12499) );
  NAND2_X1 U12522 ( .A1(n12500), .A2(n12501), .ZN(n12396) );
  NAND2_X1 U12523 ( .A1(b_16_), .A2(a_10_), .ZN(n12501) );
  INV_X1 U12524 ( .A(n12502), .ZN(n12500) );
  XOR2_X1 U12525 ( .A(n12503), .B(n12504), .Z(n12394) );
  XOR2_X1 U12526 ( .A(n12505), .B(n12506), .Z(n12503) );
  NOR2_X1 U12527 ( .A1(n8867), .A2(n12340), .ZN(n12506) );
  NAND2_X1 U12528 ( .A1(a_10_), .A2(n12502), .ZN(n12395) );
  NAND2_X1 U12529 ( .A1(n12507), .A2(n12508), .ZN(n12502) );
  INV_X1 U12530 ( .A(n12509), .ZN(n12508) );
  NOR3_X1 U12531 ( .A1(n8867), .A2(n12510), .A3(n12110), .ZN(n12509) );
  NOR2_X1 U12532 ( .A1(n12390), .A2(n12391), .ZN(n12510) );
  NAND2_X1 U12533 ( .A1(n12390), .A2(n12391), .ZN(n12507) );
  NAND2_X1 U12534 ( .A1(n12511), .A2(n12512), .ZN(n12391) );
  NAND2_X1 U12535 ( .A1(n12388), .A2(n12513), .ZN(n12512) );
  INV_X1 U12536 ( .A(n12514), .ZN(n12513) );
  NOR2_X1 U12537 ( .A1(n12387), .A2(n12386), .ZN(n12514) );
  NOR2_X1 U12538 ( .A1(n12110), .A2(n8393), .ZN(n12388) );
  NAND2_X1 U12539 ( .A1(n12386), .A2(n12387), .ZN(n12511) );
  NAND2_X1 U12540 ( .A1(n12515), .A2(n12516), .ZN(n12387) );
  NAND2_X1 U12541 ( .A1(n12384), .A2(n12517), .ZN(n12516) );
  NAND2_X1 U12542 ( .A1(n12382), .A2(n12383), .ZN(n12517) );
  NOR2_X1 U12543 ( .A1(n12110), .A2(n8996), .ZN(n12384) );
  INV_X1 U12544 ( .A(n12518), .ZN(n12515) );
  NOR2_X1 U12545 ( .A1(n12382), .A2(n12383), .ZN(n12518) );
  NOR2_X1 U12546 ( .A1(n12519), .A2(n12520), .ZN(n12383) );
  NOR3_X1 U12547 ( .A1(n9262), .A2(n12521), .A3(n12110), .ZN(n12520) );
  NOR2_X1 U12548 ( .A1(n12379), .A2(n12377), .ZN(n12521) );
  INV_X1 U12549 ( .A(n12522), .ZN(n12519) );
  NAND2_X1 U12550 ( .A1(n12377), .A2(n12379), .ZN(n12522) );
  NAND2_X1 U12551 ( .A1(n12523), .A2(n12524), .ZN(n12379) );
  INV_X1 U12552 ( .A(n12525), .ZN(n12524) );
  NOR3_X1 U12553 ( .A1(n8850), .A2(n12526), .A3(n12110), .ZN(n12525) );
  NOR2_X1 U12554 ( .A1(n12373), .A2(n12375), .ZN(n12526) );
  NAND2_X1 U12555 ( .A1(n12373), .A2(n12375), .ZN(n12523) );
  NOR2_X1 U12556 ( .A1(n12527), .A2(n12528), .ZN(n12375) );
  INV_X1 U12557 ( .A(n12529), .ZN(n12528) );
  NAND2_X1 U12558 ( .A1(n12530), .A2(n12372), .ZN(n12529) );
  NAND2_X1 U12559 ( .A1(n12370), .A2(n12371), .ZN(n12530) );
  NOR2_X1 U12560 ( .A1(n12370), .A2(n12371), .ZN(n12527) );
  NAND2_X1 U12561 ( .A1(n12531), .A2(n12532), .ZN(n12371) );
  NAND3_X1 U12562 ( .A1(a_17_), .A2(n12533), .A3(b_16_), .ZN(n12532) );
  NAND2_X1 U12563 ( .A1(n12256), .A2(n12257), .ZN(n12533) );
  INV_X1 U12564 ( .A(n12534), .ZN(n12531) );
  NOR2_X1 U12565 ( .A1(n12256), .A2(n12257), .ZN(n12534) );
  NAND2_X1 U12566 ( .A1(n12535), .A2(n12536), .ZN(n12257) );
  NAND2_X1 U12567 ( .A1(n12264), .A2(n12537), .ZN(n12536) );
  NAND2_X1 U12568 ( .A1(n12267), .A2(n12266), .ZN(n12537) );
  XNOR2_X1 U12569 ( .A(n12538), .B(n12539), .ZN(n12264) );
  XNOR2_X1 U12570 ( .A(n12540), .B(n12541), .ZN(n12539) );
  NAND2_X1 U12571 ( .A1(b_15_), .A2(a_19_), .ZN(n12541) );
  INV_X1 U12572 ( .A(n12542), .ZN(n12535) );
  NOR2_X1 U12573 ( .A1(n12266), .A2(n12267), .ZN(n12542) );
  NOR2_X1 U12574 ( .A1(n12110), .A2(n9291), .ZN(n12267) );
  NAND2_X1 U12575 ( .A1(n12543), .A2(n12544), .ZN(n12266) );
  NAND3_X1 U12576 ( .A1(a_19_), .A2(n12545), .A3(b_16_), .ZN(n12544) );
  NAND2_X1 U12577 ( .A1(n12367), .A2(n12365), .ZN(n12545) );
  INV_X1 U12578 ( .A(n12546), .ZN(n12543) );
  NOR2_X1 U12579 ( .A1(n12365), .A2(n12367), .ZN(n12546) );
  NOR2_X1 U12580 ( .A1(n12547), .A2(n12548), .ZN(n12367) );
  INV_X1 U12581 ( .A(n12549), .ZN(n12548) );
  NAND3_X1 U12582 ( .A1(a_20_), .A2(n12550), .A3(b_16_), .ZN(n12549) );
  NAND2_X1 U12583 ( .A1(n12277), .A2(n12278), .ZN(n12550) );
  NOR2_X1 U12584 ( .A1(n12277), .A2(n12278), .ZN(n12547) );
  NOR2_X1 U12585 ( .A1(n12551), .A2(n12552), .ZN(n12278) );
  NOR3_X1 U12586 ( .A1(n8759), .A2(n12553), .A3(n12110), .ZN(n12552) );
  NOR2_X1 U12587 ( .A1(n12285), .A2(n12284), .ZN(n12553) );
  INV_X1 U12588 ( .A(n12554), .ZN(n12551) );
  NAND2_X1 U12589 ( .A1(n12284), .A2(n12285), .ZN(n12554) );
  NAND2_X1 U12590 ( .A1(n12363), .A2(n12555), .ZN(n12285) );
  NAND2_X1 U12591 ( .A1(n12362), .A2(n12364), .ZN(n12555) );
  NAND2_X1 U12592 ( .A1(n12556), .A2(n12557), .ZN(n12364) );
  NAND2_X1 U12593 ( .A1(b_16_), .A2(a_22_), .ZN(n12557) );
  INV_X1 U12594 ( .A(n12558), .ZN(n12556) );
  XOR2_X1 U12595 ( .A(n12559), .B(n12560), .Z(n12362) );
  XOR2_X1 U12596 ( .A(n12561), .B(n12562), .Z(n12559) );
  NAND2_X1 U12597 ( .A1(a_22_), .A2(n12558), .ZN(n12363) );
  NAND2_X1 U12598 ( .A1(n12359), .A2(n12563), .ZN(n12558) );
  NAND2_X1 U12599 ( .A1(n12358), .A2(n12360), .ZN(n12563) );
  NAND2_X1 U12600 ( .A1(n12564), .A2(n12565), .ZN(n12360) );
  NAND2_X1 U12601 ( .A1(b_16_), .A2(a_23_), .ZN(n12565) );
  INV_X1 U12602 ( .A(n12566), .ZN(n12564) );
  XOR2_X1 U12603 ( .A(n12567), .B(n12568), .Z(n12358) );
  XOR2_X1 U12604 ( .A(n12569), .B(n12570), .Z(n12567) );
  NAND2_X1 U12605 ( .A1(a_23_), .A2(n12566), .ZN(n12359) );
  NAND2_X1 U12606 ( .A1(n12571), .A2(n12572), .ZN(n12566) );
  NAND2_X1 U12607 ( .A1(n12356), .A2(n12573), .ZN(n12572) );
  INV_X1 U12608 ( .A(n12574), .ZN(n12573) );
  NOR2_X1 U12609 ( .A1(n12354), .A2(n12355), .ZN(n12574) );
  NOR2_X1 U12610 ( .A1(n12110), .A2(n8779), .ZN(n12356) );
  NAND2_X1 U12611 ( .A1(n12354), .A2(n12355), .ZN(n12571) );
  NAND2_X1 U12612 ( .A1(n12575), .A2(n12576), .ZN(n12355) );
  NAND2_X1 U12613 ( .A1(n12352), .A2(n12577), .ZN(n12576) );
  NAND2_X1 U12614 ( .A1(n12349), .A2(n12351), .ZN(n12577) );
  NOR2_X1 U12615 ( .A1(n12110), .A2(n8788), .ZN(n12352) );
  INV_X1 U12616 ( .A(n12578), .ZN(n12575) );
  NOR2_X1 U12617 ( .A1(n12351), .A2(n12349), .ZN(n12578) );
  XNOR2_X1 U12618 ( .A(n12579), .B(n12580), .ZN(n12349) );
  XNOR2_X1 U12619 ( .A(n12581), .B(n12582), .ZN(n12580) );
  NAND2_X1 U12620 ( .A1(n12583), .A2(n12584), .ZN(n12351) );
  NAND2_X1 U12621 ( .A1(n12310), .A2(n12585), .ZN(n12584) );
  NAND2_X1 U12622 ( .A1(n12313), .A2(n12312), .ZN(n12585) );
  XNOR2_X1 U12623 ( .A(n12586), .B(n12587), .ZN(n12310) );
  XOR2_X1 U12624 ( .A(n12588), .B(n12589), .Z(n12586) );
  INV_X1 U12625 ( .A(n12590), .ZN(n12583) );
  NOR2_X1 U12626 ( .A1(n12312), .A2(n12313), .ZN(n12590) );
  NOR2_X1 U12627 ( .A1(n12110), .A2(n9344), .ZN(n12313) );
  NAND2_X1 U12628 ( .A1(n12591), .A2(n12592), .ZN(n12312) );
  NAND2_X1 U12629 ( .A1(n12320), .A2(n12593), .ZN(n12592) );
  INV_X1 U12630 ( .A(n12594), .ZN(n12593) );
  NOR2_X1 U12631 ( .A1(n12318), .A2(n12319), .ZN(n12594) );
  NOR2_X1 U12632 ( .A1(n12110), .A2(n8797), .ZN(n12320) );
  NAND2_X1 U12633 ( .A1(n12318), .A2(n12319), .ZN(n12591) );
  NAND2_X1 U12634 ( .A1(n12595), .A2(n12596), .ZN(n12319) );
  NAND2_X1 U12635 ( .A1(n12347), .A2(n12597), .ZN(n12596) );
  INV_X1 U12636 ( .A(n12598), .ZN(n12597) );
  NOR2_X1 U12637 ( .A1(n12348), .A2(n12346), .ZN(n12598) );
  NOR2_X1 U12638 ( .A1(n12110), .A2(n8314), .ZN(n12347) );
  NAND2_X1 U12639 ( .A1(n12346), .A2(n12348), .ZN(n12595) );
  NAND2_X1 U12640 ( .A1(n12599), .A2(n12600), .ZN(n12348) );
  NAND2_X1 U12641 ( .A1(n12342), .A2(n12601), .ZN(n12600) );
  INV_X1 U12642 ( .A(n12602), .ZN(n12601) );
  NOR2_X1 U12643 ( .A1(n12343), .A2(n12344), .ZN(n12602) );
  NOR2_X1 U12644 ( .A1(n12110), .A2(n9098), .ZN(n12342) );
  NAND2_X1 U12645 ( .A1(n12344), .A2(n12343), .ZN(n12599) );
  NAND2_X1 U12646 ( .A1(n12603), .A2(n12604), .ZN(n12343) );
  NAND2_X1 U12647 ( .A1(b_14_), .A2(n12605), .ZN(n12604) );
  NAND2_X1 U12648 ( .A1(n8299), .A2(n12606), .ZN(n12605) );
  NAND2_X1 U12649 ( .A1(a_31_), .A2(n12340), .ZN(n12606) );
  NAND2_X1 U12650 ( .A1(b_15_), .A2(n12607), .ZN(n12603) );
  NAND2_X1 U12651 ( .A1(n8303), .A2(n12608), .ZN(n12607) );
  NAND2_X1 U12652 ( .A1(a_30_), .A2(n12609), .ZN(n12608) );
  NOR3_X1 U12653 ( .A1(n12340), .A2(n9631), .A3(n12110), .ZN(n12344) );
  XOR2_X1 U12654 ( .A(n12610), .B(n12611), .Z(n12346) );
  XOR2_X1 U12655 ( .A(n12612), .B(n12613), .Z(n12610) );
  XOR2_X1 U12656 ( .A(n12614), .B(n12615), .Z(n12318) );
  XOR2_X1 U12657 ( .A(n12616), .B(n12617), .Z(n12614) );
  XNOR2_X1 U12658 ( .A(n12618), .B(n12619), .ZN(n12354) );
  XNOR2_X1 U12659 ( .A(n12620), .B(n12621), .ZN(n12619) );
  XNOR2_X1 U12660 ( .A(n12622), .B(n12623), .ZN(n12284) );
  XNOR2_X1 U12661 ( .A(n12624), .B(n12625), .ZN(n12623) );
  XNOR2_X1 U12662 ( .A(n12626), .B(n12627), .ZN(n12277) );
  XOR2_X1 U12663 ( .A(n12628), .B(n12629), .Z(n12626) );
  NOR2_X1 U12664 ( .A1(n8759), .A2(n12340), .ZN(n12629) );
  XOR2_X1 U12665 ( .A(n12630), .B(n12631), .Z(n12365) );
  XNOR2_X1 U12666 ( .A(n12632), .B(n12633), .ZN(n12630) );
  NOR2_X1 U12667 ( .A1(n9047), .A2(n12340), .ZN(n12633) );
  XOR2_X1 U12668 ( .A(n12634), .B(n12635), .Z(n12256) );
  XOR2_X1 U12669 ( .A(n12636), .B(n12637), .Z(n12635) );
  NAND2_X1 U12670 ( .A1(b_15_), .A2(a_18_), .ZN(n12637) );
  XNOR2_X1 U12671 ( .A(n12638), .B(n12639), .ZN(n12370) );
  XOR2_X1 U12672 ( .A(n12640), .B(n12641), .Z(n12639) );
  NAND2_X1 U12673 ( .A1(b_15_), .A2(a_17_), .ZN(n12641) );
  XNOR2_X1 U12674 ( .A(n12642), .B(n12643), .ZN(n12373) );
  XOR2_X1 U12675 ( .A(n12644), .B(n12645), .Z(n12643) );
  XNOR2_X1 U12676 ( .A(n12646), .B(n12647), .ZN(n12377) );
  XNOR2_X1 U12677 ( .A(n12648), .B(n12649), .ZN(n12646) );
  XOR2_X1 U12678 ( .A(n12650), .B(n12651), .Z(n12382) );
  NAND2_X1 U12679 ( .A1(n12652), .A2(n12653), .ZN(n12650) );
  XNOR2_X1 U12680 ( .A(n12654), .B(n12655), .ZN(n12386) );
  XOR2_X1 U12681 ( .A(n12656), .B(n12657), .Z(n12655) );
  NAND2_X1 U12682 ( .A1(b_15_), .A2(a_13_), .ZN(n12657) );
  XNOR2_X1 U12683 ( .A(n12658), .B(n12659), .ZN(n12390) );
  XOR2_X1 U12684 ( .A(n12660), .B(n12661), .Z(n12659) );
  NAND2_X1 U12685 ( .A1(b_15_), .A2(a_12_), .ZN(n12661) );
  XNOR2_X1 U12686 ( .A(n12662), .B(n12663), .ZN(n12398) );
  XOR2_X1 U12687 ( .A(n12664), .B(n12665), .Z(n12663) );
  NAND2_X1 U12688 ( .A1(b_15_), .A2(a_10_), .ZN(n12665) );
  XOR2_X1 U12689 ( .A(n12666), .B(n12667), .Z(n12414) );
  XNOR2_X1 U12690 ( .A(n12668), .B(n12669), .ZN(n12667) );
  NAND2_X1 U12691 ( .A1(b_15_), .A2(a_6_), .ZN(n12669) );
  XNOR2_X1 U12692 ( .A(n12670), .B(n12671), .ZN(n12418) );
  XNOR2_X1 U12693 ( .A(n12672), .B(n12673), .ZN(n12670) );
  NOR2_X1 U12694 ( .A1(n8938), .A2(n12340), .ZN(n12673) );
  XNOR2_X1 U12695 ( .A(n12674), .B(n12675), .ZN(n12185) );
  XNOR2_X1 U12696 ( .A(n12676), .B(n12677), .ZN(n12675) );
  NAND2_X1 U12697 ( .A1(b_15_), .A2(a_2_), .ZN(n12677) );
  NAND2_X1 U12698 ( .A1(n12678), .A2(n12679), .ZN(n12433) );
  XNOR2_X1 U12699 ( .A(n12680), .B(n12681), .ZN(n12430) );
  XOR2_X1 U12700 ( .A(n12682), .B(n12683), .Z(n12681) );
  NAND2_X1 U12701 ( .A1(b_15_), .A2(a_0_), .ZN(n12683) );
  NOR2_X1 U12702 ( .A1(n12679), .A2(n12678), .ZN(n8591) );
  NOR2_X1 U12703 ( .A1(n12684), .A2(n12685), .ZN(n12678) );
  INV_X1 U12704 ( .A(n12686), .ZN(n12685) );
  NAND3_X1 U12705 ( .A1(a_0_), .A2(n12687), .A3(b_15_), .ZN(n12686) );
  NAND2_X1 U12706 ( .A1(n12680), .A2(n12682), .ZN(n12687) );
  NOR2_X1 U12707 ( .A1(n12682), .A2(n12680), .ZN(n12684) );
  XNOR2_X1 U12708 ( .A(n12688), .B(n12689), .ZN(n12680) );
  XOR2_X1 U12709 ( .A(n12690), .B(n12691), .Z(n12689) );
  NAND2_X1 U12710 ( .A1(n12692), .A2(n12693), .ZN(n12682) );
  NAND2_X1 U12711 ( .A1(n12439), .A2(n12694), .ZN(n12693) );
  NAND2_X1 U12712 ( .A1(n12441), .A2(n12440), .ZN(n12694) );
  XNOR2_X1 U12713 ( .A(n12695), .B(n12696), .ZN(n12439) );
  XNOR2_X1 U12714 ( .A(n12697), .B(n12698), .ZN(n12696) );
  INV_X1 U12715 ( .A(n12699), .ZN(n12692) );
  NOR2_X1 U12716 ( .A1(n12440), .A2(n12441), .ZN(n12699) );
  NOR2_X1 U12717 ( .A1(n12340), .A2(n8569), .ZN(n12441) );
  NAND2_X1 U12718 ( .A1(n12700), .A2(n12701), .ZN(n12440) );
  NAND3_X1 U12719 ( .A1(a_2_), .A2(n12702), .A3(b_15_), .ZN(n12701) );
  NAND2_X1 U12720 ( .A1(n12676), .A2(n12674), .ZN(n12702) );
  INV_X1 U12721 ( .A(n12703), .ZN(n12700) );
  NOR2_X1 U12722 ( .A1(n12674), .A2(n12676), .ZN(n12703) );
  NOR2_X1 U12723 ( .A1(n12704), .A2(n12705), .ZN(n12676) );
  INV_X1 U12724 ( .A(n12706), .ZN(n12705) );
  NAND3_X1 U12725 ( .A1(a_3_), .A2(n12707), .A3(b_15_), .ZN(n12706) );
  NAND2_X1 U12726 ( .A1(n12452), .A2(n12451), .ZN(n12707) );
  NOR2_X1 U12727 ( .A1(n12451), .A2(n12452), .ZN(n12704) );
  NOR2_X1 U12728 ( .A1(n12708), .A2(n12709), .ZN(n12452) );
  NOR3_X1 U12729 ( .A1(n8439), .A2(n12710), .A3(n12340), .ZN(n12709) );
  INV_X1 U12730 ( .A(n12711), .ZN(n12710) );
  NAND2_X1 U12731 ( .A1(n12461), .A2(n12459), .ZN(n12711) );
  NOR2_X1 U12732 ( .A1(n12459), .A2(n12461), .ZN(n12708) );
  NOR2_X1 U12733 ( .A1(n12712), .A2(n12713), .ZN(n12461) );
  INV_X1 U12734 ( .A(n12714), .ZN(n12713) );
  NAND3_X1 U12735 ( .A1(a_5_), .A2(n12715), .A3(b_15_), .ZN(n12714) );
  NAND2_X1 U12736 ( .A1(n12672), .A2(n12671), .ZN(n12715) );
  NOR2_X1 U12737 ( .A1(n12671), .A2(n12672), .ZN(n12712) );
  NOR2_X1 U12738 ( .A1(n12716), .A2(n12717), .ZN(n12672) );
  NOR3_X1 U12739 ( .A1(n8430), .A2(n12718), .A3(n12340), .ZN(n12717) );
  INV_X1 U12740 ( .A(n12719), .ZN(n12718) );
  NAND2_X1 U12741 ( .A1(n12668), .A2(n12666), .ZN(n12719) );
  NOR2_X1 U12742 ( .A1(n12666), .A2(n12668), .ZN(n12716) );
  NOR2_X1 U12743 ( .A1(n12720), .A2(n12721), .ZN(n12668) );
  INV_X1 U12744 ( .A(n12722), .ZN(n12721) );
  NAND3_X1 U12745 ( .A1(a_7_), .A2(n12723), .A3(b_15_), .ZN(n12722) );
  NAND2_X1 U12746 ( .A1(n12477), .A2(n12476), .ZN(n12723) );
  NOR2_X1 U12747 ( .A1(n12476), .A2(n12477), .ZN(n12720) );
  NOR2_X1 U12748 ( .A1(n12724), .A2(n12725), .ZN(n12477) );
  NOR3_X1 U12749 ( .A1(n8968), .A2(n12726), .A3(n12340), .ZN(n12725) );
  INV_X1 U12750 ( .A(n12727), .ZN(n12726) );
  NAND2_X1 U12751 ( .A1(n12485), .A2(n12483), .ZN(n12727) );
  NOR2_X1 U12752 ( .A1(n12483), .A2(n12485), .ZN(n12724) );
  NOR2_X1 U12753 ( .A1(n12728), .A2(n12729), .ZN(n12485) );
  NOR3_X1 U12754 ( .A1(n8971), .A2(n12730), .A3(n12340), .ZN(n12729) );
  INV_X1 U12755 ( .A(n12731), .ZN(n12730) );
  NAND2_X1 U12756 ( .A1(n12493), .A2(n12492), .ZN(n12731) );
  NOR2_X1 U12757 ( .A1(n12492), .A2(n12493), .ZN(n12728) );
  NOR2_X1 U12758 ( .A1(n12732), .A2(n12733), .ZN(n12493) );
  NOR3_X1 U12759 ( .A1(n8402), .A2(n12734), .A3(n12340), .ZN(n12733) );
  NOR2_X1 U12760 ( .A1(n12664), .A2(n12662), .ZN(n12734) );
  INV_X1 U12761 ( .A(n12735), .ZN(n12732) );
  NAND2_X1 U12762 ( .A1(n12662), .A2(n12664), .ZN(n12735) );
  NAND2_X1 U12763 ( .A1(n12736), .A2(n12737), .ZN(n12664) );
  INV_X1 U12764 ( .A(n12738), .ZN(n12737) );
  NOR3_X1 U12765 ( .A1(n8867), .A2(n12739), .A3(n12340), .ZN(n12738) );
  NOR2_X1 U12766 ( .A1(n12505), .A2(n12504), .ZN(n12739) );
  NAND2_X1 U12767 ( .A1(n12504), .A2(n12505), .ZN(n12736) );
  NAND2_X1 U12768 ( .A1(n12740), .A2(n12741), .ZN(n12505) );
  INV_X1 U12769 ( .A(n12742), .ZN(n12741) );
  NOR3_X1 U12770 ( .A1(n8393), .A2(n12743), .A3(n12340), .ZN(n12742) );
  NOR2_X1 U12771 ( .A1(n12660), .A2(n12658), .ZN(n12743) );
  NAND2_X1 U12772 ( .A1(n12658), .A2(n12660), .ZN(n12740) );
  NAND2_X1 U12773 ( .A1(n12744), .A2(n12745), .ZN(n12660) );
  NAND3_X1 U12774 ( .A1(a_13_), .A2(n12746), .A3(b_15_), .ZN(n12745) );
  INV_X1 U12775 ( .A(n12747), .ZN(n12746) );
  NOR2_X1 U12776 ( .A1(n12656), .A2(n12654), .ZN(n12747) );
  NAND2_X1 U12777 ( .A1(n12654), .A2(n12656), .ZN(n12744) );
  NAND2_X1 U12778 ( .A1(n12652), .A2(n12748), .ZN(n12656) );
  NAND2_X1 U12779 ( .A1(n12651), .A2(n12653), .ZN(n12748) );
  NAND2_X1 U12780 ( .A1(n12749), .A2(n12750), .ZN(n12653) );
  NAND2_X1 U12781 ( .A1(b_15_), .A2(a_14_), .ZN(n12749) );
  XOR2_X1 U12782 ( .A(n12751), .B(n12752), .Z(n12651) );
  XOR2_X1 U12783 ( .A(n12753), .B(n12754), .Z(n12752) );
  INV_X1 U12784 ( .A(n12755), .ZN(n12652) );
  NOR2_X1 U12785 ( .A1(n12750), .A2(n9262), .ZN(n12755) );
  NAND2_X1 U12786 ( .A1(n12756), .A2(n12757), .ZN(n12750) );
  NAND2_X1 U12787 ( .A1(n12647), .A2(n12758), .ZN(n12757) );
  NAND2_X1 U12788 ( .A1(n12649), .A2(n12759), .ZN(n12758) );
  INV_X1 U12789 ( .A(n12648), .ZN(n12759) );
  XOR2_X1 U12790 ( .A(n12760), .B(n12761), .Z(n12647) );
  XNOR2_X1 U12791 ( .A(n12762), .B(n12763), .ZN(n12760) );
  NOR2_X1 U12792 ( .A1(n8376), .A2(n12609), .ZN(n12763) );
  NAND2_X1 U12793 ( .A1(n12648), .A2(n12764), .ZN(n12756) );
  NOR2_X1 U12794 ( .A1(n12765), .A2(n12766), .ZN(n12648) );
  NOR2_X1 U12795 ( .A1(n12645), .A2(n12767), .ZN(n12766) );
  NOR2_X1 U12796 ( .A1(n12644), .A2(n12642), .ZN(n12767) );
  NAND2_X1 U12797 ( .A1(b_15_), .A2(a_16_), .ZN(n12645) );
  INV_X1 U12798 ( .A(n12768), .ZN(n12765) );
  NAND2_X1 U12799 ( .A1(n12642), .A2(n12644), .ZN(n12768) );
  NAND2_X1 U12800 ( .A1(n12769), .A2(n12770), .ZN(n12644) );
  INV_X1 U12801 ( .A(n12771), .ZN(n12770) );
  NOR3_X1 U12802 ( .A1(n8371), .A2(n12772), .A3(n12340), .ZN(n12771) );
  NOR2_X1 U12803 ( .A1(n12640), .A2(n12638), .ZN(n12772) );
  NAND2_X1 U12804 ( .A1(n12638), .A2(n12640), .ZN(n12769) );
  NAND2_X1 U12805 ( .A1(n12773), .A2(n12774), .ZN(n12640) );
  NAND3_X1 U12806 ( .A1(a_18_), .A2(n12775), .A3(b_15_), .ZN(n12774) );
  INV_X1 U12807 ( .A(n12776), .ZN(n12775) );
  NOR2_X1 U12808 ( .A1(n12636), .A2(n12634), .ZN(n12776) );
  NAND2_X1 U12809 ( .A1(n12634), .A2(n12636), .ZN(n12773) );
  NAND2_X1 U12810 ( .A1(n12777), .A2(n12778), .ZN(n12636) );
  NAND3_X1 U12811 ( .A1(a_19_), .A2(n12779), .A3(b_15_), .ZN(n12778) );
  NAND2_X1 U12812 ( .A1(n12540), .A2(n12538), .ZN(n12779) );
  INV_X1 U12813 ( .A(n12780), .ZN(n12777) );
  NOR2_X1 U12814 ( .A1(n12538), .A2(n12540), .ZN(n12780) );
  NOR2_X1 U12815 ( .A1(n12781), .A2(n12782), .ZN(n12540) );
  INV_X1 U12816 ( .A(n12783), .ZN(n12782) );
  NAND3_X1 U12817 ( .A1(a_20_), .A2(n12784), .A3(b_15_), .ZN(n12783) );
  NAND2_X1 U12818 ( .A1(n12632), .A2(n12631), .ZN(n12784) );
  NOR2_X1 U12819 ( .A1(n12631), .A2(n12632), .ZN(n12781) );
  NOR2_X1 U12820 ( .A1(n12785), .A2(n12786), .ZN(n12632) );
  NOR3_X1 U12821 ( .A1(n8759), .A2(n12787), .A3(n12340), .ZN(n12786) );
  NOR2_X1 U12822 ( .A1(n12628), .A2(n12627), .ZN(n12787) );
  INV_X1 U12823 ( .A(n12788), .ZN(n12785) );
  NAND2_X1 U12824 ( .A1(n12627), .A2(n12628), .ZN(n12788) );
  NAND2_X1 U12825 ( .A1(n12789), .A2(n12790), .ZN(n12628) );
  NAND2_X1 U12826 ( .A1(n12625), .A2(n12791), .ZN(n12790) );
  INV_X1 U12827 ( .A(n12792), .ZN(n12791) );
  NOR2_X1 U12828 ( .A1(n12624), .A2(n12622), .ZN(n12792) );
  NOR2_X1 U12829 ( .A1(n12340), .A2(n12296), .ZN(n12625) );
  NAND2_X1 U12830 ( .A1(n12622), .A2(n12624), .ZN(n12789) );
  NAND2_X1 U12831 ( .A1(n12793), .A2(n12794), .ZN(n12624) );
  NAND2_X1 U12832 ( .A1(n12562), .A2(n12795), .ZN(n12794) );
  INV_X1 U12833 ( .A(n12796), .ZN(n12795) );
  NOR2_X1 U12834 ( .A1(n12561), .A2(n12560), .ZN(n12796) );
  NOR2_X1 U12835 ( .A1(n12340), .A2(n12301), .ZN(n12562) );
  NAND2_X1 U12836 ( .A1(n12560), .A2(n12561), .ZN(n12793) );
  NAND2_X1 U12837 ( .A1(n12797), .A2(n12798), .ZN(n12561) );
  NAND2_X1 U12838 ( .A1(n12570), .A2(n12799), .ZN(n12798) );
  INV_X1 U12839 ( .A(n12800), .ZN(n12799) );
  NOR2_X1 U12840 ( .A1(n12569), .A2(n12568), .ZN(n12800) );
  NOR2_X1 U12841 ( .A1(n12340), .A2(n8779), .ZN(n12570) );
  NAND2_X1 U12842 ( .A1(n12568), .A2(n12569), .ZN(n12797) );
  NAND2_X1 U12843 ( .A1(n12801), .A2(n12802), .ZN(n12569) );
  NAND2_X1 U12844 ( .A1(n12621), .A2(n12803), .ZN(n12802) );
  NAND2_X1 U12845 ( .A1(n12618), .A2(n12620), .ZN(n12803) );
  NOR2_X1 U12846 ( .A1(n12340), .A2(n8788), .ZN(n12621) );
  INV_X1 U12847 ( .A(n12804), .ZN(n12801) );
  NOR2_X1 U12848 ( .A1(n12620), .A2(n12618), .ZN(n12804) );
  XNOR2_X1 U12849 ( .A(n12805), .B(n12806), .ZN(n12618) );
  XNOR2_X1 U12850 ( .A(n12807), .B(n12808), .ZN(n12806) );
  NAND2_X1 U12851 ( .A1(n12809), .A2(n12810), .ZN(n12620) );
  NAND2_X1 U12852 ( .A1(n12579), .A2(n12811), .ZN(n12810) );
  NAND2_X1 U12853 ( .A1(n12582), .A2(n12581), .ZN(n12811) );
  XNOR2_X1 U12854 ( .A(n12812), .B(n12813), .ZN(n12579) );
  XOR2_X1 U12855 ( .A(n12814), .B(n12815), .Z(n12812) );
  INV_X1 U12856 ( .A(n12816), .ZN(n12809) );
  NOR2_X1 U12857 ( .A1(n12581), .A2(n12582), .ZN(n12816) );
  NOR2_X1 U12858 ( .A1(n12340), .A2(n9344), .ZN(n12582) );
  NAND2_X1 U12859 ( .A1(n12817), .A2(n12818), .ZN(n12581) );
  NAND2_X1 U12860 ( .A1(n12589), .A2(n12819), .ZN(n12818) );
  INV_X1 U12861 ( .A(n12820), .ZN(n12819) );
  NOR2_X1 U12862 ( .A1(n12588), .A2(n12587), .ZN(n12820) );
  NOR2_X1 U12863 ( .A1(n12340), .A2(n8797), .ZN(n12589) );
  NAND2_X1 U12864 ( .A1(n12587), .A2(n12588), .ZN(n12817) );
  NAND2_X1 U12865 ( .A1(n12821), .A2(n12822), .ZN(n12588) );
  NAND2_X1 U12866 ( .A1(n12616), .A2(n12823), .ZN(n12822) );
  INV_X1 U12867 ( .A(n12824), .ZN(n12823) );
  NOR2_X1 U12868 ( .A1(n12617), .A2(n12615), .ZN(n12824) );
  NOR2_X1 U12869 ( .A1(n12340), .A2(n8314), .ZN(n12616) );
  NAND2_X1 U12870 ( .A1(n12615), .A2(n12617), .ZN(n12821) );
  NAND2_X1 U12871 ( .A1(n12825), .A2(n12826), .ZN(n12617) );
  NAND2_X1 U12872 ( .A1(n12611), .A2(n12827), .ZN(n12826) );
  INV_X1 U12873 ( .A(n12828), .ZN(n12827) );
  NOR2_X1 U12874 ( .A1(n12612), .A2(n12613), .ZN(n12828) );
  NOR2_X1 U12875 ( .A1(n12340), .A2(n9098), .ZN(n12611) );
  NAND2_X1 U12876 ( .A1(n12613), .A2(n12612), .ZN(n12825) );
  NAND2_X1 U12877 ( .A1(n12829), .A2(n12830), .ZN(n12612) );
  NAND2_X1 U12878 ( .A1(b_13_), .A2(n12831), .ZN(n12830) );
  NAND2_X1 U12879 ( .A1(n8299), .A2(n12832), .ZN(n12831) );
  NAND2_X1 U12880 ( .A1(a_31_), .A2(n12609), .ZN(n12832) );
  NAND2_X1 U12881 ( .A1(b_14_), .A2(n12833), .ZN(n12829) );
  NAND2_X1 U12882 ( .A1(n8303), .A2(n12834), .ZN(n12833) );
  NAND2_X1 U12883 ( .A1(a_30_), .A2(n12835), .ZN(n12834) );
  NOR3_X1 U12884 ( .A1(n12340), .A2(n9631), .A3(n12609), .ZN(n12613) );
  XOR2_X1 U12885 ( .A(n12836), .B(n12837), .Z(n12615) );
  XOR2_X1 U12886 ( .A(n12838), .B(n12839), .Z(n12836) );
  XOR2_X1 U12887 ( .A(n12840), .B(n12841), .Z(n12587) );
  XOR2_X1 U12888 ( .A(n12842), .B(n12843), .Z(n12840) );
  XNOR2_X1 U12889 ( .A(n12844), .B(n12845), .ZN(n12568) );
  XNOR2_X1 U12890 ( .A(n12846), .B(n12847), .ZN(n12845) );
  XOR2_X1 U12891 ( .A(n12848), .B(n12849), .Z(n12560) );
  XOR2_X1 U12892 ( .A(n12850), .B(n12851), .Z(n12848) );
  XOR2_X1 U12893 ( .A(n12852), .B(n12853), .Z(n12622) );
  XOR2_X1 U12894 ( .A(n12854), .B(n12855), .Z(n12852) );
  XNOR2_X1 U12895 ( .A(n12856), .B(n12857), .ZN(n12627) );
  XNOR2_X1 U12896 ( .A(n12858), .B(n12859), .ZN(n12857) );
  XNOR2_X1 U12897 ( .A(n12860), .B(n12861), .ZN(n12631) );
  XOR2_X1 U12898 ( .A(n12862), .B(n12863), .Z(n12860) );
  NOR2_X1 U12899 ( .A1(n8759), .A2(n12609), .ZN(n12863) );
  XOR2_X1 U12900 ( .A(n12864), .B(n12865), .Z(n12538) );
  XNOR2_X1 U12901 ( .A(n12866), .B(n12867), .ZN(n12864) );
  NOR2_X1 U12902 ( .A1(n9047), .A2(n12609), .ZN(n12867) );
  XOR2_X1 U12903 ( .A(n12868), .B(n12869), .Z(n12634) );
  XNOR2_X1 U12904 ( .A(n12870), .B(n12871), .ZN(n12869) );
  NAND2_X1 U12905 ( .A1(b_14_), .A2(a_19_), .ZN(n12871) );
  XNOR2_X1 U12906 ( .A(n12872), .B(n12873), .ZN(n12638) );
  XOR2_X1 U12907 ( .A(n12874), .B(n12875), .Z(n12873) );
  NAND2_X1 U12908 ( .A1(b_14_), .A2(a_18_), .ZN(n12875) );
  XNOR2_X1 U12909 ( .A(n12876), .B(n12877), .ZN(n12642) );
  XNOR2_X1 U12910 ( .A(n12878), .B(n12879), .ZN(n12876) );
  NOR2_X1 U12911 ( .A1(n8371), .A2(n12609), .ZN(n12879) );
  XNOR2_X1 U12912 ( .A(n12880), .B(n12881), .ZN(n12654) );
  XOR2_X1 U12913 ( .A(n12882), .B(n12883), .Z(n12881) );
  XOR2_X1 U12914 ( .A(n12884), .B(n12885), .Z(n12658) );
  XOR2_X1 U12915 ( .A(n12886), .B(n12887), .Z(n12884) );
  XNOR2_X1 U12916 ( .A(n12888), .B(n12889), .ZN(n12504) );
  XOR2_X1 U12917 ( .A(n12890), .B(n12891), .Z(n12888) );
  XOR2_X1 U12918 ( .A(n12892), .B(n12893), .Z(n12662) );
  XOR2_X1 U12919 ( .A(n12894), .B(n12895), .Z(n12892) );
  XOR2_X1 U12920 ( .A(n12896), .B(n12897), .Z(n12492) );
  XOR2_X1 U12921 ( .A(n12898), .B(n12899), .Z(n12896) );
  XNOR2_X1 U12922 ( .A(n12900), .B(n12901), .ZN(n12483) );
  XOR2_X1 U12923 ( .A(n12902), .B(n12903), .Z(n12901) );
  XOR2_X1 U12924 ( .A(n12904), .B(n12905), .Z(n12476) );
  XOR2_X1 U12925 ( .A(n12906), .B(n12907), .Z(n12904) );
  XOR2_X1 U12926 ( .A(n12908), .B(n12909), .Z(n12666) );
  XNOR2_X1 U12927 ( .A(n12910), .B(n12911), .ZN(n12908) );
  XOR2_X1 U12928 ( .A(n12912), .B(n12913), .Z(n12671) );
  XOR2_X1 U12929 ( .A(n12914), .B(n12915), .Z(n12912) );
  XNOR2_X1 U12930 ( .A(n12916), .B(n12917), .ZN(n12459) );
  XOR2_X1 U12931 ( .A(n12918), .B(n12919), .Z(n12917) );
  XNOR2_X1 U12932 ( .A(n12920), .B(n12921), .ZN(n12451) );
  XNOR2_X1 U12933 ( .A(n12922), .B(n12923), .ZN(n12921) );
  XOR2_X1 U12934 ( .A(n12924), .B(n12925), .Z(n12674) );
  XNOR2_X1 U12935 ( .A(n12926), .B(n12927), .ZN(n12925) );
  XNOR2_X1 U12936 ( .A(n12928), .B(n12929), .ZN(n12679) );
  XNOR2_X1 U12937 ( .A(n12930), .B(n12931), .ZN(n12929) );
  XNOR2_X1 U12938 ( .A(n12932), .B(n12933), .ZN(n8536) );
  NAND2_X1 U12939 ( .A1(n8544), .A2(n8543), .ZN(n8542) );
  NOR2_X1 U12940 ( .A1(n12934), .A2(n8588), .ZN(n8543) );
  INV_X1 U12941 ( .A(n12935), .ZN(n12934) );
  NAND2_X1 U12942 ( .A1(n12936), .A2(n12937), .ZN(n12935) );
  XNOR2_X1 U12943 ( .A(n12938), .B(n12939), .ZN(n12937) );
  NOR2_X1 U12944 ( .A1(n12933), .A2(n12932), .ZN(n8544) );
  XOR2_X1 U12945 ( .A(n12940), .B(n12941), .Z(n12932) );
  XNOR2_X1 U12946 ( .A(n12942), .B(n12943), .ZN(n12940) );
  NOR2_X1 U12947 ( .A1(n8457), .A2(n12835), .ZN(n12943) );
  NAND2_X1 U12948 ( .A1(n12944), .A2(n12945), .ZN(n12933) );
  NAND2_X1 U12949 ( .A1(n12928), .A2(n12946), .ZN(n12945) );
  NAND2_X1 U12950 ( .A1(n12931), .A2(n12930), .ZN(n12946) );
  XOR2_X1 U12951 ( .A(n12947), .B(n12948), .Z(n12928) );
  XOR2_X1 U12952 ( .A(n12949), .B(n12950), .Z(n12948) );
  NAND2_X1 U12953 ( .A1(b_13_), .A2(a_1_), .ZN(n12950) );
  INV_X1 U12954 ( .A(n12951), .ZN(n12944) );
  NOR2_X1 U12955 ( .A1(n12930), .A2(n12931), .ZN(n12951) );
  NOR2_X1 U12956 ( .A1(n12609), .A2(n8457), .ZN(n12931) );
  NAND2_X1 U12957 ( .A1(n12952), .A2(n12953), .ZN(n12930) );
  NAND2_X1 U12958 ( .A1(n12691), .A2(n12954), .ZN(n12953) );
  INV_X1 U12959 ( .A(n12955), .ZN(n12954) );
  NOR2_X1 U12960 ( .A1(n12688), .A2(n12690), .ZN(n12955) );
  NOR2_X1 U12961 ( .A1(n12609), .A2(n8569), .ZN(n12691) );
  NAND2_X1 U12962 ( .A1(n12688), .A2(n12690), .ZN(n12952) );
  NOR2_X1 U12963 ( .A1(n12956), .A2(n12957), .ZN(n12690) );
  INV_X1 U12964 ( .A(n12958), .ZN(n12957) );
  NAND2_X1 U12965 ( .A1(n12695), .A2(n12959), .ZN(n12958) );
  NAND2_X1 U12966 ( .A1(n12698), .A2(n12697), .ZN(n12959) );
  XNOR2_X1 U12967 ( .A(n12960), .B(n12961), .ZN(n12695) );
  XNOR2_X1 U12968 ( .A(n12962), .B(n12963), .ZN(n12961) );
  NAND2_X1 U12969 ( .A1(b_13_), .A2(a_3_), .ZN(n12963) );
  NOR2_X1 U12970 ( .A1(n12697), .A2(n12698), .ZN(n12956) );
  NOR2_X1 U12971 ( .A1(n12609), .A2(n8448), .ZN(n12698) );
  NAND2_X1 U12972 ( .A1(n12964), .A2(n12965), .ZN(n12697) );
  NAND2_X1 U12973 ( .A1(n12927), .A2(n12966), .ZN(n12965) );
  NAND2_X1 U12974 ( .A1(n12924), .A2(n12926), .ZN(n12966) );
  NOR2_X1 U12975 ( .A1(n12609), .A2(n8900), .ZN(n12927) );
  INV_X1 U12976 ( .A(n12967), .ZN(n12964) );
  NOR2_X1 U12977 ( .A1(n12926), .A2(n12924), .ZN(n12967) );
  XOR2_X1 U12978 ( .A(n12968), .B(n12969), .Z(n12924) );
  XNOR2_X1 U12979 ( .A(n12970), .B(n12971), .ZN(n12968) );
  NOR2_X1 U12980 ( .A1(n8439), .A2(n12835), .ZN(n12971) );
  NAND2_X1 U12981 ( .A1(n12972), .A2(n12973), .ZN(n12926) );
  NAND2_X1 U12982 ( .A1(n12920), .A2(n12974), .ZN(n12973) );
  NAND2_X1 U12983 ( .A1(n12923), .A2(n12922), .ZN(n12974) );
  XOR2_X1 U12984 ( .A(n12975), .B(n12976), .Z(n12920) );
  XNOR2_X1 U12985 ( .A(n12977), .B(n12978), .ZN(n12975) );
  NOR2_X1 U12986 ( .A1(n8938), .A2(n12835), .ZN(n12978) );
  INV_X1 U12987 ( .A(n12979), .ZN(n12972) );
  NOR2_X1 U12988 ( .A1(n12922), .A2(n12923), .ZN(n12979) );
  NOR2_X1 U12989 ( .A1(n12609), .A2(n8439), .ZN(n12923) );
  NAND2_X1 U12990 ( .A1(n12980), .A2(n12981), .ZN(n12922) );
  NAND2_X1 U12991 ( .A1(n12919), .A2(n12982), .ZN(n12981) );
  INV_X1 U12992 ( .A(n12983), .ZN(n12982) );
  NOR2_X1 U12993 ( .A1(n12916), .A2(n12918), .ZN(n12983) );
  NOR2_X1 U12994 ( .A1(n12609), .A2(n8938), .ZN(n12919) );
  NAND2_X1 U12995 ( .A1(n12916), .A2(n12918), .ZN(n12980) );
  NOR2_X1 U12996 ( .A1(n12984), .A2(n12985), .ZN(n12918) );
  INV_X1 U12997 ( .A(n12986), .ZN(n12985) );
  NAND2_X1 U12998 ( .A1(n12913), .A2(n12987), .ZN(n12986) );
  NAND2_X1 U12999 ( .A1(n12915), .A2(n12914), .ZN(n12987) );
  XOR2_X1 U13000 ( .A(n12988), .B(n12989), .Z(n12913) );
  XOR2_X1 U13001 ( .A(n12990), .B(n12991), .Z(n12989) );
  NAND2_X1 U13002 ( .A1(b_13_), .A2(a_7_), .ZN(n12991) );
  NOR2_X1 U13003 ( .A1(n12914), .A2(n12915), .ZN(n12984) );
  NOR2_X1 U13004 ( .A1(n12609), .A2(n8430), .ZN(n12915) );
  NAND2_X1 U13005 ( .A1(n12992), .A2(n12993), .ZN(n12914) );
  NAND2_X1 U13006 ( .A1(n12911), .A2(n12994), .ZN(n12993) );
  INV_X1 U13007 ( .A(n12995), .ZN(n12994) );
  NOR2_X1 U13008 ( .A1(n12909), .A2(n12910), .ZN(n12995) );
  NOR2_X1 U13009 ( .A1(n12609), .A2(n8425), .ZN(n12911) );
  NAND2_X1 U13010 ( .A1(n12910), .A2(n12909), .ZN(n12992) );
  XOR2_X1 U13011 ( .A(n12996), .B(n12997), .Z(n12909) );
  XNOR2_X1 U13012 ( .A(n12998), .B(n12999), .ZN(n12997) );
  NAND2_X1 U13013 ( .A1(b_13_), .A2(a_8_), .ZN(n12999) );
  NOR2_X1 U13014 ( .A1(n13000), .A2(n13001), .ZN(n12910) );
  INV_X1 U13015 ( .A(n13002), .ZN(n13001) );
  NAND2_X1 U13016 ( .A1(n12905), .A2(n13003), .ZN(n13002) );
  NAND2_X1 U13017 ( .A1(n12907), .A2(n12906), .ZN(n13003) );
  XNOR2_X1 U13018 ( .A(n13004), .B(n13005), .ZN(n12905) );
  XNOR2_X1 U13019 ( .A(n13006), .B(n13007), .ZN(n13005) );
  NAND2_X1 U13020 ( .A1(b_13_), .A2(a_9_), .ZN(n13007) );
  NOR2_X1 U13021 ( .A1(n12906), .A2(n12907), .ZN(n13000) );
  NOR2_X1 U13022 ( .A1(n12609), .A2(n8968), .ZN(n12907) );
  NAND2_X1 U13023 ( .A1(n13008), .A2(n13009), .ZN(n12906) );
  NAND2_X1 U13024 ( .A1(n12903), .A2(n13010), .ZN(n13009) );
  INV_X1 U13025 ( .A(n13011), .ZN(n13010) );
  NOR2_X1 U13026 ( .A1(n12900), .A2(n12902), .ZN(n13011) );
  NOR2_X1 U13027 ( .A1(n12609), .A2(n8971), .ZN(n12903) );
  NAND2_X1 U13028 ( .A1(n12900), .A2(n12902), .ZN(n13008) );
  NOR2_X1 U13029 ( .A1(n13012), .A2(n13013), .ZN(n12902) );
  INV_X1 U13030 ( .A(n13014), .ZN(n13013) );
  NAND2_X1 U13031 ( .A1(n12897), .A2(n13015), .ZN(n13014) );
  NAND2_X1 U13032 ( .A1(n12899), .A2(n12898), .ZN(n13015) );
  XOR2_X1 U13033 ( .A(n13016), .B(n13017), .Z(n12897) );
  XNOR2_X1 U13034 ( .A(n13018), .B(n13019), .ZN(n13016) );
  NOR2_X1 U13035 ( .A1(n8867), .A2(n12835), .ZN(n13019) );
  NOR2_X1 U13036 ( .A1(n12898), .A2(n12899), .ZN(n13012) );
  NOR2_X1 U13037 ( .A1(n12609), .A2(n8402), .ZN(n12899) );
  NAND2_X1 U13038 ( .A1(n13020), .A2(n13021), .ZN(n12898) );
  NAND2_X1 U13039 ( .A1(n12895), .A2(n13022), .ZN(n13021) );
  NAND2_X1 U13040 ( .A1(n12893), .A2(n12894), .ZN(n13022) );
  NOR2_X1 U13041 ( .A1(n12609), .A2(n8867), .ZN(n12895) );
  INV_X1 U13042 ( .A(n13023), .ZN(n13020) );
  NOR2_X1 U13043 ( .A1(n12893), .A2(n12894), .ZN(n13023) );
  NAND2_X1 U13044 ( .A1(n13024), .A2(n13025), .ZN(n12894) );
  NAND2_X1 U13045 ( .A1(n12889), .A2(n13026), .ZN(n13025) );
  NAND2_X1 U13046 ( .A1(n12891), .A2(n12890), .ZN(n13026) );
  XOR2_X1 U13047 ( .A(n13027), .B(n13028), .Z(n12889) );
  XNOR2_X1 U13048 ( .A(n13029), .B(n13030), .ZN(n13027) );
  INV_X1 U13049 ( .A(n13031), .ZN(n13024) );
  NOR2_X1 U13050 ( .A1(n12890), .A2(n12891), .ZN(n13031) );
  NOR2_X1 U13051 ( .A1(n12609), .A2(n8393), .ZN(n12891) );
  NAND2_X1 U13052 ( .A1(n13032), .A2(n13033), .ZN(n12890) );
  NAND2_X1 U13053 ( .A1(n12887), .A2(n13034), .ZN(n13033) );
  NAND2_X1 U13054 ( .A1(n12885), .A2(n12886), .ZN(n13034) );
  NOR2_X1 U13055 ( .A1(n12609), .A2(n8996), .ZN(n12887) );
  INV_X1 U13056 ( .A(n13035), .ZN(n13032) );
  NOR2_X1 U13057 ( .A1(n12885), .A2(n12886), .ZN(n13035) );
  NAND2_X1 U13058 ( .A1(n13036), .A2(n13037), .ZN(n12886) );
  NAND2_X1 U13059 ( .A1(n13038), .A2(n12882), .ZN(n13037) );
  NAND2_X1 U13060 ( .A1(n12880), .A2(n12883), .ZN(n13038) );
  INV_X1 U13061 ( .A(n13039), .ZN(n13036) );
  NOR2_X1 U13062 ( .A1(n12883), .A2(n12880), .ZN(n13039) );
  XNOR2_X1 U13063 ( .A(n13040), .B(n13041), .ZN(n12880) );
  XOR2_X1 U13064 ( .A(n13042), .B(n13043), .Z(n13041) );
  NAND2_X1 U13065 ( .A1(b_13_), .A2(a_15_), .ZN(n13043) );
  NAND2_X1 U13066 ( .A1(n13044), .A2(n13045), .ZN(n12883) );
  NAND2_X1 U13067 ( .A1(n12754), .A2(n13046), .ZN(n13045) );
  NAND2_X1 U13068 ( .A1(n12753), .A2(n12751), .ZN(n13046) );
  NOR2_X1 U13069 ( .A1(n12609), .A2(n8850), .ZN(n12754) );
  INV_X1 U13070 ( .A(n13047), .ZN(n13044) );
  NOR2_X1 U13071 ( .A1(n12751), .A2(n12753), .ZN(n13047) );
  NOR2_X1 U13072 ( .A1(n13048), .A2(n13049), .ZN(n12753) );
  NOR3_X1 U13073 ( .A1(n8376), .A2(n13050), .A3(n12609), .ZN(n13049) );
  INV_X1 U13074 ( .A(n13051), .ZN(n13050) );
  NAND2_X1 U13075 ( .A1(n12762), .A2(n12761), .ZN(n13051) );
  NOR2_X1 U13076 ( .A1(n12761), .A2(n12762), .ZN(n13048) );
  NOR2_X1 U13077 ( .A1(n13052), .A2(n13053), .ZN(n12762) );
  INV_X1 U13078 ( .A(n13054), .ZN(n13053) );
  NAND3_X1 U13079 ( .A1(a_17_), .A2(n13055), .A3(b_14_), .ZN(n13054) );
  NAND2_X1 U13080 ( .A1(n12878), .A2(n12877), .ZN(n13055) );
  NOR2_X1 U13081 ( .A1(n12877), .A2(n12878), .ZN(n13052) );
  NOR2_X1 U13082 ( .A1(n13056), .A2(n13057), .ZN(n12878) );
  NOR3_X1 U13083 ( .A1(n9291), .A2(n13058), .A3(n12609), .ZN(n13057) );
  NOR2_X1 U13084 ( .A1(n12872), .A2(n12874), .ZN(n13058) );
  INV_X1 U13085 ( .A(n13059), .ZN(n13056) );
  NAND2_X1 U13086 ( .A1(n12872), .A2(n12874), .ZN(n13059) );
  NAND2_X1 U13087 ( .A1(n13060), .A2(n13061), .ZN(n12874) );
  NAND3_X1 U13088 ( .A1(a_19_), .A2(n13062), .A3(b_14_), .ZN(n13061) );
  NAND2_X1 U13089 ( .A1(n12870), .A2(n12868), .ZN(n13062) );
  INV_X1 U13090 ( .A(n13063), .ZN(n13060) );
  NOR2_X1 U13091 ( .A1(n12868), .A2(n12870), .ZN(n13063) );
  NOR2_X1 U13092 ( .A1(n13064), .A2(n13065), .ZN(n12870) );
  INV_X1 U13093 ( .A(n13066), .ZN(n13065) );
  NAND3_X1 U13094 ( .A1(a_20_), .A2(n13067), .A3(b_14_), .ZN(n13066) );
  NAND2_X1 U13095 ( .A1(n12865), .A2(n12866), .ZN(n13067) );
  NOR2_X1 U13096 ( .A1(n12865), .A2(n12866), .ZN(n13064) );
  NOR2_X1 U13097 ( .A1(n13068), .A2(n13069), .ZN(n12866) );
  NOR3_X1 U13098 ( .A1(n8759), .A2(n13070), .A3(n12609), .ZN(n13069) );
  NOR2_X1 U13099 ( .A1(n12862), .A2(n12861), .ZN(n13070) );
  INV_X1 U13100 ( .A(n13071), .ZN(n13068) );
  NAND2_X1 U13101 ( .A1(n12861), .A2(n12862), .ZN(n13071) );
  NAND2_X1 U13102 ( .A1(n13072), .A2(n13073), .ZN(n12862) );
  NAND2_X1 U13103 ( .A1(n12859), .A2(n13074), .ZN(n13073) );
  INV_X1 U13104 ( .A(n13075), .ZN(n13074) );
  NOR2_X1 U13105 ( .A1(n12856), .A2(n12858), .ZN(n13075) );
  NOR2_X1 U13106 ( .A1(n12609), .A2(n12296), .ZN(n12859) );
  NAND2_X1 U13107 ( .A1(n12856), .A2(n12858), .ZN(n13072) );
  NAND2_X1 U13108 ( .A1(n13076), .A2(n13077), .ZN(n12858) );
  NAND2_X1 U13109 ( .A1(n12855), .A2(n13078), .ZN(n13077) );
  INV_X1 U13110 ( .A(n13079), .ZN(n13078) );
  NOR2_X1 U13111 ( .A1(n12854), .A2(n12853), .ZN(n13079) );
  NOR2_X1 U13112 ( .A1(n12609), .A2(n12301), .ZN(n12855) );
  NAND2_X1 U13113 ( .A1(n12853), .A2(n12854), .ZN(n13076) );
  NAND2_X1 U13114 ( .A1(n13080), .A2(n13081), .ZN(n12854) );
  NAND2_X1 U13115 ( .A1(n12851), .A2(n13082), .ZN(n13081) );
  INV_X1 U13116 ( .A(n13083), .ZN(n13082) );
  NOR2_X1 U13117 ( .A1(n12849), .A2(n12850), .ZN(n13083) );
  NOR2_X1 U13118 ( .A1(n12609), .A2(n8779), .ZN(n12851) );
  NAND2_X1 U13119 ( .A1(n12849), .A2(n12850), .ZN(n13080) );
  NAND2_X1 U13120 ( .A1(n13084), .A2(n13085), .ZN(n12850) );
  NAND2_X1 U13121 ( .A1(n12847), .A2(n13086), .ZN(n13085) );
  NAND2_X1 U13122 ( .A1(n12844), .A2(n12846), .ZN(n13086) );
  NOR2_X1 U13123 ( .A1(n12609), .A2(n8788), .ZN(n12847) );
  INV_X1 U13124 ( .A(n13087), .ZN(n13084) );
  NOR2_X1 U13125 ( .A1(n12846), .A2(n12844), .ZN(n13087) );
  XNOR2_X1 U13126 ( .A(n13088), .B(n13089), .ZN(n12844) );
  XNOR2_X1 U13127 ( .A(n13090), .B(n13091), .ZN(n13089) );
  NAND2_X1 U13128 ( .A1(n13092), .A2(n13093), .ZN(n12846) );
  NAND2_X1 U13129 ( .A1(n12805), .A2(n13094), .ZN(n13093) );
  NAND2_X1 U13130 ( .A1(n12808), .A2(n12807), .ZN(n13094) );
  XNOR2_X1 U13131 ( .A(n13095), .B(n13096), .ZN(n12805) );
  XOR2_X1 U13132 ( .A(n13097), .B(n13098), .Z(n13095) );
  INV_X1 U13133 ( .A(n13099), .ZN(n13092) );
  NOR2_X1 U13134 ( .A1(n12807), .A2(n12808), .ZN(n13099) );
  NOR2_X1 U13135 ( .A1(n12609), .A2(n9344), .ZN(n12808) );
  NAND2_X1 U13136 ( .A1(n13100), .A2(n13101), .ZN(n12807) );
  NAND2_X1 U13137 ( .A1(n12815), .A2(n13102), .ZN(n13101) );
  INV_X1 U13138 ( .A(n13103), .ZN(n13102) );
  NOR2_X1 U13139 ( .A1(n12813), .A2(n12814), .ZN(n13103) );
  NOR2_X1 U13140 ( .A1(n12609), .A2(n8797), .ZN(n12815) );
  NAND2_X1 U13141 ( .A1(n12813), .A2(n12814), .ZN(n13100) );
  NAND2_X1 U13142 ( .A1(n13104), .A2(n13105), .ZN(n12814) );
  NAND2_X1 U13143 ( .A1(n12842), .A2(n13106), .ZN(n13105) );
  INV_X1 U13144 ( .A(n13107), .ZN(n13106) );
  NOR2_X1 U13145 ( .A1(n12843), .A2(n12841), .ZN(n13107) );
  NOR2_X1 U13146 ( .A1(n12609), .A2(n8314), .ZN(n12842) );
  NAND2_X1 U13147 ( .A1(n12841), .A2(n12843), .ZN(n13104) );
  NAND2_X1 U13148 ( .A1(n13108), .A2(n13109), .ZN(n12843) );
  NAND2_X1 U13149 ( .A1(n12837), .A2(n13110), .ZN(n13109) );
  INV_X1 U13150 ( .A(n13111), .ZN(n13110) );
  NOR2_X1 U13151 ( .A1(n12838), .A2(n12839), .ZN(n13111) );
  NOR2_X1 U13152 ( .A1(n12609), .A2(n9098), .ZN(n12837) );
  NAND2_X1 U13153 ( .A1(n12839), .A2(n12838), .ZN(n13108) );
  NAND2_X1 U13154 ( .A1(n13112), .A2(n13113), .ZN(n12838) );
  NAND2_X1 U13155 ( .A1(b_12_), .A2(n13114), .ZN(n13113) );
  NAND2_X1 U13156 ( .A1(n8299), .A2(n13115), .ZN(n13114) );
  NAND2_X1 U13157 ( .A1(a_31_), .A2(n12835), .ZN(n13115) );
  NAND2_X1 U13158 ( .A1(b_13_), .A2(n13116), .ZN(n13112) );
  NAND2_X1 U13159 ( .A1(n8303), .A2(n13117), .ZN(n13116) );
  NAND2_X1 U13160 ( .A1(a_30_), .A2(n13118), .ZN(n13117) );
  NOR3_X1 U13161 ( .A1(n12835), .A2(n9631), .A3(n12609), .ZN(n12839) );
  XOR2_X1 U13162 ( .A(n13119), .B(n13120), .Z(n12841) );
  XOR2_X1 U13163 ( .A(n13121), .B(n13122), .Z(n13119) );
  XOR2_X1 U13164 ( .A(n13123), .B(n13124), .Z(n12813) );
  XOR2_X1 U13165 ( .A(n13125), .B(n13126), .Z(n13123) );
  XNOR2_X1 U13166 ( .A(n13127), .B(n13128), .ZN(n12849) );
  XNOR2_X1 U13167 ( .A(n13129), .B(n13130), .ZN(n13128) );
  XOR2_X1 U13168 ( .A(n13131), .B(n13132), .Z(n12853) );
  XOR2_X1 U13169 ( .A(n13133), .B(n13134), .Z(n13131) );
  XOR2_X1 U13170 ( .A(n13135), .B(n13136), .Z(n12856) );
  XOR2_X1 U13171 ( .A(n13137), .B(n13138), .Z(n13135) );
  XNOR2_X1 U13172 ( .A(n13139), .B(n13140), .ZN(n12861) );
  XNOR2_X1 U13173 ( .A(n13141), .B(n13142), .ZN(n13140) );
  XNOR2_X1 U13174 ( .A(n13143), .B(n13144), .ZN(n12865) );
  XOR2_X1 U13175 ( .A(n13145), .B(n13146), .Z(n13143) );
  NOR2_X1 U13176 ( .A1(n8759), .A2(n12835), .ZN(n13146) );
  XOR2_X1 U13177 ( .A(n13147), .B(n13148), .Z(n12868) );
  XNOR2_X1 U13178 ( .A(n13149), .B(n13150), .ZN(n13147) );
  NOR2_X1 U13179 ( .A1(n9047), .A2(n12835), .ZN(n13150) );
  XOR2_X1 U13180 ( .A(n13151), .B(n13152), .Z(n12872) );
  XNOR2_X1 U13181 ( .A(n13153), .B(n13154), .ZN(n13152) );
  NAND2_X1 U13182 ( .A1(b_13_), .A2(a_19_), .ZN(n13154) );
  XOR2_X1 U13183 ( .A(n13155), .B(n13156), .Z(n12877) );
  XOR2_X1 U13184 ( .A(n13157), .B(n13158), .Z(n13156) );
  XNOR2_X1 U13185 ( .A(n13159), .B(n13160), .ZN(n12761) );
  XNOR2_X1 U13186 ( .A(n13161), .B(n13162), .ZN(n13159) );
  XNOR2_X1 U13187 ( .A(n13163), .B(n13164), .ZN(n12751) );
  XOR2_X1 U13188 ( .A(n13165), .B(n13166), .Z(n13163) );
  NOR2_X1 U13189 ( .A1(n8376), .A2(n12835), .ZN(n13166) );
  XOR2_X1 U13190 ( .A(n13167), .B(n13168), .Z(n12885) );
  XOR2_X1 U13191 ( .A(n13169), .B(n13170), .Z(n13168) );
  NAND2_X1 U13192 ( .A1(b_13_), .A2(a_14_), .ZN(n13170) );
  XOR2_X1 U13193 ( .A(n13171), .B(n13172), .Z(n12893) );
  XOR2_X1 U13194 ( .A(n13173), .B(n13174), .Z(n13172) );
  NAND2_X1 U13195 ( .A1(b_13_), .A2(a_12_), .ZN(n13174) );
  XOR2_X1 U13196 ( .A(n13175), .B(n13176), .Z(n12900) );
  XNOR2_X1 U13197 ( .A(n13177), .B(n13178), .ZN(n13176) );
  NAND2_X1 U13198 ( .A1(b_13_), .A2(a_10_), .ZN(n13178) );
  XOR2_X1 U13199 ( .A(n13179), .B(n13180), .Z(n12916) );
  XNOR2_X1 U13200 ( .A(n13181), .B(n13182), .ZN(n13180) );
  NAND2_X1 U13201 ( .A1(b_13_), .A2(a_6_), .ZN(n13182) );
  XNOR2_X1 U13202 ( .A(n13183), .B(n13184), .ZN(n12688) );
  XNOR2_X1 U13203 ( .A(n13185), .B(n13186), .ZN(n13183) );
  NOR2_X1 U13204 ( .A1(n8448), .A2(n12835), .ZN(n13186) );
  NOR2_X1 U13205 ( .A1(n13187), .A2(n12936), .ZN(n8588) );
  NOR2_X1 U13206 ( .A1(n13188), .A2(n13189), .ZN(n12936) );
  INV_X1 U13207 ( .A(n13190), .ZN(n13189) );
  NAND3_X1 U13208 ( .A1(a_0_), .A2(n13191), .A3(b_13_), .ZN(n13190) );
  NAND2_X1 U13209 ( .A1(n12942), .A2(n12941), .ZN(n13191) );
  NOR2_X1 U13210 ( .A1(n12941), .A2(n12942), .ZN(n13188) );
  NOR2_X1 U13211 ( .A1(n13192), .A2(n13193), .ZN(n12942) );
  NOR3_X1 U13212 ( .A1(n8569), .A2(n13194), .A3(n12835), .ZN(n13193) );
  NOR2_X1 U13213 ( .A1(n12949), .A2(n12947), .ZN(n13194) );
  INV_X1 U13214 ( .A(n13195), .ZN(n13192) );
  NAND2_X1 U13215 ( .A1(n12947), .A2(n12949), .ZN(n13195) );
  NAND2_X1 U13216 ( .A1(n13196), .A2(n13197), .ZN(n12949) );
  NAND3_X1 U13217 ( .A1(a_2_), .A2(n13198), .A3(b_13_), .ZN(n13197) );
  NAND2_X1 U13218 ( .A1(n13185), .A2(n13184), .ZN(n13198) );
  INV_X1 U13219 ( .A(n13199), .ZN(n13196) );
  NOR2_X1 U13220 ( .A1(n13184), .A2(n13185), .ZN(n13199) );
  NOR2_X1 U13221 ( .A1(n13200), .A2(n13201), .ZN(n13185) );
  NOR3_X1 U13222 ( .A1(n8900), .A2(n13202), .A3(n12835), .ZN(n13201) );
  INV_X1 U13223 ( .A(n13203), .ZN(n13202) );
  NAND2_X1 U13224 ( .A1(n12962), .A2(n12960), .ZN(n13203) );
  NOR2_X1 U13225 ( .A1(n12960), .A2(n12962), .ZN(n13200) );
  NOR2_X1 U13226 ( .A1(n13204), .A2(n13205), .ZN(n12962) );
  INV_X1 U13227 ( .A(n13206), .ZN(n13205) );
  NAND3_X1 U13228 ( .A1(a_4_), .A2(n13207), .A3(b_13_), .ZN(n13206) );
  NAND2_X1 U13229 ( .A1(n12970), .A2(n12969), .ZN(n13207) );
  NOR2_X1 U13230 ( .A1(n12969), .A2(n12970), .ZN(n13204) );
  NOR2_X1 U13231 ( .A1(n13208), .A2(n13209), .ZN(n12970) );
  INV_X1 U13232 ( .A(n13210), .ZN(n13209) );
  NAND3_X1 U13233 ( .A1(a_5_), .A2(n13211), .A3(b_13_), .ZN(n13210) );
  NAND2_X1 U13234 ( .A1(n12977), .A2(n12976), .ZN(n13211) );
  NOR2_X1 U13235 ( .A1(n12976), .A2(n12977), .ZN(n13208) );
  NOR2_X1 U13236 ( .A1(n13212), .A2(n13213), .ZN(n12977) );
  NOR3_X1 U13237 ( .A1(n8430), .A2(n13214), .A3(n12835), .ZN(n13213) );
  INV_X1 U13238 ( .A(n13215), .ZN(n13214) );
  NAND2_X1 U13239 ( .A1(n13181), .A2(n13179), .ZN(n13215) );
  NOR2_X1 U13240 ( .A1(n13179), .A2(n13181), .ZN(n13212) );
  NOR2_X1 U13241 ( .A1(n13216), .A2(n13217), .ZN(n13181) );
  NOR3_X1 U13242 ( .A1(n8425), .A2(n13218), .A3(n12835), .ZN(n13217) );
  NOR2_X1 U13243 ( .A1(n12990), .A2(n12988), .ZN(n13218) );
  INV_X1 U13244 ( .A(n13219), .ZN(n13216) );
  NAND2_X1 U13245 ( .A1(n12988), .A2(n12990), .ZN(n13219) );
  NAND2_X1 U13246 ( .A1(n13220), .A2(n13221), .ZN(n12990) );
  NAND3_X1 U13247 ( .A1(a_8_), .A2(n13222), .A3(b_13_), .ZN(n13221) );
  NAND2_X1 U13248 ( .A1(n12998), .A2(n12996), .ZN(n13222) );
  INV_X1 U13249 ( .A(n13223), .ZN(n13220) );
  NOR2_X1 U13250 ( .A1(n12996), .A2(n12998), .ZN(n13223) );
  NOR2_X1 U13251 ( .A1(n13224), .A2(n13225), .ZN(n12998) );
  NOR3_X1 U13252 ( .A1(n8971), .A2(n13226), .A3(n12835), .ZN(n13225) );
  INV_X1 U13253 ( .A(n13227), .ZN(n13226) );
  NAND2_X1 U13254 ( .A1(n13006), .A2(n13004), .ZN(n13227) );
  NOR2_X1 U13255 ( .A1(n13004), .A2(n13006), .ZN(n13224) );
  NOR2_X1 U13256 ( .A1(n13228), .A2(n13229), .ZN(n13006) );
  INV_X1 U13257 ( .A(n13230), .ZN(n13229) );
  NAND3_X1 U13258 ( .A1(a_10_), .A2(n13231), .A3(b_13_), .ZN(n13230) );
  NAND2_X1 U13259 ( .A1(n13177), .A2(n13175), .ZN(n13231) );
  NOR2_X1 U13260 ( .A1(n13175), .A2(n13177), .ZN(n13228) );
  NOR2_X1 U13261 ( .A1(n13232), .A2(n13233), .ZN(n13177) );
  INV_X1 U13262 ( .A(n13234), .ZN(n13233) );
  NAND3_X1 U13263 ( .A1(a_11_), .A2(n13235), .A3(b_13_), .ZN(n13234) );
  NAND2_X1 U13264 ( .A1(n13018), .A2(n13017), .ZN(n13235) );
  NOR2_X1 U13265 ( .A1(n13017), .A2(n13018), .ZN(n13232) );
  NOR2_X1 U13266 ( .A1(n13236), .A2(n13237), .ZN(n13018) );
  INV_X1 U13267 ( .A(n13238), .ZN(n13237) );
  NAND3_X1 U13268 ( .A1(a_12_), .A2(n13239), .A3(b_13_), .ZN(n13238) );
  NAND2_X1 U13269 ( .A1(n13171), .A2(n13173), .ZN(n13239) );
  NOR2_X1 U13270 ( .A1(n13173), .A2(n13171), .ZN(n13236) );
  XOR2_X1 U13271 ( .A(n13240), .B(n13241), .Z(n13171) );
  NAND2_X1 U13272 ( .A1(n13242), .A2(n13243), .ZN(n13240) );
  NAND2_X1 U13273 ( .A1(n13244), .A2(n13245), .ZN(n13173) );
  NAND2_X1 U13274 ( .A1(n13028), .A2(n13246), .ZN(n13245) );
  NAND2_X1 U13275 ( .A1(n13030), .A2(n13247), .ZN(n13246) );
  INV_X1 U13276 ( .A(n13029), .ZN(n13247) );
  XOR2_X1 U13277 ( .A(n13248), .B(n13249), .Z(n13028) );
  NAND2_X1 U13278 ( .A1(n13250), .A2(n13251), .ZN(n13248) );
  NAND2_X1 U13279 ( .A1(n13029), .A2(n13252), .ZN(n13244) );
  NOR2_X1 U13280 ( .A1(n13253), .A2(n13254), .ZN(n13029) );
  NOR3_X1 U13281 ( .A1(n9262), .A2(n13255), .A3(n12835), .ZN(n13254) );
  NOR2_X1 U13282 ( .A1(n13169), .A2(n13167), .ZN(n13255) );
  INV_X1 U13283 ( .A(n13256), .ZN(n13253) );
  NAND2_X1 U13284 ( .A1(n13167), .A2(n13169), .ZN(n13256) );
  NAND2_X1 U13285 ( .A1(n13257), .A2(n13258), .ZN(n13169) );
  INV_X1 U13286 ( .A(n13259), .ZN(n13258) );
  NOR3_X1 U13287 ( .A1(n8850), .A2(n13260), .A3(n12835), .ZN(n13259) );
  NOR2_X1 U13288 ( .A1(n13042), .A2(n13040), .ZN(n13260) );
  NAND2_X1 U13289 ( .A1(n13040), .A2(n13042), .ZN(n13257) );
  NAND2_X1 U13290 ( .A1(n13261), .A2(n13262), .ZN(n13042) );
  NAND3_X1 U13291 ( .A1(a_16_), .A2(n13263), .A3(b_13_), .ZN(n13262) );
  INV_X1 U13292 ( .A(n13264), .ZN(n13263) );
  NOR2_X1 U13293 ( .A1(n13165), .A2(n13164), .ZN(n13264) );
  NAND2_X1 U13294 ( .A1(n13164), .A2(n13165), .ZN(n13261) );
  NAND2_X1 U13295 ( .A1(n13265), .A2(n13266), .ZN(n13165) );
  NAND2_X1 U13296 ( .A1(n13162), .A2(n13267), .ZN(n13266) );
  NAND2_X1 U13297 ( .A1(n13161), .A2(n13268), .ZN(n13267) );
  INV_X1 U13298 ( .A(n13160), .ZN(n13268) );
  NOR2_X1 U13299 ( .A1(n12835), .A2(n8371), .ZN(n13162) );
  NAND2_X1 U13300 ( .A1(n13160), .A2(n13269), .ZN(n13265) );
  INV_X1 U13301 ( .A(n13161), .ZN(n13269) );
  NOR2_X1 U13302 ( .A1(n13270), .A2(n13271), .ZN(n13161) );
  NOR2_X1 U13303 ( .A1(n13158), .A2(n13272), .ZN(n13271) );
  NOR2_X1 U13304 ( .A1(n13157), .A2(n13155), .ZN(n13272) );
  NAND2_X1 U13305 ( .A1(b_13_), .A2(a_18_), .ZN(n13158) );
  INV_X1 U13306 ( .A(n13273), .ZN(n13270) );
  NAND2_X1 U13307 ( .A1(n13155), .A2(n13157), .ZN(n13273) );
  NAND2_X1 U13308 ( .A1(n13274), .A2(n13275), .ZN(n13157) );
  NAND3_X1 U13309 ( .A1(a_19_), .A2(n13276), .A3(b_13_), .ZN(n13275) );
  NAND2_X1 U13310 ( .A1(n13153), .A2(n13151), .ZN(n13276) );
  INV_X1 U13311 ( .A(n13277), .ZN(n13274) );
  NOR2_X1 U13312 ( .A1(n13151), .A2(n13153), .ZN(n13277) );
  NOR2_X1 U13313 ( .A1(n13278), .A2(n13279), .ZN(n13153) );
  INV_X1 U13314 ( .A(n13280), .ZN(n13279) );
  NAND3_X1 U13315 ( .A1(a_20_), .A2(n13281), .A3(b_13_), .ZN(n13280) );
  NAND2_X1 U13316 ( .A1(n13149), .A2(n13148), .ZN(n13281) );
  NOR2_X1 U13317 ( .A1(n13148), .A2(n13149), .ZN(n13278) );
  NOR2_X1 U13318 ( .A1(n13282), .A2(n13283), .ZN(n13149) );
  NOR3_X1 U13319 ( .A1(n8759), .A2(n13284), .A3(n12835), .ZN(n13283) );
  NOR2_X1 U13320 ( .A1(n13145), .A2(n13144), .ZN(n13284) );
  INV_X1 U13321 ( .A(n13285), .ZN(n13282) );
  NAND2_X1 U13322 ( .A1(n13144), .A2(n13145), .ZN(n13285) );
  NAND2_X1 U13323 ( .A1(n13286), .A2(n13287), .ZN(n13145) );
  NAND2_X1 U13324 ( .A1(n13142), .A2(n13288), .ZN(n13287) );
  INV_X1 U13325 ( .A(n13289), .ZN(n13288) );
  NOR2_X1 U13326 ( .A1(n13141), .A2(n13139), .ZN(n13289) );
  NOR2_X1 U13327 ( .A1(n12835), .A2(n12296), .ZN(n13142) );
  NAND2_X1 U13328 ( .A1(n13139), .A2(n13141), .ZN(n13286) );
  NAND2_X1 U13329 ( .A1(n13290), .A2(n13291), .ZN(n13141) );
  NAND2_X1 U13330 ( .A1(n13138), .A2(n13292), .ZN(n13291) );
  INV_X1 U13331 ( .A(n13293), .ZN(n13292) );
  NOR2_X1 U13332 ( .A1(n13137), .A2(n13136), .ZN(n13293) );
  NOR2_X1 U13333 ( .A1(n12835), .A2(n12301), .ZN(n13138) );
  NAND2_X1 U13334 ( .A1(n13136), .A2(n13137), .ZN(n13290) );
  NAND2_X1 U13335 ( .A1(n13294), .A2(n13295), .ZN(n13137) );
  NAND2_X1 U13336 ( .A1(n13134), .A2(n13296), .ZN(n13295) );
  INV_X1 U13337 ( .A(n13297), .ZN(n13296) );
  NOR2_X1 U13338 ( .A1(n13133), .A2(n13132), .ZN(n13297) );
  NOR2_X1 U13339 ( .A1(n12835), .A2(n8779), .ZN(n13134) );
  NAND2_X1 U13340 ( .A1(n13132), .A2(n13133), .ZN(n13294) );
  NAND2_X1 U13341 ( .A1(n13298), .A2(n13299), .ZN(n13133) );
  NAND2_X1 U13342 ( .A1(n13130), .A2(n13300), .ZN(n13299) );
  NAND2_X1 U13343 ( .A1(n13127), .A2(n13129), .ZN(n13300) );
  NOR2_X1 U13344 ( .A1(n12835), .A2(n8788), .ZN(n13130) );
  INV_X1 U13345 ( .A(n13301), .ZN(n13298) );
  NOR2_X1 U13346 ( .A1(n13129), .A2(n13127), .ZN(n13301) );
  XNOR2_X1 U13347 ( .A(n13302), .B(n13303), .ZN(n13127) );
  XNOR2_X1 U13348 ( .A(n13304), .B(n13305), .ZN(n13303) );
  NAND2_X1 U13349 ( .A1(n13306), .A2(n13307), .ZN(n13129) );
  NAND2_X1 U13350 ( .A1(n13088), .A2(n13308), .ZN(n13307) );
  NAND2_X1 U13351 ( .A1(n13091), .A2(n13090), .ZN(n13308) );
  XNOR2_X1 U13352 ( .A(n13309), .B(n13310), .ZN(n13088) );
  XOR2_X1 U13353 ( .A(n13311), .B(n13312), .Z(n13309) );
  INV_X1 U13354 ( .A(n13313), .ZN(n13306) );
  NOR2_X1 U13355 ( .A1(n13090), .A2(n13091), .ZN(n13313) );
  NOR2_X1 U13356 ( .A1(n12835), .A2(n9344), .ZN(n13091) );
  NAND2_X1 U13357 ( .A1(n13314), .A2(n13315), .ZN(n13090) );
  NAND2_X1 U13358 ( .A1(n13098), .A2(n13316), .ZN(n13315) );
  INV_X1 U13359 ( .A(n13317), .ZN(n13316) );
  NOR2_X1 U13360 ( .A1(n13097), .A2(n13096), .ZN(n13317) );
  NOR2_X1 U13361 ( .A1(n12835), .A2(n8797), .ZN(n13098) );
  NAND2_X1 U13362 ( .A1(n13096), .A2(n13097), .ZN(n13314) );
  NAND2_X1 U13363 ( .A1(n13318), .A2(n13319), .ZN(n13097) );
  NAND2_X1 U13364 ( .A1(n13125), .A2(n13320), .ZN(n13319) );
  INV_X1 U13365 ( .A(n13321), .ZN(n13320) );
  NOR2_X1 U13366 ( .A1(n13126), .A2(n13124), .ZN(n13321) );
  NOR2_X1 U13367 ( .A1(n12835), .A2(n8314), .ZN(n13125) );
  NAND2_X1 U13368 ( .A1(n13124), .A2(n13126), .ZN(n13318) );
  NAND2_X1 U13369 ( .A1(n13322), .A2(n13323), .ZN(n13126) );
  NAND2_X1 U13370 ( .A1(n13120), .A2(n13324), .ZN(n13323) );
  INV_X1 U13371 ( .A(n13325), .ZN(n13324) );
  NOR2_X1 U13372 ( .A1(n13121), .A2(n13122), .ZN(n13325) );
  NOR2_X1 U13373 ( .A1(n12835), .A2(n9098), .ZN(n13120) );
  NAND2_X1 U13374 ( .A1(n13122), .A2(n13121), .ZN(n13322) );
  NAND2_X1 U13375 ( .A1(n13326), .A2(n13327), .ZN(n13121) );
  NAND2_X1 U13376 ( .A1(b_11_), .A2(n13328), .ZN(n13327) );
  NAND2_X1 U13377 ( .A1(n8299), .A2(n13329), .ZN(n13328) );
  NAND2_X1 U13378 ( .A1(a_31_), .A2(n13118), .ZN(n13329) );
  NAND2_X1 U13379 ( .A1(b_12_), .A2(n13330), .ZN(n13326) );
  NAND2_X1 U13380 ( .A1(n8303), .A2(n13331), .ZN(n13330) );
  NAND2_X1 U13381 ( .A1(a_30_), .A2(n13332), .ZN(n13331) );
  NOR3_X1 U13382 ( .A1(n12835), .A2(n9631), .A3(n13118), .ZN(n13122) );
  XOR2_X1 U13383 ( .A(n13333), .B(n13334), .Z(n13124) );
  XOR2_X1 U13384 ( .A(n13335), .B(n13336), .Z(n13333) );
  XOR2_X1 U13385 ( .A(n13337), .B(n13338), .Z(n13096) );
  XOR2_X1 U13386 ( .A(n13339), .B(n13340), .Z(n13337) );
  XNOR2_X1 U13387 ( .A(n13341), .B(n13342), .ZN(n13132) );
  XNOR2_X1 U13388 ( .A(n13343), .B(n13344), .ZN(n13342) );
  XOR2_X1 U13389 ( .A(n13345), .B(n13346), .Z(n13136) );
  XOR2_X1 U13390 ( .A(n13347), .B(n13348), .Z(n13345) );
  XOR2_X1 U13391 ( .A(n13349), .B(n13350), .Z(n13139) );
  XOR2_X1 U13392 ( .A(n13351), .B(n13352), .Z(n13349) );
  XNOR2_X1 U13393 ( .A(n13353), .B(n13354), .ZN(n13144) );
  XNOR2_X1 U13394 ( .A(n13355), .B(n13356), .ZN(n13354) );
  XNOR2_X1 U13395 ( .A(n13357), .B(n13358), .ZN(n13148) );
  XOR2_X1 U13396 ( .A(n13359), .B(n13360), .Z(n13357) );
  NOR2_X1 U13397 ( .A1(n8759), .A2(n13118), .ZN(n13360) );
  XOR2_X1 U13398 ( .A(n13361), .B(n13362), .Z(n13151) );
  XNOR2_X1 U13399 ( .A(n13363), .B(n13364), .ZN(n13361) );
  NOR2_X1 U13400 ( .A1(n9047), .A2(n13118), .ZN(n13364) );
  XOR2_X1 U13401 ( .A(n13365), .B(n13366), .Z(n13155) );
  XNOR2_X1 U13402 ( .A(n13367), .B(n13368), .ZN(n13366) );
  NAND2_X1 U13403 ( .A1(b_12_), .A2(a_19_), .ZN(n13368) );
  XOR2_X1 U13404 ( .A(n13369), .B(n13370), .Z(n13160) );
  XNOR2_X1 U13405 ( .A(n13371), .B(n13372), .ZN(n13370) );
  NAND2_X1 U13406 ( .A1(b_12_), .A2(a_18_), .ZN(n13372) );
  XNOR2_X1 U13407 ( .A(n13373), .B(n13374), .ZN(n13164) );
  XNOR2_X1 U13408 ( .A(n13375), .B(n13376), .ZN(n13373) );
  XNOR2_X1 U13409 ( .A(n13377), .B(n13378), .ZN(n13040) );
  XNOR2_X1 U13410 ( .A(n13379), .B(n13380), .ZN(n13377) );
  XOR2_X1 U13411 ( .A(n13381), .B(n13382), .Z(n13167) );
  XNOR2_X1 U13412 ( .A(n13383), .B(n13384), .ZN(n13382) );
  NAND2_X1 U13413 ( .A1(b_12_), .A2(a_15_), .ZN(n13384) );
  XOR2_X1 U13414 ( .A(n13385), .B(n13386), .Z(n13017) );
  XOR2_X1 U13415 ( .A(n13387), .B(n13388), .Z(n13386) );
  XNOR2_X1 U13416 ( .A(n13389), .B(n13390), .ZN(n13175) );
  XNOR2_X1 U13417 ( .A(n13391), .B(n13392), .ZN(n13390) );
  XNOR2_X1 U13418 ( .A(n13393), .B(n13394), .ZN(n13004) );
  NOR2_X1 U13419 ( .A1(n13395), .A2(n13396), .ZN(n13394) );
  NOR2_X1 U13420 ( .A1(n13397), .A2(n13398), .ZN(n13395) );
  NOR2_X1 U13421 ( .A1(n8402), .A2(n13118), .ZN(n13398) );
  INV_X1 U13422 ( .A(n13399), .ZN(n13397) );
  XOR2_X1 U13423 ( .A(n13400), .B(n13401), .Z(n12996) );
  NAND2_X1 U13424 ( .A1(n13402), .A2(n13403), .ZN(n13400) );
  XNOR2_X1 U13425 ( .A(n13404), .B(n13405), .ZN(n12988) );
  NAND2_X1 U13426 ( .A1(n13406), .A2(n13407), .ZN(n13404) );
  XOR2_X1 U13427 ( .A(n13408), .B(n13409), .Z(n13179) );
  NAND2_X1 U13428 ( .A1(n13410), .A2(n13411), .ZN(n13408) );
  XOR2_X1 U13429 ( .A(n13412), .B(n13413), .Z(n12976) );
  NAND2_X1 U13430 ( .A1(n13414), .A2(n13415), .ZN(n13412) );
  XOR2_X1 U13431 ( .A(n13416), .B(n13417), .Z(n12969) );
  NAND2_X1 U13432 ( .A1(n13418), .A2(n13419), .ZN(n13416) );
  XOR2_X1 U13433 ( .A(n13420), .B(n13421), .Z(n12960) );
  NAND2_X1 U13434 ( .A1(n13422), .A2(n13423), .ZN(n13420) );
  XOR2_X1 U13435 ( .A(n13424), .B(n13425), .Z(n13184) );
  NAND2_X1 U13436 ( .A1(n13426), .A2(n13427), .ZN(n13424) );
  XNOR2_X1 U13437 ( .A(n13428), .B(n13429), .ZN(n12947) );
  NAND2_X1 U13438 ( .A1(n13430), .A2(n13431), .ZN(n13428) );
  XOR2_X1 U13439 ( .A(n13432), .B(n13433), .Z(n12941) );
  XOR2_X1 U13440 ( .A(n13434), .B(n13435), .Z(n13433) );
  XOR2_X1 U13441 ( .A(n12939), .B(n13436), .Z(n13187) );
  XNOR2_X1 U13442 ( .A(n13437), .B(n13438), .ZN(n12939) );
  XNOR2_X1 U13443 ( .A(n13439), .B(n13440), .ZN(n8546) );
  NAND2_X1 U13444 ( .A1(n8553), .A2(n8552), .ZN(n8551) );
  NOR2_X1 U13445 ( .A1(n13441), .A2(n8585), .ZN(n8552) );
  INV_X1 U13446 ( .A(n13442), .ZN(n13441) );
  NAND2_X1 U13447 ( .A1(n13443), .A2(n13444), .ZN(n13442) );
  INV_X1 U13448 ( .A(n13445), .ZN(n8553) );
  NAND2_X1 U13449 ( .A1(n13440), .A2(n13439), .ZN(n13445) );
  NAND2_X1 U13450 ( .A1(n13446), .A2(n13447), .ZN(n13439) );
  NAND2_X1 U13451 ( .A1(n13438), .A2(n13448), .ZN(n13447) );
  NAND2_X1 U13452 ( .A1(n13436), .A2(n13437), .ZN(n13448) );
  INV_X1 U13453 ( .A(n12938), .ZN(n13436) );
  NOR2_X1 U13454 ( .A1(n13118), .A2(n8457), .ZN(n13438) );
  NAND2_X1 U13455 ( .A1(n12938), .A2(n13449), .ZN(n13446) );
  INV_X1 U13456 ( .A(n13437), .ZN(n13449) );
  NOR2_X1 U13457 ( .A1(n13450), .A2(n13451), .ZN(n13437) );
  NOR2_X1 U13458 ( .A1(n13435), .A2(n13452), .ZN(n13451) );
  NOR2_X1 U13459 ( .A1(n13432), .A2(n13434), .ZN(n13452) );
  NAND2_X1 U13460 ( .A1(b_12_), .A2(a_1_), .ZN(n13435) );
  INV_X1 U13461 ( .A(n13453), .ZN(n13450) );
  NAND2_X1 U13462 ( .A1(n13432), .A2(n13434), .ZN(n13453) );
  NAND2_X1 U13463 ( .A1(n13430), .A2(n13454), .ZN(n13434) );
  NAND2_X1 U13464 ( .A1(n13429), .A2(n13431), .ZN(n13454) );
  NAND2_X1 U13465 ( .A1(n13455), .A2(n13456), .ZN(n13431) );
  NAND2_X1 U13466 ( .A1(b_12_), .A2(a_2_), .ZN(n13456) );
  INV_X1 U13467 ( .A(n13457), .ZN(n13455) );
  XNOR2_X1 U13468 ( .A(n13458), .B(n13459), .ZN(n13429) );
  XOR2_X1 U13469 ( .A(n13460), .B(n13461), .Z(n13459) );
  NAND2_X1 U13470 ( .A1(a_3_), .A2(b_11_), .ZN(n13461) );
  NAND2_X1 U13471 ( .A1(a_2_), .A2(n13457), .ZN(n13430) );
  NAND2_X1 U13472 ( .A1(n13426), .A2(n13462), .ZN(n13457) );
  NAND2_X1 U13473 ( .A1(n13425), .A2(n13427), .ZN(n13462) );
  NAND2_X1 U13474 ( .A1(n13463), .A2(n13464), .ZN(n13427) );
  NAND2_X1 U13475 ( .A1(b_12_), .A2(a_3_), .ZN(n13464) );
  INV_X1 U13476 ( .A(n13465), .ZN(n13463) );
  XOR2_X1 U13477 ( .A(n13466), .B(n13467), .Z(n13425) );
  XNOR2_X1 U13478 ( .A(n13468), .B(n13469), .ZN(n13467) );
  NAND2_X1 U13479 ( .A1(a_4_), .A2(b_11_), .ZN(n13469) );
  NAND2_X1 U13480 ( .A1(a_3_), .A2(n13465), .ZN(n13426) );
  NAND2_X1 U13481 ( .A1(n13422), .A2(n13470), .ZN(n13465) );
  NAND2_X1 U13482 ( .A1(n13421), .A2(n13423), .ZN(n13470) );
  NAND2_X1 U13483 ( .A1(n13471), .A2(n13472), .ZN(n13423) );
  NAND2_X1 U13484 ( .A1(b_12_), .A2(a_4_), .ZN(n13472) );
  INV_X1 U13485 ( .A(n13473), .ZN(n13471) );
  XOR2_X1 U13486 ( .A(n13474), .B(n13475), .Z(n13421) );
  XOR2_X1 U13487 ( .A(n13476), .B(n13477), .Z(n13474) );
  NOR2_X1 U13488 ( .A1(n13332), .A2(n8938), .ZN(n13477) );
  NAND2_X1 U13489 ( .A1(a_4_), .A2(n13473), .ZN(n13422) );
  NAND2_X1 U13490 ( .A1(n13418), .A2(n13478), .ZN(n13473) );
  NAND2_X1 U13491 ( .A1(n13417), .A2(n13419), .ZN(n13478) );
  NAND2_X1 U13492 ( .A1(n13479), .A2(n13480), .ZN(n13419) );
  NAND2_X1 U13493 ( .A1(b_12_), .A2(a_5_), .ZN(n13480) );
  INV_X1 U13494 ( .A(n13481), .ZN(n13479) );
  XNOR2_X1 U13495 ( .A(n13482), .B(n13483), .ZN(n13417) );
  XOR2_X1 U13496 ( .A(n13484), .B(n13485), .Z(n13483) );
  NAND2_X1 U13497 ( .A1(a_6_), .A2(b_11_), .ZN(n13485) );
  NAND2_X1 U13498 ( .A1(a_5_), .A2(n13481), .ZN(n13418) );
  NAND2_X1 U13499 ( .A1(n13414), .A2(n13486), .ZN(n13481) );
  NAND2_X1 U13500 ( .A1(n13413), .A2(n13415), .ZN(n13486) );
  NAND2_X1 U13501 ( .A1(n13487), .A2(n13488), .ZN(n13415) );
  NAND2_X1 U13502 ( .A1(b_12_), .A2(a_6_), .ZN(n13488) );
  INV_X1 U13503 ( .A(n13489), .ZN(n13487) );
  XOR2_X1 U13504 ( .A(n13490), .B(n13491), .Z(n13413) );
  XOR2_X1 U13505 ( .A(n13492), .B(n13493), .Z(n13490) );
  NOR2_X1 U13506 ( .A1(n13332), .A2(n8425), .ZN(n13493) );
  NAND2_X1 U13507 ( .A1(a_6_), .A2(n13489), .ZN(n13414) );
  NAND2_X1 U13508 ( .A1(n13410), .A2(n13494), .ZN(n13489) );
  NAND2_X1 U13509 ( .A1(n13409), .A2(n13411), .ZN(n13494) );
  NAND2_X1 U13510 ( .A1(n13495), .A2(n13496), .ZN(n13411) );
  NAND2_X1 U13511 ( .A1(b_12_), .A2(a_7_), .ZN(n13496) );
  INV_X1 U13512 ( .A(n13497), .ZN(n13495) );
  XNOR2_X1 U13513 ( .A(n13498), .B(n13499), .ZN(n13409) );
  XOR2_X1 U13514 ( .A(n13500), .B(n13501), .Z(n13499) );
  NAND2_X1 U13515 ( .A1(a_8_), .A2(b_11_), .ZN(n13501) );
  NAND2_X1 U13516 ( .A1(a_7_), .A2(n13497), .ZN(n13410) );
  NAND2_X1 U13517 ( .A1(n13406), .A2(n13502), .ZN(n13497) );
  NAND2_X1 U13518 ( .A1(n13405), .A2(n13407), .ZN(n13502) );
  NAND2_X1 U13519 ( .A1(n13503), .A2(n13504), .ZN(n13407) );
  NAND2_X1 U13520 ( .A1(b_12_), .A2(a_8_), .ZN(n13504) );
  INV_X1 U13521 ( .A(n13505), .ZN(n13503) );
  XNOR2_X1 U13522 ( .A(n13506), .B(n13507), .ZN(n13405) );
  XNOR2_X1 U13523 ( .A(n13508), .B(n13509), .ZN(n13506) );
  NOR2_X1 U13524 ( .A1(n13332), .A2(n8971), .ZN(n13509) );
  NAND2_X1 U13525 ( .A1(a_8_), .A2(n13505), .ZN(n13406) );
  NAND2_X1 U13526 ( .A1(n13402), .A2(n13510), .ZN(n13505) );
  NAND2_X1 U13527 ( .A1(n13401), .A2(n13403), .ZN(n13510) );
  NAND2_X1 U13528 ( .A1(n13511), .A2(n13512), .ZN(n13403) );
  NAND2_X1 U13529 ( .A1(b_12_), .A2(a_9_), .ZN(n13512) );
  INV_X1 U13530 ( .A(n13513), .ZN(n13511) );
  XNOR2_X1 U13531 ( .A(n13514), .B(n13515), .ZN(n13401) );
  XOR2_X1 U13532 ( .A(n13516), .B(n13517), .Z(n13515) );
  NAND2_X1 U13533 ( .A1(a_10_), .A2(b_11_), .ZN(n13517) );
  NAND2_X1 U13534 ( .A1(a_9_), .A2(n13513), .ZN(n13402) );
  NAND2_X1 U13535 ( .A1(n13518), .A2(n13519), .ZN(n13513) );
  NAND2_X1 U13536 ( .A1(n13393), .A2(n13520), .ZN(n13519) );
  NAND2_X1 U13537 ( .A1(n13399), .A2(n13521), .ZN(n13520) );
  NAND2_X1 U13538 ( .A1(b_12_), .A2(a_10_), .ZN(n13521) );
  XNOR2_X1 U13539 ( .A(n13522), .B(n13523), .ZN(n13393) );
  XNOR2_X1 U13540 ( .A(n13524), .B(n13525), .ZN(n13522) );
  INV_X1 U13541 ( .A(n13396), .ZN(n13518) );
  NOR2_X1 U13542 ( .A1(n13399), .A2(n8402), .ZN(n13396) );
  NAND2_X1 U13543 ( .A1(n13526), .A2(n13527), .ZN(n13399) );
  NAND2_X1 U13544 ( .A1(n13389), .A2(n13528), .ZN(n13527) );
  INV_X1 U13545 ( .A(n13529), .ZN(n13528) );
  NOR2_X1 U13546 ( .A1(n13392), .A2(n13391), .ZN(n13529) );
  XOR2_X1 U13547 ( .A(n13530), .B(n13531), .Z(n13389) );
  XNOR2_X1 U13548 ( .A(n13532), .B(n13533), .ZN(n13530) );
  NOR2_X1 U13549 ( .A1(n13332), .A2(n8393), .ZN(n13533) );
  NAND2_X1 U13550 ( .A1(n13391), .A2(n13392), .ZN(n13526) );
  NAND2_X1 U13551 ( .A1(b_12_), .A2(a_11_), .ZN(n13392) );
  NOR2_X1 U13552 ( .A1(n13534), .A2(n13535), .ZN(n13391) );
  NOR2_X1 U13553 ( .A1(n13387), .A2(n13536), .ZN(n13535) );
  NOR2_X1 U13554 ( .A1(n13385), .A2(n13388), .ZN(n13536) );
  INV_X1 U13555 ( .A(n13537), .ZN(n13534) );
  NAND2_X1 U13556 ( .A1(n13385), .A2(n13388), .ZN(n13537) );
  NAND2_X1 U13557 ( .A1(n13242), .A2(n13538), .ZN(n13388) );
  NAND2_X1 U13558 ( .A1(n13241), .A2(n13243), .ZN(n13538) );
  NAND2_X1 U13559 ( .A1(n13539), .A2(n13540), .ZN(n13243) );
  NAND2_X1 U13560 ( .A1(b_12_), .A2(a_13_), .ZN(n13540) );
  INV_X1 U13561 ( .A(n13541), .ZN(n13539) );
  XOR2_X1 U13562 ( .A(n13542), .B(n13543), .Z(n13241) );
  XNOR2_X1 U13563 ( .A(n13544), .B(n13545), .ZN(n13543) );
  NAND2_X1 U13564 ( .A1(a_14_), .A2(b_11_), .ZN(n13545) );
  NAND2_X1 U13565 ( .A1(a_13_), .A2(n13541), .ZN(n13242) );
  NAND2_X1 U13566 ( .A1(n13250), .A2(n13546), .ZN(n13541) );
  NAND2_X1 U13567 ( .A1(n13249), .A2(n13251), .ZN(n13546) );
  NAND2_X1 U13568 ( .A1(n13547), .A2(n13548), .ZN(n13251) );
  NAND2_X1 U13569 ( .A1(b_12_), .A2(a_14_), .ZN(n13548) );
  INV_X1 U13570 ( .A(n13549), .ZN(n13547) );
  XOR2_X1 U13571 ( .A(n13550), .B(n13551), .Z(n13249) );
  XOR2_X1 U13572 ( .A(n13552), .B(n13553), .Z(n13550) );
  NOR2_X1 U13573 ( .A1(n13332), .A2(n8850), .ZN(n13553) );
  NAND2_X1 U13574 ( .A1(a_14_), .A2(n13549), .ZN(n13250) );
  NAND2_X1 U13575 ( .A1(n13554), .A2(n13555), .ZN(n13549) );
  NAND3_X1 U13576 ( .A1(a_15_), .A2(n13556), .A3(b_12_), .ZN(n13555) );
  NAND2_X1 U13577 ( .A1(n13383), .A2(n13381), .ZN(n13556) );
  NAND2_X1 U13578 ( .A1(n13557), .A2(n13558), .ZN(n13554) );
  INV_X1 U13579 ( .A(n13383), .ZN(n13558) );
  NOR2_X1 U13580 ( .A1(n13559), .A2(n13560), .ZN(n13383) );
  INV_X1 U13581 ( .A(n13561), .ZN(n13560) );
  NAND2_X1 U13582 ( .A1(n13379), .A2(n13562), .ZN(n13561) );
  NAND2_X1 U13583 ( .A1(n13380), .A2(n13378), .ZN(n13562) );
  NOR2_X1 U13584 ( .A1(n13118), .A2(n8376), .ZN(n13379) );
  NOR2_X1 U13585 ( .A1(n13378), .A2(n13380), .ZN(n13559) );
  NOR2_X1 U13586 ( .A1(n13563), .A2(n13564), .ZN(n13380) );
  INV_X1 U13587 ( .A(n13565), .ZN(n13564) );
  NAND2_X1 U13588 ( .A1(n13376), .A2(n13566), .ZN(n13565) );
  NAND2_X1 U13589 ( .A1(n13375), .A2(n13374), .ZN(n13566) );
  NOR2_X1 U13590 ( .A1(n13118), .A2(n8371), .ZN(n13376) );
  NOR2_X1 U13591 ( .A1(n13374), .A2(n13375), .ZN(n13563) );
  NOR2_X1 U13592 ( .A1(n13567), .A2(n13568), .ZN(n13375) );
  INV_X1 U13593 ( .A(n13569), .ZN(n13568) );
  NAND3_X1 U13594 ( .A1(a_18_), .A2(n13570), .A3(b_12_), .ZN(n13569) );
  NAND2_X1 U13595 ( .A1(n13371), .A2(n13369), .ZN(n13570) );
  NOR2_X1 U13596 ( .A1(n13369), .A2(n13371), .ZN(n13567) );
  NOR2_X1 U13597 ( .A1(n13571), .A2(n13572), .ZN(n13371) );
  NOR3_X1 U13598 ( .A1(n8742), .A2(n13573), .A3(n13118), .ZN(n13572) );
  INV_X1 U13599 ( .A(n13574), .ZN(n13573) );
  NAND2_X1 U13600 ( .A1(n13367), .A2(n13365), .ZN(n13574) );
  NOR2_X1 U13601 ( .A1(n13365), .A2(n13367), .ZN(n13571) );
  NOR2_X1 U13602 ( .A1(n13575), .A2(n13576), .ZN(n13367) );
  INV_X1 U13603 ( .A(n13577), .ZN(n13576) );
  NAND3_X1 U13604 ( .A1(a_20_), .A2(n13578), .A3(b_12_), .ZN(n13577) );
  NAND2_X1 U13605 ( .A1(n13362), .A2(n13363), .ZN(n13578) );
  NOR2_X1 U13606 ( .A1(n13362), .A2(n13363), .ZN(n13575) );
  NOR2_X1 U13607 ( .A1(n13579), .A2(n13580), .ZN(n13363) );
  NOR3_X1 U13608 ( .A1(n8759), .A2(n13581), .A3(n13118), .ZN(n13580) );
  NOR2_X1 U13609 ( .A1(n13359), .A2(n13358), .ZN(n13581) );
  INV_X1 U13610 ( .A(n13582), .ZN(n13579) );
  NAND2_X1 U13611 ( .A1(n13358), .A2(n13359), .ZN(n13582) );
  NAND2_X1 U13612 ( .A1(n13583), .A2(n13584), .ZN(n13359) );
  NAND2_X1 U13613 ( .A1(n13356), .A2(n13585), .ZN(n13584) );
  INV_X1 U13614 ( .A(n13586), .ZN(n13585) );
  NOR2_X1 U13615 ( .A1(n13353), .A2(n13355), .ZN(n13586) );
  NOR2_X1 U13616 ( .A1(n13118), .A2(n12296), .ZN(n13356) );
  NAND2_X1 U13617 ( .A1(n13353), .A2(n13355), .ZN(n13583) );
  NAND2_X1 U13618 ( .A1(n13587), .A2(n13588), .ZN(n13355) );
  NAND2_X1 U13619 ( .A1(n13352), .A2(n13589), .ZN(n13588) );
  INV_X1 U13620 ( .A(n13590), .ZN(n13589) );
  NOR2_X1 U13621 ( .A1(n13351), .A2(n13350), .ZN(n13590) );
  NOR2_X1 U13622 ( .A1(n13118), .A2(n12301), .ZN(n13352) );
  NAND2_X1 U13623 ( .A1(n13350), .A2(n13351), .ZN(n13587) );
  NAND2_X1 U13624 ( .A1(n13591), .A2(n13592), .ZN(n13351) );
  NAND2_X1 U13625 ( .A1(n13348), .A2(n13593), .ZN(n13592) );
  INV_X1 U13626 ( .A(n13594), .ZN(n13593) );
  NOR2_X1 U13627 ( .A1(n13346), .A2(n13347), .ZN(n13594) );
  NOR2_X1 U13628 ( .A1(n13118), .A2(n8779), .ZN(n13348) );
  NAND2_X1 U13629 ( .A1(n13346), .A2(n13347), .ZN(n13591) );
  NAND2_X1 U13630 ( .A1(n13595), .A2(n13596), .ZN(n13347) );
  NAND2_X1 U13631 ( .A1(n13344), .A2(n13597), .ZN(n13596) );
  NAND2_X1 U13632 ( .A1(n13341), .A2(n13343), .ZN(n13597) );
  NOR2_X1 U13633 ( .A1(n13118), .A2(n8788), .ZN(n13344) );
  INV_X1 U13634 ( .A(n13598), .ZN(n13595) );
  NOR2_X1 U13635 ( .A1(n13343), .A2(n13341), .ZN(n13598) );
  XNOR2_X1 U13636 ( .A(n13599), .B(n13600), .ZN(n13341) );
  XNOR2_X1 U13637 ( .A(n13601), .B(n13602), .ZN(n13600) );
  NAND2_X1 U13638 ( .A1(n13603), .A2(n13604), .ZN(n13343) );
  NAND2_X1 U13639 ( .A1(n13302), .A2(n13605), .ZN(n13604) );
  NAND2_X1 U13640 ( .A1(n13305), .A2(n13304), .ZN(n13605) );
  XOR2_X1 U13641 ( .A(n13606), .B(n13607), .Z(n13302) );
  XNOR2_X1 U13642 ( .A(n13608), .B(n13609), .ZN(n13606) );
  INV_X1 U13643 ( .A(n13610), .ZN(n13603) );
  NOR2_X1 U13644 ( .A1(n13304), .A2(n13305), .ZN(n13610) );
  NOR2_X1 U13645 ( .A1(n13118), .A2(n9344), .ZN(n13305) );
  NAND2_X1 U13646 ( .A1(n13611), .A2(n13612), .ZN(n13304) );
  NAND2_X1 U13647 ( .A1(n13312), .A2(n13613), .ZN(n13612) );
  INV_X1 U13648 ( .A(n13614), .ZN(n13613) );
  NOR2_X1 U13649 ( .A1(n13310), .A2(n13311), .ZN(n13614) );
  NOR2_X1 U13650 ( .A1(n13118), .A2(n8797), .ZN(n13312) );
  NAND2_X1 U13651 ( .A1(n13310), .A2(n13311), .ZN(n13611) );
  NAND2_X1 U13652 ( .A1(n13615), .A2(n13616), .ZN(n13311) );
  NAND2_X1 U13653 ( .A1(n13339), .A2(n13617), .ZN(n13616) );
  INV_X1 U13654 ( .A(n13618), .ZN(n13617) );
  NOR2_X1 U13655 ( .A1(n13340), .A2(n13338), .ZN(n13618) );
  NOR2_X1 U13656 ( .A1(n13118), .A2(n8314), .ZN(n13339) );
  NAND2_X1 U13657 ( .A1(n13338), .A2(n13340), .ZN(n13615) );
  NAND2_X1 U13658 ( .A1(n13619), .A2(n13620), .ZN(n13340) );
  NAND2_X1 U13659 ( .A1(n13334), .A2(n13621), .ZN(n13620) );
  INV_X1 U13660 ( .A(n13622), .ZN(n13621) );
  NOR2_X1 U13661 ( .A1(n13335), .A2(n13336), .ZN(n13622) );
  NOR2_X1 U13662 ( .A1(n13118), .A2(n9098), .ZN(n13334) );
  NAND2_X1 U13663 ( .A1(n13336), .A2(n13335), .ZN(n13619) );
  NAND2_X1 U13664 ( .A1(n13623), .A2(n13624), .ZN(n13335) );
  NAND2_X1 U13665 ( .A1(b_10_), .A2(n13625), .ZN(n13624) );
  NAND2_X1 U13666 ( .A1(n8299), .A2(n13626), .ZN(n13625) );
  NAND2_X1 U13667 ( .A1(a_31_), .A2(n13332), .ZN(n13626) );
  NAND2_X1 U13668 ( .A1(b_11_), .A2(n13627), .ZN(n13623) );
  NAND2_X1 U13669 ( .A1(n8303), .A2(n13628), .ZN(n13627) );
  NAND2_X1 U13670 ( .A1(a_30_), .A2(n13629), .ZN(n13628) );
  NOR3_X1 U13671 ( .A1(n9631), .A2(n13332), .A3(n13118), .ZN(n13336) );
  XOR2_X1 U13672 ( .A(n13630), .B(n13631), .Z(n13338) );
  XNOR2_X1 U13673 ( .A(n13632), .B(n13633), .ZN(n13630) );
  XNOR2_X1 U13674 ( .A(n13634), .B(n13635), .ZN(n13310) );
  XNOR2_X1 U13675 ( .A(n13636), .B(n13637), .ZN(n13634) );
  XNOR2_X1 U13676 ( .A(n13638), .B(n13639), .ZN(n13346) );
  XNOR2_X1 U13677 ( .A(n13640), .B(n13641), .ZN(n13639) );
  XNOR2_X1 U13678 ( .A(n13642), .B(n13643), .ZN(n13350) );
  XNOR2_X1 U13679 ( .A(n13644), .B(n13645), .ZN(n13642) );
  XOR2_X1 U13680 ( .A(n13646), .B(n13647), .Z(n13353) );
  XOR2_X1 U13681 ( .A(n13648), .B(n13649), .Z(n13646) );
  XNOR2_X1 U13682 ( .A(n13650), .B(n13651), .ZN(n13358) );
  XNOR2_X1 U13683 ( .A(n13652), .B(n13653), .ZN(n13651) );
  XNOR2_X1 U13684 ( .A(n13654), .B(n13655), .ZN(n13362) );
  XOR2_X1 U13685 ( .A(n13656), .B(n13657), .Z(n13654) );
  XNOR2_X1 U13686 ( .A(n13658), .B(n13659), .ZN(n13365) );
  XOR2_X1 U13687 ( .A(n13660), .B(n13661), .Z(n13658) );
  XOR2_X1 U13688 ( .A(n13662), .B(n13663), .Z(n13369) );
  XOR2_X1 U13689 ( .A(n13664), .B(n13665), .Z(n13663) );
  XOR2_X1 U13690 ( .A(n13666), .B(n13667), .Z(n13374) );
  NAND2_X1 U13691 ( .A1(n13668), .A2(n13669), .ZN(n13666) );
  XNOR2_X1 U13692 ( .A(n13670), .B(n13671), .ZN(n13378) );
  XOR2_X1 U13693 ( .A(n13672), .B(n13673), .Z(n13670) );
  NOR2_X1 U13694 ( .A1(n13332), .A2(n8371), .ZN(n13673) );
  INV_X1 U13695 ( .A(n13381), .ZN(n13557) );
  XOR2_X1 U13696 ( .A(n13674), .B(n13675), .Z(n13381) );
  XOR2_X1 U13697 ( .A(n13676), .B(n13677), .Z(n13675) );
  NAND2_X1 U13698 ( .A1(a_16_), .A2(b_11_), .ZN(n13677) );
  XOR2_X1 U13699 ( .A(n13678), .B(n13679), .Z(n13385) );
  XNOR2_X1 U13700 ( .A(n13680), .B(n13681), .ZN(n13679) );
  NAND2_X1 U13701 ( .A1(a_13_), .A2(b_11_), .ZN(n13681) );
  XNOR2_X1 U13702 ( .A(n13682), .B(n13683), .ZN(n13432) );
  XOR2_X1 U13703 ( .A(n13684), .B(n13685), .Z(n13683) );
  NAND2_X1 U13704 ( .A1(a_2_), .A2(b_11_), .ZN(n13685) );
  XOR2_X1 U13705 ( .A(n13686), .B(n13687), .Z(n12938) );
  XNOR2_X1 U13706 ( .A(n13688), .B(n13689), .ZN(n13687) );
  NAND2_X1 U13707 ( .A1(a_1_), .A2(b_11_), .ZN(n13689) );
  XNOR2_X1 U13708 ( .A(n13690), .B(n13691), .ZN(n13440) );
  XNOR2_X1 U13709 ( .A(n13692), .B(n13693), .ZN(n13690) );
  NOR2_X1 U13710 ( .A1(n13332), .A2(n8457), .ZN(n13693) );
  NOR2_X1 U13711 ( .A1(n13444), .A2(n13443), .ZN(n8585) );
  NOR2_X1 U13712 ( .A1(n13694), .A2(n13695), .ZN(n13443) );
  INV_X1 U13713 ( .A(n13696), .ZN(n13695) );
  NAND3_X1 U13714 ( .A1(b_11_), .A2(n13697), .A3(a_0_), .ZN(n13696) );
  NAND2_X1 U13715 ( .A1(n13692), .A2(n13691), .ZN(n13697) );
  NOR2_X1 U13716 ( .A1(n13691), .A2(n13692), .ZN(n13694) );
  NOR2_X1 U13717 ( .A1(n13698), .A2(n13699), .ZN(n13692) );
  INV_X1 U13718 ( .A(n13700), .ZN(n13699) );
  NAND3_X1 U13719 ( .A1(b_11_), .A2(n13701), .A3(a_1_), .ZN(n13700) );
  NAND2_X1 U13720 ( .A1(n13688), .A2(n13686), .ZN(n13701) );
  NOR2_X1 U13721 ( .A1(n13686), .A2(n13688), .ZN(n13698) );
  NOR2_X1 U13722 ( .A1(n13702), .A2(n13703), .ZN(n13688) );
  NOR3_X1 U13723 ( .A1(n13332), .A2(n13704), .A3(n8448), .ZN(n13703) );
  NOR2_X1 U13724 ( .A1(n13684), .A2(n13682), .ZN(n13704) );
  INV_X1 U13725 ( .A(n13705), .ZN(n13702) );
  NAND2_X1 U13726 ( .A1(n13682), .A2(n13684), .ZN(n13705) );
  NAND2_X1 U13727 ( .A1(n13706), .A2(n13707), .ZN(n13684) );
  INV_X1 U13728 ( .A(n13708), .ZN(n13707) );
  NOR3_X1 U13729 ( .A1(n13332), .A2(n13709), .A3(n8900), .ZN(n13708) );
  NOR2_X1 U13730 ( .A1(n13460), .A2(n13458), .ZN(n13709) );
  NAND2_X1 U13731 ( .A1(n13458), .A2(n13460), .ZN(n13706) );
  NAND2_X1 U13732 ( .A1(n13710), .A2(n13711), .ZN(n13460) );
  NAND3_X1 U13733 ( .A1(b_11_), .A2(n13712), .A3(a_4_), .ZN(n13711) );
  NAND2_X1 U13734 ( .A1(n13468), .A2(n13466), .ZN(n13712) );
  INV_X1 U13735 ( .A(n13713), .ZN(n13710) );
  NOR2_X1 U13736 ( .A1(n13466), .A2(n13468), .ZN(n13713) );
  NOR2_X1 U13737 ( .A1(n13714), .A2(n13715), .ZN(n13468) );
  NOR3_X1 U13738 ( .A1(n13332), .A2(n13716), .A3(n8938), .ZN(n13715) );
  NOR2_X1 U13739 ( .A1(n13476), .A2(n13475), .ZN(n13716) );
  INV_X1 U13740 ( .A(n13717), .ZN(n13714) );
  NAND2_X1 U13741 ( .A1(n13475), .A2(n13476), .ZN(n13717) );
  NAND2_X1 U13742 ( .A1(n13718), .A2(n13719), .ZN(n13476) );
  NAND3_X1 U13743 ( .A1(b_11_), .A2(n13720), .A3(a_6_), .ZN(n13719) );
  INV_X1 U13744 ( .A(n13721), .ZN(n13720) );
  NOR2_X1 U13745 ( .A1(n13484), .A2(n13482), .ZN(n13721) );
  NAND2_X1 U13746 ( .A1(n13482), .A2(n13484), .ZN(n13718) );
  NAND2_X1 U13747 ( .A1(n13722), .A2(n13723), .ZN(n13484) );
  NAND3_X1 U13748 ( .A1(b_11_), .A2(n13724), .A3(a_7_), .ZN(n13723) );
  INV_X1 U13749 ( .A(n13725), .ZN(n13724) );
  NOR2_X1 U13750 ( .A1(n13492), .A2(n13491), .ZN(n13725) );
  NAND2_X1 U13751 ( .A1(n13491), .A2(n13492), .ZN(n13722) );
  NAND2_X1 U13752 ( .A1(n13726), .A2(n13727), .ZN(n13492) );
  NAND3_X1 U13753 ( .A1(b_11_), .A2(n13728), .A3(a_8_), .ZN(n13727) );
  INV_X1 U13754 ( .A(n13729), .ZN(n13728) );
  NOR2_X1 U13755 ( .A1(n13500), .A2(n13498), .ZN(n13729) );
  NAND2_X1 U13756 ( .A1(n13498), .A2(n13500), .ZN(n13726) );
  NAND2_X1 U13757 ( .A1(n13730), .A2(n13731), .ZN(n13500) );
  NAND3_X1 U13758 ( .A1(b_11_), .A2(n13732), .A3(a_9_), .ZN(n13731) );
  NAND2_X1 U13759 ( .A1(n13508), .A2(n13507), .ZN(n13732) );
  INV_X1 U13760 ( .A(n13733), .ZN(n13730) );
  NOR2_X1 U13761 ( .A1(n13507), .A2(n13508), .ZN(n13733) );
  NOR2_X1 U13762 ( .A1(n13734), .A2(n13735), .ZN(n13508) );
  NOR3_X1 U13763 ( .A1(n13332), .A2(n13736), .A3(n8402), .ZN(n13735) );
  INV_X1 U13764 ( .A(n13737), .ZN(n13736) );
  NAND2_X1 U13765 ( .A1(n13514), .A2(n13516), .ZN(n13737) );
  NOR2_X1 U13766 ( .A1(n13516), .A2(n13514), .ZN(n13734) );
  XOR2_X1 U13767 ( .A(n13738), .B(n13739), .Z(n13514) );
  NAND2_X1 U13768 ( .A1(n13740), .A2(n13741), .ZN(n13738) );
  NAND2_X1 U13769 ( .A1(n13742), .A2(n13743), .ZN(n13516) );
  NAND2_X1 U13770 ( .A1(n13523), .A2(n13744), .ZN(n13743) );
  NAND2_X1 U13771 ( .A1(n13525), .A2(n13745), .ZN(n13744) );
  XNOR2_X1 U13772 ( .A(n13746), .B(n13747), .ZN(n13523) );
  XOR2_X1 U13773 ( .A(n13748), .B(n13749), .Z(n13746) );
  NOR2_X1 U13774 ( .A1(n13629), .A2(n8393), .ZN(n13749) );
  INV_X1 U13775 ( .A(n13750), .ZN(n13742) );
  NOR2_X1 U13776 ( .A1(n13745), .A2(n13525), .ZN(n13750) );
  INV_X1 U13777 ( .A(n13524), .ZN(n13745) );
  NOR2_X1 U13778 ( .A1(n13751), .A2(n13752), .ZN(n13524) );
  NOR3_X1 U13779 ( .A1(n13332), .A2(n13753), .A3(n8393), .ZN(n13752) );
  INV_X1 U13780 ( .A(n13754), .ZN(n13753) );
  NAND2_X1 U13781 ( .A1(n13532), .A2(n13531), .ZN(n13754) );
  NOR2_X1 U13782 ( .A1(n13531), .A2(n13532), .ZN(n13751) );
  NOR2_X1 U13783 ( .A1(n13755), .A2(n13756), .ZN(n13532) );
  INV_X1 U13784 ( .A(n13757), .ZN(n13756) );
  NAND3_X1 U13785 ( .A1(b_11_), .A2(n13758), .A3(a_13_), .ZN(n13757) );
  NAND2_X1 U13786 ( .A1(n13680), .A2(n13678), .ZN(n13758) );
  NOR2_X1 U13787 ( .A1(n13678), .A2(n13680), .ZN(n13755) );
  NOR2_X1 U13788 ( .A1(n13759), .A2(n13760), .ZN(n13680) );
  INV_X1 U13789 ( .A(n13761), .ZN(n13760) );
  NAND3_X1 U13790 ( .A1(b_11_), .A2(n13762), .A3(a_14_), .ZN(n13761) );
  NAND2_X1 U13791 ( .A1(n13544), .A2(n13542), .ZN(n13762) );
  NOR2_X1 U13792 ( .A1(n13542), .A2(n13544), .ZN(n13759) );
  NOR2_X1 U13793 ( .A1(n13763), .A2(n13764), .ZN(n13544) );
  NOR3_X1 U13794 ( .A1(n13332), .A2(n13765), .A3(n8850), .ZN(n13764) );
  NOR2_X1 U13795 ( .A1(n13552), .A2(n13551), .ZN(n13765) );
  INV_X1 U13796 ( .A(n13766), .ZN(n13763) );
  NAND2_X1 U13797 ( .A1(n13551), .A2(n13552), .ZN(n13766) );
  NAND2_X1 U13798 ( .A1(n13767), .A2(n13768), .ZN(n13552) );
  NAND3_X1 U13799 ( .A1(b_11_), .A2(n13769), .A3(a_16_), .ZN(n13768) );
  INV_X1 U13800 ( .A(n13770), .ZN(n13769) );
  NOR2_X1 U13801 ( .A1(n13676), .A2(n13674), .ZN(n13770) );
  NAND2_X1 U13802 ( .A1(n13674), .A2(n13676), .ZN(n13767) );
  NAND2_X1 U13803 ( .A1(n13771), .A2(n13772), .ZN(n13676) );
  NAND3_X1 U13804 ( .A1(b_11_), .A2(n13773), .A3(a_17_), .ZN(n13772) );
  INV_X1 U13805 ( .A(n13774), .ZN(n13773) );
  NOR2_X1 U13806 ( .A1(n13672), .A2(n13671), .ZN(n13774) );
  NAND2_X1 U13807 ( .A1(n13671), .A2(n13672), .ZN(n13771) );
  NAND2_X1 U13808 ( .A1(n13668), .A2(n13775), .ZN(n13672) );
  NAND2_X1 U13809 ( .A1(n13667), .A2(n13669), .ZN(n13775) );
  NAND2_X1 U13810 ( .A1(n13776), .A2(n13777), .ZN(n13669) );
  NAND2_X1 U13811 ( .A1(a_18_), .A2(b_11_), .ZN(n13777) );
  XNOR2_X1 U13812 ( .A(n13778), .B(n13779), .ZN(n13667) );
  XNOR2_X1 U13813 ( .A(n13780), .B(n13781), .ZN(n13779) );
  NAND2_X1 U13814 ( .A1(a_18_), .A2(n13782), .ZN(n13668) );
  INV_X1 U13815 ( .A(n13776), .ZN(n13782) );
  NOR2_X1 U13816 ( .A1(n13783), .A2(n13784), .ZN(n13776) );
  NOR2_X1 U13817 ( .A1(n13665), .A2(n13785), .ZN(n13784) );
  NOR2_X1 U13818 ( .A1(n13664), .A2(n13662), .ZN(n13785) );
  NAND2_X1 U13819 ( .A1(b_11_), .A2(a_19_), .ZN(n13665) );
  INV_X1 U13820 ( .A(n13786), .ZN(n13783) );
  NAND2_X1 U13821 ( .A1(n13662), .A2(n13664), .ZN(n13786) );
  NAND2_X1 U13822 ( .A1(n13787), .A2(n13788), .ZN(n13664) );
  NAND2_X1 U13823 ( .A1(n13661), .A2(n13789), .ZN(n13788) );
  INV_X1 U13824 ( .A(n13790), .ZN(n13789) );
  NOR2_X1 U13825 ( .A1(n13660), .A2(n13659), .ZN(n13790) );
  NOR2_X1 U13826 ( .A1(n9047), .A2(n13332), .ZN(n13661) );
  NAND2_X1 U13827 ( .A1(n13659), .A2(n13660), .ZN(n13787) );
  NAND2_X1 U13828 ( .A1(n13791), .A2(n13792), .ZN(n13660) );
  NAND2_X1 U13829 ( .A1(n13657), .A2(n13793), .ZN(n13792) );
  INV_X1 U13830 ( .A(n13794), .ZN(n13793) );
  NOR2_X1 U13831 ( .A1(n13656), .A2(n13655), .ZN(n13794) );
  NOR2_X1 U13832 ( .A1(n8759), .A2(n13332), .ZN(n13657) );
  NAND2_X1 U13833 ( .A1(n13655), .A2(n13656), .ZN(n13791) );
  NAND2_X1 U13834 ( .A1(n13795), .A2(n13796), .ZN(n13656) );
  NAND2_X1 U13835 ( .A1(n13653), .A2(n13797), .ZN(n13796) );
  INV_X1 U13836 ( .A(n13798), .ZN(n13797) );
  NOR2_X1 U13837 ( .A1(n13652), .A2(n13650), .ZN(n13798) );
  NOR2_X1 U13838 ( .A1(n12296), .A2(n13332), .ZN(n13653) );
  NAND2_X1 U13839 ( .A1(n13650), .A2(n13652), .ZN(n13795) );
  NAND2_X1 U13840 ( .A1(n13799), .A2(n13800), .ZN(n13652) );
  NAND2_X1 U13841 ( .A1(n13649), .A2(n13801), .ZN(n13800) );
  INV_X1 U13842 ( .A(n13802), .ZN(n13801) );
  NOR2_X1 U13843 ( .A1(n13648), .A2(n13647), .ZN(n13802) );
  NOR2_X1 U13844 ( .A1(n12301), .A2(n13332), .ZN(n13649) );
  NAND2_X1 U13845 ( .A1(n13647), .A2(n13648), .ZN(n13799) );
  NAND2_X1 U13846 ( .A1(n13803), .A2(n13804), .ZN(n13648) );
  NAND2_X1 U13847 ( .A1(n13645), .A2(n13805), .ZN(n13804) );
  NAND2_X1 U13848 ( .A1(n13644), .A2(n13643), .ZN(n13805) );
  NOR2_X1 U13849 ( .A1(n8779), .A2(n13332), .ZN(n13645) );
  INV_X1 U13850 ( .A(n13806), .ZN(n13803) );
  NOR2_X1 U13851 ( .A1(n13643), .A2(n13644), .ZN(n13806) );
  NOR2_X1 U13852 ( .A1(n13807), .A2(n13808), .ZN(n13644) );
  INV_X1 U13853 ( .A(n13809), .ZN(n13808) );
  NAND2_X1 U13854 ( .A1(n13641), .A2(n13810), .ZN(n13809) );
  NAND2_X1 U13855 ( .A1(n13638), .A2(n13640), .ZN(n13810) );
  NOR2_X1 U13856 ( .A1(n8788), .A2(n13332), .ZN(n13641) );
  NOR2_X1 U13857 ( .A1(n13640), .A2(n13638), .ZN(n13807) );
  XNOR2_X1 U13858 ( .A(n13811), .B(n13812), .ZN(n13638) );
  XNOR2_X1 U13859 ( .A(n13813), .B(n13814), .ZN(n13812) );
  NAND2_X1 U13860 ( .A1(n13815), .A2(n13816), .ZN(n13640) );
  NAND2_X1 U13861 ( .A1(n13599), .A2(n13817), .ZN(n13816) );
  INV_X1 U13862 ( .A(n13818), .ZN(n13817) );
  NOR2_X1 U13863 ( .A1(n13602), .A2(n13601), .ZN(n13818) );
  XNOR2_X1 U13864 ( .A(n13819), .B(n13820), .ZN(n13599) );
  XOR2_X1 U13865 ( .A(n13821), .B(n13822), .Z(n13819) );
  NAND2_X1 U13866 ( .A1(n13601), .A2(n13602), .ZN(n13815) );
  NAND2_X1 U13867 ( .A1(a_26_), .A2(b_11_), .ZN(n13602) );
  NOR2_X1 U13868 ( .A1(n13823), .A2(n13824), .ZN(n13601) );
  INV_X1 U13869 ( .A(n13825), .ZN(n13824) );
  NAND2_X1 U13870 ( .A1(n13608), .A2(n13826), .ZN(n13825) );
  NAND2_X1 U13871 ( .A1(n13609), .A2(n13607), .ZN(n13826) );
  NOR2_X1 U13872 ( .A1(n8797), .A2(n13332), .ZN(n13608) );
  NOR2_X1 U13873 ( .A1(n13607), .A2(n13609), .ZN(n13823) );
  NOR2_X1 U13874 ( .A1(n13827), .A2(n13828), .ZN(n13609) );
  INV_X1 U13875 ( .A(n13829), .ZN(n13828) );
  NAND2_X1 U13876 ( .A1(n13636), .A2(n13830), .ZN(n13829) );
  NAND2_X1 U13877 ( .A1(n13637), .A2(n13635), .ZN(n13830) );
  NOR2_X1 U13878 ( .A1(n8314), .A2(n13332), .ZN(n13636) );
  NOR2_X1 U13879 ( .A1(n13635), .A2(n13637), .ZN(n13827) );
  NOR2_X1 U13880 ( .A1(n13831), .A2(n13832), .ZN(n13637) );
  INV_X1 U13881 ( .A(n13833), .ZN(n13832) );
  NAND2_X1 U13882 ( .A1(n13631), .A2(n13834), .ZN(n13833) );
  NAND2_X1 U13883 ( .A1(n13835), .A2(n13633), .ZN(n13834) );
  NOR2_X1 U13884 ( .A1(n9098), .A2(n13332), .ZN(n13631) );
  NOR2_X1 U13885 ( .A1(n13633), .A2(n13835), .ZN(n13831) );
  INV_X1 U13886 ( .A(n13632), .ZN(n13835) );
  NAND2_X1 U13887 ( .A1(n13836), .A2(n13837), .ZN(n13632) );
  NAND2_X1 U13888 ( .A1(b_10_), .A2(n13838), .ZN(n13837) );
  NAND2_X1 U13889 ( .A1(n8303), .A2(n13839), .ZN(n13838) );
  NAND2_X1 U13890 ( .A1(a_30_), .A2(n13840), .ZN(n13839) );
  NAND2_X1 U13891 ( .A1(b_9_), .A2(n13841), .ZN(n13836) );
  NAND2_X1 U13892 ( .A1(n8299), .A2(n13842), .ZN(n13841) );
  NAND2_X1 U13893 ( .A1(a_31_), .A2(n13629), .ZN(n13842) );
  NAND3_X1 U13894 ( .A1(n9106), .A2(b_11_), .A3(b_10_), .ZN(n13633) );
  XNOR2_X1 U13895 ( .A(n13843), .B(n13844), .ZN(n13635) );
  XOR2_X1 U13896 ( .A(n13845), .B(n13846), .Z(n13843) );
  XNOR2_X1 U13897 ( .A(n13847), .B(n13848), .ZN(n13607) );
  XOR2_X1 U13898 ( .A(n13849), .B(n13850), .Z(n13847) );
  XOR2_X1 U13899 ( .A(n13851), .B(n13852), .Z(n13643) );
  XNOR2_X1 U13900 ( .A(n13853), .B(n13854), .ZN(n13852) );
  XOR2_X1 U13901 ( .A(n13855), .B(n13856), .Z(n13647) );
  XOR2_X1 U13902 ( .A(n13857), .B(n13858), .Z(n13855) );
  XOR2_X1 U13903 ( .A(n13859), .B(n13860), .Z(n13650) );
  XOR2_X1 U13904 ( .A(n13861), .B(n13862), .Z(n13859) );
  XNOR2_X1 U13905 ( .A(n13863), .B(n13864), .ZN(n13655) );
  XNOR2_X1 U13906 ( .A(n13865), .B(n13866), .ZN(n13864) );
  XOR2_X1 U13907 ( .A(n13867), .B(n13868), .Z(n13659) );
  XOR2_X1 U13908 ( .A(n13869), .B(n13870), .Z(n13867) );
  NOR2_X1 U13909 ( .A1(n8759), .A2(n13629), .ZN(n13870) );
  XNOR2_X1 U13910 ( .A(n13871), .B(n13872), .ZN(n13662) );
  XNOR2_X1 U13911 ( .A(n13873), .B(n13874), .ZN(n13871) );
  NOR2_X1 U13912 ( .A1(n9047), .A2(n13629), .ZN(n13874) );
  XNOR2_X1 U13913 ( .A(n13875), .B(n13876), .ZN(n13671) );
  XOR2_X1 U13914 ( .A(n13877), .B(n13878), .Z(n13876) );
  NAND2_X1 U13915 ( .A1(a_18_), .A2(b_10_), .ZN(n13878) );
  XNOR2_X1 U13916 ( .A(n13879), .B(n13880), .ZN(n13674) );
  NAND2_X1 U13917 ( .A1(n13881), .A2(n13882), .ZN(n13879) );
  XNOR2_X1 U13918 ( .A(n13883), .B(n13884), .ZN(n13551) );
  NAND2_X1 U13919 ( .A1(n13885), .A2(n13886), .ZN(n13883) );
  XOR2_X1 U13920 ( .A(n13887), .B(n13888), .Z(n13542) );
  NAND2_X1 U13921 ( .A1(n13889), .A2(n13890), .ZN(n13887) );
  XOR2_X1 U13922 ( .A(n13891), .B(n13892), .Z(n13678) );
  XOR2_X1 U13923 ( .A(n13893), .B(n13894), .Z(n13892) );
  NAND2_X1 U13924 ( .A1(a_14_), .A2(b_10_), .ZN(n13894) );
  XOR2_X1 U13925 ( .A(n13895), .B(n13896), .Z(n13531) );
  NAND2_X1 U13926 ( .A1(n13897), .A2(n13898), .ZN(n13895) );
  XNOR2_X1 U13927 ( .A(n13899), .B(n13900), .ZN(n13507) );
  XOR2_X1 U13928 ( .A(n13901), .B(n13902), .Z(n13899) );
  XNOR2_X1 U13929 ( .A(n13903), .B(n13904), .ZN(n13498) );
  NAND2_X1 U13930 ( .A1(n13905), .A2(n13906), .ZN(n13903) );
  XNOR2_X1 U13931 ( .A(n13907), .B(n13908), .ZN(n13491) );
  XOR2_X1 U13932 ( .A(n13909), .B(n13910), .Z(n13907) );
  XNOR2_X1 U13933 ( .A(n13911), .B(n13912), .ZN(n13482) );
  XNOR2_X1 U13934 ( .A(n13913), .B(n13914), .ZN(n13912) );
  XOR2_X1 U13935 ( .A(n13915), .B(n13916), .Z(n13475) );
  XOR2_X1 U13936 ( .A(n13917), .B(n13918), .Z(n13915) );
  XNOR2_X1 U13937 ( .A(n13919), .B(n13920), .ZN(n13466) );
  XOR2_X1 U13938 ( .A(n13921), .B(n13922), .Z(n13919) );
  XOR2_X1 U13939 ( .A(n13923), .B(n13924), .Z(n13458) );
  XOR2_X1 U13940 ( .A(n13925), .B(n13926), .Z(n13923) );
  XOR2_X1 U13941 ( .A(n13927), .B(n13928), .Z(n13682) );
  XOR2_X1 U13942 ( .A(n13929), .B(n13930), .Z(n13927) );
  XNOR2_X1 U13943 ( .A(n13931), .B(n13932), .ZN(n13686) );
  XOR2_X1 U13944 ( .A(n13933), .B(n13934), .Z(n13931) );
  XNOR2_X1 U13945 ( .A(n13935), .B(n13936), .ZN(n13691) );
  XOR2_X1 U13946 ( .A(n13937), .B(n13938), .Z(n13935) );
  XOR2_X1 U13947 ( .A(n13939), .B(n13940), .Z(n13444) );
  XNOR2_X1 U13948 ( .A(n13941), .B(n13942), .ZN(n13939) );
  XNOR2_X1 U13949 ( .A(n8279), .B(n8280), .ZN(n8554) );
  NAND3_X1 U13950 ( .A1(n8280), .A2(n8279), .A3(n8277), .ZN(n8281) );
  NOR2_X1 U13951 ( .A1(n13943), .A2(n8583), .ZN(n8277) );
  NOR2_X1 U13952 ( .A1(n13944), .A2(n13945), .ZN(n8583) );
  INV_X1 U13953 ( .A(n13946), .ZN(n13943) );
  NAND2_X1 U13954 ( .A1(n13945), .A2(n13944), .ZN(n13946) );
  XOR2_X1 U13955 ( .A(n13947), .B(n13948), .Z(n13944) );
  XNOR2_X1 U13956 ( .A(n13949), .B(n13950), .ZN(n13947) );
  NOR2_X1 U13957 ( .A1(n13951), .A2(n13952), .ZN(n13945) );
  INV_X1 U13958 ( .A(n13953), .ZN(n13952) );
  NAND3_X1 U13959 ( .A1(b_9_), .A2(n13954), .A3(a_0_), .ZN(n13953) );
  NAND2_X1 U13960 ( .A1(n13955), .A2(n13956), .ZN(n13954) );
  NOR2_X1 U13961 ( .A1(n13955), .A2(n13956), .ZN(n13951) );
  NAND2_X1 U13962 ( .A1(n13957), .A2(n13958), .ZN(n8279) );
  NAND2_X1 U13963 ( .A1(n13942), .A2(n13959), .ZN(n13958) );
  INV_X1 U13964 ( .A(n13960), .ZN(n13959) );
  NOR2_X1 U13965 ( .A1(n13940), .A2(n13941), .ZN(n13960) );
  NOR2_X1 U13966 ( .A1(n8457), .A2(n13629), .ZN(n13942) );
  NAND2_X1 U13967 ( .A1(n13940), .A2(n13941), .ZN(n13957) );
  NAND2_X1 U13968 ( .A1(n13961), .A2(n13962), .ZN(n13941) );
  NAND2_X1 U13969 ( .A1(n13938), .A2(n13963), .ZN(n13962) );
  INV_X1 U13970 ( .A(n13964), .ZN(n13963) );
  NOR2_X1 U13971 ( .A1(n13936), .A2(n13937), .ZN(n13964) );
  NOR2_X1 U13972 ( .A1(n8569), .A2(n13629), .ZN(n13938) );
  NAND2_X1 U13973 ( .A1(n13936), .A2(n13937), .ZN(n13961) );
  NAND2_X1 U13974 ( .A1(n13965), .A2(n13966), .ZN(n13937) );
  NAND2_X1 U13975 ( .A1(n13934), .A2(n13967), .ZN(n13966) );
  INV_X1 U13976 ( .A(n13968), .ZN(n13967) );
  NOR2_X1 U13977 ( .A1(n13932), .A2(n13933), .ZN(n13968) );
  NOR2_X1 U13978 ( .A1(n8448), .A2(n13629), .ZN(n13934) );
  NAND2_X1 U13979 ( .A1(n13932), .A2(n13933), .ZN(n13965) );
  NAND2_X1 U13980 ( .A1(n13969), .A2(n13970), .ZN(n13933) );
  NAND2_X1 U13981 ( .A1(n13930), .A2(n13971), .ZN(n13970) );
  INV_X1 U13982 ( .A(n13972), .ZN(n13971) );
  NOR2_X1 U13983 ( .A1(n13928), .A2(n13929), .ZN(n13972) );
  NOR2_X1 U13984 ( .A1(n8900), .A2(n13629), .ZN(n13930) );
  NAND2_X1 U13985 ( .A1(n13928), .A2(n13929), .ZN(n13969) );
  NAND2_X1 U13986 ( .A1(n13973), .A2(n13974), .ZN(n13929) );
  NAND2_X1 U13987 ( .A1(n13926), .A2(n13975), .ZN(n13974) );
  INV_X1 U13988 ( .A(n13976), .ZN(n13975) );
  NOR2_X1 U13989 ( .A1(n13924), .A2(n13925), .ZN(n13976) );
  NOR2_X1 U13990 ( .A1(n8439), .A2(n13629), .ZN(n13926) );
  NAND2_X1 U13991 ( .A1(n13924), .A2(n13925), .ZN(n13973) );
  NAND2_X1 U13992 ( .A1(n13977), .A2(n13978), .ZN(n13925) );
  NAND2_X1 U13993 ( .A1(n13922), .A2(n13979), .ZN(n13978) );
  INV_X1 U13994 ( .A(n13980), .ZN(n13979) );
  NOR2_X1 U13995 ( .A1(n13920), .A2(n13921), .ZN(n13980) );
  NOR2_X1 U13996 ( .A1(n8938), .A2(n13629), .ZN(n13922) );
  NAND2_X1 U13997 ( .A1(n13920), .A2(n13921), .ZN(n13977) );
  NAND2_X1 U13998 ( .A1(n13981), .A2(n13982), .ZN(n13921) );
  NAND2_X1 U13999 ( .A1(n13918), .A2(n13983), .ZN(n13982) );
  INV_X1 U14000 ( .A(n13984), .ZN(n13983) );
  NOR2_X1 U14001 ( .A1(n13916), .A2(n13917), .ZN(n13984) );
  NOR2_X1 U14002 ( .A1(n8430), .A2(n13629), .ZN(n13918) );
  NAND2_X1 U14003 ( .A1(n13916), .A2(n13917), .ZN(n13981) );
  NAND2_X1 U14004 ( .A1(n13985), .A2(n13986), .ZN(n13917) );
  NAND2_X1 U14005 ( .A1(n13914), .A2(n13987), .ZN(n13986) );
  NAND2_X1 U14006 ( .A1(n13911), .A2(n13913), .ZN(n13987) );
  NOR2_X1 U14007 ( .A1(n8425), .A2(n13629), .ZN(n13914) );
  INV_X1 U14008 ( .A(n13988), .ZN(n13985) );
  NOR2_X1 U14009 ( .A1(n13913), .A2(n13911), .ZN(n13988) );
  XOR2_X1 U14010 ( .A(n13989), .B(n13990), .Z(n13911) );
  XOR2_X1 U14011 ( .A(n13991), .B(n13992), .Z(n13990) );
  NAND2_X1 U14012 ( .A1(a_8_), .A2(b_9_), .ZN(n13992) );
  NAND2_X1 U14013 ( .A1(n13993), .A2(n13994), .ZN(n13913) );
  NAND2_X1 U14014 ( .A1(n13908), .A2(n13995), .ZN(n13994) );
  NAND2_X1 U14015 ( .A1(n13910), .A2(n13909), .ZN(n13995) );
  XNOR2_X1 U14016 ( .A(n13996), .B(n13997), .ZN(n13908) );
  XNOR2_X1 U14017 ( .A(n13998), .B(n13999), .ZN(n13997) );
  INV_X1 U14018 ( .A(n14000), .ZN(n13993) );
  NOR2_X1 U14019 ( .A1(n13909), .A2(n13910), .ZN(n14000) );
  NOR2_X1 U14020 ( .A1(n8968), .A2(n13629), .ZN(n13910) );
  NAND2_X1 U14021 ( .A1(n13905), .A2(n14001), .ZN(n13909) );
  NAND2_X1 U14022 ( .A1(n13904), .A2(n13906), .ZN(n14001) );
  NAND2_X1 U14023 ( .A1(n14002), .A2(n14003), .ZN(n13906) );
  NAND2_X1 U14024 ( .A1(a_9_), .A2(b_10_), .ZN(n14003) );
  INV_X1 U14025 ( .A(n14004), .ZN(n14002) );
  XNOR2_X1 U14026 ( .A(n14005), .B(n14006), .ZN(n13904) );
  XOR2_X1 U14027 ( .A(n14007), .B(n14008), .Z(n14006) );
  NAND2_X1 U14028 ( .A1(a_10_), .A2(b_9_), .ZN(n14008) );
  NAND2_X1 U14029 ( .A1(a_9_), .A2(n14004), .ZN(n13905) );
  NAND2_X1 U14030 ( .A1(n14009), .A2(n14010), .ZN(n14004) );
  NAND2_X1 U14031 ( .A1(n13902), .A2(n14011), .ZN(n14010) );
  INV_X1 U14032 ( .A(n14012), .ZN(n14011) );
  NOR2_X1 U14033 ( .A1(n13901), .A2(n13900), .ZN(n14012) );
  NAND2_X1 U14034 ( .A1(n13900), .A2(n13901), .ZN(n14009) );
  NAND2_X1 U14035 ( .A1(n13740), .A2(n14013), .ZN(n13901) );
  NAND2_X1 U14036 ( .A1(n13739), .A2(n13741), .ZN(n14013) );
  NAND2_X1 U14037 ( .A1(n14014), .A2(n14015), .ZN(n13741) );
  NAND2_X1 U14038 ( .A1(a_11_), .A2(b_10_), .ZN(n14015) );
  XNOR2_X1 U14039 ( .A(n14016), .B(n14017), .ZN(n13739) );
  XOR2_X1 U14040 ( .A(n14018), .B(n14019), .Z(n14017) );
  NAND2_X1 U14041 ( .A1(a_12_), .A2(b_9_), .ZN(n14019) );
  INV_X1 U14042 ( .A(n14020), .ZN(n13740) );
  NOR2_X1 U14043 ( .A1(n8867), .A2(n14014), .ZN(n14020) );
  NOR2_X1 U14044 ( .A1(n14021), .A2(n14022), .ZN(n14014) );
  NOR3_X1 U14045 ( .A1(n13629), .A2(n14023), .A3(n8393), .ZN(n14022) );
  NOR2_X1 U14046 ( .A1(n13748), .A2(n13747), .ZN(n14023) );
  INV_X1 U14047 ( .A(n14024), .ZN(n14021) );
  NAND2_X1 U14048 ( .A1(n13747), .A2(n13748), .ZN(n14024) );
  NAND2_X1 U14049 ( .A1(n13897), .A2(n14025), .ZN(n13748) );
  NAND2_X1 U14050 ( .A1(n13896), .A2(n13898), .ZN(n14025) );
  NAND2_X1 U14051 ( .A1(n14026), .A2(n14027), .ZN(n13898) );
  NAND2_X1 U14052 ( .A1(a_13_), .A2(b_10_), .ZN(n14027) );
  INV_X1 U14053 ( .A(n14028), .ZN(n14026) );
  XOR2_X1 U14054 ( .A(n14029), .B(n14030), .Z(n13896) );
  XNOR2_X1 U14055 ( .A(n14031), .B(n14032), .ZN(n14030) );
  NAND2_X1 U14056 ( .A1(a_14_), .A2(b_9_), .ZN(n14032) );
  NAND2_X1 U14057 ( .A1(a_13_), .A2(n14028), .ZN(n13897) );
  NAND2_X1 U14058 ( .A1(n14033), .A2(n14034), .ZN(n14028) );
  INV_X1 U14059 ( .A(n14035), .ZN(n14034) );
  NOR3_X1 U14060 ( .A1(n13629), .A2(n14036), .A3(n9262), .ZN(n14035) );
  NOR2_X1 U14061 ( .A1(n13891), .A2(n13893), .ZN(n14036) );
  NAND2_X1 U14062 ( .A1(n13891), .A2(n13893), .ZN(n14033) );
  NAND2_X1 U14063 ( .A1(n13889), .A2(n14037), .ZN(n13893) );
  NAND2_X1 U14064 ( .A1(n13888), .A2(n13890), .ZN(n14037) );
  NAND2_X1 U14065 ( .A1(n14038), .A2(n14039), .ZN(n13890) );
  NAND2_X1 U14066 ( .A1(a_15_), .A2(b_10_), .ZN(n14039) );
  INV_X1 U14067 ( .A(n14040), .ZN(n14038) );
  XOR2_X1 U14068 ( .A(n14041), .B(n14042), .Z(n13888) );
  XNOR2_X1 U14069 ( .A(n14043), .B(n14044), .ZN(n14042) );
  NAND2_X1 U14070 ( .A1(a_16_), .A2(b_9_), .ZN(n14044) );
  NAND2_X1 U14071 ( .A1(a_15_), .A2(n14040), .ZN(n13889) );
  NAND2_X1 U14072 ( .A1(n13885), .A2(n14045), .ZN(n14040) );
  NAND2_X1 U14073 ( .A1(n13884), .A2(n13886), .ZN(n14045) );
  NAND2_X1 U14074 ( .A1(n14046), .A2(n14047), .ZN(n13886) );
  NAND2_X1 U14075 ( .A1(a_16_), .A2(b_10_), .ZN(n14047) );
  INV_X1 U14076 ( .A(n14048), .ZN(n14046) );
  XOR2_X1 U14077 ( .A(n14049), .B(n14050), .Z(n13884) );
  XOR2_X1 U14078 ( .A(n14051), .B(n14052), .Z(n14049) );
  NOR2_X1 U14079 ( .A1(n13840), .A2(n8371), .ZN(n14052) );
  NAND2_X1 U14080 ( .A1(a_16_), .A2(n14048), .ZN(n13885) );
  NAND2_X1 U14081 ( .A1(n13881), .A2(n14053), .ZN(n14048) );
  NAND2_X1 U14082 ( .A1(n13880), .A2(n13882), .ZN(n14053) );
  NAND2_X1 U14083 ( .A1(n14054), .A2(n14055), .ZN(n13882) );
  NAND2_X1 U14084 ( .A1(a_17_), .A2(b_10_), .ZN(n14055) );
  XNOR2_X1 U14085 ( .A(n14056), .B(n14057), .ZN(n13880) );
  XOR2_X1 U14086 ( .A(n14058), .B(n14059), .Z(n14057) );
  NAND2_X1 U14087 ( .A1(a_18_), .A2(b_9_), .ZN(n14059) );
  INV_X1 U14088 ( .A(n14060), .ZN(n13881) );
  NOR2_X1 U14089 ( .A1(n8371), .A2(n14054), .ZN(n14060) );
  NOR2_X1 U14090 ( .A1(n14061), .A2(n14062), .ZN(n14054) );
  NOR3_X1 U14091 ( .A1(n13629), .A2(n14063), .A3(n9291), .ZN(n14062) );
  NOR2_X1 U14092 ( .A1(n13877), .A2(n13875), .ZN(n14063) );
  INV_X1 U14093 ( .A(n14064), .ZN(n14061) );
  NAND2_X1 U14094 ( .A1(n13875), .A2(n13877), .ZN(n14064) );
  NAND2_X1 U14095 ( .A1(n14065), .A2(n14066), .ZN(n13877) );
  NAND2_X1 U14096 ( .A1(n13781), .A2(n14067), .ZN(n14066) );
  INV_X1 U14097 ( .A(n14068), .ZN(n14067) );
  NOR2_X1 U14098 ( .A1(n13778), .A2(n13780), .ZN(n14068) );
  NOR2_X1 U14099 ( .A1(n13629), .A2(n8742), .ZN(n13781) );
  NAND2_X1 U14100 ( .A1(n13778), .A2(n13780), .ZN(n14065) );
  NAND2_X1 U14101 ( .A1(n14069), .A2(n14070), .ZN(n13780) );
  NAND3_X1 U14102 ( .A1(a_20_), .A2(n14071), .A3(b_10_), .ZN(n14070) );
  NAND2_X1 U14103 ( .A1(n13873), .A2(n13872), .ZN(n14071) );
  INV_X1 U14104 ( .A(n14072), .ZN(n14069) );
  NOR2_X1 U14105 ( .A1(n13872), .A2(n13873), .ZN(n14072) );
  NOR2_X1 U14106 ( .A1(n14073), .A2(n14074), .ZN(n13873) );
  NOR3_X1 U14107 ( .A1(n8759), .A2(n14075), .A3(n13629), .ZN(n14074) );
  NOR2_X1 U14108 ( .A1(n13869), .A2(n13868), .ZN(n14075) );
  INV_X1 U14109 ( .A(n14076), .ZN(n14073) );
  NAND2_X1 U14110 ( .A1(n13868), .A2(n13869), .ZN(n14076) );
  NAND2_X1 U14111 ( .A1(n14077), .A2(n14078), .ZN(n13869) );
  NAND2_X1 U14112 ( .A1(n13866), .A2(n14079), .ZN(n14078) );
  INV_X1 U14113 ( .A(n14080), .ZN(n14079) );
  NOR2_X1 U14114 ( .A1(n13863), .A2(n13865), .ZN(n14080) );
  NOR2_X1 U14115 ( .A1(n13629), .A2(n12296), .ZN(n13866) );
  NAND2_X1 U14116 ( .A1(n13863), .A2(n13865), .ZN(n14077) );
  NAND2_X1 U14117 ( .A1(n14081), .A2(n14082), .ZN(n13865) );
  NAND2_X1 U14118 ( .A1(n13862), .A2(n14083), .ZN(n14082) );
  INV_X1 U14119 ( .A(n14084), .ZN(n14083) );
  NOR2_X1 U14120 ( .A1(n13861), .A2(n13860), .ZN(n14084) );
  NOR2_X1 U14121 ( .A1(n13629), .A2(n12301), .ZN(n13862) );
  NAND2_X1 U14122 ( .A1(n13860), .A2(n13861), .ZN(n14081) );
  NAND2_X1 U14123 ( .A1(n14085), .A2(n14086), .ZN(n13861) );
  NAND2_X1 U14124 ( .A1(n13858), .A2(n14087), .ZN(n14086) );
  INV_X1 U14125 ( .A(n14088), .ZN(n14087) );
  NOR2_X1 U14126 ( .A1(n13856), .A2(n13857), .ZN(n14088) );
  NOR2_X1 U14127 ( .A1(n13629), .A2(n8779), .ZN(n13858) );
  NAND2_X1 U14128 ( .A1(n13856), .A2(n13857), .ZN(n14085) );
  NAND2_X1 U14129 ( .A1(n14089), .A2(n14090), .ZN(n13857) );
  NAND2_X1 U14130 ( .A1(n13854), .A2(n14091), .ZN(n14090) );
  NAND2_X1 U14131 ( .A1(n13851), .A2(n13853), .ZN(n14091) );
  NOR2_X1 U14132 ( .A1(n13629), .A2(n8788), .ZN(n13854) );
  INV_X1 U14133 ( .A(n14092), .ZN(n14089) );
  NOR2_X1 U14134 ( .A1(n13853), .A2(n13851), .ZN(n14092) );
  XNOR2_X1 U14135 ( .A(n14093), .B(n14094), .ZN(n13851) );
  XNOR2_X1 U14136 ( .A(n14095), .B(n14096), .ZN(n14094) );
  NAND2_X1 U14137 ( .A1(n14097), .A2(n14098), .ZN(n13853) );
  NAND2_X1 U14138 ( .A1(n13811), .A2(n14099), .ZN(n14098) );
  NAND2_X1 U14139 ( .A1(n13814), .A2(n13813), .ZN(n14099) );
  XNOR2_X1 U14140 ( .A(n14100), .B(n14101), .ZN(n13811) );
  XOR2_X1 U14141 ( .A(n14102), .B(n14103), .Z(n14100) );
  INV_X1 U14142 ( .A(n14104), .ZN(n14097) );
  NOR2_X1 U14143 ( .A1(n13813), .A2(n13814), .ZN(n14104) );
  NOR2_X1 U14144 ( .A1(n9344), .A2(n13629), .ZN(n13814) );
  NAND2_X1 U14145 ( .A1(n14105), .A2(n14106), .ZN(n13813) );
  NAND2_X1 U14146 ( .A1(n13822), .A2(n14107), .ZN(n14106) );
  INV_X1 U14147 ( .A(n14108), .ZN(n14107) );
  NOR2_X1 U14148 ( .A1(n13820), .A2(n13821), .ZN(n14108) );
  NOR2_X1 U14149 ( .A1(n13629), .A2(n8797), .ZN(n13822) );
  NAND2_X1 U14150 ( .A1(n13820), .A2(n13821), .ZN(n14105) );
  NAND2_X1 U14151 ( .A1(n14109), .A2(n14110), .ZN(n13821) );
  NAND2_X1 U14152 ( .A1(n13849), .A2(n14111), .ZN(n14110) );
  INV_X1 U14153 ( .A(n14112), .ZN(n14111) );
  NOR2_X1 U14154 ( .A1(n13850), .A2(n13848), .ZN(n14112) );
  NOR2_X1 U14155 ( .A1(n13629), .A2(n8314), .ZN(n13849) );
  NAND2_X1 U14156 ( .A1(n13848), .A2(n13850), .ZN(n14109) );
  NAND2_X1 U14157 ( .A1(n14113), .A2(n14114), .ZN(n13850) );
  NAND2_X1 U14158 ( .A1(n13844), .A2(n14115), .ZN(n14114) );
  INV_X1 U14159 ( .A(n14116), .ZN(n14115) );
  NOR2_X1 U14160 ( .A1(n13845), .A2(n13846), .ZN(n14116) );
  NOR2_X1 U14161 ( .A1(n13629), .A2(n9098), .ZN(n13844) );
  NAND2_X1 U14162 ( .A1(n13846), .A2(n13845), .ZN(n14113) );
  NAND2_X1 U14163 ( .A1(n14117), .A2(n14118), .ZN(n13845) );
  NAND2_X1 U14164 ( .A1(b_8_), .A2(n14119), .ZN(n14118) );
  NAND2_X1 U14165 ( .A1(n8299), .A2(n14120), .ZN(n14119) );
  NAND2_X1 U14166 ( .A1(a_31_), .A2(n13840), .ZN(n14120) );
  NAND2_X1 U14167 ( .A1(b_9_), .A2(n14121), .ZN(n14117) );
  NAND2_X1 U14168 ( .A1(n8303), .A2(n14122), .ZN(n14121) );
  NAND2_X1 U14169 ( .A1(a_30_), .A2(n14123), .ZN(n14122) );
  NOR3_X1 U14170 ( .A1(n13629), .A2(n9631), .A3(n13840), .ZN(n13846) );
  XOR2_X1 U14171 ( .A(n14124), .B(n14125), .Z(n13848) );
  XOR2_X1 U14172 ( .A(n14126), .B(n14127), .Z(n14124) );
  XOR2_X1 U14173 ( .A(n14128), .B(n14129), .Z(n13820) );
  XOR2_X1 U14174 ( .A(n14130), .B(n14131), .Z(n14128) );
  XNOR2_X1 U14175 ( .A(n14132), .B(n14133), .ZN(n13856) );
  XNOR2_X1 U14176 ( .A(n14134), .B(n14135), .ZN(n14133) );
  XOR2_X1 U14177 ( .A(n14136), .B(n14137), .Z(n13860) );
  XOR2_X1 U14178 ( .A(n14138), .B(n14139), .Z(n14136) );
  XOR2_X1 U14179 ( .A(n14140), .B(n14141), .Z(n13863) );
  XOR2_X1 U14180 ( .A(n14142), .B(n14143), .Z(n14140) );
  XNOR2_X1 U14181 ( .A(n14144), .B(n14145), .ZN(n13868) );
  XNOR2_X1 U14182 ( .A(n14146), .B(n14147), .ZN(n14145) );
  XNOR2_X1 U14183 ( .A(n14148), .B(n14149), .ZN(n13872) );
  XOR2_X1 U14184 ( .A(n14150), .B(n14151), .Z(n14148) );
  XOR2_X1 U14185 ( .A(n14152), .B(n14153), .Z(n13778) );
  XOR2_X1 U14186 ( .A(n14154), .B(n14155), .Z(n14152) );
  NOR2_X1 U14187 ( .A1(n9047), .A2(n13840), .ZN(n14155) );
  XOR2_X1 U14188 ( .A(n14156), .B(n14157), .Z(n13875) );
  XNOR2_X1 U14189 ( .A(n14158), .B(n14159), .ZN(n14157) );
  NAND2_X1 U14190 ( .A1(b_9_), .A2(a_19_), .ZN(n14159) );
  XNOR2_X1 U14191 ( .A(n14160), .B(n14161), .ZN(n13891) );
  XNOR2_X1 U14192 ( .A(n14162), .B(n14163), .ZN(n14160) );
  NOR2_X1 U14193 ( .A1(n13840), .A2(n8850), .ZN(n14163) );
  XOR2_X1 U14194 ( .A(n14164), .B(n14165), .Z(n13747) );
  XOR2_X1 U14195 ( .A(n14166), .B(n14167), .Z(n14164) );
  NOR2_X1 U14196 ( .A1(n13840), .A2(n8996), .ZN(n14167) );
  XOR2_X1 U14197 ( .A(n14168), .B(n14169), .Z(n13900) );
  XOR2_X1 U14198 ( .A(n14170), .B(n14171), .Z(n14168) );
  NOR2_X1 U14199 ( .A1(n13840), .A2(n8867), .ZN(n14171) );
  XOR2_X1 U14200 ( .A(n14172), .B(n14173), .Z(n13916) );
  XNOR2_X1 U14201 ( .A(n14174), .B(n14175), .ZN(n14173) );
  NAND2_X1 U14202 ( .A1(a_7_), .A2(b_9_), .ZN(n14175) );
  XNOR2_X1 U14203 ( .A(n14176), .B(n14177), .ZN(n13920) );
  XNOR2_X1 U14204 ( .A(n14178), .B(n14179), .ZN(n14176) );
  NOR2_X1 U14205 ( .A1(n13840), .A2(n8430), .ZN(n14179) );
  XOR2_X1 U14206 ( .A(n14180), .B(n14181), .Z(n13924) );
  XNOR2_X1 U14207 ( .A(n14182), .B(n14183), .ZN(n14181) );
  NAND2_X1 U14208 ( .A1(a_5_), .A2(b_9_), .ZN(n14183) );
  XNOR2_X1 U14209 ( .A(n14184), .B(n14185), .ZN(n13928) );
  XNOR2_X1 U14210 ( .A(n14186), .B(n14187), .ZN(n14184) );
  NOR2_X1 U14211 ( .A1(n13840), .A2(n8439), .ZN(n14187) );
  XOR2_X1 U14212 ( .A(n14188), .B(n14189), .Z(n13932) );
  XNOR2_X1 U14213 ( .A(n14190), .B(n14191), .ZN(n14189) );
  NAND2_X1 U14214 ( .A1(a_3_), .A2(b_9_), .ZN(n14191) );
  XNOR2_X1 U14215 ( .A(n14192), .B(n14193), .ZN(n13936) );
  XNOR2_X1 U14216 ( .A(n14194), .B(n14195), .ZN(n14192) );
  NOR2_X1 U14217 ( .A1(n13840), .A2(n8448), .ZN(n14195) );
  XOR2_X1 U14218 ( .A(n14196), .B(n14197), .Z(n13940) );
  XNOR2_X1 U14219 ( .A(n14198), .B(n14199), .ZN(n14197) );
  NAND2_X1 U14220 ( .A1(a_1_), .A2(b_9_), .ZN(n14199) );
  XNOR2_X1 U14221 ( .A(n14200), .B(n13955), .ZN(n8280) );
  XNOR2_X1 U14222 ( .A(n14201), .B(n14202), .ZN(n13955) );
  XOR2_X1 U14223 ( .A(n14203), .B(n14204), .Z(n14201) );
  XNOR2_X1 U14224 ( .A(n13956), .B(n14205), .ZN(n14200) );
  NOR2_X1 U14225 ( .A1(n13840), .A2(n8457), .ZN(n14205) );
  NOR2_X1 U14226 ( .A1(n14206), .A2(n14207), .ZN(n13956) );
  INV_X1 U14227 ( .A(n14208), .ZN(n14207) );
  NAND3_X1 U14228 ( .A1(b_9_), .A2(n14209), .A3(a_1_), .ZN(n14208) );
  NAND2_X1 U14229 ( .A1(n14198), .A2(n14196), .ZN(n14209) );
  NOR2_X1 U14230 ( .A1(n14196), .A2(n14198), .ZN(n14206) );
  NOR2_X1 U14231 ( .A1(n14210), .A2(n14211), .ZN(n14198) );
  INV_X1 U14232 ( .A(n14212), .ZN(n14211) );
  NAND3_X1 U14233 ( .A1(b_9_), .A2(n14213), .A3(a_2_), .ZN(n14212) );
  NAND2_X1 U14234 ( .A1(n14194), .A2(n14193), .ZN(n14213) );
  NOR2_X1 U14235 ( .A1(n14193), .A2(n14194), .ZN(n14210) );
  NOR2_X1 U14236 ( .A1(n14214), .A2(n14215), .ZN(n14194) );
  NOR3_X1 U14237 ( .A1(n13840), .A2(n14216), .A3(n8900), .ZN(n14215) );
  INV_X1 U14238 ( .A(n14217), .ZN(n14216) );
  NAND2_X1 U14239 ( .A1(n14190), .A2(n14188), .ZN(n14217) );
  NOR2_X1 U14240 ( .A1(n14188), .A2(n14190), .ZN(n14214) );
  NOR2_X1 U14241 ( .A1(n14218), .A2(n14219), .ZN(n14190) );
  INV_X1 U14242 ( .A(n14220), .ZN(n14219) );
  NAND3_X1 U14243 ( .A1(b_9_), .A2(n14221), .A3(a_4_), .ZN(n14220) );
  NAND2_X1 U14244 ( .A1(n14186), .A2(n14185), .ZN(n14221) );
  NOR2_X1 U14245 ( .A1(n14185), .A2(n14186), .ZN(n14218) );
  NOR2_X1 U14246 ( .A1(n14222), .A2(n14223), .ZN(n14186) );
  NOR3_X1 U14247 ( .A1(n13840), .A2(n14224), .A3(n8938), .ZN(n14223) );
  INV_X1 U14248 ( .A(n14225), .ZN(n14224) );
  NAND2_X1 U14249 ( .A1(n14182), .A2(n14180), .ZN(n14225) );
  NOR2_X1 U14250 ( .A1(n14180), .A2(n14182), .ZN(n14222) );
  NOR2_X1 U14251 ( .A1(n14226), .A2(n14227), .ZN(n14182) );
  INV_X1 U14252 ( .A(n14228), .ZN(n14227) );
  NAND3_X1 U14253 ( .A1(b_9_), .A2(n14229), .A3(a_6_), .ZN(n14228) );
  NAND2_X1 U14254 ( .A1(n14178), .A2(n14177), .ZN(n14229) );
  NOR2_X1 U14255 ( .A1(n14177), .A2(n14178), .ZN(n14226) );
  NOR2_X1 U14256 ( .A1(n14230), .A2(n14231), .ZN(n14178) );
  INV_X1 U14257 ( .A(n14232), .ZN(n14231) );
  NAND3_X1 U14258 ( .A1(b_9_), .A2(n14233), .A3(a_7_), .ZN(n14232) );
  NAND2_X1 U14259 ( .A1(n14174), .A2(n14172), .ZN(n14233) );
  NOR2_X1 U14260 ( .A1(n14172), .A2(n14174), .ZN(n14230) );
  NOR2_X1 U14261 ( .A1(n14234), .A2(n14235), .ZN(n14174) );
  INV_X1 U14262 ( .A(n14236), .ZN(n14235) );
  NAND3_X1 U14263 ( .A1(b_9_), .A2(n14237), .A3(a_8_), .ZN(n14236) );
  NAND2_X1 U14264 ( .A1(n13989), .A2(n13991), .ZN(n14237) );
  NOR2_X1 U14265 ( .A1(n13991), .A2(n13989), .ZN(n14234) );
  XNOR2_X1 U14266 ( .A(n14238), .B(n14239), .ZN(n13989) );
  XOR2_X1 U14267 ( .A(n14240), .B(n14241), .Z(n14239) );
  NAND2_X1 U14268 ( .A1(n14242), .A2(n14243), .ZN(n13991) );
  NAND2_X1 U14269 ( .A1(n13996), .A2(n14244), .ZN(n14243) );
  NAND2_X1 U14270 ( .A1(n13999), .A2(n13998), .ZN(n14244) );
  XNOR2_X1 U14271 ( .A(n14245), .B(n14246), .ZN(n13996) );
  XOR2_X1 U14272 ( .A(n14247), .B(n14248), .Z(n14246) );
  NAND2_X1 U14273 ( .A1(n14249), .A2(n14250), .ZN(n14242) );
  INV_X1 U14274 ( .A(n13998), .ZN(n14249) );
  NAND2_X1 U14275 ( .A1(n14251), .A2(n14252), .ZN(n13998) );
  INV_X1 U14276 ( .A(n14253), .ZN(n14252) );
  NOR3_X1 U14277 ( .A1(n13840), .A2(n14254), .A3(n8402), .ZN(n14253) );
  NOR2_X1 U14278 ( .A1(n14005), .A2(n14007), .ZN(n14254) );
  NAND2_X1 U14279 ( .A1(n14005), .A2(n14007), .ZN(n14251) );
  NAND2_X1 U14280 ( .A1(n14255), .A2(n14256), .ZN(n14007) );
  NAND3_X1 U14281 ( .A1(b_9_), .A2(n14257), .A3(a_11_), .ZN(n14256) );
  INV_X1 U14282 ( .A(n14258), .ZN(n14257) );
  NOR2_X1 U14283 ( .A1(n14169), .A2(n14170), .ZN(n14258) );
  NAND2_X1 U14284 ( .A1(n14169), .A2(n14170), .ZN(n14255) );
  NAND2_X1 U14285 ( .A1(n14259), .A2(n14260), .ZN(n14170) );
  INV_X1 U14286 ( .A(n14261), .ZN(n14260) );
  NOR3_X1 U14287 ( .A1(n13840), .A2(n14262), .A3(n8393), .ZN(n14261) );
  NOR2_X1 U14288 ( .A1(n14016), .A2(n14018), .ZN(n14262) );
  NAND2_X1 U14289 ( .A1(n14016), .A2(n14018), .ZN(n14259) );
  NAND2_X1 U14290 ( .A1(n14263), .A2(n14264), .ZN(n14018) );
  NAND3_X1 U14291 ( .A1(b_9_), .A2(n14265), .A3(a_13_), .ZN(n14264) );
  INV_X1 U14292 ( .A(n14266), .ZN(n14265) );
  NOR2_X1 U14293 ( .A1(n14165), .A2(n14166), .ZN(n14266) );
  NAND2_X1 U14294 ( .A1(n14165), .A2(n14166), .ZN(n14263) );
  NAND2_X1 U14295 ( .A1(n14267), .A2(n14268), .ZN(n14166) );
  NAND3_X1 U14296 ( .A1(b_9_), .A2(n14269), .A3(a_14_), .ZN(n14268) );
  NAND2_X1 U14297 ( .A1(n14031), .A2(n14029), .ZN(n14269) );
  INV_X1 U14298 ( .A(n14270), .ZN(n14267) );
  NOR2_X1 U14299 ( .A1(n14029), .A2(n14031), .ZN(n14270) );
  NOR2_X1 U14300 ( .A1(n14271), .A2(n14272), .ZN(n14031) );
  INV_X1 U14301 ( .A(n14273), .ZN(n14272) );
  NAND3_X1 U14302 ( .A1(b_9_), .A2(n14274), .A3(a_15_), .ZN(n14273) );
  NAND2_X1 U14303 ( .A1(n14162), .A2(n14161), .ZN(n14274) );
  NOR2_X1 U14304 ( .A1(n14161), .A2(n14162), .ZN(n14271) );
  NOR2_X1 U14305 ( .A1(n14275), .A2(n14276), .ZN(n14162) );
  NOR3_X1 U14306 ( .A1(n13840), .A2(n14277), .A3(n8376), .ZN(n14276) );
  INV_X1 U14307 ( .A(n14278), .ZN(n14277) );
  NAND2_X1 U14308 ( .A1(n14043), .A2(n14041), .ZN(n14278) );
  NOR2_X1 U14309 ( .A1(n14041), .A2(n14043), .ZN(n14275) );
  NOR2_X1 U14310 ( .A1(n14279), .A2(n14280), .ZN(n14043) );
  NOR3_X1 U14311 ( .A1(n13840), .A2(n14281), .A3(n8371), .ZN(n14280) );
  NOR2_X1 U14312 ( .A1(n14050), .A2(n14051), .ZN(n14281) );
  INV_X1 U14313 ( .A(n14282), .ZN(n14279) );
  NAND2_X1 U14314 ( .A1(n14050), .A2(n14051), .ZN(n14282) );
  NAND2_X1 U14315 ( .A1(n14283), .A2(n14284), .ZN(n14051) );
  INV_X1 U14316 ( .A(n14285), .ZN(n14284) );
  NOR3_X1 U14317 ( .A1(n13840), .A2(n14286), .A3(n9291), .ZN(n14285) );
  NOR2_X1 U14318 ( .A1(n14058), .A2(n14056), .ZN(n14286) );
  NAND2_X1 U14319 ( .A1(n14056), .A2(n14058), .ZN(n14283) );
  NAND2_X1 U14320 ( .A1(n14287), .A2(n14288), .ZN(n14058) );
  NAND3_X1 U14321 ( .A1(a_19_), .A2(n14289), .A3(b_9_), .ZN(n14288) );
  NAND2_X1 U14322 ( .A1(n14156), .A2(n14158), .ZN(n14289) );
  INV_X1 U14323 ( .A(n14290), .ZN(n14287) );
  NOR2_X1 U14324 ( .A1(n14156), .A2(n14158), .ZN(n14290) );
  NOR2_X1 U14325 ( .A1(n14291), .A2(n14292), .ZN(n14158) );
  NOR3_X1 U14326 ( .A1(n9047), .A2(n14293), .A3(n13840), .ZN(n14292) );
  NOR2_X1 U14327 ( .A1(n14154), .A2(n14153), .ZN(n14293) );
  INV_X1 U14328 ( .A(n14294), .ZN(n14291) );
  NAND2_X1 U14329 ( .A1(n14153), .A2(n14154), .ZN(n14294) );
  NAND2_X1 U14330 ( .A1(n14295), .A2(n14296), .ZN(n14154) );
  NAND2_X1 U14331 ( .A1(n14151), .A2(n14297), .ZN(n14296) );
  INV_X1 U14332 ( .A(n14298), .ZN(n14297) );
  NOR2_X1 U14333 ( .A1(n14149), .A2(n14150), .ZN(n14298) );
  NOR2_X1 U14334 ( .A1(n13840), .A2(n8759), .ZN(n14151) );
  NAND2_X1 U14335 ( .A1(n14149), .A2(n14150), .ZN(n14295) );
  NAND2_X1 U14336 ( .A1(n14299), .A2(n14300), .ZN(n14150) );
  NAND2_X1 U14337 ( .A1(n14147), .A2(n14301), .ZN(n14300) );
  INV_X1 U14338 ( .A(n14302), .ZN(n14301) );
  NOR2_X1 U14339 ( .A1(n14144), .A2(n14146), .ZN(n14302) );
  NOR2_X1 U14340 ( .A1(n13840), .A2(n12296), .ZN(n14147) );
  NAND2_X1 U14341 ( .A1(n14144), .A2(n14146), .ZN(n14299) );
  NAND2_X1 U14342 ( .A1(n14303), .A2(n14304), .ZN(n14146) );
  NAND2_X1 U14343 ( .A1(n14143), .A2(n14305), .ZN(n14304) );
  INV_X1 U14344 ( .A(n14306), .ZN(n14305) );
  NOR2_X1 U14345 ( .A1(n14142), .A2(n14141), .ZN(n14306) );
  NOR2_X1 U14346 ( .A1(n13840), .A2(n12301), .ZN(n14143) );
  NAND2_X1 U14347 ( .A1(n14141), .A2(n14142), .ZN(n14303) );
  NAND2_X1 U14348 ( .A1(n14307), .A2(n14308), .ZN(n14142) );
  NAND2_X1 U14349 ( .A1(n14139), .A2(n14309), .ZN(n14308) );
  INV_X1 U14350 ( .A(n14310), .ZN(n14309) );
  NOR2_X1 U14351 ( .A1(n14137), .A2(n14138), .ZN(n14310) );
  NOR2_X1 U14352 ( .A1(n13840), .A2(n8779), .ZN(n14139) );
  NAND2_X1 U14353 ( .A1(n14137), .A2(n14138), .ZN(n14307) );
  NAND2_X1 U14354 ( .A1(n14311), .A2(n14312), .ZN(n14138) );
  NAND2_X1 U14355 ( .A1(n14135), .A2(n14313), .ZN(n14312) );
  NAND2_X1 U14356 ( .A1(n14132), .A2(n14134), .ZN(n14313) );
  NOR2_X1 U14357 ( .A1(n13840), .A2(n8788), .ZN(n14135) );
  INV_X1 U14358 ( .A(n14314), .ZN(n14311) );
  NOR2_X1 U14359 ( .A1(n14134), .A2(n14132), .ZN(n14314) );
  XNOR2_X1 U14360 ( .A(n14315), .B(n14316), .ZN(n14132) );
  XNOR2_X1 U14361 ( .A(n14317), .B(n14318), .ZN(n14316) );
  NAND2_X1 U14362 ( .A1(n14319), .A2(n14320), .ZN(n14134) );
  NAND2_X1 U14363 ( .A1(n14093), .A2(n14321), .ZN(n14320) );
  NAND2_X1 U14364 ( .A1(n14096), .A2(n14095), .ZN(n14321) );
  XNOR2_X1 U14365 ( .A(n14322), .B(n14323), .ZN(n14093) );
  XOR2_X1 U14366 ( .A(n14324), .B(n14325), .Z(n14322) );
  INV_X1 U14367 ( .A(n14326), .ZN(n14319) );
  NOR2_X1 U14368 ( .A1(n14095), .A2(n14096), .ZN(n14326) );
  NOR2_X1 U14369 ( .A1(n9344), .A2(n13840), .ZN(n14096) );
  NAND2_X1 U14370 ( .A1(n14327), .A2(n14328), .ZN(n14095) );
  NAND2_X1 U14371 ( .A1(n14103), .A2(n14329), .ZN(n14328) );
  INV_X1 U14372 ( .A(n14330), .ZN(n14329) );
  NOR2_X1 U14373 ( .A1(n14101), .A2(n14102), .ZN(n14330) );
  NOR2_X1 U14374 ( .A1(n13840), .A2(n8797), .ZN(n14103) );
  NAND2_X1 U14375 ( .A1(n14101), .A2(n14102), .ZN(n14327) );
  NAND2_X1 U14376 ( .A1(n14331), .A2(n14332), .ZN(n14102) );
  NAND2_X1 U14377 ( .A1(n14130), .A2(n14333), .ZN(n14332) );
  INV_X1 U14378 ( .A(n14334), .ZN(n14333) );
  NOR2_X1 U14379 ( .A1(n14131), .A2(n14129), .ZN(n14334) );
  NOR2_X1 U14380 ( .A1(n13840), .A2(n8314), .ZN(n14130) );
  NAND2_X1 U14381 ( .A1(n14129), .A2(n14131), .ZN(n14331) );
  NAND2_X1 U14382 ( .A1(n14335), .A2(n14336), .ZN(n14131) );
  NAND2_X1 U14383 ( .A1(n14125), .A2(n14337), .ZN(n14336) );
  INV_X1 U14384 ( .A(n14338), .ZN(n14337) );
  NOR2_X1 U14385 ( .A1(n14126), .A2(n14127), .ZN(n14338) );
  NOR2_X1 U14386 ( .A1(n13840), .A2(n9098), .ZN(n14125) );
  NAND2_X1 U14387 ( .A1(n14127), .A2(n14126), .ZN(n14335) );
  NAND2_X1 U14388 ( .A1(n14339), .A2(n14340), .ZN(n14126) );
  NAND2_X1 U14389 ( .A1(b_7_), .A2(n14341), .ZN(n14340) );
  NAND2_X1 U14390 ( .A1(n8299), .A2(n14342), .ZN(n14341) );
  NAND2_X1 U14391 ( .A1(a_31_), .A2(n14123), .ZN(n14342) );
  NAND2_X1 U14392 ( .A1(b_8_), .A2(n14343), .ZN(n14339) );
  NAND2_X1 U14393 ( .A1(n8303), .A2(n14344), .ZN(n14343) );
  NAND2_X1 U14394 ( .A1(a_30_), .A2(n14345), .ZN(n14344) );
  NOR3_X1 U14395 ( .A1(n13840), .A2(n9631), .A3(n14123), .ZN(n14127) );
  XOR2_X1 U14396 ( .A(n14346), .B(n14347), .Z(n14129) );
  XOR2_X1 U14397 ( .A(n14348), .B(n14349), .Z(n14346) );
  XOR2_X1 U14398 ( .A(n14350), .B(n14351), .Z(n14101) );
  XOR2_X1 U14399 ( .A(n14352), .B(n14353), .Z(n14350) );
  XNOR2_X1 U14400 ( .A(n14354), .B(n14355), .ZN(n14137) );
  XNOR2_X1 U14401 ( .A(n14356), .B(n14357), .ZN(n14355) );
  XOR2_X1 U14402 ( .A(n14358), .B(n14359), .Z(n14141) );
  XOR2_X1 U14403 ( .A(n14360), .B(n14361), .Z(n14358) );
  XOR2_X1 U14404 ( .A(n14362), .B(n14363), .Z(n14144) );
  XOR2_X1 U14405 ( .A(n14364), .B(n14365), .Z(n14362) );
  XNOR2_X1 U14406 ( .A(n14366), .B(n14367), .ZN(n14149) );
  XNOR2_X1 U14407 ( .A(n14368), .B(n14369), .ZN(n14367) );
  XNOR2_X1 U14408 ( .A(n14370), .B(n14371), .ZN(n14153) );
  XOR2_X1 U14409 ( .A(n14372), .B(n14373), .Z(n14371) );
  XOR2_X1 U14410 ( .A(n14374), .B(n14375), .Z(n14156) );
  XNOR2_X1 U14411 ( .A(n14376), .B(n14377), .ZN(n14374) );
  XNOR2_X1 U14412 ( .A(n14378), .B(n14379), .ZN(n14056) );
  XNOR2_X1 U14413 ( .A(n14380), .B(n14381), .ZN(n14379) );
  NAND2_X1 U14414 ( .A1(b_8_), .A2(a_19_), .ZN(n14381) );
  XNOR2_X1 U14415 ( .A(n14382), .B(n14383), .ZN(n14050) );
  NAND2_X1 U14416 ( .A1(n14384), .A2(n14385), .ZN(n14382) );
  XOR2_X1 U14417 ( .A(n14386), .B(n14387), .Z(n14041) );
  NAND2_X1 U14418 ( .A1(n14388), .A2(n14389), .ZN(n14386) );
  XOR2_X1 U14419 ( .A(n14390), .B(n14391), .Z(n14161) );
  NAND2_X1 U14420 ( .A1(n14392), .A2(n14393), .ZN(n14390) );
  XOR2_X1 U14421 ( .A(n14394), .B(n14395), .Z(n14029) );
  NAND2_X1 U14422 ( .A1(n14396), .A2(n14397), .ZN(n14394) );
  XNOR2_X1 U14423 ( .A(n14398), .B(n14399), .ZN(n14165) );
  NAND2_X1 U14424 ( .A1(n14400), .A2(n14401), .ZN(n14398) );
  XOR2_X1 U14425 ( .A(n14402), .B(n14403), .Z(n14016) );
  XNOR2_X1 U14426 ( .A(n14404), .B(n14405), .ZN(n14403) );
  XNOR2_X1 U14427 ( .A(n14406), .B(n14407), .ZN(n14169) );
  XNOR2_X1 U14428 ( .A(n14408), .B(n14409), .ZN(n14407) );
  XNOR2_X1 U14429 ( .A(n14410), .B(n14411), .ZN(n14005) );
  XNOR2_X1 U14430 ( .A(n14412), .B(n14413), .ZN(n14410) );
  XNOR2_X1 U14431 ( .A(n14414), .B(n14415), .ZN(n14172) );
  XNOR2_X1 U14432 ( .A(n14416), .B(n14417), .ZN(n14414) );
  XOR2_X1 U14433 ( .A(n14418), .B(n14419), .Z(n14177) );
  XNOR2_X1 U14434 ( .A(n14420), .B(n14421), .ZN(n14419) );
  XOR2_X1 U14435 ( .A(n14422), .B(n14423), .Z(n14180) );
  XOR2_X1 U14436 ( .A(n14424), .B(n14425), .Z(n14423) );
  XOR2_X1 U14437 ( .A(n14426), .B(n14427), .Z(n14185) );
  XNOR2_X1 U14438 ( .A(n14428), .B(n14429), .ZN(n14426) );
  XNOR2_X1 U14439 ( .A(n14430), .B(n14431), .ZN(n14188) );
  XNOR2_X1 U14440 ( .A(n14432), .B(n14433), .ZN(n14430) );
  XOR2_X1 U14441 ( .A(n14434), .B(n14435), .Z(n14193) );
  XNOR2_X1 U14442 ( .A(n14436), .B(n14437), .ZN(n14434) );
  XNOR2_X1 U14443 ( .A(n14438), .B(n14439), .ZN(n14196) );
  XOR2_X1 U14444 ( .A(n14440), .B(n14441), .Z(n14438) );
  XNOR2_X1 U14445 ( .A(n8292), .B(n8291), .ZN(n8283) );
  NAND3_X1 U14446 ( .A1(n8292), .A2(n8291), .A3(n8289), .ZN(n8293) );
  NOR2_X1 U14447 ( .A1(n14442), .A2(n8580), .ZN(n8289) );
  INV_X1 U14448 ( .A(n14443), .ZN(n8580) );
  NAND2_X1 U14449 ( .A1(n14444), .A2(n14445), .ZN(n14443) );
  NOR2_X1 U14450 ( .A1(n14445), .A2(n14444), .ZN(n14442) );
  XOR2_X1 U14451 ( .A(n14446), .B(n14447), .Z(n14444) );
  XOR2_X1 U14452 ( .A(n14448), .B(n14449), .Z(n14446) );
  NAND2_X1 U14453 ( .A1(n14450), .A2(n14451), .ZN(n14445) );
  NAND2_X1 U14454 ( .A1(n14452), .A2(n14453), .ZN(n14451) );
  NAND2_X1 U14455 ( .A1(n14454), .A2(n14455), .ZN(n14453) );
  INV_X1 U14456 ( .A(n14456), .ZN(n14450) );
  NOR2_X1 U14457 ( .A1(n14455), .A2(n14454), .ZN(n14456) );
  NAND2_X1 U14458 ( .A1(n14457), .A2(n14458), .ZN(n8291) );
  NAND2_X1 U14459 ( .A1(n13950), .A2(n14459), .ZN(n14458) );
  INV_X1 U14460 ( .A(n14460), .ZN(n14459) );
  NOR2_X1 U14461 ( .A1(n13948), .A2(n13949), .ZN(n14460) );
  NOR2_X1 U14462 ( .A1(n8457), .A2(n14123), .ZN(n13950) );
  NAND2_X1 U14463 ( .A1(n13948), .A2(n13949), .ZN(n14457) );
  NAND2_X1 U14464 ( .A1(n14461), .A2(n14462), .ZN(n13949) );
  NAND2_X1 U14465 ( .A1(n14204), .A2(n14463), .ZN(n14462) );
  INV_X1 U14466 ( .A(n14464), .ZN(n14463) );
  NOR2_X1 U14467 ( .A1(n14203), .A2(n14202), .ZN(n14464) );
  NOR2_X1 U14468 ( .A1(n8569), .A2(n14123), .ZN(n14204) );
  NAND2_X1 U14469 ( .A1(n14202), .A2(n14203), .ZN(n14461) );
  NAND2_X1 U14470 ( .A1(n14465), .A2(n14466), .ZN(n14203) );
  NAND2_X1 U14471 ( .A1(n14441), .A2(n14467), .ZN(n14466) );
  INV_X1 U14472 ( .A(n14468), .ZN(n14467) );
  NOR2_X1 U14473 ( .A1(n14439), .A2(n14440), .ZN(n14468) );
  NOR2_X1 U14474 ( .A1(n8448), .A2(n14123), .ZN(n14441) );
  NAND2_X1 U14475 ( .A1(n14439), .A2(n14440), .ZN(n14465) );
  NAND2_X1 U14476 ( .A1(n14469), .A2(n14470), .ZN(n14440) );
  NAND2_X1 U14477 ( .A1(n14437), .A2(n14471), .ZN(n14470) );
  NAND2_X1 U14478 ( .A1(n14435), .A2(n14436), .ZN(n14471) );
  NOR2_X1 U14479 ( .A1(n8900), .A2(n14123), .ZN(n14437) );
  INV_X1 U14480 ( .A(n14472), .ZN(n14469) );
  NOR2_X1 U14481 ( .A1(n14435), .A2(n14436), .ZN(n14472) );
  NOR2_X1 U14482 ( .A1(n14473), .A2(n14474), .ZN(n14436) );
  NOR2_X1 U14483 ( .A1(n14432), .A2(n14475), .ZN(n14474) );
  NOR2_X1 U14484 ( .A1(n14431), .A2(n14433), .ZN(n14475) );
  NAND2_X1 U14485 ( .A1(a_4_), .A2(b_8_), .ZN(n14432) );
  INV_X1 U14486 ( .A(n14476), .ZN(n14473) );
  NAND2_X1 U14487 ( .A1(n14431), .A2(n14433), .ZN(n14476) );
  NAND2_X1 U14488 ( .A1(n14477), .A2(n14478), .ZN(n14433) );
  NAND2_X1 U14489 ( .A1(n14429), .A2(n14479), .ZN(n14478) );
  NAND2_X1 U14490 ( .A1(n14427), .A2(n14428), .ZN(n14479) );
  NOR2_X1 U14491 ( .A1(n8938), .A2(n14123), .ZN(n14429) );
  INV_X1 U14492 ( .A(n14480), .ZN(n14477) );
  NOR2_X1 U14493 ( .A1(n14427), .A2(n14428), .ZN(n14480) );
  NOR2_X1 U14494 ( .A1(n14481), .A2(n14482), .ZN(n14428) );
  NOR2_X1 U14495 ( .A1(n14425), .A2(n14483), .ZN(n14482) );
  NOR2_X1 U14496 ( .A1(n14422), .A2(n14424), .ZN(n14483) );
  NAND2_X1 U14497 ( .A1(a_6_), .A2(b_8_), .ZN(n14425) );
  INV_X1 U14498 ( .A(n14484), .ZN(n14481) );
  NAND2_X1 U14499 ( .A1(n14422), .A2(n14424), .ZN(n14484) );
  NAND2_X1 U14500 ( .A1(n14485), .A2(n14486), .ZN(n14424) );
  NAND2_X1 U14501 ( .A1(n14421), .A2(n14487), .ZN(n14486) );
  NAND2_X1 U14502 ( .A1(n14418), .A2(n14420), .ZN(n14487) );
  NOR2_X1 U14503 ( .A1(n8425), .A2(n14123), .ZN(n14421) );
  NAND2_X1 U14504 ( .A1(n14488), .A2(n14489), .ZN(n14485) );
  INV_X1 U14505 ( .A(n14420), .ZN(n14489) );
  NAND2_X1 U14506 ( .A1(n14490), .A2(n14491), .ZN(n14420) );
  NAND2_X1 U14507 ( .A1(n14492), .A2(n14417), .ZN(n14491) );
  NAND2_X1 U14508 ( .A1(n14415), .A2(n14416), .ZN(n14492) );
  INV_X1 U14509 ( .A(n14493), .ZN(n14490) );
  NOR2_X1 U14510 ( .A1(n14415), .A2(n14416), .ZN(n14493) );
  NAND2_X1 U14511 ( .A1(n14494), .A2(n14495), .ZN(n14416) );
  NAND2_X1 U14512 ( .A1(n14241), .A2(n14496), .ZN(n14495) );
  NAND2_X1 U14513 ( .A1(n14240), .A2(n14238), .ZN(n14496) );
  NOR2_X1 U14514 ( .A1(n8971), .A2(n14123), .ZN(n14241) );
  INV_X1 U14515 ( .A(n14497), .ZN(n14494) );
  NOR2_X1 U14516 ( .A1(n14238), .A2(n14240), .ZN(n14497) );
  NOR2_X1 U14517 ( .A1(n14498), .A2(n14499), .ZN(n14240) );
  INV_X1 U14518 ( .A(n14500), .ZN(n14499) );
  NAND2_X1 U14519 ( .A1(n14248), .A2(n14501), .ZN(n14500) );
  NAND2_X1 U14520 ( .A1(n14247), .A2(n14245), .ZN(n14501) );
  NOR2_X1 U14521 ( .A1(n8402), .A2(n14123), .ZN(n14248) );
  NOR2_X1 U14522 ( .A1(n14245), .A2(n14247), .ZN(n14498) );
  NOR2_X1 U14523 ( .A1(n14502), .A2(n14503), .ZN(n14247) );
  INV_X1 U14524 ( .A(n14504), .ZN(n14503) );
  NAND2_X1 U14525 ( .A1(n14413), .A2(n14505), .ZN(n14504) );
  NAND2_X1 U14526 ( .A1(n14412), .A2(n14411), .ZN(n14505) );
  NOR2_X1 U14527 ( .A1(n8867), .A2(n14123), .ZN(n14413) );
  NOR2_X1 U14528 ( .A1(n14411), .A2(n14412), .ZN(n14502) );
  NOR2_X1 U14529 ( .A1(n14506), .A2(n14507), .ZN(n14412) );
  INV_X1 U14530 ( .A(n14508), .ZN(n14507) );
  NAND2_X1 U14531 ( .A1(n14409), .A2(n14509), .ZN(n14508) );
  NAND2_X1 U14532 ( .A1(n14406), .A2(n14408), .ZN(n14509) );
  NOR2_X1 U14533 ( .A1(n8393), .A2(n14123), .ZN(n14409) );
  NOR2_X1 U14534 ( .A1(n14408), .A2(n14406), .ZN(n14506) );
  XOR2_X1 U14535 ( .A(n14510), .B(n14511), .Z(n14406) );
  XNOR2_X1 U14536 ( .A(n14512), .B(n14513), .ZN(n14510) );
  NOR2_X1 U14537 ( .A1(n14345), .A2(n8996), .ZN(n14513) );
  NAND2_X1 U14538 ( .A1(n14514), .A2(n14515), .ZN(n14408) );
  NAND2_X1 U14539 ( .A1(n14402), .A2(n14516), .ZN(n14515) );
  NAND2_X1 U14540 ( .A1(n14405), .A2(n14404), .ZN(n14516) );
  XOR2_X1 U14541 ( .A(n14517), .B(n14518), .Z(n14402) );
  XOR2_X1 U14542 ( .A(n14519), .B(n14520), .Z(n14518) );
  NAND2_X1 U14543 ( .A1(a_14_), .A2(b_7_), .ZN(n14520) );
  INV_X1 U14544 ( .A(n14521), .ZN(n14514) );
  NOR2_X1 U14545 ( .A1(n14404), .A2(n14405), .ZN(n14521) );
  NOR2_X1 U14546 ( .A1(n8996), .A2(n14123), .ZN(n14405) );
  NAND2_X1 U14547 ( .A1(n14400), .A2(n14522), .ZN(n14404) );
  NAND2_X1 U14548 ( .A1(n14399), .A2(n14401), .ZN(n14522) );
  NAND2_X1 U14549 ( .A1(n14523), .A2(n14524), .ZN(n14401) );
  NAND2_X1 U14550 ( .A1(a_14_), .A2(b_8_), .ZN(n14524) );
  INV_X1 U14551 ( .A(n14525), .ZN(n14523) );
  XNOR2_X1 U14552 ( .A(n14526), .B(n14527), .ZN(n14399) );
  XOR2_X1 U14553 ( .A(n14528), .B(n14529), .Z(n14527) );
  NAND2_X1 U14554 ( .A1(a_15_), .A2(b_7_), .ZN(n14529) );
  NAND2_X1 U14555 ( .A1(a_14_), .A2(n14525), .ZN(n14400) );
  NAND2_X1 U14556 ( .A1(n14396), .A2(n14530), .ZN(n14525) );
  NAND2_X1 U14557 ( .A1(n14395), .A2(n14397), .ZN(n14530) );
  NAND2_X1 U14558 ( .A1(n14531), .A2(n14532), .ZN(n14397) );
  NAND2_X1 U14559 ( .A1(a_15_), .A2(b_8_), .ZN(n14532) );
  INV_X1 U14560 ( .A(n14533), .ZN(n14531) );
  XOR2_X1 U14561 ( .A(n14534), .B(n14535), .Z(n14395) );
  XOR2_X1 U14562 ( .A(n14536), .B(n14537), .Z(n14534) );
  NOR2_X1 U14563 ( .A1(n14345), .A2(n8376), .ZN(n14537) );
  NAND2_X1 U14564 ( .A1(a_15_), .A2(n14533), .ZN(n14396) );
  NAND2_X1 U14565 ( .A1(n14392), .A2(n14538), .ZN(n14533) );
  NAND2_X1 U14566 ( .A1(n14391), .A2(n14393), .ZN(n14538) );
  NAND2_X1 U14567 ( .A1(n14539), .A2(n14540), .ZN(n14393) );
  NAND2_X1 U14568 ( .A1(a_16_), .A2(b_8_), .ZN(n14540) );
  INV_X1 U14569 ( .A(n14541), .ZN(n14539) );
  XOR2_X1 U14570 ( .A(n14542), .B(n14543), .Z(n14391) );
  XNOR2_X1 U14571 ( .A(n14544), .B(n14545), .ZN(n14543) );
  NAND2_X1 U14572 ( .A1(a_17_), .A2(b_7_), .ZN(n14545) );
  NAND2_X1 U14573 ( .A1(a_16_), .A2(n14541), .ZN(n14392) );
  NAND2_X1 U14574 ( .A1(n14388), .A2(n14546), .ZN(n14541) );
  NAND2_X1 U14575 ( .A1(n14387), .A2(n14389), .ZN(n14546) );
  NAND2_X1 U14576 ( .A1(n14547), .A2(n14548), .ZN(n14389) );
  NAND2_X1 U14577 ( .A1(a_17_), .A2(b_8_), .ZN(n14548) );
  INV_X1 U14578 ( .A(n14549), .ZN(n14547) );
  XOR2_X1 U14579 ( .A(n14550), .B(n14551), .Z(n14387) );
  XOR2_X1 U14580 ( .A(n14552), .B(n14553), .Z(n14550) );
  NOR2_X1 U14581 ( .A1(n14345), .A2(n9291), .ZN(n14553) );
  NAND2_X1 U14582 ( .A1(a_17_), .A2(n14549), .ZN(n14388) );
  NAND2_X1 U14583 ( .A1(n14384), .A2(n14554), .ZN(n14549) );
  NAND2_X1 U14584 ( .A1(n14383), .A2(n14385), .ZN(n14554) );
  NAND2_X1 U14585 ( .A1(n14555), .A2(n14556), .ZN(n14385) );
  NAND2_X1 U14586 ( .A1(a_18_), .A2(b_8_), .ZN(n14556) );
  XNOR2_X1 U14587 ( .A(n14557), .B(n14558), .ZN(n14383) );
  XOR2_X1 U14588 ( .A(n14559), .B(n14560), .Z(n14558) );
  NAND2_X1 U14589 ( .A1(b_7_), .A2(a_19_), .ZN(n14560) );
  INV_X1 U14590 ( .A(n14561), .ZN(n14384) );
  NOR2_X1 U14591 ( .A1(n9291), .A2(n14555), .ZN(n14561) );
  NOR2_X1 U14592 ( .A1(n14562), .A2(n14563), .ZN(n14555) );
  NOR3_X1 U14593 ( .A1(n8742), .A2(n14564), .A3(n14123), .ZN(n14563) );
  NOR2_X1 U14594 ( .A1(n14378), .A2(n14565), .ZN(n14564) );
  INV_X1 U14595 ( .A(n14380), .ZN(n14565) );
  NOR2_X1 U14596 ( .A1(n14566), .A2(n14380), .ZN(n14562) );
  NOR2_X1 U14597 ( .A1(n14567), .A2(n14568), .ZN(n14380) );
  INV_X1 U14598 ( .A(n14569), .ZN(n14568) );
  NAND2_X1 U14599 ( .A1(n14377), .A2(n14570), .ZN(n14569) );
  NAND2_X1 U14600 ( .A1(n14376), .A2(n14375), .ZN(n14570) );
  NOR2_X1 U14601 ( .A1(n14123), .A2(n9047), .ZN(n14377) );
  NOR2_X1 U14602 ( .A1(n14375), .A2(n14376), .ZN(n14567) );
  NOR2_X1 U14603 ( .A1(n14571), .A2(n14572), .ZN(n14376) );
  NOR2_X1 U14604 ( .A1(n14373), .A2(n14573), .ZN(n14572) );
  NOR2_X1 U14605 ( .A1(n14370), .A2(n14372), .ZN(n14573) );
  NAND2_X1 U14606 ( .A1(b_8_), .A2(a_21_), .ZN(n14373) );
  INV_X1 U14607 ( .A(n14574), .ZN(n14571) );
  NAND2_X1 U14608 ( .A1(n14370), .A2(n14372), .ZN(n14574) );
  NAND2_X1 U14609 ( .A1(n14575), .A2(n14576), .ZN(n14372) );
  NAND2_X1 U14610 ( .A1(n14369), .A2(n14577), .ZN(n14576) );
  INV_X1 U14611 ( .A(n14578), .ZN(n14577) );
  NOR2_X1 U14612 ( .A1(n14368), .A2(n14366), .ZN(n14578) );
  NOR2_X1 U14613 ( .A1(n14123), .A2(n12296), .ZN(n14369) );
  NAND2_X1 U14614 ( .A1(n14366), .A2(n14368), .ZN(n14575) );
  NAND2_X1 U14615 ( .A1(n14579), .A2(n14580), .ZN(n14368) );
  NAND2_X1 U14616 ( .A1(n14365), .A2(n14581), .ZN(n14580) );
  INV_X1 U14617 ( .A(n14582), .ZN(n14581) );
  NOR2_X1 U14618 ( .A1(n14364), .A2(n14363), .ZN(n14582) );
  NOR2_X1 U14619 ( .A1(n14123), .A2(n12301), .ZN(n14365) );
  NAND2_X1 U14620 ( .A1(n14363), .A2(n14364), .ZN(n14579) );
  NAND2_X1 U14621 ( .A1(n14583), .A2(n14584), .ZN(n14364) );
  NAND2_X1 U14622 ( .A1(n14361), .A2(n14585), .ZN(n14584) );
  INV_X1 U14623 ( .A(n14586), .ZN(n14585) );
  NOR2_X1 U14624 ( .A1(n14359), .A2(n14360), .ZN(n14586) );
  NOR2_X1 U14625 ( .A1(n14123), .A2(n8779), .ZN(n14361) );
  NAND2_X1 U14626 ( .A1(n14359), .A2(n14360), .ZN(n14583) );
  NAND2_X1 U14627 ( .A1(n14587), .A2(n14588), .ZN(n14360) );
  NAND2_X1 U14628 ( .A1(n14357), .A2(n14589), .ZN(n14588) );
  NAND2_X1 U14629 ( .A1(n14354), .A2(n14356), .ZN(n14589) );
  NOR2_X1 U14630 ( .A1(n14123), .A2(n8788), .ZN(n14357) );
  INV_X1 U14631 ( .A(n14590), .ZN(n14587) );
  NOR2_X1 U14632 ( .A1(n14356), .A2(n14354), .ZN(n14590) );
  XNOR2_X1 U14633 ( .A(n14591), .B(n14592), .ZN(n14354) );
  XNOR2_X1 U14634 ( .A(n14593), .B(n14594), .ZN(n14592) );
  NAND2_X1 U14635 ( .A1(n14595), .A2(n14596), .ZN(n14356) );
  NAND2_X1 U14636 ( .A1(n14315), .A2(n14597), .ZN(n14596) );
  NAND2_X1 U14637 ( .A1(n14318), .A2(n14317), .ZN(n14597) );
  XNOR2_X1 U14638 ( .A(n14598), .B(n14599), .ZN(n14315) );
  XOR2_X1 U14639 ( .A(n14600), .B(n14601), .Z(n14598) );
  INV_X1 U14640 ( .A(n14602), .ZN(n14595) );
  NOR2_X1 U14641 ( .A1(n14317), .A2(n14318), .ZN(n14602) );
  NOR2_X1 U14642 ( .A1(n9344), .A2(n14123), .ZN(n14318) );
  NAND2_X1 U14643 ( .A1(n14603), .A2(n14604), .ZN(n14317) );
  NAND2_X1 U14644 ( .A1(n14325), .A2(n14605), .ZN(n14604) );
  INV_X1 U14645 ( .A(n14606), .ZN(n14605) );
  NOR2_X1 U14646 ( .A1(n14323), .A2(n14324), .ZN(n14606) );
  NOR2_X1 U14647 ( .A1(n14123), .A2(n8797), .ZN(n14325) );
  NAND2_X1 U14648 ( .A1(n14323), .A2(n14324), .ZN(n14603) );
  NAND2_X1 U14649 ( .A1(n14607), .A2(n14608), .ZN(n14324) );
  NAND2_X1 U14650 ( .A1(n14352), .A2(n14609), .ZN(n14608) );
  INV_X1 U14651 ( .A(n14610), .ZN(n14609) );
  NOR2_X1 U14652 ( .A1(n14353), .A2(n14351), .ZN(n14610) );
  NOR2_X1 U14653 ( .A1(n14123), .A2(n8314), .ZN(n14352) );
  NAND2_X1 U14654 ( .A1(n14351), .A2(n14353), .ZN(n14607) );
  NAND2_X1 U14655 ( .A1(n14611), .A2(n14612), .ZN(n14353) );
  NAND2_X1 U14656 ( .A1(n14347), .A2(n14613), .ZN(n14612) );
  INV_X1 U14657 ( .A(n14614), .ZN(n14613) );
  NOR2_X1 U14658 ( .A1(n14348), .A2(n14349), .ZN(n14614) );
  NOR2_X1 U14659 ( .A1(n14123), .A2(n9098), .ZN(n14347) );
  NAND2_X1 U14660 ( .A1(n14349), .A2(n14348), .ZN(n14611) );
  NAND2_X1 U14661 ( .A1(n14615), .A2(n14616), .ZN(n14348) );
  NAND2_X1 U14662 ( .A1(b_6_), .A2(n14617), .ZN(n14616) );
  NAND2_X1 U14663 ( .A1(n8299), .A2(n14618), .ZN(n14617) );
  NAND2_X1 U14664 ( .A1(a_31_), .A2(n14345), .ZN(n14618) );
  NAND2_X1 U14665 ( .A1(b_7_), .A2(n14619), .ZN(n14615) );
  NAND2_X1 U14666 ( .A1(n8303), .A2(n14620), .ZN(n14619) );
  NAND2_X1 U14667 ( .A1(a_30_), .A2(n14621), .ZN(n14620) );
  NOR3_X1 U14668 ( .A1(n14123), .A2(n9631), .A3(n14345), .ZN(n14349) );
  XOR2_X1 U14669 ( .A(n14622), .B(n14623), .Z(n14351) );
  XOR2_X1 U14670 ( .A(n14624), .B(n14625), .Z(n14622) );
  XOR2_X1 U14671 ( .A(n14626), .B(n14627), .Z(n14323) );
  XOR2_X1 U14672 ( .A(n14628), .B(n14629), .Z(n14626) );
  XNOR2_X1 U14673 ( .A(n14630), .B(n14631), .ZN(n14359) );
  XNOR2_X1 U14674 ( .A(n14632), .B(n14633), .ZN(n14631) );
  XOR2_X1 U14675 ( .A(n14634), .B(n14635), .Z(n14363) );
  XOR2_X1 U14676 ( .A(n14636), .B(n14637), .Z(n14634) );
  XOR2_X1 U14677 ( .A(n14638), .B(n14639), .Z(n14366) );
  XOR2_X1 U14678 ( .A(n14640), .B(n14641), .Z(n14638) );
  XNOR2_X1 U14679 ( .A(n14642), .B(n14643), .ZN(n14370) );
  NAND2_X1 U14680 ( .A1(n14644), .A2(n14645), .ZN(n14642) );
  XOR2_X1 U14681 ( .A(n14646), .B(n14647), .Z(n14375) );
  XOR2_X1 U14682 ( .A(n14648), .B(n14649), .Z(n14646) );
  INV_X1 U14683 ( .A(n14378), .ZN(n14566) );
  XOR2_X1 U14684 ( .A(n14650), .B(n14651), .Z(n14378) );
  XNOR2_X1 U14685 ( .A(n14652), .B(n14653), .ZN(n14651) );
  NAND2_X1 U14686 ( .A1(b_7_), .A2(a_20_), .ZN(n14653) );
  XOR2_X1 U14687 ( .A(n14654), .B(n14655), .Z(n14411) );
  XNOR2_X1 U14688 ( .A(n14656), .B(n14657), .ZN(n14654) );
  NOR2_X1 U14689 ( .A1(n14345), .A2(n8393), .ZN(n14657) );
  XOR2_X1 U14690 ( .A(n14658), .B(n14659), .Z(n14245) );
  XNOR2_X1 U14691 ( .A(n14660), .B(n14661), .ZN(n14658) );
  NOR2_X1 U14692 ( .A1(n14345), .A2(n8867), .ZN(n14661) );
  XOR2_X1 U14693 ( .A(n14662), .B(n14663), .Z(n14238) );
  XNOR2_X1 U14694 ( .A(n14664), .B(n14665), .ZN(n14662) );
  NOR2_X1 U14695 ( .A1(n14345), .A2(n8402), .ZN(n14665) );
  XNOR2_X1 U14696 ( .A(n14666), .B(n14667), .ZN(n14415) );
  XNOR2_X1 U14697 ( .A(n14668), .B(n14669), .ZN(n14666) );
  NOR2_X1 U14698 ( .A1(n14345), .A2(n8971), .ZN(n14669) );
  INV_X1 U14699 ( .A(n14418), .ZN(n14488) );
  XNOR2_X1 U14700 ( .A(n14670), .B(n14671), .ZN(n14418) );
  XNOR2_X1 U14701 ( .A(n14672), .B(n14673), .ZN(n14671) );
  NAND2_X1 U14702 ( .A1(a_8_), .A2(b_7_), .ZN(n14673) );
  XNOR2_X1 U14703 ( .A(n14674), .B(n14675), .ZN(n14422) );
  XOR2_X1 U14704 ( .A(n14676), .B(n14677), .Z(n14674) );
  XOR2_X1 U14705 ( .A(n14678), .B(n14679), .Z(n14427) );
  XNOR2_X1 U14706 ( .A(n14680), .B(n14681), .ZN(n14679) );
  XNOR2_X1 U14707 ( .A(n14682), .B(n14683), .ZN(n14431) );
  XNOR2_X1 U14708 ( .A(n14684), .B(n14685), .ZN(n14682) );
  XNOR2_X1 U14709 ( .A(n14686), .B(n14687), .ZN(n14435) );
  XOR2_X1 U14710 ( .A(n14688), .B(n14689), .Z(n14687) );
  XNOR2_X1 U14711 ( .A(n14690), .B(n14691), .ZN(n14439) );
  XNOR2_X1 U14712 ( .A(n14692), .B(n14693), .ZN(n14690) );
  XNOR2_X1 U14713 ( .A(n14694), .B(n14695), .ZN(n14202) );
  XNOR2_X1 U14714 ( .A(n14696), .B(n14697), .ZN(n14694) );
  XOR2_X1 U14715 ( .A(n14698), .B(n14699), .Z(n13948) );
  XOR2_X1 U14716 ( .A(n14700), .B(n14701), .Z(n14699) );
  XNOR2_X1 U14717 ( .A(n14702), .B(n14455), .ZN(n8292) );
  XOR2_X1 U14718 ( .A(n14703), .B(n14704), .Z(n14455) );
  XNOR2_X1 U14719 ( .A(n14705), .B(n14706), .ZN(n14704) );
  XNOR2_X1 U14720 ( .A(n14454), .B(n14452), .ZN(n14702) );
  NOR2_X1 U14721 ( .A1(n8457), .A2(n14345), .ZN(n14452) );
  NOR2_X1 U14722 ( .A1(n14707), .A2(n14708), .ZN(n14454) );
  INV_X1 U14723 ( .A(n14709), .ZN(n14708) );
  NAND2_X1 U14724 ( .A1(n14701), .A2(n14710), .ZN(n14709) );
  NAND2_X1 U14725 ( .A1(n14700), .A2(n14698), .ZN(n14710) );
  NOR2_X1 U14726 ( .A1(n8569), .A2(n14345), .ZN(n14701) );
  NOR2_X1 U14727 ( .A1(n14698), .A2(n14700), .ZN(n14707) );
  NOR2_X1 U14728 ( .A1(n14711), .A2(n14712), .ZN(n14700) );
  INV_X1 U14729 ( .A(n14713), .ZN(n14712) );
  NAND2_X1 U14730 ( .A1(n14697), .A2(n14714), .ZN(n14713) );
  NAND2_X1 U14731 ( .A1(n14695), .A2(n14696), .ZN(n14714) );
  NOR2_X1 U14732 ( .A1(n8448), .A2(n14345), .ZN(n14697) );
  NOR2_X1 U14733 ( .A1(n14695), .A2(n14696), .ZN(n14711) );
  NOR2_X1 U14734 ( .A1(n14715), .A2(n14716), .ZN(n14696) );
  INV_X1 U14735 ( .A(n14717), .ZN(n14716) );
  NAND2_X1 U14736 ( .A1(n14693), .A2(n14718), .ZN(n14717) );
  NAND2_X1 U14737 ( .A1(n14692), .A2(n14691), .ZN(n14718) );
  NOR2_X1 U14738 ( .A1(n8900), .A2(n14345), .ZN(n14693) );
  NOR2_X1 U14739 ( .A1(n14691), .A2(n14692), .ZN(n14715) );
  NOR2_X1 U14740 ( .A1(n14719), .A2(n14720), .ZN(n14692) );
  INV_X1 U14741 ( .A(n14721), .ZN(n14720) );
  NAND2_X1 U14742 ( .A1(n14689), .A2(n14722), .ZN(n14721) );
  NAND2_X1 U14743 ( .A1(n14688), .A2(n14686), .ZN(n14722) );
  NOR2_X1 U14744 ( .A1(n8439), .A2(n14345), .ZN(n14689) );
  NOR2_X1 U14745 ( .A1(n14686), .A2(n14688), .ZN(n14719) );
  NOR2_X1 U14746 ( .A1(n14723), .A2(n14724), .ZN(n14688) );
  INV_X1 U14747 ( .A(n14725), .ZN(n14724) );
  NAND2_X1 U14748 ( .A1(n14685), .A2(n14726), .ZN(n14725) );
  NAND2_X1 U14749 ( .A1(n14684), .A2(n14683), .ZN(n14726) );
  NOR2_X1 U14750 ( .A1(n8938), .A2(n14345), .ZN(n14685) );
  NOR2_X1 U14751 ( .A1(n14683), .A2(n14684), .ZN(n14723) );
  NOR2_X1 U14752 ( .A1(n14727), .A2(n14728), .ZN(n14684) );
  INV_X1 U14753 ( .A(n14729), .ZN(n14728) );
  NAND2_X1 U14754 ( .A1(n14681), .A2(n14730), .ZN(n14729) );
  NAND2_X1 U14755 ( .A1(n14678), .A2(n14680), .ZN(n14730) );
  NOR2_X1 U14756 ( .A1(n8430), .A2(n14345), .ZN(n14681) );
  NOR2_X1 U14757 ( .A1(n14680), .A2(n14678), .ZN(n14727) );
  XNOR2_X1 U14758 ( .A(n14731), .B(n14732), .ZN(n14678) );
  XOR2_X1 U14759 ( .A(n14733), .B(n14734), .Z(n14732) );
  NAND2_X1 U14760 ( .A1(n14735), .A2(n14736), .ZN(n14680) );
  NAND2_X1 U14761 ( .A1(n14675), .A2(n14737), .ZN(n14736) );
  NAND2_X1 U14762 ( .A1(n14677), .A2(n14676), .ZN(n14737) );
  INV_X1 U14763 ( .A(n14738), .ZN(n14676) );
  XOR2_X1 U14764 ( .A(n14739), .B(n14740), .Z(n14675) );
  XNOR2_X1 U14765 ( .A(n14741), .B(n14742), .ZN(n14739) );
  NAND2_X1 U14766 ( .A1(n14738), .A2(n14743), .ZN(n14735) );
  NOR2_X1 U14767 ( .A1(n14744), .A2(n14745), .ZN(n14738) );
  INV_X1 U14768 ( .A(n14746), .ZN(n14745) );
  NAND3_X1 U14769 ( .A1(b_7_), .A2(n14747), .A3(a_8_), .ZN(n14746) );
  NAND2_X1 U14770 ( .A1(n14670), .A2(n14672), .ZN(n14747) );
  NOR2_X1 U14771 ( .A1(n14670), .A2(n14672), .ZN(n14744) );
  NOR2_X1 U14772 ( .A1(n14748), .A2(n14749), .ZN(n14672) );
  INV_X1 U14773 ( .A(n14750), .ZN(n14749) );
  NAND3_X1 U14774 ( .A1(b_7_), .A2(n14751), .A3(a_9_), .ZN(n14750) );
  NAND2_X1 U14775 ( .A1(n14668), .A2(n14667), .ZN(n14751) );
  NOR2_X1 U14776 ( .A1(n14667), .A2(n14668), .ZN(n14748) );
  NOR2_X1 U14777 ( .A1(n14752), .A2(n14753), .ZN(n14668) );
  NOR3_X1 U14778 ( .A1(n14345), .A2(n14754), .A3(n8402), .ZN(n14753) );
  INV_X1 U14779 ( .A(n14755), .ZN(n14754) );
  NAND2_X1 U14780 ( .A1(n14663), .A2(n14664), .ZN(n14755) );
  NOR2_X1 U14781 ( .A1(n14663), .A2(n14664), .ZN(n14752) );
  NOR2_X1 U14782 ( .A1(n14756), .A2(n14757), .ZN(n14664) );
  INV_X1 U14783 ( .A(n14758), .ZN(n14757) );
  NAND3_X1 U14784 ( .A1(b_7_), .A2(n14759), .A3(a_11_), .ZN(n14758) );
  NAND2_X1 U14785 ( .A1(n14659), .A2(n14660), .ZN(n14759) );
  NOR2_X1 U14786 ( .A1(n14659), .A2(n14660), .ZN(n14756) );
  NOR2_X1 U14787 ( .A1(n14760), .A2(n14761), .ZN(n14660) );
  INV_X1 U14788 ( .A(n14762), .ZN(n14761) );
  NAND3_X1 U14789 ( .A1(b_7_), .A2(n14763), .A3(a_12_), .ZN(n14762) );
  NAND2_X1 U14790 ( .A1(n14655), .A2(n14656), .ZN(n14763) );
  NOR2_X1 U14791 ( .A1(n14655), .A2(n14656), .ZN(n14760) );
  NOR2_X1 U14792 ( .A1(n14764), .A2(n14765), .ZN(n14656) );
  INV_X1 U14793 ( .A(n14766), .ZN(n14765) );
  NAND3_X1 U14794 ( .A1(b_7_), .A2(n14767), .A3(a_13_), .ZN(n14766) );
  NAND2_X1 U14795 ( .A1(n14512), .A2(n14511), .ZN(n14767) );
  NOR2_X1 U14796 ( .A1(n14511), .A2(n14512), .ZN(n14764) );
  NOR2_X1 U14797 ( .A1(n14768), .A2(n14769), .ZN(n14512) );
  NOR3_X1 U14798 ( .A1(n14345), .A2(n14770), .A3(n9262), .ZN(n14769) );
  NOR2_X1 U14799 ( .A1(n14517), .A2(n14519), .ZN(n14770) );
  INV_X1 U14800 ( .A(n14771), .ZN(n14768) );
  NAND2_X1 U14801 ( .A1(n14517), .A2(n14519), .ZN(n14771) );
  NAND2_X1 U14802 ( .A1(n14772), .A2(n14773), .ZN(n14519) );
  NAND3_X1 U14803 ( .A1(b_7_), .A2(n14774), .A3(a_15_), .ZN(n14773) );
  INV_X1 U14804 ( .A(n14775), .ZN(n14774) );
  NOR2_X1 U14805 ( .A1(n14528), .A2(n14526), .ZN(n14775) );
  NAND2_X1 U14806 ( .A1(n14526), .A2(n14528), .ZN(n14772) );
  NAND2_X1 U14807 ( .A1(n14776), .A2(n14777), .ZN(n14528) );
  NAND3_X1 U14808 ( .A1(b_7_), .A2(n14778), .A3(a_16_), .ZN(n14777) );
  INV_X1 U14809 ( .A(n14779), .ZN(n14778) );
  NOR2_X1 U14810 ( .A1(n14535), .A2(n14536), .ZN(n14779) );
  NAND2_X1 U14811 ( .A1(n14535), .A2(n14536), .ZN(n14776) );
  NAND2_X1 U14812 ( .A1(n14780), .A2(n14781), .ZN(n14536) );
  NAND3_X1 U14813 ( .A1(b_7_), .A2(n14782), .A3(a_17_), .ZN(n14781) );
  NAND2_X1 U14814 ( .A1(n14542), .A2(n14544), .ZN(n14782) );
  INV_X1 U14815 ( .A(n14783), .ZN(n14780) );
  NOR2_X1 U14816 ( .A1(n14542), .A2(n14544), .ZN(n14783) );
  NOR2_X1 U14817 ( .A1(n14784), .A2(n14785), .ZN(n14544) );
  NOR3_X1 U14818 ( .A1(n14345), .A2(n14786), .A3(n9291), .ZN(n14785) );
  NOR2_X1 U14819 ( .A1(n14551), .A2(n14552), .ZN(n14786) );
  INV_X1 U14820 ( .A(n14787), .ZN(n14784) );
  NAND2_X1 U14821 ( .A1(n14551), .A2(n14552), .ZN(n14787) );
  NAND2_X1 U14822 ( .A1(n14788), .A2(n14789), .ZN(n14552) );
  INV_X1 U14823 ( .A(n14790), .ZN(n14789) );
  NOR3_X1 U14824 ( .A1(n8742), .A2(n14791), .A3(n14345), .ZN(n14790) );
  NOR2_X1 U14825 ( .A1(n14559), .A2(n14557), .ZN(n14791) );
  NAND2_X1 U14826 ( .A1(n14557), .A2(n14559), .ZN(n14788) );
  NAND2_X1 U14827 ( .A1(n14792), .A2(n14793), .ZN(n14559) );
  NAND3_X1 U14828 ( .A1(a_20_), .A2(n14794), .A3(b_7_), .ZN(n14793) );
  NAND2_X1 U14829 ( .A1(n14795), .A2(n14796), .ZN(n14794) );
  INV_X1 U14830 ( .A(n14652), .ZN(n14796) );
  INV_X1 U14831 ( .A(n14650), .ZN(n14795) );
  NAND2_X1 U14832 ( .A1(n14652), .A2(n14650), .ZN(n14792) );
  XOR2_X1 U14833 ( .A(n14797), .B(n14798), .Z(n14650) );
  XOR2_X1 U14834 ( .A(n14799), .B(n14800), .Z(n14797) );
  NOR2_X1 U14835 ( .A1(n8759), .A2(n14621), .ZN(n14800) );
  NOR2_X1 U14836 ( .A1(n14801), .A2(n14802), .ZN(n14652) );
  INV_X1 U14837 ( .A(n14803), .ZN(n14802) );
  NAND2_X1 U14838 ( .A1(n14647), .A2(n14804), .ZN(n14803) );
  NAND2_X1 U14839 ( .A1(n14649), .A2(n14648), .ZN(n14804) );
  XOR2_X1 U14840 ( .A(n14805), .B(n14806), .Z(n14647) );
  NAND2_X1 U14841 ( .A1(n14807), .A2(n14808), .ZN(n14805) );
  NOR2_X1 U14842 ( .A1(n14648), .A2(n14649), .ZN(n14801) );
  NOR2_X1 U14843 ( .A1(n14345), .A2(n8759), .ZN(n14649) );
  NAND2_X1 U14844 ( .A1(n14644), .A2(n14809), .ZN(n14648) );
  NAND2_X1 U14845 ( .A1(n14643), .A2(n14645), .ZN(n14809) );
  NAND2_X1 U14846 ( .A1(n14810), .A2(n14811), .ZN(n14645) );
  NAND2_X1 U14847 ( .A1(b_7_), .A2(a_22_), .ZN(n14811) );
  INV_X1 U14848 ( .A(n14812), .ZN(n14810) );
  XNOR2_X1 U14849 ( .A(n14813), .B(n14814), .ZN(n14643) );
  XNOR2_X1 U14850 ( .A(n14815), .B(n14816), .ZN(n14813) );
  NOR2_X1 U14851 ( .A1(n12301), .A2(n14621), .ZN(n14816) );
  NAND2_X1 U14852 ( .A1(a_22_), .A2(n14812), .ZN(n14644) );
  NAND2_X1 U14853 ( .A1(n14817), .A2(n14818), .ZN(n14812) );
  NAND2_X1 U14854 ( .A1(n14641), .A2(n14819), .ZN(n14818) );
  INV_X1 U14855 ( .A(n14820), .ZN(n14819) );
  NOR2_X1 U14856 ( .A1(n14639), .A2(n14640), .ZN(n14820) );
  NOR2_X1 U14857 ( .A1(n14345), .A2(n12301), .ZN(n14641) );
  NAND2_X1 U14858 ( .A1(n14639), .A2(n14640), .ZN(n14817) );
  NAND2_X1 U14859 ( .A1(n14821), .A2(n14822), .ZN(n14640) );
  NAND2_X1 U14860 ( .A1(n14637), .A2(n14823), .ZN(n14822) );
  INV_X1 U14861 ( .A(n14824), .ZN(n14823) );
  NOR2_X1 U14862 ( .A1(n14635), .A2(n14636), .ZN(n14824) );
  NOR2_X1 U14863 ( .A1(n14345), .A2(n8779), .ZN(n14637) );
  NAND2_X1 U14864 ( .A1(n14635), .A2(n14636), .ZN(n14821) );
  NAND2_X1 U14865 ( .A1(n14825), .A2(n14826), .ZN(n14636) );
  NAND2_X1 U14866 ( .A1(n14633), .A2(n14827), .ZN(n14826) );
  NAND2_X1 U14867 ( .A1(n14630), .A2(n14632), .ZN(n14827) );
  NOR2_X1 U14868 ( .A1(n14345), .A2(n8788), .ZN(n14633) );
  INV_X1 U14869 ( .A(n14828), .ZN(n14825) );
  NOR2_X1 U14870 ( .A1(n14632), .A2(n14630), .ZN(n14828) );
  XNOR2_X1 U14871 ( .A(n14829), .B(n14830), .ZN(n14630) );
  XNOR2_X1 U14872 ( .A(n14831), .B(n14832), .ZN(n14830) );
  NAND2_X1 U14873 ( .A1(n14833), .A2(n14834), .ZN(n14632) );
  NAND2_X1 U14874 ( .A1(n14591), .A2(n14835), .ZN(n14834) );
  NAND2_X1 U14875 ( .A1(n14594), .A2(n14593), .ZN(n14835) );
  XNOR2_X1 U14876 ( .A(n14836), .B(n14837), .ZN(n14591) );
  XOR2_X1 U14877 ( .A(n14838), .B(n14839), .Z(n14836) );
  INV_X1 U14878 ( .A(n14840), .ZN(n14833) );
  NOR2_X1 U14879 ( .A1(n14593), .A2(n14594), .ZN(n14840) );
  NOR2_X1 U14880 ( .A1(n9344), .A2(n14345), .ZN(n14594) );
  NAND2_X1 U14881 ( .A1(n14841), .A2(n14842), .ZN(n14593) );
  NAND2_X1 U14882 ( .A1(n14601), .A2(n14843), .ZN(n14842) );
  INV_X1 U14883 ( .A(n14844), .ZN(n14843) );
  NOR2_X1 U14884 ( .A1(n14599), .A2(n14600), .ZN(n14844) );
  NOR2_X1 U14885 ( .A1(n14345), .A2(n8797), .ZN(n14601) );
  NAND2_X1 U14886 ( .A1(n14599), .A2(n14600), .ZN(n14841) );
  NAND2_X1 U14887 ( .A1(n14845), .A2(n14846), .ZN(n14600) );
  NAND2_X1 U14888 ( .A1(n14628), .A2(n14847), .ZN(n14846) );
  INV_X1 U14889 ( .A(n14848), .ZN(n14847) );
  NOR2_X1 U14890 ( .A1(n14629), .A2(n14627), .ZN(n14848) );
  NOR2_X1 U14891 ( .A1(n14345), .A2(n8314), .ZN(n14628) );
  NAND2_X1 U14892 ( .A1(n14627), .A2(n14629), .ZN(n14845) );
  NAND2_X1 U14893 ( .A1(n14849), .A2(n14850), .ZN(n14629) );
  NAND2_X1 U14894 ( .A1(n14623), .A2(n14851), .ZN(n14850) );
  INV_X1 U14895 ( .A(n14852), .ZN(n14851) );
  NOR2_X1 U14896 ( .A1(n14624), .A2(n14625), .ZN(n14852) );
  NOR2_X1 U14897 ( .A1(n14345), .A2(n9098), .ZN(n14623) );
  NAND2_X1 U14898 ( .A1(n14625), .A2(n14624), .ZN(n14849) );
  NAND2_X1 U14899 ( .A1(n14853), .A2(n14854), .ZN(n14624) );
  NAND2_X1 U14900 ( .A1(b_5_), .A2(n14855), .ZN(n14854) );
  NAND2_X1 U14901 ( .A1(n8299), .A2(n14856), .ZN(n14855) );
  NAND2_X1 U14902 ( .A1(a_31_), .A2(n14621), .ZN(n14856) );
  NAND2_X1 U14903 ( .A1(b_6_), .A2(n14857), .ZN(n14853) );
  NAND2_X1 U14904 ( .A1(n8303), .A2(n14858), .ZN(n14857) );
  NAND2_X1 U14905 ( .A1(a_30_), .A2(n14859), .ZN(n14858) );
  NOR3_X1 U14906 ( .A1(n14345), .A2(n9631), .A3(n14621), .ZN(n14625) );
  XOR2_X1 U14907 ( .A(n14860), .B(n14861), .Z(n14627) );
  XOR2_X1 U14908 ( .A(n14862), .B(n14863), .Z(n14860) );
  XOR2_X1 U14909 ( .A(n14864), .B(n14865), .Z(n14599) );
  XOR2_X1 U14910 ( .A(n14866), .B(n14867), .Z(n14864) );
  XNOR2_X1 U14911 ( .A(n14868), .B(n14869), .ZN(n14635) );
  XNOR2_X1 U14912 ( .A(n14870), .B(n14871), .ZN(n14869) );
  XNOR2_X1 U14913 ( .A(n14872), .B(n14873), .ZN(n14639) );
  XNOR2_X1 U14914 ( .A(n14874), .B(n14875), .ZN(n14872) );
  NOR2_X1 U14915 ( .A1(n8779), .A2(n14621), .ZN(n14875) );
  XNOR2_X1 U14916 ( .A(n14876), .B(n14877), .ZN(n14557) );
  NAND2_X1 U14917 ( .A1(n14878), .A2(n14879), .ZN(n14876) );
  XNOR2_X1 U14918 ( .A(n14880), .B(n14881), .ZN(n14551) );
  XOR2_X1 U14919 ( .A(n14882), .B(n14883), .Z(n14880) );
  XOR2_X1 U14920 ( .A(n14884), .B(n14885), .Z(n14542) );
  XNOR2_X1 U14921 ( .A(n14886), .B(n14887), .ZN(n14884) );
  XNOR2_X1 U14922 ( .A(n14888), .B(n14889), .ZN(n14535) );
  XNOR2_X1 U14923 ( .A(n14890), .B(n14891), .ZN(n14889) );
  XNOR2_X1 U14924 ( .A(n14892), .B(n14893), .ZN(n14526) );
  XNOR2_X1 U14925 ( .A(n14894), .B(n14895), .ZN(n14893) );
  XOR2_X1 U14926 ( .A(n14896), .B(n14897), .Z(n14517) );
  XOR2_X1 U14927 ( .A(n14898), .B(n14899), .Z(n14896) );
  XOR2_X1 U14928 ( .A(n14900), .B(n14901), .Z(n14511) );
  XNOR2_X1 U14929 ( .A(n14902), .B(n14903), .ZN(n14900) );
  XOR2_X1 U14930 ( .A(n14904), .B(n14905), .Z(n14655) );
  XNOR2_X1 U14931 ( .A(n14906), .B(n14907), .ZN(n14904) );
  XOR2_X1 U14932 ( .A(n14908), .B(n14909), .Z(n14659) );
  XNOR2_X1 U14933 ( .A(n14910), .B(n14911), .ZN(n14908) );
  XNOR2_X1 U14934 ( .A(n14912), .B(n14913), .ZN(n14663) );
  XOR2_X1 U14935 ( .A(n14914), .B(n14915), .Z(n14913) );
  XNOR2_X1 U14936 ( .A(n14916), .B(n14917), .ZN(n14667) );
  XOR2_X1 U14937 ( .A(n14918), .B(n14919), .Z(n14916) );
  XNOR2_X1 U14938 ( .A(n14920), .B(n14921), .ZN(n14670) );
  XOR2_X1 U14939 ( .A(n14922), .B(n14923), .Z(n14920) );
  XNOR2_X1 U14940 ( .A(n14924), .B(n14925), .ZN(n14683) );
  XNOR2_X1 U14941 ( .A(n14926), .B(n14927), .ZN(n14924) );
  XOR2_X1 U14942 ( .A(n14928), .B(n14929), .Z(n14686) );
  XNOR2_X1 U14943 ( .A(n14930), .B(n14931), .ZN(n14929) );
  XOR2_X1 U14944 ( .A(n14932), .B(n14933), .Z(n14691) );
  XNOR2_X1 U14945 ( .A(n14934), .B(n14935), .ZN(n14933) );
  XNOR2_X1 U14946 ( .A(n14936), .B(n14937), .ZN(n14695) );
  XOR2_X1 U14947 ( .A(n14938), .B(n14939), .Z(n14936) );
  XNOR2_X1 U14948 ( .A(n14940), .B(n14941), .ZN(n14698) );
  XOR2_X1 U14949 ( .A(n14942), .B(n14943), .Z(n14940) );
  XNOR2_X1 U14950 ( .A(n8322), .B(n8323), .ZN(n8295) );
  NAND3_X1 U14951 ( .A1(n8323), .A2(n8322), .A3(n8320), .ZN(n8324) );
  NOR2_X1 U14952 ( .A1(n14944), .A2(n8577), .ZN(n8320) );
  NOR2_X1 U14953 ( .A1(n14945), .A2(n14946), .ZN(n8577) );
  INV_X1 U14954 ( .A(n14947), .ZN(n14944) );
  NAND2_X1 U14955 ( .A1(n14946), .A2(n14945), .ZN(n14947) );
  XOR2_X1 U14956 ( .A(n14948), .B(n14949), .Z(n14945) );
  XNOR2_X1 U14957 ( .A(n14950), .B(n14951), .ZN(n14948) );
  NOR2_X1 U14958 ( .A1(n14952), .A2(n14953), .ZN(n14946) );
  INV_X1 U14959 ( .A(n14954), .ZN(n14953) );
  NAND3_X1 U14960 ( .A1(b_5_), .A2(n14955), .A3(a_0_), .ZN(n14954) );
  NAND2_X1 U14961 ( .A1(n14956), .A2(n14957), .ZN(n14955) );
  NOR2_X1 U14962 ( .A1(n14957), .A2(n14956), .ZN(n14952) );
  NAND2_X1 U14963 ( .A1(n14958), .A2(n14959), .ZN(n8322) );
  NAND2_X1 U14964 ( .A1(n14449), .A2(n14960), .ZN(n14959) );
  INV_X1 U14965 ( .A(n14961), .ZN(n14960) );
  NOR2_X1 U14966 ( .A1(n14448), .A2(n14447), .ZN(n14961) );
  NOR2_X1 U14967 ( .A1(n8457), .A2(n14621), .ZN(n14449) );
  NAND2_X1 U14968 ( .A1(n14447), .A2(n14448), .ZN(n14958) );
  NAND2_X1 U14969 ( .A1(n14962), .A2(n14963), .ZN(n14448) );
  NAND2_X1 U14970 ( .A1(n14706), .A2(n14964), .ZN(n14963) );
  INV_X1 U14971 ( .A(n14965), .ZN(n14964) );
  NOR2_X1 U14972 ( .A1(n14703), .A2(n14705), .ZN(n14965) );
  NOR2_X1 U14973 ( .A1(n8569), .A2(n14621), .ZN(n14706) );
  NAND2_X1 U14974 ( .A1(n14703), .A2(n14705), .ZN(n14962) );
  NAND2_X1 U14975 ( .A1(n14966), .A2(n14967), .ZN(n14705) );
  NAND2_X1 U14976 ( .A1(n14943), .A2(n14968), .ZN(n14967) );
  INV_X1 U14977 ( .A(n14969), .ZN(n14968) );
  NOR2_X1 U14978 ( .A1(n14941), .A2(n14942), .ZN(n14969) );
  NOR2_X1 U14979 ( .A1(n8448), .A2(n14621), .ZN(n14943) );
  NAND2_X1 U14980 ( .A1(n14941), .A2(n14942), .ZN(n14966) );
  NAND2_X1 U14981 ( .A1(n14970), .A2(n14971), .ZN(n14942) );
  NAND2_X1 U14982 ( .A1(n14939), .A2(n14972), .ZN(n14971) );
  INV_X1 U14983 ( .A(n14973), .ZN(n14972) );
  NOR2_X1 U14984 ( .A1(n14938), .A2(n14937), .ZN(n14973) );
  NOR2_X1 U14985 ( .A1(n8900), .A2(n14621), .ZN(n14939) );
  NAND2_X1 U14986 ( .A1(n14937), .A2(n14938), .ZN(n14970) );
  NAND2_X1 U14987 ( .A1(n14974), .A2(n14975), .ZN(n14938) );
  NAND2_X1 U14988 ( .A1(n14935), .A2(n14976), .ZN(n14975) );
  INV_X1 U14989 ( .A(n14977), .ZN(n14976) );
  NOR2_X1 U14990 ( .A1(n14932), .A2(n14934), .ZN(n14977) );
  NOR2_X1 U14991 ( .A1(n8439), .A2(n14621), .ZN(n14935) );
  NAND2_X1 U14992 ( .A1(n14932), .A2(n14934), .ZN(n14974) );
  NAND2_X1 U14993 ( .A1(n14978), .A2(n14979), .ZN(n14934) );
  NAND2_X1 U14994 ( .A1(n14931), .A2(n14980), .ZN(n14979) );
  NAND2_X1 U14995 ( .A1(n14928), .A2(n14930), .ZN(n14980) );
  NOR2_X1 U14996 ( .A1(n8938), .A2(n14621), .ZN(n14931) );
  INV_X1 U14997 ( .A(n14981), .ZN(n14978) );
  NOR2_X1 U14998 ( .A1(n14928), .A2(n14930), .ZN(n14981) );
  NAND2_X1 U14999 ( .A1(n14982), .A2(n14983), .ZN(n14930) );
  NAND2_X1 U15000 ( .A1(n14984), .A2(n14927), .ZN(n14983) );
  NAND2_X1 U15001 ( .A1(n14925), .A2(n14926), .ZN(n14984) );
  INV_X1 U15002 ( .A(n14985), .ZN(n14982) );
  NOR2_X1 U15003 ( .A1(n14925), .A2(n14926), .ZN(n14985) );
  NAND2_X1 U15004 ( .A1(n14986), .A2(n14987), .ZN(n14926) );
  NAND2_X1 U15005 ( .A1(n14734), .A2(n14988), .ZN(n14987) );
  NAND2_X1 U15006 ( .A1(n14733), .A2(n14731), .ZN(n14988) );
  NOR2_X1 U15007 ( .A1(n8425), .A2(n14621), .ZN(n14734) );
  INV_X1 U15008 ( .A(n14989), .ZN(n14986) );
  NOR2_X1 U15009 ( .A1(n14731), .A2(n14733), .ZN(n14989) );
  NOR2_X1 U15010 ( .A1(n14990), .A2(n14991), .ZN(n14733) );
  INV_X1 U15011 ( .A(n14992), .ZN(n14991) );
  NAND2_X1 U15012 ( .A1(n14742), .A2(n14993), .ZN(n14992) );
  NAND2_X1 U15013 ( .A1(n14740), .A2(n14741), .ZN(n14993) );
  NOR2_X1 U15014 ( .A1(n8968), .A2(n14621), .ZN(n14742) );
  NOR2_X1 U15015 ( .A1(n14740), .A2(n14741), .ZN(n14990) );
  INV_X1 U15016 ( .A(n14994), .ZN(n14741) );
  NAND2_X1 U15017 ( .A1(n14995), .A2(n14996), .ZN(n14994) );
  NAND2_X1 U15018 ( .A1(n14923), .A2(n14997), .ZN(n14996) );
  INV_X1 U15019 ( .A(n14998), .ZN(n14997) );
  NOR2_X1 U15020 ( .A1(n14922), .A2(n14921), .ZN(n14998) );
  NOR2_X1 U15021 ( .A1(n8971), .A2(n14621), .ZN(n14923) );
  NAND2_X1 U15022 ( .A1(n14921), .A2(n14922), .ZN(n14995) );
  NAND2_X1 U15023 ( .A1(n14999), .A2(n15000), .ZN(n14922) );
  NAND2_X1 U15024 ( .A1(n14919), .A2(n15001), .ZN(n15000) );
  INV_X1 U15025 ( .A(n15002), .ZN(n15001) );
  NOR2_X1 U15026 ( .A1(n14917), .A2(n14918), .ZN(n15002) );
  NOR2_X1 U15027 ( .A1(n8402), .A2(n14621), .ZN(n14919) );
  NAND2_X1 U15028 ( .A1(n14917), .A2(n14918), .ZN(n14999) );
  NAND2_X1 U15029 ( .A1(n15003), .A2(n15004), .ZN(n14918) );
  NAND2_X1 U15030 ( .A1(n14915), .A2(n15005), .ZN(n15004) );
  NAND2_X1 U15031 ( .A1(n14914), .A2(n14912), .ZN(n15005) );
  NOR2_X1 U15032 ( .A1(n8867), .A2(n14621), .ZN(n14915) );
  INV_X1 U15033 ( .A(n15006), .ZN(n15003) );
  NOR2_X1 U15034 ( .A1(n14912), .A2(n14914), .ZN(n15006) );
  NOR2_X1 U15035 ( .A1(n15007), .A2(n15008), .ZN(n14914) );
  INV_X1 U15036 ( .A(n15009), .ZN(n15008) );
  NAND2_X1 U15037 ( .A1(n14911), .A2(n15010), .ZN(n15009) );
  NAND2_X1 U15038 ( .A1(n14910), .A2(n14909), .ZN(n15010) );
  NOR2_X1 U15039 ( .A1(n8393), .A2(n14621), .ZN(n14911) );
  NOR2_X1 U15040 ( .A1(n14909), .A2(n14910), .ZN(n15007) );
  NOR2_X1 U15041 ( .A1(n15011), .A2(n15012), .ZN(n14910) );
  INV_X1 U15042 ( .A(n15013), .ZN(n15012) );
  NAND2_X1 U15043 ( .A1(n14907), .A2(n15014), .ZN(n15013) );
  NAND2_X1 U15044 ( .A1(n14906), .A2(n14905), .ZN(n15014) );
  NOR2_X1 U15045 ( .A1(n8996), .A2(n14621), .ZN(n14907) );
  NOR2_X1 U15046 ( .A1(n14905), .A2(n14906), .ZN(n15011) );
  NOR2_X1 U15047 ( .A1(n15015), .A2(n15016), .ZN(n14906) );
  INV_X1 U15048 ( .A(n15017), .ZN(n15016) );
  NAND2_X1 U15049 ( .A1(n14903), .A2(n15018), .ZN(n15017) );
  NAND2_X1 U15050 ( .A1(n14901), .A2(n14902), .ZN(n15018) );
  NOR2_X1 U15051 ( .A1(n9262), .A2(n14621), .ZN(n14903) );
  NOR2_X1 U15052 ( .A1(n14901), .A2(n14902), .ZN(n15015) );
  INV_X1 U15053 ( .A(n15019), .ZN(n14902) );
  NAND2_X1 U15054 ( .A1(n15020), .A2(n15021), .ZN(n15019) );
  NAND2_X1 U15055 ( .A1(n14899), .A2(n15022), .ZN(n15021) );
  INV_X1 U15056 ( .A(n15023), .ZN(n15022) );
  NOR2_X1 U15057 ( .A1(n14898), .A2(n14897), .ZN(n15023) );
  NOR2_X1 U15058 ( .A1(n8850), .A2(n14621), .ZN(n14899) );
  NAND2_X1 U15059 ( .A1(n14897), .A2(n14898), .ZN(n15020) );
  NAND2_X1 U15060 ( .A1(n15024), .A2(n15025), .ZN(n14898) );
  NAND2_X1 U15061 ( .A1(n14895), .A2(n15026), .ZN(n15025) );
  INV_X1 U15062 ( .A(n15027), .ZN(n15026) );
  NOR2_X1 U15063 ( .A1(n14892), .A2(n14894), .ZN(n15027) );
  NOR2_X1 U15064 ( .A1(n8376), .A2(n14621), .ZN(n14895) );
  NAND2_X1 U15065 ( .A1(n14892), .A2(n14894), .ZN(n15024) );
  NAND2_X1 U15066 ( .A1(n15028), .A2(n15029), .ZN(n14894) );
  NAND2_X1 U15067 ( .A1(n14891), .A2(n15030), .ZN(n15029) );
  INV_X1 U15068 ( .A(n15031), .ZN(n15030) );
  NOR2_X1 U15069 ( .A1(n14890), .A2(n14888), .ZN(n15031) );
  NOR2_X1 U15070 ( .A1(n8371), .A2(n14621), .ZN(n14891) );
  NAND2_X1 U15071 ( .A1(n14888), .A2(n14890), .ZN(n15028) );
  NAND2_X1 U15072 ( .A1(n15032), .A2(n15033), .ZN(n14890) );
  NAND2_X1 U15073 ( .A1(n14887), .A2(n15034), .ZN(n15033) );
  INV_X1 U15074 ( .A(n15035), .ZN(n15034) );
  NOR2_X1 U15075 ( .A1(n14885), .A2(n14886), .ZN(n15035) );
  NOR2_X1 U15076 ( .A1(n9291), .A2(n14621), .ZN(n14887) );
  NAND2_X1 U15077 ( .A1(n14886), .A2(n14885), .ZN(n15032) );
  XNOR2_X1 U15078 ( .A(n15036), .B(n15037), .ZN(n14885) );
  XNOR2_X1 U15079 ( .A(n15038), .B(n15039), .ZN(n15036) );
  NOR2_X1 U15080 ( .A1(n8742), .A2(n14859), .ZN(n15039) );
  NOR2_X1 U15081 ( .A1(n15040), .A2(n15041), .ZN(n14886) );
  INV_X1 U15082 ( .A(n15042), .ZN(n15041) );
  NAND2_X1 U15083 ( .A1(n14881), .A2(n15043), .ZN(n15042) );
  NAND2_X1 U15084 ( .A1(n14883), .A2(n14882), .ZN(n15043) );
  XNOR2_X1 U15085 ( .A(n15044), .B(n15045), .ZN(n14881) );
  XOR2_X1 U15086 ( .A(n15046), .B(n15047), .Z(n15044) );
  NOR2_X1 U15087 ( .A1(n9047), .A2(n14859), .ZN(n15047) );
  NOR2_X1 U15088 ( .A1(n14882), .A2(n14883), .ZN(n15040) );
  NOR2_X1 U15089 ( .A1(n14621), .A2(n8742), .ZN(n14883) );
  NAND2_X1 U15090 ( .A1(n14878), .A2(n15048), .ZN(n14882) );
  NAND2_X1 U15091 ( .A1(n14877), .A2(n14879), .ZN(n15048) );
  NAND2_X1 U15092 ( .A1(n15049), .A2(n15050), .ZN(n14879) );
  NAND2_X1 U15093 ( .A1(b_6_), .A2(a_20_), .ZN(n15050) );
  XOR2_X1 U15094 ( .A(n15051), .B(n15052), .Z(n14877) );
  XNOR2_X1 U15095 ( .A(n15053), .B(n15054), .ZN(n15052) );
  NAND2_X1 U15096 ( .A1(b_5_), .A2(a_21_), .ZN(n15054) );
  INV_X1 U15097 ( .A(n15055), .ZN(n14878) );
  NOR2_X1 U15098 ( .A1(n9047), .A2(n15049), .ZN(n15055) );
  NOR2_X1 U15099 ( .A1(n15056), .A2(n15057), .ZN(n15049) );
  NOR3_X1 U15100 ( .A1(n8759), .A2(n15058), .A3(n14621), .ZN(n15057) );
  NOR2_X1 U15101 ( .A1(n14799), .A2(n14798), .ZN(n15058) );
  INV_X1 U15102 ( .A(n15059), .ZN(n15056) );
  NAND2_X1 U15103 ( .A1(n14798), .A2(n14799), .ZN(n15059) );
  NAND2_X1 U15104 ( .A1(n14807), .A2(n15060), .ZN(n14799) );
  NAND2_X1 U15105 ( .A1(n14806), .A2(n14808), .ZN(n15060) );
  NAND2_X1 U15106 ( .A1(n15061), .A2(n15062), .ZN(n14808) );
  NAND2_X1 U15107 ( .A1(b_6_), .A2(a_22_), .ZN(n15062) );
  XNOR2_X1 U15108 ( .A(n15063), .B(n15064), .ZN(n14806) );
  XOR2_X1 U15109 ( .A(n15065), .B(n15066), .Z(n15063) );
  NAND2_X1 U15110 ( .A1(a_22_), .A2(n15067), .ZN(n14807) );
  INV_X1 U15111 ( .A(n15061), .ZN(n15067) );
  NOR2_X1 U15112 ( .A1(n15068), .A2(n15069), .ZN(n15061) );
  NOR3_X1 U15113 ( .A1(n12301), .A2(n15070), .A3(n14621), .ZN(n15069) );
  INV_X1 U15114 ( .A(n15071), .ZN(n15070) );
  NAND2_X1 U15115 ( .A1(n14815), .A2(n14814), .ZN(n15071) );
  NOR2_X1 U15116 ( .A1(n14814), .A2(n14815), .ZN(n15068) );
  NOR2_X1 U15117 ( .A1(n15072), .A2(n15073), .ZN(n14815) );
  INV_X1 U15118 ( .A(n15074), .ZN(n15073) );
  NAND3_X1 U15119 ( .A1(a_24_), .A2(n15075), .A3(b_6_), .ZN(n15074) );
  NAND2_X1 U15120 ( .A1(n14874), .A2(n14873), .ZN(n15075) );
  NOR2_X1 U15121 ( .A1(n14873), .A2(n14874), .ZN(n15072) );
  NOR2_X1 U15122 ( .A1(n15076), .A2(n15077), .ZN(n14874) );
  INV_X1 U15123 ( .A(n15078), .ZN(n15077) );
  NAND2_X1 U15124 ( .A1(n14871), .A2(n15079), .ZN(n15078) );
  NAND2_X1 U15125 ( .A1(n14868), .A2(n14870), .ZN(n15079) );
  NOR2_X1 U15126 ( .A1(n14621), .A2(n8788), .ZN(n14871) );
  NOR2_X1 U15127 ( .A1(n14870), .A2(n14868), .ZN(n15076) );
  XNOR2_X1 U15128 ( .A(n15080), .B(n15081), .ZN(n14868) );
  XNOR2_X1 U15129 ( .A(n15082), .B(n15083), .ZN(n15081) );
  NAND2_X1 U15130 ( .A1(n15084), .A2(n15085), .ZN(n14870) );
  NAND2_X1 U15131 ( .A1(n14829), .A2(n15086), .ZN(n15085) );
  NAND2_X1 U15132 ( .A1(n14832), .A2(n14831), .ZN(n15086) );
  XNOR2_X1 U15133 ( .A(n15087), .B(n15088), .ZN(n14829) );
  XOR2_X1 U15134 ( .A(n15089), .B(n15090), .Z(n15087) );
  INV_X1 U15135 ( .A(n15091), .ZN(n15084) );
  NOR2_X1 U15136 ( .A1(n14831), .A2(n14832), .ZN(n15091) );
  NOR2_X1 U15137 ( .A1(n14621), .A2(n9344), .ZN(n14832) );
  NAND2_X1 U15138 ( .A1(n15092), .A2(n15093), .ZN(n14831) );
  NAND2_X1 U15139 ( .A1(n14839), .A2(n15094), .ZN(n15093) );
  INV_X1 U15140 ( .A(n15095), .ZN(n15094) );
  NOR2_X1 U15141 ( .A1(n14837), .A2(n14838), .ZN(n15095) );
  NOR2_X1 U15142 ( .A1(n14621), .A2(n8797), .ZN(n14839) );
  NAND2_X1 U15143 ( .A1(n14837), .A2(n14838), .ZN(n15092) );
  NAND2_X1 U15144 ( .A1(n15096), .A2(n15097), .ZN(n14838) );
  NAND2_X1 U15145 ( .A1(n14866), .A2(n15098), .ZN(n15097) );
  INV_X1 U15146 ( .A(n15099), .ZN(n15098) );
  NOR2_X1 U15147 ( .A1(n14867), .A2(n14865), .ZN(n15099) );
  NOR2_X1 U15148 ( .A1(n14621), .A2(n8314), .ZN(n14866) );
  NAND2_X1 U15149 ( .A1(n14865), .A2(n14867), .ZN(n15096) );
  NAND2_X1 U15150 ( .A1(n15100), .A2(n15101), .ZN(n14867) );
  NAND2_X1 U15151 ( .A1(n14861), .A2(n15102), .ZN(n15101) );
  INV_X1 U15152 ( .A(n15103), .ZN(n15102) );
  NOR2_X1 U15153 ( .A1(n14862), .A2(n14863), .ZN(n15103) );
  NOR2_X1 U15154 ( .A1(n14621), .A2(n9098), .ZN(n14861) );
  NAND2_X1 U15155 ( .A1(n14863), .A2(n14862), .ZN(n15100) );
  NAND2_X1 U15156 ( .A1(n15104), .A2(n15105), .ZN(n14862) );
  NAND2_X1 U15157 ( .A1(b_4_), .A2(n15106), .ZN(n15105) );
  NAND2_X1 U15158 ( .A1(n8299), .A2(n15107), .ZN(n15106) );
  NAND2_X1 U15159 ( .A1(a_31_), .A2(n14859), .ZN(n15107) );
  NAND2_X1 U15160 ( .A1(b_5_), .A2(n15108), .ZN(n15104) );
  NAND2_X1 U15161 ( .A1(n8303), .A2(n15109), .ZN(n15108) );
  NAND2_X1 U15162 ( .A1(a_30_), .A2(n15110), .ZN(n15109) );
  NOR3_X1 U15163 ( .A1(n14621), .A2(n9631), .A3(n14859), .ZN(n14863) );
  XOR2_X1 U15164 ( .A(n15111), .B(n15112), .Z(n14865) );
  XOR2_X1 U15165 ( .A(n15113), .B(n15114), .Z(n15111) );
  XOR2_X1 U15166 ( .A(n15115), .B(n15116), .Z(n14837) );
  XOR2_X1 U15167 ( .A(n15117), .B(n15118), .Z(n15115) );
  XNOR2_X1 U15168 ( .A(n15119), .B(n15120), .ZN(n14873) );
  XOR2_X1 U15169 ( .A(n15121), .B(n15122), .Z(n15120) );
  XNOR2_X1 U15170 ( .A(n15123), .B(n15124), .ZN(n14814) );
  XOR2_X1 U15171 ( .A(n15125), .B(n15126), .Z(n15123) );
  NOR2_X1 U15172 ( .A1(n8779), .A2(n14859), .ZN(n15126) );
  XOR2_X1 U15173 ( .A(n15127), .B(n15128), .Z(n14798) );
  XOR2_X1 U15174 ( .A(n15129), .B(n15130), .Z(n15127) );
  NOR2_X1 U15175 ( .A1(n12296), .A2(n14859), .ZN(n15130) );
  XNOR2_X1 U15176 ( .A(n15131), .B(n15132), .ZN(n14888) );
  XNOR2_X1 U15177 ( .A(n15133), .B(n15134), .ZN(n15131) );
  NOR2_X1 U15178 ( .A1(n14859), .A2(n9291), .ZN(n15134) );
  XNOR2_X1 U15179 ( .A(n15135), .B(n15136), .ZN(n14892) );
  XNOR2_X1 U15180 ( .A(n15137), .B(n15138), .ZN(n15135) );
  NOR2_X1 U15181 ( .A1(n14859), .A2(n8371), .ZN(n15138) );
  XNOR2_X1 U15182 ( .A(n15139), .B(n15140), .ZN(n14897) );
  XNOR2_X1 U15183 ( .A(n15141), .B(n15142), .ZN(n15139) );
  NOR2_X1 U15184 ( .A1(n14859), .A2(n8376), .ZN(n15142) );
  XOR2_X1 U15185 ( .A(n15143), .B(n15144), .Z(n14901) );
  XNOR2_X1 U15186 ( .A(n15145), .B(n15146), .ZN(n15143) );
  NOR2_X1 U15187 ( .A1(n14859), .A2(n8850), .ZN(n15146) );
  XOR2_X1 U15188 ( .A(n15147), .B(n15148), .Z(n14905) );
  XNOR2_X1 U15189 ( .A(n15149), .B(n15150), .ZN(n15147) );
  NOR2_X1 U15190 ( .A1(n14859), .A2(n9262), .ZN(n15150) );
  XOR2_X1 U15191 ( .A(n15151), .B(n15152), .Z(n14909) );
  XNOR2_X1 U15192 ( .A(n15153), .B(n15154), .ZN(n15151) );
  NOR2_X1 U15193 ( .A1(n14859), .A2(n8996), .ZN(n15154) );
  XOR2_X1 U15194 ( .A(n15155), .B(n15156), .Z(n14912) );
  XNOR2_X1 U15195 ( .A(n15157), .B(n15158), .ZN(n15155) );
  NOR2_X1 U15196 ( .A1(n14859), .A2(n8393), .ZN(n15158) );
  XNOR2_X1 U15197 ( .A(n15159), .B(n15160), .ZN(n14917) );
  XNOR2_X1 U15198 ( .A(n15161), .B(n15162), .ZN(n15159) );
  NOR2_X1 U15199 ( .A1(n14859), .A2(n8867), .ZN(n15162) );
  XNOR2_X1 U15200 ( .A(n15163), .B(n15164), .ZN(n14921) );
  XNOR2_X1 U15201 ( .A(n15165), .B(n15166), .ZN(n15163) );
  NOR2_X1 U15202 ( .A1(n14859), .A2(n8402), .ZN(n15166) );
  XOR2_X1 U15203 ( .A(n15167), .B(n15168), .Z(n14740) );
  XNOR2_X1 U15204 ( .A(n15169), .B(n15170), .ZN(n15167) );
  NOR2_X1 U15205 ( .A1(n14859), .A2(n8971), .ZN(n15170) );
  XOR2_X1 U15206 ( .A(n15171), .B(n15172), .Z(n14731) );
  XNOR2_X1 U15207 ( .A(n15173), .B(n15174), .ZN(n15171) );
  NOR2_X1 U15208 ( .A1(n14859), .A2(n8968), .ZN(n15174) );
  XNOR2_X1 U15209 ( .A(n15175), .B(n15176), .ZN(n14925) );
  XNOR2_X1 U15210 ( .A(n15177), .B(n15178), .ZN(n15175) );
  NOR2_X1 U15211 ( .A1(n14859), .A2(n8425), .ZN(n15178) );
  XOR2_X1 U15212 ( .A(n15179), .B(n15180), .Z(n14928) );
  XNOR2_X1 U15213 ( .A(n15181), .B(n15182), .ZN(n15179) );
  NOR2_X1 U15214 ( .A1(n14859), .A2(n8430), .ZN(n15182) );
  XNOR2_X1 U15215 ( .A(n15183), .B(n15184), .ZN(n14932) );
  XNOR2_X1 U15216 ( .A(n15185), .B(n15186), .ZN(n15184) );
  XNOR2_X1 U15217 ( .A(n15187), .B(n15188), .ZN(n14937) );
  XNOR2_X1 U15218 ( .A(n15189), .B(n15190), .ZN(n15187) );
  NOR2_X1 U15219 ( .A1(n14859), .A2(n8439), .ZN(n15190) );
  XNOR2_X1 U15220 ( .A(n15191), .B(n15192), .ZN(n14941) );
  XNOR2_X1 U15221 ( .A(n15193), .B(n15194), .ZN(n15191) );
  NOR2_X1 U15222 ( .A1(n14859), .A2(n8900), .ZN(n15194) );
  XNOR2_X1 U15223 ( .A(n15195), .B(n15196), .ZN(n14703) );
  XNOR2_X1 U15224 ( .A(n15197), .B(n15198), .ZN(n15195) );
  NOR2_X1 U15225 ( .A1(n14859), .A2(n8448), .ZN(n15198) );
  XNOR2_X1 U15226 ( .A(n15199), .B(n15200), .ZN(n14447) );
  XNOR2_X1 U15227 ( .A(n15201), .B(n15202), .ZN(n15199) );
  NOR2_X1 U15228 ( .A1(n14859), .A2(n8569), .ZN(n15202) );
  XNOR2_X1 U15229 ( .A(n15203), .B(n14957), .ZN(n8323) );
  XOR2_X1 U15230 ( .A(n15204), .B(n15205), .Z(n14957) );
  XNOR2_X1 U15231 ( .A(n15206), .B(n15207), .ZN(n15204) );
  XNOR2_X1 U15232 ( .A(n14956), .B(n15208), .ZN(n15203) );
  NOR2_X1 U15233 ( .A1(n14859), .A2(n8457), .ZN(n15208) );
  NOR2_X1 U15234 ( .A1(n15209), .A2(n15210), .ZN(n14956) );
  INV_X1 U15235 ( .A(n15211), .ZN(n15210) );
  NAND3_X1 U15236 ( .A1(b_5_), .A2(n15212), .A3(a_1_), .ZN(n15211) );
  NAND2_X1 U15237 ( .A1(n15200), .A2(n15201), .ZN(n15212) );
  NOR2_X1 U15238 ( .A1(n15200), .A2(n15201), .ZN(n15209) );
  NOR2_X1 U15239 ( .A1(n15213), .A2(n15214), .ZN(n15201) );
  INV_X1 U15240 ( .A(n15215), .ZN(n15214) );
  NAND3_X1 U15241 ( .A1(b_5_), .A2(n15216), .A3(a_2_), .ZN(n15215) );
  NAND2_X1 U15242 ( .A1(n15197), .A2(n15196), .ZN(n15216) );
  NOR2_X1 U15243 ( .A1(n15196), .A2(n15197), .ZN(n15213) );
  NOR2_X1 U15244 ( .A1(n15217), .A2(n15218), .ZN(n15197) );
  INV_X1 U15245 ( .A(n15219), .ZN(n15218) );
  NAND3_X1 U15246 ( .A1(b_5_), .A2(n15220), .A3(a_3_), .ZN(n15219) );
  NAND2_X1 U15247 ( .A1(n15193), .A2(n15192), .ZN(n15220) );
  NOR2_X1 U15248 ( .A1(n15192), .A2(n15193), .ZN(n15217) );
  NOR2_X1 U15249 ( .A1(n15221), .A2(n15222), .ZN(n15193) );
  INV_X1 U15250 ( .A(n15223), .ZN(n15222) );
  NAND3_X1 U15251 ( .A1(b_5_), .A2(n15224), .A3(a_4_), .ZN(n15223) );
  NAND2_X1 U15252 ( .A1(n15188), .A2(n15189), .ZN(n15224) );
  NOR2_X1 U15253 ( .A1(n15188), .A2(n15189), .ZN(n15221) );
  NOR2_X1 U15254 ( .A1(n15225), .A2(n15226), .ZN(n15189) );
  INV_X1 U15255 ( .A(n15227), .ZN(n15226) );
  NAND2_X1 U15256 ( .A1(n15183), .A2(n15228), .ZN(n15227) );
  NAND2_X1 U15257 ( .A1(n15186), .A2(n15185), .ZN(n15228) );
  XNOR2_X1 U15258 ( .A(n15229), .B(n15230), .ZN(n15183) );
  XNOR2_X1 U15259 ( .A(n15231), .B(n15232), .ZN(n15230) );
  NOR2_X1 U15260 ( .A1(n15185), .A2(n15186), .ZN(n15225) );
  NOR2_X1 U15261 ( .A1(n15233), .A2(n15234), .ZN(n15186) );
  INV_X1 U15262 ( .A(n15235), .ZN(n15234) );
  NAND3_X1 U15263 ( .A1(b_5_), .A2(n15236), .A3(a_6_), .ZN(n15235) );
  NAND2_X1 U15264 ( .A1(n15180), .A2(n15181), .ZN(n15236) );
  NOR2_X1 U15265 ( .A1(n15180), .A2(n15181), .ZN(n15233) );
  NOR2_X1 U15266 ( .A1(n15237), .A2(n15238), .ZN(n15181) );
  INV_X1 U15267 ( .A(n15239), .ZN(n15238) );
  NAND3_X1 U15268 ( .A1(b_5_), .A2(n15240), .A3(a_7_), .ZN(n15239) );
  NAND2_X1 U15269 ( .A1(n15177), .A2(n15176), .ZN(n15240) );
  NOR2_X1 U15270 ( .A1(n15176), .A2(n15177), .ZN(n15237) );
  NOR2_X1 U15271 ( .A1(n15241), .A2(n15242), .ZN(n15177) );
  NOR3_X1 U15272 ( .A1(n14859), .A2(n15243), .A3(n8968), .ZN(n15242) );
  INV_X1 U15273 ( .A(n15244), .ZN(n15243) );
  NAND2_X1 U15274 ( .A1(n15172), .A2(n15173), .ZN(n15244) );
  NOR2_X1 U15275 ( .A1(n15172), .A2(n15173), .ZN(n15241) );
  NOR2_X1 U15276 ( .A1(n15245), .A2(n15246), .ZN(n15173) );
  INV_X1 U15277 ( .A(n15247), .ZN(n15246) );
  NAND3_X1 U15278 ( .A1(b_5_), .A2(n15248), .A3(a_9_), .ZN(n15247) );
  NAND2_X1 U15279 ( .A1(n15169), .A2(n15168), .ZN(n15248) );
  NOR2_X1 U15280 ( .A1(n15168), .A2(n15169), .ZN(n15245) );
  NOR2_X1 U15281 ( .A1(n15249), .A2(n15250), .ZN(n15169) );
  NOR3_X1 U15282 ( .A1(n14859), .A2(n15251), .A3(n8402), .ZN(n15250) );
  INV_X1 U15283 ( .A(n15252), .ZN(n15251) );
  NAND2_X1 U15284 ( .A1(n15164), .A2(n15165), .ZN(n15252) );
  NOR2_X1 U15285 ( .A1(n15164), .A2(n15165), .ZN(n15249) );
  NOR2_X1 U15286 ( .A1(n15253), .A2(n15254), .ZN(n15165) );
  INV_X1 U15287 ( .A(n15255), .ZN(n15254) );
  NAND3_X1 U15288 ( .A1(b_5_), .A2(n15256), .A3(a_11_), .ZN(n15255) );
  NAND2_X1 U15289 ( .A1(n15161), .A2(n15160), .ZN(n15256) );
  NOR2_X1 U15290 ( .A1(n15160), .A2(n15161), .ZN(n15253) );
  NOR2_X1 U15291 ( .A1(n15257), .A2(n15258), .ZN(n15161) );
  NOR3_X1 U15292 ( .A1(n14859), .A2(n15259), .A3(n8393), .ZN(n15258) );
  INV_X1 U15293 ( .A(n15260), .ZN(n15259) );
  NAND2_X1 U15294 ( .A1(n15156), .A2(n15157), .ZN(n15260) );
  NOR2_X1 U15295 ( .A1(n15156), .A2(n15157), .ZN(n15257) );
  NOR2_X1 U15296 ( .A1(n15261), .A2(n15262), .ZN(n15157) );
  INV_X1 U15297 ( .A(n15263), .ZN(n15262) );
  NAND3_X1 U15298 ( .A1(b_5_), .A2(n15264), .A3(a_13_), .ZN(n15263) );
  NAND2_X1 U15299 ( .A1(n15152), .A2(n15153), .ZN(n15264) );
  NOR2_X1 U15300 ( .A1(n15152), .A2(n15153), .ZN(n15261) );
  NOR2_X1 U15301 ( .A1(n15265), .A2(n15266), .ZN(n15153) );
  INV_X1 U15302 ( .A(n15267), .ZN(n15266) );
  NAND3_X1 U15303 ( .A1(b_5_), .A2(n15268), .A3(a_14_), .ZN(n15267) );
  NAND2_X1 U15304 ( .A1(n15148), .A2(n15149), .ZN(n15268) );
  NOR2_X1 U15305 ( .A1(n15148), .A2(n15149), .ZN(n15265) );
  NOR2_X1 U15306 ( .A1(n15269), .A2(n15270), .ZN(n15149) );
  INV_X1 U15307 ( .A(n15271), .ZN(n15270) );
  NAND3_X1 U15308 ( .A1(b_5_), .A2(n15272), .A3(a_15_), .ZN(n15271) );
  NAND2_X1 U15309 ( .A1(n15145), .A2(n15144), .ZN(n15272) );
  NOR2_X1 U15310 ( .A1(n15144), .A2(n15145), .ZN(n15269) );
  NOR2_X1 U15311 ( .A1(n15273), .A2(n15274), .ZN(n15145) );
  NOR3_X1 U15312 ( .A1(n14859), .A2(n15275), .A3(n8376), .ZN(n15274) );
  INV_X1 U15313 ( .A(n15276), .ZN(n15275) );
  NAND2_X1 U15314 ( .A1(n15140), .A2(n15141), .ZN(n15276) );
  NOR2_X1 U15315 ( .A1(n15140), .A2(n15141), .ZN(n15273) );
  NOR2_X1 U15316 ( .A1(n15277), .A2(n15278), .ZN(n15141) );
  INV_X1 U15317 ( .A(n15279), .ZN(n15278) );
  NAND3_X1 U15318 ( .A1(b_5_), .A2(n15280), .A3(a_17_), .ZN(n15279) );
  NAND2_X1 U15319 ( .A1(n15137), .A2(n15136), .ZN(n15280) );
  NOR2_X1 U15320 ( .A1(n15136), .A2(n15137), .ZN(n15277) );
  NOR2_X1 U15321 ( .A1(n15281), .A2(n15282), .ZN(n15137) );
  NOR3_X1 U15322 ( .A1(n14859), .A2(n15283), .A3(n9291), .ZN(n15282) );
  INV_X1 U15323 ( .A(n15284), .ZN(n15283) );
  NAND2_X1 U15324 ( .A1(n15132), .A2(n15133), .ZN(n15284) );
  NOR2_X1 U15325 ( .A1(n15132), .A2(n15133), .ZN(n15281) );
  NOR2_X1 U15326 ( .A1(n15285), .A2(n15286), .ZN(n15133) );
  INV_X1 U15327 ( .A(n15287), .ZN(n15286) );
  NAND3_X1 U15328 ( .A1(a_19_), .A2(n15288), .A3(b_5_), .ZN(n15287) );
  NAND2_X1 U15329 ( .A1(n15038), .A2(n15037), .ZN(n15288) );
  NOR2_X1 U15330 ( .A1(n15037), .A2(n15038), .ZN(n15285) );
  NOR2_X1 U15331 ( .A1(n15289), .A2(n15290), .ZN(n15038) );
  NOR3_X1 U15332 ( .A1(n9047), .A2(n15291), .A3(n14859), .ZN(n15290) );
  NOR2_X1 U15333 ( .A1(n15045), .A2(n15046), .ZN(n15291) );
  INV_X1 U15334 ( .A(n15292), .ZN(n15289) );
  NAND2_X1 U15335 ( .A1(n15045), .A2(n15046), .ZN(n15292) );
  NAND2_X1 U15336 ( .A1(n15293), .A2(n15294), .ZN(n15046) );
  NAND3_X1 U15337 ( .A1(a_21_), .A2(n15295), .A3(b_5_), .ZN(n15294) );
  NAND2_X1 U15338 ( .A1(n15051), .A2(n15053), .ZN(n15295) );
  INV_X1 U15339 ( .A(n15296), .ZN(n15293) );
  NOR2_X1 U15340 ( .A1(n15051), .A2(n15053), .ZN(n15296) );
  NOR2_X1 U15341 ( .A1(n15297), .A2(n15298), .ZN(n15053) );
  INV_X1 U15342 ( .A(n15299), .ZN(n15298) );
  NAND3_X1 U15343 ( .A1(a_22_), .A2(n15300), .A3(b_5_), .ZN(n15299) );
  NAND2_X1 U15344 ( .A1(n15128), .A2(n15129), .ZN(n15300) );
  NOR2_X1 U15345 ( .A1(n15128), .A2(n15129), .ZN(n15297) );
  NAND2_X1 U15346 ( .A1(n15301), .A2(n15302), .ZN(n15129) );
  NAND2_X1 U15347 ( .A1(n15064), .A2(n15303), .ZN(n15302) );
  NAND2_X1 U15348 ( .A1(n15066), .A2(n15065), .ZN(n15303) );
  XOR2_X1 U15349 ( .A(n15304), .B(n15305), .Z(n15064) );
  XNOR2_X1 U15350 ( .A(n15306), .B(n15307), .ZN(n15304) );
  INV_X1 U15351 ( .A(n15308), .ZN(n15301) );
  NOR2_X1 U15352 ( .A1(n15065), .A2(n15066), .ZN(n15308) );
  NOR2_X1 U15353 ( .A1(n14859), .A2(n12301), .ZN(n15066) );
  NAND2_X1 U15354 ( .A1(n15309), .A2(n15310), .ZN(n15065) );
  NAND3_X1 U15355 ( .A1(a_24_), .A2(n15311), .A3(b_5_), .ZN(n15310) );
  INV_X1 U15356 ( .A(n15312), .ZN(n15311) );
  NOR2_X1 U15357 ( .A1(n15124), .A2(n15125), .ZN(n15312) );
  NAND2_X1 U15358 ( .A1(n15124), .A2(n15125), .ZN(n15309) );
  NAND2_X1 U15359 ( .A1(n15313), .A2(n15314), .ZN(n15125) );
  NAND2_X1 U15360 ( .A1(n15122), .A2(n15315), .ZN(n15314) );
  INV_X1 U15361 ( .A(n15316), .ZN(n15315) );
  NOR2_X1 U15362 ( .A1(n15119), .A2(n15121), .ZN(n15316) );
  NOR2_X1 U15363 ( .A1(n14859), .A2(n8788), .ZN(n15122) );
  NAND2_X1 U15364 ( .A1(n15119), .A2(n15121), .ZN(n15313) );
  NOR2_X1 U15365 ( .A1(n15317), .A2(n15318), .ZN(n15121) );
  INV_X1 U15366 ( .A(n15319), .ZN(n15318) );
  NAND2_X1 U15367 ( .A1(n15080), .A2(n15320), .ZN(n15319) );
  NAND2_X1 U15368 ( .A1(n15083), .A2(n15082), .ZN(n15320) );
  XNOR2_X1 U15369 ( .A(n15321), .B(n15322), .ZN(n15080) );
  XOR2_X1 U15370 ( .A(n15323), .B(n15324), .Z(n15321) );
  NOR2_X1 U15371 ( .A1(n8797), .A2(n15110), .ZN(n15324) );
  NOR2_X1 U15372 ( .A1(n15082), .A2(n15083), .ZN(n15317) );
  NOR2_X1 U15373 ( .A1(n14859), .A2(n9344), .ZN(n15083) );
  NAND2_X1 U15374 ( .A1(n15325), .A2(n15326), .ZN(n15082) );
  NAND2_X1 U15375 ( .A1(n15090), .A2(n15327), .ZN(n15326) );
  INV_X1 U15376 ( .A(n15328), .ZN(n15327) );
  NOR2_X1 U15377 ( .A1(n15088), .A2(n15089), .ZN(n15328) );
  NOR2_X1 U15378 ( .A1(n14859), .A2(n8797), .ZN(n15090) );
  NAND2_X1 U15379 ( .A1(n15088), .A2(n15089), .ZN(n15325) );
  NAND2_X1 U15380 ( .A1(n15329), .A2(n15330), .ZN(n15089) );
  NAND2_X1 U15381 ( .A1(n15117), .A2(n15331), .ZN(n15330) );
  INV_X1 U15382 ( .A(n15332), .ZN(n15331) );
  NOR2_X1 U15383 ( .A1(n15118), .A2(n15116), .ZN(n15332) );
  NOR2_X1 U15384 ( .A1(n14859), .A2(n8314), .ZN(n15117) );
  NAND2_X1 U15385 ( .A1(n15116), .A2(n15118), .ZN(n15329) );
  NAND2_X1 U15386 ( .A1(n15333), .A2(n15334), .ZN(n15118) );
  NAND2_X1 U15387 ( .A1(n15112), .A2(n15335), .ZN(n15334) );
  INV_X1 U15388 ( .A(n15336), .ZN(n15335) );
  NOR2_X1 U15389 ( .A1(n15113), .A2(n15114), .ZN(n15336) );
  NOR2_X1 U15390 ( .A1(n14859), .A2(n9098), .ZN(n15112) );
  NAND2_X1 U15391 ( .A1(n15114), .A2(n15113), .ZN(n15333) );
  NAND2_X1 U15392 ( .A1(n15337), .A2(n15338), .ZN(n15113) );
  NAND2_X1 U15393 ( .A1(b_3_), .A2(n15339), .ZN(n15338) );
  NAND2_X1 U15394 ( .A1(n8299), .A2(n15340), .ZN(n15339) );
  NAND2_X1 U15395 ( .A1(a_31_), .A2(n15110), .ZN(n15340) );
  NAND2_X1 U15396 ( .A1(b_4_), .A2(n15341), .ZN(n15337) );
  NAND2_X1 U15397 ( .A1(n8303), .A2(n15342), .ZN(n15341) );
  NAND2_X1 U15398 ( .A1(a_30_), .A2(n15343), .ZN(n15342) );
  NOR3_X1 U15399 ( .A1(n14859), .A2(n9631), .A3(n15110), .ZN(n15114) );
  XOR2_X1 U15400 ( .A(n15344), .B(n15345), .Z(n15116) );
  XOR2_X1 U15401 ( .A(n15346), .B(n15347), .Z(n15344) );
  XOR2_X1 U15402 ( .A(n15348), .B(n15349), .Z(n15088) );
  XOR2_X1 U15403 ( .A(n15350), .B(n15351), .Z(n15348) );
  XOR2_X1 U15404 ( .A(n15352), .B(n15353), .Z(n15119) );
  XNOR2_X1 U15405 ( .A(n15354), .B(n15355), .ZN(n15353) );
  XNOR2_X1 U15406 ( .A(n15356), .B(n15357), .ZN(n15124) );
  XNOR2_X1 U15407 ( .A(n15358), .B(n15359), .ZN(n15357) );
  XNOR2_X1 U15408 ( .A(n15360), .B(n15361), .ZN(n15128) );
  XOR2_X1 U15409 ( .A(n15362), .B(n15363), .Z(n15360) );
  XOR2_X1 U15410 ( .A(n15364), .B(n15365), .Z(n15051) );
  XOR2_X1 U15411 ( .A(n15366), .B(n15367), .Z(n15365) );
  XNOR2_X1 U15412 ( .A(n15368), .B(n15369), .ZN(n15045) );
  XNOR2_X1 U15413 ( .A(n15370), .B(n15371), .ZN(n15368) );
  XNOR2_X1 U15414 ( .A(n15372), .B(n15373), .ZN(n15037) );
  XOR2_X1 U15415 ( .A(n15374), .B(n15375), .Z(n15373) );
  XOR2_X1 U15416 ( .A(n15376), .B(n15377), .Z(n15132) );
  XNOR2_X1 U15417 ( .A(n15378), .B(n15379), .ZN(n15376) );
  XOR2_X1 U15418 ( .A(n15380), .B(n15381), .Z(n15136) );
  XOR2_X1 U15419 ( .A(n15382), .B(n15383), .Z(n15381) );
  XNOR2_X1 U15420 ( .A(n15384), .B(n15385), .ZN(n15140) );
  XOR2_X1 U15421 ( .A(n15386), .B(n15387), .Z(n15384) );
  XOR2_X1 U15422 ( .A(n15388), .B(n15389), .Z(n15144) );
  XNOR2_X1 U15423 ( .A(n15390), .B(n15391), .ZN(n15389) );
  XNOR2_X1 U15424 ( .A(n15392), .B(n15393), .ZN(n15148) );
  XOR2_X1 U15425 ( .A(n15394), .B(n15395), .Z(n15392) );
  XOR2_X1 U15426 ( .A(n15396), .B(n15397), .Z(n15152) );
  XNOR2_X1 U15427 ( .A(n15398), .B(n15399), .ZN(n15397) );
  XNOR2_X1 U15428 ( .A(n15400), .B(n15401), .ZN(n15156) );
  XOR2_X1 U15429 ( .A(n15402), .B(n15403), .Z(n15400) );
  XOR2_X1 U15430 ( .A(n15404), .B(n15405), .Z(n15160) );
  XNOR2_X1 U15431 ( .A(n15406), .B(n15407), .ZN(n15405) );
  XNOR2_X1 U15432 ( .A(n15408), .B(n15409), .ZN(n15164) );
  XOR2_X1 U15433 ( .A(n15410), .B(n15411), .Z(n15408) );
  XOR2_X1 U15434 ( .A(n15412), .B(n15413), .Z(n15168) );
  XNOR2_X1 U15435 ( .A(n15414), .B(n15415), .ZN(n15413) );
  XNOR2_X1 U15436 ( .A(n15416), .B(n15417), .ZN(n15172) );
  XOR2_X1 U15437 ( .A(n15418), .B(n15419), .Z(n15416) );
  XOR2_X1 U15438 ( .A(n15420), .B(n15421), .Z(n15176) );
  XNOR2_X1 U15439 ( .A(n15422), .B(n15423), .ZN(n15421) );
  XNOR2_X1 U15440 ( .A(n15424), .B(n15425), .ZN(n15180) );
  XOR2_X1 U15441 ( .A(n15426), .B(n15427), .Z(n15424) );
  XNOR2_X1 U15442 ( .A(n15428), .B(n15429), .ZN(n15188) );
  XOR2_X1 U15443 ( .A(n15430), .B(n15431), .Z(n15428) );
  XOR2_X1 U15444 ( .A(n15432), .B(n15433), .Z(n15192) );
  XOR2_X1 U15445 ( .A(n15434), .B(n15435), .Z(n15433) );
  XOR2_X1 U15446 ( .A(n15436), .B(n15437), .Z(n15196) );
  XNOR2_X1 U15447 ( .A(n15438), .B(n15439), .ZN(n15436) );
  XNOR2_X1 U15448 ( .A(n15440), .B(n15441), .ZN(n15200) );
  XNOR2_X1 U15449 ( .A(n15442), .B(n15443), .ZN(n15441) );
  XNOR2_X1 U15450 ( .A(n8419), .B(n8418), .ZN(n8366) );
  NAND3_X1 U15451 ( .A1(n8419), .A2(n8418), .A3(n8416), .ZN(n8420) );
  NOR2_X1 U15452 ( .A1(n15444), .A2(n8574), .ZN(n8416) );
  NOR2_X1 U15453 ( .A1(n15445), .A2(n15446), .ZN(n8574) );
  INV_X1 U15454 ( .A(n15447), .ZN(n15446) );
  XOR2_X1 U15455 ( .A(n15448), .B(n15449), .Z(n15445) );
  NOR2_X1 U15456 ( .A1(n15447), .A2(n15450), .ZN(n15444) );
  XNOR2_X1 U15457 ( .A(n15448), .B(n15449), .ZN(n15450) );
  NAND2_X1 U15458 ( .A1(n15451), .A2(n15452), .ZN(n15448) );
  NAND2_X1 U15459 ( .A1(n15453), .A2(n15454), .ZN(n15447) );
  INV_X1 U15460 ( .A(n15455), .ZN(n15454) );
  NOR3_X1 U15461 ( .A1(n15343), .A2(n15456), .A3(n8457), .ZN(n15455) );
  NOR2_X1 U15462 ( .A1(n15457), .A2(n15458), .ZN(n15456) );
  NAND2_X1 U15463 ( .A1(n15458), .A2(n15457), .ZN(n15453) );
  NAND2_X1 U15464 ( .A1(n15459), .A2(n15460), .ZN(n8418) );
  NAND2_X1 U15465 ( .A1(n14951), .A2(n15461), .ZN(n15460) );
  INV_X1 U15466 ( .A(n15462), .ZN(n15461) );
  NOR2_X1 U15467 ( .A1(n14949), .A2(n14950), .ZN(n15462) );
  NOR2_X1 U15468 ( .A1(n8457), .A2(n15110), .ZN(n14951) );
  NAND2_X1 U15469 ( .A1(n14949), .A2(n14950), .ZN(n15459) );
  NAND2_X1 U15470 ( .A1(n15463), .A2(n15464), .ZN(n14950) );
  NAND2_X1 U15471 ( .A1(n15207), .A2(n15465), .ZN(n15464) );
  NAND2_X1 U15472 ( .A1(n15205), .A2(n15206), .ZN(n15465) );
  NOR2_X1 U15473 ( .A1(n8569), .A2(n15110), .ZN(n15207) );
  INV_X1 U15474 ( .A(n15466), .ZN(n15463) );
  NOR2_X1 U15475 ( .A1(n15205), .A2(n15206), .ZN(n15466) );
  NOR2_X1 U15476 ( .A1(n15467), .A2(n15468), .ZN(n15206) );
  INV_X1 U15477 ( .A(n15469), .ZN(n15468) );
  NAND2_X1 U15478 ( .A1(n15443), .A2(n15470), .ZN(n15469) );
  NAND2_X1 U15479 ( .A1(n15471), .A2(n15440), .ZN(n15470) );
  NOR2_X1 U15480 ( .A1(n8448), .A2(n15110), .ZN(n15443) );
  NOR2_X1 U15481 ( .A1(n15440), .A2(n15471), .ZN(n15467) );
  INV_X1 U15482 ( .A(n15442), .ZN(n15471) );
  NAND2_X1 U15483 ( .A1(n15472), .A2(n15473), .ZN(n15442) );
  NAND2_X1 U15484 ( .A1(n15439), .A2(n15474), .ZN(n15473) );
  INV_X1 U15485 ( .A(n15475), .ZN(n15474) );
  NOR2_X1 U15486 ( .A1(n15437), .A2(n15438), .ZN(n15475) );
  NOR2_X1 U15487 ( .A1(n8900), .A2(n15110), .ZN(n15439) );
  NAND2_X1 U15488 ( .A1(n15437), .A2(n15438), .ZN(n15472) );
  NOR2_X1 U15489 ( .A1(n15476), .A2(n15477), .ZN(n15438) );
  INV_X1 U15490 ( .A(n15478), .ZN(n15477) );
  NAND2_X1 U15491 ( .A1(n15479), .A2(n15434), .ZN(n15478) );
  NAND2_X1 U15492 ( .A1(n15432), .A2(n15435), .ZN(n15479) );
  NOR2_X1 U15493 ( .A1(n15432), .A2(n15435), .ZN(n15476) );
  NAND2_X1 U15494 ( .A1(n15480), .A2(n15481), .ZN(n15435) );
  NAND2_X1 U15495 ( .A1(n15431), .A2(n15482), .ZN(n15481) );
  INV_X1 U15496 ( .A(n15483), .ZN(n15482) );
  NOR2_X1 U15497 ( .A1(n15430), .A2(n15429), .ZN(n15483) );
  NOR2_X1 U15498 ( .A1(n8938), .A2(n15110), .ZN(n15431) );
  NAND2_X1 U15499 ( .A1(n15429), .A2(n15430), .ZN(n15480) );
  NAND2_X1 U15500 ( .A1(n15484), .A2(n15485), .ZN(n15430) );
  NAND2_X1 U15501 ( .A1(n15232), .A2(n15486), .ZN(n15485) );
  INV_X1 U15502 ( .A(n15487), .ZN(n15486) );
  NOR2_X1 U15503 ( .A1(n15229), .A2(n15231), .ZN(n15487) );
  NOR2_X1 U15504 ( .A1(n8430), .A2(n15110), .ZN(n15232) );
  NAND2_X1 U15505 ( .A1(n15229), .A2(n15231), .ZN(n15484) );
  NAND2_X1 U15506 ( .A1(n15488), .A2(n15489), .ZN(n15231) );
  NAND2_X1 U15507 ( .A1(n15427), .A2(n15490), .ZN(n15489) );
  INV_X1 U15508 ( .A(n15491), .ZN(n15490) );
  NOR2_X1 U15509 ( .A1(n15426), .A2(n15425), .ZN(n15491) );
  NOR2_X1 U15510 ( .A1(n8425), .A2(n15110), .ZN(n15427) );
  NAND2_X1 U15511 ( .A1(n15425), .A2(n15426), .ZN(n15488) );
  NAND2_X1 U15512 ( .A1(n15492), .A2(n15493), .ZN(n15426) );
  NAND2_X1 U15513 ( .A1(n15423), .A2(n15494), .ZN(n15493) );
  INV_X1 U15514 ( .A(n15495), .ZN(n15494) );
  NOR2_X1 U15515 ( .A1(n15420), .A2(n15422), .ZN(n15495) );
  NOR2_X1 U15516 ( .A1(n8968), .A2(n15110), .ZN(n15423) );
  NAND2_X1 U15517 ( .A1(n15420), .A2(n15422), .ZN(n15492) );
  NAND2_X1 U15518 ( .A1(n15496), .A2(n15497), .ZN(n15422) );
  NAND2_X1 U15519 ( .A1(n15419), .A2(n15498), .ZN(n15497) );
  INV_X1 U15520 ( .A(n15499), .ZN(n15498) );
  NOR2_X1 U15521 ( .A1(n15418), .A2(n15417), .ZN(n15499) );
  NOR2_X1 U15522 ( .A1(n8971), .A2(n15110), .ZN(n15419) );
  NAND2_X1 U15523 ( .A1(n15417), .A2(n15418), .ZN(n15496) );
  NAND2_X1 U15524 ( .A1(n15500), .A2(n15501), .ZN(n15418) );
  NAND2_X1 U15525 ( .A1(n15415), .A2(n15502), .ZN(n15501) );
  INV_X1 U15526 ( .A(n15503), .ZN(n15502) );
  NOR2_X1 U15527 ( .A1(n15412), .A2(n15414), .ZN(n15503) );
  NOR2_X1 U15528 ( .A1(n8402), .A2(n15110), .ZN(n15415) );
  NAND2_X1 U15529 ( .A1(n15412), .A2(n15414), .ZN(n15500) );
  NAND2_X1 U15530 ( .A1(n15504), .A2(n15505), .ZN(n15414) );
  NAND2_X1 U15531 ( .A1(n15411), .A2(n15506), .ZN(n15505) );
  INV_X1 U15532 ( .A(n15507), .ZN(n15506) );
  NOR2_X1 U15533 ( .A1(n15410), .A2(n15409), .ZN(n15507) );
  NOR2_X1 U15534 ( .A1(n8867), .A2(n15110), .ZN(n15411) );
  NAND2_X1 U15535 ( .A1(n15409), .A2(n15410), .ZN(n15504) );
  NAND2_X1 U15536 ( .A1(n15508), .A2(n15509), .ZN(n15410) );
  NAND2_X1 U15537 ( .A1(n15407), .A2(n15510), .ZN(n15509) );
  INV_X1 U15538 ( .A(n15511), .ZN(n15510) );
  NOR2_X1 U15539 ( .A1(n15404), .A2(n15406), .ZN(n15511) );
  NOR2_X1 U15540 ( .A1(n8393), .A2(n15110), .ZN(n15407) );
  NAND2_X1 U15541 ( .A1(n15404), .A2(n15406), .ZN(n15508) );
  NAND2_X1 U15542 ( .A1(n15512), .A2(n15513), .ZN(n15406) );
  NAND2_X1 U15543 ( .A1(n15402), .A2(n15514), .ZN(n15513) );
  INV_X1 U15544 ( .A(n15515), .ZN(n15514) );
  NOR2_X1 U15545 ( .A1(n15403), .A2(n15401), .ZN(n15515) );
  NOR2_X1 U15546 ( .A1(n8996), .A2(n15110), .ZN(n15402) );
  NAND2_X1 U15547 ( .A1(n15401), .A2(n15403), .ZN(n15512) );
  NAND2_X1 U15548 ( .A1(n15516), .A2(n15517), .ZN(n15403) );
  NAND2_X1 U15549 ( .A1(n15399), .A2(n15518), .ZN(n15517) );
  INV_X1 U15550 ( .A(n15519), .ZN(n15518) );
  NOR2_X1 U15551 ( .A1(n15398), .A2(n15396), .ZN(n15519) );
  NOR2_X1 U15552 ( .A1(n9262), .A2(n15110), .ZN(n15399) );
  NAND2_X1 U15553 ( .A1(n15396), .A2(n15398), .ZN(n15516) );
  NAND2_X1 U15554 ( .A1(n15520), .A2(n15521), .ZN(n15398) );
  NAND2_X1 U15555 ( .A1(n15395), .A2(n15522), .ZN(n15521) );
  INV_X1 U15556 ( .A(n15523), .ZN(n15522) );
  NOR2_X1 U15557 ( .A1(n15394), .A2(n15393), .ZN(n15523) );
  NOR2_X1 U15558 ( .A1(n8850), .A2(n15110), .ZN(n15395) );
  NAND2_X1 U15559 ( .A1(n15393), .A2(n15394), .ZN(n15520) );
  NAND2_X1 U15560 ( .A1(n15524), .A2(n15525), .ZN(n15394) );
  NAND2_X1 U15561 ( .A1(n15391), .A2(n15526), .ZN(n15525) );
  INV_X1 U15562 ( .A(n15527), .ZN(n15526) );
  NOR2_X1 U15563 ( .A1(n15388), .A2(n15390), .ZN(n15527) );
  NOR2_X1 U15564 ( .A1(n8376), .A2(n15110), .ZN(n15391) );
  NAND2_X1 U15565 ( .A1(n15388), .A2(n15390), .ZN(n15524) );
  NAND2_X1 U15566 ( .A1(n15528), .A2(n15529), .ZN(n15390) );
  NAND2_X1 U15567 ( .A1(n15387), .A2(n15530), .ZN(n15529) );
  INV_X1 U15568 ( .A(n15531), .ZN(n15530) );
  NOR2_X1 U15569 ( .A1(n15386), .A2(n15385), .ZN(n15531) );
  NOR2_X1 U15570 ( .A1(n8371), .A2(n15110), .ZN(n15387) );
  NAND2_X1 U15571 ( .A1(n15385), .A2(n15386), .ZN(n15528) );
  NAND2_X1 U15572 ( .A1(n15532), .A2(n15533), .ZN(n15386) );
  NAND2_X1 U15573 ( .A1(n15383), .A2(n15534), .ZN(n15533) );
  NAND2_X1 U15574 ( .A1(n15535), .A2(n15382), .ZN(n15534) );
  INV_X1 U15575 ( .A(n15380), .ZN(n15535) );
  NOR2_X1 U15576 ( .A1(n9291), .A2(n15110), .ZN(n15383) );
  NAND2_X1 U15577 ( .A1(n15380), .A2(n15536), .ZN(n15532) );
  INV_X1 U15578 ( .A(n15382), .ZN(n15536) );
  NOR2_X1 U15579 ( .A1(n15537), .A2(n15538), .ZN(n15382) );
  INV_X1 U15580 ( .A(n15539), .ZN(n15538) );
  NAND2_X1 U15581 ( .A1(n15379), .A2(n15540), .ZN(n15539) );
  NAND2_X1 U15582 ( .A1(n15378), .A2(n15377), .ZN(n15540) );
  NOR2_X1 U15583 ( .A1(n15110), .A2(n8742), .ZN(n15379) );
  NOR2_X1 U15584 ( .A1(n15377), .A2(n15378), .ZN(n15537) );
  NOR2_X1 U15585 ( .A1(n15541), .A2(n15542), .ZN(n15378) );
  INV_X1 U15586 ( .A(n15543), .ZN(n15542) );
  NAND2_X1 U15587 ( .A1(n15375), .A2(n15544), .ZN(n15543) );
  NAND2_X1 U15588 ( .A1(n15372), .A2(n15374), .ZN(n15544) );
  NOR2_X1 U15589 ( .A1(n15110), .A2(n9047), .ZN(n15375) );
  NOR2_X1 U15590 ( .A1(n15372), .A2(n15374), .ZN(n15541) );
  NOR2_X1 U15591 ( .A1(n15545), .A2(n15546), .ZN(n15374) );
  INV_X1 U15592 ( .A(n15547), .ZN(n15546) );
  NAND2_X1 U15593 ( .A1(n15370), .A2(n15548), .ZN(n15547) );
  NAND2_X1 U15594 ( .A1(n15371), .A2(n15369), .ZN(n15548) );
  NOR2_X1 U15595 ( .A1(n15110), .A2(n8759), .ZN(n15370) );
  NOR2_X1 U15596 ( .A1(n15369), .A2(n15371), .ZN(n15545) );
  NOR2_X1 U15597 ( .A1(n15549), .A2(n15550), .ZN(n15371) );
  NOR2_X1 U15598 ( .A1(n15367), .A2(n15551), .ZN(n15550) );
  NOR2_X1 U15599 ( .A1(n15366), .A2(n15364), .ZN(n15551) );
  NAND2_X1 U15600 ( .A1(b_4_), .A2(a_22_), .ZN(n15367) );
  INV_X1 U15601 ( .A(n15552), .ZN(n15549) );
  NAND2_X1 U15602 ( .A1(n15364), .A2(n15366), .ZN(n15552) );
  NAND2_X1 U15603 ( .A1(n15553), .A2(n15554), .ZN(n15366) );
  NAND2_X1 U15604 ( .A1(n15363), .A2(n15555), .ZN(n15554) );
  INV_X1 U15605 ( .A(n15556), .ZN(n15555) );
  NOR2_X1 U15606 ( .A1(n15361), .A2(n15362), .ZN(n15556) );
  NOR2_X1 U15607 ( .A1(n15110), .A2(n12301), .ZN(n15363) );
  NAND2_X1 U15608 ( .A1(n15361), .A2(n15362), .ZN(n15553) );
  NAND2_X1 U15609 ( .A1(n15557), .A2(n15558), .ZN(n15362) );
  NAND2_X1 U15610 ( .A1(n15307), .A2(n15559), .ZN(n15558) );
  NAND2_X1 U15611 ( .A1(n15305), .A2(n15306), .ZN(n15559) );
  NOR2_X1 U15612 ( .A1(n15110), .A2(n8779), .ZN(n15307) );
  INV_X1 U15613 ( .A(n15560), .ZN(n15557) );
  NOR2_X1 U15614 ( .A1(n15305), .A2(n15306), .ZN(n15560) );
  NOR2_X1 U15615 ( .A1(n15561), .A2(n15562), .ZN(n15306) );
  INV_X1 U15616 ( .A(n15563), .ZN(n15562) );
  NAND2_X1 U15617 ( .A1(n15359), .A2(n15564), .ZN(n15563) );
  NAND2_X1 U15618 ( .A1(n15356), .A2(n15358), .ZN(n15564) );
  NOR2_X1 U15619 ( .A1(n15110), .A2(n8788), .ZN(n15359) );
  NOR2_X1 U15620 ( .A1(n15358), .A2(n15356), .ZN(n15561) );
  XOR2_X1 U15621 ( .A(n15565), .B(n15566), .Z(n15356) );
  XNOR2_X1 U15622 ( .A(n15567), .B(n15568), .ZN(n15566) );
  NAND2_X1 U15623 ( .A1(n15569), .A2(n15570), .ZN(n15358) );
  NAND2_X1 U15624 ( .A1(n15352), .A2(n15571), .ZN(n15570) );
  INV_X1 U15625 ( .A(n15572), .ZN(n15571) );
  NOR2_X1 U15626 ( .A1(n15355), .A2(n15354), .ZN(n15572) );
  XOR2_X1 U15627 ( .A(n15573), .B(n15574), .Z(n15352) );
  XNOR2_X1 U15628 ( .A(n15575), .B(n15576), .ZN(n15573) );
  NAND2_X1 U15629 ( .A1(n15354), .A2(n15355), .ZN(n15569) );
  NAND2_X1 U15630 ( .A1(b_4_), .A2(a_26_), .ZN(n15355) );
  NOR2_X1 U15631 ( .A1(n15577), .A2(n15578), .ZN(n15354) );
  NOR3_X1 U15632 ( .A1(n8797), .A2(n15579), .A3(n15110), .ZN(n15578) );
  NOR2_X1 U15633 ( .A1(n15322), .A2(n15323), .ZN(n15579) );
  INV_X1 U15634 ( .A(n15580), .ZN(n15577) );
  NAND2_X1 U15635 ( .A1(n15322), .A2(n15323), .ZN(n15580) );
  NAND2_X1 U15636 ( .A1(n15581), .A2(n15582), .ZN(n15323) );
  NAND2_X1 U15637 ( .A1(n15350), .A2(n15583), .ZN(n15582) );
  INV_X1 U15638 ( .A(n15584), .ZN(n15583) );
  NOR2_X1 U15639 ( .A1(n15351), .A2(n15349), .ZN(n15584) );
  NOR2_X1 U15640 ( .A1(n15110), .A2(n8314), .ZN(n15350) );
  NAND2_X1 U15641 ( .A1(n15349), .A2(n15351), .ZN(n15581) );
  NAND2_X1 U15642 ( .A1(n15585), .A2(n15586), .ZN(n15351) );
  NAND2_X1 U15643 ( .A1(n15345), .A2(n15587), .ZN(n15586) );
  INV_X1 U15644 ( .A(n15588), .ZN(n15587) );
  NOR2_X1 U15645 ( .A1(n15346), .A2(n15347), .ZN(n15588) );
  NOR2_X1 U15646 ( .A1(n15110), .A2(n9098), .ZN(n15345) );
  NAND2_X1 U15647 ( .A1(n15347), .A2(n15346), .ZN(n15585) );
  NAND2_X1 U15648 ( .A1(n15589), .A2(n15590), .ZN(n15346) );
  NAND2_X1 U15649 ( .A1(b_2_), .A2(n15591), .ZN(n15590) );
  NAND2_X1 U15650 ( .A1(n8299), .A2(n15592), .ZN(n15591) );
  NAND2_X1 U15651 ( .A1(a_31_), .A2(n15343), .ZN(n15592) );
  NAND2_X1 U15652 ( .A1(b_3_), .A2(n15593), .ZN(n15589) );
  NAND2_X1 U15653 ( .A1(n8303), .A2(n15594), .ZN(n15593) );
  NAND2_X1 U15654 ( .A1(a_30_), .A2(n15595), .ZN(n15594) );
  NOR3_X1 U15655 ( .A1(n15110), .A2(n9631), .A3(n15343), .ZN(n15347) );
  XOR2_X1 U15656 ( .A(n15596), .B(n15597), .Z(n15349) );
  XNOR2_X1 U15657 ( .A(n15598), .B(n15599), .ZN(n15596) );
  XNOR2_X1 U15658 ( .A(n15600), .B(n15601), .ZN(n15322) );
  XNOR2_X1 U15659 ( .A(n15602), .B(n15603), .ZN(n15600) );
  XOR2_X1 U15660 ( .A(n15604), .B(n15605), .Z(n15305) );
  NAND2_X1 U15661 ( .A1(n15606), .A2(n15607), .ZN(n15604) );
  XOR2_X1 U15662 ( .A(n15608), .B(n15609), .Z(n15361) );
  XOR2_X1 U15663 ( .A(n15610), .B(n15611), .Z(n15608) );
  NOR2_X1 U15664 ( .A1(n8779), .A2(n15343), .ZN(n15611) );
  XNOR2_X1 U15665 ( .A(n15612), .B(n15613), .ZN(n15364) );
  NAND2_X1 U15666 ( .A1(n15614), .A2(n15615), .ZN(n15612) );
  XNOR2_X1 U15667 ( .A(n15616), .B(n15617), .ZN(n15369) );
  XOR2_X1 U15668 ( .A(n15618), .B(n15619), .Z(n15616) );
  NOR2_X1 U15669 ( .A1(n12296), .A2(n15343), .ZN(n15619) );
  XOR2_X1 U15670 ( .A(n15620), .B(n15621), .Z(n15372) );
  NAND2_X1 U15671 ( .A1(n15622), .A2(n15623), .ZN(n15620) );
  XNOR2_X1 U15672 ( .A(n15624), .B(n15625), .ZN(n15377) );
  XOR2_X1 U15673 ( .A(n15626), .B(n15627), .Z(n15624) );
  NOR2_X1 U15674 ( .A1(n9047), .A2(n15343), .ZN(n15627) );
  XNOR2_X1 U15675 ( .A(n15628), .B(n15629), .ZN(n15380) );
  NAND2_X1 U15676 ( .A1(n15630), .A2(n15631), .ZN(n15628) );
  XOR2_X1 U15677 ( .A(n15632), .B(n15633), .Z(n15385) );
  XOR2_X1 U15678 ( .A(n15634), .B(n15635), .Z(n15632) );
  NOR2_X1 U15679 ( .A1(n15343), .A2(n9291), .ZN(n15635) );
  XNOR2_X1 U15680 ( .A(n15636), .B(n15637), .ZN(n15388) );
  NAND2_X1 U15681 ( .A1(n15638), .A2(n15639), .ZN(n15636) );
  XOR2_X1 U15682 ( .A(n15640), .B(n15641), .Z(n15393) );
  XOR2_X1 U15683 ( .A(n15642), .B(n15643), .Z(n15640) );
  NOR2_X1 U15684 ( .A1(n15343), .A2(n8376), .ZN(n15643) );
  XNOR2_X1 U15685 ( .A(n15644), .B(n15645), .ZN(n15396) );
  NAND2_X1 U15686 ( .A1(n15646), .A2(n15647), .ZN(n15644) );
  XOR2_X1 U15687 ( .A(n15648), .B(n15649), .Z(n15401) );
  XOR2_X1 U15688 ( .A(n15650), .B(n15651), .Z(n15648) );
  NOR2_X1 U15689 ( .A1(n15343), .A2(n9262), .ZN(n15651) );
  XNOR2_X1 U15690 ( .A(n15652), .B(n15653), .ZN(n15404) );
  NAND2_X1 U15691 ( .A1(n15654), .A2(n15655), .ZN(n15652) );
  XOR2_X1 U15692 ( .A(n15656), .B(n15657), .Z(n15409) );
  XOR2_X1 U15693 ( .A(n15658), .B(n15659), .Z(n15656) );
  NOR2_X1 U15694 ( .A1(n15343), .A2(n8393), .ZN(n15659) );
  XNOR2_X1 U15695 ( .A(n15660), .B(n15661), .ZN(n15412) );
  NAND2_X1 U15696 ( .A1(n15662), .A2(n15663), .ZN(n15660) );
  XOR2_X1 U15697 ( .A(n15664), .B(n15665), .Z(n15417) );
  XOR2_X1 U15698 ( .A(n15666), .B(n15667), .Z(n15664) );
  NOR2_X1 U15699 ( .A1(n15343), .A2(n8402), .ZN(n15667) );
  XNOR2_X1 U15700 ( .A(n15668), .B(n15669), .ZN(n15420) );
  NAND2_X1 U15701 ( .A1(n15670), .A2(n15671), .ZN(n15668) );
  XOR2_X1 U15702 ( .A(n15672), .B(n15673), .Z(n15425) );
  XOR2_X1 U15703 ( .A(n15674), .B(n15675), .Z(n15672) );
  NOR2_X1 U15704 ( .A1(n15343), .A2(n8968), .ZN(n15675) );
  XNOR2_X1 U15705 ( .A(n15676), .B(n15677), .ZN(n15229) );
  NAND2_X1 U15706 ( .A1(n15678), .A2(n15679), .ZN(n15676) );
  XOR2_X1 U15707 ( .A(n15680), .B(n15681), .Z(n15429) );
  XOR2_X1 U15708 ( .A(n15682), .B(n15683), .Z(n15680) );
  NOR2_X1 U15709 ( .A1(n15343), .A2(n8430), .ZN(n15683) );
  XNOR2_X1 U15710 ( .A(n15684), .B(n15685), .ZN(n15432) );
  NAND2_X1 U15711 ( .A1(n15686), .A2(n15687), .ZN(n15684) );
  XOR2_X1 U15712 ( .A(n15688), .B(n15689), .Z(n15437) );
  XOR2_X1 U15713 ( .A(n15690), .B(n15691), .Z(n15688) );
  NOR2_X1 U15714 ( .A1(n15343), .A2(n8439), .ZN(n15691) );
  XOR2_X1 U15715 ( .A(n15692), .B(n15693), .Z(n15440) );
  XNOR2_X1 U15716 ( .A(n15694), .B(n15695), .ZN(n15692) );
  XOR2_X1 U15717 ( .A(n15696), .B(n15697), .Z(n15205) );
  XOR2_X1 U15718 ( .A(n15698), .B(n15699), .Z(n15697) );
  NAND2_X1 U15719 ( .A1(a_2_), .A2(b_3_), .ZN(n15699) );
  XNOR2_X1 U15720 ( .A(n15700), .B(n15701), .ZN(n14949) );
  NAND2_X1 U15721 ( .A1(n15702), .A2(n15703), .ZN(n15700) );
  XOR2_X1 U15722 ( .A(n15704), .B(n15458), .Z(n8419) );
  XNOR2_X1 U15723 ( .A(n15705), .B(n15706), .ZN(n15458) );
  XOR2_X1 U15724 ( .A(n15707), .B(n15708), .Z(n15706) );
  NAND2_X1 U15725 ( .A1(a_1_), .A2(b_2_), .ZN(n15708) );
  XOR2_X1 U15726 ( .A(n15457), .B(n15709), .Z(n15704) );
  NOR2_X1 U15727 ( .A1(n15343), .A2(n8457), .ZN(n15709) );
  NAND2_X1 U15728 ( .A1(n15702), .A2(n15710), .ZN(n15457) );
  NAND2_X1 U15729 ( .A1(n15701), .A2(n15703), .ZN(n15710) );
  NAND2_X1 U15730 ( .A1(n15711), .A2(n15712), .ZN(n15703) );
  NAND2_X1 U15731 ( .A1(a_1_), .A2(b_3_), .ZN(n15712) );
  XNOR2_X1 U15732 ( .A(n15713), .B(n15714), .ZN(n15701) );
  XNOR2_X1 U15733 ( .A(n15715), .B(n15716), .ZN(n15713) );
  INV_X1 U15734 ( .A(n15717), .ZN(n15702) );
  NOR2_X1 U15735 ( .A1(n8569), .A2(n15711), .ZN(n15717) );
  NOR2_X1 U15736 ( .A1(n15718), .A2(n15719), .ZN(n15711) );
  NOR3_X1 U15737 ( .A1(n15343), .A2(n15720), .A3(n8448), .ZN(n15719) );
  INV_X1 U15738 ( .A(n15721), .ZN(n15720) );
  NAND2_X1 U15739 ( .A1(n15696), .A2(n15698), .ZN(n15721) );
  NOR2_X1 U15740 ( .A1(n15698), .A2(n15696), .ZN(n15718) );
  XOR2_X1 U15741 ( .A(n15722), .B(n15723), .Z(n15696) );
  XNOR2_X1 U15742 ( .A(n15724), .B(n15725), .ZN(n15722) );
  NAND2_X1 U15743 ( .A1(n15726), .A2(n15727), .ZN(n15698) );
  NAND2_X1 U15744 ( .A1(n15693), .A2(n15728), .ZN(n15727) );
  NAND2_X1 U15745 ( .A1(n15695), .A2(n15729), .ZN(n15728) );
  XOR2_X1 U15746 ( .A(n15730), .B(n15731), .Z(n15693) );
  XNOR2_X1 U15747 ( .A(n15732), .B(n15733), .ZN(n15730) );
  INV_X1 U15748 ( .A(n15734), .ZN(n15726) );
  NOR2_X1 U15749 ( .A1(n15729), .A2(n15695), .ZN(n15734) );
  INV_X1 U15750 ( .A(n15694), .ZN(n15729) );
  NOR2_X1 U15751 ( .A1(n15735), .A2(n15736), .ZN(n15694) );
  NOR3_X1 U15752 ( .A1(n15343), .A2(n15737), .A3(n8439), .ZN(n15736) );
  NOR2_X1 U15753 ( .A1(n15689), .A2(n15690), .ZN(n15737) );
  INV_X1 U15754 ( .A(n15738), .ZN(n15735) );
  NAND2_X1 U15755 ( .A1(n15689), .A2(n15690), .ZN(n15738) );
  NAND2_X1 U15756 ( .A1(n15686), .A2(n15739), .ZN(n15690) );
  NAND2_X1 U15757 ( .A1(n15685), .A2(n15687), .ZN(n15739) );
  NAND2_X1 U15758 ( .A1(n15740), .A2(n15741), .ZN(n15687) );
  NAND2_X1 U15759 ( .A1(a_5_), .A2(b_3_), .ZN(n15741) );
  XNOR2_X1 U15760 ( .A(n15742), .B(n15743), .ZN(n15685) );
  XNOR2_X1 U15761 ( .A(n15744), .B(n15745), .ZN(n15742) );
  NAND2_X1 U15762 ( .A1(a_5_), .A2(n15746), .ZN(n15686) );
  INV_X1 U15763 ( .A(n15740), .ZN(n15746) );
  NOR2_X1 U15764 ( .A1(n15747), .A2(n15748), .ZN(n15740) );
  NOR3_X1 U15765 ( .A1(n15343), .A2(n15749), .A3(n8430), .ZN(n15748) );
  NOR2_X1 U15766 ( .A1(n15681), .A2(n15682), .ZN(n15749) );
  INV_X1 U15767 ( .A(n15750), .ZN(n15747) );
  NAND2_X1 U15768 ( .A1(n15681), .A2(n15682), .ZN(n15750) );
  NAND2_X1 U15769 ( .A1(n15678), .A2(n15751), .ZN(n15682) );
  NAND2_X1 U15770 ( .A1(n15677), .A2(n15679), .ZN(n15751) );
  NAND2_X1 U15771 ( .A1(n15752), .A2(n15753), .ZN(n15679) );
  NAND2_X1 U15772 ( .A1(a_7_), .A2(b_3_), .ZN(n15753) );
  XNOR2_X1 U15773 ( .A(n15754), .B(n15755), .ZN(n15677) );
  XNOR2_X1 U15774 ( .A(n15756), .B(n15757), .ZN(n15754) );
  NAND2_X1 U15775 ( .A1(a_7_), .A2(n15758), .ZN(n15678) );
  INV_X1 U15776 ( .A(n15752), .ZN(n15758) );
  NOR2_X1 U15777 ( .A1(n15759), .A2(n15760), .ZN(n15752) );
  NOR3_X1 U15778 ( .A1(n15343), .A2(n15761), .A3(n8968), .ZN(n15760) );
  NOR2_X1 U15779 ( .A1(n15673), .A2(n15674), .ZN(n15761) );
  INV_X1 U15780 ( .A(n15762), .ZN(n15759) );
  NAND2_X1 U15781 ( .A1(n15673), .A2(n15674), .ZN(n15762) );
  NAND2_X1 U15782 ( .A1(n15670), .A2(n15763), .ZN(n15674) );
  NAND2_X1 U15783 ( .A1(n15669), .A2(n15671), .ZN(n15763) );
  NAND2_X1 U15784 ( .A1(n15764), .A2(n15765), .ZN(n15671) );
  NAND2_X1 U15785 ( .A1(a_9_), .A2(b_3_), .ZN(n15765) );
  INV_X1 U15786 ( .A(n15766), .ZN(n15764) );
  XNOR2_X1 U15787 ( .A(n15767), .B(n15768), .ZN(n15669) );
  XNOR2_X1 U15788 ( .A(n15769), .B(n15770), .ZN(n15767) );
  NAND2_X1 U15789 ( .A1(a_9_), .A2(n15766), .ZN(n15670) );
  NAND2_X1 U15790 ( .A1(n15771), .A2(n15772), .ZN(n15766) );
  INV_X1 U15791 ( .A(n15773), .ZN(n15772) );
  NOR3_X1 U15792 ( .A1(n15343), .A2(n15774), .A3(n8402), .ZN(n15773) );
  NOR2_X1 U15793 ( .A1(n15665), .A2(n15666), .ZN(n15774) );
  NAND2_X1 U15794 ( .A1(n15665), .A2(n15666), .ZN(n15771) );
  NAND2_X1 U15795 ( .A1(n15662), .A2(n15775), .ZN(n15666) );
  NAND2_X1 U15796 ( .A1(n15661), .A2(n15663), .ZN(n15775) );
  NAND2_X1 U15797 ( .A1(n15776), .A2(n15777), .ZN(n15663) );
  NAND2_X1 U15798 ( .A1(a_11_), .A2(b_3_), .ZN(n15777) );
  INV_X1 U15799 ( .A(n15778), .ZN(n15776) );
  XNOR2_X1 U15800 ( .A(n15779), .B(n15780), .ZN(n15661) );
  XNOR2_X1 U15801 ( .A(n15781), .B(n15782), .ZN(n15779) );
  NAND2_X1 U15802 ( .A1(a_11_), .A2(n15778), .ZN(n15662) );
  NAND2_X1 U15803 ( .A1(n15783), .A2(n15784), .ZN(n15778) );
  INV_X1 U15804 ( .A(n15785), .ZN(n15784) );
  NOR3_X1 U15805 ( .A1(n15343), .A2(n15786), .A3(n8393), .ZN(n15785) );
  NOR2_X1 U15806 ( .A1(n15657), .A2(n15658), .ZN(n15786) );
  NAND2_X1 U15807 ( .A1(n15657), .A2(n15658), .ZN(n15783) );
  NAND2_X1 U15808 ( .A1(n15654), .A2(n15787), .ZN(n15658) );
  NAND2_X1 U15809 ( .A1(n15653), .A2(n15655), .ZN(n15787) );
  NAND2_X1 U15810 ( .A1(n15788), .A2(n15789), .ZN(n15655) );
  NAND2_X1 U15811 ( .A1(a_13_), .A2(b_3_), .ZN(n15789) );
  INV_X1 U15812 ( .A(n15790), .ZN(n15788) );
  XNOR2_X1 U15813 ( .A(n15791), .B(n15792), .ZN(n15653) );
  XNOR2_X1 U15814 ( .A(n15793), .B(n15794), .ZN(n15791) );
  NAND2_X1 U15815 ( .A1(a_13_), .A2(n15790), .ZN(n15654) );
  NAND2_X1 U15816 ( .A1(n15795), .A2(n15796), .ZN(n15790) );
  INV_X1 U15817 ( .A(n15797), .ZN(n15796) );
  NOR3_X1 U15818 ( .A1(n15343), .A2(n15798), .A3(n9262), .ZN(n15797) );
  NOR2_X1 U15819 ( .A1(n15649), .A2(n15650), .ZN(n15798) );
  NAND2_X1 U15820 ( .A1(n15649), .A2(n15650), .ZN(n15795) );
  NAND2_X1 U15821 ( .A1(n15646), .A2(n15799), .ZN(n15650) );
  NAND2_X1 U15822 ( .A1(n15645), .A2(n15647), .ZN(n15799) );
  NAND2_X1 U15823 ( .A1(n15800), .A2(n15801), .ZN(n15647) );
  NAND2_X1 U15824 ( .A1(a_15_), .A2(b_3_), .ZN(n15801) );
  INV_X1 U15825 ( .A(n15802), .ZN(n15800) );
  XNOR2_X1 U15826 ( .A(n15803), .B(n15804), .ZN(n15645) );
  XNOR2_X1 U15827 ( .A(n15805), .B(n15806), .ZN(n15804) );
  NAND2_X1 U15828 ( .A1(a_15_), .A2(n15802), .ZN(n15646) );
  NAND2_X1 U15829 ( .A1(n15807), .A2(n15808), .ZN(n15802) );
  INV_X1 U15830 ( .A(n15809), .ZN(n15808) );
  NOR3_X1 U15831 ( .A1(n15343), .A2(n15810), .A3(n8376), .ZN(n15809) );
  NOR2_X1 U15832 ( .A1(n15641), .A2(n15642), .ZN(n15810) );
  NAND2_X1 U15833 ( .A1(n15641), .A2(n15642), .ZN(n15807) );
  NAND2_X1 U15834 ( .A1(n15638), .A2(n15811), .ZN(n15642) );
  NAND2_X1 U15835 ( .A1(n15637), .A2(n15639), .ZN(n15811) );
  NAND2_X1 U15836 ( .A1(n15812), .A2(n15813), .ZN(n15639) );
  NAND2_X1 U15837 ( .A1(a_17_), .A2(b_3_), .ZN(n15813) );
  INV_X1 U15838 ( .A(n15814), .ZN(n15812) );
  XNOR2_X1 U15839 ( .A(n15815), .B(n15816), .ZN(n15637) );
  XNOR2_X1 U15840 ( .A(n15817), .B(n15818), .ZN(n15816) );
  NAND2_X1 U15841 ( .A1(a_17_), .A2(n15814), .ZN(n15638) );
  NAND2_X1 U15842 ( .A1(n15819), .A2(n15820), .ZN(n15814) );
  INV_X1 U15843 ( .A(n15821), .ZN(n15820) );
  NOR3_X1 U15844 ( .A1(n15343), .A2(n15822), .A3(n9291), .ZN(n15821) );
  NOR2_X1 U15845 ( .A1(n15633), .A2(n15634), .ZN(n15822) );
  NAND2_X1 U15846 ( .A1(n15633), .A2(n15634), .ZN(n15819) );
  NAND2_X1 U15847 ( .A1(n15630), .A2(n15823), .ZN(n15634) );
  NAND2_X1 U15848 ( .A1(n15629), .A2(n15631), .ZN(n15823) );
  NAND2_X1 U15849 ( .A1(n15824), .A2(n15825), .ZN(n15631) );
  NAND2_X1 U15850 ( .A1(b_3_), .A2(a_19_), .ZN(n15825) );
  INV_X1 U15851 ( .A(n15826), .ZN(n15824) );
  XNOR2_X1 U15852 ( .A(n15827), .B(n15828), .ZN(n15629) );
  XNOR2_X1 U15853 ( .A(n15829), .B(n15830), .ZN(n15828) );
  NAND2_X1 U15854 ( .A1(a_19_), .A2(n15826), .ZN(n15630) );
  NAND2_X1 U15855 ( .A1(n15831), .A2(n15832), .ZN(n15826) );
  INV_X1 U15856 ( .A(n15833), .ZN(n15832) );
  NOR3_X1 U15857 ( .A1(n9047), .A2(n15834), .A3(n15343), .ZN(n15833) );
  NOR2_X1 U15858 ( .A1(n15625), .A2(n15626), .ZN(n15834) );
  NAND2_X1 U15859 ( .A1(n15625), .A2(n15626), .ZN(n15831) );
  NAND2_X1 U15860 ( .A1(n15622), .A2(n15835), .ZN(n15626) );
  NAND2_X1 U15861 ( .A1(n15621), .A2(n15623), .ZN(n15835) );
  NAND2_X1 U15862 ( .A1(n15836), .A2(n15837), .ZN(n15623) );
  NAND2_X1 U15863 ( .A1(b_3_), .A2(a_21_), .ZN(n15837) );
  INV_X1 U15864 ( .A(n15838), .ZN(n15836) );
  XNOR2_X1 U15865 ( .A(n15839), .B(n15840), .ZN(n15621) );
  XOR2_X1 U15866 ( .A(n15841), .B(n15842), .Z(n15840) );
  NAND2_X1 U15867 ( .A1(a_21_), .A2(n15838), .ZN(n15622) );
  NAND2_X1 U15868 ( .A1(n15843), .A2(n15844), .ZN(n15838) );
  INV_X1 U15869 ( .A(n15845), .ZN(n15844) );
  NOR3_X1 U15870 ( .A1(n12296), .A2(n15846), .A3(n15343), .ZN(n15845) );
  NOR2_X1 U15871 ( .A1(n15617), .A2(n15618), .ZN(n15846) );
  NAND2_X1 U15872 ( .A1(n15617), .A2(n15618), .ZN(n15843) );
  NAND2_X1 U15873 ( .A1(n15614), .A2(n15847), .ZN(n15618) );
  NAND2_X1 U15874 ( .A1(n15613), .A2(n15615), .ZN(n15847) );
  NAND2_X1 U15875 ( .A1(n15848), .A2(n15849), .ZN(n15615) );
  NAND2_X1 U15876 ( .A1(b_3_), .A2(a_23_), .ZN(n15849) );
  XNOR2_X1 U15877 ( .A(n15850), .B(n15851), .ZN(n15613) );
  NAND2_X1 U15878 ( .A1(n15852), .A2(n15853), .ZN(n15850) );
  INV_X1 U15879 ( .A(n15854), .ZN(n15614) );
  NOR2_X1 U15880 ( .A1(n12301), .A2(n15848), .ZN(n15854) );
  NOR2_X1 U15881 ( .A1(n15855), .A2(n15856), .ZN(n15848) );
  NOR3_X1 U15882 ( .A1(n8779), .A2(n15857), .A3(n15343), .ZN(n15856) );
  NOR2_X1 U15883 ( .A1(n15610), .A2(n15609), .ZN(n15857) );
  INV_X1 U15884 ( .A(n15858), .ZN(n15855) );
  NAND2_X1 U15885 ( .A1(n15609), .A2(n15610), .ZN(n15858) );
  NAND2_X1 U15886 ( .A1(n15606), .A2(n15859), .ZN(n15610) );
  NAND2_X1 U15887 ( .A1(n15605), .A2(n15607), .ZN(n15859) );
  NAND2_X1 U15888 ( .A1(n15860), .A2(n15861), .ZN(n15607) );
  NAND2_X1 U15889 ( .A1(b_3_), .A2(a_25_), .ZN(n15861) );
  INV_X1 U15890 ( .A(n15862), .ZN(n15860) );
  XNOR2_X1 U15891 ( .A(n15863), .B(n15864), .ZN(n15605) );
  XNOR2_X1 U15892 ( .A(n15865), .B(n15866), .ZN(n15864) );
  NOR2_X1 U15893 ( .A1(n9344), .A2(n15595), .ZN(n15866) );
  NAND2_X1 U15894 ( .A1(a_25_), .A2(n15862), .ZN(n15606) );
  NAND2_X1 U15895 ( .A1(n15867), .A2(n15868), .ZN(n15862) );
  NAND2_X1 U15896 ( .A1(n15568), .A2(n15869), .ZN(n15868) );
  INV_X1 U15897 ( .A(n15870), .ZN(n15869) );
  NOR2_X1 U15898 ( .A1(n15567), .A2(n15565), .ZN(n15870) );
  NOR2_X1 U15899 ( .A1(n15343), .A2(n9344), .ZN(n15568) );
  NAND2_X1 U15900 ( .A1(n15565), .A2(n15567), .ZN(n15867) );
  NAND2_X1 U15901 ( .A1(n15871), .A2(n15872), .ZN(n15567) );
  NAND2_X1 U15902 ( .A1(n15576), .A2(n15873), .ZN(n15872) );
  NAND2_X1 U15903 ( .A1(n15575), .A2(n15574), .ZN(n15873) );
  NOR2_X1 U15904 ( .A1(n15343), .A2(n8797), .ZN(n15576) );
  INV_X1 U15905 ( .A(n15874), .ZN(n15871) );
  NOR2_X1 U15906 ( .A1(n15574), .A2(n15575), .ZN(n15874) );
  NOR2_X1 U15907 ( .A1(n15875), .A2(n15876), .ZN(n15575) );
  INV_X1 U15908 ( .A(n15877), .ZN(n15876) );
  NAND2_X1 U15909 ( .A1(n15602), .A2(n15878), .ZN(n15877) );
  NAND2_X1 U15910 ( .A1(n15603), .A2(n15601), .ZN(n15878) );
  NOR2_X1 U15911 ( .A1(n15343), .A2(n8314), .ZN(n15602) );
  NOR2_X1 U15912 ( .A1(n15601), .A2(n15603), .ZN(n15875) );
  NOR2_X1 U15913 ( .A1(n15879), .A2(n15880), .ZN(n15603) );
  INV_X1 U15914 ( .A(n15881), .ZN(n15880) );
  NAND2_X1 U15915 ( .A1(n15597), .A2(n15882), .ZN(n15881) );
  NAND2_X1 U15916 ( .A1(n15883), .A2(n15599), .ZN(n15882) );
  NOR2_X1 U15917 ( .A1(n15343), .A2(n9098), .ZN(n15597) );
  NOR2_X1 U15918 ( .A1(n15599), .A2(n15883), .ZN(n15879) );
  INV_X1 U15919 ( .A(n15598), .ZN(n15883) );
  NAND2_X1 U15920 ( .A1(n15884), .A2(n15885), .ZN(n15598) );
  NAND2_X1 U15921 ( .A1(b_1_), .A2(n15886), .ZN(n15885) );
  NAND2_X1 U15922 ( .A1(n8299), .A2(n15887), .ZN(n15886) );
  NAND2_X1 U15923 ( .A1(a_31_), .A2(n15595), .ZN(n15887) );
  NAND2_X1 U15924 ( .A1(b_2_), .A2(n15888), .ZN(n15884) );
  NAND2_X1 U15925 ( .A1(n8303), .A2(n15889), .ZN(n15888) );
  NAND2_X1 U15926 ( .A1(a_30_), .A2(n15890), .ZN(n15889) );
  NAND3_X1 U15927 ( .A1(b_3_), .A2(n9106), .A3(b_2_), .ZN(n15599) );
  XNOR2_X1 U15928 ( .A(n15891), .B(n15892), .ZN(n15601) );
  XOR2_X1 U15929 ( .A(n15893), .B(n15894), .Z(n15891) );
  XNOR2_X1 U15930 ( .A(n15895), .B(n15896), .ZN(n15574) );
  XNOR2_X1 U15931 ( .A(n15897), .B(n15898), .ZN(n15895) );
  NAND2_X1 U15932 ( .A1(b_2_), .A2(a_28_), .ZN(n15897) );
  XNOR2_X1 U15933 ( .A(n15899), .B(n15900), .ZN(n15565) );
  NAND2_X1 U15934 ( .A1(n15901), .A2(n15902), .ZN(n15899) );
  XNOR2_X1 U15935 ( .A(n15903), .B(n15904), .ZN(n15609) );
  NAND2_X1 U15936 ( .A1(n15905), .A2(n15906), .ZN(n15903) );
  XNOR2_X1 U15937 ( .A(n15907), .B(n15908), .ZN(n15617) );
  XNOR2_X1 U15938 ( .A(n15909), .B(n15910), .ZN(n15908) );
  XNOR2_X1 U15939 ( .A(n15911), .B(n15912), .ZN(n15625) );
  XNOR2_X1 U15940 ( .A(n15913), .B(n15914), .ZN(n15911) );
  XOR2_X1 U15941 ( .A(n15915), .B(n15916), .Z(n15633) );
  XOR2_X1 U15942 ( .A(n15917), .B(n15918), .Z(n15915) );
  XNOR2_X1 U15943 ( .A(n15919), .B(n15920), .ZN(n15641) );
  XOR2_X1 U15944 ( .A(n15921), .B(n15922), .Z(n15920) );
  XNOR2_X1 U15945 ( .A(n15923), .B(n15924), .ZN(n15649) );
  XNOR2_X1 U15946 ( .A(n15925), .B(n15926), .ZN(n15923) );
  XNOR2_X1 U15947 ( .A(n15927), .B(n15928), .ZN(n15657) );
  XNOR2_X1 U15948 ( .A(n15929), .B(n15930), .ZN(n15927) );
  XNOR2_X1 U15949 ( .A(n15931), .B(n15932), .ZN(n15665) );
  XNOR2_X1 U15950 ( .A(n15933), .B(n15934), .ZN(n15931) );
  XNOR2_X1 U15951 ( .A(n15935), .B(n15936), .ZN(n15673) );
  XNOR2_X1 U15952 ( .A(n15937), .B(n15938), .ZN(n15935) );
  XNOR2_X1 U15953 ( .A(n15939), .B(n15940), .ZN(n15681) );
  XNOR2_X1 U15954 ( .A(n15941), .B(n15942), .ZN(n15939) );
  XNOR2_X1 U15955 ( .A(n15943), .B(n15944), .ZN(n15689) );
  XNOR2_X1 U15956 ( .A(n15945), .B(n15946), .ZN(n15943) );
  XNOR2_X1 U15957 ( .A(n8562), .B(n8561), .ZN(n8465) );
  XOR2_X1 U15958 ( .A(n15947), .B(n15948), .Z(n8561) );
  NOR2_X1 U15959 ( .A1(n8567), .A2(n8569), .ZN(n15948) );
  XOR2_X1 U15960 ( .A(n8570), .B(n8571), .Z(n15947) );
  NOR2_X1 U15961 ( .A1(n8457), .A2(n15890), .ZN(n8571) );
  NAND2_X1 U15962 ( .A1(n15949), .A2(n15950), .ZN(n8570) );
  NAND2_X1 U15963 ( .A1(n15951), .A2(n15952), .ZN(n15950) );
  INV_X1 U15964 ( .A(n15953), .ZN(n15952) );
  NOR2_X1 U15965 ( .A1(n15954), .A2(n15955), .ZN(n15953) );
  NAND2_X1 U15966 ( .A1(n15955), .A2(n15954), .ZN(n15949) );
  NAND2_X1 U15967 ( .A1(n15451), .A2(n15956), .ZN(n8562) );
  NAND2_X1 U15968 ( .A1(n15449), .A2(n15452), .ZN(n15956) );
  NAND2_X1 U15969 ( .A1(n15957), .A2(n15958), .ZN(n15452) );
  NAND2_X1 U15970 ( .A1(a_0_), .A2(b_2_), .ZN(n15958) );
  XOR2_X1 U15971 ( .A(n15959), .B(n15951), .Z(n15449) );
  NOR2_X1 U15972 ( .A1(n8448), .A2(n8567), .ZN(n15951) );
  XOR2_X1 U15973 ( .A(n15954), .B(n15955), .Z(n15959) );
  NAND2_X1 U15974 ( .A1(n15960), .A2(n15961), .ZN(n15954) );
  NAND2_X1 U15975 ( .A1(n15962), .A2(n15963), .ZN(n15961) );
  INV_X1 U15976 ( .A(n15964), .ZN(n15963) );
  NOR2_X1 U15977 ( .A1(n15965), .A2(n15966), .ZN(n15964) );
  NAND2_X1 U15978 ( .A1(n15966), .A2(n15965), .ZN(n15960) );
  NAND2_X1 U15979 ( .A1(a_0_), .A2(n15967), .ZN(n15451) );
  INV_X1 U15980 ( .A(n15957), .ZN(n15967) );
  NOR2_X1 U15981 ( .A1(n15968), .A2(n15969), .ZN(n15957) );
  NOR3_X1 U15982 ( .A1(n15595), .A2(n15970), .A3(n8569), .ZN(n15969) );
  INV_X1 U15983 ( .A(n15971), .ZN(n15970) );
  NAND2_X1 U15984 ( .A1(n15705), .A2(n15707), .ZN(n15971) );
  NOR2_X1 U15985 ( .A1(n15705), .A2(n15707), .ZN(n15968) );
  NAND2_X1 U15986 ( .A1(n15972), .A2(n15973), .ZN(n15707) );
  INV_X1 U15987 ( .A(n15974), .ZN(n15973) );
  NOR2_X1 U15988 ( .A1(n15975), .A2(n15716), .ZN(n15974) );
  NOR2_X1 U15989 ( .A1(n15714), .A2(n15715), .ZN(n15975) );
  NAND2_X1 U15990 ( .A1(n15715), .A2(n15714), .ZN(n15972) );
  XNOR2_X1 U15991 ( .A(n15976), .B(n15977), .ZN(n15714) );
  XOR2_X1 U15992 ( .A(n15978), .B(n15979), .Z(n15976) );
  NOR2_X1 U15993 ( .A1(n15980), .A2(n15981), .ZN(n15715) );
  INV_X1 U15994 ( .A(n15982), .ZN(n15981) );
  NAND2_X1 U15995 ( .A1(n15725), .A2(n15983), .ZN(n15982) );
  NAND2_X1 U15996 ( .A1(n15724), .A2(n15723), .ZN(n15983) );
  NOR2_X1 U15997 ( .A1(n8900), .A2(n15595), .ZN(n15725) );
  NOR2_X1 U15998 ( .A1(n15723), .A2(n15724), .ZN(n15980) );
  NOR2_X1 U15999 ( .A1(n15984), .A2(n15985), .ZN(n15724) );
  INV_X1 U16000 ( .A(n15986), .ZN(n15985) );
  NAND2_X1 U16001 ( .A1(n15733), .A2(n15987), .ZN(n15986) );
  NAND2_X1 U16002 ( .A1(n15732), .A2(n15731), .ZN(n15987) );
  NOR2_X1 U16003 ( .A1(n8439), .A2(n15595), .ZN(n15733) );
  NOR2_X1 U16004 ( .A1(n15731), .A2(n15732), .ZN(n15984) );
  NOR2_X1 U16005 ( .A1(n15988), .A2(n15989), .ZN(n15732) );
  INV_X1 U16006 ( .A(n15990), .ZN(n15989) );
  NAND2_X1 U16007 ( .A1(n15946), .A2(n15991), .ZN(n15990) );
  NAND2_X1 U16008 ( .A1(n15945), .A2(n15944), .ZN(n15991) );
  NOR2_X1 U16009 ( .A1(n8938), .A2(n15595), .ZN(n15946) );
  NOR2_X1 U16010 ( .A1(n15944), .A2(n15945), .ZN(n15988) );
  NOR2_X1 U16011 ( .A1(n15992), .A2(n15993), .ZN(n15945) );
  INV_X1 U16012 ( .A(n15994), .ZN(n15993) );
  NAND2_X1 U16013 ( .A1(n15745), .A2(n15995), .ZN(n15994) );
  NAND2_X1 U16014 ( .A1(n15744), .A2(n15743), .ZN(n15995) );
  NOR2_X1 U16015 ( .A1(n8430), .A2(n15595), .ZN(n15745) );
  NOR2_X1 U16016 ( .A1(n15743), .A2(n15744), .ZN(n15992) );
  NOR2_X1 U16017 ( .A1(n15996), .A2(n15997), .ZN(n15744) );
  INV_X1 U16018 ( .A(n15998), .ZN(n15997) );
  NAND2_X1 U16019 ( .A1(n15942), .A2(n15999), .ZN(n15998) );
  NAND2_X1 U16020 ( .A1(n15941), .A2(n15940), .ZN(n15999) );
  NOR2_X1 U16021 ( .A1(n8425), .A2(n15595), .ZN(n15942) );
  NOR2_X1 U16022 ( .A1(n15940), .A2(n15941), .ZN(n15996) );
  NOR2_X1 U16023 ( .A1(n16000), .A2(n16001), .ZN(n15941) );
  INV_X1 U16024 ( .A(n16002), .ZN(n16001) );
  NAND2_X1 U16025 ( .A1(n15757), .A2(n16003), .ZN(n16002) );
  NAND2_X1 U16026 ( .A1(n15756), .A2(n15755), .ZN(n16003) );
  NOR2_X1 U16027 ( .A1(n8968), .A2(n15595), .ZN(n15757) );
  NOR2_X1 U16028 ( .A1(n15755), .A2(n15756), .ZN(n16000) );
  NOR2_X1 U16029 ( .A1(n16004), .A2(n16005), .ZN(n15756) );
  INV_X1 U16030 ( .A(n16006), .ZN(n16005) );
  NAND2_X1 U16031 ( .A1(n15938), .A2(n16007), .ZN(n16006) );
  NAND2_X1 U16032 ( .A1(n15937), .A2(n15936), .ZN(n16007) );
  NOR2_X1 U16033 ( .A1(n8971), .A2(n15595), .ZN(n15938) );
  NOR2_X1 U16034 ( .A1(n15936), .A2(n15937), .ZN(n16004) );
  NOR2_X1 U16035 ( .A1(n16008), .A2(n16009), .ZN(n15937) );
  INV_X1 U16036 ( .A(n16010), .ZN(n16009) );
  NAND2_X1 U16037 ( .A1(n15770), .A2(n16011), .ZN(n16010) );
  NAND2_X1 U16038 ( .A1(n15769), .A2(n15768), .ZN(n16011) );
  NOR2_X1 U16039 ( .A1(n8402), .A2(n15595), .ZN(n15770) );
  NOR2_X1 U16040 ( .A1(n15768), .A2(n15769), .ZN(n16008) );
  NOR2_X1 U16041 ( .A1(n16012), .A2(n16013), .ZN(n15769) );
  INV_X1 U16042 ( .A(n16014), .ZN(n16013) );
  NAND2_X1 U16043 ( .A1(n15934), .A2(n16015), .ZN(n16014) );
  NAND2_X1 U16044 ( .A1(n15933), .A2(n15932), .ZN(n16015) );
  NOR2_X1 U16045 ( .A1(n8867), .A2(n15595), .ZN(n15934) );
  NOR2_X1 U16046 ( .A1(n15932), .A2(n15933), .ZN(n16012) );
  NOR2_X1 U16047 ( .A1(n16016), .A2(n16017), .ZN(n15933) );
  INV_X1 U16048 ( .A(n16018), .ZN(n16017) );
  NAND2_X1 U16049 ( .A1(n15782), .A2(n16019), .ZN(n16018) );
  NAND2_X1 U16050 ( .A1(n15781), .A2(n15780), .ZN(n16019) );
  NOR2_X1 U16051 ( .A1(n8393), .A2(n15595), .ZN(n15782) );
  NOR2_X1 U16052 ( .A1(n15780), .A2(n15781), .ZN(n16016) );
  NOR2_X1 U16053 ( .A1(n16020), .A2(n16021), .ZN(n15781) );
  INV_X1 U16054 ( .A(n16022), .ZN(n16021) );
  NAND2_X1 U16055 ( .A1(n15930), .A2(n16023), .ZN(n16022) );
  NAND2_X1 U16056 ( .A1(n15929), .A2(n15928), .ZN(n16023) );
  NOR2_X1 U16057 ( .A1(n8996), .A2(n15595), .ZN(n15930) );
  NOR2_X1 U16058 ( .A1(n15928), .A2(n15929), .ZN(n16020) );
  NOR2_X1 U16059 ( .A1(n16024), .A2(n16025), .ZN(n15929) );
  INV_X1 U16060 ( .A(n16026), .ZN(n16025) );
  NAND2_X1 U16061 ( .A1(n15794), .A2(n16027), .ZN(n16026) );
  NAND2_X1 U16062 ( .A1(n15793), .A2(n15792), .ZN(n16027) );
  NOR2_X1 U16063 ( .A1(n9262), .A2(n15595), .ZN(n15794) );
  NOR2_X1 U16064 ( .A1(n15792), .A2(n15793), .ZN(n16024) );
  NOR2_X1 U16065 ( .A1(n16028), .A2(n16029), .ZN(n15793) );
  INV_X1 U16066 ( .A(n16030), .ZN(n16029) );
  NAND2_X1 U16067 ( .A1(n15926), .A2(n16031), .ZN(n16030) );
  NAND2_X1 U16068 ( .A1(n15925), .A2(n15924), .ZN(n16031) );
  NOR2_X1 U16069 ( .A1(n8850), .A2(n15595), .ZN(n15926) );
  NOR2_X1 U16070 ( .A1(n15924), .A2(n15925), .ZN(n16028) );
  INV_X1 U16071 ( .A(n16032), .ZN(n15925) );
  NAND2_X1 U16072 ( .A1(n16033), .A2(n16034), .ZN(n16032) );
  NAND2_X1 U16073 ( .A1(n15806), .A2(n16035), .ZN(n16034) );
  INV_X1 U16074 ( .A(n16036), .ZN(n16035) );
  NOR2_X1 U16075 ( .A1(n15803), .A2(n15805), .ZN(n16036) );
  NOR2_X1 U16076 ( .A1(n8376), .A2(n15595), .ZN(n15806) );
  NAND2_X1 U16077 ( .A1(n15803), .A2(n15805), .ZN(n16033) );
  NAND2_X1 U16078 ( .A1(n16037), .A2(n16038), .ZN(n15805) );
  INV_X1 U16079 ( .A(n16039), .ZN(n16038) );
  NOR2_X1 U16080 ( .A1(n15922), .A2(n16040), .ZN(n16039) );
  NOR2_X1 U16081 ( .A1(n15921), .A2(n15919), .ZN(n16040) );
  NAND2_X1 U16082 ( .A1(a_17_), .A2(b_2_), .ZN(n15922) );
  NAND2_X1 U16083 ( .A1(n15919), .A2(n15921), .ZN(n16037) );
  NAND2_X1 U16084 ( .A1(n16041), .A2(n16042), .ZN(n15921) );
  NAND2_X1 U16085 ( .A1(n15818), .A2(n16043), .ZN(n16042) );
  INV_X1 U16086 ( .A(n16044), .ZN(n16043) );
  NOR2_X1 U16087 ( .A1(n15817), .A2(n15815), .ZN(n16044) );
  NOR2_X1 U16088 ( .A1(n9291), .A2(n15595), .ZN(n15818) );
  NAND2_X1 U16089 ( .A1(n15815), .A2(n15817), .ZN(n16041) );
  NAND2_X1 U16090 ( .A1(n16045), .A2(n16046), .ZN(n15817) );
  NAND2_X1 U16091 ( .A1(n15918), .A2(n16047), .ZN(n16046) );
  INV_X1 U16092 ( .A(n16048), .ZN(n16047) );
  NOR2_X1 U16093 ( .A1(n15917), .A2(n15916), .ZN(n16048) );
  NOR2_X1 U16094 ( .A1(n15595), .A2(n8742), .ZN(n15918) );
  NAND2_X1 U16095 ( .A1(n15916), .A2(n15917), .ZN(n16045) );
  NAND2_X1 U16096 ( .A1(n16049), .A2(n16050), .ZN(n15917) );
  NAND2_X1 U16097 ( .A1(n15830), .A2(n16051), .ZN(n16050) );
  INV_X1 U16098 ( .A(n16052), .ZN(n16051) );
  NOR2_X1 U16099 ( .A1(n15829), .A2(n15827), .ZN(n16052) );
  NOR2_X1 U16100 ( .A1(n15595), .A2(n9047), .ZN(n15830) );
  NAND2_X1 U16101 ( .A1(n15827), .A2(n15829), .ZN(n16049) );
  NAND2_X1 U16102 ( .A1(n16053), .A2(n16054), .ZN(n15829) );
  NAND2_X1 U16103 ( .A1(n15914), .A2(n16055), .ZN(n16054) );
  NAND2_X1 U16104 ( .A1(n15913), .A2(n15912), .ZN(n16055) );
  NOR2_X1 U16105 ( .A1(n15595), .A2(n8759), .ZN(n15914) );
  INV_X1 U16106 ( .A(n16056), .ZN(n16053) );
  NOR2_X1 U16107 ( .A1(n15912), .A2(n15913), .ZN(n16056) );
  NOR2_X1 U16108 ( .A1(n16057), .A2(n16058), .ZN(n15913) );
  NOR2_X1 U16109 ( .A1(n15842), .A2(n16059), .ZN(n16058) );
  NOR2_X1 U16110 ( .A1(n15841), .A2(n15839), .ZN(n16059) );
  NAND2_X1 U16111 ( .A1(b_2_), .A2(a_22_), .ZN(n15842) );
  INV_X1 U16112 ( .A(n16060), .ZN(n16057) );
  NAND2_X1 U16113 ( .A1(n15839), .A2(n15841), .ZN(n16060) );
  NAND2_X1 U16114 ( .A1(n16061), .A2(n16062), .ZN(n15841) );
  NAND2_X1 U16115 ( .A1(n15910), .A2(n16063), .ZN(n16062) );
  INV_X1 U16116 ( .A(n16064), .ZN(n16063) );
  NOR2_X1 U16117 ( .A1(n15909), .A2(n15907), .ZN(n16064) );
  NOR2_X1 U16118 ( .A1(n15595), .A2(n12301), .ZN(n15910) );
  NAND2_X1 U16119 ( .A1(n15907), .A2(n15909), .ZN(n16061) );
  NAND2_X1 U16120 ( .A1(n15852), .A2(n16065), .ZN(n15909) );
  NAND2_X1 U16121 ( .A1(n15851), .A2(n15853), .ZN(n16065) );
  NAND2_X1 U16122 ( .A1(n16066), .A2(n16067), .ZN(n15853) );
  NAND2_X1 U16123 ( .A1(b_2_), .A2(a_24_), .ZN(n16067) );
  INV_X1 U16124 ( .A(n16068), .ZN(n16066) );
  XOR2_X1 U16125 ( .A(n16069), .B(n16070), .Z(n15851) );
  XNOR2_X1 U16126 ( .A(n16071), .B(n16072), .ZN(n16070) );
  NAND2_X1 U16127 ( .A1(b_1_), .A2(a_25_), .ZN(n16069) );
  NAND2_X1 U16128 ( .A1(a_24_), .A2(n16068), .ZN(n15852) );
  NAND2_X1 U16129 ( .A1(n15905), .A2(n16073), .ZN(n16068) );
  NAND2_X1 U16130 ( .A1(n15904), .A2(n15906), .ZN(n16073) );
  NAND2_X1 U16131 ( .A1(n16074), .A2(n16075), .ZN(n15906) );
  NAND2_X1 U16132 ( .A1(b_2_), .A2(a_25_), .ZN(n16075) );
  XOR2_X1 U16133 ( .A(n16076), .B(n16077), .Z(n15904) );
  NOR2_X1 U16134 ( .A1(n9344), .A2(n15890), .ZN(n16077) );
  XOR2_X1 U16135 ( .A(n16078), .B(n16079), .Z(n16076) );
  NAND2_X1 U16136 ( .A1(a_25_), .A2(n16080), .ZN(n15905) );
  INV_X1 U16137 ( .A(n16074), .ZN(n16080) );
  NOR2_X1 U16138 ( .A1(n16081), .A2(n16082), .ZN(n16074) );
  NOR3_X1 U16139 ( .A1(n9344), .A2(n16083), .A3(n15595), .ZN(n16082) );
  NOR2_X1 U16140 ( .A1(n15865), .A2(n15863), .ZN(n16083) );
  INV_X1 U16141 ( .A(n16084), .ZN(n16081) );
  NAND2_X1 U16142 ( .A1(n15863), .A2(n15865), .ZN(n16084) );
  NAND2_X1 U16143 ( .A1(n15901), .A2(n16085), .ZN(n15865) );
  NAND2_X1 U16144 ( .A1(n15900), .A2(n15902), .ZN(n16085) );
  NAND2_X1 U16145 ( .A1(n16086), .A2(n16087), .ZN(n15902) );
  NAND2_X1 U16146 ( .A1(b_2_), .A2(a_27_), .ZN(n16087) );
  INV_X1 U16147 ( .A(n16088), .ZN(n16086) );
  XOR2_X1 U16148 ( .A(n16089), .B(n16090), .Z(n15900) );
  XNOR2_X1 U16149 ( .A(n16091), .B(n16092), .ZN(n16090) );
  NAND2_X1 U16150 ( .A1(b_1_), .A2(a_28_), .ZN(n16089) );
  NAND2_X1 U16151 ( .A1(a_27_), .A2(n16088), .ZN(n15901) );
  NAND2_X1 U16152 ( .A1(n16093), .A2(n16094), .ZN(n16088) );
  INV_X1 U16153 ( .A(n16095), .ZN(n16094) );
  NOR3_X1 U16154 ( .A1(n8314), .A2(n16096), .A3(n15595), .ZN(n16095) );
  NOR2_X1 U16155 ( .A1(n15896), .A2(n15898), .ZN(n16096) );
  NAND2_X1 U16156 ( .A1(n15896), .A2(n15898), .ZN(n16093) );
  NAND2_X1 U16157 ( .A1(n16097), .A2(n16098), .ZN(n15898) );
  NAND2_X1 U16158 ( .A1(n15892), .A2(n16099), .ZN(n16098) );
  INV_X1 U16159 ( .A(n16100), .ZN(n16099) );
  NOR2_X1 U16160 ( .A1(n15893), .A2(n15894), .ZN(n16100) );
  NOR2_X1 U16161 ( .A1(n15595), .A2(n9098), .ZN(n15892) );
  NAND2_X1 U16162 ( .A1(n15894), .A2(n15893), .ZN(n16097) );
  NAND2_X1 U16163 ( .A1(n16101), .A2(n16102), .ZN(n15893) );
  NAND2_X1 U16164 ( .A1(b_0_), .A2(n16103), .ZN(n16102) );
  NAND2_X1 U16165 ( .A1(n8299), .A2(n16104), .ZN(n16103) );
  NAND2_X1 U16166 ( .A1(a_31_), .A2(n15890), .ZN(n16104) );
  NAND2_X1 U16167 ( .A1(b_1_), .A2(n16106), .ZN(n16101) );
  NAND2_X1 U16168 ( .A1(n8303), .A2(n16107), .ZN(n16106) );
  NAND2_X1 U16169 ( .A1(a_30_), .A2(n8567), .ZN(n16107) );
  NOR3_X1 U16170 ( .A1(n15595), .A2(n9631), .A3(n15890), .ZN(n15894) );
  INV_X1 U16171 ( .A(n9106), .ZN(n9631) );
  XNOR2_X1 U16172 ( .A(n16109), .B(n16110), .ZN(n15896) );
  XNOR2_X1 U16173 ( .A(n16111), .B(n16112), .ZN(n16110) );
  NAND2_X1 U16174 ( .A1(b_0_), .A2(a_30_), .ZN(n16109) );
  XOR2_X1 U16175 ( .A(n16113), .B(n16114), .Z(n15863) );
  XNOR2_X1 U16176 ( .A(n16115), .B(n16116), .ZN(n16114) );
  NAND2_X1 U16177 ( .A1(b_1_), .A2(a_27_), .ZN(n16113) );
  XOR2_X1 U16178 ( .A(n16117), .B(n16118), .Z(n15907) );
  NOR2_X1 U16179 ( .A1(n8779), .A2(n15890), .ZN(n16118) );
  XOR2_X1 U16180 ( .A(n16119), .B(n16120), .Z(n16117) );
  XOR2_X1 U16181 ( .A(n16121), .B(n16122), .Z(n15839) );
  XNOR2_X1 U16182 ( .A(n16123), .B(n16124), .ZN(n16122) );
  NAND2_X1 U16183 ( .A1(b_1_), .A2(a_23_), .ZN(n16121) );
  XNOR2_X1 U16184 ( .A(n16125), .B(n16126), .ZN(n15912) );
  NOR2_X1 U16185 ( .A1(n12296), .A2(n15890), .ZN(n16126) );
  XNOR2_X1 U16186 ( .A(n16127), .B(n16128), .ZN(n16125) );
  XOR2_X1 U16187 ( .A(n16129), .B(n16130), .Z(n15827) );
  XNOR2_X1 U16188 ( .A(n16131), .B(n16132), .ZN(n16130) );
  NAND2_X1 U16189 ( .A1(b_1_), .A2(a_21_), .ZN(n16129) );
  XOR2_X1 U16190 ( .A(n16133), .B(n16134), .Z(n15916) );
  NOR2_X1 U16191 ( .A1(n9047), .A2(n15890), .ZN(n16134) );
  XOR2_X1 U16192 ( .A(n16135), .B(n16136), .Z(n16133) );
  XOR2_X1 U16193 ( .A(n16137), .B(n16138), .Z(n15815) );
  XNOR2_X1 U16194 ( .A(n16139), .B(n16140), .ZN(n16138) );
  NAND2_X1 U16195 ( .A1(b_1_), .A2(a_19_), .ZN(n16137) );
  XOR2_X1 U16196 ( .A(n16141), .B(n16142), .Z(n15919) );
  XNOR2_X1 U16197 ( .A(n16143), .B(n16144), .ZN(n16141) );
  XNOR2_X1 U16198 ( .A(n16145), .B(n16146), .ZN(n15803) );
  XNOR2_X1 U16199 ( .A(n16147), .B(n16148), .ZN(n16145) );
  XNOR2_X1 U16200 ( .A(n16149), .B(n16150), .ZN(n15924) );
  XNOR2_X1 U16201 ( .A(n16151), .B(n16152), .ZN(n16150) );
  XNOR2_X1 U16202 ( .A(n16153), .B(n16154), .ZN(n15792) );
  XOR2_X1 U16203 ( .A(n16155), .B(n16156), .Z(n16153) );
  XOR2_X1 U16204 ( .A(n16157), .B(n16158), .Z(n15928) );
  XNOR2_X1 U16205 ( .A(n16159), .B(n16160), .ZN(n16158) );
  XNOR2_X1 U16206 ( .A(n16161), .B(n16162), .ZN(n15780) );
  XOR2_X1 U16207 ( .A(n16163), .B(n16164), .Z(n16161) );
  XOR2_X1 U16208 ( .A(n16165), .B(n16166), .Z(n15932) );
  XNOR2_X1 U16209 ( .A(n16167), .B(n16168), .ZN(n16166) );
  XNOR2_X1 U16210 ( .A(n16169), .B(n16170), .ZN(n15768) );
  XOR2_X1 U16211 ( .A(n16171), .B(n16172), .Z(n16169) );
  XNOR2_X1 U16212 ( .A(n16173), .B(n16174), .ZN(n15936) );
  XOR2_X1 U16213 ( .A(n16175), .B(n16176), .Z(n16173) );
  XNOR2_X1 U16214 ( .A(n16177), .B(n16178), .ZN(n15755) );
  XOR2_X1 U16215 ( .A(n16179), .B(n16180), .Z(n16177) );
  XNOR2_X1 U16216 ( .A(n16181), .B(n16182), .ZN(n15940) );
  XOR2_X1 U16217 ( .A(n16183), .B(n16184), .Z(n16181) );
  XNOR2_X1 U16218 ( .A(n16185), .B(n16186), .ZN(n15743) );
  XOR2_X1 U16219 ( .A(n16187), .B(n16188), .Z(n16185) );
  XNOR2_X1 U16220 ( .A(n16189), .B(n16190), .ZN(n15944) );
  XOR2_X1 U16221 ( .A(n16191), .B(n16192), .Z(n16189) );
  XNOR2_X1 U16222 ( .A(n16193), .B(n16194), .ZN(n15731) );
  XOR2_X1 U16223 ( .A(n16195), .B(n16196), .Z(n16193) );
  XNOR2_X1 U16224 ( .A(n16197), .B(n16198), .ZN(n15723) );
  XOR2_X1 U16225 ( .A(n16199), .B(n16200), .Z(n16197) );
  XNOR2_X1 U16226 ( .A(n16201), .B(n15962), .ZN(n15705) );
  NOR2_X1 U16227 ( .A1(n8448), .A2(n15890), .ZN(n15962) );
  XOR2_X1 U16228 ( .A(n15965), .B(n15966), .Z(n16201) );
  NOR2_X1 U16229 ( .A1(n8900), .A2(n8567), .ZN(n15966) );
  NAND2_X1 U16230 ( .A1(n16202), .A2(n16203), .ZN(n15965) );
  NAND2_X1 U16231 ( .A1(n15977), .A2(n16204), .ZN(n16203) );
  INV_X1 U16232 ( .A(n16205), .ZN(n16204) );
  NOR2_X1 U16233 ( .A1(n15978), .A2(n15979), .ZN(n16205) );
  NOR2_X1 U16234 ( .A1(n8900), .A2(n15890), .ZN(n15977) );
  NAND2_X1 U16235 ( .A1(n15979), .A2(n15978), .ZN(n16202) );
  NAND2_X1 U16236 ( .A1(n16206), .A2(n16207), .ZN(n15978) );
  NAND2_X1 U16237 ( .A1(n16198), .A2(n16208), .ZN(n16207) );
  INV_X1 U16238 ( .A(n16209), .ZN(n16208) );
  NOR2_X1 U16239 ( .A1(n16199), .A2(n16200), .ZN(n16209) );
  NOR2_X1 U16240 ( .A1(n8439), .A2(n15890), .ZN(n16198) );
  NAND2_X1 U16241 ( .A1(n16200), .A2(n16199), .ZN(n16206) );
  NAND2_X1 U16242 ( .A1(n16210), .A2(n16211), .ZN(n16199) );
  NAND2_X1 U16243 ( .A1(n16194), .A2(n16212), .ZN(n16211) );
  INV_X1 U16244 ( .A(n16213), .ZN(n16212) );
  NOR2_X1 U16245 ( .A1(n16195), .A2(n16196), .ZN(n16213) );
  NOR2_X1 U16246 ( .A1(n8938), .A2(n15890), .ZN(n16194) );
  NAND2_X1 U16247 ( .A1(n16196), .A2(n16195), .ZN(n16210) );
  NAND2_X1 U16248 ( .A1(n16214), .A2(n16215), .ZN(n16195) );
  NAND2_X1 U16249 ( .A1(n16190), .A2(n16216), .ZN(n16215) );
  INV_X1 U16250 ( .A(n16217), .ZN(n16216) );
  NOR2_X1 U16251 ( .A1(n16191), .A2(n16192), .ZN(n16217) );
  NOR2_X1 U16252 ( .A1(n8430), .A2(n15890), .ZN(n16190) );
  NAND2_X1 U16253 ( .A1(n16192), .A2(n16191), .ZN(n16214) );
  NAND2_X1 U16254 ( .A1(n16218), .A2(n16219), .ZN(n16191) );
  NAND2_X1 U16255 ( .A1(n16186), .A2(n16220), .ZN(n16219) );
  INV_X1 U16256 ( .A(n16221), .ZN(n16220) );
  NOR2_X1 U16257 ( .A1(n16187), .A2(n16188), .ZN(n16221) );
  NOR2_X1 U16258 ( .A1(n8425), .A2(n15890), .ZN(n16186) );
  NAND2_X1 U16259 ( .A1(n16188), .A2(n16187), .ZN(n16218) );
  NAND2_X1 U16260 ( .A1(n16222), .A2(n16223), .ZN(n16187) );
  NAND2_X1 U16261 ( .A1(n16182), .A2(n16224), .ZN(n16223) );
  INV_X1 U16262 ( .A(n16225), .ZN(n16224) );
  NOR2_X1 U16263 ( .A1(n16183), .A2(n16184), .ZN(n16225) );
  NOR2_X1 U16264 ( .A1(n8968), .A2(n15890), .ZN(n16182) );
  NAND2_X1 U16265 ( .A1(n16184), .A2(n16183), .ZN(n16222) );
  NAND2_X1 U16266 ( .A1(n16226), .A2(n16227), .ZN(n16183) );
  NAND2_X1 U16267 ( .A1(n16178), .A2(n16228), .ZN(n16227) );
  INV_X1 U16268 ( .A(n16229), .ZN(n16228) );
  NOR2_X1 U16269 ( .A1(n16179), .A2(n16180), .ZN(n16229) );
  NOR2_X1 U16270 ( .A1(n8971), .A2(n15890), .ZN(n16178) );
  NAND2_X1 U16271 ( .A1(n16180), .A2(n16179), .ZN(n16226) );
  NAND2_X1 U16272 ( .A1(n16230), .A2(n16231), .ZN(n16179) );
  NAND2_X1 U16273 ( .A1(n16174), .A2(n16232), .ZN(n16231) );
  INV_X1 U16274 ( .A(n16233), .ZN(n16232) );
  NOR2_X1 U16275 ( .A1(n16175), .A2(n16176), .ZN(n16233) );
  NOR2_X1 U16276 ( .A1(n8402), .A2(n15890), .ZN(n16174) );
  NAND2_X1 U16277 ( .A1(n16176), .A2(n16175), .ZN(n16230) );
  NAND2_X1 U16278 ( .A1(n16234), .A2(n16235), .ZN(n16175) );
  NAND2_X1 U16279 ( .A1(n16170), .A2(n16236), .ZN(n16235) );
  INV_X1 U16280 ( .A(n16237), .ZN(n16236) );
  NOR2_X1 U16281 ( .A1(n16171), .A2(n16172), .ZN(n16237) );
  NOR2_X1 U16282 ( .A1(n8867), .A2(n15890), .ZN(n16170) );
  NAND2_X1 U16283 ( .A1(n16172), .A2(n16171), .ZN(n16234) );
  NAND2_X1 U16284 ( .A1(n16238), .A2(n16239), .ZN(n16171) );
  NAND2_X1 U16285 ( .A1(n16165), .A2(n16240), .ZN(n16239) );
  NAND2_X1 U16286 ( .A1(n16167), .A2(n16168), .ZN(n16240) );
  NOR2_X1 U16287 ( .A1(n8393), .A2(n15890), .ZN(n16165) );
  INV_X1 U16288 ( .A(n16241), .ZN(n16238) );
  NOR2_X1 U16289 ( .A1(n16168), .A2(n16167), .ZN(n16241) );
  NOR2_X1 U16290 ( .A1(n16242), .A2(n16243), .ZN(n16167) );
  INV_X1 U16291 ( .A(n16244), .ZN(n16243) );
  NAND2_X1 U16292 ( .A1(n16162), .A2(n16245), .ZN(n16244) );
  NAND2_X1 U16293 ( .A1(n16164), .A2(n16163), .ZN(n16245) );
  NOR2_X1 U16294 ( .A1(n8996), .A2(n15890), .ZN(n16162) );
  NOR2_X1 U16295 ( .A1(n16163), .A2(n16164), .ZN(n16242) );
  NOR2_X1 U16296 ( .A1(n16246), .A2(n16247), .ZN(n16164) );
  INV_X1 U16297 ( .A(n16248), .ZN(n16247) );
  NAND2_X1 U16298 ( .A1(n16157), .A2(n16249), .ZN(n16248) );
  NAND2_X1 U16299 ( .A1(n16159), .A2(n16160), .ZN(n16249) );
  NOR2_X1 U16300 ( .A1(n9262), .A2(n15890), .ZN(n16157) );
  NOR2_X1 U16301 ( .A1(n16160), .A2(n16159), .ZN(n16246) );
  NOR2_X1 U16302 ( .A1(n16250), .A2(n16251), .ZN(n16159) );
  INV_X1 U16303 ( .A(n16252), .ZN(n16251) );
  NAND2_X1 U16304 ( .A1(n16154), .A2(n16253), .ZN(n16252) );
  NAND2_X1 U16305 ( .A1(n16156), .A2(n16155), .ZN(n16253) );
  NOR2_X1 U16306 ( .A1(n8850), .A2(n15890), .ZN(n16154) );
  NOR2_X1 U16307 ( .A1(n16155), .A2(n16156), .ZN(n16250) );
  NOR2_X1 U16308 ( .A1(n16254), .A2(n16255), .ZN(n16156) );
  NOR2_X1 U16309 ( .A1(n16149), .A2(n16256), .ZN(n16255) );
  NOR2_X1 U16310 ( .A1(n16151), .A2(n16152), .ZN(n16256) );
  NAND2_X1 U16311 ( .A1(a_16_), .A2(b_1_), .ZN(n16149) );
  INV_X1 U16312 ( .A(n16257), .ZN(n16254) );
  NAND2_X1 U16313 ( .A1(n16152), .A2(n16151), .ZN(n16257) );
  NAND2_X1 U16314 ( .A1(n16258), .A2(n16259), .ZN(n16151) );
  NAND2_X1 U16315 ( .A1(n16146), .A2(n16260), .ZN(n16259) );
  INV_X1 U16316 ( .A(n16261), .ZN(n16260) );
  NOR2_X1 U16317 ( .A1(n16147), .A2(n16148), .ZN(n16261) );
  NOR2_X1 U16318 ( .A1(n8371), .A2(n15890), .ZN(n16146) );
  NAND2_X1 U16319 ( .A1(n16147), .A2(n16148), .ZN(n16258) );
  NOR2_X1 U16320 ( .A1(n9291), .A2(n8567), .ZN(n16148) );
  NOR2_X1 U16321 ( .A1(n16262), .A2(n16263), .ZN(n16147) );
  INV_X1 U16322 ( .A(n16264), .ZN(n16263) );
  NAND2_X1 U16323 ( .A1(n16265), .A2(n16143), .ZN(n16264) );
  NAND2_X1 U16324 ( .A1(b_0_), .A2(a_19_), .ZN(n16143) );
  NAND2_X1 U16325 ( .A1(n16142), .A2(n16144), .ZN(n16265) );
  NOR2_X1 U16326 ( .A1(n16144), .A2(n16142), .ZN(n16262) );
  NOR2_X1 U16327 ( .A1(n9291), .A2(n15890), .ZN(n16142) );
  NAND2_X1 U16328 ( .A1(n16266), .A2(n16267), .ZN(n16144) );
  INV_X1 U16329 ( .A(n16268), .ZN(n16267) );
  NOR3_X1 U16330 ( .A1(n8742), .A2(n16269), .A3(n15890), .ZN(n16268) );
  NOR2_X1 U16331 ( .A1(n16140), .A2(n16139), .ZN(n16269) );
  NAND2_X1 U16332 ( .A1(n16139), .A2(n16140), .ZN(n16266) );
  NAND2_X1 U16333 ( .A1(n16270), .A2(n16271), .ZN(n16140) );
  NAND3_X1 U16334 ( .A1(a_20_), .A2(n16272), .A3(b_1_), .ZN(n16271) );
  NAND2_X1 U16335 ( .A1(n16136), .A2(n16135), .ZN(n16272) );
  INV_X1 U16336 ( .A(n16273), .ZN(n16270) );
  NOR2_X1 U16337 ( .A1(n16135), .A2(n16136), .ZN(n16273) );
  NOR2_X1 U16338 ( .A1(n16274), .A2(n16275), .ZN(n16136) );
  NOR3_X1 U16339 ( .A1(n8759), .A2(n16276), .A3(n15890), .ZN(n16275) );
  NOR2_X1 U16340 ( .A1(n16132), .A2(n16131), .ZN(n16276) );
  INV_X1 U16341 ( .A(n16277), .ZN(n16274) );
  NAND2_X1 U16342 ( .A1(n16131), .A2(n16132), .ZN(n16277) );
  NAND2_X1 U16343 ( .A1(n16278), .A2(n16279), .ZN(n16132) );
  NAND3_X1 U16344 ( .A1(a_22_), .A2(n16280), .A3(b_1_), .ZN(n16279) );
  NAND2_X1 U16345 ( .A1(n16128), .A2(n16281), .ZN(n16280) );
  INV_X1 U16346 ( .A(n16282), .ZN(n16278) );
  NOR2_X1 U16347 ( .A1(n16281), .A2(n16128), .ZN(n16282) );
  NOR2_X1 U16348 ( .A1(n16283), .A2(n16284), .ZN(n16128) );
  NOR3_X1 U16349 ( .A1(n12301), .A2(n16285), .A3(n15890), .ZN(n16284) );
  NOR2_X1 U16350 ( .A1(n16124), .A2(n16123), .ZN(n16285) );
  INV_X1 U16351 ( .A(n16286), .ZN(n16283) );
  NAND2_X1 U16352 ( .A1(n16123), .A2(n16124), .ZN(n16286) );
  NAND2_X1 U16353 ( .A1(n16287), .A2(n16288), .ZN(n16124) );
  NAND3_X1 U16354 ( .A1(a_24_), .A2(n16289), .A3(b_1_), .ZN(n16288) );
  NAND2_X1 U16355 ( .A1(n16120), .A2(n16119), .ZN(n16289) );
  INV_X1 U16356 ( .A(n16290), .ZN(n16287) );
  NOR2_X1 U16357 ( .A1(n16119), .A2(n16120), .ZN(n16290) );
  NOR2_X1 U16358 ( .A1(n16291), .A2(n16292), .ZN(n16120) );
  NOR3_X1 U16359 ( .A1(n8788), .A2(n16293), .A3(n15890), .ZN(n16292) );
  NOR2_X1 U16360 ( .A1(n16072), .A2(n16071), .ZN(n16293) );
  INV_X1 U16361 ( .A(n16294), .ZN(n16291) );
  NAND2_X1 U16362 ( .A1(n16071), .A2(n16072), .ZN(n16294) );
  NAND2_X1 U16363 ( .A1(n16295), .A2(n16296), .ZN(n16072) );
  NAND3_X1 U16364 ( .A1(a_26_), .A2(n16297), .A3(b_1_), .ZN(n16296) );
  NAND2_X1 U16365 ( .A1(n16079), .A2(n16078), .ZN(n16297) );
  INV_X1 U16366 ( .A(n16298), .ZN(n16295) );
  NOR2_X1 U16367 ( .A1(n16078), .A2(n16079), .ZN(n16298) );
  NOR2_X1 U16368 ( .A1(n16299), .A2(n16300), .ZN(n16079) );
  NOR3_X1 U16369 ( .A1(n8797), .A2(n16301), .A3(n15890), .ZN(n16300) );
  NOR2_X1 U16370 ( .A1(n16116), .A2(n16115), .ZN(n16301) );
  INV_X1 U16371 ( .A(n16302), .ZN(n16299) );
  NAND2_X1 U16372 ( .A1(n16115), .A2(n16116), .ZN(n16302) );
  NAND2_X1 U16373 ( .A1(n16303), .A2(n16304), .ZN(n16116) );
  INV_X1 U16374 ( .A(n16305), .ZN(n16304) );
  NOR3_X1 U16375 ( .A1(n8314), .A2(n16306), .A3(n15890), .ZN(n16305) );
  NOR2_X1 U16376 ( .A1(n16092), .A2(n16091), .ZN(n16306) );
  NAND2_X1 U16377 ( .A1(n16091), .A2(n16092), .ZN(n16303) );
  NAND2_X1 U16378 ( .A1(n16112), .A2(n16307), .ZN(n16092) );
  NAND3_X1 U16379 ( .A1(b_0_), .A2(a_30_), .A3(n16111), .ZN(n16307) );
  NOR2_X1 U16380 ( .A1(n15890), .A2(n9098), .ZN(n16111) );
  NAND3_X1 U16381 ( .A1(b_1_), .A2(n9106), .A3(b_0_), .ZN(n16112) );
  NOR2_X1 U16382 ( .A1(n16108), .A2(n16105), .ZN(n9106) );
  NOR2_X1 U16383 ( .A1(n8567), .A2(n9098), .ZN(n16091) );
  NOR2_X1 U16384 ( .A1(n8567), .A2(n8314), .ZN(n16115) );
  NAND2_X1 U16385 ( .A1(b_0_), .A2(a_27_), .ZN(n16078) );
  NOR2_X1 U16386 ( .A1(n8567), .A2(n9344), .ZN(n16071) );
  NAND2_X1 U16387 ( .A1(b_0_), .A2(a_25_), .ZN(n16119) );
  NOR2_X1 U16388 ( .A1(n8567), .A2(n8779), .ZN(n16123) );
  INV_X1 U16389 ( .A(n16127), .ZN(n16281) );
  NOR2_X1 U16390 ( .A1(n8567), .A2(n12301), .ZN(n16127) );
  NOR2_X1 U16391 ( .A1(n8567), .A2(n12296), .ZN(n16131) );
  NAND2_X1 U16392 ( .A1(b_0_), .A2(a_21_), .ZN(n16135) );
  NOR2_X1 U16393 ( .A1(n8567), .A2(n9047), .ZN(n16139) );
  NOR2_X1 U16394 ( .A1(n8371), .A2(n8567), .ZN(n16152) );
  NAND2_X1 U16395 ( .A1(a_16_), .A2(b_0_), .ZN(n16155) );
  NAND2_X1 U16396 ( .A1(a_15_), .A2(b_0_), .ZN(n16160) );
  NAND2_X1 U16397 ( .A1(a_14_), .A2(b_0_), .ZN(n16163) );
  NAND2_X1 U16398 ( .A1(a_13_), .A2(b_0_), .ZN(n16168) );
  NOR2_X1 U16399 ( .A1(n8393), .A2(n8567), .ZN(n16172) );
  NOR2_X1 U16400 ( .A1(n8867), .A2(n8567), .ZN(n16176) );
  NOR2_X1 U16401 ( .A1(n8402), .A2(n8567), .ZN(n16180) );
  NOR2_X1 U16402 ( .A1(n8971), .A2(n8567), .ZN(n16184) );
  NOR2_X1 U16403 ( .A1(n8968), .A2(n8567), .ZN(n16188) );
  NOR2_X1 U16404 ( .A1(n8425), .A2(n8567), .ZN(n16192) );
  NOR2_X1 U16405 ( .A1(n8430), .A2(n8567), .ZN(n16196) );
  NOR2_X1 U16406 ( .A1(n8938), .A2(n8567), .ZN(n16200) );
  NOR2_X1 U16407 ( .A1(n8439), .A2(n8567), .ZN(n15979) );
  NAND3_X1 U16408 ( .A1(n16308), .A2(n16309), .A3(n16310), .ZN(Result_add_9_)
         );
  NAND2_X1 U16409 ( .A1(n13999), .A2(n16311), .ZN(n16310) );
  NAND3_X1 U16410 ( .A1(n16312), .A2(n8971), .A3(b_9_), .ZN(n16309) );
  NAND2_X1 U16411 ( .A1(n16313), .A2(n13840), .ZN(n16308) );
  XNOR2_X1 U16412 ( .A(n16312), .B(a_9_), .ZN(n16313) );
  XNOR2_X1 U16413 ( .A(n16314), .B(n16315), .ZN(Result_add_8_) );
  NAND2_X1 U16414 ( .A1(n16316), .A2(n14417), .ZN(n16315) );
  NAND3_X1 U16415 ( .A1(n16317), .A2(n16318), .A3(n16319), .ZN(Result_add_7_)
         );
  NAND2_X1 U16416 ( .A1(n14677), .A2(n16320), .ZN(n16319) );
  INV_X1 U16417 ( .A(n14743), .ZN(n14677) );
  NAND3_X1 U16418 ( .A1(n16321), .A2(n8425), .A3(b_7_), .ZN(n16318) );
  INV_X1 U16419 ( .A(n16320), .ZN(n16321) );
  NAND2_X1 U16420 ( .A1(n16322), .A2(n14345), .ZN(n16317) );
  XNOR2_X1 U16421 ( .A(n16320), .B(n8425), .ZN(n16322) );
  XNOR2_X1 U16422 ( .A(n16323), .B(n16324), .ZN(Result_add_6_) );
  NAND2_X1 U16423 ( .A1(n16325), .A2(n14927), .ZN(n16324) );
  NAND3_X1 U16424 ( .A1(n16326), .A2(n16327), .A3(n16328), .ZN(Result_add_5_)
         );
  NAND2_X1 U16425 ( .A1(n16329), .A2(n16330), .ZN(n16328) );
  INV_X1 U16426 ( .A(n16331), .ZN(n16327) );
  NOR3_X1 U16427 ( .A1(n16330), .A2(a_5_), .A3(n14859), .ZN(n16331) );
  NAND2_X1 U16428 ( .A1(n16332), .A2(n14859), .ZN(n16326) );
  XNOR2_X1 U16429 ( .A(n16330), .B(n8938), .ZN(n16332) );
  XNOR2_X1 U16430 ( .A(n16333), .B(n16334), .ZN(Result_add_4_) );
  NAND2_X1 U16431 ( .A1(n16335), .A2(n15434), .ZN(n16334) );
  NAND3_X1 U16432 ( .A1(n16336), .A2(n16337), .A3(n16338), .ZN(Result_add_3_)
         );
  NAND2_X1 U16433 ( .A1(n15695), .A2(n16339), .ZN(n16338) );
  INV_X1 U16434 ( .A(n16340), .ZN(n16337) );
  NOR3_X1 U16435 ( .A1(n16339), .A2(a_3_), .A3(n15343), .ZN(n16340) );
  NAND2_X1 U16436 ( .A1(n16341), .A2(n15343), .ZN(n16336) );
  XNOR2_X1 U16437 ( .A(n16339), .B(n8900), .ZN(n16341) );
  XNOR2_X1 U16438 ( .A(n8301), .B(a_31_), .ZN(Result_add_31_) );
  NAND3_X1 U16439 ( .A1(n16342), .A2(n16343), .A3(n16344), .ZN(Result_add_30_)
         );
  INV_X1 U16440 ( .A(n8306), .ZN(n16344) );
  NOR3_X1 U16441 ( .A1(n8305), .A2(n16105), .A3(n16345), .ZN(n8306) );
  NAND2_X1 U16442 ( .A1(n16346), .A2(n8305), .ZN(n16343) );
  INV_X1 U16443 ( .A(b_30_), .ZN(n8305) );
  XNOR2_X1 U16444 ( .A(a_30_), .B(n16345), .ZN(n16346) );
  NAND3_X1 U16445 ( .A1(n16345), .A2(n16105), .A3(b_30_), .ZN(n16342) );
  XNOR2_X1 U16446 ( .A(n16347), .B(n16348), .ZN(Result_add_2_) );
  NOR2_X1 U16447 ( .A1(n16349), .A2(n15716), .ZN(n16348) );
  NAND3_X1 U16448 ( .A1(n16350), .A2(n16351), .A3(n16352), .ZN(Result_add_29_)
         );
  NAND2_X1 U16449 ( .A1(n9108), .A2(n16353), .ZN(n16352) );
  NAND3_X1 U16450 ( .A1(n16354), .A2(n9098), .A3(b_29_), .ZN(n16351) );
  NAND2_X1 U16451 ( .A1(n16355), .A2(n8817), .ZN(n16350) );
  XNOR2_X1 U16452 ( .A(n16353), .B(n9098), .ZN(n16355) );
  XNOR2_X1 U16453 ( .A(n16356), .B(n16357), .ZN(Result_add_28_) );
  NOR2_X1 U16454 ( .A1(n16358), .A2(n9370), .ZN(n16357) );
  NAND3_X1 U16455 ( .A1(n16359), .A2(n16360), .A3(n16361), .ZN(Result_add_27_)
         );
  NAND2_X1 U16456 ( .A1(n9844), .A2(n16362), .ZN(n16361) );
  NAND3_X1 U16457 ( .A1(n16363), .A2(n8797), .A3(b_27_), .ZN(n16360) );
  NAND2_X1 U16458 ( .A1(n16364), .A2(n9367), .ZN(n16359) );
  XNOR2_X1 U16459 ( .A(n16363), .B(a_27_), .ZN(n16364) );
  XNOR2_X1 U16460 ( .A(n16365), .B(n16366), .ZN(Result_add_26_) );
  NAND2_X1 U16461 ( .A1(n16367), .A2(n9831), .ZN(n16366) );
  NAND3_X1 U16462 ( .A1(n16368), .A2(n16369), .A3(n16370), .ZN(Result_add_25_)
         );
  NAND2_X1 U16463 ( .A1(n10326), .A2(n16371), .ZN(n16370) );
  INV_X1 U16464 ( .A(n16372), .ZN(n16369) );
  NOR3_X1 U16465 ( .A1(n16371), .A2(a_25_), .A3(n9864), .ZN(n16372) );
  NAND2_X1 U16466 ( .A1(n16373), .A2(n9864), .ZN(n16368) );
  XNOR2_X1 U16467 ( .A(n16371), .B(n8788), .ZN(n16373) );
  XNOR2_X1 U16468 ( .A(n16374), .B(n16375), .ZN(Result_add_24_) );
  NAND2_X1 U16469 ( .A1(n16376), .A2(n10313), .ZN(n16375) );
  NAND3_X1 U16470 ( .A1(n16377), .A2(n16378), .A3(n16379), .ZN(Result_add_23_)
         );
  NAND2_X1 U16471 ( .A1(n10573), .A2(n16380), .ZN(n16379) );
  NAND3_X1 U16472 ( .A1(n16381), .A2(n12301), .A3(b_23_), .ZN(n16378) );
  NAND2_X1 U16473 ( .A1(n16382), .A2(n10358), .ZN(n16377) );
  XNOR2_X1 U16474 ( .A(n16380), .B(n12301), .ZN(n16382) );
  XNOR2_X1 U16475 ( .A(n16383), .B(n16384), .ZN(Result_add_22_) );
  NOR2_X1 U16476 ( .A1(n16385), .A2(n10892), .ZN(n16384) );
  NAND3_X1 U16477 ( .A1(n16386), .A2(n16387), .A3(n16388), .ZN(Result_add_21_)
         );
  NAND2_X1 U16478 ( .A1(n11059), .A2(n16389), .ZN(n16388) );
  INV_X1 U16479 ( .A(n16390), .ZN(n16389) );
  NAND3_X1 U16480 ( .A1(n16390), .A2(n8759), .A3(b_21_), .ZN(n16387) );
  NAND2_X1 U16481 ( .A1(n16391), .A2(n10876), .ZN(n16386) );
  XNOR2_X1 U16482 ( .A(n16390), .B(a_21_), .ZN(n16391) );
  XNOR2_X1 U16483 ( .A(n16392), .B(n16393), .ZN(Result_add_20_) );
  NOR2_X1 U16484 ( .A1(n16394), .A2(n11372), .ZN(n16393) );
  NAND2_X1 U16485 ( .A1(n16395), .A2(n16396), .ZN(Result_add_1_) );
  NAND2_X1 U16486 ( .A1(n16397), .A2(n16398), .ZN(n16396) );
  INV_X1 U16487 ( .A(n16399), .ZN(n16397) );
  NOR2_X1 U16488 ( .A1(n15955), .A2(n16400), .ZN(n16399) );
  NAND2_X1 U16489 ( .A1(n16401), .A2(n16402), .ZN(n16395) );
  XNOR2_X1 U16490 ( .A(n15890), .B(a_1_), .ZN(n16401) );
  NAND3_X1 U16491 ( .A1(n16403), .A2(n16404), .A3(n16405), .ZN(Result_add_19_)
         );
  INV_X1 U16492 ( .A(n16406), .ZN(n16405) );
  NOR2_X1 U16493 ( .A1(n11556), .A2(n16407), .ZN(n16406) );
  INV_X1 U16494 ( .A(n11787), .ZN(n11556) );
  NAND3_X1 U16495 ( .A1(n16407), .A2(n8742), .A3(b_19_), .ZN(n16404) );
  NAND2_X1 U16496 ( .A1(n16408), .A2(n11356), .ZN(n16403) );
  XNOR2_X1 U16497 ( .A(n16407), .B(a_19_), .ZN(n16408) );
  XNOR2_X1 U16498 ( .A(n16409), .B(n16410), .ZN(Result_add_18_) );
  NOR2_X1 U16499 ( .A1(n16411), .A2(n11879), .ZN(n16410) );
  NAND3_X1 U16500 ( .A1(n16412), .A2(n16413), .A3(n16414), .ZN(Result_add_17_)
         );
  INV_X1 U16501 ( .A(n16415), .ZN(n16414) );
  NOR2_X1 U16502 ( .A1(n12142), .A2(n16416), .ZN(n16415) );
  NAND3_X1 U16503 ( .A1(n16416), .A2(n8371), .A3(b_17_), .ZN(n16413) );
  NAND2_X1 U16504 ( .A1(n16417), .A2(n11859), .ZN(n16412) );
  XNOR2_X1 U16505 ( .A(n16416), .B(a_17_), .ZN(n16417) );
  XNOR2_X1 U16506 ( .A(n16418), .B(n16419), .ZN(Result_add_16_) );
  NAND2_X1 U16507 ( .A1(n16420), .A2(n12372), .ZN(n16419) );
  NAND3_X1 U16508 ( .A1(n16421), .A2(n16422), .A3(n16423), .ZN(Result_add_15_)
         );
  NAND2_X1 U16509 ( .A1(n12649), .A2(n16424), .ZN(n16423) );
  INV_X1 U16510 ( .A(n16425), .ZN(n16422) );
  NOR3_X1 U16511 ( .A1(n16424), .A2(a_15_), .A3(n12340), .ZN(n16425) );
  NAND2_X1 U16512 ( .A1(n16426), .A2(n12340), .ZN(n16421) );
  XNOR2_X1 U16513 ( .A(n16424), .B(n8850), .ZN(n16426) );
  XNOR2_X1 U16514 ( .A(n16427), .B(n16428), .ZN(Result_add_14_) );
  NAND2_X1 U16515 ( .A1(n16429), .A2(n12882), .ZN(n16428) );
  NAND3_X1 U16516 ( .A1(n16430), .A2(n16431), .A3(n16432), .ZN(Result_add_13_)
         );
  NAND2_X1 U16517 ( .A1(n13030), .A2(n16433), .ZN(n16432) );
  INV_X1 U16518 ( .A(n16434), .ZN(n16431) );
  NOR3_X1 U16519 ( .A1(n16433), .A2(a_13_), .A3(n12835), .ZN(n16434) );
  NAND2_X1 U16520 ( .A1(n16435), .A2(n12835), .ZN(n16430) );
  XNOR2_X1 U16521 ( .A(n16433), .B(n8996), .ZN(n16435) );
  XNOR2_X1 U16522 ( .A(n16436), .B(n16437), .ZN(Result_add_12_) );
  NAND2_X1 U16523 ( .A1(n16438), .A2(n13387), .ZN(n16437) );
  NAND3_X1 U16524 ( .A1(n16439), .A2(n16440), .A3(n16441), .ZN(Result_add_11_)
         );
  NAND2_X1 U16525 ( .A1(n13525), .A2(n16442), .ZN(n16441) );
  NAND3_X1 U16526 ( .A1(n16443), .A2(n8867), .A3(b_11_), .ZN(n16440) );
  NAND2_X1 U16527 ( .A1(n16444), .A2(n13332), .ZN(n16439) );
  XNOR2_X1 U16528 ( .A(n16442), .B(n8867), .ZN(n16444) );
  XNOR2_X1 U16529 ( .A(n16445), .B(n16446), .ZN(Result_add_10_) );
  NOR2_X1 U16530 ( .A1(n16447), .A2(n13902), .ZN(n16446) );
  XOR2_X1 U16531 ( .A(n16448), .B(n16449), .Z(Result_add_0_) );
  NOR2_X1 U16532 ( .A1(n16450), .A2(n8560), .ZN(n16449) );
  NOR2_X1 U16533 ( .A1(n8457), .A2(n8567), .ZN(n8560) );
  INV_X1 U16534 ( .A(b_0_), .ZN(n8567) );
  INV_X1 U16535 ( .A(a_0_), .ZN(n8457) );
  NOR2_X1 U16536 ( .A1(b_0_), .A2(a_0_), .ZN(n16450) );
  NOR2_X1 U16537 ( .A1(n16400), .A2(n16451), .ZN(n16448) );
  NOR2_X1 U16538 ( .A1(n15955), .A2(n16398), .ZN(n16451) );
  INV_X1 U16539 ( .A(n16402), .ZN(n16398) );
  NOR2_X1 U16540 ( .A1(n15716), .A2(n16452), .ZN(n16402) );
  NOR2_X1 U16541 ( .A1(n16349), .A2(n16347), .ZN(n16452) );
  NOR2_X1 U16542 ( .A1(n15695), .A2(n16453), .ZN(n16347) );
  INV_X1 U16543 ( .A(n16454), .ZN(n16453) );
  NAND2_X1 U16544 ( .A1(n16455), .A2(n16339), .ZN(n16454) );
  NAND2_X1 U16545 ( .A1(n15434), .A2(n16456), .ZN(n16339) );
  NAND2_X1 U16546 ( .A1(n16335), .A2(n16333), .ZN(n16456) );
  NAND2_X1 U16547 ( .A1(n15185), .A2(n16457), .ZN(n16333) );
  NAND2_X1 U16548 ( .A1(n16458), .A2(n16330), .ZN(n16457) );
  NAND2_X1 U16549 ( .A1(n14927), .A2(n16459), .ZN(n16330) );
  NAND2_X1 U16550 ( .A1(n16325), .A2(n16323), .ZN(n16459) );
  NAND2_X1 U16551 ( .A1(n14743), .A2(n16460), .ZN(n16323) );
  NAND2_X1 U16552 ( .A1(n16461), .A2(n16320), .ZN(n16460) );
  NAND2_X1 U16553 ( .A1(n14417), .A2(n16462), .ZN(n16320) );
  NAND2_X1 U16554 ( .A1(n16316), .A2(n16314), .ZN(n16462) );
  NAND2_X1 U16555 ( .A1(n14250), .A2(n16463), .ZN(n16314) );
  NAND2_X1 U16556 ( .A1(n16464), .A2(n16311), .ZN(n16463) );
  INV_X1 U16557 ( .A(n16312), .ZN(n16311) );
  NOR2_X1 U16558 ( .A1(n13902), .A2(n16465), .ZN(n16312) );
  NOR2_X1 U16559 ( .A1(n16447), .A2(n16445), .ZN(n16465) );
  NOR2_X1 U16560 ( .A1(n13525), .A2(n16466), .ZN(n16445) );
  NOR2_X1 U16561 ( .A1(n16467), .A2(n16443), .ZN(n16466) );
  INV_X1 U16562 ( .A(n16442), .ZN(n16443) );
  NAND2_X1 U16563 ( .A1(n13387), .A2(n16468), .ZN(n16442) );
  NAND2_X1 U16564 ( .A1(n16438), .A2(n16436), .ZN(n16468) );
  NAND2_X1 U16565 ( .A1(n13252), .A2(n16469), .ZN(n16436) );
  NAND2_X1 U16566 ( .A1(n16470), .A2(n16433), .ZN(n16469) );
  NAND2_X1 U16567 ( .A1(n12882), .A2(n16471), .ZN(n16433) );
  NAND2_X1 U16568 ( .A1(n16429), .A2(n16427), .ZN(n16471) );
  NAND2_X1 U16569 ( .A1(n12764), .A2(n16472), .ZN(n16427) );
  NAND2_X1 U16570 ( .A1(n16473), .A2(n16424), .ZN(n16472) );
  NAND2_X1 U16571 ( .A1(n12372), .A2(n16474), .ZN(n16424) );
  NAND2_X1 U16572 ( .A1(n16420), .A2(n16418), .ZN(n16474) );
  NAND2_X1 U16573 ( .A1(n12142), .A2(n16475), .ZN(n16418) );
  NAND2_X1 U16574 ( .A1(n16476), .A2(n16477), .ZN(n16475) );
  INV_X1 U16575 ( .A(n16416), .ZN(n16477) );
  NOR2_X1 U16576 ( .A1(n11879), .A2(n16478), .ZN(n16416) );
  NOR2_X1 U16577 ( .A1(n16411), .A2(n16409), .ZN(n16478) );
  NOR2_X1 U16578 ( .A1(n11787), .A2(n16479), .ZN(n16409) );
  NOR2_X1 U16579 ( .A1(n16480), .A2(n16407), .ZN(n16479) );
  NOR2_X1 U16580 ( .A1(n11372), .A2(n16481), .ZN(n16407) );
  NOR2_X1 U16581 ( .A1(n16394), .A2(n16392), .ZN(n16481) );
  NOR2_X1 U16582 ( .A1(n11059), .A2(n16482), .ZN(n16392) );
  NOR2_X1 U16583 ( .A1(n16483), .A2(n16390), .ZN(n16482) );
  NOR2_X1 U16584 ( .A1(n10892), .A2(n16484), .ZN(n16390) );
  NOR2_X1 U16585 ( .A1(n16385), .A2(n16383), .ZN(n16484) );
  NOR2_X1 U16586 ( .A1(n10573), .A2(n16485), .ZN(n16383) );
  NOR2_X1 U16587 ( .A1(n16486), .A2(n16381), .ZN(n16485) );
  INV_X1 U16588 ( .A(n16380), .ZN(n16381) );
  NAND2_X1 U16589 ( .A1(n10313), .A2(n16487), .ZN(n16380) );
  NAND2_X1 U16590 ( .A1(n16376), .A2(n16374), .ZN(n16487) );
  NAND2_X1 U16591 ( .A1(n10132), .A2(n16488), .ZN(n16374) );
  NAND2_X1 U16592 ( .A1(n16489), .A2(n16371), .ZN(n16488) );
  NAND2_X1 U16593 ( .A1(n9831), .A2(n16490), .ZN(n16371) );
  NAND2_X1 U16594 ( .A1(n16367), .A2(n16365), .ZN(n16490) );
  NAND2_X1 U16595 ( .A1(n9603), .A2(n16491), .ZN(n16365) );
  NAND2_X1 U16596 ( .A1(n16492), .A2(n16362), .ZN(n16491) );
  INV_X1 U16597 ( .A(n16363), .ZN(n16362) );
  NOR2_X1 U16598 ( .A1(n9370), .A2(n16493), .ZN(n16363) );
  NOR2_X1 U16599 ( .A1(n16358), .A2(n16356), .ZN(n16493) );
  NOR2_X1 U16600 ( .A1(n9108), .A2(n16494), .ZN(n16356) );
  NOR2_X1 U16601 ( .A1(n16495), .A2(n16354), .ZN(n16494) );
  INV_X1 U16602 ( .A(n16353), .ZN(n16354) );
  NAND2_X1 U16603 ( .A1(n16496), .A2(n16497), .ZN(n16353) );
  NAND2_X1 U16604 ( .A1(b_30_), .A2(n16498), .ZN(n16497) );
  NAND2_X1 U16605 ( .A1(n16105), .A2(n16345), .ZN(n16498) );
  INV_X1 U16606 ( .A(Result_mul_63_), .ZN(n16345) );
  INV_X1 U16607 ( .A(a_30_), .ZN(n16105) );
  NAND2_X1 U16608 ( .A1(Result_mul_63_), .A2(a_30_), .ZN(n16496) );
  NOR2_X1 U16609 ( .A1(n8301), .A2(n16108), .ZN(Result_mul_63_) );
  INV_X1 U16610 ( .A(a_31_), .ZN(n16108) );
  INV_X1 U16611 ( .A(b_31_), .ZN(n8301) );
  NOR2_X1 U16612 ( .A1(b_29_), .A2(a_29_), .ZN(n16495) );
  NOR2_X1 U16613 ( .A1(n8817), .A2(n9098), .ZN(n9108) );
  INV_X1 U16614 ( .A(b_29_), .ZN(n8817) );
  NOR2_X1 U16615 ( .A1(b_28_), .A2(a_28_), .ZN(n16358) );
  NOR2_X1 U16616 ( .A1(n9105), .A2(n8314), .ZN(n9370) );
  NAND2_X1 U16617 ( .A1(n9367), .A2(n8797), .ZN(n16492) );
  INV_X1 U16618 ( .A(n9844), .ZN(n9603) );
  NOR2_X1 U16619 ( .A1(n9367), .A2(n8797), .ZN(n9844) );
  INV_X1 U16620 ( .A(b_27_), .ZN(n9367) );
  NAND2_X1 U16621 ( .A1(n9630), .A2(n9344), .ZN(n16367) );
  INV_X1 U16622 ( .A(b_26_), .ZN(n9630) );
  NAND2_X1 U16623 ( .A1(b_26_), .A2(a_26_), .ZN(n9831) );
  NAND2_X1 U16624 ( .A1(n9864), .A2(n8788), .ZN(n16489) );
  INV_X1 U16625 ( .A(n10326), .ZN(n10132) );
  NOR2_X1 U16626 ( .A1(n9864), .A2(n8788), .ZN(n10326) );
  NAND2_X1 U16627 ( .A1(n10120), .A2(n8779), .ZN(n16376) );
  NAND2_X1 U16628 ( .A1(b_24_), .A2(a_24_), .ZN(n10313) );
  NOR2_X1 U16629 ( .A1(b_23_), .A2(a_23_), .ZN(n16486) );
  NOR2_X1 U16630 ( .A1(n10358), .A2(n12301), .ZN(n10573) );
  INV_X1 U16631 ( .A(a_23_), .ZN(n12301) );
  INV_X1 U16632 ( .A(b_23_), .ZN(n10358) );
  NOR2_X1 U16633 ( .A1(b_22_), .A2(a_22_), .ZN(n16385) );
  NOR2_X1 U16634 ( .A1(n10624), .A2(n12296), .ZN(n10892) );
  INV_X1 U16635 ( .A(a_22_), .ZN(n12296) );
  INV_X1 U16636 ( .A(b_22_), .ZN(n10624) );
  NOR2_X1 U16637 ( .A1(b_21_), .A2(a_21_), .ZN(n16483) );
  NOR2_X1 U16638 ( .A1(n10876), .A2(n8759), .ZN(n11059) );
  NOR2_X1 U16639 ( .A1(b_20_), .A2(a_20_), .ZN(n16394) );
  NOR2_X1 U16640 ( .A1(n11119), .A2(n9047), .ZN(n11372) );
  INV_X1 U16641 ( .A(b_20_), .ZN(n11119) );
  NOR2_X1 U16642 ( .A1(b_19_), .A2(a_19_), .ZN(n16480) );
  NOR2_X1 U16643 ( .A1(n11356), .A2(n8742), .ZN(n11787) );
  INV_X1 U16644 ( .A(a_19_), .ZN(n8742) );
  NOR2_X1 U16645 ( .A1(b_18_), .A2(a_18_), .ZN(n16411) );
  NOR2_X1 U16646 ( .A1(n11623), .A2(n9291), .ZN(n11879) );
  NAND2_X1 U16647 ( .A1(n11859), .A2(n8371), .ZN(n16476) );
  NAND2_X1 U16648 ( .A1(b_17_), .A2(a_17_), .ZN(n12142) );
  NAND2_X1 U16649 ( .A1(n12110), .A2(n8376), .ZN(n16420) );
  INV_X1 U16650 ( .A(a_16_), .ZN(n8376) );
  NAND2_X1 U16651 ( .A1(b_16_), .A2(a_16_), .ZN(n12372) );
  NAND2_X1 U16652 ( .A1(n12340), .A2(n8850), .ZN(n16473) );
  INV_X1 U16653 ( .A(n12649), .ZN(n12764) );
  NOR2_X1 U16654 ( .A1(n12340), .A2(n8850), .ZN(n12649) );
  NAND2_X1 U16655 ( .A1(n12609), .A2(n9262), .ZN(n16429) );
  INV_X1 U16656 ( .A(a_14_), .ZN(n9262) );
  NAND2_X1 U16657 ( .A1(b_14_), .A2(a_14_), .ZN(n12882) );
  NAND2_X1 U16658 ( .A1(n12835), .A2(n8996), .ZN(n16470) );
  INV_X1 U16659 ( .A(n13030), .ZN(n13252) );
  NOR2_X1 U16660 ( .A1(n12835), .A2(n8996), .ZN(n13030) );
  NAND2_X1 U16661 ( .A1(n13118), .A2(n8393), .ZN(n16438) );
  INV_X1 U16662 ( .A(b_12_), .ZN(n13118) );
  NAND2_X1 U16663 ( .A1(b_12_), .A2(a_12_), .ZN(n13387) );
  NOR2_X1 U16664 ( .A1(b_11_), .A2(a_11_), .ZN(n16467) );
  NOR2_X1 U16665 ( .A1(n8867), .A2(n13332), .ZN(n13525) );
  NOR2_X1 U16666 ( .A1(b_10_), .A2(a_10_), .ZN(n16447) );
  NOR2_X1 U16667 ( .A1(n8402), .A2(n13629), .ZN(n13902) );
  NAND2_X1 U16668 ( .A1(n13840), .A2(n8971), .ZN(n16464) );
  INV_X1 U16669 ( .A(n13999), .ZN(n14250) );
  NOR2_X1 U16670 ( .A1(n8971), .A2(n13840), .ZN(n13999) );
  NAND2_X1 U16671 ( .A1(n14123), .A2(n8968), .ZN(n16316) );
  INV_X1 U16672 ( .A(a_8_), .ZN(n8968) );
  NAND2_X1 U16673 ( .A1(a_8_), .A2(b_8_), .ZN(n14417) );
  NAND2_X1 U16674 ( .A1(n14345), .A2(n8425), .ZN(n16461) );
  NAND2_X1 U16675 ( .A1(a_7_), .A2(b_7_), .ZN(n14743) );
  NAND2_X1 U16676 ( .A1(n14621), .A2(n8430), .ZN(n16325) );
  INV_X1 U16677 ( .A(a_6_), .ZN(n8430) );
  NAND2_X1 U16678 ( .A1(a_6_), .A2(b_6_), .ZN(n14927) );
  NAND2_X1 U16679 ( .A1(n14859), .A2(n8938), .ZN(n16458) );
  INV_X1 U16680 ( .A(n16329), .ZN(n15185) );
  NOR2_X1 U16681 ( .A1(n8938), .A2(n14859), .ZN(n16329) );
  NAND2_X1 U16682 ( .A1(n15110), .A2(n8439), .ZN(n16335) );
  NAND2_X1 U16683 ( .A1(a_4_), .A2(b_4_), .ZN(n15434) );
  NAND2_X1 U16684 ( .A1(n15343), .A2(n8900), .ZN(n16455) );
  NOR2_X1 U16685 ( .A1(n8900), .A2(n15343), .ZN(n15695) );
  NOR2_X1 U16686 ( .A1(b_2_), .A2(a_2_), .ZN(n16349) );
  NOR2_X1 U16687 ( .A1(n8448), .A2(n15595), .ZN(n15716) );
  NOR2_X1 U16688 ( .A1(n8569), .A2(n15890), .ZN(n15955) );
  NOR2_X1 U16689 ( .A1(b_1_), .A2(a_1_), .ZN(n16400) );
endmodule

