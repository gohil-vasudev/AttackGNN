module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n670_, new_n456_, new_n170_, new_n246_, new_n266_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n655_, new_n117_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n112_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n651_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n120_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n108_, keyIn_0_14 );
not g001 ( new_n109_, N108 );
not g002 ( new_n110_, keyIn_0_7 );
and g003 ( new_n111_, new_n110_, N102 );
not g004 ( new_n112_, N102 );
and g005 ( new_n113_, new_n112_, keyIn_0_7 );
or g006 ( new_n114_, new_n111_, new_n113_, new_n109_ );
and g007 ( new_n115_, new_n114_, keyIn_0_13 );
not g008 ( new_n116_, keyIn_0_13 );
not g009 ( new_n117_, new_n111_ );
not g010 ( new_n118_, new_n113_ );
and g011 ( new_n119_, new_n117_, new_n118_, new_n116_, N108 );
or g012 ( new_n120_, new_n115_, new_n119_ );
not g013 ( new_n121_, N76 );
and g014 ( new_n122_, new_n121_, keyIn_0_5 );
not g015 ( new_n123_, keyIn_0_5 );
and g016 ( new_n124_, new_n123_, N76 );
or g017 ( new_n125_, new_n122_, new_n124_ );
and g018 ( new_n126_, new_n125_, keyIn_0_11, N82 );
not g019 ( new_n127_, keyIn_0_11 );
not g020 ( new_n128_, N82 );
or g021 ( new_n129_, new_n123_, N76 );
or g022 ( new_n130_, new_n121_, keyIn_0_5 );
and g023 ( new_n131_, new_n129_, new_n130_ );
or g024 ( new_n132_, new_n131_, new_n128_ );
and g025 ( new_n133_, new_n132_, new_n127_ );
or g026 ( new_n134_, new_n133_, new_n126_ );
not g027 ( new_n135_, keyIn_0_12 );
or g028 ( new_n136_, keyIn_0_6, N89 );
and g029 ( new_n137_, keyIn_0_6, N89 );
not g030 ( new_n138_, new_n137_ );
and g031 ( new_n139_, new_n138_, N95, new_n136_ );
and g032 ( new_n140_, new_n139_, new_n135_ );
not g033 ( new_n141_, new_n140_ );
or g034 ( new_n142_, new_n139_, new_n135_ );
and g035 ( new_n143_, new_n141_, new_n142_ );
and g036 ( new_n144_, new_n134_, new_n120_, new_n143_ );
not g037 ( new_n145_, keyIn_0_9 );
not g038 ( new_n146_, N37 );
and g039 ( new_n147_, new_n146_, keyIn_0_2 );
not g040 ( new_n148_, keyIn_0_2 );
and g041 ( new_n149_, new_n148_, N37 );
or g042 ( new_n150_, new_n147_, new_n149_ );
and g043 ( new_n151_, new_n150_, N43 );
and g044 ( new_n152_, new_n151_, new_n145_ );
not g045 ( new_n153_, N43 );
or g046 ( new_n154_, new_n148_, N37 );
or g047 ( new_n155_, new_n146_, keyIn_0_2 );
and g048 ( new_n156_, new_n154_, new_n155_ );
or g049 ( new_n157_, new_n156_, new_n153_ );
and g050 ( new_n158_, new_n157_, keyIn_0_9 );
or g051 ( new_n159_, new_n158_, new_n152_ );
not g052 ( new_n160_, N4 );
not g053 ( new_n161_, keyIn_0_0 );
and g054 ( new_n162_, new_n161_, N1 );
not g055 ( new_n163_, N1 );
and g056 ( new_n164_, new_n163_, keyIn_0_0 );
or g057 ( new_n165_, new_n162_, new_n164_, new_n160_ );
not g058 ( new_n166_, N11 );
and g059 ( new_n167_, new_n166_, N17 );
not g060 ( new_n168_, new_n167_ );
not g061 ( new_n169_, N69 );
or g062 ( new_n170_, new_n169_, N63 );
and g063 ( new_n171_, new_n165_, new_n168_, new_n170_ );
and g064 ( new_n172_, new_n159_, new_n171_ );
not g065 ( new_n173_, keyIn_0_10 );
and g066 ( new_n174_, keyIn_0_4, N50 );
not g067 ( new_n175_, keyIn_0_4 );
not g068 ( new_n176_, N50 );
and g069 ( new_n177_, new_n175_, new_n176_ );
or g070 ( new_n178_, new_n177_, new_n174_ );
and g071 ( new_n179_, new_n178_, N56 );
or g072 ( new_n180_, new_n179_, new_n173_ );
not g073 ( new_n181_, N56 );
not g074 ( new_n182_, new_n174_ );
or g075 ( new_n183_, keyIn_0_4, N50 );
and g076 ( new_n184_, new_n182_, new_n183_ );
or g077 ( new_n185_, new_n184_, new_n181_ );
or g078 ( new_n186_, new_n185_, keyIn_0_10 );
and g079 ( new_n187_, new_n180_, new_n186_ );
not g080 ( new_n188_, keyIn_0_8 );
not g081 ( new_n189_, N24 );
and g082 ( new_n190_, new_n189_, keyIn_0_1 );
not g083 ( new_n191_, keyIn_0_1 );
and g084 ( new_n192_, new_n191_, N24 );
or g085 ( new_n193_, new_n190_, new_n192_ );
and g086 ( new_n194_, new_n193_, new_n188_, N30 );
not g087 ( new_n195_, N30 );
or g088 ( new_n196_, new_n191_, N24 );
or g089 ( new_n197_, new_n189_, keyIn_0_1 );
and g090 ( new_n198_, new_n196_, new_n197_ );
or g091 ( new_n199_, new_n198_, new_n195_ );
and g092 ( new_n200_, new_n199_, keyIn_0_8 );
or g093 ( new_n201_, new_n200_, new_n194_ );
and g094 ( new_n202_, new_n201_, new_n187_ );
and g095 ( new_n203_, new_n144_, new_n172_, new_n202_, new_n108_ );
not g096 ( new_n204_, new_n203_ );
and g097 ( new_n205_, new_n144_, new_n172_, new_n202_ );
or g098 ( new_n206_, new_n205_, new_n108_ );
and g099 ( N223, new_n206_, new_n204_ );
not g100 ( new_n208_, keyIn_0_27 );
not g101 ( new_n209_, keyIn_0_21 );
not g102 ( new_n210_, keyIn_0_15 );
or g103 ( new_n211_, N223, new_n210_ );
and g104 ( new_n212_, new_n206_, new_n210_, new_n204_ );
not g105 ( new_n213_, new_n212_ );
and g106 ( new_n214_, new_n211_, new_n213_ );
or g107 ( new_n215_, new_n214_, new_n120_ );
and g108 ( new_n216_, new_n214_, new_n120_ );
not g109 ( new_n217_, new_n216_ );
and g110 ( new_n218_, new_n217_, new_n215_ );
or g111 ( new_n219_, new_n218_, new_n209_ );
and g112 ( new_n220_, new_n217_, new_n209_, new_n215_ );
not g113 ( new_n221_, new_n220_ );
not g114 ( new_n222_, N112 );
and g115 ( new_n223_, new_n222_, N108 );
and g116 ( new_n224_, new_n219_, new_n221_, new_n223_ );
and g117 ( new_n225_, new_n224_, new_n208_ );
not g118 ( new_n226_, new_n224_ );
and g119 ( new_n227_, new_n226_, keyIn_0_27 );
or g120 ( new_n228_, new_n227_, new_n225_ );
not g121 ( new_n229_, keyIn_0_26 );
not g122 ( new_n230_, keyIn_0_20 );
or g123 ( new_n231_, new_n214_, new_n170_ );
and g124 ( new_n232_, new_n214_, new_n170_ );
not g125 ( new_n233_, new_n232_ );
and g126 ( new_n234_, new_n233_, new_n231_ );
or g127 ( new_n235_, new_n234_, new_n230_ );
and g128 ( new_n236_, new_n233_, new_n231_, new_n230_ );
not g129 ( new_n237_, new_n236_ );
not g130 ( new_n238_, N73 );
and g131 ( new_n239_, new_n238_, N69 );
and g132 ( new_n240_, new_n235_, new_n237_, new_n239_ );
and g133 ( new_n241_, new_n240_, new_n229_ );
not g134 ( new_n242_, new_n240_ );
and g135 ( new_n243_, new_n242_, keyIn_0_26 );
or g136 ( new_n244_, new_n243_, new_n241_ );
not g137 ( new_n245_, N60 );
or g138 ( new_n246_, new_n214_, new_n187_ );
and g139 ( new_n247_, new_n211_, new_n187_, new_n213_ );
not g140 ( new_n248_, new_n247_ );
and g141 ( new_n249_, new_n246_, keyIn_0_19, new_n248_ );
not g142 ( new_n250_, new_n249_ );
and g143 ( new_n251_, new_n246_, new_n248_ );
or g144 ( new_n252_, new_n251_, keyIn_0_19 );
and g145 ( new_n253_, new_n252_, new_n250_ );
not g146 ( new_n254_, new_n253_ );
and g147 ( new_n255_, new_n254_, keyIn_0_25, N56, new_n245_ );
not g148 ( new_n256_, keyIn_0_25 );
or g149 ( new_n257_, new_n181_, N60 );
or g150 ( new_n258_, new_n253_, new_n257_ );
and g151 ( new_n259_, new_n258_, new_n256_ );
or g152 ( new_n260_, new_n259_, new_n255_ );
and g153 ( new_n261_, new_n260_, new_n228_, new_n244_ );
not g154 ( new_n262_, keyIn_0_22 );
not g155 ( new_n263_, N8 );
not g156 ( new_n264_, keyIn_0_16 );
or g157 ( new_n265_, new_n214_, new_n165_ );
and g158 ( new_n266_, new_n214_, new_n165_ );
not g159 ( new_n267_, new_n266_ );
and g160 ( new_n268_, new_n267_, new_n264_, new_n265_ );
not g161 ( new_n269_, new_n268_ );
and g162 ( new_n270_, new_n267_, new_n265_ );
or g163 ( new_n271_, new_n270_, new_n264_ );
and g164 ( new_n272_, new_n271_, N4, new_n263_, new_n269_ );
and g165 ( new_n273_, new_n272_, new_n262_ );
not g166 ( new_n274_, new_n272_ );
and g167 ( new_n275_, new_n274_, keyIn_0_22 );
or g168 ( new_n276_, new_n275_, new_n273_ );
not g169 ( new_n277_, N99 );
not g170 ( new_n278_, new_n143_ );
not g171 ( new_n279_, new_n214_ );
and g172 ( new_n280_, new_n279_, new_n278_ );
and g173 ( new_n281_, new_n214_, new_n143_ );
or g174 ( new_n282_, new_n280_, new_n281_ );
and g175 ( new_n283_, new_n282_, N95, new_n277_ );
not g176 ( new_n284_, new_n283_ );
not g177 ( new_n285_, N34 );
not g178 ( new_n286_, new_n194_ );
and g179 ( new_n287_, new_n193_, N30 );
or g180 ( new_n288_, new_n287_, new_n188_ );
and g181 ( new_n289_, new_n279_, new_n286_, new_n288_ );
and g182 ( new_n290_, new_n214_, new_n201_ );
or g183 ( new_n291_, new_n289_, new_n290_ );
and g184 ( new_n292_, new_n291_, N30, new_n285_ );
not g185 ( new_n293_, new_n292_ );
not g186 ( new_n294_, N86 );
not g187 ( new_n295_, new_n126_ );
and g188 ( new_n296_, new_n125_, N82 );
or g189 ( new_n297_, new_n296_, keyIn_0_11 );
and g190 ( new_n298_, new_n279_, new_n295_, new_n297_ );
and g191 ( new_n299_, new_n214_, new_n134_ );
or g192 ( new_n300_, new_n298_, new_n299_ );
and g193 ( new_n301_, new_n300_, N82, new_n294_ );
not g194 ( new_n302_, new_n301_ );
and g195 ( new_n303_, new_n293_, new_n302_, new_n284_ );
and g196 ( new_n304_, new_n276_, new_n303_ );
not g197 ( new_n305_, keyIn_0_24 );
not g198 ( new_n306_, keyIn_0_18 );
or g199 ( new_n307_, new_n214_, new_n159_ );
and g200 ( new_n308_, new_n211_, new_n159_, new_n213_ );
not g201 ( new_n309_, new_n308_ );
and g202 ( new_n310_, new_n307_, new_n306_, new_n309_ );
not g203 ( new_n311_, new_n310_ );
and g204 ( new_n312_, new_n307_, new_n309_ );
or g205 ( new_n313_, new_n312_, new_n306_ );
and g206 ( new_n314_, new_n313_, new_n311_ );
not g207 ( new_n315_, new_n314_ );
not g208 ( new_n316_, N47 );
and g209 ( new_n317_, keyIn_0_3, N43 );
not g210 ( new_n318_, new_n317_ );
or g211 ( new_n319_, keyIn_0_3, N43 );
and g212 ( new_n320_, new_n318_, new_n319_ );
not g213 ( new_n321_, new_n320_ );
and g214 ( new_n322_, new_n321_, new_n316_ );
and g215 ( new_n323_, new_n315_, new_n305_, new_n322_ );
not g216 ( new_n324_, new_n322_ );
or g217 ( new_n325_, new_n314_, new_n324_ );
and g218 ( new_n326_, new_n325_, keyIn_0_24 );
or g219 ( new_n327_, new_n326_, new_n323_ );
not g220 ( new_n328_, N21 );
or g221 ( new_n329_, new_n214_, new_n168_ );
and g222 ( new_n330_, new_n214_, new_n168_ );
not g223 ( new_n331_, new_n330_ );
and g224 ( new_n332_, new_n331_, new_n329_ );
and g225 ( new_n333_, new_n332_, keyIn_0_17 );
not g226 ( new_n334_, keyIn_0_17 );
not g227 ( new_n335_, new_n332_ );
and g228 ( new_n336_, new_n335_, new_n334_ );
or g229 ( new_n337_, new_n336_, new_n333_ );
and g230 ( new_n338_, new_n337_, N17, new_n328_ );
or g231 ( new_n339_, new_n338_, keyIn_0_23 );
not g232 ( new_n340_, keyIn_0_23 );
not g233 ( new_n341_, N17 );
not g234 ( new_n342_, new_n337_ );
or g235 ( new_n343_, new_n342_, new_n340_, new_n341_, N21 );
and g236 ( new_n344_, new_n327_, new_n339_, new_n343_ );
and g237 ( new_n345_, new_n261_, new_n344_, new_n304_ );
or g238 ( new_n346_, new_n345_, keyIn_0_28 );
and g239 ( new_n347_, new_n261_, new_n344_, keyIn_0_28, new_n304_ );
not g240 ( new_n348_, new_n347_ );
and g241 ( new_n349_, new_n346_, new_n348_ );
not g242 ( N329, new_n349_ );
not g243 ( new_n351_, keyIn_0_38 );
not g244 ( new_n352_, keyIn_0_32 );
not g245 ( new_n353_, new_n339_ );
not g246 ( new_n354_, new_n343_ );
or g247 ( new_n355_, new_n353_, new_n354_ );
or g248 ( new_n356_, new_n349_, keyIn_0_31 );
and g249 ( new_n357_, new_n346_, keyIn_0_31, new_n348_ );
not g250 ( new_n358_, new_n357_ );
and g251 ( new_n359_, new_n356_, new_n358_ );
or g252 ( new_n360_, new_n359_, new_n355_ );
and g253 ( new_n361_, new_n356_, new_n355_, new_n358_ );
not g254 ( new_n362_, new_n361_ );
and g255 ( new_n363_, new_n360_, new_n352_, new_n362_ );
not g256 ( new_n364_, new_n363_ );
and g257 ( new_n365_, new_n360_, new_n362_ );
or g258 ( new_n366_, new_n365_, new_n352_ );
not g259 ( new_n367_, N27 );
and g260 ( new_n368_, new_n337_, N17, new_n367_ );
and g261 ( new_n369_, new_n366_, new_n351_, new_n364_, new_n368_ );
not g262 ( new_n370_, new_n369_ );
and g263 ( new_n371_, new_n366_, new_n364_, new_n368_ );
or g264 ( new_n372_, new_n371_, new_n351_ );
and g265 ( new_n373_, new_n372_, new_n370_ );
not g266 ( new_n374_, keyIn_0_35 );
not g267 ( new_n375_, new_n244_ );
or g268 ( new_n376_, new_n359_, new_n375_ );
and g269 ( new_n377_, new_n356_, new_n375_, new_n358_ );
not g270 ( new_n378_, new_n377_ );
and g271 ( new_n379_, new_n376_, new_n374_, new_n378_ );
not g272 ( new_n380_, new_n379_ );
and g273 ( new_n381_, new_n376_, new_n378_ );
or g274 ( new_n382_, new_n381_, new_n374_ );
not g275 ( new_n383_, N79 );
and g276 ( new_n384_, new_n235_, new_n237_ );
and g277 ( new_n385_, new_n384_, N69, new_n383_ );
and g278 ( new_n386_, new_n385_, keyIn_0_29 );
not g279 ( new_n387_, keyIn_0_29 );
not g280 ( new_n388_, new_n385_ );
and g281 ( new_n389_, new_n388_, new_n387_ );
or g282 ( new_n390_, new_n389_, new_n386_ );
and g283 ( new_n391_, new_n382_, keyIn_0_41, new_n380_, new_n390_ );
not g284 ( new_n392_, new_n391_ );
and g285 ( new_n393_, new_n382_, new_n380_, new_n390_ );
or g286 ( new_n394_, new_n393_, keyIn_0_41 );
and g287 ( new_n395_, new_n394_, new_n392_ );
not g288 ( new_n396_, new_n228_ );
and g289 ( new_n397_, new_n356_, new_n396_, new_n358_ );
not g290 ( new_n398_, new_n397_ );
or g291 ( new_n399_, new_n359_, new_n396_ );
and g292 ( new_n400_, new_n399_, new_n398_ );
or g293 ( new_n401_, new_n400_, keyIn_0_37 );
not g294 ( new_n402_, new_n401_ );
and g295 ( new_n403_, new_n399_, keyIn_0_37, new_n398_ );
not g296 ( new_n404_, keyIn_0_30 );
not g297 ( new_n405_, N115 );
and g298 ( new_n406_, new_n219_, N108, new_n405_, new_n221_ );
or g299 ( new_n407_, new_n406_, new_n404_ );
and g300 ( new_n408_, new_n406_, new_n404_ );
not g301 ( new_n409_, new_n408_ );
and g302 ( new_n410_, new_n409_, new_n407_ );
or g303 ( new_n411_, new_n402_, keyIn_0_43, new_n403_, new_n410_ );
not g304 ( new_n412_, keyIn_0_43 );
not g305 ( new_n413_, new_n403_ );
not g306 ( new_n414_, new_n410_ );
and g307 ( new_n415_, new_n401_, new_n413_, new_n414_ );
or g308 ( new_n416_, new_n415_, new_n412_ );
and g309 ( new_n417_, new_n416_, new_n411_ );
or g310 ( new_n418_, new_n373_, new_n395_, new_n417_ );
not g311 ( new_n419_, keyIn_0_33 );
or g312 ( new_n420_, new_n359_, new_n292_ );
and g313 ( new_n421_, new_n359_, new_n292_ );
not g314 ( new_n422_, new_n421_ );
and g315 ( new_n423_, new_n422_, new_n419_, new_n420_ );
not g316 ( new_n424_, new_n423_ );
and g317 ( new_n425_, new_n422_, new_n420_ );
or g318 ( new_n426_, new_n425_, new_n419_ );
not g319 ( new_n427_, N40 );
and g320 ( new_n428_, new_n291_, N30, new_n427_ );
and g321 ( new_n429_, new_n426_, keyIn_0_39, new_n424_, new_n428_ );
not g322 ( new_n430_, new_n429_ );
not g323 ( new_n431_, keyIn_0_42 );
and g324 ( new_n432_, new_n356_, new_n283_, new_n358_ );
not g325 ( new_n433_, new_n432_ );
or g326 ( new_n434_, new_n359_, new_n283_ );
and g327 ( new_n435_, new_n434_, new_n433_ );
or g328 ( new_n436_, new_n435_, keyIn_0_36 );
and g329 ( new_n437_, new_n434_, keyIn_0_36, new_n433_ );
not g330 ( new_n438_, new_n437_ );
not g331 ( new_n439_, N105 );
and g332 ( new_n440_, new_n282_, N95, new_n439_ );
and g333 ( new_n441_, new_n436_, new_n438_, new_n440_ );
or g334 ( new_n442_, new_n441_, new_n431_ );
not g335 ( new_n443_, new_n436_ );
not g336 ( new_n444_, N95 );
not g337 ( new_n445_, new_n282_ );
or g338 ( new_n446_, new_n437_, new_n444_, N105, new_n445_ );
or g339 ( new_n447_, new_n446_, new_n443_, keyIn_0_42 );
and g340 ( new_n448_, new_n442_, new_n430_, new_n447_ );
not g341 ( new_n449_, new_n448_ );
not g342 ( new_n450_, keyIn_0_34 );
not g343 ( new_n451_, new_n260_ );
or g344 ( new_n452_, new_n359_, new_n451_ );
and g345 ( new_n453_, new_n356_, new_n451_, new_n358_ );
not g346 ( new_n454_, new_n453_ );
and g347 ( new_n455_, new_n452_, new_n450_, new_n454_ );
not g348 ( new_n456_, new_n455_ );
and g349 ( new_n457_, new_n452_, new_n454_ );
or g350 ( new_n458_, new_n457_, new_n450_ );
not g351 ( new_n459_, N66 );
and g352 ( new_n460_, new_n254_, N56, new_n459_ );
and g353 ( new_n461_, new_n458_, keyIn_0_40, new_n456_, new_n460_ );
not g354 ( new_n462_, new_n461_ );
and g355 ( new_n463_, new_n458_, new_n456_, new_n460_ );
or g356 ( new_n464_, new_n463_, keyIn_0_40 );
and g357 ( new_n465_, new_n464_, new_n462_ );
not g358 ( new_n466_, keyIn_0_39 );
and g359 ( new_n467_, new_n426_, new_n424_, new_n428_ );
not g360 ( new_n468_, new_n467_ );
and g361 ( new_n469_, new_n468_, new_n466_ );
not g362 ( new_n470_, new_n300_ );
or g363 ( new_n471_, new_n359_, new_n301_ );
and g364 ( new_n472_, new_n359_, new_n301_ );
not g365 ( new_n473_, new_n472_ );
and g366 ( new_n474_, new_n473_, new_n471_ );
or g367 ( new_n475_, new_n474_, new_n128_, N92, new_n470_ );
not g368 ( new_n476_, new_n276_ );
or g369 ( new_n477_, new_n359_, new_n476_ );
and g370 ( new_n478_, new_n359_, new_n476_ );
not g371 ( new_n479_, new_n478_ );
and g372 ( new_n480_, new_n479_, new_n477_ );
not g373 ( new_n481_, N14 );
and g374 ( new_n482_, new_n271_, N4, new_n481_, new_n269_ );
not g375 ( new_n483_, new_n482_ );
or g376 ( new_n484_, new_n480_, new_n483_ );
not g377 ( new_n485_, new_n327_ );
or g378 ( new_n486_, new_n359_, new_n485_ );
and g379 ( new_n487_, new_n359_, new_n485_ );
not g380 ( new_n488_, new_n487_ );
and g381 ( new_n489_, new_n488_, new_n486_ );
or g382 ( new_n490_, new_n489_, N53, new_n314_, new_n320_ );
and g383 ( new_n491_, new_n475_, new_n490_, new_n484_ );
not g384 ( new_n492_, new_n491_ );
or g385 ( new_n493_, new_n465_, new_n469_, new_n492_ );
or g386 ( new_n494_, new_n418_, new_n449_, new_n493_ );
and g387 ( new_n495_, new_n494_, keyIn_0_44 );
not g388 ( new_n496_, keyIn_0_44 );
not g389 ( new_n497_, new_n373_ );
not g390 ( new_n498_, new_n395_ );
not g391 ( new_n499_, new_n417_ );
and g392 ( new_n500_, new_n497_, new_n498_, new_n499_ );
not g393 ( new_n501_, new_n465_ );
or g394 ( new_n502_, new_n467_, keyIn_0_39 );
and g395 ( new_n503_, new_n502_, new_n491_ );
and g396 ( new_n504_, new_n501_, new_n448_, new_n503_ );
and g397 ( new_n505_, new_n500_, new_n504_, new_n496_ );
or g398 ( N370, new_n495_, new_n505_ );
not g399 ( new_n507_, keyIn_0_54 );
not g400 ( new_n508_, keyIn_0_45 );
and g401 ( new_n509_, new_n500_, new_n504_ );
or g402 ( new_n510_, new_n509_, new_n496_ );
not g403 ( new_n511_, new_n505_ );
and g404 ( new_n512_, new_n510_, new_n508_, new_n511_ );
not g405 ( new_n513_, new_n512_ );
and g406 ( new_n514_, new_n510_, new_n511_ );
or g407 ( new_n515_, new_n514_, new_n508_ );
and g408 ( new_n516_, new_n515_, new_n513_ );
or g409 ( new_n517_, new_n516_, new_n459_ );
or g410 ( new_n518_, new_n517_, keyIn_0_49 );
and g411 ( new_n519_, new_n517_, keyIn_0_49 );
not g412 ( new_n520_, new_n519_ );
and g413 ( new_n521_, new_n520_, new_n518_ );
and g414 ( new_n522_, N329, N60 );
and g415 ( new_n523_, N223, N50 );
or g416 ( new_n524_, new_n522_, new_n181_, new_n523_ );
or g417 ( new_n525_, new_n521_, new_n524_ );
and g418 ( new_n526_, new_n525_, new_n507_ );
not g419 ( new_n527_, keyIn_0_49 );
and g420 ( new_n528_, N370, keyIn_0_45 );
or g421 ( new_n529_, new_n528_, new_n512_ );
and g422 ( new_n530_, new_n529_, N66 );
and g423 ( new_n531_, new_n530_, new_n527_ );
or g424 ( new_n532_, new_n531_, new_n519_ );
not g425 ( new_n533_, new_n524_ );
and g426 ( new_n534_, new_n532_, keyIn_0_54, new_n533_ );
or g427 ( new_n535_, new_n526_, new_n534_ );
not g428 ( new_n536_, keyIn_0_48 );
and g429 ( new_n537_, new_n529_, new_n536_, N53 );
not g430 ( new_n538_, N53 );
or g431 ( new_n539_, new_n516_, new_n538_ );
and g432 ( new_n540_, new_n539_, keyIn_0_48 );
or g433 ( new_n541_, new_n540_, new_n537_ );
and g434 ( new_n542_, N329, N47 );
not g435 ( new_n543_, new_n542_ );
and g436 ( new_n544_, N223, N37 );
not g437 ( new_n545_, new_n544_ );
and g438 ( new_n546_, new_n543_, N43, new_n545_ );
and g439 ( new_n547_, new_n541_, keyIn_0_53, new_n546_ );
not g440 ( new_n548_, new_n547_ );
and g441 ( new_n549_, new_n541_, new_n546_ );
or g442 ( new_n550_, new_n549_, keyIn_0_53 );
and g443 ( new_n551_, new_n550_, new_n548_ );
and g444 ( new_n552_, new_n535_, new_n551_ );
not g445 ( new_n553_, new_n552_ );
not g446 ( new_n554_, keyIn_0_46 );
and g447 ( new_n555_, new_n529_, new_n554_, N27 );
or g448 ( new_n556_, new_n516_, new_n367_ );
and g449 ( new_n557_, new_n556_, keyIn_0_46 );
or g450 ( new_n558_, new_n557_, new_n555_ );
or g451 ( new_n559_, new_n349_, new_n328_ );
and g452 ( new_n560_, N223, N11 );
not g453 ( new_n561_, new_n560_ );
and g454 ( new_n562_, new_n559_, N17, new_n561_ );
and g455 ( new_n563_, new_n558_, keyIn_0_51, new_n562_ );
not g456 ( new_n564_, new_n563_ );
and g457 ( new_n565_, new_n558_, new_n562_ );
or g458 ( new_n566_, new_n565_, keyIn_0_51 );
and g459 ( new_n567_, new_n529_, keyIn_0_47, N40 );
not g460 ( new_n568_, keyIn_0_47 );
or g461 ( new_n569_, new_n516_, new_n427_ );
and g462 ( new_n570_, new_n569_, new_n568_ );
or g463 ( new_n571_, new_n570_, new_n567_ );
and g464 ( new_n572_, N329, N34 );
not g465 ( new_n573_, new_n572_ );
and g466 ( new_n574_, N223, N24 );
not g467 ( new_n575_, new_n574_ );
and g468 ( new_n576_, new_n573_, N30, new_n575_ );
and g469 ( new_n577_, new_n571_, keyIn_0_52, new_n576_ );
not g470 ( new_n578_, new_n577_ );
and g471 ( new_n579_, new_n571_, new_n576_ );
or g472 ( new_n580_, new_n579_, keyIn_0_52 );
and g473 ( new_n581_, new_n566_, new_n580_, new_n564_, new_n578_ );
not g474 ( new_n582_, new_n581_ );
not g475 ( new_n583_, keyIn_0_55 );
not g476 ( new_n584_, keyIn_0_50 );
and g477 ( new_n585_, new_n529_, N79 );
and g478 ( new_n586_, new_n585_, new_n584_ );
or g479 ( new_n587_, new_n516_, new_n383_ );
and g480 ( new_n588_, new_n587_, keyIn_0_50 );
or g481 ( new_n589_, new_n586_, new_n588_ );
and g482 ( new_n590_, N329, N73 );
and g483 ( new_n591_, N223, N63 );
or g484 ( new_n592_, new_n590_, new_n169_, new_n591_ );
not g485 ( new_n593_, new_n592_ );
and g486 ( new_n594_, new_n589_, new_n593_ );
or g487 ( new_n595_, new_n594_, new_n583_ );
and g488 ( new_n596_, new_n589_, new_n583_, new_n593_ );
not g489 ( new_n597_, new_n596_ );
and g490 ( new_n598_, new_n595_, new_n597_ );
and g491 ( new_n599_, new_n529_, N115 );
and g492 ( new_n600_, N329, N112 );
and g493 ( new_n601_, N223, N102 );
or g494 ( new_n602_, new_n599_, new_n109_, new_n600_, new_n601_ );
and g495 ( new_n603_, new_n529_, N92 );
and g496 ( new_n604_, N329, N86 );
and g497 ( new_n605_, N223, N76 );
or g498 ( new_n606_, new_n603_, new_n128_, new_n604_, new_n605_ );
and g499 ( new_n607_, new_n529_, N105 );
and g500 ( new_n608_, N329, N99 );
and g501 ( new_n609_, N223, N89 );
or g502 ( new_n610_, new_n607_, new_n444_, new_n608_, new_n609_ );
and g503 ( new_n611_, new_n602_, new_n606_, new_n610_ );
not g504 ( new_n612_, new_n611_ );
or g505 ( new_n613_, new_n598_, new_n612_ );
or g506 ( new_n614_, new_n553_, new_n613_, keyIn_0_56, new_n582_ );
not g507 ( new_n615_, keyIn_0_56 );
or g508 ( new_n616_, new_n587_, keyIn_0_50 );
or g509 ( new_n617_, new_n585_, new_n584_ );
and g510 ( new_n618_, new_n617_, new_n616_ );
or g511 ( new_n619_, new_n618_, new_n592_ );
and g512 ( new_n620_, new_n619_, keyIn_0_55 );
or g513 ( new_n621_, new_n620_, new_n596_ );
and g514 ( new_n622_, new_n581_, new_n621_, new_n611_ );
and g515 ( new_n623_, new_n622_, new_n552_ );
or g516 ( new_n624_, new_n623_, new_n615_ );
and g517 ( new_n625_, new_n624_, new_n614_ );
and g518 ( new_n626_, new_n529_, N14 );
and g519 ( new_n627_, N329, N8 );
and g520 ( new_n628_, N223, N1 );
or g521 ( new_n629_, new_n626_, new_n160_, new_n627_, new_n628_ );
not g522 ( new_n630_, new_n629_ );
or g523 ( new_n631_, new_n625_, new_n630_ );
and g524 ( new_n632_, new_n631_, keyIn_0_58 );
not g525 ( new_n633_, keyIn_0_58 );
not g526 ( new_n634_, new_n625_ );
and g527 ( new_n635_, new_n634_, new_n633_, new_n629_ );
or g528 ( N421, new_n632_, new_n635_ );
not g529 ( new_n637_, keyIn_0_61 );
and g530 ( new_n638_, new_n580_, new_n578_ );
or g531 ( new_n639_, new_n551_, keyIn_0_57 );
and g532 ( new_n640_, new_n550_, keyIn_0_57, new_n548_ );
not g533 ( new_n641_, new_n640_ );
and g534 ( new_n642_, new_n639_, keyIn_0_59, new_n638_, new_n641_ );
not g535 ( new_n643_, new_n642_ );
and g536 ( new_n644_, new_n639_, new_n638_, new_n641_ );
or g537 ( new_n645_, new_n644_, keyIn_0_59 );
and g538 ( new_n646_, new_n645_, new_n643_ );
and g539 ( new_n647_, new_n535_, new_n581_ );
not g540 ( new_n648_, new_n647_ );
or g541 ( new_n649_, new_n646_, new_n648_ );
and g542 ( new_n650_, new_n649_, new_n637_ );
not g543 ( new_n651_, new_n646_ );
and g544 ( new_n652_, new_n651_, keyIn_0_61, new_n647_ );
or g545 ( N430, new_n650_, new_n652_ );
and g546 ( new_n654_, new_n535_, new_n598_, new_n551_, new_n638_ );
or g547 ( new_n655_, new_n654_, keyIn_0_60 );
and g548 ( new_n656_, new_n551_, new_n638_ );
and g549 ( new_n657_, new_n656_, new_n535_, keyIn_0_60, new_n598_ );
not g550 ( new_n658_, new_n657_ );
and g551 ( new_n659_, new_n655_, new_n658_ );
or g552 ( new_n660_, new_n553_, new_n606_ );
and g553 ( new_n661_, new_n660_, new_n581_ );
and g554 ( new_n662_, new_n661_, new_n659_ );
and g555 ( new_n663_, new_n662_, keyIn_0_62 );
not g556 ( new_n664_, keyIn_0_62 );
not g557 ( new_n665_, new_n662_ );
and g558 ( new_n666_, new_n665_, new_n664_ );
or g559 ( N431, new_n666_, new_n663_ );
not g560 ( new_n668_, keyIn_0_63 );
not g561 ( new_n669_, new_n610_ );
and g562 ( new_n670_, new_n551_, new_n638_, new_n606_, new_n669_ );
not g563 ( new_n671_, new_n670_ );
and g564 ( new_n672_, new_n671_, new_n564_, new_n566_ );
and g565 ( new_n673_, new_n672_, new_n655_, new_n658_ );
not g566 ( new_n674_, new_n673_ );
or g567 ( new_n675_, new_n674_, new_n646_ );
and g568 ( new_n676_, new_n675_, new_n668_ );
and g569 ( new_n677_, new_n651_, keyIn_0_63, new_n673_ );
or g570 ( N432, new_n676_, new_n677_ );
endmodule