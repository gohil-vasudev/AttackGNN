module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n639_, new_n484_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n310_, new_n144_, new_n275_, new_n352_, new_n485_, new_n525_, new_n562_, new_n578_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n598_, new_n824_, new_n143_, new_n520_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n825_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n772_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n435_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n756_, new_n495_, new_n823_, new_n431_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n138_, N85 );
nand g001 ( new_n139_, new_n138_, N81 );
not g002 ( new_n140_, N81 );
nand g003 ( new_n141_, new_n140_, N85 );
not g004 ( new_n142_, N89 );
not g005 ( new_n143_, N93 );
nand g006 ( new_n144_, new_n142_, new_n143_ );
nand g007 ( new_n145_, N89, N93 );
nand g008 ( new_n146_, new_n144_, new_n139_, new_n141_, new_n145_ );
nand g009 ( new_n147_, new_n139_, new_n141_ );
nand g010 ( new_n148_, new_n144_, new_n145_ );
nand g011 ( new_n149_, new_n147_, new_n148_ );
nand g012 ( new_n150_, new_n149_, new_n146_ );
not g013 ( new_n151_, new_n150_ );
not g014 ( new_n152_, N69 );
nand g015 ( new_n153_, new_n152_, N65 );
not g016 ( new_n154_, N65 );
nand g017 ( new_n155_, new_n154_, N69 );
not g018 ( new_n156_, N73 );
not g019 ( new_n157_, N77 );
nand g020 ( new_n158_, new_n156_, new_n157_ );
nand g021 ( new_n159_, N73, N77 );
nand g022 ( new_n160_, new_n158_, new_n153_, new_n155_, new_n159_ );
nand g023 ( new_n161_, new_n153_, new_n155_ );
nand g024 ( new_n162_, new_n158_, new_n159_ );
nand g025 ( new_n163_, new_n161_, new_n162_ );
nand g026 ( new_n164_, new_n163_, new_n160_ );
nand g027 ( new_n165_, new_n151_, new_n164_ );
not g028 ( new_n166_, new_n164_ );
nand g029 ( new_n167_, new_n166_, new_n150_ );
nand g030 ( new_n168_, new_n165_, new_n167_ );
nand g031 ( new_n169_, N129, N137 );
nand g032 ( new_n170_, new_n168_, new_n169_ );
nand g033 ( new_n171_, new_n165_, new_n167_, N129, N137 );
not g034 ( new_n172_, N17 );
nand g035 ( new_n173_, new_n172_, N1 );
not g036 ( new_n174_, N1 );
nand g037 ( new_n175_, new_n174_, N17 );
not g038 ( new_n176_, N33 );
not g039 ( new_n177_, N49 );
nand g040 ( new_n178_, new_n176_, new_n177_ );
nand g041 ( new_n179_, N33, N49 );
nand g042 ( new_n180_, new_n178_, new_n173_, new_n175_, new_n179_ );
nand g043 ( new_n181_, new_n173_, new_n175_ );
nand g044 ( new_n182_, new_n178_, new_n179_ );
nand g045 ( new_n183_, new_n181_, new_n182_ );
nand g046 ( new_n184_, new_n170_, new_n171_, new_n180_, new_n183_ );
nand g047 ( new_n185_, new_n170_, new_n171_ );
nand g048 ( new_n186_, new_n183_, new_n180_ );
nand g049 ( new_n187_, new_n185_, new_n186_ );
nand g050 ( new_n188_, new_n187_, new_n184_ );
not g051 ( new_n189_, keyIn_0_23 );
not g052 ( new_n190_, keyIn_0_19 );
not g053 ( new_n191_, N9 );
not g054 ( new_n192_, N13 );
nand g055 ( new_n193_, new_n191_, new_n192_ );
nand g056 ( new_n194_, N9, N13 );
nand g057 ( new_n195_, new_n193_, new_n194_ );
nand g058 ( new_n196_, new_n195_, keyIn_0_1 );
not g059 ( new_n197_, keyIn_0_1 );
nand g060 ( new_n198_, new_n193_, new_n197_, new_n194_ );
not g061 ( new_n199_, N5 );
nand g062 ( new_n200_, new_n174_, new_n199_ );
nand g063 ( new_n201_, N1, N5 );
nand g064 ( new_n202_, new_n200_, keyIn_0_0, new_n201_ );
not g065 ( new_n203_, keyIn_0_0 );
nand g066 ( new_n204_, new_n200_, new_n201_ );
nand g067 ( new_n205_, new_n204_, new_n203_ );
nand g068 ( new_n206_, new_n205_, new_n202_ );
nand g069 ( new_n207_, new_n206_, new_n196_, new_n198_ );
nand g070 ( new_n208_, new_n196_, new_n198_ );
nand g071 ( new_n209_, new_n208_, new_n202_, new_n205_ );
nand g072 ( new_n210_, new_n207_, new_n209_, keyIn_0_12 );
not g073 ( new_n211_, keyIn_0_12 );
nand g074 ( new_n212_, new_n207_, new_n209_ );
nand g075 ( new_n213_, new_n212_, new_n211_ );
not g076 ( new_n214_, keyIn_0_14 );
not g077 ( new_n215_, N41 );
not g078 ( new_n216_, N45 );
nand g079 ( new_n217_, new_n215_, new_n216_ );
nand g080 ( new_n218_, N41, N45 );
nand g081 ( new_n219_, new_n217_, new_n218_ );
nand g082 ( new_n220_, new_n219_, keyIn_0_5 );
not g083 ( new_n221_, keyIn_0_5 );
nand g084 ( new_n222_, new_n217_, new_n221_, new_n218_ );
nand g085 ( new_n223_, new_n220_, new_n222_ );
not g086 ( new_n224_, N37 );
nand g087 ( new_n225_, new_n176_, new_n224_ );
nand g088 ( new_n226_, N33, N37 );
nand g089 ( new_n227_, new_n225_, new_n226_ );
nand g090 ( new_n228_, new_n227_, keyIn_0_4 );
not g091 ( new_n229_, keyIn_0_4 );
nand g092 ( new_n230_, new_n225_, new_n229_, new_n226_ );
nand g093 ( new_n231_, new_n228_, new_n230_ );
nand g094 ( new_n232_, new_n223_, new_n231_ );
nand g095 ( new_n233_, new_n220_, new_n228_, new_n222_, new_n230_ );
nand g096 ( new_n234_, new_n232_, new_n233_ );
nand g097 ( new_n235_, new_n234_, new_n214_ );
nand g098 ( new_n236_, new_n232_, keyIn_0_14, new_n233_ );
nand g099 ( new_n237_, new_n213_, new_n235_, new_n210_, new_n236_ );
nand g100 ( new_n238_, new_n213_, new_n210_ );
nand g101 ( new_n239_, new_n235_, new_n236_ );
nand g102 ( new_n240_, new_n238_, new_n239_ );
nand g103 ( new_n241_, new_n240_, new_n190_, new_n237_ );
nand g104 ( new_n242_, new_n240_, new_n237_ );
nand g105 ( new_n243_, new_n242_, keyIn_0_19 );
nand g106 ( new_n244_, new_n243_, new_n241_ );
nand g107 ( new_n245_, keyIn_0_7, N135, N137 );
not g108 ( new_n246_, keyIn_0_7 );
nand g109 ( new_n247_, N135, N137 );
nand g110 ( new_n248_, new_n247_, new_n246_ );
nand g111 ( new_n249_, new_n248_, new_n245_ );
nand g112 ( new_n250_, new_n244_, new_n249_ );
nand g113 ( new_n251_, new_n243_, new_n241_, new_n245_, new_n248_ );
nand g114 ( new_n252_, new_n250_, new_n251_ );
nand g115 ( new_n253_, new_n252_, keyIn_0_21 );
not g116 ( new_n254_, keyIn_0_21 );
nand g117 ( new_n255_, new_n250_, new_n254_, new_n251_ );
nand g118 ( new_n256_, new_n253_, new_n255_ );
not g119 ( new_n257_, keyIn_0_17 );
nand g120 ( new_n258_, new_n142_, N73 );
nand g121 ( new_n259_, new_n156_, N89 );
nand g122 ( new_n260_, new_n258_, new_n259_ );
nand g123 ( new_n261_, new_n260_, keyIn_0_10 );
not g124 ( new_n262_, keyIn_0_10 );
nand g125 ( new_n263_, new_n258_, new_n259_, new_n262_ );
not g126 ( new_n264_, N121 );
nand g127 ( new_n265_, new_n264_, N105 );
not g128 ( new_n266_, N105 );
nand g129 ( new_n267_, new_n266_, N121 );
nand g130 ( new_n268_, new_n265_, new_n267_ );
nand g131 ( new_n269_, new_n268_, keyIn_0_11 );
not g132 ( new_n270_, keyIn_0_11 );
nand g133 ( new_n271_, new_n265_, new_n267_, new_n270_ );
nand g134 ( new_n272_, new_n261_, new_n269_, new_n263_, new_n271_ );
nand g135 ( new_n273_, new_n261_, new_n263_ );
nand g136 ( new_n274_, new_n269_, new_n271_ );
nand g137 ( new_n275_, new_n273_, new_n274_ );
nand g138 ( new_n276_, new_n275_, new_n272_ );
nand g139 ( new_n277_, new_n276_, new_n257_ );
nand g140 ( new_n278_, new_n275_, keyIn_0_17, new_n272_ );
nand g141 ( new_n279_, new_n277_, new_n278_ );
not g142 ( new_n280_, new_n279_ );
nand g143 ( new_n281_, new_n256_, new_n280_ );
nand g144 ( new_n282_, new_n253_, new_n255_, new_n279_ );
nand g145 ( new_n283_, new_n281_, new_n189_, new_n282_ );
nand g146 ( new_n284_, new_n281_, new_n282_ );
nand g147 ( new_n285_, new_n284_, keyIn_0_23 );
nand g148 ( new_n286_, new_n285_, new_n283_ );
not g149 ( new_n287_, new_n286_ );
not g150 ( new_n288_, keyIn_0_24 );
nand g151 ( new_n289_, new_n188_, new_n288_ );
not g152 ( new_n290_, new_n188_ );
nand g153 ( new_n291_, new_n290_, keyIn_0_24 );
not g154 ( new_n292_, N101 );
nand g155 ( new_n293_, new_n292_, N97 );
not g156 ( new_n294_, N97 );
nand g157 ( new_n295_, new_n294_, N101 );
not g158 ( new_n296_, N109 );
nand g159 ( new_n297_, new_n266_, new_n296_ );
nand g160 ( new_n298_, N105, N109 );
nand g161 ( new_n299_, new_n297_, new_n293_, new_n295_, new_n298_ );
nand g162 ( new_n300_, new_n293_, new_n295_ );
nand g163 ( new_n301_, new_n297_, new_n298_ );
nand g164 ( new_n302_, new_n300_, new_n301_ );
nand g165 ( new_n303_, new_n302_, new_n299_ );
not g166 ( new_n304_, new_n303_ );
not g167 ( new_n305_, N117 );
nand g168 ( new_n306_, new_n305_, N113 );
not g169 ( new_n307_, N113 );
nand g170 ( new_n308_, new_n307_, N117 );
not g171 ( new_n309_, N125 );
nand g172 ( new_n310_, new_n264_, new_n309_ );
nand g173 ( new_n311_, N121, N125 );
nand g174 ( new_n312_, new_n310_, new_n306_, new_n308_, new_n311_ );
nand g175 ( new_n313_, new_n306_, new_n308_ );
nand g176 ( new_n314_, new_n310_, new_n311_ );
nand g177 ( new_n315_, new_n313_, new_n314_ );
nand g178 ( new_n316_, new_n315_, new_n312_ );
nand g179 ( new_n317_, new_n304_, new_n316_ );
not g180 ( new_n318_, new_n316_ );
nand g181 ( new_n319_, new_n318_, new_n303_ );
nand g182 ( new_n320_, new_n317_, new_n319_ );
nand g183 ( new_n321_, N130, N137 );
nand g184 ( new_n322_, new_n320_, new_n321_ );
nand g185 ( new_n323_, new_n317_, new_n319_, N130, N137 );
not g186 ( new_n324_, N21 );
nand g187 ( new_n325_, new_n324_, N5 );
nand g188 ( new_n326_, new_n199_, N21 );
not g189 ( new_n327_, N53 );
nand g190 ( new_n328_, new_n224_, new_n327_ );
nand g191 ( new_n329_, N37, N53 );
nand g192 ( new_n330_, new_n328_, new_n325_, new_n326_, new_n329_ );
nand g193 ( new_n331_, new_n325_, new_n326_ );
nand g194 ( new_n332_, new_n328_, new_n329_ );
nand g195 ( new_n333_, new_n331_, new_n332_ );
nand g196 ( new_n334_, new_n322_, new_n323_, new_n330_, new_n333_ );
nand g197 ( new_n335_, new_n322_, new_n323_ );
nand g198 ( new_n336_, new_n333_, new_n330_ );
nand g199 ( new_n337_, new_n335_, new_n336_ );
nand g200 ( new_n338_, new_n337_, new_n334_ );
nand g201 ( new_n339_, new_n304_, new_n164_ );
nand g202 ( new_n340_, new_n166_, new_n303_ );
nand g203 ( new_n341_, new_n339_, new_n340_ );
nand g204 ( new_n342_, N131, N137 );
nand g205 ( new_n343_, new_n341_, new_n342_ );
nand g206 ( new_n344_, new_n339_, new_n340_, N131, N137 );
not g207 ( new_n345_, N25 );
nand g208 ( new_n346_, new_n345_, N9 );
nand g209 ( new_n347_, new_n191_, N25 );
not g210 ( new_n348_, N57 );
nand g211 ( new_n349_, new_n215_, new_n348_ );
nand g212 ( new_n350_, N41, N57 );
nand g213 ( new_n351_, new_n349_, new_n346_, new_n347_, new_n350_ );
nand g214 ( new_n352_, new_n346_, new_n347_ );
nand g215 ( new_n353_, new_n349_, new_n350_ );
nand g216 ( new_n354_, new_n352_, new_n353_ );
nand g217 ( new_n355_, new_n343_, new_n344_, new_n351_, new_n354_ );
nand g218 ( new_n356_, new_n343_, new_n344_ );
nand g219 ( new_n357_, new_n354_, new_n351_ );
nand g220 ( new_n358_, new_n356_, new_n357_ );
nand g221 ( new_n359_, new_n358_, new_n355_ );
not g222 ( new_n360_, new_n359_ );
nand g223 ( new_n361_, new_n291_, new_n289_, new_n338_, new_n360_ );
nand g224 ( new_n362_, new_n290_, new_n338_, new_n359_ );
not g225 ( new_n363_, new_n338_ );
nand g226 ( new_n364_, new_n363_, new_n188_, new_n359_ );
nand g227 ( new_n365_, new_n361_, new_n362_, new_n364_ );
nand g228 ( new_n366_, new_n318_, new_n150_ );
nand g229 ( new_n367_, new_n151_, new_n316_ );
nand g230 ( new_n368_, new_n366_, new_n367_ );
nand g231 ( new_n369_, N132, N137 );
nand g232 ( new_n370_, new_n368_, new_n369_ );
nand g233 ( new_n371_, new_n366_, new_n367_, N132, N137 );
not g234 ( new_n372_, keyIn_0_15 );
not g235 ( new_n373_, N29 );
nand g236 ( new_n374_, new_n373_, N13 );
nand g237 ( new_n375_, new_n192_, N29 );
not g238 ( new_n376_, N61 );
nand g239 ( new_n377_, new_n216_, new_n376_ );
nand g240 ( new_n378_, N45, N61 );
nand g241 ( new_n379_, new_n377_, new_n374_, new_n375_, new_n378_ );
nand g242 ( new_n380_, new_n374_, new_n375_ );
nand g243 ( new_n381_, new_n377_, new_n378_ );
nand g244 ( new_n382_, new_n380_, new_n381_ );
nand g245 ( new_n383_, new_n382_, new_n372_, new_n379_ );
nand g246 ( new_n384_, new_n382_, new_n379_ );
nand g247 ( new_n385_, new_n384_, keyIn_0_15 );
nand g248 ( new_n386_, new_n370_, new_n371_, new_n383_, new_n385_ );
nand g249 ( new_n387_, new_n370_, new_n371_ );
nand g250 ( new_n388_, new_n385_, new_n383_ );
nand g251 ( new_n389_, new_n387_, new_n388_ );
nand g252 ( new_n390_, new_n389_, new_n386_ );
nand g253 ( new_n391_, new_n365_, new_n390_ );
not g254 ( new_n392_, new_n390_ );
nand g255 ( new_n393_, new_n392_, new_n188_, new_n338_, new_n359_ );
nand g256 ( new_n394_, new_n391_, new_n393_ );
nand g257 ( new_n395_, new_n172_, new_n324_ );
nand g258 ( new_n396_, N17, N21 );
nand g259 ( new_n397_, new_n395_, new_n396_ );
nand g260 ( new_n398_, new_n397_, keyIn_0_2 );
not g261 ( new_n399_, keyIn_0_2 );
nand g262 ( new_n400_, new_n395_, new_n399_, new_n396_ );
nand g263 ( new_n401_, new_n398_, new_n400_ );
nand g264 ( new_n402_, new_n345_, new_n373_ );
nand g265 ( new_n403_, N25, N29 );
nand g266 ( new_n404_, new_n402_, new_n403_ );
nand g267 ( new_n405_, new_n404_, keyIn_0_3 );
not g268 ( new_n406_, keyIn_0_3 );
nand g269 ( new_n407_, new_n402_, new_n406_, new_n403_ );
nand g270 ( new_n408_, new_n405_, new_n407_ );
nand g271 ( new_n409_, new_n401_, new_n408_ );
nand g272 ( new_n410_, new_n398_, new_n405_, new_n400_, new_n407_ );
nand g273 ( new_n411_, new_n409_, new_n410_ );
nand g274 ( new_n412_, new_n411_, keyIn_0_13 );
not g275 ( new_n413_, keyIn_0_13 );
nand g276 ( new_n414_, new_n409_, new_n413_, new_n410_ );
nand g277 ( new_n415_, new_n412_, new_n414_ );
nand g278 ( new_n416_, new_n177_, new_n327_ );
nand g279 ( new_n417_, N49, N53 );
nand g280 ( new_n418_, new_n348_, new_n376_ );
nand g281 ( new_n419_, N57, N61 );
nand g282 ( new_n420_, new_n416_, new_n418_, new_n417_, new_n419_ );
nand g283 ( new_n421_, new_n416_, new_n417_ );
nand g284 ( new_n422_, new_n418_, new_n419_ );
nand g285 ( new_n423_, new_n421_, new_n422_ );
nand g286 ( new_n424_, new_n423_, new_n420_ );
nand g287 ( new_n425_, new_n415_, new_n424_ );
not g288 ( new_n426_, new_n424_ );
nand g289 ( new_n427_, new_n412_, new_n414_, new_n426_ );
nand g290 ( new_n428_, new_n425_, N136, N137, new_n427_ );
nand g291 ( new_n429_, new_n425_, new_n427_ );
nand g292 ( new_n430_, N136, N137 );
nand g293 ( new_n431_, new_n429_, new_n430_ );
nand g294 ( new_n432_, new_n143_, N77 );
nand g295 ( new_n433_, new_n157_, N93 );
nand g296 ( new_n434_, new_n296_, new_n309_ );
nand g297 ( new_n435_, N109, N125 );
nand g298 ( new_n436_, new_n434_, new_n432_, new_n433_, new_n435_ );
nand g299 ( new_n437_, new_n432_, new_n433_ );
nand g300 ( new_n438_, new_n434_, new_n435_ );
nand g301 ( new_n439_, new_n437_, new_n438_ );
nand g302 ( new_n440_, new_n431_, new_n428_, new_n436_, new_n439_ );
nand g303 ( new_n441_, new_n431_, new_n428_ );
nand g304 ( new_n442_, new_n439_, new_n436_ );
nand g305 ( new_n443_, new_n441_, new_n442_ );
nand g306 ( new_n444_, new_n443_, new_n440_ );
nand g307 ( new_n445_, new_n287_, new_n394_, new_n444_ );
nand g308 ( new_n446_, new_n415_, new_n210_, new_n213_ );
nand g309 ( new_n447_, new_n238_, new_n412_, new_n414_ );
nand g310 ( new_n448_, new_n447_, new_n446_ );
nand g311 ( new_n449_, new_n448_, keyIn_0_18 );
not g312 ( new_n450_, keyIn_0_18 );
nand g313 ( new_n451_, new_n447_, new_n450_, new_n446_ );
nand g314 ( new_n452_, new_n449_, new_n451_ );
nand g315 ( new_n453_, keyIn_0_6, N133, N137 );
not g316 ( new_n454_, keyIn_0_6 );
nand g317 ( new_n455_, N133, N137 );
nand g318 ( new_n456_, new_n455_, new_n454_ );
nand g319 ( new_n457_, new_n456_, new_n453_ );
nand g320 ( new_n458_, new_n452_, new_n457_ );
nand g321 ( new_n459_, new_n449_, new_n451_, new_n453_, new_n456_ );
nand g322 ( new_n460_, new_n458_, new_n459_ );
nand g323 ( new_n461_, new_n460_, keyIn_0_20 );
not g324 ( new_n462_, keyIn_0_20 );
nand g325 ( new_n463_, new_n458_, new_n462_, new_n459_ );
nand g326 ( new_n464_, new_n461_, new_n463_ );
not g327 ( new_n465_, keyIn_0_16 );
nor g328 ( new_n466_, N97, N113 );
not g329 ( new_n467_, new_n466_ );
nand g330 ( new_n468_, N97, N113 );
nand g331 ( new_n469_, new_n467_, new_n468_ );
nor g332 ( new_n470_, new_n469_, keyIn_0_9 );
nand g333 ( new_n471_, new_n469_, keyIn_0_9 );
not g334 ( new_n472_, new_n471_ );
nor g335 ( new_n473_, new_n472_, new_n470_ );
nand g336 ( new_n474_, new_n140_, N65 );
nand g337 ( new_n475_, new_n154_, N81 );
nand g338 ( new_n476_, new_n474_, new_n475_ );
nand g339 ( new_n477_, new_n476_, keyIn_0_8 );
not g340 ( new_n478_, keyIn_0_8 );
nand g341 ( new_n479_, new_n474_, new_n475_, new_n478_ );
nand g342 ( new_n480_, new_n473_, new_n477_, new_n479_ );
not g343 ( new_n481_, new_n473_ );
nand g344 ( new_n482_, new_n477_, new_n479_ );
nand g345 ( new_n483_, new_n481_, new_n482_ );
nand g346 ( new_n484_, new_n483_, new_n465_, new_n480_ );
nand g347 ( new_n485_, new_n483_, new_n480_ );
nand g348 ( new_n486_, new_n485_, keyIn_0_16 );
nand g349 ( new_n487_, new_n486_, new_n484_ );
nand g350 ( new_n488_, new_n464_, new_n487_ );
nand g351 ( new_n489_, new_n461_, new_n463_, new_n484_, new_n486_ );
nand g352 ( new_n490_, new_n488_, keyIn_0_22, new_n489_ );
not g353 ( new_n491_, keyIn_0_22 );
nand g354 ( new_n492_, new_n488_, new_n489_ );
nand g355 ( new_n493_, new_n492_, new_n491_ );
nand g356 ( new_n494_, new_n493_, new_n490_ );
not g357 ( new_n495_, new_n494_ );
nand g358 ( new_n496_, new_n239_, new_n424_ );
nand g359 ( new_n497_, new_n235_, new_n236_, new_n426_ );
nand g360 ( new_n498_, new_n496_, N134, N137, new_n497_ );
nand g361 ( new_n499_, new_n496_, new_n497_ );
nand g362 ( new_n500_, N134, N137 );
nand g363 ( new_n501_, new_n499_, new_n500_ );
nand g364 ( new_n502_, new_n138_, N69 );
nand g365 ( new_n503_, new_n152_, N85 );
nand g366 ( new_n504_, new_n292_, new_n305_ );
nand g367 ( new_n505_, N101, N117 );
nand g368 ( new_n506_, new_n504_, new_n502_, new_n503_, new_n505_ );
nand g369 ( new_n507_, new_n502_, new_n503_ );
nand g370 ( new_n508_, new_n504_, new_n505_ );
nand g371 ( new_n509_, new_n507_, new_n508_ );
nand g372 ( new_n510_, new_n501_, new_n498_, new_n506_, new_n509_ );
nand g373 ( new_n511_, new_n501_, new_n498_ );
nand g374 ( new_n512_, new_n509_, new_n506_ );
nand g375 ( new_n513_, new_n511_, new_n512_ );
nand g376 ( new_n514_, new_n513_, new_n510_ );
nand g377 ( new_n515_, new_n495_, new_n514_ );
nor g378 ( new_n516_, new_n445_, new_n515_ );
not g379 ( new_n517_, new_n516_ );
nor g380 ( new_n518_, new_n517_, new_n188_ );
not g381 ( new_n519_, new_n518_ );
nand g382 ( new_n520_, new_n519_, N1 );
nand g383 ( new_n521_, new_n518_, new_n174_ );
nand g384 ( N724, new_n520_, new_n521_ );
nor g385 ( new_n523_, new_n517_, new_n338_ );
not g386 ( new_n524_, new_n523_ );
nand g387 ( new_n525_, new_n524_, N5 );
nand g388 ( new_n526_, new_n523_, new_n199_ );
nand g389 ( N725, new_n525_, new_n526_ );
nor g390 ( new_n528_, new_n517_, new_n359_ );
not g391 ( new_n529_, new_n528_ );
nand g392 ( new_n530_, new_n529_, N9 );
nand g393 ( new_n531_, new_n528_, new_n191_ );
nand g394 ( N726, new_n530_, new_n531_ );
nor g395 ( new_n533_, new_n517_, new_n390_ );
not g396 ( new_n534_, new_n533_ );
nand g397 ( new_n535_, new_n534_, N13 );
nand g398 ( new_n536_, new_n533_, new_n192_ );
nand g399 ( N727, new_n535_, new_n536_ );
not g400 ( new_n538_, new_n444_ );
nand g401 ( new_n539_, new_n286_, new_n394_, new_n538_ );
nor g402 ( new_n540_, new_n515_, new_n539_ );
not g403 ( new_n541_, new_n540_ );
nor g404 ( new_n542_, new_n541_, new_n188_ );
not g405 ( new_n543_, new_n542_ );
nand g406 ( new_n544_, new_n543_, N17 );
nand g407 ( new_n545_, new_n542_, new_n172_ );
nand g408 ( N728, new_n544_, new_n545_ );
nor g409 ( new_n547_, new_n541_, new_n338_ );
not g410 ( new_n548_, new_n547_ );
nand g411 ( new_n549_, new_n548_, N21 );
nand g412 ( new_n550_, new_n547_, new_n324_ );
nand g413 ( N729, new_n549_, new_n550_ );
nor g414 ( new_n552_, new_n541_, new_n359_ );
not g415 ( new_n553_, new_n552_ );
nand g416 ( new_n554_, new_n553_, N25 );
nand g417 ( new_n555_, new_n552_, new_n345_ );
nand g418 ( N730, new_n554_, new_n555_ );
nor g419 ( new_n557_, new_n541_, new_n390_ );
not g420 ( new_n558_, new_n557_ );
nand g421 ( new_n559_, new_n558_, N29 );
nand g422 ( new_n560_, new_n557_, new_n373_ );
nand g423 ( N731, new_n559_, new_n560_ );
not g424 ( new_n562_, new_n514_ );
nand g425 ( new_n563_, new_n494_, new_n562_ );
nor g426 ( new_n564_, new_n445_, new_n563_ );
not g427 ( new_n565_, new_n564_ );
nor g428 ( new_n566_, new_n565_, new_n188_ );
not g429 ( new_n567_, new_n566_ );
nand g430 ( new_n568_, new_n567_, N33 );
nand g431 ( new_n569_, new_n566_, new_n176_ );
nand g432 ( N732, new_n568_, new_n569_ );
nor g433 ( new_n571_, new_n565_, new_n338_ );
not g434 ( new_n572_, new_n571_ );
nand g435 ( new_n573_, new_n572_, N37 );
nand g436 ( new_n574_, new_n571_, new_n224_ );
nand g437 ( N733, new_n573_, new_n574_ );
nor g438 ( new_n576_, new_n565_, new_n359_ );
not g439 ( new_n577_, new_n576_ );
nand g440 ( new_n578_, new_n577_, N41 );
nand g441 ( new_n579_, new_n576_, new_n215_ );
nand g442 ( N734, new_n578_, new_n579_ );
nor g443 ( new_n581_, new_n565_, new_n390_ );
not g444 ( new_n582_, new_n581_ );
nand g445 ( new_n583_, new_n582_, N45 );
nand g446 ( new_n584_, new_n581_, new_n216_ );
nand g447 ( N735, new_n583_, new_n584_ );
nor g448 ( new_n586_, new_n563_, new_n539_ );
not g449 ( new_n587_, new_n586_ );
nor g450 ( new_n588_, new_n587_, new_n188_ );
not g451 ( new_n589_, new_n588_ );
nand g452 ( new_n590_, new_n589_, N49 );
nand g453 ( new_n591_, new_n588_, new_n177_ );
nand g454 ( N736, new_n590_, new_n591_ );
nor g455 ( new_n593_, new_n587_, new_n338_ );
not g456 ( new_n594_, new_n593_ );
nand g457 ( new_n595_, new_n594_, N53 );
nand g458 ( new_n596_, new_n593_, new_n327_ );
nand g459 ( N737, new_n595_, new_n596_ );
nor g460 ( new_n598_, new_n587_, new_n359_ );
not g461 ( new_n599_, new_n598_ );
nand g462 ( new_n600_, new_n599_, N57 );
nand g463 ( new_n601_, new_n598_, new_n348_ );
nand g464 ( N738, new_n600_, new_n601_ );
nor g465 ( new_n603_, new_n587_, new_n390_ );
not g466 ( new_n604_, new_n603_ );
nand g467 ( new_n605_, new_n604_, N61 );
nand g468 ( new_n606_, new_n603_, new_n376_ );
nand g469 ( N739, new_n605_, new_n606_ );
not g470 ( new_n608_, keyIn_0_52 );
not g471 ( new_n609_, keyIn_0_37 );
not g472 ( new_n610_, keyIn_0_36 );
not g473 ( new_n611_, keyIn_0_27 );
nand g474 ( new_n612_, new_n286_, new_n611_ );
nand g475 ( new_n613_, new_n285_, keyIn_0_27, new_n283_ );
nand g476 ( new_n614_, new_n612_, new_n613_ );
not g477 ( new_n615_, keyIn_0_25 );
nand g478 ( new_n616_, new_n495_, new_n615_ );
nand g479 ( new_n617_, new_n494_, keyIn_0_25 );
not g480 ( new_n618_, keyIn_0_26 );
nand g481 ( new_n619_, new_n514_, new_n618_ );
not g482 ( new_n620_, new_n619_ );
nand g483 ( new_n621_, new_n562_, keyIn_0_26 );
not g484 ( new_n622_, new_n621_ );
nor g485 ( new_n623_, new_n622_, new_n444_, new_n620_ );
nand g486 ( new_n624_, new_n616_, new_n614_, new_n617_, new_n623_ );
nand g487 ( new_n625_, new_n624_, keyIn_0_32 );
not g488 ( new_n626_, keyIn_0_32 );
nand g489 ( new_n627_, new_n617_, new_n623_ );
not g490 ( new_n628_, new_n627_ );
nand g491 ( new_n629_, new_n628_, new_n626_, new_n614_, new_n616_ );
nand g492 ( new_n630_, new_n625_, new_n629_ );
not g493 ( new_n631_, keyIn_0_31 );
nand g494 ( new_n632_, new_n285_, new_n631_, new_n283_ );
nand g495 ( new_n633_, new_n286_, keyIn_0_31 );
nand g496 ( new_n634_, new_n633_, new_n632_ );
nand g497 ( new_n635_, new_n493_, new_n444_, new_n490_, new_n514_ );
not g498 ( new_n636_, new_n635_ );
nand g499 ( new_n637_, new_n634_, new_n636_ );
nand g500 ( new_n638_, new_n637_, keyIn_0_35 );
not g501 ( new_n639_, keyIn_0_35 );
nand g502 ( new_n640_, new_n634_, new_n639_, new_n636_ );
nand g503 ( new_n641_, new_n638_, new_n640_ );
not g504 ( new_n642_, keyIn_0_33 );
not g505 ( new_n643_, keyIn_0_28 );
nand g506 ( new_n644_, new_n494_, new_n643_ );
nand g507 ( new_n645_, new_n493_, keyIn_0_28, new_n490_ );
nand g508 ( new_n646_, new_n285_, new_n283_, new_n444_, new_n514_ );
not g509 ( new_n647_, new_n646_ );
nand g510 ( new_n648_, new_n644_, new_n647_, new_n645_ );
nand g511 ( new_n649_, new_n648_, new_n642_ );
nand g512 ( new_n650_, new_n644_, new_n647_, keyIn_0_33, new_n645_ );
nand g513 ( new_n651_, new_n649_, new_n650_ );
nand g514 ( new_n652_, new_n641_, new_n651_ );
not g515 ( new_n653_, new_n652_ );
nand g516 ( new_n654_, new_n494_, keyIn_0_29 );
not g517 ( new_n655_, keyIn_0_29 );
nand g518 ( new_n656_, new_n493_, new_n655_, new_n490_ );
nand g519 ( new_n657_, new_n654_, new_n656_ );
not g520 ( new_n658_, keyIn_0_30 );
nand g521 ( new_n659_, new_n286_, new_n658_ );
nand g522 ( new_n660_, new_n285_, keyIn_0_30, new_n283_ );
nor g523 ( new_n661_, new_n538_, new_n514_ );
nand g524 ( new_n662_, new_n660_, new_n661_ );
not g525 ( new_n663_, new_n662_ );
nand g526 ( new_n664_, new_n657_, new_n663_, keyIn_0_34, new_n659_ );
not g527 ( new_n665_, keyIn_0_34 );
nand g528 ( new_n666_, new_n657_, new_n659_, new_n663_ );
nand g529 ( new_n667_, new_n666_, new_n665_ );
nand g530 ( new_n668_, new_n667_, new_n664_ );
not g531 ( new_n669_, new_n668_ );
nand g532 ( new_n670_, new_n653_, new_n610_, new_n630_, new_n669_ );
nand g533 ( new_n671_, new_n669_, new_n630_, new_n641_, new_n651_ );
nand g534 ( new_n672_, new_n671_, keyIn_0_36 );
nand g535 ( new_n673_, new_n672_, new_n670_ );
nand g536 ( new_n674_, new_n360_, new_n390_ );
nor g537 ( new_n675_, new_n674_, new_n188_, new_n363_ );
nand g538 ( new_n676_, new_n673_, new_n609_, new_n675_ );
nand g539 ( new_n677_, new_n673_, new_n675_ );
nand g540 ( new_n678_, new_n677_, keyIn_0_37 );
nand g541 ( new_n679_, new_n678_, new_n676_ );
nand g542 ( new_n680_, new_n679_, new_n495_ );
nand g543 ( new_n681_, new_n680_, keyIn_0_40 );
not g544 ( new_n682_, keyIn_0_40 );
nand g545 ( new_n683_, new_n679_, new_n682_, new_n495_ );
nand g546 ( new_n684_, new_n681_, new_n683_ );
nand g547 ( new_n685_, new_n684_, N65 );
nand g548 ( new_n686_, new_n681_, new_n154_, new_n683_ );
nand g549 ( new_n687_, new_n685_, new_n686_ );
nand g550 ( new_n688_, new_n687_, new_n608_ );
nand g551 ( new_n689_, new_n685_, keyIn_0_52, new_n686_ );
nand g552 ( N740, new_n688_, new_n689_ );
not g553 ( new_n691_, keyIn_0_53 );
not g554 ( new_n692_, keyIn_0_41 );
nand g555 ( new_n693_, new_n679_, new_n562_ );
nand g556 ( new_n694_, new_n693_, new_n692_ );
nand g557 ( new_n695_, new_n679_, keyIn_0_41, new_n562_ );
nand g558 ( new_n696_, new_n694_, new_n695_ );
nand g559 ( new_n697_, new_n696_, new_n152_ );
nand g560 ( new_n698_, new_n694_, N69, new_n695_ );
nand g561 ( new_n699_, new_n697_, new_n698_ );
nand g562 ( new_n700_, new_n699_, new_n691_ );
nand g563 ( new_n701_, new_n697_, keyIn_0_53, new_n698_ );
nand g564 ( N741, new_n700_, new_n701_ );
nand g565 ( new_n703_, new_n679_, new_n287_ );
nand g566 ( new_n704_, new_n703_, keyIn_0_42 );
not g567 ( new_n705_, keyIn_0_42 );
nand g568 ( new_n706_, new_n679_, new_n705_, new_n287_ );
nand g569 ( new_n707_, new_n704_, new_n706_ );
nand g570 ( new_n708_, new_n707_, new_n156_ );
nand g571 ( new_n709_, new_n704_, N73, new_n706_ );
nand g572 ( new_n710_, new_n708_, new_n709_ );
nand g573 ( new_n711_, new_n710_, keyIn_0_54 );
not g574 ( new_n712_, keyIn_0_54 );
nand g575 ( new_n713_, new_n708_, new_n712_, new_n709_ );
nand g576 ( N742, new_n711_, new_n713_ );
not g577 ( new_n715_, keyIn_0_55 );
nand g578 ( new_n716_, new_n679_, new_n538_ );
nand g579 ( new_n717_, new_n716_, keyIn_0_43 );
not g580 ( new_n718_, keyIn_0_43 );
nand g581 ( new_n719_, new_n679_, new_n718_, new_n538_ );
nand g582 ( new_n720_, new_n717_, new_n719_ );
nand g583 ( new_n721_, new_n720_, N77 );
nand g584 ( new_n722_, new_n717_, new_n157_, new_n719_ );
nand g585 ( new_n723_, new_n721_, new_n722_ );
nand g586 ( new_n724_, new_n723_, new_n715_ );
nand g587 ( new_n725_, new_n721_, keyIn_0_55, new_n722_ );
nand g588 ( N743, new_n724_, new_n725_ );
not g589 ( new_n727_, keyIn_0_44 );
nor g590 ( new_n728_, new_n362_, new_n390_ );
nand g591 ( new_n729_, new_n673_, new_n728_ );
nand g592 ( new_n730_, new_n729_, keyIn_0_38 );
not g593 ( new_n731_, keyIn_0_38 );
nand g594 ( new_n732_, new_n673_, new_n731_, new_n728_ );
nand g595 ( new_n733_, new_n730_, new_n495_, new_n732_ );
nand g596 ( new_n734_, new_n733_, new_n727_ );
nand g597 ( new_n735_, new_n730_, keyIn_0_44, new_n495_, new_n732_ );
nand g598 ( new_n736_, new_n734_, new_n735_ );
nand g599 ( new_n737_, new_n736_, new_n140_ );
nand g600 ( new_n738_, new_n734_, N81, new_n735_ );
nand g601 ( new_n739_, new_n737_, new_n738_ );
nand g602 ( new_n740_, new_n739_, keyIn_0_56 );
not g603 ( new_n741_, keyIn_0_56 );
nand g604 ( new_n742_, new_n737_, new_n741_, new_n738_ );
nand g605 ( N744, new_n740_, new_n742_ );
not g606 ( new_n744_, keyIn_0_57 );
nand g607 ( new_n745_, new_n730_, new_n562_, new_n732_ );
nand g608 ( new_n746_, new_n745_, keyIn_0_45 );
not g609 ( new_n747_, keyIn_0_45 );
nand g610 ( new_n748_, new_n730_, new_n747_, new_n562_, new_n732_ );
nand g611 ( new_n749_, new_n746_, new_n748_ );
nand g612 ( new_n750_, new_n749_, N85 );
nand g613 ( new_n751_, new_n746_, new_n138_, new_n748_ );
nand g614 ( new_n752_, new_n750_, new_n751_ );
nand g615 ( new_n753_, new_n752_, new_n744_ );
nand g616 ( new_n754_, new_n750_, keyIn_0_57, new_n751_ );
nand g617 ( N745, new_n753_, new_n754_ );
nand g618 ( new_n756_, new_n730_, new_n287_, new_n732_ );
nand g619 ( new_n757_, new_n756_, keyIn_0_46 );
not g620 ( new_n758_, keyIn_0_46 );
nand g621 ( new_n759_, new_n730_, new_n758_, new_n287_, new_n732_ );
nand g622 ( new_n760_, new_n757_, new_n759_ );
nand g623 ( new_n761_, new_n760_, N89 );
nand g624 ( new_n762_, new_n757_, new_n142_, new_n759_ );
nand g625 ( new_n763_, new_n761_, new_n762_ );
nand g626 ( new_n764_, new_n763_, keyIn_0_58 );
not g627 ( new_n765_, keyIn_0_58 );
nand g628 ( new_n766_, new_n761_, new_n765_, new_n762_ );
nand g629 ( N746, new_n764_, new_n766_ );
not g630 ( new_n768_, keyIn_0_59 );
nand g631 ( new_n769_, new_n730_, new_n538_, new_n732_ );
nand g632 ( new_n770_, new_n769_, keyIn_0_47 );
not g633 ( new_n771_, keyIn_0_47 );
nand g634 ( new_n772_, new_n730_, new_n771_, new_n538_, new_n732_ );
nand g635 ( new_n773_, new_n770_, new_n772_ );
nand g636 ( new_n774_, new_n773_, N93 );
nand g637 ( new_n775_, new_n770_, new_n143_, new_n772_ );
nand g638 ( new_n776_, new_n774_, new_n775_ );
nand g639 ( new_n777_, new_n776_, new_n768_ );
nand g640 ( new_n778_, new_n774_, keyIn_0_59, new_n775_ );
nand g641 ( N747, new_n777_, new_n778_ );
not g642 ( new_n780_, keyIn_0_39 );
nor g643 ( new_n781_, new_n674_, new_n290_, new_n338_ );
nand g644 ( new_n782_, new_n673_, new_n780_, new_n781_ );
nand g645 ( new_n783_, new_n673_, new_n781_ );
nand g646 ( new_n784_, new_n783_, keyIn_0_39 );
nand g647 ( new_n785_, new_n784_, new_n782_ );
nand g648 ( new_n786_, new_n785_, new_n495_ );
nand g649 ( new_n787_, new_n786_, keyIn_0_48 );
not g650 ( new_n788_, keyIn_0_48 );
nand g651 ( new_n789_, new_n785_, new_n788_, new_n495_ );
nand g652 ( new_n790_, new_n787_, new_n789_ );
nand g653 ( new_n791_, new_n790_, N97 );
nand g654 ( new_n792_, new_n787_, new_n294_, new_n789_ );
nand g655 ( new_n793_, new_n791_, new_n792_ );
nand g656 ( new_n794_, new_n793_, keyIn_0_60 );
not g657 ( new_n795_, keyIn_0_60 );
nand g658 ( new_n796_, new_n791_, new_n795_, new_n792_ );
nand g659 ( N748, new_n794_, new_n796_ );
not g660 ( new_n798_, keyIn_0_49 );
nand g661 ( new_n799_, new_n785_, new_n562_ );
nand g662 ( new_n800_, new_n799_, new_n798_ );
nand g663 ( new_n801_, new_n785_, keyIn_0_49, new_n562_ );
nand g664 ( new_n802_, new_n800_, new_n801_ );
nand g665 ( new_n803_, new_n802_, new_n292_ );
nand g666 ( new_n804_, new_n800_, N101, new_n801_ );
nand g667 ( new_n805_, new_n803_, new_n804_ );
nand g668 ( new_n806_, new_n805_, keyIn_0_61 );
not g669 ( new_n807_, keyIn_0_61 );
nand g670 ( new_n808_, new_n803_, new_n807_, new_n804_ );
nand g671 ( N749, new_n806_, new_n808_ );
not g672 ( new_n810_, keyIn_0_50 );
nand g673 ( new_n811_, new_n785_, new_n287_ );
nand g674 ( new_n812_, new_n811_, new_n810_ );
nand g675 ( new_n813_, new_n785_, keyIn_0_50, new_n287_ );
nand g676 ( new_n814_, new_n812_, new_n813_ );
nand g677 ( new_n815_, new_n814_, new_n266_ );
nand g678 ( new_n816_, new_n812_, N105, new_n813_ );
nand g679 ( new_n817_, new_n815_, new_n816_ );
nand g680 ( new_n818_, new_n817_, keyIn_0_62 );
not g681 ( new_n819_, keyIn_0_62 );
nand g682 ( new_n820_, new_n815_, new_n819_, new_n816_ );
nand g683 ( N750, new_n818_, new_n820_ );
not g684 ( new_n822_, keyIn_0_63 );
nand g685 ( new_n823_, new_n785_, new_n538_ );
nand g686 ( new_n824_, new_n823_, keyIn_0_51 );
not g687 ( new_n825_, keyIn_0_51 );
nand g688 ( new_n826_, new_n785_, new_n825_, new_n538_ );
nand g689 ( new_n827_, new_n824_, new_n826_ );
nand g690 ( new_n828_, new_n827_, new_n296_ );
nand g691 ( new_n829_, new_n824_, N109, new_n826_ );
nand g692 ( new_n830_, new_n828_, new_n829_ );
nand g693 ( new_n831_, new_n830_, new_n822_ );
nand g694 ( new_n832_, new_n828_, keyIn_0_63, new_n829_ );
nand g695 ( N751, new_n831_, new_n832_ );
not g696 ( new_n834_, new_n673_ );
nor g697 ( new_n835_, new_n834_, new_n364_, new_n390_ );
nand g698 ( new_n836_, new_n835_, new_n495_ );
nand g699 ( new_n837_, new_n836_, N113 );
nand g700 ( new_n838_, new_n835_, new_n307_, new_n495_ );
nand g701 ( N752, new_n837_, new_n838_ );
nand g702 ( new_n840_, new_n835_, new_n562_ );
nand g703 ( new_n841_, new_n840_, N117 );
nand g704 ( new_n842_, new_n835_, new_n305_, new_n562_ );
nand g705 ( N753, new_n841_, new_n842_ );
nand g706 ( new_n844_, new_n835_, new_n287_ );
nand g707 ( new_n845_, new_n844_, N121 );
nand g708 ( new_n846_, new_n835_, new_n264_, new_n287_ );
nand g709 ( N754, new_n845_, new_n846_ );
nand g710 ( new_n848_, new_n835_, new_n538_ );
nand g711 ( new_n849_, new_n848_, N125 );
nand g712 ( new_n850_, new_n835_, new_n309_, new_n538_ );
nand g713 ( N755, new_n849_, new_n850_ );
endmodule