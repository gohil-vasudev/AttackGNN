module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n1668_, new_n1359_, new_n595_, new_n1233_, new_n445_, new_n1009_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n501_, new_n1157_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1433_, new_n1517_, new_n1575_, new_n1472_, new_n1048_, new_n885_, new_n439_, new_n1532_, new_n390_, new_n743_, new_n1327_, new_n1535_, new_n566_, new_n641_, new_n386_, new_n767_, new_n401_, new_n514_, new_n1351_, new_n556_, new_n636_, new_n691_, new_n1024_, new_n670_, new_n456_, new_n1125_, new_n1590_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n1568_, new_n728_, new_n1071_, new_n1294_, new_n894_, new_n853_, new_n695_, new_n660_, new_n1311_, new_n526_, new_n908_, new_n552_, new_n678_, new_n1662_, new_n706_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n1188_, new_n1415_, new_n1390_, new_n721_, new_n504_, new_n1414_, new_n742_, new_n892_, new_n1368_, new_n472_, new_n873_, new_n1167_, new_n1530_, new_n1300_, new_n1490_, new_n774_, new_n792_, new_n1620_, new_n953_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n1580_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n1447_, new_n635_, new_n685_, new_n648_, new_n903_, new_n1595_, new_n983_, new_n822_, new_n1406_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n1054_, new_n655_, new_n1288_, new_n630_, new_n1717_, new_n385_, new_n1670_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n565_, new_n1196_, new_n1366_, new_n511_, new_n1714_, new_n1640_, new_n1285_, new_n1031_, new_n1733_, new_n1216_, new_n1632_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n1647_, new_n1713_, new_n960_, new_n1377_, new_n1522_, new_n549_, new_n491_, new_n676_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n1678_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n1463_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1424_, new_n1062_, new_n680_, new_n981_, new_n506_, new_n872_, new_n1527_, new_n1275_, new_n1277_, new_n1198_, new_n1428_, new_n1440_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n483_, new_n1004_, new_n1152_, new_n1558_, new_n394_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1735_, new_n1113_, new_n785_, new_n1501_, new_n441_, new_n477_, new_n664_, new_n600_, new_n1737_, new_n1041_, new_n1657_, new_n1562_, new_n426_, new_n1036_, new_n398_, new_n1576_, new_n1718_, new_n1333_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n1740_, new_n1395_, new_n473_, new_n1624_, new_n1147_, new_n1682_, new_n1373_, new_n1229_, new_n1422_, new_n1523_, new_n1698_, new_n1468_, new_n1679_, new_n969_, new_n835_, new_n1234_, new_n1360_, new_n378_, new_n1574_, new_n1614_, new_n621_, new_n1423_, new_n1637_, new_n1732_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1321_, new_n1690_, new_n1209_, new_n1709_, new_n347_, new_n659_, new_n700_, new_n1419_, new_n921_, new_n396_, new_n1315_, new_n1003_, new_n696_, new_n1039_, new_n1507_, new_n1439_, new_n1658_, new_n1671_, new_n1239_, new_n1365_, new_n528_, new_n952_, new_n1158_, new_n1667_, new_n729_, new_n1111_, new_n1413_, new_n1218_, new_n1385_, new_n1346_, new_n1201_, new_n559_, new_n1282_, new_n1630_, new_n762_, new_n1349_, new_n1193_, new_n1547_, new_n1437_, new_n1598_, new_n1187_, new_n1205_, new_n1154_, new_n1253_, new_n1546_, new_n1453_, new_n1256_, new_n628_, new_n1513_, new_n409_, new_n1090_, new_n1669_, new_n1489_, new_n553_, new_n745_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n834_, new_n1573_, new_n1738_, new_n1693_, new_n1171_, new_n867_, new_n954_, new_n1591_, new_n1626_, new_n1032_, new_n1545_, new_n901_, new_n688_, new_n1255_, new_n1704_, new_n410_, new_n985_, new_n851_, new_n1518_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n1712_, new_n509_, new_n661_, new_n797_, new_n1358_, new_n724_, new_n1070_, new_n1686_, new_n1416_, new_n1109_, new_n1496_, new_n672_, new_n1269_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n1600_, new_n1592_, new_n809_, new_n1631_, new_n1142_, new_n1623_, new_n604_, new_n1461_, new_n1104_, new_n1703_, new_n1511_, new_n571_, new_n1504_, new_n758_, new_n460_, new_n1267_, new_n1705_, new_n1466_, new_n1707_, new_n1716_, new_n1516_, new_n1299_, new_n1477_, new_n1079_, new_n861_, new_n1564_, new_n1656_, new_n1252_, new_n352_, new_n1553_, new_n1493_, new_n575_, new_n562_, new_n1593_, new_n944_, new_n1638_, new_n1542_, new_n1064_, new_n1065_, new_n1118_, new_n1645_, new_n493_, new_n547_, new_n1480_, new_n379_, new_n963_, new_n586_, new_n1481_, new_n1325_, new_n993_, new_n1625_, new_n1357_, new_n1191_, new_n824_, new_n1628_, new_n717_, new_n1455_, new_n403_, new_n868_, new_n1242_, new_n475_, new_n858_, new_n1612_, new_n1384_, new_n1343_, new_n936_, new_n1459_, new_n1434_, new_n1438_, new_n1016_, new_n411_, new_n673_, new_n1144_, new_n1465_, new_n666_, new_n1290_, new_n407_, new_n1519_, new_n1407_, new_n1692_, new_n1726_, new_n879_, new_n1417_, new_n1700_, new_n736_, new_n513_, new_n558_, new_n382_, new_n1370_, new_n718_, new_n1310_, new_n1710_, new_n1398_, new_n1126_, new_n546_, new_n612_, new_n1015_, new_n919_, new_n755_, new_n1040_, new_n1635_, new_n1509_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n345_, new_n499_, new_n533_, new_n1130_, new_n795_, new_n459_, new_n1441_, new_n1122_, new_n1728_, new_n1185_, new_n1240_, new_n1510_, new_n1174_, new_n968_, new_n1655_, new_n1464_, new_n613_, new_n1508_, new_n1195_, new_n417_, new_n658_, new_n837_, new_n591_, new_n801_, new_n1458_, new_n631_, new_n453_, new_n1723_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1521_, new_n1334_, new_n531_, new_n1675_, new_n593_, new_n1543_, new_n974_, new_n1565_, new_n1248_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n1454_, new_n1474_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n1430_, new_n470_, new_n769_, new_n1660_, new_n433_, new_n871_, new_n1450_, new_n992_, new_n1098_, new_n1729_, new_n732_, new_n689_, new_n933_, new_n584_, new_n815_, new_n1608_, new_n1492_, new_n1367_, new_n1619_, new_n1052_, new_n1425_, new_n857_, new_n1379_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n1471_, new_n1673_, new_n1220_, new_n989_, new_n1741_, new_n1117_, new_n1421_, new_n644_, new_n1594_, new_n836_, new_n1116_, new_n1684_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n913_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n1427_, new_n818_, new_n881_, new_n1268_, new_n1376_, new_n1381_, new_n1566_, new_n1534_, new_n684_, new_n640_, new_n1274_, new_n1665_, new_n754_, new_n653_, new_n1659_, new_n905_, new_n377_, new_n1258_, new_n1539_, new_n1643_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1391_, new_n1724_, new_n1436_, new_n567_, new_n1353_, new_n1033_, new_n576_, new_n831_, new_n791_, new_n1153_, new_n357_, new_n1339_, new_n984_, new_n780_, new_n1183_, new_n643_, new_n1316_, new_n1194_, new_n1338_, new_n1460_, new_n1230_, new_n1602_, new_n1027_, new_n610_, new_n1369_, new_n1694_, new_n843_, new_n703_, new_n698_, new_n1639_, new_n1165_, new_n1259_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1066_, new_n422_, new_n581_, new_n1664_, new_n686_, new_n934_, new_n1567_, new_n1651_, new_n770_, new_n1389_, new_n1400_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n1597_, new_n356_, new_n647_, new_n889_, new_n536_, new_n1616_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n1405_, new_n1249_, new_n1354_, new_n955_, new_n847_, new_n888_, new_n1505_, new_n1340_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1361_, new_n941_, new_n1410_, new_n738_, new_n827_, new_n1356_, new_n1363_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n1211_, new_n1412_, new_n1207_, new_n1176_, new_n1374_, new_n601_, new_n842_, new_n1552_, new_n1057_, new_n1644_, new_n1677_, new_n682_, new_n1075_, new_n812_, new_n1563_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1397_, new_n1402_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n1603_, new_n451_, new_n489_, new_n804_, new_n1342_, new_n424_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n413_, new_n1544_, new_n1382_, new_n442_, new_n677_, new_n1487_, new_n1646_, new_n642_, new_n1418_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n761_, new_n840_, new_n735_, new_n1283_, new_n898_, new_n1734_, new_n799_, new_n1304_, new_n1537_, new_n946_, new_n1108_, new_n1469_, new_n862_, new_n1606_, new_n427_, new_n532_, new_n1739_, new_n1617_, new_n418_, new_n746_, new_n1221_, new_n1585_, new_n1587_, new_n1264_, new_n1319_, new_n626_, new_n1680_, new_n1473_, new_n959_, new_n990_, new_n1629_, new_n716_, new_n701_, new_n1238_, new_n1676_, new_n1058_, new_n1162_, new_n1730_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n1696_, new_n414_, new_n1101_, new_n1250_, new_n1681_, new_n1482_, new_n1050_, new_n554_, new_n1151_, new_n844_, new_n1302_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n589_, new_n1083_, new_n759_, new_n1297_, new_n829_, new_n1257_, new_n1306_, new_n1720_, new_n988_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n1486_, new_n764_, new_n906_, new_n683_, new_n1409_, new_n1429_, new_n463_, new_n1683_, new_n1372_, new_n510_, new_n966_, new_n1685_, new_n1721_, new_n351_, new_n1184_, new_n1292_, new_n1426_, new_n517_, new_n609_, new_n961_, new_n530_, new_n890_, new_n1006_, new_n622_, new_n1706_, new_n702_, new_n833_, new_n1560_, new_n1701_, new_n715_, new_n811_, new_n1445_, new_n1371_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1622_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n1618_, new_n1652_, new_n1170_, new_n845_, new_n768_, new_n1691_, new_n773_, new_n1452_, new_n1051_, new_n899_, new_n1053_, new_n1540_, new_n1611_, new_n1708_, new_n492_, new_n1200_, new_n1533_, new_n650_, new_n750_, new_n887_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n1226_, new_n778_, new_n452_, new_n1727_, new_n381_, new_n1483_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n820_, new_n1386_, new_n771_, new_n979_, new_n508_, new_n1435_, new_n714_, new_n1280_, new_n1007_, new_n1613_, new_n1241_, new_n882_, new_n1145_, new_n1557_, new_n929_, new_n986_, new_n1159_, new_n1584_, new_n1337_, new_n1348_, new_n917_, new_n1555_, new_n1636_, new_n1322_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n541_, new_n447_, new_n1388_, new_n1550_, new_n790_, new_n1081_, new_n587_, new_n1247_, new_n1411_, new_n465_, new_n783_, new_n1380_, new_n739_, new_n996_, new_n1601_, new_n1318_, new_n846_, new_n915_, new_n488_, new_n524_, new_n349_, new_n848_, new_n1725_, new_n1245_, new_n663_, new_n1499_, new_n1497_, new_n579_, new_n1375_, new_n1711_, new_n1254_, new_n1689_, new_n438_, new_n1344_, new_n939_, new_n1393_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n1514_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n1526_, new_n397_, new_n1446_, new_n975_, new_n1199_, new_n399_, new_n1581_, new_n596_, new_n945_, new_n870_, new_n805_, new_n1420_, new_n1403_, new_n1115_, new_n1383_, new_n1231_, new_n948_, new_n1520_, new_n1055_, new_n1431_, new_n838_, new_n1609_, new_n923_, new_n1674_, new_n469_, new_n437_, new_n1085_, new_n1633_, new_n1607_, new_n794_, new_n457_, new_n1301_, new_n1128_, new_n1582_, new_n1002_, new_n1169_, new_n1702_, new_n448_, new_n384_, new_n900_, new_n1722_, new_n1329_, new_n1161_, new_n1648_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1663_, new_n1000_, new_n633_, new_n784_, new_n1273_, new_n1396_, new_n1491_, new_n1554_, new_n860_, new_n494_, new_n1160_, new_n1166_, new_n1536_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n1272_, new_n693_, new_n1287_, new_n1485_, new_n505_, new_n1462_, new_n619_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1538_, new_n1579_, new_n1289_, new_n1561_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n1095_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n1621_, new_n839_, new_n1030_, new_n485_, new_n578_, new_n525_, new_n1695_, new_n918_, new_n1586_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n1572_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n1387_, new_n719_, new_n869_, new_n1178_, new_n1525_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n520_, new_n1347_, new_n1001_, new_n825_, new_n1627_, new_n557_, new_n1642_, new_n1503_, new_n1742_, new_n507_, new_n741_, new_n806_, new_n1699_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n1286_, new_n1551_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n1650_, new_n807_, new_n1326_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n1080_, new_n583_, new_n617_, new_n1279_, new_n1467_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n916_, new_n428_, new_n487_, new_n675_, new_n1155_, new_n1186_, new_n1596_, new_n1261_, new_n1246_, new_n1488_, new_n922_, new_n387_, new_n476_, new_n987_, new_n1641_, new_n949_, new_n450_, new_n1394_, new_n1179_, new_n1088_, new_n1148_, new_n1146_, new_n569_, new_n555_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n692_, new_n502_, new_n623_, new_n446_, new_n590_, new_n826_, new_n789_, new_n1476_, new_n515_, new_n972_, new_n1634_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n1350_, new_n535_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n1736_, new_n1378_, new_n1478_, new_n1181_, new_n1093_, new_n597_, new_n1451_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1296_, new_n435_, new_n1309_, new_n1719_, new_n1010_, new_n776_, new_n687_, new_n1029_, new_n1649_, new_n1654_, new_n1515_, new_n638_, new_n523_, new_n909_, new_n1688_, new_n1571_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1610_, new_n1470_, new_n1112_, new_n1715_, new_n1156_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1475_, new_n1604_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n1731_, new_n1529_, new_n1541_, new_n645_, new_n1087_, new_n1096_, new_n723_, new_n1599_, new_n756_, new_n823_, new_n1549_, new_n1577_, new_n574_, new_n1500_, new_n928_, new_n1548_, new_n1578_, new_n1008_, new_n1687_, new_n1661_, new_n1615_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n1291_, new_n539_, new_n1399_, new_n803_, new_n1270_, new_n727_, new_n1531_, new_n1672_, new_n1589_, new_n1295_, new_n1173_, new_n704_, new_n1432_, new_n1570_, new_n1189_, new_n1197_, new_n1312_, new_n1502_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n467_, new_n404_, new_n1243_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n1666_, new_n865_, new_n358_, new_n877_, new_n1506_, new_n1583_, new_n1697_, new_n545_, new_n611_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n1556_, new_n947_, new_n994_, new_n982_, new_n1494_, new_n1449_, new_n964_, new_n1078_, new_n551_, new_n1408_, new_n455_, new_n1569_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n1605_, new_n464_, new_n1498_, new_n1588_, new_n573_, new_n765_, new_n1314_, new_n1103_;

nand g0000 ( new_n343_, N29, N42, N75 );
not g0001 ( N388, new_n343_ );
nand g0002 ( new_n345_, N29, N36, N80 );
not g0003 ( N389, new_n345_ );
nand g0004 ( new_n347_, N29, N36, N42 );
not g0005 ( N390, new_n347_ );
nand g0006 ( new_n349_, N85, N86 );
not g0007 ( N391, new_n349_ );
nand g0008 ( new_n351_, N1, N8 );
not g0009 ( new_n352_, new_n351_ );
nand g0010 ( new_n353_, new_n352_, N13, N17 );
not g0011 ( N418, new_n353_ );
not g0012 ( new_n355_, N13 );
not g0013 ( new_n356_, N17 );
nand g0014 ( new_n357_, N1, N26 );
nor g0015 ( new_n358_, new_n357_, new_n355_, new_n356_ );
nand g0016 ( N419, new_n358_, new_n347_ );
nand g0017 ( N420, N59, N75, N80 );
nand g0018 ( N421, N36, N59, N80 );
nand g0019 ( N422, N36, N42, N59 );
not g0020 ( new_n363_, keyIn_0_22 );
nor g0021 ( new_n364_, N87, N88 );
not g0022 ( new_n365_, new_n364_ );
nand g0023 ( new_n366_, new_n365_, N90 );
nand g0024 ( new_n367_, new_n366_, new_n363_ );
nand g0025 ( new_n368_, new_n365_, keyIn_0_22, N90 );
nand g0026 ( N423, new_n367_, new_n368_ );
nand g0027 ( N446, new_n358_, N390 );
not g0028 ( new_n371_, keyIn_0_0 );
nand g0029 ( new_n372_, N1, N26, N51 );
nand g0030 ( new_n373_, new_n372_, new_n371_ );
nand g0031 ( new_n374_, keyIn_0_0, N1, N26, N51 );
nand g0032 ( new_n375_, new_n373_, new_n374_ );
nand g0033 ( new_n376_, new_n375_, keyIn_0_26 );
not g0034 ( new_n377_, keyIn_0_26 );
nand g0035 ( new_n378_, new_n373_, new_n377_, new_n374_ );
nand g0036 ( new_n379_, new_n376_, new_n378_ );
not g0037 ( N447, new_n379_ );
not g0038 ( new_n381_, keyIn_0_2 );
nand g0039 ( new_n382_, new_n352_, N13, N55 );
nand g0040 ( new_n383_, new_n382_, new_n381_ );
not g0041 ( new_n384_, new_n383_ );
nor g0042 ( new_n385_, new_n382_, new_n381_ );
nor g0043 ( new_n386_, new_n384_, new_n385_ );
not g0044 ( new_n387_, new_n386_ );
nand g0045 ( new_n388_, N29, N68 );
nor g0046 ( N448, new_n387_, new_n388_ );
nand g0047 ( new_n390_, N59, N68, N74 );
nor g0048 ( N449, new_n387_, new_n390_ );
not g0049 ( new_n392_, N89 );
nor g0050 ( N450, new_n364_, new_n392_ );
not g0051 ( new_n394_, N135 );
nand g0052 ( new_n395_, N121, N126 );
not g0053 ( new_n396_, new_n395_ );
nor g0054 ( new_n397_, N121, N126 );
nor g0055 ( new_n398_, new_n396_, new_n397_ );
not g0056 ( new_n399_, new_n398_ );
not g0057 ( new_n400_, keyIn_0_6 );
nand g0058 ( new_n401_, new_n400_, N111, N116 );
not g0059 ( new_n402_, N111 );
not g0060 ( new_n403_, N116 );
nand g0061 ( new_n404_, new_n402_, new_n403_ );
nand g0062 ( new_n405_, N111, N116 );
nand g0063 ( new_n406_, new_n405_, keyIn_0_6 );
nand g0064 ( new_n407_, new_n406_, new_n401_, new_n404_ );
nand g0065 ( new_n408_, new_n399_, new_n407_ );
nand g0066 ( new_n409_, new_n398_, new_n401_, new_n404_, new_n406_ );
nand g0067 ( new_n410_, new_n408_, new_n409_ );
nand g0068 ( new_n411_, new_n410_, new_n394_ );
nand g0069 ( new_n412_, new_n408_, N135, new_n409_ );
nand g0070 ( new_n413_, new_n411_, new_n412_ );
not g0071 ( new_n414_, N130 );
not g0072 ( new_n415_, N91 );
not g0073 ( new_n416_, N96 );
nand g0074 ( new_n417_, new_n415_, new_n416_ );
nand g0075 ( new_n418_, N91, N96 );
nand g0076 ( new_n419_, new_n417_, new_n418_ );
not g0077 ( new_n420_, N101 );
not g0078 ( new_n421_, N106 );
nand g0079 ( new_n422_, new_n420_, new_n421_ );
nand g0080 ( new_n423_, N101, N106 );
nand g0081 ( new_n424_, new_n422_, new_n423_ );
nand g0082 ( new_n425_, new_n419_, new_n424_ );
nand g0083 ( new_n426_, new_n417_, new_n422_, new_n418_, new_n423_ );
nand g0084 ( new_n427_, new_n425_, new_n426_ );
nand g0085 ( new_n428_, new_n427_, new_n414_ );
nand g0086 ( new_n429_, new_n425_, N130, new_n426_ );
nand g0087 ( new_n430_, new_n428_, new_n429_ );
nand g0088 ( new_n431_, new_n413_, new_n430_ );
nand g0089 ( new_n432_, new_n411_, new_n412_, new_n428_, new_n429_ );
nand g0090 ( new_n433_, new_n431_, new_n432_ );
not g0091 ( N767, new_n433_ );
not g0092 ( new_n435_, N159 );
not g0093 ( new_n436_, N165 );
nand g0094 ( new_n437_, new_n435_, new_n436_ );
nand g0095 ( new_n438_, N159, N165 );
nand g0096 ( new_n439_, new_n437_, new_n438_ );
not g0097 ( new_n440_, N171 );
not g0098 ( new_n441_, N177 );
nand g0099 ( new_n442_, new_n440_, new_n441_ );
nand g0100 ( new_n443_, N171, N177 );
nand g0101 ( new_n444_, new_n442_, new_n443_ );
nand g0102 ( new_n445_, new_n439_, new_n444_ );
nand g0103 ( new_n446_, new_n437_, new_n442_, new_n438_, new_n443_ );
nand g0104 ( new_n447_, new_n445_, new_n446_ );
nand g0105 ( new_n448_, new_n447_, new_n414_ );
nand g0106 ( new_n449_, new_n445_, N130, new_n446_ );
nand g0107 ( new_n450_, new_n448_, new_n449_ );
not g0108 ( new_n451_, N207 );
not g0109 ( new_n452_, N183 );
not g0110 ( new_n453_, N189 );
nand g0111 ( new_n454_, new_n452_, new_n453_ );
nand g0112 ( new_n455_, N183, N189 );
nand g0113 ( new_n456_, new_n454_, new_n455_ );
not g0114 ( new_n457_, N195 );
not g0115 ( new_n458_, N201 );
nand g0116 ( new_n459_, new_n457_, new_n458_ );
nand g0117 ( new_n460_, N195, N201 );
nand g0118 ( new_n461_, new_n459_, new_n460_ );
nand g0119 ( new_n462_, new_n456_, new_n461_ );
nand g0120 ( new_n463_, new_n454_, new_n459_, new_n455_, new_n460_ );
nand g0121 ( new_n464_, new_n462_, new_n463_ );
nand g0122 ( new_n465_, new_n464_, new_n451_ );
nand g0123 ( new_n466_, new_n462_, N207, new_n463_ );
nand g0124 ( new_n467_, new_n465_, new_n466_ );
nand g0125 ( new_n468_, new_n450_, new_n467_ );
nand g0126 ( new_n469_, new_n448_, new_n465_, new_n449_, new_n466_ );
nand g0127 ( new_n470_, new_n468_, new_n469_ );
not g0128 ( N768, new_n470_ );
not g0129 ( new_n472_, keyIn_0_213 );
not g0130 ( new_n473_, keyIn_0_202 );
not g0131 ( new_n474_, keyIn_0_196 );
not g0132 ( new_n475_, keyIn_0_163 );
not g0133 ( new_n476_, keyIn_0_111 );
not g0134 ( new_n477_, keyIn_0_80 );
not g0135 ( new_n478_, keyIn_0_65 );
not g0136 ( new_n479_, keyIn_0_25 );
nand g0137 ( new_n480_, new_n375_, keyIn_0_18 );
not g0138 ( new_n481_, keyIn_0_18 );
nand g0139 ( new_n482_, new_n373_, new_n481_, new_n374_ );
nand g0140 ( new_n483_, new_n480_, new_n482_ );
nand g0141 ( new_n484_, new_n483_, new_n479_ );
nand g0142 ( new_n485_, new_n480_, keyIn_0_25, new_n482_ );
not g0143 ( new_n486_, keyIn_0_12 );
nand g0144 ( new_n487_, N59, N156 );
nand g0145 ( new_n488_, new_n487_, new_n486_ );
not g0146 ( new_n489_, new_n487_ );
nand g0147 ( new_n490_, new_n489_, keyIn_0_12 );
nand g0148 ( new_n491_, new_n490_, new_n488_ );
nand g0149 ( new_n492_, new_n491_, N17 );
not g0150 ( new_n493_, new_n492_ );
nand g0151 ( new_n494_, new_n484_, keyIn_0_35, new_n485_, new_n493_ );
not g0152 ( new_n495_, keyIn_0_35 );
nand g0153 ( new_n496_, new_n484_, new_n485_, new_n493_ );
nand g0154 ( new_n497_, new_n496_, new_n495_ );
nand g0155 ( new_n498_, new_n497_, N1, new_n494_ );
nand g0156 ( new_n499_, new_n498_, keyIn_0_46 );
not g0157 ( new_n500_, keyIn_0_46 );
nand g0158 ( new_n501_, new_n497_, new_n500_, N1, new_n494_ );
nand g0159 ( new_n502_, new_n499_, new_n501_ );
nand g0160 ( new_n503_, new_n502_, N153 );
nand g0161 ( new_n504_, new_n503_, new_n478_ );
nand g0162 ( new_n505_, new_n502_, keyIn_0_65, N153 );
nand g0163 ( new_n506_, new_n504_, new_n505_ );
nand g0164 ( new_n507_, new_n484_, new_n485_ );
not g0165 ( new_n508_, new_n507_ );
not g0166 ( new_n509_, N42 );
nand g0167 ( new_n510_, new_n356_, new_n509_ );
nand g0168 ( new_n511_, new_n510_, keyIn_0_13 );
nand g0169 ( new_n512_, N17, N42 );
nand g0170 ( new_n513_, new_n512_, keyIn_0_14 );
nor g0171 ( new_n514_, new_n512_, keyIn_0_14 );
nor g0172 ( new_n515_, keyIn_0_13, N17, N42 );
nor g0173 ( new_n516_, new_n514_, new_n515_ );
nand g0174 ( new_n517_, new_n516_, keyIn_0_24, new_n511_, new_n513_ );
not g0175 ( new_n518_, keyIn_0_24 );
not g0176 ( new_n519_, keyIn_0_14 );
nand g0177 ( new_n520_, new_n519_, N17, N42 );
not g0178 ( new_n521_, keyIn_0_13 );
nand g0179 ( new_n522_, new_n521_, new_n356_, new_n509_ );
nand g0180 ( new_n523_, new_n511_, new_n513_, new_n520_, new_n522_ );
nand g0181 ( new_n524_, new_n523_, new_n518_ );
nand g0182 ( new_n525_, new_n524_, new_n489_, new_n517_ );
not g0183 ( new_n526_, new_n525_ );
nand g0184 ( new_n527_, new_n508_, keyIn_0_34, new_n526_ );
not g0185 ( new_n528_, keyIn_0_34 );
nand g0186 ( new_n529_, new_n526_, new_n484_, new_n485_ );
nand g0187 ( new_n530_, new_n529_, new_n528_ );
not g0188 ( new_n531_, keyIn_0_28 );
nand g0189 ( new_n532_, N1, N8, N17, N51 );
nand g0190 ( new_n533_, new_n532_, keyIn_0_1 );
not g0191 ( new_n534_, keyIn_0_1 );
nand g0192 ( new_n535_, new_n352_, new_n534_, N17, N51 );
nand g0193 ( new_n536_, new_n535_, new_n533_ );
nand g0194 ( new_n537_, new_n536_, keyIn_0_19 );
not g0195 ( new_n538_, keyIn_0_19 );
nand g0196 ( new_n539_, new_n535_, new_n538_, new_n533_ );
not g0197 ( new_n540_, keyIn_0_5 );
nand g0198 ( new_n541_, N42, N59, N75 );
nand g0199 ( new_n542_, new_n541_, new_n540_ );
nand g0200 ( new_n543_, keyIn_0_5, N42, N59, N75 );
nand g0201 ( new_n544_, new_n542_, new_n543_ );
nand g0202 ( new_n545_, new_n544_, keyIn_0_21 );
not g0203 ( new_n546_, keyIn_0_21 );
nand g0204 ( new_n547_, new_n542_, new_n546_, new_n543_ );
nand g0205 ( new_n548_, new_n537_, new_n539_, new_n545_, new_n547_ );
nand g0206 ( new_n549_, new_n548_, new_n531_ );
nand g0207 ( new_n550_, new_n545_, new_n547_ );
not g0208 ( new_n551_, new_n550_ );
nand g0209 ( new_n552_, new_n551_, keyIn_0_28, new_n537_, new_n539_ );
nand g0210 ( new_n553_, new_n549_, new_n552_ );
not g0211 ( new_n554_, new_n553_ );
nand g0212 ( new_n555_, new_n530_, new_n554_, new_n527_ );
nand g0213 ( new_n556_, new_n555_, keyIn_0_37 );
not g0214 ( new_n557_, keyIn_0_37 );
nand g0215 ( new_n558_, new_n530_, new_n554_, new_n527_, new_n557_ );
nand g0216 ( new_n559_, new_n556_, new_n558_ );
nand g0217 ( new_n560_, new_n559_, N126 );
nand g0218 ( new_n561_, new_n560_, keyIn_0_66 );
not g0219 ( new_n562_, keyIn_0_66 );
nand g0220 ( new_n563_, new_n559_, new_n562_, N126 );
nand g0221 ( new_n564_, new_n561_, new_n506_, new_n477_, new_n563_ );
nand g0222 ( new_n565_, new_n561_, new_n506_, new_n563_ );
nand g0223 ( new_n566_, new_n565_, keyIn_0_80 );
not g0224 ( new_n567_, keyIn_0_50 );
not g0225 ( new_n568_, keyIn_0_4 );
nand g0226 ( new_n569_, N29, N75, N80 );
nand g0227 ( new_n570_, new_n569_, new_n568_ );
nand g0228 ( new_n571_, keyIn_0_4, N29, N75, N80 );
nand g0229 ( new_n572_, new_n570_, new_n571_ );
nand g0230 ( new_n573_, new_n508_, new_n572_ );
not g0231 ( new_n574_, new_n573_ );
nand g0232 ( new_n575_, new_n574_, N55 );
nor g0233 ( new_n576_, new_n575_, keyIn_0_33 );
nand g0234 ( new_n577_, new_n575_, keyIn_0_33 );
not g0235 ( new_n578_, new_n577_ );
not g0236 ( new_n579_, keyIn_0_23 );
not g0237 ( new_n580_, keyIn_0_8 );
nor g0238 ( new_n581_, new_n580_, N268 );
nand g0239 ( new_n582_, new_n580_, N268 );
not g0240 ( new_n583_, new_n582_ );
nor g0241 ( new_n584_, new_n583_, new_n581_ );
not g0242 ( new_n585_, new_n584_ );
nand g0243 ( new_n586_, new_n585_, new_n579_ );
nand g0244 ( new_n587_, new_n584_, keyIn_0_23 );
nand g0245 ( new_n588_, new_n586_, new_n587_ );
nor g0246 ( new_n589_, new_n578_, new_n576_, new_n588_ );
nor g0247 ( new_n590_, new_n589_, new_n567_ );
not g0248 ( new_n591_, new_n576_ );
not g0249 ( new_n592_, new_n588_ );
nand g0250 ( new_n593_, new_n591_, new_n577_, new_n592_ );
nor g0251 ( new_n594_, new_n593_, keyIn_0_50 );
nor g0252 ( new_n595_, new_n590_, new_n594_ );
nand g0253 ( new_n596_, new_n566_, new_n564_, new_n595_ );
nand g0254 ( new_n597_, new_n596_, keyIn_0_88 );
not g0255 ( new_n598_, keyIn_0_88 );
nand g0256 ( new_n599_, new_n566_, new_n598_, new_n564_, new_n595_ );
nand g0257 ( new_n600_, new_n597_, new_n458_, new_n599_ );
nand g0258 ( new_n601_, new_n600_, new_n476_ );
nand g0259 ( new_n602_, new_n597_, keyIn_0_111, new_n458_, new_n599_ );
nand g0260 ( new_n603_, new_n601_, new_n602_ );
not g0261 ( new_n604_, new_n603_ );
nand g0262 ( new_n605_, new_n597_, new_n599_ );
nand g0263 ( new_n606_, new_n605_, N201 );
nand g0264 ( new_n607_, new_n606_, keyIn_0_110 );
not g0265 ( new_n608_, keyIn_0_110 );
nand g0266 ( new_n609_, new_n605_, new_n608_, N201 );
nand g0267 ( new_n610_, new_n607_, new_n609_ );
nand g0268 ( new_n611_, new_n604_, new_n610_ );
nand g0269 ( new_n612_, new_n611_, keyIn_0_135 );
not g0270 ( new_n613_, keyIn_0_135 );
nand g0271 ( new_n614_, new_n604_, new_n610_, new_n613_ );
nand g0272 ( new_n615_, new_n612_, new_n614_ );
not g0273 ( new_n616_, new_n615_ );
nand g0274 ( new_n617_, new_n616_, N261 );
nand g0275 ( new_n618_, new_n617_, new_n475_ );
not g0276 ( new_n619_, keyIn_0_162 );
not g0277 ( new_n620_, N261 );
nand g0278 ( new_n621_, new_n615_, new_n620_ );
nand g0279 ( new_n622_, new_n621_, new_n619_ );
nand g0280 ( new_n623_, new_n615_, keyIn_0_162, new_n620_ );
nand g0281 ( new_n624_, new_n616_, keyIn_0_163, N261 );
nand g0282 ( new_n625_, new_n618_, new_n622_, new_n623_, new_n624_ );
not g0283 ( new_n626_, new_n625_ );
nand g0284 ( new_n627_, new_n626_, keyIn_0_182 );
not g0285 ( new_n628_, keyIn_0_182 );
nand g0286 ( new_n629_, new_n625_, new_n628_ );
nand g0287 ( new_n630_, new_n627_, new_n629_ );
nand g0288 ( new_n631_, new_n630_, keyIn_0_190, N219 );
not g0289 ( new_n632_, keyIn_0_190 );
nand g0290 ( new_n633_, new_n630_, N219 );
nand g0291 ( new_n634_, new_n633_, new_n632_ );
nand g0292 ( new_n635_, N121, N210 );
nand g0293 ( new_n636_, new_n635_, keyIn_0_17 );
not g0294 ( new_n637_, keyIn_0_17 );
nand g0295 ( new_n638_, new_n637_, N121, N210 );
nand g0296 ( new_n639_, new_n636_, new_n638_ );
not g0297 ( new_n640_, new_n639_ );
nand g0298 ( new_n641_, new_n634_, new_n631_, new_n640_ );
nand g0299 ( new_n642_, new_n641_, new_n474_ );
nand g0300 ( new_n643_, new_n634_, keyIn_0_196, new_n631_, new_n640_ );
nand g0301 ( new_n644_, new_n642_, new_n643_ );
nand g0302 ( new_n645_, new_n616_, keyIn_0_164, N228 );
not g0303 ( new_n646_, keyIn_0_164 );
nand g0304 ( new_n647_, new_n616_, N228 );
nand g0305 ( new_n648_, new_n647_, new_n646_ );
not g0306 ( new_n649_, keyIn_0_165 );
not g0307 ( new_n650_, keyIn_0_134 );
nand g0308 ( new_n651_, new_n610_, new_n650_ );
nand g0309 ( new_n652_, new_n607_, keyIn_0_134, new_n609_ );
nand g0310 ( new_n653_, new_n651_, new_n652_ );
nand g0311 ( new_n654_, new_n653_, N237 );
nand g0312 ( new_n655_, new_n654_, new_n649_ );
nand g0313 ( new_n656_, new_n653_, keyIn_0_165, N237 );
nand g0314 ( new_n657_, new_n648_, new_n645_, new_n655_, new_n656_ );
not g0315 ( new_n658_, new_n657_ );
nand g0316 ( new_n659_, new_n658_, keyIn_0_183 );
not g0317 ( new_n660_, keyIn_0_183 );
nand g0318 ( new_n661_, new_n657_, new_n660_ );
nand g0319 ( new_n662_, new_n659_, new_n661_ );
not g0320 ( new_n663_, keyIn_0_36 );
not g0321 ( new_n664_, keyIn_0_30 );
not g0322 ( new_n665_, keyIn_0_27 );
nand g0323 ( new_n666_, N42, N59, N68, N72 );
not g0324 ( new_n667_, new_n666_ );
nand g0325 ( new_n668_, new_n667_, keyIn_0_3 );
not g0326 ( new_n669_, keyIn_0_3 );
nand g0327 ( new_n670_, new_n666_, new_n669_ );
nand g0328 ( new_n671_, new_n386_, new_n668_, new_n670_ );
nand g0329 ( new_n672_, new_n671_, keyIn_0_20 );
not g0330 ( new_n673_, keyIn_0_20 );
nand g0331 ( new_n674_, new_n386_, new_n673_, new_n668_, new_n670_ );
nand g0332 ( new_n675_, new_n672_, new_n674_ );
nand g0333 ( new_n676_, new_n675_, N73 );
nand g0334 ( new_n677_, new_n676_, new_n665_ );
nand g0335 ( new_n678_, new_n675_, keyIn_0_27, N73 );
nand g0336 ( new_n679_, new_n677_, new_n678_ );
nand g0337 ( new_n680_, new_n679_, new_n664_ );
nand g0338 ( new_n681_, new_n677_, keyIn_0_30, new_n678_ );
nand g0339 ( new_n682_, new_n680_, new_n681_ );
nand g0340 ( new_n683_, new_n682_, new_n663_ );
nand g0341 ( new_n684_, new_n680_, keyIn_0_36, new_n681_ );
nand g0342 ( new_n685_, new_n683_, new_n684_ );
nand g0343 ( new_n686_, new_n685_, N201 );
not g0344 ( new_n687_, keyIn_0_136 );
nand g0345 ( new_n688_, new_n605_, N246 );
nand g0346 ( new_n689_, new_n688_, keyIn_0_112 );
not g0347 ( new_n690_, keyIn_0_112 );
nand g0348 ( new_n691_, new_n605_, new_n690_, N246 );
nand g0349 ( new_n692_, new_n689_, new_n691_ );
nand g0350 ( new_n693_, N255, N267 );
nand g0351 ( new_n694_, new_n692_, new_n693_ );
nand g0352 ( new_n695_, new_n694_, new_n687_ );
nand g0353 ( new_n696_, new_n692_, keyIn_0_136, new_n693_ );
nand g0354 ( new_n697_, new_n695_, new_n696_ );
nand g0355 ( new_n698_, new_n662_, new_n686_, new_n697_ );
not g0356 ( new_n699_, new_n698_ );
nand g0357 ( new_n700_, new_n644_, new_n699_ );
nand g0358 ( new_n701_, new_n700_, new_n473_ );
nand g0359 ( new_n702_, new_n644_, keyIn_0_202, new_n699_ );
nand g0360 ( new_n703_, new_n701_, new_n702_ );
nand g0361 ( new_n704_, new_n703_, new_n472_ );
nand g0362 ( new_n705_, new_n701_, keyIn_0_213, new_n702_ );
nand g0363 ( new_n706_, new_n704_, new_n705_ );
nand g0364 ( new_n707_, new_n706_, keyIn_0_224 );
not g0365 ( new_n708_, keyIn_0_224 );
nand g0366 ( new_n709_, new_n704_, new_n708_, new_n705_ );
nand g0367 ( new_n710_, new_n707_, new_n709_ );
not g0368 ( N850, new_n710_ );
not g0369 ( new_n712_, keyIn_0_238 );
not g0370 ( new_n713_, keyIn_0_221 );
not g0371 ( new_n714_, keyIn_0_199 );
not g0372 ( new_n715_, keyIn_0_193 );
not g0373 ( new_n716_, keyIn_0_184 );
nand g0374 ( new_n717_, new_n559_, N116 );
nand g0375 ( new_n718_, new_n717_, keyIn_0_62 );
not g0376 ( new_n719_, keyIn_0_62 );
nand g0377 ( new_n720_, new_n559_, new_n719_, N116 );
nand g0378 ( new_n721_, new_n718_, new_n720_ );
nand g0379 ( new_n722_, new_n502_, N146 );
nand g0380 ( new_n723_, new_n722_, keyIn_0_61 );
not g0381 ( new_n724_, keyIn_0_61 );
nand g0382 ( new_n725_, new_n502_, new_n724_, N146 );
nand g0383 ( new_n726_, new_n723_, new_n725_ );
not g0384 ( new_n727_, new_n726_ );
nand g0385 ( new_n728_, new_n721_, keyIn_0_78, new_n727_ );
not g0386 ( new_n729_, keyIn_0_78 );
nand g0387 ( new_n730_, new_n721_, new_n727_ );
nand g0388 ( new_n731_, new_n730_, new_n729_ );
not g0389 ( new_n732_, keyIn_0_48 );
nor g0390 ( new_n733_, new_n589_, new_n732_ );
nor g0391 ( new_n734_, new_n593_, keyIn_0_48 );
nor g0392 ( new_n735_, new_n733_, new_n734_ );
nand g0393 ( new_n736_, new_n731_, new_n728_, new_n735_ );
nand g0394 ( new_n737_, new_n736_, keyIn_0_86 );
not g0395 ( new_n738_, keyIn_0_86 );
nand g0396 ( new_n739_, new_n731_, new_n738_, new_n728_, new_n735_ );
nand g0397 ( new_n740_, new_n737_, new_n739_ );
nand g0398 ( new_n741_, new_n740_, new_n453_ );
nand g0399 ( new_n742_, new_n741_, keyIn_0_105 );
not g0400 ( new_n743_, keyIn_0_105 );
nand g0401 ( new_n744_, new_n740_, new_n743_, new_n453_ );
nand g0402 ( new_n745_, new_n742_, new_n744_ );
not g0403 ( new_n746_, keyIn_0_108 );
not g0404 ( new_n747_, keyIn_0_87 );
not g0405 ( new_n748_, keyIn_0_79 );
not g0406 ( new_n749_, keyIn_0_64 );
nand g0407 ( new_n750_, new_n559_, N121 );
nand g0408 ( new_n751_, new_n750_, new_n749_ );
not g0409 ( new_n752_, keyIn_0_63 );
nand g0410 ( new_n753_, new_n502_, N149 );
nand g0411 ( new_n754_, new_n753_, new_n752_ );
nand g0412 ( new_n755_, new_n559_, keyIn_0_64, N121 );
nand g0413 ( new_n756_, new_n502_, keyIn_0_63, N149 );
nand g0414 ( new_n757_, new_n755_, new_n756_ );
not g0415 ( new_n758_, new_n757_ );
nand g0416 ( new_n759_, new_n758_, new_n748_, new_n751_, new_n754_ );
nand g0417 ( new_n760_, new_n751_, new_n754_, new_n755_, new_n756_ );
nand g0418 ( new_n761_, new_n760_, keyIn_0_79 );
nor g0419 ( new_n762_, new_n589_, keyIn_0_49 );
not g0420 ( new_n763_, keyIn_0_49 );
nor g0421 ( new_n764_, new_n593_, new_n763_ );
nor g0422 ( new_n765_, new_n762_, new_n764_ );
nand g0423 ( new_n766_, new_n759_, new_n761_, new_n765_ );
nand g0424 ( new_n767_, new_n766_, new_n747_ );
nand g0425 ( new_n768_, new_n759_, new_n761_, keyIn_0_87, new_n765_ );
nand g0426 ( new_n769_, new_n767_, new_n768_ );
nand g0427 ( new_n770_, new_n769_, new_n457_ );
nand g0428 ( new_n771_, new_n770_, new_n746_ );
nand g0429 ( new_n772_, new_n769_, keyIn_0_108, new_n457_ );
nand g0430 ( new_n773_, new_n771_, new_n772_ );
not g0431 ( new_n774_, new_n773_ );
nand g0432 ( new_n775_, new_n653_, new_n745_, new_n774_ );
nand g0433 ( new_n776_, new_n775_, keyIn_0_168 );
not g0434 ( new_n777_, keyIn_0_168 );
nand g0435 ( new_n778_, new_n653_, new_n777_, new_n745_, new_n774_ );
nand g0436 ( new_n779_, new_n776_, new_n778_ );
not g0437 ( new_n780_, keyIn_0_167 );
not g0438 ( new_n781_, keyIn_0_107 );
nand g0439 ( new_n782_, new_n767_, N195, new_n768_ );
nand g0440 ( new_n783_, new_n782_, new_n781_ );
not g0441 ( new_n784_, new_n769_ );
nand g0442 ( new_n785_, new_n784_, keyIn_0_107, N195 );
nand g0443 ( new_n786_, new_n785_, new_n783_ );
nand g0444 ( new_n787_, new_n786_, keyIn_0_131 );
not g0445 ( new_n788_, keyIn_0_131 );
nand g0446 ( new_n789_, new_n785_, new_n788_, new_n783_ );
nand g0447 ( new_n790_, new_n787_, new_n745_, new_n789_ );
nand g0448 ( new_n791_, new_n790_, new_n780_ );
nand g0449 ( new_n792_, new_n787_, keyIn_0_167, new_n745_, new_n789_ );
nand g0450 ( new_n793_, new_n791_, new_n792_ );
nand g0451 ( new_n794_, new_n601_, N261, new_n602_ );
nor g0452 ( new_n795_, new_n773_, new_n794_ );
nand g0453 ( new_n796_, new_n795_, keyIn_0_139, new_n745_ );
not g0454 ( new_n797_, keyIn_0_139 );
not g0455 ( new_n798_, new_n794_ );
nand g0456 ( new_n799_, new_n745_, new_n771_, new_n798_, new_n772_ );
nand g0457 ( new_n800_, new_n799_, new_n797_ );
not g0458 ( new_n801_, keyIn_0_155 );
nand g0459 ( new_n802_, new_n737_, N189, new_n739_ );
nand g0460 ( new_n803_, new_n802_, keyIn_0_104 );
not g0461 ( new_n804_, keyIn_0_104 );
nand g0462 ( new_n805_, new_n737_, new_n804_, N189, new_n739_ );
nand g0463 ( new_n806_, new_n803_, new_n805_ );
nand g0464 ( new_n807_, new_n806_, keyIn_0_128 );
not g0465 ( new_n808_, keyIn_0_128 );
nand g0466 ( new_n809_, new_n803_, new_n808_, new_n805_ );
nand g0467 ( new_n810_, new_n807_, new_n809_ );
nand g0468 ( new_n811_, new_n810_, new_n801_ );
nand g0469 ( new_n812_, new_n807_, keyIn_0_155, new_n809_ );
nand g0470 ( new_n813_, new_n800_, new_n811_, new_n796_, new_n812_ );
not g0471 ( new_n814_, new_n813_ );
nand g0472 ( new_n815_, new_n814_, new_n779_, new_n793_ );
nand g0473 ( new_n816_, new_n815_, keyIn_0_176 );
not g0474 ( new_n817_, keyIn_0_176 );
nand g0475 ( new_n818_, new_n814_, new_n779_, new_n817_, new_n793_ );
nand g0476 ( new_n819_, new_n816_, new_n818_ );
not g0477 ( new_n820_, new_n819_ );
not g0478 ( new_n821_, keyIn_0_101 );
not g0479 ( new_n822_, keyIn_0_85 );
not g0480 ( new_n823_, keyIn_0_77 );
not g0481 ( new_n824_, keyIn_0_60 );
nand g0482 ( new_n825_, new_n559_, N111 );
nand g0483 ( new_n826_, new_n825_, new_n824_ );
nand g0484 ( new_n827_, new_n502_, N143 );
nand g0485 ( new_n828_, new_n827_, keyIn_0_59 );
nand g0486 ( new_n829_, new_n826_, new_n828_ );
not g0487 ( new_n830_, new_n829_ );
not g0488 ( new_n831_, keyIn_0_59 );
nand g0489 ( new_n832_, new_n502_, new_n831_, N143 );
nand g0490 ( new_n833_, new_n559_, keyIn_0_60, N111 );
nand g0491 ( new_n834_, new_n830_, new_n823_, new_n832_, new_n833_ );
not g0492 ( new_n835_, keyIn_0_47 );
nand g0493 ( new_n836_, new_n589_, new_n835_ );
nand g0494 ( new_n837_, new_n593_, keyIn_0_47 );
nand g0495 ( new_n838_, new_n836_, new_n837_ );
nand g0496 ( new_n839_, new_n830_, new_n832_, new_n833_ );
nand g0497 ( new_n840_, new_n839_, keyIn_0_77 );
nand g0498 ( new_n841_, new_n840_, new_n834_, new_n838_ );
nand g0499 ( new_n842_, new_n841_, new_n822_ );
nand g0500 ( new_n843_, new_n840_, keyIn_0_85, new_n834_, new_n838_ );
nand g0501 ( new_n844_, new_n842_, new_n843_ );
not g0502 ( new_n845_, new_n844_ );
nand g0503 ( new_n846_, new_n845_, N183 );
nand g0504 ( new_n847_, new_n846_, new_n821_ );
nand g0505 ( new_n848_, new_n845_, keyIn_0_101, N183 );
nand g0506 ( new_n849_, new_n847_, new_n848_ );
not g0507 ( new_n850_, new_n849_ );
not g0508 ( new_n851_, keyIn_0_102 );
nand g0509 ( new_n852_, new_n844_, new_n452_ );
nand g0510 ( new_n853_, new_n852_, new_n851_ );
nand g0511 ( new_n854_, new_n844_, keyIn_0_102, new_n452_ );
nand g0512 ( new_n855_, new_n853_, new_n854_ );
nand g0513 ( new_n856_, new_n850_, new_n855_ );
nand g0514 ( new_n857_, new_n856_, keyIn_0_126 );
not g0515 ( new_n858_, keyIn_0_126 );
nand g0516 ( new_n859_, new_n850_, new_n858_, new_n855_ );
nand g0517 ( new_n860_, new_n857_, new_n859_ );
not g0518 ( new_n861_, new_n860_ );
nand g0519 ( new_n862_, new_n820_, new_n861_ );
nand g0520 ( new_n863_, new_n862_, new_n716_ );
nand g0521 ( new_n864_, new_n820_, keyIn_0_184, new_n861_ );
nand g0522 ( new_n865_, new_n863_, new_n864_ );
nand g0523 ( new_n866_, new_n819_, new_n860_ );
nand g0524 ( new_n867_, new_n866_, keyIn_0_185 );
not g0525 ( new_n868_, keyIn_0_185 );
nand g0526 ( new_n869_, new_n819_, new_n868_, new_n860_ );
nand g0527 ( new_n870_, new_n867_, new_n869_ );
nand g0528 ( new_n871_, new_n865_, new_n870_ );
nand g0529 ( new_n872_, new_n871_, new_n715_ );
nand g0530 ( new_n873_, new_n865_, keyIn_0_193, new_n870_ );
nand g0531 ( new_n874_, new_n872_, new_n873_ );
nand g0532 ( new_n875_, new_n874_, N219 );
nand g0533 ( new_n876_, new_n875_, new_n714_ );
nand g0534 ( new_n877_, new_n874_, keyIn_0_199, N219 );
nand g0535 ( new_n878_, new_n876_, new_n877_ );
nand g0536 ( new_n879_, N106, N210 );
nand g0537 ( new_n880_, new_n878_, new_n879_ );
nand g0538 ( new_n881_, new_n880_, keyIn_0_210 );
not g0539 ( new_n882_, keyIn_0_210 );
nand g0540 ( new_n883_, new_n878_, new_n882_, new_n879_ );
nand g0541 ( new_n884_, new_n881_, new_n883_ );
not g0542 ( new_n885_, keyIn_0_153 );
nand g0543 ( new_n886_, new_n860_, N228 );
nand g0544 ( new_n887_, new_n886_, new_n885_ );
nand g0545 ( new_n888_, new_n860_, keyIn_0_153, N228 );
nand g0546 ( new_n889_, new_n887_, new_n888_ );
not g0547 ( new_n890_, keyIn_0_125 );
nand g0548 ( new_n891_, new_n850_, new_n890_ );
nand g0549 ( new_n892_, new_n849_, keyIn_0_125 );
nand g0550 ( new_n893_, new_n891_, new_n892_ );
not g0551 ( new_n894_, new_n893_ );
nand g0552 ( new_n895_, new_n894_, N237 );
nand g0553 ( new_n896_, new_n895_, keyIn_0_154 );
not g0554 ( new_n897_, keyIn_0_154 );
nand g0555 ( new_n898_, new_n894_, new_n897_, N237 );
nand g0556 ( new_n899_, new_n896_, new_n898_ );
nand g0557 ( new_n900_, new_n889_, keyIn_0_177, new_n899_ );
not g0558 ( new_n901_, keyIn_0_103 );
nand g0559 ( new_n902_, new_n845_, new_n901_, N246 );
nand g0560 ( new_n903_, new_n845_, N246 );
nand g0561 ( new_n904_, new_n903_, keyIn_0_103 );
nand g0562 ( new_n905_, new_n685_, N183 );
nand g0563 ( new_n906_, new_n905_, keyIn_0_71 );
not g0564 ( new_n907_, keyIn_0_71 );
nand g0565 ( new_n908_, new_n685_, new_n907_, N183 );
nand g0566 ( new_n909_, new_n906_, new_n908_ );
not g0567 ( new_n910_, new_n909_ );
nand g0568 ( new_n911_, new_n904_, new_n902_, new_n910_ );
nand g0569 ( new_n912_, new_n911_, keyIn_0_127 );
not g0570 ( new_n913_, keyIn_0_127 );
nand g0571 ( new_n914_, new_n904_, new_n913_, new_n902_, new_n910_ );
nand g0572 ( new_n915_, new_n912_, new_n914_ );
not g0573 ( new_n916_, keyIn_0_177 );
nand g0574 ( new_n917_, new_n889_, new_n899_ );
nand g0575 ( new_n918_, new_n917_, new_n916_ );
nand g0576 ( new_n919_, new_n918_, new_n900_, new_n915_ );
not g0577 ( new_n920_, new_n919_ );
nand g0578 ( new_n921_, new_n884_, new_n920_ );
nand g0579 ( new_n922_, new_n921_, new_n713_ );
nand g0580 ( new_n923_, new_n884_, keyIn_0_221, new_n920_ );
nand g0581 ( new_n924_, new_n922_, new_n923_ );
nand g0582 ( new_n925_, new_n924_, keyIn_0_230 );
not g0583 ( new_n926_, keyIn_0_230 );
nand g0584 ( new_n927_, new_n922_, new_n926_, new_n923_ );
nand g0585 ( new_n928_, new_n925_, new_n927_ );
nand g0586 ( new_n929_, new_n928_, new_n712_ );
nand g0587 ( new_n930_, new_n925_, keyIn_0_238, new_n927_ );
nand g0588 ( N863, new_n929_, new_n930_ );
not g0589 ( new_n932_, keyIn_0_194 );
not g0590 ( new_n933_, keyIn_0_186 );
not g0591 ( new_n934_, keyIn_0_166 );
nand g0592 ( new_n935_, new_n653_, new_n774_ );
nand g0593 ( new_n936_, new_n935_, new_n934_ );
nand g0594 ( new_n937_, new_n653_, keyIn_0_166, new_n774_ );
nand g0595 ( new_n938_, new_n936_, new_n937_ );
not g0596 ( new_n939_, keyIn_0_138 );
nor g0597 ( new_n940_, new_n795_, new_n939_ );
nor g0598 ( new_n941_, new_n773_, keyIn_0_138, new_n794_ );
nor g0599 ( new_n942_, new_n940_, new_n941_ );
not g0600 ( new_n943_, keyIn_0_158 );
nand g0601 ( new_n944_, new_n787_, new_n789_ );
not g0602 ( new_n945_, new_n944_ );
nand g0603 ( new_n946_, new_n945_, new_n943_ );
nand g0604 ( new_n947_, new_n944_, keyIn_0_158 );
nand g0605 ( new_n948_, new_n946_, new_n947_ );
nor g0606 ( new_n949_, new_n948_, new_n942_ );
nand g0607 ( new_n950_, new_n949_, new_n938_ );
nand g0608 ( new_n951_, new_n950_, keyIn_0_178 );
not g0609 ( new_n952_, keyIn_0_178 );
nand g0610 ( new_n953_, new_n949_, new_n952_, new_n938_ );
nand g0611 ( new_n954_, new_n951_, new_n953_ );
not g0612 ( new_n955_, keyIn_0_129 );
nand g0613 ( new_n956_, new_n745_, new_n806_ );
nand g0614 ( new_n957_, new_n956_, new_n955_ );
nand g0615 ( new_n958_, new_n745_, keyIn_0_129, new_n806_ );
nand g0616 ( new_n959_, new_n957_, new_n958_ );
nand g0617 ( new_n960_, new_n954_, new_n959_ );
nand g0618 ( new_n961_, new_n960_, new_n933_ );
nand g0619 ( new_n962_, new_n954_, keyIn_0_186, new_n959_ );
nand g0620 ( new_n963_, new_n961_, new_n962_ );
not g0621 ( new_n964_, new_n954_ );
not g0622 ( new_n965_, new_n959_ );
nand g0623 ( new_n966_, new_n964_, new_n965_ );
nand g0624 ( new_n967_, new_n966_, keyIn_0_187 );
not g0625 ( new_n968_, keyIn_0_187 );
nand g0626 ( new_n969_, new_n964_, new_n968_, new_n965_ );
nand g0627 ( new_n970_, new_n967_, new_n969_ );
not g0628 ( new_n971_, new_n970_ );
nand g0629 ( new_n972_, new_n971_, new_n963_ );
nand g0630 ( new_n973_, new_n972_, new_n932_ );
nand g0631 ( new_n974_, new_n971_, keyIn_0_194, new_n963_ );
nand g0632 ( new_n975_, new_n973_, new_n974_ );
nand g0633 ( new_n976_, new_n975_, N219 );
nand g0634 ( new_n977_, new_n976_, keyIn_0_200 );
not g0635 ( new_n978_, keyIn_0_200 );
nand g0636 ( new_n979_, new_n975_, new_n978_, N219 );
nand g0637 ( new_n980_, new_n977_, new_n979_ );
not g0638 ( new_n981_, keyIn_0_16 );
nand g0639 ( new_n982_, N111, N210 );
nand g0640 ( new_n983_, new_n982_, new_n981_ );
nand g0641 ( new_n984_, keyIn_0_16, N111, N210 );
nand g0642 ( new_n985_, new_n983_, new_n984_ );
not g0643 ( new_n986_, new_n985_ );
nand g0644 ( new_n987_, new_n980_, new_n986_ );
nand g0645 ( new_n988_, new_n987_, keyIn_0_211 );
not g0646 ( new_n989_, keyIn_0_211 );
nand g0647 ( new_n990_, new_n980_, new_n989_, new_n986_ );
nand g0648 ( new_n991_, new_n988_, new_n990_ );
not g0649 ( new_n992_, keyIn_0_179 );
not g0650 ( new_n993_, keyIn_0_156 );
nand g0651 ( new_n994_, new_n965_, N228 );
nand g0652 ( new_n995_, new_n994_, new_n993_ );
nand g0653 ( new_n996_, new_n965_, keyIn_0_156, N228 );
nand g0654 ( new_n997_, new_n995_, new_n996_ );
not g0655 ( new_n998_, keyIn_0_157 );
nand g0656 ( new_n999_, new_n810_, N237 );
nand g0657 ( new_n1000_, new_n999_, new_n998_ );
nand g0658 ( new_n1001_, new_n810_, keyIn_0_157, N237 );
nand g0659 ( new_n1002_, new_n1000_, new_n1001_ );
nand g0660 ( new_n1003_, new_n997_, new_n1002_ );
nand g0661 ( new_n1004_, new_n1003_, new_n992_ );
nand g0662 ( new_n1005_, new_n997_, keyIn_0_179, new_n1002_ );
nand g0663 ( new_n1006_, new_n1004_, new_n1005_ );
not g0664 ( new_n1007_, keyIn_0_130 );
not g0665 ( new_n1008_, new_n740_ );
nand g0666 ( new_n1009_, new_n1008_, keyIn_0_106, N246 );
nand g0667 ( new_n1010_, N255, N259 );
not g0668 ( new_n1011_, keyIn_0_106 );
nand g0669 ( new_n1012_, new_n1008_, N246 );
nand g0670 ( new_n1013_, new_n1012_, new_n1011_ );
nand g0671 ( new_n1014_, new_n1013_, new_n1007_, new_n1009_, new_n1010_ );
not g0672 ( new_n1015_, keyIn_0_72 );
nand g0673 ( new_n1016_, new_n685_, N189 );
nand g0674 ( new_n1017_, new_n1016_, new_n1015_ );
nand g0675 ( new_n1018_, new_n685_, keyIn_0_72, N189 );
nand g0676 ( new_n1019_, new_n1017_, new_n1018_ );
nand g0677 ( new_n1020_, new_n1013_, new_n1009_, new_n1010_ );
nand g0678 ( new_n1021_, new_n1020_, keyIn_0_130 );
nand g0679 ( new_n1022_, new_n1006_, new_n1014_, new_n1019_, new_n1021_ );
not g0680 ( new_n1023_, new_n1022_ );
nand g0681 ( new_n1024_, new_n991_, new_n1023_ );
nand g0682 ( new_n1025_, new_n1024_, keyIn_0_222 );
not g0683 ( new_n1026_, keyIn_0_222 );
nand g0684 ( new_n1027_, new_n991_, new_n1026_, new_n1023_ );
nand g0685 ( new_n1028_, new_n1025_, new_n1027_ );
nand g0686 ( new_n1029_, new_n1028_, keyIn_0_231 );
not g0687 ( new_n1030_, keyIn_0_231 );
nand g0688 ( new_n1031_, new_n1025_, new_n1030_, new_n1027_ );
nand g0689 ( new_n1032_, new_n1029_, new_n1031_ );
nand g0690 ( new_n1033_, new_n1032_, keyIn_0_239 );
not g0691 ( new_n1034_, keyIn_0_239 );
nand g0692 ( new_n1035_, new_n1029_, new_n1034_, new_n1031_ );
nand g0693 ( new_n1036_, new_n1033_, new_n1035_ );
not g0694 ( N864, new_n1036_ );
not g0695 ( new_n1038_, keyIn_0_240 );
not g0696 ( new_n1039_, keyIn_0_195 );
not g0697 ( new_n1040_, keyIn_0_188 );
nor g0698 ( new_n1041_, new_n786_, new_n773_ );
not g0699 ( new_n1042_, new_n1041_ );
nand g0700 ( new_n1043_, new_n1042_, keyIn_0_132 );
not g0701 ( new_n1044_, keyIn_0_132 );
nand g0702 ( new_n1045_, new_n1041_, new_n1044_ );
nand g0703 ( new_n1046_, new_n1043_, new_n1045_ );
not g0704 ( new_n1047_, new_n1046_ );
not g0705 ( new_n1048_, keyIn_0_180 );
not g0706 ( new_n1049_, keyIn_0_161 );
nand g0707 ( new_n1050_, new_n651_, new_n1049_, new_n652_ );
nand g0708 ( new_n1051_, new_n653_, keyIn_0_161 );
not g0709 ( new_n1052_, keyIn_0_137 );
nand g0710 ( new_n1053_, new_n798_, new_n1052_ );
nand g0711 ( new_n1054_, new_n794_, keyIn_0_137 );
nand g0712 ( new_n1055_, new_n1053_, new_n1054_ );
not g0713 ( new_n1056_, new_n1055_ );
nand g0714 ( new_n1057_, new_n1056_, new_n1051_, new_n1050_ );
nand g0715 ( new_n1058_, new_n1057_, new_n1048_ );
nand g0716 ( new_n1059_, new_n1056_, new_n1051_, keyIn_0_180, new_n1050_ );
nand g0717 ( new_n1060_, new_n1058_, new_n1059_ );
nand g0718 ( new_n1061_, new_n1060_, new_n1047_ );
nand g0719 ( new_n1062_, new_n1061_, new_n1040_ );
nand g0720 ( new_n1063_, new_n1060_, keyIn_0_188, new_n1047_ );
nand g0721 ( new_n1064_, new_n1062_, new_n1063_ );
not g0722 ( new_n1065_, new_n1060_ );
nand g0723 ( new_n1066_, new_n1065_, new_n1046_ );
nand g0724 ( new_n1067_, new_n1066_, keyIn_0_189 );
not g0725 ( new_n1068_, keyIn_0_189 );
nand g0726 ( new_n1069_, new_n1065_, new_n1068_, new_n1046_ );
nand g0727 ( new_n1070_, new_n1067_, new_n1069_ );
not g0728 ( new_n1071_, new_n1070_ );
nand g0729 ( new_n1072_, new_n1071_, new_n1064_ );
nand g0730 ( new_n1073_, new_n1072_, new_n1039_ );
nand g0731 ( new_n1074_, new_n1071_, keyIn_0_195, new_n1064_ );
nand g0732 ( new_n1075_, new_n1073_, new_n1074_ );
nand g0733 ( new_n1076_, new_n1075_, keyIn_0_201, N219 );
nand g0734 ( new_n1077_, N116, N210 );
not g0735 ( new_n1078_, keyIn_0_201 );
nand g0736 ( new_n1079_, new_n1075_, N219 );
nand g0737 ( new_n1080_, new_n1079_, new_n1078_ );
nand g0738 ( new_n1081_, new_n1080_, keyIn_0_212, new_n1076_, new_n1077_ );
not g0739 ( new_n1082_, keyIn_0_212 );
nand g0740 ( new_n1083_, new_n1080_, new_n1076_, new_n1077_ );
nand g0741 ( new_n1084_, new_n1083_, new_n1082_ );
not g0742 ( new_n1085_, keyIn_0_181 );
not g0743 ( new_n1086_, keyIn_0_159 );
nand g0744 ( new_n1087_, new_n1046_, N228 );
nand g0745 ( new_n1088_, new_n1087_, new_n1086_ );
nand g0746 ( new_n1089_, new_n1046_, keyIn_0_159, N228 );
nand g0747 ( new_n1090_, new_n1088_, new_n1089_ );
nand g0748 ( new_n1091_, new_n945_, N237 );
nand g0749 ( new_n1092_, new_n1091_, keyIn_0_160 );
not g0750 ( new_n1093_, keyIn_0_160 );
nand g0751 ( new_n1094_, new_n945_, new_n1093_, N237 );
nand g0752 ( new_n1095_, new_n1092_, new_n1094_ );
nand g0753 ( new_n1096_, new_n1090_, new_n1085_, new_n1095_ );
nand g0754 ( new_n1097_, new_n1090_, new_n1095_ );
nand g0755 ( new_n1098_, new_n1097_, keyIn_0_181 );
nand g0756 ( new_n1099_, new_n685_, N195 );
not g0757 ( new_n1100_, keyIn_0_133 );
not g0758 ( new_n1101_, keyIn_0_109 );
nand g0759 ( new_n1102_, new_n784_, N246 );
nand g0760 ( new_n1103_, new_n1102_, new_n1101_ );
nand g0761 ( new_n1104_, new_n784_, keyIn_0_109, N246 );
nand g0762 ( new_n1105_, new_n1103_, new_n1104_ );
nand g0763 ( new_n1106_, N255, N260 );
nand g0764 ( new_n1107_, new_n1105_, new_n1106_ );
nand g0765 ( new_n1108_, new_n1107_, new_n1100_ );
nand g0766 ( new_n1109_, new_n1105_, keyIn_0_133, new_n1106_ );
nand g0767 ( new_n1110_, new_n1108_, new_n1109_ );
nand g0768 ( new_n1111_, new_n1098_, new_n1096_, new_n1099_, new_n1110_ );
not g0769 ( new_n1112_, new_n1111_ );
nand g0770 ( new_n1113_, new_n1084_, new_n1081_, new_n1112_ );
nand g0771 ( new_n1114_, new_n1113_, keyIn_0_223 );
not g0772 ( new_n1115_, keyIn_0_223 );
nand g0773 ( new_n1116_, new_n1084_, new_n1115_, new_n1081_, new_n1112_ );
nand g0774 ( new_n1117_, new_n1114_, new_n1116_ );
nand g0775 ( new_n1118_, new_n1117_, keyIn_0_232 );
not g0776 ( new_n1119_, keyIn_0_232 );
nand g0777 ( new_n1120_, new_n1114_, new_n1119_, new_n1116_ );
nand g0778 ( new_n1121_, new_n1118_, new_n1120_ );
nand g0779 ( new_n1122_, new_n1121_, new_n1038_ );
nand g0780 ( new_n1123_, new_n1118_, keyIn_0_240, new_n1120_ );
nand g0781 ( N865, new_n1122_, new_n1123_ );
not g0782 ( new_n1125_, keyIn_0_241 );
not g0783 ( new_n1126_, keyIn_0_192 );
nand g0784 ( new_n1127_, new_n819_, new_n855_ );
nand g0785 ( new_n1128_, new_n1127_, keyIn_0_191 );
not g0786 ( new_n1129_, keyIn_0_191 );
nand g0787 ( new_n1130_, new_n819_, new_n1129_, new_n855_ );
nand g0788 ( new_n1131_, new_n1128_, new_n1130_ );
nand g0789 ( new_n1132_, new_n894_, keyIn_0_152 );
not g0790 ( new_n1133_, keyIn_0_152 );
nand g0791 ( new_n1134_, new_n893_, new_n1133_ );
nand g0792 ( new_n1135_, new_n1132_, new_n1134_ );
nand g0793 ( new_n1136_, new_n1131_, new_n1135_ );
nand g0794 ( new_n1137_, new_n1136_, new_n1126_ );
nand g0795 ( new_n1138_, new_n1131_, keyIn_0_192, new_n1135_ );
nand g0796 ( new_n1139_, new_n1137_, new_n1138_ );
not g0797 ( new_n1140_, keyIn_0_93 );
not g0798 ( new_n1141_, keyIn_0_74 );
nand g0799 ( new_n1142_, new_n559_, keyIn_0_53, N96 );
not g0800 ( new_n1143_, keyIn_0_53 );
nand g0801 ( new_n1144_, new_n559_, N96 );
nand g0802 ( new_n1145_, new_n1144_, new_n1143_ );
nand g0803 ( new_n1146_, N51, N138 );
nand g0804 ( new_n1147_, new_n1146_, keyIn_0_9 );
not g0805 ( new_n1148_, keyIn_0_9 );
nand g0806 ( new_n1149_, new_n1148_, N51, N138 );
nand g0807 ( new_n1150_, new_n1147_, new_n1149_ );
not g0808 ( new_n1151_, new_n1150_ );
nand g0809 ( new_n1152_, new_n1145_, new_n1141_, new_n1142_, new_n1151_ );
nand g0810 ( new_n1153_, new_n1145_, new_n1142_, new_n1151_ );
nand g0811 ( new_n1154_, new_n1153_, keyIn_0_74 );
not g0812 ( new_n1155_, keyIn_0_32 );
nand g0813 ( new_n1156_, new_n574_, N17 );
nand g0814 ( new_n1157_, new_n1156_, new_n1155_ );
not g0815 ( new_n1158_, new_n1157_ );
nor g0816 ( new_n1159_, new_n1156_, new_n1155_ );
nor g0817 ( new_n1160_, new_n1158_, new_n1159_ );
nor g0818 ( new_n1161_, new_n1160_, new_n585_ );
not g0819 ( new_n1162_, new_n1161_ );
nand g0820 ( new_n1163_, new_n1162_, keyIn_0_41 );
not g0821 ( new_n1164_, keyIn_0_41 );
nand g0822 ( new_n1165_, new_n1161_, new_n1164_ );
nand g0823 ( new_n1166_, new_n1163_, new_n1165_ );
nand g0824 ( new_n1167_, new_n508_, N55, new_n491_ );
nand g0825 ( new_n1168_, new_n1167_, keyIn_0_31 );
not g0826 ( new_n1169_, keyIn_0_31 );
nand g0827 ( new_n1170_, new_n508_, new_n1169_, N55, new_n491_ );
nand g0828 ( new_n1171_, new_n1168_, new_n1170_ );
not g0829 ( new_n1172_, new_n1171_ );
nand g0830 ( new_n1173_, new_n1172_, N146 );
nand g0831 ( new_n1174_, new_n1173_, keyIn_0_40 );
not g0832 ( new_n1175_, keyIn_0_40 );
nand g0833 ( new_n1176_, new_n1172_, new_n1175_, N146 );
nand g0834 ( new_n1177_, new_n1174_, new_n1176_ );
not g0835 ( new_n1178_, new_n1177_ );
nand g0836 ( new_n1179_, new_n1166_, new_n1178_ );
nand g0837 ( new_n1180_, new_n1179_, keyIn_0_54 );
not g0838 ( new_n1181_, keyIn_0_54 );
nand g0839 ( new_n1182_, new_n1166_, new_n1181_, new_n1178_ );
nand g0840 ( new_n1183_, new_n1180_, new_n1182_ );
not g0841 ( new_n1184_, new_n1183_ );
nand g0842 ( new_n1185_, new_n1184_, new_n1152_, new_n1154_ );
nand g0843 ( new_n1186_, new_n1185_, keyIn_0_82 );
not g0844 ( new_n1187_, keyIn_0_82 );
nand g0845 ( new_n1188_, new_n1184_, new_n1187_, new_n1152_, new_n1154_ );
nand g0846 ( new_n1189_, new_n1186_, new_n1188_ );
not g0847 ( new_n1190_, new_n1189_ );
nand g0848 ( new_n1191_, new_n1190_, new_n436_ );
nand g0849 ( new_n1192_, new_n1191_, new_n1140_ );
nand g0850 ( new_n1193_, new_n1190_, keyIn_0_93, new_n436_ );
nand g0851 ( new_n1194_, new_n1192_, new_n1193_ );
not g0852 ( new_n1195_, keyIn_0_83 );
nand g0853 ( new_n1196_, new_n1162_, keyIn_0_43 );
not g0854 ( new_n1197_, keyIn_0_43 );
nand g0855 ( new_n1198_, new_n1161_, new_n1197_ );
nand g0856 ( new_n1199_, new_n1196_, new_n1198_ );
nand g0857 ( new_n1200_, new_n1172_, N149 );
nand g0858 ( new_n1201_, new_n1200_, keyIn_0_42 );
not g0859 ( new_n1202_, keyIn_0_42 );
nand g0860 ( new_n1203_, new_n1172_, new_n1202_, N149 );
nand g0861 ( new_n1204_, new_n1201_, new_n1203_ );
not g0862 ( new_n1205_, new_n1204_ );
nand g0863 ( new_n1206_, new_n1199_, new_n1205_ );
nand g0864 ( new_n1207_, new_n1206_, keyIn_0_56 );
not g0865 ( new_n1208_, keyIn_0_56 );
nand g0866 ( new_n1209_, new_n1199_, new_n1208_, new_n1205_ );
nand g0867 ( new_n1210_, new_n1207_, new_n1209_ );
not g0868 ( new_n1211_, keyIn_0_75 );
nand g0869 ( new_n1212_, new_n559_, keyIn_0_55, N101 );
nand g0870 ( new_n1213_, N17, N138 );
nand g0871 ( new_n1214_, new_n1213_, keyIn_0_10 );
not g0872 ( new_n1215_, keyIn_0_10 );
nand g0873 ( new_n1216_, new_n1215_, N17, N138 );
nand g0874 ( new_n1217_, new_n1214_, new_n1216_ );
not g0875 ( new_n1218_, keyIn_0_55 );
nand g0876 ( new_n1219_, new_n559_, N101 );
nand g0877 ( new_n1220_, new_n1219_, new_n1218_ );
nand g0878 ( new_n1221_, new_n1220_, new_n1212_, new_n1217_ );
nand g0879 ( new_n1222_, new_n1221_, new_n1211_ );
nand g0880 ( new_n1223_, new_n1220_, keyIn_0_75, new_n1212_, new_n1217_ );
nand g0881 ( new_n1224_, new_n1222_, new_n1223_ );
nand g0882 ( new_n1225_, new_n1210_, new_n1224_ );
nand g0883 ( new_n1226_, new_n1225_, new_n1195_ );
nand g0884 ( new_n1227_, new_n1210_, keyIn_0_83, new_n1224_ );
nand g0885 ( new_n1228_, new_n1226_, new_n1227_ );
nand g0886 ( new_n1229_, new_n1228_, new_n440_ );
nand g0887 ( new_n1230_, new_n1229_, keyIn_0_96 );
not g0888 ( new_n1231_, keyIn_0_96 );
nand g0889 ( new_n1232_, new_n1228_, new_n1231_, new_n440_ );
nand g0890 ( new_n1233_, new_n1230_, new_n1232_ );
nand g0891 ( new_n1234_, new_n1194_, new_n1233_ );
not g0892 ( new_n1235_, keyIn_0_76 );
not g0893 ( new_n1236_, keyIn_0_57 );
nand g0894 ( new_n1237_, new_n559_, N106 );
nand g0895 ( new_n1238_, new_n1237_, new_n1236_ );
nand g0896 ( new_n1239_, new_n559_, keyIn_0_57, N106 );
nand g0897 ( new_n1240_, new_n1238_, new_n1239_ );
not g0898 ( new_n1241_, keyIn_0_11 );
nand g0899 ( new_n1242_, N138, N152 );
nand g0900 ( new_n1243_, new_n1242_, new_n1241_ );
nand g0901 ( new_n1244_, keyIn_0_11, N138, N152 );
nand g0902 ( new_n1245_, new_n1243_, new_n1244_ );
not g0903 ( new_n1246_, new_n1245_ );
nand g0904 ( new_n1247_, new_n1240_, new_n1246_ );
nand g0905 ( new_n1248_, new_n1247_, new_n1235_ );
nand g0906 ( new_n1249_, new_n1240_, keyIn_0_76, new_n1246_ );
nand g0907 ( new_n1250_, new_n1248_, new_n1249_ );
not g0908 ( new_n1251_, keyIn_0_58 );
not g0909 ( new_n1252_, keyIn_0_45 );
nand g0910 ( new_n1253_, new_n1162_, new_n1252_ );
nand g0911 ( new_n1254_, new_n1161_, keyIn_0_45 );
nand g0912 ( new_n1255_, new_n1253_, new_n1254_ );
not g0913 ( new_n1256_, keyIn_0_44 );
nand g0914 ( new_n1257_, new_n1172_, N153 );
nand g0915 ( new_n1258_, new_n1257_, new_n1256_ );
nand g0916 ( new_n1259_, new_n1172_, keyIn_0_44, N153 );
nand g0917 ( new_n1260_, new_n1258_, new_n1259_ );
not g0918 ( new_n1261_, new_n1260_ );
nand g0919 ( new_n1262_, new_n1255_, new_n1261_ );
nand g0920 ( new_n1263_, new_n1262_, new_n1251_ );
nand g0921 ( new_n1264_, new_n1255_, keyIn_0_58, new_n1261_ );
nand g0922 ( new_n1265_, new_n1263_, new_n1264_ );
not g0923 ( new_n1266_, new_n1265_ );
nand g0924 ( new_n1267_, new_n1266_, new_n1250_ );
nand g0925 ( new_n1268_, new_n1267_, keyIn_0_84 );
not g0926 ( new_n1269_, keyIn_0_84 );
nand g0927 ( new_n1270_, new_n1266_, new_n1269_, new_n1250_ );
nand g0928 ( new_n1271_, new_n1268_, new_n1270_ );
not g0929 ( new_n1272_, new_n1271_ );
nand g0930 ( new_n1273_, new_n1272_, new_n441_ );
nand g0931 ( new_n1274_, new_n1273_, keyIn_0_99 );
not g0932 ( new_n1275_, keyIn_0_99 );
nand g0933 ( new_n1276_, new_n1272_, new_n1275_, new_n441_ );
nand g0934 ( new_n1277_, new_n1274_, new_n1276_ );
nor g0935 ( new_n1278_, new_n1234_, new_n1277_ );
nand g0936 ( new_n1279_, new_n1139_, new_n1278_ );
nand g0937 ( new_n1280_, new_n1279_, keyIn_0_205 );
not g0938 ( new_n1281_, keyIn_0_205 );
nand g0939 ( new_n1282_, new_n1139_, new_n1281_, new_n1278_ );
nand g0940 ( new_n1283_, new_n1280_, new_n1282_ );
not g0941 ( new_n1284_, keyIn_0_171 );
not g0942 ( new_n1285_, new_n1234_ );
not g0943 ( new_n1286_, keyIn_0_122 );
not g0944 ( new_n1287_, keyIn_0_98 );
nand g0945 ( new_n1288_, new_n1271_, N177 );
nand g0946 ( new_n1289_, new_n1288_, new_n1287_ );
nand g0947 ( new_n1290_, new_n1271_, keyIn_0_98, N177 );
nand g0948 ( new_n1291_, new_n1289_, new_n1290_ );
nand g0949 ( new_n1292_, new_n1291_, new_n1286_ );
nand g0950 ( new_n1293_, new_n1289_, keyIn_0_122, new_n1290_ );
nand g0951 ( new_n1294_, new_n1292_, new_n1293_ );
not g0952 ( new_n1295_, new_n1294_ );
nand g0953 ( new_n1296_, new_n1285_, new_n1295_ );
nand g0954 ( new_n1297_, new_n1296_, new_n1284_ );
nand g0955 ( new_n1298_, new_n1285_, new_n1295_, keyIn_0_171 );
nand g0956 ( new_n1299_, new_n1297_, new_n1298_ );
not g0957 ( new_n1300_, keyIn_0_92 );
nand g0958 ( new_n1301_, new_n1189_, N165 );
nand g0959 ( new_n1302_, new_n1301_, new_n1300_ );
nand g0960 ( new_n1303_, new_n1189_, keyIn_0_92, N165 );
nand g0961 ( new_n1304_, new_n1302_, new_n1303_ );
nand g0962 ( new_n1305_, new_n1304_, keyIn_0_116 );
not g0963 ( new_n1306_, keyIn_0_116 );
nand g0964 ( new_n1307_, new_n1302_, new_n1306_, new_n1303_ );
nand g0965 ( new_n1308_, new_n1305_, new_n1307_ );
nand g0966 ( new_n1309_, new_n1308_, keyIn_0_143 );
not g0967 ( new_n1310_, keyIn_0_143 );
nand g0968 ( new_n1311_, new_n1305_, new_n1310_, new_n1307_ );
nand g0969 ( new_n1312_, new_n1309_, new_n1311_ );
not g0970 ( new_n1313_, keyIn_0_95 );
not g0971 ( new_n1314_, new_n1228_ );
nand g0972 ( new_n1315_, new_n1314_, N171 );
nand g0973 ( new_n1316_, new_n1315_, new_n1313_ );
nand g0974 ( new_n1317_, new_n1314_, keyIn_0_95, N171 );
nand g0975 ( new_n1318_, new_n1316_, new_n1317_ );
nand g0976 ( new_n1319_, new_n1318_, keyIn_0_119 );
not g0977 ( new_n1320_, keyIn_0_119 );
nand g0978 ( new_n1321_, new_n1316_, new_n1320_, new_n1317_ );
nand g0979 ( new_n1322_, new_n1319_, new_n1321_ );
not g0980 ( new_n1323_, new_n1322_ );
nand g0981 ( new_n1324_, new_n1323_, keyIn_0_170, new_n1194_ );
not g0982 ( new_n1325_, keyIn_0_170 );
nand g0983 ( new_n1326_, new_n1323_, new_n1194_ );
nand g0984 ( new_n1327_, new_n1326_, new_n1325_ );
nand g0985 ( new_n1328_, new_n1327_, new_n1312_, new_n1324_ );
nor g0986 ( new_n1329_, new_n1328_, new_n1299_ );
nand g0987 ( new_n1330_, new_n1283_, new_n1329_ );
nand g0988 ( new_n1331_, new_n1330_, keyIn_0_206 );
not g0989 ( new_n1332_, keyIn_0_206 );
nand g0990 ( new_n1333_, new_n1283_, new_n1332_, new_n1329_ );
nand g0991 ( new_n1334_, new_n1331_, new_n1333_ );
not g0992 ( new_n1335_, new_n1334_ );
not g0993 ( new_n1336_, keyIn_0_90 );
not g0994 ( new_n1337_, keyIn_0_73 );
not g0995 ( new_n1338_, keyIn_0_51 );
nand g0996 ( new_n1339_, new_n559_, N91 );
nand g0997 ( new_n1340_, new_n1339_, new_n1338_ );
nand g0998 ( new_n1341_, new_n559_, keyIn_0_51, N91 );
nand g0999 ( new_n1342_, new_n1340_, new_n1341_ );
not g1000 ( new_n1343_, keyIn_0_7 );
nand g1001 ( new_n1344_, N8, N138 );
nand g1002 ( new_n1345_, new_n1344_, new_n1343_ );
nand g1003 ( new_n1346_, keyIn_0_7, N8, N138 );
nand g1004 ( new_n1347_, new_n1345_, new_n1346_ );
not g1005 ( new_n1348_, new_n1347_ );
nand g1006 ( new_n1349_, new_n1342_, new_n1337_, new_n1348_ );
nand g1007 ( new_n1350_, new_n1342_, new_n1348_ );
nand g1008 ( new_n1351_, new_n1350_, keyIn_0_73 );
not g1009 ( new_n1352_, keyIn_0_39 );
nand g1010 ( new_n1353_, new_n1161_, new_n1352_ );
nand g1011 ( new_n1354_, new_n1162_, keyIn_0_39 );
not g1012 ( new_n1355_, keyIn_0_38 );
nand g1013 ( new_n1356_, new_n1172_, N143 );
nand g1014 ( new_n1357_, new_n1356_, new_n1355_ );
nand g1015 ( new_n1358_, new_n1172_, keyIn_0_38, N143 );
nand g1016 ( new_n1359_, new_n1357_, new_n1358_ );
not g1017 ( new_n1360_, new_n1359_ );
nand g1018 ( new_n1361_, new_n1354_, new_n1353_, new_n1360_ );
nand g1019 ( new_n1362_, new_n1361_, keyIn_0_52 );
not g1020 ( new_n1363_, keyIn_0_52 );
nand g1021 ( new_n1364_, new_n1354_, new_n1363_, new_n1353_, new_n1360_ );
nand g1022 ( new_n1365_, new_n1362_, new_n1364_ );
nand g1023 ( new_n1366_, new_n1365_, new_n1349_, new_n1351_ );
nand g1024 ( new_n1367_, new_n1366_, keyIn_0_81 );
not g1025 ( new_n1368_, keyIn_0_81 );
nand g1026 ( new_n1369_, new_n1365_, new_n1368_, new_n1349_, new_n1351_ );
nand g1027 ( new_n1370_, new_n1367_, new_n1369_ );
nand g1028 ( new_n1371_, new_n1370_, new_n435_ );
nand g1029 ( new_n1372_, new_n1371_, new_n1336_ );
nand g1030 ( new_n1373_, new_n1370_, keyIn_0_90, new_n435_ );
nand g1031 ( new_n1374_, new_n1372_, new_n1373_ );
nand g1032 ( new_n1375_, new_n1335_, keyIn_0_225, new_n1374_ );
not g1033 ( new_n1376_, keyIn_0_140 );
not g1034 ( new_n1377_, new_n1370_ );
nand g1035 ( new_n1378_, new_n1377_, N159 );
nand g1036 ( new_n1379_, new_n1378_, keyIn_0_89 );
not g1037 ( new_n1380_, keyIn_0_89 );
nand g1038 ( new_n1381_, new_n1377_, new_n1380_, N159 );
nand g1039 ( new_n1382_, new_n1379_, new_n1381_ );
not g1040 ( new_n1383_, new_n1382_ );
nand g1041 ( new_n1384_, new_n1383_, keyIn_0_113 );
not g1042 ( new_n1385_, keyIn_0_113 );
nand g1043 ( new_n1386_, new_n1382_, new_n1385_ );
nand g1044 ( new_n1387_, new_n1384_, new_n1386_ );
nand g1045 ( new_n1388_, new_n1387_, new_n1376_ );
nand g1046 ( new_n1389_, new_n1384_, keyIn_0_140, new_n1386_ );
nand g1047 ( new_n1390_, new_n1388_, new_n1389_ );
not g1048 ( new_n1391_, keyIn_0_225 );
nand g1049 ( new_n1392_, new_n1335_, new_n1374_ );
nand g1050 ( new_n1393_, new_n1392_, new_n1391_ );
nand g1051 ( new_n1394_, new_n1393_, new_n1375_, new_n1390_ );
nand g1052 ( new_n1395_, new_n1394_, keyIn_0_233 );
not g1053 ( new_n1396_, keyIn_0_233 );
nand g1054 ( new_n1397_, new_n1393_, new_n1396_, new_n1375_, new_n1390_ );
nand g1055 ( new_n1398_, new_n1395_, new_n1397_ );
nand g1056 ( new_n1399_, new_n1398_, new_n1125_ );
nand g1057 ( new_n1400_, new_n1395_, keyIn_0_241, new_n1397_ );
nand g1058 ( N866, new_n1399_, new_n1400_ );
not g1059 ( new_n1402_, keyIn_0_249 );
not g1060 ( new_n1403_, keyIn_0_245 );
not g1061 ( new_n1404_, keyIn_0_229 );
not g1062 ( new_n1405_, keyIn_0_220 );
not g1063 ( new_n1406_, keyIn_0_198 );
not g1064 ( new_n1407_, keyIn_0_123 );
nor g1065 ( new_n1408_, new_n1277_, new_n1291_ );
not g1066 ( new_n1409_, new_n1408_ );
nand g1067 ( new_n1410_, new_n1409_, new_n1407_ );
nand g1068 ( new_n1411_, new_n1408_, keyIn_0_123 );
nand g1069 ( new_n1412_, new_n1410_, new_n1411_ );
not g1070 ( new_n1413_, new_n1412_ );
nand g1071 ( new_n1414_, new_n1139_, new_n1413_ );
nand g1072 ( new_n1415_, new_n1414_, new_n1406_ );
nand g1073 ( new_n1416_, new_n1139_, keyIn_0_198, new_n1413_ );
nand g1074 ( new_n1417_, new_n1415_, new_n1416_ );
not g1075 ( new_n1418_, new_n1139_ );
nand g1076 ( new_n1419_, new_n1418_, new_n1412_ );
nand g1077 ( new_n1420_, new_n1419_, keyIn_0_197 );
not g1078 ( new_n1421_, keyIn_0_197 );
nand g1079 ( new_n1422_, new_n1418_, new_n1421_, new_n1412_ );
nand g1080 ( new_n1423_, new_n1420_, new_n1422_ );
not g1081 ( new_n1424_, new_n1423_ );
nand g1082 ( new_n1425_, new_n1424_, keyIn_0_209, new_n1417_ );
not g1083 ( new_n1426_, keyIn_0_209 );
nand g1084 ( new_n1427_, new_n1424_, new_n1417_ );
nand g1085 ( new_n1428_, new_n1427_, new_n1426_ );
nand g1086 ( new_n1429_, new_n1428_, N219, new_n1425_ );
nand g1087 ( new_n1430_, new_n1429_, new_n1405_ );
nand g1088 ( new_n1431_, new_n1428_, keyIn_0_220, N219, new_n1425_ );
nand g1089 ( new_n1432_, new_n1430_, new_n1431_ );
nand g1090 ( new_n1433_, N101, N210 );
nand g1091 ( new_n1434_, new_n1432_, new_n1404_, new_n1433_ );
nand g1092 ( new_n1435_, new_n1432_, new_n1433_ );
nand g1093 ( new_n1436_, new_n1435_, keyIn_0_229 );
not g1094 ( new_n1437_, keyIn_0_175 );
nand g1095 ( new_n1438_, new_n1413_, keyIn_0_150, N228 );
not g1096 ( new_n1439_, keyIn_0_151 );
nand g1097 ( new_n1440_, new_n1295_, N237 );
nand g1098 ( new_n1441_, new_n1440_, new_n1439_ );
nand g1099 ( new_n1442_, new_n1295_, keyIn_0_151, N237 );
nand g1100 ( new_n1443_, new_n1441_, new_n1442_ );
not g1101 ( new_n1444_, keyIn_0_150 );
nand g1102 ( new_n1445_, new_n1413_, N228 );
nand g1103 ( new_n1446_, new_n1445_, new_n1444_ );
nand g1104 ( new_n1447_, new_n1446_, new_n1438_, new_n1443_ );
nand g1105 ( new_n1448_, new_n1447_, new_n1437_ );
nand g1106 ( new_n1449_, new_n1446_, keyIn_0_175, new_n1438_, new_n1443_ );
nand g1107 ( new_n1450_, new_n1448_, new_n1449_ );
not g1108 ( new_n1451_, keyIn_0_124 );
not g1109 ( new_n1452_, keyIn_0_100 );
nand g1110 ( new_n1453_, new_n1271_, new_n1452_, N246 );
nand g1111 ( new_n1454_, new_n1271_, N246 );
nand g1112 ( new_n1455_, new_n1454_, keyIn_0_100 );
nand g1113 ( new_n1456_, new_n685_, N177 );
nand g1114 ( new_n1457_, new_n1456_, keyIn_0_70 );
not g1115 ( new_n1458_, keyIn_0_70 );
nand g1116 ( new_n1459_, new_n685_, new_n1458_, N177 );
nand g1117 ( new_n1460_, new_n1457_, new_n1459_ );
not g1118 ( new_n1461_, new_n1460_ );
nand g1119 ( new_n1462_, new_n1455_, new_n1453_, new_n1461_ );
nand g1120 ( new_n1463_, new_n1462_, new_n1451_ );
nand g1121 ( new_n1464_, new_n1455_, keyIn_0_124, new_n1453_, new_n1461_ );
nand g1122 ( new_n1465_, new_n1463_, new_n1464_ );
nand g1123 ( new_n1466_, new_n1450_, new_n1465_ );
not g1124 ( new_n1467_, new_n1466_ );
nand g1125 ( new_n1468_, new_n1436_, new_n1434_, new_n1467_ );
nand g1126 ( new_n1469_, new_n1468_, keyIn_0_237 );
not g1127 ( new_n1470_, keyIn_0_237 );
nand g1128 ( new_n1471_, new_n1436_, new_n1470_, new_n1434_, new_n1467_ );
nand g1129 ( new_n1472_, new_n1469_, new_n1471_ );
nand g1130 ( new_n1473_, new_n1472_, new_n1403_ );
nand g1131 ( new_n1474_, new_n1469_, keyIn_0_245, new_n1471_ );
nand g1132 ( new_n1475_, new_n1473_, new_n1474_ );
nand g1133 ( new_n1476_, new_n1475_, new_n1402_ );
nand g1134 ( new_n1477_, new_n1473_, keyIn_0_249, new_n1474_ );
nand g1135 ( new_n1478_, new_n1476_, new_n1477_ );
not g1136 ( N874, new_n1478_ );
not g1137 ( new_n1480_, keyIn_0_250 );
not g1138 ( new_n1481_, keyIn_0_234 );
not g1139 ( new_n1482_, keyIn_0_226 );
not g1140 ( new_n1483_, keyIn_0_114 );
nand g1141 ( new_n1484_, new_n1383_, new_n1374_ );
nand g1142 ( new_n1485_, new_n1484_, new_n1483_ );
nand g1143 ( new_n1486_, new_n1383_, keyIn_0_114, new_n1374_ );
nand g1144 ( new_n1487_, new_n1485_, new_n1486_ );
not g1145 ( new_n1488_, new_n1487_ );
nand g1146 ( new_n1489_, new_n1334_, new_n1488_ );
nand g1147 ( new_n1490_, new_n1489_, keyIn_0_214 );
not g1148 ( new_n1491_, keyIn_0_214 );
nand g1149 ( new_n1492_, new_n1334_, new_n1491_, new_n1488_ );
nand g1150 ( new_n1493_, new_n1331_, new_n1333_, new_n1487_ );
nand g1151 ( new_n1494_, new_n1493_, keyIn_0_215 );
not g1152 ( new_n1495_, keyIn_0_215 );
nand g1153 ( new_n1496_, new_n1331_, new_n1495_, new_n1333_, new_n1487_ );
nand g1154 ( new_n1497_, new_n1494_, new_n1496_ );
not g1155 ( new_n1498_, new_n1497_ );
nand g1156 ( new_n1499_, new_n1498_, new_n1482_, new_n1490_, new_n1492_ );
nand g1157 ( new_n1500_, new_n1490_, new_n1492_, new_n1494_, new_n1496_ );
nand g1158 ( new_n1501_, new_n1500_, keyIn_0_226 );
nand g1159 ( new_n1502_, new_n1499_, new_n1501_, new_n1481_, N219 );
nand g1160 ( new_n1503_, new_n1499_, new_n1501_, N219 );
nand g1161 ( new_n1504_, new_n1503_, keyIn_0_234 );
nand g1162 ( new_n1505_, new_n588_, N210 );
nand g1163 ( new_n1506_, new_n1505_, keyIn_0_29 );
not g1164 ( new_n1507_, keyIn_0_29 );
nand g1165 ( new_n1508_, new_n588_, new_n1507_, N210 );
nand g1166 ( new_n1509_, new_n1506_, new_n1508_ );
not g1167 ( new_n1510_, new_n1509_ );
nand g1168 ( new_n1511_, new_n1504_, new_n1502_, new_n1510_ );
nand g1169 ( new_n1512_, new_n1511_, keyIn_0_242 );
not g1170 ( new_n1513_, keyIn_0_242 );
nand g1171 ( new_n1514_, new_n1504_, new_n1513_, new_n1502_, new_n1510_ );
nand g1172 ( new_n1515_, new_n1512_, new_n1514_ );
not g1173 ( new_n1516_, keyIn_0_172 );
not g1174 ( new_n1517_, keyIn_0_141 );
nand g1175 ( new_n1518_, new_n1487_, N228 );
nand g1176 ( new_n1519_, new_n1518_, new_n1517_ );
nand g1177 ( new_n1520_, new_n1487_, keyIn_0_141, N228 );
nand g1178 ( new_n1521_, new_n1519_, new_n1520_ );
nand g1179 ( new_n1522_, new_n1387_, N237 );
nand g1180 ( new_n1523_, new_n1522_, keyIn_0_142 );
not g1181 ( new_n1524_, keyIn_0_142 );
nand g1182 ( new_n1525_, new_n1387_, new_n1524_, N237 );
nand g1183 ( new_n1526_, new_n1523_, new_n1525_ );
not g1184 ( new_n1527_, new_n1526_ );
nand g1185 ( new_n1528_, new_n1521_, new_n1527_ );
nand g1186 ( new_n1529_, new_n1528_, new_n1516_ );
nand g1187 ( new_n1530_, new_n1521_, keyIn_0_172, new_n1527_ );
nand g1188 ( new_n1531_, new_n1529_, new_n1530_ );
not g1189 ( new_n1532_, keyIn_0_91 );
nand g1190 ( new_n1533_, new_n1377_, new_n1532_, N246 );
nand g1191 ( new_n1534_, new_n685_, N159 );
nand g1192 ( new_n1535_, new_n1534_, keyIn_0_67 );
not g1193 ( new_n1536_, keyIn_0_67 );
nand g1194 ( new_n1537_, new_n685_, new_n1536_, N159 );
nand g1195 ( new_n1538_, new_n1535_, new_n1537_ );
nand g1196 ( new_n1539_, new_n1377_, N246 );
nand g1197 ( new_n1540_, new_n1539_, keyIn_0_91 );
nand g1198 ( new_n1541_, new_n1540_, new_n1533_, new_n1538_ );
nand g1199 ( new_n1542_, new_n1541_, keyIn_0_115 );
not g1200 ( new_n1543_, keyIn_0_115 );
nand g1201 ( new_n1544_, new_n1540_, new_n1543_, new_n1533_, new_n1538_ );
nand g1202 ( new_n1545_, new_n1542_, new_n1544_ );
nand g1203 ( new_n1546_, new_n1531_, new_n1545_ );
not g1204 ( new_n1547_, new_n1546_ );
nand g1205 ( new_n1548_, new_n1515_, new_n1547_ );
nand g1206 ( new_n1549_, new_n1548_, keyIn_0_246 );
not g1207 ( new_n1550_, keyIn_0_246 );
nand g1208 ( new_n1551_, new_n1515_, new_n1550_, new_n1547_ );
nand g1209 ( new_n1552_, new_n1549_, new_n1551_ );
nand g1210 ( new_n1553_, new_n1552_, new_n1480_ );
nand g1211 ( new_n1554_, new_n1549_, keyIn_0_250, new_n1551_ );
nand g1212 ( new_n1555_, new_n1553_, new_n1554_ );
nand g1213 ( new_n1556_, new_n1555_, keyIn_0_253 );
not g1214 ( new_n1557_, keyIn_0_253 );
nand g1215 ( new_n1558_, new_n1553_, new_n1557_, new_n1554_ );
nand g1216 ( N878, new_n1556_, new_n1558_ );
not g1217 ( new_n1560_, keyIn_0_251 );
not g1218 ( new_n1561_, keyIn_0_117 );
nand g1219 ( new_n1562_, new_n1194_, new_n1304_ );
nand g1220 ( new_n1563_, new_n1562_, new_n1561_ );
nand g1221 ( new_n1564_, new_n1194_, keyIn_0_117, new_n1304_ );
nand g1222 ( new_n1565_, new_n1563_, new_n1564_ );
not g1223 ( new_n1566_, keyIn_0_204 );
not g1224 ( new_n1567_, new_n1233_ );
nor g1225 ( new_n1568_, new_n1277_, new_n1567_ );
nand g1226 ( new_n1569_, new_n1139_, new_n1566_, new_n1568_ );
nand g1227 ( new_n1570_, new_n1139_, new_n1568_ );
nand g1228 ( new_n1571_, new_n1570_, keyIn_0_204 );
nand g1229 ( new_n1572_, new_n1295_, keyIn_0_169, new_n1233_ );
not g1230 ( new_n1573_, keyIn_0_169 );
nand g1231 ( new_n1574_, new_n1295_, new_n1233_ );
nand g1232 ( new_n1575_, new_n1574_, new_n1573_ );
nand g1233 ( new_n1576_, new_n1323_, keyIn_0_146 );
not g1234 ( new_n1577_, keyIn_0_146 );
nand g1235 ( new_n1578_, new_n1322_, new_n1577_ );
nand g1236 ( new_n1579_, new_n1575_, new_n1572_, new_n1576_, new_n1578_ );
not g1237 ( new_n1580_, new_n1579_ );
nand g1238 ( new_n1581_, new_n1571_, new_n1569_, new_n1580_ );
nand g1239 ( new_n1582_, new_n1581_, keyIn_0_207 );
not g1240 ( new_n1583_, keyIn_0_207 );
nand g1241 ( new_n1584_, new_n1571_, new_n1583_, new_n1569_, new_n1580_ );
nand g1242 ( new_n1585_, new_n1582_, new_n1565_, new_n1584_ );
nand g1243 ( new_n1586_, new_n1585_, keyIn_0_216 );
not g1244 ( new_n1587_, keyIn_0_216 );
nand g1245 ( new_n1588_, new_n1582_, new_n1587_, new_n1565_, new_n1584_ );
nand g1246 ( new_n1589_, new_n1586_, new_n1588_ );
not g1247 ( new_n1590_, keyIn_0_217 );
not g1248 ( new_n1591_, new_n1565_ );
nand g1249 ( new_n1592_, new_n1582_, new_n1584_ );
nand g1250 ( new_n1593_, new_n1592_, new_n1591_ );
nand g1251 ( new_n1594_, new_n1593_, new_n1590_ );
nand g1252 ( new_n1595_, new_n1592_, keyIn_0_217, new_n1591_ );
nand g1253 ( new_n1596_, new_n1589_, new_n1594_, new_n1595_ );
nand g1254 ( new_n1597_, new_n1596_, keyIn_0_227 );
not g1255 ( new_n1598_, keyIn_0_227 );
nand g1256 ( new_n1599_, new_n1589_, new_n1594_, new_n1598_, new_n1595_ );
nand g1257 ( new_n1600_, new_n1597_, new_n1599_ );
nand g1258 ( new_n1601_, new_n1600_, keyIn_0_235, N219 );
not g1259 ( new_n1602_, keyIn_0_15 );
nand g1260 ( new_n1603_, N91, N210 );
nand g1261 ( new_n1604_, new_n1603_, new_n1602_ );
nand g1262 ( new_n1605_, keyIn_0_15, N91, N210 );
nand g1263 ( new_n1606_, new_n1604_, new_n1605_ );
not g1264 ( new_n1607_, keyIn_0_235 );
nand g1265 ( new_n1608_, new_n1600_, N219 );
nand g1266 ( new_n1609_, new_n1608_, new_n1607_ );
nand g1267 ( new_n1610_, new_n1609_, keyIn_0_243, new_n1601_, new_n1606_ );
not g1268 ( new_n1611_, keyIn_0_243 );
nand g1269 ( new_n1612_, new_n1609_, new_n1601_, new_n1606_ );
nand g1270 ( new_n1613_, new_n1612_, new_n1611_ );
not g1271 ( new_n1614_, keyIn_0_144 );
nand g1272 ( new_n1615_, new_n1591_, new_n1614_, N228 );
nand g1273 ( new_n1616_, new_n1591_, N228 );
nand g1274 ( new_n1617_, new_n1616_, keyIn_0_144 );
nand g1275 ( new_n1618_, new_n1308_, N237 );
nand g1276 ( new_n1619_, new_n1618_, keyIn_0_145 );
not g1277 ( new_n1620_, keyIn_0_145 );
nand g1278 ( new_n1621_, new_n1308_, new_n1620_, N237 );
nand g1279 ( new_n1622_, new_n1617_, new_n1615_, new_n1619_, new_n1621_ );
nor g1280 ( new_n1623_, new_n1622_, keyIn_0_173 );
nand g1281 ( new_n1624_, new_n1622_, keyIn_0_173 );
nand g1282 ( new_n1625_, new_n1189_, N246 );
nand g1283 ( new_n1626_, new_n1625_, keyIn_0_94 );
not g1284 ( new_n1627_, keyIn_0_94 );
nand g1285 ( new_n1628_, new_n1189_, new_n1627_, N246 );
nand g1286 ( new_n1629_, new_n1626_, new_n1628_ );
nand g1287 ( new_n1630_, new_n685_, N165 );
nand g1288 ( new_n1631_, new_n1630_, keyIn_0_68 );
not g1289 ( new_n1632_, keyIn_0_68 );
nand g1290 ( new_n1633_, new_n685_, new_n1632_, N165 );
nand g1291 ( new_n1634_, new_n1631_, new_n1633_ );
nand g1292 ( new_n1635_, new_n1629_, new_n1634_ );
nand g1293 ( new_n1636_, new_n1635_, keyIn_0_118 );
not g1294 ( new_n1637_, keyIn_0_118 );
nand g1295 ( new_n1638_, new_n1629_, new_n1637_, new_n1634_ );
nand g1296 ( new_n1639_, new_n1624_, new_n1636_, new_n1638_ );
nor g1297 ( new_n1640_, new_n1639_, new_n1623_ );
nand g1298 ( new_n1641_, new_n1613_, new_n1610_, new_n1640_ );
nand g1299 ( new_n1642_, new_n1641_, keyIn_0_247 );
not g1300 ( new_n1643_, keyIn_0_247 );
nand g1301 ( new_n1644_, new_n1613_, new_n1643_, new_n1610_, new_n1640_ );
nand g1302 ( new_n1645_, new_n1642_, new_n1644_ );
nand g1303 ( new_n1646_, new_n1645_, new_n1560_ );
nand g1304 ( new_n1647_, new_n1642_, keyIn_0_251, new_n1644_ );
nand g1305 ( new_n1648_, new_n1646_, new_n1647_ );
nand g1306 ( new_n1649_, new_n1648_, keyIn_0_254 );
not g1307 ( new_n1650_, keyIn_0_254 );
nand g1308 ( new_n1651_, new_n1646_, new_n1650_, new_n1647_ );
nand g1309 ( new_n1652_, new_n1649_, new_n1651_ );
not g1310 ( N879, new_n1652_ );
not g1311 ( new_n1654_, keyIn_0_252 );
not g1312 ( new_n1655_, keyIn_0_248 );
not g1313 ( new_n1656_, keyIn_0_244 );
not g1314 ( new_n1657_, keyIn_0_236 );
not g1315 ( new_n1658_, keyIn_0_228 );
not g1316 ( new_n1659_, keyIn_0_120 );
nand g1317 ( new_n1660_, new_n1318_, new_n1233_ );
nand g1318 ( new_n1661_, new_n1660_, new_n1659_ );
nand g1319 ( new_n1662_, new_n1318_, keyIn_0_120, new_n1233_ );
nand g1320 ( new_n1663_, new_n1661_, new_n1662_ );
not g1321 ( new_n1664_, new_n1663_ );
not g1322 ( new_n1665_, keyIn_0_208 );
not g1323 ( new_n1666_, keyIn_0_203 );
not g1324 ( new_n1667_, new_n1277_ );
nand g1325 ( new_n1668_, new_n1139_, new_n1666_, new_n1667_ );
nand g1326 ( new_n1669_, new_n1139_, new_n1667_ );
nand g1327 ( new_n1670_, new_n1669_, keyIn_0_203 );
not g1328 ( new_n1671_, keyIn_0_149 );
nand g1329 ( new_n1672_, new_n1295_, new_n1671_ );
nand g1330 ( new_n1673_, new_n1294_, keyIn_0_149 );
nand g1331 ( new_n1674_, new_n1672_, new_n1673_ );
not g1332 ( new_n1675_, new_n1674_ );
nand g1333 ( new_n1676_, new_n1670_, new_n1668_, new_n1675_ );
nand g1334 ( new_n1677_, new_n1676_, new_n1665_ );
nand g1335 ( new_n1678_, new_n1670_, keyIn_0_208, new_n1668_, new_n1675_ );
nand g1336 ( new_n1679_, new_n1677_, new_n1678_ );
nand g1337 ( new_n1680_, new_n1679_, new_n1664_ );
nand g1338 ( new_n1681_, new_n1680_, keyIn_0_219 );
not g1339 ( new_n1682_, keyIn_0_219 );
nand g1340 ( new_n1683_, new_n1679_, new_n1682_, new_n1664_ );
nand g1341 ( new_n1684_, new_n1681_, new_n1683_ );
nand g1342 ( new_n1685_, new_n1677_, new_n1663_, new_n1678_ );
nand g1343 ( new_n1686_, new_n1685_, keyIn_0_218 );
not g1344 ( new_n1687_, keyIn_0_218 );
nand g1345 ( new_n1688_, new_n1677_, new_n1687_, new_n1663_, new_n1678_ );
nand g1346 ( new_n1689_, new_n1686_, new_n1688_ );
not g1347 ( new_n1690_, new_n1689_ );
nand g1348 ( new_n1691_, new_n1690_, new_n1684_ );
nand g1349 ( new_n1692_, new_n1691_, new_n1658_ );
nand g1350 ( new_n1693_, new_n1690_, new_n1684_, keyIn_0_228 );
nand g1351 ( new_n1694_, new_n1692_, new_n1657_, N219, new_n1693_ );
nand g1352 ( new_n1695_, N96, N210 );
nand g1353 ( new_n1696_, new_n1692_, N219, new_n1693_ );
nand g1354 ( new_n1697_, new_n1696_, keyIn_0_236 );
nand g1355 ( new_n1698_, new_n1697_, new_n1656_, new_n1694_, new_n1695_ );
nand g1356 ( new_n1699_, new_n1697_, new_n1694_, new_n1695_ );
nand g1357 ( new_n1700_, new_n1699_, keyIn_0_244 );
not g1358 ( new_n1701_, keyIn_0_174 );
not g1359 ( new_n1702_, keyIn_0_147 );
nand g1360 ( new_n1703_, new_n1664_, N228 );
nand g1361 ( new_n1704_, new_n1703_, new_n1702_ );
nand g1362 ( new_n1705_, new_n1664_, keyIn_0_147, N228 );
nand g1363 ( new_n1706_, new_n1704_, new_n1705_ );
nand g1364 ( new_n1707_, new_n1323_, N237 );
nand g1365 ( new_n1708_, new_n1707_, keyIn_0_148 );
not g1366 ( new_n1709_, keyIn_0_148 );
nand g1367 ( new_n1710_, new_n1323_, new_n1709_, N237 );
nand g1368 ( new_n1711_, new_n1708_, new_n1710_ );
not g1369 ( new_n1712_, new_n1711_ );
nand g1370 ( new_n1713_, new_n1706_, new_n1712_ );
nand g1371 ( new_n1714_, new_n1713_, new_n1701_ );
nand g1372 ( new_n1715_, new_n1706_, keyIn_0_174, new_n1712_ );
nand g1373 ( new_n1716_, new_n1714_, new_n1715_ );
not g1374 ( new_n1717_, keyIn_0_121 );
not g1375 ( new_n1718_, keyIn_0_97 );
nand g1376 ( new_n1719_, new_n1314_, new_n1718_, N246 );
nand g1377 ( new_n1720_, new_n685_, N171 );
nand g1378 ( new_n1721_, new_n1720_, keyIn_0_69 );
not g1379 ( new_n1722_, keyIn_0_69 );
nand g1380 ( new_n1723_, new_n685_, new_n1722_, N171 );
nand g1381 ( new_n1724_, new_n1721_, new_n1723_ );
nand g1382 ( new_n1725_, new_n1314_, N246 );
nand g1383 ( new_n1726_, new_n1725_, keyIn_0_97 );
nand g1384 ( new_n1727_, new_n1726_, new_n1719_, new_n1724_ );
nand g1385 ( new_n1728_, new_n1727_, new_n1717_ );
nand g1386 ( new_n1729_, new_n1726_, keyIn_0_121, new_n1719_, new_n1724_ );
nand g1387 ( new_n1730_, new_n1716_, new_n1728_, new_n1729_ );
not g1388 ( new_n1731_, new_n1730_ );
nand g1389 ( new_n1732_, new_n1700_, new_n1698_, new_n1731_ );
nand g1390 ( new_n1733_, new_n1732_, new_n1655_ );
nand g1391 ( new_n1734_, new_n1700_, keyIn_0_248, new_n1698_, new_n1731_ );
nand g1392 ( new_n1735_, new_n1733_, new_n1734_ );
nand g1393 ( new_n1736_, new_n1735_, new_n1654_ );
nand g1394 ( new_n1737_, new_n1733_, keyIn_0_252, new_n1734_ );
nand g1395 ( new_n1738_, new_n1736_, new_n1737_ );
nand g1396 ( new_n1739_, new_n1738_, keyIn_0_255 );
not g1397 ( new_n1740_, keyIn_0_255 );
nand g1398 ( new_n1741_, new_n1736_, new_n1740_, new_n1737_ );
nand g1399 ( new_n1742_, new_n1739_, new_n1741_ );
not g1400 ( N880, new_n1742_ );
endmodule