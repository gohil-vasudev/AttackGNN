module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX646, WX647, n3527, WX648,
         WX649, n3525, WX650, WX652, WX653, n3521, WX654, WX655, n3519, WX656,
         WX657, n3517, WX658, WX659, WX660, WX661, n3513, WX662, WX663, n3511,
         WX664, WX665, n3509, WX666, WX667, WX668, WX669, n3505, WX670, WX671,
         n3503, WX672, WX673, n3501, WX674, WX675, WX676, WX677, n3497, WX678,
         WX679, n3495, WX680, WX681, n3493, WX682, WX683, n3491, WX684, WX685,
         n3489, WX686, WX688, WX689, n3485, WX690, WX691, n3483, WX692, WX693,
         n3481, WX694, WX695, n3479, WX696, WX697, n3477, WX698, WX699, n3475,
         WX700, WX701, n3473, WX702, WX703, n3471, WX704, WX705, n3469, WX706,
         WX707, n3467, WX708, WX709, WX710, WX711, WX712, WX713, WX714, WX715,
         WX716, WX717, WX718, WX719, WX720, WX721, WX722, WX724, WX725, WX726,
         WX727, WX728, WX729, WX730, WX731, WX732, WX733, WX734, WX735, WX736,
         WX737, WX738, WX739, WX740, WX741, WX742, WX743, WX744, WX745, WX746,
         WX747, WX748, WX749, WX750, WX751, WX752, WX753, WX754, WX755, WX756,
         WX757, WX758, WX760, WX761, WX762, WX763, WX764, WX765, WX766, WX767,
         WX768, WX769, WX770, WX771, WX772, WX773, WX774, WX775, WX776, WX777,
         WX778, WX779, WX780, WX781, WX782, WX783, WX784, WX785, WX786, WX787,
         WX788, WX789, WX790, WX791, WX792, WX793, WX794, WX796, WX797, WX798,
         WX799, WX800, WX801, WX802, WX803, WX804, WX805, WX806, WX807, WX808,
         WX809, WX810, WX811, WX812, WX813, WX814, WX815, WX816, WX817, WX818,
         WX819, WX820, WX821, WX822, WX823, WX824, WX825, WX826, WX827, WX828,
         WX829, WX830, WX832, WX833, WX834, WX835, WX836, WX837, WX838, WX839,
         WX840, WX841, WX842, WX843, WX844, WX845, WX846, WX847, WX848, WX849,
         WX850, WX851, WX852, WX853, WX854, WX855, WX856, WX857, WX858, WX859,
         WX860, WX861, WX862, WX863, WX864, WX865, WX866, WX868, WX869, WX870,
         WX871, WX872, WX873, WX874, WX875, WX876, WX877, WX878, WX879, WX880,
         WX881, WX882, WX883, WX884, WX885, WX886, WX887, WX888, WX889, WX890,
         WX891, WX892, WX893, WX894, WX895, WX896, WX897, WX898, WX899, WX1264,
         WX1266, WX1268, WX1270, DFF_163_n1, WX1272, WX1274, WX1276, WX1278,
         WX1280, WX1282, WX1284, DFF_170_n1, WX1286, WX1288, WX1290, WX1292,
         WX1294, WX1296, WX1298, WX1300, WX1302, WX1304, WX1306, WX1308,
         WX1310, WX1312, WX1314, WX1316, WX1318, WX1320, WX1322, WX1324,
         WX1326, DFF_191_n1, WX1778, n8702, n4033, n8701, n4032, n8700, n4031,
         n8699, n4030, n4029, n8696, n4028, n8695, n4027, n8694, n4026, n8693,
         n4025, n8692, n4024, n8691, n4023, n8690, n4022, n8689, n4021, n8688,
         n4020, n8687, n4019, n8686, n4018, n8685, n4017, n8684, n4016, n8683,
         n4015, n8682, n4014, n8681, n4013, n8680, n4012, n4011, n8677, n4010,
         n8676, n4009, n8675, n4008, n8674, n4007, n8673, n4006, n8672, n4005,
         n8671, n4004, WX1839, n8670, n4003, WX1937, n8669, WX1939, n8668,
         WX1941, n8667, WX1943, n8666, WX1945, n8665, WX1947, n8664, WX1949,
         n8663, WX1951, n8662, WX1953, n8661, WX1955, WX1957, n8658, WX1959,
         n8657, WX1961, n8656, WX1963, n8655, WX1965, n8654, WX1967, n8653,
         WX1969, WX1970, WX1971, WX1972, WX1973, WX1974, WX1975, WX1976,
         WX1977, WX1978, WX1979, WX1980, WX1981, WX1982, WX1983, WX1984,
         WX1985, WX1986, WX1987, WX1988, WX1989, WX1990, WX1991, WX1993,
         WX1994, WX1995, WX1996, WX1997, WX1998, WX1999, WX2000, WX2001,
         WX2002, WX2003, WX2004, WX2005, WX2006, WX2007, WX2008, WX2009,
         WX2010, WX2011, WX2012, WX2013, WX2014, WX2015, WX2016, WX2017,
         WX2018, WX2019, WX2020, WX2021, WX2022, WX2023, WX2024, WX2025,
         WX2026, WX2027, WX2029, WX2030, WX2031, WX2032, WX2033, WX2034,
         WX2035, WX2036, n3783, WX2037, WX2038, WX2039, WX2040, WX2041, WX2042,
         WX2043, WX2044, n3775, WX2045, WX2046, WX2047, WX2048, WX2049, WX2050,
         WX2051, WX2052, WX2053, WX2054, WX2055, WX2056, n3763, WX2057, WX2058,
         WX2059, WX2060, WX2061, WX2062, WX2063, WX2065, WX2066, WX2067,
         WX2068, WX2069, WX2070, WX2071, WX2072, WX2073, WX2074, WX2075,
         WX2076, WX2077, WX2078, WX2079, WX2080, WX2081, WX2082, WX2083,
         WX2084, WX2085, WX2086, WX2087, WX2088, WX2089, WX2090, WX2091,
         WX2092, WX2093, WX2094, WX2095, WX2096, WX2097, WX2098, WX2099,
         WX2101, WX2102, WX2103, WX2104, WX2105, WX2106, WX2107, WX2108,
         WX2109, WX2110, WX2111, WX2112, WX2113, WX2114, WX2115, WX2116,
         WX2117, WX2118, WX2119, WX2120, WX2121, WX2122, WX2123, WX2124,
         WX2125, WX2126, WX2127, WX2128, WX2129, WX2130, WX2131, WX2132,
         WX2133, WX2134, WX2135, WX2137, WX2138, WX2139, WX2140, WX2141,
         WX2142, WX2143, WX2144, WX2145, WX2146, WX2147, WX2148, WX2149,
         WX2150, WX2151, WX2152, WX2153, WX2154, WX2155, WX2156, WX2157,
         WX2158, WX2159, WX2160, WX2161, WX2162, WX2163, WX2164, WX2165,
         WX2166, WX2167, WX2168, WX2169, WX2170, WX2171, WX2173, WX2174,
         WX2175, WX2176, WX2177, WX2178, WX2179, WX2180, WX2181, WX2182,
         WX2183, WX2184, WX2185, WX2186, WX2187, WX2188, WX2189, WX2190,
         WX2191, WX2192, WX2557, WX2559, WX2561, WX2563, DFF_355_n1, WX2565,
         WX2567, WX2569, WX2571, WX2573, WX2575, DFF_361_n1, WX2577,
         DFF_362_n1, WX2579, WX2581, WX2583, WX2585, WX2587, DFF_367_n1,
         WX2589, WX2591, WX2593, WX2595, WX2597, WX2599, WX2601, WX2603,
         WX2605, WX2607, WX2609, WX2611, DFF_379_n1, WX2613, WX2615, WX2617,
         WX2619, DFF_383_n1, WX3071, n8644, n4002, n8643, n4001, n8642, n4000,
         n8641, n3999, n8640, n3998, n8639, n3997, n8638, n3996, n8637, n3995,
         n8636, n3994, n8635, n3993, n3992, n8632, n3991, n8631, n3990, n8630,
         n3989, n8629, n3988, n8628, n3987, n8627, n3986, n8626, n3985, n8625,
         n3984, n8624, n3983, n8623, n3982, n8622, n3981, n8621, n3980, n8620,
         n3979, n8619, n3978, n8618, n3977, n8617, n3976, n8616, n3975, n3974,
         n8613, n3973, WX3132, n8612, n3972, WX3230, n8611, WX3232, n8610,
         WX3234, n8609, WX3236, n8608, WX3238, n8607, WX3240, n8606, WX3242,
         n8605, WX3244, n8604, WX3246, n8603, WX3248, n8602, WX3250, n8601,
         WX3252, n8600, WX3254, n8599, WX3256, n8598, WX3258, n8597, WX3260,
         WX3262, WX3263, WX3264, WX3265, WX3266, WX3267, WX3268, WX3269,
         WX3270, WX3271, WX3272, WX3273, WX3274, WX3275, WX3276, WX3277,
         WX3278, WX3279, WX3280, WX3281, WX3282, WX3283, WX3284, WX3285,
         WX3286, WX3287, WX3288, WX3289, WX3290, WX3291, WX3292, WX3293,
         WX3294, WX3295, WX3296, WX3298, WX3299, WX3300, WX3301, WX3302,
         WX3303, WX3304, WX3305, WX3306, WX3307, WX3308, WX3309, WX3310,
         WX3311, WX3312, WX3313, WX3314, WX3315, WX3316, WX3317, WX3318,
         WX3319, WX3320, WX3321, WX3322, WX3323, WX3324, WX3325, WX3326,
         WX3327, WX3328, WX3329, WX3330, WX3331, WX3332, WX3334, WX3335,
         WX3336, WX3337, WX3338, WX3339, WX3340, WX3341, n3739, WX3342, WX3343,
         WX3344, WX3345, n3735, WX3346, WX3347, WX3348, WX3349, WX3350, WX3351,
         WX3352, WX3353, WX3354, WX3355, WX3356, WX3357, WX3358, WX3359,
         WX3360, WX3361, WX3362, WX3363, WX3364, WX3365, WX3366, WX3367,
         WX3368, WX3370, WX3371, WX3372, WX3373, WX3374, WX3375, WX3376,
         WX3377, WX3378, WX3379, WX3380, WX3381, WX3382, WX3383, WX3384,
         WX3385, WX3386, WX3387, WX3388, WX3389, WX3390, WX3391, WX3392,
         WX3393, WX3394, WX3395, WX3396, WX3397, WX3398, WX3399, WX3400,
         WX3401, WX3402, WX3403, WX3404, WX3406, WX3407, WX3408, WX3409,
         WX3410, WX3411, WX3412, WX3413, WX3414, WX3415, WX3416, WX3417,
         WX3418, WX3419, WX3420, WX3421, WX3422, WX3423, WX3424, WX3425,
         WX3426, WX3427, WX3428, WX3429, WX3430, WX3431, WX3432, WX3433,
         WX3434, WX3435, WX3436, WX3437, WX3438, WX3440, WX3441, WX3442,
         WX3443, WX3444, WX3445, WX3446, WX3447, WX3448, WX3449, WX3450,
         WX3451, WX3452, WX3453, WX3454, WX3455, WX3456, WX3457, WX3458,
         WX3459, WX3460, WX3461, WX3462, WX3463, WX3464, WX3465, WX3466,
         WX3467, WX3468, WX3469, WX3470, WX3471, WX3472, WX3474, WX3475,
         WX3476, WX3477, WX3478, WX3479, WX3480, WX3481, WX3482, WX3483,
         WX3484, WX3485, WX3850, WX3852, WX3854, WX3856, DFF_547_n1, WX3858,
         WX3860, DFF_549_n1, WX3862, WX3864, WX3866, WX3868, WX3870, WX3872,
         WX3874, WX3876, WX3878, WX3880, DFF_559_n1, WX3882, WX3884, WX3886,
         WX3888, WX3890, WX3892, WX3894, DFF_566_n1, WX3896, WX3898, WX3900,
         WX3902, WX3904, WX3906, WX3908, WX3910, WX3912, DFF_575_n1, WX4364,
         n8586, n3971, n8585, n3970, n8584, n3969, n8583, n3968, n8582, n3967,
         n8581, n3966, n8580, n3965, n8579, n3964, n8578, n3963, n8577, n3962,
         n8576, n3961, n3960, n8573, n3959, n8572, n3958, n8571, n3957, n8570,
         n3956, n8569, n3955, n8568, n3954, n8567, n3953, n8566, n3952, n8565,
         n3951, n8564, n3950, n8563, n3949, n8562, n3948, n8561, n3947, n8560,
         n3946, n8559, n3945, n8558, n3944, n3943, n8555, n3942, WX4425, n8554,
         n3941, WX4523, n8553, WX4525, n8552, WX4527, n8551, WX4529, n8550,
         WX4531, n8549, WX4533, n8548, WX4535, n8547, WX4537, n8546, WX4539,
         n8545, WX4541, n8544, WX4543, n8543, WX4545, n8542, WX4547, n8541,
         WX4549, n8540, WX4551, WX4553, n8537, WX4555, WX4556, WX4557, WX4558,
         WX4559, WX4560, WX4561, WX4562, WX4563, WX4564, WX4565, WX4566,
         WX4567, WX4568, WX4569, WX4570, WX4571, WX4572, WX4573, WX4574,
         WX4575, WX4576, WX4577, WX4578, WX4579, WX4580, WX4581, WX4582,
         WX4583, WX4584, WX4585, WX4587, WX4588, WX4589, WX4590, WX4591,
         WX4592, WX4593, WX4594, WX4595, WX4596, WX4597, WX4598, WX4599,
         WX4600, WX4601, WX4602, WX4603, WX4604, WX4605, WX4606, WX4607,
         WX4608, WX4609, WX4610, WX4611, WX4612, WX4613, WX4614, WX4615,
         WX4616, WX4617, WX4618, WX4619, WX4621, WX4622, WX4623, WX4624, n3717,
         WX4625, WX4626, WX4627, WX4628, n3713, WX4629, WX4630, WX4631, WX4632,
         WX4633, WX4634, WX4635, WX4636, WX4637, WX4638, WX4639, WX4640,
         WX4641, WX4642, WX4643, WX4644, WX4645, WX4646, WX4647, WX4648,
         WX4649, WX4650, n3691, WX4651, WX4652, WX4653, WX4655, WX4656, WX4657,
         WX4658, WX4659, WX4660, WX4661, WX4662, WX4663, WX4664, WX4665,
         WX4666, WX4667, WX4668, WX4669, WX4670, WX4671, WX4672, WX4673,
         WX4674, WX4675, WX4676, WX4677, WX4678, WX4679, WX4680, WX4681,
         WX4682, WX4683, WX4684, WX4685, WX4686, WX4687, WX4689, WX4690,
         WX4691, WX4692, WX4693, WX4694, WX4695, WX4696, WX4697, WX4698,
         WX4699, WX4700, WX4701, WX4702, WX4703, WX4704, WX4705, WX4706,
         WX4707, WX4708, WX4709, WX4710, WX4711, WX4712, WX4713, WX4714,
         WX4715, WX4716, WX4717, WX4718, WX4719, WX4720, WX4721, WX4723,
         WX4724, WX4725, WX4726, WX4727, WX4728, WX4729, WX4730, WX4731,
         WX4732, WX4733, WX4734, WX4735, WX4736, WX4737, WX4738, WX4739,
         WX4740, WX4741, WX4742, WX4743, WX4744, WX4745, WX4746, WX4747,
         WX4748, WX4749, WX4750, WX4751, WX4752, WX4753, WX4754, WX4755,
         WX4757, WX4758, WX4759, WX4760, WX4761, WX4762, WX4763, WX4764,
         WX4765, WX4766, WX4767, WX4768, WX4769, WX4770, WX4771, WX4772,
         WX4773, WX4774, WX4775, WX4776, WX4777, WX4778, WX5143, WX5145,
         WX5147, WX5149, DFF_739_n1, WX5151, WX5153, WX5155, WX5157, WX5159,
         WX5161, WX5163, WX5165, WX5167, WX5169, WX5171, WX5173, DFF_751_n1,
         WX5175, WX5177, WX5179, WX5181, WX5183, WX5185, WX5187, WX5189,
         WX5191, WX5193, WX5195, WX5197, DFF_763_n1, WX5199, WX5201, WX5203,
         WX5205, DFF_767_n1, WX5657, n8528, n3940, n8527, n3939, n8526, n3938,
         n8525, n3937, n8524, n3936, n8523, n3935, n3934, n8520, n3933, n8519,
         n3932, n8518, n3931, n8517, n3930, n8516, n3929, n8515, n3928, n8514,
         n3927, n8513, n3926, n8512, n3925, n8511, n3924, n8510, n3923, n8509,
         n3922, n8508, n3921, n8507, n3920, n8506, n3919, n8505, n3918, n3917,
         n8502, n3916, n8501, n3915, n8500, n3914, n8499, n3913, n8498, n3912,
         n8497, n3911, WX5718, n8496, n3910, WX5816, n8495, WX5818, n8494,
         WX5820, n8493, WX5822, n8492, WX5824, n8491, WX5826, n8490, WX5828,
         n8489, WX5830, n8488, WX5832, n8487, WX5834, WX5836, n8484, WX5838,
         n8483, WX5840, n8482, WX5842, n8481, WX5844, n8480, WX5846, n8479,
         WX5848, WX5849, WX5850, WX5851, WX5852, WX5853, WX5854, WX5855,
         WX5856, WX5857, WX5858, WX5859, WX5860, WX5861, WX5862, WX5863,
         WX5864, WX5865, WX5866, WX5867, WX5868, WX5870, WX5871, WX5872,
         WX5873, WX5874, WX5875, WX5876, WX5877, WX5878, WX5879, WX5880,
         WX5881, WX5882, WX5883, WX5884, WX5885, WX5886, WX5887, WX5888,
         WX5889, WX5890, WX5891, WX5892, WX5893, WX5894, WX5895, WX5896,
         WX5897, WX5898, WX5899, WX5900, WX5901, WX5902, WX5904, WX5905,
         WX5906, WX5907, WX5908, WX5909, WX5910, WX5911, WX5912, WX5913,
         WX5914, WX5915, WX5916, WX5917, WX5918, WX5919, WX5920, WX5921,
         WX5922, WX5923, WX5924, WX5925, WX5926, WX5927, WX5928, WX5929,
         WX5930, WX5931, WX5932, WX5933, n3669, WX5934, WX5935, WX5936, WX5938,
         WX5939, WX5940, WX5941, n3661, WX5942, WX5943, WX5944, WX5945, WX5946,
         WX5947, WX5948, WX5949, WX5950, WX5951, WX5952, WX5953, WX5954,
         WX5955, WX5956, WX5957, WX5958, WX5959, WX5960, WX5961, WX5962,
         WX5963, WX5964, WX5965, WX5966, WX5967, WX5968, WX5969, WX5970,
         WX5972, WX5973, WX5974, WX5975, WX5976, WX5977, WX5978, WX5979,
         WX5980, WX5981, WX5982, WX5983, WX5984, WX5985, WX5986, WX5987,
         WX5988, WX5989, WX5990, WX5991, WX5992, WX5993, WX5994, WX5995,
         WX5996, WX5997, WX5998, WX5999, WX6000, WX6001, WX6002, WX6003,
         WX6004, WX6006, WX6007, WX6008, WX6009, WX6010, WX6011, WX6012,
         WX6013, WX6014, WX6015, WX6016, WX6017, WX6018, WX6019, WX6020,
         WX6021, WX6022, WX6023, WX6024, WX6025, WX6026, WX6027, WX6028,
         WX6029, WX6030, WX6031, WX6032, WX6033, WX6034, WX6035, WX6036,
         WX6037, WX6038, WX6040, WX6041, WX6042, WX6043, WX6044, WX6045,
         WX6046, WX6047, WX6048, WX6049, WX6050, WX6051, WX6052, WX6053,
         WX6054, WX6055, WX6056, WX6057, WX6058, WX6059, WX6060, WX6061,
         WX6062, WX6063, WX6064, WX6065, WX6066, WX6067, WX6068, WX6069,
         WX6070, WX6071, WX6436, WX6438, WX6440, WX6442, DFF_931_n1, WX6444,
         WX6446, WX6448, WX6450, WX6452, WX6454, WX6456, DFF_938_n1, WX6458,
         WX6460, WX6462, WX6464, WX6466, WX6468, WX6470, WX6472, WX6474,
         WX6476, WX6478, WX6480, WX6482, WX6484, WX6486, WX6488, WX6490,
         WX6492, WX6494, WX6496, WX6498, DFF_959_n1, WX6950, n8470, n3909,
         n3908, n8467, n3907, n8466, n3906, n8465, n3905, n8464, n3904, n8463,
         n3903, n8462, n3902, n8461, n3901, n8460, n3900, n8459, n3899, n8458,
         n3898, n8457, n3897, n8456, n3896, n8455, n3895, n8454, n3894, n8453,
         n3893, n8452, n3892, n3891, n8449, n3890, n8448, n3889, n8447, n3888,
         n8446, n3887, n8445, n3886, WX6999, n8444, n3885, n8443, n8442, n3883,
         n8441, n3882, n8440, n3881, n8439, n3880, WX7011, n8438, n3879,
         WX7109, n8437, WX7111, n8436, WX7113, n8435, WX7115, n8434, WX7117,
         WX7119, n8431, WX7121, n8430, WX7123, n8429, WX7125, n8428, WX7127,
         n8427, WX7129, n8426, WX7131, n8425, WX7133, n8424, WX7135, n8423,
         WX7137, n8422, WX7139, n8421, WX7141, WX7142, WX7143, WX7144, WX7145,
         WX7146, WX7147, WX7148, WX7149, WX7150, WX7151, WX7153, WX7154,
         WX7155, WX7156, WX7157, WX7158, WX7159, WX7160, WX7161, WX7162,
         WX7163, WX7164, WX7165, WX7166, WX7167, WX7168, WX7169, WX7170,
         WX7171, WX7172, WX7173, WX7174, WX7175, WX7176, WX7177, WX7178,
         WX7179, WX7180, WX7181, WX7182, WX7183, WX7184, WX7185, WX7187,
         WX7188, WX7189, WX7190, WX7191, WX7192, WX7193, WX7194, WX7195,
         WX7196, WX7197, WX7198, WX7199, WX7200, WX7201, WX7202, WX7203,
         WX7204, WX7205, WX7206, WX7207, WX7208, WX7209, WX7210, WX7211,
         WX7212, WX7213, WX7214, WX7215, WX7216, n3647, WX7217, WX7218, WX7219,
         WX7221, WX7222, WX7223, WX7224, n3639, WX7225, WX7226, WX7227, WX7228,
         n3635, WX7229, WX7230, WX7231, WX7232, WX7233, WX7234, WX7235, WX7236,
         WX7237, WX7238, WX7239, WX7240, WX7241, WX7242, WX7243, WX7244,
         WX7245, WX7246, WX7247, WX7248, WX7249, WX7250, WX7251, WX7252,
         WX7253, WX7255, WX7256, WX7257, WX7258, WX7259, WX7260, WX7261,
         WX7262, WX7263, WX7264, WX7265, WX7266, WX7267, WX7268, WX7269,
         WX7270, WX7271, WX7272, WX7273, WX7274, WX7275, WX7276, WX7277,
         WX7278, WX7279, WX7280, WX7281, WX7282, WX7283, WX7284, WX7285,
         WX7286, WX7287, WX7289, WX7290, WX7291, WX7292, WX7293, WX7294,
         WX7295, WX7296, WX7297, WX7298, WX7299, WX7300, WX7301, WX7302,
         WX7303, WX7304, WX7305, WX7306, WX7307, WX7308, WX7309, WX7310,
         WX7311, WX7312, WX7313, WX7314, WX7315, WX7316, WX7317, WX7318,
         WX7319, WX7320, WX7321, WX7323, WX7324, WX7325, WX7326, WX7327,
         WX7328, WX7329, WX7330, WX7331, WX7332, WX7333, WX7334, WX7335,
         WX7336, WX7337, WX7338, WX7339, WX7340, WX7341, WX7342, WX7343,
         WX7344, WX7345, WX7346, WX7347, WX7348, WX7349, WX7350, WX7351,
         WX7352, WX7353, WX7354, WX7355, WX7357, WX7358, WX7359, WX7360,
         WX7361, WX7362, WX7363, WX7364, WX7729, WX7731, WX7733, WX7735,
         WX7737, WX7739, WX7741, WX7743, WX7745, WX7747, WX7749, DFF_1130_n1,
         WX7751, WX7753, WX7755, WX7757, WX7759, DFF_1135_n1, WX7761, WX7763,
         WX7765, WX7767, WX7769, DFF_1140_n1, WX7771, WX7773, WX7775, WX7777,
         WX7779, WX7781, WX7783, WX7785, WX7787, WX7789, WX7791, DFF_1151_n1,
         WX8243, n8411, n3878, n8410, n3877, n8409, n3876, n8408, n3875, n8407,
         n3874, n8406, n3873, n8405, n3872, n8404, n3871, n8403, n3870, n8402,
         n3869, n8401, n3868, WX8266, n8400, n3867, n8399, n3865, n8396, n3864,
         n8395, n3863, n8394, n3862, n8393, n3861, n8392, n3860, n8391, n3859,
         n8390, n3858, n8389, n3857, n8388, n3856, n8387, n3855, n8386, n3854,
         n8385, n3853, n8384, n3852, n8383, n3851, n8382, n3850, n8381, n3849,
         WX8304, n3848, WX8402, n8378, WX8404, n8377, WX8406, n8376, WX8408,
         n8375, WX8410, n8374, WX8412, n8373, WX8414, n8372, WX8416, n8371,
         WX8418, n8370, WX8420, n8369, WX8422, n8368, WX8424, n8367, WX8426,
         n8366, WX8428, n8365, WX8430, n8364, WX8432, n8363, WX8434, WX8436,
         WX8437, WX8438, WX8439, WX8440, WX8441, WX8442, WX8443, WX8444,
         WX8445, WX8446, WX8447, WX8448, WX8449, WX8450, WX8451, WX8452,
         WX8453, WX8454, WX8455, WX8456, WX8457, WX8458, WX8459, WX8460,
         WX8461, WX8462, WX8463, WX8464, WX8465, WX8466, WX8467, WX8468,
         WX8470, WX8471, WX8472, WX8473, WX8474, WX8475, WX8476, WX8477,
         WX8478, WX8479, WX8480, WX8481, WX8482, WX8483, WX8484, WX8485,
         WX8486, WX8487, WX8488, WX8489, WX8490, WX8491, WX8492, WX8493,
         WX8494, WX8495, WX8496, WX8497, WX8498, WX8499, n3625, WX8500, WX8501,
         WX8502, WX8504, WX8505, WX8506, WX8507, n3617, WX8508, WX8509, WX8510,
         WX8511, n3613, WX8512, WX8513, WX8514, WX8515, WX8516, WX8517, WX8518,
         WX8519, WX8520, WX8521, WX8522, WX8523, WX8524, WX8525, WX8526,
         WX8527, WX8528, WX8529, WX8530, WX8531, WX8532, WX8533, WX8534,
         WX8535, WX8536, WX8538, WX8539, WX8540, WX8541, WX8542, WX8543,
         WX8544, WX8545, WX8546, WX8547, WX8548, WX8549, WX8550, WX8551,
         WX8552, WX8553, WX8554, WX8555, WX8556, WX8557, WX8558, WX8559,
         WX8560, WX8561, WX8562, WX8563, WX8564, WX8565, WX8566, WX8567,
         WX8568, WX8569, WX8570, WX8572, WX8573, WX8574, WX8575, WX8576,
         WX8577, WX8578, WX8579, WX8580, WX8581, WX8582, WX8583, WX8584,
         WX8585, WX8586, WX8587, WX8588, WX8589, WX8590, WX8591, WX8592,
         WX8593, WX8594, WX8595, WX8596, WX8597, WX8598, WX8599, WX8600,
         WX8601, WX8602, WX8603, WX8604, WX8606, WX8607, WX8608, WX8609,
         WX8610, WX8611, WX8612, WX8613, WX8614, WX8615, WX8616, WX8617,
         WX8618, WX8619, WX8620, WX8621, WX8622, WX8623, WX8624, WX8625,
         WX8626, WX8627, WX8628, WX8629, WX8630, WX8631, WX8632, WX8633,
         WX8634, WX8635, WX8636, WX8637, WX8638, WX8640, WX8641, WX8642,
         WX8643, WX8644, WX8645, WX8646, WX8647, WX8648, WX8649, WX8650,
         WX8651, WX8652, WX8653, WX8654, WX8655, WX8656, WX8657, WX9022,
         WX9024, WX9026, WX9028, DFF_1315_n1, WX9030, WX9032, WX9034, WX9036,
         WX9038, DFF_1320_n1, WX9040, WX9042, DFF_1322_n1, WX9044, WX9046,
         WX9048, WX9050, WX9052, DFF_1327_n1, WX9054, WX9056, WX9058, WX9060,
         WX9062, WX9064, WX9066, WX9068, WX9070, WX9072, DFF_1337_n1, WX9074,
         WX9076, WX9078, WX9080, WX9082, WX9084, DFF_1343_n1, WX9536, n8353,
         n3847, n8352, n3846, n8351, n3845, n8350, n3844, n8349, n3843, n8348,
         n3842, n8347, n3841, n8346, n3840, n3839, n8343, n3838, n8342, n3837,
         n8341, n3836, n8340, n3835, n8339, n3834, n8338, n3833, n8337, n3832,
         n8336, n3831, n8335, n3830, n8334, n3829, n8333, n3828, n8332, n3827,
         n8331, n3826, n8330, n3825, n8329, n3824, n8328, n3823, n3822, n8325,
         n3821, n8324, n3820, n8323, n3819, n8322, n3818, WX9597, n8321, n3817,
         WX9695, n8320, WX9697, n8319, WX9699, n8318, WX9701, n8317, WX9703,
         n8316, WX9705, n8315, WX9707, n8314, WX9709, n8313, WX9711, n8312,
         WX9713, n8311, WX9715, n8310, WX9717, WX9719, n8307, WX9721, n8306,
         WX9723, n8305, WX9725, n8304, WX9727, WX9728, WX9729, WX9730, WX9731,
         WX9732, WX9733, WX9734, WX9735, WX9736, WX9737, WX9738, WX9739,
         WX9740, WX9741, WX9742, WX9743, WX9744, WX9745, WX9746, WX9747,
         WX9748, WX9749, WX9750, WX9751, WX9753, WX9754, WX9755, WX9756,
         WX9757, WX9758, WX9759, WX9760, WX9761, WX9762, WX9763, WX9764,
         WX9765, WX9766, WX9767, WX9768, WX9769, WX9770, WX9771, WX9772,
         WX9773, WX9774, WX9775, WX9776, WX9777, WX9778, WX9779, WX9780,
         WX9781, WX9782, WX9783, WX9784, WX9785, WX9787, WX9788, WX9789,
         WX9790, WX9791, WX9792, WX9793, WX9794, n3591, WX9795, WX9796, WX9797,
         WX9798, WX9799, WX9800, WX9801, WX9802, WX9803, WX9804, WX9805,
         WX9806, WX9807, WX9808, WX9809, WX9810, WX9811, WX9812, WX9813,
         WX9814, WX9815, WX9816, n3569, WX9817, WX9818, WX9819, WX9821, WX9822,
         WX9823, WX9824, WX9825, WX9826, WX9827, WX9828, WX9829, WX9830,
         WX9831, WX9832, WX9833, WX9834, WX9835, WX9836, WX9837, WX9838,
         WX9839, WX9840, WX9841, WX9842, WX9843, WX9844, WX9845, WX9846,
         WX9847, WX9848, WX9849, WX9850, WX9851, WX9852, WX9853, WX9855,
         WX9856, WX9857, WX9858, WX9859, WX9860, WX9861, WX9862, WX9863,
         WX9864, WX9865, WX9866, WX9867, WX9868, WX9869, WX9870, WX9871,
         WX9872, WX9873, WX9874, WX9875, WX9876, WX9877, WX9878, WX9879,
         WX9880, WX9881, WX9882, WX9883, WX9884, WX9885, WX9886, WX9887,
         WX9889, WX9890, WX9891, WX9892, WX9893, WX9894, WX9895, WX9896,
         WX9897, WX9898, WX9899, WX9900, WX9901, WX9902, WX9903, WX9904,
         WX9905, WX9906, WX9907, WX9908, WX9909, WX9910, WX9911, WX9912,
         WX9913, WX9914, WX9915, WX9916, WX9917, WX9918, WX9919, WX9920,
         WX9921, WX9923, WX9924, WX9925, WX9926, WX9927, WX9928, WX9929,
         WX9930, WX9931, WX9932, WX9933, WX9934, WX9935, WX9936, WX9937,
         WX9938, WX9939, WX9940, WX9941, WX9942, WX9943, WX9944, WX9945,
         WX9946, WX9947, WX9948, WX9949, WX9950, WX10315, WX10317, WX10319,
         WX10321, DFF_1507_n1, WX10323, WX10325, WX10327, WX10329, WX10331,
         WX10333, WX10335, DFF_1514_n1, WX10337, WX10339, WX10341, DFF_1517_n1,
         WX10343, WX10345, DFF_1519_n1, WX10347, WX10349, WX10351, WX10353,
         WX10355, WX10357, WX10359, WX10361, WX10363, WX10365, WX10367,
         WX10369, WX10371, WX10373, WX10375, DFF_1534_n1, WX10377, DFF_1535_n1,
         WX10829, n8295, n3816, n8294, n3815, n8293, n3814, n3813, n8290,
         n3812, n8289, n3811, n8288, n3810, n8287, n3809, n8286, n3808, n8285,
         n3807, n8284, n3806, n8283, n3805, n8282, n3804, n8281, n3803, n8280,
         n3802, n8279, n3801, n8278, n3800, n8277, n3799, n8276, n3798, n8275,
         n3797, n3796, n8272, n3795, n8271, n3794, n8270, n3793, n8269, n3792,
         n8268, n3791, n8267, n3790, n8266, n3789, n8265, n3788, n8264, n3787,
         WX10890, n8263, n3786, WX10988, n8262, WX10990, n8261, WX10992, n8260,
         WX10994, n8259, WX10996, n8258, WX10998, n8257, WX11000, WX11002,
         n8254, WX11004, n8253, WX11006, n8252, WX11008, n8251, WX11010, n8250,
         WX11012, n8249, WX11014, n8248, WX11016, n8247, WX11018, n8246,
         WX11020, WX11021, WX11022, WX11023, WX11024, WX11025, WX11026,
         WX11027, WX11028, WX11029, WX11030, WX11031, WX11032, WX11033,
         WX11034, WX11036, WX11037, WX11038, WX11039, WX11040, WX11041,
         WX11042, WX11043, WX11044, WX11045, WX11046, WX11047, WX11048,
         WX11049, WX11050, WX11051, WX11052, WX11053, WX11054, WX11055,
         WX11056, WX11057, WX11058, WX11059, WX11060, WX11061, WX11062,
         WX11063, WX11064, WX11065, WX11066, WX11067, WX11068, WX11070,
         WX11071, WX11072, WX11073, WX11074, WX11075, WX11076, WX11077,
         WX11078, WX11079, WX11080, WX11081, WX11082, WX11083, WX11084,
         WX11085, WX11086, WX11087, WX11088, WX11089, WX11090, WX11091,
         WX11092, WX11093, WX11094, WX11095, WX11096, WX11097, WX11098,
         WX11099, n3547, WX11100, WX11101, WX11102, WX11104, WX11105, WX11106,
         WX11107, n3539, WX11108, WX11109, WX11110, WX11111, n3535, WX11112,
         WX11113, WX11114, WX11115, WX11116, WX11117, WX11118, WX11119,
         WX11120, WX11121, WX11122, WX11123, WX11124, WX11125, WX11126,
         WX11127, WX11128, WX11129, WX11130, WX11131, WX11132, WX11133,
         WX11134, WX11135, WX11136, WX11138, WX11139, WX11140, WX11141,
         WX11142, WX11143, WX11144, WX11145, WX11146, WX11147, WX11148,
         WX11149, WX11150, WX11151, WX11152, WX11153, WX11154, WX11155,
         WX11156, WX11157, WX11158, WX11159, WX11160, WX11161, WX11162,
         WX11163, WX11164, WX11165, WX11166, WX11167, WX11168, WX11169,
         WX11170, WX11172, WX11173, WX11174, WX11175, WX11176, WX11177,
         WX11178, WX11179, WX11180, WX11181, WX11182, WX11183, WX11184,
         WX11185, WX11186, WX11187, WX11188, WX11189, WX11190, WX11191,
         WX11192, WX11193, WX11194, WX11195, WX11196, WX11197, WX11198,
         WX11199, WX11200, WX11201, WX11202, WX11203, WX11204, WX11206,
         WX11207, WX11208, WX11209, WX11210, WX11211, WX11212, WX11213,
         WX11214, WX11215, WX11216, WX11217, WX11218, WX11219, WX11220,
         WX11221, WX11222, WX11223, WX11224, WX11225, WX11226, WX11227,
         WX11228, WX11229, WX11230, WX11231, WX11232, WX11233, WX11234,
         WX11235, WX11236, WX11237, WX11238, WX11240, WX11241, WX11242,
         WX11243, WX11608, WX11610, DFF_1697_n1, WX11612, WX11614, WX11616,
         WX11618, WX11620, WX11622, WX11624, WX11626, WX11628, WX11630,
         WX11632, WX11634, WX11636, WX11638, WX11640, WX11642, WX11644,
         DFF_1714_n1, WX11646, WX11648, WX11650, WX11652, WX11654, WX11656,
         WX11658, WX11660, WX11662, WX11664, WX11666, WX11668, WX11670, n2245,
         n2153, n3278, n2152, n2148, Tj_Trigger, Tj_OUT1, Tj_OUT2, Tj_OUT3,
         Tj_OUT4, Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         test_se_NOT, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n308, n309, n310, n311, n312, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n530,
         n2832, n2834, n2835, n2837, n2839, n2841, n2843, n2845, n2847, n2849,
         n2851, n2853, n2854, n2856, n2857, n2859, n2860, n2862, n2863, n2865,
         n2867, n2869, n2871, n2873, n2874, n2876, n2877, n2879, n2880, n2882,
         n2884, n2886, n2888, n2890, n2892, n2894, n2896, n2898, n2900, n2902,
         n2904, n2906, n2908, n2910, n2912, n2914, n2916, n2918, n2920, n2921,
         n2923, n2924, n2926, n2927, n2929, n2931, n2933, n2935, n2937, n2938,
         n2940, n2941, n2943, n2944, n2946, n2947, n2949, n2951, n2953, n2954,
         n2956, n2957, n2959, n2960, n2962, n2963, n2965, n2967, n2969, n2971,
         n2973, n2975, n2977, n2979, n2981, n2982, n2984, n2986, n2988, n2990,
         n2992, n2994, n2996, n2998, n3000, n3002, n3003, n3005, n3006, n3007,
         n3009, n3011, n3013, n3015, n3017, n3019, n3020, n3022, n3024, n3025,
         n3027, n3029, n3031, n3032, n3034, n3036, n3037, n3039, n3041, n3043,
         n3044, n3046, n3048, n3050, n3052, n3054, n3055, n3057, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3417, n3418, n3420, n3422, n3424, n3426,
         n3428, n3429, n3431, n3433, n3435, n3436, n3438, n3440, n3442, n3443,
         n3444, n3445, n3447, n3448, n3450, n3452, n3454, n3456, n3457, n3459,
         n3460, n3462, n3463, n3464, n3465, n3466, n3468, n3470, n3476, n3478,
         n3482, n3484, n3488, n3490, n3496, n3498, n3500, n3502, n3504, n3506,
         n3508, n3510, n3512, n3514, n3515, n3516, n3518, n3520, n3522, n3523,
         n3524, n3526, n3528, n3530, n3531, n3532, n3533, n3534, n3536, n3537,
         n3538, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3614, n3615, n3616, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3636, n3637, n3638, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3714, n3715, n3716, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3736, n3737, n3738, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3784, n3785, n3866, n3884,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, U3558_n1, U3871_n1, U3991_n1,
         U5716_n1, U5717_n1, U5718_n1, U5719_n1, U5720_n1, U5721_n1, U5722_n1,
         U5723_n1, U5724_n1, U5725_n1, U5726_n1, U5727_n1, U5728_n1, U5729_n1,
         U5730_n1, U5731_n1, U5732_n1, U5733_n1, U5734_n1, U5735_n1, U5736_n1,
         U5737_n1, U5738_n1, U5739_n1, U5740_n1, U5741_n1, U5742_n1, U5743_n1,
         U5744_n1, U5745_n1, U5746_n1, U5747_n1, U5748_n1, U5749_n1, U5750_n1,
         U5751_n1, U5752_n1, U5753_n1, U5754_n1, U5755_n1, U5756_n1, U5757_n1,
         U5758_n1, U5759_n1, U5760_n1, U5761_n1, U5762_n1, U5763_n1, U5764_n1,
         U5765_n1, U5766_n1, U5767_n1, U5768_n1, U5769_n1, U5770_n1, U5771_n1,
         U5772_n1, U5773_n1, U5774_n1, U5775_n1, U5776_n1, U5777_n1, U5778_n1,
         U5779_n1, U5780_n1, U5781_n1, U5782_n1, U5783_n1, U5784_n1, U5785_n1,
         U5786_n1, U5787_n1, U5788_n1, U5789_n1, U5790_n1, U5791_n1, U5792_n1,
         U5793_n1, U5794_n1, U5795_n1, U5796_n1, U5797_n1, U5798_n1, U5799_n1,
         U5800_n1, U5801_n1, U5802_n1, U5803_n1, U5804_n1, U5805_n1, U5806_n1,
         U5807_n1, U5808_n1, U5809_n1, U5810_n1, U5811_n1, U5812_n1, U5813_n1,
         U5814_n1, U5815_n1, U5816_n1, U5817_n1, U5818_n1, U5819_n1, U5820_n1,
         U5821_n1, U5822_n1, U5823_n1, U5824_n1, U5825_n1, U5826_n1, U5827_n1,
         U5828_n1, U5829_n1, U5830_n1, U5831_n1, U5832_n1, U5833_n1, U5834_n1,
         U5835_n1, U5836_n1, U5837_n1, U5838_n1, U5839_n1, U5840_n1, U5841_n1,
         U5842_n1, U5843_n1, U5844_n1, U5845_n1, U5846_n1, U5847_n1, U5848_n1,
         U5849_n1, U5850_n1, U5851_n1, U5852_n1, U5853_n1, U5854_n1, U5855_n1,
         U5856_n1, U5857_n1, U5858_n1, U5859_n1, U5860_n1, U5861_n1, U5862_n1,
         U5863_n1, U5864_n1, U5865_n1, U5866_n1, U5867_n1, U5868_n1, U5869_n1,
         U5870_n1, U5871_n1, U5872_n1, U5873_n1, U5874_n1, U5875_n1, U5876_n1,
         U5877_n1, U5878_n1, U5879_n1, U5880_n1, U5881_n1, U5882_n1, U5883_n1,
         U5884_n1, U5885_n1, U5886_n1, U5887_n1, U5888_n1, U5889_n1, U5890_n1,
         U5891_n1, U5892_n1, U5893_n1, U5894_n1, U5895_n1, U5896_n1, U5897_n1,
         U5898_n1, U5899_n1, U5900_n1, U5901_n1, U5902_n1, U5903_n1, U5904_n1,
         U5905_n1, U5906_n1, U5907_n1, U5908_n1, U5909_n1, U5910_n1, U5911_n1,
         U5912_n1, U5913_n1, U5914_n1, U5915_n1, U5916_n1, U5917_n1, U5918_n1,
         U5919_n1, U5920_n1, U5921_n1, U5922_n1, U5923_n1, U5924_n1, U5925_n1,
         U5926_n1, U5927_n1, U5928_n1, U5929_n1, U5930_n1, U5931_n1, U5932_n1,
         U5933_n1, U5934_n1, U5935_n1, U5936_n1, U5937_n1, U5938_n1, U5939_n1,
         U5940_n1, U5941_n1, U5942_n1, U5943_n1, U5944_n1, U5945_n1, U5946_n1,
         U5947_n1, U5948_n1, U5949_n1, U5950_n1, U5951_n1, U5952_n1, U5953_n1,
         U5954_n1, U5955_n1, U5956_n1, U5957_n1, U5958_n1, U5959_n1, U5960_n1,
         U5961_n1, U5962_n1, U5963_n1, U5964_n1, U5965_n1, U5966_n1, U5967_n1,
         U5968_n1, U5969_n1, U5970_n1, U5971_n1, U5972_n1, U5973_n1, U5974_n1,
         U5975_n1, U5976_n1, U5977_n1, U5978_n1, U5979_n1, U5980_n1, U5981_n1,
         U5982_n1, U5983_n1, U5984_n1, U5985_n1, U5986_n1, U5987_n1, U5988_n1,
         U5989_n1, U5990_n1, U5991_n1, U5992_n1, U5993_n1, U5994_n1, U5995_n1,
         U5996_n1, U5997_n1, U5998_n1, U5999_n1, U6000_n1, U6001_n1, U6002_n1,
         U6003_n1, U6004_n1, U6005_n1, U6006_n1, U6007_n1, U6008_n1, U6009_n1,
         U6010_n1, U6011_n1, U6012_n1, U6013_n1, U6014_n1, U6015_n1, U6016_n1,
         U6017_n1, U6018_n1, U6019_n1, U6020_n1, U6021_n1, U6022_n1, U6023_n1,
         U6024_n1, U6025_n1, U6026_n1, U6027_n1, U6028_n1, U6029_n1, U6030_n1,
         U6031_n1, U6032_n1, U6033_n1, U6034_n1, U6035_n1, U6036_n1, U6037_n1,
         U6038_n1, U6039_n1, U6040_n1, U6041_n1, U6042_n1, U6043_n1, U6044_n1,
         U6045_n1, U6046_n1, U6047_n1, U6048_n1, U6049_n1, U6050_n1, U6051_n1,
         U6052_n1, U6053_n1, U6054_n1, U6055_n1, U6056_n1, U6057_n1, U6058_n1,
         U6059_n1, U6060_n1, U6061_n1, U6062_n1, U6063_n1, U6064_n1, U6065_n1,
         U6066_n1, U6067_n1, U6068_n1, U6069_n1, U6070_n1, U6071_n1, U6072_n1,
         U6073_n1, U6074_n1, U6075_n1, U6076_n1, U6077_n1, U6078_n1, U6079_n1,
         U6080_n1, U6081_n1, U6082_n1, U6083_n1, U6084_n1, U6085_n1, U6086_n1,
         U6087_n1, U6088_n1, U6089_n1, U6090_n1, U6091_n1, U6092_n1, U6093_n1,
         U6094_n1, U6095_n1, U6096_n1, U6097_n1, U6098_n1, U6099_n1, U6100_n1,
         U6101_n1, U6102_n1, U6103_n1, U6104_n1, U6105_n1, U6106_n1, U6107_n1,
         U6108_n1, U6109_n1, U6110_n1, U6111_n1, U6112_n1, U6113_n1, U6114_n1,
         U6115_n1, U6116_n1, U6117_n1, U6118_n1, U6119_n1, U6120_n1, U6121_n1,
         U6122_n1, U6123_n1, U6124_n1, U6125_n1, U6126_n1, U6127_n1, U6128_n1,
         U6129_n1, U6130_n1, U6131_n1, U6132_n1, U6133_n1, U6134_n1, U6135_n1,
         U6136_n1, U6137_n1, U6138_n1, U6139_n1, U6140_n1, U6141_n1, U6142_n1,
         U6143_n1, U6144_n1, U6145_n1, U6146_n1, U6147_n1, U6148_n1, U6149_n1,
         U6150_n1, U6151_n1, U6152_n1, U6153_n1, U6154_n1, U6155_n1, U6156_n1,
         U6157_n1, U6158_n1, U6159_n1, U6160_n1, U6161_n1, U6162_n1, U6163_n1,
         U6164_n1, U6165_n1, U6166_n1, U6167_n1, U6168_n1, U6169_n1, U6170_n1,
         U6171_n1, U6172_n1, U6173_n1, U6174_n1, U6175_n1, U6176_n1, U6177_n1,
         U6178_n1, U6179_n1, U6180_n1, U6181_n1, U6182_n1, U6183_n1, U6184_n1,
         U6185_n1, U6186_n1, U6187_n1, U6188_n1, U6189_n1, U6190_n1, U6191_n1,
         U6192_n1, U6193_n1, U6194_n1, U6195_n1, U6196_n1, U6197_n1, U6198_n1,
         U6199_n1, U6200_n1, U6201_n1, U6202_n1, U6203_n1, U6204_n1, U6205_n1,
         U6206_n1, U6207_n1, U6208_n1, U6209_n1, U6210_n1, U6211_n1, U6212_n1,
         U6213_n1, U6214_n1, U6215_n1, U6216_n1, U6217_n1, U6218_n1, U6219_n1,
         U6220_n1, U6221_n1, U6222_n1, U6223_n1, U6224_n1, U6225_n1, U6226_n1,
         U6227_n1, U6228_n1, U6229_n1, U6230_n1, U6231_n1, U6232_n1, U6233_n1,
         U6234_n1, U6235_n1, U6236_n1, U6237_n1, U6238_n1, U6239_n1, U6240_n1,
         U6241_n1, U6242_n1, U6243_n1, U6244_n1, U6245_n1, U6246_n1, U6247_n1,
         U6248_n1, U6249_n1, U6250_n1, U6251_n1, U6252_n1, U6253_n1, U6254_n1,
         U6255_n1, U6256_n1, U6257_n1, U6258_n1, U6259_n1, U6260_n1, U6261_n1,
         U6262_n1, U6263_n1, U6264_n1, U6265_n1, U6266_n1, U6267_n1, U6268_n1,
         U6269_n1, U6270_n1, U6271_n1, U6272_n1, U6273_n1, U6274_n1, U6275_n1,
         U6276_n1, U6277_n1, U6278_n1, U6279_n1, U6280_n1, U6281_n1, U6282_n1,
         U6283_n1, U6284_n1, U6285_n1, U6286_n1, U6287_n1, U6288_n1, U6289_n1,
         U6290_n1, U6291_n1, U6292_n1, U6293_n1, U6294_n1, U6295_n1, U6296_n1,
         U6297_n1, U6298_n1, U6299_n1, U6300_n1, U6301_n1, U6302_n1, U6303_n1,
         U6304_n1, U6305_n1, U6306_n1, U6307_n1, U6308_n1, U6309_n1, U6310_n1,
         U6311_n1, U6312_n1, U6313_n1, U6314_n1, U6315_n1, U6316_n1, U6317_n1,
         U6318_n1, U6319_n1, U6320_n1, U6321_n1, U6322_n1, U6323_n1, U6324_n1,
         U6325_n1, U6326_n1, U6327_n1, U6328_n1, U6329_n1, U6330_n1, U6331_n1,
         U6332_n1, U6333_n1, U6334_n1, U6335_n1, U6336_n1, U6337_n1, U6338_n1,
         U6339_n1, U6340_n1, U6341_n1, U6342_n1, U6343_n1, U6344_n1, U6345_n1,
         U6346_n1, U6347_n1, U6348_n1, U6349_n1, U6350_n1, U6351_n1, U6352_n1,
         U6353_n1, U6354_n1, U6355_n1, U6356_n1, U6357_n1, U6358_n1, U6359_n1,
         U6360_n1, U6361_n1, U6362_n1, U6363_n1, U6364_n1, U6365_n1, U6366_n1,
         U6367_n1, U6368_n1, U6369_n1, U6370_n1, U6371_n1, U6372_n1, U6373_n1,
         U6374_n1, U6375_n1, U6376_n1, U6377_n1, U6378_n1, U6379_n1, U6380_n1,
         U6381_n1, U6382_n1, U6383_n1, U6384_n1, U6385_n1, U6386_n1, U6387_n1,
         U6388_n1, U6389_n1, U6390_n1, U6391_n1, U6392_n1, U6393_n1, U6394_n1,
         U6395_n1, U6396_n1, U6397_n1, U6398_n1, U6399_n1, U6400_n1, U6401_n1,
         U6402_n1, U6403_n1, U6404_n1, U6405_n1, U6406_n1, U6407_n1, U6408_n1,
         U6409_n1, U6410_n1, U6411_n1, U6412_n1, U6413_n1, U6414_n1, U6415_n1,
         U6416_n1, U6417_n1, U6418_n1, U6419_n1, U6420_n1, U6421_n1, U6422_n1,
         U6423_n1, U6424_n1, U6425_n1, U6426_n1, U6427_n1, U6428_n1, U6429_n1,
         U6430_n1, U6431_n1, U6432_n1, U6433_n1, U6434_n1, U6435_n1, U6436_n1,
         U6437_n1, U6438_n1, U6439_n1, U6440_n1, U6441_n1, U6442_n1, U6443_n1,
         U6444_n1, U6445_n1, U6446_n1, U6447_n1, U6448_n1, U6449_n1, U6450_n1,
         U6451_n1, U6452_n1, U6453_n1, U6454_n1, U6455_n1, U6456_n1, U6457_n1,
         U6458_n1, U6459_n1, U6460_n1, U6461_n1, U6462_n1, U6463_n1, U6464_n1,
         U6465_n1, U6466_n1, U6467_n1, U6468_n1, U6469_n1, U6470_n1, U6471_n1,
         U6472_n1, U6473_n1, U6474_n1, U6475_n1, U6476_n1, U6477_n1, U6478_n1,
         U6479_n1, U6480_n1, U6481_n1, U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n4195), .CLK(n4491), .Q(
        WX485), .QN(n3512) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n4190), .CLK(n4493), .Q(
        WX487) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n4190), .CLK(n4493), .Q(
        WX489) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n4191), .CLK(n4493), .Q(
        WX491) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n4191), .CLK(n4493), .Q(
        WX493) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n4191), .CLK(n4493), .Q(
        WX495) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n4191), .CLK(n4493), .Q(
        WX497) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n4191), .CLK(n4493), .Q(
        WX499) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n4191), .CLK(n4493), .Q(
        WX501) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n4192), .CLK(n4492), .Q(
        WX503) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n4192), .CLK(n4492), .Q(
        WX505) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n4192), .CLK(n4492), .Q(
        WX507) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n4192), .CLK(n4492), .Q(
        WX509) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n4192), .CLK(n4492), .Q(
        WX511) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(n4192), .CLK(n4492), .Q(
        WX513) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n4193), .CLK(n4492), .Q(
        WX515) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n4193), .CLK(n4492), .Q(
        WX517) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n4193), .CLK(n4492), .Q(
        test_so1) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n4193), .CLK(n4492), .Q(
        WX521) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n4193), .CLK(n4492), .Q(
        WX523) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n4193), .CLK(n4492), .Q(
        WX525) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(n4194), .CLK(n4491), .Q(
        WX527) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n4194), .CLK(n4491), .Q(
        WX529) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n4194), .CLK(n4491), .Q(
        WX531) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n4194), .CLK(n4491), .Q(
        WX533) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n4194), .CLK(n4491), .Q(
        WX535) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n4194), .CLK(n4491), .Q(
        WX537) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n4195), .CLK(n4491), .Q(
        WX539) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n4195), .CLK(n4491), .Q(
        WX541) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n4195), .CLK(n4491), .Q(
        WX543) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n4195), .CLK(n4491), .Q(
        WX545) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n4195), .CLK(n4491), .Q(
        WX547) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n4190), .CLK(n4493), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(n4190), .CLK(n4493), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(n4190), .CLK(n4493), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(n4190), .CLK(n4493), .Q(
        test_so2) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(n3652), .CLK(n4634), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(n3652), .CLK(n4634), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(n3652), .CLK(n4634), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n4189), .CLK(n4494), .Q(
        WX659) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(n4188), .CLK(n4494), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(n4188), .CLK(n4494), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(n4188), .CLK(n4494), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n4187), .CLK(n4495), .Q(
        WX667) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(n4187), .CLK(n4495), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(n4187), .CLK(n4495), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(n4186), .CLK(n4495), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n4186), .CLK(n4495), .Q(
        WX675) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(n4185), .CLK(n4496), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(n4184), .CLK(n4496), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(n4184), .CLK(n4496), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(n4183), .CLK(n4497), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(n4182), .CLK(n4497), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n4182), .CLK(n4497), .Q(
        test_so3) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(n4181), .CLK(n4498), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(n4180), .CLK(n4498), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(n4180), .CLK(n4498), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(n4179), .CLK(n4499), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(n4178), .CLK(n4499), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(n4178), .CLK(n4499), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(n4177), .CLK(n4500), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(n4176), .CLK(n4500), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(n4176), .CLK(n4500), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(n4175), .CLK(n4501), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n4174), .CLK(n4501), .Q(
        WX709), .QN(n7269) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n4174), .CLK(n4501), .Q(
        WX711), .QN(n3415) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n4173), .CLK(n4502), .Q(
        WX713) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n4189), .CLK(n4494), .Q(
        WX715), .QN(n7272) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n4189), .CLK(n4494), .Q(
        WX717) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n4189), .CLK(n4494), .Q(
        WX719) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n4189), .CLK(n4494), .Q(
        WX721) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n4189), .CLK(n4494), .Q(
        test_so4) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n4188), .CLK(n4494), .Q(
        WX725) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n4188), .CLK(n4494), .Q(
        WX727), .QN(n3454) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n4188), .CLK(n4494), .Q(
        WX729), .QN(n3460) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n4187), .CLK(n4495), .Q(
        WX731), .QN(n7278) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n4187), .CLK(n4495), .Q(
        WX733) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n4186), .CLK(n4495), .Q(
        WX735) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n4186), .CLK(n4495), .Q(
        WX737) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n4185), .CLK(n4496), .Q(
        WX739), .QN(n3447) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n4185), .CLK(n4496), .Q(
        WX741), .QN(n3457) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n4184), .CLK(n4496), .Q(
        WX743) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n4184), .CLK(n4496), .Q(
        WX745) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n4183), .CLK(n4497), .Q(
        WX747) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n4182), .CLK(n4497), .Q(
        WX749) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n4182), .CLK(n4497), .Q(
        WX751), .QN(n7287) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n4181), .CLK(n4498), .Q(
        WX753), .QN(n7265) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n4180), .CLK(n4498), .Q(
        WX755) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n4180), .CLK(n4498), .Q(
        WX757), .QN(n3478) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n4179), .CLK(n4499), .Q(
        test_so5) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n4178), .CLK(n4499), .Q(
        WX761) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n4178), .CLK(n4499), .Q(
        WX763) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n4177), .CLK(n4500), .Q(
        WX765) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n4176), .CLK(n4500), .Q(
        WX767) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n4176), .CLK(n4500), .Q(
        WX769) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n4175), .CLK(n4501), .Q(
        WX771) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n4174), .CLK(n4501), .Q(
        WX773), .QN(n3466) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n4174), .CLK(n4501), .Q(
        WX775) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n4173), .CLK(n4502), .Q(
        WX777), .QN(n7271) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n4173), .CLK(n4502), .Q(
        WX779) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n4173), .CLK(n4502), .Q(
        WX781), .QN(n7273) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n4172), .CLK(n4502), .Q(
        WX783), .QN(n7274) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n4172), .CLK(n4502), .Q(
        WX785), .QN(n7275) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n4172), .CLK(n4502), .Q(
        WX787), .QN(n7276) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n4171), .CLK(n4503), .Q(
        WX789), .QN(n7277) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n4171), .CLK(n4503), .Q(
        WX791) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n4171), .CLK(n4503), .Q(
        WX793) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n4170), .CLK(n4503), .Q(
        test_so6) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n4187), .CLK(n4495), 
        .Q(WX797), .QN(n7279) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n4186), .CLK(n4495), .Q(
        WX799), .QN(n7280) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n4186), .CLK(n4495), .Q(
        WX801), .QN(n7281) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n4185), .CLK(n4496), .Q(
        WX803), .QN(n7282) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n4185), .CLK(n4496), .Q(
        WX805) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n4184), .CLK(n4496), .Q(
        WX807), .QN(n7283) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n4183), .CLK(n4497), .Q(
        WX809), .QN(n7284) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n4183), .CLK(n4497), .Q(
        WX811), .QN(n7285) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n4182), .CLK(n4497), .Q(
        WX813), .QN(n7286) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n4181), .CLK(n4498), .Q(
        WX815) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n4181), .CLK(n4498), .Q(
        WX817), .QN(n3442) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n4180), .CLK(n4498), .Q(
        WX819), .QN(n7266) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n4179), .CLK(n4499), .Q(
        WX821) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n4179), .CLK(n4499), .Q(
        WX823), .QN(n3463) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n4178), .CLK(n4499), .Q(
        WX825), .QN(n7267) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n4177), .CLK(n4500), .Q(
        WX827), .QN(n7268) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n4177), .CLK(n4500), .Q(
        WX829), .QN(n7270) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n4176), .CLK(n4500), .Q(
        test_so7) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n4175), .CLK(n4501), 
        .Q(WX833), .QN(n7288) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n4175), .CLK(n4501), .Q(
        WX835), .QN(n3488) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n4174), .CLK(n4501), .Q(
        WX837), .QN(n3468) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n4174), .CLK(n4501), .Q(
        WX839), .QN(n3417) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n4173), .CLK(n4502), .Q(
        WX841), .QN(n3422) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n4173), .CLK(n4502), .Q(
        WX843), .QN(n3428) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n4172), .CLK(n4502), .Q(
        WX845), .QN(n3431) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n4172), .CLK(n4502), .Q(
        WX847), .QN(n3433) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n4172), .CLK(n4502), .Q(
        WX849), .QN(n3438) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n4171), .CLK(n4503), .Q(
        WX851), .QN(n3444) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n4171), .CLK(n4503), .Q(
        WX853), .QN(n3445) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n4171), .CLK(n4503), .Q(
        WX855), .QN(n3456) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n4170), .CLK(n4503), .Q(
        WX857), .QN(n3462) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n4170), .CLK(n4503), .Q(
        WX859), .QN(n3465) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n4170), .CLK(n4503), .Q(
        WX861), .QN(n3420) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n4170), .CLK(n4503), .Q(
        WX863), .QN(n3429) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n4170), .CLK(n4503), .Q(
        WX865), .QN(n3436) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n4169), .CLK(n4504), .Q(
        test_so8) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n4185), .CLK(n4496), 
        .Q(WX869), .QN(n3459) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n4184), .CLK(n4496), .Q(
        WX871), .QN(n3470) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n4183), .CLK(n4497), .Q(
        WX873), .QN(n3424) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n4183), .CLK(n4497), .Q(
        WX875), .QN(n3440) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n4182), .CLK(n4497), .Q(
        WX877), .QN(n3484) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n4181), .CLK(n4498), .Q(
        WX879), .QN(n3435) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n4181), .CLK(n4498), .Q(
        WX881), .QN(n3443) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n4180), .CLK(n4498), .Q(
        WX883), .QN(n3448) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n4179), .CLK(n4499), .Q(
        WX885), .QN(n3482) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n4179), .CLK(n4499), .Q(
        WX887), .QN(n3464) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n4178), .CLK(n4499), .Q(
        WX889), .QN(n3450) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n4177), .CLK(n4500), .Q(
        WX891), .QN(n3452) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n4177), .CLK(n4500), .Q(
        WX893), .QN(n3418) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n4176), .CLK(n4500), .Q(
        WX895), .QN(n3476) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n4175), .CLK(n4501), .Q(
        WX897), .QN(n3426) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n4175), .CLK(n4501), .Q(
        WX899), .QN(n3490) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n3655), .CLK(n4633), .Q(
        CRC_OUT_9_0) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n3655), .CLK(n4633), 
        .Q(test_so9) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n3655), .CLK(n4633), 
        .Q(CRC_OUT_9_2) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n3655), .CLK(n4633), 
        .Q(CRC_OUT_9_3), .QN(DFF_163_n1) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n3655), .CLK(n4633), 
        .Q(CRC_OUT_9_4) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n3654), .CLK(n4633), 
        .Q(CRC_OUT_9_5) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n3654), .CLK(n4633), 
        .Q(CRC_OUT_9_6) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n3654), .CLK(n4633), 
        .Q(CRC_OUT_9_7) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n3654), .CLK(n4633), 
        .Q(CRC_OUT_9_8) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n3654), .CLK(n4633), 
        .Q(CRC_OUT_9_9) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n3654), .CLK(n4633), 
        .Q(CRC_OUT_9_10), .QN(DFF_170_n1) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n3653), .CLK(n4634), .Q(CRC_OUT_9_11) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n3653), .CLK(n4634), .Q(CRC_OUT_9_12) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n3653), .CLK(n4634), .Q(CRC_OUT_9_13) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n3653), .CLK(n4634), .Q(CRC_OUT_9_14) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n3653), .CLK(n4634), .Q(CRC_OUT_9_15) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n3653), .CLK(n4634), .Q(CRC_OUT_9_16) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n3652), .CLK(n4634), .Q(CRC_OUT_9_17) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n3652), .CLK(n4634), .Q(CRC_OUT_9_18) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n3652), .CLK(n4634), .Q(test_so10) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n4169), .CLK(n4504), 
        .Q(CRC_OUT_9_20) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n4169), .CLK(n4504), .Q(CRC_OUT_9_21) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n4169), .CLK(n4504), .Q(CRC_OUT_9_22) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n4169), .CLK(n4504), .Q(CRC_OUT_9_23) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n4169), .CLK(n4504), .Q(CRC_OUT_9_24) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n4168), .CLK(n4504), .Q(CRC_OUT_9_25) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n4168), .CLK(n4504), .Q(CRC_OUT_9_26) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n4168), .CLK(n4504), .Q(CRC_OUT_9_27) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n4168), .CLK(n4504), .Q(CRC_OUT_9_28) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n4168), .CLK(n4504), .Q(CRC_OUT_9_29) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(n4168), .CLK(n4504), .Q(CRC_OUT_9_30) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n4167), .CLK(n4505), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n33), .SI(CRC_OUT_9_31), .SE(n4167), .CLK(n4505), 
        .Q(WX1778), .QN(n3496) );
  SDFFX1 DFF_193_Q_reg ( .D(n34), .SI(WX1778), .SE(n4162), .CLK(n4507), .Q(
        n8702), .QN(n4033) );
  SDFFX1 DFF_194_Q_reg ( .D(n35), .SI(n8702), .SE(n4162), .CLK(n4507), .Q(
        n8701), .QN(n4032) );
  SDFFX1 DFF_195_Q_reg ( .D(n36), .SI(n8701), .SE(n4162), .CLK(n4507), .Q(
        n8700), .QN(n4031) );
  SDFFX1 DFF_196_Q_reg ( .D(n37), .SI(n8700), .SE(n4163), .CLK(n4507), .Q(
        n8699), .QN(n4030) );
  SDFFX1 DFF_197_Q_reg ( .D(n38), .SI(n8699), .SE(n4163), .CLK(n4507), .Q(
        test_so11), .QN(n4029) );
  SDFFX1 DFF_198_Q_reg ( .D(n39), .SI(test_si12), .SE(n4163), .CLK(n4507), .Q(
        n8696), .QN(n4028) );
  SDFFX1 DFF_199_Q_reg ( .D(n40), .SI(n8696), .SE(n4163), .CLK(n4507), .Q(
        n8695), .QN(n4027) );
  SDFFX1 DFF_200_Q_reg ( .D(n41), .SI(n8695), .SE(n4163), .CLK(n4507), .Q(
        n8694), .QN(n4026) );
  SDFFX1 DFF_201_Q_reg ( .D(n42), .SI(n8694), .SE(n4163), .CLK(n4507), .Q(
        n8693), .QN(n4025) );
  SDFFX1 DFF_202_Q_reg ( .D(n43), .SI(n8693), .SE(n4164), .CLK(n4506), .Q(
        n8692), .QN(n4024) );
  SDFFX1 DFF_203_Q_reg ( .D(n44), .SI(n8692), .SE(n4164), .CLK(n4506), .Q(
        n8691), .QN(n4023) );
  SDFFX1 DFF_204_Q_reg ( .D(n45), .SI(n8691), .SE(n4164), .CLK(n4506), .Q(
        n8690), .QN(n4022) );
  SDFFX1 DFF_205_Q_reg ( .D(n46), .SI(n8690), .SE(n4164), .CLK(n4506), .Q(
        n8689), .QN(n4021) );
  SDFFX1 DFF_206_Q_reg ( .D(n47), .SI(n8689), .SE(n4164), .CLK(n4506), .Q(
        n8688), .QN(n4020) );
  SDFFX1 DFF_207_Q_reg ( .D(n48), .SI(n8688), .SE(n4164), .CLK(n4506), .Q(
        n8687), .QN(n4019) );
  SDFFX1 DFF_208_Q_reg ( .D(n49), .SI(n8687), .SE(n4165), .CLK(n4506), .Q(
        n8686), .QN(n4018) );
  SDFFX1 DFF_209_Q_reg ( .D(n50), .SI(n8686), .SE(n4165), .CLK(n4506), .Q(
        n8685), .QN(n4017) );
  SDFFX1 DFF_210_Q_reg ( .D(n51), .SI(n8685), .SE(n4165), .CLK(n4506), .Q(
        n8684), .QN(n4016) );
  SDFFX1 DFF_211_Q_reg ( .D(n52), .SI(n8684), .SE(n4165), .CLK(n4506), .Q(
        n8683), .QN(n4015) );
  SDFFX1 DFF_212_Q_reg ( .D(n53), .SI(n8683), .SE(n4165), .CLK(n4506), .Q(
        n8682), .QN(n4014) );
  SDFFX1 DFF_213_Q_reg ( .D(n54), .SI(n8682), .SE(n4165), .CLK(n4506), .Q(
        n8681), .QN(n4013) );
  SDFFX1 DFF_214_Q_reg ( .D(n55), .SI(n8681), .SE(n4166), .CLK(n4505), .Q(
        n8680), .QN(n4012) );
  SDFFX1 DFF_215_Q_reg ( .D(n56), .SI(n8680), .SE(n4166), .CLK(n4505), .Q(
        test_so12), .QN(n4011) );
  SDFFX1 DFF_216_Q_reg ( .D(n57), .SI(test_si13), .SE(n4166), .CLK(n4505), .Q(
        n8677), .QN(n4010) );
  SDFFX1 DFF_217_Q_reg ( .D(n58), .SI(n8677), .SE(n4166), .CLK(n4505), .Q(
        n8676), .QN(n4009) );
  SDFFX1 DFF_218_Q_reg ( .D(n59), .SI(n8676), .SE(n4166), .CLK(n4505), .Q(
        n8675), .QN(n4008) );
  SDFFX1 DFF_219_Q_reg ( .D(n60), .SI(n8675), .SE(n4166), .CLK(n4505), .Q(
        n8674), .QN(n4007) );
  SDFFX1 DFF_220_Q_reg ( .D(n61), .SI(n8674), .SE(n4167), .CLK(n4505), .Q(
        n8673), .QN(n4006) );
  SDFFX1 DFF_221_Q_reg ( .D(n62), .SI(n8673), .SE(n4167), .CLK(n4505), .Q(
        n8672), .QN(n4005) );
  SDFFX1 DFF_222_Q_reg ( .D(n63), .SI(n8672), .SE(n4167), .CLK(n4505), .Q(
        n8671), .QN(n4004) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n4167), .CLK(n4505), .Q(
        n8670), .QN(n4003) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n3655), .CLK(n4633), .Q(
        n8669) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n4162), .CLK(n4507), .Q(
        n8668) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n4161), .CLK(n4508), .Q(
        n8667) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n4161), .CLK(n4508), .Q(
        n8666) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n4161), .CLK(n4508), .Q(
        n8665) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n4161), .CLK(n4508), .Q(
        n8664) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n4160), .CLK(n4508), .Q(
        n8663) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n4160), .CLK(n4508), .Q(
        n8662) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n4159), .CLK(n4509), .Q(
        n8661) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n4159), .CLK(n4509), .Q(
        test_so13) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n4159), .CLK(n4509), 
        .Q(n8658) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n4159), .CLK(n4509), .Q(
        n8657) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n4158), .CLK(n4509), .Q(
        n8656) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n4158), .CLK(n4509), .Q(
        n8655), .QN(n7234) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n3665), .CLK(n4628), .Q(
        n8654) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n3656), .CLK(n4632), .Q(
        n8653) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n4157), .CLK(n4510), .Q(
        WX1970), .QN(n3172) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n4157), .CLK(n4510), .Q(
        WX1972) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n4157), .CLK(n4510), .Q(
        WX1974), .QN(n3171) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n4156), .CLK(n4510), .Q(
        WX1976), .QN(n3170) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n4156), .CLK(n4510), .Q(
        WX1978), .QN(n3169) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n4156), .CLK(n4510), .Q(
        WX1980) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n4156), .CLK(n4510), .Q(
        WX1982), .QN(n3167) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n4156), .CLK(n4510), .Q(
        WX1984), .QN(n3166) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n4156), .CLK(n4510), .Q(
        WX1986), .QN(n3165) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n4155), .CLK(n4511), .Q(
        WX1988), .QN(n3164) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n4155), .CLK(n4511), .Q(
        WX1990), .QN(n3163) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n4155), .CLK(n4511), .Q(
        test_so14) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n3656), .CLK(n4632), 
        .Q(WX1994), .QN(n3162) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n3656), .CLK(n4632), .Q(
        WX1996), .QN(n3161) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n3656), .CLK(n4632), .Q(
        WX1998), .QN(n3160) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n4154), .CLK(n4511), .Q(
        WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n4154), .CLK(n4511), .Q(
        WX2002), .QN(n2845) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n4162), .CLK(n4507), .Q(
        WX2004), .QN(n3057) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n4162), .CLK(n4507), .Q(
        WX2006), .QN(n3055) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n4161), .CLK(n4508), .Q(
        WX2008), .QN(n3054) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n4161), .CLK(n4508), .Q(
        WX2010), .QN(n3052) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n4160), .CLK(n4508), .Q(
        WX2012), .QN(n3050) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n4160), .CLK(n4508), .Q(
        WX2014), .QN(n3048) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n4160), .CLK(n4508), .Q(
        WX2016), .QN(n3046) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n4160), .CLK(n4508), .Q(
        WX2018), .QN(n3044) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n4159), .CLK(n4509), .Q(
        WX2020), .QN(n3043) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n4159), .CLK(n4509), .Q(
        WX2022), .QN(n3041) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n4158), .CLK(n4509), .Q(
        WX2024), .QN(n3039) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n4158), .CLK(n4509), .Q(
        WX2026), .QN(n3037) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n4158), .CLK(n4509), .Q(
        test_so15) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n3665), .CLK(n4628), 
        .Q(WX2030), .QN(n3034) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n3665), .CLK(n4628), .Q(
        WX2032), .QN(n3032) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n3665), .CLK(n4628), .Q(
        WX2034) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n3665), .CLK(n4628), .Q(
        WX2036), .QN(n3783) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n3664), .CLK(n4629), .Q(
        WX2038) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n3664), .CLK(n4629), .Q(
        WX2040) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n3663), .CLK(n4629), .Q(
        WX2042) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n3663), .CLK(n4629), .Q(
        WX2044), .QN(n3775) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n3662), .CLK(n4630), .Q(
        WX2046) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n3662), .CLK(n4630), .Q(
        WX2048) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n3660), .CLK(n4630), .Q(
        WX2050) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n3660), .CLK(n4630), .Q(
        WX2052) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n3659), .CLK(n4631), .Q(
        WX2054) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n4155), .CLK(n4511), .Q(
        WX2056), .QN(n3763) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n4155), .CLK(n4511), .Q(
        WX2058) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n4155), .CLK(n4511), .Q(
        WX2060) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n4154), .CLK(n4511), .Q(
        WX2062) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n4154), .CLK(n4511), .Q(
        test_so16) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n4154), .CLK(n4511), 
        .Q(WX2066) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n4154), .CLK(n4511), .Q(
        WX2068) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n4153), .CLK(n4512), .Q(
        WX2070) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n4153), .CLK(n4512), .Q(
        WX2072) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n4153), .CLK(n4512), .Q(
        WX2074) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n4153), .CLK(n4512), .Q(
        WX2076) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n4152), .CLK(n4512), .Q(
        WX2078) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n4152), .CLK(n4512), .Q(
        WX2080) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n4152), .CLK(n4512), .Q(
        WX2082) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n4151), .CLK(n4513), .Q(
        WX2084), .QN(n7239) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n4151), .CLK(n4513), .Q(
        WX2086) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n4151), .CLK(n4513), .Q(
        WX2088) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n4150), .CLK(n4513), .Q(
        WX2090) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n4158), .CLK(n4509), .Q(
        WX2092), .QN(n3036) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n4157), .CLK(n4510), .Q(
        WX2094) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n4157), .CLK(n4510), .Q(
        WX2096) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n4157), .CLK(n4510), .Q(
        WX2098), .QN(n7230) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n3664), .CLK(n4629), .Q(
        test_so17) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n3664), .CLK(n4629), 
        .Q(WX2102), .QN(n7227) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n3663), .CLK(n4629), .Q(
        WX2104), .QN(n7226) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n3663), .CLK(n4629), .Q(
        WX2106), .QN(n7224) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n3662), .CLK(n4630), .Q(
        WX2108), .QN(n3168) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n3662), .CLK(n4630), .Q(
        WX2110), .QN(n7221) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n3660), .CLK(n4630), .Q(
        WX2112), .QN(n7220) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n3660), .CLK(n4630), .Q(
        WX2114), .QN(n7218) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n3659), .CLK(n4631), .Q(
        WX2116), .QN(n7217) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n3659), .CLK(n4631), .Q(
        WX2118), .QN(n7215) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n3659), .CLK(n4631), .Q(
        WX2120) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n3658), .CLK(n4631), .Q(
        WX2122), .QN(n7212) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n3658), .CLK(n4631), .Q(
        WX2124), .QN(n7210) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n3658), .CLK(n4631), .Q(
        WX2126), .QN(n7208) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n3657), .CLK(n4632), .Q(
        WX2128), .QN(n3159) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n3657), .CLK(n4632), .Q(
        WX2130), .QN(n3389) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n3657), .CLK(n4632), .Q(
        WX2132), .QN(n3390) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n3657), .CLK(n4632), .Q(
        WX2134), .QN(n3391) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n3656), .CLK(n4632), .Q(
        test_so18) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n4153), .CLK(n4512), 
        .Q(WX2138), .QN(n3392) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n4153), .CLK(n4512), .Q(
        WX2140), .QN(n3393) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n4152), .CLK(n4512), .Q(
        WX2142), .QN(n3394) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n4152), .CLK(n4512), .Q(
        WX2144), .QN(n3395) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n4152), .CLK(n4512), .Q(
        WX2146), .QN(n3396) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n4151), .CLK(n4513), .Q(
        WX2148), .QN(n3397) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n4151), .CLK(n4513), .Q(
        WX2150), .QN(n3398) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n4151), .CLK(n4513), .Q(
        WX2152), .QN(n3399) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n4150), .CLK(n4513), .Q(
        WX2154), .QN(n3400) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n4150), .CLK(n4513), .Q(
        WX2156), .QN(n3401) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n4150), .CLK(n4513), .Q(
        WX2158), .QN(n3402) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n4150), .CLK(n4513), .Q(
        WX2160), .QN(n3191) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n4150), .CLK(n4513), .Q(
        WX2162), .QN(n3403) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n3664), .CLK(n4629), .Q(
        WX2164), .QN(n3404) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n3664), .CLK(n4629), .Q(
        WX2166), .QN(n3405) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n3663), .CLK(n4629), .Q(
        WX2168), .QN(n3406) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n3663), .CLK(n4629), .Q(
        WX2170), .QN(n3192) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n3662), .CLK(n4630), .Q(
        test_so19) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n3662), .CLK(n4630), 
        .Q(WX2174), .QN(n3407) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n3660), .CLK(n4630), .Q(
        WX2176), .QN(n3408) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n3660), .CLK(n4630), .Q(
        WX2178), .QN(n3409) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n3659), .CLK(n4631), .Q(
        WX2180), .QN(n3410) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(n3659), .CLK(n4631), .Q(
        WX2182), .QN(n3411) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n3658), .CLK(n4631), .Q(
        WX2184), .QN(n3193) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n3658), .CLK(n4631), .Q(
        WX2186), .QN(n3412) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n3658), .CLK(n4631), .Q(
        WX2188), .QN(n3413) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n3657), .CLK(n4632), .Q(
        WX2190), .QN(n3414) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n3657), .CLK(n4632), .Q(
        WX2192), .QN(n3201) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n3668), .CLK(n4627), .Q(
        CRC_OUT_8_0) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n3668), .CLK(n4627), 
        .Q(CRC_OUT_8_1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n3668), .CLK(n4627), 
        .Q(CRC_OUT_8_2) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n3668), .CLK(n4627), 
        .Q(CRC_OUT_8_3), .QN(DFF_355_n1) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n3668), .CLK(n4627), 
        .Q(CRC_OUT_8_4) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n3667), .CLK(n4627), 
        .Q(CRC_OUT_8_5) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n3667), .CLK(n4627), 
        .Q(CRC_OUT_8_6) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n3667), .CLK(n4627), 
        .Q(test_so20) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n3667), .CLK(n4627), 
        .Q(CRC_OUT_8_8) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n3667), .CLK(n4627), 
        .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n3667), .CLK(n4627), 
        .Q(CRC_OUT_8_10), .QN(DFF_362_n1) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n3666), .CLK(n4628), .Q(CRC_OUT_8_11) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n3666), .CLK(n4628), .Q(CRC_OUT_8_12) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n3666), .CLK(n4628), .Q(CRC_OUT_8_13) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n3666), .CLK(n4628), .Q(CRC_OUT_8_14) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n3666), .CLK(n4628), .Q(CRC_OUT_8_15), .QN(DFF_367_n1) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n3666), .CLK(n4628), .Q(CRC_OUT_8_16) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n3665), .CLK(n4628), .Q(CRC_OUT_8_17) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n3656), .CLK(n4632), .Q(CRC_OUT_8_18) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n4149), .CLK(n4514), .Q(CRC_OUT_8_19) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n4149), .CLK(n4514), .Q(CRC_OUT_8_20) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n4149), .CLK(n4514), .Q(CRC_OUT_8_21) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n4149), .CLK(n4514), .Q(CRC_OUT_8_22) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n4149), .CLK(n4514), .Q(CRC_OUT_8_23) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n4149), .CLK(n4514), .Q(CRC_OUT_8_24) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n4148), .CLK(n4514), .Q(test_so21) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n4148), .CLK(n4514), 
        .Q(CRC_OUT_8_26) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n4148), .CLK(n4514), .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n4148), .CLK(n4514), .Q(CRC_OUT_8_28) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n4148), .CLK(n4514), .Q(CRC_OUT_8_29) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n4148), .CLK(n4514), .Q(CRC_OUT_8_30) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n4147), .CLK(n4515), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n95), .SI(CRC_OUT_8_31), .SE(n4147), .CLK(n4515), 
        .Q(WX3071), .QN(n3498) );
  SDFFX1 DFF_385_Q_reg ( .D(n96), .SI(WX3071), .SE(n4142), .CLK(n4517), .Q(
        n8644), .QN(n4002) );
  SDFFX1 DFF_386_Q_reg ( .D(n97), .SI(n8644), .SE(n4142), .CLK(n4517), .Q(
        n8643), .QN(n4001) );
  SDFFX1 DFF_387_Q_reg ( .D(n98), .SI(n8643), .SE(n4142), .CLK(n4517), .Q(
        n8642), .QN(n4000) );
  SDFFX1 DFF_388_Q_reg ( .D(n99), .SI(n8642), .SE(n4143), .CLK(n4517), .Q(
        n8641), .QN(n3999) );
  SDFFX1 DFF_389_Q_reg ( .D(n100), .SI(n8641), .SE(n4143), .CLK(n4517), .Q(
        n8640), .QN(n3998) );
  SDFFX1 DFF_390_Q_reg ( .D(n101), .SI(n8640), .SE(n4143), .CLK(n4517), .Q(
        n8639), .QN(n3997) );
  SDFFX1 DFF_391_Q_reg ( .D(n102), .SI(n8639), .SE(n4143), .CLK(n4517), .Q(
        n8638), .QN(n3996) );
  SDFFX1 DFF_392_Q_reg ( .D(n103), .SI(n8638), .SE(n4143), .CLK(n4517), .Q(
        n8637), .QN(n3995) );
  SDFFX1 DFF_393_Q_reg ( .D(n104), .SI(n8637), .SE(n4143), .CLK(n4517), .Q(
        n8636), .QN(n3994) );
  SDFFX1 DFF_394_Q_reg ( .D(n105), .SI(n8636), .SE(n4144), .CLK(n4516), .Q(
        n8635), .QN(n3993) );
  SDFFX1 DFF_395_Q_reg ( .D(n106), .SI(n8635), .SE(n4144), .CLK(n4516), .Q(
        test_so22), .QN(n3992) );
  SDFFX1 DFF_396_Q_reg ( .D(n107), .SI(test_si23), .SE(n4144), .CLK(n4516), 
        .Q(n8632), .QN(n3991) );
  SDFFX1 DFF_397_Q_reg ( .D(n108), .SI(n8632), .SE(n4144), .CLK(n4516), .Q(
        n8631), .QN(n3990) );
  SDFFX1 DFF_398_Q_reg ( .D(n109), .SI(n8631), .SE(n4144), .CLK(n4516), .Q(
        n8630), .QN(n3989) );
  SDFFX1 DFF_399_Q_reg ( .D(n110), .SI(n8630), .SE(n4144), .CLK(n4516), .Q(
        n8629), .QN(n3988) );
  SDFFX1 DFF_400_Q_reg ( .D(n112), .SI(n8629), .SE(n4145), .CLK(n4516), .Q(
        n8628), .QN(n3987) );
  SDFFX1 DFF_401_Q_reg ( .D(n113), .SI(n8628), .SE(n4145), .CLK(n4516), .Q(
        n8627), .QN(n3986) );
  SDFFX1 DFF_402_Q_reg ( .D(n114), .SI(n8627), .SE(n4145), .CLK(n4516), .Q(
        n8626), .QN(n3985) );
  SDFFX1 DFF_403_Q_reg ( .D(n115), .SI(n8626), .SE(n4145), .CLK(n4516), .Q(
        n8625), .QN(n3984) );
  SDFFX1 DFF_404_Q_reg ( .D(n116), .SI(n8625), .SE(n4145), .CLK(n4516), .Q(
        n8624), .QN(n3983) );
  SDFFX1 DFF_405_Q_reg ( .D(n117), .SI(n8624), .SE(n4145), .CLK(n4516), .Q(
        n8623), .QN(n3982) );
  SDFFX1 DFF_406_Q_reg ( .D(n118), .SI(n8623), .SE(n4146), .CLK(n4515), .Q(
        n8622), .QN(n3981) );
  SDFFX1 DFF_407_Q_reg ( .D(n119), .SI(n8622), .SE(n4146), .CLK(n4515), .Q(
        n8621), .QN(n3980) );
  SDFFX1 DFF_408_Q_reg ( .D(n120), .SI(n8621), .SE(n4146), .CLK(n4515), .Q(
        n8620), .QN(n3979) );
  SDFFX1 DFF_409_Q_reg ( .D(n121), .SI(n8620), .SE(n4146), .CLK(n4515), .Q(
        n8619), .QN(n3978) );
  SDFFX1 DFF_410_Q_reg ( .D(n122), .SI(n8619), .SE(n4146), .CLK(n4515), .Q(
        n8618), .QN(n3977) );
  SDFFX1 DFF_411_Q_reg ( .D(n123), .SI(n8618), .SE(n4146), .CLK(n4515), .Q(
        n8617), .QN(n3976) );
  SDFFX1 DFF_412_Q_reg ( .D(n124), .SI(n8617), .SE(n4147), .CLK(n4515), .Q(
        n8616), .QN(n3975) );
  SDFFX1 DFF_413_Q_reg ( .D(n125), .SI(n8616), .SE(n4147), .CLK(n4515), .Q(
        test_so23), .QN(n3974) );
  SDFFX1 DFF_414_Q_reg ( .D(n126), .SI(test_si24), .SE(n4147), .CLK(n4515), 
        .Q(n8613), .QN(n3973) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n4147), .CLK(n4515), .Q(
        n8612), .QN(n3972) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n4037), .CLK(n4570), .Q(
        n8611), .QN(n7249) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n4037), .CLK(n4570), .Q(
        n8610), .QN(n7248) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n3768), .CLK(n4580), .Q(
        n8609), .QN(n7247) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n3672), .CLK(n4625), .Q(
        n8608), .QN(n7246) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n3670), .CLK(n4626), .Q(
        n8607), .QN(n7245) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n4035), .CLK(n4571), .Q(
        n8606), .QN(n7244) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n4034), .CLK(n4571), .Q(
        n8605), .QN(n7243) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n4034), .CLK(n4571), .Q(
        n8604), .QN(n7242) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n3884), .CLK(n4572), .Q(
        n8603), .QN(n7241) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n3884), .CLK(n4572), .Q(
        n8602), .QN(n7240) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n3866), .CLK(n4572), .Q(
        n8601), .QN(n7238) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n3866), .CLK(n4572), .Q(
        n8600), .QN(n7237) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n3784), .CLK(n4573), .Q(
        n8599), .QN(n7236) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n3784), .CLK(n4573), .Q(
        n8598), .QN(n7235) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n4046), .CLK(n4565), .Q(
        n8597), .QN(n7233) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n3670), .CLK(n4626), .Q(
        test_so24) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n3670), .CLK(n4626), 
        .Q(WX3263), .QN(n3158) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n3670), .CLK(n4626), .Q(
        WX3265), .QN(n3157) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n3670), .CLK(n4626), .Q(
        WX3267), .QN(n3156) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n4044), .CLK(n4566), .Q(
        WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n4044), .CLK(n4566), .Q(
        WX3271), .QN(n3154) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n4044), .CLK(n4566), .Q(
        WX3273), .QN(n3153) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n4044), .CLK(n4566), .Q(
        WX3275), .QN(n3152) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n4043), .CLK(n4567), .Q(
        WX3277) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n4043), .CLK(n4567), .Q(
        WX3279), .QN(n3151) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n4042), .CLK(n4567), .Q(
        WX3281) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n4042), .CLK(n4567), .Q(
        WX3283), .QN(n3149) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n4041), .CLK(n4568), .Q(
        WX3285), .QN(n3148) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n4041), .CLK(n4568), .Q(
        WX3287), .QN(n3147) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n4040), .CLK(n4568), .Q(
        WX3289), .QN(n3146) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n4039), .CLK(n4569), .Q(
        WX3291), .QN(n3145) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n4039), .CLK(n4569), .Q(
        WX3293), .QN(n3144) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n4038), .CLK(n4569), .Q(
        WX3295), .QN(n2843) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n4037), .CLK(n4570), .Q(
        test_so25) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n3768), .CLK(n4580), 
        .Q(WX3299), .QN(n3029) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n3672), .CLK(n4625), .Q(
        WX3301), .QN(n3027) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n3670), .CLK(n4626), .Q(
        WX3303), .QN(n3025) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n4035), .CLK(n4571), .Q(
        WX3305), .QN(n3024) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n4035), .CLK(n4571), .Q(
        WX3307), .QN(n3022) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n4034), .CLK(n4571), .Q(
        WX3309), .QN(n3020) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n4034), .CLK(n4571), .Q(
        WX3311), .QN(n3019) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n3884), .CLK(n4572), .Q(
        WX3313), .QN(n3017) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n3866), .CLK(n4572), .Q(
        WX3315), .QN(n3015) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n3785), .CLK(n4573), .Q(
        WX3317), .QN(n3013) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n3785), .CLK(n4573), .Q(
        WX3319), .QN(n3011) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n3784), .CLK(n4573), .Q(
        WX3321), .QN(n3009) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n4045), .CLK(n4566), .Q(
        WX3323), .QN(n3007) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n4045), .CLK(n4566), .Q(
        WX3325), .QN(n3006) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n4045), .CLK(n4566), .Q(
        WX3327) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n4045), .CLK(n4566), .Q(
        WX3329) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n4045), .CLK(n4566), .Q(
        WX3331) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n4045), .CLK(n4566), .Q(
        test_so26) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n4044), .CLK(n4566), 
        .Q(WX3335) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n4044), .CLK(n4566), .Q(
        WX3337) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n4043), .CLK(n4567), .Q(
        WX3339) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n4043), .CLK(n4567), .Q(
        WX3341), .QN(n3739) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n4043), .CLK(n4567), .Q(
        WX3343) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n4042), .CLK(n4567), .Q(
        WX3345), .QN(n3735) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n4042), .CLK(n4567), .Q(
        WX3347) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n4041), .CLK(n4568), .Q(
        WX3349) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n4040), .CLK(n4568), .Q(
        WX3351) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n4040), .CLK(n4568), .Q(
        WX3353) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n4039), .CLK(n4569), .Q(
        WX3355) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n4038), .CLK(n4569), .Q(
        WX3357) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n4038), .CLK(n4569), .Q(
        WX3359) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n4037), .CLK(n4570), .Q(
        WX3361), .QN(n3031) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n4037), .CLK(n4570), .Q(
        WX3363) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n4036), .CLK(n4570), .Q(
        WX3365) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n4036), .CLK(n4570), .Q(
        WX3367) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n4036), .CLK(n4570), .Q(
        test_so27) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n4035), .CLK(n4571), 
        .Q(WX3371) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n4034), .CLK(n4571), .Q(
        WX3373) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n3884), .CLK(n4572), .Q(
        WX3375) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n3884), .CLK(n4572), .Q(
        WX3377) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n3866), .CLK(n4572), .Q(
        WX3379) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n3785), .CLK(n4573), .Q(
        WX3381) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n3785), .CLK(n4573), .Q(
        WX3383) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n3784), .CLK(n4573), .Q(
        WX3385) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n3784), .CLK(n4573), .Q(
        WX3387) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(n3782), .CLK(n4574), .Q(
        WX3389), .QN(n7232) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n3782), .CLK(n4574), .Q(
        WX3391), .QN(n7231) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(n3782), .CLK(n4574), .Q(
        WX3393), .QN(n7229) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n3781), .CLK(n4574), .Q(
        WX3395), .QN(n7228) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n3781), .CLK(n4574), .Q(
        WX3397), .QN(n3155) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n3781), .CLK(n4574), .Q(
        WX3399), .QN(n7225) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n3780), .CLK(n4575), .Q(
        WX3401), .QN(n7223) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n3780), .CLK(n4575), .Q(
        WX3403), .QN(n7222) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n3780), .CLK(n4575), .Q(
        test_so28) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n4043), .CLK(n4567), 
        .Q(WX3407), .QN(n7219) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n4042), .CLK(n4567), .Q(
        WX3409), .QN(n3150) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n4042), .CLK(n4567), .Q(
        WX3411), .QN(n7216) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n4041), .CLK(n4568), .Q(
        WX3413), .QN(n7214) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n4040), .CLK(n4568), .Q(
        WX3415), .QN(n7213) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n4040), .CLK(n4568), .Q(
        WX3417), .QN(n7211) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n4039), .CLK(n4569), .Q(
        WX3419), .QN(n7209) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n4038), .CLK(n4569), .Q(
        WX3421), .QN(n7207) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n4038), .CLK(n4569), .Q(
        WX3423), .QN(n3363) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n4037), .CLK(n4570), .Q(
        WX3425), .QN(n3364) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n4036), .CLK(n4570), .Q(
        WX3427), .QN(n3365) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n4036), .CLK(n4570), .Q(
        WX3429), .QN(n3366) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n4036), .CLK(n4570), .Q(
        WX3431), .QN(n3367) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n4035), .CLK(n4571), .Q(
        WX3433), .QN(n3368) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n4035), .CLK(n4571), .Q(
        WX3435), .QN(n3369) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n4034), .CLK(n4571), .Q(
        WX3437), .QN(n3370) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n3884), .CLK(n4572), .Q(
        test_so29) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n3866), .CLK(n4572), 
        .Q(WX3441), .QN(n3371) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n3866), .CLK(n4572), .Q(
        WX3443), .QN(n3372) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n3785), .CLK(n4573), .Q(
        WX3445), .QN(n3373) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n3785), .CLK(n4573), .Q(
        WX3447), .QN(n3374) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n3784), .CLK(n4573), .Q(
        WX3449), .QN(n3375) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n3782), .CLK(n4574), .Q(
        WX3451), .QN(n3376) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n3782), .CLK(n4574), .Q(
        WX3453), .QN(n3188) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n3782), .CLK(n4574), .Q(
        WX3455), .QN(n3377) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n3781), .CLK(n4574), .Q(
        WX3457), .QN(n3378) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n3781), .CLK(n4574), .Q(
        WX3459), .QN(n3379) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n3781), .CLK(n4574), .Q(
        WX3461), .QN(n3380) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n3780), .CLK(n4575), .Q(
        WX3463), .QN(n3189) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n3780), .CLK(n4575), .Q(
        WX3465), .QN(n3381) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n3780), .CLK(n4575), .Q(
        WX3467), .QN(n3382) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n3779), .CLK(n4575), .Q(
        WX3469), .QN(n3383) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n3779), .CLK(n4575), .Q(
        WX3471), .QN(n3384) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n3779), .CLK(n4575), .Q(
        test_so30) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n4041), .CLK(n4568), 
        .Q(WX3475), .QN(n3385) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n4041), .CLK(n4568), .Q(
        WX3477), .QN(n3190) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n4040), .CLK(n4568), .Q(
        WX3479), .QN(n3386) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n4039), .CLK(n4569), .Q(
        WX3481), .QN(n3387) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n4039), .CLK(n4569), .Q(
        WX3483), .QN(n3388) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n4038), .CLK(n4569), .Q(
        WX3485), .QN(n3200) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n3672), .CLK(n4625), .Q(
        CRC_OUT_7_0) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n3672), .CLK(n4625), 
        .Q(CRC_OUT_7_1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n3671), .CLK(n4626), 
        .Q(CRC_OUT_7_2) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n3671), .CLK(n4626), 
        .Q(CRC_OUT_7_3), .QN(DFF_547_n1) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n3671), .CLK(n4626), 
        .Q(CRC_OUT_7_4) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n3671), .CLK(n4626), 
        .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n3671), .CLK(n4626), 
        .Q(CRC_OUT_7_6) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n3671), .CLK(n4626), 
        .Q(CRC_OUT_7_7) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n3779), .CLK(n4575), 
        .Q(CRC_OUT_7_8) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n3779), .CLK(n4575), 
        .Q(CRC_OUT_7_9) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n3779), .CLK(n4575), 
        .Q(test_so31) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n3778), .CLK(n4576), 
        .Q(CRC_OUT_7_11) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n3778), .CLK(n4576), .Q(CRC_OUT_7_12) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n3778), .CLK(n4576), .Q(CRC_OUT_7_13) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n3778), .CLK(n4576), .Q(CRC_OUT_7_14) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n3778), .CLK(n4576), .Q(CRC_OUT_7_15), .QN(DFF_559_n1) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n3778), .CLK(n4576), .Q(CRC_OUT_7_16) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n3777), .CLK(n4576), .Q(CRC_OUT_7_17) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n3777), .CLK(n4576), .Q(CRC_OUT_7_18) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n3777), .CLK(n4576), .Q(CRC_OUT_7_19) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n3777), .CLK(n4576), .Q(CRC_OUT_7_20) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n3777), .CLK(n4576), .Q(CRC_OUT_7_21) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n3777), .CLK(n4576), .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n3776), .CLK(n4577), .Q(CRC_OUT_7_23) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n3776), .CLK(n4577), .Q(CRC_OUT_7_24) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n3776), .CLK(n4577), .Q(CRC_OUT_7_25) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n3776), .CLK(n4577), .Q(CRC_OUT_7_26) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n3776), .CLK(n4577), .Q(test_so32) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n3776), .CLK(n4577), 
        .Q(CRC_OUT_7_28) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n3774), .CLK(n4577), .Q(CRC_OUT_7_29) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n3774), .CLK(n4577), .Q(CRC_OUT_7_30) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n3774), .CLK(n4577), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n158), .SI(CRC_OUT_7_31), .SE(n3774), .CLK(n4577), 
        .Q(WX4364), .QN(n3500) );
  SDFFX1 DFF_577_Q_reg ( .D(n159), .SI(WX4364), .SE(n3769), .CLK(n4580), .Q(
        n8586), .QN(n3971) );
  SDFFX1 DFF_578_Q_reg ( .D(n160), .SI(n8586), .SE(n3769), .CLK(n4580), .Q(
        n8585), .QN(n3970) );
  SDFFX1 DFF_579_Q_reg ( .D(n161), .SI(n8585), .SE(n3769), .CLK(n4580), .Q(
        n8584), .QN(n3969) );
  SDFFX1 DFF_580_Q_reg ( .D(n162), .SI(n8584), .SE(n3769), .CLK(n4580), .Q(
        n8583), .QN(n3968) );
  SDFFX1 DFF_581_Q_reg ( .D(n163), .SI(n8583), .SE(n3769), .CLK(n4580), .Q(
        n8582), .QN(n3967) );
  SDFFX1 DFF_582_Q_reg ( .D(n164), .SI(n8582), .SE(n3770), .CLK(n4579), .Q(
        n8581), .QN(n3966) );
  SDFFX1 DFF_583_Q_reg ( .D(n165), .SI(n8581), .SE(n3770), .CLK(n4579), .Q(
        n8580), .QN(n3965) );
  SDFFX1 DFF_584_Q_reg ( .D(n166), .SI(n8580), .SE(n3770), .CLK(n4579), .Q(
        n8579), .QN(n3964) );
  SDFFX1 DFF_585_Q_reg ( .D(n167), .SI(n8579), .SE(n3770), .CLK(n4579), .Q(
        n8578), .QN(n3963) );
  SDFFX1 DFF_586_Q_reg ( .D(n168), .SI(n8578), .SE(n3770), .CLK(n4579), .Q(
        n8577), .QN(n3962) );
  SDFFX1 DFF_587_Q_reg ( .D(n169), .SI(n8577), .SE(n3770), .CLK(n4579), .Q(
        n8576), .QN(n3961) );
  SDFFX1 DFF_588_Q_reg ( .D(n170), .SI(n8576), .SE(n3771), .CLK(n4579), .Q(
        test_so33), .QN(n3960) );
  SDFFX1 DFF_589_Q_reg ( .D(n171), .SI(test_si34), .SE(n3771), .CLK(n4579), 
        .Q(n8573), .QN(n3959) );
  SDFFX1 DFF_590_Q_reg ( .D(n172), .SI(n8573), .SE(n3771), .CLK(n4579), .Q(
        n8572), .QN(n3958) );
  SDFFX1 DFF_591_Q_reg ( .D(n173), .SI(n8572), .SE(n3771), .CLK(n4579), .Q(
        n8571), .QN(n3957) );
  SDFFX1 DFF_592_Q_reg ( .D(n174), .SI(n8571), .SE(n3771), .CLK(n4579), .Q(
        n8570), .QN(n3956) );
  SDFFX1 DFF_593_Q_reg ( .D(n175), .SI(n8570), .SE(n3771), .CLK(n4579), .Q(
        n8569), .QN(n3955) );
  SDFFX1 DFF_594_Q_reg ( .D(n176), .SI(n8569), .SE(n3772), .CLK(n4578), .Q(
        n8568), .QN(n3954) );
  SDFFX1 DFF_595_Q_reg ( .D(n177), .SI(n8568), .SE(n3772), .CLK(n4578), .Q(
        n8567), .QN(n3953) );
  SDFFX1 DFF_596_Q_reg ( .D(n178), .SI(n8567), .SE(n3772), .CLK(n4578), .Q(
        n8566), .QN(n3952) );
  SDFFX1 DFF_597_Q_reg ( .D(n179), .SI(n8566), .SE(n3772), .CLK(n4578), .Q(
        n8565), .QN(n3951) );
  SDFFX1 DFF_598_Q_reg ( .D(n180), .SI(n8565), .SE(n3772), .CLK(n4578), .Q(
        n8564), .QN(n3950) );
  SDFFX1 DFF_599_Q_reg ( .D(n181), .SI(n8564), .SE(n3772), .CLK(n4578), .Q(
        n8563), .QN(n3949) );
  SDFFX1 DFF_600_Q_reg ( .D(n182), .SI(n8563), .SE(n3773), .CLK(n4578), .Q(
        n8562), .QN(n3948) );
  SDFFX1 DFF_601_Q_reg ( .D(n183), .SI(n8562), .SE(n3773), .CLK(n4578), .Q(
        n8561), .QN(n3947) );
  SDFFX1 DFF_602_Q_reg ( .D(n184), .SI(n8561), .SE(n3773), .CLK(n4578), .Q(
        n8560), .QN(n3946) );
  SDFFX1 DFF_603_Q_reg ( .D(n185), .SI(n8560), .SE(n3773), .CLK(n4578), .Q(
        n8559), .QN(n3945) );
  SDFFX1 DFF_604_Q_reg ( .D(n186), .SI(n8559), .SE(n3773), .CLK(n4578), .Q(
        n8558), .QN(n3944) );
  SDFFX1 DFF_605_Q_reg ( .D(n187), .SI(n8558), .SE(n3773), .CLK(n4578), .Q(
        test_so34), .QN(n3943) );
  SDFFX1 DFF_606_Q_reg ( .D(n188), .SI(test_si35), .SE(n3774), .CLK(n4577), 
        .Q(n8555), .QN(n3942) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n3774), .CLK(n4577), .Q(
        n8554), .QN(n3941) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n3677), .CLK(n4623), .Q(
        n8553), .QN(n7206) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n3769), .CLK(n4580), .Q(
        n8552), .QN(n7205) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n3768), .CLK(n4580), .Q(
        n8551), .QN(n7204) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n3767), .CLK(n4581), .Q(
        n8550), .QN(n7203) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n3766), .CLK(n4581), .Q(
        n8549), .QN(n7202) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n3766), .CLK(n4581), .Q(
        n8548), .QN(n7201) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n3765), .CLK(n4582), .Q(
        n8547), .QN(n7200) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n3765), .CLK(n4582), .Q(
        n8546), .QN(n7199) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n3764), .CLK(n4582), .Q(
        n8545), .QN(n7198) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n3764), .CLK(n4582), .Q(
        n8544), .QN(n7197) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n3761), .CLK(n4583), .Q(
        n8543), .QN(n7196) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n3761), .CLK(n4583), .Q(
        n8542), .QN(n7195) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n3760), .CLK(n4584), .Q(
        n8541), .QN(n7194) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n3760), .CLK(n4584), .Q(
        n8540), .QN(n7193) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n4046), .CLK(n4565), .Q(
        test_so35) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n3758), .CLK(n4585), 
        .Q(n8537), .QN(n7191) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n3758), .CLK(n4585), .Q(
        WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n3757), .CLK(n4585), .Q(
        WX4558), .QN(n3142) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n3757), .CLK(n4585), .Q(
        WX4560) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n3756), .CLK(n4586), .Q(
        WX4562), .QN(n3141) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n3755), .CLK(n4586), .Q(
        WX4564) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n3755), .CLK(n4586), .Q(
        WX4566), .QN(n3139) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n3754), .CLK(n4587), .Q(
        WX4568), .QN(n3138) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n3753), .CLK(n4587), .Q(
        WX4570), .QN(n3137) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n3753), .CLK(n4587), .Q(
        WX4572), .QN(n3136) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n3752), .CLK(n4588), .Q(
        WX4574), .QN(n3135) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n3751), .CLK(n4588), .Q(
        WX4576), .QN(n3134) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n3751), .CLK(n4588), .Q(
        WX4578), .QN(n3133) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n3750), .CLK(n4589), .Q(
        WX4580), .QN(n3132) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n3749), .CLK(n4589), .Q(
        WX4582), .QN(n3131) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n3749), .CLK(n4589), .Q(
        WX4584), .QN(n3130) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n3748), .CLK(n4590), .Q(
        test_so36) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n3677), .CLK(n4623), 
        .Q(WX4588), .QN(n2841) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n3768), .CLK(n4580), .Q(
        WX4590), .QN(n3005) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n3768), .CLK(n4580), .Q(
        WX4592), .QN(n3003) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n3767), .CLK(n4581), .Q(
        WX4594), .QN(n3002) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n3767), .CLK(n4581), .Q(
        WX4596), .QN(n3000) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n3766), .CLK(n4581), .Q(
        WX4598), .QN(n2998) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n3766), .CLK(n4581), .Q(
        WX4600), .QN(n2996) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n3765), .CLK(n4582), .Q(
        WX4602), .QN(n2994) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n3764), .CLK(n4582), .Q(
        WX4604), .QN(n2992) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n3762), .CLK(n4583), .Q(
        WX4606), .QN(n2990) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n3762), .CLK(n4583), .Q(
        WX4608), .QN(n2988) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n3761), .CLK(n4583), .Q(
        WX4610), .QN(n2986) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n3761), .CLK(n4583), .Q(
        WX4612), .QN(n2984) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n3760), .CLK(n4584), .Q(
        WX4614), .QN(n2982) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n3759), .CLK(n4584), .Q(
        WX4616), .QN(n2981) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n3759), .CLK(n4584), .Q(
        WX4618), .QN(n2979) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n3758), .CLK(n4585), .Q(
        test_so37) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n3757), .CLK(n4585), 
        .Q(WX4622) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n3757), .CLK(n4585), .Q(
        WX4624), .QN(n3717) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n3756), .CLK(n4586), .Q(
        WX4626) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n3755), .CLK(n4586), .Q(
        WX4628), .QN(n3713) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n3755), .CLK(n4586), .Q(
        WX4630) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n3754), .CLK(n4587), .Q(
        WX4632) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n3753), .CLK(n4587), .Q(
        WX4634) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n3753), .CLK(n4587), .Q(
        WX4636) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n3752), .CLK(n4588), .Q(
        WX4638) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n3751), .CLK(n4588), .Q(
        WX4640) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n3751), .CLK(n4588), .Q(
        WX4642) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n3750), .CLK(n4589), .Q(
        WX4644) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n3749), .CLK(n4589), .Q(
        WX4646) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n3749), .CLK(n4589), .Q(
        WX4648) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n3748), .CLK(n4590), .Q(
        WX4650), .QN(n3691) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n3747), .CLK(n4590), .Q(
        WX4652) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n3747), .CLK(n4590), .Q(
        test_so38) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n3768), .CLK(n4580), 
        .Q(WX4656) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n3767), .CLK(n4581), .Q(
        WX4658) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n3767), .CLK(n4581), .Q(
        WX4660) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n3766), .CLK(n4581), .Q(
        WX4662) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n3765), .CLK(n4582), .Q(
        WX4664) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n3765), .CLK(n4582), .Q(
        WX4666) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n3764), .CLK(n4582), .Q(
        WX4668) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n3762), .CLK(n4583), .Q(
        WX4670) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n3762), .CLK(n4583), .Q(
        WX4672) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n3761), .CLK(n4583), .Q(
        WX4674) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n3760), .CLK(n4584), .Q(
        WX4676) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n3760), .CLK(n4584), .Q(
        WX4678) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n3759), .CLK(n4584), .Q(
        WX4680), .QN(n7192) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n3759), .CLK(n4584), .Q(
        WX4682) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n3758), .CLK(n4585), .Q(
        WX4684), .QN(n3143) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n3757), .CLK(n4585), .Q(
        WX4686), .QN(n7190) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n3756), .CLK(n4586), .Q(
        test_so39) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n3756), .CLK(n4586), 
        .Q(WX4690), .QN(n7189) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n3755), .CLK(n4586), .Q(
        WX4692), .QN(n3140) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n3754), .CLK(n4587), .Q(
        WX4694), .QN(n7188) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n3754), .CLK(n4587), .Q(
        WX4696), .QN(n7187) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n3753), .CLK(n4587), .Q(
        WX4698), .QN(n7186) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n3752), .CLK(n4588), .Q(
        WX4700), .QN(n7185) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n3752), .CLK(n4588), .Q(
        WX4702), .QN(n7184) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n3751), .CLK(n4588), .Q(
        WX4704), .QN(n7183) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n3750), .CLK(n4589), .Q(
        WX4706), .QN(n7182) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n3750), .CLK(n4589), .Q(
        WX4708), .QN(n7181) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n3749), .CLK(n4589), .Q(
        WX4710), .QN(n7180) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n3748), .CLK(n4590), .Q(
        WX4712), .QN(n7179) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n3748), .CLK(n4590), .Q(
        WX4714) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n3747), .CLK(n4590), .Q(
        WX4716), .QN(n3336) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n3747), .CLK(n4590), .Q(
        WX4718), .QN(n3337) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n3747), .CLK(n4590), .Q(
        WX4720), .QN(n3338) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n3747), .CLK(n4590), .Q(
        test_so40) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n3767), .CLK(n4581), 
        .Q(WX4724), .QN(n3339) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n3766), .CLK(n4581), .Q(
        WX4726), .QN(n3340) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n3765), .CLK(n4582), .Q(
        WX4728), .QN(n3341) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n3764), .CLK(n4582), .Q(
        WX4730), .QN(n3342) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n3764), .CLK(n4582), .Q(
        WX4732), .QN(n3343) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n3762), .CLK(n4583), .Q(
        WX4734), .QN(n3344) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n3762), .CLK(n4583), .Q(
        WX4736), .QN(n3345) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n3761), .CLK(n4583), .Q(
        WX4738), .QN(n3346) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n3760), .CLK(n4584), .Q(
        WX4740), .QN(n3347) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n3759), .CLK(n4584), .Q(
        WX4742), .QN(n3348) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n3759), .CLK(n4584), .Q(
        WX4744), .QN(n3349) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n3758), .CLK(n4585), .Q(
        WX4746), .QN(n3186) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n3758), .CLK(n4585), .Q(
        WX4748), .QN(n3350) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n3757), .CLK(n4585), .Q(
        WX4750), .QN(n3351) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n3756), .CLK(n4586), .Q(
        WX4752), .QN(n3352) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n3756), .CLK(n4586), .Q(
        WX4754), .QN(n3353) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n3755), .CLK(n4586), .Q(
        test_so41) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n3754), .CLK(n4587), 
        .Q(WX4758), .QN(n3354) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n3754), .CLK(n4587), .Q(
        WX4760), .QN(n3355) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n3753), .CLK(n4587), .Q(
        WX4762), .QN(n3356) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n3752), .CLK(n4588), .Q(
        WX4764), .QN(n3357) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n3752), .CLK(n4588), .Q(
        WX4766), .QN(n3358) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n3751), .CLK(n4588), .Q(
        WX4768), .QN(n3359) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n3750), .CLK(n4589), .Q(
        WX4770), .QN(n3187) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n3750), .CLK(n4589), .Q(
        WX4772), .QN(n3360) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n3749), .CLK(n4589), .Q(
        WX4774), .QN(n3361) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n3748), .CLK(n4590), .Q(
        WX4776), .QN(n3362) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n3748), .CLK(n4590), .Q(
        WX4778), .QN(n3199) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n3677), .CLK(n4623), .Q(
        CRC_OUT_6_0) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n3677), .CLK(n4623), 
        .Q(CRC_OUT_6_1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n3677), .CLK(n4623), 
        .Q(CRC_OUT_6_2) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n3677), .CLK(n4623), 
        .Q(CRC_OUT_6_3), .QN(DFF_739_n1) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n3676), .CLK(n4623), 
        .Q(CRC_OUT_6_4) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n3676), .CLK(n4623), 
        .Q(test_so42) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n3676), .CLK(n4623), 
        .Q(CRC_OUT_6_6) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n3676), .CLK(n4623), 
        .Q(CRC_OUT_6_7) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n3676), .CLK(n4623), 
        .Q(CRC_OUT_6_8) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n3676), .CLK(n4623), 
        .Q(CRC_OUT_6_9) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n3675), .CLK(n4624), 
        .Q(CRC_OUT_6_10) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n3675), .CLK(n4624), .Q(CRC_OUT_6_11) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n3675), .CLK(n4624), .Q(CRC_OUT_6_12) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n3675), .CLK(n4624), .Q(CRC_OUT_6_13) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n3675), .CLK(n4624), .Q(CRC_OUT_6_14) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n3675), .CLK(n4624), .Q(CRC_OUT_6_15), .QN(DFF_751_n1) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n3674), .CLK(n4624), .Q(CRC_OUT_6_16) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n3674), .CLK(n4624), .Q(CRC_OUT_6_17) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n3674), .CLK(n4624), .Q(CRC_OUT_6_18) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n3674), .CLK(n4624), .Q(CRC_OUT_6_19) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n3674), .CLK(n4624), .Q(CRC_OUT_6_20) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n3674), .CLK(n4624), .Q(CRC_OUT_6_21) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n3673), .CLK(n4625), .Q(test_so43) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n3673), .CLK(n4625), 
        .Q(CRC_OUT_6_23) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n3673), .CLK(n4625), .Q(CRC_OUT_6_24) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n3673), .CLK(n4625), .Q(CRC_OUT_6_25) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n3673), .CLK(n4625), .Q(CRC_OUT_6_26) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n3673), .CLK(n4625), .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n3672), .CLK(n4625), .Q(CRC_OUT_6_28) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n3672), .CLK(n4625), .Q(CRC_OUT_6_29) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n3746), .CLK(n4591), .Q(CRC_OUT_6_30) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n3746), .CLK(n4591), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n220), .SI(CRC_OUT_6_31), .SE(n3746), .CLK(n4591), 
        .Q(WX5657), .QN(n3502) );
  SDFFX1 DFF_769_Q_reg ( .D(n221), .SI(WX5657), .SE(n3741), .CLK(n4593), .Q(
        n8528), .QN(n3940) );
  SDFFX1 DFF_770_Q_reg ( .D(n222), .SI(n8528), .SE(n3741), .CLK(n4593), .Q(
        n8527), .QN(n3939) );
  SDFFX1 DFF_771_Q_reg ( .D(n223), .SI(n8527), .SE(n3741), .CLK(n4593), .Q(
        n8526), .QN(n3938) );
  SDFFX1 DFF_772_Q_reg ( .D(n224), .SI(n8526), .SE(n3741), .CLK(n4593), .Q(
        n8525), .QN(n3937) );
  SDFFX1 DFF_773_Q_reg ( .D(n225), .SI(n8525), .SE(n3742), .CLK(n4593), .Q(
        n8524), .QN(n3936) );
  SDFFX1 DFF_774_Q_reg ( .D(n226), .SI(n8524), .SE(n3742), .CLK(n4593), .Q(
        n8523), .QN(n3935) );
  SDFFX1 DFF_775_Q_reg ( .D(n227), .SI(n8523), .SE(n3742), .CLK(n4593), .Q(
        test_so44), .QN(n3934) );
  SDFFX1 DFF_776_Q_reg ( .D(n228), .SI(test_si45), .SE(n3742), .CLK(n4593), 
        .Q(n8520), .QN(n3933) );
  SDFFX1 DFF_777_Q_reg ( .D(n229), .SI(n8520), .SE(n3742), .CLK(n4593), .Q(
        n8519), .QN(n3932) );
  SDFFX1 DFF_778_Q_reg ( .D(n230), .SI(n8519), .SE(n3742), .CLK(n4593), .Q(
        n8518), .QN(n3931) );
  SDFFX1 DFF_779_Q_reg ( .D(n231), .SI(n8518), .SE(n3743), .CLK(n4592), .Q(
        n8517), .QN(n3930) );
  SDFFX1 DFF_780_Q_reg ( .D(n232), .SI(n8517), .SE(n3743), .CLK(n4592), .Q(
        n8516), .QN(n3929) );
  SDFFX1 DFF_781_Q_reg ( .D(n233), .SI(n8516), .SE(n3743), .CLK(n4592), .Q(
        n8515), .QN(n3928) );
  SDFFX1 DFF_782_Q_reg ( .D(n234), .SI(n8515), .SE(n3743), .CLK(n4592), .Q(
        n8514), .QN(n3927) );
  SDFFX1 DFF_783_Q_reg ( .D(n235), .SI(n8514), .SE(n3743), .CLK(n4592), .Q(
        n8513), .QN(n3926) );
  SDFFX1 DFF_784_Q_reg ( .D(n236), .SI(n8513), .SE(n3743), .CLK(n4592), .Q(
        n8512), .QN(n3925) );
  SDFFX1 DFF_785_Q_reg ( .D(n237), .SI(n8512), .SE(n3744), .CLK(n4592), .Q(
        n8511), .QN(n3924) );
  SDFFX1 DFF_786_Q_reg ( .D(n238), .SI(n8511), .SE(n3744), .CLK(n4592), .Q(
        n8510), .QN(n3923) );
  SDFFX1 DFF_787_Q_reg ( .D(n239), .SI(n8510), .SE(n3744), .CLK(n4592), .Q(
        n8509), .QN(n3922) );
  SDFFX1 DFF_788_Q_reg ( .D(n240), .SI(n8509), .SE(n3744), .CLK(n4592), .Q(
        n8508), .QN(n3921) );
  SDFFX1 DFF_789_Q_reg ( .D(n241), .SI(n8508), .SE(n3744), .CLK(n4592), .Q(
        n8507), .QN(n3920) );
  SDFFX1 DFF_790_Q_reg ( .D(n242), .SI(n8507), .SE(n3744), .CLK(n4592), .Q(
        n8506), .QN(n3919) );
  SDFFX1 DFF_791_Q_reg ( .D(n243), .SI(n8506), .SE(n3745), .CLK(n4591), .Q(
        n8505), .QN(n3918) );
  SDFFX1 DFF_792_Q_reg ( .D(n244), .SI(n8505), .SE(n3745), .CLK(n4591), .Q(
        test_so45), .QN(n3917) );
  SDFFX1 DFF_793_Q_reg ( .D(n245), .SI(test_si46), .SE(n3745), .CLK(n4591), 
        .Q(n8502), .QN(n3916) );
  SDFFX1 DFF_794_Q_reg ( .D(n246), .SI(n8502), .SE(n3745), .CLK(n4591), .Q(
        n8501), .QN(n3915) );
  SDFFX1 DFF_795_Q_reg ( .D(n247), .SI(n8501), .SE(n3745), .CLK(n4591), .Q(
        n8500), .QN(n3914) );
  SDFFX1 DFF_796_Q_reg ( .D(n248), .SI(n8500), .SE(n3745), .CLK(n4591), .Q(
        n8499), .QN(n3913) );
  SDFFX1 DFF_797_Q_reg ( .D(n249), .SI(n8499), .SE(n3746), .CLK(n4591), .Q(
        n8498), .QN(n3912) );
  SDFFX1 DFF_798_Q_reg ( .D(n250), .SI(n8498), .SE(n3746), .CLK(n4591), .Q(
        n8497), .QN(n3911) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n3746), .CLK(n4591), .Q(
        n8496), .QN(n3910) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n3678), .CLK(n4622), .Q(
        n8495), .QN(n7178) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n3741), .CLK(n4593), .Q(
        n8494), .QN(n7177) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n3740), .CLK(n4594), .Q(
        n8493), .QN(n7176) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n3740), .CLK(n4594), .Q(
        n8492), .QN(n7175) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n3740), .CLK(n4594), .Q(
        n8491), .QN(n7174) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n3738), .CLK(n4594), .Q(
        n8490), .QN(n7173) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n3738), .CLK(n4594), .Q(
        n8489), .QN(n7172) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n3738), .CLK(n4594), .Q(
        n8488), .QN(n7171) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n3737), .CLK(n4595), .Q(
        n8487), .QN(n7170) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n3737), .CLK(n4595), .Q(
        test_so46) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n3737), .CLK(n4595), 
        .Q(n8484), .QN(n7168) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n3736), .CLK(n4595), .Q(
        n8483), .QN(n7167) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n3678), .CLK(n4622), .Q(
        n8482), .QN(n7166) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n3736), .CLK(n4595), .Q(
        n8481), .QN(n7165) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n4046), .CLK(n4565), .Q(
        n8480), .QN(n7164) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n3734), .CLK(n4596), .Q(
        n8479), .QN(n7163) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n3733), .CLK(n4596), .Q(
        WX5849), .QN(n3129) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n3733), .CLK(n4596), .Q(
        WX5851), .QN(n3128) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n3732), .CLK(n4597), .Q(
        WX5853), .QN(n3127) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n3731), .CLK(n4597), .Q(
        WX5855), .QN(n3126) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n3731), .CLK(n4597), .Q(
        WX5857), .QN(n3125) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n3730), .CLK(n4598), .Q(
        WX5859), .QN(n3124) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n3729), .CLK(n4598), .Q(
        WX5861), .QN(n3123) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n3729), .CLK(n4598), .Q(
        WX5863), .QN(n3122) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n3728), .CLK(n4599), .Q(
        WX5865), .QN(n3121) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n3727), .CLK(n4599), .Q(
        WX5867), .QN(n3120) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n3727), .CLK(n4599), .Q(
        test_so47) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n3681), .CLK(n4621), 
        .Q(WX5871), .QN(n3119) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n3725), .CLK(n4600), .Q(
        WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n3725), .CLK(n4600), .Q(
        WX5875), .QN(n3117) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n3724), .CLK(n4601), .Q(
        WX5877) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n3724), .CLK(n4601), .Q(
        WX5879), .QN(n3116) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n3723), .CLK(n4601), .Q(
        WX5881), .QN(n2839) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n3741), .CLK(n4593), .Q(
        WX5883), .QN(n2977) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n3740), .CLK(n4594), .Q(
        WX5885), .QN(n2975) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n3740), .CLK(n4594), .Q(
        WX5887), .QN(n2973) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n3740), .CLK(n4594), .Q(
        WX5889), .QN(n2971) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n3738), .CLK(n4594), .Q(
        WX5891), .QN(n2969) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n3738), .CLK(n4594), .Q(
        WX5893), .QN(n2967) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n3738), .CLK(n4594), .Q(
        WX5895), .QN(n2965) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n3737), .CLK(n4595), .Q(
        WX5897), .QN(n2963) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n3737), .CLK(n4595), .Q(
        WX5899), .QN(n2962) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n3737), .CLK(n4595), .Q(
        WX5901), .QN(n2960) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n3736), .CLK(n4595), .Q(
        test_so48) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n3678), .CLK(n4622), 
        .Q(WX5905), .QN(n2957) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n3734), .CLK(n4596), .Q(
        WX5907), .QN(n2956) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n3734), .CLK(n4596), .Q(
        WX5909), .QN(n2954) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n3734), .CLK(n4596), .Q(
        WX5911), .QN(n2953) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n3733), .CLK(n4596), .Q(
        WX5913) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n3733), .CLK(n4596), .Q(
        WX5915) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n3732), .CLK(n4597), .Q(
        WX5917) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n3731), .CLK(n4597), .Q(
        WX5919) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n3731), .CLK(n4597), .Q(
        WX5921) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n3730), .CLK(n4598), .Q(
        WX5923) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n3729), .CLK(n4598), .Q(
        WX5925) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n3729), .CLK(n4598), .Q(
        WX5927) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n3728), .CLK(n4599), .Q(
        WX5929) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n3727), .CLK(n4599), .Q(
        WX5931) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n3727), .CLK(n4599), .Q(
        WX5933), .QN(n3669) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n3726), .CLK(n4600), .Q(
        WX5935) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n3726), .CLK(n4600), .Q(
        test_so49) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n3725), .CLK(n4600), 
        .Q(WX5939) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n3724), .CLK(n4601), .Q(
        WX5941), .QN(n3661) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n3723), .CLK(n4601), .Q(
        WX5943) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n3723), .CLK(n4601), .Q(
        WX5945) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n3722), .CLK(n4602), .Q(
        WX5947) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n3722), .CLK(n4602), .Q(
        WX5949) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n3722), .CLK(n4602), .Q(
        WX5951) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n3721), .CLK(n4602), .Q(
        WX5953) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n3721), .CLK(n4602), .Q(
        WX5955) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n3721), .CLK(n4602), .Q(
        WX5957) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n3720), .CLK(n4603), .Q(
        WX5959) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n3720), .CLK(n4603), .Q(
        WX5961) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n3720), .CLK(n4603), .Q(
        WX5963), .QN(n7169) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n3719), .CLK(n4603), .Q(
        WX5965) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n3736), .CLK(n4595), .Q(
        WX5967), .QN(n2959) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n3736), .CLK(n4595), .Q(
        WX5969) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n3736), .CLK(n4595), .Q(
        test_so50) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n3734), .CLK(n4596), 
        .Q(WX5973) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n3734), .CLK(n4596), .Q(
        WX5975) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n3733), .CLK(n4596), .Q(
        WX5977), .QN(n7162) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n3732), .CLK(n4597), .Q(
        WX5979), .QN(n7161) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n3732), .CLK(n4597), .Q(
        WX5981), .QN(n7160) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n3731), .CLK(n4597), .Q(
        WX5983), .QN(n7159) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n3730), .CLK(n4598), .Q(
        WX5985), .QN(n7158) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n3730), .CLK(n4598), .Q(
        WX5987), .QN(n7157) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n3729), .CLK(n4598), .Q(
        WX5989), .QN(n7156) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n3728), .CLK(n4599), .Q(
        WX5991), .QN(n7155) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n3728), .CLK(n4599), .Q(
        WX5993), .QN(n7154) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n3727), .CLK(n4599), .Q(
        WX5995), .QN(n7153) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n3726), .CLK(n4600), .Q(
        WX5997) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n3726), .CLK(n4600), .Q(
        WX5999), .QN(n7152) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n3725), .CLK(n4600), .Q(
        WX6001), .QN(n3118) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n3725), .CLK(n4600), .Q(
        WX6003), .QN(n7151) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n3724), .CLK(n4601), .Q(
        test_so51) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n3723), .CLK(n4601), 
        .Q(WX6007), .QN(n7150) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n3723), .CLK(n4601), .Q(
        WX6009), .QN(n3308) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n3722), .CLK(n4602), .Q(
        WX6011), .QN(n3309) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n3722), .CLK(n4602), .Q(
        WX6013), .QN(n3310) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n3722), .CLK(n4602), .Q(
        WX6015), .QN(n3311) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n3721), .CLK(n4602), .Q(
        WX6017), .QN(n3312) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n3721), .CLK(n4602), .Q(
        WX6019), .QN(n3313) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n3721), .CLK(n4602), .Q(
        WX6021), .QN(n3314) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n3720), .CLK(n4603), .Q(
        WX6023), .QN(n3315) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n3720), .CLK(n4603), .Q(
        WX6025), .QN(n3316) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n3720), .CLK(n4603), .Q(
        WX6027), .QN(n3317) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n3719), .CLK(n4603), .Q(
        WX6029), .QN(n3318) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n3719), .CLK(n4603), .Q(
        WX6031), .QN(n3319) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n3719), .CLK(n4603), .Q(
        WX6033), .QN(n3320) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n3719), .CLK(n4603), .Q(
        WX6035), .QN(n3321) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n3719), .CLK(n4603), .Q(
        WX6037), .QN(n3322) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n3718), .CLK(n4604), .Q(
        test_so52) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n3733), .CLK(n4596), 
        .Q(WX6041), .QN(n3323) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n3732), .CLK(n4597), .Q(
        WX6043), .QN(n3324) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n3732), .CLK(n4597), .Q(
        WX6045), .QN(n3325) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n3731), .CLK(n4597), .Q(
        WX6047), .QN(n3326) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n3730), .CLK(n4598), .Q(
        WX6049), .QN(n3184) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n3730), .CLK(n4598), .Q(
        WX6051), .QN(n3327) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n3729), .CLK(n4598), .Q(
        WX6053), .QN(n3328) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n3728), .CLK(n4599), .Q(
        WX6055), .QN(n3329) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n3728), .CLK(n4599), .Q(
        WX6057), .QN(n3330) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n3727), .CLK(n4599), .Q(
        WX6059), .QN(n3331) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n3726), .CLK(n4600), .Q(
        WX6061), .QN(n3332) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n3726), .CLK(n4600), .Q(
        WX6063), .QN(n3185) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n3725), .CLK(n4600), .Q(
        WX6065), .QN(n3333) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n3724), .CLK(n4601), .Q(
        WX6067), .QN(n3334) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n3724), .CLK(n4601), .Q(
        WX6069), .QN(n3335) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n3723), .CLK(n4601), .Q(
        WX6071), .QN(n3198) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n3682), .CLK(n4620), .Q(
        test_so53) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n3681), .CLK(n4621), 
        .Q(CRC_OUT_5_1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n3681), .CLK(n4621), 
        .Q(CRC_OUT_5_2) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n3681), .CLK(n4621), 
        .Q(CRC_OUT_5_3), .QN(DFF_931_n1) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n3681), .CLK(n4621), 
        .Q(CRC_OUT_5_4) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n3681), .CLK(n4621), 
        .Q(CRC_OUT_5_5) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n3680), .CLK(n4621), 
        .Q(CRC_OUT_5_6) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n3680), .CLK(n4621), 
        .Q(CRC_OUT_5_7) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n3680), .CLK(n4621), 
        .Q(CRC_OUT_5_8) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n3680), .CLK(n4621), 
        .Q(CRC_OUT_5_9) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n3680), .CLK(n4621), 
        .Q(CRC_OUT_5_10), .QN(DFF_938_n1) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n3680), .CLK(n4621), .Q(CRC_OUT_5_11) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n3679), .CLK(n4622), .Q(CRC_OUT_5_12) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n3679), .CLK(n4622), .Q(CRC_OUT_5_13) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n3679), .CLK(n4622), .Q(CRC_OUT_5_14) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n3679), .CLK(n4622), .Q(CRC_OUT_5_15) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n3679), .CLK(n4622), .Q(CRC_OUT_5_16) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n3679), .CLK(n4622), .Q(test_so54) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n3678), .CLK(n4622), 
        .Q(CRC_OUT_5_18) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n3678), .CLK(n4622), .Q(CRC_OUT_5_19) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n3678), .CLK(n4622), .Q(CRC_OUT_5_20) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n3718), .CLK(n4604), .Q(CRC_OUT_5_21) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n3718), .CLK(n4604), .Q(CRC_OUT_5_22) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n3718), .CLK(n4604), .Q(CRC_OUT_5_23) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n3718), .CLK(n4604), .Q(CRC_OUT_5_24) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n3718), .CLK(n4604), .Q(CRC_OUT_5_25) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n3716), .CLK(n4604), .Q(CRC_OUT_5_26) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n3716), .CLK(n4604), .Q(CRC_OUT_5_27) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n3716), .CLK(n4604), .Q(CRC_OUT_5_28) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n3716), .CLK(n4604), .Q(CRC_OUT_5_29) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n3716), .CLK(n4604), .Q(CRC_OUT_5_30) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n3716), .CLK(n4604), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n282), .SI(CRC_OUT_5_31), .SE(n3715), .CLK(n4605), 
        .Q(WX6950), .QN(n3504) );
  SDFFX1 DFF_961_Q_reg ( .D(n283), .SI(WX6950), .SE(n3709), .CLK(n4607), .Q(
        n8470), .QN(n3909) );
  SDFFX1 DFF_962_Q_reg ( .D(n284), .SI(n8470), .SE(n3709), .CLK(n4607), .Q(
        test_so55), .QN(n3908) );
  SDFFX1 DFF_963_Q_reg ( .D(n285), .SI(test_si56), .SE(n3710), .CLK(n4607), 
        .Q(n8467), .QN(n3907) );
  SDFFX1 DFF_964_Q_reg ( .D(n286), .SI(n8467), .SE(n3710), .CLK(n4607), .Q(
        n8466), .QN(n3906) );
  SDFFX1 DFF_965_Q_reg ( .D(n287), .SI(n8466), .SE(n3710), .CLK(n4607), .Q(
        n8465), .QN(n3905) );
  SDFFX1 DFF_966_Q_reg ( .D(n288), .SI(n8465), .SE(n3710), .CLK(n4607), .Q(
        n8464), .QN(n3904) );
  SDFFX1 DFF_967_Q_reg ( .D(n289), .SI(n8464), .SE(n3710), .CLK(n4607), .Q(
        n8463), .QN(n3903) );
  SDFFX1 DFF_968_Q_reg ( .D(n290), .SI(n8463), .SE(n3710), .CLK(n4607), .Q(
        n8462), .QN(n3902) );
  SDFFX1 DFF_969_Q_reg ( .D(n291), .SI(n8462), .SE(n3711), .CLK(n4606), .Q(
        n8461), .QN(n3901) );
  SDFFX1 DFF_970_Q_reg ( .D(n292), .SI(n8461), .SE(n3711), .CLK(n4606), .Q(
        n8460), .QN(n3900) );
  SDFFX1 DFF_971_Q_reg ( .D(n293), .SI(n8460), .SE(n3711), .CLK(n4606), .Q(
        n8459), .QN(n3899) );
  SDFFX1 DFF_972_Q_reg ( .D(n294), .SI(n8459), .SE(n3711), .CLK(n4606), .Q(
        n8458), .QN(n3898) );
  SDFFX1 DFF_973_Q_reg ( .D(n295), .SI(n8458), .SE(n3711), .CLK(n4606), .Q(
        n8457), .QN(n3897) );
  SDFFX1 DFF_974_Q_reg ( .D(n296), .SI(n8457), .SE(n3711), .CLK(n4606), .Q(
        n8456), .QN(n3896) );
  SDFFX1 DFF_975_Q_reg ( .D(n297), .SI(n8456), .SE(n3712), .CLK(n4606), .Q(
        n8455), .QN(n3895) );
  SDFFX1 DFF_976_Q_reg ( .D(n298), .SI(n8455), .SE(n3712), .CLK(n4606), .Q(
        n8454), .QN(n3894) );
  SDFFX1 DFF_977_Q_reg ( .D(n299), .SI(n8454), .SE(n3712), .CLK(n4606), .Q(
        n8453), .QN(n3893) );
  SDFFX1 DFF_978_Q_reg ( .D(n300), .SI(n8453), .SE(n3712), .CLK(n4606), .Q(
        n8452), .QN(n3892) );
  SDFFX1 DFF_979_Q_reg ( .D(n301), .SI(n8452), .SE(n3712), .CLK(n4606), .Q(
        test_so56), .QN(n3891) );
  SDFFX1 DFF_980_Q_reg ( .D(n302), .SI(test_si57), .SE(n3712), .CLK(n4606), 
        .Q(n8449), .QN(n3890) );
  SDFFX1 DFF_981_Q_reg ( .D(n303), .SI(n8449), .SE(n3714), .CLK(n4605), .Q(
        n8448), .QN(n3889) );
  SDFFX1 DFF_982_Q_reg ( .D(n304), .SI(n8448), .SE(n3714), .CLK(n4605), .Q(
        n8447), .QN(n3888) );
  SDFFX1 DFF_983_Q_reg ( .D(n305), .SI(n8447), .SE(n3714), .CLK(n4605), .Q(
        n8446), .QN(n3887) );
  SDFFX1 DFF_984_Q_reg ( .D(n306), .SI(n8446), .SE(n3714), .CLK(n4605), .Q(
        n8445), .QN(n3886) );
  SDFFX1 DFF_985_Q_reg ( .D(WX6999), .SI(n8445), .SE(n3714), .CLK(n4605), .Q(
        n8444), .QN(n3885) );
  SDFFX1 DFF_986_Q_reg ( .D(n308), .SI(n8444), .SE(n3714), .CLK(n4605), .Q(
        n8443) );
  SDFFX1 DFF_987_Q_reg ( .D(n309), .SI(n8443), .SE(n3715), .CLK(n4605), .Q(
        n8442), .QN(n3883) );
  SDFFX1 DFF_988_Q_reg ( .D(n310), .SI(n8442), .SE(n3715), .CLK(n4605), .Q(
        n8441), .QN(n3882) );
  SDFFX1 DFF_989_Q_reg ( .D(n311), .SI(n8441), .SE(n3715), .CLK(n4605), .Q(
        n8440), .QN(n3881) );
  SDFFX1 DFF_990_Q_reg ( .D(n312), .SI(n8440), .SE(n3715), .CLK(n4605), .Q(
        n8439), .QN(n3880) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n3715), .CLK(n4605), .Q(
        n8438), .QN(n3879) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n3682), .CLK(n4620), .Q(
        n8437), .QN(n7149) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n3709), .CLK(n4607), .Q(
        n8436), .QN(n7148) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n3709), .CLK(n4607), .Q(
        n8435), .QN(n7147) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n3708), .CLK(n4608), .Q(
        n8434), .QN(n7146) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n3682), .CLK(n4620), .Q(
        test_so57) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n3708), .CLK(n4608), 
        .Q(n8431), .QN(n7144) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n3708), .CLK(n4608), .Q(
        n8430), .QN(n7143) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n3683), .CLK(n4620), .Q(
        n8429), .QN(n7142) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n3707), .CLK(n4608), .Q(
        n8428), .QN(n7141) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n3706), .CLK(n4609), .Q(
        n8427), .QN(n7140) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n3706), .CLK(n4609), .Q(
        n8426), .QN(n7139) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n3705), .CLK(n4609), .Q(
        n8425), .QN(n7138) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n3705), .CLK(n4609), .Q(
        n8424), .QN(n7137) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n3682), .CLK(n4620), .Q(
        n8423), .QN(n7136) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n4046), .CLK(n4565), .Q(
        n8422), .QN(n7135) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n3703), .CLK(n4610), .Q(
        n8421), .QN(n7134) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n3702), .CLK(n4611), .Q(
        WX7142), .QN(n3115) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n3702), .CLK(n4611), 
        .Q(WX7144), .QN(n3114) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n3701), .CLK(n4611), 
        .Q(WX7146), .QN(n3113) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n3700), .CLK(n4612), 
        .Q(WX7148), .QN(n3112) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n3700), .CLK(n4612), 
        .Q(WX7150), .QN(n3111) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n3699), .CLK(n4612), 
        .Q(test_so58) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n3685), .CLK(n4619), 
        .Q(WX7154), .QN(n3110) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n3697), .CLK(n4613), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n3697), .CLK(n4613), 
        .Q(WX7158), .QN(n3108) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n3697), .CLK(n4613), 
        .Q(WX7160) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n3696), .CLK(n4614), 
        .Q(WX7162), .QN(n3107) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n3695), .CLK(n4614), 
        .Q(WX7164) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n3695), .CLK(n4614), 
        .Q(WX7166), .QN(n3105) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n3694), .CLK(n4615), 
        .Q(WX7168), .QN(n3104) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n3693), .CLK(n4615), 
        .Q(WX7170), .QN(n3103) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n3693), .CLK(n4615), 
        .Q(WX7172), .QN(n3102) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n3692), .CLK(n4616), 
        .Q(WX7174), .QN(n2837) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n3709), .CLK(n4607), 
        .Q(WX7176), .QN(n2951) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n3709), .CLK(n4607), 
        .Q(WX7178), .QN(n2949) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n3708), .CLK(n4608), 
        .Q(WX7180), .QN(n2947) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n3708), .CLK(n4608), 
        .Q(WX7182), .QN(n2946) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n3708), .CLK(n4608), 
        .Q(WX7184), .QN(n2944) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n3707), .CLK(n4608), 
        .Q(test_so59) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n3682), .CLK(n4620), 
        .Q(WX7188), .QN(n2941) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n3707), .CLK(n4608), 
        .Q(WX7190), .QN(n2940) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n3706), .CLK(n4609), 
        .Q(WX7192), .QN(n2938) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n3706), .CLK(n4609), 
        .Q(WX7194), .QN(n2937) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n3705), .CLK(n4609), 
        .Q(WX7196), .QN(n2935) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n3705), .CLK(n4609), 
        .Q(WX7198), .QN(n2933) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n3704), .CLK(n4610), 
        .Q(WX7200), .QN(n2931) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n3704), .CLK(n4610), 
        .Q(WX7202), .QN(n2929) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n3703), .CLK(n4610), 
        .Q(WX7204), .QN(n2927) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n3702), .CLK(n4611), 
        .Q(WX7206) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n3702), .CLK(n4611), 
        .Q(WX7208) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n3701), .CLK(n4611), 
        .Q(WX7210) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n3700), .CLK(n4612), 
        .Q(WX7212) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n3700), .CLK(n4612), 
        .Q(WX7214) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n3699), .CLK(n4612), 
        .Q(WX7216), .QN(n3647) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n3698), .CLK(n4613), 
        .Q(WX7218) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n3698), .CLK(n4613), 
        .Q(test_so60) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n3697), .CLK(n4613), 
        .Q(WX7222) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n3696), .CLK(n4614), 
        .Q(WX7224), .QN(n3639) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n3696), .CLK(n4614), 
        .Q(WX7226) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n3695), .CLK(n4614), 
        .Q(WX7228), .QN(n3635) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n3694), .CLK(n4615), 
        .Q(WX7230) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n3694), .CLK(n4615), 
        .Q(WX7232) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n3693), .CLK(n4615), 
        .Q(WX7234) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n3692), .CLK(n4616), 
        .Q(WX7236) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n3692), .CLK(n4616), 
        .Q(WX7238) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n3690), .CLK(n4616), 
        .Q(WX7240) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n3690), .CLK(n4616), 
        .Q(WX7242) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n3690), .CLK(n4616), 
        .Q(WX7244) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n3689), .CLK(n4617), 
        .Q(WX7246), .QN(n7145) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n3689), .CLK(n4617), 
        .Q(WX7248) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n3707), .CLK(n4608), 
        .Q(WX7250), .QN(n2943) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n3707), .CLK(n4608), 
        .Q(WX7252) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n3707), .CLK(n4608), 
        .Q(test_so61) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n3706), .CLK(n4609), 
        .Q(WX7256) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n3706), .CLK(n4609), 
        .Q(WX7258) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n3705), .CLK(n4609), 
        .Q(WX7260) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n3704), .CLK(n4610), 
        .Q(WX7262) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n3704), .CLK(n4610), 
        .Q(WX7264) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n3703), .CLK(n4610), 
        .Q(WX7266) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n3703), .CLK(n4610), 
        .Q(WX7268) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n3702), .CLK(n4611), 
        .Q(WX7270), .QN(n7133) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n3701), .CLK(n4611), 
        .Q(WX7272), .QN(n7132) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n3701), .CLK(n4611), 
        .Q(WX7274), .QN(n7131) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n3700), .CLK(n4612), 
        .Q(WX7276), .QN(n7130) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n3699), .CLK(n4612), 
        .Q(WX7278), .QN(n7129) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n3699), .CLK(n4612), 
        .Q(WX7280) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n3698), .CLK(n4613), 
        .Q(WX7282), .QN(n7128) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n3698), .CLK(n4613), 
        .Q(WX7284), .QN(n3109) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n3697), .CLK(n4613), 
        .Q(WX7286), .QN(n7127) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n3696), .CLK(n4614), 
        .Q(test_so62) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n3696), .CLK(n4614), 
        .Q(WX7290), .QN(n7126) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n3695), .CLK(n4614), 
        .Q(WX7292), .QN(n3106) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n3694), .CLK(n4615), 
        .Q(WX7294), .QN(n7125) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n3694), .CLK(n4615), 
        .Q(WX7296), .QN(n7124) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n3693), .CLK(n4615), 
        .Q(WX7298), .QN(n7123) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n3692), .CLK(n4616), 
        .Q(WX7300), .QN(n7122) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n3692), .CLK(n4616), 
        .Q(WX7302), .QN(n3281) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n3690), .CLK(n4616), 
        .Q(WX7304), .QN(n3282) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n3690), .CLK(n4616), 
        .Q(WX7306), .QN(n3283) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n3690), .CLK(n4616), 
        .Q(WX7308), .QN(n3284) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n3689), .CLK(n4617), 
        .Q(WX7310), .QN(n3285) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n3689), .CLK(n4617), 
        .Q(WX7312), .QN(n3286) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n3689), .CLK(n4617), 
        .Q(WX7314), .QN(n3287) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n3689), .CLK(n4617), 
        .Q(WX7316), .QN(n3288) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n3688), .CLK(n4617), 
        .Q(WX7318), .QN(n3289) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n3688), .CLK(n4617), 
        .Q(WX7320), .QN(n3290) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n3688), .CLK(n4617), 
        .Q(test_so63) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n3705), .CLK(n4609), 
        .Q(WX7324), .QN(n3291) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n3704), .CLK(n4610), 
        .Q(WX7326), .QN(n3292) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n3704), .CLK(n4610), 
        .Q(WX7328), .QN(n3293) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n3703), .CLK(n4610), 
        .Q(WX7330), .QN(n3294) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n3703), .CLK(n4610), 
        .Q(WX7332), .QN(n3182) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n3702), .CLK(n4611), 
        .Q(WX7334), .QN(n3295) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n3701), .CLK(n4611), 
        .Q(WX7336), .QN(n3296) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n3701), .CLK(n4611), 
        .Q(WX7338), .QN(n3297) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n3700), .CLK(n4612), 
        .Q(WX7340), .QN(n3298) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n3699), .CLK(n4612), 
        .Q(WX7342), .QN(n3183) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n3699), .CLK(n4612), 
        .Q(WX7344), .QN(n3299) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n3698), .CLK(n4613), 
        .Q(WX7346), .QN(n3300) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n3698), .CLK(n4613), 
        .Q(WX7348), .QN(n3301) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n3697), .CLK(n4613), 
        .Q(WX7350), .QN(n3302) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n3696), .CLK(n4614), 
        .Q(WX7352), .QN(n3303) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n3695), .CLK(n4614), 
        .Q(WX7354), .QN(n3304) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n3695), .CLK(n4614), 
        .Q(test_so64) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n3694), .CLK(n4615), 
        .Q(WX7358), .QN(n3305) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n3693), .CLK(n4615), 
        .Q(WX7360), .QN(n3306) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n3693), .CLK(n4615), 
        .Q(WX7362), .QN(n3307) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n3692), .CLK(n4616), 
        .Q(WX7364), .QN(n3197) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n3687), .CLK(n4618), 
        .Q(CRC_OUT_4_0) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n3687), .CLK(n4618), .Q(CRC_OUT_4_1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n3687), .CLK(n4618), .Q(CRC_OUT_4_2) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n3686), .CLK(n4618), .Q(CRC_OUT_4_3) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n3686), .CLK(n4618), .Q(CRC_OUT_4_4) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n3686), .CLK(n4618), .Q(CRC_OUT_4_5) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n3686), .CLK(n4618), .Q(CRC_OUT_4_6) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n3686), .CLK(n4618), .Q(CRC_OUT_4_7) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n3686), .CLK(n4618), .Q(CRC_OUT_4_8) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n3685), .CLK(n4619), .Q(CRC_OUT_4_9) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n3685), .CLK(n4619), .Q(CRC_OUT_4_10), .QN(DFF_1130_n1) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n3685), .CLK(
        n4619), .Q(CRC_OUT_4_11) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n3685), .CLK(
        n4619), .Q(test_so65) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n3685), .CLK(n4619), 
        .Q(CRC_OUT_4_13) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n3684), .CLK(
        n4619), .Q(CRC_OUT_4_14) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n3684), .CLK(
        n4619), .Q(CRC_OUT_4_15), .QN(DFF_1135_n1) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n3684), .CLK(
        n4619), .Q(CRC_OUT_4_16) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n3684), .CLK(
        n4619), .Q(CRC_OUT_4_17) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n3684), .CLK(
        n4619), .Q(CRC_OUT_4_18) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n3684), .CLK(
        n4619), .Q(CRC_OUT_4_19) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n3683), .CLK(
        n4620), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n3683), .CLK(
        n4620), .Q(CRC_OUT_4_21) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n3683), .CLK(
        n4620), .Q(CRC_OUT_4_22) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n3683), .CLK(
        n4620), .Q(CRC_OUT_4_23) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n3683), .CLK(
        n4620), .Q(CRC_OUT_4_24) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n3682), .CLK(
        n4620), .Q(CRC_OUT_4_25) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n3688), .CLK(
        n4617), .Q(CRC_OUT_4_26) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n3688), .CLK(
        n4617), .Q(CRC_OUT_4_27) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n3688), .CLK(
        n4617), .Q(CRC_OUT_4_28) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n3687), .CLK(
        n4618), .Q(test_so66) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n3687), .CLK(n4618), 
        .Q(CRC_OUT_4_30) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n3687), .CLK(
        n4618), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n344), .SI(CRC_OUT_4_31), .SE(n4140), .CLK(n4518), 
        .Q(WX8243), .QN(n3506) );
  SDFFX1 DFF_1153_Q_reg ( .D(n345), .SI(WX8243), .SE(n4140), .CLK(n4518), .Q(
        n8411), .QN(n3878) );
  SDFFX1 DFF_1154_Q_reg ( .D(n346), .SI(n8411), .SE(n4140), .CLK(n4518), .Q(
        n8410), .QN(n3877) );
  SDFFX1 DFF_1155_Q_reg ( .D(n347), .SI(n8410), .SE(n4140), .CLK(n4518), .Q(
        n8409), .QN(n3876) );
  SDFFX1 DFF_1156_Q_reg ( .D(n348), .SI(n8409), .SE(n4141), .CLK(n4518), .Q(
        n8408), .QN(n3875) );
  SDFFX1 DFF_1157_Q_reg ( .D(n349), .SI(n8408), .SE(n4141), .CLK(n4518), .Q(
        n8407), .QN(n3874) );
  SDFFX1 DFF_1158_Q_reg ( .D(n350), .SI(n8407), .SE(n4141), .CLK(n4518), .Q(
        n8406), .QN(n3873) );
  SDFFX1 DFF_1159_Q_reg ( .D(n351), .SI(n8406), .SE(n4141), .CLK(n4518), .Q(
        n8405), .QN(n3872) );
  SDFFX1 DFF_1160_Q_reg ( .D(n352), .SI(n8405), .SE(n4141), .CLK(n4518), .Q(
        n8404), .QN(n3871) );
  SDFFX1 DFF_1161_Q_reg ( .D(n353), .SI(n8404), .SE(n4141), .CLK(n4518), .Q(
        n8403), .QN(n3870) );
  SDFFX1 DFF_1162_Q_reg ( .D(n354), .SI(n8403), .SE(n4142), .CLK(n4517), .Q(
        n8402), .QN(n3869) );
  SDFFX1 DFF_1163_Q_reg ( .D(n355), .SI(n8402), .SE(n4142), .CLK(n4517), .Q(
        n8401), .QN(n3868) );
  SDFFX1 DFF_1164_Q_reg ( .D(WX8266), .SI(n8401), .SE(n4142), .CLK(n4517), .Q(
        n8400), .QN(n3867) );
  SDFFX1 DFF_1165_Q_reg ( .D(n357), .SI(n8400), .SE(n3668), .CLK(n4627), .Q(
        n8399) );
  SDFFX1 DFF_1166_Q_reg ( .D(n358), .SI(n8399), .SE(n4137), .CLK(n4520), .Q(
        test_so67), .QN(n3865) );
  SDFFX1 DFF_1167_Q_reg ( .D(n359), .SI(test_si68), .SE(n4137), .CLK(n4520), 
        .Q(n8396), .QN(n3864) );
  SDFFX1 DFF_1168_Q_reg ( .D(n360), .SI(n8396), .SE(n4137), .CLK(n4520), .Q(
        n8395), .QN(n3863) );
  SDFFX1 DFF_1169_Q_reg ( .D(n361), .SI(n8395), .SE(n4137), .CLK(n4520), .Q(
        n8394), .QN(n3862) );
  SDFFX1 DFF_1170_Q_reg ( .D(n362), .SI(n8394), .SE(n4138), .CLK(n4519), .Q(
        n8393), .QN(n3861) );
  SDFFX1 DFF_1171_Q_reg ( .D(n363), .SI(n8393), .SE(n4138), .CLK(n4519), .Q(
        n8392), .QN(n3860) );
  SDFFX1 DFF_1172_Q_reg ( .D(n364), .SI(n8392), .SE(n4138), .CLK(n4519), .Q(
        n8391), .QN(n3859) );
  SDFFX1 DFF_1173_Q_reg ( .D(n365), .SI(n8391), .SE(n4138), .CLK(n4519), .Q(
        n8390), .QN(n3858) );
  SDFFX1 DFF_1174_Q_reg ( .D(n366), .SI(n8390), .SE(n4138), .CLK(n4519), .Q(
        n8389), .QN(n3857) );
  SDFFX1 DFF_1175_Q_reg ( .D(n367), .SI(n8389), .SE(n4138), .CLK(n4519), .Q(
        n8388), .QN(n3856) );
  SDFFX1 DFF_1176_Q_reg ( .D(n368), .SI(n8388), .SE(n4139), .CLK(n4519), .Q(
        n8387), .QN(n3855) );
  SDFFX1 DFF_1177_Q_reg ( .D(n369), .SI(n8387), .SE(n4139), .CLK(n4519), .Q(
        n8386), .QN(n3854) );
  SDFFX1 DFF_1178_Q_reg ( .D(n370), .SI(n8386), .SE(n4139), .CLK(n4519), .Q(
        n8385), .QN(n3853) );
  SDFFX1 DFF_1179_Q_reg ( .D(n371), .SI(n8385), .SE(n4139), .CLK(n4519), .Q(
        n8384), .QN(n3852) );
  SDFFX1 DFF_1180_Q_reg ( .D(n372), .SI(n8384), .SE(n4139), .CLK(n4519), .Q(
        n8383), .QN(n3851) );
  SDFFX1 DFF_1181_Q_reg ( .D(n373), .SI(n8383), .SE(n4139), .CLK(n4519), .Q(
        n8382), .QN(n3850) );
  SDFFX1 DFF_1182_Q_reg ( .D(n374), .SI(n8382), .SE(n4140), .CLK(n4518), .Q(
        n8381), .QN(n3849) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n4140), .CLK(n4518), .Q(
        test_so68), .QN(n3848) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n4127), .CLK(n4525), 
        .Q(n8378), .QN(n7121) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n4127), .CLK(n4525), .Q(
        n8377), .QN(n7120) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n4107), .CLK(n4535), .Q(
        n8376), .QN(n7119) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n4126), .CLK(n4525), .Q(
        n8375), .QN(n7118) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n4125), .CLK(n4526), .Q(
        n8374), .QN(n7117) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n4125), .CLK(n4526), .Q(
        n8373), .QN(n7116) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n4123), .CLK(n4527), .Q(
        n8372), .QN(n7115) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n4123), .CLK(n4527), .Q(
        n8371), .QN(n7114) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n4122), .CLK(n4527), .Q(
        n8370), .QN(n7113) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n4122), .CLK(n4527), .Q(
        n8369), .QN(n7112) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n4121), .CLK(n4528), .Q(
        n8368), .QN(n7111) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n4121), .CLK(n4528), .Q(
        n8367), .QN(n7110) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n4119), .CLK(n4529), .Q(
        n8366), .QN(n7109) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n4119), .CLK(n4529), .Q(
        n8365), .QN(n7108) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n4137), .CLK(n4520), .Q(
        n8364), .QN(n7107) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n4136), .CLK(n4520), .Q(
        n8363), .QN(n7106) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n4136), .CLK(n4520), .Q(
        test_so69) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n4046), .CLK(n4565), 
        .Q(WX8437), .QN(n3101) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n4135), .CLK(n4521), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n4135), .CLK(n4521), 
        .Q(WX8441), .QN(n3099) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n4135), .CLK(n4521), 
        .Q(WX8443) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n4135), .CLK(n4521), 
        .Q(WX8445), .QN(n3098) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n4134), .CLK(n4521), 
        .Q(WX8447) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n4134), .CLK(n4521), 
        .Q(WX8449), .QN(n3096) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n4133), .CLK(n4522), 
        .Q(WX8451), .QN(n3095) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n4132), .CLK(n4522), 
        .Q(WX8453), .QN(n3094) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n4132), .CLK(n4522), 
        .Q(WX8455), .QN(n3093) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n4131), .CLK(n4523), 
        .Q(WX8457), .QN(n3092) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n4130), .CLK(n4523), 
        .Q(WX8459), .QN(n3091) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n4130), .CLK(n4523), 
        .Q(WX8461), .QN(n3090) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n4129), .CLK(n4524), 
        .Q(WX8463), .QN(n3089) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n4128), .CLK(n4524), 
        .Q(WX8465), .QN(n3088) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n4128), .CLK(n4524), 
        .Q(WX8467), .QN(n2835) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n4127), .CLK(n4525), 
        .Q(test_so70) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n4106), .CLK(n4535), 
        .Q(WX8471), .QN(n2924) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n4125), .CLK(n4526), 
        .Q(WX8473), .QN(n2923) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n4125), .CLK(n4526), 
        .Q(WX8475), .QN(n2921) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n4124), .CLK(n4526), 
        .Q(WX8477), .QN(n2920) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n4124), .CLK(n4526), 
        .Q(WX8479), .QN(n2918) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n4123), .CLK(n4527), 
        .Q(WX8481), .QN(n2916) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n4123), .CLK(n4527), 
        .Q(WX8483), .QN(n2914) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n4122), .CLK(n4527), 
        .Q(WX8485), .QN(n2912) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n4121), .CLK(n4528), 
        .Q(WX8487), .QN(n2910) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n4120), .CLK(n4528), 
        .Q(WX8489), .QN(n2908) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n4120), .CLK(n4528), 
        .Q(WX8491), .QN(n2906) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n4119), .CLK(n4529), 
        .Q(WX8493), .QN(n2904) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n4137), .CLK(n4520), 
        .Q(WX8495), .QN(n2902) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n4136), .CLK(n4520), 
        .Q(WX8497), .QN(n2900) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n4136), .CLK(n4520), 
        .Q(WX8499), .QN(n3625) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n4136), .CLK(n4520), 
        .Q(WX8501) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n4136), .CLK(n4520), 
        .Q(test_so71) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n4135), .CLK(n4521), 
        .Q(WX8505) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n4135), .CLK(n4521), 
        .Q(WX8507), .QN(n3617) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n4134), .CLK(n4521), 
        .Q(WX8509) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n4134), .CLK(n4521), 
        .Q(WX8511), .QN(n3613) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n4133), .CLK(n4522), 
        .Q(WX8513) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n4133), .CLK(n4522), 
        .Q(WX8515) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n4132), .CLK(n4522), 
        .Q(WX8517) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n4131), .CLK(n4523), 
        .Q(WX8519) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n4131), .CLK(n4523), 
        .Q(WX8521) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n4130), .CLK(n4523), 
        .Q(WX8523) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n4129), .CLK(n4524), 
        .Q(WX8525) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n4129), .CLK(n4524), 
        .Q(WX8527) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n4128), .CLK(n4524), 
        .Q(WX8529) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n4127), .CLK(n4525), 
        .Q(WX8531) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n4127), .CLK(n4525), 
        .Q(WX8533), .QN(n2926) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n4126), .CLK(n4525), 
        .Q(WX8535) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n4126), .CLK(n4525), 
        .Q(test_so72) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n4125), .CLK(n4526), 
        .Q(WX8539) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n4124), .CLK(n4526), 
        .Q(WX8541) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n4124), .CLK(n4526), 
        .Q(WX8543) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n4123), .CLK(n4527), 
        .Q(WX8545) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n4122), .CLK(n4527), 
        .Q(WX8547) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n4122), .CLK(n4527), 
        .Q(WX8549) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n4121), .CLK(n4528), 
        .Q(WX8551) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n4120), .CLK(n4528), 
        .Q(WX8553) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n4120), .CLK(n4528), 
        .Q(WX8555) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n4119), .CLK(n4529), 
        .Q(WX8557) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n4119), .CLK(n4529), 
        .Q(WX8559) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n4118), .CLK(n4529), 
        .Q(WX8561) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n4118), .CLK(n4529), 
        .Q(WX8563) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n4118), .CLK(n4529), 
        .Q(WX8565), .QN(n7105) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n4117), .CLK(n4530), 
        .Q(WX8567), .QN(n3100) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n4117), .CLK(n4530), 
        .Q(WX8569), .QN(n7104) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n4117), .CLK(n4530), 
        .Q(test_so73) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n4134), .CLK(n4521), 
        .Q(WX8573), .QN(n7103) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n4134), .CLK(n4521), 
        .Q(WX8575), .QN(n3097) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n4133), .CLK(n4522), 
        .Q(WX8577), .QN(n7102) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n4133), .CLK(n4522), 
        .Q(WX8579), .QN(n7101) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n4132), .CLK(n4522), 
        .Q(WX8581), .QN(n7100) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n4131), .CLK(n4523), 
        .Q(WX8583), .QN(n7099) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n4131), .CLK(n4523), 
        .Q(WX8585), .QN(n7098) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n4130), .CLK(n4523), 
        .Q(WX8587), .QN(n7097) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n4129), .CLK(n4524), 
        .Q(WX8589), .QN(n7096) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n4129), .CLK(n4524), 
        .Q(WX8591), .QN(n7095) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n4128), .CLK(n4524), 
        .Q(WX8593), .QN(n7094) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n4127), .CLK(n4525), 
        .Q(WX8595), .QN(n3254) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n4126), .CLK(n4525), 
        .Q(WX8597), .QN(n3255) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n4126), .CLK(n4525), 
        .Q(WX8599), .QN(n3256) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n4126), .CLK(n4525), 
        .Q(WX8601), .QN(n3257) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n4125), .CLK(n4526), 
        .Q(WX8603), .QN(n3258) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n4124), .CLK(n4526), 
        .Q(test_so74) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n4124), .CLK(n4526), 
        .Q(WX8607), .QN(n3259) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n4123), .CLK(n4527), 
        .Q(WX8609), .QN(n3260) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n4122), .CLK(n4527), 
        .Q(WX8611), .QN(n3261) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n4121), .CLK(n4528), 
        .Q(WX8613), .QN(n3262) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n4121), .CLK(n4528), 
        .Q(WX8615), .QN(n3263) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n4120), .CLK(n4528), 
        .Q(WX8617), .QN(n3264) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n4120), .CLK(n4528), 
        .Q(WX8619), .QN(n3265) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n4119), .CLK(n4529), 
        .Q(WX8621), .QN(n3266) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n4118), .CLK(n4529), 
        .Q(WX8623), .QN(n3267) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n4118), .CLK(n4529), 
        .Q(WX8625), .QN(n3179) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n4118), .CLK(n4529), 
        .Q(WX8627), .QN(n3268) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n4117), .CLK(n4530), 
        .Q(WX8629), .QN(n3269) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n4117), .CLK(n4530), 
        .Q(WX8631), .QN(n3270) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n4117), .CLK(n4530), 
        .Q(WX8633), .QN(n3271) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n4116), .CLK(n4530), 
        .Q(WX8635), .QN(n3180) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n4116), .CLK(n4530), 
        .Q(WX8637), .QN(n3272) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n4116), .CLK(n4530), 
        .Q(test_so75) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n4133), .CLK(n4522), 
        .Q(WX8641), .QN(n3273) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n4132), .CLK(n4522), 
        .Q(WX8643), .QN(n3274) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n4132), .CLK(n4522), 
        .Q(WX8645), .QN(n3275) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n4131), .CLK(n4523), 
        .Q(WX8647), .QN(n3276) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n4130), .CLK(n4523), 
        .Q(WX8649), .QN(n3181) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n4130), .CLK(n4523), 
        .Q(WX8651), .QN(n3277) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n4129), .CLK(n4524), 
        .Q(WX8653), .QN(n3279) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n4128), .CLK(n4524), 
        .Q(WX8655), .QN(n3280) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n4128), .CLK(n4524), 
        .Q(WX8657), .QN(n3196) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n4048), .CLK(n4564), 
        .Q(CRC_OUT_3_0) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n4048), .CLK(n4564), .Q(CRC_OUT_3_1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n4048), .CLK(n4564), .Q(CRC_OUT_3_2) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n4048), .CLK(n4564), .Q(CRC_OUT_3_3), .QN(DFF_1315_n1) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n4047), .CLK(n4565), .Q(CRC_OUT_3_4) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n4047), .CLK(n4565), .Q(CRC_OUT_3_5) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n4047), .CLK(n4565), .Q(CRC_OUT_3_6) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n4047), .CLK(n4565), .Q(test_so76) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n4047), .CLK(n4565), 
        .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n4047), .CLK(n4565), .Q(CRC_OUT_3_9) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n4046), .CLK(n4565), .Q(CRC_OUT_3_10), .QN(DFF_1322_n1) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n4116), .CLK(
        n4530), .Q(CRC_OUT_3_11) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n4116), .CLK(
        n4530), .Q(CRC_OUT_3_12) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n4116), .CLK(
        n4530), .Q(CRC_OUT_3_13) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n4115), .CLK(
        n4531), .Q(CRC_OUT_3_14) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n4115), .CLK(
        n4531), .Q(CRC_OUT_3_15), .QN(DFF_1327_n1) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n4115), .CLK(
        n4531), .Q(CRC_OUT_3_16) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n4115), .CLK(
        n4531), .Q(CRC_OUT_3_17) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n4115), .CLK(
        n4531), .Q(CRC_OUT_3_18) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n4115), .CLK(
        n4531), .Q(CRC_OUT_3_19) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n4114), .CLK(
        n4531), .Q(CRC_OUT_3_20) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n4114), .CLK(
        n4531), .Q(CRC_OUT_3_21) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n4114), .CLK(
        n4531), .Q(CRC_OUT_3_22) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n4114), .CLK(
        n4531), .Q(CRC_OUT_3_23) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n4114), .CLK(
        n4531), .Q(test_so77) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n4114), .CLK(n4531), 
        .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n4113), .CLK(
        n4532), .Q(CRC_OUT_3_26) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n4113), .CLK(
        n4532), .Q(CRC_OUT_3_27) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n4113), .CLK(
        n4532), .Q(CRC_OUT_3_28) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n4113), .CLK(
        n4532), .Q(CRC_OUT_3_29) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n4113), .CLK(
        n4532), .Q(CRC_OUT_3_30) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n4113), .CLK(
        n4532), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n406), .SI(CRC_OUT_3_31), .SE(n4112), .CLK(n4532), 
        .Q(WX9536), .QN(n3508) );
  SDFFX1 DFF_1345_Q_reg ( .D(n407), .SI(WX9536), .SE(n4107), .CLK(n4535), .Q(
        n8353), .QN(n3847) );
  SDFFX1 DFF_1346_Q_reg ( .D(n408), .SI(n8353), .SE(n4107), .CLK(n4535), .Q(
        n8352), .QN(n3846) );
  SDFFX1 DFF_1347_Q_reg ( .D(n409), .SI(n8352), .SE(n4108), .CLK(n4534), .Q(
        n8351), .QN(n3845) );
  SDFFX1 DFF_1348_Q_reg ( .D(n410), .SI(n8351), .SE(n4108), .CLK(n4534), .Q(
        n8350), .QN(n3844) );
  SDFFX1 DFF_1349_Q_reg ( .D(n411), .SI(n8350), .SE(n4108), .CLK(n4534), .Q(
        n8349), .QN(n3843) );
  SDFFX1 DFF_1350_Q_reg ( .D(n412), .SI(n8349), .SE(n4108), .CLK(n4534), .Q(
        n8348), .QN(n3842) );
  SDFFX1 DFF_1351_Q_reg ( .D(n413), .SI(n8348), .SE(n4108), .CLK(n4534), .Q(
        n8347), .QN(n3841) );
  SDFFX1 DFF_1352_Q_reg ( .D(n414), .SI(n8347), .SE(n4108), .CLK(n4534), .Q(
        n8346), .QN(n3840) );
  SDFFX1 DFF_1353_Q_reg ( .D(n415), .SI(n8346), .SE(n4109), .CLK(n4534), .Q(
        test_so78), .QN(n3839) );
  SDFFX1 DFF_1354_Q_reg ( .D(n416), .SI(test_si79), .SE(n4109), .CLK(n4534), 
        .Q(n8343), .QN(n3838) );
  SDFFX1 DFF_1355_Q_reg ( .D(n417), .SI(n8343), .SE(n4109), .CLK(n4534), .Q(
        n8342), .QN(n3837) );
  SDFFX1 DFF_1356_Q_reg ( .D(n418), .SI(n8342), .SE(n4109), .CLK(n4534), .Q(
        n8341), .QN(n3836) );
  SDFFX1 DFF_1357_Q_reg ( .D(n419), .SI(n8341), .SE(n4109), .CLK(n4534), .Q(
        n8340), .QN(n3835) );
  SDFFX1 DFF_1358_Q_reg ( .D(n420), .SI(n8340), .SE(n4109), .CLK(n4534), .Q(
        n8339), .QN(n3834) );
  SDFFX1 DFF_1359_Q_reg ( .D(n421), .SI(n8339), .SE(n4110), .CLK(n4533), .Q(
        n8338), .QN(n3833) );
  SDFFX1 DFF_1360_Q_reg ( .D(n422), .SI(n8338), .SE(n4110), .CLK(n4533), .Q(
        n8337), .QN(n3832) );
  SDFFX1 DFF_1361_Q_reg ( .D(n423), .SI(n8337), .SE(n4110), .CLK(n4533), .Q(
        n8336), .QN(n3831) );
  SDFFX1 DFF_1362_Q_reg ( .D(n424), .SI(n8336), .SE(n4110), .CLK(n4533), .Q(
        n8335), .QN(n3830) );
  SDFFX1 DFF_1363_Q_reg ( .D(n425), .SI(n8335), .SE(n4110), .CLK(n4533), .Q(
        n8334), .QN(n3829) );
  SDFFX1 DFF_1364_Q_reg ( .D(n426), .SI(n8334), .SE(n4110), .CLK(n4533), .Q(
        n8333), .QN(n3828) );
  SDFFX1 DFF_1365_Q_reg ( .D(n427), .SI(n8333), .SE(n4111), .CLK(n4533), .Q(
        n8332), .QN(n3827) );
  SDFFX1 DFF_1366_Q_reg ( .D(n428), .SI(n8332), .SE(n4111), .CLK(n4533), .Q(
        n8331), .QN(n3826) );
  SDFFX1 DFF_1367_Q_reg ( .D(n429), .SI(n8331), .SE(n4111), .CLK(n4533), .Q(
        n8330), .QN(n3825) );
  SDFFX1 DFF_1368_Q_reg ( .D(n430), .SI(n8330), .SE(n4111), .CLK(n4533), .Q(
        n8329), .QN(n3824) );
  SDFFX1 DFF_1369_Q_reg ( .D(n431), .SI(n8329), .SE(n4111), .CLK(n4533), .Q(
        n8328), .QN(n3823) );
  SDFFX1 DFF_1370_Q_reg ( .D(n432), .SI(n8328), .SE(n4111), .CLK(n4533), .Q(
        test_so79), .QN(n3822) );
  SDFFX1 DFF_1371_Q_reg ( .D(n433), .SI(test_si80), .SE(n4112), .CLK(n4532), 
        .Q(n8325), .QN(n3821) );
  SDFFX1 DFF_1372_Q_reg ( .D(n434), .SI(n8325), .SE(n4112), .CLK(n4532), .Q(
        n8324), .QN(n3820) );
  SDFFX1 DFF_1373_Q_reg ( .D(n435), .SI(n8324), .SE(n4112), .CLK(n4532), .Q(
        n8323), .QN(n3819) );
  SDFFX1 DFF_1374_Q_reg ( .D(n436), .SI(n8323), .SE(n4112), .CLK(n4532), .Q(
        n8322), .QN(n3818) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n4112), .CLK(n4532), .Q(
        n8321), .QN(n3817) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n4048), .CLK(n4564), .Q(
        n8320), .QN(n7093) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n4107), .CLK(n4535), .Q(
        n8319), .QN(n7092) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n4106), .CLK(n4535), .Q(
        n8318), .QN(n7091) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n4106), .CLK(n4535), .Q(
        n8317), .QN(n7090) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n4106), .CLK(n4535), .Q(
        n8316), .QN(n7089) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n4105), .CLK(n4536), .Q(
        n8315), .QN(n7088) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n4105), .CLK(n4536), .Q(
        n8314), .QN(n7087) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n4105), .CLK(n4536), .Q(
        n8313), .QN(n7086) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n4104), .CLK(n4536), .Q(
        n8312), .QN(n7085) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n4104), .CLK(n4536), .Q(
        n8311), .QN(n7084) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n4104), .CLK(n4536), .Q(
        n8310), .QN(n7083) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n4103), .CLK(n4537), .Q(
        test_so80) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n4103), .CLK(n4537), 
        .Q(n8307), .QN(n7081) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n4103), .CLK(n4537), .Q(
        n8306), .QN(n7080) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n4049), .CLK(n4564), .Q(
        n8305), .QN(n7079) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n4102), .CLK(n4537), .Q(
        n8304), .QN(n7078) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n4049), .CLK(n4564), .Q(
        WX9728), .QN(n3087) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n4101), .CLK(n4538), 
        .Q(WX9730) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n4101), .CLK(n4538), 
        .Q(WX9732), .QN(n3085) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n4100), .CLK(n4538), 
        .Q(WX9734), .QN(n3084) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n4099), .CLK(n4539), 
        .Q(WX9736), .QN(n3083) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n4099), .CLK(n4539), 
        .Q(WX9738), .QN(n3082) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n4098), .CLK(n4539), 
        .Q(WX9740), .QN(n3081) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n4097), .CLK(n4540), 
        .Q(WX9742), .QN(n3080) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n4097), .CLK(n4540), 
        .Q(WX9744), .QN(n3079) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n4096), .CLK(n4540), 
        .Q(WX9746), .QN(n3078) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n4095), .CLK(n4541), 
        .Q(WX9748), .QN(n3077) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n4095), .CLK(n4541), 
        .Q(WX9750), .QN(n3076) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n4094), .CLK(n4541), 
        .Q(test_so81) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n4052), .CLK(n4562), 
        .Q(WX9754), .QN(n3075) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n4092), .CLK(n4542), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n4092), .CLK(n4542), 
        .Q(WX9758), .QN(n3073) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n4092), .CLK(n4542), 
        .Q(WX9760), .QN(n2834) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n4107), .CLK(n4535), 
        .Q(WX9762), .QN(n2898) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n4107), .CLK(n4535), 
        .Q(WX9764), .QN(n2896) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n4106), .CLK(n4535), 
        .Q(WX9766), .QN(n2894) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n4106), .CLK(n4535), 
        .Q(WX9768), .QN(n2892) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n4105), .CLK(n4536), 
        .Q(WX9770), .QN(n2890) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n4105), .CLK(n4536), 
        .Q(WX9772), .QN(n2888) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n4105), .CLK(n4536), 
        .Q(WX9774), .QN(n2886) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n4104), .CLK(n4536), 
        .Q(WX9776), .QN(n2884) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n4104), .CLK(n4536), 
        .Q(WX9778), .QN(n2882) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n4104), .CLK(n4536), 
        .Q(WX9780), .QN(n2880) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n4103), .CLK(n4537), 
        .Q(WX9782), .QN(n2879) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n4103), .CLK(n4537), 
        .Q(WX9784), .QN(n2877) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n4103), .CLK(n4537), 
        .Q(test_so82) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n4048), .CLK(n4564), 
        .Q(WX9788), .QN(n2874) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n4102), .CLK(n4537), 
        .Q(WX9790), .QN(n2873) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n4102), .CLK(n4537), 
        .Q(WX9792) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n4101), .CLK(n4538), 
        .Q(WX9794), .QN(n3591) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n4101), .CLK(n4538), 
        .Q(WX9796) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n4100), .CLK(n4538), 
        .Q(WX9798) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n4099), .CLK(n4539), 
        .Q(WX9800) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n4099), .CLK(n4539), 
        .Q(WX9802) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n4098), .CLK(n4539), 
        .Q(WX9804) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n4097), .CLK(n4540), 
        .Q(WX9806) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n4097), .CLK(n4540), 
        .Q(WX9808) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n4096), .CLK(n4540), 
        .Q(WX9810) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n4095), .CLK(n4541), 
        .Q(WX9812) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n4095), .CLK(n4541), 
        .Q(WX9814) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n4094), .CLK(n4541), 
        .Q(WX9816), .QN(n3569) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n4093), .CLK(n4542), 
        .Q(WX9818) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n4093), .CLK(n4542), 
        .Q(test_so83) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n4092), .CLK(n4542), 
        .Q(WX9822) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n4091), .CLK(n4543), 
        .Q(WX9824) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n4091), .CLK(n4543), 
        .Q(WX9826) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n4091), .CLK(n4543), 
        .Q(WX9828) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n4090), .CLK(n4543), 
        .Q(WX9830) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n4090), .CLK(n4543), 
        .Q(WX9832) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n4090), .CLK(n4543), 
        .Q(WX9834) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n4089), .CLK(n4544), 
        .Q(WX9836) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n4089), .CLK(n4544), 
        .Q(WX9838) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n4089), .CLK(n4544), 
        .Q(WX9840) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n4088), .CLK(n4544), 
        .Q(WX9842) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n4088), .CLK(n4544), 
        .Q(WX9844) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n4088), .CLK(n4544), 
        .Q(WX9846), .QN(n7082) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n4087), .CLK(n4545), 
        .Q(WX9848) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n4102), .CLK(n4537), 
        .Q(WX9850), .QN(n2876) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n4102), .CLK(n4537), 
        .Q(WX9852) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n4102), .CLK(n4537), 
        .Q(test_so84) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n4101), .CLK(n4538), 
        .Q(WX9856), .QN(n7077) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n4101), .CLK(n4538), 
        .Q(WX9858), .QN(n3086) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n4100), .CLK(n4538), 
        .Q(WX9860), .QN(n7076) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n4100), .CLK(n4538), 
        .Q(WX9862), .QN(n7075) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n4099), .CLK(n4539), 
        .Q(WX9864), .QN(n7074) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n4098), .CLK(n4539), 
        .Q(WX9866), .QN(n7073) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n4098), .CLK(n4539), 
        .Q(WX9868), .QN(n7072) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n4097), .CLK(n4540), 
        .Q(WX9870), .QN(n7071) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n4096), .CLK(n4540), 
        .Q(WX9872), .QN(n7070) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n4096), .CLK(n4540), 
        .Q(WX9874), .QN(n7069) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n4095), .CLK(n4541), 
        .Q(WX9876), .QN(n7068) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n4094), .CLK(n4541), 
        .Q(WX9878), .QN(n7067) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n4094), .CLK(n4541), 
        .Q(WX9880) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n4093), .CLK(n4542), 
        .Q(WX9882), .QN(n7066) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n4093), .CLK(n4542), 
        .Q(WX9884), .QN(n3074) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n4092), .CLK(n4542), 
        .Q(WX9886), .QN(n7065) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n4091), .CLK(n4543), 
        .Q(test_so85) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n4091), .CLK(n4543), 
        .Q(WX9890), .QN(n3228) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n4091), .CLK(n4543), 
        .Q(WX9892), .QN(n3229) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n4090), .CLK(n4543), 
        .Q(WX9894), .QN(n3230) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n4090), .CLK(n4543), 
        .Q(WX9896), .QN(n3231) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n4090), .CLK(n4543), 
        .Q(WX9898), .QN(n3232) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n4089), .CLK(n4544), 
        .Q(WX9900), .QN(n3233) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n4089), .CLK(n4544), 
        .Q(WX9902), .QN(n3234) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n4089), .CLK(n4544), 
        .Q(WX9904), .QN(n3235) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n4088), .CLK(n4544), 
        .Q(WX9906), .QN(n3236) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n4088), .CLK(n4544), 
        .Q(WX9908), .QN(n3237) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n4088), .CLK(n4544), 
        .Q(WX9910), .QN(n3238) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n4087), .CLK(n4545), 
        .Q(WX9912), .QN(n3239) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n4087), .CLK(n4545), 
        .Q(WX9914), .QN(n3240) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n4087), .CLK(n4545), 
        .Q(WX9916), .QN(n3241) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n4087), .CLK(n4545), 
        .Q(WX9918), .QN(n3176) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n4087), .CLK(n4545), 
        .Q(WX9920), .QN(n3242) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n4086), .CLK(n4545), 
        .Q(test_so86) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n4100), .CLK(n4538), 
        .Q(WX9924), .QN(n3243) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n4100), .CLK(n4538), 
        .Q(WX9926), .QN(n3244) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n4099), .CLK(n4539), 
        .Q(WX9928), .QN(n3177) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n4098), .CLK(n4539), 
        .Q(WX9930), .QN(n3245) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n4098), .CLK(n4539), 
        .Q(WX9932), .QN(n3246) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n4097), .CLK(n4540), 
        .Q(WX9934), .QN(n3247) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n4096), .CLK(n4540), 
        .Q(WX9936), .QN(n3248) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n4096), .CLK(n4540), 
        .Q(WX9938), .QN(n3249) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n4095), .CLK(n4541), 
        .Q(WX9940), .QN(n3250) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n4094), .CLK(n4541), 
        .Q(WX9942), .QN(n3178) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n4094), .CLK(n4541), 
        .Q(WX9944), .QN(n3251) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n4093), .CLK(n4542), 
        .Q(WX9946), .QN(n3252) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n4093), .CLK(n4542), 
        .Q(WX9948), .QN(n3253) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n4092), .CLK(n4542), 
        .Q(WX9950), .QN(n3195) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n4052), .CLK(n4562), 
        .Q(CRC_OUT_2_0) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n4052), .CLK(
        n4562), .Q(CRC_OUT_2_1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n4052), .CLK(
        n4562), .Q(test_so87) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n4051), .CLK(n4563), 
        .Q(CRC_OUT_2_3), .QN(DFF_1507_n1) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n4051), .CLK(
        n4563), .Q(CRC_OUT_2_4) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n4051), .CLK(
        n4563), .Q(CRC_OUT_2_5) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n4051), .CLK(
        n4563), .Q(CRC_OUT_2_6) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n4051), .CLK(
        n4563), .Q(CRC_OUT_2_7) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n4051), .CLK(
        n4563), .Q(CRC_OUT_2_8) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n4050), .CLK(
        n4563), .Q(CRC_OUT_2_9) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n4050), .CLK(
        n4563), .Q(CRC_OUT_2_10), .QN(DFF_1514_n1) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n4050), .CLK(
        n4563), .Q(CRC_OUT_2_11) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n4050), .CLK(
        n4563), .Q(CRC_OUT_2_12) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n4050), .CLK(
        n4563), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n4050), .CLK(
        n4563), .Q(CRC_OUT_2_14) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n4049), .CLK(
        n4564), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n4049), .CLK(
        n4564), .Q(CRC_OUT_2_16) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n4049), .CLK(
        n4564), .Q(CRC_OUT_2_17) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n4049), .CLK(
        n4564), .Q(CRC_OUT_2_18) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n4086), .CLK(
        n4545), .Q(test_so88) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n4086), .CLK(n4545), 
        .Q(CRC_OUT_2_20) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n4086), .CLK(
        n4545), .Q(CRC_OUT_2_21) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n4086), .CLK(
        n4545), .Q(CRC_OUT_2_22) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n4086), .CLK(
        n4545), .Q(CRC_OUT_2_23) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n4085), .CLK(
        n4546), .Q(CRC_OUT_2_24) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n4085), .CLK(
        n4546), .Q(CRC_OUT_2_25) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n4085), .CLK(
        n4546), .Q(CRC_OUT_2_26) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n4085), .CLK(
        n4546), .Q(CRC_OUT_2_27) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n4085), .CLK(
        n4546), .Q(CRC_OUT_2_28) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n4085), .CLK(
        n4546), .Q(CRC_OUT_2_29) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n4084), .CLK(
        n4546), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n4084), .CLK(
        n4546), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(n468), .SI(CRC_OUT_2_31), .SE(n4084), .CLK(n4546), 
        .Q(WX10829), .QN(n3510) );
  SDFFX1 DFF_1537_Q_reg ( .D(n469), .SI(WX10829), .SE(n4079), .CLK(n4549), .Q(
        n8295), .QN(n3816) );
  SDFFX1 DFF_1538_Q_reg ( .D(n470), .SI(n8295), .SE(n4079), .CLK(n4549), .Q(
        n8294), .QN(n3815) );
  SDFFX1 DFF_1539_Q_reg ( .D(n471), .SI(n8294), .SE(n4079), .CLK(n4549), .Q(
        n8293), .QN(n3814) );
  SDFFX1 DFF_1540_Q_reg ( .D(n472), .SI(n8293), .SE(n4079), .CLK(n4549), .Q(
        test_so89), .QN(n3813) );
  SDFFX1 DFF_1541_Q_reg ( .D(n473), .SI(test_si90), .SE(n4080), .CLK(n4548), 
        .Q(n8290), .QN(n3812) );
  SDFFX1 DFF_1542_Q_reg ( .D(n474), .SI(n8290), .SE(n4080), .CLK(n4548), .Q(
        n8289), .QN(n3811) );
  SDFFX1 DFF_1543_Q_reg ( .D(n475), .SI(n8289), .SE(n4080), .CLK(n4548), .Q(
        n8288), .QN(n3810) );
  SDFFX1 DFF_1544_Q_reg ( .D(n476), .SI(n8288), .SE(n4080), .CLK(n4548), .Q(
        n8287), .QN(n3809) );
  SDFFX1 DFF_1545_Q_reg ( .D(n477), .SI(n8287), .SE(n4080), .CLK(n4548), .Q(
        n8286), .QN(n3808) );
  SDFFX1 DFF_1546_Q_reg ( .D(n478), .SI(n8286), .SE(n4080), .CLK(n4548), .Q(
        n8285), .QN(n3807) );
  SDFFX1 DFF_1547_Q_reg ( .D(n479), .SI(n8285), .SE(n4081), .CLK(n4548), .Q(
        n8284), .QN(n3806) );
  SDFFX1 DFF_1548_Q_reg ( .D(n480), .SI(n8284), .SE(n4081), .CLK(n4548), .Q(
        n8283), .QN(n3805) );
  SDFFX1 DFF_1549_Q_reg ( .D(n481), .SI(n8283), .SE(n4081), .CLK(n4548), .Q(
        n8282), .QN(n3804) );
  SDFFX1 DFF_1550_Q_reg ( .D(n482), .SI(n8282), .SE(n4081), .CLK(n4548), .Q(
        n8281), .QN(n3803) );
  SDFFX1 DFF_1551_Q_reg ( .D(n483), .SI(n8281), .SE(n4081), .CLK(n4548), .Q(
        n8280), .QN(n3802) );
  SDFFX1 DFF_1552_Q_reg ( .D(n484), .SI(n8280), .SE(n4081), .CLK(n4548), .Q(
        n8279), .QN(n3801) );
  SDFFX1 DFF_1553_Q_reg ( .D(n485), .SI(n8279), .SE(n4082), .CLK(n4547), .Q(
        n8278), .QN(n3800) );
  SDFFX1 DFF_1554_Q_reg ( .D(n486), .SI(n8278), .SE(n4082), .CLK(n4547), .Q(
        n8277), .QN(n3799) );
  SDFFX1 DFF_1555_Q_reg ( .D(n487), .SI(n8277), .SE(n4082), .CLK(n4547), .Q(
        n8276), .QN(n3798) );
  SDFFX1 DFF_1556_Q_reg ( .D(n488), .SI(n8276), .SE(n4082), .CLK(n4547), .Q(
        n8275), .QN(n3797) );
  SDFFX1 DFF_1557_Q_reg ( .D(n489), .SI(n8275), .SE(n4082), .CLK(n4547), .Q(
        test_so90), .QN(n3796) );
  SDFFX1 DFF_1558_Q_reg ( .D(n490), .SI(test_si91), .SE(n4082), .CLK(n4547), 
        .Q(n8272), .QN(n3795) );
  SDFFX1 DFF_1559_Q_reg ( .D(n491), .SI(n8272), .SE(n4083), .CLK(n4547), .Q(
        n8271), .QN(n3794) );
  SDFFX1 DFF_1560_Q_reg ( .D(n492), .SI(n8271), .SE(n4083), .CLK(n4547), .Q(
        n8270), .QN(n3793) );
  SDFFX1 DFF_1561_Q_reg ( .D(n493), .SI(n8270), .SE(n4083), .CLK(n4547), .Q(
        n8269), .QN(n3792) );
  SDFFX1 DFF_1562_Q_reg ( .D(n494), .SI(n8269), .SE(n4083), .CLK(n4547), .Q(
        n8268), .QN(n3791) );
  SDFFX1 DFF_1563_Q_reg ( .D(n495), .SI(n8268), .SE(n4083), .CLK(n4547), .Q(
        n8267), .QN(n3790) );
  SDFFX1 DFF_1564_Q_reg ( .D(n496), .SI(n8267), .SE(n4083), .CLK(n4547), .Q(
        n8266), .QN(n3789) );
  SDFFX1 DFF_1565_Q_reg ( .D(n497), .SI(n8266), .SE(n4084), .CLK(n4546), .Q(
        n8265), .QN(n3788) );
  SDFFX1 DFF_1566_Q_reg ( .D(n498), .SI(n8265), .SE(n4084), .CLK(n4546), .Q(
        n8264), .QN(n3787) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n4084), .CLK(n4546), 
        .Q(n8263), .QN(n3786) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(n4052), .CLK(n4562), 
        .Q(n8262) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(n4079), .CLK(n4549), 
        .Q(n8261) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(n4078), .CLK(n4549), 
        .Q(n8260) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(n4078), .CLK(n4549), 
        .Q(n8259) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(n4078), .CLK(n4549), 
        .Q(n8258) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(n4077), .CLK(n4550), 
        .Q(n8257) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(n4052), .CLK(n4562), 
        .Q(test_so91) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(n4077), .CLK(n4550), 
        .Q(n8254) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(n4077), .CLK(n4550), 
        .Q(n8253), .QN(n7263) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(n4053), .CLK(n4562), 
        .Q(n8252) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(n4076), .CLK(n4550), 
        .Q(n8251), .QN(n7262) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(n4075), .CLK(n4551), 
        .Q(n8250) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(n4075), .CLK(n4551), 
        .Q(n8249) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(n4074), .CLK(n4551), 
        .Q(n8248) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(n4074), .CLK(n4551), 
        .Q(n8247) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(n4073), .CLK(n4552), 
        .Q(n8246) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(n4072), .CLK(n4552), 
        .Q(WX11021), .QN(n3072) );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(n4072), .CLK(n4552), 
        .Q(WX11023), .QN(n3071) );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(n4071), .CLK(n4553), 
        .Q(WX11025), .QN(n3070) );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(n4070), .CLK(n4553), 
        .Q(WX11027), .QN(n3069) );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(n4070), .CLK(n4553), 
        .Q(WX11029), .QN(n3068) );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(n4069), .CLK(n4554), 
        .Q(WX11031), .QN(n3067) );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(n4068), .CLK(n4554), 
        .Q(WX11033), .QN(n3066) );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(n4068), .CLK(n4554), 
        .Q(test_so92) );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(n4056), .CLK(n4560), 
        .Q(WX11037), .QN(n3065) );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(n4066), .CLK(n4555), 
        .Q(WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(n4066), .CLK(n4555), 
        .Q(WX11041), .QN(n3063) );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(n4065), .CLK(n4556), 
        .Q(WX11043) );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(n4065), .CLK(n4556), 
        .Q(WX11045), .QN(n3062) );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(n4064), .CLK(n4556), 
        .Q(WX11047) );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(n4063), .CLK(n4557), 
        .Q(WX11049), .QN(n3060) );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(n4063), .CLK(n4557), 
        .Q(WX11051), .QN(n3059) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n4062), .CLK(n4557), 
        .Q(WX11053), .QN(n2832) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n4079), .CLK(n4549), 
        .Q(WX11055), .QN(n2871) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n4078), .CLK(n4549), 
        .Q(WX11057), .QN(n2869) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n4078), .CLK(n4549), 
        .Q(WX11059), .QN(n2867) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n4078), .CLK(n4549), 
        .Q(WX11061), .QN(n2865) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n4077), .CLK(n4550), 
        .Q(WX11063), .QN(n2863) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n4077), .CLK(n4550), 
        .Q(WX11065), .QN(n2862) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n4077), .CLK(n4550), 
        .Q(WX11067), .QN(n2860) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n4076), .CLK(n4550), 
        .Q(test_so93) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n4053), .CLK(n4562), 
        .Q(WX11071), .QN(n2857) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n4076), .CLK(n4550), 
        .Q(WX11073), .QN(n2856) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n4075), .CLK(n4551), 
        .Q(WX11075), .QN(n2854) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n4075), .CLK(n4551), 
        .Q(WX11077), .QN(n2853) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n4074), .CLK(n4551), 
        .Q(WX11079), .QN(n2851) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n4074), .CLK(n4551), 
        .Q(WX11081), .QN(n2849) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n4073), .CLK(n4552), 
        .Q(WX11083), .QN(n2847) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n4072), .CLK(n4552), 
        .Q(WX11085) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n4072), .CLK(n4552), 
        .Q(WX11087) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n4071), .CLK(n4553), 
        .Q(WX11089) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n4070), .CLK(n4553), 
        .Q(WX11091) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n4070), .CLK(n4553), 
        .Q(WX11093) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n4069), .CLK(n4554), 
        .Q(WX11095) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n4068), .CLK(n4554), 
        .Q(WX11097) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n4068), .CLK(n4554), 
        .Q(WX11099), .QN(n3547) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n4067), .CLK(n4555), 
        .Q(WX11101) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n4067), .CLK(n4555), 
        .Q(test_so94) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n4066), .CLK(n4555), 
        .Q(WX11105) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n4065), .CLK(n4556), 
        .Q(WX11107), .QN(n3539) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n4064), .CLK(n4556), 
        .Q(WX11109) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n4064), .CLK(n4556), 
        .Q(WX11111), .QN(n3535) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n4063), .CLK(n4557), 
        .Q(WX11113) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n4062), .CLK(n4557), 
        .Q(WX11115) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n4062), .CLK(n4557), 
        .Q(WX11117) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n4061), .CLK(n4558), 
        .Q(WX11119) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n4061), .CLK(n4558), 
        .Q(WX11121) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n4061), .CLK(n4558), 
        .Q(WX11123) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n4060), .CLK(n4558), 
        .Q(WX11125) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n4060), .CLK(n4558), 
        .Q(WX11127) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n4060), .CLK(n4558), 
        .Q(WX11129), .QN(n7264) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n4059), .CLK(n4559), 
        .Q(WX11131) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n4076), .CLK(n4550), 
        .Q(WX11133), .QN(n2859) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n4076), .CLK(n4550), 
        .Q(WX11135) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n4076), .CLK(n4550), 
        .Q(test_so95) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n4075), .CLK(n4551), 
        .Q(WX11139) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n4075), .CLK(n4551), 
        .Q(WX11141) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n4074), .CLK(n4551), 
        .Q(WX11143) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n4073), .CLK(n4552), 
        .Q(WX11145) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n4073), .CLK(n4552), 
        .Q(WX11147) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n4072), .CLK(n4552), 
        .Q(WX11149), .QN(n7261) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n4071), .CLK(n4553), 
        .Q(WX11151), .QN(n7260) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n4071), .CLK(n4553), 
        .Q(WX11153), .QN(n7259) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n4070), .CLK(n4553), 
        .Q(WX11155), .QN(n7258) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155), .SE(n4069), .CLK(n4554), 
        .Q(WX11157), .QN(n7257) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(n4069), .CLK(n4554), 
        .Q(WX11159), .QN(n7256) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(n4068), .CLK(n4554), 
        .Q(WX11161), .QN(n7255) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(n4067), .CLK(n4555), 
        .Q(WX11163) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(n4067), .CLK(n4555), 
        .Q(WX11165), .QN(n7254) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(n4066), .CLK(n4555), 
        .Q(WX11167), .QN(n3064) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(n4066), .CLK(n4555), 
        .Q(WX11169), .QN(n7253) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(n4065), .CLK(n4556), 
        .Q(test_so96) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n4064), .CLK(n4556), 
        .Q(WX11173), .QN(n7252) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n4064), .CLK(n4556), 
        .Q(WX11175), .QN(n3061) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n4063), .CLK(n4557), 
        .Q(WX11177), .QN(n7251) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n4062), .CLK(n4557), 
        .Q(WX11179), .QN(n7250) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n4062), .CLK(n4557), 
        .Q(WX11181), .QN(n3202) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n4061), .CLK(n4558), 
        .Q(WX11183), .QN(n3203) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n4061), .CLK(n4558), 
        .Q(WX11185), .QN(n3204) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n4061), .CLK(n4558), 
        .Q(WX11187), .QN(n3205) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n4060), .CLK(n4558), 
        .Q(WX11189), .QN(n3206) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n4060), .CLK(n4558), 
        .Q(WX11191), .QN(n3207) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n4060), .CLK(n4558), 
        .Q(WX11193), .QN(n3208) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n4059), .CLK(n4559), 
        .Q(WX11195), .QN(n3209) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n4059), .CLK(n4559), 
        .Q(WX11197), .QN(n3210) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n4059), .CLK(n4559), 
        .Q(WX11199), .QN(n3211) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n4059), .CLK(n4559), 
        .Q(WX11201), .QN(n3212) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n4059), .CLK(n4559), 
        .Q(WX11203), .QN(n3213) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n4058), .CLK(n4559), 
        .Q(test_so97) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n4074), .CLK(n4551), 
        .Q(WX11207), .QN(n3214) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n4073), .CLK(n4552), 
        .Q(WX11209), .QN(n3215) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n4073), .CLK(n4552), 
        .Q(WX11211), .QN(n3173) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n4072), .CLK(n4552), 
        .Q(WX11213), .QN(n3216) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n4071), .CLK(n4553), 
        .Q(WX11215), .QN(n3217) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n4071), .CLK(n4553), 
        .Q(WX11217), .QN(n3218) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n4070), .CLK(n4553), 
        .Q(WX11219), .QN(n3219) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n4069), .CLK(n4554), 
        .Q(WX11221), .QN(n3174) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n4069), .CLK(n4554), 
        .Q(WX11223), .QN(n3220) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n4068), .CLK(n4554), 
        .Q(WX11225), .QN(n3221) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n4067), .CLK(n4555), 
        .Q(WX11227), .QN(n3222) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n4067), .CLK(n4555), 
        .Q(WX11229), .QN(n3223) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n4066), .CLK(n4555), 
        .Q(WX11231), .QN(n3224) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n4065), .CLK(n4556), 
        .Q(WX11233), .QN(n3225) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n4065), .CLK(n4556), 
        .Q(WX11235), .QN(n3175) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n4064), .CLK(n4556), 
        .Q(WX11237), .QN(n3226) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n4063), .CLK(n4557), 
        .Q(test_so98) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n4063), .CLK(n4557), 
        .Q(WX11241), .QN(n3227) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n4062), .CLK(n4557), 
        .Q(WX11243), .QN(n3194) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n4057), .CLK(n4560), 
        .Q(CRC_OUT_1_0) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n4057), .CLK(
        n4560), .Q(CRC_OUT_1_1), .QN(DFF_1697_n1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n4057), .CLK(
        n4560), .Q(CRC_OUT_1_2) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n4056), .CLK(
        n4560), .Q(CRC_OUT_1_3) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n4056), .CLK(
        n4560), .Q(CRC_OUT_1_4) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n4056), .CLK(
        n4560), .Q(CRC_OUT_1_5) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n4056), .CLK(
        n4560), .Q(CRC_OUT_1_6) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n4056), .CLK(
        n4560), .Q(CRC_OUT_1_7) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n4055), .CLK(
        n4561), .Q(CRC_OUT_1_8) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n4055), .CLK(
        n4561), .Q(CRC_OUT_1_9) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n4055), .CLK(
        n4561), .Q(CRC_OUT_1_10) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n4055), .CLK(
        n4561), .Q(CRC_OUT_1_11) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n4055), .CLK(
        n4561), .Q(CRC_OUT_1_12) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n4055), .CLK(
        n4561), .Q(CRC_OUT_1_13) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n4054), .CLK(
        n4561), .Q(test_so99) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n4054), .CLK(n4561), .Q(CRC_OUT_1_15) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n4054), .CLK(
        n4561), .Q(CRC_OUT_1_16) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n4054), .CLK(
        n4561), .Q(CRC_OUT_1_17) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n4054), .CLK(
        n4561), .Q(CRC_OUT_1_18), .QN(DFF_1714_n1) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n4054), .CLK(
        n4561), .Q(CRC_OUT_1_19) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n4053), .CLK(
        n4562), .Q(CRC_OUT_1_20) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n4053), .CLK(
        n4562), .Q(CRC_OUT_1_21) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n4053), .CLK(
        n4562), .Q(CRC_OUT_1_22) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n4053), .CLK(
        n4562), .Q(CRC_OUT_1_23) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n4058), .CLK(
        n4559), .Q(CRC_OUT_1_24) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n4058), .CLK(
        n4559), .Q(CRC_OUT_1_25) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n4058), .CLK(
        n4559), .Q(CRC_OUT_1_26) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n4058), .CLK(
        n4559), .Q(CRC_OUT_1_27) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n4058), .CLK(
        n4559), .Q(CRC_OUT_1_28) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n4057), .CLK(
        n4560), .Q(CRC_OUT_1_29) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n4057), .CLK(
        n4560), .Q(CRC_OUT_1_30) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n4057), .CLK(
        n4560), .Q(test_so100) );
  NOR2X0 Trojan1 ( .IN1(WX3442), .IN2(WX5974), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(WX806), .IN2(WX782), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(WX11632), .IN2(n112), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(WX5964), .IN2(WX3324), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(WX8634), .IN2(WX3330), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n124), .IN2(n116), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(WX862), .IN2(WX7227), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(WX11616), .IN2(n485), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  INVX0 TrojanINVtest_se ( .INP(n4325), .ZN(test_se_NOT) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(test_se_NOT), .Q(Tj_Trigger) );
  INVX0 U3578 ( .INP(TM1), .ZN(n3514) );
  INVX0 U3579 ( .INP(TM1), .ZN(n3515) );
  INVX0 U3580 ( .INP(TM1), .ZN(n3516) );
  INVX0 U3581 ( .INP(TM1), .ZN(n3518) );
  NBUFFX2 U3582 ( .INP(n3616), .Z(n3588) );
  NBUFFX2 U3583 ( .INP(n3616), .Z(n3589) );
  NBUFFX2 U3584 ( .INP(n3614), .Z(n3598) );
  NBUFFX2 U3585 ( .INP(n3614), .Z(n3600) );
  NBUFFX2 U3586 ( .INP(n3612), .Z(n3601) );
  NBUFFX2 U3587 ( .INP(n3612), .Z(n3602) );
  NBUFFX2 U3588 ( .INP(n3612), .Z(n3603) );
  NBUFFX2 U3589 ( .INP(n3612), .Z(n3604) );
  NBUFFX2 U3590 ( .INP(n3612), .Z(n3605) );
  NBUFFX2 U3591 ( .INP(n3611), .Z(n3609) );
  NBUFFX2 U3592 ( .INP(n3615), .Z(n3590) );
  NBUFFX2 U3593 ( .INP(n3615), .Z(n3592) );
  NBUFFX2 U3594 ( .INP(n3615), .Z(n3593) );
  NBUFFX2 U3595 ( .INP(n3614), .Z(n3599) );
  NBUFFX2 U3596 ( .INP(n3615), .Z(n3594) );
  NBUFFX2 U3597 ( .INP(n3615), .Z(n3595) );
  NBUFFX2 U3598 ( .INP(n3614), .Z(n3596) );
  NBUFFX2 U3599 ( .INP(n3614), .Z(n3597) );
  NBUFFX2 U3600 ( .INP(n3611), .Z(n3606) );
  NBUFFX2 U3601 ( .INP(n3611), .Z(n3607) );
  NBUFFX2 U3602 ( .INP(n3611), .Z(n3608) );
  NBUFFX2 U3603 ( .INP(n3616), .Z(n3587) );
  NBUFFX2 U3604 ( .INP(n4663), .Z(n4494) );
  NBUFFX2 U3605 ( .INP(n4663), .Z(n4492) );
  NBUFFX2 U3606 ( .INP(n4663), .Z(n4493) );
  NBUFFX2 U3607 ( .INP(n4663), .Z(n4491) );
  NBUFFX2 U3608 ( .INP(n4649), .Z(n4561) );
  NBUFFX2 U3609 ( .INP(n4650), .Z(n4559) );
  NBUFFX2 U3610 ( .INP(n4650), .Z(n4558) );
  NBUFFX2 U3611 ( .INP(n4650), .Z(n4557) );
  NBUFFX2 U3612 ( .INP(n4650), .Z(n4556) );
  NBUFFX2 U3613 ( .INP(n4650), .Z(n4555) );
  NBUFFX2 U3614 ( .INP(n4649), .Z(n4560) );
  NBUFFX2 U3615 ( .INP(n4651), .Z(n4554) );
  NBUFFX2 U3616 ( .INP(n4651), .Z(n4553) );
  NBUFFX2 U3617 ( .INP(n4651), .Z(n4552) );
  NBUFFX2 U3618 ( .INP(n4651), .Z(n4551) );
  NBUFFX2 U3619 ( .INP(n4651), .Z(n4550) );
  NBUFFX2 U3620 ( .INP(n4652), .Z(n4547) );
  NBUFFX2 U3621 ( .INP(n4652), .Z(n4548) );
  NBUFFX2 U3622 ( .INP(n4652), .Z(n4549) );
  NBUFFX2 U3623 ( .INP(n4652), .Z(n4546) );
  NBUFFX2 U3624 ( .INP(n4649), .Z(n4563) );
  NBUFFX2 U3625 ( .INP(n4652), .Z(n4545) );
  NBUFFX2 U3626 ( .INP(n4653), .Z(n4544) );
  NBUFFX2 U3627 ( .INP(n4653), .Z(n4543) );
  NBUFFX2 U3628 ( .INP(n4653), .Z(n4542) );
  NBUFFX2 U3629 ( .INP(n4649), .Z(n4562) );
  NBUFFX2 U3630 ( .INP(n4653), .Z(n4541) );
  NBUFFX2 U3631 ( .INP(n4653), .Z(n4540) );
  NBUFFX2 U3632 ( .INP(n4654), .Z(n4539) );
  NBUFFX2 U3633 ( .INP(n4654), .Z(n4538) );
  NBUFFX2 U3634 ( .INP(n4654), .Z(n4537) );
  NBUFFX2 U3635 ( .INP(n4654), .Z(n4536) );
  NBUFFX2 U3636 ( .INP(n4655), .Z(n4533) );
  NBUFFX2 U3637 ( .INP(n4655), .Z(n4534) );
  NBUFFX2 U3638 ( .INP(n4655), .Z(n4532) );
  NBUFFX2 U3639 ( .INP(n4655), .Z(n4531) );
  NBUFFX2 U3640 ( .INP(n4649), .Z(n4564) );
  NBUFFX2 U3641 ( .INP(n4655), .Z(n4530) );
  NBUFFX2 U3642 ( .INP(n4657), .Z(n4524) );
  NBUFFX2 U3643 ( .INP(n4657), .Z(n4523) );
  NBUFFX2 U3644 ( .INP(n4657), .Z(n4522) );
  NBUFFX2 U3645 ( .INP(n4657), .Z(n4521) );
  NBUFFX2 U3646 ( .INP(n4656), .Z(n4529) );
  NBUFFX2 U3647 ( .INP(n4656), .Z(n4528) );
  NBUFFX2 U3648 ( .INP(n4656), .Z(n4527) );
  NBUFFX2 U3649 ( .INP(n4656), .Z(n4526) );
  NBUFFX2 U3650 ( .INP(n4654), .Z(n4535) );
  NBUFFX2 U3651 ( .INP(n4656), .Z(n4525) );
  NBUFFX2 U3652 ( .INP(n4658), .Z(n4519) );
  NBUFFX2 U3653 ( .INP(n4657), .Z(n4520) );
  NBUFFX2 U3654 ( .INP(n4658), .Z(n4518) );
  NBUFFX2 U3655 ( .INP(n4638), .Z(n4618) );
  NBUFFX2 U3656 ( .INP(n4638), .Z(n4617) );
  NBUFFX2 U3657 ( .INP(n4638), .Z(n4616) );
  NBUFFX2 U3658 ( .INP(n4638), .Z(n4615) );
  NBUFFX2 U3659 ( .INP(n4639), .Z(n4614) );
  NBUFFX2 U3660 ( .INP(n4639), .Z(n4613) );
  NBUFFX2 U3661 ( .INP(n4638), .Z(n4619) );
  NBUFFX2 U3662 ( .INP(n4639), .Z(n4612) );
  NBUFFX2 U3663 ( .INP(n4639), .Z(n4611) );
  NBUFFX2 U3664 ( .INP(n4639), .Z(n4610) );
  NBUFFX2 U3665 ( .INP(n4640), .Z(n4609) );
  NBUFFX2 U3666 ( .INP(n4640), .Z(n4608) );
  NBUFFX2 U3667 ( .INP(n4640), .Z(n4606) );
  NBUFFX2 U3668 ( .INP(n4640), .Z(n4607) );
  NBUFFX2 U3669 ( .INP(n4640), .Z(n4605) );
  NBUFFX2 U3670 ( .INP(n4637), .Z(n4620) );
  NBUFFX2 U3671 ( .INP(n4641), .Z(n4604) );
  NBUFFX2 U3672 ( .INP(n4641), .Z(n4603) );
  NBUFFX2 U3673 ( .INP(n4641), .Z(n4602) );
  NBUFFX2 U3674 ( .INP(n4641), .Z(n4601) );
  NBUFFX2 U3675 ( .INP(n4641), .Z(n4600) );
  NBUFFX2 U3676 ( .INP(n4637), .Z(n4621) );
  NBUFFX2 U3677 ( .INP(n4642), .Z(n4599) );
  NBUFFX2 U3678 ( .INP(n4642), .Z(n4598) );
  NBUFFX2 U3679 ( .INP(n4642), .Z(n4597) );
  NBUFFX2 U3680 ( .INP(n4642), .Z(n4596) );
  NBUFFX2 U3681 ( .INP(n4642), .Z(n4595) );
  NBUFFX2 U3682 ( .INP(n4643), .Z(n4594) );
  NBUFFX2 U3683 ( .INP(n4637), .Z(n4622) );
  NBUFFX2 U3684 ( .INP(n4643), .Z(n4592) );
  NBUFFX2 U3685 ( .INP(n4643), .Z(n4593) );
  NBUFFX2 U3686 ( .INP(n4643), .Z(n4591) );
  NBUFFX2 U3687 ( .INP(n4637), .Z(n4624) );
  NBUFFX2 U3688 ( .INP(n4643), .Z(n4590) );
  NBUFFX2 U3689 ( .INP(n4644), .Z(n4589) );
  NBUFFX2 U3690 ( .INP(n4644), .Z(n4588) );
  NBUFFX2 U3691 ( .INP(n4644), .Z(n4587) );
  NBUFFX2 U3692 ( .INP(n4644), .Z(n4586) );
  NBUFFX2 U3693 ( .INP(n4644), .Z(n4585) );
  NBUFFX2 U3694 ( .INP(n4645), .Z(n4584) );
  NBUFFX2 U3695 ( .INP(n4645), .Z(n4583) );
  NBUFFX2 U3696 ( .INP(n4645), .Z(n4582) );
  NBUFFX2 U3697 ( .INP(n4645), .Z(n4581) );
  NBUFFX2 U3698 ( .INP(n4637), .Z(n4623) );
  NBUFFX2 U3699 ( .INP(n4646), .Z(n4578) );
  NBUFFX2 U3700 ( .INP(n4646), .Z(n4579) );
  NBUFFX2 U3701 ( .INP(n4646), .Z(n4577) );
  NBUFFX2 U3702 ( .INP(n4646), .Z(n4576) );
  NBUFFX2 U3703 ( .INP(n4646), .Z(n4575) );
  NBUFFX2 U3704 ( .INP(n4647), .Z(n4574) );
  NBUFFX2 U3705 ( .INP(n4648), .Z(n4569) );
  NBUFFX2 U3706 ( .INP(n4648), .Z(n4568) );
  NBUFFX2 U3707 ( .INP(n4648), .Z(n4567) );
  NBUFFX2 U3708 ( .INP(n4648), .Z(n4566) );
  NBUFFX2 U3709 ( .INP(n4648), .Z(n4565) );
  NBUFFX2 U3710 ( .INP(n4647), .Z(n4573) );
  NBUFFX2 U3711 ( .INP(n4647), .Z(n4572) );
  NBUFFX2 U3712 ( .INP(n4647), .Z(n4571) );
  NBUFFX2 U3713 ( .INP(n4636), .Z(n4626) );
  NBUFFX2 U3714 ( .INP(n4636), .Z(n4625) );
  NBUFFX2 U3715 ( .INP(n4645), .Z(n4580) );
  NBUFFX2 U3716 ( .INP(n4647), .Z(n4570) );
  NBUFFX2 U3717 ( .INP(n4658), .Z(n4516) );
  NBUFFX2 U3718 ( .INP(n4658), .Z(n4517) );
  NBUFFX2 U3719 ( .INP(n4658), .Z(n4515) );
  NBUFFX2 U3720 ( .INP(n4659), .Z(n4514) );
  NBUFFX2 U3721 ( .INP(n4636), .Z(n4627) );
  NBUFFX2 U3722 ( .INP(n4659), .Z(n4513) );
  NBUFFX2 U3723 ( .INP(n4659), .Z(n4512) );
  NBUFFX2 U3724 ( .INP(n4635), .Z(n4631) );
  NBUFFX2 U3725 ( .INP(n4635), .Z(n4630) );
  NBUFFX2 U3726 ( .INP(n4636), .Z(n4629) );
  NBUFFX2 U3727 ( .INP(n4659), .Z(n4511) );
  NBUFFX2 U3728 ( .INP(n4659), .Z(n4510) );
  NBUFFX2 U3729 ( .INP(n4635), .Z(n4632) );
  NBUFFX2 U3730 ( .INP(n4636), .Z(n4628) );
  NBUFFX2 U3731 ( .INP(n4660), .Z(n4509) );
  NBUFFX2 U3732 ( .INP(n4660), .Z(n4508) );
  NBUFFX2 U3733 ( .INP(n4660), .Z(n4506) );
  NBUFFX2 U3734 ( .INP(n4660), .Z(n4507) );
  NBUFFX2 U3735 ( .INP(n4660), .Z(n4505) );
  NBUFFX2 U3736 ( .INP(n4635), .Z(n4633) );
  NBUFFX2 U3737 ( .INP(n4661), .Z(n4504) );
  NBUFFX2 U3738 ( .INP(n4661), .Z(n4503) );
  NBUFFX2 U3739 ( .INP(n4661), .Z(n4502) );
  NBUFFX2 U3740 ( .INP(n4661), .Z(n4501) );
  NBUFFX2 U3741 ( .INP(n4661), .Z(n4500) );
  NBUFFX2 U3742 ( .INP(n4662), .Z(n4499) );
  NBUFFX2 U3743 ( .INP(n4662), .Z(n4498) );
  NBUFFX2 U3744 ( .INP(n4662), .Z(n4497) );
  NBUFFX2 U3745 ( .INP(n4662), .Z(n4496) );
  NBUFFX2 U3746 ( .INP(n4662), .Z(n4495) );
  NBUFFX2 U3747 ( .INP(n4635), .Z(n4634) );
  NBUFFX2 U3748 ( .INP(n3611), .Z(n3610) );
  NBUFFX2 U3749 ( .INP(n3650), .Z(n3628) );
  NBUFFX2 U3750 ( .INP(n3648), .Z(n3636) );
  NBUFFX2 U3751 ( .INP(n3648), .Z(n3637) );
  NBUFFX2 U3752 ( .INP(n3648), .Z(n3638) );
  NBUFFX2 U3753 ( .INP(n3648), .Z(n3640) );
  NBUFFX2 U3754 ( .INP(n3646), .Z(n3644) );
  NBUFFX2 U3755 ( .INP(n3649), .Z(n3630) );
  NBUFFX2 U3756 ( .INP(n3649), .Z(n3631) );
  NBUFFX2 U3757 ( .INP(n3649), .Z(n3632) );
  NBUFFX2 U3758 ( .INP(n3649), .Z(n3629) );
  NBUFFX2 U3759 ( .INP(n3648), .Z(n3634) );
  NBUFFX2 U3760 ( .INP(n3649), .Z(n3633) );
  NBUFFX2 U3761 ( .INP(n3646), .Z(n3641) );
  NBUFFX2 U3762 ( .INP(n3646), .Z(n3642) );
  NBUFFX2 U3763 ( .INP(n3646), .Z(n3643) );
  NBUFFX2 U3764 ( .INP(n3651), .Z(n3620) );
  NBUFFX2 U3765 ( .INP(n3651), .Z(n3622) );
  NBUFFX2 U3766 ( .INP(n3651), .Z(n3621) );
  NBUFFX2 U3767 ( .INP(n3650), .Z(n3627) );
  NBUFFX2 U3768 ( .INP(n3650), .Z(n3626) );
  NBUFFX2 U3769 ( .INP(n3650), .Z(n3623) );
  NBUFFX2 U3770 ( .INP(n3650), .Z(n3624) );
  NBUFFX2 U3771 ( .INP(n3646), .Z(n3645) );
  NBUFFX2 U3772 ( .INP(n3522), .Z(n3534) );
  NBUFFX2 U3773 ( .INP(n3526), .Z(n3553) );
  NBUFFX2 U3774 ( .INP(n3526), .Z(n3552) );
  NBUFFX2 U3775 ( .INP(n3523), .Z(n3544) );
  NBUFFX2 U3776 ( .INP(n3523), .Z(n3543) );
  NBUFFX2 U3777 ( .INP(n3523), .Z(n3542) );
  NBUFFX2 U3778 ( .INP(n3523), .Z(n3541) );
  NBUFFX2 U3779 ( .INP(n3522), .Z(n3540) );
  NBUFFX2 U3780 ( .INP(n3524), .Z(n3551) );
  NBUFFX2 U3781 ( .INP(n3524), .Z(n3550) );
  NBUFFX2 U3782 ( .INP(n3524), .Z(n3549) );
  NBUFFX2 U3783 ( .INP(n3524), .Z(n3548) );
  NBUFFX2 U3784 ( .INP(n3524), .Z(n3546) );
  NBUFFX2 U3785 ( .INP(n3523), .Z(n3545) );
  NBUFFX2 U3786 ( .INP(n3522), .Z(n3536) );
  NBUFFX2 U3787 ( .INP(n3522), .Z(n3537) );
  NBUFFX2 U3788 ( .INP(n3522), .Z(n3538) );
  NBUFFX2 U3789 ( .INP(n3559), .Z(n3583) );
  NBUFFX2 U3790 ( .INP(n3559), .Z(n3582) );
  NBUFFX2 U3791 ( .INP(n3559), .Z(n3581) );
  NBUFFX2 U3792 ( .INP(n3555), .Z(n3561) );
  NBUFFX2 U3793 ( .INP(n3555), .Z(n3560) );
  NBUFFX2 U3794 ( .INP(n3558), .Z(n3580) );
  NBUFFX2 U3795 ( .INP(n3558), .Z(n3579) );
  NBUFFX2 U3796 ( .INP(n3558), .Z(n3578) );
  NBUFFX2 U3797 ( .INP(n3558), .Z(n3577) );
  NBUFFX2 U3798 ( .INP(n3557), .Z(n3572) );
  NBUFFX2 U3799 ( .INP(n3557), .Z(n3571) );
  NBUFFX2 U3800 ( .INP(n3556), .Z(n3570) );
  NBUFFX2 U3801 ( .INP(n3556), .Z(n3568) );
  NBUFFX2 U3802 ( .INP(n3556), .Z(n3567) );
  NBUFFX2 U3803 ( .INP(n3556), .Z(n3566) );
  NBUFFX2 U3804 ( .INP(n3556), .Z(n3565) );
  NBUFFX2 U3805 ( .INP(n3555), .Z(n3564) );
  NBUFFX2 U3806 ( .INP(n3555), .Z(n3563) );
  NBUFFX2 U3807 ( .INP(n3555), .Z(n3562) );
  NBUFFX2 U3808 ( .INP(n3558), .Z(n3576) );
  NBUFFX2 U3809 ( .INP(n3557), .Z(n3575) );
  NBUFFX2 U3810 ( .INP(n3557), .Z(n3574) );
  NBUFFX2 U3811 ( .INP(n3557), .Z(n3573) );
  NBUFFX2 U3812 ( .INP(n3520), .Z(n3533) );
  NBUFFX2 U3813 ( .INP(n3520), .Z(n3532) );
  NBUFFX2 U3814 ( .INP(n3520), .Z(n3531) );
  NBUFFX2 U3815 ( .INP(n3520), .Z(n3530) );
  NBUFFX2 U3816 ( .INP(n3520), .Z(n3528) );
  NBUFFX2 U3817 ( .INP(n3526), .Z(n3554) );
  NBUFFX2 U3818 ( .INP(n3559), .Z(n3584) );
  NBUFFX2 U3819 ( .INP(n4694), .Z(n3520) );
  NBUFFX2 U3820 ( .INP(n4694), .Z(n3522) );
  NBUFFX2 U3821 ( .INP(n4694), .Z(n3523) );
  NBUFFX2 U3822 ( .INP(n4694), .Z(n3524) );
  NBUFFX2 U3823 ( .INP(n4694), .Z(n3526) );
  NBUFFX2 U3824 ( .INP(n2148), .Z(n3555) );
  NBUFFX2 U3825 ( .INP(n2148), .Z(n3556) );
  NBUFFX2 U3826 ( .INP(n2148), .Z(n3557) );
  NBUFFX2 U3827 ( .INP(n2148), .Z(n3558) );
  NBUFFX2 U3828 ( .INP(n2148), .Z(n3559) );
  NBUFFX2 U3829 ( .INP(n2152), .Z(n3585) );
  NBUFFX2 U3830 ( .INP(n2152), .Z(n3586) );
  NBUFFX2 U3831 ( .INP(n3585), .Z(n3611) );
  NBUFFX2 U3832 ( .INP(n3585), .Z(n3612) );
  NBUFFX2 U3833 ( .INP(n3585), .Z(n3614) );
  NBUFFX2 U3834 ( .INP(n3586), .Z(n3615) );
  NBUFFX2 U3835 ( .INP(n3586), .Z(n3616) );
  NBUFFX2 U3836 ( .INP(n2153), .Z(n3618) );
  NBUFFX2 U3837 ( .INP(n2153), .Z(n3619) );
  NBUFFX2 U3838 ( .INP(n3618), .Z(n3646) );
  NBUFFX2 U3839 ( .INP(n3618), .Z(n3648) );
  NBUFFX2 U3840 ( .INP(n3618), .Z(n3649) );
  NBUFFX2 U3841 ( .INP(n3619), .Z(n3650) );
  NBUFFX2 U3842 ( .INP(n3619), .Z(n3651) );
  NBUFFX2 U3843 ( .INP(n4292), .Z(n3652) );
  NBUFFX2 U3844 ( .INP(n4291), .Z(n3653) );
  NBUFFX2 U3845 ( .INP(n4291), .Z(n3654) );
  NBUFFX2 U3846 ( .INP(n4291), .Z(n3655) );
  NBUFFX2 U3847 ( .INP(n4290), .Z(n3656) );
  NBUFFX2 U3848 ( .INP(n4290), .Z(n3657) );
  NBUFFX2 U3849 ( .INP(n4290), .Z(n3658) );
  NBUFFX2 U3850 ( .INP(n4289), .Z(n3659) );
  NBUFFX2 U3851 ( .INP(n4289), .Z(n3660) );
  NBUFFX2 U3852 ( .INP(n4289), .Z(n3662) );
  NBUFFX2 U3853 ( .INP(n4288), .Z(n3663) );
  NBUFFX2 U3854 ( .INP(n4288), .Z(n3664) );
  NBUFFX2 U3855 ( .INP(n4288), .Z(n3665) );
  NBUFFX2 U3856 ( .INP(n4287), .Z(n3666) );
  NBUFFX2 U3857 ( .INP(n4287), .Z(n3667) );
  NBUFFX2 U3858 ( .INP(n4287), .Z(n3668) );
  NBUFFX2 U3859 ( .INP(n4286), .Z(n3670) );
  NBUFFX2 U3860 ( .INP(n4286), .Z(n3671) );
  NBUFFX2 U3861 ( .INP(n4286), .Z(n3672) );
  NBUFFX2 U3862 ( .INP(n4285), .Z(n3673) );
  NBUFFX2 U3863 ( .INP(n4285), .Z(n3674) );
  NBUFFX2 U3864 ( .INP(n4285), .Z(n3675) );
  NBUFFX2 U3865 ( .INP(n4284), .Z(n3676) );
  NBUFFX2 U3866 ( .INP(n4284), .Z(n3677) );
  NBUFFX2 U3867 ( .INP(n4284), .Z(n3678) );
  NBUFFX2 U3868 ( .INP(n4283), .Z(n3679) );
  NBUFFX2 U3869 ( .INP(n4283), .Z(n3680) );
  NBUFFX2 U3870 ( .INP(n4283), .Z(n3681) );
  NBUFFX2 U3872 ( .INP(n4282), .Z(n3682) );
  NBUFFX2 U3873 ( .INP(n4282), .Z(n3683) );
  NBUFFX2 U3874 ( .INP(n4282), .Z(n3684) );
  NBUFFX2 U3875 ( .INP(n4281), .Z(n3685) );
  NBUFFX2 U3876 ( .INP(n4281), .Z(n3686) );
  NBUFFX2 U3877 ( .INP(n4281), .Z(n3687) );
  NBUFFX2 U3878 ( .INP(n4280), .Z(n3688) );
  NBUFFX2 U3879 ( .INP(n4280), .Z(n3689) );
  NBUFFX2 U3880 ( .INP(n4280), .Z(n3690) );
  NBUFFX2 U3881 ( .INP(n4279), .Z(n3692) );
  NBUFFX2 U3882 ( .INP(n4279), .Z(n3693) );
  NBUFFX2 U3883 ( .INP(n4279), .Z(n3694) );
  NBUFFX2 U3884 ( .INP(n4278), .Z(n3695) );
  NBUFFX2 U3885 ( .INP(n4278), .Z(n3696) );
  NBUFFX2 U3886 ( .INP(n4278), .Z(n3697) );
  NBUFFX2 U3887 ( .INP(n4277), .Z(n3698) );
  NBUFFX2 U3888 ( .INP(n4277), .Z(n3699) );
  NBUFFX2 U3889 ( .INP(n4277), .Z(n3700) );
  NBUFFX2 U3890 ( .INP(n4276), .Z(n3701) );
  NBUFFX2 U3891 ( .INP(n4276), .Z(n3702) );
  NBUFFX2 U3892 ( .INP(n4276), .Z(n3703) );
  NBUFFX2 U3893 ( .INP(n4275), .Z(n3704) );
  NBUFFX2 U3894 ( .INP(n4275), .Z(n3705) );
  NBUFFX2 U3895 ( .INP(n4275), .Z(n3706) );
  NBUFFX2 U3896 ( .INP(n4274), .Z(n3707) );
  NBUFFX2 U3897 ( .INP(n4274), .Z(n3708) );
  NBUFFX2 U3898 ( .INP(n4274), .Z(n3709) );
  NBUFFX2 U3899 ( .INP(n4273), .Z(n3710) );
  NBUFFX2 U3900 ( .INP(n4273), .Z(n3711) );
  NBUFFX2 U3901 ( .INP(n4273), .Z(n3712) );
  NBUFFX2 U3902 ( .INP(n4272), .Z(n3714) );
  NBUFFX2 U3903 ( .INP(n4272), .Z(n3715) );
  NBUFFX2 U3904 ( .INP(n4272), .Z(n3716) );
  NBUFFX2 U3905 ( .INP(n4271), .Z(n3718) );
  NBUFFX2 U3906 ( .INP(n4271), .Z(n3719) );
  NBUFFX2 U3907 ( .INP(n4271), .Z(n3720) );
  NBUFFX2 U3908 ( .INP(n4270), .Z(n3721) );
  NBUFFX2 U3909 ( .INP(n4270), .Z(n3722) );
  NBUFFX2 U3910 ( .INP(n4270), .Z(n3723) );
  NBUFFX2 U3911 ( .INP(n4269), .Z(n3724) );
  NBUFFX2 U3912 ( .INP(n4269), .Z(n3725) );
  NBUFFX2 U3913 ( .INP(n4269), .Z(n3726) );
  NBUFFX2 U3914 ( .INP(n4268), .Z(n3727) );
  NBUFFX2 U3915 ( .INP(n4268), .Z(n3728) );
  NBUFFX2 U3916 ( .INP(n4268), .Z(n3729) );
  NBUFFX2 U3917 ( .INP(n4267), .Z(n3730) );
  NBUFFX2 U3918 ( .INP(n4267), .Z(n3731) );
  NBUFFX2 U3919 ( .INP(n4267), .Z(n3732) );
  NBUFFX2 U3920 ( .INP(n4266), .Z(n3733) );
  NBUFFX2 U3921 ( .INP(n4266), .Z(n3734) );
  NBUFFX2 U3922 ( .INP(n4266), .Z(n3736) );
  NBUFFX2 U3923 ( .INP(n4265), .Z(n3737) );
  NBUFFX2 U3924 ( .INP(n4265), .Z(n3738) );
  NBUFFX2 U3925 ( .INP(n4265), .Z(n3740) );
  NBUFFX2 U3926 ( .INP(n4264), .Z(n3741) );
  NBUFFX2 U3927 ( .INP(n4264), .Z(n3742) );
  NBUFFX2 U3928 ( .INP(n4264), .Z(n3743) );
  NBUFFX2 U3929 ( .INP(n4263), .Z(n3744) );
  NBUFFX2 U3930 ( .INP(n4263), .Z(n3745) );
  NBUFFX2 U3931 ( .INP(n4263), .Z(n3746) );
  NBUFFX2 U3932 ( .INP(n4262), .Z(n3747) );
  NBUFFX2 U3933 ( .INP(n4262), .Z(n3748) );
  NBUFFX2 U3934 ( .INP(n4262), .Z(n3749) );
  NBUFFX2 U3935 ( .INP(n4261), .Z(n3750) );
  NBUFFX2 U3936 ( .INP(n4261), .Z(n3751) );
  NBUFFX2 U3937 ( .INP(n4261), .Z(n3752) );
  NBUFFX2 U3938 ( .INP(n4260), .Z(n3753) );
  NBUFFX2 U3939 ( .INP(n4260), .Z(n3754) );
  NBUFFX2 U3940 ( .INP(n4260), .Z(n3755) );
  NBUFFX2 U3941 ( .INP(n4259), .Z(n3756) );
  NBUFFX2 U3942 ( .INP(n4259), .Z(n3757) );
  NBUFFX2 U3943 ( .INP(n4259), .Z(n3758) );
  NBUFFX2 U3944 ( .INP(n4258), .Z(n3759) );
  NBUFFX2 U3945 ( .INP(n4258), .Z(n3760) );
  NBUFFX2 U3946 ( .INP(n4258), .Z(n3761) );
  NBUFFX2 U3947 ( .INP(n4257), .Z(n3762) );
  NBUFFX2 U3948 ( .INP(n4257), .Z(n3764) );
  NBUFFX2 U3949 ( .INP(n4257), .Z(n3765) );
  NBUFFX2 U3950 ( .INP(n4256), .Z(n3766) );
  NBUFFX2 U3951 ( .INP(n4256), .Z(n3767) );
  NBUFFX2 U3952 ( .INP(n4256), .Z(n3768) );
  NBUFFX2 U3953 ( .INP(n4255), .Z(n3769) );
  NBUFFX2 U3954 ( .INP(n4255), .Z(n3770) );
  NBUFFX2 U3955 ( .INP(n4255), .Z(n3771) );
  NBUFFX2 U3956 ( .INP(n4254), .Z(n3772) );
  NBUFFX2 U3957 ( .INP(n4254), .Z(n3773) );
  NBUFFX2 U3958 ( .INP(n4254), .Z(n3774) );
  NBUFFX2 U3959 ( .INP(n4253), .Z(n3776) );
  NBUFFX2 U3960 ( .INP(n4253), .Z(n3777) );
  NBUFFX2 U3961 ( .INP(n4253), .Z(n3778) );
  NBUFFX2 U3962 ( .INP(n4252), .Z(n3779) );
  NBUFFX2 U3963 ( .INP(n4252), .Z(n3780) );
  NBUFFX2 U3964 ( .INP(n4252), .Z(n3781) );
  NBUFFX2 U3965 ( .INP(n4251), .Z(n3782) );
  NBUFFX2 U3966 ( .INP(n4251), .Z(n3784) );
  NBUFFX2 U3967 ( .INP(n4251), .Z(n3785) );
  NBUFFX2 U3968 ( .INP(n4250), .Z(n3866) );
  NBUFFX2 U3969 ( .INP(n4250), .Z(n3884) );
  NBUFFX2 U3970 ( .INP(n4250), .Z(n4034) );
  NBUFFX2 U3971 ( .INP(n4249), .Z(n4035) );
  NBUFFX2 U3972 ( .INP(n4249), .Z(n4036) );
  NBUFFX2 U3973 ( .INP(n4249), .Z(n4037) );
  NBUFFX2 U3974 ( .INP(n4248), .Z(n4038) );
  NBUFFX2 U3975 ( .INP(n4248), .Z(n4039) );
  NBUFFX2 U3976 ( .INP(n4248), .Z(n4040) );
  NBUFFX2 U3977 ( .INP(n4247), .Z(n4041) );
  NBUFFX2 U3978 ( .INP(n4247), .Z(n4042) );
  NBUFFX2 U3979 ( .INP(n4247), .Z(n4043) );
  NBUFFX2 U3980 ( .INP(n4246), .Z(n4044) );
  NBUFFX2 U3981 ( .INP(n4246), .Z(n4045) );
  NBUFFX2 U3982 ( .INP(n4246), .Z(n4046) );
  NBUFFX2 U3983 ( .INP(n4245), .Z(n4047) );
  NBUFFX2 U3984 ( .INP(n4245), .Z(n4048) );
  NBUFFX2 U3985 ( .INP(n4245), .Z(n4049) );
  NBUFFX2 U3986 ( .INP(n4244), .Z(n4050) );
  NBUFFX2 U3987 ( .INP(n4244), .Z(n4051) );
  NBUFFX2 U3988 ( .INP(n4244), .Z(n4052) );
  NBUFFX2 U3989 ( .INP(n4243), .Z(n4053) );
  NBUFFX2 U3990 ( .INP(n4243), .Z(n4054) );
  NBUFFX2 U3992 ( .INP(n4243), .Z(n4055) );
  NBUFFX2 U3993 ( .INP(n4242), .Z(n4056) );
  NBUFFX2 U3994 ( .INP(n4242), .Z(n4057) );
  NBUFFX2 U3995 ( .INP(n4242), .Z(n4058) );
  NBUFFX2 U3996 ( .INP(n4241), .Z(n4059) );
  NBUFFX2 U3997 ( .INP(n4241), .Z(n4060) );
  NBUFFX2 U3998 ( .INP(n4241), .Z(n4061) );
  NBUFFX2 U3999 ( .INP(n4240), .Z(n4062) );
  NBUFFX2 U4000 ( .INP(n4240), .Z(n4063) );
  NBUFFX2 U4001 ( .INP(n4240), .Z(n4064) );
  NBUFFX2 U4002 ( .INP(n4239), .Z(n4065) );
  NBUFFX2 U4003 ( .INP(n4239), .Z(n4066) );
  NBUFFX2 U4004 ( .INP(n4239), .Z(n4067) );
  NBUFFX2 U4005 ( .INP(n4238), .Z(n4068) );
  NBUFFX2 U4006 ( .INP(n4238), .Z(n4069) );
  NBUFFX2 U4007 ( .INP(n4238), .Z(n4070) );
  NBUFFX2 U4008 ( .INP(n4237), .Z(n4071) );
  NBUFFX2 U4009 ( .INP(n4237), .Z(n4072) );
  NBUFFX2 U4010 ( .INP(n4237), .Z(n4073) );
  NBUFFX2 U4011 ( .INP(n4236), .Z(n4074) );
  NBUFFX2 U4012 ( .INP(n4236), .Z(n4075) );
  NBUFFX2 U4013 ( .INP(n4236), .Z(n4076) );
  NBUFFX2 U4014 ( .INP(n4235), .Z(n4077) );
  NBUFFX2 U4015 ( .INP(n4235), .Z(n4078) );
  NBUFFX2 U4016 ( .INP(n4235), .Z(n4079) );
  NBUFFX2 U4017 ( .INP(n4234), .Z(n4080) );
  NBUFFX2 U4018 ( .INP(n4234), .Z(n4081) );
  NBUFFX2 U4019 ( .INP(n4234), .Z(n4082) );
  NBUFFX2 U4020 ( .INP(n4233), .Z(n4083) );
  NBUFFX2 U4021 ( .INP(n4233), .Z(n4084) );
  NBUFFX2 U4022 ( .INP(n4233), .Z(n4085) );
  NBUFFX2 U4023 ( .INP(n4232), .Z(n4086) );
  NBUFFX2 U4024 ( .INP(n4232), .Z(n4087) );
  NBUFFX2 U4025 ( .INP(n4232), .Z(n4088) );
  NBUFFX2 U4026 ( .INP(n4231), .Z(n4089) );
  NBUFFX2 U4027 ( .INP(n4231), .Z(n4090) );
  NBUFFX2 U4028 ( .INP(n4231), .Z(n4091) );
  NBUFFX2 U4029 ( .INP(n4230), .Z(n4092) );
  NBUFFX2 U4030 ( .INP(n4230), .Z(n4093) );
  NBUFFX2 U4031 ( .INP(n4230), .Z(n4094) );
  NBUFFX2 U4032 ( .INP(n4229), .Z(n4095) );
  NBUFFX2 U4033 ( .INP(n4229), .Z(n4096) );
  NBUFFX2 U4034 ( .INP(n4229), .Z(n4097) );
  NBUFFX2 U4035 ( .INP(n4228), .Z(n4098) );
  NBUFFX2 U4036 ( .INP(n4228), .Z(n4099) );
  NBUFFX2 U4037 ( .INP(n4228), .Z(n4100) );
  NBUFFX2 U4038 ( .INP(n4227), .Z(n4101) );
  NBUFFX2 U4039 ( .INP(n4227), .Z(n4102) );
  NBUFFX2 U4040 ( .INP(n4227), .Z(n4103) );
  NBUFFX2 U4041 ( .INP(n4226), .Z(n4104) );
  NBUFFX2 U4042 ( .INP(n4226), .Z(n4105) );
  NBUFFX2 U4043 ( .INP(n4226), .Z(n4106) );
  NBUFFX2 U4044 ( .INP(n4225), .Z(n4107) );
  NBUFFX2 U4045 ( .INP(n4225), .Z(n4108) );
  NBUFFX2 U4046 ( .INP(n4225), .Z(n4109) );
  NBUFFX2 U4047 ( .INP(n4224), .Z(n4110) );
  NBUFFX2 U4048 ( .INP(n4224), .Z(n4111) );
  NBUFFX2 U4049 ( .INP(n4224), .Z(n4112) );
  NBUFFX2 U4050 ( .INP(n4223), .Z(n4113) );
  NBUFFX2 U4051 ( .INP(n4223), .Z(n4114) );
  NBUFFX2 U4052 ( .INP(n4223), .Z(n4115) );
  NBUFFX2 U4053 ( .INP(n4222), .Z(n4116) );
  NBUFFX2 U4054 ( .INP(n4222), .Z(n4117) );
  NBUFFX2 U4055 ( .INP(n4222), .Z(n4118) );
  NBUFFX2 U4056 ( .INP(n4221), .Z(n4119) );
  NBUFFX2 U4057 ( .INP(n4221), .Z(n4120) );
  NBUFFX2 U4058 ( .INP(n4221), .Z(n4121) );
  NBUFFX2 U4059 ( .INP(n4220), .Z(n4122) );
  NBUFFX2 U4060 ( .INP(n4220), .Z(n4123) );
  NBUFFX2 U4061 ( .INP(n4220), .Z(n4124) );
  NBUFFX2 U4062 ( .INP(n4219), .Z(n4125) );
  NBUFFX2 U4063 ( .INP(n4219), .Z(n4126) );
  NBUFFX2 U4064 ( .INP(n4219), .Z(n4127) );
  NBUFFX2 U4065 ( .INP(n4218), .Z(n4128) );
  NBUFFX2 U4066 ( .INP(n4218), .Z(n4129) );
  NBUFFX2 U4067 ( .INP(n4218), .Z(n4130) );
  NBUFFX2 U4068 ( .INP(n4217), .Z(n4131) );
  NBUFFX2 U4069 ( .INP(n4217), .Z(n4132) );
  NBUFFX2 U4070 ( .INP(n4217), .Z(n4133) );
  NBUFFX2 U4071 ( .INP(n4216), .Z(n4134) );
  NBUFFX2 U4072 ( .INP(n4216), .Z(n4135) );
  NBUFFX2 U4073 ( .INP(n4216), .Z(n4136) );
  NBUFFX2 U4074 ( .INP(n4215), .Z(n4137) );
  NBUFFX2 U4075 ( .INP(n4215), .Z(n4138) );
  NBUFFX2 U4076 ( .INP(n4215), .Z(n4139) );
  NBUFFX2 U4077 ( .INP(n4214), .Z(n4140) );
  NBUFFX2 U4078 ( .INP(n4214), .Z(n4141) );
  NBUFFX2 U4079 ( .INP(n4214), .Z(n4142) );
  NBUFFX2 U4080 ( .INP(n4213), .Z(n4143) );
  NBUFFX2 U4081 ( .INP(n4213), .Z(n4144) );
  NBUFFX2 U4082 ( .INP(n4213), .Z(n4145) );
  NBUFFX2 U4083 ( .INP(n4212), .Z(n4146) );
  NBUFFX2 U4084 ( .INP(n4212), .Z(n4147) );
  NBUFFX2 U4085 ( .INP(n4212), .Z(n4148) );
  NBUFFX2 U4086 ( .INP(n4211), .Z(n4149) );
  NBUFFX2 U4087 ( .INP(n4211), .Z(n4150) );
  NBUFFX2 U4088 ( .INP(n4211), .Z(n4151) );
  NBUFFX2 U4089 ( .INP(n4210), .Z(n4152) );
  NBUFFX2 U4090 ( .INP(n4210), .Z(n4153) );
  NBUFFX2 U4091 ( .INP(n4210), .Z(n4154) );
  NBUFFX2 U4092 ( .INP(n4209), .Z(n4155) );
  NBUFFX2 U4093 ( .INP(n4209), .Z(n4156) );
  NBUFFX2 U4094 ( .INP(n4209), .Z(n4157) );
  NBUFFX2 U4095 ( .INP(n4208), .Z(n4158) );
  NBUFFX2 U4096 ( .INP(n4208), .Z(n4159) );
  NBUFFX2 U4097 ( .INP(n4208), .Z(n4160) );
  NBUFFX2 U4098 ( .INP(n4207), .Z(n4161) );
  NBUFFX2 U4099 ( .INP(n4207), .Z(n4162) );
  NBUFFX2 U4100 ( .INP(n4207), .Z(n4163) );
  NBUFFX2 U4101 ( .INP(n4206), .Z(n4164) );
  NBUFFX2 U4102 ( .INP(n4206), .Z(n4165) );
  NBUFFX2 U4103 ( .INP(n4206), .Z(n4166) );
  NBUFFX2 U4104 ( .INP(n4205), .Z(n4167) );
  NBUFFX2 U4105 ( .INP(n4205), .Z(n4168) );
  NBUFFX2 U4106 ( .INP(n4205), .Z(n4169) );
  NBUFFX2 U4107 ( .INP(n4204), .Z(n4170) );
  NBUFFX2 U4108 ( .INP(n4204), .Z(n4171) );
  NBUFFX2 U4109 ( .INP(n4204), .Z(n4172) );
  NBUFFX2 U4110 ( .INP(n4203), .Z(n4173) );
  NBUFFX2 U4111 ( .INP(n4203), .Z(n4174) );
  NBUFFX2 U4112 ( .INP(n4203), .Z(n4175) );
  NBUFFX2 U4113 ( .INP(n4202), .Z(n4176) );
  NBUFFX2 U4114 ( .INP(n4202), .Z(n4177) );
  NBUFFX2 U4115 ( .INP(n4202), .Z(n4178) );
  NBUFFX2 U4116 ( .INP(n4201), .Z(n4179) );
  NBUFFX2 U4117 ( .INP(n4201), .Z(n4180) );
  NBUFFX2 U4118 ( .INP(n4201), .Z(n4181) );
  NBUFFX2 U4119 ( .INP(n4200), .Z(n4182) );
  NBUFFX2 U4120 ( .INP(n4200), .Z(n4183) );
  NBUFFX2 U4121 ( .INP(n4200), .Z(n4184) );
  NBUFFX2 U4122 ( .INP(n4199), .Z(n4185) );
  NBUFFX2 U4123 ( .INP(n4199), .Z(n4186) );
  NBUFFX2 U4124 ( .INP(n4199), .Z(n4187) );
  NBUFFX2 U4125 ( .INP(n4198), .Z(n4188) );
  NBUFFX2 U4126 ( .INP(n4198), .Z(n4189) );
  NBUFFX2 U4127 ( .INP(n4198), .Z(n4190) );
  NBUFFX2 U4128 ( .INP(n4197), .Z(n4191) );
  NBUFFX2 U4129 ( .INP(n4197), .Z(n4192) );
  NBUFFX2 U4130 ( .INP(n4197), .Z(n4193) );
  NBUFFX2 U4131 ( .INP(n4196), .Z(n4194) );
  NBUFFX2 U4132 ( .INP(n4196), .Z(n4195) );
  NBUFFX2 U4133 ( .INP(n4325), .Z(n4196) );
  NBUFFX2 U4134 ( .INP(n4324), .Z(n4197) );
  NBUFFX2 U4135 ( .INP(n4324), .Z(n4198) );
  NBUFFX2 U4136 ( .INP(n4324), .Z(n4199) );
  NBUFFX2 U4137 ( .INP(n4323), .Z(n4200) );
  NBUFFX2 U4138 ( .INP(n4323), .Z(n4201) );
  NBUFFX2 U4139 ( .INP(n4323), .Z(n4202) );
  NBUFFX2 U4140 ( .INP(n4322), .Z(n4203) );
  NBUFFX2 U4141 ( .INP(n4322), .Z(n4204) );
  NBUFFX2 U4142 ( .INP(n4322), .Z(n4205) );
  NBUFFX2 U4143 ( .INP(n4321), .Z(n4206) );
  NBUFFX2 U4144 ( .INP(n4321), .Z(n4207) );
  NBUFFX2 U4145 ( .INP(n4321), .Z(n4208) );
  NBUFFX2 U4146 ( .INP(n4320), .Z(n4209) );
  NBUFFX2 U4147 ( .INP(n4320), .Z(n4210) );
  NBUFFX2 U4148 ( .INP(n4320), .Z(n4211) );
  NBUFFX2 U4149 ( .INP(n4319), .Z(n4212) );
  NBUFFX2 U4150 ( .INP(n4319), .Z(n4213) );
  NBUFFX2 U4151 ( .INP(n4319), .Z(n4214) );
  NBUFFX2 U4152 ( .INP(n4318), .Z(n4215) );
  NBUFFX2 U4153 ( .INP(n4318), .Z(n4216) );
  NBUFFX2 U4154 ( .INP(n4318), .Z(n4217) );
  NBUFFX2 U4155 ( .INP(n4317), .Z(n4218) );
  NBUFFX2 U4156 ( .INP(n4317), .Z(n4219) );
  NBUFFX2 U4157 ( .INP(n4317), .Z(n4220) );
  NBUFFX2 U4158 ( .INP(n4316), .Z(n4221) );
  NBUFFX2 U4159 ( .INP(n4316), .Z(n4222) );
  NBUFFX2 U4160 ( .INP(n4316), .Z(n4223) );
  NBUFFX2 U4161 ( .INP(n4315), .Z(n4224) );
  NBUFFX2 U4162 ( .INP(n4315), .Z(n4225) );
  NBUFFX2 U4163 ( .INP(n4315), .Z(n4226) );
  NBUFFX2 U4164 ( .INP(n4314), .Z(n4227) );
  NBUFFX2 U4165 ( .INP(n4314), .Z(n4228) );
  NBUFFX2 U4166 ( .INP(n4314), .Z(n4229) );
  NBUFFX2 U4167 ( .INP(n4313), .Z(n4230) );
  NBUFFX2 U4168 ( .INP(n4313), .Z(n4231) );
  NBUFFX2 U4169 ( .INP(n4313), .Z(n4232) );
  NBUFFX2 U4170 ( .INP(n4312), .Z(n4233) );
  NBUFFX2 U4171 ( .INP(n4312), .Z(n4234) );
  NBUFFX2 U4172 ( .INP(n4312), .Z(n4235) );
  NBUFFX2 U4173 ( .INP(n4311), .Z(n4236) );
  NBUFFX2 U4174 ( .INP(n4311), .Z(n4237) );
  NBUFFX2 U4175 ( .INP(n4311), .Z(n4238) );
  NBUFFX2 U4176 ( .INP(n4310), .Z(n4239) );
  NBUFFX2 U4177 ( .INP(n4310), .Z(n4240) );
  NBUFFX2 U4178 ( .INP(n4310), .Z(n4241) );
  NBUFFX2 U4179 ( .INP(n4309), .Z(n4242) );
  NBUFFX2 U4180 ( .INP(n4309), .Z(n4243) );
  NBUFFX2 U4181 ( .INP(n4309), .Z(n4244) );
  NBUFFX2 U4182 ( .INP(n4308), .Z(n4245) );
  NBUFFX2 U4183 ( .INP(n4308), .Z(n4246) );
  NBUFFX2 U4184 ( .INP(n4308), .Z(n4247) );
  NBUFFX2 U4185 ( .INP(n4307), .Z(n4248) );
  NBUFFX2 U4186 ( .INP(n4307), .Z(n4249) );
  NBUFFX2 U4187 ( .INP(n4307), .Z(n4250) );
  NBUFFX2 U4188 ( .INP(n4306), .Z(n4251) );
  NBUFFX2 U4189 ( .INP(n4306), .Z(n4252) );
  NBUFFX2 U4190 ( .INP(n4306), .Z(n4253) );
  NBUFFX2 U4191 ( .INP(n4305), .Z(n4254) );
  NBUFFX2 U4192 ( .INP(n4305), .Z(n4255) );
  NBUFFX2 U4193 ( .INP(n4305), .Z(n4256) );
  NBUFFX2 U4194 ( .INP(n4304), .Z(n4257) );
  NBUFFX2 U4195 ( .INP(n4304), .Z(n4258) );
  NBUFFX2 U4196 ( .INP(n4304), .Z(n4259) );
  NBUFFX2 U4197 ( .INP(n4303), .Z(n4260) );
  NBUFFX2 U4198 ( .INP(n4303), .Z(n4261) );
  NBUFFX2 U4199 ( .INP(n4303), .Z(n4262) );
  NBUFFX2 U4200 ( .INP(n4302), .Z(n4263) );
  NBUFFX2 U4201 ( .INP(n4302), .Z(n4264) );
  NBUFFX2 U4202 ( .INP(n4302), .Z(n4265) );
  NBUFFX2 U4203 ( .INP(n4301), .Z(n4266) );
  NBUFFX2 U4204 ( .INP(n4301), .Z(n4267) );
  NBUFFX2 U4205 ( .INP(n4301), .Z(n4268) );
  NBUFFX2 U4206 ( .INP(n4300), .Z(n4269) );
  NBUFFX2 U4207 ( .INP(n4300), .Z(n4270) );
  NBUFFX2 U4208 ( .INP(n4300), .Z(n4271) );
  NBUFFX2 U4209 ( .INP(n4299), .Z(n4272) );
  NBUFFX2 U4210 ( .INP(n4299), .Z(n4273) );
  NBUFFX2 U4211 ( .INP(n4299), .Z(n4274) );
  NBUFFX2 U4212 ( .INP(n4298), .Z(n4275) );
  NBUFFX2 U4213 ( .INP(n4298), .Z(n4276) );
  NBUFFX2 U4214 ( .INP(n4298), .Z(n4277) );
  NBUFFX2 U4215 ( .INP(n4297), .Z(n4278) );
  NBUFFX2 U4216 ( .INP(n4297), .Z(n4279) );
  NBUFFX2 U4217 ( .INP(n4297), .Z(n4280) );
  NBUFFX2 U4218 ( .INP(n4296), .Z(n4281) );
  NBUFFX2 U4219 ( .INP(n4296), .Z(n4282) );
  NBUFFX2 U4220 ( .INP(n4296), .Z(n4283) );
  NBUFFX2 U4221 ( .INP(n4295), .Z(n4284) );
  NBUFFX2 U4222 ( .INP(n4295), .Z(n4285) );
  NBUFFX2 U4223 ( .INP(n4295), .Z(n4286) );
  NBUFFX2 U4224 ( .INP(n4294), .Z(n4287) );
  NBUFFX2 U4225 ( .INP(n4294), .Z(n4288) );
  NBUFFX2 U4226 ( .INP(n4294), .Z(n4289) );
  NBUFFX2 U4227 ( .INP(n4293), .Z(n4290) );
  NBUFFX2 U4228 ( .INP(n4293), .Z(n4291) );
  NBUFFX2 U4229 ( .INP(n4293), .Z(n4292) );
  NBUFFX2 U4230 ( .INP(n4336), .Z(n4293) );
  NBUFFX2 U4231 ( .INP(n4336), .Z(n4294) );
  NBUFFX2 U4232 ( .INP(n4336), .Z(n4295) );
  NBUFFX2 U4233 ( .INP(n4335), .Z(n4296) );
  NBUFFX2 U4234 ( .INP(n4335), .Z(n4297) );
  NBUFFX2 U4235 ( .INP(n4335), .Z(n4298) );
  NBUFFX2 U4236 ( .INP(n4334), .Z(n4299) );
  NBUFFX2 U4237 ( .INP(n4334), .Z(n4300) );
  NBUFFX2 U4238 ( .INP(n4334), .Z(n4301) );
  NBUFFX2 U4239 ( .INP(n4333), .Z(n4302) );
  NBUFFX2 U4240 ( .INP(n4333), .Z(n4303) );
  NBUFFX2 U4241 ( .INP(n4333), .Z(n4304) );
  NBUFFX2 U4242 ( .INP(n4332), .Z(n4305) );
  NBUFFX2 U4243 ( .INP(n4332), .Z(n4306) );
  NBUFFX2 U4244 ( .INP(n4332), .Z(n4307) );
  NBUFFX2 U4245 ( .INP(n4331), .Z(n4308) );
  NBUFFX2 U4246 ( .INP(n4331), .Z(n4309) );
  NBUFFX2 U4247 ( .INP(n4331), .Z(n4310) );
  NBUFFX2 U4248 ( .INP(n4330), .Z(n4311) );
  NBUFFX2 U4249 ( .INP(n4330), .Z(n4312) );
  NBUFFX2 U4250 ( .INP(n4330), .Z(n4313) );
  NBUFFX2 U4251 ( .INP(n4329), .Z(n4314) );
  NBUFFX2 U4252 ( .INP(n4329), .Z(n4315) );
  NBUFFX2 U4253 ( .INP(n4329), .Z(n4316) );
  NBUFFX2 U4254 ( .INP(n4328), .Z(n4317) );
  NBUFFX2 U4255 ( .INP(n4328), .Z(n4318) );
  NBUFFX2 U4256 ( .INP(n4328), .Z(n4319) );
  NBUFFX2 U4257 ( .INP(n4327), .Z(n4320) );
  NBUFFX2 U4258 ( .INP(n4327), .Z(n4321) );
  NBUFFX2 U4259 ( .INP(n4327), .Z(n4322) );
  NBUFFX2 U4260 ( .INP(n4326), .Z(n4323) );
  NBUFFX2 U4261 ( .INP(n4326), .Z(n4324) );
  NBUFFX2 U4262 ( .INP(n4326), .Z(n4325) );
  NBUFFX2 U4263 ( .INP(n4340), .Z(n4326) );
  NBUFFX2 U4264 ( .INP(n4340), .Z(n4327) );
  NBUFFX2 U4265 ( .INP(n4339), .Z(n4328) );
  NBUFFX2 U4266 ( .INP(n4339), .Z(n4329) );
  NBUFFX2 U4267 ( .INP(n4339), .Z(n4330) );
  NBUFFX2 U4268 ( .INP(n4338), .Z(n4331) );
  NBUFFX2 U4269 ( .INP(n4338), .Z(n4332) );
  NBUFFX2 U4270 ( .INP(n4338), .Z(n4333) );
  NBUFFX2 U4271 ( .INP(n4337), .Z(n4334) );
  NBUFFX2 U4272 ( .INP(n4337), .Z(n4335) );
  NBUFFX2 U4273 ( .INP(n4337), .Z(n4336) );
  NBUFFX2 U4274 ( .INP(test_se), .Z(n4337) );
  NBUFFX2 U4275 ( .INP(test_se), .Z(n4338) );
  NBUFFX2 U4276 ( .INP(test_se), .Z(n4339) );
  NBUFFX2 U4277 ( .INP(test_se), .Z(n4340) );
  NBUFFX2 U4278 ( .INP(n4403), .Z(n4341) );
  NBUFFX2 U4279 ( .INP(n4403), .Z(n4342) );
  NBUFFX2 U4280 ( .INP(n4402), .Z(n4343) );
  NBUFFX2 U4281 ( .INP(n4402), .Z(n4344) );
  NBUFFX2 U4282 ( .INP(n4402), .Z(n4345) );
  NBUFFX2 U4283 ( .INP(n4401), .Z(n4346) );
  NBUFFX2 U4284 ( .INP(n4401), .Z(n4347) );
  NBUFFX2 U4285 ( .INP(n4401), .Z(n4348) );
  NBUFFX2 U4286 ( .INP(n4400), .Z(n4349) );
  NBUFFX2 U4287 ( .INP(n4400), .Z(n4350) );
  NBUFFX2 U4288 ( .INP(n4400), .Z(n4351) );
  NBUFFX2 U4289 ( .INP(n4399), .Z(n4352) );
  NBUFFX2 U4290 ( .INP(n4399), .Z(n4353) );
  NBUFFX2 U4291 ( .INP(n4399), .Z(n4354) );
  NBUFFX2 U4292 ( .INP(n4398), .Z(n4355) );
  NBUFFX2 U4293 ( .INP(n4398), .Z(n4356) );
  NBUFFX2 U4294 ( .INP(n4398), .Z(n4357) );
  NBUFFX2 U4295 ( .INP(n4397), .Z(n4358) );
  NBUFFX2 U4296 ( .INP(n4397), .Z(n4359) );
  NBUFFX2 U4297 ( .INP(n4397), .Z(n4360) );
  NBUFFX2 U4298 ( .INP(n4396), .Z(n4361) );
  NBUFFX2 U4299 ( .INP(n4396), .Z(n4362) );
  NBUFFX2 U4300 ( .INP(n4396), .Z(n4363) );
  NBUFFX2 U4301 ( .INP(n4395), .Z(n4364) );
  NBUFFX2 U4302 ( .INP(n4395), .Z(n4365) );
  NBUFFX2 U4303 ( .INP(n4395), .Z(n4366) );
  NBUFFX2 U4304 ( .INP(n4394), .Z(n4367) );
  NBUFFX2 U4305 ( .INP(n4394), .Z(n4368) );
  NBUFFX2 U4306 ( .INP(n4394), .Z(n4369) );
  NBUFFX2 U4307 ( .INP(n4393), .Z(n4370) );
  NBUFFX2 U4308 ( .INP(n4393), .Z(n4371) );
  NBUFFX2 U4309 ( .INP(n4393), .Z(n4372) );
  NBUFFX2 U4310 ( .INP(n4392), .Z(n4373) );
  NBUFFX2 U4311 ( .INP(n4392), .Z(n4374) );
  NBUFFX2 U4312 ( .INP(n4392), .Z(n4375) );
  NBUFFX2 U4313 ( .INP(n4391), .Z(n4376) );
  NBUFFX2 U4314 ( .INP(n4391), .Z(n4377) );
  NBUFFX2 U4315 ( .INP(n4391), .Z(n4378) );
  NBUFFX2 U4316 ( .INP(n4390), .Z(n4379) );
  NBUFFX2 U4317 ( .INP(n4390), .Z(n4380) );
  NBUFFX2 U4318 ( .INP(n4390), .Z(n4381) );
  NBUFFX2 U4319 ( .INP(n4389), .Z(n4382) );
  NBUFFX2 U4320 ( .INP(n4389), .Z(n4383) );
  NBUFFX2 U4321 ( .INP(n4389), .Z(n4384) );
  NBUFFX2 U4322 ( .INP(n4388), .Z(n4385) );
  NBUFFX2 U4323 ( .INP(n4388), .Z(n4386) );
  NBUFFX2 U4324 ( .INP(n4388), .Z(n4387) );
  NBUFFX2 U4325 ( .INP(n4409), .Z(n4388) );
  NBUFFX2 U4326 ( .INP(n4408), .Z(n4389) );
  NBUFFX2 U4327 ( .INP(n4408), .Z(n4390) );
  NBUFFX2 U4328 ( .INP(n4408), .Z(n4391) );
  NBUFFX2 U4329 ( .INP(n4407), .Z(n4392) );
  NBUFFX2 U4330 ( .INP(n4407), .Z(n4393) );
  NBUFFX2 U4331 ( .INP(n4407), .Z(n4394) );
  NBUFFX2 U4332 ( .INP(n4406), .Z(n4395) );
  NBUFFX2 U4333 ( .INP(n4406), .Z(n4396) );
  NBUFFX2 U4334 ( .INP(n4406), .Z(n4397) );
  NBUFFX2 U4335 ( .INP(n4405), .Z(n4398) );
  NBUFFX2 U4336 ( .INP(n4405), .Z(n4399) );
  NBUFFX2 U4337 ( .INP(n4405), .Z(n4400) );
  NBUFFX2 U4338 ( .INP(n4404), .Z(n4401) );
  NBUFFX2 U4339 ( .INP(n4404), .Z(n4402) );
  NBUFFX2 U4340 ( .INP(n4404), .Z(n4403) );
  NBUFFX2 U4341 ( .INP(RESET), .Z(n4404) );
  NBUFFX2 U4342 ( .INP(RESET), .Z(n4405) );
  NBUFFX2 U4343 ( .INP(RESET), .Z(n4406) );
  NBUFFX2 U4344 ( .INP(RESET), .Z(n4407) );
  NBUFFX2 U4345 ( .INP(RESET), .Z(n4408) );
  NBUFFX2 U4346 ( .INP(RESET), .Z(n4409) );
  INVX0 U4347 ( .INP(n4341), .ZN(n4410) );
  INVX0 U4348 ( .INP(n4341), .ZN(n4411) );
  INVX0 U4349 ( .INP(n4341), .ZN(n4412) );
  INVX0 U4350 ( .INP(n4341), .ZN(n4413) );
  INVX0 U4351 ( .INP(n4341), .ZN(n4414) );
  INVX0 U4352 ( .INP(n4341), .ZN(n4415) );
  INVX0 U4353 ( .INP(n4341), .ZN(n4416) );
  INVX0 U4354 ( .INP(n4341), .ZN(n4417) );
  INVX0 U4355 ( .INP(n4342), .ZN(n4418) );
  INVX0 U4356 ( .INP(n4342), .ZN(n4419) );
  INVX0 U4357 ( .INP(n4342), .ZN(n4420) );
  INVX0 U4358 ( .INP(n4342), .ZN(n4421) );
  INVX0 U4359 ( .INP(n4342), .ZN(n4422) );
  INVX0 U4360 ( .INP(n4342), .ZN(n4423) );
  INVX0 U4361 ( .INP(n4342), .ZN(n4424) );
  INVX0 U4362 ( .INP(n4342), .ZN(n4425) );
  INVX0 U4363 ( .INP(n4343), .ZN(n4426) );
  INVX0 U4364 ( .INP(n4343), .ZN(n4427) );
  INVX0 U4365 ( .INP(n4343), .ZN(n4428) );
  INVX0 U4366 ( .INP(n4343), .ZN(n4429) );
  INVX0 U4367 ( .INP(n4343), .ZN(n4430) );
  INVX0 U4368 ( .INP(n4343), .ZN(n4431) );
  INVX0 U4369 ( .INP(n4343), .ZN(n4432) );
  INVX0 U4370 ( .INP(n4343), .ZN(n4433) );
  INVX0 U4371 ( .INP(n4344), .ZN(n4434) );
  INVX0 U4372 ( .INP(n4344), .ZN(n4435) );
  INVX0 U4373 ( .INP(n4344), .ZN(n4436) );
  INVX0 U4374 ( .INP(n4344), .ZN(n4437) );
  INVX0 U4375 ( .INP(n4344), .ZN(n4438) );
  INVX0 U4376 ( .INP(n4344), .ZN(n4439) );
  INVX0 U4377 ( .INP(n4344), .ZN(n4440) );
  INVX0 U4378 ( .INP(n4344), .ZN(n4441) );
  INVX0 U4379 ( .INP(n4345), .ZN(n4442) );
  INVX0 U4380 ( .INP(n4345), .ZN(n4443) );
  INVX0 U4381 ( .INP(n4345), .ZN(n4444) );
  INVX0 U4382 ( .INP(n4345), .ZN(n4445) );
  INVX0 U4383 ( .INP(n4345), .ZN(n4446) );
  INVX0 U4384 ( .INP(n4345), .ZN(n4447) );
  INVX0 U4385 ( .INP(n4345), .ZN(n4448) );
  INVX0 U4386 ( .INP(n4345), .ZN(n4449) );
  INVX0 U4387 ( .INP(n4346), .ZN(n4450) );
  INVX0 U4388 ( .INP(n4346), .ZN(n4451) );
  INVX0 U4389 ( .INP(n4346), .ZN(n4452) );
  INVX0 U4390 ( .INP(n4346), .ZN(n4453) );
  INVX0 U4391 ( .INP(n4346), .ZN(n4454) );
  INVX0 U4392 ( .INP(n4346), .ZN(n4455) );
  INVX0 U4393 ( .INP(n4346), .ZN(n4456) );
  INVX0 U4394 ( .INP(n4347), .ZN(n4457) );
  INVX0 U4395 ( .INP(n4347), .ZN(n4458) );
  INVX0 U4396 ( .INP(n4347), .ZN(n4459) );
  INVX0 U4397 ( .INP(n4347), .ZN(n4460) );
  INVX0 U4398 ( .INP(n4347), .ZN(n4461) );
  INVX0 U4399 ( .INP(n4347), .ZN(n4462) );
  INVX0 U4400 ( .INP(n4347), .ZN(n4463) );
  INVX0 U4401 ( .INP(n4347), .ZN(n4464) );
  INVX0 U4402 ( .INP(n4348), .ZN(n4465) );
  INVX0 U4403 ( .INP(n4348), .ZN(n4466) );
  INVX0 U4404 ( .INP(n4348), .ZN(n4467) );
  INVX0 U4405 ( .INP(n4348), .ZN(n4468) );
  INVX0 U4406 ( .INP(n4348), .ZN(n4469) );
  INVX0 U4407 ( .INP(n4348), .ZN(n4470) );
  INVX0 U4408 ( .INP(n4348), .ZN(n4471) );
  INVX0 U4409 ( .INP(n4348), .ZN(n4472) );
  INVX0 U4410 ( .INP(n4349), .ZN(n4473) );
  INVX0 U4411 ( .INP(n4349), .ZN(n4474) );
  INVX0 U4412 ( .INP(n4349), .ZN(n4475) );
  INVX0 U4413 ( .INP(n4349), .ZN(n4476) );
  INVX0 U4414 ( .INP(n4349), .ZN(n4477) );
  INVX0 U4415 ( .INP(n4349), .ZN(n4478) );
  INVX0 U4416 ( .INP(n4349), .ZN(n4479) );
  INVX0 U4417 ( .INP(n4349), .ZN(n4480) );
  INVX0 U4418 ( .INP(n4350), .ZN(n4481) );
  INVX0 U4419 ( .INP(n4350), .ZN(n4482) );
  INVX0 U4420 ( .INP(n4350), .ZN(n4483) );
  INVX0 U4421 ( .INP(n4350), .ZN(n4484) );
  INVX0 U4422 ( .INP(n4350), .ZN(n4485) );
  INVX0 U4423 ( .INP(n4350), .ZN(n4486) );
  INVX0 U4424 ( .INP(n4350), .ZN(n4487) );
  INVX0 U4425 ( .INP(n4350), .ZN(n4488) );
  INVX0 U4426 ( .INP(n4351), .ZN(n4489) );
  INVX0 U4427 ( .INP(n4351), .ZN(n4490) );
  NBUFFX2 U4428 ( .INP(n4673), .Z(n4635) );
  NBUFFX2 U4429 ( .INP(n4673), .Z(n4636) );
  NBUFFX2 U4430 ( .INP(n4672), .Z(n4637) );
  NBUFFX2 U4431 ( .INP(n4672), .Z(n4638) );
  NBUFFX2 U4432 ( .INP(n4672), .Z(n4639) );
  NBUFFX2 U4433 ( .INP(n4671), .Z(n4640) );
  NBUFFX2 U4434 ( .INP(n4671), .Z(n4641) );
  NBUFFX2 U4435 ( .INP(n4671), .Z(n4642) );
  NBUFFX2 U4436 ( .INP(n4670), .Z(n4643) );
  NBUFFX2 U4437 ( .INP(n4670), .Z(n4644) );
  NBUFFX2 U4438 ( .INP(n4670), .Z(n4645) );
  NBUFFX2 U4439 ( .INP(n4669), .Z(n4646) );
  NBUFFX2 U4440 ( .INP(n4669), .Z(n4647) );
  NBUFFX2 U4441 ( .INP(n4669), .Z(n4648) );
  NBUFFX2 U4442 ( .INP(n4668), .Z(n4649) );
  NBUFFX2 U4443 ( .INP(n4668), .Z(n4650) );
  NBUFFX2 U4444 ( .INP(n4668), .Z(n4651) );
  NBUFFX2 U4445 ( .INP(n4667), .Z(n4652) );
  NBUFFX2 U4446 ( .INP(n4667), .Z(n4653) );
  NBUFFX2 U4447 ( .INP(n4667), .Z(n4654) );
  NBUFFX2 U4448 ( .INP(n4666), .Z(n4655) );
  NBUFFX2 U4449 ( .INP(n4666), .Z(n4656) );
  NBUFFX2 U4450 ( .INP(n4666), .Z(n4657) );
  NBUFFX2 U4451 ( .INP(n4665), .Z(n4658) );
  NBUFFX2 U4452 ( .INP(n4665), .Z(n4659) );
  NBUFFX2 U4453 ( .INP(n4665), .Z(n4660) );
  NBUFFX2 U4454 ( .INP(n4664), .Z(n4661) );
  NBUFFX2 U4455 ( .INP(n4664), .Z(n4662) );
  NBUFFX2 U4456 ( .INP(n4664), .Z(n4663) );
  NBUFFX2 U4457 ( .INP(CK), .Z(n4664) );
  NBUFFX2 U4458 ( .INP(CK), .Z(n4665) );
  NBUFFX2 U4459 ( .INP(n4673), .Z(n4666) );
  NBUFFX2 U4460 ( .INP(CK), .Z(n4667) );
  NBUFFX2 U4461 ( .INP(n4669), .Z(n4668) );
  NBUFFX2 U4462 ( .INP(CK), .Z(n4669) );
  NBUFFX2 U4463 ( .INP(n4664), .Z(n4670) );
  NBUFFX2 U4464 ( .INP(n4665), .Z(n4671) );
  NBUFFX2 U4465 ( .INP(n4667), .Z(n4672) );
  NBUFFX2 U4466 ( .INP(n4504), .Z(n4673) );
  AND2X1 U4467 ( .IN1(n4385), .IN2(n3518), .Q(n3278) );
  INVX0 U4468 ( .INP(n4674), .ZN(WX9789) );
  OR2X1 U4469 ( .IN1(n4410), .IN2(n7078), .Q(n4674) );
  INVX0 U4470 ( .INP(n4675), .ZN(WX9787) );
  OR2X1 U4471 ( .IN1(n4423), .IN2(n7079), .Q(n4675) );
  INVX0 U4472 ( .INP(n4676), .ZN(WX9785) );
  OR2X1 U4473 ( .IN1(n4423), .IN2(n7080), .Q(n4676) );
  INVX0 U4474 ( .INP(n4677), .ZN(WX9783) );
  OR2X1 U4475 ( .IN1(n4422), .IN2(n7081), .Q(n4677) );
  AND2X1 U4476 ( .IN1(test_so80), .IN2(n4364), .Q(WX9781) );
  INVX0 U4477 ( .INP(n4678), .ZN(WX9779) );
  OR2X1 U4478 ( .IN1(n4422), .IN2(n7083), .Q(n4678) );
  INVX0 U4479 ( .INP(n4679), .ZN(WX9777) );
  OR2X1 U4480 ( .IN1(n4422), .IN2(n7084), .Q(n4679) );
  INVX0 U4481 ( .INP(n4680), .ZN(WX9775) );
  OR2X1 U4482 ( .IN1(n4422), .IN2(n7085), .Q(n4680) );
  INVX0 U4483 ( .INP(n4681), .ZN(WX9773) );
  OR2X1 U4484 ( .IN1(n4422), .IN2(n7086), .Q(n4681) );
  INVX0 U4485 ( .INP(n4682), .ZN(WX9771) );
  OR2X1 U4486 ( .IN1(n4422), .IN2(n7087), .Q(n4682) );
  INVX0 U4487 ( .INP(n4683), .ZN(WX9769) );
  OR2X1 U4488 ( .IN1(n4422), .IN2(n7088), .Q(n4683) );
  INVX0 U4489 ( .INP(n4684), .ZN(WX9767) );
  OR2X1 U4490 ( .IN1(n4422), .IN2(n7089), .Q(n4684) );
  INVX0 U4491 ( .INP(n4685), .ZN(WX9765) );
  OR2X1 U4492 ( .IN1(n4422), .IN2(n7090), .Q(n4685) );
  INVX0 U4493 ( .INP(n4686), .ZN(WX9763) );
  OR2X1 U4494 ( .IN1(n4422), .IN2(n7091), .Q(n4686) );
  INVX0 U4495 ( .INP(n4687), .ZN(WX9761) );
  OR2X1 U4496 ( .IN1(n4422), .IN2(n7092), .Q(n4687) );
  INVX0 U4497 ( .INP(n4688), .ZN(WX9759) );
  OR2X1 U4498 ( .IN1(n4422), .IN2(n7093), .Q(n4688) );
  OR4X1 U4499 ( .IN1(n4689), .IN2(n4690), .IN3(n4691), .IN4(n4692), .Q(WX9757)
         );
  AND2X1 U4500 ( .IN1(n3630), .IN2(n4693), .Q(n4692) );
  AND2X1 U4501 ( .IN1(n3543), .IN2(n4695), .Q(n4691) );
  AND2X1 U4502 ( .IN1(n3589), .IN2(CRC_OUT_2_0), .Q(n4690) );
  AND2X1 U4503 ( .IN1(n436), .IN2(n3584), .Q(n4689) );
  INVX0 U4504 ( .INP(n4696), .ZN(n436) );
  OR2X1 U4505 ( .IN1(n4422), .IN2(n3817), .Q(n4696) );
  OR4X1 U4506 ( .IN1(n4697), .IN2(n4698), .IN3(n4699), .IN4(n4700), .Q(WX9755)
         );
  AND2X1 U4507 ( .IN1(n3640), .IN2(n4701), .Q(n4700) );
  AND2X1 U4508 ( .IN1(n4702), .IN2(n3528), .Q(n4699) );
  AND2X1 U4509 ( .IN1(n3604), .IN2(CRC_OUT_2_1), .Q(n4698) );
  AND2X1 U4510 ( .IN1(n435), .IN2(n3584), .Q(n4697) );
  INVX0 U4511 ( .INP(n4703), .ZN(n435) );
  OR2X1 U4512 ( .IN1(n4421), .IN2(n3818), .Q(n4703) );
  OR4X1 U4513 ( .IN1(n4704), .IN2(n4705), .IN3(n4706), .IN4(n4707), .Q(WX9753)
         );
  AND2X1 U4514 ( .IN1(n4708), .IN2(n3624), .Q(n4707) );
  AND2X1 U4515 ( .IN1(n3543), .IN2(n4709), .Q(n4706) );
  AND2X1 U4516 ( .IN1(test_so87), .IN2(n3587), .Q(n4705) );
  AND2X1 U4517 ( .IN1(n434), .IN2(n3584), .Q(n4704) );
  INVX0 U4518 ( .INP(n4710), .ZN(n434) );
  OR2X1 U4519 ( .IN1(n4421), .IN2(n3819), .Q(n4710) );
  OR4X1 U4520 ( .IN1(n4711), .IN2(n4712), .IN3(n4713), .IN4(n4714), .Q(WX9751)
         );
  AND2X1 U4521 ( .IN1(n3634), .IN2(n4715), .Q(n4714) );
  AND2X1 U4522 ( .IN1(n4716), .IN2(n3528), .Q(n4713) );
  AND2X1 U4523 ( .IN1(n3599), .IN2(CRC_OUT_2_3), .Q(n4712) );
  AND2X1 U4524 ( .IN1(n433), .IN2(n3583), .Q(n4711) );
  INVX0 U4525 ( .INP(n4717), .ZN(n433) );
  OR2X1 U4526 ( .IN1(n4421), .IN2(n3820), .Q(n4717) );
  OR4X1 U4527 ( .IN1(n4718), .IN2(n4719), .IN3(n4720), .IN4(n4721), .Q(WX9749)
         );
  AND2X1 U4528 ( .IN1(n4722), .IN2(n3624), .Q(n4721) );
  AND2X1 U4529 ( .IN1(n3543), .IN2(n4723), .Q(n4720) );
  AND2X1 U4530 ( .IN1(n3599), .IN2(CRC_OUT_2_4), .Q(n4719) );
  AND2X1 U4531 ( .IN1(n432), .IN2(n3583), .Q(n4718) );
  INVX0 U4532 ( .INP(n4724), .ZN(n432) );
  OR2X1 U4533 ( .IN1(n4421), .IN2(n3821), .Q(n4724) );
  OR4X1 U4534 ( .IN1(n4725), .IN2(n4726), .IN3(n4727), .IN4(n4728), .Q(WX9747)
         );
  AND2X1 U4535 ( .IN1(n3634), .IN2(n4729), .Q(n4728) );
  AND2X1 U4536 ( .IN1(n3543), .IN2(n4730), .Q(n4727) );
  AND2X1 U4537 ( .IN1(n3599), .IN2(CRC_OUT_2_5), .Q(n4726) );
  AND2X1 U4538 ( .IN1(n431), .IN2(n3583), .Q(n4725) );
  INVX0 U4539 ( .INP(n4731), .ZN(n431) );
  OR2X1 U4540 ( .IN1(n4421), .IN2(n3822), .Q(n4731) );
  OR4X1 U4541 ( .IN1(n4732), .IN2(n4733), .IN3(n4734), .IN4(n4735), .Q(WX9745)
         );
  AND2X1 U4542 ( .IN1(n4736), .IN2(n3626), .Q(n4735) );
  AND2X1 U4543 ( .IN1(n3543), .IN2(n4737), .Q(n4734) );
  AND2X1 U4544 ( .IN1(n3599), .IN2(CRC_OUT_2_6), .Q(n4733) );
  AND2X1 U4545 ( .IN1(n430), .IN2(n3583), .Q(n4732) );
  INVX0 U4546 ( .INP(n4738), .ZN(n430) );
  OR2X1 U4547 ( .IN1(n4421), .IN2(n3823), .Q(n4738) );
  OR4X1 U4548 ( .IN1(n4739), .IN2(n4740), .IN3(n4741), .IN4(n4742), .Q(WX9743)
         );
  AND2X1 U4549 ( .IN1(n3634), .IN2(n4743), .Q(n4742) );
  AND2X1 U4550 ( .IN1(n3543), .IN2(n4744), .Q(n4741) );
  AND2X1 U4551 ( .IN1(n3599), .IN2(CRC_OUT_2_7), .Q(n4740) );
  AND2X1 U4552 ( .IN1(n429), .IN2(n3583), .Q(n4739) );
  INVX0 U4553 ( .INP(n4745), .ZN(n429) );
  OR2X1 U4554 ( .IN1(n4421), .IN2(n3824), .Q(n4745) );
  OR4X1 U4555 ( .IN1(n4746), .IN2(n4747), .IN3(n4748), .IN4(n4749), .Q(WX9741)
         );
  AND2X1 U4556 ( .IN1(n4750), .IN2(n3626), .Q(n4749) );
  AND2X1 U4557 ( .IN1(n3543), .IN2(n4751), .Q(n4748) );
  AND2X1 U4558 ( .IN1(n3600), .IN2(CRC_OUT_2_8), .Q(n4747) );
  AND2X1 U4559 ( .IN1(n428), .IN2(n3583), .Q(n4746) );
  INVX0 U4560 ( .INP(n4752), .ZN(n428) );
  OR2X1 U4561 ( .IN1(n4421), .IN2(n3825), .Q(n4752) );
  OR4X1 U4562 ( .IN1(n4753), .IN2(n4754), .IN3(n4755), .IN4(n4756), .Q(WX9739)
         );
  AND2X1 U4563 ( .IN1(n3634), .IN2(n4757), .Q(n4756) );
  AND2X1 U4564 ( .IN1(n3543), .IN2(n4758), .Q(n4755) );
  AND2X1 U4565 ( .IN1(n3600), .IN2(CRC_OUT_2_9), .Q(n4754) );
  AND2X1 U4566 ( .IN1(n427), .IN2(n3583), .Q(n4753) );
  INVX0 U4567 ( .INP(n4759), .ZN(n427) );
  OR2X1 U4568 ( .IN1(n4421), .IN2(n3826), .Q(n4759) );
  OR4X1 U4569 ( .IN1(n4760), .IN2(n4761), .IN3(n4762), .IN4(n4763), .Q(WX9737)
         );
  AND2X1 U4570 ( .IN1(n3634), .IN2(n4764), .Q(n4763) );
  AND2X1 U4571 ( .IN1(n3543), .IN2(n4765), .Q(n4762) );
  AND2X1 U4572 ( .IN1(n3600), .IN2(CRC_OUT_2_10), .Q(n4761) );
  AND2X1 U4573 ( .IN1(n426), .IN2(n3583), .Q(n4760) );
  INVX0 U4574 ( .INP(n4766), .ZN(n426) );
  OR2X1 U4575 ( .IN1(n4421), .IN2(n3827), .Q(n4766) );
  OR4X1 U4576 ( .IN1(n4767), .IN2(n4768), .IN3(n4769), .IN4(n4770), .Q(WX9735)
         );
  AND2X1 U4577 ( .IN1(n3634), .IN2(n4771), .Q(n4770) );
  AND2X1 U4578 ( .IN1(n3543), .IN2(n4772), .Q(n4769) );
  AND2X1 U4579 ( .IN1(n3600), .IN2(CRC_OUT_2_11), .Q(n4768) );
  AND2X1 U4580 ( .IN1(n425), .IN2(n3583), .Q(n4767) );
  INVX0 U4581 ( .INP(n4773), .ZN(n425) );
  OR2X1 U4582 ( .IN1(n4421), .IN2(n3828), .Q(n4773) );
  OR4X1 U4583 ( .IN1(n4774), .IN2(n4775), .IN3(n4776), .IN4(n4777), .Q(WX9733)
         );
  AND2X1 U4584 ( .IN1(n3634), .IN2(n4778), .Q(n4777) );
  AND2X1 U4585 ( .IN1(n3543), .IN2(n4779), .Q(n4776) );
  AND2X1 U4586 ( .IN1(n3600), .IN2(CRC_OUT_2_12), .Q(n4775) );
  AND2X1 U4587 ( .IN1(n424), .IN2(n3583), .Q(n4774) );
  INVX0 U4588 ( .INP(n4780), .ZN(n424) );
  OR2X1 U4589 ( .IN1(n4421), .IN2(n3829), .Q(n4780) );
  OR4X1 U4590 ( .IN1(n4781), .IN2(n4782), .IN3(n4783), .IN4(n4784), .Q(WX9731)
         );
  AND2X1 U4591 ( .IN1(n3634), .IN2(n4785), .Q(n4784) );
  AND2X1 U4592 ( .IN1(n3543), .IN2(n4786), .Q(n4783) );
  AND2X1 U4593 ( .IN1(n3600), .IN2(CRC_OUT_2_13), .Q(n4782) );
  AND2X1 U4594 ( .IN1(n423), .IN2(n3583), .Q(n4781) );
  INVX0 U4595 ( .INP(n4787), .ZN(n423) );
  OR2X1 U4596 ( .IN1(n4421), .IN2(n3830), .Q(n4787) );
  OR4X1 U4597 ( .IN1(n4788), .IN2(n4789), .IN3(n4790), .IN4(n4791), .Q(WX9729)
         );
  AND2X1 U4598 ( .IN1(n3634), .IN2(n4792), .Q(n4791) );
  AND2X1 U4599 ( .IN1(n4793), .IN2(n3530), .Q(n4790) );
  AND2X1 U4600 ( .IN1(n3600), .IN2(CRC_OUT_2_14), .Q(n4789) );
  AND2X1 U4601 ( .IN1(n422), .IN2(n3583), .Q(n4788) );
  INVX0 U4602 ( .INP(n4794), .ZN(n422) );
  OR2X1 U4603 ( .IN1(n4420), .IN2(n3831), .Q(n4794) );
  OR4X1 U4604 ( .IN1(n4795), .IN2(n4796), .IN3(n4797), .IN4(n4798), .Q(WX9727)
         );
  AND2X1 U4605 ( .IN1(n3634), .IN2(n4799), .Q(n4798) );
  AND2X1 U4606 ( .IN1(n3542), .IN2(n4800), .Q(n4797) );
  AND2X1 U4607 ( .IN1(n3600), .IN2(CRC_OUT_2_15), .Q(n4796) );
  AND2X1 U4608 ( .IN1(n421), .IN2(n3582), .Q(n4795) );
  INVX0 U4609 ( .INP(n4801), .ZN(n421) );
  OR2X1 U4610 ( .IN1(n4420), .IN2(n3832), .Q(n4801) );
  OR4X1 U4611 ( .IN1(n4802), .IN2(n4803), .IN3(n4804), .IN4(n4805), .Q(WX9725)
         );
  AND2X1 U4612 ( .IN1(n3634), .IN2(n4806), .Q(n4805) );
  AND2X1 U4613 ( .IN1(n4807), .IN2(n3530), .Q(n4804) );
  AND2X1 U4614 ( .IN1(n3600), .IN2(CRC_OUT_2_16), .Q(n4803) );
  AND2X1 U4615 ( .IN1(n420), .IN2(n3582), .Q(n4802) );
  INVX0 U4616 ( .INP(n4808), .ZN(n420) );
  OR2X1 U4617 ( .IN1(n4420), .IN2(n3833), .Q(n4808) );
  OR4X1 U4618 ( .IN1(n4809), .IN2(n4810), .IN3(n4811), .IN4(n4812), .Q(WX9723)
         );
  AND2X1 U4619 ( .IN1(n3636), .IN2(n4813), .Q(n4812) );
  AND2X1 U4620 ( .IN1(n3542), .IN2(n4814), .Q(n4811) );
  AND2X1 U4621 ( .IN1(n3600), .IN2(CRC_OUT_2_17), .Q(n4810) );
  AND2X1 U4622 ( .IN1(n419), .IN2(n3582), .Q(n4809) );
  INVX0 U4623 ( .INP(n4815), .ZN(n419) );
  OR2X1 U4624 ( .IN1(n4420), .IN2(n3834), .Q(n4815) );
  OR4X1 U4625 ( .IN1(n4816), .IN2(n4817), .IN3(n4818), .IN4(n4819), .Q(WX9721)
         );
  AND2X1 U4626 ( .IN1(n3636), .IN2(n4820), .Q(n4819) );
  AND2X1 U4627 ( .IN1(n4821), .IN2(n3530), .Q(n4818) );
  AND2X1 U4628 ( .IN1(n3600), .IN2(CRC_OUT_2_18), .Q(n4817) );
  AND2X1 U4629 ( .IN1(n418), .IN2(n3582), .Q(n4816) );
  INVX0 U4630 ( .INP(n4822), .ZN(n418) );
  OR2X1 U4631 ( .IN1(n4420), .IN2(n3835), .Q(n4822) );
  OR4X1 U4632 ( .IN1(n4823), .IN2(n4824), .IN3(n4825), .IN4(n4826), .Q(WX9719)
         );
  AND2X1 U4633 ( .IN1(n4827), .IN2(n3628), .Q(n4826) );
  AND2X1 U4634 ( .IN1(n3542), .IN2(n4828), .Q(n4825) );
  AND2X1 U4635 ( .IN1(test_so88), .IN2(n3587), .Q(n4824) );
  AND2X1 U4636 ( .IN1(n417), .IN2(n3582), .Q(n4823) );
  INVX0 U4637 ( .INP(n4829), .ZN(n417) );
  OR2X1 U4638 ( .IN1(n4420), .IN2(n3836), .Q(n4829) );
  OR4X1 U4639 ( .IN1(n4830), .IN2(n4831), .IN3(n4832), .IN4(n4833), .Q(WX9717)
         );
  AND2X1 U4640 ( .IN1(n3636), .IN2(n4834), .Q(n4833) );
  AND2X1 U4641 ( .IN1(n4835), .IN2(n3530), .Q(n4832) );
  AND2X1 U4642 ( .IN1(n3600), .IN2(CRC_OUT_2_20), .Q(n4831) );
  AND2X1 U4643 ( .IN1(n416), .IN2(n3582), .Q(n4830) );
  INVX0 U4644 ( .INP(n4836), .ZN(n416) );
  OR2X1 U4645 ( .IN1(n4420), .IN2(n3837), .Q(n4836) );
  OR4X1 U4646 ( .IN1(n4837), .IN2(n4838), .IN3(n4839), .IN4(n4840), .Q(WX9715)
         );
  AND2X1 U4647 ( .IN1(n4841), .IN2(n3627), .Q(n4840) );
  AND2X1 U4648 ( .IN1(n3542), .IN2(n4842), .Q(n4839) );
  AND2X1 U4649 ( .IN1(n3600), .IN2(CRC_OUT_2_21), .Q(n4838) );
  AND2X1 U4650 ( .IN1(n415), .IN2(n3582), .Q(n4837) );
  INVX0 U4651 ( .INP(n4843), .ZN(n415) );
  OR2X1 U4652 ( .IN1(n4420), .IN2(n3838), .Q(n4843) );
  OR4X1 U4653 ( .IN1(n4844), .IN2(n4845), .IN3(n4846), .IN4(n4847), .Q(WX9713)
         );
  AND2X1 U4654 ( .IN1(n3636), .IN2(n4848), .Q(n4847) );
  AND2X1 U4655 ( .IN1(n3542), .IN2(n4849), .Q(n4846) );
  AND2X1 U4656 ( .IN1(n3601), .IN2(CRC_OUT_2_22), .Q(n4845) );
  AND2X1 U4657 ( .IN1(n414), .IN2(n3582), .Q(n4844) );
  INVX0 U4658 ( .INP(n4850), .ZN(n414) );
  OR2X1 U4659 ( .IN1(n4420), .IN2(n3839), .Q(n4850) );
  OR4X1 U4660 ( .IN1(n4851), .IN2(n4852), .IN3(n4853), .IN4(n4854), .Q(WX9711)
         );
  AND2X1 U4661 ( .IN1(n4855), .IN2(n3628), .Q(n4854) );
  AND2X1 U4662 ( .IN1(n3542), .IN2(n4856), .Q(n4853) );
  AND2X1 U4663 ( .IN1(n3601), .IN2(CRC_OUT_2_23), .Q(n4852) );
  AND2X1 U4664 ( .IN1(n413), .IN2(n3582), .Q(n4851) );
  INVX0 U4665 ( .INP(n4857), .ZN(n413) );
  OR2X1 U4666 ( .IN1(n4420), .IN2(n3840), .Q(n4857) );
  OR4X1 U4667 ( .IN1(n4858), .IN2(n4859), .IN3(n4860), .IN4(n4861), .Q(WX9709)
         );
  AND2X1 U4668 ( .IN1(n3636), .IN2(n4862), .Q(n4861) );
  AND2X1 U4669 ( .IN1(n3542), .IN2(n4863), .Q(n4860) );
  AND2X1 U4670 ( .IN1(n3601), .IN2(CRC_OUT_2_24), .Q(n4859) );
  AND2X1 U4671 ( .IN1(n412), .IN2(n3582), .Q(n4858) );
  INVX0 U4672 ( .INP(n4864), .ZN(n412) );
  OR2X1 U4673 ( .IN1(n4420), .IN2(n3841), .Q(n4864) );
  OR4X1 U4674 ( .IN1(n4865), .IN2(n4866), .IN3(n4867), .IN4(n4868), .Q(WX9707)
         );
  AND2X1 U4675 ( .IN1(n4869), .IN2(n3627), .Q(n4868) );
  AND2X1 U4676 ( .IN1(n3542), .IN2(n4870), .Q(n4867) );
  AND2X1 U4677 ( .IN1(n3601), .IN2(CRC_OUT_2_25), .Q(n4866) );
  AND2X1 U4678 ( .IN1(n411), .IN2(n3582), .Q(n4865) );
  INVX0 U4679 ( .INP(n4871), .ZN(n411) );
  OR2X1 U4680 ( .IN1(n4420), .IN2(n3842), .Q(n4871) );
  OR4X1 U4681 ( .IN1(n4872), .IN2(n4873), .IN3(n4874), .IN4(n4875), .Q(WX9705)
         );
  AND2X1 U4682 ( .IN1(n3636), .IN2(n4876), .Q(n4875) );
  AND2X1 U4683 ( .IN1(n3542), .IN2(n4877), .Q(n4874) );
  AND2X1 U4684 ( .IN1(n3601), .IN2(CRC_OUT_2_26), .Q(n4873) );
  AND2X1 U4685 ( .IN1(n410), .IN2(n3582), .Q(n4872) );
  INVX0 U4686 ( .INP(n4878), .ZN(n410) );
  OR2X1 U4687 ( .IN1(n4420), .IN2(n3843), .Q(n4878) );
  OR4X1 U4688 ( .IN1(n4879), .IN2(n4880), .IN3(n4881), .IN4(n4882), .Q(WX9703)
         );
  AND2X1 U4689 ( .IN1(n3636), .IN2(n4883), .Q(n4882) );
  AND2X1 U4690 ( .IN1(n3542), .IN2(n4884), .Q(n4881) );
  AND2X1 U4691 ( .IN1(n3601), .IN2(CRC_OUT_2_27), .Q(n4880) );
  AND2X1 U4692 ( .IN1(n409), .IN2(n3581), .Q(n4879) );
  INVX0 U4693 ( .INP(n4885), .ZN(n409) );
  OR2X1 U4694 ( .IN1(n4419), .IN2(n3844), .Q(n4885) );
  OR4X1 U4695 ( .IN1(n4886), .IN2(n4887), .IN3(n4888), .IN4(n4889), .Q(WX9701)
         );
  AND2X1 U4696 ( .IN1(n3636), .IN2(n4890), .Q(n4889) );
  AND2X1 U4697 ( .IN1(n3542), .IN2(n4891), .Q(n4888) );
  AND2X1 U4698 ( .IN1(n3601), .IN2(CRC_OUT_2_28), .Q(n4887) );
  AND2X1 U4699 ( .IN1(n408), .IN2(n3581), .Q(n4886) );
  INVX0 U4700 ( .INP(n4892), .ZN(n408) );
  OR2X1 U4701 ( .IN1(n4419), .IN2(n3845), .Q(n4892) );
  OR4X1 U4702 ( .IN1(n4893), .IN2(n4894), .IN3(n4895), .IN4(n4896), .Q(WX9699)
         );
  AND2X1 U4703 ( .IN1(n3636), .IN2(n4897), .Q(n4896) );
  AND2X1 U4704 ( .IN1(n3542), .IN2(n4898), .Q(n4895) );
  AND2X1 U4705 ( .IN1(n3601), .IN2(CRC_OUT_2_29), .Q(n4894) );
  AND2X1 U4706 ( .IN1(n407), .IN2(n3581), .Q(n4893) );
  INVX0 U4707 ( .INP(n4899), .ZN(n407) );
  OR2X1 U4708 ( .IN1(n4419), .IN2(n3846), .Q(n4899) );
  OR4X1 U4709 ( .IN1(n4900), .IN2(n4901), .IN3(n4902), .IN4(n4903), .Q(WX9697)
         );
  AND2X1 U4710 ( .IN1(n3636), .IN2(n4904), .Q(n4903) );
  AND2X1 U4711 ( .IN1(n3542), .IN2(n4905), .Q(n4902) );
  AND2X1 U4712 ( .IN1(n3601), .IN2(CRC_OUT_2_30), .Q(n4901) );
  AND2X1 U4713 ( .IN1(n406), .IN2(n3581), .Q(n4900) );
  INVX0 U4714 ( .INP(n4906), .ZN(n406) );
  OR2X1 U4715 ( .IN1(n4419), .IN2(n3847), .Q(n4906) );
  OR4X1 U4716 ( .IN1(n4907), .IN2(n4908), .IN3(n4909), .IN4(n4910), .Q(WX9695)
         );
  AND2X1 U4717 ( .IN1(n3636), .IN2(n4911), .Q(n4910) );
  AND2X1 U4718 ( .IN1(n4912), .IN2(n3532), .Q(n4909) );
  AND2X1 U4719 ( .IN1(n2245), .IN2(WX9536), .Q(n4908) );
  AND2X1 U4720 ( .IN1(n3601), .IN2(CRC_OUT_2_31), .Q(n4907) );
  AND2X1 U4721 ( .IN1(n3508), .IN2(n4364), .Q(WX9597) );
  AND2X1 U4722 ( .IN1(n4913), .IN2(n4364), .Q(WX9084) );
  XOR2X1 U4723 ( .IN1(CRC_OUT_3_30), .IN2(n3254), .Q(n4913) );
  AND2X1 U4724 ( .IN1(n4914), .IN2(n4364), .Q(WX9082) );
  XOR2X1 U4725 ( .IN1(CRC_OUT_3_29), .IN2(n3255), .Q(n4914) );
  AND2X1 U4726 ( .IN1(n4915), .IN2(n4364), .Q(WX9080) );
  XOR2X1 U4727 ( .IN1(CRC_OUT_3_28), .IN2(n3256), .Q(n4915) );
  AND2X1 U4728 ( .IN1(n4916), .IN2(n4364), .Q(WX9078) );
  XOR2X1 U4729 ( .IN1(CRC_OUT_3_27), .IN2(n3257), .Q(n4916) );
  AND2X1 U4730 ( .IN1(n4917), .IN2(n4364), .Q(WX9076) );
  XOR2X1 U4731 ( .IN1(CRC_OUT_3_26), .IN2(n3258), .Q(n4917) );
  AND2X1 U4732 ( .IN1(n4918), .IN2(n4364), .Q(WX9074) );
  XOR2X1 U4733 ( .IN1(test_so74), .IN2(DFF_1337_n1), .Q(n4918) );
  AND2X1 U4734 ( .IN1(n4919), .IN2(n4364), .Q(WX9072) );
  XOR2X1 U4735 ( .IN1(test_so77), .IN2(n3259), .Q(n4919) );
  AND2X1 U4736 ( .IN1(n4920), .IN2(n4363), .Q(WX9070) );
  XOR2X1 U4737 ( .IN1(CRC_OUT_3_23), .IN2(n3260), .Q(n4920) );
  AND2X1 U4738 ( .IN1(n4921), .IN2(n4363), .Q(WX9068) );
  XOR2X1 U4739 ( .IN1(CRC_OUT_3_22), .IN2(n3261), .Q(n4921) );
  AND2X1 U4740 ( .IN1(n4922), .IN2(n4363), .Q(WX9066) );
  XOR2X1 U4741 ( .IN1(CRC_OUT_3_21), .IN2(n3262), .Q(n4922) );
  AND2X1 U4742 ( .IN1(n4923), .IN2(n4363), .Q(WX9064) );
  XOR2X1 U4743 ( .IN1(CRC_OUT_3_20), .IN2(n3263), .Q(n4923) );
  AND2X1 U4744 ( .IN1(n4924), .IN2(n4363), .Q(WX9062) );
  XOR2X1 U4745 ( .IN1(CRC_OUT_3_19), .IN2(n3264), .Q(n4924) );
  AND2X1 U4746 ( .IN1(n4925), .IN2(n4363), .Q(WX9060) );
  XOR2X1 U4747 ( .IN1(CRC_OUT_3_18), .IN2(n3265), .Q(n4925) );
  AND2X1 U4748 ( .IN1(n4926), .IN2(n4363), .Q(WX9058) );
  XOR2X1 U4749 ( .IN1(CRC_OUT_3_17), .IN2(n3266), .Q(n4926) );
  AND2X1 U4750 ( .IN1(n4927), .IN2(n4363), .Q(WX9056) );
  XOR2X1 U4751 ( .IN1(CRC_OUT_3_16), .IN2(n3267), .Q(n4927) );
  AND2X1 U4752 ( .IN1(n4928), .IN2(n4363), .Q(WX9054) );
  XOR3X1 U4753 ( .IN1(n3179), .IN2(DFF_1343_n1), .IN3(DFF_1327_n1), .Q(n4928)
         );
  AND2X1 U4754 ( .IN1(n4929), .IN2(n4362), .Q(WX9052) );
  XOR2X1 U4755 ( .IN1(CRC_OUT_3_14), .IN2(n3268), .Q(n4929) );
  AND2X1 U4756 ( .IN1(n4930), .IN2(n4362), .Q(WX9050) );
  XOR2X1 U4757 ( .IN1(CRC_OUT_3_13), .IN2(n3269), .Q(n4930) );
  AND2X1 U4758 ( .IN1(n4931), .IN2(n4362), .Q(WX9048) );
  XOR2X1 U4759 ( .IN1(CRC_OUT_3_12), .IN2(n3270), .Q(n4931) );
  AND2X1 U4760 ( .IN1(n4932), .IN2(n4362), .Q(WX9046) );
  XOR2X1 U4761 ( .IN1(CRC_OUT_3_11), .IN2(n3271), .Q(n4932) );
  AND2X1 U4762 ( .IN1(n4933), .IN2(n4362), .Q(WX9044) );
  XOR3X1 U4763 ( .IN1(n3180), .IN2(DFF_1343_n1), .IN3(DFF_1322_n1), .Q(n4933)
         );
  AND2X1 U4764 ( .IN1(n4934), .IN2(n4362), .Q(WX9042) );
  XOR2X1 U4765 ( .IN1(CRC_OUT_3_9), .IN2(n3272), .Q(n4934) );
  AND2X1 U4766 ( .IN1(n4935), .IN2(n4362), .Q(WX9040) );
  XOR2X1 U4767 ( .IN1(test_so75), .IN2(DFF_1320_n1), .Q(n4935) );
  AND2X1 U4768 ( .IN1(n4936), .IN2(n4362), .Q(WX9038) );
  XOR2X1 U4769 ( .IN1(test_so76), .IN2(n3273), .Q(n4936) );
  AND2X1 U4770 ( .IN1(n4937), .IN2(n4362), .Q(WX9036) );
  XOR2X1 U4771 ( .IN1(CRC_OUT_3_6), .IN2(n3274), .Q(n4937) );
  AND2X1 U4772 ( .IN1(n4938), .IN2(n4361), .Q(WX9034) );
  XOR2X1 U4773 ( .IN1(CRC_OUT_3_5), .IN2(n3275), .Q(n4938) );
  AND2X1 U4774 ( .IN1(n4939), .IN2(n4361), .Q(WX9032) );
  XOR2X1 U4775 ( .IN1(CRC_OUT_3_4), .IN2(n3276), .Q(n4939) );
  AND2X1 U4776 ( .IN1(n4940), .IN2(n4361), .Q(WX9030) );
  XOR3X1 U4777 ( .IN1(n3181), .IN2(DFF_1343_n1), .IN3(DFF_1315_n1), .Q(n4940)
         );
  AND2X1 U4778 ( .IN1(n4941), .IN2(n4361), .Q(WX9028) );
  XOR2X1 U4779 ( .IN1(CRC_OUT_3_2), .IN2(n3277), .Q(n4941) );
  AND2X1 U4780 ( .IN1(n4942), .IN2(n4361), .Q(WX9026) );
  XOR2X1 U4781 ( .IN1(CRC_OUT_3_1), .IN2(n3279), .Q(n4942) );
  AND2X1 U4782 ( .IN1(n4943), .IN2(n4361), .Q(WX9024) );
  XOR2X1 U4783 ( .IN1(CRC_OUT_3_0), .IN2(n3280), .Q(n4943) );
  AND2X1 U4784 ( .IN1(n4944), .IN2(n4361), .Q(WX9022) );
  XOR2X1 U4785 ( .IN1(n3196), .IN2(CRC_OUT_3_31), .Q(n4944) );
  INVX0 U4786 ( .INP(n4945), .ZN(WX8496) );
  OR2X1 U4787 ( .IN1(n4419), .IN2(n7106), .Q(n4945) );
  INVX0 U4788 ( .INP(n4946), .ZN(WX8494) );
  OR2X1 U4789 ( .IN1(n4419), .IN2(n7107), .Q(n4946) );
  INVX0 U4790 ( .INP(n4947), .ZN(WX8492) );
  OR2X1 U4791 ( .IN1(n4419), .IN2(n7108), .Q(n4947) );
  INVX0 U4792 ( .INP(n4948), .ZN(WX8490) );
  OR2X1 U4793 ( .IN1(n4419), .IN2(n7109), .Q(n4948) );
  INVX0 U4794 ( .INP(n4949), .ZN(WX8488) );
  OR2X1 U4795 ( .IN1(n4419), .IN2(n7110), .Q(n4949) );
  INVX0 U4796 ( .INP(n4950), .ZN(WX8486) );
  OR2X1 U4797 ( .IN1(n4419), .IN2(n7111), .Q(n4950) );
  INVX0 U4798 ( .INP(n4951), .ZN(WX8484) );
  OR2X1 U4799 ( .IN1(n4419), .IN2(n7112), .Q(n4951) );
  INVX0 U4800 ( .INP(n4952), .ZN(WX8482) );
  OR2X1 U4801 ( .IN1(n4419), .IN2(n7113), .Q(n4952) );
  INVX0 U4802 ( .INP(n4953), .ZN(WX8480) );
  OR2X1 U4803 ( .IN1(n4419), .IN2(n7114), .Q(n4953) );
  INVX0 U4804 ( .INP(n4954), .ZN(WX8478) );
  OR2X1 U4805 ( .IN1(n4418), .IN2(n7115), .Q(n4954) );
  INVX0 U4806 ( .INP(n4955), .ZN(WX8476) );
  OR2X1 U4807 ( .IN1(n4418), .IN2(n7116), .Q(n4955) );
  INVX0 U4808 ( .INP(n4956), .ZN(WX8474) );
  OR2X1 U4809 ( .IN1(n4418), .IN2(n7117), .Q(n4956) );
  INVX0 U4810 ( .INP(n4957), .ZN(WX8472) );
  OR2X1 U4811 ( .IN1(n4418), .IN2(n7118), .Q(n4957) );
  INVX0 U4812 ( .INP(n4958), .ZN(WX8470) );
  OR2X1 U4813 ( .IN1(n4418), .IN2(n7119), .Q(n4958) );
  INVX0 U4814 ( .INP(n4959), .ZN(WX8468) );
  OR2X1 U4815 ( .IN1(n4418), .IN2(n7120), .Q(n4959) );
  INVX0 U4816 ( .INP(n4960), .ZN(WX8466) );
  OR2X1 U4817 ( .IN1(n4418), .IN2(n7121), .Q(n4960) );
  OR4X1 U4818 ( .IN1(n4961), .IN2(n4962), .IN3(n4963), .IN4(n4964), .Q(WX8464)
         );
  AND2X1 U4819 ( .IN1(n3541), .IN2(n4965), .Q(n4964) );
  AND2X1 U4820 ( .IN1(n3636), .IN2(n4695), .Q(n4963) );
  XNOR3X1 U4821 ( .IN1(n3195), .IN2(n3073), .IN3(n4966), .Q(n4695) );
  XOR2X1 U4822 ( .IN1(WX9822), .IN2(n7065), .Q(n4966) );
  AND2X1 U4823 ( .IN1(n3601), .IN2(CRC_OUT_3_0), .Q(n4962) );
  AND2X1 U4824 ( .IN1(n374), .IN2(n3581), .Q(n4961) );
  INVX0 U4825 ( .INP(n4967), .ZN(n374) );
  OR2X1 U4826 ( .IN1(n4418), .IN2(n3848), .Q(n4967) );
  OR4X1 U4827 ( .IN1(n4968), .IN2(n4969), .IN3(n4970), .IN4(n4971), .Q(WX8462)
         );
  AND2X1 U4828 ( .IN1(n3541), .IN2(n4972), .Q(n4971) );
  AND2X1 U4829 ( .IN1(n4702), .IN2(n3626), .Q(n4970) );
  XOR3X1 U4830 ( .IN1(n3253), .IN2(n3074), .IN3(n4973), .Q(n4702) );
  XOR2X1 U4831 ( .IN1(WX9756), .IN2(test_so83), .Q(n4973) );
  AND2X1 U4832 ( .IN1(n3601), .IN2(CRC_OUT_3_1), .Q(n4969) );
  AND2X1 U4833 ( .IN1(n373), .IN2(n3581), .Q(n4968) );
  INVX0 U4834 ( .INP(n4974), .ZN(n373) );
  OR2X1 U4835 ( .IN1(n4418), .IN2(n3849), .Q(n4974) );
  OR4X1 U4836 ( .IN1(n4975), .IN2(n4976), .IN3(n4977), .IN4(n4978), .Q(WX8460)
         );
  AND2X1 U4837 ( .IN1(n3541), .IN2(n4979), .Q(n4978) );
  AND2X1 U4838 ( .IN1(n3636), .IN2(n4709), .Q(n4977) );
  XNOR3X1 U4839 ( .IN1(n3252), .IN2(n3075), .IN3(n4980), .Q(n4709) );
  XOR2X1 U4840 ( .IN1(WX9818), .IN2(n7066), .Q(n4980) );
  AND2X1 U4841 ( .IN1(n3601), .IN2(CRC_OUT_3_2), .Q(n4976) );
  AND2X1 U4842 ( .IN1(n372), .IN2(n3581), .Q(n4975) );
  INVX0 U4843 ( .INP(n4981), .ZN(n372) );
  OR2X1 U4844 ( .IN1(n4418), .IN2(n3850), .Q(n4981) );
  OR4X1 U4845 ( .IN1(n4982), .IN2(n4983), .IN3(n4984), .IN4(n4985), .Q(WX8458)
         );
  AND2X1 U4846 ( .IN1(n3541), .IN2(n4986), .Q(n4985) );
  AND2X1 U4847 ( .IN1(n4716), .IN2(n3624), .Q(n4984) );
  XOR3X1 U4848 ( .IN1(n3569), .IN2(n3251), .IN3(n4987), .Q(n4716) );
  XOR2X1 U4849 ( .IN1(WX9880), .IN2(test_so81), .Q(n4987) );
  AND2X1 U4850 ( .IN1(n3602), .IN2(CRC_OUT_3_3), .Q(n4983) );
  AND2X1 U4851 ( .IN1(n371), .IN2(n3581), .Q(n4982) );
  INVX0 U4852 ( .INP(n4988), .ZN(n371) );
  OR2X1 U4853 ( .IN1(n4418), .IN2(n3851), .Q(n4988) );
  OR4X1 U4854 ( .IN1(n4989), .IN2(n4990), .IN3(n4991), .IN4(n4992), .Q(WX8456)
         );
  AND2X1 U4855 ( .IN1(n3541), .IN2(n4993), .Q(n4992) );
  AND2X1 U4856 ( .IN1(n3637), .IN2(n4723), .Q(n4991) );
  XNOR3X1 U4857 ( .IN1(n3178), .IN2(n3076), .IN3(n4994), .Q(n4723) );
  XOR2X1 U4858 ( .IN1(WX9814), .IN2(n7067), .Q(n4994) );
  AND2X1 U4859 ( .IN1(n3602), .IN2(CRC_OUT_3_4), .Q(n4990) );
  AND2X1 U4860 ( .IN1(n370), .IN2(n3581), .Q(n4989) );
  INVX0 U4861 ( .INP(n4995), .ZN(n370) );
  OR2X1 U4862 ( .IN1(n4418), .IN2(n3852), .Q(n4995) );
  OR4X1 U4863 ( .IN1(n4996), .IN2(n4997), .IN3(n4998), .IN4(n4999), .Q(WX8454)
         );
  AND2X1 U4864 ( .IN1(n3541), .IN2(n5000), .Q(n4999) );
  AND2X1 U4865 ( .IN1(n3637), .IN2(n4730), .Q(n4998) );
  XNOR3X1 U4866 ( .IN1(n3250), .IN2(n3077), .IN3(n5001), .Q(n4730) );
  XOR2X1 U4867 ( .IN1(WX9812), .IN2(n7068), .Q(n5001) );
  AND2X1 U4868 ( .IN1(n3602), .IN2(CRC_OUT_3_5), .Q(n4997) );
  AND2X1 U4869 ( .IN1(n369), .IN2(n3581), .Q(n4996) );
  INVX0 U4870 ( .INP(n5002), .ZN(n369) );
  OR2X1 U4871 ( .IN1(n4418), .IN2(n3853), .Q(n5002) );
  OR4X1 U4872 ( .IN1(n5003), .IN2(n5004), .IN3(n5005), .IN4(n5006), .Q(WX8452)
         );
  AND2X1 U4873 ( .IN1(n3541), .IN2(n5007), .Q(n5006) );
  AND2X1 U4874 ( .IN1(n3637), .IN2(n4737), .Q(n5005) );
  XNOR3X1 U4875 ( .IN1(n3249), .IN2(n3078), .IN3(n5008), .Q(n4737) );
  XOR2X1 U4876 ( .IN1(WX9810), .IN2(n7069), .Q(n5008) );
  AND2X1 U4877 ( .IN1(n3602), .IN2(CRC_OUT_3_6), .Q(n5004) );
  AND2X1 U4878 ( .IN1(n368), .IN2(n3581), .Q(n5003) );
  INVX0 U4879 ( .INP(n5009), .ZN(n368) );
  OR2X1 U4880 ( .IN1(n4417), .IN2(n3854), .Q(n5009) );
  OR4X1 U4881 ( .IN1(n5010), .IN2(n5011), .IN3(n5012), .IN4(n5013), .Q(WX8450)
         );
  AND2X1 U4882 ( .IN1(n3541), .IN2(n5014), .Q(n5013) );
  AND2X1 U4883 ( .IN1(n3637), .IN2(n4744), .Q(n5012) );
  XNOR3X1 U4884 ( .IN1(n3248), .IN2(n3079), .IN3(n5015), .Q(n4744) );
  XOR2X1 U4885 ( .IN1(WX9808), .IN2(n7070), .Q(n5015) );
  AND2X1 U4886 ( .IN1(test_so76), .IN2(n3588), .Q(n5011) );
  AND2X1 U4887 ( .IN1(n367), .IN2(n3581), .Q(n5010) );
  INVX0 U4888 ( .INP(n5016), .ZN(n367) );
  OR2X1 U4889 ( .IN1(n4417), .IN2(n3855), .Q(n5016) );
  OR4X1 U4890 ( .IN1(n5017), .IN2(n5018), .IN3(n5019), .IN4(n5020), .Q(WX8448)
         );
  AND2X1 U4891 ( .IN1(n3541), .IN2(n5021), .Q(n5020) );
  AND2X1 U4892 ( .IN1(n3637), .IN2(n4751), .Q(n5019) );
  XNOR3X1 U4893 ( .IN1(n3247), .IN2(n3080), .IN3(n5022), .Q(n4751) );
  XOR2X1 U4894 ( .IN1(WX9806), .IN2(n7071), .Q(n5022) );
  AND2X1 U4895 ( .IN1(n3602), .IN2(CRC_OUT_3_8), .Q(n5018) );
  AND2X1 U4896 ( .IN1(n366), .IN2(n3580), .Q(n5017) );
  INVX0 U4897 ( .INP(n5023), .ZN(n366) );
  OR2X1 U4898 ( .IN1(n4417), .IN2(n3856), .Q(n5023) );
  OR4X1 U4899 ( .IN1(n5024), .IN2(n5025), .IN3(n5026), .IN4(n5027), .Q(WX8446)
         );
  AND2X1 U4900 ( .IN1(n5028), .IN2(n3533), .Q(n5027) );
  AND2X1 U4901 ( .IN1(n3637), .IN2(n4758), .Q(n5026) );
  XNOR3X1 U4902 ( .IN1(n3246), .IN2(n3081), .IN3(n5029), .Q(n4758) );
  XOR2X1 U4903 ( .IN1(WX9804), .IN2(n7072), .Q(n5029) );
  AND2X1 U4904 ( .IN1(n3602), .IN2(CRC_OUT_3_9), .Q(n5025) );
  AND2X1 U4905 ( .IN1(n365), .IN2(n3580), .Q(n5024) );
  INVX0 U4906 ( .INP(n5030), .ZN(n365) );
  OR2X1 U4907 ( .IN1(n4417), .IN2(n3857), .Q(n5030) );
  OR4X1 U4908 ( .IN1(n5031), .IN2(n5032), .IN3(n5033), .IN4(n5034), .Q(WX8444)
         );
  AND2X1 U4909 ( .IN1(n3541), .IN2(n5035), .Q(n5034) );
  AND2X1 U4910 ( .IN1(n3637), .IN2(n4765), .Q(n5033) );
  XNOR3X1 U4911 ( .IN1(n3245), .IN2(n3082), .IN3(n5036), .Q(n4765) );
  XOR2X1 U4912 ( .IN1(WX9802), .IN2(n7073), .Q(n5036) );
  AND2X1 U4913 ( .IN1(n3602), .IN2(CRC_OUT_3_10), .Q(n5032) );
  AND2X1 U4914 ( .IN1(n364), .IN2(n3580), .Q(n5031) );
  INVX0 U4915 ( .INP(n5037), .ZN(n364) );
  OR2X1 U4916 ( .IN1(n4417), .IN2(n3858), .Q(n5037) );
  OR4X1 U4917 ( .IN1(n5038), .IN2(n5039), .IN3(n5040), .IN4(n5041), .Q(WX8442)
         );
  AND2X1 U4918 ( .IN1(n5042), .IN2(n3533), .Q(n5041) );
  AND2X1 U4919 ( .IN1(n3637), .IN2(n4772), .Q(n5040) );
  XNOR3X1 U4920 ( .IN1(n3177), .IN2(n3083), .IN3(n5043), .Q(n4772) );
  XOR2X1 U4921 ( .IN1(WX9800), .IN2(n7074), .Q(n5043) );
  AND2X1 U4922 ( .IN1(n3602), .IN2(CRC_OUT_3_11), .Q(n5039) );
  AND2X1 U4923 ( .IN1(n363), .IN2(n3580), .Q(n5038) );
  INVX0 U4924 ( .INP(n5044), .ZN(n363) );
  OR2X1 U4925 ( .IN1(n4417), .IN2(n3859), .Q(n5044) );
  OR4X1 U4926 ( .IN1(n5045), .IN2(n5046), .IN3(n5047), .IN4(n5048), .Q(WX8440)
         );
  AND2X1 U4927 ( .IN1(n3541), .IN2(n5049), .Q(n5048) );
  AND2X1 U4928 ( .IN1(n3637), .IN2(n4779), .Q(n5047) );
  XNOR3X1 U4929 ( .IN1(n3244), .IN2(n3084), .IN3(n5050), .Q(n4779) );
  XOR2X1 U4930 ( .IN1(WX9798), .IN2(n7075), .Q(n5050) );
  AND2X1 U4931 ( .IN1(n3602), .IN2(CRC_OUT_3_12), .Q(n5046) );
  AND2X1 U4932 ( .IN1(n362), .IN2(n3580), .Q(n5045) );
  INVX0 U4933 ( .INP(n5051), .ZN(n362) );
  OR2X1 U4934 ( .IN1(n4417), .IN2(n3860), .Q(n5051) );
  OR4X1 U4935 ( .IN1(n5052), .IN2(n5053), .IN3(n5054), .IN4(n5055), .Q(WX8438)
         );
  AND2X1 U4936 ( .IN1(n5056), .IN2(n3533), .Q(n5055) );
  AND2X1 U4937 ( .IN1(n3637), .IN2(n4786), .Q(n5054) );
  XNOR3X1 U4938 ( .IN1(n3243), .IN2(n3085), .IN3(n5057), .Q(n4786) );
  XOR2X1 U4939 ( .IN1(WX9796), .IN2(n7076), .Q(n5057) );
  AND2X1 U4940 ( .IN1(n3602), .IN2(CRC_OUT_3_13), .Q(n5053) );
  AND2X1 U4941 ( .IN1(n361), .IN2(n3580), .Q(n5052) );
  INVX0 U4942 ( .INP(n5058), .ZN(n361) );
  OR2X1 U4943 ( .IN1(n4417), .IN2(n3861), .Q(n5058) );
  OR4X1 U4944 ( .IN1(n5059), .IN2(n5060), .IN3(n5061), .IN4(n5062), .Q(WX8436)
         );
  AND2X1 U4945 ( .IN1(n3541), .IN2(n5063), .Q(n5062) );
  AND2X1 U4946 ( .IN1(n4793), .IN2(n3624), .Q(n5061) );
  XOR3X1 U4947 ( .IN1(n3591), .IN2(n3086), .IN3(n5064), .Q(n4793) );
  XOR2X1 U4948 ( .IN1(WX9730), .IN2(test_so86), .Q(n5064) );
  AND2X1 U4949 ( .IN1(n3602), .IN2(CRC_OUT_3_14), .Q(n5060) );
  AND2X1 U4950 ( .IN1(n360), .IN2(n3580), .Q(n5059) );
  INVX0 U4951 ( .INP(n5065), .ZN(n360) );
  OR2X1 U4952 ( .IN1(n4417), .IN2(n3862), .Q(n5065) );
  OR4X1 U4953 ( .IN1(n5066), .IN2(n5067), .IN3(n5068), .IN4(n5069), .Q(WX8434)
         );
  AND2X1 U4954 ( .IN1(n5070), .IN2(n3532), .Q(n5069) );
  AND2X1 U4955 ( .IN1(n3637), .IN2(n4800), .Q(n5068) );
  XNOR3X1 U4956 ( .IN1(n3242), .IN2(n3087), .IN3(n5071), .Q(n4800) );
  XOR2X1 U4957 ( .IN1(WX9792), .IN2(n7077), .Q(n5071) );
  AND2X1 U4958 ( .IN1(n3602), .IN2(CRC_OUT_3_15), .Q(n5067) );
  AND2X1 U4959 ( .IN1(n359), .IN2(n3580), .Q(n5066) );
  INVX0 U4960 ( .INP(n5072), .ZN(n359) );
  OR2X1 U4961 ( .IN1(n4417), .IN2(n3863), .Q(n5072) );
  OR4X1 U4962 ( .IN1(n5073), .IN2(n5074), .IN3(n5075), .IN4(n5076), .Q(WX8432)
         );
  AND2X1 U4963 ( .IN1(n3541), .IN2(n5077), .Q(n5076) );
  AND2X1 U4964 ( .IN1(n4807), .IN2(n3623), .Q(n5075) );
  XOR3X1 U4965 ( .IN1(n2873), .IN2(TM1), .IN3(n5078), .Q(n4807) );
  XNOR3X1 U4966 ( .IN1(test_so84), .IN2(n7078), .IN3(n3176), .Q(n5078) );
  AND2X1 U4967 ( .IN1(n3602), .IN2(CRC_OUT_3_16), .Q(n5074) );
  AND2X1 U4968 ( .IN1(n358), .IN2(n3580), .Q(n5073) );
  INVX0 U4969 ( .INP(n5079), .ZN(n358) );
  OR2X1 U4970 ( .IN1(n4417), .IN2(n3864), .Q(n5079) );
  OR4X1 U4971 ( .IN1(n5080), .IN2(n5081), .IN3(n5082), .IN4(n5083), .Q(WX8430)
         );
  AND2X1 U4972 ( .IN1(n3540), .IN2(n5084), .Q(n5083) );
  AND2X1 U4973 ( .IN1(n3637), .IN2(n4814), .Q(n5082) );
  XOR3X1 U4974 ( .IN1(n2874), .IN2(n3516), .IN3(n5085), .Q(n4814) );
  XOR3X1 U4975 ( .IN1(n7079), .IN2(n3241), .IN3(WX9852), .Q(n5085) );
  AND2X1 U4976 ( .IN1(n3603), .IN2(CRC_OUT_3_17), .Q(n5081) );
  AND2X1 U4977 ( .IN1(n357), .IN2(n3580), .Q(n5080) );
  INVX0 U4978 ( .INP(n5086), .ZN(n357) );
  OR2X1 U4979 ( .IN1(n4417), .IN2(n3865), .Q(n5086) );
  OR4X1 U4980 ( .IN1(n5087), .IN2(n5088), .IN3(n5089), .IN4(n5090), .Q(WX8428)
         );
  AND2X1 U4981 ( .IN1(n3540), .IN2(n5091), .Q(n5090) );
  AND2X1 U4982 ( .IN1(n4821), .IN2(n3623), .Q(n5089) );
  XOR3X1 U4983 ( .IN1(n2876), .IN2(TM1), .IN3(n5092), .Q(n4821) );
  XNOR3X1 U4984 ( .IN1(test_so82), .IN2(n7080), .IN3(n3240), .Q(n5092) );
  AND2X1 U4985 ( .IN1(n3603), .IN2(CRC_OUT_3_18), .Q(n5088) );
  AND2X1 U4986 ( .IN1(WX8266), .IN2(n3580), .Q(n5087) );
  OR4X1 U4987 ( .IN1(n5093), .IN2(n5094), .IN3(n5095), .IN4(n5096), .Q(WX8426)
         );
  AND2X1 U4988 ( .IN1(n3540), .IN2(n5097), .Q(n5096) );
  AND2X1 U4989 ( .IN1(n3637), .IN2(n4828), .Q(n5095) );
  XOR3X1 U4990 ( .IN1(n2877), .IN2(n3515), .IN3(n5098), .Q(n4828) );
  XOR3X1 U4991 ( .IN1(n7081), .IN2(n3239), .IN3(WX9848), .Q(n5098) );
  AND2X1 U4992 ( .IN1(n3603), .IN2(CRC_OUT_3_19), .Q(n5094) );
  AND2X1 U4993 ( .IN1(n355), .IN2(n3580), .Q(n5093) );
  INVX0 U4994 ( .INP(n5099), .ZN(n355) );
  OR2X1 U4995 ( .IN1(n4417), .IN2(n3867), .Q(n5099) );
  OR4X1 U4996 ( .IN1(n5100), .IN2(n5101), .IN3(n5102), .IN4(n5103), .Q(WX8424)
         );
  AND2X1 U4997 ( .IN1(n3540), .IN2(n5104), .Q(n5103) );
  AND2X1 U4998 ( .IN1(n4835), .IN2(n3623), .Q(n5102) );
  XOR3X1 U4999 ( .IN1(n2879), .IN2(TM1), .IN3(n5105), .Q(n4835) );
  XNOR3X1 U5000 ( .IN1(test_so80), .IN2(n7082), .IN3(n3238), .Q(n5105) );
  AND2X1 U5001 ( .IN1(n3603), .IN2(CRC_OUT_3_20), .Q(n5101) );
  AND2X1 U5002 ( .IN1(n354), .IN2(n3579), .Q(n5100) );
  INVX0 U5003 ( .INP(n5106), .ZN(n354) );
  OR2X1 U5004 ( .IN1(n4416), .IN2(n3868), .Q(n5106) );
  OR4X1 U5005 ( .IN1(n5107), .IN2(n5108), .IN3(n5109), .IN4(n5110), .Q(WX8422)
         );
  AND2X1 U5006 ( .IN1(n3540), .IN2(n5111), .Q(n5110) );
  AND2X1 U5007 ( .IN1(n3638), .IN2(n4842), .Q(n5109) );
  XOR3X1 U5008 ( .IN1(n2880), .IN2(n3514), .IN3(n5112), .Q(n4842) );
  XOR3X1 U5009 ( .IN1(n7083), .IN2(n3237), .IN3(WX9844), .Q(n5112) );
  AND2X1 U5010 ( .IN1(n3603), .IN2(CRC_OUT_3_21), .Q(n5108) );
  AND2X1 U5011 ( .IN1(n353), .IN2(n3579), .Q(n5107) );
  INVX0 U5012 ( .INP(n5113), .ZN(n353) );
  OR2X1 U5013 ( .IN1(n4416), .IN2(n3869), .Q(n5113) );
  OR4X1 U5014 ( .IN1(n5114), .IN2(n5115), .IN3(n5116), .IN4(n5117), .Q(WX8420)
         );
  AND2X1 U5015 ( .IN1(n3540), .IN2(n5118), .Q(n5117) );
  AND2X1 U5016 ( .IN1(n3638), .IN2(n4849), .Q(n5116) );
  XOR3X1 U5017 ( .IN1(n2882), .IN2(n3518), .IN3(n5119), .Q(n4849) );
  XOR3X1 U5018 ( .IN1(n7084), .IN2(n3236), .IN3(WX9842), .Q(n5119) );
  AND2X1 U5019 ( .IN1(n3603), .IN2(CRC_OUT_3_22), .Q(n5115) );
  AND2X1 U5020 ( .IN1(n352), .IN2(n3579), .Q(n5114) );
  INVX0 U5021 ( .INP(n5120), .ZN(n352) );
  OR2X1 U5022 ( .IN1(n4416), .IN2(n3870), .Q(n5120) );
  OR4X1 U5023 ( .IN1(n5121), .IN2(n5122), .IN3(n5123), .IN4(n5124), .Q(WX8418)
         );
  AND2X1 U5024 ( .IN1(n3540), .IN2(n5125), .Q(n5124) );
  AND2X1 U5025 ( .IN1(n3638), .IN2(n4856), .Q(n5123) );
  XOR3X1 U5026 ( .IN1(n2884), .IN2(n3516), .IN3(n5126), .Q(n4856) );
  XOR3X1 U5027 ( .IN1(n7085), .IN2(n3235), .IN3(WX9840), .Q(n5126) );
  AND2X1 U5028 ( .IN1(n3603), .IN2(CRC_OUT_3_23), .Q(n5122) );
  AND2X1 U5029 ( .IN1(n351), .IN2(n3579), .Q(n5121) );
  INVX0 U5030 ( .INP(n5127), .ZN(n351) );
  OR2X1 U5031 ( .IN1(n4416), .IN2(n3871), .Q(n5127) );
  OR4X1 U5032 ( .IN1(n5128), .IN2(n5129), .IN3(n5130), .IN4(n5131), .Q(WX8416)
         );
  AND2X1 U5033 ( .IN1(n3540), .IN2(n5132), .Q(n5131) );
  AND2X1 U5034 ( .IN1(n3638), .IN2(n4863), .Q(n5130) );
  XOR3X1 U5035 ( .IN1(n2886), .IN2(n3515), .IN3(n5133), .Q(n4863) );
  XOR3X1 U5036 ( .IN1(n7086), .IN2(n3234), .IN3(WX9838), .Q(n5133) );
  AND2X1 U5037 ( .IN1(test_so77), .IN2(n3587), .Q(n5129) );
  AND2X1 U5038 ( .IN1(n350), .IN2(n3579), .Q(n5128) );
  INVX0 U5039 ( .INP(n5134), .ZN(n350) );
  OR2X1 U5040 ( .IN1(n4416), .IN2(n3872), .Q(n5134) );
  OR4X1 U5041 ( .IN1(n5135), .IN2(n5136), .IN3(n5137), .IN4(n5138), .Q(WX8414)
         );
  AND2X1 U5042 ( .IN1(n3540), .IN2(n5139), .Q(n5138) );
  AND2X1 U5043 ( .IN1(n3638), .IN2(n4870), .Q(n5137) );
  XOR3X1 U5044 ( .IN1(n2888), .IN2(n3514), .IN3(n5140), .Q(n4870) );
  XOR3X1 U5045 ( .IN1(n7087), .IN2(n3233), .IN3(WX9836), .Q(n5140) );
  AND2X1 U5046 ( .IN1(n3603), .IN2(CRC_OUT_3_25), .Q(n5136) );
  AND2X1 U5047 ( .IN1(n349), .IN2(n3579), .Q(n5135) );
  INVX0 U5048 ( .INP(n5141), .ZN(n349) );
  OR2X1 U5049 ( .IN1(n4416), .IN2(n3873), .Q(n5141) );
  OR4X1 U5050 ( .IN1(n5142), .IN2(n5143), .IN3(n5144), .IN4(n5145), .Q(WX8412)
         );
  AND2X1 U5051 ( .IN1(n5146), .IN2(n3533), .Q(n5145) );
  AND2X1 U5052 ( .IN1(n3638), .IN2(n4877), .Q(n5144) );
  XOR3X1 U5053 ( .IN1(n2890), .IN2(n3518), .IN3(n5147), .Q(n4877) );
  XOR3X1 U5054 ( .IN1(n7088), .IN2(n3232), .IN3(WX9834), .Q(n5147) );
  AND2X1 U5055 ( .IN1(n3603), .IN2(CRC_OUT_3_26), .Q(n5143) );
  AND2X1 U5056 ( .IN1(n348), .IN2(n3579), .Q(n5142) );
  INVX0 U5057 ( .INP(n5148), .ZN(n348) );
  OR2X1 U5058 ( .IN1(n4416), .IN2(n3874), .Q(n5148) );
  OR4X1 U5059 ( .IN1(n5149), .IN2(n5150), .IN3(n5151), .IN4(n5152), .Q(WX8410)
         );
  AND2X1 U5060 ( .IN1(n3540), .IN2(n5153), .Q(n5152) );
  AND2X1 U5061 ( .IN1(n3638), .IN2(n4884), .Q(n5151) );
  XOR3X1 U5062 ( .IN1(n2892), .IN2(n3516), .IN3(n5154), .Q(n4884) );
  XOR3X1 U5063 ( .IN1(n7089), .IN2(n3231), .IN3(WX9832), .Q(n5154) );
  AND2X1 U5064 ( .IN1(n3603), .IN2(CRC_OUT_3_27), .Q(n5150) );
  AND2X1 U5065 ( .IN1(n347), .IN2(n3579), .Q(n5149) );
  INVX0 U5066 ( .INP(n5155), .ZN(n347) );
  OR2X1 U5067 ( .IN1(n4416), .IN2(n3875), .Q(n5155) );
  OR4X1 U5068 ( .IN1(n5156), .IN2(n5157), .IN3(n5158), .IN4(n5159), .Q(WX8408)
         );
  AND2X1 U5069 ( .IN1(n5160), .IN2(n3534), .Q(n5159) );
  AND2X1 U5070 ( .IN1(n3638), .IN2(n4891), .Q(n5158) );
  XOR3X1 U5071 ( .IN1(n2894), .IN2(n3515), .IN3(n5161), .Q(n4891) );
  XOR3X1 U5072 ( .IN1(n7090), .IN2(n3230), .IN3(WX9830), .Q(n5161) );
  AND2X1 U5073 ( .IN1(n3603), .IN2(CRC_OUT_3_28), .Q(n5157) );
  AND2X1 U5074 ( .IN1(n346), .IN2(n3579), .Q(n5156) );
  INVX0 U5075 ( .INP(n5162), .ZN(n346) );
  OR2X1 U5076 ( .IN1(n4416), .IN2(n3876), .Q(n5162) );
  OR4X1 U5077 ( .IN1(n5163), .IN2(n5164), .IN3(n5165), .IN4(n5166), .Q(WX8406)
         );
  AND2X1 U5078 ( .IN1(n3540), .IN2(n5167), .Q(n5166) );
  AND2X1 U5079 ( .IN1(n3638), .IN2(n4898), .Q(n5165) );
  XOR3X1 U5080 ( .IN1(n2896), .IN2(n3514), .IN3(n5168), .Q(n4898) );
  XOR3X1 U5081 ( .IN1(n7091), .IN2(n3229), .IN3(WX9828), .Q(n5168) );
  AND2X1 U5082 ( .IN1(n3603), .IN2(CRC_OUT_3_29), .Q(n5164) );
  AND2X1 U5083 ( .IN1(n345), .IN2(n3579), .Q(n5163) );
  INVX0 U5084 ( .INP(n5169), .ZN(n345) );
  OR2X1 U5085 ( .IN1(n4416), .IN2(n3877), .Q(n5169) );
  OR4X1 U5086 ( .IN1(n5170), .IN2(n5171), .IN3(n5172), .IN4(n5173), .Q(WX8404)
         );
  AND2X1 U5087 ( .IN1(n5174), .IN2(n3533), .Q(n5173) );
  AND2X1 U5088 ( .IN1(n3638), .IN2(n4905), .Q(n5172) );
  XOR3X1 U5089 ( .IN1(n2898), .IN2(n3518), .IN3(n5175), .Q(n4905) );
  XOR3X1 U5090 ( .IN1(n7092), .IN2(n3228), .IN3(WX9826), .Q(n5175) );
  AND2X1 U5091 ( .IN1(n3603), .IN2(CRC_OUT_3_30), .Q(n5171) );
  AND2X1 U5092 ( .IN1(n344), .IN2(n3579), .Q(n5170) );
  INVX0 U5093 ( .INP(n5176), .ZN(n344) );
  OR2X1 U5094 ( .IN1(n4416), .IN2(n3878), .Q(n5176) );
  OR4X1 U5095 ( .IN1(n5177), .IN2(n5178), .IN3(n5179), .IN4(n5180), .Q(WX8402)
         );
  AND2X1 U5096 ( .IN1(n3540), .IN2(n5181), .Q(n5180) );
  AND2X1 U5097 ( .IN1(n4912), .IN2(n3623), .Q(n5179) );
  XOR3X1 U5098 ( .IN1(n2834), .IN2(TM1), .IN3(n5182), .Q(n4912) );
  XOR3X1 U5099 ( .IN1(test_so85), .IN2(n7093), .IN3(WX9824), .Q(n5182) );
  AND2X1 U5100 ( .IN1(n2245), .IN2(WX8243), .Q(n5178) );
  AND2X1 U5101 ( .IN1(n3604), .IN2(CRC_OUT_3_31), .Q(n5177) );
  AND2X1 U5102 ( .IN1(n3506), .IN2(n4361), .Q(WX8304) );
  AND2X1 U5103 ( .IN1(n5183), .IN2(n8399), .Q(WX8266) );
  AND2X1 U5104 ( .IN1(n5184), .IN2(n4361), .Q(WX7791) );
  XOR2X1 U5105 ( .IN1(CRC_OUT_4_30), .IN2(n3281), .Q(n5184) );
  AND2X1 U5106 ( .IN1(n5185), .IN2(n4360), .Q(WX7789) );
  XOR2X1 U5107 ( .IN1(test_so66), .IN2(n3282), .Q(n5185) );
  AND2X1 U5108 ( .IN1(n5186), .IN2(n4360), .Q(WX7787) );
  XOR2X1 U5109 ( .IN1(CRC_OUT_4_28), .IN2(n3283), .Q(n5186) );
  AND2X1 U5110 ( .IN1(n5187), .IN2(n4360), .Q(WX7785) );
  XOR2X1 U5111 ( .IN1(CRC_OUT_4_27), .IN2(n3284), .Q(n5187) );
  AND2X1 U5112 ( .IN1(n5188), .IN2(n5183), .Q(WX7783) );
  XOR2X1 U5113 ( .IN1(CRC_OUT_4_26), .IN2(n3285), .Q(n5188) );
  AND2X1 U5114 ( .IN1(n5189), .IN2(n4360), .Q(WX7781) );
  XOR2X1 U5115 ( .IN1(CRC_OUT_4_25), .IN2(n3286), .Q(n5189) );
  AND2X1 U5116 ( .IN1(n5190), .IN2(n4360), .Q(WX7779) );
  XOR2X1 U5117 ( .IN1(CRC_OUT_4_24), .IN2(n3287), .Q(n5190) );
  AND2X1 U5118 ( .IN1(n5191), .IN2(n4360), .Q(WX7777) );
  XOR2X1 U5119 ( .IN1(CRC_OUT_4_23), .IN2(n3288), .Q(n5191) );
  AND2X1 U5120 ( .IN1(n5192), .IN2(n4360), .Q(WX7775) );
  XOR2X1 U5121 ( .IN1(CRC_OUT_4_22), .IN2(n3289), .Q(n5192) );
  AND2X1 U5122 ( .IN1(n5193), .IN2(n4360), .Q(WX7773) );
  XOR2X1 U5123 ( .IN1(CRC_OUT_4_21), .IN2(n3290), .Q(n5193) );
  AND2X1 U5124 ( .IN1(n5194), .IN2(n4360), .Q(WX7771) );
  XOR2X1 U5125 ( .IN1(test_so63), .IN2(DFF_1140_n1), .Q(n5194) );
  AND2X1 U5126 ( .IN1(n5195), .IN2(n4359), .Q(WX7769) );
  XOR2X1 U5127 ( .IN1(CRC_OUT_4_19), .IN2(n3291), .Q(n5195) );
  AND2X1 U5128 ( .IN1(n5196), .IN2(n4359), .Q(WX7767) );
  XOR2X1 U5129 ( .IN1(CRC_OUT_4_18), .IN2(n3292), .Q(n5196) );
  AND2X1 U5130 ( .IN1(n5197), .IN2(n4359), .Q(WX7765) );
  XOR2X1 U5131 ( .IN1(CRC_OUT_4_17), .IN2(n3293), .Q(n5197) );
  AND2X1 U5132 ( .IN1(n5198), .IN2(n4359), .Q(WX7763) );
  XOR2X1 U5133 ( .IN1(CRC_OUT_4_16), .IN2(n3294), .Q(n5198) );
  AND2X1 U5134 ( .IN1(n5199), .IN2(n4359), .Q(WX7761) );
  XOR3X1 U5135 ( .IN1(n3182), .IN2(DFF_1151_n1), .IN3(DFF_1135_n1), .Q(n5199)
         );
  AND2X1 U5136 ( .IN1(n5200), .IN2(n4359), .Q(WX7759) );
  XOR2X1 U5137 ( .IN1(CRC_OUT_4_14), .IN2(n3295), .Q(n5200) );
  AND2X1 U5138 ( .IN1(n5201), .IN2(n4359), .Q(WX7757) );
  XOR2X1 U5139 ( .IN1(CRC_OUT_4_13), .IN2(n3296), .Q(n5201) );
  AND2X1 U5140 ( .IN1(n5202), .IN2(n4359), .Q(WX7755) );
  XOR2X1 U5141 ( .IN1(test_so65), .IN2(n3297), .Q(n5202) );
  AND2X1 U5142 ( .IN1(n5203), .IN2(n4359), .Q(WX7753) );
  XOR2X1 U5143 ( .IN1(CRC_OUT_4_11), .IN2(n3298), .Q(n5203) );
  AND2X1 U5144 ( .IN1(n5204), .IN2(n4358), .Q(WX7751) );
  XOR3X1 U5145 ( .IN1(n3183), .IN2(DFF_1151_n1), .IN3(DFF_1130_n1), .Q(n5204)
         );
  AND2X1 U5146 ( .IN1(n5205), .IN2(n4358), .Q(WX7749) );
  XOR2X1 U5147 ( .IN1(CRC_OUT_4_9), .IN2(n3299), .Q(n5205) );
  AND2X1 U5148 ( .IN1(n5206), .IN2(n4358), .Q(WX7747) );
  XOR2X1 U5149 ( .IN1(CRC_OUT_4_8), .IN2(n3300), .Q(n5206) );
  AND2X1 U5150 ( .IN1(n5207), .IN2(n4358), .Q(WX7745) );
  XOR2X1 U5151 ( .IN1(CRC_OUT_4_7), .IN2(n3301), .Q(n5207) );
  AND2X1 U5152 ( .IN1(n5208), .IN2(n4358), .Q(WX7743) );
  XOR2X1 U5153 ( .IN1(CRC_OUT_4_6), .IN2(n3302), .Q(n5208) );
  AND2X1 U5154 ( .IN1(n5209), .IN2(n4358), .Q(WX7741) );
  XOR2X1 U5155 ( .IN1(CRC_OUT_4_5), .IN2(n3303), .Q(n5209) );
  AND2X1 U5156 ( .IN1(n5210), .IN2(n4358), .Q(WX7739) );
  XOR2X1 U5157 ( .IN1(CRC_OUT_4_4), .IN2(n3304), .Q(n5210) );
  AND2X1 U5158 ( .IN1(n5211), .IN2(n4354), .Q(WX7737) );
  XOR3X1 U5159 ( .IN1(test_so64), .IN2(DFF_1151_n1), .IN3(CRC_OUT_4_3), .Q(
        n5211) );
  AND2X1 U5160 ( .IN1(n5212), .IN2(n4351), .Q(WX7735) );
  XOR2X1 U5161 ( .IN1(CRC_OUT_4_2), .IN2(n3305), .Q(n5212) );
  AND2X1 U5162 ( .IN1(n5213), .IN2(n4351), .Q(WX7733) );
  XOR2X1 U5163 ( .IN1(CRC_OUT_4_1), .IN2(n3306), .Q(n5213) );
  AND2X1 U5164 ( .IN1(n5214), .IN2(n4351), .Q(WX7731) );
  XOR2X1 U5165 ( .IN1(CRC_OUT_4_0), .IN2(n3307), .Q(n5214) );
  AND2X1 U5166 ( .IN1(n5215), .IN2(n4351), .Q(WX7729) );
  XOR2X1 U5167 ( .IN1(n3197), .IN2(CRC_OUT_4_31), .Q(n5215) );
  INVX0 U5168 ( .INP(n5216), .ZN(WX7203) );
  OR2X1 U5169 ( .IN1(n4416), .IN2(n7134), .Q(n5216) );
  INVX0 U5170 ( .INP(n5217), .ZN(WX7201) );
  OR2X1 U5171 ( .IN1(n4415), .IN2(n7135), .Q(n5217) );
  INVX0 U5172 ( .INP(n5218), .ZN(WX7199) );
  OR2X1 U5173 ( .IN1(n4415), .IN2(n7136), .Q(n5218) );
  INVX0 U5174 ( .INP(n5219), .ZN(WX7197) );
  OR2X1 U5175 ( .IN1(n4415), .IN2(n7137), .Q(n5219) );
  INVX0 U5176 ( .INP(n5220), .ZN(WX7195) );
  OR2X1 U5177 ( .IN1(n4415), .IN2(n7138), .Q(n5220) );
  INVX0 U5178 ( .INP(n5221), .ZN(WX7193) );
  OR2X1 U5179 ( .IN1(n4415), .IN2(n7139), .Q(n5221) );
  INVX0 U5180 ( .INP(n5222), .ZN(WX7191) );
  OR2X1 U5181 ( .IN1(n4415), .IN2(n7140), .Q(n5222) );
  INVX0 U5182 ( .INP(n5223), .ZN(WX7189) );
  OR2X1 U5183 ( .IN1(n4415), .IN2(n7141), .Q(n5223) );
  INVX0 U5184 ( .INP(n5224), .ZN(WX7187) );
  OR2X1 U5185 ( .IN1(n4415), .IN2(n7142), .Q(n5224) );
  INVX0 U5186 ( .INP(n5225), .ZN(WX7185) );
  OR2X1 U5187 ( .IN1(n4415), .IN2(n7143), .Q(n5225) );
  INVX0 U5188 ( .INP(n5226), .ZN(WX7183) );
  OR2X1 U5189 ( .IN1(n4415), .IN2(n7144), .Q(n5226) );
  AND2X1 U5190 ( .IN1(test_so57), .IN2(n4351), .Q(WX7181) );
  INVX0 U5191 ( .INP(n5227), .ZN(WX7179) );
  OR2X1 U5192 ( .IN1(n4415), .IN2(n7146), .Q(n5227) );
  INVX0 U5193 ( .INP(n5228), .ZN(WX7177) );
  OR2X1 U5194 ( .IN1(n4415), .IN2(n7147), .Q(n5228) );
  INVX0 U5195 ( .INP(n5229), .ZN(WX7175) );
  OR2X1 U5196 ( .IN1(n4415), .IN2(n7148), .Q(n5229) );
  INVX0 U5197 ( .INP(n5230), .ZN(WX7173) );
  OR2X1 U5198 ( .IN1(n4414), .IN2(n7149), .Q(n5230) );
  OR4X1 U5199 ( .IN1(n5231), .IN2(n5232), .IN3(n5233), .IN4(n5234), .Q(WX7171)
         );
  AND2X1 U5200 ( .IN1(n3540), .IN2(n5235), .Q(n5234) );
  AND2X1 U5201 ( .IN1(n3638), .IN2(n4965), .Q(n5233) );
  XNOR3X1 U5202 ( .IN1(n3196), .IN2(n3088), .IN3(n5236), .Q(n4965) );
  XOR2X1 U5203 ( .IN1(WX8529), .IN2(n7094), .Q(n5236) );
  AND2X1 U5204 ( .IN1(n3604), .IN2(CRC_OUT_4_0), .Q(n5232) );
  AND2X1 U5205 ( .IN1(n312), .IN2(n3579), .Q(n5231) );
  INVX0 U5206 ( .INP(n5237), .ZN(n312) );
  OR2X1 U5207 ( .IN1(n4414), .IN2(n3879), .Q(n5237) );
  OR4X1 U5208 ( .IN1(n5238), .IN2(n5239), .IN3(n5240), .IN4(n5241), .Q(WX7169)
         );
  AND2X1 U5209 ( .IN1(n3538), .IN2(n5242), .Q(n5241) );
  AND2X1 U5210 ( .IN1(n3638), .IN2(n4972), .Q(n5240) );
  XNOR3X1 U5211 ( .IN1(n3280), .IN2(n3089), .IN3(n5243), .Q(n4972) );
  XOR2X1 U5212 ( .IN1(WX8527), .IN2(n7095), .Q(n5243) );
  AND2X1 U5213 ( .IN1(n3604), .IN2(CRC_OUT_4_1), .Q(n5239) );
  AND2X1 U5214 ( .IN1(n311), .IN2(n3578), .Q(n5238) );
  INVX0 U5215 ( .INP(n5244), .ZN(n311) );
  OR2X1 U5216 ( .IN1(n4414), .IN2(n3880), .Q(n5244) );
  OR4X1 U5217 ( .IN1(n5245), .IN2(n5246), .IN3(n5247), .IN4(n5248), .Q(WX7167)
         );
  AND2X1 U5218 ( .IN1(n3538), .IN2(n5249), .Q(n5248) );
  AND2X1 U5219 ( .IN1(n3638), .IN2(n4979), .Q(n5247) );
  XNOR3X1 U5220 ( .IN1(n3279), .IN2(n3090), .IN3(n5250), .Q(n4979) );
  XOR2X1 U5221 ( .IN1(WX8525), .IN2(n7096), .Q(n5250) );
  AND2X1 U5222 ( .IN1(n3604), .IN2(CRC_OUT_4_2), .Q(n5246) );
  AND2X1 U5223 ( .IN1(n310), .IN2(n3578), .Q(n5245) );
  INVX0 U5224 ( .INP(n5251), .ZN(n310) );
  OR2X1 U5225 ( .IN1(n4414), .IN2(n3881), .Q(n5251) );
  OR4X1 U5226 ( .IN1(n5252), .IN2(n5253), .IN3(n5254), .IN4(n5255), .Q(WX7165)
         );
  AND2X1 U5227 ( .IN1(n3538), .IN2(n5256), .Q(n5255) );
  AND2X1 U5228 ( .IN1(n3640), .IN2(n4986), .Q(n5254) );
  XNOR3X1 U5229 ( .IN1(n3277), .IN2(n3091), .IN3(n5257), .Q(n4986) );
  XOR2X1 U5230 ( .IN1(WX8523), .IN2(n7097), .Q(n5257) );
  AND2X1 U5231 ( .IN1(n3604), .IN2(CRC_OUT_4_3), .Q(n5253) );
  AND2X1 U5232 ( .IN1(n309), .IN2(n3578), .Q(n5252) );
  INVX0 U5233 ( .INP(n5258), .ZN(n309) );
  OR2X1 U5234 ( .IN1(n4414), .IN2(n3882), .Q(n5258) );
  OR4X1 U5235 ( .IN1(n5259), .IN2(n5260), .IN3(n5261), .IN4(n5262), .Q(WX7163)
         );
  AND2X1 U5236 ( .IN1(n5263), .IN2(n3531), .Q(n5262) );
  AND2X1 U5237 ( .IN1(n3640), .IN2(n4993), .Q(n5261) );
  XNOR3X1 U5238 ( .IN1(n3181), .IN2(n3092), .IN3(n5264), .Q(n4993) );
  XOR2X1 U5239 ( .IN1(WX8521), .IN2(n7098), .Q(n5264) );
  AND2X1 U5240 ( .IN1(n3604), .IN2(CRC_OUT_4_4), .Q(n5260) );
  AND2X1 U5241 ( .IN1(n308), .IN2(n3578), .Q(n5259) );
  INVX0 U5242 ( .INP(n5265), .ZN(n308) );
  OR2X1 U5243 ( .IN1(n4414), .IN2(n3883), .Q(n5265) );
  OR4X1 U5244 ( .IN1(n5266), .IN2(n5267), .IN3(n5268), .IN4(n5269), .Q(WX7161)
         );
  AND2X1 U5245 ( .IN1(n3538), .IN2(n5270), .Q(n5269) );
  AND2X1 U5246 ( .IN1(n3640), .IN2(n5000), .Q(n5268) );
  XNOR3X1 U5247 ( .IN1(n3276), .IN2(n3093), .IN3(n5271), .Q(n5000) );
  XOR2X1 U5248 ( .IN1(WX8519), .IN2(n7099), .Q(n5271) );
  AND2X1 U5249 ( .IN1(n3604), .IN2(CRC_OUT_4_5), .Q(n5267) );
  AND2X1 U5250 ( .IN1(WX6999), .IN2(n3578), .Q(n5266) );
  OR4X1 U5251 ( .IN1(n5272), .IN2(n5273), .IN3(n5274), .IN4(n5275), .Q(WX7159)
         );
  AND2X1 U5252 ( .IN1(n5276), .IN2(n3531), .Q(n5275) );
  AND2X1 U5253 ( .IN1(n3640), .IN2(n5007), .Q(n5274) );
  XNOR3X1 U5254 ( .IN1(n3275), .IN2(n3094), .IN3(n5277), .Q(n5007) );
  XOR2X1 U5255 ( .IN1(WX8517), .IN2(n7100), .Q(n5277) );
  AND2X1 U5256 ( .IN1(n3604), .IN2(CRC_OUT_4_6), .Q(n5273) );
  AND2X1 U5257 ( .IN1(n306), .IN2(n3578), .Q(n5272) );
  INVX0 U5258 ( .INP(n5278), .ZN(n306) );
  OR2X1 U5259 ( .IN1(n4414), .IN2(n3885), .Q(n5278) );
  OR4X1 U5260 ( .IN1(n5279), .IN2(n5280), .IN3(n5281), .IN4(n5282), .Q(WX7157)
         );
  AND2X1 U5261 ( .IN1(n3538), .IN2(n5283), .Q(n5282) );
  AND2X1 U5262 ( .IN1(n3640), .IN2(n5014), .Q(n5281) );
  XNOR3X1 U5263 ( .IN1(n3274), .IN2(n3095), .IN3(n5284), .Q(n5014) );
  XOR2X1 U5264 ( .IN1(WX8515), .IN2(n7101), .Q(n5284) );
  AND2X1 U5265 ( .IN1(n3604), .IN2(CRC_OUT_4_7), .Q(n5280) );
  AND2X1 U5266 ( .IN1(n305), .IN2(n3578), .Q(n5279) );
  INVX0 U5267 ( .INP(n5285), .ZN(n305) );
  OR2X1 U5268 ( .IN1(n4414), .IN2(n3886), .Q(n5285) );
  OR4X1 U5269 ( .IN1(n5286), .IN2(n5287), .IN3(n5288), .IN4(n5289), .Q(WX7155)
         );
  AND2X1 U5270 ( .IN1(n5290), .IN2(n3530), .Q(n5289) );
  AND2X1 U5271 ( .IN1(n3640), .IN2(n5021), .Q(n5288) );
  XNOR3X1 U5272 ( .IN1(n3273), .IN2(n3096), .IN3(n5291), .Q(n5021) );
  XOR2X1 U5273 ( .IN1(WX8513), .IN2(n7102), .Q(n5291) );
  AND2X1 U5274 ( .IN1(n3604), .IN2(CRC_OUT_4_8), .Q(n5287) );
  AND2X1 U5275 ( .IN1(n304), .IN2(n3578), .Q(n5286) );
  INVX0 U5276 ( .INP(n5292), .ZN(n304) );
  OR2X1 U5277 ( .IN1(n4414), .IN2(n3887), .Q(n5292) );
  OR4X1 U5278 ( .IN1(n5293), .IN2(n5294), .IN3(n5295), .IN4(n5296), .Q(WX7153)
         );
  AND2X1 U5279 ( .IN1(n3538), .IN2(n5297), .Q(n5296) );
  AND2X1 U5280 ( .IN1(n5028), .IN2(n3622), .Q(n5295) );
  XOR3X1 U5281 ( .IN1(n3613), .IN2(n3097), .IN3(n5298), .Q(n5028) );
  XOR2X1 U5282 ( .IN1(WX8447), .IN2(test_so75), .Q(n5298) );
  AND2X1 U5283 ( .IN1(n3604), .IN2(CRC_OUT_4_9), .Q(n5294) );
  AND2X1 U5284 ( .IN1(n303), .IN2(n3578), .Q(n5293) );
  INVX0 U5285 ( .INP(n5299), .ZN(n303) );
  OR2X1 U5286 ( .IN1(n4414), .IN2(n3888), .Q(n5299) );
  OR4X1 U5287 ( .IN1(n5300), .IN2(n5301), .IN3(n5302), .IN4(n5303), .Q(WX7151)
         );
  AND2X1 U5288 ( .IN1(n5304), .IN2(n3530), .Q(n5303) );
  AND2X1 U5289 ( .IN1(n3640), .IN2(n5035), .Q(n5302) );
  XNOR3X1 U5290 ( .IN1(n3272), .IN2(n3098), .IN3(n5305), .Q(n5035) );
  XOR2X1 U5291 ( .IN1(WX8509), .IN2(n7103), .Q(n5305) );
  AND2X1 U5292 ( .IN1(n3604), .IN2(CRC_OUT_4_10), .Q(n5301) );
  AND2X1 U5293 ( .IN1(n302), .IN2(n3578), .Q(n5300) );
  INVX0 U5294 ( .INP(n5306), .ZN(n302) );
  OR2X1 U5295 ( .IN1(n4414), .IN2(n3889), .Q(n5306) );
  OR4X1 U5296 ( .IN1(n5307), .IN2(n5308), .IN3(n5309), .IN4(n5310), .Q(WX7149)
         );
  AND2X1 U5297 ( .IN1(n3538), .IN2(n5311), .Q(n5310) );
  AND2X1 U5298 ( .IN1(n5042), .IN2(n3622), .Q(n5309) );
  XOR3X1 U5299 ( .IN1(n3617), .IN2(n3180), .IN3(n5312), .Q(n5042) );
  XOR2X1 U5300 ( .IN1(WX8443), .IN2(test_so73), .Q(n5312) );
  AND2X1 U5301 ( .IN1(n3605), .IN2(CRC_OUT_4_11), .Q(n5308) );
  AND2X1 U5302 ( .IN1(n301), .IN2(n3578), .Q(n5307) );
  INVX0 U5303 ( .INP(n5313), .ZN(n301) );
  OR2X1 U5304 ( .IN1(n4414), .IN2(n3890), .Q(n5313) );
  OR4X1 U5305 ( .IN1(n5314), .IN2(n5315), .IN3(n5316), .IN4(n5317), .Q(WX7147)
         );
  AND2X1 U5306 ( .IN1(n3538), .IN2(n5318), .Q(n5317) );
  AND2X1 U5307 ( .IN1(n3640), .IN2(n5049), .Q(n5316) );
  XNOR3X1 U5308 ( .IN1(n3271), .IN2(n3099), .IN3(n5319), .Q(n5049) );
  XOR2X1 U5309 ( .IN1(WX8505), .IN2(n7104), .Q(n5319) );
  AND2X1 U5310 ( .IN1(test_so65), .IN2(n3587), .Q(n5315) );
  AND2X1 U5311 ( .IN1(n300), .IN2(n3578), .Q(n5314) );
  INVX0 U5312 ( .INP(n5320), .ZN(n300) );
  OR2X1 U5313 ( .IN1(n4414), .IN2(n3891), .Q(n5320) );
  OR4X1 U5314 ( .IN1(n5321), .IN2(n5322), .IN3(n5323), .IN4(n5324), .Q(WX7145)
         );
  AND2X1 U5315 ( .IN1(n3538), .IN2(n5325), .Q(n5324) );
  AND2X1 U5316 ( .IN1(n5056), .IN2(n3622), .Q(n5323) );
  XOR3X1 U5317 ( .IN1(n3270), .IN2(n3100), .IN3(n5326), .Q(n5056) );
  XOR2X1 U5318 ( .IN1(WX8439), .IN2(test_so71), .Q(n5326) );
  AND2X1 U5319 ( .IN1(n3605), .IN2(CRC_OUT_4_13), .Q(n5322) );
  AND2X1 U5320 ( .IN1(n299), .IN2(n3577), .Q(n5321) );
  INVX0 U5321 ( .INP(n5327), .ZN(n299) );
  OR2X1 U5322 ( .IN1(n4413), .IN2(n3892), .Q(n5327) );
  OR4X1 U5323 ( .IN1(n5328), .IN2(n5329), .IN3(n5330), .IN4(n5331), .Q(WX7143)
         );
  AND2X1 U5324 ( .IN1(n3534), .IN2(n5332), .Q(n5331) );
  AND2X1 U5325 ( .IN1(n3640), .IN2(n5063), .Q(n5330) );
  XNOR3X1 U5326 ( .IN1(n3269), .IN2(n3101), .IN3(n5333), .Q(n5063) );
  XOR2X1 U5327 ( .IN1(WX8501), .IN2(n7105), .Q(n5333) );
  AND2X1 U5328 ( .IN1(n3605), .IN2(CRC_OUT_4_14), .Q(n5329) );
  AND2X1 U5329 ( .IN1(n298), .IN2(n3577), .Q(n5328) );
  INVX0 U5330 ( .INP(n5334), .ZN(n298) );
  OR2X1 U5331 ( .IN1(n4413), .IN2(n3893), .Q(n5334) );
  OR4X1 U5332 ( .IN1(n5335), .IN2(n5336), .IN3(n5337), .IN4(n5338), .Q(WX7141)
         );
  AND2X1 U5333 ( .IN1(n3534), .IN2(n5339), .Q(n5338) );
  AND2X1 U5334 ( .IN1(n5070), .IN2(n3622), .Q(n5337) );
  XOR3X1 U5335 ( .IN1(n3625), .IN2(n3268), .IN3(n5340), .Q(n5070) );
  XOR2X1 U5336 ( .IN1(WX8563), .IN2(test_so69), .Q(n5340) );
  AND2X1 U5337 ( .IN1(n3605), .IN2(CRC_OUT_4_15), .Q(n5336) );
  AND2X1 U5338 ( .IN1(n297), .IN2(n3577), .Q(n5335) );
  INVX0 U5339 ( .INP(n5341), .ZN(n297) );
  OR2X1 U5340 ( .IN1(n4413), .IN2(n3894), .Q(n5341) );
  OR4X1 U5341 ( .IN1(n5342), .IN2(n5343), .IN3(n5344), .IN4(n5345), .Q(WX7139)
         );
  AND2X1 U5342 ( .IN1(n3534), .IN2(n5346), .Q(n5345) );
  AND2X1 U5343 ( .IN1(n3640), .IN2(n5077), .Q(n5344) );
  XOR3X1 U5344 ( .IN1(n2900), .IN2(n3516), .IN3(n5347), .Q(n5077) );
  XOR3X1 U5345 ( .IN1(n7106), .IN2(n3179), .IN3(WX8561), .Q(n5347) );
  AND2X1 U5346 ( .IN1(n3605), .IN2(CRC_OUT_4_16), .Q(n5343) );
  AND2X1 U5347 ( .IN1(n296), .IN2(n3577), .Q(n5342) );
  INVX0 U5348 ( .INP(n5348), .ZN(n296) );
  OR2X1 U5349 ( .IN1(n4413), .IN2(n3895), .Q(n5348) );
  OR4X1 U5350 ( .IN1(n5349), .IN2(n5350), .IN3(n5351), .IN4(n5352), .Q(WX7137)
         );
  AND2X1 U5351 ( .IN1(n3534), .IN2(n5353), .Q(n5352) );
  AND2X1 U5352 ( .IN1(n3640), .IN2(n5084), .Q(n5351) );
  XOR3X1 U5353 ( .IN1(n2902), .IN2(n3515), .IN3(n5354), .Q(n5084) );
  XOR3X1 U5354 ( .IN1(n7107), .IN2(n3267), .IN3(WX8559), .Q(n5354) );
  AND2X1 U5355 ( .IN1(n3605), .IN2(CRC_OUT_4_17), .Q(n5350) );
  AND2X1 U5356 ( .IN1(n295), .IN2(n3577), .Q(n5349) );
  INVX0 U5357 ( .INP(n5355), .ZN(n295) );
  OR2X1 U5358 ( .IN1(n4413), .IN2(n3896), .Q(n5355) );
  OR4X1 U5359 ( .IN1(n5356), .IN2(n5357), .IN3(n5358), .IN4(n5359), .Q(WX7135)
         );
  AND2X1 U5360 ( .IN1(n3534), .IN2(n5360), .Q(n5359) );
  AND2X1 U5361 ( .IN1(n3640), .IN2(n5091), .Q(n5358) );
  XOR3X1 U5362 ( .IN1(n2904), .IN2(n3514), .IN3(n5361), .Q(n5091) );
  XOR3X1 U5363 ( .IN1(n7108), .IN2(n3266), .IN3(WX8557), .Q(n5361) );
  AND2X1 U5364 ( .IN1(n3605), .IN2(CRC_OUT_4_18), .Q(n5357) );
  AND2X1 U5365 ( .IN1(n294), .IN2(n3577), .Q(n5356) );
  INVX0 U5366 ( .INP(n5362), .ZN(n294) );
  OR2X1 U5367 ( .IN1(n4413), .IN2(n3897), .Q(n5362) );
  OR4X1 U5368 ( .IN1(n5363), .IN2(n5364), .IN3(n5365), .IN4(n5366), .Q(WX7133)
         );
  AND2X1 U5369 ( .IN1(n3536), .IN2(n5367), .Q(n5366) );
  AND2X1 U5370 ( .IN1(n3641), .IN2(n5097), .Q(n5365) );
  XOR3X1 U5371 ( .IN1(n2906), .IN2(n3518), .IN3(n5368), .Q(n5097) );
  XOR3X1 U5372 ( .IN1(n7109), .IN2(n3265), .IN3(WX8555), .Q(n5368) );
  AND2X1 U5373 ( .IN1(n3605), .IN2(CRC_OUT_4_19), .Q(n5364) );
  AND2X1 U5374 ( .IN1(n293), .IN2(n3577), .Q(n5363) );
  INVX0 U5375 ( .INP(n5369), .ZN(n293) );
  OR2X1 U5376 ( .IN1(n4413), .IN2(n3898), .Q(n5369) );
  OR4X1 U5377 ( .IN1(n5370), .IN2(n5371), .IN3(n5372), .IN4(n5373), .Q(WX7131)
         );
  AND2X1 U5378 ( .IN1(n3534), .IN2(n5374), .Q(n5373) );
  AND2X1 U5379 ( .IN1(n3641), .IN2(n5104), .Q(n5372) );
  XOR3X1 U5380 ( .IN1(n2908), .IN2(n3516), .IN3(n5375), .Q(n5104) );
  XOR3X1 U5381 ( .IN1(n7110), .IN2(n3264), .IN3(WX8553), .Q(n5375) );
  AND2X1 U5382 ( .IN1(n3605), .IN2(CRC_OUT_4_20), .Q(n5371) );
  AND2X1 U5383 ( .IN1(n292), .IN2(n3577), .Q(n5370) );
  INVX0 U5384 ( .INP(n5376), .ZN(n292) );
  OR2X1 U5385 ( .IN1(n4413), .IN2(n3899), .Q(n5376) );
  OR4X1 U5386 ( .IN1(n5377), .IN2(n5378), .IN3(n5379), .IN4(n5380), .Q(WX7129)
         );
  AND2X1 U5387 ( .IN1(n5381), .IN2(n3532), .Q(n5380) );
  AND2X1 U5388 ( .IN1(n3641), .IN2(n5111), .Q(n5379) );
  XOR3X1 U5389 ( .IN1(n2910), .IN2(n3515), .IN3(n5382), .Q(n5111) );
  XOR3X1 U5390 ( .IN1(n7111), .IN2(n3263), .IN3(WX8551), .Q(n5382) );
  AND2X1 U5391 ( .IN1(n3605), .IN2(CRC_OUT_4_21), .Q(n5378) );
  AND2X1 U5392 ( .IN1(n291), .IN2(n3577), .Q(n5377) );
  INVX0 U5393 ( .INP(n5383), .ZN(n291) );
  OR2X1 U5394 ( .IN1(n4413), .IN2(n3900), .Q(n5383) );
  OR4X1 U5395 ( .IN1(n5384), .IN2(n5385), .IN3(n5386), .IN4(n5387), .Q(WX7127)
         );
  AND2X1 U5396 ( .IN1(n3534), .IN2(n5388), .Q(n5387) );
  AND2X1 U5397 ( .IN1(n3641), .IN2(n5118), .Q(n5386) );
  XOR3X1 U5398 ( .IN1(n2912), .IN2(n3514), .IN3(n5389), .Q(n5118) );
  XOR3X1 U5399 ( .IN1(n7112), .IN2(n3262), .IN3(WX8549), .Q(n5389) );
  AND2X1 U5400 ( .IN1(n3605), .IN2(CRC_OUT_4_22), .Q(n5385) );
  AND2X1 U5401 ( .IN1(n290), .IN2(n3577), .Q(n5384) );
  INVX0 U5402 ( .INP(n5390), .ZN(n290) );
  OR2X1 U5403 ( .IN1(n4413), .IN2(n3901), .Q(n5390) );
  OR4X1 U5404 ( .IN1(n5391), .IN2(n5392), .IN3(n5393), .IN4(n5394), .Q(WX7125)
         );
  AND2X1 U5405 ( .IN1(n5395), .IN2(n3533), .Q(n5394) );
  AND2X1 U5406 ( .IN1(n3641), .IN2(n5125), .Q(n5393) );
  XOR3X1 U5407 ( .IN1(n2914), .IN2(n3518), .IN3(n5396), .Q(n5125) );
  XOR3X1 U5408 ( .IN1(n7113), .IN2(n3261), .IN3(WX8547), .Q(n5396) );
  AND2X1 U5409 ( .IN1(n3605), .IN2(CRC_OUT_4_23), .Q(n5392) );
  AND2X1 U5410 ( .IN1(n289), .IN2(n3577), .Q(n5391) );
  INVX0 U5411 ( .INP(n5397), .ZN(n289) );
  OR2X1 U5412 ( .IN1(n4413), .IN2(n3902), .Q(n5397) );
  OR4X1 U5413 ( .IN1(n5398), .IN2(n5399), .IN3(n5400), .IN4(n5401), .Q(WX7123)
         );
  AND2X1 U5414 ( .IN1(n3534), .IN2(n5402), .Q(n5401) );
  AND2X1 U5415 ( .IN1(n3641), .IN2(n5132), .Q(n5400) );
  XOR3X1 U5416 ( .IN1(n2916), .IN2(n3516), .IN3(n5403), .Q(n5132) );
  XOR3X1 U5417 ( .IN1(n7114), .IN2(n3260), .IN3(WX8545), .Q(n5403) );
  AND2X1 U5418 ( .IN1(n3605), .IN2(CRC_OUT_4_24), .Q(n5399) );
  AND2X1 U5419 ( .IN1(n288), .IN2(n3577), .Q(n5398) );
  INVX0 U5420 ( .INP(n5404), .ZN(n288) );
  OR2X1 U5421 ( .IN1(n4413), .IN2(n3903), .Q(n5404) );
  OR4X1 U5422 ( .IN1(n5405), .IN2(n5406), .IN3(n5407), .IN4(n5408), .Q(WX7121)
         );
  AND2X1 U5423 ( .IN1(n5409), .IN2(n3533), .Q(n5408) );
  AND2X1 U5424 ( .IN1(n3641), .IN2(n5139), .Q(n5407) );
  XOR3X1 U5425 ( .IN1(n2918), .IN2(n3515), .IN3(n5410), .Q(n5139) );
  XOR3X1 U5426 ( .IN1(n7115), .IN2(n3259), .IN3(WX8543), .Q(n5410) );
  AND2X1 U5427 ( .IN1(n3606), .IN2(CRC_OUT_4_25), .Q(n5406) );
  AND2X1 U5428 ( .IN1(n287), .IN2(n3576), .Q(n5405) );
  INVX0 U5429 ( .INP(n5411), .ZN(n287) );
  OR2X1 U5430 ( .IN1(n4413), .IN2(n3904), .Q(n5411) );
  OR4X1 U5431 ( .IN1(n5412), .IN2(n5413), .IN3(n5414), .IN4(n5415), .Q(WX7119)
         );
  AND2X1 U5432 ( .IN1(n3536), .IN2(n5416), .Q(n5415) );
  AND2X1 U5433 ( .IN1(n5146), .IN2(n3622), .Q(n5414) );
  XOR3X1 U5434 ( .IN1(n2920), .IN2(TM1), .IN3(n5417), .Q(n5146) );
  XOR3X1 U5435 ( .IN1(test_so74), .IN2(n7116), .IN3(WX8541), .Q(n5417) );
  AND2X1 U5436 ( .IN1(n3606), .IN2(CRC_OUT_4_26), .Q(n5413) );
  AND2X1 U5437 ( .IN1(n286), .IN2(n3576), .Q(n5412) );
  INVX0 U5438 ( .INP(n5418), .ZN(n286) );
  OR2X1 U5439 ( .IN1(n4412), .IN2(n3905), .Q(n5418) );
  OR4X1 U5440 ( .IN1(n5419), .IN2(n5420), .IN3(n5421), .IN4(n5422), .Q(WX7117)
         );
  AND2X1 U5441 ( .IN1(n5423), .IN2(n3534), .Q(n5422) );
  AND2X1 U5442 ( .IN1(n3641), .IN2(n5153), .Q(n5421) );
  XOR3X1 U5443 ( .IN1(n2921), .IN2(n3514), .IN3(n5424), .Q(n5153) );
  XOR3X1 U5444 ( .IN1(n7117), .IN2(n3258), .IN3(WX8539), .Q(n5424) );
  AND2X1 U5445 ( .IN1(n3606), .IN2(CRC_OUT_4_27), .Q(n5420) );
  AND2X1 U5446 ( .IN1(n285), .IN2(n3576), .Q(n5419) );
  INVX0 U5447 ( .INP(n5425), .ZN(n285) );
  OR2X1 U5448 ( .IN1(n4412), .IN2(n3906), .Q(n5425) );
  OR4X1 U5449 ( .IN1(n5426), .IN2(n5427), .IN3(n5428), .IN4(n5429), .Q(WX7115)
         );
  AND2X1 U5450 ( .IN1(n3536), .IN2(n5430), .Q(n5429) );
  AND2X1 U5451 ( .IN1(n5160), .IN2(n3622), .Q(n5428) );
  XOR3X1 U5452 ( .IN1(n2923), .IN2(TM1), .IN3(n5431), .Q(n5160) );
  XNOR3X1 U5453 ( .IN1(test_so72), .IN2(n7118), .IN3(n3257), .Q(n5431) );
  AND2X1 U5454 ( .IN1(n3606), .IN2(CRC_OUT_4_28), .Q(n5427) );
  AND2X1 U5455 ( .IN1(n284), .IN2(n3576), .Q(n5426) );
  INVX0 U5456 ( .INP(n5432), .ZN(n284) );
  OR2X1 U5457 ( .IN1(n4412), .IN2(n3907), .Q(n5432) );
  OR4X1 U5458 ( .IN1(n5433), .IN2(n5434), .IN3(n5435), .IN4(n5436), .Q(WX7113)
         );
  AND2X1 U5459 ( .IN1(n3536), .IN2(n5437), .Q(n5436) );
  AND2X1 U5460 ( .IN1(n3641), .IN2(n5167), .Q(n5435) );
  XOR3X1 U5461 ( .IN1(n2924), .IN2(n3518), .IN3(n5438), .Q(n5167) );
  XOR3X1 U5462 ( .IN1(n7119), .IN2(n3256), .IN3(WX8535), .Q(n5438) );
  AND2X1 U5463 ( .IN1(test_so66), .IN2(n3587), .Q(n5434) );
  AND2X1 U5464 ( .IN1(n283), .IN2(n3576), .Q(n5433) );
  INVX0 U5465 ( .INP(n5439), .ZN(n283) );
  OR2X1 U5466 ( .IN1(n4412), .IN2(n3908), .Q(n5439) );
  OR4X1 U5467 ( .IN1(n5440), .IN2(n5441), .IN3(n5442), .IN4(n5443), .Q(WX7111)
         );
  AND2X1 U5468 ( .IN1(n3536), .IN2(n5444), .Q(n5443) );
  AND2X1 U5469 ( .IN1(n5174), .IN2(n3622), .Q(n5442) );
  XOR3X1 U5470 ( .IN1(n2926), .IN2(TM1), .IN3(n5445), .Q(n5174) );
  XNOR3X1 U5471 ( .IN1(test_so70), .IN2(n7120), .IN3(n3255), .Q(n5445) );
  AND2X1 U5472 ( .IN1(n3606), .IN2(CRC_OUT_4_30), .Q(n5441) );
  AND2X1 U5473 ( .IN1(n282), .IN2(n3576), .Q(n5440) );
  INVX0 U5474 ( .INP(n5446), .ZN(n282) );
  OR2X1 U5475 ( .IN1(n4412), .IN2(n3909), .Q(n5446) );
  OR4X1 U5476 ( .IN1(n5447), .IN2(n5448), .IN3(n5449), .IN4(n5450), .Q(WX7109)
         );
  AND2X1 U5477 ( .IN1(n3536), .IN2(n5451), .Q(n5450) );
  AND2X1 U5478 ( .IN1(n3641), .IN2(n5181), .Q(n5449) );
  XOR3X1 U5479 ( .IN1(n2835), .IN2(n3516), .IN3(n5452), .Q(n5181) );
  XOR3X1 U5480 ( .IN1(n7121), .IN2(n3254), .IN3(WX8531), .Q(n5452) );
  AND2X1 U5481 ( .IN1(n2245), .IN2(WX6950), .Q(n5448) );
  AND2X1 U5482 ( .IN1(n3606), .IN2(CRC_OUT_4_31), .Q(n5447) );
  OR4X1 U5483 ( .IN1(n5453), .IN2(n5454), .IN3(n5455), .IN4(n5456), .Q(WX706)
         );
  AND2X1 U5484 ( .IN1(n3536), .IN2(n5457), .Q(n5456) );
  AND2X1 U5485 ( .IN1(n5458), .IN2(n3622), .Q(n5455) );
  AND2X1 U5486 ( .IN1(n3606), .IN2(CRC_OUT_9_0), .Q(n5454) );
  AND2X1 U5487 ( .IN1(WX544), .IN2(n3576), .Q(n5453) );
  OR4X1 U5488 ( .IN1(n5459), .IN2(n5460), .IN3(n5461), .IN4(n5462), .Q(WX704)
         );
  AND2X1 U5489 ( .IN1(n3536), .IN2(n5463), .Q(n5462) );
  AND2X1 U5490 ( .IN1(n3641), .IN2(n5464), .Q(n5461) );
  AND2X1 U5491 ( .IN1(test_so9), .IN2(n3588), .Q(n5460) );
  AND2X1 U5492 ( .IN1(WX542), .IN2(n3576), .Q(n5459) );
  OR4X1 U5493 ( .IN1(n5465), .IN2(n5466), .IN3(n5467), .IN4(n5468), .Q(WX702)
         );
  AND2X1 U5494 ( .IN1(n5469), .IN2(n3532), .Q(n5468) );
  AND2X1 U5495 ( .IN1(n3641), .IN2(n5470), .Q(n5467) );
  AND2X1 U5496 ( .IN1(n3606), .IN2(CRC_OUT_9_2), .Q(n5466) );
  AND2X1 U5497 ( .IN1(WX540), .IN2(n3576), .Q(n5465) );
  AND2X1 U5498 ( .IN1(n3504), .IN2(n4351), .Q(WX7011) );
  OR4X1 U5499 ( .IN1(n5471), .IN2(n5472), .IN3(n5473), .IN4(n5474), .Q(WX700)
         );
  AND2X1 U5500 ( .IN1(n3536), .IN2(n5475), .Q(n5474) );
  AND2X1 U5501 ( .IN1(n3641), .IN2(n5476), .Q(n5473) );
  AND2X1 U5502 ( .IN1(n3606), .IN2(CRC_OUT_9_3), .Q(n5472) );
  AND2X1 U5503 ( .IN1(WX538), .IN2(n3576), .Q(n5471) );
  AND2X1 U5504 ( .IN1(n5183), .IN2(n8443), .Q(WX6999) );
  OR4X1 U5505 ( .IN1(n5477), .IN2(n5478), .IN3(n5479), .IN4(n5480), .Q(WX698)
         );
  AND2X1 U5506 ( .IN1(n3536), .IN2(n5481), .Q(n5480) );
  AND2X1 U5507 ( .IN1(n5482), .IN2(n3622), .Q(n5479) );
  AND2X1 U5508 ( .IN1(n3606), .IN2(CRC_OUT_9_4), .Q(n5478) );
  AND2X1 U5509 ( .IN1(WX536), .IN2(n3576), .Q(n5477) );
  OR4X1 U5510 ( .IN1(n5483), .IN2(n5484), .IN3(n5485), .IN4(n5486), .Q(WX696)
         );
  AND2X1 U5511 ( .IN1(n3536), .IN2(n5487), .Q(n5486) );
  AND2X1 U5512 ( .IN1(n3642), .IN2(n5488), .Q(n5485) );
  AND2X1 U5513 ( .IN1(n3606), .IN2(CRC_OUT_9_5), .Q(n5484) );
  AND2X1 U5514 ( .IN1(WX534), .IN2(n3576), .Q(n5483) );
  OR4X1 U5515 ( .IN1(n5489), .IN2(n5490), .IN3(n5491), .IN4(n5492), .Q(WX694)
         );
  AND2X1 U5516 ( .IN1(n5493), .IN2(n3532), .Q(n5492) );
  AND2X1 U5517 ( .IN1(n3642), .IN2(n5494), .Q(n5491) );
  AND2X1 U5518 ( .IN1(n3606), .IN2(CRC_OUT_9_6), .Q(n5490) );
  AND2X1 U5519 ( .IN1(WX532), .IN2(n3575), .Q(n5489) );
  OR4X1 U5520 ( .IN1(n5495), .IN2(n5496), .IN3(n5497), .IN4(n5498), .Q(WX692)
         );
  AND2X1 U5521 ( .IN1(n3536), .IN2(n5499), .Q(n5498) );
  AND2X1 U5522 ( .IN1(n3642), .IN2(n5500), .Q(n5497) );
  AND2X1 U5523 ( .IN1(n3606), .IN2(CRC_OUT_9_7), .Q(n5496) );
  AND2X1 U5524 ( .IN1(WX530), .IN2(n3575), .Q(n5495) );
  OR4X1 U5525 ( .IN1(n5501), .IN2(n5502), .IN3(n5503), .IN4(n5504), .Q(WX690)
         );
  AND2X1 U5526 ( .IN1(n3537), .IN2(n5505), .Q(n5504) );
  AND2X1 U5527 ( .IN1(n3642), .IN2(n5506), .Q(n5503) );
  AND2X1 U5528 ( .IN1(n3607), .IN2(CRC_OUT_9_8), .Q(n5502) );
  AND2X1 U5529 ( .IN1(WX528), .IN2(n3575), .Q(n5501) );
  OR4X1 U5530 ( .IN1(n5507), .IN2(n5508), .IN3(n5509), .IN4(n5510), .Q(WX688)
         );
  AND2X1 U5531 ( .IN1(n3537), .IN2(n5511), .Q(n5510) );
  AND2X1 U5532 ( .IN1(n3642), .IN2(n5512), .Q(n5509) );
  AND2X1 U5533 ( .IN1(n3607), .IN2(CRC_OUT_9_9), .Q(n5508) );
  AND2X1 U5534 ( .IN1(WX526), .IN2(n3575), .Q(n5507) );
  OR4X1 U5535 ( .IN1(n5513), .IN2(n5514), .IN3(n5515), .IN4(n5516), .Q(WX686)
         );
  AND2X1 U5536 ( .IN1(n5517), .IN2(n3531), .Q(n5516) );
  AND2X1 U5537 ( .IN1(n5518), .IN2(n3621), .Q(n5515) );
  AND2X1 U5538 ( .IN1(n3607), .IN2(CRC_OUT_9_10), .Q(n5514) );
  AND2X1 U5539 ( .IN1(WX524), .IN2(n3575), .Q(n5513) );
  OR4X1 U5540 ( .IN1(n5519), .IN2(n5520), .IN3(n5521), .IN4(n5522), .Q(WX684)
         );
  AND2X1 U5541 ( .IN1(n3537), .IN2(n5523), .Q(n5522) );
  AND2X1 U5542 ( .IN1(n3642), .IN2(n5524), .Q(n5521) );
  AND2X1 U5543 ( .IN1(n3607), .IN2(CRC_OUT_9_11), .Q(n5520) );
  AND2X1 U5544 ( .IN1(WX522), .IN2(n3575), .Q(n5519) );
  OR4X1 U5545 ( .IN1(n5525), .IN2(n5526), .IN3(n5527), .IN4(n5528), .Q(WX682)
         );
  AND2X1 U5546 ( .IN1(n3537), .IN2(n5529), .Q(n5528) );
  AND2X1 U5547 ( .IN1(n3642), .IN2(n5530), .Q(n5527) );
  AND2X1 U5548 ( .IN1(n3607), .IN2(CRC_OUT_9_12), .Q(n5526) );
  AND2X1 U5549 ( .IN1(WX520), .IN2(n3575), .Q(n5525) );
  OR4X1 U5550 ( .IN1(n5531), .IN2(n5532), .IN3(n5533), .IN4(n5534), .Q(WX680)
         );
  AND2X1 U5551 ( .IN1(n3537), .IN2(n5535), .Q(n5534) );
  AND2X1 U5552 ( .IN1(n3642), .IN2(n5536), .Q(n5533) );
  AND2X1 U5553 ( .IN1(n3607), .IN2(CRC_OUT_9_13), .Q(n5532) );
  AND2X1 U5554 ( .IN1(WX518), .IN2(n3575), .Q(n5531) );
  OR4X1 U5555 ( .IN1(n5537), .IN2(n5538), .IN3(n5539), .IN4(n5540), .Q(WX678)
         );
  AND2X1 U5556 ( .IN1(n3537), .IN2(n5541), .Q(n5540) );
  AND2X1 U5557 ( .IN1(n5542), .IN2(n3621), .Q(n5539) );
  AND2X1 U5558 ( .IN1(n3607), .IN2(CRC_OUT_9_14), .Q(n5538) );
  AND2X1 U5559 ( .IN1(WX516), .IN2(n3575), .Q(n5537) );
  OR4X1 U5560 ( .IN1(n5543), .IN2(n5544), .IN3(n5545), .IN4(n5546), .Q(WX676)
         );
  AND2X1 U5561 ( .IN1(n3537), .IN2(n5547), .Q(n5546) );
  AND2X1 U5562 ( .IN1(n3642), .IN2(n5548), .Q(n5545) );
  AND2X1 U5563 ( .IN1(n3607), .IN2(CRC_OUT_9_15), .Q(n5544) );
  AND2X1 U5564 ( .IN1(WX514), .IN2(n3575), .Q(n5543) );
  OR4X1 U5565 ( .IN1(n5549), .IN2(n5550), .IN3(n5551), .IN4(n5552), .Q(WX674)
         );
  AND2X1 U5566 ( .IN1(n5553), .IN2(n3531), .Q(n5552) );
  AND2X1 U5567 ( .IN1(n3642), .IN2(n5554), .Q(n5551) );
  AND2X1 U5568 ( .IN1(n3607), .IN2(CRC_OUT_9_16), .Q(n5550) );
  AND2X1 U5569 ( .IN1(WX512), .IN2(n3575), .Q(n5549) );
  OR4X1 U5570 ( .IN1(n5555), .IN2(n5556), .IN3(n5557), .IN4(n5558), .Q(WX672)
         );
  AND2X1 U5571 ( .IN1(n3537), .IN2(n5559), .Q(n5558) );
  AND2X1 U5572 ( .IN1(n3642), .IN2(n5560), .Q(n5557) );
  AND2X1 U5573 ( .IN1(n3607), .IN2(CRC_OUT_9_17), .Q(n5556) );
  AND2X1 U5574 ( .IN1(WX510), .IN2(n3575), .Q(n5555) );
  OR4X1 U5575 ( .IN1(n5561), .IN2(n5562), .IN3(n5563), .IN4(n5564), .Q(WX670)
         );
  AND2X1 U5576 ( .IN1(n3537), .IN2(n5565), .Q(n5564) );
  AND2X1 U5577 ( .IN1(n5566), .IN2(n3621), .Q(n5563) );
  AND2X1 U5578 ( .IN1(n3607), .IN2(CRC_OUT_9_18), .Q(n5562) );
  AND2X1 U5579 ( .IN1(WX508), .IN2(n3574), .Q(n5561) );
  OR4X1 U5580 ( .IN1(n5567), .IN2(n5568), .IN3(n5569), .IN4(n5570), .Q(WX668)
         );
  AND2X1 U5581 ( .IN1(n3537), .IN2(n5571), .Q(n5570) );
  AND2X1 U5582 ( .IN1(n3642), .IN2(n5572), .Q(n5569) );
  AND2X1 U5583 ( .IN1(test_so10), .IN2(n3587), .Q(n5568) );
  AND2X1 U5584 ( .IN1(WX506), .IN2(n3574), .Q(n5567) );
  OR4X1 U5585 ( .IN1(n5573), .IN2(n5574), .IN3(n5575), .IN4(n5576), .Q(WX666)
         );
  AND2X1 U5586 ( .IN1(n5577), .IN2(n3530), .Q(n5576) );
  AND2X1 U5587 ( .IN1(n3642), .IN2(n5578), .Q(n5575) );
  AND2X1 U5588 ( .IN1(n3607), .IN2(CRC_OUT_9_20), .Q(n5574) );
  AND2X1 U5589 ( .IN1(WX504), .IN2(n3574), .Q(n5573) );
  OR4X1 U5590 ( .IN1(n5579), .IN2(n5580), .IN3(n5581), .IN4(n5582), .Q(WX664)
         );
  AND2X1 U5591 ( .IN1(n3537), .IN2(n5583), .Q(n5582) );
  AND2X1 U5592 ( .IN1(n3643), .IN2(n5584), .Q(n5581) );
  AND2X1 U5593 ( .IN1(n3607), .IN2(CRC_OUT_9_21), .Q(n5580) );
  AND2X1 U5594 ( .IN1(WX502), .IN2(n3574), .Q(n5579) );
  OR4X1 U5595 ( .IN1(n5585), .IN2(n5586), .IN3(n5587), .IN4(n5588), .Q(WX662)
         );
  AND2X1 U5596 ( .IN1(n3537), .IN2(n5589), .Q(n5588) );
  AND2X1 U5597 ( .IN1(n5590), .IN2(n3621), .Q(n5587) );
  AND2X1 U5598 ( .IN1(n3608), .IN2(CRC_OUT_9_22), .Q(n5586) );
  AND2X1 U5599 ( .IN1(WX500), .IN2(n3574), .Q(n5585) );
  OR4X1 U5600 ( .IN1(n5591), .IN2(n5592), .IN3(n5593), .IN4(n5594), .Q(WX660)
         );
  AND2X1 U5601 ( .IN1(n3537), .IN2(n5595), .Q(n5594) );
  AND2X1 U5602 ( .IN1(n3643), .IN2(n5596), .Q(n5593) );
  AND2X1 U5603 ( .IN1(n3608), .IN2(CRC_OUT_9_23), .Q(n5592) );
  AND2X1 U5604 ( .IN1(WX498), .IN2(n3574), .Q(n5591) );
  OR4X1 U5605 ( .IN1(n5597), .IN2(n5598), .IN3(n5599), .IN4(n5600), .Q(WX658)
         );
  AND2X1 U5606 ( .IN1(n5601), .IN2(n3530), .Q(n5600) );
  AND2X1 U5607 ( .IN1(n3643), .IN2(n5602), .Q(n5599) );
  AND2X1 U5608 ( .IN1(n3608), .IN2(CRC_OUT_9_24), .Q(n5598) );
  AND2X1 U5609 ( .IN1(WX496), .IN2(n3574), .Q(n5597) );
  OR4X1 U5610 ( .IN1(n5603), .IN2(n5604), .IN3(n5605), .IN4(n5606), .Q(WX656)
         );
  AND2X1 U5611 ( .IN1(n3538), .IN2(n5607), .Q(n5606) );
  AND2X1 U5612 ( .IN1(n3643), .IN2(n5608), .Q(n5605) );
  AND2X1 U5613 ( .IN1(n3608), .IN2(CRC_OUT_9_25), .Q(n5604) );
  AND2X1 U5614 ( .IN1(WX494), .IN2(n3574), .Q(n5603) );
  OR4X1 U5615 ( .IN1(n5609), .IN2(n5610), .IN3(n5611), .IN4(n5612), .Q(WX654)
         );
  AND2X1 U5616 ( .IN1(n3538), .IN2(n5613), .Q(n5612) );
  AND2X1 U5617 ( .IN1(n3643), .IN2(n5614), .Q(n5611) );
  AND2X1 U5618 ( .IN1(n3608), .IN2(CRC_OUT_9_26), .Q(n5610) );
  AND2X1 U5619 ( .IN1(WX492), .IN2(n3574), .Q(n5609) );
  OR4X1 U5620 ( .IN1(n5615), .IN2(n5616), .IN3(n5617), .IN4(n5618), .Q(WX652)
         );
  AND2X1 U5621 ( .IN1(n3538), .IN2(n5619), .Q(n5618) );
  AND2X1 U5622 ( .IN1(n3643), .IN2(n5620), .Q(n5617) );
  AND2X1 U5623 ( .IN1(n3608), .IN2(CRC_OUT_9_27), .Q(n5616) );
  AND2X1 U5624 ( .IN1(WX490), .IN2(n3574), .Q(n5615) );
  OR4X1 U5625 ( .IN1(n5621), .IN2(n5622), .IN3(n5623), .IN4(n5624), .Q(WX650)
         );
  AND2X1 U5626 ( .IN1(n5625), .IN2(n3528), .Q(n5624) );
  AND2X1 U5627 ( .IN1(n5626), .IN2(n3621), .Q(n5623) );
  AND2X1 U5628 ( .IN1(n3608), .IN2(CRC_OUT_9_28), .Q(n5622) );
  AND2X1 U5629 ( .IN1(WX488), .IN2(n3574), .Q(n5621) );
  AND2X1 U5630 ( .IN1(n5627), .IN2(n4352), .Q(WX6498) );
  XOR2X1 U5631 ( .IN1(CRC_OUT_5_30), .IN2(n3308), .Q(n5627) );
  AND2X1 U5632 ( .IN1(n5628), .IN2(n4352), .Q(WX6496) );
  XOR2X1 U5633 ( .IN1(CRC_OUT_5_29), .IN2(n3309), .Q(n5628) );
  AND2X1 U5634 ( .IN1(n5629), .IN2(n4352), .Q(WX6494) );
  XOR2X1 U5635 ( .IN1(CRC_OUT_5_28), .IN2(n3310), .Q(n5629) );
  AND2X1 U5636 ( .IN1(n5630), .IN2(n4352), .Q(WX6492) );
  XOR2X1 U5637 ( .IN1(CRC_OUT_5_27), .IN2(n3311), .Q(n5630) );
  AND2X1 U5638 ( .IN1(n5631), .IN2(n4352), .Q(WX6490) );
  XOR2X1 U5639 ( .IN1(CRC_OUT_5_26), .IN2(n3312), .Q(n5631) );
  AND2X1 U5640 ( .IN1(n5632), .IN2(n4352), .Q(WX6488) );
  XOR2X1 U5641 ( .IN1(CRC_OUT_5_25), .IN2(n3313), .Q(n5632) );
  AND2X1 U5642 ( .IN1(n5633), .IN2(n4352), .Q(WX6486) );
  XOR2X1 U5643 ( .IN1(CRC_OUT_5_24), .IN2(n3314), .Q(n5633) );
  AND2X1 U5644 ( .IN1(n5634), .IN2(n5183), .Q(WX6484) );
  INVX0 U5645 ( .INP(n5635), .ZN(n5183) );
  OR2X1 U5646 ( .IN1(Tj_Trigger), .IN2(n4410), .Q(n5635) );
  XOR2X1 U5647 ( .IN1(CRC_OUT_5_23), .IN2(n3315), .Q(n5634) );
  AND2X1 U5648 ( .IN1(n5636), .IN2(n4352), .Q(WX6482) );
  XOR2X1 U5649 ( .IN1(CRC_OUT_5_22), .IN2(n3316), .Q(n5636) );
  AND2X1 U5650 ( .IN1(n5637), .IN2(n4352), .Q(WX6480) );
  XOR2X1 U5651 ( .IN1(CRC_OUT_5_21), .IN2(n3317), .Q(n5637) );
  OR4X1 U5652 ( .IN1(n5638), .IN2(n5639), .IN3(n5640), .IN4(n5641), .Q(WX648)
         );
  AND2X1 U5653 ( .IN1(n3538), .IN2(n5642), .Q(n5641) );
  AND2X1 U5654 ( .IN1(n3643), .IN2(n5643), .Q(n5640) );
  AND2X1 U5655 ( .IN1(n3608), .IN2(CRC_OUT_9_29), .Q(n5639) );
  AND2X1 U5656 ( .IN1(WX486), .IN2(n3574), .Q(n5638) );
  AND2X1 U5657 ( .IN1(n5644), .IN2(n4353), .Q(WX6478) );
  XOR2X1 U5658 ( .IN1(CRC_OUT_5_20), .IN2(n3318), .Q(n5644) );
  AND2X1 U5659 ( .IN1(n5645), .IN2(n4353), .Q(WX6476) );
  XOR2X1 U5660 ( .IN1(CRC_OUT_5_19), .IN2(n3319), .Q(n5645) );
  AND2X1 U5661 ( .IN1(n5646), .IN2(n4353), .Q(WX6474) );
  XOR2X1 U5662 ( .IN1(CRC_OUT_5_18), .IN2(n3320), .Q(n5646) );
  AND2X1 U5663 ( .IN1(n5647), .IN2(n4353), .Q(WX6472) );
  XOR2X1 U5664 ( .IN1(test_so54), .IN2(n3321), .Q(n5647) );
  AND2X1 U5665 ( .IN1(n5648), .IN2(n4353), .Q(WX6470) );
  XOR2X1 U5666 ( .IN1(CRC_OUT_5_16), .IN2(n3322), .Q(n5648) );
  AND2X1 U5667 ( .IN1(n5649), .IN2(n4353), .Q(WX6468) );
  XOR3X1 U5668 ( .IN1(test_so52), .IN2(DFF_959_n1), .IN3(CRC_OUT_5_15), .Q(
        n5649) );
  AND2X1 U5669 ( .IN1(n5650), .IN2(n4353), .Q(WX6466) );
  XOR2X1 U5670 ( .IN1(CRC_OUT_5_14), .IN2(n3323), .Q(n5650) );
  AND2X1 U5671 ( .IN1(n5651), .IN2(n4353), .Q(WX6464) );
  XOR2X1 U5672 ( .IN1(CRC_OUT_5_13), .IN2(n3324), .Q(n5651) );
  AND2X1 U5673 ( .IN1(n5652), .IN2(n4353), .Q(WX6462) );
  XOR2X1 U5674 ( .IN1(CRC_OUT_5_12), .IN2(n3325), .Q(n5652) );
  AND2X1 U5675 ( .IN1(n5653), .IN2(n4354), .Q(WX6460) );
  XOR2X1 U5676 ( .IN1(CRC_OUT_5_11), .IN2(n3326), .Q(n5653) );
  OR4X1 U5677 ( .IN1(n5654), .IN2(n5655), .IN3(n5656), .IN4(n5657), .Q(WX646)
         );
  AND2X1 U5678 ( .IN1(n3554), .IN2(n5658), .Q(n5657) );
  AND2X1 U5679 ( .IN1(n3643), .IN2(n5659), .Q(n5656) );
  AND2X1 U5680 ( .IN1(n3608), .IN2(CRC_OUT_9_30), .Q(n5655) );
  AND2X1 U5681 ( .IN1(WX484), .IN2(n3573), .Q(n5654) );
  AND2X1 U5682 ( .IN1(n5660), .IN2(n4354), .Q(WX6458) );
  XOR3X1 U5683 ( .IN1(n3184), .IN2(DFF_959_n1), .IN3(DFF_938_n1), .Q(n5660) );
  AND2X1 U5684 ( .IN1(n5661), .IN2(n4354), .Q(WX6456) );
  XOR2X1 U5685 ( .IN1(CRC_OUT_5_9), .IN2(n3327), .Q(n5661) );
  AND2X1 U5686 ( .IN1(n5662), .IN2(n4354), .Q(WX6454) );
  XOR2X1 U5687 ( .IN1(CRC_OUT_5_8), .IN2(n3328), .Q(n5662) );
  AND2X1 U5688 ( .IN1(n5663), .IN2(n4354), .Q(WX6452) );
  XOR2X1 U5689 ( .IN1(CRC_OUT_5_7), .IN2(n3329), .Q(n5663) );
  AND2X1 U5690 ( .IN1(n5664), .IN2(n4354), .Q(WX6450) );
  XOR2X1 U5691 ( .IN1(CRC_OUT_5_6), .IN2(n3330), .Q(n5664) );
  AND2X1 U5692 ( .IN1(n5665), .IN2(n4354), .Q(WX6448) );
  XOR2X1 U5693 ( .IN1(CRC_OUT_5_5), .IN2(n3331), .Q(n5665) );
  AND2X1 U5694 ( .IN1(n5666), .IN2(n4354), .Q(WX6446) );
  XOR2X1 U5695 ( .IN1(CRC_OUT_5_4), .IN2(n3332), .Q(n5666) );
  AND2X1 U5696 ( .IN1(n5667), .IN2(n4355), .Q(WX6444) );
  XOR3X1 U5697 ( .IN1(n3185), .IN2(DFF_959_n1), .IN3(DFF_931_n1), .Q(n5667) );
  AND2X1 U5698 ( .IN1(n5668), .IN2(n4355), .Q(WX6442) );
  XOR2X1 U5699 ( .IN1(CRC_OUT_5_2), .IN2(n3333), .Q(n5668) );
  AND2X1 U5700 ( .IN1(n5669), .IN2(n4355), .Q(WX6440) );
  XOR2X1 U5701 ( .IN1(CRC_OUT_5_1), .IN2(n3334), .Q(n5669) );
  OR4X1 U5702 ( .IN1(n5670), .IN2(n5671), .IN3(n5672), .IN4(n5673), .Q(WX644)
         );
  AND2X1 U5703 ( .IN1(n3554), .IN2(n5674), .Q(n5673) );
  AND2X1 U5704 ( .IN1(n3643), .IN2(n5675), .Q(n5672) );
  AND2X1 U5705 ( .IN1(n2245), .IN2(WX485), .Q(n5671) );
  AND2X1 U5706 ( .IN1(n3608), .IN2(CRC_OUT_9_31), .Q(n5670) );
  AND2X1 U5707 ( .IN1(n5676), .IN2(n4355), .Q(WX6438) );
  XOR2X1 U5708 ( .IN1(test_so53), .IN2(n3335), .Q(n5676) );
  AND2X1 U5709 ( .IN1(n5677), .IN2(n4355), .Q(WX6436) );
  XOR2X1 U5710 ( .IN1(n3198), .IN2(CRC_OUT_5_31), .Q(n5677) );
  INVX0 U5711 ( .INP(n5678), .ZN(WX5910) );
  OR2X1 U5712 ( .IN1(n4412), .IN2(n7163), .Q(n5678) );
  INVX0 U5713 ( .INP(n5679), .ZN(WX5908) );
  OR2X1 U5714 ( .IN1(n4412), .IN2(n7164), .Q(n5679) );
  INVX0 U5715 ( .INP(n5680), .ZN(WX5906) );
  OR2X1 U6483 ( .IN1(n4412), .IN2(n7165), .Q(n5680) );
  INVX0 U6484 ( .INP(n5681), .ZN(WX5904) );
  OR2X1 U6485 ( .IN1(n4412), .IN2(n7166), .Q(n5681) );
  INVX0 U6486 ( .INP(n5682), .ZN(WX5902) );
  OR2X1 U6487 ( .IN1(n4412), .IN2(n7167), .Q(n5682) );
  INVX0 U6488 ( .INP(n5683), .ZN(WX5900) );
  OR2X1 U6489 ( .IN1(n4412), .IN2(n7168), .Q(n5683) );
  AND2X1 U6490 ( .IN1(test_so46), .IN2(n4355), .Q(WX5898) );
  INVX0 U6491 ( .INP(n5684), .ZN(WX5896) );
  OR2X1 U6492 ( .IN1(n4412), .IN2(n7170), .Q(n5684) );
  INVX0 U6493 ( .INP(n5685), .ZN(WX5894) );
  OR2X1 U6494 ( .IN1(n4411), .IN2(n7171), .Q(n5685) );
  INVX0 U6495 ( .INP(n5686), .ZN(WX5892) );
  OR2X1 U6496 ( .IN1(n4411), .IN2(n7172), .Q(n5686) );
  INVX0 U6497 ( .INP(n5687), .ZN(WX5890) );
  OR2X1 U6498 ( .IN1(n4411), .IN2(n7173), .Q(n5687) );
  INVX0 U6499 ( .INP(n5688), .ZN(WX5888) );
  OR2X1 U6500 ( .IN1(n4411), .IN2(n7174), .Q(n5688) );
  INVX0 U6501 ( .INP(n5689), .ZN(WX5886) );
  OR2X1 U6502 ( .IN1(n4411), .IN2(n7175), .Q(n5689) );
  INVX0 U6503 ( .INP(n5690), .ZN(WX5884) );
  OR2X1 U6504 ( .IN1(n4411), .IN2(n7176), .Q(n5690) );
  INVX0 U6505 ( .INP(n5691), .ZN(WX5882) );
  OR2X1 U6506 ( .IN1(n4411), .IN2(n7177), .Q(n5691) );
  INVX0 U6507 ( .INP(n5692), .ZN(WX5880) );
  OR2X1 U6508 ( .IN1(n4411), .IN2(n7178), .Q(n5692) );
  OR4X1 U6509 ( .IN1(n5693), .IN2(n5694), .IN3(n5695), .IN4(n5696), .Q(WX5878)
         );
  AND2X1 U6510 ( .IN1(n3554), .IN2(n5697), .Q(n5696) );
  AND2X1 U6511 ( .IN1(n3643), .IN2(n5235), .Q(n5695) );
  XNOR3X1 U6512 ( .IN1(n3197), .IN2(n3102), .IN3(n5698), .Q(n5235) );
  XOR2X1 U6513 ( .IN1(WX7236), .IN2(n7122), .Q(n5698) );
  AND2X1 U6514 ( .IN1(test_so53), .IN2(n3588), .Q(n5694) );
  AND2X1 U6515 ( .IN1(n250), .IN2(n3573), .Q(n5693) );
  INVX0 U6516 ( .INP(n5699), .ZN(n250) );
  OR2X1 U6517 ( .IN1(n4411), .IN2(n3910), .Q(n5699) );
  OR4X1 U6518 ( .IN1(n5700), .IN2(n5701), .IN3(n5702), .IN4(n5703), .Q(WX5876)
         );
  AND2X1 U6519 ( .IN1(n5704), .IN2(n3528), .Q(n5703) );
  AND2X1 U6520 ( .IN1(n3643), .IN2(n5242), .Q(n5702) );
  XNOR3X1 U6521 ( .IN1(n3307), .IN2(n3103), .IN3(n5705), .Q(n5242) );
  XOR2X1 U6522 ( .IN1(WX7234), .IN2(n7123), .Q(n5705) );
  AND2X1 U6523 ( .IN1(n3608), .IN2(CRC_OUT_5_1), .Q(n5701) );
  AND2X1 U6524 ( .IN1(n249), .IN2(n3573), .Q(n5700) );
  INVX0 U6525 ( .INP(n5706), .ZN(n249) );
  OR2X1 U6526 ( .IN1(n4412), .IN2(n3911), .Q(n5706) );
  OR4X1 U6527 ( .IN1(n5707), .IN2(n5708), .IN3(n5709), .IN4(n5710), .Q(WX5874)
         );
  AND2X1 U6528 ( .IN1(n3554), .IN2(n5711), .Q(n5710) );
  AND2X1 U6529 ( .IN1(n3643), .IN2(n5249), .Q(n5709) );
  XNOR3X1 U6530 ( .IN1(n3306), .IN2(n3104), .IN3(n5712), .Q(n5249) );
  XOR2X1 U6531 ( .IN1(WX7232), .IN2(n7124), .Q(n5712) );
  AND2X1 U6532 ( .IN1(n3608), .IN2(CRC_OUT_5_2), .Q(n5708) );
  AND2X1 U6533 ( .IN1(n248), .IN2(n3573), .Q(n5707) );
  INVX0 U6534 ( .INP(n5713), .ZN(n248) );
  OR2X1 U6535 ( .IN1(n4411), .IN2(n3912), .Q(n5713) );
  OR4X1 U6536 ( .IN1(n5714), .IN2(n5715), .IN3(n5716), .IN4(n5717), .Q(WX5872)
         );
  AND2X1 U6537 ( .IN1(n5718), .IN2(n3528), .Q(n5717) );
  AND2X1 U6538 ( .IN1(n3643), .IN2(n5256), .Q(n5716) );
  XNOR3X1 U6539 ( .IN1(n3305), .IN2(n3105), .IN3(n5719), .Q(n5256) );
  XOR2X1 U6540 ( .IN1(WX7230), .IN2(n7125), .Q(n5719) );
  AND2X1 U6541 ( .IN1(n3608), .IN2(CRC_OUT_5_3), .Q(n5715) );
  AND2X1 U6542 ( .IN1(n247), .IN2(n3573), .Q(n5714) );
  INVX0 U6543 ( .INP(n5720), .ZN(n247) );
  OR2X1 U6544 ( .IN1(n4411), .IN2(n3913), .Q(n5720) );
  OR4X1 U6545 ( .IN1(n5721), .IN2(n5722), .IN3(n5723), .IN4(n5724), .Q(WX5870)
         );
  AND2X1 U6546 ( .IN1(n3554), .IN2(n5725), .Q(n5724) );
  AND2X1 U6547 ( .IN1(n5263), .IN2(n3621), .Q(n5723) );
  XOR3X1 U6548 ( .IN1(n3635), .IN2(n3106), .IN3(n5726), .Q(n5263) );
  XOR2X1 U6549 ( .IN1(WX7164), .IN2(test_so64), .Q(n5726) );
  AND2X1 U6550 ( .IN1(n3609), .IN2(CRC_OUT_5_4), .Q(n5722) );
  AND2X1 U6551 ( .IN1(n246), .IN2(n3573), .Q(n5721) );
  INVX0 U6552 ( .INP(n5727), .ZN(n246) );
  OR2X1 U6553 ( .IN1(n4411), .IN2(n3914), .Q(n5727) );
  OR4X1 U6554 ( .IN1(n5728), .IN2(n5729), .IN3(n5730), .IN4(n5731), .Q(WX5868)
         );
  AND2X1 U6555 ( .IN1(n5732), .IN2(n3528), .Q(n5731) );
  AND2X1 U6556 ( .IN1(n3644), .IN2(n5270), .Q(n5730) );
  XNOR3X1 U6557 ( .IN1(n3304), .IN2(n3107), .IN3(n5733), .Q(n5270) );
  XOR2X1 U6558 ( .IN1(WX7226), .IN2(n7126), .Q(n5733) );
  AND2X1 U6559 ( .IN1(n3609), .IN2(CRC_OUT_5_5), .Q(n5729) );
  AND2X1 U6560 ( .IN1(n245), .IN2(n3573), .Q(n5728) );
  INVX0 U6561 ( .INP(n5734), .ZN(n245) );
  OR2X1 U6562 ( .IN1(n4411), .IN2(n3915), .Q(n5734) );
  OR4X1 U6563 ( .IN1(n5735), .IN2(n5736), .IN3(n5737), .IN4(n5738), .Q(WX5866)
         );
  AND2X1 U6564 ( .IN1(n3554), .IN2(n5739), .Q(n5738) );
  AND2X1 U6565 ( .IN1(n5276), .IN2(n3621), .Q(n5737) );
  XOR3X1 U6566 ( .IN1(n3639), .IN2(n3303), .IN3(n5740), .Q(n5276) );
  XOR2X1 U6567 ( .IN1(WX7160), .IN2(test_so62), .Q(n5740) );
  AND2X1 U6568 ( .IN1(n3609), .IN2(CRC_OUT_5_6), .Q(n5736) );
  AND2X1 U6569 ( .IN1(n244), .IN2(n3573), .Q(n5735) );
  INVX0 U6570 ( .INP(n5741), .ZN(n244) );
  OR2X1 U6571 ( .IN1(n4410), .IN2(n3916), .Q(n5741) );
  OR4X1 U6572 ( .IN1(n5742), .IN2(n5743), .IN3(n5744), .IN4(n5745), .Q(WX5864)
         );
  AND2X1 U6573 ( .IN1(n3554), .IN2(n5746), .Q(n5745) );
  AND2X1 U6574 ( .IN1(n3644), .IN2(n5283), .Q(n5744) );
  XNOR3X1 U6575 ( .IN1(n3302), .IN2(n3108), .IN3(n5747), .Q(n5283) );
  XOR2X1 U6576 ( .IN1(WX7222), .IN2(n7127), .Q(n5747) );
  AND2X1 U6577 ( .IN1(n3609), .IN2(CRC_OUT_5_7), .Q(n5743) );
  AND2X1 U6578 ( .IN1(n243), .IN2(n3573), .Q(n5742) );
  INVX0 U6579 ( .INP(n5748), .ZN(n243) );
  OR2X1 U6580 ( .IN1(n4410), .IN2(n3917), .Q(n5748) );
  OR4X1 U6581 ( .IN1(n5749), .IN2(n5750), .IN3(n5751), .IN4(n5752), .Q(WX5862)
         );
  AND2X1 U6582 ( .IN1(n3553), .IN2(n5753), .Q(n5752) );
  AND2X1 U6583 ( .IN1(n5290), .IN2(n3620), .Q(n5751) );
  XOR3X1 U6584 ( .IN1(n3301), .IN2(n3109), .IN3(n5754), .Q(n5290) );
  XOR2X1 U6585 ( .IN1(WX7156), .IN2(test_so60), .Q(n5754) );
  AND2X1 U6586 ( .IN1(n3609), .IN2(CRC_OUT_5_8), .Q(n5750) );
  AND2X1 U6587 ( .IN1(n242), .IN2(n3573), .Q(n5749) );
  INVX0 U6588 ( .INP(n5755), .ZN(n242) );
  OR2X1 U6589 ( .IN1(n4410), .IN2(n3918), .Q(n5755) );
  OR4X1 U6590 ( .IN1(n5756), .IN2(n5757), .IN3(n5758), .IN4(n5759), .Q(WX5860)
         );
  AND2X1 U6591 ( .IN1(n3553), .IN2(n5760), .Q(n5759) );
  AND2X1 U6592 ( .IN1(n3644), .IN2(n5297), .Q(n5758) );
  XNOR3X1 U6593 ( .IN1(n3300), .IN2(n3110), .IN3(n5761), .Q(n5297) );
  XOR2X1 U6594 ( .IN1(WX7218), .IN2(n7128), .Q(n5761) );
  AND2X1 U6595 ( .IN1(n3609), .IN2(CRC_OUT_5_9), .Q(n5757) );
  AND2X1 U6596 ( .IN1(n241), .IN2(n3573), .Q(n5756) );
  INVX0 U6597 ( .INP(n5762), .ZN(n241) );
  OR2X1 U6598 ( .IN1(n4410), .IN2(n3919), .Q(n5762) );
  OR4X1 U6599 ( .IN1(n5763), .IN2(n5764), .IN3(n5765), .IN4(n5766), .Q(WX5858)
         );
  AND2X1 U6600 ( .IN1(n3553), .IN2(n5767), .Q(n5766) );
  AND2X1 U6601 ( .IN1(n5304), .IN2(n3620), .Q(n5765) );
  XOR3X1 U6602 ( .IN1(n3647), .IN2(n3299), .IN3(n5768), .Q(n5304) );
  XOR2X1 U6603 ( .IN1(WX7280), .IN2(test_so58), .Q(n5768) );
  AND2X1 U6604 ( .IN1(n3609), .IN2(CRC_OUT_5_10), .Q(n5764) );
  AND2X1 U6605 ( .IN1(n240), .IN2(n3573), .Q(n5763) );
  INVX0 U6606 ( .INP(n5769), .ZN(n240) );
  OR2X1 U6607 ( .IN1(n4410), .IN2(n3920), .Q(n5769) );
  OR4X1 U6608 ( .IN1(n5770), .IN2(n5771), .IN3(n5772), .IN4(n5773), .Q(WX5856)
         );
  AND2X1 U6609 ( .IN1(n3553), .IN2(n5774), .Q(n5773) );
  AND2X1 U6610 ( .IN1(n3644), .IN2(n5311), .Q(n5772) );
  XNOR3X1 U6611 ( .IN1(n3183), .IN2(n3111), .IN3(n5775), .Q(n5311) );
  XOR2X1 U6612 ( .IN1(WX7214), .IN2(n7129), .Q(n5775) );
  AND2X1 U6613 ( .IN1(n3609), .IN2(CRC_OUT_5_11), .Q(n5771) );
  AND2X1 U6614 ( .IN1(n239), .IN2(n3572), .Q(n5770) );
  INVX0 U6615 ( .INP(n5776), .ZN(n239) );
  OR2X1 U6616 ( .IN1(n4410), .IN2(n3921), .Q(n5776) );
  OR4X1 U6617 ( .IN1(n5777), .IN2(n5778), .IN3(n5779), .IN4(n5780), .Q(WX5854)
         );
  AND2X1 U6618 ( .IN1(n3553), .IN2(n5781), .Q(n5780) );
  AND2X1 U6619 ( .IN1(n3644), .IN2(n5318), .Q(n5779) );
  XNOR3X1 U6620 ( .IN1(n3298), .IN2(n3112), .IN3(n5782), .Q(n5318) );
  XOR2X1 U6621 ( .IN1(WX7212), .IN2(n7130), .Q(n5782) );
  AND2X1 U6622 ( .IN1(n3609), .IN2(CRC_OUT_5_12), .Q(n5778) );
  AND2X1 U6623 ( .IN1(n238), .IN2(n3572), .Q(n5777) );
  INVX0 U6624 ( .INP(n5783), .ZN(n238) );
  OR2X1 U6625 ( .IN1(n4410), .IN2(n3922), .Q(n5783) );
  OR4X1 U6626 ( .IN1(n5784), .IN2(n5785), .IN3(n5786), .IN4(n5787), .Q(WX5852)
         );
  AND2X1 U6627 ( .IN1(n3553), .IN2(n5788), .Q(n5787) );
  AND2X1 U6628 ( .IN1(n3644), .IN2(n5325), .Q(n5786) );
  XNOR3X1 U6629 ( .IN1(n3297), .IN2(n3113), .IN3(n5789), .Q(n5325) );
  XOR2X1 U6630 ( .IN1(WX7210), .IN2(n7131), .Q(n5789) );
  AND2X1 U6631 ( .IN1(n3609), .IN2(CRC_OUT_5_13), .Q(n5785) );
  AND2X1 U6632 ( .IN1(n237), .IN2(n3572), .Q(n5784) );
  INVX0 U6633 ( .INP(n5790), .ZN(n237) );
  OR2X1 U6634 ( .IN1(n4410), .IN2(n3923), .Q(n5790) );
  OR4X1 U6635 ( .IN1(n5791), .IN2(n5792), .IN3(n5793), .IN4(n5794), .Q(WX5850)
         );
  AND2X1 U6636 ( .IN1(n3553), .IN2(n5795), .Q(n5794) );
  AND2X1 U6637 ( .IN1(n3644), .IN2(n5332), .Q(n5793) );
  XNOR3X1 U6638 ( .IN1(n3296), .IN2(n3114), .IN3(n5796), .Q(n5332) );
  XOR2X1 U6639 ( .IN1(WX7208), .IN2(n7132), .Q(n5796) );
  AND2X1 U6640 ( .IN1(n3609), .IN2(CRC_OUT_5_14), .Q(n5792) );
  AND2X1 U6641 ( .IN1(n236), .IN2(n3572), .Q(n5791) );
  INVX0 U6642 ( .INP(n5797), .ZN(n236) );
  OR2X1 U6643 ( .IN1(n4410), .IN2(n3924), .Q(n5797) );
  OR4X1 U6644 ( .IN1(n5798), .IN2(n5799), .IN3(n5800), .IN4(n5801), .Q(WX5848)
         );
  AND2X1 U6645 ( .IN1(n3553), .IN2(n5802), .Q(n5801) );
  AND2X1 U6646 ( .IN1(n3644), .IN2(n5339), .Q(n5800) );
  XNOR3X1 U6647 ( .IN1(n3295), .IN2(n3115), .IN3(n5803), .Q(n5339) );
  XOR2X1 U6648 ( .IN1(WX7206), .IN2(n7133), .Q(n5803) );
  AND2X1 U6649 ( .IN1(n3609), .IN2(CRC_OUT_5_15), .Q(n5799) );
  AND2X1 U6650 ( .IN1(n235), .IN2(n3572), .Q(n5798) );
  INVX0 U6651 ( .INP(n5804), .ZN(n235) );
  OR2X1 U6652 ( .IN1(n4410), .IN2(n3925), .Q(n5804) );
  OR4X1 U6653 ( .IN1(n5805), .IN2(n5806), .IN3(n5807), .IN4(n5808), .Q(WX5846)
         );
  AND2X1 U6654 ( .IN1(n5809), .IN2(n3531), .Q(n5808) );
  AND2X1 U6655 ( .IN1(n3644), .IN2(n5346), .Q(n5807) );
  XOR3X1 U6656 ( .IN1(n2927), .IN2(n3515), .IN3(n5810), .Q(n5346) );
  XOR3X1 U6657 ( .IN1(n7134), .IN2(n3182), .IN3(WX7268), .Q(n5810) );
  AND2X1 U6658 ( .IN1(n3609), .IN2(CRC_OUT_5_16), .Q(n5806) );
  AND2X1 U6659 ( .IN1(n234), .IN2(n3572), .Q(n5805) );
  INVX0 U6660 ( .INP(n5811), .ZN(n234) );
  OR2X1 U6661 ( .IN1(n4410), .IN2(n3926), .Q(n5811) );
  OR4X1 U6662 ( .IN1(n5812), .IN2(n5813), .IN3(n5814), .IN4(n5815), .Q(WX5844)
         );
  AND2X1 U6663 ( .IN1(n3553), .IN2(n5816), .Q(n5815) );
  AND2X1 U6664 ( .IN1(n3644), .IN2(n5353), .Q(n5814) );
  XOR3X1 U6665 ( .IN1(n2929), .IN2(n3514), .IN3(n5817), .Q(n5353) );
  XOR3X1 U6666 ( .IN1(n7135), .IN2(n3294), .IN3(WX7266), .Q(n5817) );
  AND2X1 U6667 ( .IN1(test_so54), .IN2(n3587), .Q(n5813) );
  AND2X1 U6668 ( .IN1(n233), .IN2(n3572), .Q(n5812) );
  INVX0 U6669 ( .INP(n5818), .ZN(n233) );
  OR2X1 U6670 ( .IN1(n4416), .IN2(n3927), .Q(n5818) );
  OR4X1 U6671 ( .IN1(n5819), .IN2(n5820), .IN3(n5821), .IN4(n5822), .Q(WX5842)
         );
  AND2X1 U6672 ( .IN1(n5823), .IN2(n3531), .Q(n5822) );
  AND2X1 U6673 ( .IN1(n3644), .IN2(n5360), .Q(n5821) );
  XOR3X1 U6674 ( .IN1(n2931), .IN2(n3518), .IN3(n5824), .Q(n5360) );
  XOR3X1 U6675 ( .IN1(n7136), .IN2(n3293), .IN3(WX7264), .Q(n5824) );
  AND2X1 U6676 ( .IN1(n3610), .IN2(CRC_OUT_5_18), .Q(n5820) );
  AND2X1 U6677 ( .IN1(n232), .IN2(n3572), .Q(n5819) );
  INVX0 U6678 ( .INP(n5825), .ZN(n232) );
  OR2X1 U6679 ( .IN1(n4429), .IN2(n3928), .Q(n5825) );
  OR4X1 U6680 ( .IN1(n5826), .IN2(n5827), .IN3(n5828), .IN4(n5829), .Q(WX5840)
         );
  AND2X1 U6681 ( .IN1(n3553), .IN2(n5830), .Q(n5829) );
  AND2X1 U6682 ( .IN1(n3644), .IN2(n5367), .Q(n5828) );
  XOR3X1 U6683 ( .IN1(n2933), .IN2(n3516), .IN3(n5831), .Q(n5367) );
  XOR3X1 U6684 ( .IN1(n7137), .IN2(n3292), .IN3(WX7262), .Q(n5831) );
  AND2X1 U6685 ( .IN1(n3610), .IN2(CRC_OUT_5_19), .Q(n5827) );
  AND2X1 U6686 ( .IN1(n231), .IN2(n3572), .Q(n5826) );
  INVX0 U6687 ( .INP(n5832), .ZN(n231) );
  OR2X1 U6688 ( .IN1(n4429), .IN2(n3929), .Q(n5832) );
  OR4X1 U6689 ( .IN1(n5833), .IN2(n5834), .IN3(n5835), .IN4(n5836), .Q(WX5838)
         );
  AND2X1 U6690 ( .IN1(n5837), .IN2(n3531), .Q(n5836) );
  AND2X1 U6691 ( .IN1(n3644), .IN2(n5374), .Q(n5835) );
  XOR3X1 U6692 ( .IN1(n2935), .IN2(n3515), .IN3(n5838), .Q(n5374) );
  XOR3X1 U6693 ( .IN1(n7138), .IN2(n3291), .IN3(WX7260), .Q(n5838) );
  AND2X1 U6694 ( .IN1(n3610), .IN2(CRC_OUT_5_20), .Q(n5834) );
  AND2X1 U6695 ( .IN1(n230), .IN2(n3572), .Q(n5833) );
  INVX0 U6696 ( .INP(n5839), .ZN(n230) );
  OR2X1 U6697 ( .IN1(n4429), .IN2(n3930), .Q(n5839) );
  OR4X1 U6698 ( .IN1(n5840), .IN2(n5841), .IN3(n5842), .IN4(n5843), .Q(WX5836)
         );
  AND2X1 U6699 ( .IN1(n3553), .IN2(n5844), .Q(n5843) );
  AND2X1 U6700 ( .IN1(n5381), .IN2(n3620), .Q(n5842) );
  XOR3X1 U6701 ( .IN1(n2937), .IN2(TM1), .IN3(n5845), .Q(n5381) );
  XOR3X1 U6702 ( .IN1(test_so63), .IN2(n7139), .IN3(WX7258), .Q(n5845) );
  AND2X1 U6703 ( .IN1(n3594), .IN2(CRC_OUT_5_21), .Q(n5841) );
  AND2X1 U6704 ( .IN1(n229), .IN2(n3572), .Q(n5840) );
  INVX0 U6705 ( .INP(n5846), .ZN(n229) );
  OR2X1 U6706 ( .IN1(n4429), .IN2(n3931), .Q(n5846) );
  OR4X1 U6707 ( .IN1(n5847), .IN2(n5848), .IN3(n5849), .IN4(n5850), .Q(WX5834)
         );
  AND2X1 U6708 ( .IN1(n5851), .IN2(n3531), .Q(n5850) );
  AND2X1 U6709 ( .IN1(n3645), .IN2(n5388), .Q(n5849) );
  XOR3X1 U6710 ( .IN1(n2938), .IN2(n3514), .IN3(n5852), .Q(n5388) );
  XOR3X1 U6711 ( .IN1(n7140), .IN2(n3290), .IN3(WX7256), .Q(n5852) );
  AND2X1 U6712 ( .IN1(n3588), .IN2(CRC_OUT_5_22), .Q(n5848) );
  AND2X1 U6713 ( .IN1(n228), .IN2(n3572), .Q(n5847) );
  INVX0 U6714 ( .INP(n5853), .ZN(n228) );
  OR2X1 U6715 ( .IN1(n4430), .IN2(n3932), .Q(n5853) );
  OR4X1 U6716 ( .IN1(n5854), .IN2(n5855), .IN3(n5856), .IN4(n5857), .Q(WX5832)
         );
  AND2X1 U6717 ( .IN1(n3553), .IN2(n5858), .Q(n5857) );
  AND2X1 U6718 ( .IN1(n5395), .IN2(n3620), .Q(n5856) );
  XOR3X1 U6719 ( .IN1(n2940), .IN2(TM1), .IN3(n5859), .Q(n5395) );
  XNOR3X1 U6720 ( .IN1(test_so61), .IN2(n7141), .IN3(n3289), .Q(n5859) );
  AND2X1 U6721 ( .IN1(n3590), .IN2(CRC_OUT_5_23), .Q(n5855) );
  AND2X1 U6722 ( .IN1(n227), .IN2(n3571), .Q(n5854) );
  INVX0 U6723 ( .INP(n5860), .ZN(n227) );
  OR2X1 U6724 ( .IN1(n4430), .IN2(n3933), .Q(n5860) );
  OR4X1 U6725 ( .IN1(n5861), .IN2(n5862), .IN3(n5863), .IN4(n5864), .Q(WX5830)
         );
  AND2X1 U6726 ( .IN1(n3553), .IN2(n5865), .Q(n5864) );
  AND2X1 U6727 ( .IN1(n3645), .IN2(n5402), .Q(n5863) );
  XOR3X1 U6728 ( .IN1(n2941), .IN2(n3518), .IN3(n5866), .Q(n5402) );
  XOR3X1 U6729 ( .IN1(n7142), .IN2(n3288), .IN3(WX7252), .Q(n5866) );
  AND2X1 U6730 ( .IN1(n3588), .IN2(CRC_OUT_5_24), .Q(n5862) );
  AND2X1 U6731 ( .IN1(n226), .IN2(n3571), .Q(n5861) );
  INVX0 U6732 ( .INP(n5867), .ZN(n226) );
  OR2X1 U6733 ( .IN1(n4430), .IN2(n3934), .Q(n5867) );
  OR4X1 U6734 ( .IN1(n5868), .IN2(n5869), .IN3(n5870), .IN4(n5871), .Q(WX5828)
         );
  AND2X1 U6735 ( .IN1(n3552), .IN2(n5872), .Q(n5871) );
  AND2X1 U6736 ( .IN1(n5409), .IN2(n3620), .Q(n5870) );
  XOR3X1 U6737 ( .IN1(n2943), .IN2(TM1), .IN3(n5873), .Q(n5409) );
  XNOR3X1 U6738 ( .IN1(test_so59), .IN2(n7143), .IN3(n3287), .Q(n5873) );
  AND2X1 U6739 ( .IN1(n3589), .IN2(CRC_OUT_5_25), .Q(n5869) );
  AND2X1 U6740 ( .IN1(n225), .IN2(n3571), .Q(n5868) );
  INVX0 U6741 ( .INP(n5874), .ZN(n225) );
  OR2X1 U6742 ( .IN1(n4430), .IN2(n3935), .Q(n5874) );
  OR4X1 U6743 ( .IN1(n5875), .IN2(n5876), .IN3(n5877), .IN4(n5878), .Q(WX5826)
         );
  AND2X1 U6744 ( .IN1(n3552), .IN2(n5879), .Q(n5878) );
  AND2X1 U6745 ( .IN1(n3645), .IN2(n5416), .Q(n5877) );
  XOR3X1 U6746 ( .IN1(n2944), .IN2(n3516), .IN3(n5880), .Q(n5416) );
  XOR3X1 U6747 ( .IN1(n7144), .IN2(n3286), .IN3(WX7248), .Q(n5880) );
  AND2X1 U6748 ( .IN1(n3588), .IN2(CRC_OUT_5_26), .Q(n5876) );
  AND2X1 U6749 ( .IN1(n224), .IN2(n3571), .Q(n5875) );
  INVX0 U6750 ( .INP(n5881), .ZN(n224) );
  OR2X1 U6751 ( .IN1(n4430), .IN2(n3936), .Q(n5881) );
  OR4X1 U6752 ( .IN1(n5882), .IN2(n5883), .IN3(n5884), .IN4(n5885), .Q(WX5824)
         );
  AND2X1 U6753 ( .IN1(n3552), .IN2(n5886), .Q(n5885) );
  AND2X1 U6754 ( .IN1(n5423), .IN2(n3620), .Q(n5884) );
  XOR3X1 U6755 ( .IN1(n2946), .IN2(TM1), .IN3(n5887), .Q(n5423) );
  XNOR3X1 U6756 ( .IN1(test_so57), .IN2(n7145), .IN3(n3285), .Q(n5887) );
  AND2X1 U6757 ( .IN1(n3589), .IN2(CRC_OUT_5_27), .Q(n5883) );
  AND2X1 U6758 ( .IN1(n223), .IN2(n3571), .Q(n5882) );
  INVX0 U6759 ( .INP(n5888), .ZN(n223) );
  OR2X1 U6760 ( .IN1(n4430), .IN2(n3937), .Q(n5888) );
  OR4X1 U6761 ( .IN1(n5889), .IN2(n5890), .IN3(n5891), .IN4(n5892), .Q(WX5822)
         );
  AND2X1 U6762 ( .IN1(n3552), .IN2(n5893), .Q(n5892) );
  AND2X1 U6763 ( .IN1(n3645), .IN2(n5430), .Q(n5891) );
  XOR3X1 U6764 ( .IN1(n2947), .IN2(n3515), .IN3(n5894), .Q(n5430) );
  XOR3X1 U6765 ( .IN1(n7146), .IN2(n3284), .IN3(WX7244), .Q(n5894) );
  AND2X1 U6766 ( .IN1(n3588), .IN2(CRC_OUT_5_28), .Q(n5890) );
  AND2X1 U6767 ( .IN1(n222), .IN2(n3571), .Q(n5889) );
  INVX0 U6768 ( .INP(n5895), .ZN(n222) );
  OR2X1 U6769 ( .IN1(n4430), .IN2(n3938), .Q(n5895) );
  OR4X1 U6770 ( .IN1(n5896), .IN2(n5897), .IN3(n5898), .IN4(n5899), .Q(WX5820)
         );
  AND2X1 U6771 ( .IN1(n3552), .IN2(n5900), .Q(n5899) );
  AND2X1 U6772 ( .IN1(n3645), .IN2(n5437), .Q(n5898) );
  XOR3X1 U6773 ( .IN1(n2949), .IN2(n3514), .IN3(n5901), .Q(n5437) );
  XOR3X1 U6774 ( .IN1(n7147), .IN2(n3283), .IN3(WX7242), .Q(n5901) );
  AND2X1 U6775 ( .IN1(n3589), .IN2(CRC_OUT_5_29), .Q(n5897) );
  AND2X1 U6776 ( .IN1(n221), .IN2(n3571), .Q(n5896) );
  INVX0 U6777 ( .INP(n5902), .ZN(n221) );
  OR2X1 U6778 ( .IN1(n4430), .IN2(n3939), .Q(n5902) );
  OR4X1 U6779 ( .IN1(n5903), .IN2(n5904), .IN3(n5905), .IN4(n5906), .Q(WX5818)
         );
  AND2X1 U6780 ( .IN1(n3552), .IN2(n5907), .Q(n5906) );
  AND2X1 U6781 ( .IN1(n3645), .IN2(n5444), .Q(n5905) );
  XOR3X1 U6782 ( .IN1(n2951), .IN2(n3518), .IN3(n5908), .Q(n5444) );
  XOR3X1 U6783 ( .IN1(n7148), .IN2(n3282), .IN3(WX7240), .Q(n5908) );
  AND2X1 U6784 ( .IN1(n3588), .IN2(CRC_OUT_5_30), .Q(n5904) );
  AND2X1 U6785 ( .IN1(n220), .IN2(n3571), .Q(n5903) );
  INVX0 U6786 ( .INP(n5909), .ZN(n220) );
  OR2X1 U6787 ( .IN1(n4430), .IN2(n3940), .Q(n5909) );
  OR4X1 U6788 ( .IN1(n5910), .IN2(n5911), .IN3(n5912), .IN4(n5913), .Q(WX5816)
         );
  AND2X1 U6789 ( .IN1(n3552), .IN2(n5914), .Q(n5913) );
  AND2X1 U6790 ( .IN1(n3645), .IN2(n5451), .Q(n5912) );
  XOR3X1 U6791 ( .IN1(n2837), .IN2(n3516), .IN3(n5915), .Q(n5451) );
  XOR3X1 U6792 ( .IN1(n7149), .IN2(n3281), .IN3(WX7238), .Q(n5915) );
  AND2X1 U6793 ( .IN1(n2245), .IN2(WX5657), .Q(n5911) );
  AND2X1 U6794 ( .IN1(n3590), .IN2(CRC_OUT_5_31), .Q(n5910) );
  AND2X1 U6795 ( .IN1(n3502), .IN2(n4355), .Q(WX5718) );
  AND2X1 U6796 ( .IN1(n3512), .IN2(n4355), .Q(WX546) );
  AND2X1 U6797 ( .IN1(n5916), .IN2(n4355), .Q(WX5205) );
  XOR2X1 U6798 ( .IN1(CRC_OUT_6_30), .IN2(n3336), .Q(n5916) );
  AND2X1 U6799 ( .IN1(n5917), .IN2(n4356), .Q(WX5203) );
  XOR2X1 U6800 ( .IN1(CRC_OUT_6_29), .IN2(n3337), .Q(n5917) );
  AND2X1 U6801 ( .IN1(n5918), .IN2(n4356), .Q(WX5201) );
  XOR2X1 U6802 ( .IN1(CRC_OUT_6_28), .IN2(n3338), .Q(n5918) );
  AND2X1 U6803 ( .IN1(n5919), .IN2(n4356), .Q(WX5199) );
  XOR2X1 U6804 ( .IN1(test_so40), .IN2(DFF_763_n1), .Q(n5919) );
  AND2X1 U6805 ( .IN1(n5920), .IN2(n4356), .Q(WX5197) );
  XOR2X1 U6806 ( .IN1(CRC_OUT_6_26), .IN2(n3339), .Q(n5920) );
  AND2X1 U6807 ( .IN1(n5921), .IN2(n4356), .Q(WX5195) );
  XOR2X1 U6808 ( .IN1(CRC_OUT_6_25), .IN2(n3340), .Q(n5921) );
  AND2X1 U6809 ( .IN1(n5922), .IN2(n4356), .Q(WX5193) );
  XOR2X1 U6810 ( .IN1(CRC_OUT_6_24), .IN2(n3341), .Q(n5922) );
  AND2X1 U6811 ( .IN1(n5923), .IN2(n4356), .Q(WX5191) );
  XOR2X1 U6812 ( .IN1(CRC_OUT_6_23), .IN2(n3342), .Q(n5923) );
  AND2X1 U6813 ( .IN1(n5924), .IN2(n4356), .Q(WX5189) );
  XOR2X1 U6814 ( .IN1(test_so43), .IN2(n3343), .Q(n5924) );
  AND2X1 U6815 ( .IN1(n5925), .IN2(n4356), .Q(WX5187) );
  XOR2X1 U6816 ( .IN1(CRC_OUT_6_21), .IN2(n3344), .Q(n5925) );
  AND2X1 U6817 ( .IN1(n5926), .IN2(n4357), .Q(WX5185) );
  XOR2X1 U6818 ( .IN1(CRC_OUT_6_20), .IN2(n3345), .Q(n5926) );
  AND2X1 U6819 ( .IN1(n5927), .IN2(n4357), .Q(WX5183) );
  XOR2X1 U6820 ( .IN1(CRC_OUT_6_19), .IN2(n3346), .Q(n5927) );
  AND2X1 U6821 ( .IN1(n5928), .IN2(n4357), .Q(WX5181) );
  XOR2X1 U6822 ( .IN1(CRC_OUT_6_18), .IN2(n3347), .Q(n5928) );
  AND2X1 U6823 ( .IN1(n5929), .IN2(n4357), .Q(WX5179) );
  XOR2X1 U6824 ( .IN1(CRC_OUT_6_17), .IN2(n3348), .Q(n5929) );
  AND2X1 U6825 ( .IN1(n5930), .IN2(n4357), .Q(WX5177) );
  XOR2X1 U6826 ( .IN1(CRC_OUT_6_16), .IN2(n3349), .Q(n5930) );
  AND2X1 U6827 ( .IN1(n5931), .IN2(n4357), .Q(WX5175) );
  XOR3X1 U6828 ( .IN1(n3186), .IN2(DFF_767_n1), .IN3(DFF_751_n1), .Q(n5931) );
  AND2X1 U6829 ( .IN1(n5932), .IN2(n4357), .Q(WX5173) );
  XOR2X1 U6830 ( .IN1(CRC_OUT_6_14), .IN2(n3350), .Q(n5932) );
  AND2X1 U6831 ( .IN1(n5933), .IN2(n4357), .Q(WX5171) );
  XOR2X1 U6832 ( .IN1(CRC_OUT_6_13), .IN2(n3351), .Q(n5933) );
  AND2X1 U6833 ( .IN1(n5934), .IN2(n4357), .Q(WX5169) );
  XOR2X1 U6834 ( .IN1(CRC_OUT_6_12), .IN2(n3352), .Q(n5934) );
  AND2X1 U6835 ( .IN1(n5935), .IN2(n4358), .Q(WX5167) );
  XOR2X1 U6836 ( .IN1(CRC_OUT_6_11), .IN2(n3353), .Q(n5935) );
  AND2X1 U6837 ( .IN1(n5936), .IN2(n4358), .Q(WX5165) );
  XOR3X1 U6838 ( .IN1(test_so41), .IN2(DFF_767_n1), .IN3(CRC_OUT_6_10), .Q(
        n5936) );
  AND2X1 U6839 ( .IN1(n5937), .IN2(n4381), .Q(WX5163) );
  XOR2X1 U6840 ( .IN1(CRC_OUT_6_9), .IN2(n3354), .Q(n5937) );
  AND2X1 U6841 ( .IN1(n5938), .IN2(n4375), .Q(WX5161) );
  XOR2X1 U6842 ( .IN1(CRC_OUT_6_8), .IN2(n3355), .Q(n5938) );
  AND2X1 U6843 ( .IN1(n5939), .IN2(n4375), .Q(WX5159) );
  XOR2X1 U6844 ( .IN1(CRC_OUT_6_7), .IN2(n3356), .Q(n5939) );
  AND2X1 U6845 ( .IN1(n5940), .IN2(n4376), .Q(WX5157) );
  XOR2X1 U6846 ( .IN1(CRC_OUT_6_6), .IN2(n3357), .Q(n5940) );
  AND2X1 U6847 ( .IN1(n5941), .IN2(n4376), .Q(WX5155) );
  XOR2X1 U6848 ( .IN1(test_so42), .IN2(n3358), .Q(n5941) );
  AND2X1 U6849 ( .IN1(n5942), .IN2(n4376), .Q(WX5153) );
  XOR2X1 U6850 ( .IN1(CRC_OUT_6_4), .IN2(n3359), .Q(n5942) );
  AND2X1 U6851 ( .IN1(n5943), .IN2(n4376), .Q(WX5151) );
  XOR3X1 U6852 ( .IN1(n3187), .IN2(DFF_767_n1), .IN3(DFF_739_n1), .Q(n5943) );
  AND2X1 U6853 ( .IN1(n5944), .IN2(n4376), .Q(WX5149) );
  XOR2X1 U6854 ( .IN1(CRC_OUT_6_2), .IN2(n3360), .Q(n5944) );
  AND2X1 U6855 ( .IN1(n5945), .IN2(n4376), .Q(WX5147) );
  XOR2X1 U6856 ( .IN1(CRC_OUT_6_1), .IN2(n3361), .Q(n5945) );
  AND2X1 U6857 ( .IN1(n5946), .IN2(n4376), .Q(WX5145) );
  XOR2X1 U6858 ( .IN1(CRC_OUT_6_0), .IN2(n3362), .Q(n5946) );
  AND2X1 U6859 ( .IN1(n5947), .IN2(n4376), .Q(WX5143) );
  XOR2X1 U6860 ( .IN1(n3199), .IN2(CRC_OUT_6_31), .Q(n5947) );
  INVX0 U6861 ( .INP(n5948), .ZN(WX4617) );
  OR2X1 U6862 ( .IN1(n4430), .IN2(n7191), .Q(n5948) );
  AND2X1 U6863 ( .IN1(test_so35), .IN2(n4376), .Q(WX4615) );
  INVX0 U6864 ( .INP(n5949), .ZN(WX4613) );
  OR2X1 U6865 ( .IN1(n4430), .IN2(n7193), .Q(n5949) );
  INVX0 U6866 ( .INP(n5950), .ZN(WX4611) );
  OR2X1 U6867 ( .IN1(n4430), .IN2(n7194), .Q(n5950) );
  INVX0 U6868 ( .INP(n5951), .ZN(WX4609) );
  OR2X1 U6869 ( .IN1(n4430), .IN2(n7195), .Q(n5951) );
  INVX0 U6870 ( .INP(n5952), .ZN(WX4607) );
  OR2X1 U6871 ( .IN1(n4431), .IN2(n7196), .Q(n5952) );
  INVX0 U6872 ( .INP(n5953), .ZN(WX4605) );
  OR2X1 U6873 ( .IN1(n4431), .IN2(n7197), .Q(n5953) );
  INVX0 U6874 ( .INP(n5954), .ZN(WX4603) );
  OR2X1 U6875 ( .IN1(n4431), .IN2(n7198), .Q(n5954) );
  INVX0 U6876 ( .INP(n5955), .ZN(WX4601) );
  OR2X1 U6877 ( .IN1(n4431), .IN2(n7199), .Q(n5955) );
  INVX0 U6878 ( .INP(n5956), .ZN(WX4599) );
  OR2X1 U6879 ( .IN1(n4431), .IN2(n7200), .Q(n5956) );
  INVX0 U6880 ( .INP(n5957), .ZN(WX4597) );
  OR2X1 U6881 ( .IN1(n4431), .IN2(n7201), .Q(n5957) );
  INVX0 U6882 ( .INP(n5958), .ZN(WX4595) );
  OR2X1 U6883 ( .IN1(n4431), .IN2(n7202), .Q(n5958) );
  INVX0 U6884 ( .INP(n5959), .ZN(WX4593) );
  OR2X1 U6885 ( .IN1(n4431), .IN2(n7203), .Q(n5959) );
  INVX0 U6886 ( .INP(n5960), .ZN(WX4591) );
  OR2X1 U6887 ( .IN1(n4431), .IN2(n7204), .Q(n5960) );
  INVX0 U6888 ( .INP(n5961), .ZN(WX4589) );
  OR2X1 U6889 ( .IN1(n4431), .IN2(n7205), .Q(n5961) );
  INVX0 U6890 ( .INP(n5962), .ZN(WX4587) );
  OR2X1 U6891 ( .IN1(n4431), .IN2(n7206), .Q(n5962) );
  OR4X1 U6892 ( .IN1(n5963), .IN2(n5964), .IN3(n5965), .IN4(n5966), .Q(WX4585)
         );
  AND2X1 U6893 ( .IN1(n5967), .IN2(n3532), .Q(n5966) );
  AND2X1 U6894 ( .IN1(n3645), .IN2(n5697), .Q(n5965) );
  XNOR3X1 U6895 ( .IN1(n3198), .IN2(n3116), .IN3(n5968), .Q(n5697) );
  XOR2X1 U6896 ( .IN1(WX5943), .IN2(n7150), .Q(n5968) );
  AND2X1 U6897 ( .IN1(n3588), .IN2(CRC_OUT_6_0), .Q(n5964) );
  AND2X1 U6898 ( .IN1(n188), .IN2(n3571), .Q(n5963) );
  INVX0 U6899 ( .INP(n5969), .ZN(n188) );
  OR2X1 U6900 ( .IN1(n4431), .IN2(n3941), .Q(n5969) );
  OR4X1 U6901 ( .IN1(n5970), .IN2(n5971), .IN3(n5972), .IN4(n5973), .Q(WX4583)
         );
  AND2X1 U6902 ( .IN1(n3552), .IN2(n5974), .Q(n5973) );
  AND2X1 U6903 ( .IN1(n5704), .IN2(n3620), .Q(n5972) );
  XOR3X1 U6904 ( .IN1(n3661), .IN2(n3335), .IN3(n5975), .Q(n5704) );
  XOR2X1 U6905 ( .IN1(WX5877), .IN2(test_so51), .Q(n5975) );
  AND2X1 U6906 ( .IN1(n3589), .IN2(CRC_OUT_6_1), .Q(n5971) );
  AND2X1 U6907 ( .IN1(n187), .IN2(n3571), .Q(n5970) );
  INVX0 U6908 ( .INP(n5976), .ZN(n187) );
  OR2X1 U6909 ( .IN1(n4431), .IN2(n3942), .Q(n5976) );
  OR4X1 U6910 ( .IN1(n5977), .IN2(n5978), .IN3(n5979), .IN4(n5980), .Q(WX4581)
         );
  AND2X1 U6911 ( .IN1(n3552), .IN2(n5981), .Q(n5980) );
  AND2X1 U6912 ( .IN1(n3645), .IN2(n5711), .Q(n5979) );
  XNOR3X1 U6913 ( .IN1(n3334), .IN2(n3117), .IN3(n5982), .Q(n5711) );
  XOR2X1 U6914 ( .IN1(WX5939), .IN2(n7151), .Q(n5982) );
  AND2X1 U6915 ( .IN1(n3588), .IN2(CRC_OUT_6_2), .Q(n5978) );
  AND2X1 U6916 ( .IN1(n186), .IN2(n3571), .Q(n5977) );
  INVX0 U6917 ( .INP(n5983), .ZN(n186) );
  OR2X1 U6918 ( .IN1(n4432), .IN2(n3943), .Q(n5983) );
  OR4X1 U6919 ( .IN1(n5984), .IN2(n5985), .IN3(n5986), .IN4(n5987), .Q(WX4579)
         );
  AND2X1 U6920 ( .IN1(n3552), .IN2(n5988), .Q(n5987) );
  AND2X1 U6921 ( .IN1(n5718), .IN2(n3620), .Q(n5986) );
  XOR3X1 U6922 ( .IN1(n3333), .IN2(n3118), .IN3(n5989), .Q(n5718) );
  XOR2X1 U6923 ( .IN1(WX5873), .IN2(test_so49), .Q(n5989) );
  AND2X1 U6924 ( .IN1(n3589), .IN2(CRC_OUT_6_3), .Q(n5985) );
  AND2X1 U6925 ( .IN1(n185), .IN2(n3571), .Q(n5984) );
  INVX0 U6926 ( .INP(n5990), .ZN(n185) );
  OR2X1 U6927 ( .IN1(n4432), .IN2(n3944), .Q(n5990) );
  OR4X1 U6928 ( .IN1(n5991), .IN2(n5992), .IN3(n5993), .IN4(n5994), .Q(WX4577)
         );
  AND2X1 U6929 ( .IN1(n3552), .IN2(n5995), .Q(n5994) );
  AND2X1 U6930 ( .IN1(n3628), .IN2(n5725), .Q(n5993) );
  XNOR3X1 U6931 ( .IN1(n3185), .IN2(n3119), .IN3(n5996), .Q(n5725) );
  XOR2X1 U6932 ( .IN1(WX5935), .IN2(n7152), .Q(n5996) );
  AND2X1 U6933 ( .IN1(n3589), .IN2(CRC_OUT_6_4), .Q(n5992) );
  AND2X1 U6934 ( .IN1(n184), .IN2(n3570), .Q(n5991) );
  INVX0 U6935 ( .INP(n5997), .ZN(n184) );
  OR2X1 U6936 ( .IN1(n4432), .IN2(n3945), .Q(n5997) );
  OR4X1 U6937 ( .IN1(n5998), .IN2(n5999), .IN3(n6000), .IN4(n6001), .Q(WX4575)
         );
  AND2X1 U6938 ( .IN1(n3552), .IN2(n6002), .Q(n6001) );
  AND2X1 U6939 ( .IN1(n5732), .IN2(n3620), .Q(n6000) );
  XOR3X1 U6940 ( .IN1(n3669), .IN2(n3332), .IN3(n6003), .Q(n5732) );
  XOR2X1 U6941 ( .IN1(WX5997), .IN2(test_so47), .Q(n6003) );
  AND2X1 U6942 ( .IN1(test_so42), .IN2(n3587), .Q(n5999) );
  AND2X1 U6943 ( .IN1(n183), .IN2(n3570), .Q(n5998) );
  INVX0 U6944 ( .INP(n6004), .ZN(n183) );
  OR2X1 U6945 ( .IN1(n4432), .IN2(n3946), .Q(n6004) );
  OR4X1 U6946 ( .IN1(n6005), .IN2(n6006), .IN3(n6007), .IN4(n6008), .Q(WX4573)
         );
  AND2X1 U6947 ( .IN1(n3552), .IN2(n6009), .Q(n6008) );
  AND2X1 U6948 ( .IN1(n3630), .IN2(n5739), .Q(n6007) );
  XNOR3X1 U6949 ( .IN1(n3331), .IN2(n3120), .IN3(n6010), .Q(n5739) );
  XOR2X1 U6950 ( .IN1(WX5931), .IN2(n7153), .Q(n6010) );
  AND2X1 U6951 ( .IN1(n3589), .IN2(CRC_OUT_6_6), .Q(n6006) );
  AND2X1 U6952 ( .IN1(n182), .IN2(n3570), .Q(n6005) );
  INVX0 U6953 ( .INP(n6011), .ZN(n182) );
  OR2X1 U6954 ( .IN1(n4432), .IN2(n3947), .Q(n6011) );
  OR4X1 U6955 ( .IN1(n6012), .IN2(n6013), .IN3(n6014), .IN4(n6015), .Q(WX4571)
         );
  AND2X1 U6956 ( .IN1(n3551), .IN2(n6016), .Q(n6015) );
  AND2X1 U6957 ( .IN1(n3628), .IN2(n5746), .Q(n6014) );
  XNOR3X1 U6958 ( .IN1(n3330), .IN2(n3121), .IN3(n6017), .Q(n5746) );
  XOR2X1 U6959 ( .IN1(WX5929), .IN2(n7154), .Q(n6017) );
  AND2X1 U6960 ( .IN1(n3589), .IN2(CRC_OUT_6_7), .Q(n6013) );
  AND2X1 U6961 ( .IN1(n181), .IN2(n3570), .Q(n6012) );
  INVX0 U6962 ( .INP(n6018), .ZN(n181) );
  OR2X1 U6963 ( .IN1(n4432), .IN2(n3948), .Q(n6018) );
  OR4X1 U6964 ( .IN1(n6019), .IN2(n6020), .IN3(n6021), .IN4(n6022), .Q(WX4569)
         );
  AND2X1 U6965 ( .IN1(n3551), .IN2(n6023), .Q(n6022) );
  AND2X1 U6966 ( .IN1(n3628), .IN2(n5753), .Q(n6021) );
  XNOR3X1 U6967 ( .IN1(n3329), .IN2(n3122), .IN3(n6024), .Q(n5753) );
  XOR2X1 U6968 ( .IN1(WX5927), .IN2(n7155), .Q(n6024) );
  AND2X1 U6969 ( .IN1(n3592), .IN2(CRC_OUT_6_8), .Q(n6020) );
  AND2X1 U6970 ( .IN1(n180), .IN2(n3570), .Q(n6019) );
  INVX0 U6971 ( .INP(n6025), .ZN(n180) );
  OR2X1 U6972 ( .IN1(n4432), .IN2(n3949), .Q(n6025) );
  OR4X1 U6973 ( .IN1(n6026), .IN2(n6027), .IN3(n6028), .IN4(n6029), .Q(WX4567)
         );
  AND2X1 U6974 ( .IN1(n3551), .IN2(n6030), .Q(n6029) );
  AND2X1 U6975 ( .IN1(n3629), .IN2(n5760), .Q(n6028) );
  XNOR3X1 U6976 ( .IN1(n3328), .IN2(n3123), .IN3(n6031), .Q(n5760) );
  XOR2X1 U6977 ( .IN1(WX5925), .IN2(n7156), .Q(n6031) );
  AND2X1 U6978 ( .IN1(n3589), .IN2(CRC_OUT_6_9), .Q(n6027) );
  AND2X1 U6979 ( .IN1(n179), .IN2(n3570), .Q(n6026) );
  INVX0 U6980 ( .INP(n6032), .ZN(n179) );
  OR2X1 U6981 ( .IN1(n4432), .IN2(n3950), .Q(n6032) );
  OR4X1 U6982 ( .IN1(n6033), .IN2(n6034), .IN3(n6035), .IN4(n6036), .Q(WX4565)
         );
  AND2X1 U6983 ( .IN1(n3551), .IN2(n6037), .Q(n6036) );
  AND2X1 U6984 ( .IN1(n3629), .IN2(n5767), .Q(n6035) );
  XNOR3X1 U6985 ( .IN1(n3327), .IN2(n3124), .IN3(n6038), .Q(n5767) );
  XOR2X1 U6986 ( .IN1(WX5923), .IN2(n7157), .Q(n6038) );
  AND2X1 U6987 ( .IN1(n3590), .IN2(CRC_OUT_6_10), .Q(n6034) );
  AND2X1 U6988 ( .IN1(n178), .IN2(n3570), .Q(n6033) );
  INVX0 U6989 ( .INP(n6039), .ZN(n178) );
  OR2X1 U6990 ( .IN1(n4432), .IN2(n3951), .Q(n6039) );
  OR4X1 U6991 ( .IN1(n6040), .IN2(n6041), .IN3(n6042), .IN4(n6043), .Q(WX4563)
         );
  AND2X1 U6992 ( .IN1(n6044), .IN2(n3534), .Q(n6043) );
  AND2X1 U6993 ( .IN1(n3628), .IN2(n5774), .Q(n6042) );
  XNOR3X1 U6994 ( .IN1(n3184), .IN2(n3125), .IN3(n6045), .Q(n5774) );
  XOR2X1 U6995 ( .IN1(WX5921), .IN2(n7158), .Q(n6045) );
  AND2X1 U6996 ( .IN1(n3589), .IN2(CRC_OUT_6_11), .Q(n6041) );
  AND2X1 U6997 ( .IN1(n177), .IN2(n3570), .Q(n6040) );
  INVX0 U6998 ( .INP(n6046), .ZN(n177) );
  OR2X1 U6999 ( .IN1(n4432), .IN2(n3952), .Q(n6046) );
  OR4X1 U7000 ( .IN1(n6047), .IN2(n6048), .IN3(n6049), .IN4(n6050), .Q(WX4561)
         );
  AND2X1 U7001 ( .IN1(n3551), .IN2(n6051), .Q(n6050) );
  AND2X1 U7002 ( .IN1(n3629), .IN2(n5781), .Q(n6049) );
  XNOR3X1 U7003 ( .IN1(n3326), .IN2(n3126), .IN3(n6052), .Q(n5781) );
  XOR2X1 U7004 ( .IN1(WX5919), .IN2(n7159), .Q(n6052) );
  AND2X1 U7005 ( .IN1(n3590), .IN2(CRC_OUT_6_12), .Q(n6048) );
  AND2X1 U7006 ( .IN1(n176), .IN2(n3570), .Q(n6047) );
  INVX0 U7007 ( .INP(n6053), .ZN(n176) );
  OR2X1 U7008 ( .IN1(n4432), .IN2(n3953), .Q(n6053) );
  OR4X1 U7009 ( .IN1(n6054), .IN2(n6055), .IN3(n6056), .IN4(n6057), .Q(WX4559)
         );
  AND2X1 U7010 ( .IN1(n6058), .IN2(n3534), .Q(n6057) );
  AND2X1 U7011 ( .IN1(n3629), .IN2(n5788), .Q(n6056) );
  XNOR3X1 U7012 ( .IN1(n3325), .IN2(n3127), .IN3(n6059), .Q(n5788) );
  XOR2X1 U7013 ( .IN1(WX5917), .IN2(n7160), .Q(n6059) );
  AND2X1 U7014 ( .IN1(n3589), .IN2(CRC_OUT_6_13), .Q(n6055) );
  AND2X1 U7015 ( .IN1(n175), .IN2(n3570), .Q(n6054) );
  INVX0 U7016 ( .INP(n6060), .ZN(n175) );
  OR2X1 U7017 ( .IN1(n4432), .IN2(n3954), .Q(n6060) );
  OR4X1 U7018 ( .IN1(n6061), .IN2(n6062), .IN3(n6063), .IN4(n6064), .Q(WX4557)
         );
  AND2X1 U7019 ( .IN1(n3551), .IN2(n6065), .Q(n6064) );
  AND2X1 U7020 ( .IN1(n3628), .IN2(n5795), .Q(n6063) );
  XNOR3X1 U7021 ( .IN1(n3324), .IN2(n3128), .IN3(n6066), .Q(n5795) );
  XOR2X1 U7022 ( .IN1(WX5915), .IN2(n7161), .Q(n6066) );
  AND2X1 U7023 ( .IN1(n3592), .IN2(CRC_OUT_6_14), .Q(n6062) );
  AND2X1 U7024 ( .IN1(n174), .IN2(n3570), .Q(n6061) );
  INVX0 U7025 ( .INP(n6067), .ZN(n174) );
  OR2X1 U7026 ( .IN1(n4433), .IN2(n3955), .Q(n6067) );
  OR4X1 U7027 ( .IN1(n6068), .IN2(n6069), .IN3(n6070), .IN4(n6071), .Q(WX4555)
         );
  AND2X1 U7028 ( .IN1(n6072), .IN2(n3532), .Q(n6071) );
  AND2X1 U7029 ( .IN1(n3629), .IN2(n5802), .Q(n6070) );
  XNOR3X1 U7030 ( .IN1(n3323), .IN2(n3129), .IN3(n6073), .Q(n5802) );
  XOR2X1 U7031 ( .IN1(WX5913), .IN2(n7162), .Q(n6073) );
  AND2X1 U7032 ( .IN1(n3589), .IN2(CRC_OUT_6_15), .Q(n6069) );
  AND2X1 U7033 ( .IN1(n173), .IN2(n3570), .Q(n6068) );
  INVX0 U7034 ( .INP(n6074), .ZN(n173) );
  OR2X1 U7035 ( .IN1(n4433), .IN2(n3956), .Q(n6074) );
  OR4X1 U7036 ( .IN1(n6075), .IN2(n6076), .IN3(n6077), .IN4(n6078), .Q(WX4553)
         );
  AND2X1 U7037 ( .IN1(n3551), .IN2(n6079), .Q(n6078) );
  AND2X1 U7038 ( .IN1(n5809), .IN2(n3620), .Q(n6077) );
  XOR3X1 U7039 ( .IN1(n2953), .IN2(TM1), .IN3(n6080), .Q(n5809) );
  XOR3X1 U7040 ( .IN1(test_so52), .IN2(n7163), .IN3(WX5975), .Q(n6080) );
  AND2X1 U7041 ( .IN1(n3590), .IN2(CRC_OUT_6_16), .Q(n6076) );
  AND2X1 U7042 ( .IN1(n172), .IN2(n3568), .Q(n6075) );
  INVX0 U7043 ( .INP(n6081), .ZN(n172) );
  OR2X1 U7044 ( .IN1(n4433), .IN2(n3957), .Q(n6081) );
  OR4X1 U7045 ( .IN1(n6082), .IN2(n6083), .IN3(n6084), .IN4(n6085), .Q(WX4551)
         );
  AND2X1 U7046 ( .IN1(n6086), .IN2(n3532), .Q(n6085) );
  AND2X1 U7047 ( .IN1(n3628), .IN2(n5816), .Q(n6084) );
  XOR3X1 U7048 ( .IN1(n2954), .IN2(n3515), .IN3(n6087), .Q(n5816) );
  XOR3X1 U7049 ( .IN1(n7164), .IN2(n3322), .IN3(WX5973), .Q(n6087) );
  AND2X1 U7050 ( .IN1(n3590), .IN2(CRC_OUT_6_17), .Q(n6083) );
  AND2X1 U7051 ( .IN1(n171), .IN2(n3568), .Q(n6082) );
  INVX0 U7052 ( .INP(n6088), .ZN(n171) );
  OR2X1 U7053 ( .IN1(n4433), .IN2(n3958), .Q(n6088) );
  OR4X1 U7054 ( .IN1(n6089), .IN2(n6090), .IN3(n6091), .IN4(n6092), .Q(WX4549)
         );
  AND2X1 U7055 ( .IN1(n3551), .IN2(n6093), .Q(n6092) );
  AND2X1 U7056 ( .IN1(n5823), .IN2(n3623), .Q(n6091) );
  XOR3X1 U7057 ( .IN1(n2956), .IN2(TM1), .IN3(n6094), .Q(n5823) );
  XNOR3X1 U7058 ( .IN1(test_so50), .IN2(n7165), .IN3(n3321), .Q(n6094) );
  AND2X1 U7059 ( .IN1(n3590), .IN2(CRC_OUT_6_18), .Q(n6090) );
  AND2X1 U7060 ( .IN1(n170), .IN2(n3568), .Q(n6089) );
  INVX0 U7061 ( .INP(n6095), .ZN(n170) );
  OR2X1 U7062 ( .IN1(n4433), .IN2(n3959), .Q(n6095) );
  OR4X1 U7063 ( .IN1(n6096), .IN2(n6097), .IN3(n6098), .IN4(n6099), .Q(WX4547)
         );
  AND2X1 U7064 ( .IN1(n3551), .IN2(n6100), .Q(n6099) );
  AND2X1 U7065 ( .IN1(n3628), .IN2(n5830), .Q(n6098) );
  XOR3X1 U7066 ( .IN1(n2957), .IN2(n3514), .IN3(n6101), .Q(n5830) );
  XOR3X1 U7067 ( .IN1(n7166), .IN2(n3320), .IN3(WX5969), .Q(n6101) );
  AND2X1 U7068 ( .IN1(n3590), .IN2(CRC_OUT_6_19), .Q(n6097) );
  AND2X1 U7069 ( .IN1(n169), .IN2(n3568), .Q(n6096) );
  INVX0 U7070 ( .INP(n6102), .ZN(n169) );
  OR2X1 U7071 ( .IN1(n4433), .IN2(n3960), .Q(n6102) );
  OR4X1 U7072 ( .IN1(n6103), .IN2(n6104), .IN3(n6105), .IN4(n6106), .Q(WX4545)
         );
  AND2X1 U7073 ( .IN1(n3551), .IN2(n6107), .Q(n6106) );
  AND2X1 U7074 ( .IN1(n5837), .IN2(n3620), .Q(n6105) );
  XOR3X1 U7075 ( .IN1(n2959), .IN2(TM1), .IN3(n6108), .Q(n5837) );
  XNOR3X1 U7076 ( .IN1(test_so48), .IN2(n7167), .IN3(n3319), .Q(n6108) );
  AND2X1 U7077 ( .IN1(n3590), .IN2(CRC_OUT_6_20), .Q(n6104) );
  AND2X1 U7078 ( .IN1(n168), .IN2(n3568), .Q(n6103) );
  INVX0 U7079 ( .INP(n6109), .ZN(n168) );
  OR2X1 U7080 ( .IN1(n4433), .IN2(n3961), .Q(n6109) );
  OR4X1 U7081 ( .IN1(n6110), .IN2(n6111), .IN3(n6112), .IN4(n6113), .Q(WX4543)
         );
  AND2X1 U7082 ( .IN1(n3551), .IN2(n6114), .Q(n6113) );
  AND2X1 U7083 ( .IN1(n3629), .IN2(n5844), .Q(n6112) );
  XOR3X1 U7084 ( .IN1(n2960), .IN2(n3518), .IN3(n6115), .Q(n5844) );
  XOR3X1 U7085 ( .IN1(n7168), .IN2(n3318), .IN3(WX5965), .Q(n6115) );
  AND2X1 U7086 ( .IN1(n3590), .IN2(CRC_OUT_6_21), .Q(n6111) );
  AND2X1 U7087 ( .IN1(n167), .IN2(n3568), .Q(n6110) );
  INVX0 U7088 ( .INP(n6116), .ZN(n167) );
  OR2X1 U7089 ( .IN1(n4433), .IN2(n3962), .Q(n6116) );
  OR4X1 U7090 ( .IN1(n6117), .IN2(n6118), .IN3(n6119), .IN4(n6120), .Q(WX4541)
         );
  AND2X1 U7091 ( .IN1(n3551), .IN2(n6121), .Q(n6120) );
  AND2X1 U7092 ( .IN1(n5851), .IN2(n3620), .Q(n6119) );
  XOR3X1 U7093 ( .IN1(n2962), .IN2(TM1), .IN3(n6122), .Q(n5851) );
  XNOR3X1 U7094 ( .IN1(test_so46), .IN2(n7169), .IN3(n3317), .Q(n6122) );
  AND2X1 U7095 ( .IN1(test_so43), .IN2(n3587), .Q(n6118) );
  AND2X1 U7096 ( .IN1(n166), .IN2(n3568), .Q(n6117) );
  INVX0 U7097 ( .INP(n6123), .ZN(n166) );
  OR2X1 U7098 ( .IN1(n4433), .IN2(n3963), .Q(n6123) );
  OR4X1 U7099 ( .IN1(n6124), .IN2(n6125), .IN3(n6126), .IN4(n6127), .Q(WX4539)
         );
  AND2X1 U7100 ( .IN1(n3551), .IN2(n6128), .Q(n6127) );
  AND2X1 U7101 ( .IN1(n3629), .IN2(n5858), .Q(n6126) );
  XOR3X1 U7102 ( .IN1(n2963), .IN2(n3516), .IN3(n6129), .Q(n5858) );
  XOR3X1 U7103 ( .IN1(n7170), .IN2(n3316), .IN3(WX5961), .Q(n6129) );
  AND2X1 U7104 ( .IN1(n3592), .IN2(CRC_OUT_6_23), .Q(n6125) );
  AND2X1 U7105 ( .IN1(n165), .IN2(n3568), .Q(n6124) );
  INVX0 U7106 ( .INP(n6130), .ZN(n165) );
  OR2X1 U7107 ( .IN1(n4433), .IN2(n3964), .Q(n6130) );
  OR4X1 U7108 ( .IN1(n6131), .IN2(n6132), .IN3(n6133), .IN4(n6134), .Q(WX4537)
         );
  AND2X1 U7109 ( .IN1(n3550), .IN2(n6135), .Q(n6134) );
  AND2X1 U7110 ( .IN1(n3629), .IN2(n5865), .Q(n6133) );
  XOR3X1 U7111 ( .IN1(n2965), .IN2(n3515), .IN3(n6136), .Q(n5865) );
  XOR3X1 U7112 ( .IN1(n7171), .IN2(n3315), .IN3(WX5959), .Q(n6136) );
  AND2X1 U7113 ( .IN1(n3590), .IN2(CRC_OUT_6_24), .Q(n6132) );
  AND2X1 U7114 ( .IN1(n164), .IN2(n3568), .Q(n6131) );
  INVX0 U7115 ( .INP(n6137), .ZN(n164) );
  OR2X1 U7116 ( .IN1(n4433), .IN2(n3965), .Q(n6137) );
  OR4X1 U7117 ( .IN1(n6138), .IN2(n6139), .IN3(n6140), .IN4(n6141), .Q(WX4535)
         );
  AND2X1 U7118 ( .IN1(n3550), .IN2(n6142), .Q(n6141) );
  AND2X1 U7119 ( .IN1(n3629), .IN2(n5872), .Q(n6140) );
  XOR3X1 U7120 ( .IN1(n2967), .IN2(n3514), .IN3(n6143), .Q(n5872) );
  XOR3X1 U7121 ( .IN1(n7172), .IN2(n3314), .IN3(WX5957), .Q(n6143) );
  AND2X1 U7122 ( .IN1(n3592), .IN2(CRC_OUT_6_25), .Q(n6139) );
  AND2X1 U7123 ( .IN1(n163), .IN2(n3568), .Q(n6138) );
  INVX0 U7124 ( .INP(n6144), .ZN(n163) );
  OR2X1 U7125 ( .IN1(n4433), .IN2(n3966), .Q(n6144) );
  OR4X1 U7126 ( .IN1(n6145), .IN2(n6146), .IN3(n6147), .IN4(n6148), .Q(WX4533)
         );
  AND2X1 U7127 ( .IN1(n3550), .IN2(n6149), .Q(n6148) );
  AND2X1 U7128 ( .IN1(n3629), .IN2(n5879), .Q(n6147) );
  XOR3X1 U7129 ( .IN1(n2969), .IN2(n3518), .IN3(n6150), .Q(n5879) );
  XOR3X1 U7130 ( .IN1(n7173), .IN2(n3313), .IN3(WX5955), .Q(n6150) );
  AND2X1 U7131 ( .IN1(n3590), .IN2(CRC_OUT_6_26), .Q(n6146) );
  AND2X1 U7132 ( .IN1(n162), .IN2(n3568), .Q(n6145) );
  INVX0 U7133 ( .INP(n6151), .ZN(n162) );
  OR2X1 U7134 ( .IN1(n4433), .IN2(n3967), .Q(n6151) );
  OR4X1 U7135 ( .IN1(n6152), .IN2(n6153), .IN3(n6154), .IN4(n6155), .Q(WX4531)
         );
  AND2X1 U7136 ( .IN1(n3550), .IN2(n6156), .Q(n6155) );
  AND2X1 U7137 ( .IN1(n3629), .IN2(n5886), .Q(n6154) );
  XOR3X1 U7138 ( .IN1(n2971), .IN2(n3516), .IN3(n6157), .Q(n5886) );
  XOR3X1 U7139 ( .IN1(n7174), .IN2(n3312), .IN3(WX5953), .Q(n6157) );
  AND2X1 U7140 ( .IN1(n3592), .IN2(CRC_OUT_6_27), .Q(n6153) );
  AND2X1 U7141 ( .IN1(n161), .IN2(n3568), .Q(n6152) );
  INVX0 U7142 ( .INP(n6158), .ZN(n161) );
  OR2X1 U7143 ( .IN1(n4434), .IN2(n3968), .Q(n6158) );
  OR4X1 U7144 ( .IN1(n6159), .IN2(n6160), .IN3(n6161), .IN4(n6162), .Q(WX4529)
         );
  AND2X1 U7145 ( .IN1(n6163), .IN2(n3528), .Q(n6162) );
  AND2X1 U7146 ( .IN1(n3630), .IN2(n5893), .Q(n6161) );
  XOR3X1 U7147 ( .IN1(n2973), .IN2(n3515), .IN3(n6164), .Q(n5893) );
  XOR3X1 U7148 ( .IN1(n7175), .IN2(n3311), .IN3(WX5951), .Q(n6164) );
  AND2X1 U7149 ( .IN1(n3590), .IN2(CRC_OUT_6_28), .Q(n6160) );
  AND2X1 U7150 ( .IN1(n160), .IN2(n3567), .Q(n6159) );
  INVX0 U7151 ( .INP(n6165), .ZN(n160) );
  OR2X1 U7152 ( .IN1(n4434), .IN2(n3969), .Q(n6165) );
  OR4X1 U7153 ( .IN1(n6166), .IN2(n6167), .IN3(n6168), .IN4(n6169), .Q(WX4527)
         );
  AND2X1 U7154 ( .IN1(n3550), .IN2(n6170), .Q(n6169) );
  AND2X1 U7155 ( .IN1(n3629), .IN2(n5900), .Q(n6168) );
  XOR3X1 U7156 ( .IN1(n2975), .IN2(n3514), .IN3(n6171), .Q(n5900) );
  XOR3X1 U7157 ( .IN1(n7176), .IN2(n3310), .IN3(WX5949), .Q(n6171) );
  AND2X1 U7158 ( .IN1(n3593), .IN2(CRC_OUT_6_29), .Q(n6167) );
  AND2X1 U7159 ( .IN1(n159), .IN2(n3567), .Q(n6166) );
  INVX0 U7160 ( .INP(n6172), .ZN(n159) );
  OR2X1 U7161 ( .IN1(n4434), .IN2(n3970), .Q(n6172) );
  OR4X1 U7162 ( .IN1(n6173), .IN2(n6174), .IN3(n6175), .IN4(n6176), .Q(WX4525)
         );
  AND2X1 U7163 ( .IN1(n6177), .IN2(n3528), .Q(n6176) );
  AND2X1 U7164 ( .IN1(n3630), .IN2(n5907), .Q(n6175) );
  XOR3X1 U7165 ( .IN1(n2977), .IN2(n3518), .IN3(n6178), .Q(n5907) );
  XOR3X1 U7166 ( .IN1(n7177), .IN2(n3309), .IN3(WX5947), .Q(n6178) );
  AND2X1 U7167 ( .IN1(n3592), .IN2(CRC_OUT_6_30), .Q(n6174) );
  AND2X1 U7168 ( .IN1(n158), .IN2(n3567), .Q(n6173) );
  INVX0 U7169 ( .INP(n6179), .ZN(n158) );
  OR2X1 U7170 ( .IN1(n4434), .IN2(n3971), .Q(n6179) );
  OR4X1 U7171 ( .IN1(n6180), .IN2(n6181), .IN3(n6182), .IN4(n6183), .Q(WX4523)
         );
  AND2X1 U7172 ( .IN1(n3550), .IN2(n6184), .Q(n6183) );
  AND2X1 U7173 ( .IN1(n3630), .IN2(n5914), .Q(n6182) );
  XOR3X1 U7174 ( .IN1(n2839), .IN2(n3516), .IN3(n6185), .Q(n5914) );
  XOR3X1 U7175 ( .IN1(n7178), .IN2(n3308), .IN3(WX5945), .Q(n6185) );
  AND2X1 U7176 ( .IN1(n2245), .IN2(WX4364), .Q(n6181) );
  AND2X1 U7177 ( .IN1(n3592), .IN2(CRC_OUT_6_31), .Q(n6180) );
  AND2X1 U7178 ( .IN1(n3500), .IN2(n4377), .Q(WX4425) );
  AND2X1 U7179 ( .IN1(n6186), .IN2(n4377), .Q(WX3912) );
  XOR2X1 U7180 ( .IN1(CRC_OUT_7_30), .IN2(n3363), .Q(n6186) );
  AND2X1 U7181 ( .IN1(n6187), .IN2(n4377), .Q(WX3910) );
  XOR2X1 U7182 ( .IN1(CRC_OUT_7_29), .IN2(n3364), .Q(n6187) );
  AND2X1 U7183 ( .IN1(n6188), .IN2(n4377), .Q(WX3908) );
  XOR2X1 U7184 ( .IN1(CRC_OUT_7_28), .IN2(n3365), .Q(n6188) );
  AND2X1 U7185 ( .IN1(n6189), .IN2(n4377), .Q(WX3906) );
  XOR2X1 U7186 ( .IN1(test_so32), .IN2(n3366), .Q(n6189) );
  AND2X1 U7187 ( .IN1(n6190), .IN2(n4377), .Q(WX3904) );
  XOR2X1 U7188 ( .IN1(CRC_OUT_7_26), .IN2(n3367), .Q(n6190) );
  AND2X1 U7189 ( .IN1(n6191), .IN2(n4377), .Q(WX3902) );
  XOR2X1 U7190 ( .IN1(CRC_OUT_7_25), .IN2(n3368), .Q(n6191) );
  AND2X1 U7191 ( .IN1(n6192), .IN2(n4377), .Q(WX3900) );
  XOR2X1 U7192 ( .IN1(CRC_OUT_7_24), .IN2(n3369), .Q(n6192) );
  AND2X1 U7193 ( .IN1(n6193), .IN2(n4377), .Q(WX3898) );
  XOR2X1 U7194 ( .IN1(CRC_OUT_7_23), .IN2(n3370), .Q(n6193) );
  AND2X1 U7195 ( .IN1(n6194), .IN2(n4378), .Q(WX3896) );
  XOR2X1 U7196 ( .IN1(test_so29), .IN2(DFF_566_n1), .Q(n6194) );
  AND2X1 U7197 ( .IN1(n6195), .IN2(n4378), .Q(WX3894) );
  XOR2X1 U7198 ( .IN1(CRC_OUT_7_21), .IN2(n3371), .Q(n6195) );
  AND2X1 U7199 ( .IN1(n6196), .IN2(n4378), .Q(WX3892) );
  XOR2X1 U7200 ( .IN1(CRC_OUT_7_20), .IN2(n3372), .Q(n6196) );
  AND2X1 U7201 ( .IN1(n6197), .IN2(n4378), .Q(WX3890) );
  XOR2X1 U7202 ( .IN1(CRC_OUT_7_19), .IN2(n3373), .Q(n6197) );
  AND2X1 U7203 ( .IN1(n6198), .IN2(n4378), .Q(WX3888) );
  XOR2X1 U7204 ( .IN1(CRC_OUT_7_18), .IN2(n3374), .Q(n6198) );
  AND2X1 U7205 ( .IN1(n6199), .IN2(n4378), .Q(WX3886) );
  XOR2X1 U7206 ( .IN1(CRC_OUT_7_17), .IN2(n3375), .Q(n6199) );
  AND2X1 U7207 ( .IN1(n6200), .IN2(n4378), .Q(WX3884) );
  XOR2X1 U7208 ( .IN1(CRC_OUT_7_16), .IN2(n3376), .Q(n6200) );
  AND2X1 U7209 ( .IN1(n6201), .IN2(n4378), .Q(WX3882) );
  XOR3X1 U7210 ( .IN1(n3188), .IN2(DFF_575_n1), .IN3(DFF_559_n1), .Q(n6201) );
  AND2X1 U7211 ( .IN1(n6202), .IN2(n4378), .Q(WX3880) );
  XOR2X1 U7212 ( .IN1(CRC_OUT_7_14), .IN2(n3377), .Q(n6202) );
  AND2X1 U7213 ( .IN1(n6203), .IN2(n4379), .Q(WX3878) );
  XOR2X1 U7214 ( .IN1(CRC_OUT_7_13), .IN2(n3378), .Q(n6203) );
  AND2X1 U7215 ( .IN1(n6204), .IN2(n4379), .Q(WX3876) );
  XOR2X1 U7216 ( .IN1(CRC_OUT_7_12), .IN2(n3379), .Q(n6204) );
  AND2X1 U7217 ( .IN1(n6205), .IN2(n4379), .Q(WX3874) );
  XOR2X1 U7218 ( .IN1(CRC_OUT_7_11), .IN2(n3380), .Q(n6205) );
  AND2X1 U7219 ( .IN1(n6206), .IN2(n4379), .Q(WX3872) );
  XOR3X1 U7220 ( .IN1(test_so31), .IN2(n3189), .IN3(CRC_OUT_7_31), .Q(n6206)
         );
  AND2X1 U7221 ( .IN1(n6207), .IN2(n4379), .Q(WX3870) );
  XOR2X1 U7222 ( .IN1(CRC_OUT_7_9), .IN2(n3381), .Q(n6207) );
  AND2X1 U7223 ( .IN1(n6208), .IN2(n4379), .Q(WX3868) );
  XOR2X1 U7224 ( .IN1(CRC_OUT_7_8), .IN2(n3382), .Q(n6208) );
  AND2X1 U7225 ( .IN1(n6209), .IN2(n4379), .Q(WX3866) );
  XOR2X1 U7226 ( .IN1(CRC_OUT_7_7), .IN2(n3383), .Q(n6209) );
  AND2X1 U7227 ( .IN1(n6210), .IN2(n4379), .Q(WX3864) );
  XOR2X1 U7228 ( .IN1(CRC_OUT_7_6), .IN2(n3384), .Q(n6210) );
  AND2X1 U7229 ( .IN1(n6211), .IN2(n4379), .Q(WX3862) );
  XOR2X1 U7230 ( .IN1(test_so30), .IN2(DFF_549_n1), .Q(n6211) );
  AND2X1 U7231 ( .IN1(n6212), .IN2(n4380), .Q(WX3860) );
  XOR2X1 U7232 ( .IN1(CRC_OUT_7_4), .IN2(n3385), .Q(n6212) );
  AND2X1 U7233 ( .IN1(n6213), .IN2(n4380), .Q(WX3858) );
  XOR3X1 U7234 ( .IN1(n3190), .IN2(DFF_575_n1), .IN3(DFF_547_n1), .Q(n6213) );
  AND2X1 U7235 ( .IN1(n6214), .IN2(n4380), .Q(WX3856) );
  XOR2X1 U7236 ( .IN1(CRC_OUT_7_2), .IN2(n3386), .Q(n6214) );
  AND2X1 U7237 ( .IN1(n6215), .IN2(n4380), .Q(WX3854) );
  XOR2X1 U7238 ( .IN1(CRC_OUT_7_1), .IN2(n3387), .Q(n6215) );
  AND2X1 U7239 ( .IN1(n6216), .IN2(n4380), .Q(WX3852) );
  XOR2X1 U7240 ( .IN1(CRC_OUT_7_0), .IN2(n3388), .Q(n6216) );
  AND2X1 U7241 ( .IN1(n6217), .IN2(n4380), .Q(WX3850) );
  XOR2X1 U7242 ( .IN1(n3200), .IN2(CRC_OUT_7_31), .Q(n6217) );
  AND2X1 U7243 ( .IN1(test_so24), .IN2(n4380), .Q(WX3324) );
  INVX0 U7244 ( .INP(n6218), .ZN(WX3322) );
  OR2X1 U7245 ( .IN1(n4434), .IN2(n7233), .Q(n6218) );
  INVX0 U7246 ( .INP(n6219), .ZN(WX3320) );
  OR2X1 U7247 ( .IN1(n4434), .IN2(n7235), .Q(n6219) );
  INVX0 U7248 ( .INP(n6220), .ZN(WX3318) );
  OR2X1 U7249 ( .IN1(n4434), .IN2(n7236), .Q(n6220) );
  INVX0 U7250 ( .INP(n6221), .ZN(WX3316) );
  OR2X1 U7251 ( .IN1(n4434), .IN2(n7237), .Q(n6221) );
  INVX0 U7252 ( .INP(n6222), .ZN(WX3314) );
  OR2X1 U7253 ( .IN1(n4434), .IN2(n7238), .Q(n6222) );
  INVX0 U7254 ( .INP(n6223), .ZN(WX3312) );
  OR2X1 U7255 ( .IN1(n4434), .IN2(n7240), .Q(n6223) );
  INVX0 U7256 ( .INP(n6224), .ZN(WX3310) );
  OR2X1 U7257 ( .IN1(n4434), .IN2(n7241), .Q(n6224) );
  INVX0 U7258 ( .INP(n6225), .ZN(WX3308) );
  OR2X1 U7259 ( .IN1(n4434), .IN2(n7242), .Q(n6225) );
  INVX0 U7260 ( .INP(n6226), .ZN(WX3306) );
  OR2X1 U7261 ( .IN1(n4434), .IN2(n7243), .Q(n6226) );
  INVX0 U7262 ( .INP(n6227), .ZN(WX3304) );
  OR2X1 U7263 ( .IN1(n4435), .IN2(n7244), .Q(n6227) );
  INVX0 U7264 ( .INP(n6228), .ZN(WX3302) );
  OR2X1 U7265 ( .IN1(n4435), .IN2(n7245), .Q(n6228) );
  INVX0 U7266 ( .INP(n6229), .ZN(WX3300) );
  OR2X1 U7267 ( .IN1(n4435), .IN2(n7246), .Q(n6229) );
  INVX0 U7268 ( .INP(n6230), .ZN(WX3298) );
  OR2X1 U7269 ( .IN1(n4435), .IN2(n7247), .Q(n6230) );
  INVX0 U7270 ( .INP(n6231), .ZN(WX3296) );
  OR2X1 U7271 ( .IN1(n4435), .IN2(n7248), .Q(n6231) );
  INVX0 U7272 ( .INP(n6232), .ZN(WX3294) );
  OR2X1 U7273 ( .IN1(n4435), .IN2(n7249), .Q(n6232) );
  OR4X1 U7274 ( .IN1(n6233), .IN2(n6234), .IN3(n6235), .IN4(n6236), .Q(WX3292)
         );
  AND2X1 U7275 ( .IN1(n3550), .IN2(n6237), .Q(n6236) );
  AND2X1 U7276 ( .IN1(n5967), .IN2(n3621), .Q(n6235) );
  XOR3X1 U7277 ( .IN1(n3691), .IN2(n3199), .IN3(n6238), .Q(n5967) );
  XOR2X1 U7278 ( .IN1(WX4714), .IN2(test_so36), .Q(n6238) );
  AND2X1 U7279 ( .IN1(n3592), .IN2(CRC_OUT_7_0), .Q(n6234) );
  AND2X1 U7280 ( .IN1(n126), .IN2(n3567), .Q(n6233) );
  INVX0 U7281 ( .INP(n6239), .ZN(n126) );
  OR2X1 U7282 ( .IN1(n4435), .IN2(n3972), .Q(n6239) );
  OR4X1 U7283 ( .IN1(n6240), .IN2(n6241), .IN3(n6242), .IN4(n6243), .Q(WX3290)
         );
  AND2X1 U7284 ( .IN1(n3550), .IN2(n6244), .Q(n6243) );
  AND2X1 U7285 ( .IN1(n3630), .IN2(n5974), .Q(n6242) );
  XNOR3X1 U7286 ( .IN1(n3362), .IN2(n3130), .IN3(n6245), .Q(n5974) );
  XOR2X1 U7287 ( .IN1(WX4648), .IN2(n7179), .Q(n6245) );
  AND2X1 U7288 ( .IN1(n3592), .IN2(CRC_OUT_7_1), .Q(n6241) );
  AND2X1 U7289 ( .IN1(n125), .IN2(n3567), .Q(n6240) );
  INVX0 U7290 ( .INP(n6246), .ZN(n125) );
  OR2X1 U7291 ( .IN1(n4435), .IN2(n3973), .Q(n6246) );
  OR4X1 U7292 ( .IN1(n6247), .IN2(n6248), .IN3(n6249), .IN4(n6250), .Q(WX3288)
         );
  AND2X1 U7293 ( .IN1(n3550), .IN2(n6251), .Q(n6250) );
  AND2X1 U7294 ( .IN1(n3630), .IN2(n5981), .Q(n6249) );
  XNOR3X1 U7295 ( .IN1(n3361), .IN2(n3131), .IN3(n6252), .Q(n5981) );
  XOR2X1 U7296 ( .IN1(WX4646), .IN2(n7180), .Q(n6252) );
  AND2X1 U7297 ( .IN1(n3592), .IN2(CRC_OUT_7_2), .Q(n6248) );
  AND2X1 U7298 ( .IN1(n124), .IN2(n3567), .Q(n6247) );
  INVX0 U7299 ( .INP(n6253), .ZN(n124) );
  OR2X1 U7300 ( .IN1(n4435), .IN2(n3974), .Q(n6253) );
  OR4X1 U7301 ( .IN1(n6254), .IN2(n6255), .IN3(n6256), .IN4(n6257), .Q(WX3286)
         );
  AND2X1 U7302 ( .IN1(n3550), .IN2(n6258), .Q(n6257) );
  AND2X1 U7303 ( .IN1(n3630), .IN2(n5988), .Q(n6256) );
  XNOR3X1 U7304 ( .IN1(n3360), .IN2(n3132), .IN3(n6259), .Q(n5988) );
  XOR2X1 U7305 ( .IN1(WX4644), .IN2(n7181), .Q(n6259) );
  AND2X1 U7306 ( .IN1(n3593), .IN2(CRC_OUT_7_3), .Q(n6255) );
  AND2X1 U7307 ( .IN1(n123), .IN2(n3567), .Q(n6254) );
  INVX0 U7308 ( .INP(n6260), .ZN(n123) );
  OR2X1 U7309 ( .IN1(n4435), .IN2(n3975), .Q(n6260) );
  OR4X1 U7310 ( .IN1(n6261), .IN2(n6262), .IN3(n6263), .IN4(n6264), .Q(WX3284)
         );
  AND2X1 U7311 ( .IN1(n3550), .IN2(n6265), .Q(n6264) );
  AND2X1 U7312 ( .IN1(n3630), .IN2(n5995), .Q(n6263) );
  XNOR3X1 U7313 ( .IN1(n3187), .IN2(n3133), .IN3(n6266), .Q(n5995) );
  XOR2X1 U7314 ( .IN1(WX4642), .IN2(n7182), .Q(n6266) );
  AND2X1 U7315 ( .IN1(n3592), .IN2(CRC_OUT_7_4), .Q(n6262) );
  AND2X1 U7316 ( .IN1(n122), .IN2(n3567), .Q(n6261) );
  INVX0 U7317 ( .INP(n6267), .ZN(n122) );
  OR2X1 U7318 ( .IN1(n4435), .IN2(n3976), .Q(n6267) );
  OR4X1 U7319 ( .IN1(n6268), .IN2(n6269), .IN3(n6270), .IN4(n6271), .Q(WX3282)
         );
  AND2X1 U7320 ( .IN1(n3550), .IN2(n6272), .Q(n6271) );
  AND2X1 U7321 ( .IN1(n3630), .IN2(n6002), .Q(n6270) );
  XNOR3X1 U7322 ( .IN1(n3359), .IN2(n3134), .IN3(n6273), .Q(n6002) );
  XOR2X1 U7323 ( .IN1(WX4640), .IN2(n7183), .Q(n6273) );
  AND2X1 U7324 ( .IN1(n3593), .IN2(CRC_OUT_7_5), .Q(n6269) );
  AND2X1 U7325 ( .IN1(n121), .IN2(n3567), .Q(n6268) );
  INVX0 U7326 ( .INP(n6274), .ZN(n121) );
  OR2X1 U7327 ( .IN1(n4435), .IN2(n3977), .Q(n6274) );
  OR4X1 U7328 ( .IN1(n6275), .IN2(n6276), .IN3(n6277), .IN4(n6278), .Q(WX3280)
         );
  AND2X1 U7329 ( .IN1(n6279), .IN2(n3531), .Q(n6278) );
  AND2X1 U7330 ( .IN1(n3630), .IN2(n6009), .Q(n6277) );
  XNOR3X1 U7331 ( .IN1(n3358), .IN2(n3135), .IN3(n6280), .Q(n6009) );
  XOR2X1 U7332 ( .IN1(WX4638), .IN2(n7184), .Q(n6280) );
  AND2X1 U7333 ( .IN1(n3592), .IN2(CRC_OUT_7_6), .Q(n6276) );
  AND2X1 U7334 ( .IN1(n120), .IN2(n3567), .Q(n6275) );
  INVX0 U7335 ( .INP(n6281), .ZN(n120) );
  OR2X1 U7336 ( .IN1(n4435), .IN2(n3978), .Q(n6281) );
  OR4X1 U7337 ( .IN1(n6282), .IN2(n6283), .IN3(n6284), .IN4(n6285), .Q(WX3278)
         );
  AND2X1 U7338 ( .IN1(n3550), .IN2(n6286), .Q(n6285) );
  AND2X1 U7339 ( .IN1(n3630), .IN2(n6016), .Q(n6284) );
  XNOR3X1 U7340 ( .IN1(n3357), .IN2(n3136), .IN3(n6287), .Q(n6016) );
  XOR2X1 U7341 ( .IN1(WX4636), .IN2(n7185), .Q(n6287) );
  AND2X1 U7342 ( .IN1(n3592), .IN2(CRC_OUT_7_7), .Q(n6283) );
  AND2X1 U7343 ( .IN1(n119), .IN2(n3567), .Q(n6282) );
  INVX0 U7344 ( .INP(n6288), .ZN(n119) );
  OR2X1 U7345 ( .IN1(n4436), .IN2(n3979), .Q(n6288) );
  OR4X1 U7346 ( .IN1(n6289), .IN2(n6290), .IN3(n6291), .IN4(n6292), .Q(WX3276)
         );
  AND2X1 U7347 ( .IN1(n6293), .IN2(n3532), .Q(n6292) );
  AND2X1 U7348 ( .IN1(n3630), .IN2(n6023), .Q(n6291) );
  XNOR3X1 U7349 ( .IN1(n3356), .IN2(n3137), .IN3(n6294), .Q(n6023) );
  XOR2X1 U7350 ( .IN1(WX4634), .IN2(n7186), .Q(n6294) );
  AND2X1 U7351 ( .IN1(n3593), .IN2(CRC_OUT_7_8), .Q(n6290) );
  AND2X1 U7352 ( .IN1(n118), .IN2(n3567), .Q(n6289) );
  INVX0 U7353 ( .INP(n6295), .ZN(n118) );
  OR2X1 U7354 ( .IN1(n4436), .IN2(n3980), .Q(n6295) );
  OR4X1 U7355 ( .IN1(n6296), .IN2(n6297), .IN3(n6298), .IN4(n6299), .Q(WX3274)
         );
  AND2X1 U7356 ( .IN1(n3549), .IN2(n6300), .Q(n6299) );
  AND2X1 U7357 ( .IN1(n3631), .IN2(n6030), .Q(n6298) );
  XNOR3X1 U7358 ( .IN1(n3355), .IN2(n3138), .IN3(n6301), .Q(n6030) );
  XOR2X1 U7359 ( .IN1(WX4632), .IN2(n7187), .Q(n6301) );
  AND2X1 U7360 ( .IN1(n3593), .IN2(CRC_OUT_7_9), .Q(n6297) );
  AND2X1 U7361 ( .IN1(n117), .IN2(n3566), .Q(n6296) );
  INVX0 U7362 ( .INP(n6302), .ZN(n117) );
  OR2X1 U7363 ( .IN1(n4436), .IN2(n3981), .Q(n6302) );
  OR4X1 U7364 ( .IN1(n6303), .IN2(n6304), .IN3(n6305), .IN4(n6306), .Q(WX3272)
         );
  AND2X1 U7365 ( .IN1(n3549), .IN2(n6307), .Q(n6306) );
  AND2X1 U7366 ( .IN1(n3631), .IN2(n6037), .Q(n6305) );
  XNOR3X1 U7367 ( .IN1(n3354), .IN2(n3139), .IN3(n6308), .Q(n6037) );
  XOR2X1 U7368 ( .IN1(WX4630), .IN2(n7188), .Q(n6308) );
  AND2X1 U7369 ( .IN1(test_so31), .IN2(n3588), .Q(n6304) );
  AND2X1 U7370 ( .IN1(n116), .IN2(n3566), .Q(n6303) );
  INVX0 U7371 ( .INP(n6309), .ZN(n116) );
  OR2X1 U7372 ( .IN1(n4429), .IN2(n3982), .Q(n6309) );
  OR4X1 U7373 ( .IN1(n6310), .IN2(n6311), .IN3(n6312), .IN4(n6313), .Q(WX3270)
         );
  AND2X1 U7374 ( .IN1(n3549), .IN2(n6314), .Q(n6313) );
  AND2X1 U7375 ( .IN1(n6044), .IN2(n3621), .Q(n6312) );
  XOR3X1 U7376 ( .IN1(n3713), .IN2(n3140), .IN3(n6315), .Q(n6044) );
  XOR2X1 U7377 ( .IN1(WX4564), .IN2(test_so41), .Q(n6315) );
  AND2X1 U7378 ( .IN1(n3593), .IN2(CRC_OUT_7_11), .Q(n6311) );
  AND2X1 U7379 ( .IN1(n115), .IN2(n3566), .Q(n6310) );
  INVX0 U7380 ( .INP(n6316), .ZN(n115) );
  OR2X1 U7381 ( .IN1(n4429), .IN2(n3983), .Q(n6316) );
  OR4X1 U7382 ( .IN1(n6317), .IN2(n6318), .IN3(n6319), .IN4(n6320), .Q(WX3268)
         );
  AND2X1 U7383 ( .IN1(n6321), .IN2(n3532), .Q(n6320) );
  AND2X1 U7384 ( .IN1(n3631), .IN2(n6051), .Q(n6319) );
  XNOR3X1 U7385 ( .IN1(n3353), .IN2(n3141), .IN3(n6322), .Q(n6051) );
  XOR2X1 U7386 ( .IN1(WX4626), .IN2(n7189), .Q(n6322) );
  AND2X1 U7387 ( .IN1(n3593), .IN2(CRC_OUT_7_12), .Q(n6318) );
  AND2X1 U7388 ( .IN1(n114), .IN2(n3566), .Q(n6317) );
  INVX0 U7389 ( .INP(n6323), .ZN(n114) );
  OR2X1 U7390 ( .IN1(n4429), .IN2(n3984), .Q(n6323) );
  OR4X1 U7391 ( .IN1(n6324), .IN2(n6325), .IN3(n6326), .IN4(n6327), .Q(WX3266)
         );
  AND2X1 U7392 ( .IN1(n3549), .IN2(n6328), .Q(n6327) );
  AND2X1 U7393 ( .IN1(n6058), .IN2(n3621), .Q(n6326) );
  XOR3X1 U7394 ( .IN1(n3717), .IN2(n3352), .IN3(n6329), .Q(n6058) );
  XOR2X1 U7395 ( .IN1(WX4560), .IN2(test_so39), .Q(n6329) );
  AND2X1 U7396 ( .IN1(n3593), .IN2(CRC_OUT_7_13), .Q(n6325) );
  AND2X1 U7397 ( .IN1(n113), .IN2(n3566), .Q(n6324) );
  INVX0 U7398 ( .INP(n6330), .ZN(n113) );
  OR2X1 U7399 ( .IN1(n4429), .IN2(n3985), .Q(n6330) );
  OR4X1 U7400 ( .IN1(n6331), .IN2(n6332), .IN3(n6333), .IN4(n6334), .Q(WX3264)
         );
  AND2X1 U7401 ( .IN1(n3549), .IN2(n6335), .Q(n6334) );
  AND2X1 U7402 ( .IN1(n3631), .IN2(n6065), .Q(n6333) );
  XNOR3X1 U7403 ( .IN1(n3351), .IN2(n3142), .IN3(n6336), .Q(n6065) );
  XOR2X1 U7404 ( .IN1(WX4622), .IN2(n7190), .Q(n6336) );
  AND2X1 U7405 ( .IN1(n3593), .IN2(CRC_OUT_7_14), .Q(n6332) );
  AND2X1 U7406 ( .IN1(n112), .IN2(n3566), .Q(n6331) );
  INVX0 U7407 ( .INP(n6337), .ZN(n112) );
  OR2X1 U7408 ( .IN1(n4429), .IN2(n3986), .Q(n6337) );
  OR4X1 U7409 ( .IN1(n6338), .IN2(n6339), .IN3(n6340), .IN4(n6341), .Q(WX3262)
         );
  AND2X1 U7410 ( .IN1(n3549), .IN2(n6342), .Q(n6341) );
  AND2X1 U7411 ( .IN1(n6072), .IN2(n3621), .Q(n6340) );
  XOR3X1 U7412 ( .IN1(n3350), .IN2(n3143), .IN3(n6343), .Q(n6072) );
  XOR2X1 U7413 ( .IN1(WX4556), .IN2(test_so37), .Q(n6343) );
  AND2X1 U7414 ( .IN1(n3593), .IN2(CRC_OUT_7_15), .Q(n6339) );
  AND2X1 U7415 ( .IN1(n110), .IN2(n3566), .Q(n6338) );
  INVX0 U7416 ( .INP(n6344), .ZN(n110) );
  OR2X1 U7417 ( .IN1(n4429), .IN2(n3987), .Q(n6344) );
  OR4X1 U7418 ( .IN1(n6345), .IN2(n6346), .IN3(n6347), .IN4(n6348), .Q(WX3260)
         );
  AND2X1 U7419 ( .IN1(n6349), .IN2(n3533), .Q(n6348) );
  AND2X1 U7420 ( .IN1(n3631), .IN2(n6079), .Q(n6347) );
  XOR3X1 U7421 ( .IN1(n2979), .IN2(n3515), .IN3(n6350), .Q(n6079) );
  XOR3X1 U7422 ( .IN1(n7191), .IN2(n3186), .IN3(WX4682), .Q(n6350) );
  AND2X1 U7423 ( .IN1(n3593), .IN2(CRC_OUT_7_16), .Q(n6346) );
  AND2X1 U7424 ( .IN1(n109), .IN2(n3566), .Q(n6345) );
  INVX0 U7425 ( .INP(n6351), .ZN(n109) );
  OR2X1 U7426 ( .IN1(n4429), .IN2(n3988), .Q(n6351) );
  OR4X1 U7427 ( .IN1(n6352), .IN2(n6353), .IN3(n6354), .IN4(n6355), .Q(WX3258)
         );
  AND2X1 U7428 ( .IN1(n3549), .IN2(n6356), .Q(n6355) );
  AND2X1 U7429 ( .IN1(n6086), .IN2(n3621), .Q(n6354) );
  XOR3X1 U7430 ( .IN1(n2981), .IN2(TM1), .IN3(n6357), .Q(n6086) );
  XNOR3X1 U7431 ( .IN1(test_so35), .IN2(n7192), .IN3(n3349), .Q(n6357) );
  AND2X1 U7432 ( .IN1(n3593), .IN2(CRC_OUT_7_17), .Q(n6353) );
  AND2X1 U7433 ( .IN1(n108), .IN2(n3566), .Q(n6352) );
  INVX0 U7434 ( .INP(n6358), .ZN(n108) );
  OR2X1 U7435 ( .IN1(n4429), .IN2(n3989), .Q(n6358) );
  OR4X1 U7436 ( .IN1(n6359), .IN2(n6360), .IN3(n6361), .IN4(n6362), .Q(WX3256)
         );
  AND2X1 U7437 ( .IN1(n3549), .IN2(n6363), .Q(n6362) );
  AND2X1 U7438 ( .IN1(n3631), .IN2(n6093), .Q(n6361) );
  XOR3X1 U7439 ( .IN1(n2982), .IN2(n3514), .IN3(n6364), .Q(n6093) );
  XOR3X1 U7440 ( .IN1(n7193), .IN2(n3348), .IN3(WX4678), .Q(n6364) );
  AND2X1 U7441 ( .IN1(n3594), .IN2(CRC_OUT_7_18), .Q(n6360) );
  AND2X1 U7442 ( .IN1(n107), .IN2(n3566), .Q(n6359) );
  INVX0 U7443 ( .INP(n6365), .ZN(n107) );
  OR2X1 U7444 ( .IN1(n4429), .IN2(n3990), .Q(n6365) );
  OR4X1 U7445 ( .IN1(n6366), .IN2(n6367), .IN3(n6368), .IN4(n6369), .Q(WX3254)
         );
  AND2X1 U7446 ( .IN1(n3549), .IN2(n6370), .Q(n6369) );
  AND2X1 U7447 ( .IN1(n3631), .IN2(n6100), .Q(n6368) );
  XOR3X1 U7448 ( .IN1(n2984), .IN2(n3518), .IN3(n6371), .Q(n6100) );
  XOR3X1 U7449 ( .IN1(n7194), .IN2(n3347), .IN3(WX4676), .Q(n6371) );
  AND2X1 U7450 ( .IN1(n3593), .IN2(CRC_OUT_7_19), .Q(n6367) );
  AND2X1 U7451 ( .IN1(n106), .IN2(n3566), .Q(n6366) );
  INVX0 U7452 ( .INP(n6372), .ZN(n106) );
  OR2X1 U7453 ( .IN1(n4428), .IN2(n3991), .Q(n6372) );
  OR4X1 U7454 ( .IN1(n6373), .IN2(n6374), .IN3(n6375), .IN4(n6376), .Q(WX3252)
         );
  AND2X1 U7455 ( .IN1(n3549), .IN2(n6377), .Q(n6376) );
  AND2X1 U7456 ( .IN1(n3631), .IN2(n6107), .Q(n6375) );
  XOR3X1 U7457 ( .IN1(n2986), .IN2(n3516), .IN3(n6378), .Q(n6107) );
  XOR3X1 U7458 ( .IN1(n7195), .IN2(n3346), .IN3(WX4674), .Q(n6378) );
  AND2X1 U7459 ( .IN1(n3594), .IN2(CRC_OUT_7_20), .Q(n6374) );
  AND2X1 U7460 ( .IN1(n105), .IN2(n3566), .Q(n6373) );
  INVX0 U7461 ( .INP(n6379), .ZN(n105) );
  OR2X1 U7462 ( .IN1(n4428), .IN2(n3992), .Q(n6379) );
  OR4X1 U7463 ( .IN1(n6380), .IN2(n6381), .IN3(n6382), .IN4(n6383), .Q(WX3250)
         );
  AND2X1 U7464 ( .IN1(n3549), .IN2(n6384), .Q(n6383) );
  AND2X1 U7465 ( .IN1(n3631), .IN2(n6114), .Q(n6382) );
  XOR3X1 U7466 ( .IN1(n2988), .IN2(n3515), .IN3(n6385), .Q(n6114) );
  XOR3X1 U7467 ( .IN1(n7196), .IN2(n3345), .IN3(WX4672), .Q(n6385) );
  AND2X1 U7468 ( .IN1(n3594), .IN2(CRC_OUT_7_21), .Q(n6381) );
  AND2X1 U7469 ( .IN1(n104), .IN2(n3565), .Q(n6380) );
  INVX0 U7470 ( .INP(n6386), .ZN(n104) );
  OR2X1 U7471 ( .IN1(n4428), .IN2(n3993), .Q(n6386) );
  OR4X1 U7472 ( .IN1(n6387), .IN2(n6388), .IN3(n6389), .IN4(n6390), .Q(WX3248)
         );
  AND2X1 U7473 ( .IN1(n3549), .IN2(n6391), .Q(n6390) );
  AND2X1 U7474 ( .IN1(n3631), .IN2(n6121), .Q(n6389) );
  XOR3X1 U7475 ( .IN1(n2990), .IN2(n3514), .IN3(n6392), .Q(n6121) );
  XOR3X1 U7476 ( .IN1(n7197), .IN2(n3344), .IN3(WX4670), .Q(n6392) );
  AND2X1 U7477 ( .IN1(n3594), .IN2(CRC_OUT_7_22), .Q(n6388) );
  AND2X1 U7478 ( .IN1(n103), .IN2(n3565), .Q(n6387) );
  INVX0 U7479 ( .INP(n6393), .ZN(n103) );
  OR2X1 U7480 ( .IN1(n4428), .IN2(n3994), .Q(n6393) );
  OR4X1 U7481 ( .IN1(n6394), .IN2(n6395), .IN3(n6396), .IN4(n6397), .Q(WX3246)
         );
  AND2X1 U7482 ( .IN1(n6398), .IN2(n3534), .Q(n6397) );
  AND2X1 U7483 ( .IN1(n3634), .IN2(n6128), .Q(n6396) );
  XOR3X1 U7484 ( .IN1(n2992), .IN2(n3518), .IN3(n6399), .Q(n6128) );
  XOR3X1 U7485 ( .IN1(n7198), .IN2(n3343), .IN3(WX4668), .Q(n6399) );
  AND2X1 U7486 ( .IN1(n3599), .IN2(CRC_OUT_7_23), .Q(n6395) );
  AND2X1 U7487 ( .IN1(n102), .IN2(n3565), .Q(n6394) );
  INVX0 U7488 ( .INP(n6400), .ZN(n102) );
  OR2X1 U7489 ( .IN1(n4428), .IN2(n3995), .Q(n6400) );
  OR4X1 U7490 ( .IN1(n6401), .IN2(n6402), .IN3(n6403), .IN4(n6404), .Q(WX3244)
         );
  AND2X1 U7491 ( .IN1(n3548), .IN2(n6405), .Q(n6404) );
  AND2X1 U7492 ( .IN1(n3631), .IN2(n6135), .Q(n6403) );
  XOR3X1 U7493 ( .IN1(n2994), .IN2(n3516), .IN3(n6406), .Q(n6135) );
  XOR3X1 U7494 ( .IN1(n7199), .IN2(n3342), .IN3(WX4666), .Q(n6406) );
  AND2X1 U7495 ( .IN1(n3594), .IN2(CRC_OUT_7_24), .Q(n6402) );
  AND2X1 U7496 ( .IN1(n101), .IN2(n3565), .Q(n6401) );
  INVX0 U7497 ( .INP(n6407), .ZN(n101) );
  OR2X1 U7498 ( .IN1(n4428), .IN2(n3996), .Q(n6407) );
  OR4X1 U7499 ( .IN1(n6408), .IN2(n6409), .IN3(n6410), .IN4(n6411), .Q(WX3242)
         );
  AND2X1 U7500 ( .IN1(n3548), .IN2(n6412), .Q(n6411) );
  AND2X1 U7501 ( .IN1(n3631), .IN2(n6142), .Q(n6410) );
  XOR3X1 U7502 ( .IN1(n2996), .IN2(n3515), .IN3(n6413), .Q(n6142) );
  XOR3X1 U7503 ( .IN1(n7200), .IN2(n3341), .IN3(WX4664), .Q(n6413) );
  AND2X1 U7504 ( .IN1(n3594), .IN2(CRC_OUT_7_25), .Q(n6409) );
  AND2X1 U7505 ( .IN1(n100), .IN2(n3565), .Q(n6408) );
  INVX0 U7506 ( .INP(n6414), .ZN(n100) );
  OR2X1 U7507 ( .IN1(n4428), .IN2(n3997), .Q(n6414) );
  OR4X1 U7508 ( .IN1(n6415), .IN2(n6416), .IN3(n6417), .IN4(n6418), .Q(WX3240)
         );
  AND2X1 U7509 ( .IN1(n6419), .IN2(n3533), .Q(n6418) );
  AND2X1 U7510 ( .IN1(n3631), .IN2(n6149), .Q(n6417) );
  XOR3X1 U7511 ( .IN1(n2998), .IN2(n3514), .IN3(n6420), .Q(n6149) );
  XOR3X1 U7512 ( .IN1(n7201), .IN2(n3340), .IN3(WX4662), .Q(n6420) );
  AND2X1 U7513 ( .IN1(n3594), .IN2(CRC_OUT_7_26), .Q(n6416) );
  AND2X1 U7514 ( .IN1(n99), .IN2(n3565), .Q(n6415) );
  INVX0 U7515 ( .INP(n6421), .ZN(n99) );
  OR2X1 U7516 ( .IN1(n4428), .IN2(n3998), .Q(n6421) );
  OR4X1 U7517 ( .IN1(n6422), .IN2(n6423), .IN3(n6424), .IN4(n6425), .Q(WX3238)
         );
  AND2X1 U7518 ( .IN1(n3548), .IN2(n6426), .Q(n6425) );
  AND2X1 U7519 ( .IN1(n3632), .IN2(n6156), .Q(n6424) );
  XOR3X1 U7520 ( .IN1(n3000), .IN2(n3518), .IN3(n6427), .Q(n6156) );
  XOR3X1 U7521 ( .IN1(n7202), .IN2(n3339), .IN3(WX4660), .Q(n6427) );
  AND2X1 U7522 ( .IN1(test_so32), .IN2(n3587), .Q(n6423) );
  AND2X1 U7523 ( .IN1(n98), .IN2(n3565), .Q(n6422) );
  INVX0 U7524 ( .INP(n6428), .ZN(n98) );
  OR2X1 U7525 ( .IN1(n4428), .IN2(n3999), .Q(n6428) );
  OR4X1 U7526 ( .IN1(n6429), .IN2(n6430), .IN3(n6431), .IN4(n6432), .Q(WX3236)
         );
  AND2X1 U7527 ( .IN1(n3548), .IN2(n6433), .Q(n6432) );
  AND2X1 U7528 ( .IN1(n6163), .IN2(n3622), .Q(n6431) );
  XOR3X1 U7529 ( .IN1(n3002), .IN2(TM1), .IN3(n6434), .Q(n6163) );
  XOR3X1 U7530 ( .IN1(test_so40), .IN2(n7203), .IN3(WX4658), .Q(n6434) );
  AND2X1 U7531 ( .IN1(n3594), .IN2(CRC_OUT_7_28), .Q(n6430) );
  AND2X1 U7532 ( .IN1(n97), .IN2(n3565), .Q(n6429) );
  INVX0 U7533 ( .INP(n6435), .ZN(n97) );
  OR2X1 U7534 ( .IN1(n4428), .IN2(n4000), .Q(n6435) );
  OR4X1 U7535 ( .IN1(n6436), .IN2(n6437), .IN3(n6438), .IN4(n6439), .Q(WX3234)
         );
  AND2X1 U7536 ( .IN1(n3548), .IN2(n6440), .Q(n6439) );
  AND2X1 U7537 ( .IN1(n3632), .IN2(n6170), .Q(n6438) );
  XOR3X1 U7538 ( .IN1(n3003), .IN2(n3516), .IN3(n6441), .Q(n6170) );
  XOR3X1 U7539 ( .IN1(n7204), .IN2(n3338), .IN3(WX4656), .Q(n6441) );
  AND2X1 U7540 ( .IN1(n3594), .IN2(CRC_OUT_7_29), .Q(n6437) );
  AND2X1 U7541 ( .IN1(n96), .IN2(n3565), .Q(n6436) );
  INVX0 U7542 ( .INP(n6442), .ZN(n96) );
  OR2X1 U7543 ( .IN1(n4428), .IN2(n4001), .Q(n6442) );
  OR4X1 U7544 ( .IN1(n6443), .IN2(n6444), .IN3(n6445), .IN4(n6446), .Q(WX3232)
         );
  AND2X1 U7545 ( .IN1(n6447), .IN2(n3533), .Q(n6446) );
  AND2X1 U7546 ( .IN1(n6177), .IN2(n3622), .Q(n6445) );
  XOR3X1 U7547 ( .IN1(n3005), .IN2(TM1), .IN3(n6448), .Q(n6177) );
  XNOR3X1 U7548 ( .IN1(test_so38), .IN2(n7205), .IN3(n3337), .Q(n6448) );
  AND2X1 U7549 ( .IN1(n3594), .IN2(CRC_OUT_7_30), .Q(n6444) );
  AND2X1 U7550 ( .IN1(n95), .IN2(n3565), .Q(n6443) );
  INVX0 U7551 ( .INP(n6449), .ZN(n95) );
  OR2X1 U7552 ( .IN1(n4428), .IN2(n4002), .Q(n6449) );
  OR4X1 U7553 ( .IN1(n6450), .IN2(n6451), .IN3(n6452), .IN4(n6453), .Q(WX3230)
         );
  AND2X1 U7554 ( .IN1(n3548), .IN2(n6454), .Q(n6453) );
  AND2X1 U7555 ( .IN1(n3632), .IN2(n6184), .Q(n6452) );
  XOR3X1 U7556 ( .IN1(n2841), .IN2(n3515), .IN3(n6455), .Q(n6184) );
  XOR3X1 U7557 ( .IN1(n7206), .IN2(n3336), .IN3(WX4652), .Q(n6455) );
  AND2X1 U7558 ( .IN1(n2245), .IN2(WX3071), .Q(n6451) );
  AND2X1 U7559 ( .IN1(n3594), .IN2(CRC_OUT_7_31), .Q(n6450) );
  AND2X1 U7560 ( .IN1(n3498), .IN2(n4380), .Q(WX3132) );
  AND2X1 U7561 ( .IN1(n6456), .IN2(n4380), .Q(WX2619) );
  XOR2X1 U7562 ( .IN1(CRC_OUT_8_30), .IN2(n3389), .Q(n6456) );
  AND2X1 U7563 ( .IN1(n6457), .IN2(n4381), .Q(WX2617) );
  XOR2X1 U7564 ( .IN1(CRC_OUT_8_29), .IN2(n3390), .Q(n6457) );
  AND2X1 U7565 ( .IN1(n6458), .IN2(n4381), .Q(WX2615) );
  XOR2X1 U7566 ( .IN1(CRC_OUT_8_28), .IN2(n3391), .Q(n6458) );
  AND2X1 U7567 ( .IN1(n6459), .IN2(n4381), .Q(WX2613) );
  XOR2X1 U7568 ( .IN1(test_so18), .IN2(DFF_379_n1), .Q(n6459) );
  AND2X1 U7569 ( .IN1(n6460), .IN2(n4381), .Q(WX2611) );
  XOR2X1 U7570 ( .IN1(CRC_OUT_8_26), .IN2(n3392), .Q(n6460) );
  AND2X1 U7571 ( .IN1(n6461), .IN2(n4381), .Q(WX2609) );
  XOR2X1 U7572 ( .IN1(test_so21), .IN2(n3393), .Q(n6461) );
  AND2X1 U7573 ( .IN1(n6462), .IN2(n4381), .Q(WX2607) );
  XOR2X1 U7574 ( .IN1(CRC_OUT_8_24), .IN2(n3394), .Q(n6462) );
  AND2X1 U7575 ( .IN1(n6463), .IN2(n4381), .Q(WX2605) );
  XOR2X1 U7576 ( .IN1(CRC_OUT_8_23), .IN2(n3395), .Q(n6463) );
  AND2X1 U7577 ( .IN1(n6464), .IN2(n4381), .Q(WX2603) );
  XOR2X1 U7578 ( .IN1(CRC_OUT_8_22), .IN2(n3396), .Q(n6464) );
  AND2X1 U7579 ( .IN1(n6465), .IN2(n4382), .Q(WX2601) );
  XOR2X1 U7580 ( .IN1(CRC_OUT_8_21), .IN2(n3397), .Q(n6465) );
  AND2X1 U7581 ( .IN1(n6466), .IN2(n4382), .Q(WX2599) );
  XOR2X1 U7582 ( .IN1(CRC_OUT_8_20), .IN2(n3398), .Q(n6466) );
  AND2X1 U7583 ( .IN1(n6467), .IN2(n4382), .Q(WX2597) );
  XOR2X1 U7584 ( .IN1(CRC_OUT_8_19), .IN2(n3399), .Q(n6467) );
  AND2X1 U7585 ( .IN1(n6468), .IN2(n4382), .Q(WX2595) );
  XOR2X1 U7586 ( .IN1(CRC_OUT_8_18), .IN2(n3400), .Q(n6468) );
  AND2X1 U7587 ( .IN1(n6469), .IN2(n4382), .Q(WX2593) );
  XOR2X1 U7588 ( .IN1(CRC_OUT_8_17), .IN2(n3401), .Q(n6469) );
  AND2X1 U7589 ( .IN1(n6470), .IN2(n4382), .Q(WX2591) );
  XOR2X1 U7590 ( .IN1(CRC_OUT_8_16), .IN2(n3402), .Q(n6470) );
  AND2X1 U7591 ( .IN1(n6471), .IN2(n4382), .Q(WX2589) );
  XOR3X1 U7592 ( .IN1(n3191), .IN2(DFF_383_n1), .IN3(DFF_367_n1), .Q(n6471) );
  AND2X1 U7593 ( .IN1(n6472), .IN2(n4382), .Q(WX2587) );
  XOR2X1 U7594 ( .IN1(CRC_OUT_8_14), .IN2(n3403), .Q(n6472) );
  AND2X1 U7595 ( .IN1(n6473), .IN2(n4383), .Q(WX2585) );
  XOR2X1 U7596 ( .IN1(CRC_OUT_8_13), .IN2(n3404), .Q(n6473) );
  AND2X1 U7597 ( .IN1(n6474), .IN2(n4382), .Q(WX2583) );
  XOR2X1 U7598 ( .IN1(CRC_OUT_8_12), .IN2(n3405), .Q(n6474) );
  AND2X1 U7599 ( .IN1(n6475), .IN2(n4384), .Q(WX2581) );
  XOR2X1 U7600 ( .IN1(CRC_OUT_8_11), .IN2(n3406), .Q(n6475) );
  AND2X1 U7601 ( .IN1(n6476), .IN2(n4383), .Q(WX2579) );
  XOR3X1 U7602 ( .IN1(n3192), .IN2(DFF_383_n1), .IN3(DFF_362_n1), .Q(n6476) );
  AND2X1 U7603 ( .IN1(n6477), .IN2(n4383), .Q(WX2577) );
  XOR2X1 U7604 ( .IN1(test_so19), .IN2(DFF_361_n1), .Q(n6477) );
  AND2X1 U7605 ( .IN1(n6478), .IN2(n4383), .Q(WX2575) );
  XOR2X1 U7606 ( .IN1(CRC_OUT_8_8), .IN2(n3407), .Q(n6478) );
  AND2X1 U7607 ( .IN1(n6479), .IN2(n4383), .Q(WX2573) );
  XOR2X1 U7608 ( .IN1(test_so20), .IN2(n3408), .Q(n6479) );
  AND2X1 U7609 ( .IN1(n6480), .IN2(n4384), .Q(WX2571) );
  XOR2X1 U7610 ( .IN1(CRC_OUT_8_6), .IN2(n3409), .Q(n6480) );
  AND2X1 U7611 ( .IN1(n6481), .IN2(n4383), .Q(WX2569) );
  XOR2X1 U7612 ( .IN1(CRC_OUT_8_5), .IN2(n3410), .Q(n6481) );
  AND2X1 U7613 ( .IN1(n6482), .IN2(n4384), .Q(WX2567) );
  XOR2X1 U7614 ( .IN1(CRC_OUT_8_4), .IN2(n3411), .Q(n6482) );
  AND2X1 U7615 ( .IN1(n6483), .IN2(n4383), .Q(WX2565) );
  XOR3X1 U7616 ( .IN1(n3193), .IN2(DFF_383_n1), .IN3(DFF_355_n1), .Q(n6483) );
  AND2X1 U7617 ( .IN1(n6484), .IN2(n4384), .Q(WX2563) );
  XOR2X1 U7618 ( .IN1(CRC_OUT_8_2), .IN2(n3412), .Q(n6484) );
  AND2X1 U7619 ( .IN1(n6485), .IN2(n4384), .Q(WX2561) );
  XOR2X1 U7620 ( .IN1(CRC_OUT_8_1), .IN2(n3413), .Q(n6485) );
  AND2X1 U7621 ( .IN1(n6486), .IN2(n4384), .Q(WX2559) );
  XOR2X1 U7622 ( .IN1(CRC_OUT_8_0), .IN2(n3414), .Q(n6486) );
  AND2X1 U7623 ( .IN1(n6487), .IN2(n4384), .Q(WX2557) );
  XOR2X1 U7624 ( .IN1(n3201), .IN2(CRC_OUT_8_31), .Q(n6487) );
  AND2X1 U7625 ( .IN1(n4386), .IN2(n8653), .Q(WX2031) );
  AND2X1 U7626 ( .IN1(n4386), .IN2(n8654), .Q(WX2029) );
  INVX0 U7627 ( .INP(n6488), .ZN(WX2027) );
  OR2X1 U7628 ( .IN1(n4428), .IN2(n7234), .Q(n6488) );
  AND2X1 U7629 ( .IN1(n4386), .IN2(n8656), .Q(WX2025) );
  AND2X1 U7630 ( .IN1(n4387), .IN2(n8657), .Q(WX2023) );
  AND2X1 U7631 ( .IN1(n4386), .IN2(n8658), .Q(WX2021) );
  AND2X1 U7632 ( .IN1(test_so13), .IN2(n4383), .Q(WX2019) );
  AND2X1 U7633 ( .IN1(n4386), .IN2(n8661), .Q(WX2017) );
  AND2X1 U7634 ( .IN1(n4386), .IN2(n8662), .Q(WX2015) );
  AND2X1 U7635 ( .IN1(n4387), .IN2(n8663), .Q(WX2013) );
  AND2X1 U7636 ( .IN1(n4387), .IN2(n8664), .Q(WX2011) );
  AND2X1 U7637 ( .IN1(n4387), .IN2(n8665), .Q(WX2009) );
  AND2X1 U7638 ( .IN1(n4387), .IN2(n8666), .Q(WX2007) );
  AND2X1 U7639 ( .IN1(n4387), .IN2(n8667), .Q(WX2005) );
  AND2X1 U7640 ( .IN1(n4387), .IN2(n8668), .Q(WX2003) );
  AND2X1 U7641 ( .IN1(n4387), .IN2(n8669), .Q(WX2001) );
  OR4X1 U7642 ( .IN1(n6489), .IN2(n6490), .IN3(n6491), .IN4(n6492), .Q(WX1999)
         );
  AND2X1 U7643 ( .IN1(n3632), .IN2(n6237), .Q(n6492) );
  XNOR3X1 U7644 ( .IN1(n3200), .IN2(n3144), .IN3(n6493), .Q(n6237) );
  XOR2X1 U7645 ( .IN1(WX3357), .IN2(n7207), .Q(n6493) );
  AND2X1 U7646 ( .IN1(n5458), .IN2(n3533), .Q(n6491) );
  XOR3X1 U7647 ( .IN1(n3201), .IN2(n3159), .IN3(n6494), .Q(n5458) );
  XOR2X1 U7648 ( .IN1(WX2000), .IN2(test_so16), .Q(n6494) );
  AND2X1 U7649 ( .IN1(n3594), .IN2(CRC_OUT_8_0), .Q(n6490) );
  AND2X1 U7650 ( .IN1(n63), .IN2(n3565), .Q(n6489) );
  INVX0 U7651 ( .INP(n6495), .ZN(n63) );
  OR2X1 U7652 ( .IN1(n4427), .IN2(n4003), .Q(n6495) );
  OR4X1 U7653 ( .IN1(n6496), .IN2(n6497), .IN3(n6498), .IN4(n6499), .Q(WX1997)
         );
  AND2X1 U7654 ( .IN1(n3632), .IN2(n6244), .Q(n6499) );
  XNOR3X1 U7655 ( .IN1(n3388), .IN2(n3145), .IN3(n6500), .Q(n6244) );
  XOR2X1 U7656 ( .IN1(WX3355), .IN2(n7209), .Q(n6500) );
  AND2X1 U7657 ( .IN1(n3548), .IN2(n5464), .Q(n6498) );
  XNOR3X1 U7658 ( .IN1(n3414), .IN2(n3160), .IN3(n6501), .Q(n5464) );
  XOR2X1 U7659 ( .IN1(WX2062), .IN2(n7208), .Q(n6501) );
  AND2X1 U7660 ( .IN1(n3595), .IN2(CRC_OUT_8_1), .Q(n6497) );
  AND2X1 U7661 ( .IN1(n62), .IN2(n3565), .Q(n6496) );
  INVX0 U7662 ( .INP(n6502), .ZN(n62) );
  OR2X1 U7663 ( .IN1(n4427), .IN2(n4004), .Q(n6502) );
  OR4X1 U7664 ( .IN1(n6503), .IN2(n6504), .IN3(n6505), .IN4(n6506), .Q(WX1995)
         );
  AND2X1 U7665 ( .IN1(n3632), .IN2(n6251), .Q(n6506) );
  XNOR3X1 U7666 ( .IN1(n3387), .IN2(n3146), .IN3(n6507), .Q(n6251) );
  XOR2X1 U7667 ( .IN1(WX3353), .IN2(n7211), .Q(n6507) );
  AND2X1 U7668 ( .IN1(n3548), .IN2(n5470), .Q(n6505) );
  XNOR3X1 U7669 ( .IN1(n3413), .IN2(n3161), .IN3(n6508), .Q(n5470) );
  XOR2X1 U7670 ( .IN1(WX2060), .IN2(n7210), .Q(n6508) );
  AND2X1 U7671 ( .IN1(n3595), .IN2(CRC_OUT_8_2), .Q(n6504) );
  AND2X1 U7672 ( .IN1(n61), .IN2(n3564), .Q(n6503) );
  INVX0 U7673 ( .INP(n6509), .ZN(n61) );
  OR2X1 U7674 ( .IN1(n4427), .IN2(n4005), .Q(n6509) );
  OR4X1 U7675 ( .IN1(n6510), .IN2(n6511), .IN3(n6512), .IN4(n6513), .Q(WX1993)
         );
  AND2X1 U7676 ( .IN1(n3632), .IN2(n6258), .Q(n6513) );
  XNOR3X1 U7677 ( .IN1(n3386), .IN2(n3147), .IN3(n6514), .Q(n6258) );
  XOR2X1 U7678 ( .IN1(WX3351), .IN2(n7213), .Q(n6514) );
  AND2X1 U7679 ( .IN1(n3548), .IN2(n5476), .Q(n6512) );
  XNOR3X1 U7680 ( .IN1(n3412), .IN2(n3162), .IN3(n6515), .Q(n5476) );
  XOR2X1 U7681 ( .IN1(WX2058), .IN2(n7212), .Q(n6515) );
  AND2X1 U7682 ( .IN1(n3595), .IN2(CRC_OUT_8_3), .Q(n6511) );
  AND2X1 U7683 ( .IN1(n60), .IN2(n3564), .Q(n6510) );
  INVX0 U7684 ( .INP(n6516), .ZN(n60) );
  OR2X1 U7685 ( .IN1(n4427), .IN2(n4006), .Q(n6516) );
  OR4X1 U7686 ( .IN1(n6517), .IN2(n6518), .IN3(n6519), .IN4(n6520), .Q(WX1991)
         );
  AND2X1 U7687 ( .IN1(n3632), .IN2(n6265), .Q(n6520) );
  XNOR3X1 U7688 ( .IN1(n3190), .IN2(n3148), .IN3(n6521), .Q(n6265) );
  XOR2X1 U7689 ( .IN1(WX3349), .IN2(n7214), .Q(n6521) );
  AND2X1 U7690 ( .IN1(n5482), .IN2(n3533), .Q(n6519) );
  XOR3X1 U7691 ( .IN1(n3763), .IN2(n3193), .IN3(n6522), .Q(n5482) );
  XOR2X1 U7692 ( .IN1(WX2120), .IN2(test_so14), .Q(n6522) );
  AND2X1 U7693 ( .IN1(n3595), .IN2(CRC_OUT_8_4), .Q(n6518) );
  AND2X1 U7694 ( .IN1(n59), .IN2(n3564), .Q(n6517) );
  INVX0 U7695 ( .INP(n6523), .ZN(n59) );
  OR2X1 U7696 ( .IN1(n4427), .IN2(n4007), .Q(n6523) );
  OR4X1 U7697 ( .IN1(n6524), .IN2(n6525), .IN3(n6526), .IN4(n6527), .Q(WX1989)
         );
  AND2X1 U7698 ( .IN1(n3632), .IN2(n6272), .Q(n6527) );
  XNOR3X1 U7699 ( .IN1(n3385), .IN2(n3149), .IN3(n6528), .Q(n6272) );
  XOR2X1 U7700 ( .IN1(WX3347), .IN2(n7216), .Q(n6528) );
  AND2X1 U7701 ( .IN1(n3548), .IN2(n5488), .Q(n6526) );
  XNOR3X1 U7702 ( .IN1(n3411), .IN2(n3163), .IN3(n6529), .Q(n5488) );
  XOR2X1 U7703 ( .IN1(WX2054), .IN2(n7215), .Q(n6529) );
  AND2X1 U7704 ( .IN1(n3595), .IN2(CRC_OUT_8_5), .Q(n6525) );
  AND2X1 U7705 ( .IN1(n58), .IN2(n3564), .Q(n6524) );
  INVX0 U7706 ( .INP(n6530), .ZN(n58) );
  OR2X1 U7707 ( .IN1(n4427), .IN2(n4008), .Q(n6530) );
  OR4X1 U7708 ( .IN1(n6531), .IN2(n6532), .IN3(n6533), .IN4(n6534), .Q(WX1987)
         );
  AND2X1 U7709 ( .IN1(n6279), .IN2(n3623), .Q(n6534) );
  XOR3X1 U7710 ( .IN1(n3735), .IN2(n3150), .IN3(n6535), .Q(n6279) );
  XOR2X1 U7711 ( .IN1(WX3281), .IN2(test_so30), .Q(n6535) );
  AND2X1 U7712 ( .IN1(n3548), .IN2(n5494), .Q(n6533) );
  XNOR3X1 U7713 ( .IN1(n3410), .IN2(n3164), .IN3(n6536), .Q(n5494) );
  XOR2X1 U7714 ( .IN1(WX2052), .IN2(n7217), .Q(n6536) );
  AND2X1 U7715 ( .IN1(n3595), .IN2(CRC_OUT_8_6), .Q(n6532) );
  AND2X1 U7716 ( .IN1(n57), .IN2(n3564), .Q(n6531) );
  INVX0 U7717 ( .INP(n6537), .ZN(n57) );
  OR2X1 U7718 ( .IN1(n4427), .IN2(n4009), .Q(n6537) );
  OR4X1 U7719 ( .IN1(n6538), .IN2(n6539), .IN3(n6540), .IN4(n6541), .Q(WX1985)
         );
  AND2X1 U7720 ( .IN1(n3632), .IN2(n6286), .Q(n6541) );
  XNOR3X1 U7721 ( .IN1(n3384), .IN2(n3151), .IN3(n6542), .Q(n6286) );
  XOR2X1 U7722 ( .IN1(WX3343), .IN2(n7219), .Q(n6542) );
  AND2X1 U7723 ( .IN1(n3548), .IN2(n5500), .Q(n6540) );
  XNOR3X1 U7724 ( .IN1(n3409), .IN2(n3165), .IN3(n6543), .Q(n5500) );
  XOR2X1 U7725 ( .IN1(WX2050), .IN2(n7218), .Q(n6543) );
  AND2X1 U7726 ( .IN1(test_so20), .IN2(n3587), .Q(n6539) );
  AND2X1 U7727 ( .IN1(n56), .IN2(n3564), .Q(n6538) );
  INVX0 U7728 ( .INP(n6544), .ZN(n56) );
  OR2X1 U7729 ( .IN1(n4427), .IN2(n4010), .Q(n6544) );
  OR4X1 U7730 ( .IN1(n6545), .IN2(n6546), .IN3(n6547), .IN4(n6548), .Q(WX1983)
         );
  AND2X1 U7731 ( .IN1(n6293), .IN2(n3623), .Q(n6548) );
  XOR3X1 U7732 ( .IN1(n3739), .IN2(n3383), .IN3(n6549), .Q(n6293) );
  XOR2X1 U7733 ( .IN1(WX3277), .IN2(test_so28), .Q(n6549) );
  AND2X1 U7734 ( .IN1(n3548), .IN2(n5506), .Q(n6547) );
  XNOR3X1 U7735 ( .IN1(n3408), .IN2(n3166), .IN3(n6550), .Q(n5506) );
  XOR2X1 U7736 ( .IN1(WX2048), .IN2(n7220), .Q(n6550) );
  AND2X1 U7737 ( .IN1(n3595), .IN2(CRC_OUT_8_8), .Q(n6546) );
  AND2X1 U7738 ( .IN1(n55), .IN2(n3564), .Q(n6545) );
  INVX0 U7739 ( .INP(n6551), .ZN(n55) );
  OR2X1 U7740 ( .IN1(n4427), .IN2(n4011), .Q(n6551) );
  OR4X1 U7741 ( .IN1(n6552), .IN2(n6553), .IN3(n6554), .IN4(n6555), .Q(WX1981)
         );
  AND2X1 U7742 ( .IN1(n3632), .IN2(n6300), .Q(n6555) );
  XNOR3X1 U7743 ( .IN1(n3382), .IN2(n3152), .IN3(n6556), .Q(n6300) );
  XOR2X1 U7744 ( .IN1(WX3339), .IN2(n7222), .Q(n6556) );
  AND2X1 U7745 ( .IN1(n3546), .IN2(n5512), .Q(n6554) );
  XNOR3X1 U7746 ( .IN1(n3407), .IN2(n3167), .IN3(n6557), .Q(n5512) );
  XOR2X1 U7747 ( .IN1(WX2046), .IN2(n7221), .Q(n6557) );
  AND2X1 U7748 ( .IN1(n3595), .IN2(CRC_OUT_8_9), .Q(n6553) );
  AND2X1 U7749 ( .IN1(n54), .IN2(n3564), .Q(n6552) );
  INVX0 U7750 ( .INP(n6558), .ZN(n54) );
  OR2X1 U7751 ( .IN1(n4427), .IN2(n4012), .Q(n6558) );
  OR4X1 U7752 ( .IN1(n6559), .IN2(n6560), .IN3(n6561), .IN4(n6562), .Q(WX1979)
         );
  AND2X1 U7753 ( .IN1(n3632), .IN2(n6307), .Q(n6562) );
  XNOR3X1 U7754 ( .IN1(n3381), .IN2(n3153), .IN3(n6563), .Q(n6307) );
  XOR2X1 U7755 ( .IN1(WX3337), .IN2(n7223), .Q(n6563) );
  AND2X1 U7756 ( .IN1(n5518), .IN2(n3532), .Q(n6561) );
  XOR3X1 U7757 ( .IN1(n3775), .IN2(n3168), .IN3(n6564), .Q(n5518) );
  XOR2X1 U7758 ( .IN1(WX1980), .IN2(test_so19), .Q(n6564) );
  AND2X1 U7759 ( .IN1(n3595), .IN2(CRC_OUT_8_10), .Q(n6560) );
  AND2X1 U7760 ( .IN1(n53), .IN2(n3564), .Q(n6559) );
  INVX0 U7761 ( .INP(n6565), .ZN(n53) );
  OR2X1 U7762 ( .IN1(n4427), .IN2(n4013), .Q(n6565) );
  OR4X1 U7763 ( .IN1(n6566), .IN2(n6567), .IN3(n6568), .IN4(n6569), .Q(WX1977)
         );
  AND2X1 U7764 ( .IN1(n3632), .IN2(n6314), .Q(n6569) );
  XNOR3X1 U7765 ( .IN1(n3189), .IN2(n3154), .IN3(n6570), .Q(n6314) );
  XOR2X1 U7766 ( .IN1(WX3335), .IN2(n7225), .Q(n6570) );
  AND2X1 U7767 ( .IN1(n3546), .IN2(n5524), .Q(n6568) );
  XNOR3X1 U7768 ( .IN1(n3192), .IN2(n3169), .IN3(n6571), .Q(n5524) );
  XOR2X1 U7769 ( .IN1(WX2042), .IN2(n7224), .Q(n6571) );
  AND2X1 U7770 ( .IN1(n3595), .IN2(CRC_OUT_8_11), .Q(n6567) );
  AND2X1 U7771 ( .IN1(n52), .IN2(n3564), .Q(n6566) );
  INVX0 U7772 ( .INP(n6572), .ZN(n52) );
  OR2X1 U7773 ( .IN1(n4427), .IN2(n4014), .Q(n6572) );
  OR4X1 U7774 ( .IN1(n6573), .IN2(n6574), .IN3(n6575), .IN4(n6576), .Q(WX1975)
         );
  AND2X1 U7775 ( .IN1(n6321), .IN2(n3623), .Q(n6576) );
  XOR3X1 U7776 ( .IN1(n3380), .IN2(n3155), .IN3(n6577), .Q(n6321) );
  XOR2X1 U7777 ( .IN1(WX3269), .IN2(test_so26), .Q(n6577) );
  AND2X1 U7778 ( .IN1(n3546), .IN2(n5530), .Q(n6575) );
  XNOR3X1 U7779 ( .IN1(n3406), .IN2(n3170), .IN3(n6578), .Q(n5530) );
  XOR2X1 U7780 ( .IN1(WX2040), .IN2(n7226), .Q(n6578) );
  AND2X1 U7781 ( .IN1(n3595), .IN2(CRC_OUT_8_12), .Q(n6574) );
  AND2X1 U7782 ( .IN1(n51), .IN2(n3564), .Q(n6573) );
  INVX0 U7783 ( .INP(n6579), .ZN(n51) );
  OR2X1 U7784 ( .IN1(n4427), .IN2(n4015), .Q(n6579) );
  OR4X1 U7785 ( .IN1(n6580), .IN2(n6581), .IN3(n6582), .IN4(n6583), .Q(WX1973)
         );
  AND2X1 U7786 ( .IN1(n3633), .IN2(n6328), .Q(n6583) );
  XNOR3X1 U7787 ( .IN1(n3379), .IN2(n3156), .IN3(n6584), .Q(n6328) );
  XOR2X1 U7788 ( .IN1(WX3331), .IN2(n7228), .Q(n6584) );
  AND2X1 U7789 ( .IN1(n3546), .IN2(n5536), .Q(n6582) );
  XNOR3X1 U7790 ( .IN1(n3405), .IN2(n3171), .IN3(n6585), .Q(n5536) );
  XOR2X1 U7791 ( .IN1(WX2038), .IN2(n7227), .Q(n6585) );
  AND2X1 U7792 ( .IN1(n3595), .IN2(CRC_OUT_8_13), .Q(n6581) );
  AND2X1 U7793 ( .IN1(n50), .IN2(n3564), .Q(n6580) );
  INVX0 U7794 ( .INP(n6586), .ZN(n50) );
  OR2X1 U7795 ( .IN1(n4426), .IN2(n4016), .Q(n6586) );
  OR4X1 U7796 ( .IN1(n6587), .IN2(n6588), .IN3(n6589), .IN4(n6590), .Q(WX1971)
         );
  AND2X1 U7797 ( .IN1(n3633), .IN2(n6335), .Q(n6590) );
  XNOR3X1 U7798 ( .IN1(n3378), .IN2(n3157), .IN3(n6591), .Q(n6335) );
  XOR2X1 U7799 ( .IN1(WX3329), .IN2(n7229), .Q(n6591) );
  AND2X1 U7800 ( .IN1(n5542), .IN2(n3531), .Q(n6589) );
  XOR3X1 U7801 ( .IN1(n3783), .IN2(n3404), .IN3(n6592), .Q(n5542) );
  XOR2X1 U7802 ( .IN1(WX1972), .IN2(test_so17), .Q(n6592) );
  AND2X1 U7803 ( .IN1(n3595), .IN2(CRC_OUT_8_14), .Q(n6588) );
  AND2X1 U7804 ( .IN1(n49), .IN2(n3563), .Q(n6587) );
  INVX0 U7805 ( .INP(n6593), .ZN(n49) );
  OR2X1 U7806 ( .IN1(n4426), .IN2(n4017), .Q(n6593) );
  OR4X1 U7807 ( .IN1(n6594), .IN2(n6595), .IN3(n6596), .IN4(n6597), .Q(WX1969)
         );
  AND2X1 U7808 ( .IN1(n3633), .IN2(n6342), .Q(n6597) );
  XNOR3X1 U7809 ( .IN1(n3377), .IN2(n3158), .IN3(n6598), .Q(n6342) );
  XOR2X1 U7810 ( .IN1(WX3327), .IN2(n7231), .Q(n6598) );
  AND2X1 U7811 ( .IN1(n3546), .IN2(n5548), .Q(n6596) );
  XNOR3X1 U7812 ( .IN1(n3403), .IN2(n3172), .IN3(n6599), .Q(n5548) );
  XOR2X1 U7813 ( .IN1(WX2034), .IN2(n7230), .Q(n6599) );
  AND2X1 U7814 ( .IN1(n3596), .IN2(CRC_OUT_8_15), .Q(n6595) );
  AND2X1 U7815 ( .IN1(n48), .IN2(n3563), .Q(n6594) );
  INVX0 U7816 ( .INP(n6600), .ZN(n48) );
  OR2X1 U7817 ( .IN1(n4426), .IN2(n4018), .Q(n6600) );
  OR4X1 U7818 ( .IN1(n6601), .IN2(n6602), .IN3(n6603), .IN4(n6604), .Q(WX1967)
         );
  AND2X1 U7819 ( .IN1(n6349), .IN2(n3623), .Q(n6604) );
  XOR3X1 U7820 ( .IN1(n3006), .IN2(TM1), .IN3(n6605), .Q(n6349) );
  XNOR3X1 U7821 ( .IN1(test_so24), .IN2(n7232), .IN3(n3188), .Q(n6605) );
  AND2X1 U7822 ( .IN1(n3546), .IN2(n5554), .Q(n6603) );
  XOR3X1 U7823 ( .IN1(n3032), .IN2(n3514), .IN3(n6606), .Q(n5554) );
  XNOR3X1 U7824 ( .IN1(n8653), .IN2(n3191), .IN3(WX2096), .Q(n6606) );
  AND2X1 U7825 ( .IN1(n3596), .IN2(CRC_OUT_8_16), .Q(n6602) );
  AND2X1 U7826 ( .IN1(n47), .IN2(n3563), .Q(n6601) );
  INVX0 U7827 ( .INP(n6607), .ZN(n47) );
  OR2X1 U7828 ( .IN1(n4426), .IN2(n4019), .Q(n6607) );
  OR4X1 U7829 ( .IN1(n6608), .IN2(n6609), .IN3(n6610), .IN4(n6611), .Q(WX1965)
         );
  AND2X1 U7830 ( .IN1(n3633), .IN2(n6356), .Q(n6611) );
  XOR3X1 U7831 ( .IN1(n3007), .IN2(n3518), .IN3(n6612), .Q(n6356) );
  XOR3X1 U7832 ( .IN1(n7233), .IN2(n3376), .IN3(WX3387), .Q(n6612) );
  AND2X1 U7833 ( .IN1(n3546), .IN2(n5560), .Q(n6610) );
  XOR3X1 U7834 ( .IN1(n3034), .IN2(n3516), .IN3(n6613), .Q(n5560) );
  XNOR3X1 U7835 ( .IN1(n8654), .IN2(n3402), .IN3(WX2094), .Q(n6613) );
  AND2X1 U7836 ( .IN1(n3596), .IN2(CRC_OUT_8_17), .Q(n6609) );
  AND2X1 U7837 ( .IN1(n46), .IN2(n3563), .Q(n6608) );
  INVX0 U7838 ( .INP(n6614), .ZN(n46) );
  OR2X1 U7839 ( .IN1(n4426), .IN2(n4020), .Q(n6614) );
  OR4X1 U7840 ( .IN1(n6615), .IN2(n6616), .IN3(n6617), .IN4(n6618), .Q(WX1963)
         );
  AND2X1 U7841 ( .IN1(n3633), .IN2(n6363), .Q(n6618) );
  XOR3X1 U7842 ( .IN1(n3009), .IN2(n3515), .IN3(n6619), .Q(n6363) );
  XOR3X1 U7843 ( .IN1(n7235), .IN2(n3375), .IN3(WX3385), .Q(n6619) );
  AND2X1 U7844 ( .IN1(n5566), .IN2(n3532), .Q(n6617) );
  XOR3X1 U7845 ( .IN1(n3036), .IN2(TM1), .IN3(n6620), .Q(n5566) );
  XNOR3X1 U7846 ( .IN1(test_so15), .IN2(n7234), .IN3(n3401), .Q(n6620) );
  AND2X1 U7847 ( .IN1(n3596), .IN2(CRC_OUT_8_18), .Q(n6616) );
  AND2X1 U7848 ( .IN1(n45), .IN2(n3563), .Q(n6615) );
  INVX0 U7849 ( .INP(n6621), .ZN(n45) );
  OR2X1 U7850 ( .IN1(n4426), .IN2(n4021), .Q(n6621) );
  OR4X1 U7851 ( .IN1(n6622), .IN2(n6623), .IN3(n6624), .IN4(n6625), .Q(WX1961)
         );
  AND2X1 U7852 ( .IN1(n3633), .IN2(n6370), .Q(n6625) );
  XOR3X1 U7853 ( .IN1(n3011), .IN2(n3514), .IN3(n6626), .Q(n6370) );
  XOR3X1 U7854 ( .IN1(n7236), .IN2(n3374), .IN3(WX3383), .Q(n6626) );
  AND2X1 U7855 ( .IN1(n3546), .IN2(n5572), .Q(n6624) );
  XOR3X1 U7856 ( .IN1(n3037), .IN2(n3518), .IN3(n6627), .Q(n5572) );
  XNOR3X1 U7857 ( .IN1(n8656), .IN2(n3400), .IN3(WX2090), .Q(n6627) );
  AND2X1 U7858 ( .IN1(n3596), .IN2(CRC_OUT_8_19), .Q(n6623) );
  AND2X1 U7859 ( .IN1(n44), .IN2(n3563), .Q(n6622) );
  INVX0 U7860 ( .INP(n6628), .ZN(n44) );
  OR2X1 U7861 ( .IN1(n4426), .IN2(n4022), .Q(n6628) );
  OR4X1 U7862 ( .IN1(n6629), .IN2(n6630), .IN3(n6631), .IN4(n6632), .Q(WX1959)
         );
  AND2X1 U7863 ( .IN1(n3633), .IN2(n6377), .Q(n6632) );
  XOR3X1 U7864 ( .IN1(n3013), .IN2(n3516), .IN3(n6633), .Q(n6377) );
  XOR3X1 U7865 ( .IN1(n7237), .IN2(n3373), .IN3(WX3381), .Q(n6633) );
  AND2X1 U7866 ( .IN1(n3546), .IN2(n5578), .Q(n6631) );
  XOR3X1 U7867 ( .IN1(n3039), .IN2(n3515), .IN3(n6634), .Q(n5578) );
  XNOR3X1 U7868 ( .IN1(n8657), .IN2(n3399), .IN3(WX2088), .Q(n6634) );
  AND2X1 U7869 ( .IN1(n3596), .IN2(CRC_OUT_8_20), .Q(n6630) );
  AND2X1 U7870 ( .IN1(n43), .IN2(n3563), .Q(n6629) );
  INVX0 U7871 ( .INP(n6635), .ZN(n43) );
  OR2X1 U7872 ( .IN1(n4426), .IN2(n4023), .Q(n6635) );
  OR4X1 U7873 ( .IN1(n6636), .IN2(n6637), .IN3(n6638), .IN4(n6639), .Q(WX1957)
         );
  AND2X1 U7874 ( .IN1(n3633), .IN2(n6384), .Q(n6639) );
  XOR3X1 U7875 ( .IN1(n3015), .IN2(n3514), .IN3(n6640), .Q(n6384) );
  XOR3X1 U7876 ( .IN1(n7238), .IN2(n3372), .IN3(WX3379), .Q(n6640) );
  AND2X1 U7877 ( .IN1(n3546), .IN2(n5584), .Q(n6638) );
  XOR3X1 U7878 ( .IN1(n3041), .IN2(n3518), .IN3(n6641), .Q(n5584) );
  XNOR3X1 U7879 ( .IN1(n8658), .IN2(n3398), .IN3(WX2086), .Q(n6641) );
  AND2X1 U7880 ( .IN1(n3596), .IN2(CRC_OUT_8_21), .Q(n6637) );
  AND2X1 U7881 ( .IN1(n42), .IN2(n3563), .Q(n6636) );
  INVX0 U7882 ( .INP(n6642), .ZN(n42) );
  OR2X1 U7883 ( .IN1(n4426), .IN2(n4024), .Q(n6642) );
  OR4X1 U7884 ( .IN1(n6643), .IN2(n6644), .IN3(n6645), .IN4(n6646), .Q(WX1955)
         );
  AND2X1 U7885 ( .IN1(n3633), .IN2(n6391), .Q(n6646) );
  XOR3X1 U7886 ( .IN1(n3017), .IN2(n3516), .IN3(n6647), .Q(n6391) );
  XOR3X1 U7887 ( .IN1(n7240), .IN2(n3371), .IN3(WX3377), .Q(n6647) );
  AND2X1 U7888 ( .IN1(n5590), .IN2(n3531), .Q(n6645) );
  XOR3X1 U7889 ( .IN1(n3043), .IN2(TM1), .IN3(n6648), .Q(n5590) );
  XNOR3X1 U7890 ( .IN1(test_so13), .IN2(n7239), .IN3(n3397), .Q(n6648) );
  AND2X1 U7891 ( .IN1(n3596), .IN2(CRC_OUT_8_22), .Q(n6644) );
  AND2X1 U7892 ( .IN1(n41), .IN2(n3563), .Q(n6643) );
  INVX0 U7893 ( .INP(n6649), .ZN(n41) );
  OR2X1 U7894 ( .IN1(n4426), .IN2(n4025), .Q(n6649) );
  OR4X1 U7895 ( .IN1(n6650), .IN2(n6651), .IN3(n6652), .IN4(n6653), .Q(WX1953)
         );
  AND2X1 U7896 ( .IN1(n6398), .IN2(n3623), .Q(n6653) );
  XOR3X1 U7897 ( .IN1(n3019), .IN2(TM1), .IN3(n6654), .Q(n6398) );
  XOR3X1 U7898 ( .IN1(test_so29), .IN2(n7241), .IN3(WX3375), .Q(n6654) );
  AND2X1 U7899 ( .IN1(n3546), .IN2(n5596), .Q(n6652) );
  XOR3X1 U7900 ( .IN1(n3044), .IN2(n3515), .IN3(n6655), .Q(n5596) );
  XNOR3X1 U7901 ( .IN1(n8661), .IN2(n3396), .IN3(WX2082), .Q(n6655) );
  AND2X1 U7902 ( .IN1(n3596), .IN2(CRC_OUT_8_23), .Q(n6651) );
  AND2X1 U7903 ( .IN1(n40), .IN2(n3563), .Q(n6650) );
  INVX0 U7904 ( .INP(n6656), .ZN(n40) );
  OR2X1 U7905 ( .IN1(n4426), .IN2(n4026), .Q(n6656) );
  OR4X1 U7906 ( .IN1(n6657), .IN2(n6658), .IN3(n6659), .IN4(n6660), .Q(WX1951)
         );
  AND2X1 U7907 ( .IN1(n3633), .IN2(n6405), .Q(n6660) );
  XOR3X1 U7908 ( .IN1(n3020), .IN2(n3514), .IN3(n6661), .Q(n6405) );
  XOR3X1 U7909 ( .IN1(n7242), .IN2(n3370), .IN3(WX3373), .Q(n6661) );
  AND2X1 U7910 ( .IN1(n3546), .IN2(n5602), .Q(n6659) );
  XOR3X1 U7911 ( .IN1(n3046), .IN2(n3518), .IN3(n6662), .Q(n5602) );
  XNOR3X1 U7912 ( .IN1(n8662), .IN2(n3395), .IN3(WX2080), .Q(n6662) );
  AND2X1 U7913 ( .IN1(n3596), .IN2(CRC_OUT_8_24), .Q(n6658) );
  AND2X1 U7914 ( .IN1(n39), .IN2(n3563), .Q(n6657) );
  INVX0 U7915 ( .INP(n6663), .ZN(n39) );
  OR2X1 U7916 ( .IN1(n4426), .IN2(n4027), .Q(n6663) );
  OR4X1 U7917 ( .IN1(n6664), .IN2(n6665), .IN3(n6666), .IN4(n6667), .Q(WX1949)
         );
  AND2X1 U7918 ( .IN1(n3633), .IN2(n6412), .Q(n6667) );
  XOR3X1 U7919 ( .IN1(n3022), .IN2(n3516), .IN3(n6668), .Q(n6412) );
  XOR3X1 U7920 ( .IN1(n7243), .IN2(n3369), .IN3(WX3371), .Q(n6668) );
  AND2X1 U7921 ( .IN1(n3546), .IN2(n5608), .Q(n6666) );
  XOR3X1 U7922 ( .IN1(n3048), .IN2(n3515), .IN3(n6669), .Q(n5608) );
  XNOR3X1 U7923 ( .IN1(n8663), .IN2(n3394), .IN3(WX2078), .Q(n6669) );
  AND2X1 U7924 ( .IN1(test_so21), .IN2(n3588), .Q(n6665) );
  AND2X1 U7925 ( .IN1(n38), .IN2(n3563), .Q(n6664) );
  INVX0 U7926 ( .INP(n6670), .ZN(n38) );
  OR2X1 U7927 ( .IN1(n4426), .IN2(n4028), .Q(n6670) );
  OR4X1 U7928 ( .IN1(n6671), .IN2(n6672), .IN3(n6673), .IN4(n6674), .Q(WX1947)
         );
  AND2X1 U7929 ( .IN1(n6419), .IN2(n3623), .Q(n6674) );
  XOR3X1 U7930 ( .IN1(n3024), .IN2(TM1), .IN3(n6675), .Q(n6419) );
  XNOR3X1 U7931 ( .IN1(test_so27), .IN2(n7244), .IN3(n3368), .Q(n6675) );
  AND2X1 U7932 ( .IN1(n3545), .IN2(n5614), .Q(n6673) );
  XOR3X1 U7933 ( .IN1(n3050), .IN2(n3514), .IN3(n6676), .Q(n5614) );
  XNOR3X1 U7934 ( .IN1(n8664), .IN2(n3393), .IN3(WX2076), .Q(n6676) );
  AND2X1 U7935 ( .IN1(n3596), .IN2(CRC_OUT_8_26), .Q(n6672) );
  AND2X1 U7936 ( .IN1(n37), .IN2(n3562), .Q(n6671) );
  INVX0 U7937 ( .INP(n6677), .ZN(n37) );
  OR2X1 U7938 ( .IN1(n4425), .IN2(n4029), .Q(n6677) );
  OR4X1 U7939 ( .IN1(n6678), .IN2(n6679), .IN3(n6680), .IN4(n6681), .Q(WX1945)
         );
  AND2X1 U7940 ( .IN1(n3629), .IN2(n6426), .Q(n6681) );
  XOR3X1 U7941 ( .IN1(n3025), .IN2(n3518), .IN3(n6682), .Q(n6426) );
  XOR3X1 U7942 ( .IN1(n7245), .IN2(n3367), .IN3(WX3367), .Q(n6682) );
  AND2X1 U7943 ( .IN1(n3545), .IN2(n5620), .Q(n6680) );
  XOR3X1 U7944 ( .IN1(n3052), .IN2(n3516), .IN3(n6683), .Q(n5620) );
  XNOR3X1 U7945 ( .IN1(n8665), .IN2(n3392), .IN3(WX2074), .Q(n6683) );
  AND2X1 U7946 ( .IN1(n3596), .IN2(CRC_OUT_8_27), .Q(n6679) );
  AND2X1 U7947 ( .IN1(n36), .IN2(n3562), .Q(n6678) );
  INVX0 U7948 ( .INP(n6684), .ZN(n36) );
  OR2X1 U7949 ( .IN1(n4425), .IN2(n4030), .Q(n6684) );
  OR4X1 U7950 ( .IN1(n6685), .IN2(n6686), .IN3(n6687), .IN4(n6688), .Q(WX1943)
         );
  AND2X1 U7951 ( .IN1(n3634), .IN2(n6433), .Q(n6688) );
  XOR3X1 U7952 ( .IN1(n3027), .IN2(n3515), .IN3(n6689), .Q(n6433) );
  XOR3X1 U7953 ( .IN1(n7246), .IN2(n3366), .IN3(WX3365), .Q(n6689) );
  AND2X1 U7954 ( .IN1(n5626), .IN2(n3531), .Q(n6687) );
  XOR3X1 U7955 ( .IN1(n3054), .IN2(TM1), .IN3(n6690), .Q(n5626) );
  XNOR3X1 U7956 ( .IN1(test_so18), .IN2(n8666), .IN3(WX2072), .Q(n6690) );
  AND2X1 U7957 ( .IN1(n3596), .IN2(CRC_OUT_8_28), .Q(n6686) );
  AND2X1 U7958 ( .IN1(n35), .IN2(n3562), .Q(n6685) );
  INVX0 U7959 ( .INP(n6691), .ZN(n35) );
  OR2X1 U7960 ( .IN1(n4425), .IN2(n4031), .Q(n6691) );
  OR4X1 U7961 ( .IN1(n6692), .IN2(n6693), .IN3(n6694), .IN4(n6695), .Q(WX1941)
         );
  AND2X1 U7962 ( .IN1(n3633), .IN2(n6440), .Q(n6695) );
  XOR3X1 U7963 ( .IN1(n3029), .IN2(n3514), .IN3(n6696), .Q(n6440) );
  XOR3X1 U7964 ( .IN1(n7247), .IN2(n3365), .IN3(WX3363), .Q(n6696) );
  AND2X1 U7965 ( .IN1(n3545), .IN2(n5643), .Q(n6694) );
  XOR3X1 U7966 ( .IN1(n3055), .IN2(n3518), .IN3(n6697), .Q(n5643) );
  XNOR3X1 U7967 ( .IN1(n8667), .IN2(n3391), .IN3(WX2070), .Q(n6697) );
  AND2X1 U7968 ( .IN1(n3597), .IN2(CRC_OUT_8_29), .Q(n6693) );
  AND2X1 U7969 ( .IN1(n34), .IN2(n3562), .Q(n6692) );
  INVX0 U7970 ( .INP(n6698), .ZN(n34) );
  OR2X1 U7971 ( .IN1(n4425), .IN2(n4032), .Q(n6698) );
  OR4X1 U7972 ( .IN1(n6699), .IN2(n6700), .IN3(n6701), .IN4(n6702), .Q(WX1939)
         );
  AND2X1 U7973 ( .IN1(n6447), .IN2(n3624), .Q(n6702) );
  XOR3X1 U7974 ( .IN1(n3031), .IN2(TM1), .IN3(n6703), .Q(n6447) );
  XNOR3X1 U7975 ( .IN1(test_so25), .IN2(n7248), .IN3(n3364), .Q(n6703) );
  AND2X1 U7976 ( .IN1(n3545), .IN2(n5659), .Q(n6701) );
  XOR3X1 U7977 ( .IN1(n3057), .IN2(n3516), .IN3(n6704), .Q(n5659) );
  XNOR3X1 U7978 ( .IN1(n8668), .IN2(n3390), .IN3(WX2068), .Q(n6704) );
  AND2X1 U7979 ( .IN1(n3597), .IN2(CRC_OUT_8_30), .Q(n6700) );
  AND2X1 U7980 ( .IN1(n33), .IN2(n3562), .Q(n6699) );
  INVX0 U7981 ( .INP(n6705), .ZN(n33) );
  OR2X1 U7982 ( .IN1(n4425), .IN2(n4033), .Q(n6705) );
  OR4X1 U7983 ( .IN1(n6706), .IN2(n6707), .IN3(n6708), .IN4(n6709), .Q(WX1937)
         );
  AND2X1 U7984 ( .IN1(n3545), .IN2(n5675), .Q(n6709) );
  XOR3X1 U7985 ( .IN1(n2845), .IN2(n3515), .IN3(n6710), .Q(n5675) );
  XNOR3X1 U7986 ( .IN1(n8669), .IN2(n3389), .IN3(WX2066), .Q(n6710) );
  AND2X1 U7987 ( .IN1(n3633), .IN2(n6454), .Q(n6708) );
  XOR3X1 U7988 ( .IN1(n2843), .IN2(n3514), .IN3(n6711), .Q(n6454) );
  XOR3X1 U7989 ( .IN1(n7249), .IN2(n3363), .IN3(WX3359), .Q(n6711) );
  AND2X1 U7990 ( .IN1(n2245), .IN2(WX1778), .Q(n6707) );
  AND2X1 U7991 ( .IN1(n3597), .IN2(CRC_OUT_8_31), .Q(n6706) );
  AND2X1 U7992 ( .IN1(n3496), .IN2(n4383), .Q(WX1839) );
  AND2X1 U7993 ( .IN1(n6712), .IN2(n4375), .Q(WX1326) );
  XOR2X1 U7994 ( .IN1(CRC_OUT_9_30), .IN2(n3468), .Q(n6712) );
  AND2X1 U7995 ( .IN1(n6713), .IN2(n4375), .Q(WX1324) );
  XOR2X1 U7996 ( .IN1(CRC_OUT_9_29), .IN2(n3417), .Q(n6713) );
  AND2X1 U7997 ( .IN1(n6714), .IN2(n4375), .Q(WX1322) );
  XOR2X1 U7998 ( .IN1(CRC_OUT_9_28), .IN2(n3422), .Q(n6714) );
  AND2X1 U7999 ( .IN1(n6715), .IN2(n4375), .Q(WX1320) );
  XOR2X1 U8000 ( .IN1(CRC_OUT_9_27), .IN2(n3428), .Q(n6715) );
  AND2X1 U8001 ( .IN1(n6716), .IN2(n4375), .Q(WX1318) );
  XOR2X1 U8002 ( .IN1(CRC_OUT_9_26), .IN2(n3431), .Q(n6716) );
  AND2X1 U8003 ( .IN1(n6717), .IN2(n4375), .Q(WX1316) );
  XOR2X1 U8004 ( .IN1(CRC_OUT_9_25), .IN2(n3433), .Q(n6717) );
  AND2X1 U8005 ( .IN1(n6718), .IN2(n4374), .Q(WX1314) );
  XOR2X1 U8006 ( .IN1(CRC_OUT_9_24), .IN2(n3438), .Q(n6718) );
  AND2X1 U8007 ( .IN1(n6719), .IN2(n4374), .Q(WX1312) );
  XOR2X1 U8008 ( .IN1(CRC_OUT_9_23), .IN2(n3444), .Q(n6719) );
  AND2X1 U8009 ( .IN1(n6720), .IN2(n4374), .Q(WX1310) );
  XOR2X1 U8010 ( .IN1(CRC_OUT_9_22), .IN2(n3445), .Q(n6720) );
  AND2X1 U8011 ( .IN1(n6721), .IN2(n4374), .Q(WX1308) );
  XOR2X1 U8012 ( .IN1(CRC_OUT_9_21), .IN2(n3456), .Q(n6721) );
  AND2X1 U8013 ( .IN1(n6722), .IN2(n4374), .Q(WX1306) );
  XOR2X1 U8014 ( .IN1(CRC_OUT_9_20), .IN2(n3462), .Q(n6722) );
  AND2X1 U8015 ( .IN1(n6723), .IN2(n4374), .Q(WX1304) );
  XOR2X1 U8016 ( .IN1(test_so10), .IN2(n3465), .Q(n6723) );
  AND2X1 U8017 ( .IN1(n6724), .IN2(n4374), .Q(WX1302) );
  XOR2X1 U8018 ( .IN1(CRC_OUT_9_18), .IN2(n3420), .Q(n6724) );
  AND2X1 U8019 ( .IN1(n6725), .IN2(n4374), .Q(WX1300) );
  XOR2X1 U8020 ( .IN1(CRC_OUT_9_17), .IN2(n3429), .Q(n6725) );
  AND2X1 U8021 ( .IN1(n6726), .IN2(n4374), .Q(WX1298) );
  XOR2X1 U8022 ( .IN1(CRC_OUT_9_16), .IN2(n3436), .Q(n6726) );
  AND2X1 U8023 ( .IN1(n6727), .IN2(n4373), .Q(WX1296) );
  XOR3X1 U8024 ( .IN1(test_so8), .IN2(DFF_191_n1), .IN3(CRC_OUT_9_15), .Q(
        n6727) );
  AND2X1 U8025 ( .IN1(n6728), .IN2(n4373), .Q(WX1294) );
  XOR2X1 U8026 ( .IN1(CRC_OUT_9_14), .IN2(n3459), .Q(n6728) );
  AND2X1 U8027 ( .IN1(n6729), .IN2(n4373), .Q(WX1292) );
  XOR2X1 U8028 ( .IN1(CRC_OUT_9_13), .IN2(n3470), .Q(n6729) );
  AND2X1 U8029 ( .IN1(n6730), .IN2(n4373), .Q(WX1290) );
  XOR2X1 U8030 ( .IN1(CRC_OUT_9_12), .IN2(n3424), .Q(n6730) );
  AND2X1 U8031 ( .IN1(n6731), .IN2(n4373), .Q(WX1288) );
  XOR2X1 U8032 ( .IN1(CRC_OUT_9_11), .IN2(n3440), .Q(n6731) );
  AND2X1 U8033 ( .IN1(n6732), .IN2(n4373), .Q(WX1286) );
  XOR3X1 U8034 ( .IN1(n3484), .IN2(DFF_191_n1), .IN3(DFF_170_n1), .Q(n6732) );
  AND2X1 U8035 ( .IN1(n6733), .IN2(n4373), .Q(WX1284) );
  XOR2X1 U8036 ( .IN1(CRC_OUT_9_9), .IN2(n3435), .Q(n6733) );
  AND2X1 U8037 ( .IN1(n6734), .IN2(n4373), .Q(WX1282) );
  XOR2X1 U8038 ( .IN1(CRC_OUT_9_8), .IN2(n3443), .Q(n6734) );
  AND2X1 U8039 ( .IN1(n6735), .IN2(n4373), .Q(WX1280) );
  XOR2X1 U8040 ( .IN1(CRC_OUT_9_7), .IN2(n3448), .Q(n6735) );
  AND2X1 U8041 ( .IN1(n6736), .IN2(n4372), .Q(WX1278) );
  XOR2X1 U8042 ( .IN1(CRC_OUT_9_6), .IN2(n3482), .Q(n6736) );
  AND2X1 U8043 ( .IN1(n6737), .IN2(n4372), .Q(WX1276) );
  XOR2X1 U8044 ( .IN1(CRC_OUT_9_5), .IN2(n3464), .Q(n6737) );
  AND2X1 U8045 ( .IN1(n6738), .IN2(n4372), .Q(WX1274) );
  XOR2X1 U8046 ( .IN1(CRC_OUT_9_4), .IN2(n3450), .Q(n6738) );
  AND2X1 U8047 ( .IN1(n6739), .IN2(n4372), .Q(WX1272) );
  XOR3X1 U8048 ( .IN1(n3452), .IN2(DFF_191_n1), .IN3(DFF_163_n1), .Q(n6739) );
  AND2X1 U8049 ( .IN1(n6740), .IN2(n4372), .Q(WX1270) );
  XOR2X1 U8050 ( .IN1(CRC_OUT_9_2), .IN2(n3418), .Q(n6740) );
  AND2X1 U8051 ( .IN1(n6741), .IN2(n4372), .Q(WX1268) );
  XOR2X1 U8052 ( .IN1(test_so9), .IN2(n3476), .Q(n6741) );
  AND2X1 U8053 ( .IN1(n6742), .IN2(n4372), .Q(WX1266) );
  XOR2X1 U8054 ( .IN1(CRC_OUT_9_0), .IN2(n3426), .Q(n6742) );
  AND2X1 U8055 ( .IN1(n6743), .IN2(n4372), .Q(WX1264) );
  XOR2X1 U8056 ( .IN1(n3490), .IN2(CRC_OUT_9_31), .Q(n6743) );
  AND2X1 U8057 ( .IN1(n6744), .IN2(n4372), .Q(WX11670) );
  XOR2X1 U8058 ( .IN1(CRC_OUT_1_30), .IN2(n3202), .Q(n6744) );
  AND2X1 U8059 ( .IN1(n6745), .IN2(n4371), .Q(WX11668) );
  XOR2X1 U8060 ( .IN1(CRC_OUT_1_29), .IN2(n3203), .Q(n6745) );
  AND2X1 U8061 ( .IN1(n6746), .IN2(n4371), .Q(WX11666) );
  XOR2X1 U8062 ( .IN1(CRC_OUT_1_28), .IN2(n3204), .Q(n6746) );
  AND2X1 U8063 ( .IN1(n6747), .IN2(n4371), .Q(WX11664) );
  XOR2X1 U8064 ( .IN1(CRC_OUT_1_27), .IN2(n3205), .Q(n6747) );
  AND2X1 U8065 ( .IN1(n6748), .IN2(n4371), .Q(WX11662) );
  XOR2X1 U8066 ( .IN1(CRC_OUT_1_26), .IN2(n3206), .Q(n6748) );
  AND2X1 U8067 ( .IN1(n6749), .IN2(n4371), .Q(WX11660) );
  XOR2X1 U8068 ( .IN1(CRC_OUT_1_25), .IN2(n3207), .Q(n6749) );
  AND2X1 U8069 ( .IN1(n6750), .IN2(n4371), .Q(WX11658) );
  XOR2X1 U8070 ( .IN1(CRC_OUT_1_24), .IN2(n3208), .Q(n6750) );
  AND2X1 U8071 ( .IN1(n6751), .IN2(n4371), .Q(WX11656) );
  XOR2X1 U8072 ( .IN1(CRC_OUT_1_23), .IN2(n3209), .Q(n6751) );
  AND2X1 U8073 ( .IN1(n6752), .IN2(n4371), .Q(WX11654) );
  XOR2X1 U8074 ( .IN1(CRC_OUT_1_22), .IN2(n3210), .Q(n6752) );
  AND2X1 U8075 ( .IN1(n6753), .IN2(n4371), .Q(WX11652) );
  XOR2X1 U8076 ( .IN1(CRC_OUT_1_21), .IN2(n3211), .Q(n6753) );
  AND2X1 U8077 ( .IN1(n6754), .IN2(n4370), .Q(WX11650) );
  XOR2X1 U8078 ( .IN1(CRC_OUT_1_20), .IN2(n3212), .Q(n6754) );
  AND2X1 U8079 ( .IN1(n6755), .IN2(n4370), .Q(WX11648) );
  XOR2X1 U8080 ( .IN1(CRC_OUT_1_19), .IN2(n3213), .Q(n6755) );
  AND2X1 U8081 ( .IN1(n6756), .IN2(n4370), .Q(WX11646) );
  XOR2X1 U8082 ( .IN1(test_so97), .IN2(DFF_1714_n1), .Q(n6756) );
  AND2X1 U8083 ( .IN1(n6757), .IN2(n4370), .Q(WX11644) );
  XOR2X1 U8084 ( .IN1(CRC_OUT_1_17), .IN2(n3214), .Q(n6757) );
  AND2X1 U8085 ( .IN1(n6758), .IN2(n4370), .Q(WX11642) );
  XOR2X1 U8086 ( .IN1(CRC_OUT_1_16), .IN2(n3215), .Q(n6758) );
  AND2X1 U8087 ( .IN1(n6759), .IN2(n4370), .Q(WX11640) );
  XOR3X1 U8088 ( .IN1(test_so100), .IN2(n3173), .IN3(CRC_OUT_1_15), .Q(n6759)
         );
  AND2X1 U8089 ( .IN1(n6760), .IN2(n4370), .Q(WX11638) );
  XOR2X1 U8090 ( .IN1(test_so99), .IN2(n3216), .Q(n6760) );
  AND2X1 U8091 ( .IN1(n6761), .IN2(n4370), .Q(WX11636) );
  XOR2X1 U8092 ( .IN1(CRC_OUT_1_13), .IN2(n3217), .Q(n6761) );
  AND2X1 U8093 ( .IN1(n6762), .IN2(n4370), .Q(WX11634) );
  XOR2X1 U8094 ( .IN1(CRC_OUT_1_12), .IN2(n3218), .Q(n6762) );
  AND2X1 U8095 ( .IN1(n6763), .IN2(n4369), .Q(WX11632) );
  XOR2X1 U8096 ( .IN1(CRC_OUT_1_11), .IN2(n3219), .Q(n6763) );
  AND2X1 U8097 ( .IN1(n6764), .IN2(n4369), .Q(WX11630) );
  XOR3X1 U8098 ( .IN1(test_so100), .IN2(n3174), .IN3(CRC_OUT_1_10), .Q(n6764)
         );
  AND2X1 U8099 ( .IN1(n6765), .IN2(n4369), .Q(WX11628) );
  XOR2X1 U8100 ( .IN1(CRC_OUT_1_9), .IN2(n3220), .Q(n6765) );
  AND2X1 U8101 ( .IN1(n6766), .IN2(n4369), .Q(WX11626) );
  XOR2X1 U8102 ( .IN1(CRC_OUT_1_8), .IN2(n3221), .Q(n6766) );
  AND2X1 U8103 ( .IN1(n6767), .IN2(n4369), .Q(WX11624) );
  XOR2X1 U8104 ( .IN1(CRC_OUT_1_7), .IN2(n3222), .Q(n6767) );
  AND2X1 U8105 ( .IN1(n6768), .IN2(n4369), .Q(WX11622) );
  XOR2X1 U8106 ( .IN1(CRC_OUT_1_6), .IN2(n3223), .Q(n6768) );
  AND2X1 U8107 ( .IN1(n6769), .IN2(n4369), .Q(WX11620) );
  XOR2X1 U8108 ( .IN1(CRC_OUT_1_5), .IN2(n3224), .Q(n6769) );
  AND2X1 U8109 ( .IN1(n6770), .IN2(n4369), .Q(WX11618) );
  XOR2X1 U8110 ( .IN1(CRC_OUT_1_4), .IN2(n3225), .Q(n6770) );
  AND2X1 U8111 ( .IN1(n6771), .IN2(n4369), .Q(WX11616) );
  XOR3X1 U8112 ( .IN1(test_so100), .IN2(n3175), .IN3(CRC_OUT_1_3), .Q(n6771)
         );
  AND2X1 U8113 ( .IN1(n6772), .IN2(n4368), .Q(WX11614) );
  XOR2X1 U8114 ( .IN1(CRC_OUT_1_2), .IN2(n3226), .Q(n6772) );
  AND2X1 U8115 ( .IN1(n6773), .IN2(n4368), .Q(WX11612) );
  XOR2X1 U8116 ( .IN1(test_so98), .IN2(DFF_1697_n1), .Q(n6773) );
  AND2X1 U8117 ( .IN1(n6774), .IN2(n4368), .Q(WX11610) );
  XOR2X1 U8118 ( .IN1(CRC_OUT_1_0), .IN2(n3227), .Q(n6774) );
  AND2X1 U8119 ( .IN1(n6775), .IN2(n4368), .Q(WX11608) );
  XOR2X1 U8120 ( .IN1(test_so100), .IN2(n3194), .Q(n6775) );
  AND2X1 U8121 ( .IN1(n4385), .IN2(n8246), .Q(WX11082) );
  AND2X1 U8122 ( .IN1(n4385), .IN2(n8247), .Q(WX11080) );
  AND2X1 U8123 ( .IN1(n4384), .IN2(n8248), .Q(WX11078) );
  AND2X1 U8124 ( .IN1(n4385), .IN2(n8249), .Q(WX11076) );
  AND2X1 U8125 ( .IN1(n4384), .IN2(n8250), .Q(WX11074) );
  INVX0 U8126 ( .INP(n6776), .ZN(WX11072) );
  OR2X1 U8127 ( .IN1(n4425), .IN2(n7262), .Q(n6776) );
  AND2X1 U8128 ( .IN1(n4386), .IN2(n8252), .Q(WX11070) );
  INVX0 U8129 ( .INP(n6777), .ZN(WX11068) );
  OR2X1 U8130 ( .IN1(n4425), .IN2(n7263), .Q(n6777) );
  AND2X1 U8131 ( .IN1(n4385), .IN2(n8254), .Q(WX11066) );
  AND2X1 U8132 ( .IN1(test_so91), .IN2(n4368), .Q(WX11064) );
  AND2X1 U8133 ( .IN1(n4385), .IN2(n8257), .Q(WX11062) );
  AND2X1 U8134 ( .IN1(n4386), .IN2(n8258), .Q(WX11060) );
  AND2X1 U8135 ( .IN1(n4386), .IN2(n8259), .Q(WX11058) );
  AND2X1 U8136 ( .IN1(n4385), .IN2(n8260), .Q(WX11056) );
  AND2X1 U8137 ( .IN1(n4385), .IN2(n8261), .Q(WX11054) );
  AND2X1 U8138 ( .IN1(n4385), .IN2(n8262), .Q(WX11052) );
  OR4X1 U8139 ( .IN1(n6778), .IN2(n6779), .IN3(n6780), .IN4(n6781), .Q(WX11050) );
  AND2X1 U8140 ( .IN1(n498), .IN2(n3562), .Q(n6781) );
  INVX0 U8141 ( .INP(n6782), .ZN(n498) );
  OR2X1 U8142 ( .IN1(n4425), .IN2(n3786), .Q(n6782) );
  AND2X1 U8143 ( .IN1(n3545), .IN2(n4693), .Q(n6780) );
  XNOR3X1 U8144 ( .IN1(n3194), .IN2(n3059), .IN3(n6783), .Q(n4693) );
  XOR2X1 U8145 ( .IN1(WX11115), .IN2(n7250), .Q(n6783) );
  AND2X1 U8146 ( .IN1(n3597), .IN2(CRC_OUT_1_0), .Q(n6779) );
  AND2X1 U8147 ( .IN1(DATA_0_0), .IN2(n3623), .Q(n6778) );
  OR4X1 U8148 ( .IN1(n6784), .IN2(n6785), .IN3(n6786), .IN4(n6787), .Q(WX11048) );
  AND2X1 U8149 ( .IN1(n497), .IN2(n3562), .Q(n6787) );
  INVX0 U8150 ( .INP(n6788), .ZN(n497) );
  OR2X1 U8151 ( .IN1(n4425), .IN2(n3787), .Q(n6788) );
  AND2X1 U8152 ( .IN1(n3545), .IN2(n4701), .Q(n6786) );
  XNOR3X1 U8153 ( .IN1(n3227), .IN2(n3060), .IN3(n6789), .Q(n4701) );
  XOR2X1 U8154 ( .IN1(WX11113), .IN2(n7251), .Q(n6789) );
  AND2X1 U8155 ( .IN1(n3597), .IN2(CRC_OUT_1_1), .Q(n6785) );
  AND2X1 U8156 ( .IN1(DATA_0_1), .IN2(n3624), .Q(n6784) );
  OR4X1 U8157 ( .IN1(n6790), .IN2(n6791), .IN3(n6792), .IN4(n6793), .Q(WX11046) );
  AND2X1 U8158 ( .IN1(n496), .IN2(n3562), .Q(n6793) );
  INVX0 U8159 ( .INP(n6794), .ZN(n496) );
  OR2X1 U8160 ( .IN1(n4425), .IN2(n3788), .Q(n6794) );
  AND2X1 U8161 ( .IN1(n4708), .IN2(n3530), .Q(n6792) );
  XOR3X1 U8162 ( .IN1(n3535), .IN2(n3061), .IN3(n6795), .Q(n4708) );
  XOR2X1 U8163 ( .IN1(WX11047), .IN2(test_so98), .Q(n6795) );
  AND2X1 U8164 ( .IN1(n3597), .IN2(CRC_OUT_1_2), .Q(n6791) );
  AND2X1 U8165 ( .IN1(DATA_0_2), .IN2(n3626), .Q(n6790) );
  OR4X1 U8166 ( .IN1(n6796), .IN2(n6797), .IN3(n6798), .IN4(n6799), .Q(WX11044) );
  AND2X1 U8167 ( .IN1(n495), .IN2(n3562), .Q(n6799) );
  INVX0 U8168 ( .INP(n6800), .ZN(n495) );
  OR2X1 U8169 ( .IN1(n4425), .IN2(n3789), .Q(n6800) );
  AND2X1 U8170 ( .IN1(n3545), .IN2(n4715), .Q(n6798) );
  XNOR3X1 U8171 ( .IN1(n3226), .IN2(n3062), .IN3(n6801), .Q(n4715) );
  XOR2X1 U8172 ( .IN1(WX11109), .IN2(n7252), .Q(n6801) );
  AND2X1 U8173 ( .IN1(n3597), .IN2(CRC_OUT_1_3), .Q(n6797) );
  AND2X1 U8174 ( .IN1(DATA_0_3), .IN2(n3626), .Q(n6796) );
  OR4X1 U8175 ( .IN1(n6802), .IN2(n6803), .IN3(n6804), .IN4(n6805), .Q(WX11042) );
  AND2X1 U8176 ( .IN1(n494), .IN2(n3562), .Q(n6805) );
  INVX0 U8177 ( .INP(n6806), .ZN(n494) );
  OR2X1 U8178 ( .IN1(n4425), .IN2(n3790), .Q(n6806) );
  AND2X1 U8179 ( .IN1(n4722), .IN2(n3530), .Q(n6804) );
  XOR3X1 U8180 ( .IN1(n3539), .IN2(n3175), .IN3(n6807), .Q(n4722) );
  XOR2X1 U8181 ( .IN1(WX11043), .IN2(test_so96), .Q(n6807) );
  AND2X1 U8182 ( .IN1(n3597), .IN2(CRC_OUT_1_4), .Q(n6803) );
  AND2X1 U8183 ( .IN1(DATA_0_4), .IN2(n3626), .Q(n6802) );
  OR4X1 U8184 ( .IN1(n6808), .IN2(n6809), .IN3(n6810), .IN4(n6811), .Q(WX11040) );
  AND2X1 U8185 ( .IN1(n493), .IN2(n3562), .Q(n6811) );
  INVX0 U8186 ( .INP(n6812), .ZN(n493) );
  OR2X1 U8187 ( .IN1(n4425), .IN2(n3791), .Q(n6812) );
  AND2X1 U8188 ( .IN1(n3545), .IN2(n4729), .Q(n6810) );
  XNOR3X1 U8189 ( .IN1(n3225), .IN2(n3063), .IN3(n6813), .Q(n4729) );
  XOR2X1 U8190 ( .IN1(WX11105), .IN2(n7253), .Q(n6813) );
  AND2X1 U8191 ( .IN1(n3597), .IN2(CRC_OUT_1_5), .Q(n6809) );
  AND2X1 U8192 ( .IN1(DATA_0_5), .IN2(n3626), .Q(n6808) );
  OR4X1 U8193 ( .IN1(n6814), .IN2(n6815), .IN3(n6816), .IN4(n6817), .Q(WX11038) );
  AND2X1 U8194 ( .IN1(n492), .IN2(n3562), .Q(n6817) );
  INVX0 U8195 ( .INP(n6818), .ZN(n492) );
  OR2X1 U8196 ( .IN1(n4424), .IN2(n3792), .Q(n6818) );
  AND2X1 U8197 ( .IN1(n4736), .IN2(n3530), .Q(n6816) );
  XOR3X1 U8198 ( .IN1(n3224), .IN2(n3064), .IN3(n6819), .Q(n4736) );
  XOR2X1 U8199 ( .IN1(WX11039), .IN2(test_so94), .Q(n6819) );
  AND2X1 U8200 ( .IN1(n3597), .IN2(CRC_OUT_1_6), .Q(n6815) );
  AND2X1 U8201 ( .IN1(DATA_0_6), .IN2(n3626), .Q(n6814) );
  OR4X1 U8202 ( .IN1(n6820), .IN2(n6821), .IN3(n6822), .IN4(n6823), .Q(WX11036) );
  AND2X1 U8203 ( .IN1(n491), .IN2(n3561), .Q(n6823) );
  INVX0 U8204 ( .INP(n6824), .ZN(n491) );
  OR2X1 U8205 ( .IN1(n4424), .IN2(n3793), .Q(n6824) );
  AND2X1 U8206 ( .IN1(n3545), .IN2(n4743), .Q(n6822) );
  XNOR3X1 U8207 ( .IN1(n3223), .IN2(n3065), .IN3(n6825), .Q(n4743) );
  XOR2X1 U8208 ( .IN1(WX11101), .IN2(n7254), .Q(n6825) );
  AND2X1 U8209 ( .IN1(n3597), .IN2(CRC_OUT_1_7), .Q(n6821) );
  AND2X1 U8210 ( .IN1(DATA_0_7), .IN2(n3627), .Q(n6820) );
  OR4X1 U8211 ( .IN1(n6826), .IN2(n6827), .IN3(n6828), .IN4(n6829), .Q(WX11034) );
  AND2X1 U8212 ( .IN1(n490), .IN2(n3561), .Q(n6829) );
  INVX0 U8213 ( .INP(n6830), .ZN(n490) );
  OR2X1 U8214 ( .IN1(n4424), .IN2(n3794), .Q(n6830) );
  AND2X1 U8215 ( .IN1(n4750), .IN2(n3530), .Q(n6828) );
  XOR3X1 U8216 ( .IN1(n3547), .IN2(n3222), .IN3(n6831), .Q(n4750) );
  XOR2X1 U8217 ( .IN1(WX11163), .IN2(test_so92), .Q(n6831) );
  AND2X1 U8218 ( .IN1(n3597), .IN2(CRC_OUT_1_8), .Q(n6827) );
  AND2X1 U8219 ( .IN1(DATA_0_8), .IN2(n3627), .Q(n6826) );
  OR4X1 U8220 ( .IN1(n6832), .IN2(n6833), .IN3(n6834), .IN4(n6835), .Q(WX11032) );
  AND2X1 U8221 ( .IN1(n489), .IN2(n3561), .Q(n6835) );
  INVX0 U8222 ( .INP(n6836), .ZN(n489) );
  OR2X1 U8223 ( .IN1(n4424), .IN2(n3795), .Q(n6836) );
  AND2X1 U8224 ( .IN1(n3545), .IN2(n4757), .Q(n6834) );
  XNOR3X1 U8225 ( .IN1(n3221), .IN2(n3066), .IN3(n6837), .Q(n4757) );
  XOR2X1 U8226 ( .IN1(WX11097), .IN2(n7255), .Q(n6837) );
  AND2X1 U8227 ( .IN1(n3597), .IN2(CRC_OUT_1_9), .Q(n6833) );
  AND2X1 U8228 ( .IN1(DATA_0_9), .IN2(n3627), .Q(n6832) );
  OR4X1 U8229 ( .IN1(n6838), .IN2(n6839), .IN3(n6840), .IN4(n6841), .Q(WX11030) );
  AND2X1 U8230 ( .IN1(n488), .IN2(n3561), .Q(n6841) );
  INVX0 U8231 ( .INP(n6842), .ZN(n488) );
  OR2X1 U8232 ( .IN1(n4424), .IN2(n3796), .Q(n6842) );
  AND2X1 U8233 ( .IN1(n3545), .IN2(n4764), .Q(n6840) );
  XNOR3X1 U8234 ( .IN1(n3220), .IN2(n3067), .IN3(n6843), .Q(n4764) );
  XOR2X1 U8235 ( .IN1(WX11095), .IN2(n7256), .Q(n6843) );
  AND2X1 U8236 ( .IN1(n3598), .IN2(CRC_OUT_1_10), .Q(n6839) );
  AND2X1 U8237 ( .IN1(DATA_0_10), .IN2(n3627), .Q(n6838) );
  OR4X1 U8238 ( .IN1(n6844), .IN2(n6845), .IN3(n6846), .IN4(n6847), .Q(WX11028) );
  AND2X1 U8239 ( .IN1(n487), .IN2(n3561), .Q(n6847) );
  INVX0 U8240 ( .INP(n6848), .ZN(n487) );
  OR2X1 U8241 ( .IN1(n4424), .IN2(n3797), .Q(n6848) );
  AND2X1 U8242 ( .IN1(n3545), .IN2(n4771), .Q(n6846) );
  XNOR3X1 U8243 ( .IN1(n3174), .IN2(n3068), .IN3(n6849), .Q(n4771) );
  XOR2X1 U8244 ( .IN1(WX11093), .IN2(n7257), .Q(n6849) );
  AND2X1 U8245 ( .IN1(n3598), .IN2(CRC_OUT_1_11), .Q(n6845) );
  AND2X1 U8246 ( .IN1(DATA_0_11), .IN2(n3624), .Q(n6844) );
  OR4X1 U8247 ( .IN1(n6850), .IN2(n6851), .IN3(n6852), .IN4(n6853), .Q(WX11026) );
  AND2X1 U8248 ( .IN1(n486), .IN2(n3561), .Q(n6853) );
  INVX0 U8249 ( .INP(n6854), .ZN(n486) );
  OR2X1 U8250 ( .IN1(n4424), .IN2(n3798), .Q(n6854) );
  AND2X1 U8251 ( .IN1(n3544), .IN2(n4778), .Q(n6852) );
  XNOR3X1 U8252 ( .IN1(n3219), .IN2(n3069), .IN3(n6855), .Q(n4778) );
  XOR2X1 U8253 ( .IN1(WX11091), .IN2(n7258), .Q(n6855) );
  AND2X1 U8254 ( .IN1(n3598), .IN2(CRC_OUT_1_12), .Q(n6851) );
  AND2X1 U8255 ( .IN1(DATA_0_12), .IN2(n3627), .Q(n6850) );
  OR4X1 U8256 ( .IN1(n6856), .IN2(n6857), .IN3(n6858), .IN4(n6859), .Q(WX11024) );
  AND2X1 U8257 ( .IN1(n485), .IN2(n3561), .Q(n6859) );
  INVX0 U8258 ( .INP(n6860), .ZN(n485) );
  OR2X1 U8259 ( .IN1(n4424), .IN2(n3799), .Q(n6860) );
  AND2X1 U8260 ( .IN1(n3544), .IN2(n4785), .Q(n6858) );
  XNOR3X1 U8261 ( .IN1(n3218), .IN2(n3070), .IN3(n6861), .Q(n4785) );
  XOR2X1 U8262 ( .IN1(WX11089), .IN2(n7259), .Q(n6861) );
  AND2X1 U8263 ( .IN1(n3598), .IN2(CRC_OUT_1_13), .Q(n6857) );
  AND2X1 U8264 ( .IN1(DATA_0_13), .IN2(n3627), .Q(n6856) );
  OR4X1 U8265 ( .IN1(n6862), .IN2(n6863), .IN3(n6864), .IN4(n6865), .Q(WX11022) );
  AND2X1 U8266 ( .IN1(n484), .IN2(n3561), .Q(n6865) );
  INVX0 U8267 ( .INP(n6866), .ZN(n484) );
  OR2X1 U8268 ( .IN1(n4424), .IN2(n3800), .Q(n6866) );
  AND2X1 U8269 ( .IN1(n3544), .IN2(n4792), .Q(n6864) );
  XNOR3X1 U8270 ( .IN1(n3217), .IN2(n3071), .IN3(n6867), .Q(n4792) );
  XOR2X1 U8271 ( .IN1(WX11087), .IN2(n7260), .Q(n6867) );
  AND2X1 U8272 ( .IN1(test_so99), .IN2(n3587), .Q(n6863) );
  AND2X1 U8273 ( .IN1(DATA_0_14), .IN2(n3628), .Q(n6862) );
  OR4X1 U8274 ( .IN1(n6868), .IN2(n6869), .IN3(n6870), .IN4(n6871), .Q(WX11020) );
  AND2X1 U8275 ( .IN1(n483), .IN2(n3561), .Q(n6871) );
  INVX0 U8276 ( .INP(n6872), .ZN(n483) );
  OR2X1 U8277 ( .IN1(n4424), .IN2(n3801), .Q(n6872) );
  AND2X1 U8278 ( .IN1(n3544), .IN2(n4799), .Q(n6870) );
  XNOR3X1 U8279 ( .IN1(n3216), .IN2(n3072), .IN3(n6873), .Q(n4799) );
  XOR2X1 U8280 ( .IN1(WX11085), .IN2(n7261), .Q(n6873) );
  AND2X1 U8281 ( .IN1(n3598), .IN2(CRC_OUT_1_15), .Q(n6869) );
  AND2X1 U8282 ( .IN1(DATA_0_15), .IN2(n3628), .Q(n6868) );
  OR4X1 U8283 ( .IN1(n6874), .IN2(n6875), .IN3(n6876), .IN4(n6877), .Q(WX11018) );
  AND2X1 U8284 ( .IN1(n482), .IN2(n3561), .Q(n6877) );
  INVX0 U8285 ( .INP(n6878), .ZN(n482) );
  OR2X1 U8286 ( .IN1(n4424), .IN2(n3802), .Q(n6878) );
  AND2X1 U8287 ( .IN1(n3544), .IN2(n4806), .Q(n6876) );
  XOR3X1 U8288 ( .IN1(n2847), .IN2(n3518), .IN3(n6879), .Q(n4806) );
  XNOR3X1 U8289 ( .IN1(n8246), .IN2(n3173), .IN3(WX11147), .Q(n6879) );
  AND2X1 U8290 ( .IN1(n3598), .IN2(CRC_OUT_1_16), .Q(n6875) );
  AND2X1 U8291 ( .IN1(DATA_0_16), .IN2(n3627), .Q(n6874) );
  OR4X1 U8292 ( .IN1(n6880), .IN2(n6881), .IN3(n6882), .IN4(n6883), .Q(WX11016) );
  AND2X1 U8293 ( .IN1(n481), .IN2(n3561), .Q(n6883) );
  INVX0 U8294 ( .INP(n6884), .ZN(n481) );
  OR2X1 U8295 ( .IN1(n4424), .IN2(n3803), .Q(n6884) );
  AND2X1 U8296 ( .IN1(n3544), .IN2(n4813), .Q(n6882) );
  XOR3X1 U8297 ( .IN1(n2849), .IN2(n3516), .IN3(n6885), .Q(n4813) );
  XNOR3X1 U8298 ( .IN1(n8247), .IN2(n3215), .IN3(WX11145), .Q(n6885) );
  AND2X1 U8299 ( .IN1(n3598), .IN2(CRC_OUT_1_17), .Q(n6881) );
  AND2X1 U8300 ( .IN1(DATA_0_17), .IN2(n3628), .Q(n6880) );
  OR4X1 U8301 ( .IN1(n6886), .IN2(n6887), .IN3(n6888), .IN4(n6889), .Q(WX11014) );
  AND2X1 U8302 ( .IN1(n480), .IN2(n3561), .Q(n6889) );
  INVX0 U8303 ( .INP(n6890), .ZN(n480) );
  OR2X1 U8304 ( .IN1(n4424), .IN2(n3804), .Q(n6890) );
  AND2X1 U8305 ( .IN1(n3544), .IN2(n4820), .Q(n6888) );
  XOR3X1 U8306 ( .IN1(n2851), .IN2(n3515), .IN3(n6891), .Q(n4820) );
  XNOR3X1 U8307 ( .IN1(n8248), .IN2(n3214), .IN3(WX11143), .Q(n6891) );
  AND2X1 U8308 ( .IN1(n3598), .IN2(CRC_OUT_1_18), .Q(n6887) );
  AND2X1 U8309 ( .IN1(DATA_0_18), .IN2(n3626), .Q(n6886) );
  OR4X1 U8310 ( .IN1(n6892), .IN2(n6893), .IN3(n6894), .IN4(n6895), .Q(WX11012) );
  AND2X1 U8311 ( .IN1(n479), .IN2(n3560), .Q(n6895) );
  INVX0 U8312 ( .INP(n6896), .ZN(n479) );
  OR2X1 U8313 ( .IN1(n4423), .IN2(n3805), .Q(n6896) );
  AND2X1 U8314 ( .IN1(n4827), .IN2(n3528), .Q(n6894) );
  XOR3X1 U8315 ( .IN1(n2853), .IN2(TM1), .IN3(n6897), .Q(n4827) );
  XNOR3X1 U8316 ( .IN1(test_so97), .IN2(n8249), .IN3(WX11141), .Q(n6897) );
  AND2X1 U8317 ( .IN1(n3598), .IN2(CRC_OUT_1_19), .Q(n6893) );
  AND2X1 U8318 ( .IN1(DATA_0_19), .IN2(n3624), .Q(n6892) );
  OR4X1 U8319 ( .IN1(n6898), .IN2(n6899), .IN3(n6900), .IN4(n6901), .Q(WX11010) );
  AND2X1 U8320 ( .IN1(n478), .IN2(n3560), .Q(n6901) );
  INVX0 U8321 ( .INP(n6902), .ZN(n478) );
  OR2X1 U8322 ( .IN1(n4423), .IN2(n3806), .Q(n6902) );
  AND2X1 U8323 ( .IN1(n3544), .IN2(n4834), .Q(n6900) );
  XOR3X1 U8324 ( .IN1(n2854), .IN2(n3514), .IN3(n6903), .Q(n4834) );
  XNOR3X1 U8325 ( .IN1(n8250), .IN2(n3213), .IN3(WX11139), .Q(n6903) );
  AND2X1 U8326 ( .IN1(n3598), .IN2(CRC_OUT_1_20), .Q(n6899) );
  AND2X1 U8327 ( .IN1(DATA_0_20), .IN2(n3628), .Q(n6898) );
  OR4X1 U8328 ( .IN1(n6904), .IN2(n6905), .IN3(n6906), .IN4(n6907), .Q(WX11008) );
  AND2X1 U8329 ( .IN1(n477), .IN2(n3560), .Q(n6907) );
  INVX0 U8330 ( .INP(n6908), .ZN(n477) );
  OR2X1 U8331 ( .IN1(n4423), .IN2(n3807), .Q(n6908) );
  AND2X1 U8332 ( .IN1(n4841), .IN2(n3528), .Q(n6906) );
  XOR3X1 U8333 ( .IN1(n2856), .IN2(TM1), .IN3(n6909), .Q(n4841) );
  XNOR3X1 U8334 ( .IN1(test_so95), .IN2(n7262), .IN3(n3212), .Q(n6909) );
  AND2X1 U8335 ( .IN1(n3598), .IN2(CRC_OUT_1_21), .Q(n6905) );
  AND2X1 U8336 ( .IN1(DATA_0_21), .IN2(n3626), .Q(n6904) );
  OR4X1 U8337 ( .IN1(n6910), .IN2(n6911), .IN3(n6912), .IN4(n6913), .Q(WX11006) );
  AND2X1 U8338 ( .IN1(n476), .IN2(n3560), .Q(n6913) );
  INVX0 U8339 ( .INP(n6914), .ZN(n476) );
  OR2X1 U8340 ( .IN1(n4423), .IN2(n3808), .Q(n6914) );
  AND2X1 U8341 ( .IN1(n3544), .IN2(n4848), .Q(n6912) );
  XOR3X1 U8342 ( .IN1(n2857), .IN2(n3518), .IN3(n6915), .Q(n4848) );
  XNOR3X1 U8343 ( .IN1(n8252), .IN2(n3211), .IN3(WX11135), .Q(n6915) );
  AND2X1 U8344 ( .IN1(n3598), .IN2(CRC_OUT_1_22), .Q(n6911) );
  AND2X1 U8345 ( .IN1(DATA_0_22), .IN2(n3627), .Q(n6910) );
  OR4X1 U8346 ( .IN1(n6916), .IN2(n6917), .IN3(n6918), .IN4(n6919), .Q(WX11004) );
  AND2X1 U8347 ( .IN1(n475), .IN2(n3560), .Q(n6919) );
  INVX0 U8348 ( .INP(n6920), .ZN(n475) );
  OR2X1 U8349 ( .IN1(n4423), .IN2(n3809), .Q(n6920) );
  AND2X1 U8350 ( .IN1(n4855), .IN2(n3528), .Q(n6918) );
  XOR3X1 U8351 ( .IN1(n2859), .IN2(TM1), .IN3(n6921), .Q(n4855) );
  XNOR3X1 U8352 ( .IN1(test_so93), .IN2(n7263), .IN3(n3210), .Q(n6921) );
  AND2X1 U8353 ( .IN1(n3598), .IN2(CRC_OUT_1_23), .Q(n6917) );
  AND2X1 U8354 ( .IN1(DATA_0_23), .IN2(n3624), .Q(n6916) );
  OR4X1 U8355 ( .IN1(n6922), .IN2(n6923), .IN3(n6924), .IN4(n6925), .Q(WX11002) );
  AND2X1 U8356 ( .IN1(n474), .IN2(n3560), .Q(n6925) );
  INVX0 U8357 ( .INP(n6926), .ZN(n474) );
  OR2X1 U8358 ( .IN1(n4423), .IN2(n3810), .Q(n6926) );
  AND2X1 U8359 ( .IN1(n3544), .IN2(n4862), .Q(n6924) );
  XOR3X1 U8360 ( .IN1(n2860), .IN2(n3516), .IN3(n6927), .Q(n4862) );
  XNOR3X1 U8361 ( .IN1(n8254), .IN2(n3209), .IN3(WX11131), .Q(n6927) );
  AND2X1 U8362 ( .IN1(n3599), .IN2(CRC_OUT_1_24), .Q(n6923) );
  AND2X1 U8363 ( .IN1(DATA_0_24), .IN2(n3626), .Q(n6922) );
  OR4X1 U8364 ( .IN1(n6928), .IN2(n6929), .IN3(n6930), .IN4(n6931), .Q(WX11000) );
  AND2X1 U8365 ( .IN1(n473), .IN2(n3560), .Q(n6931) );
  INVX0 U8366 ( .INP(n6932), .ZN(n473) );
  OR2X1 U8367 ( .IN1(n4423), .IN2(n3811), .Q(n6932) );
  AND2X1 U8368 ( .IN1(n4869), .IN2(n3528), .Q(n6930) );
  XOR3X1 U8369 ( .IN1(n2862), .IN2(TM1), .IN3(n6933), .Q(n4869) );
  XNOR3X1 U8370 ( .IN1(test_so91), .IN2(n7264), .IN3(n3208), .Q(n6933) );
  AND2X1 U8371 ( .IN1(n3599), .IN2(CRC_OUT_1_25), .Q(n6929) );
  AND2X1 U8372 ( .IN1(DATA_0_25), .IN2(n3627), .Q(n6928) );
  OR4X1 U8373 ( .IN1(n6934), .IN2(n6935), .IN3(n6936), .IN4(n6937), .Q(WX10998) );
  AND2X1 U8374 ( .IN1(n472), .IN2(n3560), .Q(n6937) );
  INVX0 U8375 ( .INP(n6938), .ZN(n472) );
  OR2X1 U8376 ( .IN1(n4423), .IN2(n3812), .Q(n6938) );
  AND2X1 U8377 ( .IN1(n3544), .IN2(n4876), .Q(n6936) );
  XOR3X1 U8378 ( .IN1(n2863), .IN2(n3515), .IN3(n6939), .Q(n4876) );
  XNOR3X1 U8379 ( .IN1(n8257), .IN2(n3207), .IN3(WX11127), .Q(n6939) );
  AND2X1 U8380 ( .IN1(n3599), .IN2(CRC_OUT_1_26), .Q(n6935) );
  AND2X1 U8381 ( .IN1(DATA_0_26), .IN2(n3627), .Q(n6934) );
  OR4X1 U8382 ( .IN1(n6940), .IN2(n6941), .IN3(n6942), .IN4(n6943), .Q(WX10996) );
  AND2X1 U8383 ( .IN1(n471), .IN2(n3560), .Q(n6943) );
  INVX0 U8384 ( .INP(n6944), .ZN(n471) );
  OR2X1 U8385 ( .IN1(n4423), .IN2(n3813), .Q(n6944) );
  AND2X1 U8386 ( .IN1(n3544), .IN2(n4883), .Q(n6942) );
  XOR3X1 U8387 ( .IN1(n2865), .IN2(n3514), .IN3(n6945), .Q(n4883) );
  XNOR3X1 U8388 ( .IN1(n8258), .IN2(n3206), .IN3(WX11125), .Q(n6945) );
  AND2X1 U8389 ( .IN1(n3599), .IN2(CRC_OUT_1_27), .Q(n6941) );
  AND2X1 U8390 ( .IN1(DATA_0_27), .IN2(n3626), .Q(n6940) );
  OR4X1 U8391 ( .IN1(n6946), .IN2(n6947), .IN3(n6948), .IN4(n6949), .Q(WX10994) );
  AND2X1 U8392 ( .IN1(n470), .IN2(n3560), .Q(n6949) );
  INVX0 U8393 ( .INP(n6950), .ZN(n470) );
  OR2X1 U8394 ( .IN1(n4423), .IN2(n3814), .Q(n6950) );
  AND2X1 U8395 ( .IN1(n3544), .IN2(n4890), .Q(n6948) );
  XOR3X1 U8396 ( .IN1(n2867), .IN2(n3518), .IN3(n6951), .Q(n4890) );
  XNOR3X1 U8397 ( .IN1(n8259), .IN2(n3205), .IN3(WX11123), .Q(n6951) );
  AND2X1 U8398 ( .IN1(n3599), .IN2(CRC_OUT_1_28), .Q(n6947) );
  AND2X1 U8399 ( .IN1(DATA_0_28), .IN2(n3624), .Q(n6946) );
  OR4X1 U8400 ( .IN1(n6952), .IN2(n6953), .IN3(n6954), .IN4(n6955), .Q(WX10992) );
  AND2X1 U8401 ( .IN1(n469), .IN2(n3560), .Q(n6955) );
  INVX0 U8402 ( .INP(n6956), .ZN(n469) );
  OR2X1 U8403 ( .IN1(n4423), .IN2(n3815), .Q(n6956) );
  AND2X1 U8404 ( .IN1(n3543), .IN2(n4897), .Q(n6954) );
  XOR3X1 U8405 ( .IN1(n2869), .IN2(n3516), .IN3(n6957), .Q(n4897) );
  XNOR3X1 U8406 ( .IN1(n8260), .IN2(n3204), .IN3(WX11121), .Q(n6957) );
  AND2X1 U8407 ( .IN1(n3599), .IN2(CRC_OUT_1_29), .Q(n6953) );
  AND2X1 U8408 ( .IN1(DATA_0_29), .IN2(n3624), .Q(n6952) );
  OR4X1 U8409 ( .IN1(n6958), .IN2(n6959), .IN3(n6960), .IN4(n6961), .Q(WX10990) );
  AND2X1 U8410 ( .IN1(n468), .IN2(n3560), .Q(n6961) );
  AND2X1 U8411 ( .IN1(TM0), .IN2(TM1), .Q(n2148) );
  INVX0 U8412 ( .INP(n6962), .ZN(n468) );
  OR2X1 U8413 ( .IN1(n4432), .IN2(n3816), .Q(n6962) );
  AND2X1 U8414 ( .IN1(n3549), .IN2(n4904), .Q(n6960) );
  XOR3X1 U8415 ( .IN1(n2871), .IN2(n3515), .IN3(n6963), .Q(n4904) );
  XNOR3X1 U8416 ( .IN1(n8261), .IN2(n3203), .IN3(WX11119), .Q(n6963) );
  AND2X1 U8417 ( .IN1(n3599), .IN2(CRC_OUT_1_30), .Q(n6959) );
  AND2X1 U8418 ( .IN1(DATA_0_30), .IN2(n3624), .Q(n6958) );
  OR4X1 U8419 ( .IN1(n6964), .IN2(n6965), .IN3(n6966), .IN4(n6967), .Q(WX10988) );
  AND2X1 U8420 ( .IN1(DATA_0_31), .IN2(n3622), .Q(n6967) );
  AND2X1 U8421 ( .IN1(n3536), .IN2(n4911), .Q(n6966) );
  XOR3X1 U8422 ( .IN1(n2832), .IN2(n3514), .IN3(n6968), .Q(n4911) );
  XNOR3X1 U8423 ( .IN1(n8262), .IN2(n3202), .IN3(WX11117), .Q(n6968) );
  AND3X1 U8424 ( .IN1(n530), .IN2(n4387), .IN3(TM1), .Q(n4694) );
  AND2X1 U8425 ( .IN1(n2245), .IN2(WX10829), .Q(n6965) );
  AND2X1 U8426 ( .IN1(test_so100), .IN2(n3588), .Q(n6964) );
  AND2X1 U8427 ( .IN1(n3510), .IN2(n4368), .Q(WX10890) );
  AND2X1 U8428 ( .IN1(n6969), .IN2(n4368), .Q(WX10377) );
  XOR2X1 U8429 ( .IN1(test_so85), .IN2(DFF_1534_n1), .Q(n6969) );
  AND2X1 U8430 ( .IN1(n6970), .IN2(n4368), .Q(WX10375) );
  XOR2X1 U8431 ( .IN1(CRC_OUT_2_29), .IN2(n3228), .Q(n6970) );
  AND2X1 U8432 ( .IN1(n6971), .IN2(n4368), .Q(WX10373) );
  XOR2X1 U8433 ( .IN1(CRC_OUT_2_28), .IN2(n3229), .Q(n6971) );
  AND2X1 U8434 ( .IN1(n6972), .IN2(n4367), .Q(WX10371) );
  XOR2X1 U8435 ( .IN1(CRC_OUT_2_27), .IN2(n3230), .Q(n6972) );
  AND2X1 U8436 ( .IN1(n6973), .IN2(n4367), .Q(WX10369) );
  XOR2X1 U8437 ( .IN1(CRC_OUT_2_26), .IN2(n3231), .Q(n6973) );
  AND2X1 U8438 ( .IN1(n6974), .IN2(n4367), .Q(WX10367) );
  XOR2X1 U8439 ( .IN1(CRC_OUT_2_25), .IN2(n3232), .Q(n6974) );
  AND2X1 U8440 ( .IN1(n6975), .IN2(n4367), .Q(WX10365) );
  XOR2X1 U8441 ( .IN1(CRC_OUT_2_24), .IN2(n3233), .Q(n6975) );
  AND2X1 U8442 ( .IN1(n6976), .IN2(n4367), .Q(WX10363) );
  XOR2X1 U8443 ( .IN1(CRC_OUT_2_23), .IN2(n3234), .Q(n6976) );
  AND2X1 U8444 ( .IN1(n6977), .IN2(n4367), .Q(WX10361) );
  XOR2X1 U8445 ( .IN1(CRC_OUT_2_22), .IN2(n3235), .Q(n6977) );
  AND2X1 U8446 ( .IN1(n6978), .IN2(n4367), .Q(WX10359) );
  XOR2X1 U8447 ( .IN1(CRC_OUT_2_21), .IN2(n3236), .Q(n6978) );
  AND2X1 U8448 ( .IN1(n6979), .IN2(n4367), .Q(WX10357) );
  XOR2X1 U8449 ( .IN1(CRC_OUT_2_20), .IN2(n3237), .Q(n6979) );
  AND2X1 U8450 ( .IN1(n6980), .IN2(n4367), .Q(WX10355) );
  XOR2X1 U8451 ( .IN1(test_so88), .IN2(n3238), .Q(n6980) );
  AND2X1 U8452 ( .IN1(n6981), .IN2(n4366), .Q(WX10353) );
  XOR2X1 U8453 ( .IN1(CRC_OUT_2_18), .IN2(n3239), .Q(n6981) );
  AND2X1 U8454 ( .IN1(n6982), .IN2(n4366), .Q(WX10351) );
  XOR2X1 U8455 ( .IN1(CRC_OUT_2_17), .IN2(n3240), .Q(n6982) );
  AND2X1 U8456 ( .IN1(n6983), .IN2(n4366), .Q(WX10349) );
  XOR2X1 U8457 ( .IN1(CRC_OUT_2_16), .IN2(n3241), .Q(n6983) );
  AND2X1 U8458 ( .IN1(n6984), .IN2(n4366), .Q(WX10347) );
  XOR3X1 U8459 ( .IN1(n3176), .IN2(DFF_1535_n1), .IN3(DFF_1519_n1), .Q(n6984)
         );
  AND2X1 U8460 ( .IN1(n6985), .IN2(n4366), .Q(WX10345) );
  XOR2X1 U8461 ( .IN1(CRC_OUT_2_14), .IN2(n3242), .Q(n6985) );
  AND2X1 U8462 ( .IN1(n6986), .IN2(n4366), .Q(WX10343) );
  XOR2X1 U8463 ( .IN1(test_so86), .IN2(DFF_1517_n1), .Q(n6986) );
  AND2X1 U8464 ( .IN1(n6987), .IN2(n4366), .Q(WX10341) );
  XOR2X1 U8465 ( .IN1(CRC_OUT_2_12), .IN2(n3243), .Q(n6987) );
  AND2X1 U8466 ( .IN1(n6988), .IN2(n4366), .Q(WX10339) );
  XOR2X1 U8467 ( .IN1(CRC_OUT_2_11), .IN2(n3244), .Q(n6988) );
  AND2X1 U8468 ( .IN1(n6989), .IN2(n4366), .Q(WX10337) );
  XOR3X1 U8469 ( .IN1(n3177), .IN2(DFF_1535_n1), .IN3(DFF_1514_n1), .Q(n6989)
         );
  AND2X1 U8470 ( .IN1(n6990), .IN2(n4365), .Q(WX10335) );
  XOR2X1 U8471 ( .IN1(CRC_OUT_2_9), .IN2(n3245), .Q(n6990) );
  AND2X1 U8472 ( .IN1(n6991), .IN2(n4365), .Q(WX10333) );
  XOR2X1 U8473 ( .IN1(CRC_OUT_2_8), .IN2(n3246), .Q(n6991) );
  AND2X1 U8474 ( .IN1(n6992), .IN2(n4365), .Q(WX10331) );
  XOR2X1 U8475 ( .IN1(CRC_OUT_2_7), .IN2(n3247), .Q(n6992) );
  AND2X1 U8476 ( .IN1(n6993), .IN2(n4365), .Q(WX10329) );
  XOR2X1 U8477 ( .IN1(CRC_OUT_2_6), .IN2(n3248), .Q(n6993) );
  AND2X1 U8478 ( .IN1(n6994), .IN2(n4365), .Q(WX10327) );
  XOR2X1 U8479 ( .IN1(CRC_OUT_2_5), .IN2(n3249), .Q(n6994) );
  AND2X1 U8480 ( .IN1(n6995), .IN2(n4365), .Q(WX10325) );
  XOR2X1 U8481 ( .IN1(CRC_OUT_2_4), .IN2(n3250), .Q(n6995) );
  AND2X1 U8482 ( .IN1(n6996), .IN2(n4365), .Q(WX10323) );
  XOR3X1 U8483 ( .IN1(n3178), .IN2(DFF_1535_n1), .IN3(DFF_1507_n1), .Q(n6996)
         );
  AND2X1 U8484 ( .IN1(n6997), .IN2(n4365), .Q(WX10321) );
  XOR2X1 U8485 ( .IN1(test_so87), .IN2(n3251), .Q(n6997) );
  AND2X1 U8486 ( .IN1(n6998), .IN2(n4375), .Q(WX10319) );
  XOR2X1 U8487 ( .IN1(CRC_OUT_2_1), .IN2(n3252), .Q(n6998) );
  AND2X1 U8488 ( .IN1(n6999), .IN2(n4351), .Q(WX10317) );
  XOR2X1 U8489 ( .IN1(CRC_OUT_2_0), .IN2(n3253), .Q(n6999) );
  AND2X1 U8490 ( .IN1(n7000), .IN2(n4365), .Q(WX10315) );
  XOR2X1 U8491 ( .IN1(n3195), .IN2(CRC_OUT_2_31), .Q(n7000) );
  XOR2X1 U8492 ( .IN1(n7001), .IN2(n5511), .Q(DATA_9_9) );
  XOR3X1 U8493 ( .IN1(n3442), .IN2(n530), .IN3(n7002), .Q(n5511) );
  XNOR3X1 U8494 ( .IN1(n7265), .IN2(n3485), .IN3(n3443), .Q(n7002) );
  AND2X1 U8495 ( .IN1(TM0), .IN2(WX529), .Q(n7001) );
  XOR2X1 U8496 ( .IN1(n7003), .IN2(n5505), .Q(DATA_9_8) );
  XOR3X1 U8497 ( .IN1(n3448), .IN2(n530), .IN3(n7004), .Q(n5505) );
  XOR3X1 U8498 ( .IN1(n7266), .IN2(n3483), .IN3(WX755), .Q(n7004) );
  AND2X1 U8499 ( .IN1(TM0), .IN2(WX531), .Q(n7003) );
  XOR2X1 U8500 ( .IN1(n7005), .IN2(n5499), .Q(DATA_9_7) );
  XOR3X1 U8501 ( .IN1(n3478), .IN2(n530), .IN3(n7006), .Q(n5499) );
  XOR3X1 U8502 ( .IN1(n3482), .IN2(n3481), .IN3(WX821), .Q(n7006) );
  AND2X1 U8503 ( .IN1(TM0), .IN2(WX533), .Q(n7005) );
  XOR2X1 U8504 ( .IN1(n5493), .IN2(n7007), .Q(DATA_9_6) );
  AND2X1 U8505 ( .IN1(TM0), .IN2(WX535), .Q(n7007) );
  XOR3X1 U8506 ( .IN1(n3463), .IN2(TM0), .IN3(n7008), .Q(n5493) );
  XNOR3X1 U8507 ( .IN1(test_so5), .IN2(n3479), .IN3(n3464), .Q(n7008) );
  XOR2X1 U8508 ( .IN1(n7009), .IN2(n5487), .Q(DATA_9_5) );
  XOR3X1 U8509 ( .IN1(n3450), .IN2(n530), .IN3(n7010), .Q(n5487) );
  XOR3X1 U8510 ( .IN1(n7267), .IN2(n3477), .IN3(WX761), .Q(n7010) );
  AND2X1 U8511 ( .IN1(TM0), .IN2(WX537), .Q(n7009) );
  XOR2X1 U8512 ( .IN1(n7011), .IN2(n5481), .Q(DATA_9_4) );
  XOR3X1 U8513 ( .IN1(n3452), .IN2(n530), .IN3(n7012), .Q(n5481) );
  XOR3X1 U8514 ( .IN1(n7268), .IN2(n3475), .IN3(WX763), .Q(n7012) );
  AND2X1 U8515 ( .IN1(TM0), .IN2(WX539), .Q(n7011) );
  XOR2X1 U8516 ( .IN1(n7013), .IN2(n5674), .Q(DATA_9_31) );
  XOR3X1 U8517 ( .IN1(n3466), .IN2(n3518), .IN3(n7014), .Q(n5674) );
  XNOR3X1 U8518 ( .IN1(n7269), .IN2(n3529), .IN3(n3468), .Q(n7014) );
  AND2X1 U8519 ( .IN1(TM0), .IN2(WX485), .Q(n7013) );
  XOR2X1 U8520 ( .IN1(n7015), .IN2(n5658), .Q(DATA_9_30) );
  XOR3X1 U8521 ( .IN1(n3415), .IN2(n3516), .IN3(n7016), .Q(n5658) );
  XOR3X1 U8522 ( .IN1(n3527), .IN2(n3417), .IN3(WX775), .Q(n7016) );
  AND2X1 U8523 ( .IN1(TM0), .IN2(WX487), .Q(n7015) );
  XOR2X1 U8524 ( .IN1(n7017), .IN2(n5475), .Q(DATA_9_3) );
  XOR3X1 U8525 ( .IN1(n3418), .IN2(n530), .IN3(n7018), .Q(n5475) );
  XOR3X1 U8526 ( .IN1(n7270), .IN2(n3473), .IN3(WX765), .Q(n7018) );
  AND2X1 U8527 ( .IN1(TM0), .IN2(WX541), .Q(n7017) );
  XOR2X1 U8528 ( .IN1(n7019), .IN2(n5642), .Q(DATA_9_29) );
  XOR3X1 U8529 ( .IN1(n3422), .IN2(n3515), .IN3(n7020), .Q(n5642) );
  XOR3X1 U8530 ( .IN1(n7271), .IN2(n3525), .IN3(WX713), .Q(n7020) );
  AND2X1 U8531 ( .IN1(TM0), .IN2(WX489), .Q(n7019) );
  XOR2X1 U8532 ( .IN1(n5625), .IN2(n7021), .Q(DATA_9_28) );
  AND2X1 U8533 ( .IN1(TM0), .IN2(WX491), .Q(n7021) );
  XOR3X1 U8534 ( .IN1(n3428), .IN2(TM1), .IN3(n7022), .Q(n5625) );
  XOR3X1 U8535 ( .IN1(test_so2), .IN2(n7272), .IN3(WX779), .Q(n7022) );
  XOR2X1 U8536 ( .IN1(n7023), .IN2(n5619), .Q(DATA_9_27) );
  XOR3X1 U8537 ( .IN1(n3431), .IN2(n3514), .IN3(n7024), .Q(n5619) );
  XOR3X1 U8538 ( .IN1(n7273), .IN2(n3521), .IN3(WX717), .Q(n7024) );
  AND2X1 U8539 ( .IN1(TM0), .IN2(WX493), .Q(n7023) );
  XOR2X1 U8540 ( .IN1(n7025), .IN2(n5613), .Q(DATA_9_26) );
  XOR3X1 U8541 ( .IN1(n3433), .IN2(n3518), .IN3(n7026), .Q(n5613) );
  XOR3X1 U8542 ( .IN1(n7274), .IN2(n3519), .IN3(WX719), .Q(n7026) );
  AND2X1 U8543 ( .IN1(TM0), .IN2(WX495), .Q(n7025) );
  XOR2X1 U8544 ( .IN1(n7027), .IN2(n5607), .Q(DATA_9_25) );
  XOR3X1 U8545 ( .IN1(n3438), .IN2(n3516), .IN3(n7028), .Q(n5607) );
  XOR3X1 U8546 ( .IN1(n7275), .IN2(n3517), .IN3(WX721), .Q(n7028) );
  AND2X1 U8547 ( .IN1(TM0), .IN2(WX497), .Q(n7027) );
  XOR2X1 U8548 ( .IN1(n5601), .IN2(n7029), .Q(DATA_9_24) );
  AND2X1 U8549 ( .IN1(TM0), .IN2(WX499), .Q(n7029) );
  XOR3X1 U8550 ( .IN1(n3444), .IN2(TM1), .IN3(n7030), .Q(n5601) );
  XOR3X1 U8551 ( .IN1(test_so4), .IN2(n7276), .IN3(WX659), .Q(n7030) );
  XOR2X1 U8552 ( .IN1(n7031), .IN2(n5595), .Q(DATA_9_23) );
  XOR3X1 U8553 ( .IN1(n3445), .IN2(n3515), .IN3(n7032), .Q(n5595) );
  XOR3X1 U8554 ( .IN1(n7277), .IN2(n3513), .IN3(WX725), .Q(n7032) );
  AND2X1 U8555 ( .IN1(TM0), .IN2(WX501), .Q(n7031) );
  XOR2X1 U8556 ( .IN1(n7033), .IN2(n5589), .Q(DATA_9_22) );
  XOR3X1 U8557 ( .IN1(n3454), .IN2(n3514), .IN3(n7034), .Q(n5589) );
  XOR3X1 U8558 ( .IN1(n3511), .IN2(n3456), .IN3(WX791), .Q(n7034) );
  AND2X1 U8559 ( .IN1(TM0), .IN2(WX503), .Q(n7033) );
  XOR2X1 U8560 ( .IN1(n7035), .IN2(n5583), .Q(DATA_9_21) );
  XOR3X1 U8561 ( .IN1(n3460), .IN2(n3518), .IN3(n7036), .Q(n5583) );
  XOR3X1 U8562 ( .IN1(n3509), .IN2(n3462), .IN3(WX793), .Q(n7036) );
  AND2X1 U8563 ( .IN1(TM0), .IN2(WX505), .Q(n7035) );
  XOR2X1 U8564 ( .IN1(n5577), .IN2(n7037), .Q(DATA_9_20) );
  AND2X1 U8565 ( .IN1(TM0), .IN2(WX507), .Q(n7037) );
  XOR3X1 U8566 ( .IN1(n3465), .IN2(TM1), .IN3(n7038), .Q(n5577) );
  XOR3X1 U8567 ( .IN1(test_so6), .IN2(n7278), .IN3(WX667), .Q(n7038) );
  XOR2X1 U8568 ( .IN1(n5469), .IN2(n7039), .Q(DATA_9_2) );
  AND2X1 U8569 ( .IN1(TM0), .IN2(WX543), .Q(n7039) );
  XOR3X1 U8570 ( .IN1(n3471), .IN2(TM0), .IN3(n7040), .Q(n5469) );
  XOR3X1 U8571 ( .IN1(test_so7), .IN2(n3476), .IN3(WX767), .Q(n7040) );
  XOR2X1 U8572 ( .IN1(n7041), .IN2(n5571), .Q(DATA_9_19) );
  XOR3X1 U8573 ( .IN1(n3420), .IN2(n3516), .IN3(n7042), .Q(n5571) );
  XOR3X1 U8574 ( .IN1(n7279), .IN2(n3505), .IN3(WX733), .Q(n7042) );
  AND2X1 U8575 ( .IN1(TM0), .IN2(WX509), .Q(n7041) );
  XOR2X1 U8576 ( .IN1(n7043), .IN2(n5565), .Q(DATA_9_18) );
  XOR3X1 U8577 ( .IN1(n3429), .IN2(n3515), .IN3(n7044), .Q(n5565) );
  XOR3X1 U8578 ( .IN1(n7280), .IN2(n3503), .IN3(WX735), .Q(n7044) );
  AND2X1 U8579 ( .IN1(TM0), .IN2(WX511), .Q(n7043) );
  XOR2X1 U8580 ( .IN1(n7045), .IN2(n5559), .Q(DATA_9_17) );
  XOR3X1 U8581 ( .IN1(n3436), .IN2(n3514), .IN3(n7046), .Q(n5559) );
  XOR3X1 U8582 ( .IN1(n7281), .IN2(n3501), .IN3(WX737), .Q(n7046) );
  AND2X1 U8583 ( .IN1(TM0), .IN2(WX513), .Q(n7045) );
  XOR2X1 U8584 ( .IN1(n5553), .IN2(n7047), .Q(DATA_9_16) );
  AND2X1 U8585 ( .IN1(TM0), .IN2(WX515), .Q(n7047) );
  XOR3X1 U8586 ( .IN1(n3447), .IN2(TM1), .IN3(n7048), .Q(n5553) );
  XOR3X1 U8587 ( .IN1(test_so8), .IN2(n7282), .IN3(WX675), .Q(n7048) );
  XOR2X1 U8588 ( .IN1(n7049), .IN2(n5547), .Q(DATA_9_15) );
  XOR3X1 U8589 ( .IN1(n3457), .IN2(n530), .IN3(n7050), .Q(n5547) );
  XOR3X1 U8590 ( .IN1(n3497), .IN2(n3459), .IN3(WX805), .Q(n7050) );
  AND2X1 U8591 ( .IN1(TM0), .IN2(WX517), .Q(n7049) );
  XOR2X1 U8592 ( .IN1(n7051), .IN2(n5541), .Q(DATA_9_14) );
  XOR3X1 U8593 ( .IN1(n3470), .IN2(n530), .IN3(n7052), .Q(n5541) );
  XOR3X1 U8594 ( .IN1(n7283), .IN2(n3495), .IN3(WX743), .Q(n7052) );
  AND2X1 U8595 ( .IN1(test_so1), .IN2(TM0), .Q(n7051) );
  XOR2X1 U8596 ( .IN1(n7053), .IN2(n5535), .Q(DATA_9_13) );
  XOR3X1 U8597 ( .IN1(n3424), .IN2(n530), .IN3(n7054), .Q(n5535) );
  XOR3X1 U8598 ( .IN1(n7284), .IN2(n3493), .IN3(WX745), .Q(n7054) );
  AND2X1 U8599 ( .IN1(TM0), .IN2(WX521), .Q(n7053) );
  XOR2X1 U8600 ( .IN1(n7055), .IN2(n5529), .Q(DATA_9_12) );
  XOR3X1 U8601 ( .IN1(n3440), .IN2(n530), .IN3(n7056), .Q(n5529) );
  XOR3X1 U8602 ( .IN1(n7285), .IN2(n3491), .IN3(WX747), .Q(n7056) );
  AND2X1 U8603 ( .IN1(TM0), .IN2(WX523), .Q(n7055) );
  XOR2X1 U8604 ( .IN1(n7057), .IN2(n5523), .Q(DATA_9_11) );
  XOR3X1 U8605 ( .IN1(n3484), .IN2(n530), .IN3(n7058), .Q(n5523) );
  XOR3X1 U8606 ( .IN1(n7286), .IN2(n3489), .IN3(WX749), .Q(n7058) );
  AND2X1 U8607 ( .IN1(TM0), .IN2(WX525), .Q(n7057) );
  XOR2X1 U8608 ( .IN1(n5517), .IN2(n7059), .Q(DATA_9_10) );
  AND2X1 U8609 ( .IN1(TM0), .IN2(WX527), .Q(n7059) );
  XOR3X1 U8610 ( .IN1(n3435), .IN2(TM0), .IN3(n7060), .Q(n5517) );
  XOR3X1 U8611 ( .IN1(test_so3), .IN2(n7287), .IN3(WX815), .Q(n7060) );
  XOR2X1 U8612 ( .IN1(n7061), .IN2(n5463), .Q(DATA_9_1) );
  XOR3X1 U8613 ( .IN1(n3426), .IN2(n530), .IN3(n7062), .Q(n5463) );
  XOR3X1 U8614 ( .IN1(n7288), .IN2(n3469), .IN3(WX769), .Q(n7062) );
  AND2X1 U8615 ( .IN1(TM0), .IN2(WX545), .Q(n7061) );
  XOR2X1 U8616 ( .IN1(n7063), .IN2(n5457), .Q(DATA_9_0) );
  XOR3X1 U8617 ( .IN1(n3467), .IN2(n530), .IN3(n7064), .Q(n5457) );
  XOR3X1 U8618 ( .IN1(n3490), .IN2(n3488), .IN3(WX771), .Q(n7064) );
  INVX0 U8619 ( .INP(TM0), .ZN(n530) );
  AND2X1 U8620 ( .IN1(TM0), .IN2(WX547), .Q(n7063) );
  AND2X1 U3558_U2 ( .IN1(n3584), .IN2(U3558_n1), .Q(n2245) );
  INVX0 U3558_U1 ( .INP(n4447), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(TM0), .ZN(U3871_n1) );
  AND2X1 U3871_U1 ( .IN1(n3278), .IN2(U3871_n1), .Q(n2153) );
  INVX0 U3991_U2 ( .INP(n530), .ZN(U3991_n1) );
  AND2X1 U3991_U1 ( .IN1(n3278), .IN2(U3991_n1), .Q(n2152) );
  AND2X1 U5716_U2 ( .IN1(WX547), .IN2(U5716_n1), .Q(WX544) );
  INVX0 U5716_U1 ( .INP(n4451), .ZN(U5716_n1) );
  AND2X1 U5717_U2 ( .IN1(WX545), .IN2(U5717_n1), .Q(WX542) );
  INVX0 U5717_U1 ( .INP(n4436), .ZN(U5717_n1) );
  AND2X1 U5718_U2 ( .IN1(WX543), .IN2(U5718_n1), .Q(WX540) );
  INVX0 U5718_U1 ( .INP(n4471), .ZN(U5718_n1) );
  AND2X1 U5719_U2 ( .IN1(WX541), .IN2(U5719_n1), .Q(WX538) );
  INVX0 U5719_U1 ( .INP(n4466), .ZN(U5719_n1) );
  AND2X1 U5720_U2 ( .IN1(WX539), .IN2(U5720_n1), .Q(WX536) );
  INVX0 U5720_U1 ( .INP(n4461), .ZN(U5720_n1) );
  AND2X1 U5721_U2 ( .IN1(WX537), .IN2(U5721_n1), .Q(WX534) );
  INVX0 U5721_U1 ( .INP(n4461), .ZN(U5721_n1) );
  AND2X1 U5722_U2 ( .IN1(WX535), .IN2(U5722_n1), .Q(WX532) );
  INVX0 U5722_U1 ( .INP(n4461), .ZN(U5722_n1) );
  AND2X1 U5723_U2 ( .IN1(WX533), .IN2(U5723_n1), .Q(WX530) );
  INVX0 U5723_U1 ( .INP(n4461), .ZN(U5723_n1) );
  AND2X1 U5724_U2 ( .IN1(WX531), .IN2(U5724_n1), .Q(WX528) );
  INVX0 U5724_U1 ( .INP(n4461), .ZN(U5724_n1) );
  AND2X1 U5725_U2 ( .IN1(WX529), .IN2(U5725_n1), .Q(WX526) );
  INVX0 U5725_U1 ( .INP(n4461), .ZN(U5725_n1) );
  AND2X1 U5726_U2 ( .IN1(WX527), .IN2(U5726_n1), .Q(WX524) );
  INVX0 U5726_U1 ( .INP(n4461), .ZN(U5726_n1) );
  AND2X1 U5727_U2 ( .IN1(WX525), .IN2(U5727_n1), .Q(WX522) );
  INVX0 U5727_U1 ( .INP(n4462), .ZN(U5727_n1) );
  AND2X1 U5728_U2 ( .IN1(WX523), .IN2(U5728_n1), .Q(WX520) );
  INVX0 U5728_U1 ( .INP(n4462), .ZN(U5728_n1) );
  AND2X1 U5729_U2 ( .IN1(WX521), .IN2(U5729_n1), .Q(WX518) );
  INVX0 U5729_U1 ( .INP(n4462), .ZN(U5729_n1) );
  AND2X1 U5730_U2 ( .IN1(test_so1), .IN2(U5730_n1), .Q(WX516) );
  INVX0 U5730_U1 ( .INP(n4462), .ZN(U5730_n1) );
  AND2X1 U5731_U2 ( .IN1(WX517), .IN2(U5731_n1), .Q(WX514) );
  INVX0 U5731_U1 ( .INP(n4462), .ZN(U5731_n1) );
  AND2X1 U5732_U2 ( .IN1(WX515), .IN2(U5732_n1), .Q(WX512) );
  INVX0 U5732_U1 ( .INP(n4462), .ZN(U5732_n1) );
  AND2X1 U5733_U2 ( .IN1(WX513), .IN2(U5733_n1), .Q(WX510) );
  INVX0 U5733_U1 ( .INP(n4462), .ZN(U5733_n1) );
  AND2X1 U5734_U2 ( .IN1(WX511), .IN2(U5734_n1), .Q(WX508) );
  INVX0 U5734_U1 ( .INP(n4462), .ZN(U5734_n1) );
  AND2X1 U5735_U2 ( .IN1(WX509), .IN2(U5735_n1), .Q(WX506) );
  INVX0 U5735_U1 ( .INP(n4462), .ZN(U5735_n1) );
  AND2X1 U5736_U2 ( .IN1(WX507), .IN2(U5736_n1), .Q(WX504) );
  INVX0 U5736_U1 ( .INP(n4462), .ZN(U5736_n1) );
  AND2X1 U5737_U2 ( .IN1(WX505), .IN2(U5737_n1), .Q(WX502) );
  INVX0 U5737_U1 ( .INP(n4462), .ZN(U5737_n1) );
  AND2X1 U5738_U2 ( .IN1(WX503), .IN2(U5738_n1), .Q(WX500) );
  INVX0 U5738_U1 ( .INP(n4462), .ZN(U5738_n1) );
  AND2X1 U5739_U2 ( .IN1(WX501), .IN2(U5739_n1), .Q(WX498) );
  INVX0 U5739_U1 ( .INP(n4462), .ZN(U5739_n1) );
  AND2X1 U5740_U2 ( .IN1(WX499), .IN2(U5740_n1), .Q(WX496) );
  INVX0 U5740_U1 ( .INP(n4462), .ZN(U5740_n1) );
  AND2X1 U5741_U2 ( .IN1(WX497), .IN2(U5741_n1), .Q(WX494) );
  INVX0 U5741_U1 ( .INP(n4463), .ZN(U5741_n1) );
  AND2X1 U5742_U2 ( .IN1(WX495), .IN2(U5742_n1), .Q(WX492) );
  INVX0 U5742_U1 ( .INP(n4463), .ZN(U5742_n1) );
  AND2X1 U5743_U2 ( .IN1(WX493), .IN2(U5743_n1), .Q(WX490) );
  INVX0 U5743_U1 ( .INP(n4463), .ZN(U5743_n1) );
  AND2X1 U5744_U2 ( .IN1(WX491), .IN2(U5744_n1), .Q(WX488) );
  INVX0 U5744_U1 ( .INP(n4463), .ZN(U5744_n1) );
  AND2X1 U5745_U2 ( .IN1(WX489), .IN2(U5745_n1), .Q(WX486) );
  INVX0 U5745_U1 ( .INP(n4463), .ZN(U5745_n1) );
  AND2X1 U5746_U2 ( .IN1(WX487), .IN2(U5746_n1), .Q(WX484) );
  INVX0 U5746_U1 ( .INP(n4463), .ZN(U5746_n1) );
  AND2X1 U5747_U2 ( .IN1(WX5939), .IN2(U5747_n1), .Q(WX6002) );
  INVX0 U5747_U1 ( .INP(n4463), .ZN(U5747_n1) );
  AND2X1 U5748_U2 ( .IN1(test_so49), .IN2(U5748_n1), .Q(WX6000) );
  INVX0 U5748_U1 ( .INP(n4463), .ZN(U5748_n1) );
  AND2X1 U5749_U2 ( .IN1(WX5935), .IN2(U5749_n1), .Q(WX5998) );
  INVX0 U5749_U1 ( .INP(n4463), .ZN(U5749_n1) );
  AND2X1 U5750_U2 ( .IN1(WX5933), .IN2(U5750_n1), .Q(WX5996) );
  INVX0 U5750_U1 ( .INP(n4463), .ZN(U5750_n1) );
  AND2X1 U5751_U2 ( .IN1(WX5931), .IN2(U5751_n1), .Q(WX5994) );
  INVX0 U5751_U1 ( .INP(n4463), .ZN(U5751_n1) );
  AND2X1 U5752_U2 ( .IN1(WX3269), .IN2(U5752_n1), .Q(WX3332) );
  INVX0 U5752_U1 ( .INP(n4463), .ZN(U5752_n1) );
  AND2X1 U5753_U2 ( .IN1(WX3265), .IN2(U5753_n1), .Q(WX3328) );
  INVX0 U5753_U1 ( .INP(n4463), .ZN(U5753_n1) );
  AND2X1 U5754_U2 ( .IN1(WX3263), .IN2(U5754_n1), .Q(WX3326) );
  INVX0 U5754_U1 ( .INP(n4463), .ZN(U5754_n1) );
  AND2X1 U5755_U2 ( .IN1(WX11179), .IN2(U5755_n1), .Q(WX11242) );
  INVX0 U5755_U1 ( .INP(n4464), .ZN(U5755_n1) );
  AND2X1 U5756_U2 ( .IN1(WX11177), .IN2(U5756_n1), .Q(WX11240) );
  INVX0 U5756_U1 ( .INP(n4464), .ZN(U5756_n1) );
  AND2X1 U5757_U2 ( .IN1(WX11175), .IN2(U5757_n1), .Q(WX11238) );
  INVX0 U5757_U1 ( .INP(n4464), .ZN(U5757_n1) );
  AND2X1 U5758_U2 ( .IN1(WX11173), .IN2(U5758_n1), .Q(WX11236) );
  INVX0 U5758_U1 ( .INP(n4464), .ZN(U5758_n1) );
  AND2X1 U5759_U2 ( .IN1(test_so96), .IN2(U5759_n1), .Q(WX11234) );
  INVX0 U5759_U1 ( .INP(n4464), .ZN(U5759_n1) );
  AND2X1 U5760_U2 ( .IN1(WX11169), .IN2(U5760_n1), .Q(WX11232) );
  INVX0 U5760_U1 ( .INP(n4464), .ZN(U5760_n1) );
  AND2X1 U5761_U2 ( .IN1(WX11167), .IN2(U5761_n1), .Q(WX11230) );
  INVX0 U5761_U1 ( .INP(n4464), .ZN(U5761_n1) );
  AND2X1 U5762_U2 ( .IN1(WX11165), .IN2(U5762_n1), .Q(WX11228) );
  INVX0 U5762_U1 ( .INP(n4464), .ZN(U5762_n1) );
  AND2X1 U5763_U2 ( .IN1(WX11163), .IN2(U5763_n1), .Q(WX11226) );
  INVX0 U5763_U1 ( .INP(n4464), .ZN(U5763_n1) );
  AND2X1 U5764_U2 ( .IN1(WX11161), .IN2(U5764_n1), .Q(WX11224) );
  INVX0 U5764_U1 ( .INP(n4464), .ZN(U5764_n1) );
  AND2X1 U5765_U2 ( .IN1(WX11159), .IN2(U5765_n1), .Q(WX11222) );
  INVX0 U5765_U1 ( .INP(n4464), .ZN(U5765_n1) );
  AND2X1 U5766_U2 ( .IN1(WX11157), .IN2(U5766_n1), .Q(WX11220) );
  INVX0 U5766_U1 ( .INP(n4464), .ZN(U5766_n1) );
  AND2X1 U5767_U2 ( .IN1(WX11155), .IN2(U5767_n1), .Q(WX11218) );
  INVX0 U5767_U1 ( .INP(n4464), .ZN(U5767_n1) );
  AND2X1 U5768_U2 ( .IN1(WX11153), .IN2(U5768_n1), .Q(WX11216) );
  INVX0 U5768_U1 ( .INP(n4464), .ZN(U5768_n1) );
  AND2X1 U5769_U2 ( .IN1(WX11151), .IN2(U5769_n1), .Q(WX11214) );
  INVX0 U5769_U1 ( .INP(n4465), .ZN(U5769_n1) );
  AND2X1 U5770_U2 ( .IN1(WX11149), .IN2(U5770_n1), .Q(WX11212) );
  INVX0 U5770_U1 ( .INP(n4465), .ZN(U5770_n1) );
  AND2X1 U5771_U2 ( .IN1(WX11147), .IN2(U5771_n1), .Q(WX11210) );
  INVX0 U5771_U1 ( .INP(n4465), .ZN(U5771_n1) );
  AND2X1 U5772_U2 ( .IN1(WX11145), .IN2(U5772_n1), .Q(WX11208) );
  INVX0 U5772_U1 ( .INP(n4465), .ZN(U5772_n1) );
  AND2X1 U5773_U2 ( .IN1(WX11143), .IN2(U5773_n1), .Q(WX11206) );
  INVX0 U5773_U1 ( .INP(n4465), .ZN(U5773_n1) );
  AND2X1 U5774_U2 ( .IN1(WX11141), .IN2(U5774_n1), .Q(WX11204) );
  INVX0 U5774_U1 ( .INP(n4465), .ZN(U5774_n1) );
  AND2X1 U5775_U2 ( .IN1(WX11139), .IN2(U5775_n1), .Q(WX11202) );
  INVX0 U5775_U1 ( .INP(n4465), .ZN(U5775_n1) );
  AND2X1 U5776_U2 ( .IN1(test_so95), .IN2(U5776_n1), .Q(WX11200) );
  INVX0 U5776_U1 ( .INP(n4465), .ZN(U5776_n1) );
  AND2X1 U5777_U2 ( .IN1(WX11135), .IN2(U5777_n1), .Q(WX11198) );
  INVX0 U5777_U1 ( .INP(n4465), .ZN(U5777_n1) );
  AND2X1 U5778_U2 ( .IN1(WX11133), .IN2(U5778_n1), .Q(WX11196) );
  INVX0 U5778_U1 ( .INP(n4465), .ZN(U5778_n1) );
  AND2X1 U5779_U2 ( .IN1(WX11131), .IN2(U5779_n1), .Q(WX11194) );
  INVX0 U5779_U1 ( .INP(n4465), .ZN(U5779_n1) );
  AND2X1 U5780_U2 ( .IN1(WX11129), .IN2(U5780_n1), .Q(WX11192) );
  INVX0 U5780_U1 ( .INP(n4465), .ZN(U5780_n1) );
  AND2X1 U5781_U2 ( .IN1(WX11127), .IN2(U5781_n1), .Q(WX11190) );
  INVX0 U5781_U1 ( .INP(n4465), .ZN(U5781_n1) );
  AND2X1 U5782_U2 ( .IN1(WX11125), .IN2(U5782_n1), .Q(WX11188) );
  INVX0 U5782_U1 ( .INP(n4465), .ZN(U5782_n1) );
  AND2X1 U5783_U2 ( .IN1(WX11123), .IN2(U5783_n1), .Q(WX11186) );
  INVX0 U5783_U1 ( .INP(n4466), .ZN(U5783_n1) );
  AND2X1 U5784_U2 ( .IN1(WX11121), .IN2(U5784_n1), .Q(WX11184) );
  INVX0 U5784_U1 ( .INP(n4466), .ZN(U5784_n1) );
  AND2X1 U5785_U2 ( .IN1(WX11119), .IN2(U5785_n1), .Q(WX11182) );
  INVX0 U5785_U1 ( .INP(n4466), .ZN(U5785_n1) );
  AND2X1 U5786_U2 ( .IN1(WX11117), .IN2(U5786_n1), .Q(WX11180) );
  INVX0 U5786_U1 ( .INP(n4466), .ZN(U5786_n1) );
  AND2X1 U5787_U2 ( .IN1(WX11115), .IN2(U5787_n1), .Q(WX11178) );
  INVX0 U5787_U1 ( .INP(n4466), .ZN(U5787_n1) );
  AND2X1 U5788_U2 ( .IN1(WX11113), .IN2(U5788_n1), .Q(WX11176) );
  INVX0 U5788_U1 ( .INP(n4466), .ZN(U5788_n1) );
  AND2X1 U5789_U2 ( .IN1(WX11111), .IN2(U5789_n1), .Q(WX11174) );
  INVX0 U5789_U1 ( .INP(n4466), .ZN(U5789_n1) );
  AND2X1 U5790_U2 ( .IN1(WX11109), .IN2(U5790_n1), .Q(WX11172) );
  INVX0 U5790_U1 ( .INP(n4466), .ZN(U5790_n1) );
  AND2X1 U5791_U2 ( .IN1(WX11107), .IN2(U5791_n1), .Q(WX11170) );
  INVX0 U5791_U1 ( .INP(n4466), .ZN(U5791_n1) );
  AND2X1 U5792_U2 ( .IN1(WX11105), .IN2(U5792_n1), .Q(WX11168) );
  INVX0 U5792_U1 ( .INP(n4466), .ZN(U5792_n1) );
  AND2X1 U5793_U2 ( .IN1(test_so94), .IN2(U5793_n1), .Q(WX11166) );
  INVX0 U5793_U1 ( .INP(n4466), .ZN(U5793_n1) );
  AND2X1 U5794_U2 ( .IN1(WX11101), .IN2(U5794_n1), .Q(WX11164) );
  INVX0 U5794_U1 ( .INP(n4466), .ZN(U5794_n1) );
  AND2X1 U5795_U2 ( .IN1(WX11099), .IN2(U5795_n1), .Q(WX11162) );
  INVX0 U5795_U1 ( .INP(n4466), .ZN(U5795_n1) );
  AND2X1 U5796_U2 ( .IN1(WX11097), .IN2(U5796_n1), .Q(WX11160) );
  INVX0 U5796_U1 ( .INP(n4467), .ZN(U5796_n1) );
  AND2X1 U5797_U2 ( .IN1(WX11095), .IN2(U5797_n1), .Q(WX11158) );
  INVX0 U5797_U1 ( .INP(n4467), .ZN(U5797_n1) );
  AND2X1 U5798_U2 ( .IN1(WX11093), .IN2(U5798_n1), .Q(WX11156) );
  INVX0 U5798_U1 ( .INP(n4467), .ZN(U5798_n1) );
  AND2X1 U5799_U2 ( .IN1(WX11091), .IN2(U5799_n1), .Q(WX11154) );
  INVX0 U5799_U1 ( .INP(n4467), .ZN(U5799_n1) );
  AND2X1 U5800_U2 ( .IN1(WX11089), .IN2(U5800_n1), .Q(WX11152) );
  INVX0 U5800_U1 ( .INP(n4467), .ZN(U5800_n1) );
  AND2X1 U5801_U2 ( .IN1(WX11087), .IN2(U5801_n1), .Q(WX11150) );
  INVX0 U5801_U1 ( .INP(n4467), .ZN(U5801_n1) );
  AND2X1 U5802_U2 ( .IN1(WX11085), .IN2(U5802_n1), .Q(WX11148) );
  INVX0 U5802_U1 ( .INP(n4467), .ZN(U5802_n1) );
  AND2X1 U5803_U2 ( .IN1(WX11083), .IN2(U5803_n1), .Q(WX11146) );
  INVX0 U5803_U1 ( .INP(n4467), .ZN(U5803_n1) );
  AND2X1 U5804_U2 ( .IN1(WX11081), .IN2(U5804_n1), .Q(WX11144) );
  INVX0 U5804_U1 ( .INP(n4467), .ZN(U5804_n1) );
  AND2X1 U5805_U2 ( .IN1(WX11079), .IN2(U5805_n1), .Q(WX11142) );
  INVX0 U5805_U1 ( .INP(n4467), .ZN(U5805_n1) );
  AND2X1 U5806_U2 ( .IN1(WX11077), .IN2(U5806_n1), .Q(WX11140) );
  INVX0 U5806_U1 ( .INP(n4467), .ZN(U5806_n1) );
  AND2X1 U5807_U2 ( .IN1(WX11075), .IN2(U5807_n1), .Q(WX11138) );
  INVX0 U5807_U1 ( .INP(n4467), .ZN(U5807_n1) );
  AND2X1 U5808_U2 ( .IN1(WX11073), .IN2(U5808_n1), .Q(WX11136) );
  INVX0 U5808_U1 ( .INP(n4467), .ZN(U5808_n1) );
  AND2X1 U5809_U2 ( .IN1(WX11071), .IN2(U5809_n1), .Q(WX11134) );
  INVX0 U5809_U1 ( .INP(n4467), .ZN(U5809_n1) );
  AND2X1 U5810_U2 ( .IN1(test_so93), .IN2(U5810_n1), .Q(WX11132) );
  INVX0 U5810_U1 ( .INP(n4468), .ZN(U5810_n1) );
  AND2X1 U5811_U2 ( .IN1(WX11067), .IN2(U5811_n1), .Q(WX11130) );
  INVX0 U5811_U1 ( .INP(n4468), .ZN(U5811_n1) );
  AND2X1 U5812_U2 ( .IN1(WX11065), .IN2(U5812_n1), .Q(WX11128) );
  INVX0 U5812_U1 ( .INP(n4468), .ZN(U5812_n1) );
  AND2X1 U5813_U2 ( .IN1(WX11063), .IN2(U5813_n1), .Q(WX11126) );
  INVX0 U5813_U1 ( .INP(n4468), .ZN(U5813_n1) );
  AND2X1 U5814_U2 ( .IN1(WX11061), .IN2(U5814_n1), .Q(WX11124) );
  INVX0 U5814_U1 ( .INP(n4468), .ZN(U5814_n1) );
  AND2X1 U5815_U2 ( .IN1(WX11059), .IN2(U5815_n1), .Q(WX11122) );
  INVX0 U5815_U1 ( .INP(n4468), .ZN(U5815_n1) );
  AND2X1 U5816_U2 ( .IN1(WX11057), .IN2(U5816_n1), .Q(WX11120) );
  INVX0 U5816_U1 ( .INP(n4468), .ZN(U5816_n1) );
  AND2X1 U5817_U2 ( .IN1(WX11055), .IN2(U5817_n1), .Q(WX11118) );
  INVX0 U5817_U1 ( .INP(n4468), .ZN(U5817_n1) );
  AND2X1 U5818_U2 ( .IN1(WX11053), .IN2(U5818_n1), .Q(WX11116) );
  INVX0 U5818_U1 ( .INP(n4468), .ZN(U5818_n1) );
  AND2X1 U5819_U2 ( .IN1(WX11051), .IN2(U5819_n1), .Q(WX11114) );
  INVX0 U5819_U1 ( .INP(n4468), .ZN(U5819_n1) );
  AND2X1 U5820_U2 ( .IN1(WX11049), .IN2(U5820_n1), .Q(WX11112) );
  INVX0 U5820_U1 ( .INP(n4468), .ZN(U5820_n1) );
  AND2X1 U5821_U2 ( .IN1(WX11047), .IN2(U5821_n1), .Q(WX11110) );
  INVX0 U5821_U1 ( .INP(n4468), .ZN(U5821_n1) );
  AND2X1 U5822_U2 ( .IN1(WX11045), .IN2(U5822_n1), .Q(WX11108) );
  INVX0 U5822_U1 ( .INP(n4468), .ZN(U5822_n1) );
  AND2X1 U5823_U2 ( .IN1(WX11043), .IN2(U5823_n1), .Q(WX11106) );
  INVX0 U5823_U1 ( .INP(n4468), .ZN(U5823_n1) );
  AND2X1 U5824_U2 ( .IN1(WX11041), .IN2(U5824_n1), .Q(WX11104) );
  INVX0 U5824_U1 ( .INP(n4469), .ZN(U5824_n1) );
  AND2X1 U5825_U2 ( .IN1(WX11039), .IN2(U5825_n1), .Q(WX11102) );
  INVX0 U5825_U1 ( .INP(n4469), .ZN(U5825_n1) );
  AND2X1 U5826_U2 ( .IN1(WX11037), .IN2(U5826_n1), .Q(WX11100) );
  INVX0 U5826_U1 ( .INP(n4469), .ZN(U5826_n1) );
  AND2X1 U5827_U2 ( .IN1(test_so92), .IN2(U5827_n1), .Q(WX11098) );
  INVX0 U5827_U1 ( .INP(n4469), .ZN(U5827_n1) );
  AND2X1 U5828_U2 ( .IN1(WX11033), .IN2(U5828_n1), .Q(WX11096) );
  INVX0 U5828_U1 ( .INP(n4469), .ZN(U5828_n1) );
  AND2X1 U5829_U2 ( .IN1(WX11031), .IN2(U5829_n1), .Q(WX11094) );
  INVX0 U5829_U1 ( .INP(n4469), .ZN(U5829_n1) );
  AND2X1 U5830_U2 ( .IN1(WX11029), .IN2(U5830_n1), .Q(WX11092) );
  INVX0 U5830_U1 ( .INP(n4469), .ZN(U5830_n1) );
  AND2X1 U5831_U2 ( .IN1(WX11027), .IN2(U5831_n1), .Q(WX11090) );
  INVX0 U5831_U1 ( .INP(n4469), .ZN(U5831_n1) );
  AND2X1 U5832_U2 ( .IN1(WX11025), .IN2(U5832_n1), .Q(WX11088) );
  INVX0 U5832_U1 ( .INP(n4469), .ZN(U5832_n1) );
  AND2X1 U5833_U2 ( .IN1(WX11023), .IN2(U5833_n1), .Q(WX11086) );
  INVX0 U5833_U1 ( .INP(n4469), .ZN(U5833_n1) );
  AND2X1 U5834_U2 ( .IN1(WX11021), .IN2(U5834_n1), .Q(WX11084) );
  INVX0 U5834_U1 ( .INP(n4469), .ZN(U5834_n1) );
  AND2X1 U5835_U2 ( .IN1(WX9886), .IN2(U5835_n1), .Q(WX9949) );
  INVX0 U5835_U1 ( .INP(n4469), .ZN(U5835_n1) );
  AND2X1 U5836_U2 ( .IN1(WX9884), .IN2(U5836_n1), .Q(WX9947) );
  INVX0 U5836_U1 ( .INP(n4469), .ZN(U5836_n1) );
  AND2X1 U5837_U2 ( .IN1(WX9882), .IN2(U5837_n1), .Q(WX9945) );
  INVX0 U5837_U1 ( .INP(n4469), .ZN(U5837_n1) );
  AND2X1 U5838_U2 ( .IN1(WX9880), .IN2(U5838_n1), .Q(WX9943) );
  INVX0 U5838_U1 ( .INP(n4470), .ZN(U5838_n1) );
  AND2X1 U5839_U2 ( .IN1(WX9878), .IN2(U5839_n1), .Q(WX9941) );
  INVX0 U5839_U1 ( .INP(n4470), .ZN(U5839_n1) );
  AND2X1 U5840_U2 ( .IN1(WX9876), .IN2(U5840_n1), .Q(WX9939) );
  INVX0 U5840_U1 ( .INP(n4470), .ZN(U5840_n1) );
  AND2X1 U5841_U2 ( .IN1(WX9874), .IN2(U5841_n1), .Q(WX9937) );
  INVX0 U5841_U1 ( .INP(n4470), .ZN(U5841_n1) );
  AND2X1 U5842_U2 ( .IN1(WX9872), .IN2(U5842_n1), .Q(WX9935) );
  INVX0 U5842_U1 ( .INP(n4470), .ZN(U5842_n1) );
  AND2X1 U5843_U2 ( .IN1(WX9870), .IN2(U5843_n1), .Q(WX9933) );
  INVX0 U5843_U1 ( .INP(n4470), .ZN(U5843_n1) );
  AND2X1 U5844_U2 ( .IN1(WX9868), .IN2(U5844_n1), .Q(WX9931) );
  INVX0 U5844_U1 ( .INP(n4470), .ZN(U5844_n1) );
  AND2X1 U5845_U2 ( .IN1(WX9866), .IN2(U5845_n1), .Q(WX9929) );
  INVX0 U5845_U1 ( .INP(n4470), .ZN(U5845_n1) );
  AND2X1 U5846_U2 ( .IN1(WX9864), .IN2(U5846_n1), .Q(WX9927) );
  INVX0 U5846_U1 ( .INP(n4470), .ZN(U5846_n1) );
  AND2X1 U5847_U2 ( .IN1(WX9862), .IN2(U5847_n1), .Q(WX9925) );
  INVX0 U5847_U1 ( .INP(n4470), .ZN(U5847_n1) );
  AND2X1 U5848_U2 ( .IN1(WX9860), .IN2(U5848_n1), .Q(WX9923) );
  INVX0 U5848_U1 ( .INP(n4470), .ZN(U5848_n1) );
  AND2X1 U5849_U2 ( .IN1(WX9858), .IN2(U5849_n1), .Q(WX9921) );
  INVX0 U5849_U1 ( .INP(n4470), .ZN(U5849_n1) );
  AND2X1 U5850_U2 ( .IN1(WX9856), .IN2(U5850_n1), .Q(WX9919) );
  INVX0 U5850_U1 ( .INP(n4470), .ZN(U5850_n1) );
  AND2X1 U5851_U2 ( .IN1(test_so84), .IN2(U5851_n1), .Q(WX9917) );
  INVX0 U5851_U1 ( .INP(n4470), .ZN(U5851_n1) );
  AND2X1 U5852_U2 ( .IN1(WX9852), .IN2(U5852_n1), .Q(WX9915) );
  INVX0 U5852_U1 ( .INP(n4471), .ZN(U5852_n1) );
  AND2X1 U5853_U2 ( .IN1(WX9850), .IN2(U5853_n1), .Q(WX9913) );
  INVX0 U5853_U1 ( .INP(n4471), .ZN(U5853_n1) );
  AND2X1 U5854_U2 ( .IN1(WX9848), .IN2(U5854_n1), .Q(WX9911) );
  INVX0 U5854_U1 ( .INP(n4471), .ZN(U5854_n1) );
  AND2X1 U5855_U2 ( .IN1(WX9846), .IN2(U5855_n1), .Q(WX9909) );
  INVX0 U5855_U1 ( .INP(n4471), .ZN(U5855_n1) );
  AND2X1 U5856_U2 ( .IN1(WX9844), .IN2(U5856_n1), .Q(WX9907) );
  INVX0 U5856_U1 ( .INP(n4471), .ZN(U5856_n1) );
  AND2X1 U5857_U2 ( .IN1(WX9842), .IN2(U5857_n1), .Q(WX9905) );
  INVX0 U5857_U1 ( .INP(n4456), .ZN(U5857_n1) );
  AND2X1 U5858_U2 ( .IN1(WX9840), .IN2(U5858_n1), .Q(WX9903) );
  INVX0 U5858_U1 ( .INP(n4451), .ZN(U5858_n1) );
  AND2X1 U5859_U2 ( .IN1(WX9838), .IN2(U5859_n1), .Q(WX9901) );
  INVX0 U5859_U1 ( .INP(n4451), .ZN(U5859_n1) );
  AND2X1 U5860_U2 ( .IN1(WX9836), .IN2(U5860_n1), .Q(WX9899) );
  INVX0 U5860_U1 ( .INP(n4451), .ZN(U5860_n1) );
  AND2X1 U5861_U2 ( .IN1(WX9834), .IN2(U5861_n1), .Q(WX9897) );
  INVX0 U5861_U1 ( .INP(n4451), .ZN(U5861_n1) );
  AND2X1 U5862_U2 ( .IN1(WX9832), .IN2(U5862_n1), .Q(WX9895) );
  INVX0 U5862_U1 ( .INP(n4451), .ZN(U5862_n1) );
  AND2X1 U5863_U2 ( .IN1(WX9830), .IN2(U5863_n1), .Q(WX9893) );
  INVX0 U5863_U1 ( .INP(n4452), .ZN(U5863_n1) );
  AND2X1 U5864_U2 ( .IN1(WX9828), .IN2(U5864_n1), .Q(WX9891) );
  INVX0 U5864_U1 ( .INP(n4452), .ZN(U5864_n1) );
  AND2X1 U5865_U2 ( .IN1(WX9826), .IN2(U5865_n1), .Q(WX9889) );
  INVX0 U5865_U1 ( .INP(n4452), .ZN(U5865_n1) );
  AND2X1 U5866_U2 ( .IN1(WX9824), .IN2(U5866_n1), .Q(WX9887) );
  INVX0 U5866_U1 ( .INP(n4452), .ZN(U5866_n1) );
  AND2X1 U5867_U2 ( .IN1(WX9822), .IN2(U5867_n1), .Q(WX9885) );
  INVX0 U5867_U1 ( .INP(n4452), .ZN(U5867_n1) );
  AND2X1 U5868_U2 ( .IN1(test_so83), .IN2(U5868_n1), .Q(WX9883) );
  INVX0 U5868_U1 ( .INP(n4452), .ZN(U5868_n1) );
  AND2X1 U5869_U2 ( .IN1(WX9818), .IN2(U5869_n1), .Q(WX9881) );
  INVX0 U5869_U1 ( .INP(n4452), .ZN(U5869_n1) );
  AND2X1 U5870_U2 ( .IN1(WX9816), .IN2(U5870_n1), .Q(WX9879) );
  INVX0 U5870_U1 ( .INP(n4452), .ZN(U5870_n1) );
  AND2X1 U5871_U2 ( .IN1(WX9814), .IN2(U5871_n1), .Q(WX9877) );
  INVX0 U5871_U1 ( .INP(n4452), .ZN(U5871_n1) );
  AND2X1 U5872_U2 ( .IN1(WX9812), .IN2(U5872_n1), .Q(WX9875) );
  INVX0 U5872_U1 ( .INP(n4452), .ZN(U5872_n1) );
  AND2X1 U5873_U2 ( .IN1(WX9810), .IN2(U5873_n1), .Q(WX9873) );
  INVX0 U5873_U1 ( .INP(n4452), .ZN(U5873_n1) );
  AND2X1 U5874_U2 ( .IN1(WX9808), .IN2(U5874_n1), .Q(WX9871) );
  INVX0 U5874_U1 ( .INP(n4452), .ZN(U5874_n1) );
  AND2X1 U5875_U2 ( .IN1(WX9806), .IN2(U5875_n1), .Q(WX9869) );
  INVX0 U5875_U1 ( .INP(n4452), .ZN(U5875_n1) );
  AND2X1 U5876_U2 ( .IN1(WX9804), .IN2(U5876_n1), .Q(WX9867) );
  INVX0 U5876_U1 ( .INP(n4452), .ZN(U5876_n1) );
  AND2X1 U5877_U2 ( .IN1(WX9802), .IN2(U5877_n1), .Q(WX9865) );
  INVX0 U5877_U1 ( .INP(n4453), .ZN(U5877_n1) );
  AND2X1 U5878_U2 ( .IN1(WX9800), .IN2(U5878_n1), .Q(WX9863) );
  INVX0 U5878_U1 ( .INP(n4453), .ZN(U5878_n1) );
  AND2X1 U5879_U2 ( .IN1(WX9798), .IN2(U5879_n1), .Q(WX9861) );
  INVX0 U5879_U1 ( .INP(n4453), .ZN(U5879_n1) );
  AND2X1 U5880_U2 ( .IN1(WX9796), .IN2(U5880_n1), .Q(WX9859) );
  INVX0 U5880_U1 ( .INP(n4453), .ZN(U5880_n1) );
  AND2X1 U5881_U2 ( .IN1(WX9794), .IN2(U5881_n1), .Q(WX9857) );
  INVX0 U5881_U1 ( .INP(n4453), .ZN(U5881_n1) );
  AND2X1 U5882_U2 ( .IN1(WX9792), .IN2(U5882_n1), .Q(WX9855) );
  INVX0 U5882_U1 ( .INP(n4453), .ZN(U5882_n1) );
  AND2X1 U5883_U2 ( .IN1(WX9790), .IN2(U5883_n1), .Q(WX9853) );
  INVX0 U5883_U1 ( .INP(n4453), .ZN(U5883_n1) );
  AND2X1 U5884_U2 ( .IN1(WX9788), .IN2(U5884_n1), .Q(WX9851) );
  INVX0 U5884_U1 ( .INP(n4453), .ZN(U5884_n1) );
  AND2X1 U5885_U2 ( .IN1(test_so82), .IN2(U5885_n1), .Q(WX9849) );
  INVX0 U5885_U1 ( .INP(n4453), .ZN(U5885_n1) );
  AND2X1 U5886_U2 ( .IN1(WX9784), .IN2(U5886_n1), .Q(WX9847) );
  INVX0 U5886_U1 ( .INP(n4453), .ZN(U5886_n1) );
  AND2X1 U5887_U2 ( .IN1(WX9782), .IN2(U5887_n1), .Q(WX9845) );
  INVX0 U5887_U1 ( .INP(n4453), .ZN(U5887_n1) );
  AND2X1 U5888_U2 ( .IN1(WX9780), .IN2(U5888_n1), .Q(WX9843) );
  INVX0 U5888_U1 ( .INP(n4453), .ZN(U5888_n1) );
  AND2X1 U5889_U2 ( .IN1(WX9778), .IN2(U5889_n1), .Q(WX9841) );
  INVX0 U5889_U1 ( .INP(n4453), .ZN(U5889_n1) );
  AND2X1 U5890_U2 ( .IN1(WX9776), .IN2(U5890_n1), .Q(WX9839) );
  INVX0 U5890_U1 ( .INP(n4453), .ZN(U5890_n1) );
  AND2X1 U5891_U2 ( .IN1(WX9774), .IN2(U5891_n1), .Q(WX9837) );
  INVX0 U5891_U1 ( .INP(n4454), .ZN(U5891_n1) );
  AND2X1 U5892_U2 ( .IN1(WX9772), .IN2(U5892_n1), .Q(WX9835) );
  INVX0 U5892_U1 ( .INP(n4454), .ZN(U5892_n1) );
  AND2X1 U5893_U2 ( .IN1(WX9770), .IN2(U5893_n1), .Q(WX9833) );
  INVX0 U5893_U1 ( .INP(n4454), .ZN(U5893_n1) );
  AND2X1 U5894_U2 ( .IN1(WX9768), .IN2(U5894_n1), .Q(WX9831) );
  INVX0 U5894_U1 ( .INP(n4454), .ZN(U5894_n1) );
  AND2X1 U5895_U2 ( .IN1(WX9766), .IN2(U5895_n1), .Q(WX9829) );
  INVX0 U5895_U1 ( .INP(n4454), .ZN(U5895_n1) );
  AND2X1 U5896_U2 ( .IN1(WX9764), .IN2(U5896_n1), .Q(WX9827) );
  INVX0 U5896_U1 ( .INP(n4454), .ZN(U5896_n1) );
  AND2X1 U5897_U2 ( .IN1(WX9762), .IN2(U5897_n1), .Q(WX9825) );
  INVX0 U5897_U1 ( .INP(n4454), .ZN(U5897_n1) );
  AND2X1 U5898_U2 ( .IN1(WX9760), .IN2(U5898_n1), .Q(WX9823) );
  INVX0 U5898_U1 ( .INP(n4454), .ZN(U5898_n1) );
  AND2X1 U5899_U2 ( .IN1(WX9758), .IN2(U5899_n1), .Q(WX9821) );
  INVX0 U5899_U1 ( .INP(n4454), .ZN(U5899_n1) );
  AND2X1 U5900_U2 ( .IN1(WX9756), .IN2(U5900_n1), .Q(WX9819) );
  INVX0 U5900_U1 ( .INP(n4454), .ZN(U5900_n1) );
  AND2X1 U5901_U2 ( .IN1(WX9754), .IN2(U5901_n1), .Q(WX9817) );
  INVX0 U5901_U1 ( .INP(n4454), .ZN(U5901_n1) );
  AND2X1 U5902_U2 ( .IN1(test_so81), .IN2(U5902_n1), .Q(WX9815) );
  INVX0 U5902_U1 ( .INP(n4454), .ZN(U5902_n1) );
  AND2X1 U5903_U2 ( .IN1(WX9750), .IN2(U5903_n1), .Q(WX9813) );
  INVX0 U5903_U1 ( .INP(n4454), .ZN(U5903_n1) );
  AND2X1 U5904_U2 ( .IN1(WX9748), .IN2(U5904_n1), .Q(WX9811) );
  INVX0 U5904_U1 ( .INP(n4454), .ZN(U5904_n1) );
  AND2X1 U5905_U2 ( .IN1(WX9746), .IN2(U5905_n1), .Q(WX9809) );
  INVX0 U5905_U1 ( .INP(n4455), .ZN(U5905_n1) );
  AND2X1 U5906_U2 ( .IN1(WX9744), .IN2(U5906_n1), .Q(WX9807) );
  INVX0 U5906_U1 ( .INP(n4455), .ZN(U5906_n1) );
  AND2X1 U5907_U2 ( .IN1(WX9742), .IN2(U5907_n1), .Q(WX9805) );
  INVX0 U5907_U1 ( .INP(n4455), .ZN(U5907_n1) );
  AND2X1 U5908_U2 ( .IN1(WX9740), .IN2(U5908_n1), .Q(WX9803) );
  INVX0 U5908_U1 ( .INP(n4455), .ZN(U5908_n1) );
  AND2X1 U5909_U2 ( .IN1(WX9738), .IN2(U5909_n1), .Q(WX9801) );
  INVX0 U5909_U1 ( .INP(n4455), .ZN(U5909_n1) );
  AND2X1 U5910_U2 ( .IN1(WX9736), .IN2(U5910_n1), .Q(WX9799) );
  INVX0 U5910_U1 ( .INP(n4455), .ZN(U5910_n1) );
  AND2X1 U5911_U2 ( .IN1(WX9734), .IN2(U5911_n1), .Q(WX9797) );
  INVX0 U5911_U1 ( .INP(n4455), .ZN(U5911_n1) );
  AND2X1 U5912_U2 ( .IN1(WX9732), .IN2(U5912_n1), .Q(WX9795) );
  INVX0 U5912_U1 ( .INP(n4455), .ZN(U5912_n1) );
  AND2X1 U5913_U2 ( .IN1(WX9730), .IN2(U5913_n1), .Q(WX9793) );
  INVX0 U5913_U1 ( .INP(n4455), .ZN(U5913_n1) );
  AND2X1 U5914_U2 ( .IN1(WX9728), .IN2(U5914_n1), .Q(WX9791) );
  INVX0 U5914_U1 ( .INP(n4455), .ZN(U5914_n1) );
  AND2X1 U5915_U2 ( .IN1(WX8593), .IN2(U5915_n1), .Q(WX8656) );
  INVX0 U5915_U1 ( .INP(n4455), .ZN(U5915_n1) );
  AND2X1 U5916_U2 ( .IN1(WX8591), .IN2(U5916_n1), .Q(WX8654) );
  INVX0 U5916_U1 ( .INP(n4455), .ZN(U5916_n1) );
  AND2X1 U5917_U2 ( .IN1(WX8589), .IN2(U5917_n1), .Q(WX8652) );
  INVX0 U5917_U1 ( .INP(n4455), .ZN(U5917_n1) );
  AND2X1 U5918_U2 ( .IN1(WX8587), .IN2(U5918_n1), .Q(WX8650) );
  INVX0 U5918_U1 ( .INP(n4455), .ZN(U5918_n1) );
  AND2X1 U5919_U2 ( .IN1(WX8585), .IN2(U5919_n1), .Q(WX8648) );
  INVX0 U5919_U1 ( .INP(n4456), .ZN(U5919_n1) );
  AND2X1 U5920_U2 ( .IN1(WX8583), .IN2(U5920_n1), .Q(WX8646) );
  INVX0 U5920_U1 ( .INP(n4456), .ZN(U5920_n1) );
  AND2X1 U5921_U2 ( .IN1(WX8581), .IN2(U5921_n1), .Q(WX8644) );
  INVX0 U5921_U1 ( .INP(n4456), .ZN(U5921_n1) );
  AND2X1 U5922_U2 ( .IN1(WX8579), .IN2(U5922_n1), .Q(WX8642) );
  INVX0 U5922_U1 ( .INP(n4456), .ZN(U5922_n1) );
  AND2X1 U5923_U2 ( .IN1(WX8577), .IN2(U5923_n1), .Q(WX8640) );
  INVX0 U5923_U1 ( .INP(n4456), .ZN(U5923_n1) );
  AND2X1 U5924_U2 ( .IN1(WX8575), .IN2(U5924_n1), .Q(WX8638) );
  INVX0 U5924_U1 ( .INP(n4456), .ZN(U5924_n1) );
  AND2X1 U5925_U2 ( .IN1(WX8573), .IN2(U5925_n1), .Q(WX8636) );
  INVX0 U5925_U1 ( .INP(n4456), .ZN(U5925_n1) );
  AND2X1 U5926_U2 ( .IN1(test_so73), .IN2(U5926_n1), .Q(WX8634) );
  INVX0 U5926_U1 ( .INP(n4456), .ZN(U5926_n1) );
  AND2X1 U5927_U2 ( .IN1(WX8569), .IN2(U5927_n1), .Q(WX8632) );
  INVX0 U5927_U1 ( .INP(n4456), .ZN(U5927_n1) );
  AND2X1 U5928_U2 ( .IN1(WX8567), .IN2(U5928_n1), .Q(WX8630) );
  INVX0 U5928_U1 ( .INP(n4456), .ZN(U5928_n1) );
  AND2X1 U5929_U2 ( .IN1(WX8565), .IN2(U5929_n1), .Q(WX8628) );
  INVX0 U5929_U1 ( .INP(n4456), .ZN(U5929_n1) );
  AND2X1 U5930_U2 ( .IN1(WX8563), .IN2(U5930_n1), .Q(WX8626) );
  INVX0 U5930_U1 ( .INP(n4456), .ZN(U5930_n1) );
  AND2X1 U5931_U2 ( .IN1(WX8561), .IN2(U5931_n1), .Q(WX8624) );
  INVX0 U5931_U1 ( .INP(n4456), .ZN(U5931_n1) );
  AND2X1 U5932_U2 ( .IN1(WX8559), .IN2(U5932_n1), .Q(WX8622) );
  INVX0 U5932_U1 ( .INP(n4457), .ZN(U5932_n1) );
  AND2X1 U5933_U2 ( .IN1(WX8557), .IN2(U5933_n1), .Q(WX8620) );
  INVX0 U5933_U1 ( .INP(n4457), .ZN(U5933_n1) );
  AND2X1 U5934_U2 ( .IN1(WX8555), .IN2(U5934_n1), .Q(WX8618) );
  INVX0 U5934_U1 ( .INP(n4457), .ZN(U5934_n1) );
  AND2X1 U5935_U2 ( .IN1(WX8553), .IN2(U5935_n1), .Q(WX8616) );
  INVX0 U5935_U1 ( .INP(n4457), .ZN(U5935_n1) );
  AND2X1 U5936_U2 ( .IN1(WX8551), .IN2(U5936_n1), .Q(WX8614) );
  INVX0 U5936_U1 ( .INP(n4457), .ZN(U5936_n1) );
  AND2X1 U5937_U2 ( .IN1(WX8549), .IN2(U5937_n1), .Q(WX8612) );
  INVX0 U5937_U1 ( .INP(n4457), .ZN(U5937_n1) );
  AND2X1 U5938_U2 ( .IN1(WX8547), .IN2(U5938_n1), .Q(WX8610) );
  INVX0 U5938_U1 ( .INP(n4457), .ZN(U5938_n1) );
  AND2X1 U5939_U2 ( .IN1(WX8545), .IN2(U5939_n1), .Q(WX8608) );
  INVX0 U5939_U1 ( .INP(n4457), .ZN(U5939_n1) );
  AND2X1 U5940_U2 ( .IN1(WX8543), .IN2(U5940_n1), .Q(WX8606) );
  INVX0 U5940_U1 ( .INP(n4457), .ZN(U5940_n1) );
  AND2X1 U5941_U2 ( .IN1(WX8541), .IN2(U5941_n1), .Q(WX8604) );
  INVX0 U5941_U1 ( .INP(n4457), .ZN(U5941_n1) );
  AND2X1 U5942_U2 ( .IN1(WX8539), .IN2(U5942_n1), .Q(WX8602) );
  INVX0 U5942_U1 ( .INP(n4457), .ZN(U5942_n1) );
  AND2X1 U5943_U2 ( .IN1(test_so72), .IN2(U5943_n1), .Q(WX8600) );
  INVX0 U5943_U1 ( .INP(n4457), .ZN(U5943_n1) );
  AND2X1 U5944_U2 ( .IN1(WX8535), .IN2(U5944_n1), .Q(WX8598) );
  INVX0 U5944_U1 ( .INP(n4457), .ZN(U5944_n1) );
  AND2X1 U5945_U2 ( .IN1(WX8533), .IN2(U5945_n1), .Q(WX8596) );
  INVX0 U5945_U1 ( .INP(n4457), .ZN(U5945_n1) );
  AND2X1 U5946_U2 ( .IN1(WX8531), .IN2(U5946_n1), .Q(WX8594) );
  INVX0 U5946_U1 ( .INP(n4458), .ZN(U5946_n1) );
  AND2X1 U5947_U2 ( .IN1(WX8529), .IN2(U5947_n1), .Q(WX8592) );
  INVX0 U5947_U1 ( .INP(n4458), .ZN(U5947_n1) );
  AND2X1 U5948_U2 ( .IN1(WX8527), .IN2(U5948_n1), .Q(WX8590) );
  INVX0 U5948_U1 ( .INP(n4458), .ZN(U5948_n1) );
  AND2X1 U5949_U2 ( .IN1(WX8525), .IN2(U5949_n1), .Q(WX8588) );
  INVX0 U5949_U1 ( .INP(n4458), .ZN(U5949_n1) );
  AND2X1 U5950_U2 ( .IN1(WX8523), .IN2(U5950_n1), .Q(WX8586) );
  INVX0 U5950_U1 ( .INP(n4458), .ZN(U5950_n1) );
  AND2X1 U5951_U2 ( .IN1(WX8521), .IN2(U5951_n1), .Q(WX8584) );
  INVX0 U5951_U1 ( .INP(n4458), .ZN(U5951_n1) );
  AND2X1 U5952_U2 ( .IN1(WX8519), .IN2(U5952_n1), .Q(WX8582) );
  INVX0 U5952_U1 ( .INP(n4458), .ZN(U5952_n1) );
  AND2X1 U5953_U2 ( .IN1(WX8517), .IN2(U5953_n1), .Q(WX8580) );
  INVX0 U5953_U1 ( .INP(n4458), .ZN(U5953_n1) );
  AND2X1 U5954_U2 ( .IN1(WX8515), .IN2(U5954_n1), .Q(WX8578) );
  INVX0 U5954_U1 ( .INP(n4458), .ZN(U5954_n1) );
  AND2X1 U5955_U2 ( .IN1(WX8513), .IN2(U5955_n1), .Q(WX8576) );
  INVX0 U5955_U1 ( .INP(n4458), .ZN(U5955_n1) );
  AND2X1 U5956_U2 ( .IN1(WX8511), .IN2(U5956_n1), .Q(WX8574) );
  INVX0 U5956_U1 ( .INP(n4458), .ZN(U5956_n1) );
  AND2X1 U5957_U2 ( .IN1(WX8509), .IN2(U5957_n1), .Q(WX8572) );
  INVX0 U5957_U1 ( .INP(n4458), .ZN(U5957_n1) );
  AND2X1 U5958_U2 ( .IN1(WX8507), .IN2(U5958_n1), .Q(WX8570) );
  INVX0 U5958_U1 ( .INP(n4458), .ZN(U5958_n1) );
  AND2X1 U5959_U2 ( .IN1(WX8505), .IN2(U5959_n1), .Q(WX8568) );
  INVX0 U5959_U1 ( .INP(n4458), .ZN(U5959_n1) );
  AND2X1 U5960_U2 ( .IN1(test_so71), .IN2(U5960_n1), .Q(WX8566) );
  INVX0 U5960_U1 ( .INP(n4459), .ZN(U5960_n1) );
  AND2X1 U5961_U2 ( .IN1(WX8501), .IN2(U5961_n1), .Q(WX8564) );
  INVX0 U5961_U1 ( .INP(n4459), .ZN(U5961_n1) );
  AND2X1 U5962_U2 ( .IN1(WX8499), .IN2(U5962_n1), .Q(WX8562) );
  INVX0 U5962_U1 ( .INP(n4459), .ZN(U5962_n1) );
  AND2X1 U5963_U2 ( .IN1(WX8497), .IN2(U5963_n1), .Q(WX8560) );
  INVX0 U5963_U1 ( .INP(n4459), .ZN(U5963_n1) );
  AND2X1 U5964_U2 ( .IN1(WX8495), .IN2(U5964_n1), .Q(WX8558) );
  INVX0 U5964_U1 ( .INP(n4459), .ZN(U5964_n1) );
  AND2X1 U5965_U2 ( .IN1(WX8493), .IN2(U5965_n1), .Q(WX8556) );
  INVX0 U5965_U1 ( .INP(n4459), .ZN(U5965_n1) );
  AND2X1 U5966_U2 ( .IN1(WX8491), .IN2(U5966_n1), .Q(WX8554) );
  INVX0 U5966_U1 ( .INP(n4459), .ZN(U5966_n1) );
  AND2X1 U5967_U2 ( .IN1(WX8489), .IN2(U5967_n1), .Q(WX8552) );
  INVX0 U5967_U1 ( .INP(n4459), .ZN(U5967_n1) );
  AND2X1 U5968_U2 ( .IN1(WX8487), .IN2(U5968_n1), .Q(WX8550) );
  INVX0 U5968_U1 ( .INP(n4459), .ZN(U5968_n1) );
  AND2X1 U5969_U2 ( .IN1(WX8485), .IN2(U5969_n1), .Q(WX8548) );
  INVX0 U5969_U1 ( .INP(n4459), .ZN(U5969_n1) );
  AND2X1 U5970_U2 ( .IN1(WX8483), .IN2(U5970_n1), .Q(WX8546) );
  INVX0 U5970_U1 ( .INP(n4459), .ZN(U5970_n1) );
  AND2X1 U5971_U2 ( .IN1(WX8481), .IN2(U5971_n1), .Q(WX8544) );
  INVX0 U5971_U1 ( .INP(n4459), .ZN(U5971_n1) );
  AND2X1 U5972_U2 ( .IN1(WX8479), .IN2(U5972_n1), .Q(WX8542) );
  INVX0 U5972_U1 ( .INP(n4459), .ZN(U5972_n1) );
  AND2X1 U5973_U2 ( .IN1(WX8477), .IN2(U5973_n1), .Q(WX8540) );
  INVX0 U5973_U1 ( .INP(n4459), .ZN(U5973_n1) );
  AND2X1 U5974_U2 ( .IN1(WX8475), .IN2(U5974_n1), .Q(WX8538) );
  INVX0 U5974_U1 ( .INP(n4460), .ZN(U5974_n1) );
  AND2X1 U5975_U2 ( .IN1(WX8473), .IN2(U5975_n1), .Q(WX8536) );
  INVX0 U5975_U1 ( .INP(n4460), .ZN(U5975_n1) );
  AND2X1 U5976_U2 ( .IN1(WX8471), .IN2(U5976_n1), .Q(WX8534) );
  INVX0 U5976_U1 ( .INP(n4460), .ZN(U5976_n1) );
  AND2X1 U5977_U2 ( .IN1(test_so70), .IN2(U5977_n1), .Q(WX8532) );
  INVX0 U5977_U1 ( .INP(n4460), .ZN(U5977_n1) );
  AND2X1 U5978_U2 ( .IN1(WX8467), .IN2(U5978_n1), .Q(WX8530) );
  INVX0 U5978_U1 ( .INP(n4460), .ZN(U5978_n1) );
  AND2X1 U5979_U2 ( .IN1(WX8465), .IN2(U5979_n1), .Q(WX8528) );
  INVX0 U5979_U1 ( .INP(n4460), .ZN(U5979_n1) );
  AND2X1 U5980_U2 ( .IN1(WX8463), .IN2(U5980_n1), .Q(WX8526) );
  INVX0 U5980_U1 ( .INP(n4460), .ZN(U5980_n1) );
  AND2X1 U5981_U2 ( .IN1(WX8461), .IN2(U5981_n1), .Q(WX8524) );
  INVX0 U5981_U1 ( .INP(n4460), .ZN(U5981_n1) );
  AND2X1 U5982_U2 ( .IN1(WX8459), .IN2(U5982_n1), .Q(WX8522) );
  INVX0 U5982_U1 ( .INP(n4460), .ZN(U5982_n1) );
  AND2X1 U5983_U2 ( .IN1(WX8457), .IN2(U5983_n1), .Q(WX8520) );
  INVX0 U5983_U1 ( .INP(n4460), .ZN(U5983_n1) );
  AND2X1 U5984_U2 ( .IN1(WX8455), .IN2(U5984_n1), .Q(WX8518) );
  INVX0 U5984_U1 ( .INP(n4460), .ZN(U5984_n1) );
  AND2X1 U5985_U2 ( .IN1(WX8453), .IN2(U5985_n1), .Q(WX8516) );
  INVX0 U5985_U1 ( .INP(n4460), .ZN(U5985_n1) );
  AND2X1 U5986_U2 ( .IN1(WX8451), .IN2(U5986_n1), .Q(WX8514) );
  INVX0 U5986_U1 ( .INP(n4460), .ZN(U5986_n1) );
  AND2X1 U5987_U2 ( .IN1(WX8449), .IN2(U5987_n1), .Q(WX8512) );
  INVX0 U5987_U1 ( .INP(n4460), .ZN(U5987_n1) );
  AND2X1 U5988_U2 ( .IN1(WX8447), .IN2(U5988_n1), .Q(WX8510) );
  INVX0 U5988_U1 ( .INP(n4461), .ZN(U5988_n1) );
  AND2X1 U5989_U2 ( .IN1(WX8445), .IN2(U5989_n1), .Q(WX8508) );
  INVX0 U5989_U1 ( .INP(n4461), .ZN(U5989_n1) );
  AND2X1 U5990_U2 ( .IN1(WX8443), .IN2(U5990_n1), .Q(WX8506) );
  INVX0 U5990_U1 ( .INP(n4461), .ZN(U5990_n1) );
  AND2X1 U5991_U2 ( .IN1(WX8441), .IN2(U5991_n1), .Q(WX8504) );
  INVX0 U5991_U1 ( .INP(n4461), .ZN(U5991_n1) );
  AND2X1 U5992_U2 ( .IN1(WX8439), .IN2(U5992_n1), .Q(WX8502) );
  INVX0 U5992_U1 ( .INP(n4461), .ZN(U5992_n1) );
  AND2X1 U5993_U2 ( .IN1(WX8437), .IN2(U5993_n1), .Q(WX8500) );
  INVX0 U5993_U1 ( .INP(n4461), .ZN(U5993_n1) );
  AND2X1 U5994_U2 ( .IN1(test_so69), .IN2(U5994_n1), .Q(WX8498) );
  INVX0 U5994_U1 ( .INP(n4461), .ZN(U5994_n1) );
  AND2X1 U5995_U2 ( .IN1(WX7300), .IN2(U5995_n1), .Q(WX7363) );
  INVX0 U5995_U1 ( .INP(n4486), .ZN(U5995_n1) );
  AND2X1 U5996_U2 ( .IN1(WX7298), .IN2(U5996_n1), .Q(WX7361) );
  INVX0 U5996_U1 ( .INP(n4481), .ZN(U5996_n1) );
  AND2X1 U5997_U2 ( .IN1(WX7296), .IN2(U5997_n1), .Q(WX7359) );
  INVX0 U5997_U1 ( .INP(n4481), .ZN(U5997_n1) );
  AND2X1 U5998_U2 ( .IN1(WX7294), .IN2(U5998_n1), .Q(WX7357) );
  INVX0 U5998_U1 ( .INP(n4481), .ZN(U5998_n1) );
  AND2X1 U5999_U2 ( .IN1(WX7292), .IN2(U5999_n1), .Q(WX7355) );
  INVX0 U5999_U1 ( .INP(n4481), .ZN(U5999_n1) );
  AND2X1 U6000_U2 ( .IN1(WX7290), .IN2(U6000_n1), .Q(WX7353) );
  INVX0 U6000_U1 ( .INP(n4481), .ZN(U6000_n1) );
  AND2X1 U6001_U2 ( .IN1(test_so62), .IN2(U6001_n1), .Q(WX7351) );
  INVX0 U6001_U1 ( .INP(n4481), .ZN(U6001_n1) );
  AND2X1 U6002_U2 ( .IN1(WX7286), .IN2(U6002_n1), .Q(WX7349) );
  INVX0 U6002_U1 ( .INP(n4481), .ZN(U6002_n1) );
  AND2X1 U6003_U2 ( .IN1(WX7284), .IN2(U6003_n1), .Q(WX7347) );
  INVX0 U6003_U1 ( .INP(n4481), .ZN(U6003_n1) );
  AND2X1 U6004_U2 ( .IN1(WX7282), .IN2(U6004_n1), .Q(WX7345) );
  INVX0 U6004_U1 ( .INP(n4481), .ZN(U6004_n1) );
  AND2X1 U6005_U2 ( .IN1(WX7280), .IN2(U6005_n1), .Q(WX7343) );
  INVX0 U6005_U1 ( .INP(n4481), .ZN(U6005_n1) );
  AND2X1 U6006_U2 ( .IN1(WX7278), .IN2(U6006_n1), .Q(WX7341) );
  INVX0 U6006_U1 ( .INP(n4482), .ZN(U6006_n1) );
  AND2X1 U6007_U2 ( .IN1(WX7276), .IN2(U6007_n1), .Q(WX7339) );
  INVX0 U6007_U1 ( .INP(n4482), .ZN(U6007_n1) );
  AND2X1 U6008_U2 ( .IN1(WX7274), .IN2(U6008_n1), .Q(WX7337) );
  INVX0 U6008_U1 ( .INP(n4482), .ZN(U6008_n1) );
  AND2X1 U6009_U2 ( .IN1(WX7272), .IN2(U6009_n1), .Q(WX7335) );
  INVX0 U6009_U1 ( .INP(n4482), .ZN(U6009_n1) );
  AND2X1 U6010_U2 ( .IN1(WX7270), .IN2(U6010_n1), .Q(WX7333) );
  INVX0 U6010_U1 ( .INP(n4482), .ZN(U6010_n1) );
  AND2X1 U6011_U2 ( .IN1(WX7268), .IN2(U6011_n1), .Q(WX7331) );
  INVX0 U6011_U1 ( .INP(n4482), .ZN(U6011_n1) );
  AND2X1 U6012_U2 ( .IN1(WX7266), .IN2(U6012_n1), .Q(WX7329) );
  INVX0 U6012_U1 ( .INP(n4482), .ZN(U6012_n1) );
  AND2X1 U6013_U2 ( .IN1(WX7264), .IN2(U6013_n1), .Q(WX7327) );
  INVX0 U6013_U1 ( .INP(n4482), .ZN(U6013_n1) );
  AND2X1 U6014_U2 ( .IN1(WX7262), .IN2(U6014_n1), .Q(WX7325) );
  INVX0 U6014_U1 ( .INP(n4482), .ZN(U6014_n1) );
  AND2X1 U6015_U2 ( .IN1(WX7260), .IN2(U6015_n1), .Q(WX7323) );
  INVX0 U6015_U1 ( .INP(n4482), .ZN(U6015_n1) );
  AND2X1 U6016_U2 ( .IN1(WX7258), .IN2(U6016_n1), .Q(WX7321) );
  INVX0 U6016_U1 ( .INP(n4482), .ZN(U6016_n1) );
  AND2X1 U6017_U2 ( .IN1(WX7256), .IN2(U6017_n1), .Q(WX7319) );
  INVX0 U6017_U1 ( .INP(n4482), .ZN(U6017_n1) );
  AND2X1 U6018_U2 ( .IN1(test_so61), .IN2(U6018_n1), .Q(WX7317) );
  INVX0 U6018_U1 ( .INP(n4482), .ZN(U6018_n1) );
  AND2X1 U6019_U2 ( .IN1(WX7252), .IN2(U6019_n1), .Q(WX7315) );
  INVX0 U6019_U1 ( .INP(n4482), .ZN(U6019_n1) );
  AND2X1 U6020_U2 ( .IN1(WX7250), .IN2(U6020_n1), .Q(WX7313) );
  INVX0 U6020_U1 ( .INP(n4483), .ZN(U6020_n1) );
  AND2X1 U6021_U2 ( .IN1(WX7248), .IN2(U6021_n1), .Q(WX7311) );
  INVX0 U6021_U1 ( .INP(n4483), .ZN(U6021_n1) );
  AND2X1 U6022_U2 ( .IN1(WX7246), .IN2(U6022_n1), .Q(WX7309) );
  INVX0 U6022_U1 ( .INP(n4483), .ZN(U6022_n1) );
  AND2X1 U6023_U2 ( .IN1(WX7244), .IN2(U6023_n1), .Q(WX7307) );
  INVX0 U6023_U1 ( .INP(n4483), .ZN(U6023_n1) );
  AND2X1 U6024_U2 ( .IN1(WX7242), .IN2(U6024_n1), .Q(WX7305) );
  INVX0 U6024_U1 ( .INP(n4483), .ZN(U6024_n1) );
  AND2X1 U6025_U2 ( .IN1(WX7240), .IN2(U6025_n1), .Q(WX7303) );
  INVX0 U6025_U1 ( .INP(n4483), .ZN(U6025_n1) );
  AND2X1 U6026_U2 ( .IN1(WX7238), .IN2(U6026_n1), .Q(WX7301) );
  INVX0 U6026_U1 ( .INP(n4483), .ZN(U6026_n1) );
  AND2X1 U6027_U2 ( .IN1(WX7236), .IN2(U6027_n1), .Q(WX7299) );
  INVX0 U6027_U1 ( .INP(n4483), .ZN(U6027_n1) );
  AND2X1 U6028_U2 ( .IN1(WX7234), .IN2(U6028_n1), .Q(WX7297) );
  INVX0 U6028_U1 ( .INP(n4483), .ZN(U6028_n1) );
  AND2X1 U6029_U2 ( .IN1(WX7232), .IN2(U6029_n1), .Q(WX7295) );
  INVX0 U6029_U1 ( .INP(n4483), .ZN(U6029_n1) );
  AND2X1 U6030_U2 ( .IN1(WX7230), .IN2(U6030_n1), .Q(WX7293) );
  INVX0 U6030_U1 ( .INP(n4483), .ZN(U6030_n1) );
  AND2X1 U6031_U2 ( .IN1(WX7228), .IN2(U6031_n1), .Q(WX7291) );
  INVX0 U6031_U1 ( .INP(n4483), .ZN(U6031_n1) );
  AND2X1 U6032_U2 ( .IN1(WX7226), .IN2(U6032_n1), .Q(WX7289) );
  INVX0 U6032_U1 ( .INP(n4483), .ZN(U6032_n1) );
  AND2X1 U6033_U2 ( .IN1(WX7224), .IN2(U6033_n1), .Q(WX7287) );
  INVX0 U6033_U1 ( .INP(n4483), .ZN(U6033_n1) );
  AND2X1 U6034_U2 ( .IN1(WX7222), .IN2(U6034_n1), .Q(WX7285) );
  INVX0 U6034_U1 ( .INP(n4484), .ZN(U6034_n1) );
  AND2X1 U6035_U2 ( .IN1(test_so60), .IN2(U6035_n1), .Q(WX7283) );
  INVX0 U6035_U1 ( .INP(n4484), .ZN(U6035_n1) );
  AND2X1 U6036_U2 ( .IN1(WX7218), .IN2(U6036_n1), .Q(WX7281) );
  INVX0 U6036_U1 ( .INP(n4484), .ZN(U6036_n1) );
  AND2X1 U6037_U2 ( .IN1(WX7216), .IN2(U6037_n1), .Q(WX7279) );
  INVX0 U6037_U1 ( .INP(n4484), .ZN(U6037_n1) );
  AND2X1 U6038_U2 ( .IN1(WX7214), .IN2(U6038_n1), .Q(WX7277) );
  INVX0 U6038_U1 ( .INP(n4484), .ZN(U6038_n1) );
  AND2X1 U6039_U2 ( .IN1(WX7212), .IN2(U6039_n1), .Q(WX7275) );
  INVX0 U6039_U1 ( .INP(n4484), .ZN(U6039_n1) );
  AND2X1 U6040_U2 ( .IN1(WX7210), .IN2(U6040_n1), .Q(WX7273) );
  INVX0 U6040_U1 ( .INP(n4484), .ZN(U6040_n1) );
  AND2X1 U6041_U2 ( .IN1(WX7208), .IN2(U6041_n1), .Q(WX7271) );
  INVX0 U6041_U1 ( .INP(n4484), .ZN(U6041_n1) );
  AND2X1 U6042_U2 ( .IN1(WX7206), .IN2(U6042_n1), .Q(WX7269) );
  INVX0 U6042_U1 ( .INP(n4484), .ZN(U6042_n1) );
  AND2X1 U6043_U2 ( .IN1(WX7204), .IN2(U6043_n1), .Q(WX7267) );
  INVX0 U6043_U1 ( .INP(n4484), .ZN(U6043_n1) );
  AND2X1 U6044_U2 ( .IN1(WX7202), .IN2(U6044_n1), .Q(WX7265) );
  INVX0 U6044_U1 ( .INP(n4484), .ZN(U6044_n1) );
  AND2X1 U6045_U2 ( .IN1(WX7200), .IN2(U6045_n1), .Q(WX7263) );
  INVX0 U6045_U1 ( .INP(n4484), .ZN(U6045_n1) );
  AND2X1 U6046_U2 ( .IN1(WX7198), .IN2(U6046_n1), .Q(WX7261) );
  INVX0 U6046_U1 ( .INP(n4484), .ZN(U6046_n1) );
  AND2X1 U6047_U2 ( .IN1(WX7196), .IN2(U6047_n1), .Q(WX7259) );
  INVX0 U6047_U1 ( .INP(n4484), .ZN(U6047_n1) );
  AND2X1 U6048_U2 ( .IN1(WX7194), .IN2(U6048_n1), .Q(WX7257) );
  INVX0 U6048_U1 ( .INP(n4485), .ZN(U6048_n1) );
  AND2X1 U6049_U2 ( .IN1(WX7192), .IN2(U6049_n1), .Q(WX7255) );
  INVX0 U6049_U1 ( .INP(n4485), .ZN(U6049_n1) );
  AND2X1 U6050_U2 ( .IN1(WX7190), .IN2(U6050_n1), .Q(WX7253) );
  INVX0 U6050_U1 ( .INP(n4485), .ZN(U6050_n1) );
  AND2X1 U6051_U2 ( .IN1(WX7188), .IN2(U6051_n1), .Q(WX7251) );
  INVX0 U6051_U1 ( .INP(n4485), .ZN(U6051_n1) );
  AND2X1 U6052_U2 ( .IN1(test_so59), .IN2(U6052_n1), .Q(WX7249) );
  INVX0 U6052_U1 ( .INP(n4485), .ZN(U6052_n1) );
  AND2X1 U6053_U2 ( .IN1(WX7184), .IN2(U6053_n1), .Q(WX7247) );
  INVX0 U6053_U1 ( .INP(n4485), .ZN(U6053_n1) );
  AND2X1 U6054_U2 ( .IN1(WX7182), .IN2(U6054_n1), .Q(WX7245) );
  INVX0 U6054_U1 ( .INP(n4485), .ZN(U6054_n1) );
  AND2X1 U6055_U2 ( .IN1(WX7180), .IN2(U6055_n1), .Q(WX7243) );
  INVX0 U6055_U1 ( .INP(n4485), .ZN(U6055_n1) );
  AND2X1 U6056_U2 ( .IN1(WX7178), .IN2(U6056_n1), .Q(WX7241) );
  INVX0 U6056_U1 ( .INP(n4485), .ZN(U6056_n1) );
  AND2X1 U6057_U2 ( .IN1(WX7176), .IN2(U6057_n1), .Q(WX7239) );
  INVX0 U6057_U1 ( .INP(n4485), .ZN(U6057_n1) );
  AND2X1 U6058_U2 ( .IN1(WX7174), .IN2(U6058_n1), .Q(WX7237) );
  INVX0 U6058_U1 ( .INP(n4485), .ZN(U6058_n1) );
  AND2X1 U6059_U2 ( .IN1(WX7172), .IN2(U6059_n1), .Q(WX7235) );
  INVX0 U6059_U1 ( .INP(n4485), .ZN(U6059_n1) );
  AND2X1 U6060_U2 ( .IN1(WX7170), .IN2(U6060_n1), .Q(WX7233) );
  INVX0 U6060_U1 ( .INP(n4485), .ZN(U6060_n1) );
  AND2X1 U6061_U2 ( .IN1(WX7168), .IN2(U6061_n1), .Q(WX7231) );
  INVX0 U6061_U1 ( .INP(n4485), .ZN(U6061_n1) );
  AND2X1 U6062_U2 ( .IN1(WX7166), .IN2(U6062_n1), .Q(WX7229) );
  INVX0 U6062_U1 ( .INP(n4486), .ZN(U6062_n1) );
  AND2X1 U6063_U2 ( .IN1(WX7164), .IN2(U6063_n1), .Q(WX7227) );
  INVX0 U6063_U1 ( .INP(n4486), .ZN(U6063_n1) );
  AND2X1 U6064_U2 ( .IN1(WX7162), .IN2(U6064_n1), .Q(WX7225) );
  INVX0 U6064_U1 ( .INP(n4486), .ZN(U6064_n1) );
  AND2X1 U6065_U2 ( .IN1(WX7160), .IN2(U6065_n1), .Q(WX7223) );
  INVX0 U6065_U1 ( .INP(n4486), .ZN(U6065_n1) );
  AND2X1 U6066_U2 ( .IN1(WX7158), .IN2(U6066_n1), .Q(WX7221) );
  INVX0 U6066_U1 ( .INP(n4486), .ZN(U6066_n1) );
  AND2X1 U6067_U2 ( .IN1(WX7156), .IN2(U6067_n1), .Q(WX7219) );
  INVX0 U6067_U1 ( .INP(n4486), .ZN(U6067_n1) );
  AND2X1 U6068_U2 ( .IN1(WX7154), .IN2(U6068_n1), .Q(WX7217) );
  INVX0 U6068_U1 ( .INP(n4486), .ZN(U6068_n1) );
  AND2X1 U6069_U2 ( .IN1(test_so58), .IN2(U6069_n1), .Q(WX7215) );
  INVX0 U6069_U1 ( .INP(n4486), .ZN(U6069_n1) );
  AND2X1 U6070_U2 ( .IN1(WX7150), .IN2(U6070_n1), .Q(WX7213) );
  INVX0 U6070_U1 ( .INP(n4486), .ZN(U6070_n1) );
  AND2X1 U6071_U2 ( .IN1(WX7148), .IN2(U6071_n1), .Q(WX7211) );
  INVX0 U6071_U1 ( .INP(n4486), .ZN(U6071_n1) );
  AND2X1 U6072_U2 ( .IN1(WX7146), .IN2(U6072_n1), .Q(WX7209) );
  INVX0 U6072_U1 ( .INP(n4486), .ZN(U6072_n1) );
  AND2X1 U6073_U2 ( .IN1(WX7144), .IN2(U6073_n1), .Q(WX7207) );
  INVX0 U6073_U1 ( .INP(n4486), .ZN(U6073_n1) );
  AND2X1 U6074_U2 ( .IN1(WX7142), .IN2(U6074_n1), .Q(WX7205) );
  INVX0 U6074_U1 ( .INP(n4486), .ZN(U6074_n1) );
  AND2X1 U6075_U2 ( .IN1(WX6007), .IN2(U6075_n1), .Q(WX6070) );
  INVX0 U6075_U1 ( .INP(n4487), .ZN(U6075_n1) );
  AND2X1 U6076_U2 ( .IN1(test_so51), .IN2(U6076_n1), .Q(WX6068) );
  INVX0 U6076_U1 ( .INP(n4487), .ZN(U6076_n1) );
  AND2X1 U6077_U2 ( .IN1(WX6003), .IN2(U6077_n1), .Q(WX6066) );
  INVX0 U6077_U1 ( .INP(n4487), .ZN(U6077_n1) );
  AND2X1 U6078_U2 ( .IN1(WX6001), .IN2(U6078_n1), .Q(WX6064) );
  INVX0 U6078_U1 ( .INP(n4487), .ZN(U6078_n1) );
  AND2X1 U6079_U2 ( .IN1(WX5999), .IN2(U6079_n1), .Q(WX6062) );
  INVX0 U6079_U1 ( .INP(n4487), .ZN(U6079_n1) );
  AND2X1 U6080_U2 ( .IN1(WX5997), .IN2(U6080_n1), .Q(WX6060) );
  INVX0 U6080_U1 ( .INP(n4487), .ZN(U6080_n1) );
  AND2X1 U6081_U2 ( .IN1(WX5995), .IN2(U6081_n1), .Q(WX6058) );
  INVX0 U6081_U1 ( .INP(n4487), .ZN(U6081_n1) );
  AND2X1 U6082_U2 ( .IN1(WX5993), .IN2(U6082_n1), .Q(WX6056) );
  INVX0 U6082_U1 ( .INP(n4487), .ZN(U6082_n1) );
  AND2X1 U6083_U2 ( .IN1(WX5991), .IN2(U6083_n1), .Q(WX6054) );
  INVX0 U6083_U1 ( .INP(n4487), .ZN(U6083_n1) );
  AND2X1 U6084_U2 ( .IN1(WX5989), .IN2(U6084_n1), .Q(WX6052) );
  INVX0 U6084_U1 ( .INP(n4487), .ZN(U6084_n1) );
  AND2X1 U6085_U2 ( .IN1(WX5987), .IN2(U6085_n1), .Q(WX6050) );
  INVX0 U6085_U1 ( .INP(n4487), .ZN(U6085_n1) );
  AND2X1 U6086_U2 ( .IN1(WX5985), .IN2(U6086_n1), .Q(WX6048) );
  INVX0 U6086_U1 ( .INP(n4487), .ZN(U6086_n1) );
  AND2X1 U6087_U2 ( .IN1(WX5983), .IN2(U6087_n1), .Q(WX6046) );
  INVX0 U6087_U1 ( .INP(n4487), .ZN(U6087_n1) );
  AND2X1 U6088_U2 ( .IN1(WX5981), .IN2(U6088_n1), .Q(WX6044) );
  INVX0 U6088_U1 ( .INP(n4487), .ZN(U6088_n1) );
  AND2X1 U6089_U2 ( .IN1(WX5979), .IN2(U6089_n1), .Q(WX6042) );
  INVX0 U6089_U1 ( .INP(n4488), .ZN(U6089_n1) );
  AND2X1 U6090_U2 ( .IN1(WX5977), .IN2(U6090_n1), .Q(WX6040) );
  INVX0 U6090_U1 ( .INP(n4488), .ZN(U6090_n1) );
  AND2X1 U6091_U2 ( .IN1(WX5975), .IN2(U6091_n1), .Q(WX6038) );
  INVX0 U6091_U1 ( .INP(n4488), .ZN(U6091_n1) );
  AND2X1 U6092_U2 ( .IN1(WX5973), .IN2(U6092_n1), .Q(WX6036) );
  INVX0 U6092_U1 ( .INP(n4488), .ZN(U6092_n1) );
  AND2X1 U6093_U2 ( .IN1(test_so50), .IN2(U6093_n1), .Q(WX6034) );
  INVX0 U6093_U1 ( .INP(n4488), .ZN(U6093_n1) );
  AND2X1 U6094_U2 ( .IN1(WX5969), .IN2(U6094_n1), .Q(WX6032) );
  INVX0 U6094_U1 ( .INP(n4488), .ZN(U6094_n1) );
  AND2X1 U6095_U2 ( .IN1(WX5967), .IN2(U6095_n1), .Q(WX6030) );
  INVX0 U6095_U1 ( .INP(n4488), .ZN(U6095_n1) );
  AND2X1 U6096_U2 ( .IN1(WX5965), .IN2(U6096_n1), .Q(WX6028) );
  INVX0 U6096_U1 ( .INP(n4488), .ZN(U6096_n1) );
  AND2X1 U6097_U2 ( .IN1(WX5963), .IN2(U6097_n1), .Q(WX6026) );
  INVX0 U6097_U1 ( .INP(n4488), .ZN(U6097_n1) );
  AND2X1 U6098_U2 ( .IN1(WX5961), .IN2(U6098_n1), .Q(WX6024) );
  INVX0 U6098_U1 ( .INP(n4488), .ZN(U6098_n1) );
  AND2X1 U6099_U2 ( .IN1(WX5959), .IN2(U6099_n1), .Q(WX6022) );
  INVX0 U6099_U1 ( .INP(n4488), .ZN(U6099_n1) );
  AND2X1 U6100_U2 ( .IN1(WX5957), .IN2(U6100_n1), .Q(WX6020) );
  INVX0 U6100_U1 ( .INP(n4488), .ZN(U6100_n1) );
  AND2X1 U6101_U2 ( .IN1(WX5955), .IN2(U6101_n1), .Q(WX6018) );
  INVX0 U6101_U1 ( .INP(n4488), .ZN(U6101_n1) );
  AND2X1 U6102_U2 ( .IN1(WX5953), .IN2(U6102_n1), .Q(WX6016) );
  INVX0 U6102_U1 ( .INP(n4488), .ZN(U6102_n1) );
  AND2X1 U6103_U2 ( .IN1(WX5951), .IN2(U6103_n1), .Q(WX6014) );
  INVX0 U6103_U1 ( .INP(n4489), .ZN(U6103_n1) );
  AND2X1 U6104_U2 ( .IN1(WX5949), .IN2(U6104_n1), .Q(WX6012) );
  INVX0 U6104_U1 ( .INP(n4489), .ZN(U6104_n1) );
  AND2X1 U6105_U2 ( .IN1(WX5947), .IN2(U6105_n1), .Q(WX6010) );
  INVX0 U6105_U1 ( .INP(n4489), .ZN(U6105_n1) );
  AND2X1 U6106_U2 ( .IN1(WX5945), .IN2(U6106_n1), .Q(WX6008) );
  INVX0 U6106_U1 ( .INP(n4489), .ZN(U6106_n1) );
  AND2X1 U6107_U2 ( .IN1(WX5943), .IN2(U6107_n1), .Q(WX6006) );
  INVX0 U6107_U1 ( .INP(n4489), .ZN(U6107_n1) );
  AND2X1 U6108_U2 ( .IN1(WX5941), .IN2(U6108_n1), .Q(WX6004) );
  INVX0 U6108_U1 ( .INP(n4489), .ZN(U6108_n1) );
  AND2X1 U6109_U2 ( .IN1(WX5929), .IN2(U6109_n1), .Q(WX5992) );
  INVX0 U6109_U1 ( .INP(n4489), .ZN(U6109_n1) );
  AND2X1 U6110_U2 ( .IN1(WX5927), .IN2(U6110_n1), .Q(WX5990) );
  INVX0 U6110_U1 ( .INP(n4489), .ZN(U6110_n1) );
  AND2X1 U6111_U2 ( .IN1(WX5925), .IN2(U6111_n1), .Q(WX5988) );
  INVX0 U6111_U1 ( .INP(n4489), .ZN(U6111_n1) );
  AND2X1 U6112_U2 ( .IN1(WX5923), .IN2(U6112_n1), .Q(WX5986) );
  INVX0 U6112_U1 ( .INP(n4489), .ZN(U6112_n1) );
  AND2X1 U6113_U2 ( .IN1(WX5921), .IN2(U6113_n1), .Q(WX5984) );
  INVX0 U6113_U1 ( .INP(n4489), .ZN(U6113_n1) );
  AND2X1 U6114_U2 ( .IN1(WX5919), .IN2(U6114_n1), .Q(WX5982) );
  INVX0 U6114_U1 ( .INP(n4489), .ZN(U6114_n1) );
  AND2X1 U6115_U2 ( .IN1(WX5917), .IN2(U6115_n1), .Q(WX5980) );
  INVX0 U6115_U1 ( .INP(n4489), .ZN(U6115_n1) );
  AND2X1 U6116_U2 ( .IN1(WX5915), .IN2(U6116_n1), .Q(WX5978) );
  INVX0 U6116_U1 ( .INP(n4489), .ZN(U6116_n1) );
  AND2X1 U6117_U2 ( .IN1(WX5913), .IN2(U6117_n1), .Q(WX5976) );
  INVX0 U6117_U1 ( .INP(n4490), .ZN(U6117_n1) );
  AND2X1 U6118_U2 ( .IN1(WX5911), .IN2(U6118_n1), .Q(WX5974) );
  INVX0 U6118_U1 ( .INP(n4490), .ZN(U6118_n1) );
  AND2X1 U6119_U2 ( .IN1(WX5909), .IN2(U6119_n1), .Q(WX5972) );
  INVX0 U6119_U1 ( .INP(n4490), .ZN(U6119_n1) );
  AND2X1 U6120_U2 ( .IN1(WX5907), .IN2(U6120_n1), .Q(WX5970) );
  INVX0 U6120_U1 ( .INP(n4490), .ZN(U6120_n1) );
  AND2X1 U6121_U2 ( .IN1(WX5905), .IN2(U6121_n1), .Q(WX5968) );
  INVX0 U6121_U1 ( .INP(n4490), .ZN(U6121_n1) );
  AND2X1 U6122_U2 ( .IN1(test_so48), .IN2(U6122_n1), .Q(WX5966) );
  INVX0 U6122_U1 ( .INP(n4490), .ZN(U6122_n1) );
  AND2X1 U6123_U2 ( .IN1(WX5901), .IN2(U6123_n1), .Q(WX5964) );
  INVX0 U6123_U1 ( .INP(n4490), .ZN(U6123_n1) );
  AND2X1 U6124_U2 ( .IN1(WX5899), .IN2(U6124_n1), .Q(WX5962) );
  INVX0 U6124_U1 ( .INP(n4490), .ZN(U6124_n1) );
  AND2X1 U6125_U2 ( .IN1(WX5897), .IN2(U6125_n1), .Q(WX5960) );
  INVX0 U6125_U1 ( .INP(n4490), .ZN(U6125_n1) );
  AND2X1 U6126_U2 ( .IN1(WX5895), .IN2(U6126_n1), .Q(WX5958) );
  INVX0 U6126_U1 ( .INP(n4490), .ZN(U6126_n1) );
  AND2X1 U6127_U2 ( .IN1(WX5893), .IN2(U6127_n1), .Q(WX5956) );
  INVX0 U6127_U1 ( .INP(n4490), .ZN(U6127_n1) );
  AND2X1 U6128_U2 ( .IN1(WX5891), .IN2(U6128_n1), .Q(WX5954) );
  INVX0 U6128_U1 ( .INP(n4490), .ZN(U6128_n1) );
  AND2X1 U6129_U2 ( .IN1(WX5889), .IN2(U6129_n1), .Q(WX5952) );
  INVX0 U6129_U1 ( .INP(n4490), .ZN(U6129_n1) );
  AND2X1 U6130_U2 ( .IN1(WX5887), .IN2(U6130_n1), .Q(WX5950) );
  INVX0 U6130_U1 ( .INP(n4490), .ZN(U6130_n1) );
  AND2X1 U6131_U2 ( .IN1(WX5885), .IN2(U6131_n1), .Q(WX5948) );
  INVX0 U6131_U1 ( .INP(n4479), .ZN(U6131_n1) );
  AND2X1 U6132_U2 ( .IN1(WX5883), .IN2(U6132_n1), .Q(WX5946) );
  INVX0 U6132_U1 ( .INP(n4480), .ZN(U6132_n1) );
  AND2X1 U6133_U2 ( .IN1(WX5881), .IN2(U6133_n1), .Q(WX5944) );
  INVX0 U6133_U1 ( .INP(n4476), .ZN(U6133_n1) );
  AND2X1 U6134_U2 ( .IN1(WX5879), .IN2(U6134_n1), .Q(WX5942) );
  INVX0 U6134_U1 ( .INP(n4471), .ZN(U6134_n1) );
  AND2X1 U6135_U2 ( .IN1(WX5877), .IN2(U6135_n1), .Q(WX5940) );
  INVX0 U6135_U1 ( .INP(n4471), .ZN(U6135_n1) );
  AND2X1 U6136_U2 ( .IN1(WX5875), .IN2(U6136_n1), .Q(WX5938) );
  INVX0 U6136_U1 ( .INP(n4471), .ZN(U6136_n1) );
  AND2X1 U6137_U2 ( .IN1(WX5873), .IN2(U6137_n1), .Q(WX5936) );
  INVX0 U6137_U1 ( .INP(n4471), .ZN(U6137_n1) );
  AND2X1 U6138_U2 ( .IN1(WX5871), .IN2(U6138_n1), .Q(WX5934) );
  INVX0 U6138_U1 ( .INP(n4471), .ZN(U6138_n1) );
  AND2X1 U6139_U2 ( .IN1(test_so47), .IN2(U6139_n1), .Q(WX5932) );
  INVX0 U6139_U1 ( .INP(n4471), .ZN(U6139_n1) );
  AND2X1 U6140_U2 ( .IN1(WX5867), .IN2(U6140_n1), .Q(WX5930) );
  INVX0 U6140_U1 ( .INP(n4471), .ZN(U6140_n1) );
  AND2X1 U6141_U2 ( .IN1(WX5865), .IN2(U6141_n1), .Q(WX5928) );
  INVX0 U6141_U1 ( .INP(n4471), .ZN(U6141_n1) );
  AND2X1 U6142_U2 ( .IN1(WX5863), .IN2(U6142_n1), .Q(WX5926) );
  INVX0 U6142_U1 ( .INP(n4472), .ZN(U6142_n1) );
  AND2X1 U6143_U2 ( .IN1(WX5861), .IN2(U6143_n1), .Q(WX5924) );
  INVX0 U6143_U1 ( .INP(n4472), .ZN(U6143_n1) );
  AND2X1 U6144_U2 ( .IN1(WX5859), .IN2(U6144_n1), .Q(WX5922) );
  INVX0 U6144_U1 ( .INP(n4472), .ZN(U6144_n1) );
  AND2X1 U6145_U2 ( .IN1(WX5857), .IN2(U6145_n1), .Q(WX5920) );
  INVX0 U6145_U1 ( .INP(n4472), .ZN(U6145_n1) );
  AND2X1 U6146_U2 ( .IN1(WX5855), .IN2(U6146_n1), .Q(WX5918) );
  INVX0 U6146_U1 ( .INP(n4472), .ZN(U6146_n1) );
  AND2X1 U6147_U2 ( .IN1(WX5853), .IN2(U6147_n1), .Q(WX5916) );
  INVX0 U6147_U1 ( .INP(n4472), .ZN(U6147_n1) );
  AND2X1 U6148_U2 ( .IN1(WX5851), .IN2(U6148_n1), .Q(WX5914) );
  INVX0 U6148_U1 ( .INP(n4472), .ZN(U6148_n1) );
  AND2X1 U6149_U2 ( .IN1(WX5849), .IN2(U6149_n1), .Q(WX5912) );
  INVX0 U6149_U1 ( .INP(n4472), .ZN(U6149_n1) );
  AND2X1 U6150_U2 ( .IN1(WX4714), .IN2(U6150_n1), .Q(WX4777) );
  INVX0 U6150_U1 ( .INP(n4472), .ZN(U6150_n1) );
  AND2X1 U6151_U2 ( .IN1(WX4712), .IN2(U6151_n1), .Q(WX4775) );
  INVX0 U6151_U1 ( .INP(n4472), .ZN(U6151_n1) );
  AND2X1 U6152_U2 ( .IN1(WX4710), .IN2(U6152_n1), .Q(WX4773) );
  INVX0 U6152_U1 ( .INP(n4472), .ZN(U6152_n1) );
  AND2X1 U6153_U2 ( .IN1(WX4708), .IN2(U6153_n1), .Q(WX4771) );
  INVX0 U6153_U1 ( .INP(n4472), .ZN(U6153_n1) );
  AND2X1 U6154_U2 ( .IN1(WX4706), .IN2(U6154_n1), .Q(WX4769) );
  INVX0 U6154_U1 ( .INP(n4472), .ZN(U6154_n1) );
  AND2X1 U6155_U2 ( .IN1(WX4704), .IN2(U6155_n1), .Q(WX4767) );
  INVX0 U6155_U1 ( .INP(n4472), .ZN(U6155_n1) );
  AND2X1 U6156_U2 ( .IN1(WX4702), .IN2(U6156_n1), .Q(WX4765) );
  INVX0 U6156_U1 ( .INP(n4473), .ZN(U6156_n1) );
  AND2X1 U6157_U2 ( .IN1(WX4700), .IN2(U6157_n1), .Q(WX4763) );
  INVX0 U6157_U1 ( .INP(n4473), .ZN(U6157_n1) );
  AND2X1 U6158_U2 ( .IN1(WX4698), .IN2(U6158_n1), .Q(WX4761) );
  INVX0 U6158_U1 ( .INP(n4473), .ZN(U6158_n1) );
  AND2X1 U6159_U2 ( .IN1(WX4696), .IN2(U6159_n1), .Q(WX4759) );
  INVX0 U6159_U1 ( .INP(n4473), .ZN(U6159_n1) );
  AND2X1 U6160_U2 ( .IN1(WX4694), .IN2(U6160_n1), .Q(WX4757) );
  INVX0 U6160_U1 ( .INP(n4473), .ZN(U6160_n1) );
  AND2X1 U6161_U2 ( .IN1(WX4692), .IN2(U6161_n1), .Q(WX4755) );
  INVX0 U6161_U1 ( .INP(n4473), .ZN(U6161_n1) );
  AND2X1 U6162_U2 ( .IN1(WX4690), .IN2(U6162_n1), .Q(WX4753) );
  INVX0 U6162_U1 ( .INP(n4473), .ZN(U6162_n1) );
  AND2X1 U6163_U2 ( .IN1(test_so39), .IN2(U6163_n1), .Q(WX4751) );
  INVX0 U6163_U1 ( .INP(n4473), .ZN(U6163_n1) );
  AND2X1 U6164_U2 ( .IN1(WX4686), .IN2(U6164_n1), .Q(WX4749) );
  INVX0 U6164_U1 ( .INP(n4473), .ZN(U6164_n1) );
  AND2X1 U6165_U2 ( .IN1(WX4684), .IN2(U6165_n1), .Q(WX4747) );
  INVX0 U6165_U1 ( .INP(n4473), .ZN(U6165_n1) );
  AND2X1 U6166_U2 ( .IN1(WX4682), .IN2(U6166_n1), .Q(WX4745) );
  INVX0 U6166_U1 ( .INP(n4473), .ZN(U6166_n1) );
  AND2X1 U6167_U2 ( .IN1(WX4680), .IN2(U6167_n1), .Q(WX4743) );
  INVX0 U6167_U1 ( .INP(n4473), .ZN(U6167_n1) );
  AND2X1 U6168_U2 ( .IN1(WX4678), .IN2(U6168_n1), .Q(WX4741) );
  INVX0 U6168_U1 ( .INP(n4473), .ZN(U6168_n1) );
  AND2X1 U6169_U2 ( .IN1(WX4676), .IN2(U6169_n1), .Q(WX4739) );
  INVX0 U6169_U1 ( .INP(n4473), .ZN(U6169_n1) );
  AND2X1 U6170_U2 ( .IN1(WX4674), .IN2(U6170_n1), .Q(WX4737) );
  INVX0 U6170_U1 ( .INP(n4474), .ZN(U6170_n1) );
  AND2X1 U6171_U2 ( .IN1(WX4672), .IN2(U6171_n1), .Q(WX4735) );
  INVX0 U6171_U1 ( .INP(n4474), .ZN(U6171_n1) );
  AND2X1 U6172_U2 ( .IN1(WX4670), .IN2(U6172_n1), .Q(WX4733) );
  INVX0 U6172_U1 ( .INP(n4474), .ZN(U6172_n1) );
  AND2X1 U6173_U2 ( .IN1(WX4668), .IN2(U6173_n1), .Q(WX4731) );
  INVX0 U6173_U1 ( .INP(n4474), .ZN(U6173_n1) );
  AND2X1 U6174_U2 ( .IN1(WX4666), .IN2(U6174_n1), .Q(WX4729) );
  INVX0 U6174_U1 ( .INP(n4474), .ZN(U6174_n1) );
  AND2X1 U6175_U2 ( .IN1(WX4664), .IN2(U6175_n1), .Q(WX4727) );
  INVX0 U6175_U1 ( .INP(n4474), .ZN(U6175_n1) );
  AND2X1 U6176_U2 ( .IN1(WX4662), .IN2(U6176_n1), .Q(WX4725) );
  INVX0 U6176_U1 ( .INP(n4474), .ZN(U6176_n1) );
  AND2X1 U6177_U2 ( .IN1(WX4660), .IN2(U6177_n1), .Q(WX4723) );
  INVX0 U6177_U1 ( .INP(n4474), .ZN(U6177_n1) );
  AND2X1 U6178_U2 ( .IN1(WX4658), .IN2(U6178_n1), .Q(WX4721) );
  INVX0 U6178_U1 ( .INP(n4474), .ZN(U6178_n1) );
  AND2X1 U6179_U2 ( .IN1(WX4656), .IN2(U6179_n1), .Q(WX4719) );
  INVX0 U6179_U1 ( .INP(n4474), .ZN(U6179_n1) );
  AND2X1 U6180_U2 ( .IN1(test_so38), .IN2(U6180_n1), .Q(WX4717) );
  INVX0 U6180_U1 ( .INP(n4474), .ZN(U6180_n1) );
  AND2X1 U6181_U2 ( .IN1(WX4652), .IN2(U6181_n1), .Q(WX4715) );
  INVX0 U6181_U1 ( .INP(n4474), .ZN(U6181_n1) );
  AND2X1 U6182_U2 ( .IN1(WX4650), .IN2(U6182_n1), .Q(WX4713) );
  INVX0 U6182_U1 ( .INP(n4474), .ZN(U6182_n1) );
  AND2X1 U6183_U2 ( .IN1(WX4648), .IN2(U6183_n1), .Q(WX4711) );
  INVX0 U6183_U1 ( .INP(n4474), .ZN(U6183_n1) );
  AND2X1 U6184_U2 ( .IN1(WX4646), .IN2(U6184_n1), .Q(WX4709) );
  INVX0 U6184_U1 ( .INP(n4475), .ZN(U6184_n1) );
  AND2X1 U6185_U2 ( .IN1(WX4644), .IN2(U6185_n1), .Q(WX4707) );
  INVX0 U6185_U1 ( .INP(n4475), .ZN(U6185_n1) );
  AND2X1 U6186_U2 ( .IN1(WX4642), .IN2(U6186_n1), .Q(WX4705) );
  INVX0 U6186_U1 ( .INP(n4475), .ZN(U6186_n1) );
  AND2X1 U6187_U2 ( .IN1(WX4640), .IN2(U6187_n1), .Q(WX4703) );
  INVX0 U6187_U1 ( .INP(n4475), .ZN(U6187_n1) );
  AND2X1 U6188_U2 ( .IN1(WX4638), .IN2(U6188_n1), .Q(WX4701) );
  INVX0 U6188_U1 ( .INP(n4475), .ZN(U6188_n1) );
  AND2X1 U6189_U2 ( .IN1(WX4636), .IN2(U6189_n1), .Q(WX4699) );
  INVX0 U6189_U1 ( .INP(n4475), .ZN(U6189_n1) );
  AND2X1 U6190_U2 ( .IN1(WX4634), .IN2(U6190_n1), .Q(WX4697) );
  INVX0 U6190_U1 ( .INP(n4475), .ZN(U6190_n1) );
  AND2X1 U6191_U2 ( .IN1(WX4632), .IN2(U6191_n1), .Q(WX4695) );
  INVX0 U6191_U1 ( .INP(n4475), .ZN(U6191_n1) );
  AND2X1 U6192_U2 ( .IN1(WX4630), .IN2(U6192_n1), .Q(WX4693) );
  INVX0 U6192_U1 ( .INP(n4475), .ZN(U6192_n1) );
  AND2X1 U6193_U2 ( .IN1(WX4628), .IN2(U6193_n1), .Q(WX4691) );
  INVX0 U6193_U1 ( .INP(n4475), .ZN(U6193_n1) );
  AND2X1 U6194_U2 ( .IN1(WX4626), .IN2(U6194_n1), .Q(WX4689) );
  INVX0 U6194_U1 ( .INP(n4475), .ZN(U6194_n1) );
  AND2X1 U6195_U2 ( .IN1(WX4624), .IN2(U6195_n1), .Q(WX4687) );
  INVX0 U6195_U1 ( .INP(n4475), .ZN(U6195_n1) );
  AND2X1 U6196_U2 ( .IN1(WX4622), .IN2(U6196_n1), .Q(WX4685) );
  INVX0 U6196_U1 ( .INP(n4475), .ZN(U6196_n1) );
  AND2X1 U6197_U2 ( .IN1(test_so37), .IN2(U6197_n1), .Q(WX4683) );
  INVX0 U6197_U1 ( .INP(n4475), .ZN(U6197_n1) );
  AND2X1 U6198_U2 ( .IN1(WX4618), .IN2(U6198_n1), .Q(WX4681) );
  INVX0 U6198_U1 ( .INP(n4476), .ZN(U6198_n1) );
  AND2X1 U6199_U2 ( .IN1(WX4616), .IN2(U6199_n1), .Q(WX4679) );
  INVX0 U6199_U1 ( .INP(n4476), .ZN(U6199_n1) );
  AND2X1 U6200_U2 ( .IN1(WX4614), .IN2(U6200_n1), .Q(WX4677) );
  INVX0 U6200_U1 ( .INP(n4476), .ZN(U6200_n1) );
  AND2X1 U6201_U2 ( .IN1(WX4612), .IN2(U6201_n1), .Q(WX4675) );
  INVX0 U6201_U1 ( .INP(n4476), .ZN(U6201_n1) );
  AND2X1 U6202_U2 ( .IN1(WX4610), .IN2(U6202_n1), .Q(WX4673) );
  INVX0 U6202_U1 ( .INP(n4476), .ZN(U6202_n1) );
  AND2X1 U6203_U2 ( .IN1(WX4608), .IN2(U6203_n1), .Q(WX4671) );
  INVX0 U6203_U1 ( .INP(n4476), .ZN(U6203_n1) );
  AND2X1 U6204_U2 ( .IN1(WX4606), .IN2(U6204_n1), .Q(WX4669) );
  INVX0 U6204_U1 ( .INP(n4476), .ZN(U6204_n1) );
  AND2X1 U6205_U2 ( .IN1(WX4604), .IN2(U6205_n1), .Q(WX4667) );
  INVX0 U6205_U1 ( .INP(n4476), .ZN(U6205_n1) );
  AND2X1 U6206_U2 ( .IN1(WX4602), .IN2(U6206_n1), .Q(WX4665) );
  INVX0 U6206_U1 ( .INP(n4476), .ZN(U6206_n1) );
  AND2X1 U6207_U2 ( .IN1(WX4600), .IN2(U6207_n1), .Q(WX4663) );
  INVX0 U6207_U1 ( .INP(n4476), .ZN(U6207_n1) );
  AND2X1 U6208_U2 ( .IN1(WX4598), .IN2(U6208_n1), .Q(WX4661) );
  INVX0 U6208_U1 ( .INP(n4476), .ZN(U6208_n1) );
  AND2X1 U6209_U2 ( .IN1(WX4596), .IN2(U6209_n1), .Q(WX4659) );
  INVX0 U6209_U1 ( .INP(n4476), .ZN(U6209_n1) );
  AND2X1 U6210_U2 ( .IN1(WX4594), .IN2(U6210_n1), .Q(WX4657) );
  INVX0 U6210_U1 ( .INP(n4476), .ZN(U6210_n1) );
  AND2X1 U6211_U2 ( .IN1(WX4592), .IN2(U6211_n1), .Q(WX4655) );
  INVX0 U6211_U1 ( .INP(n4477), .ZN(U6211_n1) );
  AND2X1 U6212_U2 ( .IN1(WX4590), .IN2(U6212_n1), .Q(WX4653) );
  INVX0 U6212_U1 ( .INP(n4477), .ZN(U6212_n1) );
  AND2X1 U6213_U2 ( .IN1(WX4588), .IN2(U6213_n1), .Q(WX4651) );
  INVX0 U6213_U1 ( .INP(n4477), .ZN(U6213_n1) );
  AND2X1 U6214_U2 ( .IN1(test_so36), .IN2(U6214_n1), .Q(WX4649) );
  INVX0 U6214_U1 ( .INP(n4477), .ZN(U6214_n1) );
  AND2X1 U6215_U2 ( .IN1(WX4584), .IN2(U6215_n1), .Q(WX4647) );
  INVX0 U6215_U1 ( .INP(n4477), .ZN(U6215_n1) );
  AND2X1 U6216_U2 ( .IN1(WX4582), .IN2(U6216_n1), .Q(WX4645) );
  INVX0 U6216_U1 ( .INP(n4477), .ZN(U6216_n1) );
  AND2X1 U6217_U2 ( .IN1(WX4580), .IN2(U6217_n1), .Q(WX4643) );
  INVX0 U6217_U1 ( .INP(n4477), .ZN(U6217_n1) );
  AND2X1 U6218_U2 ( .IN1(WX4578), .IN2(U6218_n1), .Q(WX4641) );
  INVX0 U6218_U1 ( .INP(n4477), .ZN(U6218_n1) );
  AND2X1 U6219_U2 ( .IN1(WX4576), .IN2(U6219_n1), .Q(WX4639) );
  INVX0 U6219_U1 ( .INP(n4477), .ZN(U6219_n1) );
  AND2X1 U6220_U2 ( .IN1(WX4574), .IN2(U6220_n1), .Q(WX4637) );
  INVX0 U6220_U1 ( .INP(n4477), .ZN(U6220_n1) );
  AND2X1 U6221_U2 ( .IN1(WX4572), .IN2(U6221_n1), .Q(WX4635) );
  INVX0 U6221_U1 ( .INP(n4477), .ZN(U6221_n1) );
  AND2X1 U6222_U2 ( .IN1(WX4570), .IN2(U6222_n1), .Q(WX4633) );
  INVX0 U6222_U1 ( .INP(n4477), .ZN(U6222_n1) );
  AND2X1 U6223_U2 ( .IN1(WX4568), .IN2(U6223_n1), .Q(WX4631) );
  INVX0 U6223_U1 ( .INP(n4477), .ZN(U6223_n1) );
  AND2X1 U6224_U2 ( .IN1(WX4566), .IN2(U6224_n1), .Q(WX4629) );
  INVX0 U6224_U1 ( .INP(n4477), .ZN(U6224_n1) );
  AND2X1 U6225_U2 ( .IN1(WX4564), .IN2(U6225_n1), .Q(WX4627) );
  INVX0 U6225_U1 ( .INP(n4478), .ZN(U6225_n1) );
  AND2X1 U6226_U2 ( .IN1(WX4562), .IN2(U6226_n1), .Q(WX4625) );
  INVX0 U6226_U1 ( .INP(n4478), .ZN(U6226_n1) );
  AND2X1 U6227_U2 ( .IN1(WX4560), .IN2(U6227_n1), .Q(WX4623) );
  INVX0 U6227_U1 ( .INP(n4478), .ZN(U6227_n1) );
  AND2X1 U6228_U2 ( .IN1(WX4558), .IN2(U6228_n1), .Q(WX4621) );
  INVX0 U6228_U1 ( .INP(n4478), .ZN(U6228_n1) );
  AND2X1 U6229_U2 ( .IN1(WX4556), .IN2(U6229_n1), .Q(WX4619) );
  INVX0 U6229_U1 ( .INP(n4478), .ZN(U6229_n1) );
  AND2X1 U6230_U2 ( .IN1(WX3421), .IN2(U6230_n1), .Q(WX3484) );
  INVX0 U6230_U1 ( .INP(n4478), .ZN(U6230_n1) );
  AND2X1 U6231_U2 ( .IN1(WX3419), .IN2(U6231_n1), .Q(WX3482) );
  INVX0 U6231_U1 ( .INP(n4478), .ZN(U6231_n1) );
  AND2X1 U6232_U2 ( .IN1(WX3417), .IN2(U6232_n1), .Q(WX3480) );
  INVX0 U6232_U1 ( .INP(n4478), .ZN(U6232_n1) );
  AND2X1 U6233_U2 ( .IN1(WX3415), .IN2(U6233_n1), .Q(WX3478) );
  INVX0 U6233_U1 ( .INP(n4478), .ZN(U6233_n1) );
  AND2X1 U6234_U2 ( .IN1(WX3413), .IN2(U6234_n1), .Q(WX3476) );
  INVX0 U6234_U1 ( .INP(n4478), .ZN(U6234_n1) );
  AND2X1 U6235_U2 ( .IN1(WX3411), .IN2(U6235_n1), .Q(WX3474) );
  INVX0 U6235_U1 ( .INP(n4478), .ZN(U6235_n1) );
  AND2X1 U6236_U2 ( .IN1(WX3409), .IN2(U6236_n1), .Q(WX3472) );
  INVX0 U6236_U1 ( .INP(n4478), .ZN(U6236_n1) );
  AND2X1 U6237_U2 ( .IN1(WX3407), .IN2(U6237_n1), .Q(WX3470) );
  INVX0 U6237_U1 ( .INP(n4478), .ZN(U6237_n1) );
  AND2X1 U6238_U2 ( .IN1(test_so28), .IN2(U6238_n1), .Q(WX3468) );
  INVX0 U6238_U1 ( .INP(n4478), .ZN(U6238_n1) );
  AND2X1 U6239_U2 ( .IN1(WX3403), .IN2(U6239_n1), .Q(WX3466) );
  INVX0 U6239_U1 ( .INP(n4479), .ZN(U6239_n1) );
  AND2X1 U6240_U2 ( .IN1(WX3401), .IN2(U6240_n1), .Q(WX3464) );
  INVX0 U6240_U1 ( .INP(n4479), .ZN(U6240_n1) );
  AND2X1 U6241_U2 ( .IN1(WX3399), .IN2(U6241_n1), .Q(WX3462) );
  INVX0 U6241_U1 ( .INP(n4479), .ZN(U6241_n1) );
  AND2X1 U6242_U2 ( .IN1(WX3397), .IN2(U6242_n1), .Q(WX3460) );
  INVX0 U6242_U1 ( .INP(n4479), .ZN(U6242_n1) );
  AND2X1 U6243_U2 ( .IN1(WX3395), .IN2(U6243_n1), .Q(WX3458) );
  INVX0 U6243_U1 ( .INP(n4479), .ZN(U6243_n1) );
  AND2X1 U6244_U2 ( .IN1(WX3393), .IN2(U6244_n1), .Q(WX3456) );
  INVX0 U6244_U1 ( .INP(n4479), .ZN(U6244_n1) );
  AND2X1 U6245_U2 ( .IN1(WX3391), .IN2(U6245_n1), .Q(WX3454) );
  INVX0 U6245_U1 ( .INP(n4479), .ZN(U6245_n1) );
  AND2X1 U6246_U2 ( .IN1(WX3389), .IN2(U6246_n1), .Q(WX3452) );
  INVX0 U6246_U1 ( .INP(n4479), .ZN(U6246_n1) );
  AND2X1 U6247_U2 ( .IN1(WX3387), .IN2(U6247_n1), .Q(WX3450) );
  INVX0 U6247_U1 ( .INP(n4479), .ZN(U6247_n1) );
  AND2X1 U6248_U2 ( .IN1(WX3385), .IN2(U6248_n1), .Q(WX3448) );
  INVX0 U6248_U1 ( .INP(n4479), .ZN(U6248_n1) );
  AND2X1 U6249_U2 ( .IN1(WX3383), .IN2(U6249_n1), .Q(WX3446) );
  INVX0 U6249_U1 ( .INP(n4479), .ZN(U6249_n1) );
  AND2X1 U6250_U2 ( .IN1(WX3381), .IN2(U6250_n1), .Q(WX3444) );
  INVX0 U6250_U1 ( .INP(n4479), .ZN(U6250_n1) );
  AND2X1 U6251_U2 ( .IN1(WX3379), .IN2(U6251_n1), .Q(WX3442) );
  INVX0 U6251_U1 ( .INP(n4479), .ZN(U6251_n1) );
  AND2X1 U6252_U2 ( .IN1(WX3377), .IN2(U6252_n1), .Q(WX3440) );
  INVX0 U6252_U1 ( .INP(n4479), .ZN(U6252_n1) );
  AND2X1 U6253_U2 ( .IN1(WX3375), .IN2(U6253_n1), .Q(WX3438) );
  INVX0 U6253_U1 ( .INP(n4480), .ZN(U6253_n1) );
  AND2X1 U6254_U2 ( .IN1(WX3373), .IN2(U6254_n1), .Q(WX3436) );
  INVX0 U6254_U1 ( .INP(n4480), .ZN(U6254_n1) );
  AND2X1 U6255_U2 ( .IN1(WX3371), .IN2(U6255_n1), .Q(WX3434) );
  INVX0 U6255_U1 ( .INP(n4480), .ZN(U6255_n1) );
  AND2X1 U6256_U2 ( .IN1(test_so27), .IN2(U6256_n1), .Q(WX3432) );
  INVX0 U6256_U1 ( .INP(n4480), .ZN(U6256_n1) );
  AND2X1 U6257_U2 ( .IN1(WX3367), .IN2(U6257_n1), .Q(WX3430) );
  INVX0 U6257_U1 ( .INP(n4480), .ZN(U6257_n1) );
  AND2X1 U6258_U2 ( .IN1(WX3365), .IN2(U6258_n1), .Q(WX3428) );
  INVX0 U6258_U1 ( .INP(n4480), .ZN(U6258_n1) );
  AND2X1 U6259_U2 ( .IN1(WX3363), .IN2(U6259_n1), .Q(WX3426) );
  INVX0 U6259_U1 ( .INP(n4480), .ZN(U6259_n1) );
  AND2X1 U6260_U2 ( .IN1(WX3361), .IN2(U6260_n1), .Q(WX3424) );
  INVX0 U6260_U1 ( .INP(n4480), .ZN(U6260_n1) );
  AND2X1 U6261_U2 ( .IN1(WX3359), .IN2(U6261_n1), .Q(WX3422) );
  INVX0 U6261_U1 ( .INP(n4480), .ZN(U6261_n1) );
  AND2X1 U6262_U2 ( .IN1(WX3357), .IN2(U6262_n1), .Q(WX3420) );
  INVX0 U6262_U1 ( .INP(n4480), .ZN(U6262_n1) );
  AND2X1 U6263_U2 ( .IN1(WX3355), .IN2(U6263_n1), .Q(WX3418) );
  INVX0 U6263_U1 ( .INP(n4480), .ZN(U6263_n1) );
  AND2X1 U6264_U2 ( .IN1(WX3353), .IN2(U6264_n1), .Q(WX3416) );
  INVX0 U6264_U1 ( .INP(n4480), .ZN(U6264_n1) );
  AND2X1 U6265_U2 ( .IN1(WX3351), .IN2(U6265_n1), .Q(WX3414) );
  INVX0 U6265_U1 ( .INP(n4480), .ZN(U6265_n1) );
  AND2X1 U6266_U2 ( .IN1(WX3349), .IN2(U6266_n1), .Q(WX3412) );
  INVX0 U6266_U1 ( .INP(n4480), .ZN(U6266_n1) );
  AND2X1 U6267_U2 ( .IN1(WX3347), .IN2(U6267_n1), .Q(WX3410) );
  INVX0 U6267_U1 ( .INP(n4481), .ZN(U6267_n1) );
  AND2X1 U6268_U2 ( .IN1(WX3345), .IN2(U6268_n1), .Q(WX3408) );
  INVX0 U6268_U1 ( .INP(n4481), .ZN(U6268_n1) );
  AND2X1 U6269_U2 ( .IN1(WX3343), .IN2(U6269_n1), .Q(WX3406) );
  INVX0 U6269_U1 ( .INP(n4481), .ZN(U6269_n1) );
  AND2X1 U6270_U2 ( .IN1(WX3341), .IN2(U6270_n1), .Q(WX3404) );
  INVX0 U6270_U1 ( .INP(n4481), .ZN(U6270_n1) );
  AND2X1 U6271_U2 ( .IN1(WX3339), .IN2(U6271_n1), .Q(WX3402) );
  INVX0 U6271_U1 ( .INP(n4443), .ZN(U6271_n1) );
  AND2X1 U6272_U2 ( .IN1(WX3337), .IN2(U6272_n1), .Q(WX3400) );
  INVX0 U6272_U1 ( .INP(n4443), .ZN(U6272_n1) );
  AND2X1 U6273_U2 ( .IN1(WX3335), .IN2(U6273_n1), .Q(WX3398) );
  INVX0 U6273_U1 ( .INP(n4443), .ZN(U6273_n1) );
  AND2X1 U6274_U2 ( .IN1(test_so26), .IN2(U6274_n1), .Q(WX3396) );
  INVX0 U6274_U1 ( .INP(n4443), .ZN(U6274_n1) );
  AND2X1 U6275_U2 ( .IN1(WX3331), .IN2(U6275_n1), .Q(WX3394) );
  INVX0 U6275_U1 ( .INP(n4443), .ZN(U6275_n1) );
  AND2X1 U6276_U2 ( .IN1(WX3329), .IN2(U6276_n1), .Q(WX3392) );
  INVX0 U6276_U1 ( .INP(n4443), .ZN(U6276_n1) );
  AND2X1 U6277_U2 ( .IN1(WX3327), .IN2(U6277_n1), .Q(WX3390) );
  INVX0 U6277_U1 ( .INP(n4443), .ZN(U6277_n1) );
  AND2X1 U6278_U2 ( .IN1(WX3325), .IN2(U6278_n1), .Q(WX3388) );
  INVX0 U6278_U1 ( .INP(n4443), .ZN(U6278_n1) );
  AND2X1 U6279_U2 ( .IN1(WX3323), .IN2(U6279_n1), .Q(WX3386) );
  INVX0 U6279_U1 ( .INP(n4443), .ZN(U6279_n1) );
  AND2X1 U6280_U2 ( .IN1(WX3321), .IN2(U6280_n1), .Q(WX3384) );
  INVX0 U6280_U1 ( .INP(n4443), .ZN(U6280_n1) );
  AND2X1 U6281_U2 ( .IN1(WX3319), .IN2(U6281_n1), .Q(WX3382) );
  INVX0 U6281_U1 ( .INP(n4443), .ZN(U6281_n1) );
  AND2X1 U6282_U2 ( .IN1(WX3317), .IN2(U6282_n1), .Q(WX3380) );
  INVX0 U6282_U1 ( .INP(n4443), .ZN(U6282_n1) );
  AND2X1 U6283_U2 ( .IN1(WX3315), .IN2(U6283_n1), .Q(WX3378) );
  INVX0 U6283_U1 ( .INP(n4443), .ZN(U6283_n1) );
  AND2X1 U6284_U2 ( .IN1(WX3313), .IN2(U6284_n1), .Q(WX3376) );
  INVX0 U6284_U1 ( .INP(n4443), .ZN(U6284_n1) );
  AND2X1 U6285_U2 ( .IN1(WX3311), .IN2(U6285_n1), .Q(WX3374) );
  INVX0 U6285_U1 ( .INP(n4442), .ZN(U6285_n1) );
  AND2X1 U6286_U2 ( .IN1(WX3309), .IN2(U6286_n1), .Q(WX3372) );
  INVX0 U6286_U1 ( .INP(n4442), .ZN(U6286_n1) );
  AND2X1 U6287_U2 ( .IN1(WX3307), .IN2(U6287_n1), .Q(WX3370) );
  INVX0 U6287_U1 ( .INP(n4442), .ZN(U6287_n1) );
  AND2X1 U6288_U2 ( .IN1(WX3305), .IN2(U6288_n1), .Q(WX3368) );
  INVX0 U6288_U1 ( .INP(n4442), .ZN(U6288_n1) );
  AND2X1 U6289_U2 ( .IN1(WX3303), .IN2(U6289_n1), .Q(WX3366) );
  INVX0 U6289_U1 ( .INP(n4442), .ZN(U6289_n1) );
  AND2X1 U6290_U2 ( .IN1(WX3301), .IN2(U6290_n1), .Q(WX3364) );
  INVX0 U6290_U1 ( .INP(n4442), .ZN(U6290_n1) );
  AND2X1 U6291_U2 ( .IN1(WX3299), .IN2(U6291_n1), .Q(WX3362) );
  INVX0 U6291_U1 ( .INP(n4442), .ZN(U6291_n1) );
  AND2X1 U6292_U2 ( .IN1(test_so25), .IN2(U6292_n1), .Q(WX3360) );
  INVX0 U6292_U1 ( .INP(n4442), .ZN(U6292_n1) );
  AND2X1 U6293_U2 ( .IN1(WX3295), .IN2(U6293_n1), .Q(WX3358) );
  INVX0 U6293_U1 ( .INP(n4442), .ZN(U6293_n1) );
  AND2X1 U6294_U2 ( .IN1(WX3293), .IN2(U6294_n1), .Q(WX3356) );
  INVX0 U6294_U1 ( .INP(n4442), .ZN(U6294_n1) );
  AND2X1 U6295_U2 ( .IN1(WX3291), .IN2(U6295_n1), .Q(WX3354) );
  INVX0 U6295_U1 ( .INP(n4442), .ZN(U6295_n1) );
  AND2X1 U6296_U2 ( .IN1(WX3289), .IN2(U6296_n1), .Q(WX3352) );
  INVX0 U6296_U1 ( .INP(n4442), .ZN(U6296_n1) );
  AND2X1 U6297_U2 ( .IN1(WX3287), .IN2(U6297_n1), .Q(WX3350) );
  INVX0 U6297_U1 ( .INP(n4442), .ZN(U6297_n1) );
  AND2X1 U6298_U2 ( .IN1(WX3285), .IN2(U6298_n1), .Q(WX3348) );
  INVX0 U6298_U1 ( .INP(n4442), .ZN(U6298_n1) );
  AND2X1 U6299_U2 ( .IN1(WX3283), .IN2(U6299_n1), .Q(WX3346) );
  INVX0 U6299_U1 ( .INP(n4441), .ZN(U6299_n1) );
  AND2X1 U6300_U2 ( .IN1(WX3281), .IN2(U6300_n1), .Q(WX3344) );
  INVX0 U6300_U1 ( .INP(n4441), .ZN(U6300_n1) );
  AND2X1 U6301_U2 ( .IN1(WX3279), .IN2(U6301_n1), .Q(WX3342) );
  INVX0 U6301_U1 ( .INP(n4441), .ZN(U6301_n1) );
  AND2X1 U6302_U2 ( .IN1(WX3277), .IN2(U6302_n1), .Q(WX3340) );
  INVX0 U6302_U1 ( .INP(n4441), .ZN(U6302_n1) );
  AND2X1 U6303_U2 ( .IN1(WX3275), .IN2(U6303_n1), .Q(WX3338) );
  INVX0 U6303_U1 ( .INP(n4441), .ZN(U6303_n1) );
  AND2X1 U6304_U2 ( .IN1(WX3273), .IN2(U6304_n1), .Q(WX3336) );
  INVX0 U6304_U1 ( .INP(n4441), .ZN(U6304_n1) );
  AND2X1 U6305_U2 ( .IN1(WX3271), .IN2(U6305_n1), .Q(WX3334) );
  INVX0 U6305_U1 ( .INP(n4441), .ZN(U6305_n1) );
  AND2X1 U6306_U2 ( .IN1(WX3267), .IN2(U6306_n1), .Q(WX3330) );
  INVX0 U6306_U1 ( .INP(n4441), .ZN(U6306_n1) );
  AND2X1 U6307_U2 ( .IN1(WX2128), .IN2(U6307_n1), .Q(WX2191) );
  INVX0 U6307_U1 ( .INP(n4441), .ZN(U6307_n1) );
  AND2X1 U6308_U2 ( .IN1(WX2126), .IN2(U6308_n1), .Q(WX2189) );
  INVX0 U6308_U1 ( .INP(n4441), .ZN(U6308_n1) );
  AND2X1 U6309_U2 ( .IN1(WX2124), .IN2(U6309_n1), .Q(WX2187) );
  INVX0 U6309_U1 ( .INP(n4441), .ZN(U6309_n1) );
  AND2X1 U6310_U2 ( .IN1(WX2122), .IN2(U6310_n1), .Q(WX2185) );
  INVX0 U6310_U1 ( .INP(n4441), .ZN(U6310_n1) );
  AND2X1 U6311_U2 ( .IN1(WX2120), .IN2(U6311_n1), .Q(WX2183) );
  INVX0 U6311_U1 ( .INP(n4441), .ZN(U6311_n1) );
  AND2X1 U6312_U2 ( .IN1(WX2118), .IN2(U6312_n1), .Q(WX2181) );
  INVX0 U6312_U1 ( .INP(n4441), .ZN(U6312_n1) );
  AND2X1 U6313_U2 ( .IN1(WX2116), .IN2(U6313_n1), .Q(WX2179) );
  INVX0 U6313_U1 ( .INP(n4440), .ZN(U6313_n1) );
  AND2X1 U6314_U2 ( .IN1(WX2114), .IN2(U6314_n1), .Q(WX2177) );
  INVX0 U6314_U1 ( .INP(n4440), .ZN(U6314_n1) );
  AND2X1 U6315_U2 ( .IN1(WX2112), .IN2(U6315_n1), .Q(WX2175) );
  INVX0 U6315_U1 ( .INP(n4440), .ZN(U6315_n1) );
  AND2X1 U6316_U2 ( .IN1(WX2110), .IN2(U6316_n1), .Q(WX2173) );
  INVX0 U6316_U1 ( .INP(n4440), .ZN(U6316_n1) );
  AND2X1 U6317_U2 ( .IN1(WX2108), .IN2(U6317_n1), .Q(WX2171) );
  INVX0 U6317_U1 ( .INP(n4440), .ZN(U6317_n1) );
  AND2X1 U6318_U2 ( .IN1(WX2106), .IN2(U6318_n1), .Q(WX2169) );
  INVX0 U6318_U1 ( .INP(n4440), .ZN(U6318_n1) );
  AND2X1 U6319_U2 ( .IN1(WX2104), .IN2(U6319_n1), .Q(WX2167) );
  INVX0 U6319_U1 ( .INP(n4440), .ZN(U6319_n1) );
  AND2X1 U6320_U2 ( .IN1(WX2102), .IN2(U6320_n1), .Q(WX2165) );
  INVX0 U6320_U1 ( .INP(n4440), .ZN(U6320_n1) );
  AND2X1 U6321_U2 ( .IN1(test_so17), .IN2(U6321_n1), .Q(WX2163) );
  INVX0 U6321_U1 ( .INP(n4440), .ZN(U6321_n1) );
  AND2X1 U6322_U2 ( .IN1(WX2098), .IN2(U6322_n1), .Q(WX2161) );
  INVX0 U6322_U1 ( .INP(n4440), .ZN(U6322_n1) );
  AND2X1 U6323_U2 ( .IN1(WX2096), .IN2(U6323_n1), .Q(WX2159) );
  INVX0 U6323_U1 ( .INP(n4440), .ZN(U6323_n1) );
  AND2X1 U6324_U2 ( .IN1(WX2094), .IN2(U6324_n1), .Q(WX2157) );
  INVX0 U6324_U1 ( .INP(n4440), .ZN(U6324_n1) );
  AND2X1 U6325_U2 ( .IN1(WX2092), .IN2(U6325_n1), .Q(WX2155) );
  INVX0 U6325_U1 ( .INP(n4440), .ZN(U6325_n1) );
  AND2X1 U6326_U2 ( .IN1(WX2090), .IN2(U6326_n1), .Q(WX2153) );
  INVX0 U6326_U1 ( .INP(n4439), .ZN(U6326_n1) );
  AND2X1 U6327_U2 ( .IN1(WX2088), .IN2(U6327_n1), .Q(WX2151) );
  INVX0 U6327_U1 ( .INP(n4439), .ZN(U6327_n1) );
  AND2X1 U6328_U2 ( .IN1(WX2086), .IN2(U6328_n1), .Q(WX2149) );
  INVX0 U6328_U1 ( .INP(n4439), .ZN(U6328_n1) );
  AND2X1 U6329_U2 ( .IN1(WX2084), .IN2(U6329_n1), .Q(WX2147) );
  INVX0 U6329_U1 ( .INP(n4439), .ZN(U6329_n1) );
  AND2X1 U6330_U2 ( .IN1(WX2082), .IN2(U6330_n1), .Q(WX2145) );
  INVX0 U6330_U1 ( .INP(n4439), .ZN(U6330_n1) );
  AND2X1 U6331_U2 ( .IN1(WX2080), .IN2(U6331_n1), .Q(WX2143) );
  INVX0 U6331_U1 ( .INP(n4439), .ZN(U6331_n1) );
  AND2X1 U6332_U2 ( .IN1(WX2078), .IN2(U6332_n1), .Q(WX2141) );
  INVX0 U6332_U1 ( .INP(n4439), .ZN(U6332_n1) );
  AND2X1 U6333_U2 ( .IN1(WX2076), .IN2(U6333_n1), .Q(WX2139) );
  INVX0 U6333_U1 ( .INP(n4439), .ZN(U6333_n1) );
  AND2X1 U6334_U2 ( .IN1(WX2074), .IN2(U6334_n1), .Q(WX2137) );
  INVX0 U6334_U1 ( .INP(n4439), .ZN(U6334_n1) );
  AND2X1 U6335_U2 ( .IN1(WX2072), .IN2(U6335_n1), .Q(WX2135) );
  INVX0 U6335_U1 ( .INP(n4439), .ZN(U6335_n1) );
  AND2X1 U6336_U2 ( .IN1(WX2070), .IN2(U6336_n1), .Q(WX2133) );
  INVX0 U6336_U1 ( .INP(n4439), .ZN(U6336_n1) );
  AND2X1 U6337_U2 ( .IN1(WX2068), .IN2(U6337_n1), .Q(WX2131) );
  INVX0 U6337_U1 ( .INP(n4439), .ZN(U6337_n1) );
  AND2X1 U6338_U2 ( .IN1(WX2066), .IN2(U6338_n1), .Q(WX2129) );
  INVX0 U6338_U1 ( .INP(n4439), .ZN(U6338_n1) );
  AND2X1 U6339_U2 ( .IN1(test_so16), .IN2(U6339_n1), .Q(WX2127) );
  INVX0 U6339_U1 ( .INP(n4439), .ZN(U6339_n1) );
  AND2X1 U6340_U2 ( .IN1(WX2062), .IN2(U6340_n1), .Q(WX2125) );
  INVX0 U6340_U1 ( .INP(n4438), .ZN(U6340_n1) );
  AND2X1 U6341_U2 ( .IN1(WX2060), .IN2(U6341_n1), .Q(WX2123) );
  INVX0 U6341_U1 ( .INP(n4438), .ZN(U6341_n1) );
  AND2X1 U6342_U2 ( .IN1(WX2058), .IN2(U6342_n1), .Q(WX2121) );
  INVX0 U6342_U1 ( .INP(n4438), .ZN(U6342_n1) );
  AND2X1 U6343_U2 ( .IN1(WX2056), .IN2(U6343_n1), .Q(WX2119) );
  INVX0 U6343_U1 ( .INP(n4438), .ZN(U6343_n1) );
  AND2X1 U6344_U2 ( .IN1(WX2054), .IN2(U6344_n1), .Q(WX2117) );
  INVX0 U6344_U1 ( .INP(n4438), .ZN(U6344_n1) );
  AND2X1 U6345_U2 ( .IN1(WX2052), .IN2(U6345_n1), .Q(WX2115) );
  INVX0 U6345_U1 ( .INP(n4438), .ZN(U6345_n1) );
  AND2X1 U6346_U2 ( .IN1(WX2050), .IN2(U6346_n1), .Q(WX2113) );
  INVX0 U6346_U1 ( .INP(n4438), .ZN(U6346_n1) );
  AND2X1 U6347_U2 ( .IN1(WX2048), .IN2(U6347_n1), .Q(WX2111) );
  INVX0 U6347_U1 ( .INP(n4438), .ZN(U6347_n1) );
  AND2X1 U6348_U2 ( .IN1(WX2046), .IN2(U6348_n1), .Q(WX2109) );
  INVX0 U6348_U1 ( .INP(n4438), .ZN(U6348_n1) );
  AND2X1 U6349_U2 ( .IN1(WX2044), .IN2(U6349_n1), .Q(WX2107) );
  INVX0 U6349_U1 ( .INP(n4438), .ZN(U6349_n1) );
  AND2X1 U6350_U2 ( .IN1(WX2042), .IN2(U6350_n1), .Q(WX2105) );
  INVX0 U6350_U1 ( .INP(n4438), .ZN(U6350_n1) );
  AND2X1 U6351_U2 ( .IN1(WX2040), .IN2(U6351_n1), .Q(WX2103) );
  INVX0 U6351_U1 ( .INP(n4438), .ZN(U6351_n1) );
  AND2X1 U6352_U2 ( .IN1(WX2038), .IN2(U6352_n1), .Q(WX2101) );
  INVX0 U6352_U1 ( .INP(n4438), .ZN(U6352_n1) );
  AND2X1 U6353_U2 ( .IN1(WX2036), .IN2(U6353_n1), .Q(WX2099) );
  INVX0 U6353_U1 ( .INP(n4438), .ZN(U6353_n1) );
  AND2X1 U6354_U2 ( .IN1(WX2034), .IN2(U6354_n1), .Q(WX2097) );
  INVX0 U6354_U1 ( .INP(n4437), .ZN(U6354_n1) );
  AND2X1 U6355_U2 ( .IN1(WX2032), .IN2(U6355_n1), .Q(WX2095) );
  INVX0 U6355_U1 ( .INP(n4437), .ZN(U6355_n1) );
  AND2X1 U6356_U2 ( .IN1(WX2030), .IN2(U6356_n1), .Q(WX2093) );
  INVX0 U6356_U1 ( .INP(n4437), .ZN(U6356_n1) );
  AND2X1 U6357_U2 ( .IN1(test_so15), .IN2(U6357_n1), .Q(WX2091) );
  INVX0 U6357_U1 ( .INP(n4437), .ZN(U6357_n1) );
  AND2X1 U6358_U2 ( .IN1(WX2026), .IN2(U6358_n1), .Q(WX2089) );
  INVX0 U6358_U1 ( .INP(n4437), .ZN(U6358_n1) );
  AND2X1 U6359_U2 ( .IN1(WX2024), .IN2(U6359_n1), .Q(WX2087) );
  INVX0 U6359_U1 ( .INP(n4437), .ZN(U6359_n1) );
  AND2X1 U6360_U2 ( .IN1(WX2022), .IN2(U6360_n1), .Q(WX2085) );
  INVX0 U6360_U1 ( .INP(n4437), .ZN(U6360_n1) );
  AND2X1 U6361_U2 ( .IN1(WX2020), .IN2(U6361_n1), .Q(WX2083) );
  INVX0 U6361_U1 ( .INP(n4437), .ZN(U6361_n1) );
  AND2X1 U6362_U2 ( .IN1(WX2018), .IN2(U6362_n1), .Q(WX2081) );
  INVX0 U6362_U1 ( .INP(n4437), .ZN(U6362_n1) );
  AND2X1 U6363_U2 ( .IN1(WX2016), .IN2(U6363_n1), .Q(WX2079) );
  INVX0 U6363_U1 ( .INP(n4437), .ZN(U6363_n1) );
  AND2X1 U6364_U2 ( .IN1(WX2014), .IN2(U6364_n1), .Q(WX2077) );
  INVX0 U6364_U1 ( .INP(n4437), .ZN(U6364_n1) );
  AND2X1 U6365_U2 ( .IN1(WX2012), .IN2(U6365_n1), .Q(WX2075) );
  INVX0 U6365_U1 ( .INP(n4437), .ZN(U6365_n1) );
  AND2X1 U6366_U2 ( .IN1(WX2010), .IN2(U6366_n1), .Q(WX2073) );
  INVX0 U6366_U1 ( .INP(n4437), .ZN(U6366_n1) );
  AND2X1 U6367_U2 ( .IN1(WX2008), .IN2(U6367_n1), .Q(WX2071) );
  INVX0 U6367_U1 ( .INP(n4437), .ZN(U6367_n1) );
  AND2X1 U6368_U2 ( .IN1(WX2006), .IN2(U6368_n1), .Q(WX2069) );
  INVX0 U6368_U1 ( .INP(n4436), .ZN(U6368_n1) );
  AND2X1 U6369_U2 ( .IN1(WX2004), .IN2(U6369_n1), .Q(WX2067) );
  INVX0 U6369_U1 ( .INP(n4436), .ZN(U6369_n1) );
  AND2X1 U6370_U2 ( .IN1(WX2002), .IN2(U6370_n1), .Q(WX2065) );
  INVX0 U6370_U1 ( .INP(n4436), .ZN(U6370_n1) );
  AND2X1 U6371_U2 ( .IN1(WX2000), .IN2(U6371_n1), .Q(WX2063) );
  INVX0 U6371_U1 ( .INP(n4436), .ZN(U6371_n1) );
  AND2X1 U6372_U2 ( .IN1(WX1998), .IN2(U6372_n1), .Q(WX2061) );
  INVX0 U6372_U1 ( .INP(n4436), .ZN(U6372_n1) );
  AND2X1 U6373_U2 ( .IN1(WX1996), .IN2(U6373_n1), .Q(WX2059) );
  INVX0 U6373_U1 ( .INP(n4436), .ZN(U6373_n1) );
  AND2X1 U6374_U2 ( .IN1(WX1994), .IN2(U6374_n1), .Q(WX2057) );
  INVX0 U6374_U1 ( .INP(n4436), .ZN(U6374_n1) );
  AND2X1 U6375_U2 ( .IN1(test_so14), .IN2(U6375_n1), .Q(WX2055) );
  INVX0 U6375_U1 ( .INP(n4436), .ZN(U6375_n1) );
  AND2X1 U6376_U2 ( .IN1(WX1990), .IN2(U6376_n1), .Q(WX2053) );
  INVX0 U6376_U1 ( .INP(n4436), .ZN(U6376_n1) );
  AND2X1 U6377_U2 ( .IN1(WX1988), .IN2(U6377_n1), .Q(WX2051) );
  INVX0 U6377_U1 ( .INP(n4440), .ZN(U6377_n1) );
  AND2X1 U6378_U2 ( .IN1(WX1986), .IN2(U6378_n1), .Q(WX2049) );
  INVX0 U6378_U1 ( .INP(n4451), .ZN(U6378_n1) );
  AND2X1 U6379_U2 ( .IN1(WX1984), .IN2(U6379_n1), .Q(WX2047) );
  INVX0 U6379_U1 ( .INP(n4451), .ZN(U6379_n1) );
  AND2X1 U6380_U2 ( .IN1(WX1982), .IN2(U6380_n1), .Q(WX2045) );
  INVX0 U6380_U1 ( .INP(n4451), .ZN(U6380_n1) );
  AND2X1 U6381_U2 ( .IN1(WX1980), .IN2(U6381_n1), .Q(WX2043) );
  INVX0 U6381_U1 ( .INP(n4451), .ZN(U6381_n1) );
  AND2X1 U6382_U2 ( .IN1(WX1978), .IN2(U6382_n1), .Q(WX2041) );
  INVX0 U6382_U1 ( .INP(n4451), .ZN(U6382_n1) );
  AND2X1 U6383_U2 ( .IN1(WX1976), .IN2(U6383_n1), .Q(WX2039) );
  INVX0 U6383_U1 ( .INP(n4451), .ZN(U6383_n1) );
  AND2X1 U6384_U2 ( .IN1(WX1974), .IN2(U6384_n1), .Q(WX2037) );
  INVX0 U6384_U1 ( .INP(n4451), .ZN(U6384_n1) );
  AND2X1 U6385_U2 ( .IN1(WX1972), .IN2(U6385_n1), .Q(WX2035) );
  INVX0 U6385_U1 ( .INP(n4451), .ZN(U6385_n1) );
  AND2X1 U6386_U2 ( .IN1(WX1970), .IN2(U6386_n1), .Q(WX2033) );
  INVX0 U6386_U1 ( .INP(n4450), .ZN(U6386_n1) );
  AND2X1 U6387_U2 ( .IN1(WX835), .IN2(U6387_n1), .Q(WX898) );
  INVX0 U6387_U1 ( .INP(n4450), .ZN(U6387_n1) );
  AND2X1 U6388_U2 ( .IN1(WX833), .IN2(U6388_n1), .Q(WX896) );
  INVX0 U6388_U1 ( .INP(n4450), .ZN(U6388_n1) );
  AND2X1 U6389_U2 ( .IN1(test_so7), .IN2(U6389_n1), .Q(WX894) );
  INVX0 U6389_U1 ( .INP(n4450), .ZN(U6389_n1) );
  AND2X1 U6390_U2 ( .IN1(WX829), .IN2(U6390_n1), .Q(WX892) );
  INVX0 U6390_U1 ( .INP(n4450), .ZN(U6390_n1) );
  AND2X1 U6391_U2 ( .IN1(WX827), .IN2(U6391_n1), .Q(WX890) );
  INVX0 U6391_U1 ( .INP(n4450), .ZN(U6391_n1) );
  AND2X1 U6392_U2 ( .IN1(WX825), .IN2(U6392_n1), .Q(WX888) );
  INVX0 U6392_U1 ( .INP(n4450), .ZN(U6392_n1) );
  AND2X1 U6393_U2 ( .IN1(WX823), .IN2(U6393_n1), .Q(WX886) );
  INVX0 U6393_U1 ( .INP(n4450), .ZN(U6393_n1) );
  AND2X1 U6394_U2 ( .IN1(WX821), .IN2(U6394_n1), .Q(WX884) );
  INVX0 U6394_U1 ( .INP(n4450), .ZN(U6394_n1) );
  AND2X1 U6395_U2 ( .IN1(WX819), .IN2(U6395_n1), .Q(WX882) );
  INVX0 U6395_U1 ( .INP(n4450), .ZN(U6395_n1) );
  AND2X1 U6396_U2 ( .IN1(WX817), .IN2(U6396_n1), .Q(WX880) );
  INVX0 U6396_U1 ( .INP(n4450), .ZN(U6396_n1) );
  AND2X1 U6397_U2 ( .IN1(WX815), .IN2(U6397_n1), .Q(WX878) );
  INVX0 U6397_U1 ( .INP(n4450), .ZN(U6397_n1) );
  AND2X1 U6398_U2 ( .IN1(WX813), .IN2(U6398_n1), .Q(WX876) );
  INVX0 U6398_U1 ( .INP(n4450), .ZN(U6398_n1) );
  AND2X1 U6399_U2 ( .IN1(WX811), .IN2(U6399_n1), .Q(WX874) );
  INVX0 U6399_U1 ( .INP(n4450), .ZN(U6399_n1) );
  AND2X1 U6400_U2 ( .IN1(WX809), .IN2(U6400_n1), .Q(WX872) );
  INVX0 U6400_U1 ( .INP(n4449), .ZN(U6400_n1) );
  AND2X1 U6401_U2 ( .IN1(WX807), .IN2(U6401_n1), .Q(WX870) );
  INVX0 U6401_U1 ( .INP(n4449), .ZN(U6401_n1) );
  AND2X1 U6402_U2 ( .IN1(WX805), .IN2(U6402_n1), .Q(WX868) );
  INVX0 U6402_U1 ( .INP(n4449), .ZN(U6402_n1) );
  AND2X1 U6403_U2 ( .IN1(WX803), .IN2(U6403_n1), .Q(WX866) );
  INVX0 U6403_U1 ( .INP(n4449), .ZN(U6403_n1) );
  AND2X1 U6404_U2 ( .IN1(WX801), .IN2(U6404_n1), .Q(WX864) );
  INVX0 U6404_U1 ( .INP(n4449), .ZN(U6404_n1) );
  AND2X1 U6405_U2 ( .IN1(WX799), .IN2(U6405_n1), .Q(WX862) );
  INVX0 U6405_U1 ( .INP(n4449), .ZN(U6405_n1) );
  AND2X1 U6406_U2 ( .IN1(WX797), .IN2(U6406_n1), .Q(WX860) );
  INVX0 U6406_U1 ( .INP(n4449), .ZN(U6406_n1) );
  AND2X1 U6407_U2 ( .IN1(test_so6), .IN2(U6407_n1), .Q(WX858) );
  INVX0 U6407_U1 ( .INP(n4449), .ZN(U6407_n1) );
  AND2X1 U6408_U2 ( .IN1(WX793), .IN2(U6408_n1), .Q(WX856) );
  INVX0 U6408_U1 ( .INP(n4449), .ZN(U6408_n1) );
  AND2X1 U6409_U2 ( .IN1(WX791), .IN2(U6409_n1), .Q(WX854) );
  INVX0 U6409_U1 ( .INP(n4449), .ZN(U6409_n1) );
  AND2X1 U6410_U2 ( .IN1(WX789), .IN2(U6410_n1), .Q(WX852) );
  INVX0 U6410_U1 ( .INP(n4449), .ZN(U6410_n1) );
  AND2X1 U6411_U2 ( .IN1(WX787), .IN2(U6411_n1), .Q(WX850) );
  INVX0 U6411_U1 ( .INP(n4449), .ZN(U6411_n1) );
  AND2X1 U6412_U2 ( .IN1(WX785), .IN2(U6412_n1), .Q(WX848) );
  INVX0 U6412_U1 ( .INP(n4449), .ZN(U6412_n1) );
  AND2X1 U6413_U2 ( .IN1(WX783), .IN2(U6413_n1), .Q(WX846) );
  INVX0 U6413_U1 ( .INP(n4449), .ZN(U6413_n1) );
  AND2X1 U6414_U2 ( .IN1(WX781), .IN2(U6414_n1), .Q(WX844) );
  INVX0 U6414_U1 ( .INP(n4448), .ZN(U6414_n1) );
  AND2X1 U6415_U2 ( .IN1(WX779), .IN2(U6415_n1), .Q(WX842) );
  INVX0 U6415_U1 ( .INP(n4448), .ZN(U6415_n1) );
  AND2X1 U6416_U2 ( .IN1(WX777), .IN2(U6416_n1), .Q(WX840) );
  INVX0 U6416_U1 ( .INP(n4448), .ZN(U6416_n1) );
  AND2X1 U6417_U2 ( .IN1(WX775), .IN2(U6417_n1), .Q(WX838) );
  INVX0 U6417_U1 ( .INP(n4448), .ZN(U6417_n1) );
  AND2X1 U6418_U2 ( .IN1(WX773), .IN2(U6418_n1), .Q(WX836) );
  INVX0 U6418_U1 ( .INP(n4448), .ZN(U6418_n1) );
  AND2X1 U6419_U2 ( .IN1(WX771), .IN2(U6419_n1), .Q(WX834) );
  INVX0 U6419_U1 ( .INP(n4448), .ZN(U6419_n1) );
  AND2X1 U6420_U2 ( .IN1(WX769), .IN2(U6420_n1), .Q(WX832) );
  INVX0 U6420_U1 ( .INP(n4448), .ZN(U6420_n1) );
  AND2X1 U6421_U2 ( .IN1(WX767), .IN2(U6421_n1), .Q(WX830) );
  INVX0 U6421_U1 ( .INP(n4448), .ZN(U6421_n1) );
  AND2X1 U6422_U2 ( .IN1(WX765), .IN2(U6422_n1), .Q(WX828) );
  INVX0 U6422_U1 ( .INP(n4448), .ZN(U6422_n1) );
  AND2X1 U6423_U2 ( .IN1(WX763), .IN2(U6423_n1), .Q(WX826) );
  INVX0 U6423_U1 ( .INP(n4448), .ZN(U6423_n1) );
  AND2X1 U6424_U2 ( .IN1(WX761), .IN2(U6424_n1), .Q(WX824) );
  INVX0 U6424_U1 ( .INP(n4448), .ZN(U6424_n1) );
  AND2X1 U6425_U2 ( .IN1(test_so5), .IN2(U6425_n1), .Q(WX822) );
  INVX0 U6425_U1 ( .INP(n4448), .ZN(U6425_n1) );
  AND2X1 U6426_U2 ( .IN1(WX757), .IN2(U6426_n1), .Q(WX820) );
  INVX0 U6426_U1 ( .INP(n4448), .ZN(U6426_n1) );
  AND2X1 U6427_U2 ( .IN1(WX755), .IN2(U6427_n1), .Q(WX818) );
  INVX0 U6427_U1 ( .INP(n4448), .ZN(U6427_n1) );
  AND2X1 U6428_U2 ( .IN1(WX753), .IN2(U6428_n1), .Q(WX816) );
  INVX0 U6428_U1 ( .INP(n4447), .ZN(U6428_n1) );
  AND2X1 U6429_U2 ( .IN1(WX751), .IN2(U6429_n1), .Q(WX814) );
  INVX0 U6429_U1 ( .INP(n4447), .ZN(U6429_n1) );
  AND2X1 U6430_U2 ( .IN1(WX749), .IN2(U6430_n1), .Q(WX812) );
  INVX0 U6430_U1 ( .INP(n4447), .ZN(U6430_n1) );
  AND2X1 U6431_U2 ( .IN1(WX747), .IN2(U6431_n1), .Q(WX810) );
  INVX0 U6431_U1 ( .INP(n4447), .ZN(U6431_n1) );
  AND2X1 U6432_U2 ( .IN1(WX745), .IN2(U6432_n1), .Q(WX808) );
  INVX0 U6432_U1 ( .INP(n4447), .ZN(U6432_n1) );
  AND2X1 U6433_U2 ( .IN1(WX743), .IN2(U6433_n1), .Q(WX806) );
  INVX0 U6433_U1 ( .INP(n4447), .ZN(U6433_n1) );
  AND2X1 U6434_U2 ( .IN1(WX741), .IN2(U6434_n1), .Q(WX804) );
  INVX0 U6434_U1 ( .INP(n4447), .ZN(U6434_n1) );
  AND2X1 U6435_U2 ( .IN1(WX739), .IN2(U6435_n1), .Q(WX802) );
  INVX0 U6435_U1 ( .INP(n4447), .ZN(U6435_n1) );
  AND2X1 U6436_U2 ( .IN1(WX737), .IN2(U6436_n1), .Q(WX800) );
  INVX0 U6436_U1 ( .INP(n4447), .ZN(U6436_n1) );
  AND2X1 U6437_U2 ( .IN1(WX735), .IN2(U6437_n1), .Q(WX798) );
  INVX0 U6437_U1 ( .INP(n4447), .ZN(U6437_n1) );
  AND2X1 U6438_U2 ( .IN1(WX733), .IN2(U6438_n1), .Q(WX796) );
  INVX0 U6438_U1 ( .INP(n4447), .ZN(U6438_n1) );
  AND2X1 U6439_U2 ( .IN1(WX731), .IN2(U6439_n1), .Q(WX794) );
  INVX0 U6439_U1 ( .INP(n4447), .ZN(U6439_n1) );
  AND2X1 U6440_U2 ( .IN1(WX729), .IN2(U6440_n1), .Q(WX792) );
  INVX0 U6440_U1 ( .INP(n4447), .ZN(U6440_n1) );
  AND2X1 U6441_U2 ( .IN1(WX727), .IN2(U6441_n1), .Q(WX790) );
  INVX0 U6441_U1 ( .INP(n4446), .ZN(U6441_n1) );
  AND2X1 U6442_U2 ( .IN1(WX725), .IN2(U6442_n1), .Q(WX788) );
  INVX0 U6442_U1 ( .INP(n4446), .ZN(U6442_n1) );
  AND2X1 U6443_U2 ( .IN1(test_so4), .IN2(U6443_n1), .Q(WX786) );
  INVX0 U6443_U1 ( .INP(n4446), .ZN(U6443_n1) );
  AND2X1 U6444_U2 ( .IN1(WX721), .IN2(U6444_n1), .Q(WX784) );
  INVX0 U6444_U1 ( .INP(n4446), .ZN(U6444_n1) );
  AND2X1 U6445_U2 ( .IN1(WX719), .IN2(U6445_n1), .Q(WX782) );
  INVX0 U6445_U1 ( .INP(n4446), .ZN(U6445_n1) );
  AND2X1 U6446_U2 ( .IN1(WX717), .IN2(U6446_n1), .Q(WX780) );
  INVX0 U6446_U1 ( .INP(n4446), .ZN(U6446_n1) );
  AND2X1 U6447_U2 ( .IN1(WX715), .IN2(U6447_n1), .Q(WX778) );
  INVX0 U6447_U1 ( .INP(n4446), .ZN(U6447_n1) );
  AND2X1 U6448_U2 ( .IN1(WX713), .IN2(U6448_n1), .Q(WX776) );
  INVX0 U6448_U1 ( .INP(n4446), .ZN(U6448_n1) );
  AND2X1 U6449_U2 ( .IN1(WX711), .IN2(U6449_n1), .Q(WX774) );
  INVX0 U6449_U1 ( .INP(n4446), .ZN(U6449_n1) );
  AND2X1 U6450_U2 ( .IN1(WX709), .IN2(U6450_n1), .Q(WX772) );
  INVX0 U6450_U1 ( .INP(n4446), .ZN(U6450_n1) );
  AND2X1 U6451_U2 ( .IN1(WX707), .IN2(U6451_n1), .Q(WX770) );
  INVX0 U6451_U1 ( .INP(n4446), .ZN(U6451_n1) );
  AND2X1 U6452_U2 ( .IN1(WX705), .IN2(U6452_n1), .Q(WX768) );
  INVX0 U6452_U1 ( .INP(n4446), .ZN(U6452_n1) );
  AND2X1 U6453_U2 ( .IN1(WX703), .IN2(U6453_n1), .Q(WX766) );
  INVX0 U6453_U1 ( .INP(n4446), .ZN(U6453_n1) );
  AND2X1 U6454_U2 ( .IN1(WX701), .IN2(U6454_n1), .Q(WX764) );
  INVX0 U6454_U1 ( .INP(n4446), .ZN(U6454_n1) );
  AND2X1 U6455_U2 ( .IN1(WX699), .IN2(U6455_n1), .Q(WX762) );
  INVX0 U6455_U1 ( .INP(n4445), .ZN(U6455_n1) );
  AND2X1 U6456_U2 ( .IN1(WX697), .IN2(U6456_n1), .Q(WX760) );
  INVX0 U6456_U1 ( .INP(n4445), .ZN(U6456_n1) );
  AND2X1 U6457_U2 ( .IN1(WX695), .IN2(U6457_n1), .Q(WX758) );
  INVX0 U6457_U1 ( .INP(n4445), .ZN(U6457_n1) );
  AND2X1 U6458_U2 ( .IN1(WX693), .IN2(U6458_n1), .Q(WX756) );
  INVX0 U6458_U1 ( .INP(n4445), .ZN(U6458_n1) );
  AND2X1 U6459_U2 ( .IN1(WX691), .IN2(U6459_n1), .Q(WX754) );
  INVX0 U6459_U1 ( .INP(n4445), .ZN(U6459_n1) );
  AND2X1 U6460_U2 ( .IN1(WX689), .IN2(U6460_n1), .Q(WX752) );
  INVX0 U6460_U1 ( .INP(n4445), .ZN(U6460_n1) );
  AND2X1 U6461_U2 ( .IN1(test_so3), .IN2(U6461_n1), .Q(WX750) );
  INVX0 U6461_U1 ( .INP(n4445), .ZN(U6461_n1) );
  AND2X1 U6462_U2 ( .IN1(WX685), .IN2(U6462_n1), .Q(WX748) );
  INVX0 U6462_U1 ( .INP(n4445), .ZN(U6462_n1) );
  AND2X1 U6463_U2 ( .IN1(WX683), .IN2(U6463_n1), .Q(WX746) );
  INVX0 U6463_U1 ( .INP(n4445), .ZN(U6463_n1) );
  AND2X1 U6464_U2 ( .IN1(WX681), .IN2(U6464_n1), .Q(WX744) );
  INVX0 U6464_U1 ( .INP(n4445), .ZN(U6464_n1) );
  AND2X1 U6465_U2 ( .IN1(WX679), .IN2(U6465_n1), .Q(WX742) );
  INVX0 U6465_U1 ( .INP(n4445), .ZN(U6465_n1) );
  AND2X1 U6466_U2 ( .IN1(WX677), .IN2(U6466_n1), .Q(WX740) );
  INVX0 U6466_U1 ( .INP(n4445), .ZN(U6466_n1) );
  AND2X1 U6467_U2 ( .IN1(WX675), .IN2(U6467_n1), .Q(WX738) );
  INVX0 U6467_U1 ( .INP(n4445), .ZN(U6467_n1) );
  AND2X1 U6468_U2 ( .IN1(WX673), .IN2(U6468_n1), .Q(WX736) );
  INVX0 U6468_U1 ( .INP(n4445), .ZN(U6468_n1) );
  AND2X1 U6469_U2 ( .IN1(WX671), .IN2(U6469_n1), .Q(WX734) );
  INVX0 U6469_U1 ( .INP(n4444), .ZN(U6469_n1) );
  AND2X1 U6470_U2 ( .IN1(WX669), .IN2(U6470_n1), .Q(WX732) );
  INVX0 U6470_U1 ( .INP(n4444), .ZN(U6470_n1) );
  AND2X1 U6471_U2 ( .IN1(WX667), .IN2(U6471_n1), .Q(WX730) );
  INVX0 U6471_U1 ( .INP(n4444), .ZN(U6471_n1) );
  AND2X1 U6472_U2 ( .IN1(WX665), .IN2(U6472_n1), .Q(WX728) );
  INVX0 U6472_U1 ( .INP(n4444), .ZN(U6472_n1) );
  AND2X1 U6473_U2 ( .IN1(WX663), .IN2(U6473_n1), .Q(WX726) );
  INVX0 U6473_U1 ( .INP(n4444), .ZN(U6473_n1) );
  AND2X1 U6474_U2 ( .IN1(WX661), .IN2(U6474_n1), .Q(WX724) );
  INVX0 U6474_U1 ( .INP(n4444), .ZN(U6474_n1) );
  AND2X1 U6475_U2 ( .IN1(WX659), .IN2(U6475_n1), .Q(WX722) );
  INVX0 U6475_U1 ( .INP(n4444), .ZN(U6475_n1) );
  AND2X1 U6476_U2 ( .IN1(WX657), .IN2(U6476_n1), .Q(WX720) );
  INVX0 U6476_U1 ( .INP(n4444), .ZN(U6476_n1) );
  AND2X1 U6477_U2 ( .IN1(WX655), .IN2(U6477_n1), .Q(WX718) );
  INVX0 U6477_U1 ( .INP(n4444), .ZN(U6477_n1) );
  AND2X1 U6478_U2 ( .IN1(WX653), .IN2(U6478_n1), .Q(WX716) );
  INVX0 U6478_U1 ( .INP(n4444), .ZN(U6478_n1) );
  AND2X1 U6479_U2 ( .IN1(test_so2), .IN2(U6479_n1), .Q(WX714) );
  INVX0 U6479_U1 ( .INP(n4444), .ZN(U6479_n1) );
  AND2X1 U6480_U2 ( .IN1(WX649), .IN2(U6480_n1), .Q(WX712) );
  INVX0 U6480_U1 ( .INP(n4444), .ZN(U6480_n1) );
  AND2X1 U6481_U2 ( .IN1(WX647), .IN2(U6481_n1), .Q(WX710) );
  INVX0 U6481_U1 ( .INP(n4444), .ZN(U6481_n1) );
  AND2X1 U6482_U2 ( .IN1(WX645), .IN2(U6482_n1), .Q(WX708) );
  INVX0 U6482_U1 ( .INP(n4444), .ZN(U6482_n1) );
endmodule

