module rs232 ( sys_clk, sys_rst_l, uart_XMIT_dataH, xmitH, xmit_dataH_7_, 
        xmit_dataH_6_, xmit_dataH_5_, xmit_dataH_4_, xmit_dataH_3_, 
        xmit_dataH_2_, xmit_dataH_1_, xmit_dataH_0_, xmit_doneH, 
        uart_REC_dataH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_, rec_dataH_4_, 
        rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_, rec_readyH, 
        test_mode, test_se, test_si, test_so );
  input sys_clk, sys_rst_l, xmitH, xmit_dataH_7_, xmit_dataH_6_, xmit_dataH_5_,
         xmit_dataH_4_, xmit_dataH_3_, xmit_dataH_2_, xmit_dataH_1_,
         xmit_dataH_0_, uart_REC_dataH, test_mode, test_se, test_si;
  output uart_XMIT_dataH, xmit_doneH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_,
         rec_dataH_4_, rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_,
         rec_readyH, test_so;
  wire   rec_dataH_temp_6, rec_dataH_temp_5, rec_dataH_temp_4,
         rec_dataH_temp_3, rec_dataH_temp_2, rec_dataH_temp_1,
         rec_dataH_temp_0, iCTRL, xmit_doneH_temp, iXMIT_CRTL, iRECEIVER_CTRL,
         iRECEIVER_state_CTRL, iRECEIVER_bitCell_CTRL, n400, n401, n402, n403,
         iRECEIVER_next_state_2_, iRECEIVER_state_0_, iRECEIVER_state_1_,
         iRECEIVER_state_2_, iXMIT_state_CTRL, iXMIT_N_CTRL_1_,
         iXMIT_N_CTRL_2_, iXMIT_xmit_CTRL, iXMIT_N24, iXMIT_xmit_ShiftRegH_7_,
         iXMIT_xmit_ShiftRegH_6_, iXMIT_xmit_ShiftRegH_5_, iXMIT_N28,
         iXMIT_N27, iXMIT_N26, iXMIT_N25, iXMIT_N46, iXMIT_N45, iXMIT_N44,
         iXMIT_N29, iXMIT_state_0_, iXMIT_state_1_, iXMIT_state_2_, n241, n245,
         n238, n242, n246, n239, rec_dataH_rec_7, rec_dataH_rec_6,
         rec_dataH_rec_5, rec_dataH_rec_4, rec_dataH_rec_3, rec_dataH_rec_2,
         rec_dataH_rec_1, rec_dataH_rec_0, n370, n371, n187, n186, n185, n184,
         n183, n182, n181, n180, n179, n178, n177, n176, n175, n174, n173,
         n172, n171, n170, n169, n168, n167, n166, n164, n163, n162, n161,
         test_point_DOUT, n160, n159, n157, n156, n155, n154, n153, n152, n150,
         n149, n148, n147, n146, n145, n143, n142, n141, n140, n139, n138,
         n136, n135, n134, n133, n132, n131, n129, n128, n127, n126, n125,
         n124, n397, n398, n399, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705;

  AND2X4 TrojanU303 ( .IN1(iCTRL), .IN2(xmit_doneH_temp), .Q(xmit_doneH) );
  OR2X1 TrojanU302 ( .IN1(iXMIT_CRTL), .IN2(iRECEIVER_CTRL), .Q(iCTRL) );
  OR2X1 TrojanU301 ( .IN1(iRECEIVER_state_CTRL), .IN2(iRECEIVER_bitCell_CTRL), 
        .Q(iRECEIVER_CTRL) );
  NAND4X1 TrojanU300 ( .IN1(n400), .IN2(n401), .IN3(n402), .IN4(n403), .QN(
        iRECEIVER_bitCell_CTRL) );
  NAND4X1 TrojanU297 ( .IN1(iRECEIVER_next_state_2_), .IN2(iRECEIVER_state_0_), 
        .IN3(iRECEIVER_state_1_), .IN4(iRECEIVER_state_2_), .QN(
        iRECEIVER_state_CTRL) );
  OR4X4 TrojanU296 ( .IN1(iXMIT_state_CTRL), .IN2(iXMIT_N_CTRL_1_), .IN3(
        iXMIT_N_CTRL_2_), .IN4(iXMIT_xmit_CTRL), .Q(iXMIT_CRTL) );
  NAND4X1 TrojanU295 ( .IN1(iXMIT_N24), .IN2(iXMIT_xmit_ShiftRegH_7_), .IN3(
        iXMIT_xmit_ShiftRegH_6_), .IN4(iXMIT_xmit_ShiftRegH_5_), .QN(
        iXMIT_xmit_CTRL) );
  NAND4X1 TrojanU294 ( .IN1(iXMIT_N28), .IN2(iXMIT_N27), .IN3(iXMIT_N26), 
        .IN4(iXMIT_N25), .QN(iXMIT_N_CTRL_2_) );
  NAND4X1 TrojanU293 ( .IN1(iXMIT_N46), .IN2(iXMIT_N45), .IN3(iXMIT_N44), 
        .IN4(iXMIT_N29), .QN(iXMIT_N_CTRL_1_) );
  NAND4X1 TrojanU292 ( .IN1(n397), .IN2(iXMIT_state_0_), .IN3(iXMIT_state_1_), 
        .IN4(iXMIT_state_2_), .QN(iXMIT_state_CTRL) );
  INVX32 TrojanU290 ( .INP(n370), .ZN(n371) );
  NAND2X4 TrojanU289 ( .IN1(1'b1), .IN2(test_mode), .QN(n370) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_2_ ( .D(n187), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n700) );
  DFFARX1 iXMIT_state_reg_0_ ( .D(n186), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_0_), .QN(n239) );
  DFFARX1 iXMIT_state_reg_2_ ( .D(n185), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_2_), .QN(n242) );
  DFFARX1 iXMIT_state_reg_1_ ( .D(n184), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_1_), .QN(n246) );
  DFFARX1 iXMIT_bitCountH_reg_0_ ( .D(n183), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n697), .QN(n398) );
  DFFARX1 iXMIT_bitCountH_reg_1_ ( .D(n182), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n698), .QN(n405) );
  DFFARX1 iXMIT_bitCountH_reg_2_ ( .D(n181), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n696), .QN(n410) );
  DFFARX1 iXMIT_bitCountH_reg_3_ ( .D(n180), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n695) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_7_ ( .D(n179), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_7_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_6_ ( .D(n178), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_6_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_5_ ( .D(n177), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_5_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_4_ ( .D(n176), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n684) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_3_ ( .D(n175), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n685) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_2_ ( .D(n174), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n686) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_1_ ( .D(n173), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n687) );
  DFFARX1 iXMIT_xmit_doneH_reg ( .D(n172), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(xmit_doneH_temp) );
  DFFARX1 iRECEIVER_state_reg_1_ ( .D(n171), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_1_), .QN(n241) );
  DFFASX1 iRECEIVER_state_reg_0_ ( .D(n170), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(iRECEIVER_state_0_), .QN(n245) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_0_ ( .D(n169), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n690), .QN(n399) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_1_ ( .D(n168), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n705), .QN(n407) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_2_ ( .D(n167), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n703) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_3_ ( .D(n166), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n704), .QN(n414) );
  DFFARX1 iRECEIVER_state_reg_2_ ( .D(n164), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_2_), .QN(n238) );
  DFFARX1 iRECEIVER_rec_readyH_reg ( .D(n163), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(rec_readyH) );
  DFFARX1 iRECEIVER_par_dataH_reg_7_ ( .D(n162), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_7) );
  DFFARX1 rec_dataH_temp_reg_7_ ( .D(n161), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(test_so) );
  DFFARX1 rec_dataH_reg_7_ ( .D(n160), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_7_) );
  DFFARX1 iRECEIVER_par_dataH_reg_6_ ( .D(n159), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_6) );
  DFFARX1 rec_dataH_temp_reg_6_ ( .D(n157), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_6) );
  DFFARX1 rec_dataH_reg_6_ ( .D(n156), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_6_) );
  DFFARX1 iRECEIVER_par_dataH_reg_5_ ( .D(n155), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_5) );
  DFFARX1 rec_dataH_temp_reg_5_ ( .D(n154), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_5) );
  DFFARX1 rec_dataH_reg_5_ ( .D(n153), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_5_) );
  DFFARX1 iRECEIVER_par_dataH_reg_4_ ( .D(n152), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_4) );
  DFFARX1 rec_dataH_temp_reg_4_ ( .D(n150), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_4) );
  DFFARX1 rec_dataH_reg_4_ ( .D(n149), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_4_) );
  DFFARX1 iRECEIVER_par_dataH_reg_3_ ( .D(n148), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_3) );
  DFFARX1 rec_dataH_temp_reg_3_ ( .D(n147), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_3) );
  DFFARX1 rec_dataH_reg_3_ ( .D(n146), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_3_) );
  DFFARX1 iRECEIVER_par_dataH_reg_2_ ( .D(n145), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_2) );
  DFFARX1 rec_dataH_temp_reg_2_ ( .D(n143), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_2) );
  DFFARX1 rec_dataH_reg_2_ ( .D(n142), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_2_) );
  DFFARX1 iRECEIVER_par_dataH_reg_1_ ( .D(n141), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_1) );
  DFFARX1 rec_dataH_temp_reg_1_ ( .D(n140), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_1) );
  DFFARX1 rec_dataH_reg_1_ ( .D(n139), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_1_) );
  DFFARX1 iRECEIVER_par_dataH_reg_0_ ( .D(n138), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_0) );
  DFFARX1 rec_dataH_temp_reg_0_ ( .D(n136), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_0) );
  DFFARX1 rec_dataH_reg_0_ ( .D(n135), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_0_) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_3_ ( .D(n134), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n691), .QN(n416) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_0_ ( .D(n133), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n693), .QN(n404) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_1_ ( .D(n132), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n692), .QN(n406) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_2_ ( .D(n131), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n694), .QN(n409) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_3_ ( .D(n129), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n699), .QN(n411) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_0_ ( .D(n128), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n702), .QN(n413) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_1_ ( .D(n127), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n701), .QN(n415) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_0_ ( .D(n126), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n408) );
  DFFASX1 iRECEIVER_rec_datSyncH_reg ( .D(n125), .CLK(sys_clk), .SETB(
        sys_rst_l), .Q(n688) );
  DFFASX1 iRECEIVER_rec_datH_reg ( .D(n124), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(n689), .QN(n412) );
  DFFARX1 TrojaniDatasend_reg_1 ( .D(n127), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n400) );
  DFFARX1 TrojaniDatasend_reg_2 ( .D(n126), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n401) );
  DFFASX1 TrojaniDatasend_reg_3 ( .D(n125), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(n402) );
  DFFASX1 TrojaniDatasend_reg_4 ( .D(n124), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(n403) );
  MUX21X2 TrojanU291 ( .IN1(rec_readyH), .IN2(sys_clk), .S(n371), .Q(
        test_point_DOUT) );
  OR3X1 U545 ( .IN1(n417), .IN2(n418), .IN3(n419), .Q(uart_XMIT_dataH) );
  AND2X1 U546 ( .IN1(n246), .IN2(n242), .Q(n419) );
  AND2X1 U547 ( .IN1(n420), .IN2(n408), .Q(n418) );
  OR2X1 U548 ( .IN1(iXMIT_state_0_), .IN2(iXMIT_state_2_), .Q(n420) );
  OR2X1 U549 ( .IN1(n421), .IN2(n422), .Q(n187) );
  AND2X1 U550 ( .IN1(test_se), .IN2(n701), .Q(n422) );
  AND2X1 U551 ( .IN1(iXMIT_N28), .IN2(n423), .Q(n421) );
  OR2X1 U552 ( .IN1(n424), .IN2(n425), .Q(n186) );
  AND2X1 U553 ( .IN1(n426), .IN2(n423), .Q(n425) );
  OR2X1 U554 ( .IN1(n427), .IN2(n428), .Q(n426) );
  AND3X1 U555 ( .IN1(n429), .IN2(iXMIT_state_1_), .IN3(n430), .Q(n428) );
  OR2X1 U556 ( .IN1(n431), .IN2(iXMIT_state_0_), .Q(n430) );
  AND2X1 U557 ( .IN1(n432), .IN2(iXMIT_state_2_), .Q(n427) );
  OR2X1 U558 ( .IN1(n239), .IN2(n433), .Q(n432) );
  AND2X1 U559 ( .IN1(n695), .IN2(test_se), .Q(n424) );
  OR2X1 U560 ( .IN1(n434), .IN2(n435), .Q(n185) );
  AND2X1 U561 ( .IN1(n397), .IN2(n423), .Q(n435) );
  OR2X1 U562 ( .IN1(n436), .IN2(n437), .Q(n397) );
  AND2X1 U563 ( .IN1(n438), .IN2(iXMIT_state_1_), .Q(n437) );
  INVX0 U564 ( .INP(n439), .ZN(n438) );
  AND2X1 U565 ( .IN1(n417), .IN2(n433), .Q(n436) );
  AND2X1 U566 ( .IN1(test_se), .IN2(iXMIT_state_1_), .Q(n434) );
  OR2X1 U567 ( .IN1(n440), .IN2(n441), .Q(n184) );
  AND2X1 U568 ( .IN1(n442), .IN2(n423), .Q(n441) );
  OR2X1 U569 ( .IN1(n443), .IN2(n444), .Q(n442) );
  AND2X1 U570 ( .IN1(test_se), .IN2(iXMIT_state_0_), .Q(n440) );
  OR3X1 U571 ( .IN1(n445), .IN2(n446), .IN3(n447), .Q(n183) );
  AND2X1 U572 ( .IN1(test_se), .IN2(n699), .Q(n447) );
  AND2X1 U573 ( .IN1(n697), .IN2(n448), .Q(n446) );
  OR2X1 U574 ( .IN1(n449), .IN2(n450), .Q(n182) );
  AND2X1 U575 ( .IN1(n697), .IN2(n451), .Q(n450) );
  OR2X1 U576 ( .IN1(n452), .IN2(test_se), .Q(n451) );
  AND2X1 U577 ( .IN1(n453), .IN2(n405), .Q(n452) );
  AND2X1 U578 ( .IN1(n698), .IN2(n454), .Q(n449) );
  OR2X1 U579 ( .IN1(n445), .IN2(n448), .Q(n454) );
  AND2X1 U580 ( .IN1(n398), .IN2(n455), .Q(n445) );
  OR3X1 U581 ( .IN1(n456), .IN2(n457), .IN3(n458), .Q(n181) );
  AND2X1 U582 ( .IN1(n698), .IN2(test_se), .Q(n458) );
  AND2X1 U583 ( .IN1(n696), .IN2(n448), .Q(n457) );
  AND2X1 U584 ( .IN1(iXMIT_N45), .IN2(n455), .Q(n456) );
  OR3X1 U585 ( .IN1(n459), .IN2(n460), .IN3(n461), .Q(n180) );
  AND2X1 U586 ( .IN1(n696), .IN2(test_se), .Q(n461) );
  AND2X1 U587 ( .IN1(n448), .IN2(n695), .Q(n460) );
  AND3X1 U588 ( .IN1(n423), .IN2(n462), .IN3(n463), .Q(n448) );
  AND2X1 U589 ( .IN1(n455), .IN2(iXMIT_N46), .Q(n459) );
  AND2X1 U590 ( .IN1(n423), .IN2(n453), .Q(n455) );
  INVX0 U591 ( .INP(n462), .ZN(n453) );
  OR3X1 U592 ( .IN1(n246), .IN2(n239), .IN3(n429), .Q(n462) );
  OR2X1 U593 ( .IN1(n464), .IN2(n465), .Q(n429) );
  AND4X1 U594 ( .IN1(n695), .IN2(n405), .IN3(n398), .IN4(n410), .Q(n464) );
  OR2X1 U595 ( .IN1(n466), .IN2(n467), .Q(n179) );
  AND2X1 U596 ( .IN1(n468), .IN2(n423), .Q(n467) );
  OR3X1 U597 ( .IN1(n469), .IN2(n470), .IN3(n471), .Q(n468) );
  AND2X1 U598 ( .IN1(xmit_dataH_7_), .IN2(n444), .Q(n470) );
  AND2X1 U599 ( .IN1(n472), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n469) );
  AND2X1 U600 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n466) );
  OR2X1 U601 ( .IN1(n473), .IN2(n474), .Q(n178) );
  AND2X1 U602 ( .IN1(n475), .IN2(n423), .Q(n474) );
  OR3X1 U603 ( .IN1(n476), .IN2(n477), .IN3(n478), .Q(n475) );
  AND2X1 U604 ( .IN1(xmit_dataH_6_), .IN2(n479), .Q(n478) );
  AND2X1 U605 ( .IN1(n472), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n477) );
  AND2X1 U606 ( .IN1(n471), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n476) );
  AND2X1 U607 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n473) );
  OR2X1 U608 ( .IN1(n480), .IN2(n481), .Q(n177) );
  AND2X1 U609 ( .IN1(n482), .IN2(n423), .Q(n481) );
  OR3X1 U610 ( .IN1(n483), .IN2(n484), .IN3(n485), .Q(n482) );
  AND2X1 U611 ( .IN1(xmit_dataH_5_), .IN2(n479), .Q(n485) );
  AND2X1 U612 ( .IN1(n472), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n484) );
  AND2X1 U613 ( .IN1(n471), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n483) );
  AND2X1 U614 ( .IN1(n684), .IN2(test_se), .Q(n480) );
  OR2X1 U615 ( .IN1(n486), .IN2(n487), .Q(n176) );
  AND2X1 U616 ( .IN1(n488), .IN2(n423), .Q(n487) );
  OR3X1 U617 ( .IN1(n489), .IN2(n490), .IN3(n491), .Q(n488) );
  AND2X1 U618 ( .IN1(xmit_dataH_4_), .IN2(n479), .Q(n491) );
  AND2X1 U619 ( .IN1(n684), .IN2(n472), .Q(n490) );
  AND2X1 U620 ( .IN1(n471), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n489) );
  AND2X1 U621 ( .IN1(n685), .IN2(test_se), .Q(n486) );
  OR2X1 U622 ( .IN1(n492), .IN2(n493), .Q(n175) );
  AND2X1 U623 ( .IN1(n494), .IN2(n423), .Q(n493) );
  OR3X1 U624 ( .IN1(n495), .IN2(n496), .IN3(n497), .Q(n494) );
  AND2X1 U625 ( .IN1(xmit_dataH_3_), .IN2(n479), .Q(n497) );
  AND2X1 U626 ( .IN1(n685), .IN2(n472), .Q(n496) );
  AND2X1 U627 ( .IN1(n684), .IN2(n471), .Q(n495) );
  AND2X1 U628 ( .IN1(n686), .IN2(test_se), .Q(n492) );
  OR2X1 U629 ( .IN1(n498), .IN2(n499), .Q(n174) );
  AND2X1 U630 ( .IN1(n500), .IN2(n423), .Q(n499) );
  OR3X1 U631 ( .IN1(n501), .IN2(n502), .IN3(n503), .Q(n500) );
  AND2X1 U632 ( .IN1(xmit_dataH_2_), .IN2(n479), .Q(n503) );
  AND2X1 U633 ( .IN1(n686), .IN2(n472), .Q(n502) );
  AND2X1 U634 ( .IN1(n685), .IN2(n471), .Q(n501) );
  AND2X1 U635 ( .IN1(n687), .IN2(test_se), .Q(n498) );
  OR2X1 U636 ( .IN1(n504), .IN2(n505), .Q(n173) );
  AND2X1 U637 ( .IN1(n506), .IN2(n423), .Q(n505) );
  OR3X1 U638 ( .IN1(n507), .IN2(n508), .IN3(n509), .Q(n506) );
  AND2X1 U639 ( .IN1(xmit_dataH_1_), .IN2(n479), .Q(n509) );
  AND2X1 U640 ( .IN1(n687), .IN2(n472), .Q(n508) );
  AND2X1 U641 ( .IN1(n686), .IN2(n471), .Q(n507) );
  AND2X1 U642 ( .IN1(test_se), .IN2(n408), .Q(n504) );
  OR2X1 U643 ( .IN1(n510), .IN2(n511), .Q(n172) );
  AND2X1 U644 ( .IN1(n512), .IN2(n423), .Q(n511) );
  OR2X1 U645 ( .IN1(n513), .IN2(n514), .Q(n512) );
  INVX0 U646 ( .INP(n463), .ZN(n514) );
  OR3X1 U647 ( .IN1(xmitH), .IN2(iXMIT_state_2_), .IN3(iXMIT_state_1_), .Q(
        n463) );
  AND2X1 U648 ( .IN1(n431), .IN2(n417), .Q(n513) );
  INVX0 U649 ( .INP(n433), .ZN(n431) );
  OR2X1 U650 ( .IN1(n515), .IN2(n411), .Q(n433) );
  AND2X1 U651 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n510) );
  OR3X1 U652 ( .IN1(n516), .IN2(n517), .IN3(n518), .Q(n171) );
  AND3X1 U653 ( .IN1(n519), .IN2(n423), .IN3(n245), .Q(n517) );
  OR2X1 U654 ( .IN1(n520), .IN2(n412), .Q(n519) );
  AND2X1 U655 ( .IN1(n521), .IN2(iRECEIVER_state_1_), .Q(n520) );
  AND2X1 U656 ( .IN1(n522), .IN2(iRECEIVER_state_0_), .Q(n516) );
  OR3X1 U657 ( .IN1(n523), .IN2(n524), .IN3(test_se), .Q(n522) );
  AND3X1 U658 ( .IN1(n238), .IN2(n412), .IN3(n241), .Q(n524) );
  AND2X1 U659 ( .IN1(n525), .IN2(iRECEIVER_state_1_), .Q(n523) );
  OR2X1 U660 ( .IN1(n526), .IN2(n527), .Q(n170) );
  AND2X1 U661 ( .IN1(n528), .IN2(n423), .Q(n527) );
  OR3X1 U662 ( .IN1(n529), .IN2(n530), .IN3(iRECEIVER_state_2_), .Q(n528) );
  AND2X1 U663 ( .IN1(n531), .IN2(iRECEIVER_state_1_), .Q(n530) );
  OR2X1 U664 ( .IN1(n532), .IN2(n533), .Q(n531) );
  AND2X1 U665 ( .IN1(n534), .IN2(iRECEIVER_state_0_), .Q(n532) );
  OR2X1 U666 ( .IN1(n535), .IN2(n525), .Q(n534) );
  AND4X1 U667 ( .IN1(n691), .IN2(n409), .IN3(n404), .IN4(n406), .Q(n535) );
  AND2X1 U668 ( .IN1(n241), .IN2(n689), .Q(n529) );
  AND2X1 U669 ( .IN1(n691), .IN2(test_se), .Q(n526) );
  OR2X1 U670 ( .IN1(n536), .IN2(n537), .Q(n169) );
  AND2X1 U671 ( .IN1(test_si), .IN2(test_se), .Q(n537) );
  AND2X1 U672 ( .IN1(n538), .IN2(n399), .Q(n536) );
  OR2X1 U673 ( .IN1(n539), .IN2(n540), .Q(n168) );
  AND3X1 U674 ( .IN1(n538), .IN2(n705), .IN3(n399), .Q(n540) );
  AND2X1 U675 ( .IN1(n690), .IN2(n541), .Q(n539) );
  OR2X1 U676 ( .IN1(n542), .IN2(test_se), .Q(n541) );
  AND2X1 U677 ( .IN1(n543), .IN2(n407), .Q(n542) );
  OR2X1 U678 ( .IN1(n544), .IN2(n545), .Q(n167) );
  AND2X1 U679 ( .IN1(n705), .IN2(test_se), .Q(n545) );
  AND3X1 U680 ( .IN1(n546), .IN2(n547), .IN3(n538), .Q(n544) );
  OR2X1 U681 ( .IN1(n548), .IN2(n703), .Q(n546) );
  AND2X1 U682 ( .IN1(n690), .IN2(n705), .Q(n548) );
  OR2X1 U683 ( .IN1(n549), .IN2(n550), .Q(n166) );
  AND2X1 U684 ( .IN1(n703), .IN2(test_se), .Q(n550) );
  AND2X1 U685 ( .IN1(n538), .IN2(n551), .Q(n549) );
  OR2X1 U686 ( .IN1(n552), .IN2(n553), .Q(n551) );
  AND2X1 U687 ( .IN1(n554), .IN2(n414), .Q(n553) );
  AND2X1 U688 ( .IN1(n704), .IN2(n547), .Q(n552) );
  INVX0 U689 ( .INP(n554), .ZN(n547) );
  AND3X1 U690 ( .IN1(n703), .IN2(n705), .IN3(n690), .Q(n554) );
  AND2X1 U691 ( .IN1(n423), .IN2(n543), .Q(n538) );
  AND4X1 U692 ( .IN1(n555), .IN2(n238), .IN3(iRECEIVER_state_1_), .IN4(n556), 
        .Q(n543) );
  OR2X1 U693 ( .IN1(n521), .IN2(iRECEIVER_state_0_), .Q(n556) );
  INVX0 U694 ( .INP(n533), .ZN(n521) );
  AND4X1 U695 ( .IN1(n407), .IN2(n703), .IN3(n399), .IN4(n414), .Q(n533) );
  OR2X1 U696 ( .IN1(n557), .IN2(iRECEIVER_next_state_2_), .Q(n164) );
  AND2X1 U697 ( .IN1(test_se), .IN2(iRECEIVER_state_1_), .Q(n557) );
  OR2X1 U698 ( .IN1(n558), .IN2(n559), .Q(n163) );
  AND2X1 U699 ( .IN1(n688), .IN2(test_se), .Q(n559) );
  AND2X1 U700 ( .IN1(n560), .IN2(n423), .Q(n558) );
  OR2X1 U701 ( .IN1(n561), .IN2(n562), .Q(n560) );
  AND2X1 U702 ( .IN1(iRECEIVER_state_2_), .IN2(iRECEIVER_state_0_), .Q(n561)
         );
  OR3X1 U703 ( .IN1(n563), .IN2(n564), .IN3(n565), .Q(n162) );
  AND2X1 U704 ( .IN1(rec_dataH_rec_6), .IN2(test_se), .Q(n565) );
  AND2X1 U705 ( .IN1(n518), .IN2(n689), .Q(n564) );
  AND2X1 U706 ( .IN1(rec_dataH_rec_7), .IN2(n566), .Q(n563) );
  OR2X1 U707 ( .IN1(n567), .IN2(n568), .Q(n161) );
  AND2X1 U708 ( .IN1(rec_dataH_temp_6), .IN2(test_se), .Q(n568) );
  AND2X1 U709 ( .IN1(rec_dataH_rec_7), .IN2(n423), .Q(n567) );
  OR2X1 U710 ( .IN1(n569), .IN2(n570), .Q(n160) );
  AND2X1 U711 ( .IN1(rec_dataH_6_), .IN2(test_se), .Q(n570) );
  AND2X1 U712 ( .IN1(test_so), .IN2(n423), .Q(n569) );
  OR3X1 U713 ( .IN1(n571), .IN2(n572), .IN3(n573), .Q(n159) );
  AND2X1 U714 ( .IN1(rec_dataH_rec_5), .IN2(test_se), .Q(n573) );
  AND2X1 U715 ( .IN1(n518), .IN2(rec_dataH_rec_7), .Q(n572) );
  AND2X1 U716 ( .IN1(rec_dataH_rec_6), .IN2(n566), .Q(n571) );
  OR2X1 U717 ( .IN1(n574), .IN2(n575), .Q(n157) );
  AND2X1 U718 ( .IN1(rec_dataH_temp_5), .IN2(test_se), .Q(n575) );
  AND2X1 U719 ( .IN1(rec_dataH_rec_6), .IN2(n423), .Q(n574) );
  OR2X1 U720 ( .IN1(n576), .IN2(n577), .Q(n156) );
  AND2X1 U721 ( .IN1(rec_dataH_5_), .IN2(test_se), .Q(n577) );
  AND2X1 U722 ( .IN1(rec_dataH_temp_6), .IN2(n423), .Q(n576) );
  OR3X1 U723 ( .IN1(n578), .IN2(n579), .IN3(n580), .Q(n155) );
  AND2X1 U724 ( .IN1(rec_dataH_rec_4), .IN2(test_se), .Q(n580) );
  AND2X1 U725 ( .IN1(rec_dataH_rec_6), .IN2(n518), .Q(n579) );
  AND2X1 U726 ( .IN1(rec_dataH_rec_5), .IN2(n566), .Q(n578) );
  OR2X1 U727 ( .IN1(n581), .IN2(n582), .Q(n154) );
  AND2X1 U728 ( .IN1(rec_dataH_temp_4), .IN2(test_se), .Q(n582) );
  AND2X1 U729 ( .IN1(rec_dataH_rec_5), .IN2(n423), .Q(n581) );
  OR2X1 U730 ( .IN1(n583), .IN2(n584), .Q(n153) );
  AND2X1 U731 ( .IN1(rec_dataH_4_), .IN2(test_se), .Q(n584) );
  AND2X1 U732 ( .IN1(rec_dataH_temp_5), .IN2(n423), .Q(n583) );
  OR3X1 U733 ( .IN1(n585), .IN2(n586), .IN3(n587), .Q(n152) );
  AND2X1 U734 ( .IN1(rec_dataH_rec_3), .IN2(test_se), .Q(n587) );
  AND2X1 U735 ( .IN1(rec_dataH_rec_5), .IN2(n518), .Q(n586) );
  AND2X1 U736 ( .IN1(rec_dataH_rec_4), .IN2(n566), .Q(n585) );
  OR2X1 U737 ( .IN1(n588), .IN2(n589), .Q(n150) );
  AND2X1 U738 ( .IN1(rec_dataH_temp_3), .IN2(test_se), .Q(n589) );
  AND2X1 U739 ( .IN1(rec_dataH_rec_4), .IN2(n423), .Q(n588) );
  OR2X1 U740 ( .IN1(n590), .IN2(n591), .Q(n149) );
  AND2X1 U741 ( .IN1(rec_dataH_3_), .IN2(test_se), .Q(n591) );
  AND2X1 U742 ( .IN1(rec_dataH_temp_4), .IN2(n423), .Q(n590) );
  OR3X1 U743 ( .IN1(n592), .IN2(n593), .IN3(n594), .Q(n148) );
  AND2X1 U744 ( .IN1(rec_dataH_rec_2), .IN2(test_se), .Q(n594) );
  AND2X1 U745 ( .IN1(rec_dataH_rec_4), .IN2(n518), .Q(n593) );
  AND2X1 U746 ( .IN1(rec_dataH_rec_3), .IN2(n566), .Q(n592) );
  OR2X1 U747 ( .IN1(n595), .IN2(n596), .Q(n147) );
  AND2X1 U748 ( .IN1(rec_dataH_temp_2), .IN2(test_se), .Q(n596) );
  AND2X1 U749 ( .IN1(rec_dataH_rec_3), .IN2(n423), .Q(n595) );
  OR2X1 U750 ( .IN1(n597), .IN2(n598), .Q(n146) );
  AND2X1 U751 ( .IN1(rec_dataH_2_), .IN2(test_se), .Q(n598) );
  AND2X1 U752 ( .IN1(rec_dataH_temp_3), .IN2(n423), .Q(n597) );
  OR3X1 U753 ( .IN1(n599), .IN2(n600), .IN3(n601), .Q(n145) );
  AND2X1 U754 ( .IN1(rec_dataH_rec_1), .IN2(test_se), .Q(n601) );
  AND2X1 U755 ( .IN1(rec_dataH_rec_3), .IN2(n518), .Q(n600) );
  AND2X1 U756 ( .IN1(rec_dataH_rec_2), .IN2(n566), .Q(n599) );
  OR2X1 U757 ( .IN1(n602), .IN2(n603), .Q(n143) );
  AND2X1 U758 ( .IN1(rec_dataH_temp_1), .IN2(test_se), .Q(n603) );
  AND2X1 U759 ( .IN1(rec_dataH_rec_2), .IN2(n423), .Q(n602) );
  OR2X1 U760 ( .IN1(n604), .IN2(n605), .Q(n142) );
  AND2X1 U761 ( .IN1(rec_dataH_1_), .IN2(test_se), .Q(n605) );
  AND2X1 U762 ( .IN1(rec_dataH_temp_2), .IN2(n423), .Q(n604) );
  OR3X1 U763 ( .IN1(n606), .IN2(n607), .IN3(n608), .Q(n141) );
  AND2X1 U764 ( .IN1(rec_dataH_rec_0), .IN2(test_se), .Q(n608) );
  AND2X1 U765 ( .IN1(rec_dataH_rec_2), .IN2(n518), .Q(n607) );
  AND2X1 U766 ( .IN1(rec_dataH_rec_1), .IN2(n566), .Q(n606) );
  OR2X1 U767 ( .IN1(n609), .IN2(n610), .Q(n140) );
  AND2X1 U768 ( .IN1(rec_dataH_temp_0), .IN2(test_se), .Q(n610) );
  AND2X1 U769 ( .IN1(rec_dataH_rec_1), .IN2(n423), .Q(n609) );
  OR2X1 U770 ( .IN1(n611), .IN2(n612), .Q(n139) );
  AND2X1 U771 ( .IN1(rec_dataH_0_), .IN2(test_se), .Q(n612) );
  AND2X1 U772 ( .IN1(rec_dataH_temp_1), .IN2(n423), .Q(n611) );
  OR3X1 U773 ( .IN1(n613), .IN2(n614), .IN3(n615), .Q(n138) );
  AND2X1 U774 ( .IN1(n704), .IN2(test_se), .Q(n615) );
  AND2X1 U775 ( .IN1(rec_dataH_rec_1), .IN2(n518), .Q(n614) );
  AND2X1 U776 ( .IN1(rec_dataH_rec_0), .IN2(n566), .Q(n613) );
  INVX0 U777 ( .INP(n616), .ZN(n566) );
  OR2X1 U778 ( .IN1(test_se), .IN2(n617), .Q(n616) );
  OR2X1 U779 ( .IN1(n618), .IN2(n619), .Q(n136) );
  AND2X1 U780 ( .IN1(rec_dataH_7_), .IN2(test_se), .Q(n619) );
  AND2X1 U781 ( .IN1(rec_dataH_rec_0), .IN2(n423), .Q(n618) );
  OR2X1 U782 ( .IN1(n620), .IN2(n621), .Q(n135) );
  AND2X1 U783 ( .IN1(xmit_doneH_temp), .IN2(test_se), .Q(n621) );
  AND2X1 U784 ( .IN1(rec_dataH_temp_0), .IN2(n423), .Q(n620) );
  OR2X1 U785 ( .IN1(n622), .IN2(n623), .Q(n134) );
  AND2X1 U786 ( .IN1(n691), .IN2(n624), .Q(n623) );
  OR3X1 U787 ( .IN1(n625), .IN2(n626), .IN3(n627), .Q(n624) );
  AND2X1 U788 ( .IN1(n518), .IN2(n409), .Q(n626) );
  AND2X1 U789 ( .IN1(n694), .IN2(n628), .Q(n622) );
  OR2X1 U790 ( .IN1(n629), .IN2(test_se), .Q(n628) );
  AND4X1 U791 ( .IN1(n692), .IN2(n693), .IN3(n518), .IN4(n416), .Q(n629) );
  OR3X1 U792 ( .IN1(n625), .IN2(n630), .IN3(n631), .Q(n133) );
  AND2X1 U793 ( .IN1(rec_readyH), .IN2(test_se), .Q(n631) );
  AND2X1 U794 ( .IN1(n632), .IN2(n693), .Q(n630) );
  OR2X1 U795 ( .IN1(n633), .IN2(n634), .Q(n132) );
  AND2X1 U796 ( .IN1(n692), .IN2(n635), .Q(n634) );
  OR2X1 U797 ( .IN1(n625), .IN2(n632), .Q(n635) );
  AND2X1 U798 ( .IN1(n404), .IN2(n518), .Q(n625) );
  AND2X1 U799 ( .IN1(n693), .IN2(n636), .Q(n633) );
  OR2X1 U800 ( .IN1(n637), .IN2(test_se), .Q(n636) );
  AND2X1 U801 ( .IN1(n617), .IN2(n406), .Q(n637) );
  OR2X1 U802 ( .IN1(n638), .IN2(n639), .Q(n131) );
  AND2X1 U803 ( .IN1(n694), .IN2(n627), .Q(n639) );
  OR2X1 U804 ( .IN1(n640), .IN2(n632), .Q(n627) );
  INVX0 U805 ( .INP(n641), .ZN(n632) );
  OR3X1 U806 ( .IN1(n617), .IN2(n562), .IN3(test_se), .Q(n641) );
  AND3X1 U807 ( .IN1(n241), .IN2(n689), .IN3(n238), .Q(n562) );
  AND2X1 U808 ( .IN1(n518), .IN2(n406), .Q(n640) );
  AND2X1 U809 ( .IN1(n423), .IN2(n617), .Q(n518) );
  AND2X1 U810 ( .IN1(n692), .IN2(n642), .Q(n638) );
  OR2X1 U811 ( .IN1(n643), .IN2(test_se), .Q(n642) );
  AND2X1 U812 ( .IN1(n617), .IN2(n644), .Q(n643) );
  OR2X1 U813 ( .IN1(n645), .IN2(n646), .Q(n644) );
  AND2X1 U814 ( .IN1(n694), .IN2(n404), .Q(n646) );
  AND2X1 U815 ( .IN1(n693), .IN2(n409), .Q(n645) );
  AND2X1 U816 ( .IN1(n245), .IN2(iRECEIVER_state_2_), .Q(n617) );
  OR2X1 U817 ( .IN1(n647), .IN2(n648), .Q(n129) );
  AND2X1 U818 ( .IN1(test_se), .IN2(n700), .Q(n648) );
  AND2X1 U819 ( .IN1(iXMIT_N29), .IN2(n423), .Q(n647) );
  OR2X1 U820 ( .IN1(n649), .IN2(n650), .Q(n128) );
  AND2X1 U821 ( .IN1(iXMIT_N26), .IN2(n423), .Q(n650) );
  AND2X1 U822 ( .IN1(test_se), .IN2(iRECEIVER_state_2_), .Q(n649) );
  OR2X1 U823 ( .IN1(n651), .IN2(n652), .Q(n127) );
  AND2X1 U824 ( .IN1(test_se), .IN2(n702), .Q(n652) );
  AND2X1 U825 ( .IN1(iXMIT_N27), .IN2(n423), .Q(n651) );
  OR2X1 U826 ( .IN1(n653), .IN2(n654), .Q(n126) );
  AND2X1 U827 ( .IN1(n655), .IN2(n423), .Q(n654) );
  OR3X1 U828 ( .IN1(n656), .IN2(n657), .IN3(n658), .Q(n655) );
  AND2X1 U829 ( .IN1(xmit_dataH_0_), .IN2(n479), .Q(n658) );
  AND2X1 U830 ( .IN1(n472), .IN2(n408), .Q(n657) );
  AND2X1 U831 ( .IN1(n687), .IN2(n471), .Q(n656) );
  INVX0 U832 ( .INP(n659), .ZN(n471) );
  OR2X1 U833 ( .IN1(n479), .IN2(n472), .Q(n659) );
  INVX0 U834 ( .INP(n444), .ZN(n472) );
  OR2X1 U835 ( .IN1(n660), .IN2(n479), .Q(n444) );
  AND2X1 U836 ( .IN1(n239), .IN2(iXMIT_state_2_), .Q(n660) );
  AND3X1 U837 ( .IN1(n242), .IN2(n246), .IN3(xmitH), .Q(n479) );
  AND2X1 U838 ( .IN1(test_se), .IN2(iXMIT_state_2_), .Q(n653) );
  OR2X1 U839 ( .IN1(n661), .IN2(n662), .Q(n125) );
  AND2X1 U840 ( .IN1(n689), .IN2(test_se), .Q(n662) );
  AND2X1 U841 ( .IN1(uart_REC_dataH), .IN2(n423), .Q(n661) );
  OR2X1 U842 ( .IN1(n663), .IN2(n664), .Q(n124) );
  AND2X1 U843 ( .IN1(rec_dataH_rec_7), .IN2(test_se), .Q(n664) );
  AND2X1 U844 ( .IN1(n688), .IN2(n423), .Q(n663) );
  INVX0 U845 ( .INP(test_se), .ZN(n423) );
  OR2X1 U846 ( .IN1(n665), .IN2(n666), .Q(iXMIT_N46) );
  INVX0 U847 ( .INP(n667), .ZN(n666) );
  OR2X1 U848 ( .IN1(n668), .IN2(n695), .Q(n667) );
  AND2X1 U849 ( .IN1(n695), .IN2(n668), .Q(n665) );
  AND2X1 U850 ( .IN1(n668), .IN2(n669), .Q(iXMIT_N45) );
  OR2X1 U851 ( .IN1(n696), .IN2(n670), .Q(n669) );
  AND2X1 U852 ( .IN1(n697), .IN2(n698), .Q(n670) );
  OR3X1 U853 ( .IN1(n398), .IN2(n405), .IN3(n410), .Q(n668) );
  OR2X1 U854 ( .IN1(n671), .IN2(n672), .Q(iXMIT_N44) );
  AND2X1 U855 ( .IN1(n698), .IN2(n398), .Q(n672) );
  AND2X1 U856 ( .IN1(n697), .IN2(n405), .Q(n671) );
  AND2X1 U857 ( .IN1(n673), .IN2(iXMIT_N25), .Q(iXMIT_N29) );
  AND2X1 U858 ( .IN1(n673), .IN2(iXMIT_N24), .Q(iXMIT_N28) );
  OR2X1 U859 ( .IN1(n674), .IN2(n675), .Q(iXMIT_N27) );
  AND2X1 U860 ( .IN1(iXMIT_N26), .IN2(n701), .Q(n675) );
  AND3X1 U861 ( .IN1(n702), .IN2(n673), .IN3(n415), .Q(n674) );
  AND2X1 U862 ( .IN1(n413), .IN2(n673), .Q(iXMIT_N26) );
  OR2X1 U863 ( .IN1(n417), .IN2(n443), .Q(n673) );
  AND2X1 U864 ( .IN1(n439), .IN2(iXMIT_state_1_), .Q(n443) );
  OR2X1 U865 ( .IN1(n239), .IN2(n465), .Q(n439) );
  INVX0 U866 ( .INP(n676), .ZN(n465) );
  AND4X1 U867 ( .IN1(n700), .IN2(n699), .IN3(n413), .IN4(n701), .Q(n676) );
  AND2X1 U868 ( .IN1(iXMIT_state_2_), .IN2(iXMIT_state_0_), .Q(n417) );
  OR2X1 U869 ( .IN1(n677), .IN2(n678), .Q(iXMIT_N25) );
  AND2X1 U870 ( .IN1(n679), .IN2(n411), .Q(n678) );
  AND2X1 U871 ( .IN1(n699), .IN2(n515), .Q(n677) );
  AND2X1 U872 ( .IN1(n515), .IN2(n680), .Q(iXMIT_N24) );
  OR2X1 U873 ( .IN1(n700), .IN2(n681), .Q(n680) );
  AND2X1 U874 ( .IN1(n702), .IN2(n701), .Q(n681) );
  INVX0 U875 ( .INP(n679), .ZN(n515) );
  AND3X1 U876 ( .IN1(n702), .IN2(n701), .IN3(n700), .Q(n679) );
  AND2X1 U877 ( .IN1(iRECEIVER_state_1_), .IN2(n682), .Q(
        iRECEIVER_next_state_2_) );
  INVX0 U878 ( .INP(n555), .ZN(n682) );
  OR2X1 U879 ( .IN1(n245), .IN2(n525), .Q(n555) );
  INVX0 U880 ( .INP(n683), .ZN(n525) );
  AND4X1 U881 ( .IN1(n705), .IN2(n704), .IN3(n399), .IN4(n703), .Q(n683) );
endmodule

