module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n1132_, new_n500_, new_n898_, new_n1163_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n1162_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1151_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n1145_, new_n657_, new_n1150_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1159_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n1147_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n1154_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n1032_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n775_, new_n371_, new_n886_, new_n509_, new_n1096_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n1160_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n918_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n468_, new_n1122_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n597_, new_n978_, new_n1092_, new_n408_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n651_, new_n433_, new_n1164_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n226_, new_n802_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n202_, keyIn_0_72 );
not g001 ( new_n203_, keyIn_0_64 );
not g002 ( new_n204_, keyIn_0_45 );
not g003 ( new_n205_, N93 );
nand g004 ( new_n206_, new_n205_, N89 );
not g005 ( new_n207_, N89 );
nand g006 ( new_n208_, new_n207_, N93 );
nand g007 ( new_n209_, new_n206_, new_n208_ );
nand g008 ( new_n210_, new_n209_, keyIn_0_11 );
not g009 ( new_n211_, keyIn_0_11 );
nand g010 ( new_n212_, new_n206_, new_n208_, new_n211_ );
nand g011 ( new_n213_, new_n210_, new_n212_ );
not g012 ( new_n214_, N81 );
not g013 ( new_n215_, N85 );
nand g014 ( new_n216_, new_n214_, new_n215_ );
nand g015 ( new_n217_, N81, N85 );
nand g016 ( new_n218_, new_n216_, new_n217_ );
nand g017 ( new_n219_, new_n218_, keyIn_0_10 );
not g018 ( new_n220_, keyIn_0_10 );
nand g019 ( new_n221_, new_n216_, new_n220_, new_n217_ );
nand g020 ( new_n222_, new_n219_, new_n221_ );
nand g021 ( new_n223_, new_n213_, new_n222_ );
nand g022 ( new_n224_, new_n210_, new_n219_, new_n212_, new_n221_ );
nand g023 ( new_n225_, new_n223_, new_n224_ );
nand g024 ( new_n226_, new_n225_, new_n204_ );
nand g025 ( new_n227_, new_n223_, keyIn_0_45, new_n224_ );
nand g026 ( new_n228_, new_n226_, new_n227_ );
not g027 ( new_n229_, keyIn_0_44 );
not g028 ( new_n230_, keyIn_0_9 );
not g029 ( new_n231_, N77 );
nand g030 ( new_n232_, new_n231_, N73 );
not g031 ( new_n233_, N73 );
nand g032 ( new_n234_, new_n233_, N77 );
nand g033 ( new_n235_, new_n232_, new_n234_ );
nand g034 ( new_n236_, new_n235_, new_n230_ );
nand g035 ( new_n237_, new_n232_, new_n234_, keyIn_0_9 );
nand g036 ( new_n238_, new_n236_, new_n237_ );
not g037 ( new_n239_, N69 );
nand g038 ( new_n240_, new_n239_, N65 );
not g039 ( new_n241_, N65 );
nand g040 ( new_n242_, new_n241_, N69 );
nand g041 ( new_n243_, new_n240_, new_n242_, keyIn_0_8 );
not g042 ( new_n244_, keyIn_0_8 );
nand g043 ( new_n245_, new_n240_, new_n242_ );
nand g044 ( new_n246_, new_n245_, new_n244_ );
nand g045 ( new_n247_, new_n238_, new_n243_, new_n246_ );
nand g046 ( new_n248_, new_n246_, new_n243_ );
nand g047 ( new_n249_, new_n248_, new_n236_, new_n237_ );
nand g048 ( new_n250_, new_n247_, new_n249_ );
nand g049 ( new_n251_, new_n250_, new_n229_ );
nand g050 ( new_n252_, new_n247_, new_n249_, keyIn_0_44 );
nand g051 ( new_n253_, new_n251_, new_n252_ );
nand g052 ( new_n254_, new_n253_, new_n228_ );
nand g053 ( new_n255_, new_n251_, new_n226_, new_n227_, new_n252_ );
nand g054 ( new_n256_, new_n254_, new_n255_ );
nand g055 ( new_n257_, new_n256_, keyIn_0_60 );
not g056 ( new_n258_, keyIn_0_60 );
nand g057 ( new_n259_, new_n254_, new_n258_, new_n255_ );
nand g058 ( new_n260_, new_n257_, new_n259_ );
nand g059 ( new_n261_, N129, N137 );
nand g060 ( new_n262_, new_n261_, keyIn_0_16 );
not g061 ( new_n263_, keyIn_0_16 );
nand g062 ( new_n264_, new_n263_, N129, N137 );
nand g063 ( new_n265_, new_n262_, new_n264_ );
nand g064 ( new_n266_, new_n260_, new_n265_ );
nand g065 ( new_n267_, new_n257_, new_n259_, new_n262_, new_n264_ );
nand g066 ( new_n268_, new_n266_, new_n267_ );
nand g067 ( new_n269_, new_n268_, new_n203_ );
nand g068 ( new_n270_, new_n266_, keyIn_0_64, new_n267_ );
nand g069 ( new_n271_, new_n269_, new_n270_ );
not g070 ( new_n272_, keyIn_0_48 );
nor g071 ( new_n273_, N33, N49 );
not g072 ( new_n274_, new_n273_ );
nand g073 ( new_n275_, N33, N49 );
nand g074 ( new_n276_, new_n274_, new_n275_ );
nand g075 ( new_n277_, new_n276_, keyIn_0_25 );
not g076 ( new_n278_, new_n277_ );
nor g077 ( new_n279_, new_n276_, keyIn_0_25 );
nor g078 ( new_n280_, new_n278_, new_n279_ );
not g079 ( new_n281_, new_n280_ );
not g080 ( new_n282_, N17 );
nand g081 ( new_n283_, new_n282_, N1 );
not g082 ( new_n284_, N1 );
nand g083 ( new_n285_, new_n284_, N17 );
nand g084 ( new_n286_, new_n283_, new_n285_ );
nand g085 ( new_n287_, new_n286_, keyIn_0_24 );
not g086 ( new_n288_, keyIn_0_24 );
nand g087 ( new_n289_, new_n283_, new_n285_, new_n288_ );
nand g088 ( new_n290_, new_n287_, new_n289_ );
nand g089 ( new_n291_, new_n281_, new_n290_ );
nand g090 ( new_n292_, new_n280_, new_n287_, new_n289_ );
nand g091 ( new_n293_, new_n291_, new_n292_ );
nand g092 ( new_n294_, new_n293_, new_n272_ );
nand g093 ( new_n295_, new_n291_, keyIn_0_48, new_n292_ );
nand g094 ( new_n296_, new_n294_, new_n295_ );
nand g095 ( new_n297_, new_n271_, new_n296_ );
nand g096 ( new_n298_, new_n269_, new_n270_, new_n294_, new_n295_ );
nand g097 ( new_n299_, new_n297_, new_n298_ );
nand g098 ( new_n300_, new_n299_, new_n202_ );
nand g099 ( new_n301_, new_n297_, keyIn_0_72, new_n298_ );
nand g100 ( new_n302_, new_n300_, new_n301_ );
not g101 ( new_n303_, new_n302_ );
not g102 ( new_n304_, keyIn_0_112 );
not g103 ( new_n305_, keyIn_0_89 );
not g104 ( new_n306_, keyIn_0_65 );
not g105 ( new_n307_, keyIn_0_61 );
not g106 ( new_n308_, keyIn_0_47 );
not g107 ( new_n309_, N117 );
nand g108 ( new_n310_, new_n309_, N113 );
not g109 ( new_n311_, N113 );
nand g110 ( new_n312_, new_n311_, N117 );
nand g111 ( new_n313_, new_n310_, new_n312_ );
nand g112 ( new_n314_, new_n313_, keyIn_0_14 );
not g113 ( new_n315_, keyIn_0_14 );
nand g114 ( new_n316_, new_n310_, new_n312_, new_n315_ );
nand g115 ( new_n317_, new_n314_, new_n316_ );
not g116 ( new_n318_, N125 );
nand g117 ( new_n319_, new_n318_, N121 );
not g118 ( new_n320_, N121 );
nand g119 ( new_n321_, new_n320_, N125 );
nand g120 ( new_n322_, new_n319_, new_n321_ );
nand g121 ( new_n323_, new_n322_, keyIn_0_15 );
not g122 ( new_n324_, keyIn_0_15 );
nand g123 ( new_n325_, new_n319_, new_n321_, new_n324_ );
nand g124 ( new_n326_, new_n323_, new_n325_ );
nand g125 ( new_n327_, new_n317_, new_n326_ );
nand g126 ( new_n328_, new_n314_, new_n323_, new_n316_, new_n325_ );
nand g127 ( new_n329_, new_n327_, new_n328_ );
nand g128 ( new_n330_, new_n329_, new_n308_ );
nand g129 ( new_n331_, new_n327_, keyIn_0_47, new_n328_ );
nand g130 ( new_n332_, new_n330_, new_n331_ );
not g131 ( new_n333_, new_n332_ );
not g132 ( new_n334_, keyIn_0_46 );
not g133 ( new_n335_, N101 );
nand g134 ( new_n336_, new_n335_, N97 );
not g135 ( new_n337_, N97 );
nand g136 ( new_n338_, new_n337_, N101 );
nand g137 ( new_n339_, new_n336_, new_n338_ );
nand g138 ( new_n340_, new_n339_, keyIn_0_12 );
not g139 ( new_n341_, keyIn_0_12 );
nand g140 ( new_n342_, new_n336_, new_n338_, new_n341_ );
nand g141 ( new_n343_, new_n340_, new_n342_ );
nand g142 ( new_n344_, new_n343_, keyIn_0_13 );
not g143 ( new_n345_, keyIn_0_13 );
nand g144 ( new_n346_, new_n340_, new_n345_, new_n342_ );
nand g145 ( new_n347_, new_n344_, new_n346_ );
not g146 ( new_n348_, N105 );
nor g147 ( new_n349_, new_n348_, N109 );
not g148 ( new_n350_, N109 );
nor g149 ( new_n351_, new_n350_, N105 );
nor g150 ( new_n352_, new_n349_, new_n351_ );
nand g151 ( new_n353_, new_n347_, new_n352_ );
not g152 ( new_n354_, new_n352_ );
nand g153 ( new_n355_, new_n344_, new_n346_, new_n354_ );
nand g154 ( new_n356_, new_n353_, new_n355_ );
nand g155 ( new_n357_, new_n356_, new_n334_ );
nand g156 ( new_n358_, new_n353_, keyIn_0_46, new_n355_ );
nand g157 ( new_n359_, new_n357_, new_n358_ );
nand g158 ( new_n360_, new_n359_, new_n333_ );
nand g159 ( new_n361_, new_n357_, new_n332_, new_n358_ );
nand g160 ( new_n362_, new_n360_, new_n361_ );
nand g161 ( new_n363_, new_n362_, new_n307_ );
nand g162 ( new_n364_, new_n360_, keyIn_0_61, new_n361_ );
nand g163 ( new_n365_, new_n363_, new_n364_ );
not g164 ( new_n366_, keyIn_0_17 );
nand g165 ( new_n367_, N130, N137 );
nand g166 ( new_n368_, new_n367_, new_n366_ );
nand g167 ( new_n369_, keyIn_0_17, N130, N137 );
nand g168 ( new_n370_, new_n368_, new_n369_ );
not g169 ( new_n371_, new_n370_ );
nand g170 ( new_n372_, new_n365_, new_n371_ );
nand g171 ( new_n373_, new_n363_, new_n364_, new_n370_ );
nand g172 ( new_n374_, new_n372_, new_n373_ );
nand g173 ( new_n375_, new_n374_, new_n306_ );
nand g174 ( new_n376_, new_n372_, keyIn_0_65, new_n373_ );
nand g175 ( new_n377_, new_n375_, new_n376_ );
nor g176 ( new_n378_, N5, N21 );
not g177 ( new_n379_, new_n378_ );
nand g178 ( new_n380_, N5, N21 );
nand g179 ( new_n381_, new_n379_, new_n380_ );
nand g180 ( new_n382_, new_n381_, keyIn_0_26 );
not g181 ( new_n383_, new_n382_ );
nor g182 ( new_n384_, new_n381_, keyIn_0_26 );
nor g183 ( new_n385_, new_n383_, new_n384_ );
not g184 ( new_n386_, new_n385_ );
not g185 ( new_n387_, N53 );
nand g186 ( new_n388_, new_n387_, N37 );
not g187 ( new_n389_, N37 );
nand g188 ( new_n390_, new_n389_, N53 );
nand g189 ( new_n391_, new_n388_, new_n390_ );
nand g190 ( new_n392_, new_n391_, keyIn_0_27 );
not g191 ( new_n393_, keyIn_0_27 );
nand g192 ( new_n394_, new_n388_, new_n390_, new_n393_ );
nand g193 ( new_n395_, new_n392_, new_n394_ );
nand g194 ( new_n396_, new_n386_, new_n395_ );
nand g195 ( new_n397_, new_n385_, new_n392_, new_n394_ );
nand g196 ( new_n398_, new_n396_, new_n397_ );
nand g197 ( new_n399_, new_n398_, keyIn_0_49 );
not g198 ( new_n400_, keyIn_0_49 );
nand g199 ( new_n401_, new_n396_, new_n400_, new_n397_ );
nand g200 ( new_n402_, new_n399_, new_n401_ );
nand g201 ( new_n403_, new_n377_, new_n402_ );
nand g202 ( new_n404_, new_n375_, new_n376_, new_n399_, new_n401_ );
nand g203 ( new_n405_, new_n403_, new_n404_ );
nand g204 ( new_n406_, new_n405_, keyIn_0_73 );
not g205 ( new_n407_, keyIn_0_73 );
nand g206 ( new_n408_, new_n403_, new_n407_, new_n404_ );
nand g207 ( new_n409_, new_n406_, new_n408_ );
nand g208 ( new_n410_, new_n409_, new_n305_ );
not g209 ( new_n411_, keyIn_0_67 );
not g210 ( new_n412_, keyIn_0_63 );
nand g211 ( new_n413_, new_n332_, new_n228_ );
nand g212 ( new_n414_, new_n330_, new_n226_, new_n331_, new_n227_ );
nand g213 ( new_n415_, new_n413_, new_n414_ );
nand g214 ( new_n416_, new_n415_, new_n412_ );
nand g215 ( new_n417_, new_n413_, keyIn_0_63, new_n414_ );
nand g216 ( new_n418_, new_n416_, new_n417_ );
not g217 ( new_n419_, keyIn_0_19 );
nand g218 ( new_n420_, N132, N137 );
nand g219 ( new_n421_, new_n420_, new_n419_ );
nand g220 ( new_n422_, keyIn_0_19, N132, N137 );
nand g221 ( new_n423_, new_n421_, new_n422_ );
nand g222 ( new_n424_, new_n418_, new_n423_ );
nand g223 ( new_n425_, new_n416_, new_n417_, new_n421_, new_n422_ );
nand g224 ( new_n426_, new_n424_, new_n425_ );
nand g225 ( new_n427_, new_n426_, new_n411_ );
nand g226 ( new_n428_, new_n424_, keyIn_0_67, new_n425_ );
nand g227 ( new_n429_, new_n427_, new_n428_ );
nor g228 ( new_n430_, N45, N61 );
not g229 ( new_n431_, new_n430_ );
nand g230 ( new_n432_, N45, N61 );
nand g231 ( new_n433_, new_n431_, new_n432_ );
nand g232 ( new_n434_, new_n433_, keyIn_0_31 );
not g233 ( new_n435_, new_n434_ );
nor g234 ( new_n436_, new_n433_, keyIn_0_31 );
nor g235 ( new_n437_, new_n435_, new_n436_ );
not g236 ( new_n438_, new_n437_ );
not g237 ( new_n439_, N29 );
nand g238 ( new_n440_, new_n439_, N13 );
not g239 ( new_n441_, N13 );
nand g240 ( new_n442_, new_n441_, N29 );
nand g241 ( new_n443_, new_n440_, new_n442_ );
nand g242 ( new_n444_, new_n443_, keyIn_0_30 );
not g243 ( new_n445_, keyIn_0_30 );
nand g244 ( new_n446_, new_n440_, new_n442_, new_n445_ );
nand g245 ( new_n447_, new_n444_, new_n446_ );
nand g246 ( new_n448_, new_n438_, new_n447_ );
nand g247 ( new_n449_, new_n437_, new_n444_, new_n446_ );
nand g248 ( new_n450_, new_n448_, new_n449_ );
nand g249 ( new_n451_, new_n450_, keyIn_0_51 );
not g250 ( new_n452_, keyIn_0_51 );
nand g251 ( new_n453_, new_n448_, new_n452_, new_n449_ );
nand g252 ( new_n454_, new_n451_, new_n453_ );
nand g253 ( new_n455_, new_n429_, new_n454_ );
nand g254 ( new_n456_, new_n427_, new_n428_, new_n451_, new_n453_ );
nand g255 ( new_n457_, new_n455_, new_n456_ );
nand g256 ( new_n458_, new_n457_, keyIn_0_75 );
not g257 ( new_n459_, keyIn_0_75 );
nand g258 ( new_n460_, new_n455_, new_n459_, new_n456_ );
nand g259 ( new_n461_, new_n458_, keyIn_0_91, new_n460_ );
not g260 ( new_n462_, keyIn_0_91 );
nand g261 ( new_n463_, new_n458_, new_n460_ );
nand g262 ( new_n464_, new_n463_, new_n462_ );
nand g263 ( new_n465_, new_n464_, new_n303_, new_n461_ );
not g264 ( new_n466_, new_n465_ );
nand g265 ( new_n467_, new_n466_, new_n410_ );
nand g266 ( new_n468_, new_n406_, keyIn_0_89, new_n408_ );
not g267 ( new_n469_, keyIn_0_74 );
not g268 ( new_n470_, keyIn_0_66 );
not g269 ( new_n471_, keyIn_0_62 );
not g270 ( new_n472_, new_n253_ );
nand g271 ( new_n473_, new_n359_, new_n472_ );
nand g272 ( new_n474_, new_n357_, new_n358_, new_n253_ );
nand g273 ( new_n475_, new_n473_, new_n474_ );
nand g274 ( new_n476_, new_n475_, new_n471_ );
nand g275 ( new_n477_, new_n473_, keyIn_0_62, new_n474_ );
nand g276 ( new_n478_, new_n476_, new_n477_ );
not g277 ( new_n479_, keyIn_0_18 );
nand g278 ( new_n480_, N131, N137 );
nand g279 ( new_n481_, new_n480_, new_n479_ );
nand g280 ( new_n482_, keyIn_0_18, N131, N137 );
nand g281 ( new_n483_, new_n481_, new_n482_ );
nand g282 ( new_n484_, new_n478_, new_n483_ );
nand g283 ( new_n485_, new_n476_, new_n477_, new_n481_, new_n482_ );
nand g284 ( new_n486_, new_n484_, new_n485_ );
nand g285 ( new_n487_, new_n486_, new_n470_ );
nand g286 ( new_n488_, new_n484_, keyIn_0_66, new_n485_ );
nand g287 ( new_n489_, new_n487_, new_n488_ );
not g288 ( new_n490_, N25 );
nand g289 ( new_n491_, new_n490_, N9 );
not g290 ( new_n492_, N9 );
nand g291 ( new_n493_, new_n492_, N25 );
nand g292 ( new_n494_, new_n491_, new_n493_ );
nand g293 ( new_n495_, new_n494_, keyIn_0_28 );
not g294 ( new_n496_, keyIn_0_28 );
nand g295 ( new_n497_, new_n491_, new_n493_, new_n496_ );
nand g296 ( new_n498_, new_n495_, new_n497_ );
not g297 ( new_n499_, N57 );
nand g298 ( new_n500_, new_n499_, N41 );
not g299 ( new_n501_, N41 );
nand g300 ( new_n502_, new_n501_, N57 );
nand g301 ( new_n503_, new_n500_, new_n502_ );
nand g302 ( new_n504_, new_n503_, keyIn_0_29 );
not g303 ( new_n505_, keyIn_0_29 );
nand g304 ( new_n506_, new_n500_, new_n502_, new_n505_ );
nand g305 ( new_n507_, new_n504_, new_n506_ );
nand g306 ( new_n508_, new_n498_, new_n507_ );
nand g307 ( new_n509_, new_n495_, new_n504_, new_n497_, new_n506_ );
nand g308 ( new_n510_, new_n508_, new_n509_ );
nand g309 ( new_n511_, new_n510_, keyIn_0_50 );
not g310 ( new_n512_, keyIn_0_50 );
nand g311 ( new_n513_, new_n508_, new_n512_, new_n509_ );
nand g312 ( new_n514_, new_n511_, new_n513_ );
nand g313 ( new_n515_, new_n489_, new_n514_ );
nand g314 ( new_n516_, new_n487_, new_n488_, new_n511_, new_n513_ );
nand g315 ( new_n517_, new_n515_, new_n516_ );
nand g316 ( new_n518_, new_n517_, new_n469_ );
nand g317 ( new_n519_, new_n515_, keyIn_0_74, new_n516_ );
nand g318 ( new_n520_, new_n518_, new_n519_ );
nand g319 ( new_n521_, new_n520_, keyIn_0_90 );
not g320 ( new_n522_, keyIn_0_90 );
nand g321 ( new_n523_, new_n518_, new_n522_, new_n519_ );
nand g322 ( new_n524_, new_n521_, new_n468_, new_n523_ );
nor g323 ( new_n525_, new_n467_, new_n524_ );
nor g324 ( new_n526_, new_n525_, keyIn_0_107 );
nand g325 ( new_n527_, new_n463_, keyIn_0_85 );
not g326 ( new_n528_, keyIn_0_85 );
nand g327 ( new_n529_, new_n458_, new_n528_, new_n460_ );
nand g328 ( new_n530_, new_n527_, new_n529_ );
not g329 ( new_n531_, keyIn_0_83 );
nand g330 ( new_n532_, new_n302_, new_n531_ );
nand g331 ( new_n533_, new_n300_, keyIn_0_83, new_n301_ );
nand g332 ( new_n534_, new_n532_, new_n533_ );
nand g333 ( new_n535_, new_n534_, new_n530_, new_n518_, new_n519_ );
nand g334 ( new_n536_, new_n409_, keyIn_0_84 );
not g335 ( new_n537_, keyIn_0_84 );
nand g336 ( new_n538_, new_n406_, new_n537_, new_n408_ );
nand g337 ( new_n539_, new_n536_, new_n538_ );
nor g338 ( new_n540_, new_n539_, new_n535_, keyIn_0_105 );
not g339 ( new_n541_, keyIn_0_105 );
nor g340 ( new_n542_, new_n539_, new_n535_ );
nor g341 ( new_n543_, new_n542_, new_n541_ );
nor g342 ( new_n544_, new_n526_, new_n543_, new_n540_ );
not g343 ( new_n545_, keyIn_0_104 );
nand g344 ( new_n546_, new_n409_, keyIn_0_81 );
not g345 ( new_n547_, keyIn_0_81 );
nand g346 ( new_n548_, new_n406_, new_n547_, new_n408_ );
nand g347 ( new_n549_, new_n546_, new_n548_ );
not g348 ( new_n550_, keyIn_0_82 );
not g349 ( new_n551_, new_n520_ );
nand g350 ( new_n552_, new_n551_, new_n550_ );
nand g351 ( new_n553_, new_n520_, keyIn_0_82 );
not g352 ( new_n554_, new_n553_ );
not g353 ( new_n555_, new_n463_ );
nand g354 ( new_n556_, new_n302_, keyIn_0_80 );
not g355 ( new_n557_, keyIn_0_80 );
nand g356 ( new_n558_, new_n300_, new_n557_, new_n301_ );
nand g357 ( new_n559_, new_n556_, new_n558_ );
nand g358 ( new_n560_, new_n559_, new_n555_ );
nor g359 ( new_n561_, new_n554_, new_n560_ );
nand g360 ( new_n562_, new_n561_, new_n545_, new_n549_, new_n552_ );
not g361 ( new_n563_, keyIn_0_88 );
nand g362 ( new_n564_, new_n463_, new_n563_ );
nand g363 ( new_n565_, new_n458_, keyIn_0_88, new_n460_ );
nand g364 ( new_n566_, new_n564_, new_n565_ );
nand g365 ( new_n567_, new_n300_, keyIn_0_86, new_n301_ );
not g366 ( new_n568_, keyIn_0_86 );
nand g367 ( new_n569_, new_n302_, new_n568_ );
nand g368 ( new_n570_, new_n569_, new_n567_ );
nor g369 ( new_n571_, new_n570_, new_n409_ );
nand g370 ( new_n572_, new_n520_, keyIn_0_87 );
not g371 ( new_n573_, keyIn_0_87 );
nand g372 ( new_n574_, new_n551_, new_n573_ );
nand g373 ( new_n575_, new_n574_, new_n571_, new_n566_, new_n572_ );
nand g374 ( new_n576_, new_n575_, keyIn_0_106 );
not g375 ( new_n577_, keyIn_0_106 );
not g376 ( new_n578_, new_n566_ );
nor g377 ( new_n579_, new_n578_, new_n409_, new_n570_ );
nand g378 ( new_n580_, new_n579_, new_n577_, new_n572_, new_n574_ );
nand g379 ( new_n581_, new_n576_, new_n580_ );
not g380 ( new_n582_, new_n524_ );
nand g381 ( new_n583_, new_n582_, keyIn_0_107, new_n410_, new_n466_ );
not g382 ( new_n584_, new_n560_ );
nand g383 ( new_n585_, new_n584_, new_n549_, new_n552_, new_n553_ );
nand g384 ( new_n586_, new_n585_, keyIn_0_104 );
nand g385 ( new_n587_, new_n586_, new_n583_ );
not g386 ( new_n588_, new_n587_ );
nand g387 ( new_n589_, new_n544_, new_n588_, new_n562_, new_n581_ );
nand g388 ( new_n590_, new_n589_, new_n304_ );
nand g389 ( new_n591_, new_n581_, new_n562_ );
not g390 ( new_n592_, new_n591_ );
nand g391 ( new_n593_, new_n592_, keyIn_0_112, new_n544_, new_n588_ );
not g392 ( new_n594_, keyIn_0_70 );
not g393 ( new_n595_, keyIn_0_42 );
nand g394 ( new_n596_, new_n389_, N33 );
not g395 ( new_n597_, N33 );
nand g396 ( new_n598_, new_n597_, N37 );
nand g397 ( new_n599_, new_n596_, new_n598_ );
nand g398 ( new_n600_, new_n599_, keyIn_0_4 );
not g399 ( new_n601_, keyIn_0_4 );
nand g400 ( new_n602_, new_n596_, new_n598_, new_n601_ );
nand g401 ( new_n603_, new_n600_, new_n602_ );
not g402 ( new_n604_, N45 );
nand g403 ( new_n605_, new_n604_, N41 );
nand g404 ( new_n606_, new_n501_, N45 );
nand g405 ( new_n607_, new_n605_, new_n606_ );
nand g406 ( new_n608_, new_n607_, keyIn_0_5 );
not g407 ( new_n609_, keyIn_0_5 );
nand g408 ( new_n610_, new_n605_, new_n606_, new_n609_ );
nand g409 ( new_n611_, new_n603_, new_n608_, new_n610_ );
nand g410 ( new_n612_, new_n608_, new_n610_ );
nand g411 ( new_n613_, new_n612_, new_n600_, new_n602_ );
nand g412 ( new_n614_, new_n611_, new_n613_ );
nand g413 ( new_n615_, new_n614_, new_n595_ );
nand g414 ( new_n616_, new_n611_, new_n613_, keyIn_0_42 );
nand g415 ( new_n617_, new_n615_, new_n616_ );
not g416 ( new_n618_, keyIn_0_40 );
not g417 ( new_n619_, N5 );
nand g418 ( new_n620_, new_n619_, N1 );
nand g419 ( new_n621_, new_n284_, N5 );
nand g420 ( new_n622_, new_n620_, new_n621_ );
nand g421 ( new_n623_, new_n622_, keyIn_0_0 );
not g422 ( new_n624_, keyIn_0_0 );
nand g423 ( new_n625_, new_n620_, new_n621_, new_n624_ );
nand g424 ( new_n626_, new_n623_, new_n625_ );
not g425 ( new_n627_, keyIn_0_1 );
nand g426 ( new_n628_, new_n441_, N9 );
nand g427 ( new_n629_, new_n492_, N13 );
nand g428 ( new_n630_, new_n628_, new_n629_ );
nand g429 ( new_n631_, new_n630_, new_n627_ );
nand g430 ( new_n632_, new_n628_, new_n629_, keyIn_0_1 );
nand g431 ( new_n633_, new_n626_, new_n631_, new_n632_ );
nand g432 ( new_n634_, new_n631_, new_n632_ );
nand g433 ( new_n635_, new_n634_, new_n623_, new_n625_ );
nand g434 ( new_n636_, new_n633_, new_n635_, new_n618_ );
nand g435 ( new_n637_, new_n633_, new_n635_ );
nand g436 ( new_n638_, new_n637_, keyIn_0_40 );
nand g437 ( new_n639_, new_n617_, new_n636_, new_n638_ );
nand g438 ( new_n640_, new_n638_, new_n636_ );
nand g439 ( new_n641_, new_n640_, new_n615_, new_n616_ );
nand g440 ( new_n642_, new_n639_, new_n641_ );
nand g441 ( new_n643_, new_n642_, keyIn_0_58 );
not g442 ( new_n644_, keyIn_0_58 );
nand g443 ( new_n645_, new_n639_, new_n641_, new_n644_ );
nand g444 ( new_n646_, keyIn_0_22, N135, N137 );
not g445 ( new_n647_, keyIn_0_22 );
nand g446 ( new_n648_, N135, N137 );
nand g447 ( new_n649_, new_n648_, new_n647_ );
nand g448 ( new_n650_, new_n649_, new_n646_ );
nand g449 ( new_n651_, new_n643_, new_n645_, new_n650_ );
nand g450 ( new_n652_, new_n643_, new_n645_ );
nand g451 ( new_n653_, new_n652_, new_n646_, new_n649_ );
nand g452 ( new_n654_, new_n653_, new_n651_ );
nand g453 ( new_n655_, new_n654_, new_n594_ );
nand g454 ( new_n656_, new_n653_, keyIn_0_70, new_n651_ );
not g455 ( new_n657_, keyIn_0_54 );
nand g456 ( new_n658_, new_n207_, N73 );
nand g457 ( new_n659_, new_n233_, N89 );
nand g458 ( new_n660_, new_n658_, new_n659_ );
nand g459 ( new_n661_, new_n660_, keyIn_0_36 );
not g460 ( new_n662_, keyIn_0_36 );
nand g461 ( new_n663_, new_n658_, new_n659_, new_n662_ );
nand g462 ( new_n664_, new_n661_, new_n663_ );
nand g463 ( new_n665_, new_n320_, N105 );
nand g464 ( new_n666_, new_n348_, N121 );
nand g465 ( new_n667_, new_n665_, new_n666_ );
nand g466 ( new_n668_, new_n667_, keyIn_0_37 );
not g467 ( new_n669_, keyIn_0_37 );
nand g468 ( new_n670_, new_n665_, new_n666_, new_n669_ );
nand g469 ( new_n671_, new_n668_, new_n670_ );
nand g470 ( new_n672_, new_n664_, new_n671_ );
nand g471 ( new_n673_, new_n661_, new_n668_, new_n663_, new_n670_ );
nand g472 ( new_n674_, new_n672_, new_n673_ );
nand g473 ( new_n675_, new_n674_, new_n657_ );
nand g474 ( new_n676_, new_n672_, keyIn_0_54, new_n673_ );
nand g475 ( new_n677_, new_n675_, new_n676_ );
nand g476 ( new_n678_, new_n655_, new_n656_, new_n677_ );
nand g477 ( new_n679_, new_n655_, new_n656_ );
nand g478 ( new_n680_, new_n679_, new_n675_, new_n676_ );
nand g479 ( new_n681_, new_n680_, new_n678_ );
nand g480 ( new_n682_, new_n681_, keyIn_0_78 );
not g481 ( new_n683_, keyIn_0_78 );
nand g482 ( new_n684_, new_n680_, new_n683_, new_n678_ );
nand g483 ( new_n685_, new_n682_, new_n684_ );
not g484 ( new_n686_, new_n685_ );
not g485 ( new_n687_, keyIn_0_71 );
not g486 ( new_n688_, keyIn_0_59 );
not g487 ( new_n689_, N61 );
nand g488 ( new_n690_, new_n689_, N57 );
nand g489 ( new_n691_, new_n499_, N61 );
nand g490 ( new_n692_, new_n690_, new_n691_ );
nand g491 ( new_n693_, new_n692_, keyIn_0_7 );
not g492 ( new_n694_, keyIn_0_7 );
nand g493 ( new_n695_, new_n690_, new_n691_, new_n694_ );
nand g494 ( new_n696_, new_n693_, new_n695_ );
nand g495 ( new_n697_, new_n387_, N49 );
not g496 ( new_n698_, N49 );
nand g497 ( new_n699_, new_n698_, N53 );
nand g498 ( new_n700_, new_n697_, new_n699_ );
nand g499 ( new_n701_, new_n700_, keyIn_0_6 );
not g500 ( new_n702_, keyIn_0_6 );
nand g501 ( new_n703_, new_n697_, new_n699_, new_n702_ );
nand g502 ( new_n704_, new_n696_, new_n701_, new_n703_ );
nand g503 ( new_n705_, new_n701_, new_n703_ );
nand g504 ( new_n706_, new_n705_, new_n693_, new_n695_ );
nand g505 ( new_n707_, new_n704_, new_n706_ );
nand g506 ( new_n708_, new_n707_, keyIn_0_43 );
not g507 ( new_n709_, keyIn_0_43 );
nand g508 ( new_n710_, new_n704_, new_n706_, new_n709_ );
nand g509 ( new_n711_, new_n708_, new_n710_ );
not g510 ( new_n712_, keyIn_0_41 );
not g511 ( new_n713_, N21 );
nand g512 ( new_n714_, new_n713_, N17 );
nand g513 ( new_n715_, new_n282_, N21 );
nand g514 ( new_n716_, new_n714_, new_n715_ );
nand g515 ( new_n717_, new_n716_, keyIn_0_2 );
not g516 ( new_n718_, keyIn_0_2 );
nand g517 ( new_n719_, new_n714_, new_n715_, new_n718_ );
nand g518 ( new_n720_, new_n717_, new_n719_ );
nand g519 ( new_n721_, new_n439_, N25 );
nand g520 ( new_n722_, new_n490_, N29 );
nand g521 ( new_n723_, new_n721_, new_n722_ );
nand g522 ( new_n724_, new_n723_, keyIn_0_3 );
not g523 ( new_n725_, keyIn_0_3 );
nand g524 ( new_n726_, new_n721_, new_n722_, new_n725_ );
nand g525 ( new_n727_, new_n724_, new_n726_ );
nand g526 ( new_n728_, new_n720_, new_n727_ );
nand g527 ( new_n729_, new_n717_, new_n724_, new_n719_, new_n726_ );
nand g528 ( new_n730_, new_n728_, new_n729_ );
nand g529 ( new_n731_, new_n730_, new_n712_ );
nand g530 ( new_n732_, new_n728_, keyIn_0_41, new_n729_ );
nand g531 ( new_n733_, new_n711_, new_n731_, new_n732_ );
nand g532 ( new_n734_, new_n731_, new_n732_ );
nand g533 ( new_n735_, new_n734_, new_n708_, new_n710_ );
nand g534 ( new_n736_, new_n733_, new_n735_ );
nand g535 ( new_n737_, new_n736_, new_n688_ );
nand g536 ( new_n738_, new_n733_, keyIn_0_59, new_n735_ );
not g537 ( new_n739_, keyIn_0_23 );
nand g538 ( new_n740_, new_n739_, N136, N137 );
nand g539 ( new_n741_, N136, N137 );
nand g540 ( new_n742_, new_n741_, keyIn_0_23 );
nand g541 ( new_n743_, new_n742_, new_n740_ );
nand g542 ( new_n744_, new_n737_, new_n738_, new_n743_ );
nand g543 ( new_n745_, new_n737_, new_n738_ );
nand g544 ( new_n746_, new_n745_, new_n740_, new_n742_ );
nand g545 ( new_n747_, new_n746_, new_n744_ );
nand g546 ( new_n748_, new_n747_, new_n687_ );
nand g547 ( new_n749_, new_n746_, keyIn_0_71, new_n744_ );
nor g548 ( new_n750_, N77, N93 );
not g549 ( new_n751_, new_n750_ );
nand g550 ( new_n752_, N77, N93 );
nand g551 ( new_n753_, new_n751_, new_n752_ );
nand g552 ( new_n754_, new_n753_, keyIn_0_38 );
not g553 ( new_n755_, new_n754_ );
nor g554 ( new_n756_, new_n753_, keyIn_0_38 );
nor g555 ( new_n757_, new_n755_, new_n756_ );
not g556 ( new_n758_, new_n757_ );
nand g557 ( new_n759_, new_n318_, N109 );
nand g558 ( new_n760_, new_n350_, N125 );
nand g559 ( new_n761_, new_n759_, new_n760_ );
nand g560 ( new_n762_, new_n761_, keyIn_0_39 );
not g561 ( new_n763_, keyIn_0_39 );
nand g562 ( new_n764_, new_n759_, new_n760_, new_n763_ );
nand g563 ( new_n765_, new_n762_, new_n764_ );
nand g564 ( new_n766_, new_n758_, new_n765_ );
nand g565 ( new_n767_, new_n757_, new_n762_, new_n764_ );
nand g566 ( new_n768_, new_n766_, new_n767_ );
nand g567 ( new_n769_, new_n768_, keyIn_0_55 );
not g568 ( new_n770_, keyIn_0_55 );
nand g569 ( new_n771_, new_n766_, new_n770_, new_n767_ );
nand g570 ( new_n772_, new_n769_, new_n771_ );
nand g571 ( new_n773_, new_n748_, new_n749_, new_n772_ );
nand g572 ( new_n774_, new_n748_, new_n749_ );
not g573 ( new_n775_, new_n772_ );
nand g574 ( new_n776_, new_n774_, new_n775_ );
nand g575 ( new_n777_, new_n776_, new_n773_ );
nand g576 ( new_n778_, new_n777_, keyIn_0_79 );
not g577 ( new_n779_, keyIn_0_79 );
nand g578 ( new_n780_, new_n776_, new_n779_, new_n773_ );
nand g579 ( new_n781_, new_n686_, new_n778_, new_n780_ );
not g580 ( new_n782_, keyIn_0_76 );
not g581 ( new_n783_, keyIn_0_68 );
nand g582 ( new_n784_, new_n640_, new_n734_ );
nand g583 ( new_n785_, new_n638_, new_n731_, new_n636_, new_n732_ );
nand g584 ( new_n786_, new_n784_, new_n785_ );
nand g585 ( new_n787_, new_n786_, keyIn_0_56 );
not g586 ( new_n788_, keyIn_0_56 );
nand g587 ( new_n789_, new_n784_, new_n788_, new_n785_ );
nand g588 ( new_n790_, new_n787_, new_n789_ );
not g589 ( new_n791_, keyIn_0_20 );
nand g590 ( new_n792_, N133, N137 );
nand g591 ( new_n793_, new_n792_, new_n791_ );
nand g592 ( new_n794_, keyIn_0_20, N133, N137 );
nand g593 ( new_n795_, new_n793_, new_n794_ );
nand g594 ( new_n796_, new_n790_, new_n795_ );
nand g595 ( new_n797_, new_n787_, new_n789_, new_n793_, new_n794_ );
nand g596 ( new_n798_, new_n796_, new_n797_ );
nand g597 ( new_n799_, new_n798_, new_n783_ );
nand g598 ( new_n800_, new_n796_, keyIn_0_68, new_n797_ );
nand g599 ( new_n801_, new_n799_, new_n800_ );
nand g600 ( new_n802_, new_n214_, N65 );
nand g601 ( new_n803_, new_n241_, N81 );
nand g602 ( new_n804_, new_n802_, new_n803_ );
nand g603 ( new_n805_, new_n804_, keyIn_0_32 );
not g604 ( new_n806_, keyIn_0_32 );
nand g605 ( new_n807_, new_n802_, new_n803_, new_n806_ );
nand g606 ( new_n808_, new_n805_, new_n807_ );
nand g607 ( new_n809_, new_n311_, N97 );
nand g608 ( new_n810_, new_n337_, N113 );
nand g609 ( new_n811_, new_n809_, new_n810_ );
nand g610 ( new_n812_, new_n811_, keyIn_0_33 );
not g611 ( new_n813_, keyIn_0_33 );
nand g612 ( new_n814_, new_n809_, new_n810_, new_n813_ );
nand g613 ( new_n815_, new_n812_, new_n814_ );
nand g614 ( new_n816_, new_n808_, new_n815_ );
nand g615 ( new_n817_, new_n805_, new_n812_, new_n807_, new_n814_ );
nand g616 ( new_n818_, new_n816_, new_n817_ );
nand g617 ( new_n819_, new_n818_, keyIn_0_52 );
not g618 ( new_n820_, keyIn_0_52 );
nand g619 ( new_n821_, new_n816_, new_n820_, new_n817_ );
nand g620 ( new_n822_, new_n819_, new_n821_ );
nand g621 ( new_n823_, new_n801_, new_n822_ );
nand g622 ( new_n824_, new_n799_, new_n800_, new_n819_, new_n821_ );
nand g623 ( new_n825_, new_n823_, new_n824_ );
nand g624 ( new_n826_, new_n825_, new_n782_ );
nand g625 ( new_n827_, new_n823_, keyIn_0_76, new_n824_ );
nand g626 ( new_n828_, new_n826_, new_n827_ );
not g627 ( new_n829_, keyIn_0_69 );
not g628 ( new_n830_, keyIn_0_57 );
nand g629 ( new_n831_, new_n617_, new_n711_ );
nand g630 ( new_n832_, new_n615_, new_n708_, new_n616_, new_n710_ );
nand g631 ( new_n833_, new_n831_, new_n832_ );
nand g632 ( new_n834_, new_n833_, new_n830_ );
nand g633 ( new_n835_, new_n831_, keyIn_0_57, new_n832_ );
nand g634 ( new_n836_, new_n834_, new_n835_ );
nand g635 ( new_n837_, N134, N137 );
nand g636 ( new_n838_, new_n837_, keyIn_0_21 );
not g637 ( new_n839_, keyIn_0_21 );
nand g638 ( new_n840_, new_n839_, N134, N137 );
nand g639 ( new_n841_, new_n838_, new_n840_ );
nand g640 ( new_n842_, new_n836_, new_n841_ );
nand g641 ( new_n843_, new_n834_, new_n835_, new_n838_, new_n840_ );
nand g642 ( new_n844_, new_n842_, new_n843_ );
nand g643 ( new_n845_, new_n844_, new_n829_ );
nand g644 ( new_n846_, new_n842_, keyIn_0_69, new_n843_ );
nor g645 ( new_n847_, N69, N85 );
not g646 ( new_n848_, new_n847_ );
nand g647 ( new_n849_, N69, N85 );
nand g648 ( new_n850_, new_n848_, new_n849_ );
nand g649 ( new_n851_, new_n850_, keyIn_0_34 );
not g650 ( new_n852_, new_n851_ );
nor g651 ( new_n853_, new_n850_, keyIn_0_34 );
nor g652 ( new_n854_, new_n852_, new_n853_ );
not g653 ( new_n855_, new_n854_ );
nor g654 ( new_n856_, N101, N117 );
not g655 ( new_n857_, new_n856_ );
nand g656 ( new_n858_, N101, N117 );
nand g657 ( new_n859_, new_n857_, new_n858_ );
nand g658 ( new_n860_, new_n859_, keyIn_0_35 );
not g659 ( new_n861_, new_n860_ );
nor g660 ( new_n862_, new_n859_, keyIn_0_35 );
nor g661 ( new_n863_, new_n861_, new_n862_ );
not g662 ( new_n864_, new_n863_ );
nand g663 ( new_n865_, new_n855_, new_n864_ );
nand g664 ( new_n866_, new_n854_, new_n863_ );
nand g665 ( new_n867_, new_n865_, new_n866_ );
nand g666 ( new_n868_, new_n867_, keyIn_0_53 );
not g667 ( new_n869_, keyIn_0_53 );
nand g668 ( new_n870_, new_n865_, new_n869_, new_n866_ );
nand g669 ( new_n871_, new_n868_, new_n870_ );
nand g670 ( new_n872_, new_n845_, new_n846_, new_n871_ );
nand g671 ( new_n873_, new_n845_, new_n846_ );
nand g672 ( new_n874_, new_n873_, new_n868_, new_n870_ );
nand g673 ( new_n875_, new_n874_, new_n872_ );
nand g674 ( new_n876_, new_n875_, keyIn_0_77 );
not g675 ( new_n877_, keyIn_0_77 );
nand g676 ( new_n878_, new_n874_, new_n877_, new_n872_ );
nand g677 ( new_n879_, new_n828_, new_n876_, new_n878_ );
nor g678 ( new_n880_, new_n781_, new_n879_ );
nand g679 ( new_n881_, new_n590_, keyIn_0_114, new_n593_, new_n880_ );
not g680 ( new_n882_, keyIn_0_114 );
nand g681 ( new_n883_, new_n590_, new_n593_, new_n880_ );
nand g682 ( new_n884_, new_n883_, new_n882_ );
nand g683 ( new_n885_, new_n884_, new_n303_, new_n881_ );
nand g684 ( new_n886_, new_n885_, N1 );
nand g685 ( new_n887_, new_n884_, new_n284_, new_n303_, new_n881_ );
nand g686 ( N724, new_n886_, new_n887_ );
not g687 ( new_n889_, new_n409_ );
nand g688 ( new_n890_, new_n884_, new_n889_, new_n881_ );
nand g689 ( new_n891_, new_n890_, N5 );
nand g690 ( new_n892_, new_n884_, new_n619_, new_n889_, new_n881_ );
nand g691 ( N725, new_n891_, new_n892_ );
nand g692 ( new_n894_, new_n884_, new_n551_, new_n881_ );
nand g693 ( new_n895_, new_n894_, N9 );
nand g694 ( new_n896_, new_n884_, new_n492_, new_n551_, new_n881_ );
nand g695 ( N726, new_n895_, new_n896_ );
nand g696 ( new_n898_, new_n884_, new_n555_, new_n881_ );
nand g697 ( new_n899_, new_n898_, N13 );
nand g698 ( new_n900_, new_n884_, new_n441_, new_n555_, new_n881_ );
nand g699 ( N727, new_n899_, new_n900_ );
not g700 ( new_n902_, keyIn_0_115 );
nand g701 ( new_n903_, new_n778_, new_n780_ );
nand g702 ( new_n904_, new_n685_, new_n903_ );
nor g703 ( new_n905_, new_n904_, new_n879_ );
nand g704 ( new_n906_, new_n590_, new_n902_, new_n593_, new_n905_ );
nand g705 ( new_n907_, new_n590_, new_n593_, new_n905_ );
nand g706 ( new_n908_, new_n907_, keyIn_0_115 );
nand g707 ( new_n909_, new_n908_, new_n303_, new_n906_ );
nand g708 ( new_n910_, new_n909_, N17 );
nand g709 ( new_n911_, new_n908_, new_n282_, new_n303_, new_n906_ );
nand g710 ( N728, new_n910_, new_n911_ );
nand g711 ( new_n913_, new_n908_, new_n889_, new_n906_ );
nand g712 ( new_n914_, new_n913_, N21 );
nand g713 ( new_n915_, new_n908_, new_n713_, new_n889_, new_n906_ );
nand g714 ( N729, new_n914_, new_n915_ );
nand g715 ( new_n917_, new_n908_, new_n551_, new_n906_ );
nand g716 ( new_n918_, new_n917_, N25 );
nand g717 ( new_n919_, new_n908_, new_n490_, new_n551_, new_n906_ );
nand g718 ( N730, new_n918_, new_n919_ );
nand g719 ( new_n921_, new_n908_, new_n555_, new_n906_ );
nand g720 ( new_n922_, new_n921_, N29 );
nand g721 ( new_n923_, new_n908_, new_n439_, new_n555_, new_n906_ );
nand g722 ( N731, new_n922_, new_n923_ );
not g723 ( new_n925_, keyIn_0_116 );
nand g724 ( new_n926_, new_n876_, new_n878_ );
nand g725 ( new_n927_, new_n926_, new_n826_, new_n827_ );
nor g726 ( new_n928_, new_n781_, new_n927_ );
nand g727 ( new_n929_, new_n590_, new_n593_, new_n928_ );
nand g728 ( new_n930_, new_n929_, new_n925_ );
nand g729 ( new_n931_, new_n590_, keyIn_0_116, new_n593_, new_n928_ );
nand g730 ( new_n932_, new_n930_, new_n931_ );
nand g731 ( new_n933_, new_n932_, new_n303_ );
nand g732 ( new_n934_, new_n933_, N33 );
nand g733 ( new_n935_, new_n932_, new_n597_, new_n303_ );
nand g734 ( N732, new_n934_, new_n935_ );
nand g735 ( new_n937_, new_n932_, new_n889_ );
nand g736 ( new_n938_, new_n937_, N37 );
nand g737 ( new_n939_, new_n932_, new_n389_, new_n889_ );
nand g738 ( N733, new_n938_, new_n939_ );
nand g739 ( new_n941_, new_n932_, new_n551_ );
nand g740 ( new_n942_, new_n941_, N41 );
nand g741 ( new_n943_, new_n932_, new_n501_, new_n551_ );
nand g742 ( N734, new_n942_, new_n943_ );
nand g743 ( new_n945_, new_n932_, new_n555_ );
nand g744 ( new_n946_, new_n945_, N45 );
nand g745 ( new_n947_, new_n932_, new_n604_, new_n555_ );
nand g746 ( N735, new_n946_, new_n947_ );
not g747 ( new_n949_, keyIn_0_117 );
nor g748 ( new_n950_, new_n904_, new_n927_ );
nand g749 ( new_n951_, new_n590_, new_n593_, new_n950_ );
nand g750 ( new_n952_, new_n951_, new_n949_ );
nand g751 ( new_n953_, new_n590_, keyIn_0_117, new_n593_, new_n950_ );
nand g752 ( new_n954_, new_n952_, new_n953_ );
nand g753 ( new_n955_, new_n954_, new_n303_ );
nand g754 ( new_n956_, new_n955_, N49 );
nand g755 ( new_n957_, new_n954_, new_n698_, new_n303_ );
nand g756 ( N736, new_n956_, new_n957_ );
nand g757 ( new_n959_, new_n954_, new_n889_ );
nand g758 ( new_n960_, new_n959_, N53 );
nand g759 ( new_n961_, new_n954_, new_n387_, new_n889_ );
nand g760 ( N737, new_n960_, new_n961_ );
nand g761 ( new_n963_, new_n954_, new_n551_ );
nand g762 ( new_n964_, new_n963_, N57 );
nand g763 ( new_n965_, new_n954_, new_n499_, new_n551_ );
nand g764 ( N738, new_n964_, new_n965_ );
nand g765 ( new_n967_, new_n954_, new_n555_ );
nand g766 ( new_n968_, new_n967_, keyIn_0_122 );
not g767 ( new_n969_, keyIn_0_122 );
nand g768 ( new_n970_, new_n954_, new_n969_, new_n555_ );
nand g769 ( new_n971_, new_n968_, new_n970_ );
nand g770 ( new_n972_, new_n971_, new_n689_ );
nand g771 ( new_n973_, new_n968_, N61, new_n970_ );
nand g772 ( N739, new_n972_, new_n973_ );
not g773 ( new_n975_, keyIn_0_109 );
not g774 ( new_n976_, keyIn_0_97 );
nand g775 ( new_n977_, new_n778_, new_n976_, new_n780_ );
nand g776 ( new_n978_, new_n903_, keyIn_0_97 );
nand g777 ( new_n979_, new_n686_, new_n978_, new_n977_ );
not g778 ( new_n980_, keyIn_0_96 );
nand g779 ( new_n981_, new_n926_, new_n980_ );
nand g780 ( new_n982_, new_n876_, keyIn_0_96, new_n878_ );
nand g781 ( new_n983_, new_n981_, new_n982_ );
not g782 ( new_n984_, keyIn_0_95 );
nand g783 ( new_n985_, new_n828_, new_n984_ );
nand g784 ( new_n986_, new_n826_, keyIn_0_95, new_n827_ );
nand g785 ( new_n987_, new_n985_, new_n986_ );
nand g786 ( new_n988_, new_n983_, new_n987_ );
nor g787 ( new_n989_, new_n988_, new_n979_, new_n975_ );
nor g788 ( new_n990_, new_n988_, new_n979_ );
nor g789 ( new_n991_, new_n990_, keyIn_0_109 );
nor g790 ( new_n992_, new_n991_, new_n989_ );
not g791 ( new_n993_, keyIn_0_108 );
not g792 ( new_n994_, keyIn_0_92 );
nand g793 ( new_n995_, new_n828_, new_n994_ );
not g794 ( new_n996_, new_n995_ );
nand g795 ( new_n997_, new_n826_, keyIn_0_92, new_n827_ );
nand g796 ( new_n998_, new_n903_, new_n997_ );
nor g797 ( new_n999_, new_n996_, new_n998_ );
nand g798 ( new_n1000_, new_n926_, keyIn_0_93 );
not g799 ( new_n1001_, keyIn_0_93 );
nand g800 ( new_n1002_, new_n876_, new_n1001_, new_n878_ );
nand g801 ( new_n1003_, new_n1000_, new_n1002_ );
nand g802 ( new_n1004_, new_n685_, keyIn_0_94 );
not g803 ( new_n1005_, keyIn_0_94 );
nand g804 ( new_n1006_, new_n682_, new_n1005_, new_n684_ );
nand g805 ( new_n1007_, new_n1004_, new_n1006_ );
nand g806 ( new_n1008_, new_n999_, new_n1007_, new_n1003_ );
nand g807 ( new_n1009_, new_n1008_, new_n993_ );
nand g808 ( new_n1010_, new_n999_, new_n1007_, keyIn_0_108, new_n1003_ );
nand g809 ( new_n1011_, new_n1009_, new_n1010_ );
not g810 ( new_n1012_, new_n1011_ );
not g811 ( new_n1013_, keyIn_0_111 );
not g812 ( new_n1014_, keyIn_0_101 );
nand g813 ( new_n1015_, new_n876_, new_n1014_, new_n878_ );
nand g814 ( new_n1016_, new_n903_, keyIn_0_103 );
not g815 ( new_n1017_, keyIn_0_103 );
nand g816 ( new_n1018_, new_n778_, new_n1017_, new_n780_ );
nand g817 ( new_n1019_, new_n1016_, new_n1015_, new_n1018_ );
not g818 ( new_n1020_, new_n1019_ );
nand g819 ( new_n1021_, new_n686_, keyIn_0_102 );
not g820 ( new_n1022_, keyIn_0_102 );
nand g821 ( new_n1023_, new_n685_, new_n1022_ );
nand g822 ( new_n1024_, new_n1021_, new_n1023_ );
nand g823 ( new_n1025_, new_n926_, keyIn_0_101 );
nand g824 ( new_n1026_, new_n1025_, new_n828_ );
not g825 ( new_n1027_, new_n1026_ );
nand g826 ( new_n1028_, new_n1024_, new_n1020_, new_n1027_ );
nand g827 ( new_n1029_, new_n1028_, new_n1013_ );
nand g828 ( new_n1030_, new_n1024_, new_n1020_, keyIn_0_111, new_n1027_ );
nand g829 ( new_n1031_, new_n1029_, new_n1030_ );
not g830 ( new_n1032_, keyIn_0_99 );
nand g831 ( new_n1033_, new_n682_, new_n1032_, new_n684_ );
nand g832 ( new_n1034_, new_n685_, keyIn_0_99 );
not g833 ( new_n1035_, keyIn_0_100 );
nand g834 ( new_n1036_, new_n778_, new_n1035_, new_n780_ );
nand g835 ( new_n1037_, new_n1034_, new_n1033_, new_n1036_ );
not g836 ( new_n1038_, keyIn_0_98 );
nand g837 ( new_n1039_, new_n828_, new_n1038_ );
nand g838 ( new_n1040_, new_n826_, keyIn_0_98, new_n827_ );
nand g839 ( new_n1041_, new_n1039_, new_n1040_ );
nand g840 ( new_n1042_, new_n903_, keyIn_0_100 );
nand g841 ( new_n1043_, new_n1041_, new_n926_, new_n1042_ );
nor g842 ( new_n1044_, new_n1043_, new_n1037_ );
nor g843 ( new_n1045_, new_n1044_, keyIn_0_110 );
not g844 ( new_n1046_, keyIn_0_110 );
nor g845 ( new_n1047_, new_n1043_, new_n1037_, new_n1046_ );
nor g846 ( new_n1048_, new_n1045_, new_n1047_ );
nand g847 ( new_n1049_, new_n992_, new_n1012_, new_n1048_, new_n1031_ );
nand g848 ( new_n1050_, new_n1049_, keyIn_0_113 );
not g849 ( new_n1051_, keyIn_0_113 );
nor g850 ( new_n1052_, new_n1011_, new_n991_, new_n989_ );
nand g851 ( new_n1053_, new_n1052_, new_n1051_, new_n1031_, new_n1048_ );
nand g852 ( new_n1054_, new_n1050_, new_n1053_ );
nand g853 ( new_n1055_, new_n551_, new_n463_ );
nor g854 ( new_n1056_, new_n1055_, new_n889_, new_n302_ );
nand g855 ( new_n1057_, new_n1054_, new_n1056_ );
nand g856 ( new_n1058_, new_n1057_, keyIn_0_118 );
not g857 ( new_n1059_, keyIn_0_118 );
nand g858 ( new_n1060_, new_n1054_, new_n1059_, new_n1056_ );
nand g859 ( new_n1061_, new_n1058_, new_n1060_ );
nand g860 ( new_n1062_, new_n1061_, new_n828_ );
nand g861 ( new_n1063_, new_n1062_, keyIn_0_123 );
not g862 ( new_n1064_, keyIn_0_123 );
nand g863 ( new_n1065_, new_n1061_, new_n1064_, new_n828_ );
nand g864 ( new_n1066_, new_n1063_, new_n1065_ );
nand g865 ( new_n1067_, new_n1066_, N65 );
nand g866 ( new_n1068_, new_n1063_, new_n241_, new_n1065_ );
nand g867 ( N740, new_n1067_, new_n1068_ );
not g868 ( new_n1070_, keyIn_0_124 );
nand g869 ( new_n1071_, new_n1061_, new_n926_ );
nand g870 ( new_n1072_, new_n1071_, new_n1070_ );
nand g871 ( new_n1073_, new_n1061_, keyIn_0_124, new_n926_ );
nand g872 ( new_n1074_, new_n1072_, new_n1073_ );
nand g873 ( new_n1075_, new_n1074_, new_n239_ );
nand g874 ( new_n1076_, new_n1072_, N69, new_n1073_ );
nand g875 ( N741, new_n1075_, new_n1076_ );
not g876 ( new_n1078_, keyIn_0_125 );
nand g877 ( new_n1079_, new_n1061_, new_n686_ );
nand g878 ( new_n1080_, new_n1079_, new_n1078_ );
nand g879 ( new_n1081_, new_n1061_, keyIn_0_125, new_n686_ );
nand g880 ( new_n1082_, new_n1080_, new_n1081_ );
nand g881 ( new_n1083_, new_n1082_, N73 );
nand g882 ( new_n1084_, new_n1080_, new_n233_, new_n1081_ );
nand g883 ( N742, new_n1083_, new_n1084_ );
not g884 ( new_n1086_, keyIn_0_126 );
nand g885 ( new_n1087_, new_n1061_, new_n903_ );
nand g886 ( new_n1088_, new_n1087_, new_n1086_ );
nand g887 ( new_n1089_, new_n1061_, keyIn_0_126, new_n903_ );
nand g888 ( new_n1090_, new_n1088_, new_n1089_ );
nand g889 ( new_n1091_, new_n1090_, new_n231_ );
nand g890 ( new_n1092_, new_n1088_, N77, new_n1089_ );
nand g891 ( N743, new_n1091_, new_n1092_ );
nand g892 ( new_n1094_, new_n409_, new_n520_, new_n555_, new_n303_ );
not g893 ( new_n1095_, new_n1094_ );
nand g894 ( new_n1096_, new_n1054_, new_n1095_ );
nand g895 ( new_n1097_, new_n1096_, keyIn_0_119 );
not g896 ( new_n1098_, keyIn_0_119 );
nand g897 ( new_n1099_, new_n1054_, new_n1098_, new_n1095_ );
nand g898 ( new_n1100_, new_n1097_, new_n1099_ );
nand g899 ( new_n1101_, new_n1100_, new_n828_ );
nand g900 ( new_n1102_, new_n1101_, keyIn_0_127 );
not g901 ( new_n1103_, keyIn_0_127 );
nand g902 ( new_n1104_, new_n1100_, new_n1103_, new_n828_ );
nand g903 ( new_n1105_, new_n1102_, new_n1104_ );
nand g904 ( new_n1106_, new_n1105_, N81 );
nand g905 ( new_n1107_, new_n1102_, new_n214_, new_n1104_ );
nand g906 ( N744, new_n1106_, new_n1107_ );
nand g907 ( new_n1109_, new_n1100_, new_n926_ );
nand g908 ( new_n1110_, new_n1109_, N85 );
nand g909 ( new_n1111_, new_n1100_, new_n215_, new_n926_ );
nand g910 ( N745, new_n1110_, new_n1111_ );
nand g911 ( new_n1113_, new_n1100_, new_n686_ );
nand g912 ( new_n1114_, new_n1113_, N89 );
nand g913 ( new_n1115_, new_n1100_, new_n207_, new_n686_ );
nand g914 ( N746, new_n1114_, new_n1115_ );
nand g915 ( new_n1117_, new_n1100_, new_n903_ );
nand g916 ( new_n1118_, new_n1117_, N93 );
nand g917 ( new_n1119_, new_n1100_, new_n205_, new_n903_ );
nand g918 ( N747, new_n1118_, new_n1119_ );
not g919 ( new_n1121_, keyIn_0_120 );
nand g920 ( new_n1122_, new_n889_, new_n302_ );
nor g921 ( new_n1123_, new_n1055_, new_n1122_ );
nand g922 ( new_n1124_, new_n1054_, new_n1123_ );
nand g923 ( new_n1125_, new_n1124_, new_n1121_ );
nand g924 ( new_n1126_, new_n1054_, keyIn_0_120, new_n1123_ );
nand g925 ( new_n1127_, new_n1125_, new_n1126_ );
nand g926 ( new_n1128_, new_n1127_, new_n828_ );
nand g927 ( new_n1129_, new_n1128_, N97 );
nand g928 ( new_n1130_, new_n1127_, new_n337_, new_n828_ );
nand g929 ( N748, new_n1129_, new_n1130_ );
nand g930 ( new_n1132_, new_n1127_, new_n926_ );
nand g931 ( new_n1133_, new_n1132_, N101 );
nand g932 ( new_n1134_, new_n1127_, new_n335_, new_n926_ );
nand g933 ( N749, new_n1133_, new_n1134_ );
nand g934 ( new_n1136_, new_n1127_, new_n686_ );
nand g935 ( new_n1137_, new_n1136_, N105 );
nand g936 ( new_n1138_, new_n1127_, new_n348_, new_n686_ );
nand g937 ( N750, new_n1137_, new_n1138_ );
nand g938 ( new_n1140_, new_n1127_, new_n903_ );
nand g939 ( new_n1141_, new_n1140_, N109 );
nand g940 ( new_n1142_, new_n1127_, new_n350_, new_n903_ );
nand g941 ( N751, new_n1141_, new_n1142_ );
nor g942 ( new_n1144_, new_n1122_, new_n463_, new_n551_ );
nand g943 ( new_n1145_, new_n1054_, new_n1144_ );
nand g944 ( new_n1146_, new_n1145_, keyIn_0_121 );
not g945 ( new_n1147_, keyIn_0_121 );
nand g946 ( new_n1148_, new_n1054_, new_n1147_, new_n1144_ );
nand g947 ( new_n1149_, new_n1146_, new_n1148_ );
nand g948 ( new_n1150_, new_n1149_, new_n828_ );
nand g949 ( new_n1151_, new_n1150_, N113 );
nand g950 ( new_n1152_, new_n1149_, new_n311_, new_n828_ );
nand g951 ( N752, new_n1151_, new_n1152_ );
nand g952 ( new_n1154_, new_n1149_, new_n926_ );
nand g953 ( new_n1155_, new_n1154_, N117 );
nand g954 ( new_n1156_, new_n1149_, new_n309_, new_n926_ );
nand g955 ( N753, new_n1155_, new_n1156_ );
nand g956 ( new_n1158_, new_n1149_, new_n686_ );
nand g957 ( new_n1159_, new_n1158_, N121 );
nand g958 ( new_n1160_, new_n1149_, new_n320_, new_n686_ );
nand g959 ( N754, new_n1159_, new_n1160_ );
nand g960 ( new_n1162_, new_n1149_, new_n903_ );
nand g961 ( new_n1163_, new_n1162_, N125 );
nand g962 ( new_n1164_, new_n1149_, new_n318_, new_n903_ );
nand g963 ( N755, new_n1163_, new_n1164_ );
endmodule