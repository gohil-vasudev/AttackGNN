module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n170_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n735_, new_n500_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n716_, new_n701_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n628_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n724_, new_n176_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n310_, new_n275_, new_n352_, new_n575_, new_n562_, new_n525_, new_n578_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n407_, new_n666_, new_n480_, new_n625_, new_n730_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n662_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n307_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n727_, new_n375_, new_n294_, new_n627_, new_n704_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n697_, new_n185_, new_n709_, new_n373_, new_n540_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n573_, new_n405_;

not g000 ( new_n151_, N75 );
nand g001 ( new_n152_, N29, N42 );
nor g002 ( N388, new_n152_, new_n151_ );
not g003 ( new_n154_, N80 );
nand g004 ( new_n155_, N29, N36 );
nor g005 ( N389, new_n155_, new_n154_ );
not g006 ( new_n157_, N42 );
nor g007 ( N390, new_n155_, new_n157_ );
nand g008 ( new_n159_, N85, N86 );
not g009 ( N391, new_n159_ );
not g010 ( new_n161_, N17 );
not g011 ( new_n162_, N13 );
nand g012 ( new_n163_, N1, N8 );
nor g013 ( new_n164_, new_n163_, new_n162_ );
not g014 ( new_n165_, new_n164_ );
nor g015 ( N418, new_n165_, new_n161_ );
not g016 ( new_n167_, N390 );
nand g017 ( new_n168_, N1, N26 );
nand g018 ( new_n169_, N13, N17 );
nor g019 ( new_n170_, new_n168_, new_n169_ );
nand g020 ( N419, new_n167_, new_n170_ );
nand g021 ( new_n172_, N59, N75 );
not g022 ( new_n173_, new_n172_ );
nand g023 ( N420, new_n173_, N80 );
nand g024 ( new_n175_, N36, N59 );
not g025 ( new_n176_, new_n175_ );
nand g026 ( N421, new_n176_, N80 );
nand g027 ( N422, new_n176_, N42 );
not g028 ( new_n179_, N90 );
nor g029 ( new_n180_, N87, N88 );
nor g030 ( N423, new_n180_, new_n179_ );
nand g031 ( N446, new_n170_, N390 );
not g032 ( new_n183_, new_n168_ );
nand g033 ( new_n184_, new_n183_, N51 );
nand g034 ( new_n185_, new_n184_, keyIn_0_0 );
not g035 ( new_n186_, keyIn_0_0 );
not g036 ( new_n187_, N51 );
nor g037 ( new_n188_, new_n168_, new_n187_ );
nand g038 ( new_n189_, new_n188_, new_n186_ );
nand g039 ( N447, new_n185_, new_n189_ );
not g040 ( new_n191_, N55 );
nor g041 ( new_n192_, new_n165_, new_n191_ );
not g042 ( new_n193_, new_n192_ );
nand g043 ( new_n194_, N29, N68 );
nor g044 ( N448, new_n193_, new_n194_ );
not g045 ( new_n196_, N74 );
nand g046 ( new_n197_, N59, N68 );
nor g047 ( new_n198_, new_n193_, new_n197_ );
not g048 ( new_n199_, new_n198_ );
nor g049 ( N449, new_n199_, new_n196_ );
not g050 ( new_n201_, N89 );
nor g051 ( N450, new_n180_, new_n201_ );
xor g052 ( new_n203_, N111, N116 );
xnor g053 ( new_n204_, N121, N126 );
xnor g054 ( new_n205_, new_n203_, new_n204_ );
nor g055 ( new_n206_, new_n205_, N135 );
xor g056 ( new_n207_, new_n206_, keyIn_0_21 );
nand g057 ( new_n208_, new_n205_, N135 );
nand g058 ( new_n209_, new_n207_, new_n208_ );
xnor g059 ( new_n210_, N91, N96 );
xnor g060 ( new_n211_, N101, N106 );
xnor g061 ( new_n212_, new_n210_, new_n211_ );
xnor g062 ( new_n213_, new_n212_, N130 );
xnor g063 ( N767, new_n209_, new_n213_ );
xnor g064 ( new_n215_, N195, N201 );
nand g065 ( new_n216_, keyIn_0_6, N183 );
xnor g066 ( new_n217_, new_n215_, new_n216_ );
not g067 ( new_n218_, N189 );
nor g068 ( new_n219_, keyIn_0_6, N183 );
nor g069 ( new_n220_, new_n219_, new_n218_ );
xnor g070 ( new_n221_, new_n217_, new_n220_ );
xnor g071 ( new_n222_, new_n221_, N207 );
xnor g072 ( new_n223_, N159, N165 );
xnor g073 ( new_n224_, N171, N177 );
xnor g074 ( new_n225_, new_n223_, new_n224_ );
xnor g075 ( new_n226_, new_n225_, N130 );
xnor g076 ( N768, new_n222_, new_n226_ );
not g077 ( new_n228_, N261 );
not g078 ( new_n229_, N201 );
xnor g079 ( new_n230_, N447, keyIn_0_8 );
nand g080 ( new_n231_, new_n230_, keyIn_0_12 );
not g081 ( new_n232_, keyIn_0_12 );
not g082 ( new_n233_, keyIn_0_8 );
nand g083 ( new_n234_, N447, new_n233_ );
xnor g084 ( new_n235_, new_n188_, keyIn_0_0 );
nand g085 ( new_n236_, new_n235_, keyIn_0_8 );
nand g086 ( new_n237_, new_n236_, new_n234_ );
nand g087 ( new_n238_, new_n237_, new_n232_ );
nand g088 ( new_n239_, new_n231_, new_n238_ );
nand g089 ( new_n240_, N17, N42 );
xnor g090 ( new_n241_, new_n240_, keyIn_0_5 );
nor g091 ( new_n242_, N17, N42 );
xnor g092 ( new_n243_, new_n242_, keyIn_0_4 );
not g093 ( new_n244_, new_n243_ );
nand g094 ( new_n245_, new_n244_, new_n241_ );
nor g095 ( new_n246_, new_n245_, keyIn_0_11 );
nand g096 ( new_n247_, new_n245_, keyIn_0_11 );
nand g097 ( new_n248_, N59, N156 );
not g098 ( new_n249_, new_n248_ );
nand g099 ( new_n250_, new_n247_, new_n249_ );
nor g100 ( new_n251_, new_n250_, new_n246_ );
nand g101 ( new_n252_, new_n239_, new_n251_ );
nand g102 ( new_n253_, new_n252_, keyIn_0_15 );
not g103 ( new_n254_, keyIn_0_15 );
xnor g104 ( new_n255_, new_n237_, keyIn_0_12 );
not g105 ( new_n256_, new_n246_ );
not g106 ( new_n257_, keyIn_0_11 );
not g107 ( new_n258_, new_n241_ );
nor g108 ( new_n259_, new_n258_, new_n243_ );
nor g109 ( new_n260_, new_n259_, new_n257_ );
nor g110 ( new_n261_, new_n260_, new_n248_ );
nand g111 ( new_n262_, new_n261_, new_n256_ );
nor g112 ( new_n263_, new_n255_, new_n262_ );
nand g113 ( new_n264_, new_n263_, new_n254_ );
nand g114 ( new_n265_, new_n264_, new_n253_ );
nand g115 ( new_n266_, N17, N51 );
nor g116 ( new_n267_, new_n163_, new_n266_ );
xor g117 ( new_n268_, new_n267_, keyIn_0_1 );
not g118 ( new_n269_, new_n268_ );
nand g119 ( new_n270_, new_n269_, keyIn_0_9 );
nand g120 ( new_n271_, N42, N59 );
nor g121 ( new_n272_, new_n271_, new_n151_ );
xor g122 ( new_n273_, new_n272_, keyIn_0_2 );
not g123 ( new_n274_, new_n273_ );
nand g124 ( new_n275_, new_n274_, keyIn_0_10 );
nand g125 ( new_n276_, new_n270_, new_n275_ );
not g126 ( new_n277_, keyIn_0_9 );
nand g127 ( new_n278_, new_n268_, new_n277_ );
not g128 ( new_n279_, keyIn_0_10 );
nand g129 ( new_n280_, new_n273_, new_n279_ );
nand g130 ( new_n281_, new_n278_, new_n280_ );
nor g131 ( new_n282_, new_n276_, new_n281_ );
xnor g132 ( new_n283_, new_n282_, keyIn_0_13 );
nand g133 ( new_n284_, new_n265_, new_n283_ );
xnor g134 ( new_n285_, new_n284_, keyIn_0_17 );
nand g135 ( new_n286_, new_n285_, N126 );
not g136 ( new_n287_, keyIn_0_18 );
not g137 ( new_n288_, keyIn_0_16 );
xor g138 ( new_n289_, new_n248_, keyIn_0_3 );
not g139 ( new_n290_, new_n289_ );
nor g140 ( new_n291_, new_n290_, new_n161_ );
nand g141 ( new_n292_, new_n239_, new_n291_ );
nand g142 ( new_n293_, new_n292_, new_n288_ );
not g143 ( new_n294_, new_n293_ );
not g144 ( new_n295_, new_n291_ );
nor g145 ( new_n296_, new_n255_, new_n295_ );
nand g146 ( new_n297_, new_n296_, keyIn_0_16 );
nand g147 ( new_n298_, new_n297_, N1 );
nor g148 ( new_n299_, new_n298_, new_n294_ );
nand g149 ( new_n300_, new_n299_, new_n287_ );
not g150 ( new_n301_, N1 );
nor g151 ( new_n302_, new_n292_, new_n288_ );
nor g152 ( new_n303_, new_n302_, new_n301_ );
nand g153 ( new_n304_, new_n303_, new_n293_ );
nand g154 ( new_n305_, new_n304_, keyIn_0_18 );
nand g155 ( new_n306_, new_n300_, new_n305_ );
nand g156 ( new_n307_, new_n306_, N153 );
nand g157 ( new_n308_, new_n286_, new_n307_ );
xnor g158 ( new_n309_, new_n308_, keyIn_0_27 );
not g159 ( new_n310_, keyIn_0_14 );
nand g160 ( new_n311_, N29, N75 );
nor g161 ( new_n312_, new_n311_, new_n154_ );
nand g162 ( new_n313_, new_n239_, new_n312_ );
nor g163 ( new_n314_, new_n313_, new_n191_ );
nor g164 ( new_n315_, new_n314_, new_n310_ );
not g165 ( new_n316_, N268 );
nand g166 ( new_n317_, new_n314_, new_n310_ );
nand g167 ( new_n318_, new_n317_, new_n316_ );
nor g168 ( new_n319_, new_n318_, new_n315_ );
not g169 ( new_n320_, new_n319_ );
nand g170 ( new_n321_, new_n309_, new_n320_ );
xor g171 ( new_n322_, new_n321_, keyIn_0_30 );
nand g172 ( new_n323_, new_n322_, new_n229_ );
xnor g173 ( new_n324_, new_n323_, keyIn_0_35 );
nor g174 ( new_n325_, new_n322_, new_n229_ );
not g175 ( new_n326_, new_n325_ );
nand g176 ( new_n327_, new_n324_, new_n326_ );
nand g177 ( new_n328_, new_n327_, new_n228_ );
not g178 ( new_n329_, N219 );
nand g179 ( new_n330_, new_n324_, N261 );
nor g180 ( new_n331_, new_n330_, new_n325_ );
nor g181 ( new_n332_, new_n331_, new_n329_ );
nand g182 ( new_n333_, new_n332_, new_n328_ );
not g183 ( new_n334_, N228 );
nor g184 ( new_n335_, new_n327_, new_n334_ );
nand g185 ( new_n336_, new_n325_, N237 );
not g186 ( new_n337_, N246 );
nor g187 ( new_n338_, new_n322_, new_n337_ );
not g188 ( new_n339_, N73 );
nand g189 ( new_n340_, N42, N72 );
nor g190 ( new_n341_, new_n340_, new_n339_ );
nand g191 ( new_n342_, new_n198_, new_n341_ );
not g192 ( new_n343_, new_n342_ );
nand g193 ( new_n344_, new_n343_, N201 );
not g194 ( new_n345_, keyIn_0_7 );
nand g195 ( new_n346_, N121, N210 );
nor g196 ( new_n347_, new_n346_, new_n345_ );
nand g197 ( new_n348_, new_n346_, new_n345_ );
nand g198 ( new_n349_, N255, N267 );
nand g199 ( new_n350_, new_n348_, new_n349_ );
nor g200 ( new_n351_, new_n350_, new_n347_ );
nand g201 ( new_n352_, new_n344_, new_n351_ );
nor g202 ( new_n353_, new_n338_, new_n352_ );
nand g203 ( new_n354_, new_n353_, new_n336_ );
nor g204 ( new_n355_, new_n335_, new_n354_ );
nand g205 ( N850, new_n333_, new_n355_ );
not g206 ( new_n357_, keyIn_0_28 );
not g207 ( new_n358_, keyIn_0_23 );
nand g208 ( new_n359_, new_n285_, N116 );
xnor g209 ( new_n360_, new_n359_, new_n358_ );
not g210 ( new_n361_, keyIn_0_22 );
nand g211 ( new_n362_, new_n306_, N146 );
xnor g212 ( new_n363_, new_n362_, new_n361_ );
nor g213 ( new_n364_, new_n360_, new_n363_ );
nand g214 ( new_n365_, new_n364_, keyIn_0_25 );
not g215 ( new_n366_, keyIn_0_25 );
nand g216 ( new_n367_, new_n359_, keyIn_0_23 );
not g217 ( new_n368_, N116 );
not g218 ( new_n369_, keyIn_0_17 );
xnor g219 ( new_n370_, new_n284_, new_n369_ );
nor g220 ( new_n371_, new_n370_, new_n368_ );
nand g221 ( new_n372_, new_n371_, new_n358_ );
nand g222 ( new_n373_, new_n372_, new_n367_ );
xnor g223 ( new_n374_, new_n362_, keyIn_0_22 );
nand g224 ( new_n375_, new_n373_, new_n374_ );
nand g225 ( new_n376_, new_n375_, new_n366_ );
nand g226 ( new_n377_, new_n365_, new_n376_ );
xor g227 ( new_n378_, new_n319_, keyIn_0_20 );
not g228 ( new_n379_, new_n378_ );
nand g229 ( new_n380_, new_n377_, new_n379_ );
xnor g230 ( new_n381_, new_n380_, new_n357_ );
nand g231 ( new_n382_, new_n381_, N189 );
xnor g232 ( new_n383_, new_n382_, keyIn_0_31 );
xnor g233 ( new_n384_, new_n383_, keyIn_0_36 );
nand g234 ( new_n385_, new_n384_, keyIn_0_39 );
not g235 ( new_n386_, keyIn_0_26 );
not g236 ( new_n387_, keyIn_0_24 );
nand g237 ( new_n388_, new_n285_, N121 );
nor g238 ( new_n389_, new_n388_, new_n387_ );
nand g239 ( new_n390_, new_n388_, new_n387_ );
nand g240 ( new_n391_, new_n306_, N149 );
nand g241 ( new_n392_, new_n390_, new_n391_ );
nor g242 ( new_n393_, new_n392_, new_n389_ );
nand g243 ( new_n394_, new_n393_, new_n386_ );
nor g244 ( new_n395_, new_n393_, new_n386_ );
nor g245 ( new_n396_, new_n395_, new_n319_ );
nand g246 ( new_n397_, new_n396_, new_n394_ );
xnor g247 ( new_n398_, new_n397_, keyIn_0_29 );
nor g248 ( new_n399_, new_n398_, N195 );
xnor g249 ( new_n400_, new_n399_, keyIn_0_34 );
nand g250 ( new_n401_, new_n380_, keyIn_0_28 );
xnor g251 ( new_n402_, new_n375_, keyIn_0_25 );
nor g252 ( new_n403_, new_n402_, new_n378_ );
nand g253 ( new_n404_, new_n403_, new_n357_ );
nand g254 ( new_n405_, new_n404_, new_n401_ );
nand g255 ( new_n406_, new_n405_, new_n218_ );
nand g256 ( new_n407_, new_n406_, keyIn_0_32 );
not g257 ( new_n408_, keyIn_0_32 );
nor g258 ( new_n409_, new_n381_, N189 );
nand g259 ( new_n410_, new_n409_, new_n408_ );
nand g260 ( new_n411_, new_n410_, new_n407_ );
nor g261 ( new_n412_, new_n411_, new_n330_ );
nand g262 ( new_n413_, new_n412_, new_n400_ );
nand g263 ( new_n414_, new_n413_, keyIn_0_38 );
nand g264 ( new_n415_, new_n385_, new_n414_ );
not g265 ( new_n416_, keyIn_0_39 );
not g266 ( new_n417_, keyIn_0_36 );
xnor g267 ( new_n418_, new_n383_, new_n417_ );
nand g268 ( new_n419_, new_n418_, new_n416_ );
not g269 ( new_n420_, keyIn_0_38 );
not g270 ( new_n421_, keyIn_0_34 );
xnor g271 ( new_n422_, new_n399_, new_n421_ );
not g272 ( new_n423_, new_n330_ );
xnor g273 ( new_n424_, new_n406_, new_n408_ );
nand g274 ( new_n425_, new_n423_, new_n424_ );
nor g275 ( new_n426_, new_n425_, new_n422_ );
nand g276 ( new_n427_, new_n426_, new_n420_ );
nand g277 ( new_n428_, new_n419_, new_n427_ );
nor g278 ( new_n429_, new_n415_, new_n428_ );
not g279 ( new_n430_, keyIn_0_40 );
nand g280 ( new_n431_, new_n398_, N195 );
xnor g281 ( new_n432_, new_n431_, keyIn_0_33 );
nand g282 ( new_n433_, new_n432_, keyIn_0_37 );
not g283 ( new_n434_, keyIn_0_37 );
not g284 ( new_n435_, keyIn_0_33 );
nand g285 ( new_n436_, new_n431_, new_n435_ );
not g286 ( new_n437_, N195 );
not g287 ( new_n438_, keyIn_0_29 );
xnor g288 ( new_n439_, new_n397_, new_n438_ );
nor g289 ( new_n440_, new_n439_, new_n437_ );
nand g290 ( new_n441_, new_n440_, keyIn_0_33 );
nand g291 ( new_n442_, new_n441_, new_n436_ );
nand g292 ( new_n443_, new_n442_, new_n434_ );
nand g293 ( new_n444_, new_n433_, new_n443_ );
nand g294 ( new_n445_, new_n444_, new_n424_ );
nor g295 ( new_n446_, new_n445_, new_n430_ );
not g296 ( new_n447_, keyIn_0_41 );
nand g297 ( new_n448_, new_n424_, new_n325_ );
nor g298 ( new_n449_, new_n448_, new_n422_ );
nand g299 ( new_n450_, new_n449_, new_n447_ );
nor g300 ( new_n451_, new_n411_, new_n326_ );
nand g301 ( new_n452_, new_n451_, new_n400_ );
nand g302 ( new_n453_, new_n452_, keyIn_0_41 );
nand g303 ( new_n454_, new_n450_, new_n453_ );
nand g304 ( new_n455_, new_n445_, new_n430_ );
nand g305 ( new_n456_, new_n454_, new_n455_ );
nor g306 ( new_n457_, new_n456_, new_n446_ );
nand g307 ( new_n458_, new_n457_, new_n429_ );
xnor g308 ( new_n459_, new_n458_, keyIn_0_42 );
nand g309 ( new_n460_, new_n285_, N111 );
not g310 ( new_n461_, new_n460_ );
nand g311 ( new_n462_, new_n306_, N143 );
xnor g312 ( new_n463_, new_n319_, keyIn_0_19 );
nand g313 ( new_n464_, new_n463_, new_n462_ );
nor g314 ( new_n465_, new_n464_, new_n461_ );
not g315 ( new_n466_, new_n465_ );
nor g316 ( new_n467_, new_n466_, N183 );
nand g317 ( new_n468_, new_n466_, N183 );
not g318 ( new_n469_, new_n468_ );
nor g319 ( new_n470_, new_n469_, new_n467_ );
nand g320 ( new_n471_, new_n459_, new_n470_ );
nor g321 ( new_n472_, new_n459_, new_n470_ );
nor g322 ( new_n473_, new_n472_, new_n329_ );
nand g323 ( new_n474_, new_n473_, new_n471_ );
not g324 ( new_n475_, new_n470_ );
nor g325 ( new_n476_, new_n475_, new_n334_ );
nand g326 ( new_n477_, new_n469_, N237 );
nor g327 ( new_n478_, new_n465_, new_n337_ );
nand g328 ( new_n479_, new_n343_, N183 );
nand g329 ( new_n480_, N106, N210 );
nand g330 ( new_n481_, new_n479_, new_n480_ );
nor g331 ( new_n482_, new_n478_, new_n481_ );
nand g332 ( new_n483_, new_n477_, new_n482_ );
nor g333 ( new_n484_, new_n476_, new_n483_ );
nand g334 ( N863, new_n474_, new_n484_ );
not g335 ( new_n486_, new_n444_ );
nor g336 ( new_n487_, new_n423_, new_n325_ );
not g337 ( new_n488_, new_n487_ );
nand g338 ( new_n489_, new_n488_, new_n400_ );
nand g339 ( new_n490_, new_n489_, new_n486_ );
nor g340 ( new_n491_, new_n383_, new_n411_ );
nor g341 ( new_n492_, new_n490_, new_n491_ );
nand g342 ( new_n493_, new_n490_, new_n491_ );
nand g343 ( new_n494_, new_n493_, N219 );
nor g344 ( new_n495_, new_n494_, new_n492_ );
nand g345 ( new_n496_, N111, N210 );
not g346 ( new_n497_, new_n496_ );
nor g347 ( new_n498_, new_n495_, new_n497_ );
xnor g348 ( new_n499_, new_n498_, keyIn_0_50 );
not g349 ( new_n500_, N237 );
nor g350 ( new_n501_, new_n418_, new_n500_ );
nand g351 ( new_n502_, new_n491_, N228 );
nor g352 ( new_n503_, new_n405_, new_n337_ );
nand g353 ( new_n504_, new_n343_, N189 );
nand g354 ( new_n505_, N255, N259 );
nand g355 ( new_n506_, new_n504_, new_n505_ );
nor g356 ( new_n507_, new_n503_, new_n506_ );
nand g357 ( new_n508_, new_n502_, new_n507_ );
nor g358 ( new_n509_, new_n501_, new_n508_ );
nand g359 ( N864, new_n499_, new_n509_ );
nor g360 ( new_n511_, new_n422_, new_n432_ );
not g361 ( new_n512_, new_n511_ );
nand g362 ( new_n513_, new_n512_, new_n487_ );
nor g363 ( new_n514_, new_n489_, new_n432_ );
nor g364 ( new_n515_, new_n514_, new_n329_ );
nand g365 ( new_n516_, new_n515_, new_n513_ );
nor g366 ( new_n517_, new_n486_, new_n500_ );
nand g367 ( new_n518_, new_n511_, N228 );
nor g368 ( new_n519_, new_n439_, new_n337_ );
nand g369 ( new_n520_, new_n343_, N195 );
nand g370 ( new_n521_, N255, N260 );
nand g371 ( new_n522_, N116, N210 );
nand g372 ( new_n523_, new_n521_, new_n522_ );
not g373 ( new_n524_, new_n523_ );
nand g374 ( new_n525_, new_n520_, new_n524_ );
nor g375 ( new_n526_, new_n519_, new_n525_ );
nand g376 ( new_n527_, new_n518_, new_n526_ );
nor g377 ( new_n528_, new_n517_, new_n527_ );
nand g378 ( N865, new_n516_, new_n528_ );
not g379 ( new_n530_, keyIn_0_48 );
not g380 ( new_n531_, new_n467_ );
nand g381 ( new_n532_, new_n459_, new_n531_ );
nand g382 ( new_n533_, new_n532_, keyIn_0_43 );
not g383 ( new_n534_, keyIn_0_43 );
not g384 ( new_n535_, keyIn_0_42 );
xnor g385 ( new_n536_, new_n458_, new_n535_ );
nor g386 ( new_n537_, new_n536_, new_n467_ );
nand g387 ( new_n538_, new_n537_, new_n534_ );
nand g388 ( new_n539_, new_n538_, new_n533_ );
nand g389 ( new_n540_, new_n539_, new_n468_ );
xnor g390 ( new_n541_, new_n540_, keyIn_0_44 );
nand g391 ( new_n542_, new_n285_, N96 );
nor g392 ( new_n543_, new_n290_, new_n191_ );
nand g393 ( new_n544_, new_n239_, new_n543_ );
not g394 ( new_n545_, new_n544_ );
nand g395 ( new_n546_, new_n545_, N146 );
not g396 ( new_n547_, new_n546_ );
nor g397 ( new_n548_, new_n161_, N268 );
not g398 ( new_n549_, new_n548_ );
nor g399 ( new_n550_, new_n313_, new_n549_ );
not g400 ( new_n551_, new_n550_ );
nand g401 ( new_n552_, N51, N138 );
nand g402 ( new_n553_, new_n551_, new_n552_ );
nor g403 ( new_n554_, new_n553_, new_n547_ );
nand g404 ( new_n555_, new_n542_, new_n554_ );
nor g405 ( new_n556_, new_n555_, N165 );
nand g406 ( new_n557_, new_n285_, N101 );
nand g407 ( new_n558_, new_n545_, N149 );
not g408 ( new_n559_, new_n558_ );
nand g409 ( new_n560_, N17, N138 );
nand g410 ( new_n561_, new_n551_, new_n560_ );
nor g411 ( new_n562_, new_n561_, new_n559_ );
nand g412 ( new_n563_, new_n557_, new_n562_ );
nor g413 ( new_n564_, new_n563_, N171 );
nor g414 ( new_n565_, new_n556_, new_n564_ );
not g415 ( new_n566_, new_n565_ );
nand g416 ( new_n567_, new_n285_, N106 );
nand g417 ( new_n568_, new_n545_, N153 );
not g418 ( new_n569_, new_n568_ );
nand g419 ( new_n570_, N138, N152 );
nand g420 ( new_n571_, new_n551_, new_n570_ );
nor g421 ( new_n572_, new_n571_, new_n569_ );
nand g422 ( new_n573_, new_n567_, new_n572_ );
nor g423 ( new_n574_, new_n573_, N177 );
nor g424 ( new_n575_, new_n566_, new_n574_ );
nand g425 ( new_n576_, new_n541_, new_n575_ );
nor g426 ( new_n577_, new_n576_, keyIn_0_47 );
not g427 ( new_n578_, new_n577_ );
not g428 ( new_n579_, keyIn_0_47 );
not g429 ( new_n580_, keyIn_0_44 );
xnor g430 ( new_n581_, new_n540_, new_n580_ );
not g431 ( new_n582_, new_n575_ );
nor g432 ( new_n583_, new_n581_, new_n582_ );
nor g433 ( new_n584_, new_n583_, new_n579_ );
nand g434 ( new_n585_, new_n573_, N177 );
nand g435 ( new_n586_, new_n563_, N171 );
nand g436 ( new_n587_, new_n585_, new_n586_ );
nand g437 ( new_n588_, new_n565_, new_n587_ );
nand g438 ( new_n589_, new_n555_, N165 );
nand g439 ( new_n590_, new_n588_, new_n589_ );
nor g440 ( new_n591_, new_n584_, new_n590_ );
nand g441 ( new_n592_, new_n591_, new_n578_ );
nand g442 ( new_n593_, new_n592_, new_n530_ );
nand g443 ( new_n594_, new_n576_, keyIn_0_47 );
not g444 ( new_n595_, new_n590_ );
nand g445 ( new_n596_, new_n594_, new_n595_ );
nor g446 ( new_n597_, new_n596_, new_n577_ );
nand g447 ( new_n598_, new_n597_, keyIn_0_48 );
nand g448 ( new_n599_, new_n593_, new_n598_ );
not g449 ( new_n600_, N159 );
nand g450 ( new_n601_, new_n285_, N91 );
nand g451 ( new_n602_, new_n545_, N143 );
not g452 ( new_n603_, new_n602_ );
nand g453 ( new_n604_, N8, N138 );
nand g454 ( new_n605_, new_n551_, new_n604_ );
nor g455 ( new_n606_, new_n605_, new_n603_ );
nand g456 ( new_n607_, new_n601_, new_n606_ );
not g457 ( new_n608_, new_n607_ );
nand g458 ( new_n609_, new_n608_, new_n600_ );
nand g459 ( new_n610_, new_n599_, new_n609_ );
nand g460 ( new_n611_, new_n607_, N159 );
nand g461 ( N866, new_n610_, new_n611_ );
not g462 ( new_n613_, keyIn_0_55 );
not g463 ( new_n614_, new_n574_ );
nand g464 ( new_n615_, new_n614_, new_n585_ );
not g465 ( new_n616_, new_n615_ );
nand g466 ( new_n617_, new_n541_, new_n616_ );
xnor g467 ( new_n618_, new_n617_, keyIn_0_46 );
nand g468 ( new_n619_, new_n581_, new_n615_ );
xnor g469 ( new_n620_, new_n619_, keyIn_0_45 );
nor g470 ( new_n621_, new_n618_, new_n620_ );
nand g471 ( new_n622_, new_n621_, keyIn_0_49 );
nor g472 ( new_n623_, new_n621_, keyIn_0_49 );
nor g473 ( new_n624_, new_n623_, new_n329_ );
nand g474 ( new_n625_, new_n624_, new_n622_ );
xnor g475 ( new_n626_, new_n625_, keyIn_0_53 );
nand g476 ( new_n627_, N101, N210 );
nand g477 ( new_n628_, new_n626_, new_n627_ );
nand g478 ( new_n629_, new_n628_, new_n613_ );
nor g479 ( new_n630_, new_n628_, new_n613_ );
nand g480 ( new_n631_, new_n616_, N228 );
nor g481 ( new_n632_, new_n585_, new_n500_ );
nand g482 ( new_n633_, new_n573_, N246 );
nand g483 ( new_n634_, new_n343_, N177 );
nand g484 ( new_n635_, new_n633_, new_n634_ );
nor g485 ( new_n636_, new_n632_, new_n635_ );
nand g486 ( new_n637_, new_n631_, new_n636_ );
nor g487 ( new_n638_, new_n630_, new_n637_ );
nand g488 ( new_n639_, new_n638_, new_n629_ );
xor g489 ( new_n640_, new_n639_, keyIn_0_57 );
xnor g490 ( new_n641_, new_n640_, keyIn_0_59 );
xor g491 ( N874, new_n641_, keyIn_0_61 );
not g492 ( new_n643_, keyIn_0_63 );
not g493 ( new_n644_, keyIn_0_58 );
not g494 ( new_n645_, keyIn_0_56 );
not g495 ( new_n646_, keyIn_0_54 );
nand g496 ( new_n647_, new_n609_, new_n611_ );
not g497 ( new_n648_, new_n647_ );
nand g498 ( new_n649_, new_n599_, new_n648_ );
nand g499 ( new_n650_, new_n649_, keyIn_0_52 );
xnor g500 ( new_n651_, new_n597_, new_n530_ );
nand g501 ( new_n652_, new_n651_, new_n647_ );
nand g502 ( new_n653_, new_n652_, keyIn_0_51 );
nand g503 ( new_n654_, new_n653_, new_n650_ );
not g504 ( new_n655_, new_n654_ );
nor g505 ( new_n656_, new_n652_, keyIn_0_51 );
nor g506 ( new_n657_, new_n649_, keyIn_0_52 );
nor g507 ( new_n658_, new_n656_, new_n657_ );
nand g508 ( new_n659_, new_n655_, new_n658_ );
nand g509 ( new_n660_, new_n659_, new_n646_ );
not g510 ( new_n661_, keyIn_0_51 );
nor g511 ( new_n662_, new_n599_, new_n648_ );
nand g512 ( new_n663_, new_n662_, new_n661_ );
not g513 ( new_n664_, keyIn_0_52 );
nor g514 ( new_n665_, new_n651_, new_n647_ );
nand g515 ( new_n666_, new_n665_, new_n664_ );
nand g516 ( new_n667_, new_n666_, new_n663_ );
nor g517 ( new_n668_, new_n667_, new_n654_ );
nand g518 ( new_n669_, new_n668_, keyIn_0_54 );
nand g519 ( new_n670_, new_n660_, new_n669_ );
nand g520 ( new_n671_, new_n670_, N219 );
xnor g521 ( new_n672_, new_n671_, new_n645_ );
nand g522 ( new_n673_, N210, N268 );
not g523 ( new_n674_, new_n673_ );
nor g524 ( new_n675_, new_n672_, new_n674_ );
nor g525 ( new_n676_, new_n675_, new_n644_ );
not g526 ( new_n677_, new_n676_ );
nand g527 ( new_n678_, new_n671_, keyIn_0_56 );
xnor g528 ( new_n679_, new_n668_, new_n646_ );
nor g529 ( new_n680_, new_n679_, new_n329_ );
nand g530 ( new_n681_, new_n680_, new_n645_ );
nand g531 ( new_n682_, new_n681_, new_n678_ );
nand g532 ( new_n683_, new_n682_, new_n673_ );
nor g533 ( new_n684_, new_n683_, keyIn_0_58 );
nor g534 ( new_n685_, new_n647_, new_n334_ );
nor g535 ( new_n686_, new_n611_, new_n500_ );
nand g536 ( new_n687_, new_n607_, N246 );
nand g537 ( new_n688_, new_n343_, N159 );
nand g538 ( new_n689_, new_n687_, new_n688_ );
nor g539 ( new_n690_, new_n686_, new_n689_ );
not g540 ( new_n691_, new_n690_ );
nor g541 ( new_n692_, new_n691_, new_n685_ );
not g542 ( new_n693_, new_n692_ );
nor g543 ( new_n694_, new_n684_, new_n693_ );
nand g544 ( new_n695_, new_n694_, new_n677_ );
nand g545 ( new_n696_, new_n695_, keyIn_0_60 );
not g546 ( new_n697_, keyIn_0_60 );
nand g547 ( new_n698_, new_n675_, new_n644_ );
nand g548 ( new_n699_, new_n698_, new_n692_ );
nor g549 ( new_n700_, new_n699_, new_n676_ );
nand g550 ( new_n701_, new_n700_, new_n697_ );
nand g551 ( new_n702_, new_n701_, new_n696_ );
xnor g552 ( new_n703_, new_n702_, keyIn_0_62 );
nand g553 ( new_n704_, new_n703_, new_n643_ );
not g554 ( new_n705_, keyIn_0_62 );
nand g555 ( new_n706_, new_n702_, new_n705_ );
xnor g556 ( new_n707_, new_n695_, new_n697_ );
nand g557 ( new_n708_, new_n707_, keyIn_0_62 );
nand g558 ( new_n709_, new_n708_, new_n706_ );
nand g559 ( new_n710_, new_n709_, keyIn_0_63 );
nand g560 ( N878, new_n704_, new_n710_ );
not g561 ( new_n712_, new_n564_ );
nand g562 ( new_n713_, new_n541_, new_n614_ );
nand g563 ( new_n714_, new_n713_, new_n585_ );
nand g564 ( new_n715_, new_n714_, new_n712_ );
nand g565 ( new_n716_, new_n715_, new_n586_ );
not g566 ( new_n717_, new_n589_ );
nor g567 ( new_n718_, new_n717_, new_n556_ );
nand g568 ( new_n719_, new_n716_, new_n718_ );
nor g569 ( new_n720_, new_n716_, new_n718_ );
nor g570 ( new_n721_, new_n720_, new_n329_ );
nand g571 ( new_n722_, new_n721_, new_n719_ );
not g572 ( new_n723_, new_n718_ );
nor g573 ( new_n724_, new_n723_, new_n334_ );
nand g574 ( new_n725_, new_n717_, N237 );
nand g575 ( new_n726_, new_n555_, N246 );
not g576 ( new_n727_, N165 );
nor g577 ( new_n728_, new_n342_, new_n727_ );
nand g578 ( new_n729_, N91, N210 );
not g579 ( new_n730_, new_n729_ );
nor g580 ( new_n731_, new_n728_, new_n730_ );
nand g581 ( new_n732_, new_n726_, new_n731_ );
not g582 ( new_n733_, new_n732_ );
nand g583 ( new_n734_, new_n725_, new_n733_ );
nor g584 ( new_n735_, new_n724_, new_n734_ );
nand g585 ( N879, new_n722_, new_n735_ );
not g586 ( new_n737_, new_n586_ );
nor g587 ( new_n738_, new_n737_, new_n564_ );
nand g588 ( new_n739_, new_n714_, new_n738_ );
nor g589 ( new_n740_, new_n714_, new_n738_ );
nor g590 ( new_n741_, new_n740_, new_n329_ );
nand g591 ( new_n742_, new_n741_, new_n739_ );
not g592 ( new_n743_, new_n738_ );
nor g593 ( new_n744_, new_n743_, new_n334_ );
nand g594 ( new_n745_, new_n737_, N237 );
nand g595 ( new_n746_, new_n563_, N246 );
not g596 ( new_n747_, N171 );
nor g597 ( new_n748_, new_n342_, new_n747_ );
nand g598 ( new_n749_, N96, N210 );
not g599 ( new_n750_, new_n749_ );
nor g600 ( new_n751_, new_n748_, new_n750_ );
nand g601 ( new_n752_, new_n746_, new_n751_ );
not g602 ( new_n753_, new_n752_ );
nand g603 ( new_n754_, new_n745_, new_n753_ );
nor g604 ( new_n755_, new_n744_, new_n754_ );
nand g605 ( N880, new_n742_, new_n755_ );
endmodule