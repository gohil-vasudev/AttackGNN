module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n851_, new_n878_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n108_, keyIn_0_10 );
not g001 ( new_n109_, N56 );
and g002 ( new_n110_, keyIn_0_4, N50 );
not g003 ( new_n111_, new_n110_ );
or g004 ( new_n112_, keyIn_0_4, N50 );
and g005 ( new_n113_, new_n111_, new_n112_ );
or g006 ( new_n114_, new_n113_, new_n109_ );
and g007 ( new_n115_, new_n114_, new_n108_ );
not g008 ( new_n116_, new_n115_ );
or g009 ( new_n117_, new_n114_, new_n108_ );
and g010 ( new_n118_, new_n116_, new_n117_ );
not g011 ( new_n119_, keyIn_0_11 );
not g012 ( new_n120_, N82 );
not g013 ( new_n121_, keyIn_0_5 );
or g014 ( new_n122_, new_n121_, N76 );
not g015 ( new_n123_, N76 );
or g016 ( new_n124_, new_n123_, keyIn_0_5 );
and g017 ( new_n125_, new_n122_, new_n124_ );
or g018 ( new_n126_, new_n125_, new_n120_ );
or g019 ( new_n127_, new_n126_, new_n119_ );
and g020 ( new_n128_, new_n123_, keyIn_0_5 );
and g021 ( new_n129_, new_n121_, N76 );
or g022 ( new_n130_, new_n128_, new_n129_ );
and g023 ( new_n131_, new_n130_, N82 );
or g024 ( new_n132_, new_n131_, keyIn_0_11 );
and g025 ( new_n133_, new_n127_, new_n132_ );
or g026 ( new_n134_, keyIn_0_6, N89 );
and g027 ( new_n135_, keyIn_0_6, N89 );
not g028 ( new_n136_, new_n135_ );
and g029 ( new_n137_, new_n136_, N95 );
and g030 ( new_n138_, new_n137_, new_n134_ );
or g031 ( new_n139_, new_n138_, keyIn_0_12 );
not g032 ( new_n140_, keyIn_0_12 );
not g033 ( new_n141_, new_n134_ );
not g034 ( new_n142_, N95 );
or g035 ( new_n143_, new_n135_, new_n142_ );
or g036 ( new_n144_, new_n143_, new_n141_ );
or g037 ( new_n145_, new_n144_, new_n140_ );
and g038 ( new_n146_, new_n139_, new_n145_ );
or g039 ( new_n147_, new_n133_, new_n146_ );
or g040 ( new_n148_, new_n147_, new_n118_ );
not g041 ( new_n149_, N30 );
not g042 ( new_n150_, keyIn_0_1 );
or g043 ( new_n151_, new_n150_, N24 );
not g044 ( new_n152_, N24 );
or g045 ( new_n153_, new_n152_, keyIn_0_1 );
and g046 ( new_n154_, new_n151_, new_n153_ );
or g047 ( new_n155_, new_n154_, new_n149_ );
or g048 ( new_n156_, new_n155_, keyIn_0_8 );
not g049 ( new_n157_, keyIn_0_8 );
and g050 ( new_n158_, new_n152_, keyIn_0_1 );
and g051 ( new_n159_, new_n150_, N24 );
or g052 ( new_n160_, new_n158_, new_n159_ );
and g053 ( new_n161_, new_n160_, N30 );
or g054 ( new_n162_, new_n161_, new_n157_ );
and g055 ( new_n163_, new_n156_, new_n162_ );
not g056 ( new_n164_, N1 );
and g057 ( new_n165_, new_n164_, keyIn_0_0 );
not g058 ( new_n166_, new_n165_ );
or g059 ( new_n167_, new_n164_, keyIn_0_0 );
and g060 ( new_n168_, new_n167_, N4 );
and g061 ( new_n169_, new_n168_, new_n166_ );
not g062 ( new_n170_, N63 );
and g063 ( new_n171_, new_n170_, N69 );
not g064 ( new_n172_, N11 );
and g065 ( new_n173_, new_n172_, N17 );
or g066 ( new_n174_, new_n171_, new_n173_ );
or g067 ( new_n175_, new_n169_, new_n174_ );
or g068 ( new_n176_, new_n163_, new_n175_ );
not g069 ( new_n177_, N102 );
and g070 ( new_n178_, new_n177_, keyIn_0_7 );
not g071 ( new_n179_, N108 );
not g072 ( new_n180_, keyIn_0_7 );
and g073 ( new_n181_, new_n180_, N102 );
or g074 ( new_n182_, new_n181_, new_n179_ );
or g075 ( new_n183_, new_n182_, new_n178_ );
or g076 ( new_n184_, new_n183_, keyIn_0_13 );
not g077 ( new_n185_, keyIn_0_13 );
not g078 ( new_n186_, new_n178_ );
or g079 ( new_n187_, new_n177_, keyIn_0_7 );
and g080 ( new_n188_, new_n187_, N108 );
and g081 ( new_n189_, new_n188_, new_n186_ );
or g082 ( new_n190_, new_n189_, new_n185_ );
and g083 ( new_n191_, new_n184_, new_n190_ );
not g084 ( new_n192_, N43 );
not g085 ( new_n193_, keyIn_0_2 );
or g086 ( new_n194_, new_n193_, N37 );
not g087 ( new_n195_, N37 );
or g088 ( new_n196_, new_n195_, keyIn_0_2 );
and g089 ( new_n197_, new_n194_, new_n196_ );
or g090 ( new_n198_, new_n197_, new_n192_ );
or g091 ( new_n199_, new_n198_, keyIn_0_9 );
not g092 ( new_n200_, keyIn_0_9 );
and g093 ( new_n201_, new_n195_, keyIn_0_2 );
and g094 ( new_n202_, new_n193_, N37 );
or g095 ( new_n203_, new_n201_, new_n202_ );
and g096 ( new_n204_, new_n203_, N43 );
or g097 ( new_n205_, new_n204_, new_n200_ );
and g098 ( new_n206_, new_n199_, new_n205_ );
or g099 ( new_n207_, new_n206_, new_n191_ );
or g100 ( new_n208_, new_n207_, new_n176_ );
or g101 ( new_n209_, new_n208_, new_n148_ );
or g102 ( new_n210_, new_n209_, keyIn_0_14 );
not g103 ( new_n211_, keyIn_0_14 );
not g104 ( new_n212_, new_n118_ );
and g105 ( new_n213_, new_n131_, keyIn_0_11 );
and g106 ( new_n214_, new_n126_, new_n119_ );
or g107 ( new_n215_, new_n214_, new_n213_ );
and g108 ( new_n216_, new_n144_, new_n140_ );
not g109 ( new_n217_, new_n145_ );
or g110 ( new_n218_, new_n217_, new_n216_ );
and g111 ( new_n219_, new_n218_, new_n215_ );
and g112 ( new_n220_, new_n219_, new_n212_ );
and g113 ( new_n221_, new_n161_, new_n157_ );
and g114 ( new_n222_, new_n155_, keyIn_0_8 );
or g115 ( new_n223_, new_n222_, new_n221_ );
not g116 ( new_n224_, new_n175_ );
and g117 ( new_n225_, new_n223_, new_n224_ );
and g118 ( new_n226_, new_n189_, new_n185_ );
and g119 ( new_n227_, new_n183_, keyIn_0_13 );
or g120 ( new_n228_, new_n227_, new_n226_ );
and g121 ( new_n229_, new_n204_, new_n200_ );
and g122 ( new_n230_, new_n198_, keyIn_0_9 );
or g123 ( new_n231_, new_n230_, new_n229_ );
and g124 ( new_n232_, new_n231_, new_n228_ );
and g125 ( new_n233_, new_n225_, new_n232_ );
and g126 ( new_n234_, new_n233_, new_n220_ );
or g127 ( new_n235_, new_n234_, new_n211_ );
and g128 ( N223, new_n210_, new_n235_ );
not g129 ( new_n237_, keyIn_0_28 );
not g130 ( new_n238_, keyIn_0_16 );
not g131 ( new_n239_, new_n169_ );
not g132 ( new_n240_, keyIn_0_15 );
and g133 ( new_n241_, new_n234_, new_n211_ );
and g134 ( new_n242_, new_n209_, keyIn_0_14 );
or g135 ( new_n243_, new_n242_, new_n241_ );
and g136 ( new_n244_, new_n243_, new_n240_ );
and g137 ( new_n245_, N223, keyIn_0_15 );
or g138 ( new_n246_, new_n244_, new_n245_ );
and g139 ( new_n247_, new_n246_, new_n239_ );
or g140 ( new_n248_, N223, keyIn_0_15 );
or g141 ( new_n249_, new_n243_, new_n240_ );
and g142 ( new_n250_, new_n248_, new_n249_ );
and g143 ( new_n251_, new_n250_, new_n169_ );
or g144 ( new_n252_, new_n247_, new_n251_ );
or g145 ( new_n253_, new_n252_, new_n238_ );
or g146 ( new_n254_, new_n250_, new_n169_ );
or g147 ( new_n255_, new_n246_, new_n239_ );
and g148 ( new_n256_, new_n255_, new_n254_ );
or g149 ( new_n257_, new_n256_, keyIn_0_16 );
and g150 ( new_n258_, new_n253_, new_n257_ );
not g151 ( new_n259_, N8 );
and g152 ( new_n260_, new_n259_, N4 );
not g153 ( new_n261_, new_n260_ );
or g154 ( new_n262_, new_n258_, new_n261_ );
and g155 ( new_n263_, new_n262_, keyIn_0_22 );
not g156 ( new_n264_, keyIn_0_22 );
and g157 ( new_n265_, new_n256_, keyIn_0_16 );
and g158 ( new_n266_, new_n252_, new_n238_ );
or g159 ( new_n267_, new_n266_, new_n265_ );
and g160 ( new_n268_, new_n267_, new_n260_ );
and g161 ( new_n269_, new_n268_, new_n264_ );
or g162 ( new_n270_, new_n263_, new_n269_ );
and g163 ( new_n271_, new_n246_, new_n231_ );
and g164 ( new_n272_, new_n250_, new_n206_ );
or g165 ( new_n273_, new_n271_, new_n272_ );
or g166 ( new_n274_, new_n273_, keyIn_0_18 );
not g167 ( new_n275_, keyIn_0_18 );
or g168 ( new_n276_, new_n250_, new_n206_ );
or g169 ( new_n277_, new_n246_, new_n231_ );
and g170 ( new_n278_, new_n277_, new_n276_ );
or g171 ( new_n279_, new_n278_, new_n275_ );
and g172 ( new_n280_, new_n274_, new_n279_ );
not g173 ( new_n281_, N47 );
and g174 ( new_n282_, keyIn_0_3, N43 );
not g175 ( new_n283_, new_n282_ );
or g176 ( new_n284_, keyIn_0_3, N43 );
and g177 ( new_n285_, new_n283_, new_n284_ );
not g178 ( new_n286_, new_n285_ );
and g179 ( new_n287_, new_n286_, new_n281_ );
not g180 ( new_n288_, new_n287_ );
or g181 ( new_n289_, new_n280_, new_n288_ );
and g182 ( new_n290_, new_n289_, keyIn_0_24 );
not g183 ( new_n291_, keyIn_0_24 );
and g184 ( new_n292_, new_n278_, new_n275_ );
and g185 ( new_n293_, new_n273_, keyIn_0_18 );
or g186 ( new_n294_, new_n293_, new_n292_ );
and g187 ( new_n295_, new_n294_, new_n287_ );
and g188 ( new_n296_, new_n295_, new_n291_ );
or g189 ( new_n297_, new_n290_, new_n296_ );
and g190 ( new_n298_, new_n270_, new_n297_ );
and g191 ( new_n299_, new_n246_, new_n228_ );
and g192 ( new_n300_, new_n250_, new_n191_ );
or g193 ( new_n301_, new_n299_, new_n300_ );
and g194 ( new_n302_, new_n301_, keyIn_0_21 );
not g195 ( new_n303_, keyIn_0_21 );
or g196 ( new_n304_, new_n250_, new_n191_ );
or g197 ( new_n305_, new_n246_, new_n228_ );
and g198 ( new_n306_, new_n305_, new_n304_ );
and g199 ( new_n307_, new_n306_, new_n303_ );
or g200 ( new_n308_, new_n302_, new_n307_ );
not g201 ( new_n309_, N112 );
and g202 ( new_n310_, new_n309_, N108 );
not g203 ( new_n311_, new_n310_ );
or g204 ( new_n312_, new_n308_, new_n311_ );
and g205 ( new_n313_, new_n312_, keyIn_0_27 );
not g206 ( new_n314_, keyIn_0_27 );
or g207 ( new_n315_, new_n306_, new_n303_ );
or g208 ( new_n316_, new_n301_, keyIn_0_21 );
and g209 ( new_n317_, new_n316_, new_n315_ );
and g210 ( new_n318_, new_n317_, new_n310_ );
and g211 ( new_n319_, new_n318_, new_n314_ );
or g212 ( new_n320_, new_n313_, new_n319_ );
not g213 ( new_n321_, keyIn_0_25 );
not g214 ( new_n322_, keyIn_0_19 );
and g215 ( new_n323_, new_n246_, new_n212_ );
and g216 ( new_n324_, new_n250_, new_n118_ );
or g217 ( new_n325_, new_n323_, new_n324_ );
or g218 ( new_n326_, new_n325_, new_n322_ );
or g219 ( new_n327_, new_n250_, new_n118_ );
or g220 ( new_n328_, new_n246_, new_n212_ );
and g221 ( new_n329_, new_n328_, new_n327_ );
or g222 ( new_n330_, new_n329_, keyIn_0_19 );
and g223 ( new_n331_, new_n326_, new_n330_ );
not g224 ( new_n332_, N60 );
and g225 ( new_n333_, new_n332_, N56 );
not g226 ( new_n334_, new_n333_ );
or g227 ( new_n335_, new_n331_, new_n334_ );
and g228 ( new_n336_, new_n335_, new_n321_ );
and g229 ( new_n337_, new_n329_, keyIn_0_19 );
and g230 ( new_n338_, new_n325_, new_n322_ );
or g231 ( new_n339_, new_n338_, new_n337_ );
and g232 ( new_n340_, new_n339_, new_n333_ );
and g233 ( new_n341_, new_n340_, keyIn_0_25 );
or g234 ( new_n342_, new_n336_, new_n341_ );
and g235 ( new_n343_, new_n342_, new_n320_ );
and g236 ( new_n344_, new_n298_, new_n343_ );
not g237 ( new_n345_, N17 );
not g238 ( new_n346_, keyIn_0_17 );
not g239 ( new_n347_, new_n173_ );
and g240 ( new_n348_, new_n246_, new_n347_ );
and g241 ( new_n349_, new_n250_, new_n173_ );
or g242 ( new_n350_, new_n348_, new_n349_ );
or g243 ( new_n351_, new_n350_, new_n346_ );
or g244 ( new_n352_, new_n250_, new_n173_ );
or g245 ( new_n353_, new_n246_, new_n347_ );
and g246 ( new_n354_, new_n353_, new_n352_ );
or g247 ( new_n355_, new_n354_, keyIn_0_17 );
and g248 ( new_n356_, new_n351_, new_n355_ );
or g249 ( new_n357_, new_n356_, new_n345_ );
or g250 ( new_n358_, new_n357_, N21 );
and g251 ( new_n359_, new_n358_, keyIn_0_23 );
not g252 ( new_n360_, keyIn_0_23 );
not g253 ( new_n361_, N21 );
and g254 ( new_n362_, new_n354_, keyIn_0_17 );
and g255 ( new_n363_, new_n350_, new_n346_ );
or g256 ( new_n364_, new_n363_, new_n362_ );
and g257 ( new_n365_, new_n364_, N17 );
and g258 ( new_n366_, new_n365_, new_n361_ );
and g259 ( new_n367_, new_n366_, new_n360_ );
or g260 ( new_n368_, new_n359_, new_n367_ );
not g261 ( new_n369_, keyIn_0_20 );
not g262 ( new_n370_, new_n171_ );
and g263 ( new_n371_, new_n246_, new_n370_ );
and g264 ( new_n372_, new_n250_, new_n171_ );
or g265 ( new_n373_, new_n371_, new_n372_ );
or g266 ( new_n374_, new_n373_, new_n369_ );
or g267 ( new_n375_, new_n250_, new_n171_ );
or g268 ( new_n376_, new_n246_, new_n370_ );
and g269 ( new_n377_, new_n376_, new_n375_ );
or g270 ( new_n378_, new_n377_, keyIn_0_20 );
and g271 ( new_n379_, new_n374_, new_n378_ );
not g272 ( new_n380_, N73 );
and g273 ( new_n381_, new_n380_, N69 );
not g274 ( new_n382_, new_n381_ );
or g275 ( new_n383_, new_n379_, new_n382_ );
and g276 ( new_n384_, new_n383_, keyIn_0_26 );
not g277 ( new_n385_, keyIn_0_26 );
and g278 ( new_n386_, new_n377_, keyIn_0_20 );
and g279 ( new_n387_, new_n373_, new_n369_ );
or g280 ( new_n388_, new_n387_, new_n386_ );
and g281 ( new_n389_, new_n388_, new_n381_ );
and g282 ( new_n390_, new_n389_, new_n385_ );
or g283 ( new_n391_, new_n384_, new_n390_ );
not g284 ( new_n392_, N34 );
and g285 ( new_n393_, new_n246_, new_n223_ );
and g286 ( new_n394_, new_n250_, new_n163_ );
or g287 ( new_n395_, new_n393_, new_n394_ );
and g288 ( new_n396_, new_n395_, N30 );
and g289 ( new_n397_, new_n396_, new_n392_ );
not g290 ( new_n398_, new_n397_ );
not g291 ( new_n399_, N99 );
and g292 ( new_n400_, new_n246_, new_n218_ );
and g293 ( new_n401_, new_n250_, new_n146_ );
or g294 ( new_n402_, new_n400_, new_n401_ );
and g295 ( new_n403_, new_n402_, N95 );
and g296 ( new_n404_, new_n403_, new_n399_ );
not g297 ( new_n405_, new_n404_ );
and g298 ( new_n406_, new_n246_, new_n215_ );
and g299 ( new_n407_, new_n250_, new_n133_ );
or g300 ( new_n408_, new_n406_, new_n407_ );
not g301 ( new_n409_, N86 );
and g302 ( new_n410_, new_n409_, N82 );
and g303 ( new_n411_, new_n408_, new_n410_ );
not g304 ( new_n412_, new_n411_ );
and g305 ( new_n413_, new_n405_, new_n412_ );
and g306 ( new_n414_, new_n413_, new_n398_ );
and g307 ( new_n415_, new_n391_, new_n414_ );
and g308 ( new_n416_, new_n368_, new_n415_ );
and g309 ( new_n417_, new_n344_, new_n416_ );
and g310 ( new_n418_, new_n417_, new_n237_ );
not g311 ( new_n419_, new_n418_ );
or g312 ( new_n420_, new_n417_, new_n237_ );
and g313 ( N329, new_n419_, new_n420_ );
not g314 ( new_n422_, keyIn_0_37 );
not g315 ( new_n423_, keyIn_0_31 );
or g316 ( new_n424_, new_n268_, new_n264_ );
or g317 ( new_n425_, new_n262_, keyIn_0_22 );
and g318 ( new_n426_, new_n425_, new_n424_ );
or g319 ( new_n427_, new_n295_, new_n291_ );
or g320 ( new_n428_, new_n289_, keyIn_0_24 );
and g321 ( new_n429_, new_n428_, new_n427_ );
or g322 ( new_n430_, new_n426_, new_n429_ );
or g323 ( new_n431_, new_n318_, new_n314_ );
or g324 ( new_n432_, new_n312_, keyIn_0_27 );
and g325 ( new_n433_, new_n432_, new_n431_ );
or g326 ( new_n434_, new_n340_, keyIn_0_25 );
or g327 ( new_n435_, new_n335_, new_n321_ );
and g328 ( new_n436_, new_n435_, new_n434_ );
or g329 ( new_n437_, new_n433_, new_n436_ );
or g330 ( new_n438_, new_n430_, new_n437_ );
or g331 ( new_n439_, new_n366_, new_n360_ );
or g332 ( new_n440_, new_n358_, keyIn_0_23 );
and g333 ( new_n441_, new_n440_, new_n439_ );
or g334 ( new_n442_, new_n389_, new_n385_ );
or g335 ( new_n443_, new_n383_, keyIn_0_26 );
and g336 ( new_n444_, new_n443_, new_n442_ );
not g337 ( new_n445_, new_n414_ );
or g338 ( new_n446_, new_n444_, new_n445_ );
or g339 ( new_n447_, new_n446_, new_n441_ );
or g340 ( new_n448_, new_n438_, new_n447_ );
and g341 ( new_n449_, new_n448_, keyIn_0_28 );
or g342 ( new_n450_, new_n449_, new_n418_ );
and g343 ( new_n451_, new_n450_, new_n423_ );
and g344 ( new_n452_, N329, keyIn_0_31 );
or g345 ( new_n453_, new_n451_, new_n452_ );
and g346 ( new_n454_, new_n453_, new_n320_ );
or g347 ( new_n455_, N329, keyIn_0_31 );
or g348 ( new_n456_, new_n450_, new_n423_ );
and g349 ( new_n457_, new_n456_, new_n455_ );
and g350 ( new_n458_, new_n457_, new_n433_ );
or g351 ( new_n459_, new_n454_, new_n458_ );
not g352 ( new_n460_, new_n459_ );
and g353 ( new_n461_, new_n460_, new_n422_ );
and g354 ( new_n462_, new_n459_, keyIn_0_37 );
not g355 ( new_n463_, N115 );
and g356 ( new_n464_, new_n463_, N108 );
and g357 ( new_n465_, new_n317_, new_n464_ );
not g358 ( new_n466_, new_n465_ );
and g359 ( new_n467_, new_n466_, keyIn_0_30 );
not g360 ( new_n468_, new_n467_ );
or g361 ( new_n469_, new_n466_, keyIn_0_30 );
and g362 ( new_n470_, new_n468_, new_n469_ );
or g363 ( new_n471_, new_n462_, new_n470_ );
or g364 ( new_n472_, new_n471_, new_n461_ );
and g365 ( new_n473_, new_n472_, keyIn_0_43 );
not g366 ( new_n474_, new_n473_ );
or g367 ( new_n475_, new_n472_, keyIn_0_43 );
and g368 ( new_n476_, new_n474_, new_n475_ );
not g369 ( new_n477_, new_n476_ );
not g370 ( new_n478_, keyIn_0_40 );
not g371 ( new_n479_, keyIn_0_34 );
or g372 ( new_n480_, new_n457_, new_n342_ );
or g373 ( new_n481_, new_n453_, new_n436_ );
and g374 ( new_n482_, new_n481_, new_n480_ );
and g375 ( new_n483_, new_n482_, new_n479_ );
and g376 ( new_n484_, new_n453_, new_n436_ );
and g377 ( new_n485_, new_n457_, new_n342_ );
or g378 ( new_n486_, new_n484_, new_n485_ );
and g379 ( new_n487_, new_n486_, keyIn_0_34 );
not g380 ( new_n488_, N66 );
and g381 ( new_n489_, new_n488_, N56 );
and g382 ( new_n490_, new_n339_, new_n489_ );
not g383 ( new_n491_, new_n490_ );
or g384 ( new_n492_, new_n487_, new_n491_ );
or g385 ( new_n493_, new_n492_, new_n483_ );
and g386 ( new_n494_, new_n493_, new_n478_ );
not g387 ( new_n495_, new_n483_ );
or g388 ( new_n496_, new_n482_, new_n479_ );
and g389 ( new_n497_, new_n496_, new_n490_ );
and g390 ( new_n498_, new_n497_, new_n495_ );
and g391 ( new_n499_, new_n498_, keyIn_0_40 );
or g392 ( new_n500_, new_n494_, new_n499_ );
not g393 ( new_n501_, keyIn_0_41 );
not g394 ( new_n502_, keyIn_0_35 );
or g395 ( new_n503_, new_n457_, new_n391_ );
or g396 ( new_n504_, new_n453_, new_n444_ );
and g397 ( new_n505_, new_n504_, new_n503_ );
and g398 ( new_n506_, new_n505_, new_n502_ );
and g399 ( new_n507_, new_n453_, new_n444_ );
and g400 ( new_n508_, new_n457_, new_n391_ );
or g401 ( new_n509_, new_n507_, new_n508_ );
and g402 ( new_n510_, new_n509_, keyIn_0_35 );
not g403 ( new_n511_, keyIn_0_29 );
not g404 ( new_n512_, N79 );
and g405 ( new_n513_, new_n512_, N69 );
and g406 ( new_n514_, new_n388_, new_n513_ );
not g407 ( new_n515_, new_n514_ );
and g408 ( new_n516_, new_n515_, new_n511_ );
and g409 ( new_n517_, new_n514_, keyIn_0_29 );
or g410 ( new_n518_, new_n516_, new_n517_ );
not g411 ( new_n519_, new_n518_ );
or g412 ( new_n520_, new_n510_, new_n519_ );
or g413 ( new_n521_, new_n520_, new_n506_ );
and g414 ( new_n522_, new_n521_, new_n501_ );
not g415 ( new_n523_, new_n506_ );
or g416 ( new_n524_, new_n505_, new_n502_ );
and g417 ( new_n525_, new_n524_, new_n518_ );
and g418 ( new_n526_, new_n525_, new_n523_ );
and g419 ( new_n527_, new_n526_, keyIn_0_41 );
or g420 ( new_n528_, new_n522_, new_n527_ );
and g421 ( new_n529_, new_n500_, new_n528_ );
and g422 ( new_n530_, new_n529_, new_n477_ );
not g423 ( new_n531_, keyIn_0_36 );
or g424 ( new_n532_, new_n457_, new_n404_ );
or g425 ( new_n533_, new_n453_, new_n405_ );
and g426 ( new_n534_, new_n533_, new_n532_ );
and g427 ( new_n535_, new_n534_, new_n531_ );
and g428 ( new_n536_, new_n453_, new_n405_ );
and g429 ( new_n537_, new_n457_, new_n404_ );
or g430 ( new_n538_, new_n536_, new_n537_ );
and g431 ( new_n539_, new_n538_, keyIn_0_36 );
not g432 ( new_n540_, N105 );
and g433 ( new_n541_, new_n403_, new_n540_ );
not g434 ( new_n542_, new_n541_ );
or g435 ( new_n543_, new_n539_, new_n542_ );
or g436 ( new_n544_, new_n543_, new_n535_ );
and g437 ( new_n545_, new_n544_, keyIn_0_42 );
not g438 ( new_n546_, new_n545_ );
or g439 ( new_n547_, new_n544_, keyIn_0_42 );
or g440 ( new_n548_, new_n457_, new_n397_ );
or g441 ( new_n549_, new_n453_, new_n398_ );
and g442 ( new_n550_, new_n549_, new_n548_ );
and g443 ( new_n551_, new_n550_, keyIn_0_33 );
not g444 ( new_n552_, new_n551_ );
or g445 ( new_n553_, new_n550_, keyIn_0_33 );
not g446 ( new_n554_, N40 );
and g447 ( new_n555_, new_n396_, new_n554_ );
and g448 ( new_n556_, new_n553_, new_n555_ );
and g449 ( new_n557_, new_n556_, new_n552_ );
or g450 ( new_n558_, new_n557_, keyIn_0_39 );
and g451 ( new_n559_, new_n547_, new_n558_ );
and g452 ( new_n560_, new_n559_, new_n546_ );
not g453 ( new_n561_, keyIn_0_38 );
not g454 ( new_n562_, keyIn_0_32 );
or g455 ( new_n563_, new_n457_, new_n368_ );
or g456 ( new_n564_, new_n453_, new_n441_ );
and g457 ( new_n565_, new_n564_, new_n563_ );
and g458 ( new_n566_, new_n565_, new_n562_ );
and g459 ( new_n567_, new_n453_, new_n441_ );
and g460 ( new_n568_, new_n457_, new_n368_ );
or g461 ( new_n569_, new_n567_, new_n568_ );
and g462 ( new_n570_, new_n569_, keyIn_0_32 );
not g463 ( new_n571_, N27 );
and g464 ( new_n572_, new_n365_, new_n571_ );
not g465 ( new_n573_, new_n572_ );
or g466 ( new_n574_, new_n570_, new_n573_ );
or g467 ( new_n575_, new_n574_, new_n566_ );
or g468 ( new_n576_, new_n575_, new_n561_ );
and g469 ( new_n577_, new_n453_, new_n429_ );
and g470 ( new_n578_, new_n457_, new_n297_ );
or g471 ( new_n579_, new_n577_, new_n578_ );
not g472 ( new_n580_, N53 );
and g473 ( new_n581_, new_n286_, new_n580_ );
and g474 ( new_n582_, new_n294_, new_n581_ );
and g475 ( new_n583_, new_n579_, new_n582_ );
or g476 ( new_n584_, new_n453_, new_n412_ );
and g477 ( new_n585_, new_n453_, new_n412_ );
not g478 ( new_n586_, new_n585_ );
not g479 ( new_n587_, N92 );
and g480 ( new_n588_, new_n587_, N82 );
and g481 ( new_n589_, new_n408_, new_n588_ );
and g482 ( new_n590_, new_n586_, new_n589_ );
and g483 ( new_n591_, new_n590_, new_n584_ );
and g484 ( new_n592_, new_n453_, new_n426_ );
and g485 ( new_n593_, new_n457_, new_n270_ );
or g486 ( new_n594_, new_n592_, new_n593_ );
not g487 ( new_n595_, N14 );
and g488 ( new_n596_, new_n595_, N4 );
and g489 ( new_n597_, new_n267_, new_n596_ );
and g490 ( new_n598_, new_n594_, new_n597_ );
or g491 ( new_n599_, new_n591_, new_n598_ );
or g492 ( new_n600_, new_n599_, new_n583_ );
not g493 ( new_n601_, new_n600_ );
and g494 ( new_n602_, new_n576_, new_n601_ );
not g495 ( new_n603_, keyIn_0_39 );
not g496 ( new_n604_, keyIn_0_33 );
and g497 ( new_n605_, new_n453_, new_n398_ );
and g498 ( new_n606_, new_n457_, new_n397_ );
or g499 ( new_n607_, new_n605_, new_n606_ );
and g500 ( new_n608_, new_n607_, new_n604_ );
not g501 ( new_n609_, new_n555_ );
or g502 ( new_n610_, new_n608_, new_n609_ );
or g503 ( new_n611_, new_n610_, new_n551_ );
or g504 ( new_n612_, new_n611_, new_n603_ );
not g505 ( new_n613_, new_n566_ );
or g506 ( new_n614_, new_n565_, new_n562_ );
and g507 ( new_n615_, new_n614_, new_n572_ );
and g508 ( new_n616_, new_n615_, new_n613_ );
or g509 ( new_n617_, new_n616_, keyIn_0_38 );
and g510 ( new_n618_, new_n612_, new_n617_ );
and g511 ( new_n619_, new_n602_, new_n618_ );
and g512 ( new_n620_, new_n619_, new_n560_ );
and g513 ( new_n621_, new_n530_, new_n620_ );
and g514 ( new_n622_, new_n621_, keyIn_0_44 );
not g515 ( new_n623_, new_n622_ );
or g516 ( new_n624_, new_n621_, keyIn_0_44 );
and g517 ( N370, new_n623_, new_n624_ );
not g518 ( new_n626_, keyIn_0_56 );
not g519 ( new_n627_, keyIn_0_51 );
not g520 ( new_n628_, keyIn_0_46 );
not g521 ( new_n629_, keyIn_0_45 );
or g522 ( new_n630_, N370, new_n629_ );
not g523 ( new_n631_, keyIn_0_44 );
or g524 ( new_n632_, new_n498_, keyIn_0_40 );
not g525 ( new_n633_, new_n499_ );
and g526 ( new_n634_, new_n633_, new_n632_ );
or g527 ( new_n635_, new_n526_, keyIn_0_41 );
or g528 ( new_n636_, new_n521_, new_n501_ );
and g529 ( new_n637_, new_n636_, new_n635_ );
or g530 ( new_n638_, new_n634_, new_n637_ );
or g531 ( new_n639_, new_n638_, new_n476_ );
not g532 ( new_n640_, keyIn_0_42 );
not g533 ( new_n641_, new_n535_ );
or g534 ( new_n642_, new_n534_, new_n531_ );
and g535 ( new_n643_, new_n642_, new_n541_ );
and g536 ( new_n644_, new_n643_, new_n641_ );
and g537 ( new_n645_, new_n644_, new_n640_ );
and g538 ( new_n646_, new_n611_, new_n603_ );
or g539 ( new_n647_, new_n646_, new_n645_ );
or g540 ( new_n648_, new_n647_, new_n545_ );
and g541 ( new_n649_, new_n616_, keyIn_0_38 );
or g542 ( new_n650_, new_n649_, new_n600_ );
and g543 ( new_n651_, new_n557_, keyIn_0_39 );
and g544 ( new_n652_, new_n575_, new_n561_ );
or g545 ( new_n653_, new_n652_, new_n651_ );
or g546 ( new_n654_, new_n653_, new_n650_ );
or g547 ( new_n655_, new_n648_, new_n654_ );
or g548 ( new_n656_, new_n639_, new_n655_ );
and g549 ( new_n657_, new_n656_, new_n631_ );
or g550 ( new_n658_, new_n657_, new_n622_ );
or g551 ( new_n659_, new_n658_, keyIn_0_45 );
and g552 ( new_n660_, new_n659_, new_n630_ );
and g553 ( new_n661_, new_n660_, N27 );
and g554 ( new_n662_, new_n661_, new_n628_ );
not g555 ( new_n663_, new_n662_ );
or g556 ( new_n664_, new_n661_, new_n628_ );
and g557 ( new_n665_, new_n663_, new_n664_ );
and g558 ( new_n666_, N329, N21 );
and g559 ( new_n667_, N223, N11 );
or g560 ( new_n668_, new_n667_, new_n345_ );
or g561 ( new_n669_, new_n666_, new_n668_ );
or g562 ( new_n670_, new_n665_, new_n669_ );
and g563 ( new_n671_, new_n670_, new_n627_ );
not g564 ( new_n672_, new_n671_ );
or g565 ( new_n673_, new_n670_, new_n627_ );
and g566 ( new_n674_, new_n672_, new_n673_ );
not g567 ( new_n675_, keyIn_0_47 );
and g568 ( new_n676_, new_n658_, keyIn_0_45 );
and g569 ( new_n677_, N370, new_n629_ );
or g570 ( new_n678_, new_n676_, new_n677_ );
or g571 ( new_n679_, new_n678_, new_n554_ );
and g572 ( new_n680_, new_n679_, new_n675_ );
and g573 ( new_n681_, new_n660_, N40 );
and g574 ( new_n682_, new_n681_, keyIn_0_47 );
or g575 ( new_n683_, new_n680_, new_n682_ );
and g576 ( new_n684_, N329, N34 );
and g577 ( new_n685_, N223, N24 );
or g578 ( new_n686_, new_n685_, new_n149_ );
or g579 ( new_n687_, new_n684_, new_n686_ );
not g580 ( new_n688_, new_n687_ );
and g581 ( new_n689_, new_n683_, new_n688_ );
and g582 ( new_n690_, new_n689_, keyIn_0_52 );
not g583 ( new_n691_, new_n690_ );
or g584 ( new_n692_, new_n689_, keyIn_0_52 );
and g585 ( new_n693_, new_n691_, new_n692_ );
and g586 ( new_n694_, new_n674_, new_n693_ );
or g587 ( new_n695_, new_n678_, new_n580_ );
or g588 ( new_n696_, new_n695_, keyIn_0_48 );
not g589 ( new_n697_, keyIn_0_48 );
and g590 ( new_n698_, new_n660_, N53 );
or g591 ( new_n699_, new_n698_, new_n697_ );
and g592 ( new_n700_, new_n696_, new_n699_ );
and g593 ( new_n701_, N329, N47 );
and g594 ( new_n702_, N223, N37 );
or g595 ( new_n703_, new_n702_, new_n192_ );
or g596 ( new_n704_, new_n701_, new_n703_ );
or g597 ( new_n705_, new_n700_, new_n704_ );
and g598 ( new_n706_, new_n705_, keyIn_0_53 );
not g599 ( new_n707_, keyIn_0_53 );
and g600 ( new_n708_, new_n698_, new_n697_ );
and g601 ( new_n709_, new_n695_, keyIn_0_48 );
or g602 ( new_n710_, new_n709_, new_n708_ );
not g603 ( new_n711_, new_n704_ );
and g604 ( new_n712_, new_n710_, new_n711_ );
and g605 ( new_n713_, new_n712_, new_n707_ );
or g606 ( new_n714_, new_n706_, new_n713_ );
or g607 ( new_n715_, new_n678_, new_n488_ );
or g608 ( new_n716_, new_n715_, keyIn_0_49 );
not g609 ( new_n717_, keyIn_0_49 );
and g610 ( new_n718_, new_n660_, N66 );
or g611 ( new_n719_, new_n718_, new_n717_ );
and g612 ( new_n720_, new_n716_, new_n719_ );
and g613 ( new_n721_, N329, N60 );
and g614 ( new_n722_, N223, N50 );
or g615 ( new_n723_, new_n722_, new_n109_ );
or g616 ( new_n724_, new_n721_, new_n723_ );
or g617 ( new_n725_, new_n720_, new_n724_ );
or g618 ( new_n726_, new_n725_, keyIn_0_54 );
not g619 ( new_n727_, keyIn_0_54 );
and g620 ( new_n728_, new_n718_, new_n717_ );
and g621 ( new_n729_, new_n715_, keyIn_0_49 );
or g622 ( new_n730_, new_n729_, new_n728_ );
not g623 ( new_n731_, new_n724_ );
and g624 ( new_n732_, new_n730_, new_n731_ );
or g625 ( new_n733_, new_n732_, new_n727_ );
and g626 ( new_n734_, new_n726_, new_n733_ );
and g627 ( new_n735_, new_n714_, new_n734_ );
not g628 ( new_n736_, keyIn_0_50 );
or g629 ( new_n737_, new_n678_, new_n512_ );
and g630 ( new_n738_, new_n737_, new_n736_ );
not g631 ( new_n739_, new_n738_ );
or g632 ( new_n740_, new_n737_, new_n736_ );
and g633 ( new_n741_, N329, N73 );
not g634 ( new_n742_, new_n741_ );
and g635 ( new_n743_, N223, N63 );
not g636 ( new_n744_, new_n743_ );
and g637 ( new_n745_, new_n744_, N69 );
and g638 ( new_n746_, new_n742_, new_n745_ );
and g639 ( new_n747_, new_n740_, new_n746_ );
and g640 ( new_n748_, new_n747_, new_n739_ );
or g641 ( new_n749_, new_n748_, keyIn_0_55 );
not g642 ( new_n750_, keyIn_0_55 );
and g643 ( new_n751_, new_n660_, N79 );
and g644 ( new_n752_, new_n751_, keyIn_0_50 );
not g645 ( new_n753_, new_n746_ );
or g646 ( new_n754_, new_n752_, new_n753_ );
or g647 ( new_n755_, new_n754_, new_n738_ );
or g648 ( new_n756_, new_n755_, new_n750_ );
and g649 ( new_n757_, new_n749_, new_n756_ );
and g650 ( new_n758_, new_n660_, N92 );
and g651 ( new_n759_, N329, N86 );
and g652 ( new_n760_, N223, N76 );
or g653 ( new_n761_, new_n760_, new_n120_ );
or g654 ( new_n762_, new_n759_, new_n761_ );
or g655 ( new_n763_, new_n758_, new_n762_ );
and g656 ( new_n764_, new_n660_, N105 );
and g657 ( new_n765_, N329, N99 );
and g658 ( new_n766_, N223, N89 );
or g659 ( new_n767_, new_n766_, new_n142_ );
or g660 ( new_n768_, new_n765_, new_n767_ );
or g661 ( new_n769_, new_n764_, new_n768_ );
and g662 ( new_n770_, new_n660_, N115 );
and g663 ( new_n771_, N329, N112 );
and g664 ( new_n772_, N223, N102 );
or g665 ( new_n773_, new_n772_, new_n179_ );
or g666 ( new_n774_, new_n771_, new_n773_ );
or g667 ( new_n775_, new_n770_, new_n774_ );
and g668 ( new_n776_, new_n769_, new_n775_ );
and g669 ( new_n777_, new_n776_, new_n763_ );
and g670 ( new_n778_, new_n757_, new_n777_ );
and g671 ( new_n779_, new_n735_, new_n778_ );
and g672 ( new_n780_, new_n779_, new_n694_ );
and g673 ( new_n781_, new_n780_, new_n626_ );
not g674 ( new_n782_, new_n781_ );
or g675 ( new_n783_, new_n780_, new_n626_ );
and g676 ( new_n784_, new_n782_, new_n783_ );
and g677 ( new_n785_, new_n660_, N14 );
and g678 ( new_n786_, N329, N8 );
not g679 ( new_n787_, N4 );
and g680 ( new_n788_, N223, N1 );
or g681 ( new_n789_, new_n788_, new_n787_ );
or g682 ( new_n790_, new_n786_, new_n789_ );
or g683 ( new_n791_, new_n785_, new_n790_ );
not g684 ( new_n792_, new_n791_ );
or g685 ( new_n793_, new_n784_, new_n792_ );
and g686 ( new_n794_, new_n793_, keyIn_0_58 );
not g687 ( new_n795_, keyIn_0_58 );
not g688 ( new_n796_, new_n694_ );
or g689 ( new_n797_, new_n712_, new_n707_ );
or g690 ( new_n798_, new_n705_, keyIn_0_53 );
and g691 ( new_n799_, new_n798_, new_n797_ );
and g692 ( new_n800_, new_n732_, new_n727_ );
and g693 ( new_n801_, new_n725_, keyIn_0_54 );
or g694 ( new_n802_, new_n801_, new_n800_ );
or g695 ( new_n803_, new_n802_, new_n799_ );
and g696 ( new_n804_, new_n755_, new_n750_ );
and g697 ( new_n805_, new_n748_, keyIn_0_55 );
or g698 ( new_n806_, new_n805_, new_n804_ );
not g699 ( new_n807_, new_n777_ );
or g700 ( new_n808_, new_n806_, new_n807_ );
or g701 ( new_n809_, new_n803_, new_n808_ );
or g702 ( new_n810_, new_n809_, new_n796_ );
and g703 ( new_n811_, new_n810_, keyIn_0_56 );
or g704 ( new_n812_, new_n811_, new_n781_ );
and g705 ( new_n813_, new_n812_, new_n791_ );
and g706 ( new_n814_, new_n813_, new_n795_ );
or g707 ( N421, new_n794_, new_n814_ );
not g708 ( new_n816_, keyIn_0_61 );
not g709 ( new_n817_, keyIn_0_59 );
not g710 ( new_n818_, keyIn_0_57 );
and g711 ( new_n819_, new_n799_, new_n818_ );
not g712 ( new_n820_, keyIn_0_52 );
or g713 ( new_n821_, new_n681_, keyIn_0_47 );
or g714 ( new_n822_, new_n679_, new_n675_ );
and g715 ( new_n823_, new_n822_, new_n821_ );
or g716 ( new_n824_, new_n823_, new_n687_ );
and g717 ( new_n825_, new_n824_, new_n820_ );
or g718 ( new_n826_, new_n825_, new_n690_ );
and g719 ( new_n827_, new_n714_, keyIn_0_57 );
or g720 ( new_n828_, new_n827_, new_n826_ );
or g721 ( new_n829_, new_n828_, new_n819_ );
or g722 ( new_n830_, new_n829_, new_n817_ );
not g723 ( new_n831_, new_n819_ );
or g724 ( new_n832_, new_n799_, new_n818_ );
and g725 ( new_n833_, new_n832_, new_n693_ );
and g726 ( new_n834_, new_n833_, new_n831_ );
or g727 ( new_n835_, new_n834_, keyIn_0_59 );
and g728 ( new_n836_, new_n830_, new_n835_ );
and g729 ( new_n837_, new_n694_, new_n734_ );
not g730 ( new_n838_, new_n837_ );
or g731 ( new_n839_, new_n836_, new_n838_ );
and g732 ( new_n840_, new_n839_, new_n816_ );
and g733 ( new_n841_, new_n834_, keyIn_0_59 );
and g734 ( new_n842_, new_n829_, new_n817_ );
or g735 ( new_n843_, new_n842_, new_n841_ );
and g736 ( new_n844_, new_n843_, new_n837_ );
and g737 ( new_n845_, new_n844_, keyIn_0_61 );
or g738 ( N430, new_n840_, new_n845_ );
or g739 ( new_n847_, new_n826_, new_n757_ );
or g740 ( new_n848_, new_n803_, new_n847_ );
or g741 ( new_n849_, new_n848_, keyIn_0_60 );
not g742 ( new_n850_, keyIn_0_60 );
and g743 ( new_n851_, new_n693_, new_n806_ );
and g744 ( new_n852_, new_n851_, new_n735_ );
or g745 ( new_n853_, new_n852_, new_n850_ );
and g746 ( new_n854_, new_n849_, new_n853_ );
not g747 ( new_n855_, new_n763_ );
and g748 ( new_n856_, new_n735_, new_n855_ );
or g749 ( new_n857_, new_n796_, new_n856_ );
or g750 ( new_n858_, new_n854_, new_n857_ );
not g751 ( new_n859_, new_n858_ );
and g752 ( new_n860_, new_n859_, keyIn_0_62 );
not g753 ( new_n861_, keyIn_0_62 );
and g754 ( new_n862_, new_n858_, new_n861_ );
or g755 ( N431, new_n860_, new_n862_ );
not g756 ( new_n864_, keyIn_0_63 );
or g757 ( new_n865_, new_n855_, new_n769_ );
or g758 ( new_n866_, new_n799_, new_n865_ );
or g759 ( new_n867_, new_n866_, new_n826_ );
and g760 ( new_n868_, new_n867_, new_n674_ );
not g761 ( new_n869_, new_n868_ );
or g762 ( new_n870_, new_n854_, new_n869_ );
or g763 ( new_n871_, new_n870_, new_n836_ );
and g764 ( new_n872_, new_n871_, new_n864_ );
and g765 ( new_n873_, new_n852_, new_n850_ );
and g766 ( new_n874_, new_n848_, keyIn_0_60 );
or g767 ( new_n875_, new_n874_, new_n873_ );
and g768 ( new_n876_, new_n875_, new_n868_ );
and g769 ( new_n877_, new_n876_, new_n843_ );
and g770 ( new_n878_, new_n877_, keyIn_0_63 );
or g771 ( N432, new_n872_, new_n878_ );
endmodule