module add_mul_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        operation, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218;

  OR2_X1 U113 ( .A1(n105), .A2(n106), .ZN(Result_7_) );
  AND2_X1 U114 ( .A1(operation), .A2(n107), .ZN(n106) );
  AND2_X1 U115 ( .A1(n108), .A2(n109), .ZN(n105) );
  XNOR2_X1 U116 ( .A(n110), .B(a_3_), .ZN(n108) );
  OR2_X1 U117 ( .A1(n111), .A2(n112), .ZN(Result_6_) );
  AND2_X1 U118 ( .A1(n113), .A2(operation), .ZN(n112) );
  XOR2_X1 U119 ( .A(n114), .B(n115), .Z(n113) );
  AND2_X1 U120 ( .A1(b_2_), .A2(a_3_), .ZN(n115) );
  AND2_X1 U121 ( .A1(n116), .A2(n109), .ZN(n111) );
  XOR2_X1 U122 ( .A(n107), .B(n117), .Z(n116) );
  XNOR2_X1 U123 ( .A(n118), .B(a_2_), .ZN(n117) );
  OR2_X1 U124 ( .A1(n119), .A2(n120), .ZN(Result_5_) );
  AND2_X1 U125 ( .A1(n121), .A2(operation), .ZN(n120) );
  XOR2_X1 U126 ( .A(n122), .B(n123), .Z(n121) );
  XNOR2_X1 U127 ( .A(n124), .B(n125), .ZN(n123) );
  AND2_X1 U128 ( .A1(n126), .A2(n109), .ZN(n119) );
  OR3_X1 U129 ( .A1(n127), .A2(n128), .A3(n129), .ZN(n126) );
  AND2_X1 U130 ( .A1(n130), .A2(n131), .ZN(n129) );
  AND2_X1 U131 ( .A1(n132), .A2(n133), .ZN(n128) );
  XNOR2_X1 U132 ( .A(n131), .B(n134), .ZN(n132) );
  INV_X1 U133 ( .A(n135), .ZN(n127) );
  OR3_X1 U134 ( .A1(n131), .A2(a_1_), .A3(n133), .ZN(n135) );
  OR2_X1 U135 ( .A1(n136), .A2(n137), .ZN(Result_4_) );
  AND2_X1 U136 ( .A1(n138), .A2(operation), .ZN(n137) );
  XNOR2_X1 U137 ( .A(n139), .B(n140), .ZN(n138) );
  XOR2_X1 U138 ( .A(n141), .B(n142), .Z(n140) );
  AND2_X1 U139 ( .A1(n143), .A2(n109), .ZN(n136) );
  XOR2_X1 U140 ( .A(n144), .B(n145), .Z(n143) );
  XNOR2_X1 U141 ( .A(n146), .B(a_0_), .ZN(n145) );
  OR2_X1 U142 ( .A1(n147), .A2(n130), .ZN(n144) );
  AND2_X1 U143 ( .A1(n148), .A2(n131), .ZN(n147) );
  OR3_X1 U144 ( .A1(n149), .A2(n150), .A3(n151), .ZN(n131) );
  AND2_X1 U145 ( .A1(n114), .A2(a_3_), .ZN(n151) );
  AND2_X1 U146 ( .A1(b_2_), .A2(n107), .ZN(n150) );
  AND2_X1 U147 ( .A1(a_3_), .A2(b_3_), .ZN(n107) );
  OR2_X1 U148 ( .A1(a_1_), .A2(b_1_), .ZN(n148) );
  AND2_X1 U149 ( .A1(operation), .A2(n152), .ZN(Result_3_) );
  XOR2_X1 U150 ( .A(n153), .B(n154), .Z(n152) );
  AND2_X1 U151 ( .A1(n155), .A2(operation), .ZN(Result_2_) );
  XOR2_X1 U152 ( .A(n156), .B(n157), .Z(n155) );
  AND3_X1 U153 ( .A1(n158), .A2(n159), .A3(operation), .ZN(Result_1_) );
  INV_X1 U154 ( .A(n160), .ZN(n158) );
  AND2_X1 U155 ( .A1(n161), .A2(n162), .ZN(n160) );
  OR2_X1 U156 ( .A1(n157), .A2(n156), .ZN(n161) );
  INV_X1 U157 ( .A(n163), .ZN(Result_0_) );
  OR2_X1 U158 ( .A1(n109), .A2(n164), .ZN(n163) );
  AND3_X1 U159 ( .A1(n165), .A2(n159), .A3(n166), .ZN(n164) );
  OR2_X1 U160 ( .A1(n167), .A2(n168), .ZN(n166) );
  OR3_X1 U161 ( .A1(n157), .A2(n156), .A3(n162), .ZN(n159) );
  OR2_X1 U162 ( .A1(n169), .A2(n170), .ZN(n162) );
  INV_X1 U163 ( .A(n165), .ZN(n170) );
  AND2_X1 U164 ( .A1(n171), .A2(n172), .ZN(n169) );
  OR2_X1 U165 ( .A1(n173), .A2(n174), .ZN(n172) );
  XNOR2_X1 U166 ( .A(n173), .B(n174), .ZN(n156) );
  OR2_X1 U167 ( .A1(n154), .A2(n153), .ZN(n157) );
  OR2_X1 U168 ( .A1(n175), .A2(n176), .ZN(n153) );
  AND2_X1 U169 ( .A1(n142), .A2(n141), .ZN(n176) );
  AND2_X1 U170 ( .A1(n139), .A2(n177), .ZN(n175) );
  OR2_X1 U171 ( .A1(n141), .A2(n142), .ZN(n177) );
  OR2_X1 U172 ( .A1(n110), .A2(n168), .ZN(n142) );
  OR2_X1 U173 ( .A1(n178), .A2(n179), .ZN(n141) );
  AND2_X1 U174 ( .A1(n122), .A2(n125), .ZN(n179) );
  AND2_X1 U175 ( .A1(n180), .A2(n124), .ZN(n178) );
  INV_X1 U176 ( .A(n181), .ZN(n124) );
  AND2_X1 U177 ( .A1(n182), .A2(n183), .ZN(n181) );
  OR2_X1 U178 ( .A1(n184), .A2(n149), .ZN(n182) );
  AND2_X1 U179 ( .A1(a_3_), .A2(b_1_), .ZN(n184) );
  OR2_X1 U180 ( .A1(n125), .A2(n122), .ZN(n180) );
  OR2_X1 U181 ( .A1(n110), .A2(n134), .ZN(n122) );
  INV_X1 U182 ( .A(b_3_), .ZN(n110) );
  INV_X1 U183 ( .A(n185), .ZN(n125) );
  AND3_X1 U184 ( .A1(a_3_), .A2(b_2_), .A3(n114), .ZN(n185) );
  AND2_X1 U185 ( .A1(b_3_), .A2(a_2_), .ZN(n114) );
  XNOR2_X1 U186 ( .A(n186), .B(n187), .ZN(n139) );
  XNOR2_X1 U187 ( .A(n188), .B(n183), .ZN(n186) );
  XNOR2_X1 U188 ( .A(n189), .B(n190), .ZN(n154) );
  XNOR2_X1 U189 ( .A(n191), .B(n192), .ZN(n189) );
  OR3_X1 U190 ( .A1(n171), .A2(n173), .A3(n174), .ZN(n165) );
  OR2_X1 U191 ( .A1(n193), .A2(n194), .ZN(n174) );
  AND2_X1 U192 ( .A1(n192), .A2(n191), .ZN(n194) );
  AND2_X1 U193 ( .A1(n190), .A2(n195), .ZN(n193) );
  OR2_X1 U194 ( .A1(n191), .A2(n192), .ZN(n195) );
  OR2_X1 U195 ( .A1(n196), .A2(n197), .ZN(n192) );
  AND2_X1 U196 ( .A1(n187), .A2(n183), .ZN(n197) );
  AND2_X1 U197 ( .A1(n198), .A2(n188), .ZN(n196) );
  OR2_X1 U198 ( .A1(n199), .A2(n200), .ZN(n188) );
  INV_X1 U199 ( .A(n201), .ZN(n199) );
  OR2_X1 U200 ( .A1(n202), .A2(n203), .ZN(n201) );
  AND2_X1 U201 ( .A1(a_2_), .A2(b_1_), .ZN(n202) );
  OR2_X1 U202 ( .A1(n183), .A2(n187), .ZN(n198) );
  OR2_X1 U203 ( .A1(n118), .A2(n134), .ZN(n187) );
  INV_X1 U204 ( .A(n204), .ZN(n183) );
  AND3_X1 U205 ( .A1(a_3_), .A2(b_1_), .A3(n149), .ZN(n204) );
  AND2_X1 U206 ( .A1(a_2_), .A2(b_2_), .ZN(n149) );
  OR2_X1 U207 ( .A1(n118), .A2(n168), .ZN(n191) );
  INV_X1 U208 ( .A(b_2_), .ZN(n118) );
  XOR2_X1 U209 ( .A(n205), .B(n200), .Z(n190) );
  OR2_X1 U210 ( .A1(n206), .A2(n207), .ZN(n205) );
  INV_X1 U211 ( .A(n208), .ZN(n206) );
  OR2_X1 U212 ( .A1(n130), .A2(n209), .ZN(n208) );
  XOR2_X1 U213 ( .A(n210), .B(n211), .Z(n173) );
  XNOR2_X1 U214 ( .A(n212), .B(n213), .ZN(n210) );
  XNOR2_X1 U215 ( .A(n214), .B(n167), .ZN(n171) );
  OR2_X1 U216 ( .A1(n215), .A2(n216), .ZN(n167) );
  AND2_X1 U217 ( .A1(n211), .A2(n213), .ZN(n216) );
  AND2_X1 U218 ( .A1(n217), .A2(n218), .ZN(n215) );
  OR2_X1 U219 ( .A1(n213), .A2(n211), .ZN(n218) );
  OR2_X1 U220 ( .A1(n134), .A2(n146), .ZN(n211) );
  INV_X1 U221 ( .A(a_1_), .ZN(n134) );
  OR2_X1 U222 ( .A1(n133), .A2(n168), .ZN(n213) );
  INV_X1 U223 ( .A(b_1_), .ZN(n133) );
  INV_X1 U224 ( .A(n212), .ZN(n217) );
  OR2_X1 U225 ( .A1(n207), .A2(n200), .ZN(n212) );
  AND3_X1 U226 ( .A1(a_2_), .A2(b_1_), .A3(n203), .ZN(n200) );
  AND2_X1 U227 ( .A1(a_3_), .A2(b_0_), .ZN(n203) );
  AND2_X1 U228 ( .A1(n130), .A2(n209), .ZN(n207) );
  AND2_X1 U229 ( .A1(a_2_), .A2(b_0_), .ZN(n209) );
  AND2_X1 U230 ( .A1(a_1_), .A2(b_1_), .ZN(n130) );
  OR2_X1 U231 ( .A1(n146), .A2(n168), .ZN(n214) );
  INV_X1 U232 ( .A(a_0_), .ZN(n168) );
  INV_X1 U233 ( .A(b_0_), .ZN(n146) );
  INV_X1 U234 ( .A(operation), .ZN(n109) );
endmodule

