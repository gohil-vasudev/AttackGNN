module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n762_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n583_, new_n239_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n801_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n108_, keyIn_0_8 );
not g001 ( new_n109_, N24 );
and g002 ( new_n110_, new_n108_, new_n109_ );
and g003 ( new_n111_, new_n110_, N30 );
not g004 ( new_n112_, new_n111_ );
and g005 ( new_n113_, new_n109_, N30 );
or g006 ( new_n114_, new_n113_, new_n108_ );
and g007 ( new_n115_, new_n112_, new_n114_ );
not g008 ( new_n116_, N17 );
not g009 ( new_n117_, keyIn_0_7 );
or g010 ( new_n118_, new_n117_, N11 );
or g011 ( new_n119_, new_n118_, new_n116_ );
not g012 ( new_n120_, N11 );
and g013 ( new_n121_, new_n120_, N17 );
or g014 ( new_n122_, new_n121_, keyIn_0_7 );
and g015 ( new_n123_, new_n119_, new_n122_ );
not g016 ( new_n124_, keyIn_0_2 );
not g017 ( new_n125_, N37 );
and g018 ( new_n126_, new_n124_, new_n125_ );
and g019 ( new_n127_, keyIn_0_2, N37 );
or g020 ( new_n128_, new_n126_, new_n127_ );
and g021 ( new_n129_, new_n128_, N43 );
or g022 ( new_n130_, new_n123_, new_n129_ );
or g023 ( new_n131_, new_n130_, new_n115_ );
not g024 ( new_n132_, keyIn_0_10 );
not g025 ( new_n133_, N108 );
or g026 ( new_n134_, new_n133_, N102 );
and g027 ( new_n135_, new_n134_, new_n132_ );
not g028 ( new_n136_, N102 );
and g029 ( new_n137_, new_n136_, keyIn_0_10 );
and g030 ( new_n138_, new_n137_, N108 );
or g031 ( new_n139_, new_n135_, new_n138_ );
not g032 ( new_n140_, N4 );
or g033 ( new_n141_, new_n140_, N1 );
not g034 ( new_n142_, new_n141_ );
not g035 ( new_n143_, N50 );
and g036 ( new_n144_, new_n143_, N56 );
not g037 ( new_n145_, N76 );
and g038 ( new_n146_, new_n145_, N82 );
or g039 ( new_n147_, new_n144_, new_n146_ );
or g040 ( new_n148_, new_n147_, new_n142_ );
or g041 ( new_n149_, new_n148_, new_n139_ );
not g042 ( new_n150_, keyIn_0_9 );
not g043 ( new_n151_, N69 );
or g044 ( new_n152_, new_n151_, N63 );
and g045 ( new_n153_, new_n152_, new_n150_ );
not g046 ( new_n154_, N63 );
and g047 ( new_n155_, new_n154_, keyIn_0_9 );
and g048 ( new_n156_, new_n155_, N69 );
or g049 ( new_n157_, new_n153_, new_n156_ );
or g050 ( new_n158_, keyIn_0_5, N89 );
and g051 ( new_n159_, keyIn_0_5, N89 );
not g052 ( new_n160_, new_n159_ );
and g053 ( new_n161_, new_n160_, N95 );
and g054 ( new_n162_, new_n161_, new_n158_ );
or g055 ( new_n163_, new_n157_, new_n162_ );
or g056 ( new_n164_, new_n149_, new_n163_ );
or g057 ( new_n165_, new_n164_, new_n131_ );
and g058 ( new_n166_, new_n165_, keyIn_0_20 );
not g059 ( new_n167_, keyIn_0_20 );
not g060 ( new_n168_, new_n115_ );
and g061 ( new_n169_, new_n120_, keyIn_0_7 );
and g062 ( new_n170_, new_n169_, N17 );
or g063 ( new_n171_, new_n116_, N11 );
and g064 ( new_n172_, new_n171_, new_n117_ );
or g065 ( new_n173_, new_n172_, new_n170_ );
not g066 ( new_n174_, N43 );
or g067 ( new_n175_, keyIn_0_2, N37 );
not g068 ( new_n176_, new_n127_ );
and g069 ( new_n177_, new_n176_, new_n175_ );
or g070 ( new_n178_, new_n177_, new_n174_ );
and g071 ( new_n179_, new_n173_, new_n178_ );
and g072 ( new_n180_, new_n179_, new_n168_ );
and g073 ( new_n181_, new_n136_, N108 );
or g074 ( new_n182_, new_n181_, keyIn_0_10 );
or g075 ( new_n183_, new_n132_, N102 );
or g076 ( new_n184_, new_n183_, new_n133_ );
and g077 ( new_n185_, new_n184_, new_n182_ );
not g078 ( new_n186_, N56 );
or g079 ( new_n187_, new_n186_, N50 );
not g080 ( new_n188_, N82 );
or g081 ( new_n189_, new_n188_, N76 );
and g082 ( new_n190_, new_n187_, new_n189_ );
and g083 ( new_n191_, new_n190_, new_n141_ );
and g084 ( new_n192_, new_n185_, new_n191_ );
and g085 ( new_n193_, new_n154_, N69 );
or g086 ( new_n194_, new_n193_, keyIn_0_9 );
or g087 ( new_n195_, new_n150_, N63 );
or g088 ( new_n196_, new_n195_, new_n151_ );
and g089 ( new_n197_, new_n196_, new_n194_ );
not g090 ( new_n198_, new_n158_ );
not g091 ( new_n199_, N95 );
or g092 ( new_n200_, new_n159_, new_n199_ );
or g093 ( new_n201_, new_n200_, new_n198_ );
and g094 ( new_n202_, new_n197_, new_n201_ );
and g095 ( new_n203_, new_n192_, new_n202_ );
and g096 ( new_n204_, new_n203_, new_n180_ );
and g097 ( new_n205_, new_n204_, new_n167_ );
or g098 ( N223, new_n166_, new_n205_ );
not g099 ( new_n207_, keyIn_0_38 );
not g100 ( new_n208_, keyIn_0_21 );
and g101 ( new_n209_, new_n165_, keyIn_0_18 );
not g102 ( new_n210_, keyIn_0_18 );
and g103 ( new_n211_, new_n204_, new_n210_ );
or g104 ( new_n212_, new_n209_, new_n211_ );
and g105 ( new_n213_, new_n212_, new_n173_ );
or g106 ( new_n214_, new_n204_, new_n210_ );
not g107 ( new_n215_, new_n211_ );
and g108 ( new_n216_, new_n215_, new_n214_ );
and g109 ( new_n217_, new_n216_, new_n123_ );
or g110 ( new_n218_, new_n213_, new_n217_ );
and g111 ( new_n219_, new_n218_, new_n208_ );
or g112 ( new_n220_, new_n216_, new_n123_ );
or g113 ( new_n221_, new_n212_, new_n173_ );
and g114 ( new_n222_, new_n221_, new_n220_ );
and g115 ( new_n223_, new_n222_, keyIn_0_21 );
or g116 ( new_n224_, new_n219_, new_n223_ );
not g117 ( new_n225_, N21 );
and g118 ( new_n226_, new_n225_, N17 );
not g119 ( new_n227_, new_n226_ );
or g120 ( new_n228_, new_n224_, new_n227_ );
or g121 ( new_n229_, new_n228_, keyIn_0_29 );
not g122 ( new_n230_, keyIn_0_29 );
or g123 ( new_n231_, new_n222_, keyIn_0_21 );
or g124 ( new_n232_, new_n218_, new_n208_ );
and g125 ( new_n233_, new_n232_, new_n231_ );
and g126 ( new_n234_, new_n233_, new_n226_ );
or g127 ( new_n235_, new_n234_, new_n230_ );
and g128 ( new_n236_, new_n229_, new_n235_ );
and g129 ( new_n237_, new_n212_, new_n201_ );
and g130 ( new_n238_, new_n216_, new_n162_ );
or g131 ( new_n239_, new_n237_, new_n238_ );
not g132 ( new_n240_, N99 );
and g133 ( new_n241_, new_n240_, N95 );
and g134 ( new_n242_, new_n239_, new_n241_ );
not g135 ( new_n243_, new_n242_ );
and g136 ( new_n244_, new_n212_, new_n185_ );
and g137 ( new_n245_, new_n139_, new_n210_ );
or g138 ( new_n246_, new_n244_, new_n245_ );
not g139 ( new_n247_, N112 );
and g140 ( new_n248_, new_n247_, N108 );
not g141 ( new_n249_, new_n248_ );
and g142 ( new_n250_, new_n249_, keyIn_0_17 );
not g143 ( new_n251_, new_n250_ );
or g144 ( new_n252_, new_n249_, keyIn_0_17 );
and g145 ( new_n253_, new_n251_, new_n252_ );
and g146 ( new_n254_, new_n246_, new_n253_ );
not g147 ( new_n255_, new_n254_ );
and g148 ( new_n256_, new_n243_, new_n255_ );
not g149 ( new_n257_, new_n256_ );
and g150 ( new_n258_, new_n212_, new_n187_ );
and g151 ( new_n259_, new_n216_, new_n144_ );
or g152 ( new_n260_, new_n258_, new_n259_ );
not g153 ( new_n261_, N60 );
and g154 ( new_n262_, new_n261_, N56 );
and g155 ( new_n263_, new_n262_, keyIn_0_13 );
not g156 ( new_n264_, new_n263_ );
or g157 ( new_n265_, new_n262_, keyIn_0_13 );
and g158 ( new_n266_, new_n264_, new_n265_ );
and g159 ( new_n267_, new_n260_, new_n266_ );
and g160 ( new_n268_, new_n212_, new_n168_ );
and g161 ( new_n269_, new_n115_, new_n210_ );
or g162 ( new_n270_, new_n268_, new_n269_ );
not g163 ( new_n271_, N34 );
not g164 ( new_n272_, N30 );
and g165 ( new_n273_, new_n272_, keyIn_0_1 );
not g166 ( new_n274_, new_n273_ );
or g167 ( new_n275_, new_n272_, keyIn_0_1 );
and g168 ( new_n276_, new_n274_, new_n275_ );
and g169 ( new_n277_, new_n276_, new_n271_ );
and g170 ( new_n278_, new_n270_, new_n277_ );
or g171 ( new_n279_, new_n267_, new_n278_ );
and g172 ( new_n280_, new_n212_, new_n189_ );
and g173 ( new_n281_, new_n216_, new_n146_ );
or g174 ( new_n282_, new_n280_, new_n281_ );
not g175 ( new_n283_, N86 );
and g176 ( new_n284_, new_n283_, N82 );
and g177 ( new_n285_, new_n282_, new_n284_ );
and g178 ( new_n286_, new_n212_, new_n197_ );
and g179 ( new_n287_, new_n216_, new_n157_ );
or g180 ( new_n288_, new_n286_, new_n287_ );
not g181 ( new_n289_, N73 );
and g182 ( new_n290_, keyIn_0_4, N69 );
not g183 ( new_n291_, new_n290_ );
or g184 ( new_n292_, keyIn_0_4, N69 );
and g185 ( new_n293_, new_n291_, new_n292_ );
not g186 ( new_n294_, new_n293_ );
and g187 ( new_n295_, new_n294_, new_n289_ );
and g188 ( new_n296_, new_n288_, new_n295_ );
or g189 ( new_n297_, new_n285_, new_n296_ );
or g190 ( new_n298_, new_n297_, new_n279_ );
or g191 ( new_n299_, new_n298_, new_n257_ );
or g192 ( new_n300_, new_n212_, new_n141_ );
or g193 ( new_n301_, new_n216_, new_n142_ );
and g194 ( new_n302_, new_n300_, new_n301_ );
not g195 ( new_n303_, N8 );
and g196 ( new_n304_, new_n140_, keyIn_0_0 );
not g197 ( new_n305_, new_n304_ );
or g198 ( new_n306_, new_n140_, keyIn_0_0 );
and g199 ( new_n307_, new_n305_, new_n306_ );
not g200 ( new_n308_, new_n307_ );
and g201 ( new_n309_, new_n308_, new_n303_ );
not g202 ( new_n310_, new_n309_ );
and g203 ( new_n311_, new_n310_, keyIn_0_6 );
not g204 ( new_n312_, new_n311_ );
or g205 ( new_n313_, new_n310_, keyIn_0_6 );
and g206 ( new_n314_, new_n312_, new_n313_ );
not g207 ( new_n315_, new_n314_ );
or g208 ( new_n316_, new_n302_, new_n315_ );
and g209 ( new_n317_, new_n316_, keyIn_0_27 );
not g210 ( new_n318_, keyIn_0_27 );
and g211 ( new_n319_, new_n216_, new_n142_ );
and g212 ( new_n320_, new_n212_, new_n141_ );
or g213 ( new_n321_, new_n320_, new_n319_ );
and g214 ( new_n322_, new_n321_, new_n314_ );
and g215 ( new_n323_, new_n322_, new_n318_ );
or g216 ( new_n324_, new_n317_, new_n323_ );
not g217 ( new_n325_, keyIn_0_30 );
or g218 ( new_n326_, new_n212_, new_n178_ );
or g219 ( new_n327_, new_n216_, new_n129_ );
and g220 ( new_n328_, new_n326_, new_n327_ );
not g221 ( new_n329_, N47 );
and g222 ( new_n330_, new_n174_, keyIn_0_3 );
not g223 ( new_n331_, new_n330_ );
or g224 ( new_n332_, new_n174_, keyIn_0_3 );
and g225 ( new_n333_, new_n331_, new_n332_ );
not g226 ( new_n334_, new_n333_ );
and g227 ( new_n335_, new_n334_, new_n329_ );
not g228 ( new_n336_, new_n335_ );
and g229 ( new_n337_, new_n336_, keyIn_0_12 );
not g230 ( new_n338_, new_n337_ );
or g231 ( new_n339_, new_n336_, keyIn_0_12 );
and g232 ( new_n340_, new_n338_, new_n339_ );
not g233 ( new_n341_, new_n340_ );
or g234 ( new_n342_, new_n328_, new_n341_ );
or g235 ( new_n343_, new_n342_, new_n325_ );
and g236 ( new_n344_, new_n216_, new_n129_ );
and g237 ( new_n345_, new_n212_, new_n178_ );
or g238 ( new_n346_, new_n345_, new_n344_ );
and g239 ( new_n347_, new_n346_, new_n340_ );
or g240 ( new_n348_, new_n347_, keyIn_0_30 );
and g241 ( new_n349_, new_n343_, new_n348_ );
or g242 ( new_n350_, new_n324_, new_n349_ );
or g243 ( new_n351_, new_n299_, new_n350_ );
or g244 ( new_n352_, new_n351_, new_n236_ );
and g245 ( new_n353_, new_n352_, keyIn_0_32 );
not g246 ( new_n354_, keyIn_0_32 );
and g247 ( new_n355_, new_n234_, new_n230_ );
and g248 ( new_n356_, new_n228_, keyIn_0_29 );
or g249 ( new_n357_, new_n356_, new_n355_ );
not g250 ( new_n358_, new_n267_ );
not g251 ( new_n359_, new_n278_ );
and g252 ( new_n360_, new_n358_, new_n359_ );
not g253 ( new_n361_, new_n285_ );
not g254 ( new_n362_, new_n296_ );
and g255 ( new_n363_, new_n361_, new_n362_ );
and g256 ( new_n364_, new_n363_, new_n360_ );
and g257 ( new_n365_, new_n364_, new_n256_ );
or g258 ( new_n366_, new_n322_, new_n318_ );
not g259 ( new_n367_, new_n323_ );
and g260 ( new_n368_, new_n367_, new_n366_ );
and g261 ( new_n369_, new_n347_, keyIn_0_30 );
and g262 ( new_n370_, new_n342_, new_n325_ );
or g263 ( new_n371_, new_n370_, new_n369_ );
and g264 ( new_n372_, new_n368_, new_n371_ );
and g265 ( new_n373_, new_n365_, new_n372_ );
and g266 ( new_n374_, new_n373_, new_n357_ );
and g267 ( new_n375_, new_n374_, new_n354_ );
or g268 ( new_n376_, new_n353_, new_n375_ );
and g269 ( new_n377_, new_n376_, new_n207_ );
or g270 ( new_n378_, new_n374_, new_n354_ );
or g271 ( new_n379_, new_n352_, keyIn_0_32 );
and g272 ( new_n380_, new_n379_, new_n378_ );
and g273 ( new_n381_, new_n380_, keyIn_0_38 );
or g274 ( N329, new_n377_, new_n381_ );
not g275 ( new_n383_, keyIn_0_48 );
not g276 ( new_n384_, keyIn_0_46 );
not g277 ( new_n385_, keyIn_0_37 );
and g278 ( new_n386_, new_n376_, new_n385_ );
and g279 ( new_n387_, new_n380_, keyIn_0_37 );
or g280 ( new_n388_, new_n386_, new_n387_ );
and g281 ( new_n389_, new_n388_, new_n296_ );
or g282 ( new_n390_, new_n380_, keyIn_0_37 );
or g283 ( new_n391_, new_n376_, new_n385_ );
and g284 ( new_n392_, new_n390_, new_n391_ );
and g285 ( new_n393_, new_n392_, new_n362_ );
or g286 ( new_n394_, new_n389_, new_n393_ );
and g287 ( new_n395_, new_n394_, keyIn_0_42 );
not g288 ( new_n396_, keyIn_0_42 );
or g289 ( new_n397_, new_n392_, new_n362_ );
or g290 ( new_n398_, new_n388_, new_n296_ );
and g291 ( new_n399_, new_n398_, new_n397_ );
and g292 ( new_n400_, new_n399_, new_n396_ );
or g293 ( new_n401_, new_n395_, new_n400_ );
not g294 ( new_n402_, keyIn_0_35 );
not g295 ( new_n403_, new_n286_ );
not g296 ( new_n404_, new_n287_ );
and g297 ( new_n405_, new_n403_, new_n404_ );
not g298 ( new_n406_, keyIn_0_14 );
not g299 ( new_n407_, N79 );
and g300 ( new_n408_, new_n294_, new_n407_ );
not g301 ( new_n409_, new_n408_ );
and g302 ( new_n410_, new_n409_, new_n406_ );
and g303 ( new_n411_, new_n408_, keyIn_0_14 );
or g304 ( new_n412_, new_n410_, new_n411_ );
or g305 ( new_n413_, new_n405_, new_n412_ );
and g306 ( new_n414_, new_n413_, new_n402_ );
not g307 ( new_n415_, new_n414_ );
or g308 ( new_n416_, new_n413_, new_n402_ );
and g309 ( new_n417_, new_n415_, new_n416_ );
and g310 ( new_n418_, new_n401_, new_n417_ );
and g311 ( new_n419_, new_n418_, new_n384_ );
not g312 ( new_n420_, new_n419_ );
or g313 ( new_n421_, new_n418_, new_n384_ );
not g314 ( new_n422_, keyIn_0_40 );
or g315 ( new_n423_, new_n392_, new_n357_ );
or g316 ( new_n424_, new_n388_, new_n236_ );
and g317 ( new_n425_, new_n424_, new_n423_ );
and g318 ( new_n426_, new_n425_, new_n422_ );
and g319 ( new_n427_, new_n388_, new_n236_ );
and g320 ( new_n428_, new_n392_, new_n357_ );
or g321 ( new_n429_, new_n427_, new_n428_ );
and g322 ( new_n430_, new_n429_, keyIn_0_40 );
not g323 ( new_n431_, keyIn_0_33 );
not g324 ( new_n432_, N27 );
and g325 ( new_n433_, new_n432_, N17 );
and g326 ( new_n434_, new_n233_, new_n433_ );
not g327 ( new_n435_, new_n434_ );
and g328 ( new_n436_, new_n435_, new_n431_ );
and g329 ( new_n437_, new_n434_, keyIn_0_33 );
or g330 ( new_n438_, new_n436_, new_n437_ );
or g331 ( new_n439_, new_n430_, new_n438_ );
or g332 ( new_n440_, new_n439_, new_n426_ );
and g333 ( new_n441_, new_n388_, new_n278_ );
and g334 ( new_n442_, new_n392_, new_n359_ );
or g335 ( new_n443_, new_n441_, new_n442_ );
not g336 ( new_n444_, keyIn_0_34 );
not g337 ( new_n445_, new_n268_ );
not g338 ( new_n446_, new_n269_ );
and g339 ( new_n447_, new_n445_, new_n446_ );
not g340 ( new_n448_, keyIn_0_11 );
not g341 ( new_n449_, N40 );
and g342 ( new_n450_, new_n276_, new_n449_ );
not g343 ( new_n451_, new_n450_ );
and g344 ( new_n452_, new_n451_, new_n448_ );
and g345 ( new_n453_, new_n450_, keyIn_0_11 );
or g346 ( new_n454_, new_n452_, new_n453_ );
or g347 ( new_n455_, new_n447_, new_n454_ );
and g348 ( new_n456_, new_n455_, new_n444_ );
not g349 ( new_n457_, new_n456_ );
or g350 ( new_n458_, new_n455_, new_n444_ );
and g351 ( new_n459_, new_n457_, new_n458_ );
not g352 ( new_n460_, new_n459_ );
and g353 ( new_n461_, new_n443_, new_n460_ );
not g354 ( new_n462_, new_n461_ );
or g355 ( new_n463_, new_n388_, new_n267_ );
or g356 ( new_n464_, new_n392_, new_n358_ );
and g357 ( new_n465_, new_n463_, new_n464_ );
not g358 ( new_n466_, N66 );
and g359 ( new_n467_, new_n466_, N56 );
and g360 ( new_n468_, new_n260_, new_n467_ );
not g361 ( new_n469_, new_n468_ );
or g362 ( new_n470_, new_n465_, new_n469_ );
or g363 ( new_n471_, new_n388_, new_n285_ );
or g364 ( new_n472_, new_n392_, new_n361_ );
and g365 ( new_n473_, new_n471_, new_n472_ );
not g366 ( new_n474_, N92 );
and g367 ( new_n475_, new_n474_, N82 );
and g368 ( new_n476_, new_n475_, keyIn_0_15 );
not g369 ( new_n477_, new_n476_ );
or g370 ( new_n478_, new_n475_, keyIn_0_15 );
and g371 ( new_n479_, new_n477_, new_n478_ );
and g372 ( new_n480_, new_n282_, new_n479_ );
not g373 ( new_n481_, new_n480_ );
and g374 ( new_n482_, new_n481_, keyIn_0_36 );
not g375 ( new_n483_, new_n482_ );
or g376 ( new_n484_, new_n481_, keyIn_0_36 );
and g377 ( new_n485_, new_n483_, new_n484_ );
not g378 ( new_n486_, new_n485_ );
or g379 ( new_n487_, new_n473_, new_n486_ );
and g380 ( new_n488_, new_n470_, new_n487_ );
and g381 ( new_n489_, new_n488_, new_n462_ );
and g382 ( new_n490_, new_n440_, new_n489_ );
and g383 ( new_n491_, new_n421_, new_n490_ );
and g384 ( new_n492_, new_n491_, new_n420_ );
not g385 ( new_n493_, keyIn_0_45 );
and g386 ( new_n494_, new_n388_, new_n349_ );
and g387 ( new_n495_, new_n392_, new_n371_ );
or g388 ( new_n496_, new_n494_, new_n495_ );
or g389 ( new_n497_, new_n496_, keyIn_0_41 );
not g390 ( new_n498_, keyIn_0_41 );
or g391 ( new_n499_, new_n392_, new_n371_ );
or g392 ( new_n500_, new_n388_, new_n349_ );
and g393 ( new_n501_, new_n500_, new_n499_ );
or g394 ( new_n502_, new_n501_, new_n498_ );
and g395 ( new_n503_, new_n497_, new_n502_ );
not g396 ( new_n504_, N53 );
and g397 ( new_n505_, new_n334_, new_n504_ );
and g398 ( new_n506_, new_n346_, new_n505_ );
not g399 ( new_n507_, new_n506_ );
or g400 ( new_n508_, new_n503_, new_n507_ );
and g401 ( new_n509_, new_n508_, new_n493_ );
and g402 ( new_n510_, new_n501_, new_n498_ );
and g403 ( new_n511_, new_n496_, keyIn_0_41 );
or g404 ( new_n512_, new_n511_, new_n510_ );
and g405 ( new_n513_, new_n512_, new_n506_ );
and g406 ( new_n514_, new_n513_, keyIn_0_45 );
or g407 ( new_n515_, new_n509_, new_n514_ );
not g408 ( new_n516_, keyIn_0_47 );
and g409 ( new_n517_, new_n392_, new_n243_ );
and g410 ( new_n518_, new_n388_, new_n242_ );
or g411 ( new_n519_, new_n518_, new_n517_ );
not g412 ( new_n520_, new_n239_ );
not g413 ( new_n521_, keyIn_0_16 );
not g414 ( new_n522_, N105 );
and g415 ( new_n523_, new_n522_, N95 );
not g416 ( new_n524_, new_n523_ );
and g417 ( new_n525_, new_n524_, new_n521_ );
and g418 ( new_n526_, new_n523_, keyIn_0_16 );
or g419 ( new_n527_, new_n525_, new_n526_ );
or g420 ( new_n528_, new_n520_, new_n527_ );
not g421 ( new_n529_, new_n528_ );
and g422 ( new_n530_, new_n519_, new_n529_ );
not g423 ( new_n531_, new_n530_ );
and g424 ( new_n532_, new_n531_, new_n516_ );
and g425 ( new_n533_, new_n530_, keyIn_0_47 );
or g426 ( new_n534_, new_n532_, new_n533_ );
or g427 ( new_n535_, new_n392_, new_n255_ );
or g428 ( new_n536_, new_n388_, new_n254_ );
and g429 ( new_n537_, new_n536_, new_n535_ );
and g430 ( new_n538_, new_n537_, keyIn_0_43 );
not g431 ( new_n539_, keyIn_0_43 );
and g432 ( new_n540_, new_n388_, new_n254_ );
and g433 ( new_n541_, new_n392_, new_n255_ );
or g434 ( new_n542_, new_n540_, new_n541_ );
and g435 ( new_n543_, new_n542_, new_n539_ );
not g436 ( new_n544_, keyIn_0_31 );
not g437 ( new_n545_, N115 );
and g438 ( new_n546_, new_n545_, N108 );
and g439 ( new_n547_, new_n246_, new_n546_ );
not g440 ( new_n548_, new_n547_ );
and g441 ( new_n549_, new_n548_, new_n544_ );
and g442 ( new_n550_, new_n547_, keyIn_0_31 );
or g443 ( new_n551_, new_n549_, new_n550_ );
not g444 ( new_n552_, new_n551_ );
or g445 ( new_n553_, new_n543_, new_n552_ );
or g446 ( new_n554_, new_n553_, new_n538_ );
or g447 ( new_n555_, new_n392_, new_n368_ );
or g448 ( new_n556_, new_n388_, new_n324_ );
and g449 ( new_n557_, new_n556_, new_n555_ );
and g450 ( new_n558_, new_n557_, keyIn_0_39 );
not g451 ( new_n559_, keyIn_0_39 );
and g452 ( new_n560_, new_n388_, new_n324_ );
and g453 ( new_n561_, new_n392_, new_n368_ );
or g454 ( new_n562_, new_n560_, new_n561_ );
and g455 ( new_n563_, new_n562_, new_n559_ );
not g456 ( new_n564_, keyIn_0_28 );
not g457 ( new_n565_, N14 );
and g458 ( new_n566_, new_n308_, new_n565_ );
and g459 ( new_n567_, new_n321_, new_n566_ );
not g460 ( new_n568_, new_n567_ );
and g461 ( new_n569_, new_n568_, new_n564_ );
and g462 ( new_n570_, new_n567_, keyIn_0_28 );
or g463 ( new_n571_, new_n569_, new_n570_ );
not g464 ( new_n572_, new_n571_ );
or g465 ( new_n573_, new_n563_, new_n572_ );
or g466 ( new_n574_, new_n573_, new_n558_ );
and g467 ( new_n575_, new_n554_, new_n574_ );
and g468 ( new_n576_, new_n575_, new_n534_ );
and g469 ( new_n577_, new_n515_, new_n576_ );
and g470 ( new_n578_, new_n577_, new_n492_ );
not g471 ( new_n579_, new_n578_ );
and g472 ( new_n580_, new_n579_, new_n383_ );
and g473 ( new_n581_, new_n578_, keyIn_0_48 );
or g474 ( N370, new_n580_, new_n581_ );
not g475 ( new_n583_, keyIn_0_49 );
or g476 ( new_n584_, new_n578_, keyIn_0_48 );
not g477 ( new_n585_, new_n581_ );
and g478 ( new_n586_, new_n585_, new_n584_ );
and g479 ( new_n587_, new_n586_, new_n583_ );
not g480 ( new_n588_, new_n587_ );
or g481 ( new_n589_, new_n586_, new_n583_ );
and g482 ( new_n590_, new_n589_, N105 );
and g483 ( new_n591_, new_n590_, new_n588_ );
and g484 ( new_n592_, new_n591_, keyIn_0_52 );
not g485 ( new_n593_, new_n592_ );
or g486 ( new_n594_, new_n591_, keyIn_0_52 );
and g487 ( new_n595_, new_n593_, new_n594_ );
and g488 ( new_n596_, new_n376_, N99 );
and g489 ( new_n597_, new_n165_, keyIn_0_19 );
not g490 ( new_n598_, keyIn_0_19 );
and g491 ( new_n599_, new_n204_, new_n598_ );
or g492 ( new_n600_, new_n597_, new_n599_ );
not g493 ( new_n601_, new_n600_ );
and g494 ( new_n602_, new_n601_, N89 );
or g495 ( new_n603_, new_n602_, new_n199_ );
or g496 ( new_n604_, new_n596_, new_n603_ );
or g497 ( new_n605_, new_n595_, new_n604_ );
and g498 ( new_n606_, new_n605_, keyIn_0_55 );
not g499 ( new_n607_, new_n606_ );
or g500 ( new_n608_, new_n605_, keyIn_0_55 );
and g501 ( new_n609_, new_n607_, new_n608_ );
not g502 ( new_n610_, keyIn_0_50 );
and g503 ( new_n611_, new_n589_, N66 );
and g504 ( new_n612_, new_n611_, new_n588_ );
and g505 ( new_n613_, new_n612_, new_n610_ );
and g506 ( new_n614_, N370, keyIn_0_49 );
or g507 ( new_n615_, new_n614_, new_n466_ );
or g508 ( new_n616_, new_n615_, new_n587_ );
and g509 ( new_n617_, new_n616_, keyIn_0_50 );
and g510 ( new_n618_, new_n376_, N60 );
not g511 ( new_n619_, new_n618_ );
not g512 ( new_n620_, keyIn_0_24 );
and g513 ( new_n621_, new_n601_, N50 );
and g514 ( new_n622_, new_n621_, new_n620_ );
not g515 ( new_n623_, new_n622_ );
or g516 ( new_n624_, new_n621_, new_n620_ );
and g517 ( new_n625_, new_n624_, N56 );
and g518 ( new_n626_, new_n625_, new_n623_ );
and g519 ( new_n627_, new_n619_, new_n626_ );
not g520 ( new_n628_, new_n627_ );
or g521 ( new_n629_, new_n617_, new_n628_ );
or g522 ( new_n630_, new_n629_, new_n613_ );
or g523 ( new_n631_, new_n614_, new_n504_ );
or g524 ( new_n632_, new_n631_, new_n587_ );
and g525 ( new_n633_, new_n376_, N47 );
and g526 ( new_n634_, new_n601_, N37 );
not g527 ( new_n635_, new_n634_ );
and g528 ( new_n636_, new_n635_, keyIn_0_23 );
not g529 ( new_n637_, new_n636_ );
or g530 ( new_n638_, new_n635_, keyIn_0_23 );
and g531 ( new_n639_, new_n637_, new_n638_ );
or g532 ( new_n640_, new_n639_, new_n174_ );
or g533 ( new_n641_, new_n633_, new_n640_ );
not g534 ( new_n642_, new_n641_ );
and g535 ( new_n643_, new_n632_, new_n642_ );
not g536 ( new_n644_, new_n643_ );
and g537 ( new_n645_, new_n630_, new_n644_ );
not g538 ( new_n646_, keyIn_0_56 );
and g539 ( new_n647_, new_n589_, N115 );
and g540 ( new_n648_, new_n647_, new_n588_ );
not g541 ( new_n649_, new_n648_ );
not g542 ( new_n650_, keyIn_0_44 );
and g543 ( new_n651_, new_n376_, N112 );
not g544 ( new_n652_, new_n651_ );
and g545 ( new_n653_, new_n652_, new_n650_ );
and g546 ( new_n654_, new_n651_, keyIn_0_44 );
or g547 ( new_n655_, new_n653_, new_n654_ );
and g548 ( new_n656_, new_n601_, N102 );
or g549 ( new_n657_, new_n656_, new_n133_ );
not g550 ( new_n658_, new_n657_ );
and g551 ( new_n659_, new_n655_, new_n658_ );
and g552 ( new_n660_, new_n649_, new_n659_ );
and g553 ( new_n661_, new_n660_, new_n646_ );
not g554 ( new_n662_, new_n661_ );
or g555 ( new_n663_, new_n660_, new_n646_ );
and g556 ( new_n664_, new_n662_, new_n663_ );
or g557 ( new_n665_, new_n614_, new_n432_ );
or g558 ( new_n666_, new_n665_, new_n587_ );
and g559 ( new_n667_, new_n376_, N21 );
not g560 ( new_n668_, new_n667_ );
not g561 ( new_n669_, keyIn_0_22 );
and g562 ( new_n670_, new_n601_, N11 );
and g563 ( new_n671_, new_n670_, new_n669_ );
not g564 ( new_n672_, new_n671_ );
or g565 ( new_n673_, new_n670_, new_n669_ );
and g566 ( new_n674_, new_n673_, N17 );
and g567 ( new_n675_, new_n674_, new_n672_ );
and g568 ( new_n676_, new_n668_, new_n675_ );
and g569 ( new_n677_, new_n666_, new_n676_ );
or g570 ( new_n678_, new_n614_, new_n449_ );
or g571 ( new_n679_, new_n678_, new_n587_ );
and g572 ( new_n680_, new_n376_, N34 );
and g573 ( new_n681_, new_n601_, N24 );
or g574 ( new_n682_, new_n681_, new_n272_ );
or g575 ( new_n683_, new_n680_, new_n682_ );
not g576 ( new_n684_, new_n683_ );
and g577 ( new_n685_, new_n679_, new_n684_ );
or g578 ( new_n686_, new_n677_, new_n685_ );
or g579 ( new_n687_, new_n664_, new_n686_ );
not g580 ( new_n688_, keyIn_0_54 );
or g581 ( new_n689_, new_n614_, new_n474_ );
or g582 ( new_n690_, new_n689_, new_n587_ );
and g583 ( new_n691_, new_n376_, N86 );
not g584 ( new_n692_, new_n691_ );
not g585 ( new_n693_, keyIn_0_26 );
and g586 ( new_n694_, new_n601_, N76 );
not g587 ( new_n695_, new_n694_ );
and g588 ( new_n696_, new_n695_, new_n693_ );
and g589 ( new_n697_, new_n694_, keyIn_0_26 );
or g590 ( new_n698_, new_n696_, new_n697_ );
and g591 ( new_n699_, new_n698_, N82 );
and g592 ( new_n700_, new_n692_, new_n699_ );
and g593 ( new_n701_, new_n690_, new_n700_ );
or g594 ( new_n702_, new_n701_, new_n688_ );
and g595 ( new_n703_, new_n589_, N92 );
and g596 ( new_n704_, new_n703_, new_n588_ );
not g597 ( new_n705_, new_n700_ );
or g598 ( new_n706_, new_n704_, new_n705_ );
or g599 ( new_n707_, new_n706_, keyIn_0_54 );
and g600 ( new_n708_, new_n702_, new_n707_ );
and g601 ( new_n709_, new_n589_, N79 );
and g602 ( new_n710_, new_n709_, new_n588_ );
not g603 ( new_n711_, new_n710_ );
and g604 ( new_n712_, new_n711_, keyIn_0_51 );
not g605 ( new_n713_, keyIn_0_51 );
and g606 ( new_n714_, new_n710_, new_n713_ );
or g607 ( new_n715_, new_n712_, new_n714_ );
and g608 ( new_n716_, new_n376_, N73 );
not g609 ( new_n717_, new_n716_ );
not g610 ( new_n718_, keyIn_0_25 );
and g611 ( new_n719_, new_n601_, N63 );
not g612 ( new_n720_, new_n719_ );
and g613 ( new_n721_, new_n720_, new_n718_ );
and g614 ( new_n722_, new_n719_, keyIn_0_25 );
or g615 ( new_n723_, new_n721_, new_n722_ );
and g616 ( new_n724_, new_n723_, N69 );
and g617 ( new_n725_, new_n717_, new_n724_ );
and g618 ( new_n726_, new_n715_, new_n725_ );
or g619 ( new_n727_, new_n726_, new_n708_ );
or g620 ( new_n728_, new_n687_, new_n727_ );
not g621 ( new_n729_, new_n728_ );
and g622 ( new_n730_, new_n729_, new_n645_ );
and g623 ( new_n731_, new_n730_, new_n609_ );
and g624 ( new_n732_, new_n731_, keyIn_0_58 );
not g625 ( new_n733_, keyIn_0_58 );
not g626 ( new_n734_, new_n609_ );
not g627 ( new_n735_, new_n613_ );
or g628 ( new_n736_, new_n612_, new_n610_ );
and g629 ( new_n737_, new_n736_, new_n627_ );
and g630 ( new_n738_, new_n737_, new_n735_ );
or g631 ( new_n739_, new_n738_, new_n643_ );
or g632 ( new_n740_, new_n728_, new_n739_ );
or g633 ( new_n741_, new_n740_, new_n734_ );
and g634 ( new_n742_, new_n741_, new_n733_ );
or g635 ( new_n743_, new_n732_, new_n742_ );
not g636 ( new_n744_, keyIn_0_53 );
and g637 ( new_n745_, new_n589_, N14 );
and g638 ( new_n746_, new_n745_, new_n588_ );
and g639 ( new_n747_, new_n376_, N8 );
and g640 ( new_n748_, new_n601_, N1 );
or g641 ( new_n749_, new_n748_, new_n140_ );
or g642 ( new_n750_, new_n747_, new_n749_ );
or g643 ( new_n751_, new_n746_, new_n750_ );
and g644 ( new_n752_, new_n751_, new_n744_ );
not g645 ( new_n753_, new_n752_ );
or g646 ( new_n754_, new_n751_, new_n744_ );
and g647 ( new_n755_, new_n753_, new_n754_ );
not g648 ( new_n756_, new_n755_ );
or g649 ( new_n757_, new_n756_, keyIn_0_57 );
not g650 ( new_n758_, keyIn_0_57 );
or g651 ( new_n759_, new_n755_, new_n758_ );
and g652 ( new_n760_, new_n757_, new_n759_ );
and g653 ( N421, new_n743_, new_n760_ );
not g654 ( new_n762_, keyIn_0_62 );
not g655 ( new_n763_, new_n685_ );
and g656 ( new_n764_, new_n763_, new_n643_ );
not g657 ( new_n765_, new_n764_ );
and g658 ( new_n766_, new_n765_, keyIn_0_60 );
not g659 ( new_n767_, new_n766_ );
or g660 ( new_n768_, new_n765_, keyIn_0_60 );
and g661 ( new_n769_, new_n767_, new_n768_ );
not g662 ( new_n770_, new_n769_ );
not g663 ( new_n771_, new_n686_ );
and g664 ( new_n772_, new_n630_, new_n771_ );
and g665 ( new_n773_, new_n770_, new_n772_ );
not g666 ( new_n774_, new_n773_ );
or g667 ( new_n775_, new_n774_, new_n762_ );
or g668 ( new_n776_, new_n773_, keyIn_0_62 );
and g669 ( N430, new_n775_, new_n776_ );
not g670 ( new_n778_, keyIn_0_59 );
and g671 ( new_n779_, new_n708_, new_n778_ );
not g672 ( new_n780_, new_n779_ );
or g673 ( new_n781_, new_n708_, new_n778_ );
and g674 ( new_n782_, new_n781_, new_n645_ );
and g675 ( new_n783_, new_n782_, new_n780_ );
and g676 ( new_n784_, new_n783_, keyIn_0_61 );
not g677 ( new_n785_, keyIn_0_61 );
and g678 ( new_n786_, new_n706_, keyIn_0_54 );
and g679 ( new_n787_, new_n701_, new_n688_ );
or g680 ( new_n788_, new_n787_, new_n786_ );
and g681 ( new_n789_, new_n788_, keyIn_0_59 );
or g682 ( new_n790_, new_n789_, new_n739_ );
or g683 ( new_n791_, new_n790_, new_n779_ );
and g684 ( new_n792_, new_n791_, new_n785_ );
and g685 ( new_n793_, new_n726_, new_n763_ );
and g686 ( new_n794_, new_n793_, new_n645_ );
or g687 ( new_n795_, new_n794_, new_n686_ );
or g688 ( new_n796_, new_n792_, new_n795_ );
or g689 ( new_n797_, new_n796_, new_n784_ );
or g690 ( new_n798_, new_n797_, keyIn_0_63 );
not g691 ( new_n799_, keyIn_0_63 );
not g692 ( new_n800_, new_n784_ );
or g693 ( new_n801_, new_n783_, keyIn_0_61 );
not g694 ( new_n802_, new_n795_ );
and g695 ( new_n803_, new_n801_, new_n802_ );
and g696 ( new_n804_, new_n803_, new_n800_ );
or g697 ( new_n805_, new_n804_, new_n799_ );
and g698 ( N431, new_n798_, new_n805_ );
and g699 ( new_n807_, new_n644_, new_n763_ );
and g700 ( new_n808_, new_n788_, new_n807_ );
and g701 ( new_n809_, new_n734_, new_n808_ );
or g702 ( new_n810_, new_n769_, new_n677_ );
or g703 ( new_n811_, new_n810_, new_n794_ );
or g704 ( N432, new_n811_, new_n809_ );
endmodule