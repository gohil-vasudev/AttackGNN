module add_mul_mix_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_, 
        c_9_, c_10_, c_11_, c_12_, c_13_, c_14_, c_15_, d_0_, d_1_, d_2_, d_3_, 
        d_4_, d_5_, d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, 
        d_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_, c_9_, c_10_,
         c_11_, c_12_, c_13_, c_14_, c_15_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_,
         d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, d_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001;

  XOR2_X2 U1948 ( .A(n3274), .B(n3275), .Z(n3015) );
  XOR2_X2 U1949 ( .A(n3903), .B(n3904), .Z(n2117) );
  XOR2_X2 U1950 ( .A(n3905), .B(n3906), .Z(n2459) );
  XNOR2_X2 U1951 ( .A(n2525), .B(n2526), .ZN(n2229) );
  XOR2_X2 U1952 ( .A(n3396), .B(n3397), .Z(n3140) );
  XOR2_X2 U1953 ( .A(n3797), .B(n3798), .Z(n3523) );
  XOR2_X2 U1954 ( .A(n3144), .B(n3145), .Z(n2893) );
  XNOR2_X2 U1955 ( .A(n2213), .B(n2307), .ZN(n1955) );
  XOR2_X2 U1956 ( .A(n2413), .B(n2414), .Z(n2200) );
  INV_X1 U1957 ( .A(n3269), .ZN(n1916) );
  XOR2_X2 U1958 ( .A(n3891), .B(n3892), .Z(n2165) );
  XOR2_X2 U1959 ( .A(n3895), .B(n3896), .Z(n2149) );
  XNOR2_X2 U1960 ( .A(n3887), .B(n3888), .ZN(n2182) );
  XOR2_X2 U1961 ( .A(n3899), .B(n3900), .Z(n2133) );
  XOR2_X2 U1962 ( .A(n3907), .B(n3908), .Z(n2026) );
  INV_X1 U1963 ( .A(n2362), .ZN(n1917) );
  XOR2_X2 U1964 ( .A(n3957), .B(n3958), .Z(n3711) );
  XOR2_X2 U1965 ( .A(n3913), .B(n3916), .Z(n2095) );
  INV_X1 U1966 ( .A(n3391), .ZN(n1918) );
  XOR2_X1 U1967 ( .A(n1919), .B(n1920), .Z(Result_9_) );
  AND2_X1 U1968 ( .A1(n1921), .A2(n1922), .ZN(n1920) );
  XOR2_X1 U1969 ( .A(n1923), .B(n1924), .Z(Result_8_) );
  AND2_X1 U1970 ( .A1(n1925), .A2(n1926), .ZN(n1924) );
  XOR2_X1 U1971 ( .A(n1927), .B(n1928), .Z(Result_7_) );
  AND2_X1 U1972 ( .A1(n1929), .A2(n1930), .ZN(n1928) );
  XOR2_X1 U1973 ( .A(n1931), .B(n1932), .Z(Result_6_) );
  AND2_X1 U1974 ( .A1(n1933), .A2(n1934), .ZN(n1932) );
  XOR2_X1 U1975 ( .A(n1935), .B(n1936), .Z(Result_5_) );
  AND2_X1 U1976 ( .A1(n1937), .A2(n1938), .ZN(n1936) );
  XOR2_X1 U1977 ( .A(n1939), .B(n1940), .Z(Result_4_) );
  AND2_X1 U1978 ( .A1(n1941), .A2(n1942), .ZN(n1940) );
  XOR2_X1 U1979 ( .A(n1943), .B(n1944), .Z(Result_3_) );
  AND2_X1 U1980 ( .A1(n1945), .A2(n1946), .ZN(n1944) );
  NOR2_X1 U1981 ( .A1(n1947), .A2(n1948), .ZN(Result_31_) );
  NAND2_X1 U1982 ( .A1(n1949), .A2(n1950), .ZN(Result_30_) );
  NAND2_X1 U1983 ( .A1(n1951), .A2(n1952), .ZN(n1950) );
  NAND2_X1 U1984 ( .A1(n1953), .A2(n1954), .ZN(n1952) );
  NAND2_X1 U1985 ( .A1(n1955), .A2(n1956), .ZN(n1954) );
  NAND2_X1 U1986 ( .A1(n1957), .A2(n1958), .ZN(n1949) );
  NAND2_X1 U1987 ( .A1(n1959), .A2(n1960), .ZN(n1958) );
  NAND2_X1 U1988 ( .A1(n1961), .A2(n1948), .ZN(n1960) );
  XOR2_X1 U1989 ( .A(n1962), .B(n1963), .Z(Result_2_) );
  AND2_X1 U1990 ( .A1(n1964), .A2(n1965), .ZN(n1963) );
  XNOR2_X1 U1991 ( .A(n1966), .B(n1967), .ZN(Result_29_) );
  XNOR2_X1 U1992 ( .A(n1968), .B(n1969), .ZN(n1967) );
  XOR2_X1 U1993 ( .A(n1970), .B(n1971), .Z(Result_28_) );
  XOR2_X1 U1994 ( .A(n1972), .B(n1973), .Z(n1971) );
  XOR2_X1 U1995 ( .A(n1974), .B(n1975), .Z(Result_27_) );
  XOR2_X1 U1996 ( .A(n1976), .B(n1977), .Z(n1974) );
  XNOR2_X1 U1997 ( .A(n1978), .B(n1979), .ZN(Result_26_) );
  NAND2_X1 U1998 ( .A1(n1980), .A2(n1981), .ZN(n1978) );
  XOR2_X1 U1999 ( .A(n1982), .B(n1983), .Z(Result_25_) );
  XOR2_X1 U2000 ( .A(n1984), .B(n1985), .Z(n1982) );
  XNOR2_X1 U2001 ( .A(n1986), .B(n1987), .ZN(Result_24_) );
  NAND2_X1 U2002 ( .A1(n1988), .A2(n1989), .ZN(n1986) );
  XOR2_X1 U2003 ( .A(n1990), .B(n1991), .Z(Result_23_) );
  XOR2_X1 U2004 ( .A(n1992), .B(n1993), .Z(n1990) );
  XNOR2_X1 U2005 ( .A(n1994), .B(n1995), .ZN(Result_22_) );
  NAND2_X1 U2006 ( .A1(n1996), .A2(n1997), .ZN(n1994) );
  XOR2_X1 U2007 ( .A(n1998), .B(n1999), .Z(Result_21_) );
  XOR2_X1 U2008 ( .A(n2000), .B(n2001), .Z(n1998) );
  XNOR2_X1 U2009 ( .A(n2002), .B(n2003), .ZN(Result_20_) );
  NAND2_X1 U2010 ( .A1(n2004), .A2(n2005), .ZN(n2002) );
  XNOR2_X1 U2011 ( .A(n2006), .B(n2007), .ZN(Result_1_) );
  NOR2_X1 U2012 ( .A1(n2008), .A2(n2009), .ZN(n2007) );
  XOR2_X1 U2013 ( .A(n2010), .B(n2011), .Z(Result_19_) );
  XOR2_X1 U2014 ( .A(n2012), .B(n2013), .Z(n2010) );
  XNOR2_X1 U2015 ( .A(n2014), .B(n2015), .ZN(Result_18_) );
  NAND2_X1 U2016 ( .A1(n2016), .A2(n2017), .ZN(n2014) );
  XNOR2_X1 U2017 ( .A(n2018), .B(n2019), .ZN(Result_17_) );
  NAND2_X1 U2018 ( .A1(n2020), .A2(n2021), .ZN(n2018) );
  XOR2_X1 U2019 ( .A(n2022), .B(n2023), .Z(Result_16_) );
  XOR2_X1 U2020 ( .A(n2024), .B(n2025), .Z(n2022) );
  NOR2_X1 U2021 ( .A1(n2026), .A2(n1948), .ZN(n2025) );
  XOR2_X1 U2022 ( .A(n2027), .B(n2028), .Z(Result_15_) );
  NOR2_X1 U2023 ( .A1(n2029), .A2(n2030), .ZN(Result_14_) );
  NOR2_X1 U2024 ( .A1(n2031), .A2(n2032), .ZN(n2030) );
  AND2_X1 U2025 ( .A1(n2027), .A2(n2028), .ZN(n2031) );
  XNOR2_X1 U2026 ( .A(n2029), .B(n2033), .ZN(Result_13_) );
  NAND2_X1 U2027 ( .A1(n2034), .A2(n2035), .ZN(n2033) );
  NAND2_X1 U2028 ( .A1(n2036), .A2(n2037), .ZN(n2035) );
  INV_X1 U2029 ( .A(n2038), .ZN(n2037) );
  NAND2_X1 U2030 ( .A1(n2039), .A2(n2040), .ZN(n2036) );
  XOR2_X1 U2031 ( .A(n2041), .B(n2042), .Z(Result_12_) );
  XNOR2_X1 U2032 ( .A(n2043), .B(n2044), .ZN(Result_11_) );
  NAND2_X1 U2033 ( .A1(n2045), .A2(n2046), .ZN(n2044) );
  XNOR2_X1 U2034 ( .A(n2047), .B(n2048), .ZN(Result_10_) );
  NAND2_X1 U2035 ( .A1(n2049), .A2(n2050), .ZN(n2047) );
  NAND2_X1 U2036 ( .A1(n2051), .A2(n2052), .ZN(Result_0_) );
  NAND2_X1 U2037 ( .A1(n2053), .A2(n2054), .ZN(n2052) );
  NOR2_X1 U2038 ( .A1(n2009), .A2(n2055), .ZN(n2051) );
  NOR2_X1 U2039 ( .A1(n2006), .A2(n2008), .ZN(n2055) );
  AND2_X1 U2040 ( .A1(n2056), .A2(n2057), .ZN(n2008) );
  XOR2_X1 U2041 ( .A(n2054), .B(n2058), .Z(n2056) );
  NAND2_X1 U2042 ( .A1(n2053), .A2(n2059), .ZN(n2058) );
  AND2_X1 U2043 ( .A1(n1965), .A2(n2060), .ZN(n2006) );
  NAND2_X1 U2044 ( .A1(n1964), .A2(n1962), .ZN(n2060) );
  NAND2_X1 U2045 ( .A1(n1946), .A2(n2061), .ZN(n1962) );
  NAND2_X1 U2046 ( .A1(n1945), .A2(n1943), .ZN(n2061) );
  NAND2_X1 U2047 ( .A1(n1942), .A2(n2062), .ZN(n1943) );
  NAND2_X1 U2048 ( .A1(n1941), .A2(n1939), .ZN(n2062) );
  NAND2_X1 U2049 ( .A1(n1938), .A2(n2063), .ZN(n1939) );
  NAND2_X1 U2050 ( .A1(n1937), .A2(n1935), .ZN(n2063) );
  NAND2_X1 U2051 ( .A1(n1934), .A2(n2064), .ZN(n1935) );
  NAND2_X1 U2052 ( .A1(n1933), .A2(n1931), .ZN(n2064) );
  NAND2_X1 U2053 ( .A1(n1930), .A2(n2065), .ZN(n1931) );
  NAND2_X1 U2054 ( .A1(n1929), .A2(n1927), .ZN(n2065) );
  NAND2_X1 U2055 ( .A1(n1926), .A2(n2066), .ZN(n1927) );
  NAND2_X1 U2056 ( .A1(n1925), .A2(n1923), .ZN(n2066) );
  NAND2_X1 U2057 ( .A1(n1922), .A2(n2067), .ZN(n1923) );
  NAND2_X1 U2058 ( .A1(n1921), .A2(n1919), .ZN(n2067) );
  NAND2_X1 U2059 ( .A1(n2049), .A2(n2068), .ZN(n1919) );
  NAND2_X1 U2060 ( .A1(n2048), .A2(n2050), .ZN(n2068) );
  NAND2_X1 U2061 ( .A1(n2069), .A2(n2070), .ZN(n2050) );
  XOR2_X1 U2062 ( .A(n2071), .B(n2072), .Z(n2069) );
  NAND2_X1 U2063 ( .A1(n2045), .A2(n2073), .ZN(n2048) );
  NAND2_X1 U2064 ( .A1(n2043), .A2(n2046), .ZN(n2073) );
  NAND2_X1 U2065 ( .A1(n2074), .A2(n2075), .ZN(n2046) );
  NAND2_X1 U2066 ( .A1(n2076), .A2(n2070), .ZN(n2075) );
  NAND2_X1 U2067 ( .A1(n2077), .A2(n2078), .ZN(n2076) );
  NAND2_X1 U2068 ( .A1(n2079), .A2(n2080), .ZN(n2074) );
  AND2_X1 U2069 ( .A1(n2042), .A2(n2041), .ZN(n2043) );
  NAND2_X1 U2070 ( .A1(n2081), .A2(n2082), .ZN(n2041) );
  NAND2_X1 U2071 ( .A1(n2029), .A2(n2038), .ZN(n2082) );
  AND2_X1 U2072 ( .A1(n2083), .A2(n2028), .ZN(n2029) );
  XNOR2_X1 U2073 ( .A(n2084), .B(n2085), .ZN(n2028) );
  XOR2_X1 U2074 ( .A(n2086), .B(n2087), .Z(n2085) );
  NAND2_X1 U2075 ( .A1(n1957), .A2(n2053), .ZN(n2087) );
  AND2_X1 U2076 ( .A1(n2027), .A2(n2032), .ZN(n2083) );
  XOR2_X1 U2077 ( .A(n2040), .B(n2039), .Z(n2032) );
  NAND2_X1 U2078 ( .A1(n2088), .A2(n2089), .ZN(n2027) );
  NAND2_X1 U2079 ( .A1(n2090), .A2(n1951), .ZN(n2089) );
  NOR2_X1 U2080 ( .A1(n2091), .A2(n2026), .ZN(n2090) );
  NOR2_X1 U2081 ( .A1(n2023), .A2(n2024), .ZN(n2091) );
  NAND2_X1 U2082 ( .A1(n2023), .A2(n2024), .ZN(n2088) );
  NAND2_X1 U2083 ( .A1(n2020), .A2(n2092), .ZN(n2024) );
  NAND2_X1 U2084 ( .A1(n2019), .A2(n2021), .ZN(n2092) );
  NAND2_X1 U2085 ( .A1(n2093), .A2(n2094), .ZN(n2021) );
  NAND2_X1 U2086 ( .A1(n1951), .A2(n2095), .ZN(n2094) );
  INV_X1 U2087 ( .A(n2096), .ZN(n2093) );
  XOR2_X1 U2088 ( .A(n2097), .B(n2098), .Z(n2019) );
  XNOR2_X1 U2089 ( .A(n2099), .B(n2100), .ZN(n2097) );
  NAND2_X1 U2090 ( .A1(n1917), .A2(n1957), .ZN(n2099) );
  NAND2_X1 U2091 ( .A1(n2095), .A2(n2096), .ZN(n2020) );
  NAND2_X1 U2092 ( .A1(n2016), .A2(n2102), .ZN(n2096) );
  NAND2_X1 U2093 ( .A1(n2015), .A2(n2017), .ZN(n2102) );
  NAND2_X1 U2094 ( .A1(n2103), .A2(n2104), .ZN(n2017) );
  NAND2_X1 U2095 ( .A1(n1951), .A2(n1917), .ZN(n2104) );
  INV_X1 U2096 ( .A(n2105), .ZN(n2103) );
  XNOR2_X1 U2097 ( .A(n2106), .B(n2107), .ZN(n2015) );
  XNOR2_X1 U2098 ( .A(n2108), .B(n2109), .ZN(n2107) );
  NAND2_X1 U2099 ( .A1(n1917), .A2(n2105), .ZN(n2016) );
  NAND2_X1 U2100 ( .A1(n2110), .A2(n2111), .ZN(n2105) );
  NAND2_X1 U2101 ( .A1(n2011), .A2(n2112), .ZN(n2111) );
  OR2_X1 U2102 ( .A1(n2012), .A2(n2013), .ZN(n2112) );
  XOR2_X1 U2103 ( .A(n2113), .B(n2114), .Z(n2011) );
  XNOR2_X1 U2104 ( .A(n2115), .B(n2116), .ZN(n2113) );
  NAND2_X1 U2105 ( .A1(n2117), .A2(n1957), .ZN(n2115) );
  NAND2_X1 U2106 ( .A1(n2013), .A2(n2012), .ZN(n2110) );
  NAND2_X1 U2107 ( .A1(n2004), .A2(n2118), .ZN(n2012) );
  NAND2_X1 U2108 ( .A1(n2003), .A2(n2005), .ZN(n2118) );
  NAND2_X1 U2109 ( .A1(n2119), .A2(n2120), .ZN(n2005) );
  NAND2_X1 U2110 ( .A1(n1951), .A2(n2117), .ZN(n2120) );
  INV_X1 U2111 ( .A(n2121), .ZN(n2119) );
  XNOR2_X1 U2112 ( .A(n2122), .B(n2123), .ZN(n2003) );
  XNOR2_X1 U2113 ( .A(n2124), .B(n2125), .ZN(n2123) );
  NAND2_X1 U2114 ( .A1(n2117), .A2(n2121), .ZN(n2004) );
  NAND2_X1 U2115 ( .A1(n2126), .A2(n2127), .ZN(n2121) );
  NAND2_X1 U2116 ( .A1(n1999), .A2(n2128), .ZN(n2127) );
  OR2_X1 U2117 ( .A1(n2000), .A2(n2001), .ZN(n2128) );
  XOR2_X1 U2118 ( .A(n2129), .B(n2130), .Z(n1999) );
  XNOR2_X1 U2119 ( .A(n2131), .B(n2132), .ZN(n2129) );
  NAND2_X1 U2120 ( .A1(n2133), .A2(n1957), .ZN(n2131) );
  NAND2_X1 U2121 ( .A1(n2001), .A2(n2000), .ZN(n2126) );
  NAND2_X1 U2122 ( .A1(n1996), .A2(n2134), .ZN(n2000) );
  NAND2_X1 U2123 ( .A1(n1995), .A2(n1997), .ZN(n2134) );
  NAND2_X1 U2124 ( .A1(n2135), .A2(n2136), .ZN(n1997) );
  NAND2_X1 U2125 ( .A1(n1951), .A2(n2133), .ZN(n2136) );
  INV_X1 U2126 ( .A(n2137), .ZN(n2135) );
  XNOR2_X1 U2127 ( .A(n2138), .B(n2139), .ZN(n1995) );
  XNOR2_X1 U2128 ( .A(n2140), .B(n2141), .ZN(n2139) );
  NAND2_X1 U2129 ( .A1(n2133), .A2(n2137), .ZN(n1996) );
  NAND2_X1 U2130 ( .A1(n2142), .A2(n2143), .ZN(n2137) );
  NAND2_X1 U2131 ( .A1(n1991), .A2(n2144), .ZN(n2143) );
  OR2_X1 U2132 ( .A1(n1992), .A2(n1993), .ZN(n2144) );
  XOR2_X1 U2133 ( .A(n2145), .B(n2146), .Z(n1991) );
  XNOR2_X1 U2134 ( .A(n2147), .B(n2148), .ZN(n2145) );
  NAND2_X1 U2135 ( .A1(n2149), .A2(n1957), .ZN(n2147) );
  NAND2_X1 U2136 ( .A1(n1993), .A2(n1992), .ZN(n2142) );
  NAND2_X1 U2137 ( .A1(n1988), .A2(n2150), .ZN(n1992) );
  NAND2_X1 U2138 ( .A1(n1987), .A2(n1989), .ZN(n2150) );
  NAND2_X1 U2139 ( .A1(n2151), .A2(n2152), .ZN(n1989) );
  NAND2_X1 U2140 ( .A1(n1951), .A2(n2149), .ZN(n2152) );
  INV_X1 U2141 ( .A(n2153), .ZN(n2151) );
  XNOR2_X1 U2142 ( .A(n2154), .B(n2155), .ZN(n1987) );
  XNOR2_X1 U2143 ( .A(n2156), .B(n2157), .ZN(n2155) );
  NAND2_X1 U2144 ( .A1(n2149), .A2(n2153), .ZN(n1988) );
  NAND2_X1 U2145 ( .A1(n2158), .A2(n2159), .ZN(n2153) );
  NAND2_X1 U2146 ( .A1(n1983), .A2(n2160), .ZN(n2159) );
  OR2_X1 U2147 ( .A1(n1984), .A2(n1985), .ZN(n2160) );
  XOR2_X1 U2148 ( .A(n2161), .B(n2162), .Z(n1983) );
  XNOR2_X1 U2149 ( .A(n2163), .B(n2164), .ZN(n2161) );
  NAND2_X1 U2150 ( .A1(n2165), .A2(n1957), .ZN(n2163) );
  NAND2_X1 U2151 ( .A1(n1985), .A2(n1984), .ZN(n2158) );
  NAND2_X1 U2152 ( .A1(n1980), .A2(n2166), .ZN(n1984) );
  NAND2_X1 U2153 ( .A1(n1979), .A2(n1981), .ZN(n2166) );
  NAND2_X1 U2154 ( .A1(n2167), .A2(n2168), .ZN(n1981) );
  NAND2_X1 U2155 ( .A1(n1951), .A2(n2165), .ZN(n2168) );
  INV_X1 U2156 ( .A(n2169), .ZN(n2167) );
  XOR2_X1 U2157 ( .A(n2170), .B(n2171), .Z(n1979) );
  XOR2_X1 U2158 ( .A(n2172), .B(n2173), .Z(n2170) );
  NAND2_X1 U2159 ( .A1(n2165), .A2(n2169), .ZN(n1980) );
  NAND2_X1 U2160 ( .A1(n2174), .A2(n2175), .ZN(n2169) );
  NAND2_X1 U2161 ( .A1(n1975), .A2(n2176), .ZN(n2175) );
  NAND2_X1 U2162 ( .A1(n1977), .A2(n1976), .ZN(n2176) );
  INV_X1 U2163 ( .A(n2177), .ZN(n1977) );
  XOR2_X1 U2164 ( .A(n2178), .B(n2179), .Z(n1975) );
  XNOR2_X1 U2165 ( .A(n2180), .B(n2181), .ZN(n2178) );
  NAND2_X1 U2166 ( .A1(n2182), .A2(n1957), .ZN(n2180) );
  NAND2_X1 U2167 ( .A1(n2183), .A2(n2177), .ZN(n2174) );
  NAND2_X1 U2168 ( .A1(n2184), .A2(n2185), .ZN(n2177) );
  NAND2_X1 U2169 ( .A1(n1973), .A2(n2186), .ZN(n2185) );
  NAND2_X1 U2170 ( .A1(n1972), .A2(n1970), .ZN(n2186) );
  NOR2_X1 U2171 ( .A1(n1948), .A2(n2187), .ZN(n1973) );
  OR2_X1 U2172 ( .A1(n1970), .A2(n1972), .ZN(n2184) );
  AND2_X1 U2173 ( .A1(n2188), .A2(n2189), .ZN(n1972) );
  NAND2_X1 U2174 ( .A1(n1969), .A2(n2190), .ZN(n2189) );
  OR2_X1 U2175 ( .A1(n1968), .A2(n1966), .ZN(n2190) );
  AND2_X1 U2176 ( .A1(n2191), .A2(n1951), .ZN(n1969) );
  NAND2_X1 U2177 ( .A1(n1966), .A2(n1968), .ZN(n2188) );
  NAND2_X1 U2178 ( .A1(n2192), .A2(n2193), .ZN(n1968) );
  NAND2_X1 U2179 ( .A1(n2194), .A2(n1957), .ZN(n2193) );
  NOR2_X1 U2180 ( .A1(n2195), .A2(n2196), .ZN(n2194) );
  NOR2_X1 U2181 ( .A1(n2197), .A2(n2198), .ZN(n2195) );
  NAND2_X1 U2182 ( .A1(n2199), .A2(n2200), .ZN(n2192) );
  NOR2_X1 U2183 ( .A1(n2201), .A2(n1947), .ZN(n2199) );
  NOR2_X1 U2184 ( .A1(n2202), .A2(n1955), .ZN(n2201) );
  NOR2_X1 U2185 ( .A1(n1948), .A2(n2203), .ZN(n1966) );
  XOR2_X1 U2186 ( .A(n2204), .B(n2205), .Z(n1970) );
  XNOR2_X1 U2187 ( .A(n2206), .B(n2207), .ZN(n2205) );
  INV_X1 U2188 ( .A(n1976), .ZN(n2183) );
  NAND2_X1 U2189 ( .A1(n1951), .A2(n2208), .ZN(n1976) );
  NOR2_X1 U2190 ( .A1(n1948), .A2(n2209), .ZN(n1985) );
  NOR2_X1 U2191 ( .A1(n1948), .A2(n2210), .ZN(n1993) );
  NOR2_X1 U2192 ( .A1(n1948), .A2(n2211), .ZN(n2001) );
  NOR2_X1 U2193 ( .A1(n1948), .A2(n2212), .ZN(n2013) );
  INV_X1 U2194 ( .A(n1951), .ZN(n1948) );
  NOR2_X1 U2195 ( .A1(n2213), .A2(n2214), .ZN(n1951) );
  NOR2_X1 U2196 ( .A1(c_15_), .A2(d_15_), .ZN(n2214) );
  XNOR2_X1 U2197 ( .A(n2215), .B(n2216), .ZN(n2023) );
  XOR2_X1 U2198 ( .A(n2217), .B(n2218), .Z(n2216) );
  NAND2_X1 U2199 ( .A1(n2095), .A2(n1957), .ZN(n2218) );
  NOR2_X1 U2200 ( .A1(n2219), .A2(n2220), .ZN(n2081) );
  INV_X1 U2201 ( .A(n2034), .ZN(n2219) );
  NAND2_X1 U2202 ( .A1(n2221), .A2(n2038), .ZN(n2034) );
  NOR2_X1 U2203 ( .A1(n2220), .A2(n2222), .ZN(n2038) );
  AND2_X1 U2204 ( .A1(n2223), .A2(n2224), .ZN(n2222) );
  NOR2_X1 U2205 ( .A1(n2224), .A2(n2223), .ZN(n2220) );
  XNOR2_X1 U2206 ( .A(n2225), .B(n2226), .ZN(n2223) );
  XNOR2_X1 U2207 ( .A(n2227), .B(n2228), .ZN(n2225) );
  NAND2_X1 U2208 ( .A1(n2229), .A2(n2053), .ZN(n2227) );
  NAND2_X1 U2209 ( .A1(n2230), .A2(n2231), .ZN(n2224) );
  NAND2_X1 U2210 ( .A1(n2232), .A2(n2233), .ZN(n2231) );
  NAND2_X1 U2211 ( .A1(n2234), .A2(n2235), .ZN(n2233) );
  OR2_X1 U2212 ( .A1(n2235), .A2(n2234), .ZN(n2230) );
  AND2_X1 U2213 ( .A1(n2040), .A2(n2039), .ZN(n2221) );
  XNOR2_X1 U2214 ( .A(n2235), .B(n2236), .ZN(n2039) );
  XOR2_X1 U2215 ( .A(n2232), .B(n2234), .Z(n2236) );
  NOR2_X1 U2216 ( .A1(n2198), .A2(n2026), .ZN(n2234) );
  AND2_X1 U2217 ( .A1(n2237), .A2(n2238), .ZN(n2232) );
  NAND2_X1 U2218 ( .A1(n2239), .A2(n2200), .ZN(n2238) );
  NOR2_X1 U2219 ( .A1(n2240), .A2(n2241), .ZN(n2239) );
  NOR2_X1 U2220 ( .A1(n2242), .A2(n2243), .ZN(n2240) );
  NAND2_X1 U2221 ( .A1(n2242), .A2(n2243), .ZN(n2237) );
  XNOR2_X1 U2222 ( .A(n2244), .B(n2245), .ZN(n2235) );
  XNOR2_X1 U2223 ( .A(n2246), .B(n2247), .ZN(n2244) );
  NAND2_X1 U2224 ( .A1(n2248), .A2(n2249), .ZN(n2040) );
  NAND2_X1 U2225 ( .A1(n2250), .A2(n1957), .ZN(n2249) );
  INV_X1 U2226 ( .A(n1955), .ZN(n1957) );
  NOR2_X1 U2227 ( .A1(n2251), .A2(n2026), .ZN(n2250) );
  NOR2_X1 U2228 ( .A1(n2084), .A2(n2086), .ZN(n2251) );
  NAND2_X1 U2229 ( .A1(n2084), .A2(n2086), .ZN(n2248) );
  NAND2_X1 U2230 ( .A1(n2252), .A2(n2253), .ZN(n2086) );
  NAND2_X1 U2231 ( .A1(n2254), .A2(n2095), .ZN(n2253) );
  NOR2_X1 U2232 ( .A1(n2255), .A2(n1955), .ZN(n2254) );
  NOR2_X1 U2233 ( .A1(n2215), .A2(n2217), .ZN(n2255) );
  NAND2_X1 U2234 ( .A1(n2215), .A2(n2217), .ZN(n2252) );
  NAND2_X1 U2235 ( .A1(n2256), .A2(n2257), .ZN(n2217) );
  NAND2_X1 U2236 ( .A1(n2258), .A2(n2101), .ZN(n2257) );
  NOR2_X1 U2237 ( .A1(n2259), .A2(n1955), .ZN(n2258) );
  NOR2_X1 U2238 ( .A1(n2098), .A2(n2100), .ZN(n2259) );
  NAND2_X1 U2239 ( .A1(n2098), .A2(n2100), .ZN(n2256) );
  NAND2_X1 U2240 ( .A1(n2260), .A2(n2261), .ZN(n2100) );
  NAND2_X1 U2241 ( .A1(n2109), .A2(n2262), .ZN(n2261) );
  OR2_X1 U2242 ( .A1(n2108), .A2(n2106), .ZN(n2262) );
  NOR2_X1 U2243 ( .A1(n2212), .A2(n1955), .ZN(n2109) );
  NAND2_X1 U2244 ( .A1(n2106), .A2(n2108), .ZN(n2260) );
  NAND2_X1 U2245 ( .A1(n2263), .A2(n2264), .ZN(n2108) );
  NAND2_X1 U2246 ( .A1(n2265), .A2(n2117), .ZN(n2264) );
  NOR2_X1 U2247 ( .A1(n2266), .A2(n1955), .ZN(n2265) );
  NOR2_X1 U2248 ( .A1(n2114), .A2(n2116), .ZN(n2266) );
  NAND2_X1 U2249 ( .A1(n2114), .A2(n2116), .ZN(n2263) );
  NAND2_X1 U2250 ( .A1(n2267), .A2(n2268), .ZN(n2116) );
  NAND2_X1 U2251 ( .A1(n2125), .A2(n2269), .ZN(n2268) );
  OR2_X1 U2252 ( .A1(n2124), .A2(n2122), .ZN(n2269) );
  NOR2_X1 U2253 ( .A1(n2211), .A2(n1955), .ZN(n2125) );
  NAND2_X1 U2254 ( .A1(n2122), .A2(n2124), .ZN(n2267) );
  NAND2_X1 U2255 ( .A1(n2270), .A2(n2271), .ZN(n2124) );
  NAND2_X1 U2256 ( .A1(n2272), .A2(n2133), .ZN(n2271) );
  NOR2_X1 U2257 ( .A1(n2273), .A2(n1955), .ZN(n2272) );
  NOR2_X1 U2258 ( .A1(n2130), .A2(n2132), .ZN(n2273) );
  NAND2_X1 U2259 ( .A1(n2130), .A2(n2132), .ZN(n2270) );
  NAND2_X1 U2260 ( .A1(n2274), .A2(n2275), .ZN(n2132) );
  NAND2_X1 U2261 ( .A1(n2141), .A2(n2276), .ZN(n2275) );
  OR2_X1 U2262 ( .A1(n2140), .A2(n2138), .ZN(n2276) );
  NOR2_X1 U2263 ( .A1(n2210), .A2(n1955), .ZN(n2141) );
  NAND2_X1 U2264 ( .A1(n2138), .A2(n2140), .ZN(n2274) );
  NAND2_X1 U2265 ( .A1(n2277), .A2(n2278), .ZN(n2140) );
  NAND2_X1 U2266 ( .A1(n2279), .A2(n2149), .ZN(n2278) );
  NOR2_X1 U2267 ( .A1(n2280), .A2(n1955), .ZN(n2279) );
  NOR2_X1 U2268 ( .A1(n2146), .A2(n2148), .ZN(n2280) );
  NAND2_X1 U2269 ( .A1(n2146), .A2(n2148), .ZN(n2277) );
  NAND2_X1 U2270 ( .A1(n2281), .A2(n2282), .ZN(n2148) );
  NAND2_X1 U2271 ( .A1(n2157), .A2(n2283), .ZN(n2282) );
  OR2_X1 U2272 ( .A1(n2156), .A2(n2154), .ZN(n2283) );
  NOR2_X1 U2273 ( .A1(n2209), .A2(n1955), .ZN(n2157) );
  NAND2_X1 U2274 ( .A1(n2154), .A2(n2156), .ZN(n2281) );
  NAND2_X1 U2275 ( .A1(n2284), .A2(n2285), .ZN(n2156) );
  NAND2_X1 U2276 ( .A1(n2286), .A2(n2165), .ZN(n2285) );
  NOR2_X1 U2277 ( .A1(n2287), .A2(n1955), .ZN(n2286) );
  NOR2_X1 U2278 ( .A1(n2162), .A2(n2164), .ZN(n2287) );
  NAND2_X1 U2279 ( .A1(n2162), .A2(n2164), .ZN(n2284) );
  NAND2_X1 U2280 ( .A1(n2288), .A2(n2289), .ZN(n2164) );
  NAND2_X1 U2281 ( .A1(n2173), .A2(n2290), .ZN(n2289) );
  OR2_X1 U2282 ( .A1(n2172), .A2(n2171), .ZN(n2290) );
  NOR2_X1 U2283 ( .A1(n2291), .A2(n1955), .ZN(n2173) );
  NAND2_X1 U2284 ( .A1(n2171), .A2(n2172), .ZN(n2288) );
  NAND2_X1 U2285 ( .A1(n2292), .A2(n2293), .ZN(n2172) );
  NAND2_X1 U2286 ( .A1(n2294), .A2(n2182), .ZN(n2293) );
  NOR2_X1 U2287 ( .A1(n2295), .A2(n1955), .ZN(n2294) );
  NOR2_X1 U2288 ( .A1(n2179), .A2(n2181), .ZN(n2295) );
  NAND2_X1 U2289 ( .A1(n2179), .A2(n2181), .ZN(n2292) );
  NAND2_X1 U2290 ( .A1(n2296), .A2(n2297), .ZN(n2181) );
  NAND2_X1 U2291 ( .A1(n2204), .A2(n2298), .ZN(n2297) );
  NAND2_X1 U2292 ( .A1(n2206), .A2(n2207), .ZN(n2298) );
  NOR2_X1 U2293 ( .A1(n2203), .A2(n1955), .ZN(n2204) );
  OR2_X1 U2294 ( .A1(n2207), .A2(n2206), .ZN(n2296) );
  AND2_X1 U2295 ( .A1(n2299), .A2(n2300), .ZN(n2206) );
  NAND2_X1 U2296 ( .A1(n2301), .A2(n2200), .ZN(n2300) );
  NOR2_X1 U2297 ( .A1(n2302), .A2(n2196), .ZN(n2301) );
  NOR2_X1 U2298 ( .A1(n2197), .A2(n2303), .ZN(n2302) );
  NAND2_X1 U2299 ( .A1(n2304), .A2(n2229), .ZN(n2299) );
  NOR2_X1 U2300 ( .A1(n2305), .A2(n1947), .ZN(n2304) );
  NOR2_X1 U2301 ( .A1(n2202), .A2(n2198), .ZN(n2305) );
  NAND2_X1 U2302 ( .A1(n2191), .A2(n2200), .ZN(n2207) );
  NOR2_X1 U2303 ( .A1(n1955), .A2(n2306), .ZN(n2191) );
  XOR2_X1 U2304 ( .A(d_14_), .B(c_14_), .Z(n2307) );
  XNOR2_X1 U2305 ( .A(n2308), .B(n2309), .ZN(n2179) );
  XNOR2_X1 U2306 ( .A(n2310), .B(n2311), .ZN(n2309) );
  XOR2_X1 U2307 ( .A(n2312), .B(n2313), .Z(n2171) );
  XNOR2_X1 U2308 ( .A(n2314), .B(n2315), .ZN(n2312) );
  NAND2_X1 U2309 ( .A1(n2200), .A2(n2182), .ZN(n2314) );
  XNOR2_X1 U2310 ( .A(n2316), .B(n2317), .ZN(n2162) );
  XNOR2_X1 U2311 ( .A(n2318), .B(n2319), .ZN(n2317) );
  XOR2_X1 U2312 ( .A(n2320), .B(n2321), .Z(n2154) );
  XNOR2_X1 U2313 ( .A(n2322), .B(n2323), .ZN(n2320) );
  NAND2_X1 U2314 ( .A1(n2200), .A2(n2165), .ZN(n2322) );
  XNOR2_X1 U2315 ( .A(n2324), .B(n2325), .ZN(n2146) );
  XNOR2_X1 U2316 ( .A(n2326), .B(n2327), .ZN(n2325) );
  XOR2_X1 U2317 ( .A(n2328), .B(n2329), .Z(n2138) );
  XNOR2_X1 U2318 ( .A(n2330), .B(n2331), .ZN(n2328) );
  NAND2_X1 U2319 ( .A1(n2200), .A2(n2149), .ZN(n2330) );
  XNOR2_X1 U2320 ( .A(n2332), .B(n2333), .ZN(n2130) );
  XNOR2_X1 U2321 ( .A(n2334), .B(n2335), .ZN(n2333) );
  XOR2_X1 U2322 ( .A(n2336), .B(n2337), .Z(n2122) );
  XNOR2_X1 U2323 ( .A(n2338), .B(n2339), .ZN(n2336) );
  NAND2_X1 U2324 ( .A1(n2200), .A2(n2133), .ZN(n2338) );
  XNOR2_X1 U2325 ( .A(n2340), .B(n2341), .ZN(n2114) );
  XNOR2_X1 U2326 ( .A(n2342), .B(n2343), .ZN(n2341) );
  XOR2_X1 U2327 ( .A(n2344), .B(n2345), .Z(n2106) );
  XNOR2_X1 U2328 ( .A(n2346), .B(n2347), .ZN(n2344) );
  NAND2_X1 U2329 ( .A1(n2200), .A2(n2117), .ZN(n2346) );
  XNOR2_X1 U2330 ( .A(n2348), .B(n2349), .ZN(n2098) );
  XNOR2_X1 U2331 ( .A(n2350), .B(n2351), .ZN(n2349) );
  XOR2_X1 U2332 ( .A(n2352), .B(n2353), .Z(n2215) );
  XNOR2_X1 U2333 ( .A(n2354), .B(n2355), .ZN(n2352) );
  NAND2_X1 U2334 ( .A1(n2200), .A2(n2101), .ZN(n2354) );
  XNOR2_X1 U2335 ( .A(n2242), .B(n2356), .ZN(n2084) );
  XOR2_X1 U2336 ( .A(n2243), .B(n2357), .Z(n2356) );
  NAND2_X1 U2337 ( .A1(n2200), .A2(n2095), .ZN(n2357) );
  NAND2_X1 U2338 ( .A1(n2358), .A2(n2359), .ZN(n2243) );
  NAND2_X1 U2339 ( .A1(n2360), .A2(n2200), .ZN(n2359) );
  NOR2_X1 U2340 ( .A1(n2361), .A2(n2362), .ZN(n2360) );
  NOR2_X1 U2341 ( .A1(n2353), .A2(n2355), .ZN(n2361) );
  NAND2_X1 U2342 ( .A1(n2353), .A2(n2355), .ZN(n2358) );
  NAND2_X1 U2343 ( .A1(n2363), .A2(n2364), .ZN(n2355) );
  NAND2_X1 U2344 ( .A1(n2351), .A2(n2365), .ZN(n2364) );
  OR2_X1 U2345 ( .A1(n2350), .A2(n2348), .ZN(n2365) );
  NOR2_X1 U2346 ( .A1(n2198), .A2(n2212), .ZN(n2351) );
  NAND2_X1 U2347 ( .A1(n2348), .A2(n2350), .ZN(n2363) );
  NAND2_X1 U2348 ( .A1(n2366), .A2(n2367), .ZN(n2350) );
  NAND2_X1 U2349 ( .A1(n2368), .A2(n2200), .ZN(n2367) );
  NOR2_X1 U2350 ( .A1(n2369), .A2(n2370), .ZN(n2368) );
  NOR2_X1 U2351 ( .A1(n2345), .A2(n2347), .ZN(n2369) );
  NAND2_X1 U2352 ( .A1(n2345), .A2(n2347), .ZN(n2366) );
  NAND2_X1 U2353 ( .A1(n2371), .A2(n2372), .ZN(n2347) );
  NAND2_X1 U2354 ( .A1(n2343), .A2(n2373), .ZN(n2372) );
  OR2_X1 U2355 ( .A1(n2342), .A2(n2340), .ZN(n2373) );
  NOR2_X1 U2356 ( .A1(n2198), .A2(n2211), .ZN(n2343) );
  NAND2_X1 U2357 ( .A1(n2340), .A2(n2342), .ZN(n2371) );
  NAND2_X1 U2358 ( .A1(n2374), .A2(n2375), .ZN(n2342) );
  NAND2_X1 U2359 ( .A1(n2376), .A2(n2200), .ZN(n2375) );
  NOR2_X1 U2360 ( .A1(n2377), .A2(n2378), .ZN(n2376) );
  NOR2_X1 U2361 ( .A1(n2337), .A2(n2339), .ZN(n2377) );
  NAND2_X1 U2362 ( .A1(n2337), .A2(n2339), .ZN(n2374) );
  NAND2_X1 U2363 ( .A1(n2379), .A2(n2380), .ZN(n2339) );
  NAND2_X1 U2364 ( .A1(n2335), .A2(n2381), .ZN(n2380) );
  OR2_X1 U2365 ( .A1(n2334), .A2(n2332), .ZN(n2381) );
  NOR2_X1 U2366 ( .A1(n2198), .A2(n2210), .ZN(n2335) );
  NAND2_X1 U2367 ( .A1(n2332), .A2(n2334), .ZN(n2379) );
  NAND2_X1 U2368 ( .A1(n2382), .A2(n2383), .ZN(n2334) );
  NAND2_X1 U2369 ( .A1(n2384), .A2(n2200), .ZN(n2383) );
  NOR2_X1 U2370 ( .A1(n2385), .A2(n2386), .ZN(n2384) );
  NOR2_X1 U2371 ( .A1(n2329), .A2(n2331), .ZN(n2385) );
  NAND2_X1 U2372 ( .A1(n2329), .A2(n2331), .ZN(n2382) );
  NAND2_X1 U2373 ( .A1(n2387), .A2(n2388), .ZN(n2331) );
  NAND2_X1 U2374 ( .A1(n2327), .A2(n2389), .ZN(n2388) );
  OR2_X1 U2375 ( .A1(n2326), .A2(n2324), .ZN(n2389) );
  NOR2_X1 U2376 ( .A1(n2198), .A2(n2209), .ZN(n2327) );
  NAND2_X1 U2377 ( .A1(n2324), .A2(n2326), .ZN(n2387) );
  NAND2_X1 U2378 ( .A1(n2390), .A2(n2391), .ZN(n2326) );
  NAND2_X1 U2379 ( .A1(n2392), .A2(n2200), .ZN(n2391) );
  NOR2_X1 U2380 ( .A1(n2393), .A2(n2394), .ZN(n2392) );
  NOR2_X1 U2381 ( .A1(n2321), .A2(n2323), .ZN(n2393) );
  NAND2_X1 U2382 ( .A1(n2321), .A2(n2323), .ZN(n2390) );
  NAND2_X1 U2383 ( .A1(n2395), .A2(n2396), .ZN(n2323) );
  NAND2_X1 U2384 ( .A1(n2319), .A2(n2397), .ZN(n2396) );
  OR2_X1 U2385 ( .A1(n2318), .A2(n2316), .ZN(n2397) );
  NOR2_X1 U2386 ( .A1(n2198), .A2(n2291), .ZN(n2319) );
  NAND2_X1 U2387 ( .A1(n2316), .A2(n2318), .ZN(n2395) );
  NAND2_X1 U2388 ( .A1(n2398), .A2(n2399), .ZN(n2318) );
  NAND2_X1 U2389 ( .A1(n2400), .A2(n2200), .ZN(n2399) );
  NOR2_X1 U2390 ( .A1(n2401), .A2(n2187), .ZN(n2400) );
  NOR2_X1 U2391 ( .A1(n2313), .A2(n2315), .ZN(n2401) );
  NAND2_X1 U2392 ( .A1(n2313), .A2(n2315), .ZN(n2398) );
  NAND2_X1 U2393 ( .A1(n2402), .A2(n2403), .ZN(n2315) );
  NAND2_X1 U2394 ( .A1(n2308), .A2(n2404), .ZN(n2403) );
  NAND2_X1 U2395 ( .A1(n2310), .A2(n2311), .ZN(n2404) );
  NOR2_X1 U2396 ( .A1(n2198), .A2(n2203), .ZN(n2308) );
  INV_X1 U2397 ( .A(n2200), .ZN(n2198) );
  OR2_X1 U2398 ( .A1(n2311), .A2(n2310), .ZN(n2402) );
  AND2_X1 U2399 ( .A1(n2405), .A2(n2406), .ZN(n2310) );
  NAND2_X1 U2400 ( .A1(n2407), .A2(n2229), .ZN(n2406) );
  NOR2_X1 U2401 ( .A1(n2408), .A2(n2196), .ZN(n2407) );
  NOR2_X1 U2402 ( .A1(n2197), .A2(n2409), .ZN(n2408) );
  NAND2_X1 U2403 ( .A1(n2410), .A2(n1961), .ZN(n2405) );
  NOR2_X1 U2404 ( .A1(n2411), .A2(n2409), .ZN(n2410) );
  NOR2_X1 U2405 ( .A1(n2202), .A2(n2303), .ZN(n2411) );
  NAND2_X1 U2406 ( .A1(n2412), .A2(n2200), .ZN(n2311) );
  XOR2_X1 U2407 ( .A(d_13_), .B(c_13_), .Z(n2414) );
  NOR2_X1 U2408 ( .A1(n2306), .A2(n2303), .ZN(n2412) );
  XNOR2_X1 U2409 ( .A(n2415), .B(n2416), .ZN(n2313) );
  XNOR2_X1 U2410 ( .A(n2417), .B(n2418), .ZN(n2416) );
  XOR2_X1 U2411 ( .A(n2419), .B(n2420), .Z(n2316) );
  XNOR2_X1 U2412 ( .A(n2421), .B(n2422), .ZN(n2419) );
  NAND2_X1 U2413 ( .A1(n2229), .A2(n2182), .ZN(n2421) );
  XOR2_X1 U2414 ( .A(n2423), .B(n2424), .Z(n2321) );
  XOR2_X1 U2415 ( .A(n2425), .B(n2426), .Z(n2423) );
  XOR2_X1 U2416 ( .A(n2427), .B(n2428), .Z(n2324) );
  XNOR2_X1 U2417 ( .A(n2429), .B(n2430), .ZN(n2427) );
  NAND2_X1 U2418 ( .A1(n2229), .A2(n2165), .ZN(n2429) );
  XNOR2_X1 U2419 ( .A(n2431), .B(n2432), .ZN(n2329) );
  XNOR2_X1 U2420 ( .A(n2433), .B(n2434), .ZN(n2432) );
  XOR2_X1 U2421 ( .A(n2435), .B(n2436), .Z(n2332) );
  XNOR2_X1 U2422 ( .A(n2437), .B(n2438), .ZN(n2435) );
  NAND2_X1 U2423 ( .A1(n2229), .A2(n2149), .ZN(n2437) );
  XOR2_X1 U2424 ( .A(n2439), .B(n2440), .Z(n2337) );
  XOR2_X1 U2425 ( .A(n2441), .B(n2442), .Z(n2439) );
  XOR2_X1 U2426 ( .A(n2443), .B(n2444), .Z(n2340) );
  XNOR2_X1 U2427 ( .A(n2445), .B(n2446), .ZN(n2443) );
  NAND2_X1 U2428 ( .A1(n2229), .A2(n2133), .ZN(n2445) );
  XNOR2_X1 U2429 ( .A(n2447), .B(n2448), .ZN(n2345) );
  XNOR2_X1 U2430 ( .A(n2449), .B(n2450), .ZN(n2448) );
  XOR2_X1 U2431 ( .A(n2451), .B(n2452), .Z(n2348) );
  XNOR2_X1 U2432 ( .A(n2453), .B(n2454), .ZN(n2451) );
  NAND2_X1 U2433 ( .A1(n2229), .A2(n2117), .ZN(n2453) );
  XNOR2_X1 U2434 ( .A(n2455), .B(n2456), .ZN(n2353) );
  XOR2_X1 U2435 ( .A(n2457), .B(n2458), .Z(n2456) );
  NAND2_X1 U2436 ( .A1(n2229), .A2(n2459), .ZN(n2458) );
  XNOR2_X1 U2437 ( .A(n2460), .B(n2461), .ZN(n2242) );
  XNOR2_X1 U2438 ( .A(n2462), .B(n2463), .ZN(n2461) );
  XOR2_X1 U2439 ( .A(n2080), .B(n2079), .Z(n2042) );
  NAND2_X1 U2440 ( .A1(n2464), .A2(n2465), .ZN(n2045) );
  AND2_X1 U2441 ( .A1(n2070), .A2(n2080), .ZN(n2465) );
  NAND2_X1 U2442 ( .A1(n2466), .A2(n2467), .ZN(n2080) );
  NAND2_X1 U2443 ( .A1(n2468), .A2(n2229), .ZN(n2467) );
  NOR2_X1 U2444 ( .A1(n2469), .A2(n2026), .ZN(n2468) );
  NOR2_X1 U2445 ( .A1(n2226), .A2(n2228), .ZN(n2469) );
  NAND2_X1 U2446 ( .A1(n2226), .A2(n2228), .ZN(n2466) );
  NAND2_X1 U2447 ( .A1(n2470), .A2(n2471), .ZN(n2228) );
  NAND2_X1 U2448 ( .A1(n2247), .A2(n2472), .ZN(n2471) );
  NAND2_X1 U2449 ( .A1(n2246), .A2(n2245), .ZN(n2472) );
  NOR2_X1 U2450 ( .A1(n2303), .A2(n2241), .ZN(n2247) );
  OR2_X1 U2451 ( .A1(n2245), .A2(n2246), .ZN(n2470) );
  AND2_X1 U2452 ( .A1(n2473), .A2(n2474), .ZN(n2246) );
  NAND2_X1 U2453 ( .A1(n2463), .A2(n2475), .ZN(n2474) );
  OR2_X1 U2454 ( .A1(n2462), .A2(n2460), .ZN(n2475) );
  NOR2_X1 U2455 ( .A1(n2303), .A2(n2362), .ZN(n2463) );
  NAND2_X1 U2456 ( .A1(n2460), .A2(n2462), .ZN(n2473) );
  NAND2_X1 U2457 ( .A1(n2476), .A2(n2477), .ZN(n2462) );
  NAND2_X1 U2458 ( .A1(n2478), .A2(n2229), .ZN(n2477) );
  NOR2_X1 U2459 ( .A1(n2479), .A2(n2212), .ZN(n2478) );
  NOR2_X1 U2460 ( .A1(n2455), .A2(n2457), .ZN(n2479) );
  NAND2_X1 U2461 ( .A1(n2455), .A2(n2457), .ZN(n2476) );
  NAND2_X1 U2462 ( .A1(n2480), .A2(n2481), .ZN(n2457) );
  NAND2_X1 U2463 ( .A1(n2482), .A2(n2229), .ZN(n2481) );
  NOR2_X1 U2464 ( .A1(n2483), .A2(n2370), .ZN(n2482) );
  NOR2_X1 U2465 ( .A1(n2452), .A2(n2454), .ZN(n2483) );
  NAND2_X1 U2466 ( .A1(n2452), .A2(n2454), .ZN(n2480) );
  NAND2_X1 U2467 ( .A1(n2484), .A2(n2485), .ZN(n2454) );
  NAND2_X1 U2468 ( .A1(n2450), .A2(n2486), .ZN(n2485) );
  OR2_X1 U2469 ( .A1(n2449), .A2(n2447), .ZN(n2486) );
  NOR2_X1 U2470 ( .A1(n2303), .A2(n2211), .ZN(n2450) );
  NAND2_X1 U2471 ( .A1(n2447), .A2(n2449), .ZN(n2484) );
  NAND2_X1 U2472 ( .A1(n2487), .A2(n2488), .ZN(n2449) );
  NAND2_X1 U2473 ( .A1(n2489), .A2(n2229), .ZN(n2488) );
  NOR2_X1 U2474 ( .A1(n2490), .A2(n2378), .ZN(n2489) );
  NOR2_X1 U2475 ( .A1(n2444), .A2(n2446), .ZN(n2490) );
  NAND2_X1 U2476 ( .A1(n2444), .A2(n2446), .ZN(n2487) );
  NAND2_X1 U2477 ( .A1(n2491), .A2(n2492), .ZN(n2446) );
  NAND2_X1 U2478 ( .A1(n2442), .A2(n2493), .ZN(n2492) );
  OR2_X1 U2479 ( .A1(n2441), .A2(n2440), .ZN(n2493) );
  NOR2_X1 U2480 ( .A1(n2303), .A2(n2210), .ZN(n2442) );
  NAND2_X1 U2481 ( .A1(n2440), .A2(n2441), .ZN(n2491) );
  NAND2_X1 U2482 ( .A1(n2494), .A2(n2495), .ZN(n2441) );
  NAND2_X1 U2483 ( .A1(n2496), .A2(n2229), .ZN(n2495) );
  NOR2_X1 U2484 ( .A1(n2497), .A2(n2386), .ZN(n2496) );
  NOR2_X1 U2485 ( .A1(n2436), .A2(n2438), .ZN(n2497) );
  NAND2_X1 U2486 ( .A1(n2436), .A2(n2438), .ZN(n2494) );
  NAND2_X1 U2487 ( .A1(n2498), .A2(n2499), .ZN(n2438) );
  NAND2_X1 U2488 ( .A1(n2434), .A2(n2500), .ZN(n2499) );
  OR2_X1 U2489 ( .A1(n2433), .A2(n2431), .ZN(n2500) );
  NOR2_X1 U2490 ( .A1(n2303), .A2(n2209), .ZN(n2434) );
  NAND2_X1 U2491 ( .A1(n2431), .A2(n2433), .ZN(n2498) );
  NAND2_X1 U2492 ( .A1(n2501), .A2(n2502), .ZN(n2433) );
  NAND2_X1 U2493 ( .A1(n2503), .A2(n2229), .ZN(n2502) );
  NOR2_X1 U2494 ( .A1(n2504), .A2(n2394), .ZN(n2503) );
  NOR2_X1 U2495 ( .A1(n2428), .A2(n2430), .ZN(n2504) );
  NAND2_X1 U2496 ( .A1(n2428), .A2(n2430), .ZN(n2501) );
  NAND2_X1 U2497 ( .A1(n2505), .A2(n2506), .ZN(n2430) );
  NAND2_X1 U2498 ( .A1(n2426), .A2(n2507), .ZN(n2506) );
  OR2_X1 U2499 ( .A1(n2425), .A2(n2424), .ZN(n2507) );
  NOR2_X1 U2500 ( .A1(n2303), .A2(n2291), .ZN(n2426) );
  NAND2_X1 U2501 ( .A1(n2424), .A2(n2425), .ZN(n2505) );
  NAND2_X1 U2502 ( .A1(n2508), .A2(n2509), .ZN(n2425) );
  NAND2_X1 U2503 ( .A1(n2510), .A2(n2229), .ZN(n2509) );
  NOR2_X1 U2504 ( .A1(n2511), .A2(n2187), .ZN(n2510) );
  NOR2_X1 U2505 ( .A1(n2420), .A2(n2422), .ZN(n2511) );
  NAND2_X1 U2506 ( .A1(n2420), .A2(n2422), .ZN(n2508) );
  NAND2_X1 U2507 ( .A1(n2512), .A2(n2513), .ZN(n2422) );
  NAND2_X1 U2508 ( .A1(n2415), .A2(n2514), .ZN(n2513) );
  NAND2_X1 U2509 ( .A1(n2418), .A2(n2417), .ZN(n2514) );
  NOR2_X1 U2510 ( .A1(n2303), .A2(n2203), .ZN(n2415) );
  INV_X1 U2511 ( .A(n2229), .ZN(n2303) );
  OR2_X1 U2512 ( .A1(n2417), .A2(n2418), .ZN(n2512) );
  AND2_X1 U2513 ( .A1(n2515), .A2(n2516), .ZN(n2418) );
  NAND2_X1 U2514 ( .A1(n2517), .A2(n2518), .ZN(n2516) );
  NAND2_X1 U2515 ( .A1(n1953), .A2(n2519), .ZN(n2518) );
  NAND2_X1 U2516 ( .A1(n2520), .A2(n1956), .ZN(n2519) );
  NAND2_X1 U2517 ( .A1(n2521), .A2(n2522), .ZN(n2515) );
  NAND2_X1 U2518 ( .A1(n1959), .A2(n2523), .ZN(n2522) );
  NAND2_X1 U2519 ( .A1(n1961), .A2(n2409), .ZN(n2523) );
  NAND2_X1 U2520 ( .A1(n2524), .A2(n2229), .ZN(n2417) );
  XNOR2_X1 U2521 ( .A(c_12_), .B(d_12_), .ZN(n2525) );
  NOR2_X1 U2522 ( .A1(n2306), .A2(n2409), .ZN(n2524) );
  XNOR2_X1 U2523 ( .A(n2527), .B(n2528), .ZN(n2420) );
  XNOR2_X1 U2524 ( .A(n2529), .B(n2530), .ZN(n2528) );
  XOR2_X1 U2525 ( .A(n2531), .B(n2532), .Z(n2424) );
  XNOR2_X1 U2526 ( .A(n2533), .B(n2534), .ZN(n2531) );
  NAND2_X1 U2527 ( .A1(n2182), .A2(n2517), .ZN(n2533) );
  XNOR2_X1 U2528 ( .A(n2535), .B(n2536), .ZN(n2428) );
  XNOR2_X1 U2529 ( .A(n2537), .B(n2538), .ZN(n2536) );
  XOR2_X1 U2530 ( .A(n2539), .B(n2540), .Z(n2431) );
  XNOR2_X1 U2531 ( .A(n2541), .B(n2542), .ZN(n2539) );
  NAND2_X1 U2532 ( .A1(n2165), .A2(n2517), .ZN(n2541) );
  XNOR2_X1 U2533 ( .A(n2543), .B(n2544), .ZN(n2436) );
  XNOR2_X1 U2534 ( .A(n2545), .B(n2546), .ZN(n2544) );
  XOR2_X1 U2535 ( .A(n2547), .B(n2548), .Z(n2440) );
  XNOR2_X1 U2536 ( .A(n2549), .B(n2550), .ZN(n2547) );
  NAND2_X1 U2537 ( .A1(n2149), .A2(n2517), .ZN(n2549) );
  XNOR2_X1 U2538 ( .A(n2551), .B(n2552), .ZN(n2444) );
  XNOR2_X1 U2539 ( .A(n2553), .B(n2554), .ZN(n2552) );
  XOR2_X1 U2540 ( .A(n2555), .B(n2556), .Z(n2447) );
  XNOR2_X1 U2541 ( .A(n2557), .B(n2558), .ZN(n2555) );
  NAND2_X1 U2542 ( .A1(n2133), .A2(n2517), .ZN(n2557) );
  XNOR2_X1 U2543 ( .A(n2559), .B(n2560), .ZN(n2452) );
  XNOR2_X1 U2544 ( .A(n2561), .B(n2562), .ZN(n2560) );
  XOR2_X1 U2545 ( .A(n2563), .B(n2564), .Z(n2455) );
  XOR2_X1 U2546 ( .A(n2565), .B(n2566), .Z(n2563) );
  XOR2_X1 U2547 ( .A(n2567), .B(n2568), .Z(n2460) );
  XNOR2_X1 U2548 ( .A(n2569), .B(n2570), .ZN(n2567) );
  NAND2_X1 U2549 ( .A1(n2459), .A2(n2517), .ZN(n2569) );
  XOR2_X1 U2550 ( .A(n2571), .B(n2572), .Z(n2245) );
  XOR2_X1 U2551 ( .A(n2573), .B(n2574), .Z(n2572) );
  NAND2_X1 U2552 ( .A1(n1917), .A2(n2517), .ZN(n2574) );
  XNOR2_X1 U2553 ( .A(n2575), .B(n2576), .ZN(n2226) );
  XOR2_X1 U2554 ( .A(n2577), .B(n2578), .Z(n2576) );
  NAND2_X1 U2555 ( .A1(n2095), .A2(n2517), .ZN(n2578) );
  INV_X1 U2556 ( .A(n2579), .ZN(n2070) );
  NOR2_X1 U2557 ( .A1(n2580), .A2(n2581), .ZN(n2464) );
  INV_X1 U2558 ( .A(n2079), .ZN(n2581) );
  XOR2_X1 U2559 ( .A(n2582), .B(n2583), .Z(n2079) );
  XNOR2_X1 U2560 ( .A(n2584), .B(n2585), .ZN(n2583) );
  AND2_X1 U2561 ( .A1(n2078), .A2(n2077), .ZN(n2580) );
  NAND2_X1 U2562 ( .A1(n2586), .A2(n2579), .ZN(n2049) );
  NOR2_X1 U2563 ( .A1(n2078), .A2(n2077), .ZN(n2579) );
  XNOR2_X1 U2564 ( .A(n2587), .B(n2588), .ZN(n2077) );
  XOR2_X1 U2565 ( .A(n2589), .B(n2590), .Z(n2587) );
  NOR2_X1 U2566 ( .A1(n2026), .A2(n2520), .ZN(n2590) );
  NAND2_X1 U2567 ( .A1(n2591), .A2(n2592), .ZN(n2078) );
  NAND2_X1 U2568 ( .A1(n2582), .A2(n2593), .ZN(n2592) );
  NAND2_X1 U2569 ( .A1(n2585), .A2(n2584), .ZN(n2593) );
  XOR2_X1 U2570 ( .A(n2594), .B(n2595), .Z(n2582) );
  XNOR2_X1 U2571 ( .A(n2596), .B(n2597), .ZN(n2594) );
  OR2_X1 U2572 ( .A1(n2584), .A2(n2585), .ZN(n2591) );
  NOR2_X1 U2573 ( .A1(n2409), .A2(n2026), .ZN(n2585) );
  NAND2_X1 U2574 ( .A1(n2598), .A2(n2599), .ZN(n2584) );
  NAND2_X1 U2575 ( .A1(n2600), .A2(n2095), .ZN(n2599) );
  NOR2_X1 U2576 ( .A1(n2601), .A2(n2409), .ZN(n2600) );
  NOR2_X1 U2577 ( .A1(n2575), .A2(n2577), .ZN(n2601) );
  NAND2_X1 U2578 ( .A1(n2575), .A2(n2577), .ZN(n2598) );
  NAND2_X1 U2579 ( .A1(n2602), .A2(n2603), .ZN(n2577) );
  NAND2_X1 U2580 ( .A1(n2604), .A2(n2101), .ZN(n2603) );
  NOR2_X1 U2581 ( .A1(n2605), .A2(n2409), .ZN(n2604) );
  NOR2_X1 U2582 ( .A1(n2571), .A2(n2573), .ZN(n2605) );
  NAND2_X1 U2583 ( .A1(n2571), .A2(n2573), .ZN(n2602) );
  NAND2_X1 U2584 ( .A1(n2606), .A2(n2607), .ZN(n2573) );
  NAND2_X1 U2585 ( .A1(n2608), .A2(n2459), .ZN(n2607) );
  NOR2_X1 U2586 ( .A1(n2609), .A2(n2409), .ZN(n2608) );
  NOR2_X1 U2587 ( .A1(n2568), .A2(n2570), .ZN(n2609) );
  NAND2_X1 U2588 ( .A1(n2568), .A2(n2570), .ZN(n2606) );
  NAND2_X1 U2589 ( .A1(n2610), .A2(n2611), .ZN(n2570) );
  NAND2_X1 U2590 ( .A1(n2565), .A2(n2612), .ZN(n2611) );
  OR2_X1 U2591 ( .A1(n2566), .A2(n2564), .ZN(n2612) );
  NOR2_X1 U2592 ( .A1(n2370), .A2(n2409), .ZN(n2565) );
  NAND2_X1 U2593 ( .A1(n2564), .A2(n2566), .ZN(n2610) );
  NAND2_X1 U2594 ( .A1(n2613), .A2(n2614), .ZN(n2566) );
  NAND2_X1 U2595 ( .A1(n2562), .A2(n2615), .ZN(n2614) );
  OR2_X1 U2596 ( .A1(n2561), .A2(n2559), .ZN(n2615) );
  NOR2_X1 U2597 ( .A1(n2211), .A2(n2409), .ZN(n2562) );
  NAND2_X1 U2598 ( .A1(n2559), .A2(n2561), .ZN(n2613) );
  NAND2_X1 U2599 ( .A1(n2616), .A2(n2617), .ZN(n2561) );
  NAND2_X1 U2600 ( .A1(n2618), .A2(n2133), .ZN(n2617) );
  NOR2_X1 U2601 ( .A1(n2619), .A2(n2409), .ZN(n2618) );
  NOR2_X1 U2602 ( .A1(n2556), .A2(n2558), .ZN(n2619) );
  NAND2_X1 U2603 ( .A1(n2556), .A2(n2558), .ZN(n2616) );
  NAND2_X1 U2604 ( .A1(n2620), .A2(n2621), .ZN(n2558) );
  NAND2_X1 U2605 ( .A1(n2554), .A2(n2622), .ZN(n2621) );
  OR2_X1 U2606 ( .A1(n2553), .A2(n2551), .ZN(n2622) );
  NOR2_X1 U2607 ( .A1(n2210), .A2(n2409), .ZN(n2554) );
  NAND2_X1 U2608 ( .A1(n2551), .A2(n2553), .ZN(n2620) );
  NAND2_X1 U2609 ( .A1(n2623), .A2(n2624), .ZN(n2553) );
  NAND2_X1 U2610 ( .A1(n2625), .A2(n2149), .ZN(n2624) );
  NOR2_X1 U2611 ( .A1(n2626), .A2(n2409), .ZN(n2625) );
  NOR2_X1 U2612 ( .A1(n2548), .A2(n2550), .ZN(n2626) );
  NAND2_X1 U2613 ( .A1(n2548), .A2(n2550), .ZN(n2623) );
  NAND2_X1 U2614 ( .A1(n2627), .A2(n2628), .ZN(n2550) );
  NAND2_X1 U2615 ( .A1(n2546), .A2(n2629), .ZN(n2628) );
  OR2_X1 U2616 ( .A1(n2545), .A2(n2543), .ZN(n2629) );
  NOR2_X1 U2617 ( .A1(n2209), .A2(n2409), .ZN(n2546) );
  NAND2_X1 U2618 ( .A1(n2543), .A2(n2545), .ZN(n2627) );
  NAND2_X1 U2619 ( .A1(n2630), .A2(n2631), .ZN(n2545) );
  NAND2_X1 U2620 ( .A1(n2632), .A2(n2165), .ZN(n2631) );
  NOR2_X1 U2621 ( .A1(n2633), .A2(n2409), .ZN(n2632) );
  NOR2_X1 U2622 ( .A1(n2540), .A2(n2542), .ZN(n2633) );
  NAND2_X1 U2623 ( .A1(n2540), .A2(n2542), .ZN(n2630) );
  NAND2_X1 U2624 ( .A1(n2634), .A2(n2635), .ZN(n2542) );
  NAND2_X1 U2625 ( .A1(n2538), .A2(n2636), .ZN(n2635) );
  OR2_X1 U2626 ( .A1(n2537), .A2(n2535), .ZN(n2636) );
  NOR2_X1 U2627 ( .A1(n2291), .A2(n2409), .ZN(n2538) );
  NAND2_X1 U2628 ( .A1(n2535), .A2(n2537), .ZN(n2634) );
  NAND2_X1 U2629 ( .A1(n2637), .A2(n2638), .ZN(n2537) );
  NAND2_X1 U2630 ( .A1(n2639), .A2(n2182), .ZN(n2638) );
  NOR2_X1 U2631 ( .A1(n2640), .A2(n2409), .ZN(n2639) );
  NOR2_X1 U2632 ( .A1(n2532), .A2(n2534), .ZN(n2640) );
  NAND2_X1 U2633 ( .A1(n2532), .A2(n2534), .ZN(n2637) );
  NAND2_X1 U2634 ( .A1(n2641), .A2(n2642), .ZN(n2534) );
  NAND2_X1 U2635 ( .A1(n2527), .A2(n2643), .ZN(n2642) );
  NAND2_X1 U2636 ( .A1(n2530), .A2(n2529), .ZN(n2643) );
  NOR2_X1 U2637 ( .A1(n2203), .A2(n2409), .ZN(n2527) );
  OR2_X1 U2638 ( .A1(n2529), .A2(n2530), .ZN(n2641) );
  AND2_X1 U2639 ( .A1(n2644), .A2(n2645), .ZN(n2530) );
  NAND2_X1 U2640 ( .A1(n2521), .A2(n2646), .ZN(n2645) );
  NAND2_X1 U2641 ( .A1(n1953), .A2(n2647), .ZN(n2646) );
  NAND2_X1 U2642 ( .A1(n2648), .A2(n1956), .ZN(n2647) );
  NAND2_X1 U2643 ( .A1(n2649), .A2(n2650), .ZN(n2644) );
  NAND2_X1 U2644 ( .A1(n1959), .A2(n2651), .ZN(n2650) );
  NAND2_X1 U2645 ( .A1(n1961), .A2(n2520), .ZN(n2651) );
  NAND2_X1 U2646 ( .A1(n2652), .A2(n2653), .ZN(n2529) );
  INV_X1 U2647 ( .A(n2306), .ZN(n2653) );
  NOR2_X1 U2648 ( .A1(n2520), .A2(n2409), .ZN(n2652) );
  INV_X1 U2649 ( .A(n2517), .ZN(n2409) );
  XOR2_X1 U2650 ( .A(n2654), .B(n2655), .Z(n2517) );
  XOR2_X1 U2651 ( .A(d_11_), .B(c_11_), .Z(n2655) );
  XNOR2_X1 U2652 ( .A(n2656), .B(n2657), .ZN(n2532) );
  XNOR2_X1 U2653 ( .A(n2658), .B(n2659), .ZN(n2657) );
  XOR2_X1 U2654 ( .A(n2660), .B(n2661), .Z(n2535) );
  XNOR2_X1 U2655 ( .A(n2662), .B(n2663), .ZN(n2660) );
  NAND2_X1 U2656 ( .A1(n2182), .A2(n2521), .ZN(n2662) );
  XOR2_X1 U2657 ( .A(n2664), .B(n2665), .Z(n2540) );
  XOR2_X1 U2658 ( .A(n2666), .B(n2667), .Z(n2664) );
  XOR2_X1 U2659 ( .A(n2668), .B(n2669), .Z(n2543) );
  XOR2_X1 U2660 ( .A(n2670), .B(n2671), .Z(n2668) );
  NOR2_X1 U2661 ( .A1(n2520), .A2(n2394), .ZN(n2671) );
  XOR2_X1 U2662 ( .A(n2672), .B(n2673), .Z(n2548) );
  XOR2_X1 U2663 ( .A(n2674), .B(n2675), .Z(n2672) );
  XOR2_X1 U2664 ( .A(n2676), .B(n2677), .Z(n2551) );
  XOR2_X1 U2665 ( .A(n2678), .B(n2679), .Z(n2676) );
  NOR2_X1 U2666 ( .A1(n2520), .A2(n2386), .ZN(n2679) );
  XNOR2_X1 U2667 ( .A(n2680), .B(n2681), .ZN(n2556) );
  XNOR2_X1 U2668 ( .A(n2682), .B(n2683), .ZN(n2681) );
  XOR2_X1 U2669 ( .A(n2684), .B(n2685), .Z(n2559) );
  XOR2_X1 U2670 ( .A(n2686), .B(n2687), .Z(n2684) );
  NOR2_X1 U2671 ( .A1(n2520), .A2(n2378), .ZN(n2687) );
  XNOR2_X1 U2672 ( .A(n2688), .B(n2689), .ZN(n2564) );
  XOR2_X1 U2673 ( .A(n2690), .B(n2691), .Z(n2689) );
  NAND2_X1 U2674 ( .A1(n2521), .A2(n2692), .ZN(n2691) );
  XNOR2_X1 U2675 ( .A(n2693), .B(n2694), .ZN(n2568) );
  XNOR2_X1 U2676 ( .A(n2695), .B(n2696), .ZN(n2694) );
  XNOR2_X1 U2677 ( .A(n2697), .B(n2698), .ZN(n2571) );
  XNOR2_X1 U2678 ( .A(n2699), .B(n2700), .ZN(n2697) );
  XNOR2_X1 U2679 ( .A(n2701), .B(n2702), .ZN(n2575) );
  XNOR2_X1 U2680 ( .A(n2703), .B(n2704), .ZN(n2701) );
  XOR2_X1 U2681 ( .A(n2072), .B(n2705), .Z(n2586) );
  NAND2_X1 U2682 ( .A1(n2706), .A2(n2707), .ZN(n1921) );
  OR2_X1 U2683 ( .A1(n2072), .A2(n2705), .ZN(n2707) );
  XOR2_X1 U2684 ( .A(n2708), .B(n2709), .Z(n2706) );
  NAND2_X1 U2685 ( .A1(n2710), .A2(n2711), .ZN(n1922) );
  XOR2_X1 U2686 ( .A(n2712), .B(n2709), .Z(n2711) );
  NOR2_X1 U2687 ( .A1(n2705), .A2(n2072), .ZN(n2710) );
  XNOR2_X1 U2688 ( .A(n2713), .B(n2714), .ZN(n2072) );
  XOR2_X1 U2689 ( .A(n2715), .B(n2716), .Z(n2713) );
  NOR2_X1 U2690 ( .A1(n2026), .A2(n2648), .ZN(n2716) );
  INV_X1 U2691 ( .A(n2071), .ZN(n2705) );
  NAND2_X1 U2692 ( .A1(n2717), .A2(n2718), .ZN(n2071) );
  NAND2_X1 U2693 ( .A1(n2719), .A2(n2521), .ZN(n2718) );
  NOR2_X1 U2694 ( .A1(n2720), .A2(n2026), .ZN(n2719) );
  NOR2_X1 U2695 ( .A1(n2589), .A2(n2588), .ZN(n2720) );
  NAND2_X1 U2696 ( .A1(n2588), .A2(n2589), .ZN(n2717) );
  NAND2_X1 U2697 ( .A1(n2721), .A2(n2722), .ZN(n2589) );
  NAND2_X1 U2698 ( .A1(n2597), .A2(n2723), .ZN(n2722) );
  NAND2_X1 U2699 ( .A1(n2596), .A2(n2595), .ZN(n2723) );
  NOR2_X1 U2700 ( .A1(n2241), .A2(n2520), .ZN(n2597) );
  OR2_X1 U2701 ( .A1(n2595), .A2(n2596), .ZN(n2721) );
  AND2_X1 U2702 ( .A1(n2724), .A2(n2725), .ZN(n2596) );
  NAND2_X1 U2703 ( .A1(n2703), .A2(n2726), .ZN(n2725) );
  NAND2_X1 U2704 ( .A1(n2704), .A2(n2702), .ZN(n2726) );
  NOR2_X1 U2705 ( .A1(n2362), .A2(n2520), .ZN(n2703) );
  OR2_X1 U2706 ( .A1(n2702), .A2(n2704), .ZN(n2724) );
  AND2_X1 U2707 ( .A1(n2727), .A2(n2728), .ZN(n2704) );
  NAND2_X1 U2708 ( .A1(n2700), .A2(n2729), .ZN(n2728) );
  NAND2_X1 U2709 ( .A1(n2699), .A2(n2698), .ZN(n2729) );
  NOR2_X1 U2710 ( .A1(n2212), .A2(n2520), .ZN(n2700) );
  OR2_X1 U2711 ( .A1(n2698), .A2(n2699), .ZN(n2727) );
  AND2_X1 U2712 ( .A1(n2730), .A2(n2731), .ZN(n2699) );
  NAND2_X1 U2713 ( .A1(n2696), .A2(n2732), .ZN(n2731) );
  OR2_X1 U2714 ( .A1(n2695), .A2(n2693), .ZN(n2732) );
  NOR2_X1 U2715 ( .A1(n2520), .A2(n2370), .ZN(n2696) );
  NAND2_X1 U2716 ( .A1(n2693), .A2(n2695), .ZN(n2730) );
  NAND2_X1 U2717 ( .A1(n2733), .A2(n2734), .ZN(n2695) );
  NAND2_X1 U2718 ( .A1(n2735), .A2(n2521), .ZN(n2734) );
  NOR2_X1 U2719 ( .A1(n2736), .A2(n2211), .ZN(n2735) );
  NOR2_X1 U2720 ( .A1(n2688), .A2(n2690), .ZN(n2736) );
  NAND2_X1 U2721 ( .A1(n2688), .A2(n2690), .ZN(n2733) );
  NAND2_X1 U2722 ( .A1(n2737), .A2(n2738), .ZN(n2690) );
  NAND2_X1 U2723 ( .A1(n2739), .A2(n2133), .ZN(n2738) );
  NOR2_X1 U2724 ( .A1(n2740), .A2(n2520), .ZN(n2739) );
  NOR2_X1 U2725 ( .A1(n2685), .A2(n2686), .ZN(n2740) );
  NAND2_X1 U2726 ( .A1(n2685), .A2(n2686), .ZN(n2737) );
  NAND2_X1 U2727 ( .A1(n2741), .A2(n2742), .ZN(n2686) );
  NAND2_X1 U2728 ( .A1(n2683), .A2(n2743), .ZN(n2742) );
  OR2_X1 U2729 ( .A1(n2680), .A2(n2682), .ZN(n2743) );
  NOR2_X1 U2730 ( .A1(n2520), .A2(n2210), .ZN(n2683) );
  NAND2_X1 U2731 ( .A1(n2680), .A2(n2682), .ZN(n2741) );
  NAND2_X1 U2732 ( .A1(n2744), .A2(n2745), .ZN(n2682) );
  NAND2_X1 U2733 ( .A1(n2746), .A2(n2149), .ZN(n2745) );
  NOR2_X1 U2734 ( .A1(n2747), .A2(n2520), .ZN(n2746) );
  NOR2_X1 U2735 ( .A1(n2677), .A2(n2678), .ZN(n2747) );
  NAND2_X1 U2736 ( .A1(n2677), .A2(n2678), .ZN(n2744) );
  NAND2_X1 U2737 ( .A1(n2748), .A2(n2749), .ZN(n2678) );
  NAND2_X1 U2738 ( .A1(n2675), .A2(n2750), .ZN(n2749) );
  OR2_X1 U2739 ( .A1(n2673), .A2(n2674), .ZN(n2750) );
  NOR2_X1 U2740 ( .A1(n2520), .A2(n2209), .ZN(n2675) );
  NAND2_X1 U2741 ( .A1(n2673), .A2(n2674), .ZN(n2748) );
  NAND2_X1 U2742 ( .A1(n2751), .A2(n2752), .ZN(n2674) );
  NAND2_X1 U2743 ( .A1(n2753), .A2(n2165), .ZN(n2752) );
  NOR2_X1 U2744 ( .A1(n2754), .A2(n2520), .ZN(n2753) );
  NOR2_X1 U2745 ( .A1(n2669), .A2(n2670), .ZN(n2754) );
  NAND2_X1 U2746 ( .A1(n2669), .A2(n2670), .ZN(n2751) );
  NAND2_X1 U2747 ( .A1(n2755), .A2(n2756), .ZN(n2670) );
  NAND2_X1 U2748 ( .A1(n2667), .A2(n2757), .ZN(n2756) );
  OR2_X1 U2749 ( .A1(n2665), .A2(n2666), .ZN(n2757) );
  NOR2_X1 U2750 ( .A1(n2520), .A2(n2291), .ZN(n2667) );
  NAND2_X1 U2751 ( .A1(n2665), .A2(n2666), .ZN(n2755) );
  NAND2_X1 U2752 ( .A1(n2758), .A2(n2759), .ZN(n2666) );
  NAND2_X1 U2753 ( .A1(n2760), .A2(n2182), .ZN(n2759) );
  NOR2_X1 U2754 ( .A1(n2761), .A2(n2520), .ZN(n2760) );
  NOR2_X1 U2755 ( .A1(n2661), .A2(n2663), .ZN(n2761) );
  NAND2_X1 U2756 ( .A1(n2661), .A2(n2663), .ZN(n2758) );
  NAND2_X1 U2757 ( .A1(n2762), .A2(n2763), .ZN(n2663) );
  NAND2_X1 U2758 ( .A1(n2656), .A2(n2764), .ZN(n2763) );
  NAND2_X1 U2759 ( .A1(n2659), .A2(n2658), .ZN(n2764) );
  NOR2_X1 U2760 ( .A1(n2520), .A2(n2203), .ZN(n2656) );
  OR2_X1 U2761 ( .A1(n2658), .A2(n2659), .ZN(n2762) );
  AND2_X1 U2762 ( .A1(n2765), .A2(n2766), .ZN(n2659) );
  NAND2_X1 U2763 ( .A1(n2649), .A2(n2767), .ZN(n2766) );
  NAND2_X1 U2764 ( .A1(n1953), .A2(n2768), .ZN(n2767) );
  NAND2_X1 U2765 ( .A1(n2769), .A2(n1956), .ZN(n2768) );
  NAND2_X1 U2766 ( .A1(n2770), .A2(n2771), .ZN(n2765) );
  NAND2_X1 U2767 ( .A1(n1959), .A2(n2772), .ZN(n2771) );
  NAND2_X1 U2768 ( .A1(n1961), .A2(n2648), .ZN(n2772) );
  NAND2_X1 U2769 ( .A1(n2773), .A2(n2649), .ZN(n2658) );
  NOR2_X1 U2770 ( .A1(n2306), .A2(n2520), .ZN(n2773) );
  INV_X1 U2771 ( .A(n2521), .ZN(n2520) );
  XOR2_X1 U2772 ( .A(n2774), .B(n2775), .Z(n2521) );
  XOR2_X1 U2773 ( .A(d_10_), .B(c_10_), .Z(n2775) );
  XNOR2_X1 U2774 ( .A(n2776), .B(n2777), .ZN(n2661) );
  XNOR2_X1 U2775 ( .A(n2778), .B(n2779), .ZN(n2777) );
  XOR2_X1 U2776 ( .A(n2780), .B(n2781), .Z(n2665) );
  XNOR2_X1 U2777 ( .A(n2782), .B(n2783), .ZN(n2780) );
  NAND2_X1 U2778 ( .A1(n2182), .A2(n2649), .ZN(n2782) );
  XNOR2_X1 U2779 ( .A(n2784), .B(n2785), .ZN(n2669) );
  XNOR2_X1 U2780 ( .A(n2786), .B(n2787), .ZN(n2785) );
  XOR2_X1 U2781 ( .A(n2788), .B(n2789), .Z(n2673) );
  XOR2_X1 U2782 ( .A(n2790), .B(n2791), .Z(n2788) );
  NOR2_X1 U2783 ( .A1(n2648), .A2(n2394), .ZN(n2791) );
  XNOR2_X1 U2784 ( .A(n2792), .B(n2793), .ZN(n2677) );
  XNOR2_X1 U2785 ( .A(n2794), .B(n2795), .ZN(n2793) );
  XOR2_X1 U2786 ( .A(n2796), .B(n2797), .Z(n2680) );
  XOR2_X1 U2787 ( .A(n2798), .B(n2799), .Z(n2796) );
  NOR2_X1 U2788 ( .A1(n2648), .A2(n2386), .ZN(n2799) );
  XNOR2_X1 U2789 ( .A(n2800), .B(n2801), .ZN(n2685) );
  XNOR2_X1 U2790 ( .A(n2802), .B(n2803), .ZN(n2801) );
  XOR2_X1 U2791 ( .A(n2804), .B(n2805), .Z(n2688) );
  XOR2_X1 U2792 ( .A(n2806), .B(n2807), .Z(n2804) );
  XOR2_X1 U2793 ( .A(n2808), .B(n2809), .Z(n2693) );
  XOR2_X1 U2794 ( .A(n2810), .B(n2811), .Z(n2808) );
  NOR2_X1 U2795 ( .A1(n2211), .A2(n2648), .ZN(n2811) );
  XOR2_X1 U2796 ( .A(n2812), .B(n2813), .Z(n2698) );
  XOR2_X1 U2797 ( .A(n2814), .B(n2815), .Z(n2813) );
  NAND2_X1 U2798 ( .A1(n2649), .A2(n2117), .ZN(n2815) );
  XOR2_X1 U2799 ( .A(n2816), .B(n2817), .Z(n2702) );
  XOR2_X1 U2800 ( .A(n2818), .B(n2819), .Z(n2817) );
  NAND2_X1 U2801 ( .A1(n2459), .A2(n2649), .ZN(n2819) );
  XOR2_X1 U2802 ( .A(n2820), .B(n2821), .Z(n2595) );
  XOR2_X1 U2803 ( .A(n2822), .B(n2823), .Z(n2821) );
  NAND2_X1 U2804 ( .A1(n1917), .A2(n2649), .ZN(n2823) );
  XOR2_X1 U2805 ( .A(n2824), .B(n2825), .Z(n2588) );
  XOR2_X1 U2806 ( .A(n2826), .B(n2827), .Z(n2824) );
  NOR2_X1 U2807 ( .A1(n2648), .A2(n2241), .ZN(n2827) );
  NAND2_X1 U2808 ( .A1(n2828), .A2(n2829), .ZN(n1925) );
  NAND2_X1 U2809 ( .A1(n2709), .A2(n2712), .ZN(n2829) );
  NAND2_X1 U2810 ( .A1(n2830), .A2(n2709), .ZN(n1926) );
  XNOR2_X1 U2811 ( .A(n2831), .B(n2832), .ZN(n2709) );
  XNOR2_X1 U2812 ( .A(n2833), .B(n2834), .ZN(n2832) );
  NOR2_X1 U2813 ( .A1(n2708), .A2(n2828), .ZN(n2830) );
  XOR2_X1 U2814 ( .A(n2835), .B(n2836), .Z(n2828) );
  INV_X1 U2815 ( .A(n2712), .ZN(n2708) );
  NAND2_X1 U2816 ( .A1(n2837), .A2(n2838), .ZN(n2712) );
  NAND2_X1 U2817 ( .A1(n2839), .A2(n2649), .ZN(n2838) );
  NOR2_X1 U2818 ( .A1(n2840), .A2(n2026), .ZN(n2839) );
  NOR2_X1 U2819 ( .A1(n2714), .A2(n2715), .ZN(n2840) );
  NAND2_X1 U2820 ( .A1(n2714), .A2(n2715), .ZN(n2837) );
  NAND2_X1 U2821 ( .A1(n2841), .A2(n2842), .ZN(n2715) );
  NAND2_X1 U2822 ( .A1(n2843), .A2(n2095), .ZN(n2842) );
  NOR2_X1 U2823 ( .A1(n2844), .A2(n2648), .ZN(n2843) );
  NOR2_X1 U2824 ( .A1(n2825), .A2(n2826), .ZN(n2844) );
  NAND2_X1 U2825 ( .A1(n2825), .A2(n2826), .ZN(n2841) );
  NAND2_X1 U2826 ( .A1(n2845), .A2(n2846), .ZN(n2826) );
  NAND2_X1 U2827 ( .A1(n2847), .A2(n2101), .ZN(n2846) );
  NOR2_X1 U2828 ( .A1(n2848), .A2(n2648), .ZN(n2847) );
  NOR2_X1 U2829 ( .A1(n2822), .A2(n2820), .ZN(n2848) );
  NAND2_X1 U2830 ( .A1(n2820), .A2(n2822), .ZN(n2845) );
  NAND2_X1 U2831 ( .A1(n2849), .A2(n2850), .ZN(n2822) );
  NAND2_X1 U2832 ( .A1(n2851), .A2(n2459), .ZN(n2850) );
  NOR2_X1 U2833 ( .A1(n2852), .A2(n2648), .ZN(n2851) );
  NOR2_X1 U2834 ( .A1(n2818), .A2(n2816), .ZN(n2852) );
  NAND2_X1 U2835 ( .A1(n2816), .A2(n2818), .ZN(n2849) );
  NAND2_X1 U2836 ( .A1(n2853), .A2(n2854), .ZN(n2818) );
  NAND2_X1 U2837 ( .A1(n2855), .A2(n2649), .ZN(n2854) );
  NOR2_X1 U2838 ( .A1(n2856), .A2(n2370), .ZN(n2855) );
  NOR2_X1 U2839 ( .A1(n2814), .A2(n2812), .ZN(n2856) );
  NAND2_X1 U2840 ( .A1(n2812), .A2(n2814), .ZN(n2853) );
  NAND2_X1 U2841 ( .A1(n2857), .A2(n2858), .ZN(n2814) );
  NAND2_X1 U2842 ( .A1(n2859), .A2(n2649), .ZN(n2858) );
  NOR2_X1 U2843 ( .A1(n2860), .A2(n2211), .ZN(n2859) );
  NOR2_X1 U2844 ( .A1(n2810), .A2(n2809), .ZN(n2860) );
  NAND2_X1 U2845 ( .A1(n2809), .A2(n2810), .ZN(n2857) );
  NAND2_X1 U2846 ( .A1(n2861), .A2(n2862), .ZN(n2810) );
  NAND2_X1 U2847 ( .A1(n2807), .A2(n2863), .ZN(n2862) );
  OR2_X1 U2848 ( .A1(n2805), .A2(n2806), .ZN(n2863) );
  NOR2_X1 U2849 ( .A1(n2378), .A2(n2648), .ZN(n2807) );
  NAND2_X1 U2850 ( .A1(n2805), .A2(n2806), .ZN(n2861) );
  NAND2_X1 U2851 ( .A1(n2864), .A2(n2865), .ZN(n2806) );
  NAND2_X1 U2852 ( .A1(n2803), .A2(n2866), .ZN(n2865) );
  OR2_X1 U2853 ( .A1(n2800), .A2(n2802), .ZN(n2866) );
  NOR2_X1 U2854 ( .A1(n2648), .A2(n2210), .ZN(n2803) );
  NAND2_X1 U2855 ( .A1(n2800), .A2(n2802), .ZN(n2864) );
  NAND2_X1 U2856 ( .A1(n2867), .A2(n2868), .ZN(n2802) );
  NAND2_X1 U2857 ( .A1(n2869), .A2(n2149), .ZN(n2868) );
  NOR2_X1 U2858 ( .A1(n2870), .A2(n2648), .ZN(n2869) );
  NOR2_X1 U2859 ( .A1(n2797), .A2(n2798), .ZN(n2870) );
  NAND2_X1 U2860 ( .A1(n2797), .A2(n2798), .ZN(n2867) );
  NAND2_X1 U2861 ( .A1(n2871), .A2(n2872), .ZN(n2798) );
  NAND2_X1 U2862 ( .A1(n2795), .A2(n2873), .ZN(n2872) );
  OR2_X1 U2863 ( .A1(n2792), .A2(n2794), .ZN(n2873) );
  NOR2_X1 U2864 ( .A1(n2648), .A2(n2209), .ZN(n2795) );
  NAND2_X1 U2865 ( .A1(n2792), .A2(n2794), .ZN(n2871) );
  NAND2_X1 U2866 ( .A1(n2874), .A2(n2875), .ZN(n2794) );
  NAND2_X1 U2867 ( .A1(n2876), .A2(n2165), .ZN(n2875) );
  NOR2_X1 U2868 ( .A1(n2877), .A2(n2648), .ZN(n2876) );
  NOR2_X1 U2869 ( .A1(n2789), .A2(n2790), .ZN(n2877) );
  NAND2_X1 U2870 ( .A1(n2789), .A2(n2790), .ZN(n2874) );
  NAND2_X1 U2871 ( .A1(n2878), .A2(n2879), .ZN(n2790) );
  NAND2_X1 U2872 ( .A1(n2787), .A2(n2880), .ZN(n2879) );
  OR2_X1 U2873 ( .A1(n2784), .A2(n2786), .ZN(n2880) );
  NOR2_X1 U2874 ( .A1(n2648), .A2(n2291), .ZN(n2787) );
  NAND2_X1 U2875 ( .A1(n2784), .A2(n2786), .ZN(n2878) );
  NAND2_X1 U2876 ( .A1(n2881), .A2(n2882), .ZN(n2786) );
  NAND2_X1 U2877 ( .A1(n2883), .A2(n2182), .ZN(n2882) );
  NOR2_X1 U2878 ( .A1(n2884), .A2(n2648), .ZN(n2883) );
  NOR2_X1 U2879 ( .A1(n2781), .A2(n2783), .ZN(n2884) );
  NAND2_X1 U2880 ( .A1(n2781), .A2(n2783), .ZN(n2881) );
  NAND2_X1 U2881 ( .A1(n2885), .A2(n2886), .ZN(n2783) );
  NAND2_X1 U2882 ( .A1(n2776), .A2(n2887), .ZN(n2886) );
  NAND2_X1 U2883 ( .A1(n2779), .A2(n2778), .ZN(n2887) );
  NOR2_X1 U2884 ( .A1(n2648), .A2(n2203), .ZN(n2776) );
  OR2_X1 U2885 ( .A1(n2778), .A2(n2779), .ZN(n2885) );
  AND2_X1 U2886 ( .A1(n2888), .A2(n2889), .ZN(n2779) );
  NAND2_X1 U2887 ( .A1(n2770), .A2(n2890), .ZN(n2889) );
  NAND2_X1 U2888 ( .A1(n1953), .A2(n2891), .ZN(n2890) );
  NAND2_X1 U2889 ( .A1(n2892), .A2(n1956), .ZN(n2891) );
  NAND2_X1 U2890 ( .A1(n2893), .A2(n2894), .ZN(n2888) );
  NAND2_X1 U2891 ( .A1(n1959), .A2(n2895), .ZN(n2894) );
  NAND2_X1 U2892 ( .A1(n1961), .A2(n2769), .ZN(n2895) );
  NAND2_X1 U2893 ( .A1(n2896), .A2(n2770), .ZN(n2778) );
  NOR2_X1 U2894 ( .A1(n2306), .A2(n2648), .ZN(n2896) );
  INV_X1 U2895 ( .A(n2649), .ZN(n2648) );
  XOR2_X1 U2896 ( .A(n2897), .B(n2898), .Z(n2649) );
  XOR2_X1 U2897 ( .A(d_9_), .B(c_9_), .Z(n2898) );
  XNOR2_X1 U2898 ( .A(n2899), .B(n2900), .ZN(n2781) );
  XNOR2_X1 U2899 ( .A(n2901), .B(n2902), .ZN(n2900) );
  XOR2_X1 U2900 ( .A(n2903), .B(n2904), .Z(n2784) );
  XNOR2_X1 U2901 ( .A(n2905), .B(n2906), .ZN(n2903) );
  NAND2_X1 U2902 ( .A1(n2182), .A2(n2770), .ZN(n2905) );
  XOR2_X1 U2903 ( .A(n2907), .B(n2908), .Z(n2789) );
  XOR2_X1 U2904 ( .A(n2909), .B(n2910), .Z(n2907) );
  XOR2_X1 U2905 ( .A(n2911), .B(n2912), .Z(n2792) );
  XOR2_X1 U2906 ( .A(n2913), .B(n2914), .Z(n2911) );
  NOR2_X1 U2907 ( .A1(n2769), .A2(n2394), .ZN(n2914) );
  XNOR2_X1 U2908 ( .A(n2915), .B(n2916), .ZN(n2797) );
  XNOR2_X1 U2909 ( .A(n2917), .B(n2918), .ZN(n2916) );
  XOR2_X1 U2910 ( .A(n2919), .B(n2920), .Z(n2800) );
  XOR2_X1 U2911 ( .A(n2921), .B(n2922), .Z(n2919) );
  NOR2_X1 U2912 ( .A1(n2769), .A2(n2386), .ZN(n2922) );
  XNOR2_X1 U2913 ( .A(n2923), .B(n2924), .ZN(n2805) );
  XOR2_X1 U2914 ( .A(n2925), .B(n2926), .Z(n2924) );
  NAND2_X1 U2915 ( .A1(n2770), .A2(n2927), .ZN(n2926) );
  XNOR2_X1 U2916 ( .A(n2928), .B(n2929), .ZN(n2809) );
  XNOR2_X1 U2917 ( .A(n2930), .B(n2931), .ZN(n2929) );
  XNOR2_X1 U2918 ( .A(n2932), .B(n2933), .ZN(n2812) );
  XNOR2_X1 U2919 ( .A(n2934), .B(n2935), .ZN(n2932) );
  XNOR2_X1 U2920 ( .A(n2936), .B(n2937), .ZN(n2816) );
  XNOR2_X1 U2921 ( .A(n2938), .B(n2939), .ZN(n2936) );
  XNOR2_X1 U2922 ( .A(n2940), .B(n2941), .ZN(n2820) );
  XNOR2_X1 U2923 ( .A(n2942), .B(n2943), .ZN(n2941) );
  XOR2_X1 U2924 ( .A(n2944), .B(n2945), .Z(n2825) );
  XOR2_X1 U2925 ( .A(n2946), .B(n2947), .Z(n2944) );
  NOR2_X1 U2926 ( .A1(n2769), .A2(n2362), .ZN(n2947) );
  XNOR2_X1 U2927 ( .A(n2948), .B(n2949), .ZN(n2714) );
  XOR2_X1 U2928 ( .A(n2950), .B(n2951), .Z(n2949) );
  NAND2_X1 U2929 ( .A1(n2095), .A2(n2770), .ZN(n2951) );
  NAND2_X1 U2930 ( .A1(n2952), .A2(n2953), .ZN(n1929) );
  NAND2_X1 U2931 ( .A1(n2835), .A2(n2954), .ZN(n2953) );
  NAND2_X1 U2932 ( .A1(n2955), .A2(n2835), .ZN(n1930) );
  XOR2_X1 U2933 ( .A(n2956), .B(n2957), .Z(n2835) );
  XOR2_X1 U2934 ( .A(n2958), .B(n2959), .Z(n2956) );
  NOR2_X1 U2935 ( .A1(n2026), .A2(n2892), .ZN(n2959) );
  NOR2_X1 U2936 ( .A1(n2836), .A2(n2952), .ZN(n2955) );
  XNOR2_X1 U2937 ( .A(n2960), .B(n2961), .ZN(n2952) );
  INV_X1 U2938 ( .A(n2954), .ZN(n2836) );
  NAND2_X1 U2939 ( .A1(n2962), .A2(n2963), .ZN(n2954) );
  NAND2_X1 U2940 ( .A1(n2834), .A2(n2964), .ZN(n2963) );
  OR2_X1 U2941 ( .A1(n2831), .A2(n2833), .ZN(n2964) );
  NOR2_X1 U2942 ( .A1(n2769), .A2(n2026), .ZN(n2834) );
  NAND2_X1 U2943 ( .A1(n2831), .A2(n2833), .ZN(n2962) );
  NAND2_X1 U2944 ( .A1(n2965), .A2(n2966), .ZN(n2833) );
  NAND2_X1 U2945 ( .A1(n2967), .A2(n2095), .ZN(n2966) );
  NOR2_X1 U2946 ( .A1(n2968), .A2(n2769), .ZN(n2967) );
  NOR2_X1 U2947 ( .A1(n2950), .A2(n2948), .ZN(n2968) );
  NAND2_X1 U2948 ( .A1(n2948), .A2(n2950), .ZN(n2965) );
  NAND2_X1 U2949 ( .A1(n2969), .A2(n2970), .ZN(n2950) );
  NAND2_X1 U2950 ( .A1(n2971), .A2(n2101), .ZN(n2970) );
  NOR2_X1 U2951 ( .A1(n2972), .A2(n2769), .ZN(n2971) );
  NOR2_X1 U2952 ( .A1(n2946), .A2(n2945), .ZN(n2972) );
  NAND2_X1 U2953 ( .A1(n2945), .A2(n2946), .ZN(n2969) );
  NAND2_X1 U2954 ( .A1(n2973), .A2(n2974), .ZN(n2946) );
  NAND2_X1 U2955 ( .A1(n2943), .A2(n2975), .ZN(n2974) );
  OR2_X1 U2956 ( .A1(n2942), .A2(n2940), .ZN(n2975) );
  NOR2_X1 U2957 ( .A1(n2212), .A2(n2769), .ZN(n2943) );
  NAND2_X1 U2958 ( .A1(n2940), .A2(n2942), .ZN(n2973) );
  NAND2_X1 U2959 ( .A1(n2976), .A2(n2977), .ZN(n2942) );
  NAND2_X1 U2960 ( .A1(n2938), .A2(n2978), .ZN(n2977) );
  NAND2_X1 U2961 ( .A1(n2939), .A2(n2937), .ZN(n2978) );
  NOR2_X1 U2962 ( .A1(n2769), .A2(n2370), .ZN(n2938) );
  OR2_X1 U2963 ( .A1(n2937), .A2(n2939), .ZN(n2976) );
  AND2_X1 U2964 ( .A1(n2979), .A2(n2980), .ZN(n2939) );
  NAND2_X1 U2965 ( .A1(n2935), .A2(n2981), .ZN(n2980) );
  NAND2_X1 U2966 ( .A1(n2934), .A2(n2933), .ZN(n2981) );
  NOR2_X1 U2967 ( .A1(n2769), .A2(n2211), .ZN(n2935) );
  OR2_X1 U2968 ( .A1(n2933), .A2(n2934), .ZN(n2979) );
  AND2_X1 U2969 ( .A1(n2982), .A2(n2983), .ZN(n2934) );
  NAND2_X1 U2970 ( .A1(n2931), .A2(n2984), .ZN(n2983) );
  OR2_X1 U2971 ( .A1(n2930), .A2(n2928), .ZN(n2984) );
  NOR2_X1 U2972 ( .A1(n2378), .A2(n2769), .ZN(n2931) );
  NAND2_X1 U2973 ( .A1(n2928), .A2(n2930), .ZN(n2982) );
  NAND2_X1 U2974 ( .A1(n2985), .A2(n2986), .ZN(n2930) );
  NAND2_X1 U2975 ( .A1(n2987), .A2(n2770), .ZN(n2986) );
  NOR2_X1 U2976 ( .A1(n2988), .A2(n2210), .ZN(n2987) );
  NOR2_X1 U2977 ( .A1(n2923), .A2(n2925), .ZN(n2988) );
  NAND2_X1 U2978 ( .A1(n2923), .A2(n2925), .ZN(n2985) );
  NAND2_X1 U2979 ( .A1(n2989), .A2(n2990), .ZN(n2925) );
  NAND2_X1 U2980 ( .A1(n2991), .A2(n2149), .ZN(n2990) );
  NOR2_X1 U2981 ( .A1(n2992), .A2(n2769), .ZN(n2991) );
  NOR2_X1 U2982 ( .A1(n2920), .A2(n2921), .ZN(n2992) );
  NAND2_X1 U2983 ( .A1(n2920), .A2(n2921), .ZN(n2989) );
  NAND2_X1 U2984 ( .A1(n2993), .A2(n2994), .ZN(n2921) );
  NAND2_X1 U2985 ( .A1(n2918), .A2(n2995), .ZN(n2994) );
  OR2_X1 U2986 ( .A1(n2915), .A2(n2917), .ZN(n2995) );
  NOR2_X1 U2987 ( .A1(n2769), .A2(n2209), .ZN(n2918) );
  NAND2_X1 U2988 ( .A1(n2915), .A2(n2917), .ZN(n2993) );
  NAND2_X1 U2989 ( .A1(n2996), .A2(n2997), .ZN(n2917) );
  NAND2_X1 U2990 ( .A1(n2998), .A2(n2165), .ZN(n2997) );
  NOR2_X1 U2991 ( .A1(n2999), .A2(n2769), .ZN(n2998) );
  NOR2_X1 U2992 ( .A1(n2912), .A2(n2913), .ZN(n2999) );
  NAND2_X1 U2993 ( .A1(n2912), .A2(n2913), .ZN(n2996) );
  NAND2_X1 U2994 ( .A1(n3000), .A2(n3001), .ZN(n2913) );
  NAND2_X1 U2995 ( .A1(n2910), .A2(n3002), .ZN(n3001) );
  OR2_X1 U2996 ( .A1(n2908), .A2(n2909), .ZN(n3002) );
  NOR2_X1 U2997 ( .A1(n2769), .A2(n2291), .ZN(n2910) );
  NAND2_X1 U2998 ( .A1(n2908), .A2(n2909), .ZN(n3000) );
  NAND2_X1 U2999 ( .A1(n3003), .A2(n3004), .ZN(n2909) );
  NAND2_X1 U3000 ( .A1(n3005), .A2(n2182), .ZN(n3004) );
  NOR2_X1 U3001 ( .A1(n3006), .A2(n2769), .ZN(n3005) );
  NOR2_X1 U3002 ( .A1(n2904), .A2(n2906), .ZN(n3006) );
  NAND2_X1 U3003 ( .A1(n2904), .A2(n2906), .ZN(n3003) );
  NAND2_X1 U3004 ( .A1(n3007), .A2(n3008), .ZN(n2906) );
  NAND2_X1 U3005 ( .A1(n2899), .A2(n3009), .ZN(n3008) );
  NAND2_X1 U3006 ( .A1(n2902), .A2(n2901), .ZN(n3009) );
  NOR2_X1 U3007 ( .A1(n2769), .A2(n2203), .ZN(n2899) );
  OR2_X1 U3008 ( .A1(n2901), .A2(n2902), .ZN(n3007) );
  AND2_X1 U3009 ( .A1(n3010), .A2(n3011), .ZN(n2902) );
  NAND2_X1 U3010 ( .A1(n2893), .A2(n3012), .ZN(n3011) );
  NAND2_X1 U3011 ( .A1(n1953), .A2(n3013), .ZN(n3012) );
  NAND2_X1 U3012 ( .A1(n3014), .A2(n1956), .ZN(n3013) );
  NAND2_X1 U3013 ( .A1(n3015), .A2(n3016), .ZN(n3010) );
  NAND2_X1 U3014 ( .A1(n1959), .A2(n3017), .ZN(n3016) );
  NAND2_X1 U3015 ( .A1(n1961), .A2(n2892), .ZN(n3017) );
  NAND2_X1 U3016 ( .A1(n3018), .A2(n2893), .ZN(n2901) );
  NOR2_X1 U3017 ( .A1(n2306), .A2(n2769), .ZN(n3018) );
  INV_X1 U3018 ( .A(n2770), .ZN(n2769) );
  XOR2_X1 U3019 ( .A(n3019), .B(n3020), .Z(n2770) );
  XOR2_X1 U3020 ( .A(d_8_), .B(c_8_), .Z(n3020) );
  XNOR2_X1 U3021 ( .A(n3021), .B(n3022), .ZN(n2904) );
  XNOR2_X1 U3022 ( .A(n3023), .B(n3024), .ZN(n3022) );
  XOR2_X1 U3023 ( .A(n3025), .B(n3026), .Z(n2908) );
  XNOR2_X1 U3024 ( .A(n3027), .B(n3028), .ZN(n3025) );
  NAND2_X1 U3025 ( .A1(n2893), .A2(n2182), .ZN(n3027) );
  XNOR2_X1 U3026 ( .A(n3029), .B(n3030), .ZN(n2912) );
  XNOR2_X1 U3027 ( .A(n3031), .B(n3032), .ZN(n3030) );
  XOR2_X1 U3028 ( .A(n3033), .B(n3034), .Z(n2915) );
  XOR2_X1 U3029 ( .A(n3035), .B(n3036), .Z(n3033) );
  NOR2_X1 U3030 ( .A1(n2892), .A2(n2394), .ZN(n3036) );
  XNOR2_X1 U3031 ( .A(n3037), .B(n3038), .ZN(n2920) );
  XNOR2_X1 U3032 ( .A(n3039), .B(n3040), .ZN(n3038) );
  XOR2_X1 U3033 ( .A(n3041), .B(n3042), .Z(n2923) );
  XOR2_X1 U3034 ( .A(n3043), .B(n3044), .Z(n3041) );
  XOR2_X1 U3035 ( .A(n3045), .B(n3046), .Z(n2928) );
  XOR2_X1 U3036 ( .A(n3047), .B(n3048), .Z(n3045) );
  NOR2_X1 U3037 ( .A1(n2210), .A2(n2892), .ZN(n3048) );
  XOR2_X1 U3038 ( .A(n3049), .B(n3050), .Z(n2933) );
  XOR2_X1 U3039 ( .A(n3051), .B(n3052), .Z(n3050) );
  NAND2_X1 U3040 ( .A1(n2133), .A2(n2893), .ZN(n3052) );
  XOR2_X1 U3041 ( .A(n3053), .B(n3054), .Z(n2937) );
  XOR2_X1 U3042 ( .A(n3055), .B(n3056), .Z(n3054) );
  NAND2_X1 U3043 ( .A1(n2893), .A2(n2692), .ZN(n3056) );
  XNOR2_X1 U3044 ( .A(n3057), .B(n3058), .ZN(n2940) );
  XOR2_X1 U3045 ( .A(n3059), .B(n3060), .Z(n3058) );
  NAND2_X1 U3046 ( .A1(n2893), .A2(n2117), .ZN(n3060) );
  XNOR2_X1 U3047 ( .A(n3061), .B(n3062), .ZN(n2945) );
  XOR2_X1 U3048 ( .A(n3063), .B(n3064), .Z(n3062) );
  NAND2_X1 U3049 ( .A1(n2459), .A2(n2893), .ZN(n3064) );
  XNOR2_X1 U3050 ( .A(n3065), .B(n3066), .ZN(n2948) );
  XOR2_X1 U3051 ( .A(n3067), .B(n3068), .Z(n3066) );
  NAND2_X1 U3052 ( .A1(n1917), .A2(n2893), .ZN(n3068) );
  XNOR2_X1 U3053 ( .A(n3069), .B(n3070), .ZN(n2831) );
  XOR2_X1 U3054 ( .A(n3071), .B(n3072), .Z(n3070) );
  NAND2_X1 U3055 ( .A1(n2095), .A2(n2893), .ZN(n3072) );
  NAND2_X1 U3056 ( .A1(n3073), .A2(n3074), .ZN(n1933) );
  OR2_X1 U3057 ( .A1(n2961), .A2(n2960), .ZN(n3074) );
  XNOR2_X1 U3058 ( .A(n3075), .B(n3076), .ZN(n3073) );
  NAND2_X1 U3059 ( .A1(n3077), .A2(n3078), .ZN(n1934) );
  XOR2_X1 U3060 ( .A(n3075), .B(n3076), .Z(n3078) );
  NOR2_X1 U3061 ( .A1(n2960), .A2(n2961), .ZN(n3077) );
  XOR2_X1 U3062 ( .A(n3079), .B(n3080), .Z(n2961) );
  XOR2_X1 U3063 ( .A(n3081), .B(n3082), .Z(n3080) );
  NAND2_X1 U3064 ( .A1(n3015), .A2(n2053), .ZN(n3082) );
  AND2_X1 U3065 ( .A1(n3083), .A2(n3084), .ZN(n2960) );
  NAND2_X1 U3066 ( .A1(n3085), .A2(n2893), .ZN(n3084) );
  NOR2_X1 U3067 ( .A1(n3086), .A2(n2026), .ZN(n3085) );
  NOR2_X1 U3068 ( .A1(n2958), .A2(n2957), .ZN(n3086) );
  NAND2_X1 U3069 ( .A1(n2957), .A2(n2958), .ZN(n3083) );
  NAND2_X1 U3070 ( .A1(n3087), .A2(n3088), .ZN(n2958) );
  NAND2_X1 U3071 ( .A1(n3089), .A2(n2095), .ZN(n3088) );
  NOR2_X1 U3072 ( .A1(n3090), .A2(n2892), .ZN(n3089) );
  NOR2_X1 U3073 ( .A1(n3069), .A2(n3071), .ZN(n3090) );
  NAND2_X1 U3074 ( .A1(n3069), .A2(n3071), .ZN(n3087) );
  NAND2_X1 U3075 ( .A1(n3091), .A2(n3092), .ZN(n3071) );
  NAND2_X1 U3076 ( .A1(n3093), .A2(n2101), .ZN(n3092) );
  NOR2_X1 U3077 ( .A1(n3094), .A2(n2892), .ZN(n3093) );
  NOR2_X1 U3078 ( .A1(n3065), .A2(n3067), .ZN(n3094) );
  NAND2_X1 U3079 ( .A1(n3065), .A2(n3067), .ZN(n3091) );
  NAND2_X1 U3080 ( .A1(n3095), .A2(n3096), .ZN(n3067) );
  NAND2_X1 U3081 ( .A1(n3097), .A2(n2459), .ZN(n3096) );
  NOR2_X1 U3082 ( .A1(n3098), .A2(n2892), .ZN(n3097) );
  NOR2_X1 U3083 ( .A1(n3061), .A2(n3063), .ZN(n3098) );
  NAND2_X1 U3084 ( .A1(n3061), .A2(n3063), .ZN(n3095) );
  NAND2_X1 U3085 ( .A1(n3099), .A2(n3100), .ZN(n3063) );
  NAND2_X1 U3086 ( .A1(n3101), .A2(n2893), .ZN(n3100) );
  NOR2_X1 U3087 ( .A1(n3102), .A2(n2370), .ZN(n3101) );
  NOR2_X1 U3088 ( .A1(n3059), .A2(n3057), .ZN(n3102) );
  NAND2_X1 U3089 ( .A1(n3057), .A2(n3059), .ZN(n3099) );
  NAND2_X1 U3090 ( .A1(n3103), .A2(n3104), .ZN(n3059) );
  NAND2_X1 U3091 ( .A1(n3105), .A2(n2893), .ZN(n3104) );
  NOR2_X1 U3092 ( .A1(n3106), .A2(n2211), .ZN(n3105) );
  NOR2_X1 U3093 ( .A1(n3055), .A2(n3053), .ZN(n3106) );
  NAND2_X1 U3094 ( .A1(n3053), .A2(n3055), .ZN(n3103) );
  NAND2_X1 U3095 ( .A1(n3107), .A2(n3108), .ZN(n3055) );
  NAND2_X1 U3096 ( .A1(n3109), .A2(n2133), .ZN(n3108) );
  NOR2_X1 U3097 ( .A1(n3110), .A2(n2892), .ZN(n3109) );
  NOR2_X1 U3098 ( .A1(n3051), .A2(n3049), .ZN(n3110) );
  NAND2_X1 U3099 ( .A1(n3049), .A2(n3051), .ZN(n3107) );
  NAND2_X1 U3100 ( .A1(n3111), .A2(n3112), .ZN(n3051) );
  NAND2_X1 U3101 ( .A1(n3113), .A2(n2893), .ZN(n3112) );
  NOR2_X1 U3102 ( .A1(n3114), .A2(n2210), .ZN(n3113) );
  NOR2_X1 U3103 ( .A1(n3047), .A2(n3046), .ZN(n3114) );
  NAND2_X1 U3104 ( .A1(n3046), .A2(n3047), .ZN(n3111) );
  NAND2_X1 U3105 ( .A1(n3115), .A2(n3116), .ZN(n3047) );
  NAND2_X1 U3106 ( .A1(n3044), .A2(n3117), .ZN(n3116) );
  OR2_X1 U3107 ( .A1(n3042), .A2(n3043), .ZN(n3117) );
  NOR2_X1 U3108 ( .A1(n2386), .A2(n2892), .ZN(n3044) );
  NAND2_X1 U3109 ( .A1(n3042), .A2(n3043), .ZN(n3115) );
  NAND2_X1 U3110 ( .A1(n3118), .A2(n3119), .ZN(n3043) );
  NAND2_X1 U3111 ( .A1(n3040), .A2(n3120), .ZN(n3119) );
  OR2_X1 U3112 ( .A1(n3037), .A2(n3039), .ZN(n3120) );
  NOR2_X1 U3113 ( .A1(n2892), .A2(n2209), .ZN(n3040) );
  NAND2_X1 U3114 ( .A1(n3037), .A2(n3039), .ZN(n3118) );
  NAND2_X1 U3115 ( .A1(n3121), .A2(n3122), .ZN(n3039) );
  NAND2_X1 U3116 ( .A1(n3123), .A2(n2165), .ZN(n3122) );
  NOR2_X1 U3117 ( .A1(n3124), .A2(n2892), .ZN(n3123) );
  NOR2_X1 U3118 ( .A1(n3034), .A2(n3035), .ZN(n3124) );
  NAND2_X1 U3119 ( .A1(n3034), .A2(n3035), .ZN(n3121) );
  NAND2_X1 U3120 ( .A1(n3125), .A2(n3126), .ZN(n3035) );
  NAND2_X1 U3121 ( .A1(n3032), .A2(n3127), .ZN(n3126) );
  OR2_X1 U3122 ( .A1(n3029), .A2(n3031), .ZN(n3127) );
  NOR2_X1 U3123 ( .A1(n2892), .A2(n2291), .ZN(n3032) );
  NAND2_X1 U3124 ( .A1(n3029), .A2(n3031), .ZN(n3125) );
  NAND2_X1 U3125 ( .A1(n3128), .A2(n3129), .ZN(n3031) );
  NAND2_X1 U3126 ( .A1(n3130), .A2(n2893), .ZN(n3129) );
  NOR2_X1 U3127 ( .A1(n3131), .A2(n2187), .ZN(n3130) );
  NOR2_X1 U3128 ( .A1(n3026), .A2(n3028), .ZN(n3131) );
  NAND2_X1 U3129 ( .A1(n3026), .A2(n3028), .ZN(n3128) );
  NAND2_X1 U3130 ( .A1(n3132), .A2(n3133), .ZN(n3028) );
  NAND2_X1 U3131 ( .A1(n3021), .A2(n3134), .ZN(n3133) );
  NAND2_X1 U3132 ( .A1(n3024), .A2(n3023), .ZN(n3134) );
  NOR2_X1 U3133 ( .A1(n2892), .A2(n2203), .ZN(n3021) );
  OR2_X1 U3134 ( .A1(n3023), .A2(n3024), .ZN(n3132) );
  AND2_X1 U3135 ( .A1(n3135), .A2(n3136), .ZN(n3024) );
  NAND2_X1 U3136 ( .A1(n3015), .A2(n3137), .ZN(n3136) );
  NAND2_X1 U3137 ( .A1(n1953), .A2(n3138), .ZN(n3137) );
  NAND2_X1 U3138 ( .A1(n3139), .A2(n1956), .ZN(n3138) );
  NAND2_X1 U3139 ( .A1(n3140), .A2(n3141), .ZN(n3135) );
  NAND2_X1 U3140 ( .A1(n1959), .A2(n3142), .ZN(n3141) );
  NAND2_X1 U3141 ( .A1(n1961), .A2(n3014), .ZN(n3142) );
  NAND2_X1 U3142 ( .A1(n3143), .A2(n3015), .ZN(n3023) );
  NOR2_X1 U3143 ( .A1(n2306), .A2(n2892), .ZN(n3143) );
  INV_X1 U3144 ( .A(n2893), .ZN(n2892) );
  XOR2_X1 U3145 ( .A(d_7_), .B(c_7_), .Z(n3145) );
  XNOR2_X1 U3146 ( .A(n3146), .B(n3147), .ZN(n3026) );
  XNOR2_X1 U3147 ( .A(n3148), .B(n3149), .ZN(n3147) );
  XOR2_X1 U3148 ( .A(n3150), .B(n3151), .Z(n3029) );
  XNOR2_X1 U3149 ( .A(n3152), .B(n3153), .ZN(n3150) );
  NAND2_X1 U3150 ( .A1(n3015), .A2(n2182), .ZN(n3152) );
  XNOR2_X1 U3151 ( .A(n3154), .B(n3155), .ZN(n3034) );
  XNOR2_X1 U3152 ( .A(n3156), .B(n3157), .ZN(n3155) );
  XOR2_X1 U3153 ( .A(n3158), .B(n3159), .Z(n3037) );
  XOR2_X1 U3154 ( .A(n3160), .B(n3161), .Z(n3158) );
  NOR2_X1 U3155 ( .A1(n3014), .A2(n2394), .ZN(n3161) );
  XNOR2_X1 U3156 ( .A(n3162), .B(n3163), .ZN(n3042) );
  XOR2_X1 U3157 ( .A(n3164), .B(n3165), .Z(n3163) );
  NAND2_X1 U3158 ( .A1(n3015), .A2(n3166), .ZN(n3165) );
  XNOR2_X1 U3159 ( .A(n3167), .B(n3168), .ZN(n3046) );
  XNOR2_X1 U3160 ( .A(n3169), .B(n3170), .ZN(n3168) );
  XNOR2_X1 U3161 ( .A(n3171), .B(n3172), .ZN(n3049) );
  XNOR2_X1 U3162 ( .A(n3173), .B(n3174), .ZN(n3171) );
  XOR2_X1 U3163 ( .A(n3175), .B(n3176), .Z(n3053) );
  XNOR2_X1 U3164 ( .A(n3177), .B(n3178), .ZN(n3175) );
  NAND2_X1 U3165 ( .A1(n2133), .A2(n3015), .ZN(n3177) );
  XOR2_X1 U3166 ( .A(n3179), .B(n3180), .Z(n3057) );
  XOR2_X1 U3167 ( .A(n3181), .B(n3182), .Z(n3180) );
  XNOR2_X1 U3168 ( .A(n3183), .B(n3184), .ZN(n3061) );
  XNOR2_X1 U3169 ( .A(n3185), .B(n3186), .ZN(n3184) );
  XNOR2_X1 U3170 ( .A(n3187), .B(n3188), .ZN(n3065) );
  NAND2_X1 U3171 ( .A1(n3189), .A2(n3190), .ZN(n3187) );
  XNOR2_X1 U3172 ( .A(n3191), .B(n3192), .ZN(n3069) );
  XOR2_X1 U3173 ( .A(n3193), .B(n3194), .Z(n3192) );
  NAND2_X1 U3174 ( .A1(n1917), .A2(n3015), .ZN(n3194) );
  XNOR2_X1 U3175 ( .A(n3195), .B(n3196), .ZN(n2957) );
  XOR2_X1 U3176 ( .A(n3197), .B(n3198), .Z(n3196) );
  NAND2_X1 U3177 ( .A1(n2095), .A2(n3015), .ZN(n3198) );
  NAND2_X1 U3178 ( .A1(n3199), .A2(n3200), .ZN(n1937) );
  NAND2_X1 U3179 ( .A1(n3076), .A2(n3075), .ZN(n3200) );
  XOR2_X1 U3180 ( .A(n3201), .B(n3202), .Z(n3199) );
  NAND2_X1 U3181 ( .A1(n3203), .A2(n3204), .ZN(n1938) );
  XOR2_X1 U3182 ( .A(n3205), .B(n3202), .Z(n3204) );
  INV_X1 U3183 ( .A(n3206), .ZN(n3202) );
  AND2_X1 U3184 ( .A1(n3075), .A2(n3076), .ZN(n3203) );
  XNOR2_X1 U3185 ( .A(n3207), .B(n3208), .ZN(n3076) );
  XOR2_X1 U3186 ( .A(n3209), .B(n3210), .Z(n3208) );
  NAND2_X1 U3187 ( .A1(n3140), .A2(n2053), .ZN(n3210) );
  NAND2_X1 U3188 ( .A1(n3211), .A2(n3212), .ZN(n3075) );
  NAND2_X1 U3189 ( .A1(n3213), .A2(n3015), .ZN(n3212) );
  NOR2_X1 U3190 ( .A1(n3214), .A2(n2026), .ZN(n3213) );
  NOR2_X1 U3191 ( .A1(n3081), .A2(n3079), .ZN(n3214) );
  NAND2_X1 U3192 ( .A1(n3079), .A2(n3081), .ZN(n3211) );
  NAND2_X1 U3193 ( .A1(n3215), .A2(n3216), .ZN(n3081) );
  NAND2_X1 U3194 ( .A1(n3217), .A2(n2095), .ZN(n3216) );
  NOR2_X1 U3195 ( .A1(n3218), .A2(n3014), .ZN(n3217) );
  NOR2_X1 U3196 ( .A1(n3195), .A2(n3197), .ZN(n3218) );
  NAND2_X1 U3197 ( .A1(n3195), .A2(n3197), .ZN(n3215) );
  NAND2_X1 U3198 ( .A1(n3219), .A2(n3220), .ZN(n3197) );
  NAND2_X1 U3199 ( .A1(n3221), .A2(n2101), .ZN(n3220) );
  NOR2_X1 U3200 ( .A1(n3222), .A2(n3014), .ZN(n3221) );
  NOR2_X1 U3201 ( .A1(n3193), .A2(n3191), .ZN(n3222) );
  NAND2_X1 U3202 ( .A1(n3191), .A2(n3193), .ZN(n3219) );
  NAND2_X1 U3203 ( .A1(n3189), .A2(n3223), .ZN(n3193) );
  NAND2_X1 U3204 ( .A1(n3188), .A2(n3190), .ZN(n3223) );
  NAND2_X1 U3205 ( .A1(n3224), .A2(n3225), .ZN(n3190) );
  NAND2_X1 U3206 ( .A1(n2459), .A2(n3015), .ZN(n3225) );
  INV_X1 U3207 ( .A(n3226), .ZN(n3224) );
  XNOR2_X1 U3208 ( .A(n3227), .B(n3228), .ZN(n3188) );
  XOR2_X1 U3209 ( .A(n3229), .B(n3230), .Z(n3228) );
  NAND2_X1 U3210 ( .A1(n3140), .A2(n2117), .ZN(n3230) );
  NAND2_X1 U3211 ( .A1(n2459), .A2(n3226), .ZN(n3189) );
  NAND2_X1 U3212 ( .A1(n3231), .A2(n3232), .ZN(n3226) );
  NAND2_X1 U3213 ( .A1(n3186), .A2(n3233), .ZN(n3232) );
  OR2_X1 U3214 ( .A1(n3183), .A2(n3185), .ZN(n3233) );
  NOR2_X1 U3215 ( .A1(n3014), .A2(n2370), .ZN(n3186) );
  NAND2_X1 U3216 ( .A1(n3183), .A2(n3185), .ZN(n3231) );
  NAND2_X1 U3217 ( .A1(n3234), .A2(n3235), .ZN(n3185) );
  NAND2_X1 U3218 ( .A1(n3182), .A2(n3236), .ZN(n3235) );
  NAND2_X1 U3219 ( .A1(n3181), .A2(n3179), .ZN(n3236) );
  NOR2_X1 U3220 ( .A1(n3014), .A2(n2211), .ZN(n3182) );
  OR2_X1 U3221 ( .A1(n3179), .A2(n3181), .ZN(n3234) );
  AND2_X1 U3222 ( .A1(n3237), .A2(n3238), .ZN(n3181) );
  NAND2_X1 U3223 ( .A1(n3239), .A2(n2133), .ZN(n3238) );
  NOR2_X1 U3224 ( .A1(n3240), .A2(n3014), .ZN(n3239) );
  NOR2_X1 U3225 ( .A1(n3176), .A2(n3178), .ZN(n3240) );
  NAND2_X1 U3226 ( .A1(n3176), .A2(n3178), .ZN(n3237) );
  NAND2_X1 U3227 ( .A1(n3241), .A2(n3242), .ZN(n3178) );
  NAND2_X1 U3228 ( .A1(n3174), .A2(n3243), .ZN(n3242) );
  NAND2_X1 U3229 ( .A1(n3173), .A2(n3172), .ZN(n3243) );
  NOR2_X1 U3230 ( .A1(n3014), .A2(n2210), .ZN(n3174) );
  OR2_X1 U3231 ( .A1(n3172), .A2(n3173), .ZN(n3241) );
  AND2_X1 U3232 ( .A1(n3244), .A2(n3245), .ZN(n3173) );
  NAND2_X1 U3233 ( .A1(n3170), .A2(n3246), .ZN(n3245) );
  OR2_X1 U3234 ( .A1(n3169), .A2(n3167), .ZN(n3246) );
  NOR2_X1 U3235 ( .A1(n2386), .A2(n3014), .ZN(n3170) );
  NAND2_X1 U3236 ( .A1(n3167), .A2(n3169), .ZN(n3244) );
  NAND2_X1 U3237 ( .A1(n3247), .A2(n3248), .ZN(n3169) );
  NAND2_X1 U3238 ( .A1(n3249), .A2(n3015), .ZN(n3248) );
  NOR2_X1 U3239 ( .A1(n3250), .A2(n2209), .ZN(n3249) );
  NOR2_X1 U3240 ( .A1(n3162), .A2(n3164), .ZN(n3250) );
  NAND2_X1 U3241 ( .A1(n3162), .A2(n3164), .ZN(n3247) );
  NAND2_X1 U3242 ( .A1(n3251), .A2(n3252), .ZN(n3164) );
  NAND2_X1 U3243 ( .A1(n3253), .A2(n2165), .ZN(n3252) );
  NOR2_X1 U3244 ( .A1(n3254), .A2(n3014), .ZN(n3253) );
  NOR2_X1 U3245 ( .A1(n3159), .A2(n3160), .ZN(n3254) );
  NAND2_X1 U3246 ( .A1(n3159), .A2(n3160), .ZN(n3251) );
  NAND2_X1 U3247 ( .A1(n3255), .A2(n3256), .ZN(n3160) );
  NAND2_X1 U3248 ( .A1(n3157), .A2(n3257), .ZN(n3256) );
  OR2_X1 U3249 ( .A1(n3154), .A2(n3156), .ZN(n3257) );
  NOR2_X1 U3250 ( .A1(n3014), .A2(n2291), .ZN(n3157) );
  NAND2_X1 U3251 ( .A1(n3154), .A2(n3156), .ZN(n3255) );
  NAND2_X1 U3252 ( .A1(n3258), .A2(n3259), .ZN(n3156) );
  NAND2_X1 U3253 ( .A1(n3260), .A2(n3015), .ZN(n3259) );
  NOR2_X1 U3254 ( .A1(n3261), .A2(n2187), .ZN(n3260) );
  NOR2_X1 U3255 ( .A1(n3151), .A2(n3153), .ZN(n3261) );
  NAND2_X1 U3256 ( .A1(n3151), .A2(n3153), .ZN(n3258) );
  NAND2_X1 U3257 ( .A1(n3262), .A2(n3263), .ZN(n3153) );
  NAND2_X1 U3258 ( .A1(n3146), .A2(n3264), .ZN(n3263) );
  NAND2_X1 U3259 ( .A1(n3149), .A2(n3148), .ZN(n3264) );
  NOR2_X1 U3260 ( .A1(n3014), .A2(n2203), .ZN(n3146) );
  OR2_X1 U3261 ( .A1(n3148), .A2(n3149), .ZN(n3262) );
  AND2_X1 U3262 ( .A1(n3265), .A2(n3266), .ZN(n3149) );
  NAND2_X1 U3263 ( .A1(n3140), .A2(n3267), .ZN(n3266) );
  NAND2_X1 U3264 ( .A1(n1953), .A2(n3268), .ZN(n3267) );
  NAND2_X1 U3265 ( .A1(n3269), .A2(n1956), .ZN(n3268) );
  NAND2_X1 U3266 ( .A1(n1916), .A2(n3271), .ZN(n3265) );
  NAND2_X1 U3267 ( .A1(n1959), .A2(n3272), .ZN(n3271) );
  NAND2_X1 U3268 ( .A1(n1961), .A2(n3139), .ZN(n3272) );
  NAND2_X1 U3269 ( .A1(n3273), .A2(n3140), .ZN(n3148) );
  NOR2_X1 U3270 ( .A1(n2306), .A2(n3014), .ZN(n3273) );
  INV_X1 U3271 ( .A(n3015), .ZN(n3014) );
  XOR2_X1 U3272 ( .A(d_6_), .B(c_6_), .Z(n3275) );
  XNOR2_X1 U3273 ( .A(n3276), .B(n3277), .ZN(n3151) );
  XNOR2_X1 U3274 ( .A(n3278), .B(n3279), .ZN(n3277) );
  XOR2_X1 U3275 ( .A(n3280), .B(n3281), .Z(n3154) );
  XNOR2_X1 U3276 ( .A(n3282), .B(n3283), .ZN(n3280) );
  NAND2_X1 U3277 ( .A1(n3140), .A2(n2182), .ZN(n3282) );
  XNOR2_X1 U3278 ( .A(n3284), .B(n3285), .ZN(n3159) );
  XNOR2_X1 U3279 ( .A(n3286), .B(n3287), .ZN(n3285) );
  XOR2_X1 U3280 ( .A(n3288), .B(n3289), .Z(n3162) );
  XOR2_X1 U3281 ( .A(n3290), .B(n3291), .Z(n3288) );
  XOR2_X1 U3282 ( .A(n3292), .B(n3293), .Z(n3167) );
  XOR2_X1 U3283 ( .A(n3294), .B(n3295), .Z(n3292) );
  NOR2_X1 U3284 ( .A1(n2209), .A2(n3139), .ZN(n3295) );
  XOR2_X1 U3285 ( .A(n3296), .B(n3297), .Z(n3172) );
  XOR2_X1 U3286 ( .A(n3298), .B(n3299), .Z(n3297) );
  NAND2_X1 U3287 ( .A1(n2149), .A2(n3140), .ZN(n3299) );
  XNOR2_X1 U3288 ( .A(n3300), .B(n3301), .ZN(n3176) );
  XOR2_X1 U3289 ( .A(n3302), .B(n3303), .Z(n3301) );
  NAND2_X1 U3290 ( .A1(n3140), .A2(n2927), .ZN(n3303) );
  XNOR2_X1 U3291 ( .A(n3304), .B(n3305), .ZN(n3179) );
  XOR2_X1 U3292 ( .A(n3306), .B(n3307), .Z(n3304) );
  NOR2_X1 U3293 ( .A1(n3139), .A2(n2378), .ZN(n3307) );
  XOR2_X1 U3294 ( .A(n3308), .B(n3309), .Z(n3183) );
  XOR2_X1 U3295 ( .A(n3310), .B(n3311), .Z(n3308) );
  NOR2_X1 U3296 ( .A1(n2211), .A2(n3139), .ZN(n3311) );
  XNOR2_X1 U3297 ( .A(n3312), .B(n3313), .ZN(n3191) );
  XOR2_X1 U3298 ( .A(n3314), .B(n3315), .Z(n3313) );
  NAND2_X1 U3299 ( .A1(n2459), .A2(n3140), .ZN(n3315) );
  XNOR2_X1 U3300 ( .A(n3316), .B(n3317), .ZN(n3195) );
  XOR2_X1 U3301 ( .A(n3318), .B(n3319), .Z(n3317) );
  NAND2_X1 U3302 ( .A1(n1917), .A2(n3140), .ZN(n3319) );
  XNOR2_X1 U3303 ( .A(n3320), .B(n3321), .ZN(n3079) );
  XOR2_X1 U3304 ( .A(n3322), .B(n3323), .Z(n3321) );
  NAND2_X1 U3305 ( .A1(n2095), .A2(n3140), .ZN(n3323) );
  NAND2_X1 U3306 ( .A1(n3324), .A2(n3325), .ZN(n1941) );
  NAND2_X1 U3307 ( .A1(n3206), .A2(n3201), .ZN(n3325) );
  NAND2_X1 U3308 ( .A1(n3326), .A2(n3206), .ZN(n1942) );
  XNOR2_X1 U3309 ( .A(n3327), .B(n3328), .ZN(n3206) );
  XOR2_X1 U3310 ( .A(n3329), .B(n3330), .Z(n3328) );
  NAND2_X1 U3311 ( .A1(n1916), .A2(n2053), .ZN(n3330) );
  NOR2_X1 U3312 ( .A1(n3205), .A2(n3324), .ZN(n3326) );
  XOR2_X1 U3313 ( .A(n3331), .B(n3332), .Z(n3324) );
  INV_X1 U3314 ( .A(n3333), .ZN(n3332) );
  INV_X1 U3315 ( .A(n3201), .ZN(n3205) );
  NAND2_X1 U3316 ( .A1(n3334), .A2(n3335), .ZN(n3201) );
  NAND2_X1 U3317 ( .A1(n3336), .A2(n3140), .ZN(n3335) );
  NOR2_X1 U3318 ( .A1(n3337), .A2(n2026), .ZN(n3336) );
  NOR2_X1 U3319 ( .A1(n3207), .A2(n3209), .ZN(n3337) );
  NAND2_X1 U3320 ( .A1(n3207), .A2(n3209), .ZN(n3334) );
  NAND2_X1 U3321 ( .A1(n3338), .A2(n3339), .ZN(n3209) );
  NAND2_X1 U3322 ( .A1(n3340), .A2(n2095), .ZN(n3339) );
  NOR2_X1 U3323 ( .A1(n3341), .A2(n3139), .ZN(n3340) );
  NOR2_X1 U3324 ( .A1(n3320), .A2(n3322), .ZN(n3341) );
  NAND2_X1 U3325 ( .A1(n3320), .A2(n3322), .ZN(n3338) );
  NAND2_X1 U3326 ( .A1(n3342), .A2(n3343), .ZN(n3322) );
  NAND2_X1 U3327 ( .A1(n3344), .A2(n2101), .ZN(n3343) );
  NOR2_X1 U3328 ( .A1(n3345), .A2(n3139), .ZN(n3344) );
  NOR2_X1 U3329 ( .A1(n3318), .A2(n3316), .ZN(n3345) );
  NAND2_X1 U3330 ( .A1(n3316), .A2(n3318), .ZN(n3342) );
  NAND2_X1 U3331 ( .A1(n3346), .A2(n3347), .ZN(n3318) );
  NAND2_X1 U3332 ( .A1(n3348), .A2(n2459), .ZN(n3347) );
  NOR2_X1 U3333 ( .A1(n3349), .A2(n3139), .ZN(n3348) );
  NOR2_X1 U3334 ( .A1(n3312), .A2(n3314), .ZN(n3349) );
  NAND2_X1 U3335 ( .A1(n3312), .A2(n3314), .ZN(n3346) );
  NAND2_X1 U3336 ( .A1(n3350), .A2(n3351), .ZN(n3314) );
  NAND2_X1 U3337 ( .A1(n3352), .A2(n3140), .ZN(n3351) );
  NOR2_X1 U3338 ( .A1(n3353), .A2(n2370), .ZN(n3352) );
  NOR2_X1 U3339 ( .A1(n3229), .A2(n3227), .ZN(n3353) );
  NAND2_X1 U3340 ( .A1(n3227), .A2(n3229), .ZN(n3350) );
  NAND2_X1 U3341 ( .A1(n3354), .A2(n3355), .ZN(n3229) );
  NAND2_X1 U3342 ( .A1(n3356), .A2(n3140), .ZN(n3355) );
  NOR2_X1 U3343 ( .A1(n3357), .A2(n2211), .ZN(n3356) );
  NOR2_X1 U3344 ( .A1(n3309), .A2(n3310), .ZN(n3357) );
  NAND2_X1 U3345 ( .A1(n3309), .A2(n3310), .ZN(n3354) );
  NAND2_X1 U3346 ( .A1(n3358), .A2(n3359), .ZN(n3310) );
  NAND2_X1 U3347 ( .A1(n3360), .A2(n2133), .ZN(n3359) );
  NOR2_X1 U3348 ( .A1(n3361), .A2(n3139), .ZN(n3360) );
  NOR2_X1 U3349 ( .A1(n3306), .A2(n3305), .ZN(n3361) );
  NAND2_X1 U3350 ( .A1(n3305), .A2(n3306), .ZN(n3358) );
  NAND2_X1 U3351 ( .A1(n3362), .A2(n3363), .ZN(n3306) );
  NAND2_X1 U3352 ( .A1(n3364), .A2(n3140), .ZN(n3363) );
  NOR2_X1 U3353 ( .A1(n3365), .A2(n2210), .ZN(n3364) );
  NOR2_X1 U3354 ( .A1(n3302), .A2(n3300), .ZN(n3365) );
  NAND2_X1 U3355 ( .A1(n3300), .A2(n3302), .ZN(n3362) );
  NAND2_X1 U3356 ( .A1(n3366), .A2(n3367), .ZN(n3302) );
  NAND2_X1 U3357 ( .A1(n3368), .A2(n2149), .ZN(n3367) );
  NOR2_X1 U3358 ( .A1(n3369), .A2(n3139), .ZN(n3368) );
  NOR2_X1 U3359 ( .A1(n3298), .A2(n3296), .ZN(n3369) );
  NAND2_X1 U3360 ( .A1(n3296), .A2(n3298), .ZN(n3366) );
  NAND2_X1 U3361 ( .A1(n3370), .A2(n3371), .ZN(n3298) );
  NAND2_X1 U3362 ( .A1(n3372), .A2(n3140), .ZN(n3371) );
  NOR2_X1 U3363 ( .A1(n3373), .A2(n2209), .ZN(n3372) );
  NOR2_X1 U3364 ( .A1(n3294), .A2(n3293), .ZN(n3373) );
  NAND2_X1 U3365 ( .A1(n3293), .A2(n3294), .ZN(n3370) );
  NAND2_X1 U3366 ( .A1(n3374), .A2(n3375), .ZN(n3294) );
  NAND2_X1 U3367 ( .A1(n3290), .A2(n3376), .ZN(n3375) );
  OR2_X1 U3368 ( .A1(n3289), .A2(n3291), .ZN(n3376) );
  NOR2_X1 U3369 ( .A1(n3139), .A2(n2394), .ZN(n3290) );
  NAND2_X1 U3370 ( .A1(n3289), .A2(n3291), .ZN(n3374) );
  NAND2_X1 U3371 ( .A1(n3377), .A2(n3378), .ZN(n3291) );
  NAND2_X1 U3372 ( .A1(n3287), .A2(n3379), .ZN(n3378) );
  OR2_X1 U3373 ( .A1(n3284), .A2(n3286), .ZN(n3379) );
  NOR2_X1 U3374 ( .A1(n3139), .A2(n2291), .ZN(n3287) );
  NAND2_X1 U3375 ( .A1(n3284), .A2(n3286), .ZN(n3377) );
  NAND2_X1 U3376 ( .A1(n3380), .A2(n3381), .ZN(n3286) );
  NAND2_X1 U3377 ( .A1(n3382), .A2(n3140), .ZN(n3381) );
  NOR2_X1 U3378 ( .A1(n3383), .A2(n2187), .ZN(n3382) );
  NOR2_X1 U3379 ( .A1(n3281), .A2(n3283), .ZN(n3383) );
  NAND2_X1 U3380 ( .A1(n3281), .A2(n3283), .ZN(n3380) );
  NAND2_X1 U3381 ( .A1(n3384), .A2(n3385), .ZN(n3283) );
  NAND2_X1 U3382 ( .A1(n3276), .A2(n3386), .ZN(n3385) );
  NAND2_X1 U3383 ( .A1(n3279), .A2(n3278), .ZN(n3386) );
  NOR2_X1 U3384 ( .A1(n3139), .A2(n2203), .ZN(n3276) );
  OR2_X1 U3385 ( .A1(n3278), .A2(n3279), .ZN(n3384) );
  AND2_X1 U3386 ( .A1(n3387), .A2(n3388), .ZN(n3279) );
  NAND2_X1 U3387 ( .A1(n1916), .A2(n3389), .ZN(n3388) );
  NAND2_X1 U3388 ( .A1(n1953), .A2(n3390), .ZN(n3389) );
  NAND2_X1 U3389 ( .A1(n3391), .A2(n1956), .ZN(n3390) );
  NAND2_X1 U3390 ( .A1(n1918), .A2(n3393), .ZN(n3387) );
  NAND2_X1 U3391 ( .A1(n1959), .A2(n3394), .ZN(n3393) );
  NAND2_X1 U3392 ( .A1(n1961), .A2(n3269), .ZN(n3394) );
  NAND2_X1 U3393 ( .A1(n3395), .A2(n1916), .ZN(n3278) );
  NOR2_X1 U3394 ( .A1(n2306), .A2(n3139), .ZN(n3395) );
  INV_X1 U3395 ( .A(n3140), .ZN(n3139) );
  XOR2_X1 U3396 ( .A(d_5_), .B(c_5_), .Z(n3397) );
  XNOR2_X1 U3397 ( .A(n3398), .B(n3399), .ZN(n3281) );
  XNOR2_X1 U3398 ( .A(n3400), .B(n3401), .ZN(n3399) );
  XOR2_X1 U3399 ( .A(n3402), .B(n3403), .Z(n3284) );
  XNOR2_X1 U3400 ( .A(n3404), .B(n3405), .ZN(n3402) );
  NAND2_X1 U3401 ( .A1(n1916), .A2(n2182), .ZN(n3404) );
  XNOR2_X1 U3402 ( .A(n3406), .B(n3407), .ZN(n3289) );
  XOR2_X1 U3403 ( .A(n3408), .B(n3409), .Z(n3407) );
  NAND2_X1 U3404 ( .A1(n1916), .A2(n2208), .ZN(n3409) );
  XNOR2_X1 U3405 ( .A(n3410), .B(n3411), .ZN(n3293) );
  XOR2_X1 U3406 ( .A(n3412), .B(n3413), .Z(n3411) );
  NAND2_X1 U3407 ( .A1(n1916), .A2(n2165), .ZN(n3413) );
  XNOR2_X1 U3408 ( .A(n3414), .B(n3415), .ZN(n3296) );
  XNOR2_X1 U3409 ( .A(n3416), .B(n3417), .ZN(n3414) );
  XNOR2_X1 U3410 ( .A(n3418), .B(n3419), .ZN(n3300) );
  NAND2_X1 U3411 ( .A1(n3420), .A2(n3421), .ZN(n3418) );
  XNOR2_X1 U3412 ( .A(n3422), .B(n3423), .ZN(n3305) );
  XOR2_X1 U3413 ( .A(n3424), .B(n3425), .Z(n3423) );
  NAND2_X1 U3414 ( .A1(n1916), .A2(n2927), .ZN(n3425) );
  XNOR2_X1 U3415 ( .A(n3426), .B(n3427), .ZN(n3309) );
  XOR2_X1 U3416 ( .A(n3428), .B(n3429), .Z(n3427) );
  NAND2_X1 U3417 ( .A1(n2133), .A2(n1916), .ZN(n3429) );
  XNOR2_X1 U3418 ( .A(n3430), .B(n3431), .ZN(n3227) );
  XOR2_X1 U3419 ( .A(n3432), .B(n3433), .Z(n3431) );
  NAND2_X1 U3420 ( .A1(n1916), .A2(n2692), .ZN(n3433) );
  XNOR2_X1 U3421 ( .A(n3434), .B(n3435), .ZN(n3312) );
  XOR2_X1 U3422 ( .A(n3436), .B(n3437), .Z(n3435) );
  NAND2_X1 U3423 ( .A1(n1916), .A2(n2117), .ZN(n3437) );
  XNOR2_X1 U3424 ( .A(n3438), .B(n3439), .ZN(n3316) );
  XOR2_X1 U3425 ( .A(n3440), .B(n3441), .Z(n3439) );
  NAND2_X1 U3426 ( .A1(n2459), .A2(n3270), .ZN(n3441) );
  XNOR2_X1 U3427 ( .A(n3442), .B(n3443), .ZN(n3320) );
  XOR2_X1 U3428 ( .A(n3444), .B(n3445), .Z(n3443) );
  NAND2_X1 U3429 ( .A1(n1917), .A2(n3270), .ZN(n3445) );
  XOR2_X1 U3430 ( .A(n3446), .B(n3447), .Z(n3207) );
  XOR2_X1 U3431 ( .A(n3448), .B(n3449), .Z(n3446) );
  NOR2_X1 U3432 ( .A1(n3269), .A2(n2241), .ZN(n3449) );
  NAND2_X1 U3433 ( .A1(n3450), .A2(n3451), .ZN(n1945) );
  NAND2_X1 U3434 ( .A1(n3333), .A2(n3331), .ZN(n3451) );
  NAND2_X1 U3435 ( .A1(n3452), .A2(n3333), .ZN(n1946) );
  XOR2_X1 U3436 ( .A(n3453), .B(n3454), .Z(n3333) );
  XOR2_X1 U3437 ( .A(n3455), .B(n3456), .Z(n3453) );
  NOR2_X1 U3438 ( .A1(n2026), .A2(n3391), .ZN(n3456) );
  NOR2_X1 U3439 ( .A1(n3457), .A2(n3450), .ZN(n3452) );
  XOR2_X1 U3440 ( .A(n3458), .B(n3459), .Z(n3450) );
  INV_X1 U3441 ( .A(n3331), .ZN(n3457) );
  NAND2_X1 U3442 ( .A1(n3460), .A2(n3461), .ZN(n3331) );
  NAND2_X1 U3443 ( .A1(n3462), .A2(n3270), .ZN(n3461) );
  NOR2_X1 U3444 ( .A1(n3463), .A2(n2026), .ZN(n3462) );
  NOR2_X1 U3445 ( .A1(n3329), .A2(n3327), .ZN(n3463) );
  NAND2_X1 U3446 ( .A1(n3327), .A2(n3329), .ZN(n3460) );
  NAND2_X1 U3447 ( .A1(n3464), .A2(n3465), .ZN(n3329) );
  NAND2_X1 U3448 ( .A1(n3466), .A2(n2095), .ZN(n3465) );
  NOR2_X1 U3449 ( .A1(n3467), .A2(n3269), .ZN(n3466) );
  NOR2_X1 U3450 ( .A1(n3448), .A2(n3447), .ZN(n3467) );
  NAND2_X1 U3451 ( .A1(n3447), .A2(n3448), .ZN(n3464) );
  NAND2_X1 U3452 ( .A1(n3468), .A2(n3469), .ZN(n3448) );
  NAND2_X1 U3453 ( .A1(n3470), .A2(n2101), .ZN(n3469) );
  NOR2_X1 U3454 ( .A1(n3471), .A2(n3269), .ZN(n3470) );
  NOR2_X1 U3455 ( .A1(n3444), .A2(n3442), .ZN(n3471) );
  NAND2_X1 U3456 ( .A1(n3442), .A2(n3444), .ZN(n3468) );
  NAND2_X1 U3457 ( .A1(n3472), .A2(n3473), .ZN(n3444) );
  NAND2_X1 U3458 ( .A1(n3474), .A2(n2459), .ZN(n3473) );
  NOR2_X1 U3459 ( .A1(n3475), .A2(n3269), .ZN(n3474) );
  NOR2_X1 U3460 ( .A1(n3438), .A2(n3440), .ZN(n3475) );
  NAND2_X1 U3461 ( .A1(n3438), .A2(n3440), .ZN(n3472) );
  NAND2_X1 U3462 ( .A1(n3476), .A2(n3477), .ZN(n3440) );
  NAND2_X1 U3463 ( .A1(n3478), .A2(n3270), .ZN(n3477) );
  NOR2_X1 U3464 ( .A1(n3479), .A2(n2370), .ZN(n3478) );
  NOR2_X1 U3465 ( .A1(n3436), .A2(n3434), .ZN(n3479) );
  NAND2_X1 U3466 ( .A1(n3434), .A2(n3436), .ZN(n3476) );
  NAND2_X1 U3467 ( .A1(n3480), .A2(n3481), .ZN(n3436) );
  NAND2_X1 U3468 ( .A1(n3482), .A2(n3270), .ZN(n3481) );
  NOR2_X1 U3469 ( .A1(n3483), .A2(n2211), .ZN(n3482) );
  NOR2_X1 U3470 ( .A1(n3430), .A2(n3432), .ZN(n3483) );
  NAND2_X1 U3471 ( .A1(n3430), .A2(n3432), .ZN(n3480) );
  NAND2_X1 U3472 ( .A1(n3484), .A2(n3485), .ZN(n3432) );
  NAND2_X1 U3473 ( .A1(n3486), .A2(n2133), .ZN(n3485) );
  NOR2_X1 U3474 ( .A1(n3487), .A2(n3269), .ZN(n3486) );
  NOR2_X1 U3475 ( .A1(n3428), .A2(n3426), .ZN(n3487) );
  NAND2_X1 U3476 ( .A1(n3426), .A2(n3428), .ZN(n3484) );
  NAND2_X1 U3477 ( .A1(n3488), .A2(n3489), .ZN(n3428) );
  NAND2_X1 U3478 ( .A1(n3490), .A2(n3270), .ZN(n3489) );
  NOR2_X1 U3479 ( .A1(n3491), .A2(n2210), .ZN(n3490) );
  NOR2_X1 U3480 ( .A1(n3422), .A2(n3424), .ZN(n3491) );
  NAND2_X1 U3481 ( .A1(n3422), .A2(n3424), .ZN(n3488) );
  NAND2_X1 U3482 ( .A1(n3420), .A2(n3492), .ZN(n3424) );
  NAND2_X1 U3483 ( .A1(n3419), .A2(n3421), .ZN(n3492) );
  NAND2_X1 U3484 ( .A1(n3493), .A2(n3494), .ZN(n3421) );
  NAND2_X1 U3485 ( .A1(n2149), .A2(n3270), .ZN(n3494) );
  INV_X1 U3486 ( .A(n3495), .ZN(n3493) );
  XNOR2_X1 U3487 ( .A(n3496), .B(n3497), .ZN(n3419) );
  XOR2_X1 U3488 ( .A(n3498), .B(n3499), .Z(n3497) );
  NAND2_X1 U3489 ( .A1(n1918), .A2(n3166), .ZN(n3499) );
  NAND2_X1 U3490 ( .A1(n2149), .A2(n3495), .ZN(n3420) );
  NAND2_X1 U3491 ( .A1(n3500), .A2(n3501), .ZN(n3495) );
  NAND2_X1 U3492 ( .A1(n3417), .A2(n3502), .ZN(n3501) );
  NAND2_X1 U3493 ( .A1(n3416), .A2(n3415), .ZN(n3502) );
  NOR2_X1 U3494 ( .A1(n3269), .A2(n2209), .ZN(n3417) );
  OR2_X1 U3495 ( .A1(n3415), .A2(n3416), .ZN(n3500) );
  AND2_X1 U3496 ( .A1(n3503), .A2(n3504), .ZN(n3416) );
  NAND2_X1 U3497 ( .A1(n3505), .A2(n3270), .ZN(n3504) );
  NOR2_X1 U3498 ( .A1(n3506), .A2(n2394), .ZN(n3505) );
  NOR2_X1 U3499 ( .A1(n3410), .A2(n3412), .ZN(n3506) );
  NAND2_X1 U3500 ( .A1(n3410), .A2(n3412), .ZN(n3503) );
  NAND2_X1 U3501 ( .A1(n3507), .A2(n3508), .ZN(n3412) );
  NAND2_X1 U3502 ( .A1(n3509), .A2(n3270), .ZN(n3508) );
  NOR2_X1 U3503 ( .A1(n3510), .A2(n2291), .ZN(n3509) );
  NOR2_X1 U3504 ( .A1(n3406), .A2(n3408), .ZN(n3510) );
  NAND2_X1 U3505 ( .A1(n3406), .A2(n3408), .ZN(n3507) );
  NAND2_X1 U3506 ( .A1(n3511), .A2(n3512), .ZN(n3408) );
  NAND2_X1 U3507 ( .A1(n3513), .A2(n3270), .ZN(n3512) );
  NOR2_X1 U3508 ( .A1(n3514), .A2(n2187), .ZN(n3513) );
  NOR2_X1 U3509 ( .A1(n3403), .A2(n3405), .ZN(n3514) );
  NAND2_X1 U3510 ( .A1(n3403), .A2(n3405), .ZN(n3511) );
  NAND2_X1 U3511 ( .A1(n3515), .A2(n3516), .ZN(n3405) );
  NAND2_X1 U3512 ( .A1(n3398), .A2(n3517), .ZN(n3516) );
  NAND2_X1 U3513 ( .A1(n3401), .A2(n3400), .ZN(n3517) );
  NOR2_X1 U3514 ( .A1(n3269), .A2(n2203), .ZN(n3398) );
  OR2_X1 U3515 ( .A1(n3400), .A2(n3401), .ZN(n3515) );
  AND2_X1 U3516 ( .A1(n3518), .A2(n3519), .ZN(n3401) );
  NAND2_X1 U3517 ( .A1(n1918), .A2(n3520), .ZN(n3519) );
  NAND2_X1 U3518 ( .A1(n1953), .A2(n3521), .ZN(n3520) );
  NAND2_X1 U3519 ( .A1(n3522), .A2(n1956), .ZN(n3521) );
  NAND2_X1 U3520 ( .A1(n3523), .A2(n3524), .ZN(n3518) );
  NAND2_X1 U3521 ( .A1(n1959), .A2(n3525), .ZN(n3524) );
  NAND2_X1 U3522 ( .A1(n1961), .A2(n3391), .ZN(n3525) );
  NAND2_X1 U3523 ( .A1(n3526), .A2(n1918), .ZN(n3400) );
  NOR2_X1 U3524 ( .A1(n2306), .A2(n3269), .ZN(n3526) );
  INV_X1 U3525 ( .A(n3270), .ZN(n3269) );
  XOR2_X1 U3526 ( .A(n3527), .B(n3528), .Z(n3270) );
  XOR2_X1 U3527 ( .A(d_4_), .B(c_4_), .Z(n3528) );
  XOR2_X1 U3528 ( .A(n3529), .B(n3530), .Z(n3403) );
  XNOR2_X1 U3529 ( .A(n3531), .B(n3532), .ZN(n3530) );
  NAND2_X1 U3530 ( .A1(n1918), .A2(n3533), .ZN(n3529) );
  XNOR2_X1 U3531 ( .A(n3534), .B(n3535), .ZN(n3406) );
  NAND2_X1 U3532 ( .A1(n3536), .A2(n3537), .ZN(n3534) );
  XNOR2_X1 U3533 ( .A(n3538), .B(n3539), .ZN(n3410) );
  XOR2_X1 U3534 ( .A(n3540), .B(n3541), .Z(n3539) );
  NAND2_X1 U3535 ( .A1(n1918), .A2(n2208), .ZN(n3541) );
  XOR2_X1 U3536 ( .A(n3542), .B(n3543), .Z(n3415) );
  XOR2_X1 U3537 ( .A(n3544), .B(n3545), .Z(n3543) );
  NAND2_X1 U3538 ( .A1(n1918), .A2(n2165), .ZN(n3545) );
  XNOR2_X1 U3539 ( .A(n3546), .B(n3547), .ZN(n3422) );
  XOR2_X1 U3540 ( .A(n3548), .B(n3549), .Z(n3547) );
  NAND2_X1 U3541 ( .A1(n1918), .A2(n2149), .ZN(n3549) );
  XNOR2_X1 U3542 ( .A(n3550), .B(n3551), .ZN(n3426) );
  XOR2_X1 U3543 ( .A(n3552), .B(n3553), .Z(n3551) );
  NAND2_X1 U3544 ( .A1(n1918), .A2(n2927), .ZN(n3553) );
  XNOR2_X1 U3545 ( .A(n3554), .B(n3555), .ZN(n3430) );
  XOR2_X1 U3546 ( .A(n3556), .B(n3557), .Z(n3555) );
  NAND2_X1 U3547 ( .A1(n2133), .A2(n1918), .ZN(n3557) );
  XNOR2_X1 U3548 ( .A(n3558), .B(n3559), .ZN(n3434) );
  XOR2_X1 U3549 ( .A(n3560), .B(n3561), .Z(n3559) );
  NAND2_X1 U3550 ( .A1(n1918), .A2(n2692), .ZN(n3561) );
  XNOR2_X1 U3551 ( .A(n3562), .B(n3563), .ZN(n3438) );
  XOR2_X1 U3552 ( .A(n3564), .B(n3565), .Z(n3563) );
  NAND2_X1 U3553 ( .A1(n1918), .A2(n2117), .ZN(n3565) );
  XNOR2_X1 U3554 ( .A(n3566), .B(n3567), .ZN(n3442) );
  XOR2_X1 U3555 ( .A(n3568), .B(n3569), .Z(n3567) );
  NAND2_X1 U3556 ( .A1(n2459), .A2(n1918), .ZN(n3569) );
  XNOR2_X1 U3557 ( .A(n3570), .B(n3571), .ZN(n3447) );
  NAND2_X1 U3558 ( .A1(n3572), .A2(n3573), .ZN(n3570) );
  XOR2_X1 U3559 ( .A(n3574), .B(n3575), .Z(n3327) );
  XOR2_X1 U3560 ( .A(n3576), .B(n3577), .Z(n3574) );
  NOR2_X1 U3561 ( .A1(n3391), .A2(n2241), .ZN(n3577) );
  NAND2_X1 U3562 ( .A1(n3578), .A2(n3579), .ZN(n1964) );
  NAND2_X1 U3563 ( .A1(n3580), .A2(n3458), .ZN(n3579) );
  INV_X1 U3564 ( .A(n3459), .ZN(n3580) );
  XNOR2_X1 U3565 ( .A(n3581), .B(n3582), .ZN(n3578) );
  NAND2_X1 U3566 ( .A1(n3583), .A2(n3584), .ZN(n1965) );
  AND2_X1 U3567 ( .A1(n2057), .A2(n3458), .ZN(n3584) );
  NAND2_X1 U3568 ( .A1(n3585), .A2(n3586), .ZN(n3458) );
  NAND2_X1 U3569 ( .A1(n3587), .A2(n1918), .ZN(n3586) );
  NOR2_X1 U3570 ( .A1(n3588), .A2(n2026), .ZN(n3587) );
  NOR2_X1 U3571 ( .A1(n3455), .A2(n3454), .ZN(n3588) );
  NAND2_X1 U3572 ( .A1(n3454), .A2(n3455), .ZN(n3585) );
  NAND2_X1 U3573 ( .A1(n3589), .A2(n3590), .ZN(n3455) );
  NAND2_X1 U3574 ( .A1(n3591), .A2(n2095), .ZN(n3590) );
  NOR2_X1 U3575 ( .A1(n3592), .A2(n3391), .ZN(n3591) );
  NOR2_X1 U3576 ( .A1(n3575), .A2(n3576), .ZN(n3592) );
  NAND2_X1 U3577 ( .A1(n3575), .A2(n3576), .ZN(n3589) );
  NAND2_X1 U3578 ( .A1(n3572), .A2(n3593), .ZN(n3576) );
  NAND2_X1 U3579 ( .A1(n3571), .A2(n3573), .ZN(n3593) );
  NAND2_X1 U3580 ( .A1(n3594), .A2(n3595), .ZN(n3573) );
  NAND2_X1 U3581 ( .A1(n1917), .A2(n3392), .ZN(n3595) );
  INV_X1 U3582 ( .A(n3596), .ZN(n3594) );
  XNOR2_X1 U3583 ( .A(n3597), .B(n3598), .ZN(n3571) );
  XNOR2_X1 U3584 ( .A(n3599), .B(n3600), .ZN(n3597) );
  NAND2_X1 U3585 ( .A1(n1917), .A2(n3596), .ZN(n3572) );
  NAND2_X1 U3586 ( .A1(n3601), .A2(n3602), .ZN(n3596) );
  NAND2_X1 U3587 ( .A1(n3603), .A2(n2459), .ZN(n3602) );
  NOR2_X1 U3588 ( .A1(n3604), .A2(n3391), .ZN(n3603) );
  NOR2_X1 U3589 ( .A1(n3566), .A2(n3568), .ZN(n3604) );
  NAND2_X1 U3590 ( .A1(n3566), .A2(n3568), .ZN(n3601) );
  NAND2_X1 U3591 ( .A1(n3605), .A2(n3606), .ZN(n3568) );
  NAND2_X1 U3592 ( .A1(n3607), .A2(n3392), .ZN(n3606) );
  NOR2_X1 U3593 ( .A1(n3608), .A2(n2370), .ZN(n3607) );
  NOR2_X1 U3594 ( .A1(n3564), .A2(n3562), .ZN(n3608) );
  NAND2_X1 U3595 ( .A1(n3562), .A2(n3564), .ZN(n3605) );
  NAND2_X1 U3596 ( .A1(n3609), .A2(n3610), .ZN(n3564) );
  NAND2_X1 U3597 ( .A1(n3611), .A2(n3392), .ZN(n3610) );
  NOR2_X1 U3598 ( .A1(n3612), .A2(n2211), .ZN(n3611) );
  NOR2_X1 U3599 ( .A1(n3558), .A2(n3560), .ZN(n3612) );
  NAND2_X1 U3600 ( .A1(n3558), .A2(n3560), .ZN(n3609) );
  NAND2_X1 U3601 ( .A1(n3613), .A2(n3614), .ZN(n3560) );
  NAND2_X1 U3602 ( .A1(n3615), .A2(n2133), .ZN(n3614) );
  NOR2_X1 U3603 ( .A1(n3616), .A2(n3391), .ZN(n3615) );
  NOR2_X1 U3604 ( .A1(n3556), .A2(n3554), .ZN(n3616) );
  NAND2_X1 U3605 ( .A1(n3554), .A2(n3556), .ZN(n3613) );
  NAND2_X1 U3606 ( .A1(n3617), .A2(n3618), .ZN(n3556) );
  NAND2_X1 U3607 ( .A1(n3619), .A2(n3392), .ZN(n3618) );
  NOR2_X1 U3608 ( .A1(n3620), .A2(n2210), .ZN(n3619) );
  NOR2_X1 U3609 ( .A1(n3550), .A2(n3552), .ZN(n3620) );
  NAND2_X1 U3610 ( .A1(n3550), .A2(n3552), .ZN(n3617) );
  NAND2_X1 U3611 ( .A1(n3621), .A2(n3622), .ZN(n3552) );
  NAND2_X1 U3612 ( .A1(n3623), .A2(n3392), .ZN(n3622) );
  NOR2_X1 U3613 ( .A1(n3624), .A2(n2386), .ZN(n3623) );
  NOR2_X1 U3614 ( .A1(n3548), .A2(n3546), .ZN(n3624) );
  NAND2_X1 U3615 ( .A1(n3546), .A2(n3548), .ZN(n3621) );
  NAND2_X1 U3616 ( .A1(n3625), .A2(n3626), .ZN(n3548) );
  NAND2_X1 U3617 ( .A1(n3627), .A2(n3392), .ZN(n3626) );
  NOR2_X1 U3618 ( .A1(n3628), .A2(n2209), .ZN(n3627) );
  NOR2_X1 U3619 ( .A1(n3496), .A2(n3498), .ZN(n3628) );
  NAND2_X1 U3620 ( .A1(n3496), .A2(n3498), .ZN(n3625) );
  NAND2_X1 U3621 ( .A1(n3629), .A2(n3630), .ZN(n3498) );
  NAND2_X1 U3622 ( .A1(n3631), .A2(n3392), .ZN(n3630) );
  NOR2_X1 U3623 ( .A1(n3632), .A2(n2394), .ZN(n3631) );
  NOR2_X1 U3624 ( .A1(n3544), .A2(n3542), .ZN(n3632) );
  NAND2_X1 U3625 ( .A1(n3542), .A2(n3544), .ZN(n3629) );
  NAND2_X1 U3626 ( .A1(n3633), .A2(n3634), .ZN(n3544) );
  NAND2_X1 U3627 ( .A1(n3635), .A2(n3392), .ZN(n3634) );
  NOR2_X1 U3628 ( .A1(n3636), .A2(n2291), .ZN(n3635) );
  NOR2_X1 U3629 ( .A1(n3540), .A2(n3538), .ZN(n3636) );
  NAND2_X1 U3630 ( .A1(n3538), .A2(n3540), .ZN(n3633) );
  NAND2_X1 U3631 ( .A1(n3536), .A2(n3637), .ZN(n3540) );
  NAND2_X1 U3632 ( .A1(n3535), .A2(n3537), .ZN(n3637) );
  NAND2_X1 U3633 ( .A1(n3638), .A2(n3639), .ZN(n3537) );
  NAND2_X1 U3634 ( .A1(n1918), .A2(n2182), .ZN(n3639) );
  INV_X1 U3635 ( .A(n3640), .ZN(n3638) );
  XOR2_X1 U3636 ( .A(n3641), .B(n3642), .Z(n3535) );
  XNOR2_X1 U3637 ( .A(n3643), .B(n3644), .ZN(n3642) );
  NAND2_X1 U3638 ( .A1(n3523), .A2(n3533), .ZN(n3641) );
  NAND2_X1 U3639 ( .A1(n2182), .A2(n3640), .ZN(n3536) );
  NAND2_X1 U3640 ( .A1(n3645), .A2(n3646), .ZN(n3640) );
  NAND2_X1 U3641 ( .A1(n3647), .A2(n3392), .ZN(n3646) );
  NOR2_X1 U3642 ( .A1(n3648), .A2(n2203), .ZN(n3647) );
  NOR2_X1 U3643 ( .A1(n3531), .A2(n3532), .ZN(n3648) );
  NAND2_X1 U3644 ( .A1(n3531), .A2(n3532), .ZN(n3645) );
  NAND2_X1 U3645 ( .A1(n3649), .A2(n3650), .ZN(n3532) );
  NAND2_X1 U3646 ( .A1(n3523), .A2(n3651), .ZN(n3650) );
  NAND2_X1 U3647 ( .A1(n1953), .A2(n3652), .ZN(n3651) );
  NAND2_X1 U3648 ( .A1(n1956), .A2(n3653), .ZN(n3652) );
  NAND2_X1 U3649 ( .A1(n3654), .A2(n3655), .ZN(n3649) );
  NAND2_X1 U3650 ( .A1(n1959), .A2(n3656), .ZN(n3655) );
  NAND2_X1 U3651 ( .A1(n1961), .A2(n3522), .ZN(n3656) );
  AND2_X1 U3652 ( .A1(n3657), .A2(n3523), .ZN(n3531) );
  NOR2_X1 U3653 ( .A1(n2306), .A2(n3391), .ZN(n3657) );
  INV_X1 U3654 ( .A(n3392), .ZN(n3391) );
  XOR2_X1 U3655 ( .A(n3658), .B(n3659), .Z(n3392) );
  XOR2_X1 U3656 ( .A(d_3_), .B(c_3_), .Z(n3659) );
  XNOR2_X1 U3657 ( .A(n3660), .B(n3661), .ZN(n3538) );
  NAND2_X1 U3658 ( .A1(n3662), .A2(n3663), .ZN(n3660) );
  XOR2_X1 U3659 ( .A(n3664), .B(n3665), .Z(n3542) );
  XOR2_X1 U3660 ( .A(n3666), .B(n3667), .Z(n3664) );
  XNOR2_X1 U3661 ( .A(n3668), .B(n3669), .ZN(n3496) );
  NAND2_X1 U3662 ( .A1(n3670), .A2(n3671), .ZN(n3668) );
  XOR2_X1 U3663 ( .A(n3672), .B(n3673), .Z(n3546) );
  XOR2_X1 U3664 ( .A(n3674), .B(n3675), .Z(n3672) );
  XNOR2_X1 U3665 ( .A(n3676), .B(n3677), .ZN(n3550) );
  NAND2_X1 U3666 ( .A1(n3678), .A2(n3679), .ZN(n3676) );
  XOR2_X1 U3667 ( .A(n3680), .B(n3681), .Z(n3554) );
  XOR2_X1 U3668 ( .A(n3682), .B(n3683), .Z(n3680) );
  XNOR2_X1 U3669 ( .A(n3684), .B(n3685), .ZN(n3558) );
  NAND2_X1 U3670 ( .A1(n3686), .A2(n3687), .ZN(n3684) );
  XOR2_X1 U3671 ( .A(n3688), .B(n3689), .Z(n3562) );
  XOR2_X1 U3672 ( .A(n3690), .B(n3691), .Z(n3688) );
  XNOR2_X1 U3673 ( .A(n3692), .B(n3693), .ZN(n3566) );
  NAND2_X1 U3674 ( .A1(n3694), .A2(n3695), .ZN(n3692) );
  XNOR2_X1 U3675 ( .A(n3696), .B(n3697), .ZN(n3575) );
  NAND2_X1 U3676 ( .A1(n3698), .A2(n3699), .ZN(n3696) );
  XNOR2_X1 U3677 ( .A(n3700), .B(n3701), .ZN(n3454) );
  XNOR2_X1 U3678 ( .A(n3702), .B(n3703), .ZN(n3700) );
  NOR2_X1 U3679 ( .A1(n3704), .A2(n3459), .ZN(n3583) );
  XOR2_X1 U3680 ( .A(n3705), .B(n3706), .Z(n3459) );
  NAND2_X1 U3681 ( .A1(n3707), .A2(n3708), .ZN(n3705) );
  NOR2_X1 U3682 ( .A1(n3582), .A2(n3581), .ZN(n3704) );
  AND2_X1 U3683 ( .A1(n3709), .A2(n3710), .ZN(n2009) );
  NOR2_X1 U3684 ( .A1(n3711), .A2(n2026), .ZN(n3710) );
  NOR2_X1 U3685 ( .A1(n2054), .A2(n2057), .ZN(n3709) );
  NAND2_X1 U3686 ( .A1(n3582), .A2(n3581), .ZN(n2057) );
  NAND2_X1 U3687 ( .A1(n3707), .A2(n3712), .ZN(n3581) );
  NAND2_X1 U3688 ( .A1(n3706), .A2(n3708), .ZN(n3712) );
  NAND2_X1 U3689 ( .A1(n3713), .A2(n3714), .ZN(n3708) );
  NAND2_X1 U3690 ( .A1(n3523), .A2(n2053), .ZN(n3714) );
  INV_X1 U3691 ( .A(n3715), .ZN(n3713) );
  XOR2_X1 U3692 ( .A(n3716), .B(n3717), .Z(n3706) );
  NOR2_X1 U3693 ( .A1(n3711), .A2(n2362), .ZN(n3717) );
  XOR2_X1 U3694 ( .A(n3718), .B(n3719), .Z(n3716) );
  NAND2_X1 U3695 ( .A1(n2053), .A2(n3715), .ZN(n3707) );
  NAND2_X1 U3696 ( .A1(n3720), .A2(n3721), .ZN(n3715) );
  NAND2_X1 U3697 ( .A1(n3703), .A2(n3722), .ZN(n3721) );
  NAND2_X1 U3698 ( .A1(n3702), .A2(n3701), .ZN(n3722) );
  NOR2_X1 U3699 ( .A1(n2241), .A2(n3522), .ZN(n3703) );
  OR2_X1 U3700 ( .A1(n3701), .A2(n3702), .ZN(n3720) );
  AND2_X1 U3701 ( .A1(n3698), .A2(n3723), .ZN(n3702) );
  NAND2_X1 U3702 ( .A1(n3697), .A2(n3699), .ZN(n3723) );
  NAND2_X1 U3703 ( .A1(n3724), .A2(n3725), .ZN(n3699) );
  NAND2_X1 U3704 ( .A1(n1917), .A2(n3523), .ZN(n3725) );
  INV_X1 U3705 ( .A(n3726), .ZN(n3724) );
  XOR2_X1 U3706 ( .A(n3727), .B(n3728), .Z(n3697) );
  NOR2_X1 U3707 ( .A1(n3653), .A2(n2212), .ZN(n3728) );
  XOR2_X1 U3708 ( .A(n3729), .B(n3730), .Z(n3727) );
  NAND2_X1 U3709 ( .A1(n1917), .A2(n3726), .ZN(n3698) );
  NAND2_X1 U3710 ( .A1(n3731), .A2(n3732), .ZN(n3726) );
  NAND2_X1 U3711 ( .A1(n3600), .A2(n3733), .ZN(n3732) );
  NAND2_X1 U3712 ( .A1(n3599), .A2(n3598), .ZN(n3733) );
  NOR2_X1 U3713 ( .A1(n2212), .A2(n3522), .ZN(n3600) );
  OR2_X1 U3714 ( .A1(n3598), .A2(n3599), .ZN(n3731) );
  AND2_X1 U3715 ( .A1(n3694), .A2(n3734), .ZN(n3599) );
  NAND2_X1 U3716 ( .A1(n3693), .A2(n3695), .ZN(n3734) );
  NAND2_X1 U3717 ( .A1(n3735), .A2(n3736), .ZN(n3695) );
  NAND2_X1 U3718 ( .A1(n3523), .A2(n2117), .ZN(n3736) );
  INV_X1 U3719 ( .A(n3737), .ZN(n3735) );
  XOR2_X1 U3720 ( .A(n3738), .B(n3739), .Z(n3693) );
  NOR2_X1 U3721 ( .A1(n2211), .A2(n3653), .ZN(n3739) );
  XOR2_X1 U3722 ( .A(n3740), .B(n3741), .Z(n3738) );
  NAND2_X1 U3723 ( .A1(n2117), .A2(n3737), .ZN(n3694) );
  NAND2_X1 U3724 ( .A1(n3742), .A2(n3743), .ZN(n3737) );
  NAND2_X1 U3725 ( .A1(n3691), .A2(n3744), .ZN(n3743) );
  OR2_X1 U3726 ( .A1(n3690), .A2(n3689), .ZN(n3744) );
  NOR2_X1 U3727 ( .A1(n3522), .A2(n2211), .ZN(n3691) );
  NAND2_X1 U3728 ( .A1(n3689), .A2(n3690), .ZN(n3742) );
  NAND2_X1 U3729 ( .A1(n3686), .A2(n3745), .ZN(n3690) );
  NAND2_X1 U3730 ( .A1(n3685), .A2(n3687), .ZN(n3745) );
  NAND2_X1 U3731 ( .A1(n3746), .A2(n3747), .ZN(n3687) );
  NAND2_X1 U3732 ( .A1(n2133), .A2(n3523), .ZN(n3747) );
  INV_X1 U3733 ( .A(n3748), .ZN(n3746) );
  XOR2_X1 U3734 ( .A(n3749), .B(n3750), .Z(n3685) );
  NOR2_X1 U3735 ( .A1(n2210), .A2(n3653), .ZN(n3750) );
  XOR2_X1 U3736 ( .A(n3751), .B(n3752), .Z(n3749) );
  NAND2_X1 U3737 ( .A1(n2133), .A2(n3748), .ZN(n3686) );
  NAND2_X1 U3738 ( .A1(n3753), .A2(n3754), .ZN(n3748) );
  NAND2_X1 U3739 ( .A1(n3683), .A2(n3755), .ZN(n3754) );
  OR2_X1 U3740 ( .A1(n3682), .A2(n3681), .ZN(n3755) );
  NOR2_X1 U3741 ( .A1(n3522), .A2(n2210), .ZN(n3683) );
  NAND2_X1 U3742 ( .A1(n3681), .A2(n3682), .ZN(n3753) );
  NAND2_X1 U3743 ( .A1(n3678), .A2(n3756), .ZN(n3682) );
  NAND2_X1 U3744 ( .A1(n3677), .A2(n3679), .ZN(n3756) );
  NAND2_X1 U3745 ( .A1(n3757), .A2(n3758), .ZN(n3679) );
  NAND2_X1 U3746 ( .A1(n3523), .A2(n2149), .ZN(n3758) );
  INV_X1 U3747 ( .A(n3759), .ZN(n3757) );
  XOR2_X1 U3748 ( .A(n3760), .B(n3761), .Z(n3677) );
  NOR2_X1 U3749 ( .A1(n2209), .A2(n3653), .ZN(n3761) );
  XOR2_X1 U3750 ( .A(n3762), .B(n3763), .Z(n3760) );
  NAND2_X1 U3751 ( .A1(n2149), .A2(n3759), .ZN(n3678) );
  NAND2_X1 U3752 ( .A1(n3764), .A2(n3765), .ZN(n3759) );
  NAND2_X1 U3753 ( .A1(n3675), .A2(n3766), .ZN(n3765) );
  OR2_X1 U3754 ( .A1(n3674), .A2(n3673), .ZN(n3766) );
  NOR2_X1 U3755 ( .A1(n3522), .A2(n2209), .ZN(n3675) );
  NAND2_X1 U3756 ( .A1(n3673), .A2(n3674), .ZN(n3764) );
  NAND2_X1 U3757 ( .A1(n3670), .A2(n3767), .ZN(n3674) );
  NAND2_X1 U3758 ( .A1(n3669), .A2(n3671), .ZN(n3767) );
  NAND2_X1 U3759 ( .A1(n3768), .A2(n3769), .ZN(n3671) );
  NAND2_X1 U3760 ( .A1(n3523), .A2(n2165), .ZN(n3769) );
  INV_X1 U3761 ( .A(n3770), .ZN(n3768) );
  XOR2_X1 U3762 ( .A(n3771), .B(n3772), .Z(n3669) );
  XNOR2_X1 U3763 ( .A(n3773), .B(n3774), .ZN(n3772) );
  NAND2_X1 U3764 ( .A1(n3654), .A2(n2208), .ZN(n3771) );
  NAND2_X1 U3765 ( .A1(n2165), .A2(n3770), .ZN(n3670) );
  NAND2_X1 U3766 ( .A1(n3775), .A2(n3776), .ZN(n3770) );
  NAND2_X1 U3767 ( .A1(n3667), .A2(n3777), .ZN(n3776) );
  OR2_X1 U3768 ( .A1(n3666), .A2(n3665), .ZN(n3777) );
  NOR2_X1 U3769 ( .A1(n3522), .A2(n2291), .ZN(n3667) );
  NAND2_X1 U3770 ( .A1(n3665), .A2(n3666), .ZN(n3775) );
  NAND2_X1 U3771 ( .A1(n3662), .A2(n3778), .ZN(n3666) );
  NAND2_X1 U3772 ( .A1(n3661), .A2(n3663), .ZN(n3778) );
  NAND2_X1 U3773 ( .A1(n3779), .A2(n3780), .ZN(n3663) );
  NAND2_X1 U3774 ( .A1(n3523), .A2(n2182), .ZN(n3780) );
  INV_X1 U3775 ( .A(n3781), .ZN(n3779) );
  XNOR2_X1 U3776 ( .A(n3782), .B(n3783), .ZN(n3661) );
  NAND2_X1 U3777 ( .A1(n3784), .A2(n3785), .ZN(n3782) );
  NAND2_X1 U3778 ( .A1(n2182), .A2(n3781), .ZN(n3662) );
  NAND2_X1 U3779 ( .A1(n3786), .A2(n3787), .ZN(n3781) );
  NAND2_X1 U3780 ( .A1(n3788), .A2(n3523), .ZN(n3787) );
  NOR2_X1 U3781 ( .A1(n3789), .A2(n2203), .ZN(n3788) );
  NOR2_X1 U3782 ( .A1(n3644), .A2(n3643), .ZN(n3789) );
  NAND2_X1 U3783 ( .A1(n3644), .A2(n3643), .ZN(n3786) );
  NAND2_X1 U3784 ( .A1(n3790), .A2(n3791), .ZN(n3643) );
  NAND2_X1 U3785 ( .A1(n3792), .A2(n3654), .ZN(n3791) );
  NOR2_X1 U3786 ( .A1(n3793), .A2(n2196), .ZN(n3792) );
  NOR2_X1 U3787 ( .A1(n2197), .A2(n3711), .ZN(n3793) );
  INV_X1 U3788 ( .A(n1953), .ZN(n2197) );
  NAND2_X1 U3789 ( .A1(n1956), .A2(n1947), .ZN(n1953) );
  NAND2_X1 U3790 ( .A1(n3794), .A2(n1961), .ZN(n3790) );
  NOR2_X1 U3791 ( .A1(n3795), .A2(n3711), .ZN(n3794) );
  NOR2_X1 U3792 ( .A1(n2202), .A2(n3653), .ZN(n3795) );
  INV_X1 U3793 ( .A(n1959), .ZN(n2202) );
  NAND2_X1 U3794 ( .A1(n2196), .A2(n1961), .ZN(n1959) );
  AND2_X1 U3795 ( .A1(n3796), .A2(n3654), .ZN(n3644) );
  NOR2_X1 U3796 ( .A1(n2306), .A2(n3522), .ZN(n3796) );
  INV_X1 U3797 ( .A(n3523), .ZN(n3522) );
  XOR2_X1 U3798 ( .A(d_2_), .B(c_2_), .Z(n3798) );
  NAND2_X1 U3799 ( .A1(n1961), .A2(n1956), .ZN(n2306) );
  INV_X1 U3800 ( .A(n2196), .ZN(n1956) );
  INV_X1 U3801 ( .A(n1947), .ZN(n1961) );
  XOR2_X1 U3802 ( .A(n3799), .B(n3800), .Z(n3665) );
  XOR2_X1 U3803 ( .A(n3801), .B(n3802), .Z(n3799) );
  XNOR2_X1 U3804 ( .A(n3803), .B(n3804), .ZN(n3673) );
  XNOR2_X1 U3805 ( .A(n3805), .B(n3806), .ZN(n3804) );
  XNOR2_X1 U3806 ( .A(n3807), .B(n3808), .ZN(n3681) );
  XOR2_X1 U3807 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR2_X1 U3808 ( .A(n3811), .B(n3812), .Z(n3689) );
  XOR2_X1 U3809 ( .A(n3813), .B(n3814), .Z(n3811) );
  XOR2_X1 U3810 ( .A(n3815), .B(n3816), .Z(n3598) );
  XOR2_X1 U3811 ( .A(n3817), .B(n3818), .Z(n3816) );
  XNOR2_X1 U3812 ( .A(n3819), .B(n3820), .ZN(n3701) );
  XOR2_X1 U3813 ( .A(n3821), .B(n3822), .Z(n3819) );
  INV_X1 U3814 ( .A(n2026), .ZN(n2053) );
  XOR2_X1 U3815 ( .A(n3823), .B(n3824), .Z(n3582) );
  NOR2_X1 U3816 ( .A1(n3825), .A2(n3826), .ZN(n3824) );
  INV_X1 U3817 ( .A(n3827), .ZN(n3826) );
  NOR2_X1 U3818 ( .A1(n3828), .A2(n3829), .ZN(n3825) );
  NAND2_X1 U3819 ( .A1(n3827), .A2(n3830), .ZN(n2054) );
  NAND2_X1 U3820 ( .A1(n3831), .A2(n3823), .ZN(n3830) );
  NAND2_X1 U3821 ( .A1(n3832), .A2(n3833), .ZN(n3823) );
  NAND2_X1 U3822 ( .A1(n3834), .A2(n2101), .ZN(n3833) );
  NOR2_X1 U3823 ( .A1(n3835), .A2(n3711), .ZN(n3834) );
  NOR2_X1 U3824 ( .A1(n3718), .A2(n3719), .ZN(n3835) );
  NAND2_X1 U3825 ( .A1(n3718), .A2(n3719), .ZN(n3832) );
  NAND2_X1 U3826 ( .A1(n3836), .A2(n3837), .ZN(n3719) );
  NAND2_X1 U3827 ( .A1(n3820), .A2(n3838), .ZN(n3837) );
  OR2_X1 U3828 ( .A1(n3821), .A2(n3822), .ZN(n3838) );
  NOR2_X1 U3829 ( .A1(n2362), .A2(n3653), .ZN(n3820) );
  INV_X1 U3830 ( .A(n2101), .ZN(n2362) );
  XOR2_X1 U3831 ( .A(n3839), .B(n3840), .Z(n2101) );
  XOR2_X1 U3832 ( .A(b_2_), .B(a_2_), .Z(n3840) );
  NAND2_X1 U3833 ( .A1(n3822), .A2(n3821), .ZN(n3836) );
  NAND2_X1 U3834 ( .A1(n3841), .A2(n3842), .ZN(n3821) );
  NAND2_X1 U3835 ( .A1(n3843), .A2(n2459), .ZN(n3842) );
  NOR2_X1 U3836 ( .A1(n3844), .A2(n3653), .ZN(n3843) );
  NOR2_X1 U3837 ( .A1(n3730), .A2(n3729), .ZN(n3844) );
  NAND2_X1 U3838 ( .A1(n3730), .A2(n3729), .ZN(n3841) );
  NAND2_X1 U3839 ( .A1(n3845), .A2(n3846), .ZN(n3729) );
  NAND2_X1 U3840 ( .A1(n3815), .A2(n3847), .ZN(n3846) );
  NAND2_X1 U3841 ( .A1(n3818), .A2(n3848), .ZN(n3847) );
  INV_X1 U3842 ( .A(n3849), .ZN(n3818) );
  NOR2_X1 U3843 ( .A1(n3653), .A2(n2370), .ZN(n3815) );
  NAND2_X1 U3844 ( .A1(n3817), .A2(n3849), .ZN(n3845) );
  NAND2_X1 U3845 ( .A1(n3850), .A2(n3851), .ZN(n3849) );
  NAND2_X1 U3846 ( .A1(n3852), .A2(n3654), .ZN(n3851) );
  NOR2_X1 U3847 ( .A1(n3853), .A2(n2211), .ZN(n3852) );
  INV_X1 U3848 ( .A(n2692), .ZN(n2211) );
  NOR2_X1 U3849 ( .A1(n3740), .A2(n3741), .ZN(n3853) );
  NAND2_X1 U3850 ( .A1(n3740), .A2(n3741), .ZN(n3850) );
  NAND2_X1 U3851 ( .A1(n3854), .A2(n3855), .ZN(n3741) );
  NAND2_X1 U3852 ( .A1(n3812), .A2(n3856), .ZN(n3855) );
  OR2_X1 U3853 ( .A1(n3813), .A2(n3814), .ZN(n3856) );
  NOR2_X1 U3854 ( .A1(n3653), .A2(n2378), .ZN(n3812) );
  NAND2_X1 U3855 ( .A1(n3814), .A2(n3813), .ZN(n3854) );
  NAND2_X1 U3856 ( .A1(n3857), .A2(n3858), .ZN(n3813) );
  NAND2_X1 U3857 ( .A1(n3859), .A2(n3654), .ZN(n3858) );
  NOR2_X1 U3858 ( .A1(n3860), .A2(n2210), .ZN(n3859) );
  NOR2_X1 U3859 ( .A1(n3752), .A2(n3751), .ZN(n3860) );
  NAND2_X1 U3860 ( .A1(n3752), .A2(n3751), .ZN(n3857) );
  NAND2_X1 U3861 ( .A1(n3861), .A2(n3862), .ZN(n3751) );
  NAND2_X1 U3862 ( .A1(n3807), .A2(n3863), .ZN(n3862) );
  NAND2_X1 U3863 ( .A1(n3810), .A2(n3864), .ZN(n3863) );
  INV_X1 U3864 ( .A(n3865), .ZN(n3810) );
  NOR2_X1 U3865 ( .A1(n3653), .A2(n2386), .ZN(n3807) );
  NAND2_X1 U3866 ( .A1(n3809), .A2(n3865), .ZN(n3861) );
  NAND2_X1 U3867 ( .A1(n3866), .A2(n3867), .ZN(n3865) );
  NAND2_X1 U3868 ( .A1(n3868), .A2(n3654), .ZN(n3867) );
  NOR2_X1 U3869 ( .A1(n3869), .A2(n2209), .ZN(n3868) );
  INV_X1 U3870 ( .A(n3166), .ZN(n2209) );
  NOR2_X1 U3871 ( .A1(n3762), .A2(n3763), .ZN(n3869) );
  NAND2_X1 U3872 ( .A1(n3762), .A2(n3763), .ZN(n3866) );
  NAND2_X1 U3873 ( .A1(n3870), .A2(n3871), .ZN(n3763) );
  NAND2_X1 U3874 ( .A1(n3803), .A2(n3872), .ZN(n3871) );
  OR2_X1 U3875 ( .A1(n3806), .A2(n3805), .ZN(n3872) );
  NOR2_X1 U3876 ( .A1(n3653), .A2(n2394), .ZN(n3803) );
  NAND2_X1 U3877 ( .A1(n3805), .A2(n3806), .ZN(n3870) );
  NAND2_X1 U3878 ( .A1(n3873), .A2(n3874), .ZN(n3806) );
  NAND2_X1 U3879 ( .A1(n3875), .A2(n3654), .ZN(n3874) );
  NOR2_X1 U3880 ( .A1(n3876), .A2(n2291), .ZN(n3875) );
  NOR2_X1 U3881 ( .A1(n3774), .A2(n3773), .ZN(n3876) );
  NAND2_X1 U3882 ( .A1(n3774), .A2(n3773), .ZN(n3873) );
  NAND2_X1 U3883 ( .A1(n3877), .A2(n3878), .ZN(n3773) );
  NAND2_X1 U3884 ( .A1(n3800), .A2(n3879), .ZN(n3878) );
  OR2_X1 U3885 ( .A1(n3801), .A2(n3802), .ZN(n3879) );
  NOR2_X1 U3886 ( .A1(n3653), .A2(n2187), .ZN(n3800) );
  NAND2_X1 U3887 ( .A1(n3802), .A2(n3801), .ZN(n3877) );
  NAND2_X1 U3888 ( .A1(n3880), .A2(n3785), .ZN(n3801) );
  NAND2_X1 U3889 ( .A1(n3881), .A2(n3784), .ZN(n3785) );
  NOR2_X1 U3890 ( .A1(n1947), .A2(n3653), .ZN(n3881) );
  NAND2_X1 U3891 ( .A1(n3882), .A2(n3883), .ZN(n1947) );
  OR2_X1 U3892 ( .A1(b_15_), .A2(a_15_), .ZN(n3882) );
  NAND2_X1 U3893 ( .A1(n3783), .A2(n3784), .ZN(n3880) );
  NOR2_X1 U3894 ( .A1(n2196), .A2(n3711), .ZN(n3784) );
  XOR2_X1 U3895 ( .A(n3883), .B(n3884), .Z(n2196) );
  XOR2_X1 U3896 ( .A(b_14_), .B(a_14_), .Z(n3884) );
  NOR2_X1 U3897 ( .A1(n3653), .A2(n2203), .ZN(n3783) );
  NOR2_X1 U3898 ( .A1(n2203), .A2(n3711), .ZN(n3802) );
  INV_X1 U3899 ( .A(n3533), .ZN(n2203) );
  XOR2_X1 U3900 ( .A(n3885), .B(n3886), .Z(n3533) );
  XOR2_X1 U3901 ( .A(b_13_), .B(a_13_), .Z(n3886) );
  NOR2_X1 U3902 ( .A1(n2187), .A2(n3711), .ZN(n3774) );
  INV_X1 U3903 ( .A(n2182), .ZN(n2187) );
  XNOR2_X1 U3904 ( .A(a_12_), .B(b_12_), .ZN(n3887) );
  NOR2_X1 U3905 ( .A1(n2291), .A2(n3711), .ZN(n3805) );
  INV_X1 U3906 ( .A(n2208), .ZN(n2291) );
  XOR2_X1 U3907 ( .A(n3889), .B(n3890), .Z(n2208) );
  XOR2_X1 U3908 ( .A(b_11_), .B(a_11_), .Z(n3890) );
  NOR2_X1 U3909 ( .A1(n2394), .A2(n3711), .ZN(n3762) );
  INV_X1 U3910 ( .A(n2165), .ZN(n2394) );
  XOR2_X1 U3911 ( .A(b_10_), .B(a_10_), .Z(n3892) );
  INV_X1 U3912 ( .A(n3864), .ZN(n3809) );
  NAND2_X1 U3913 ( .A1(n3166), .A2(n2059), .ZN(n3864) );
  XOR2_X1 U3914 ( .A(n3893), .B(n3894), .Z(n3166) );
  XOR2_X1 U3915 ( .A(b_9_), .B(a_9_), .Z(n3894) );
  NOR2_X1 U3916 ( .A1(n2386), .A2(n3711), .ZN(n3752) );
  INV_X1 U3917 ( .A(n2149), .ZN(n2386) );
  XOR2_X1 U3918 ( .A(b_8_), .B(a_8_), .Z(n3896) );
  NOR2_X1 U3919 ( .A1(n2210), .A2(n3711), .ZN(n3814) );
  INV_X1 U3920 ( .A(n2927), .ZN(n2210) );
  XOR2_X1 U3921 ( .A(n3897), .B(n3898), .Z(n2927) );
  XOR2_X1 U3922 ( .A(b_7_), .B(a_7_), .Z(n3898) );
  NOR2_X1 U3923 ( .A1(n2378), .A2(n3711), .ZN(n3740) );
  INV_X1 U3924 ( .A(n2133), .ZN(n2378) );
  XOR2_X1 U3925 ( .A(b_6_), .B(a_6_), .Z(n3900) );
  INV_X1 U3926 ( .A(n3848), .ZN(n3817) );
  NAND2_X1 U3927 ( .A1(n2692), .A2(n2059), .ZN(n3848) );
  INV_X1 U3928 ( .A(n3711), .ZN(n2059) );
  XOR2_X1 U3929 ( .A(n3901), .B(n3902), .Z(n2692) );
  XOR2_X1 U3930 ( .A(b_5_), .B(a_5_), .Z(n3902) );
  NOR2_X1 U3931 ( .A1(n2370), .A2(n3711), .ZN(n3730) );
  INV_X1 U3932 ( .A(n2117), .ZN(n2370) );
  XOR2_X1 U3933 ( .A(b_4_), .B(a_4_), .Z(n3904) );
  NOR2_X1 U3934 ( .A1(n2212), .A2(n3711), .ZN(n3822) );
  INV_X1 U3935 ( .A(n2459), .ZN(n2212) );
  XOR2_X1 U3936 ( .A(b_3_), .B(a_3_), .Z(n3906) );
  NOR2_X1 U3937 ( .A1(n2241), .A2(n3653), .ZN(n3718) );
  OR2_X1 U3938 ( .A1(n2095), .A2(n3828), .ZN(n3831) );
  NAND2_X1 U3939 ( .A1(n3829), .A2(n3828), .ZN(n3827) );
  NOR2_X1 U3940 ( .A1(n3653), .A2(n2026), .ZN(n3828) );
  XOR2_X1 U3941 ( .A(b_0_), .B(a_0_), .Z(n3908) );
  NAND2_X1 U3942 ( .A1(n3909), .A2(n3910), .ZN(n3907) );
  NAND2_X1 U3943 ( .A1(n3911), .A2(n3912), .ZN(n3910) );
  INV_X1 U3944 ( .A(b_1_), .ZN(n3912) );
  NAND2_X1 U3945 ( .A1(a_1_), .A2(n3913), .ZN(n3911) );
  OR2_X1 U3946 ( .A1(n3913), .A2(a_1_), .ZN(n3909) );
  INV_X1 U3947 ( .A(n3654), .ZN(n3653) );
  XOR2_X1 U3948 ( .A(n3914), .B(n3915), .Z(n3654) );
  XOR2_X1 U3949 ( .A(d_1_), .B(c_1_), .Z(n3915) );
  NOR2_X1 U3950 ( .A1(n3711), .A2(n2241), .ZN(n3829) );
  INV_X1 U3951 ( .A(n2095), .ZN(n2241) );
  XOR2_X1 U3952 ( .A(b_1_), .B(a_1_), .Z(n3916) );
  NAND2_X1 U3953 ( .A1(n3917), .A2(n3918), .ZN(n3913) );
  NAND2_X1 U3954 ( .A1(b_2_), .A2(n3919), .ZN(n3918) );
  OR2_X1 U3955 ( .A1(n3839), .A2(a_2_), .ZN(n3919) );
  NAND2_X1 U3956 ( .A1(a_2_), .A2(n3839), .ZN(n3917) );
  NAND2_X1 U3957 ( .A1(n3920), .A2(n3921), .ZN(n3839) );
  NAND2_X1 U3958 ( .A1(b_3_), .A2(n3922), .ZN(n3921) );
  OR2_X1 U3959 ( .A1(n3905), .A2(a_3_), .ZN(n3922) );
  NAND2_X1 U3960 ( .A1(a_3_), .A2(n3905), .ZN(n3920) );
  NAND2_X1 U3961 ( .A1(n3923), .A2(n3924), .ZN(n3905) );
  NAND2_X1 U3962 ( .A1(b_4_), .A2(n3925), .ZN(n3924) );
  OR2_X1 U3963 ( .A1(n3903), .A2(a_4_), .ZN(n3925) );
  NAND2_X1 U3964 ( .A1(a_4_), .A2(n3903), .ZN(n3923) );
  NAND2_X1 U3965 ( .A1(n3926), .A2(n3927), .ZN(n3903) );
  NAND2_X1 U3966 ( .A1(b_5_), .A2(n3928), .ZN(n3927) );
  OR2_X1 U3967 ( .A1(n3901), .A2(a_5_), .ZN(n3928) );
  NAND2_X1 U3968 ( .A1(a_5_), .A2(n3901), .ZN(n3926) );
  NAND2_X1 U3969 ( .A1(n3929), .A2(n3930), .ZN(n3901) );
  NAND2_X1 U3970 ( .A1(b_6_), .A2(n3931), .ZN(n3930) );
  OR2_X1 U3971 ( .A1(n3899), .A2(a_6_), .ZN(n3931) );
  NAND2_X1 U3972 ( .A1(a_6_), .A2(n3899), .ZN(n3929) );
  NAND2_X1 U3973 ( .A1(n3932), .A2(n3933), .ZN(n3899) );
  NAND2_X1 U3974 ( .A1(b_7_), .A2(n3934), .ZN(n3933) );
  OR2_X1 U3975 ( .A1(n3897), .A2(a_7_), .ZN(n3934) );
  NAND2_X1 U3976 ( .A1(a_7_), .A2(n3897), .ZN(n3932) );
  NAND2_X1 U3977 ( .A1(n3935), .A2(n3936), .ZN(n3897) );
  NAND2_X1 U3978 ( .A1(b_8_), .A2(n3937), .ZN(n3936) );
  OR2_X1 U3979 ( .A1(n3895), .A2(a_8_), .ZN(n3937) );
  NAND2_X1 U3980 ( .A1(a_8_), .A2(n3895), .ZN(n3935) );
  NAND2_X1 U3981 ( .A1(n3938), .A2(n3939), .ZN(n3895) );
  NAND2_X1 U3982 ( .A1(b_9_), .A2(n3940), .ZN(n3939) );
  OR2_X1 U3983 ( .A1(n3893), .A2(a_9_), .ZN(n3940) );
  NAND2_X1 U3984 ( .A1(a_9_), .A2(n3893), .ZN(n3938) );
  NAND2_X1 U3985 ( .A1(n3941), .A2(n3942), .ZN(n3893) );
  NAND2_X1 U3986 ( .A1(b_10_), .A2(n3943), .ZN(n3942) );
  OR2_X1 U3987 ( .A1(n3891), .A2(a_10_), .ZN(n3943) );
  NAND2_X1 U3988 ( .A1(a_10_), .A2(n3891), .ZN(n3941) );
  NAND2_X1 U3989 ( .A1(n3944), .A2(n3945), .ZN(n3891) );
  NAND2_X1 U3990 ( .A1(b_11_), .A2(n3946), .ZN(n3945) );
  OR2_X1 U3991 ( .A1(n3889), .A2(a_11_), .ZN(n3946) );
  NAND2_X1 U3992 ( .A1(a_11_), .A2(n3889), .ZN(n3944) );
  NAND2_X1 U3993 ( .A1(n3947), .A2(n3948), .ZN(n3889) );
  NAND2_X1 U3994 ( .A1(b_12_), .A2(n3949), .ZN(n3948) );
  OR2_X1 U3995 ( .A1(n3888), .A2(a_12_), .ZN(n3949) );
  NAND2_X1 U3996 ( .A1(a_12_), .A2(n3888), .ZN(n3947) );
  NAND2_X1 U3997 ( .A1(n3950), .A2(n3951), .ZN(n3888) );
  NAND2_X1 U3998 ( .A1(b_13_), .A2(n3952), .ZN(n3951) );
  OR2_X1 U3999 ( .A1(n3885), .A2(a_13_), .ZN(n3952) );
  NAND2_X1 U4000 ( .A1(a_13_), .A2(n3885), .ZN(n3950) );
  NAND2_X1 U4001 ( .A1(n3953), .A2(n3954), .ZN(n3885) );
  NAND2_X1 U4002 ( .A1(b_14_), .A2(n3955), .ZN(n3954) );
  OR2_X1 U4003 ( .A1(a_14_), .A2(n3956), .ZN(n3955) );
  NAND2_X1 U4004 ( .A1(a_14_), .A2(n3956), .ZN(n3953) );
  INV_X1 U4005 ( .A(n3883), .ZN(n3956) );
  NAND2_X1 U4006 ( .A1(b_15_), .A2(a_15_), .ZN(n3883) );
  XOR2_X1 U4007 ( .A(d_0_), .B(c_0_), .Z(n3958) );
  NAND2_X1 U4008 ( .A1(n3959), .A2(n3960), .ZN(n3957) );
  NAND2_X1 U4009 ( .A1(n3961), .A2(n3962), .ZN(n3960) );
  INV_X1 U4010 ( .A(d_1_), .ZN(n3962) );
  NAND2_X1 U4011 ( .A1(c_1_), .A2(n3914), .ZN(n3961) );
  OR2_X1 U4012 ( .A1(n3914), .A2(c_1_), .ZN(n3959) );
  NAND2_X1 U4013 ( .A1(n3963), .A2(n3964), .ZN(n3914) );
  NAND2_X1 U4014 ( .A1(d_2_), .A2(n3965), .ZN(n3964) );
  OR2_X1 U4015 ( .A1(n3797), .A2(c_2_), .ZN(n3965) );
  NAND2_X1 U4016 ( .A1(c_2_), .A2(n3797), .ZN(n3963) );
  NAND2_X1 U4017 ( .A1(n3966), .A2(n3967), .ZN(n3797) );
  NAND2_X1 U4018 ( .A1(d_3_), .A2(n3968), .ZN(n3967) );
  OR2_X1 U4019 ( .A1(n3658), .A2(c_3_), .ZN(n3968) );
  NAND2_X1 U4020 ( .A1(c_3_), .A2(n3658), .ZN(n3966) );
  NAND2_X1 U4021 ( .A1(n3969), .A2(n3970), .ZN(n3658) );
  NAND2_X1 U4022 ( .A1(d_4_), .A2(n3971), .ZN(n3970) );
  OR2_X1 U4023 ( .A1(n3527), .A2(c_4_), .ZN(n3971) );
  NAND2_X1 U4024 ( .A1(c_4_), .A2(n3527), .ZN(n3969) );
  NAND2_X1 U4025 ( .A1(n3972), .A2(n3973), .ZN(n3527) );
  NAND2_X1 U4026 ( .A1(d_5_), .A2(n3974), .ZN(n3973) );
  OR2_X1 U4027 ( .A1(n3396), .A2(c_5_), .ZN(n3974) );
  NAND2_X1 U4028 ( .A1(c_5_), .A2(n3396), .ZN(n3972) );
  NAND2_X1 U4029 ( .A1(n3975), .A2(n3976), .ZN(n3396) );
  NAND2_X1 U4030 ( .A1(d_6_), .A2(n3977), .ZN(n3976) );
  OR2_X1 U4031 ( .A1(n3274), .A2(c_6_), .ZN(n3977) );
  NAND2_X1 U4032 ( .A1(c_6_), .A2(n3274), .ZN(n3975) );
  NAND2_X1 U4033 ( .A1(n3978), .A2(n3979), .ZN(n3274) );
  NAND2_X1 U4034 ( .A1(d_7_), .A2(n3980), .ZN(n3979) );
  OR2_X1 U4035 ( .A1(n3144), .A2(c_7_), .ZN(n3980) );
  NAND2_X1 U4036 ( .A1(c_7_), .A2(n3144), .ZN(n3978) );
  NAND2_X1 U4037 ( .A1(n3981), .A2(n3982), .ZN(n3144) );
  NAND2_X1 U4038 ( .A1(d_8_), .A2(n3983), .ZN(n3982) );
  OR2_X1 U4039 ( .A1(n3019), .A2(c_8_), .ZN(n3983) );
  NAND2_X1 U4040 ( .A1(c_8_), .A2(n3019), .ZN(n3981) );
  NAND2_X1 U4041 ( .A1(n3984), .A2(n3985), .ZN(n3019) );
  NAND2_X1 U4042 ( .A1(d_9_), .A2(n3986), .ZN(n3985) );
  OR2_X1 U4043 ( .A1(n2897), .A2(c_9_), .ZN(n3986) );
  NAND2_X1 U4044 ( .A1(c_9_), .A2(n2897), .ZN(n3984) );
  NAND2_X1 U4045 ( .A1(n3987), .A2(n3988), .ZN(n2897) );
  NAND2_X1 U4046 ( .A1(d_10_), .A2(n3989), .ZN(n3988) );
  OR2_X1 U4047 ( .A1(n2774), .A2(c_10_), .ZN(n3989) );
  NAND2_X1 U4048 ( .A1(c_10_), .A2(n2774), .ZN(n3987) );
  NAND2_X1 U4049 ( .A1(n3990), .A2(n3991), .ZN(n2774) );
  NAND2_X1 U4050 ( .A1(d_11_), .A2(n3992), .ZN(n3991) );
  OR2_X1 U4051 ( .A1(n2654), .A2(c_11_), .ZN(n3992) );
  NAND2_X1 U4052 ( .A1(c_11_), .A2(n2654), .ZN(n3990) );
  NAND2_X1 U4053 ( .A1(n3993), .A2(n3994), .ZN(n2654) );
  NAND2_X1 U4054 ( .A1(d_12_), .A2(n3995), .ZN(n3994) );
  OR2_X1 U4055 ( .A1(n2526), .A2(c_12_), .ZN(n3995) );
  NAND2_X1 U4056 ( .A1(c_12_), .A2(n2526), .ZN(n3993) );
  NAND2_X1 U4057 ( .A1(n3996), .A2(n3997), .ZN(n2526) );
  NAND2_X1 U4058 ( .A1(d_13_), .A2(n3998), .ZN(n3997) );
  OR2_X1 U4059 ( .A1(n2413), .A2(c_13_), .ZN(n3998) );
  NAND2_X1 U4060 ( .A1(c_13_), .A2(n2413), .ZN(n3996) );
  NAND2_X1 U4061 ( .A1(n3999), .A2(n4000), .ZN(n2413) );
  NAND2_X1 U4062 ( .A1(d_14_), .A2(n4001), .ZN(n4000) );
  OR2_X1 U4063 ( .A1(c_14_), .A2(n2213), .ZN(n4001) );
  NAND2_X1 U4064 ( .A1(c_14_), .A2(n2213), .ZN(n3999) );
  AND2_X1 U4065 ( .A1(d_15_), .A2(c_15_), .ZN(n2213) );
endmodule

