module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n894_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n735_, new_n500_, new_n898_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n124_, new_n326_, new_n554_, new_n903_, new_n164_, new_n230_, new_n281_, new_n430_, new_n844_, new_n482_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n875_, new_n506_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n882_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n851_, new_n878_, new_n543_, new_n113_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n529_, new_n323_, new_n884_, new_n259_, new_n362_, new_n809_, new_n654_, new_n880_, new_n227_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n617_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n826_, new_n591_, new_n837_, new_n801_, new_n789_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n857_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n904_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n881_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, N85 );
and g001 ( new_n107_, new_n106_, N81 );
not g002 ( new_n108_, N81 );
and g003 ( new_n109_, new_n108_, N85 );
or g004 ( new_n110_, new_n107_, new_n109_ );
and g005 ( new_n111_, N89, N93 );
not g006 ( new_n112_, N89 );
not g007 ( new_n113_, N93 );
and g008 ( new_n114_, new_n112_, new_n113_ );
or g009 ( new_n115_, new_n114_, new_n111_ );
and g010 ( new_n116_, new_n110_, new_n115_ );
not g011 ( new_n117_, new_n116_ );
or g012 ( new_n118_, new_n110_, new_n115_ );
and g013 ( new_n119_, new_n117_, new_n118_ );
not g014 ( new_n120_, new_n119_ );
not g015 ( new_n121_, N69 );
and g016 ( new_n122_, new_n121_, N65 );
not g017 ( new_n123_, N65 );
and g018 ( new_n124_, new_n123_, N69 );
or g019 ( new_n125_, new_n122_, new_n124_ );
and g020 ( new_n126_, N73, N77 );
not g021 ( new_n127_, N73 );
not g022 ( new_n128_, N77 );
and g023 ( new_n129_, new_n127_, new_n128_ );
or g024 ( new_n130_, new_n129_, new_n126_ );
and g025 ( new_n131_, new_n125_, new_n130_ );
not g026 ( new_n132_, new_n131_ );
or g027 ( new_n133_, new_n125_, new_n130_ );
and g028 ( new_n134_, new_n132_, new_n133_ );
and g029 ( new_n135_, new_n120_, new_n134_ );
not g030 ( new_n136_, new_n134_ );
and g031 ( new_n137_, new_n136_, new_n119_ );
or g032 ( new_n138_, new_n135_, new_n137_ );
and g033 ( new_n139_, N129, N137 );
not g034 ( new_n140_, new_n139_ );
and g035 ( new_n141_, new_n138_, new_n140_ );
not g036 ( new_n142_, new_n141_ );
or g037 ( new_n143_, new_n138_, new_n140_ );
and g038 ( new_n144_, new_n142_, new_n143_ );
not g039 ( new_n145_, N17 );
and g040 ( new_n146_, new_n145_, N1 );
not g041 ( new_n147_, N1 );
and g042 ( new_n148_, new_n147_, N17 );
or g043 ( new_n149_, new_n146_, new_n148_ );
and g044 ( new_n150_, N33, N49 );
not g045 ( new_n151_, N33 );
not g046 ( new_n152_, N49 );
and g047 ( new_n153_, new_n151_, new_n152_ );
or g048 ( new_n154_, new_n153_, new_n150_ );
and g049 ( new_n155_, new_n149_, new_n154_ );
not g050 ( new_n156_, new_n155_ );
or g051 ( new_n157_, new_n149_, new_n154_ );
and g052 ( new_n158_, new_n156_, new_n157_ );
not g053 ( new_n159_, new_n158_ );
and g054 ( new_n160_, new_n159_, keyIn_0_9 );
not g055 ( new_n161_, new_n160_ );
or g056 ( new_n162_, new_n159_, keyIn_0_9 );
and g057 ( new_n163_, new_n161_, new_n162_ );
or g058 ( new_n164_, new_n144_, new_n163_ );
and g059 ( new_n165_, new_n144_, new_n163_ );
not g060 ( new_n166_, new_n165_ );
and g061 ( new_n167_, new_n166_, new_n164_ );
not g062 ( new_n168_, keyIn_0_19 );
and g063 ( new_n169_, N105, N109 );
not g064 ( new_n170_, N105 );
not g065 ( new_n171_, N109 );
and g066 ( new_n172_, new_n170_, new_n171_ );
or g067 ( new_n173_, new_n172_, new_n169_ );
and g068 ( new_n174_, new_n173_, keyIn_0_3 );
not g069 ( new_n175_, new_n174_ );
or g070 ( new_n176_, new_n173_, keyIn_0_3 );
and g071 ( new_n177_, new_n175_, new_n176_ );
not g072 ( new_n178_, N101 );
and g073 ( new_n179_, new_n178_, N97 );
not g074 ( new_n180_, N97 );
and g075 ( new_n181_, new_n180_, N101 );
or g076 ( new_n182_, new_n179_, new_n181_ );
not g077 ( new_n183_, new_n182_ );
or g078 ( new_n184_, new_n177_, new_n183_ );
and g079 ( new_n185_, new_n177_, new_n183_ );
not g080 ( new_n186_, new_n185_ );
and g081 ( new_n187_, new_n186_, new_n184_ );
not g082 ( new_n188_, new_n187_ );
and g083 ( new_n189_, N113, N117 );
not g084 ( new_n190_, N113 );
not g085 ( new_n191_, N117 );
and g086 ( new_n192_, new_n190_, new_n191_ );
or g087 ( new_n193_, new_n192_, new_n189_ );
and g088 ( new_n194_, new_n193_, keyIn_0_4 );
not g089 ( new_n195_, new_n194_ );
or g090 ( new_n196_, new_n193_, keyIn_0_4 );
and g091 ( new_n197_, new_n195_, new_n196_ );
not g092 ( new_n198_, new_n197_ );
and g093 ( new_n199_, N121, N125 );
not g094 ( new_n200_, N121 );
not g095 ( new_n201_, N125 );
and g096 ( new_n202_, new_n200_, new_n201_ );
or g097 ( new_n203_, new_n202_, new_n199_ );
and g098 ( new_n204_, new_n198_, new_n203_ );
not g099 ( new_n205_, new_n204_ );
or g100 ( new_n206_, new_n198_, new_n203_ );
and g101 ( new_n207_, new_n205_, new_n206_ );
and g102 ( new_n208_, new_n207_, new_n188_ );
not g103 ( new_n209_, new_n207_ );
and g104 ( new_n210_, new_n209_, new_n187_ );
or g105 ( new_n211_, new_n210_, new_n208_ );
and g106 ( new_n212_, N130, N137 );
not g107 ( new_n213_, new_n212_ );
and g108 ( new_n214_, new_n211_, new_n213_ );
not g109 ( new_n215_, new_n214_ );
or g110 ( new_n216_, new_n211_, new_n213_ );
and g111 ( new_n217_, new_n215_, new_n216_ );
not g112 ( new_n218_, new_n217_ );
and g113 ( new_n219_, N5, N21 );
not g114 ( new_n220_, N5 );
not g115 ( new_n221_, N21 );
and g116 ( new_n222_, new_n220_, new_n221_ );
or g117 ( new_n223_, new_n222_, new_n219_ );
and g118 ( new_n224_, N37, N53 );
not g119 ( new_n225_, N37 );
not g120 ( new_n226_, N53 );
and g121 ( new_n227_, new_n225_, new_n226_ );
or g122 ( new_n228_, new_n227_, new_n224_ );
and g123 ( new_n229_, new_n223_, new_n228_ );
not g124 ( new_n230_, new_n229_ );
or g125 ( new_n231_, new_n223_, new_n228_ );
and g126 ( new_n232_, new_n230_, new_n231_ );
not g127 ( new_n233_, new_n232_ );
and g128 ( new_n234_, new_n218_, new_n233_ );
and g129 ( new_n235_, new_n217_, new_n232_ );
or g130 ( new_n236_, new_n234_, new_n235_ );
not g131 ( new_n237_, new_n236_ );
and g132 ( new_n238_, new_n209_, new_n119_ );
and g133 ( new_n239_, new_n207_, new_n120_ );
or g134 ( new_n240_, new_n238_, new_n239_ );
and g135 ( new_n241_, N132, N137 );
not g136 ( new_n242_, new_n241_ );
and g137 ( new_n243_, new_n240_, new_n242_ );
not g138 ( new_n244_, new_n243_ );
or g139 ( new_n245_, new_n240_, new_n242_ );
and g140 ( new_n246_, new_n244_, new_n245_ );
not g141 ( new_n247_, new_n246_ );
and g142 ( new_n248_, N13, N29 );
not g143 ( new_n249_, N13 );
not g144 ( new_n250_, N29 );
and g145 ( new_n251_, new_n249_, new_n250_ );
or g146 ( new_n252_, new_n251_, new_n248_ );
and g147 ( new_n253_, N45, N61 );
not g148 ( new_n254_, N45 );
not g149 ( new_n255_, N61 );
and g150 ( new_n256_, new_n254_, new_n255_ );
or g151 ( new_n257_, new_n256_, new_n253_ );
and g152 ( new_n258_, new_n252_, new_n257_ );
not g153 ( new_n259_, new_n258_ );
or g154 ( new_n260_, new_n252_, new_n257_ );
and g155 ( new_n261_, new_n259_, new_n260_ );
not g156 ( new_n262_, new_n261_ );
and g157 ( new_n263_, new_n247_, new_n262_ );
and g158 ( new_n264_, new_n246_, new_n261_ );
or g159 ( new_n265_, new_n263_, new_n264_ );
and g160 ( new_n266_, new_n237_, new_n265_ );
and g161 ( new_n267_, new_n188_, new_n134_ );
and g162 ( new_n268_, new_n187_, new_n136_ );
or g163 ( new_n269_, new_n267_, new_n268_ );
and g164 ( new_n270_, N131, N137 );
not g165 ( new_n271_, new_n270_ );
and g166 ( new_n272_, new_n269_, new_n271_ );
not g167 ( new_n273_, new_n272_ );
or g168 ( new_n274_, new_n269_, new_n271_ );
and g169 ( new_n275_, new_n273_, new_n274_ );
not g170 ( new_n276_, new_n275_ );
and g171 ( new_n277_, N41, N57 );
not g172 ( new_n278_, N41 );
not g173 ( new_n279_, N57 );
and g174 ( new_n280_, new_n278_, new_n279_ );
or g175 ( new_n281_, new_n280_, new_n277_ );
and g176 ( new_n282_, new_n281_, keyIn_0_6 );
not g177 ( new_n283_, new_n282_ );
or g178 ( new_n284_, new_n281_, keyIn_0_6 );
and g179 ( new_n285_, new_n283_, new_n284_ );
not g180 ( new_n286_, new_n285_ );
and g181 ( new_n287_, N9, N25 );
not g182 ( new_n288_, N9 );
not g183 ( new_n289_, N25 );
and g184 ( new_n290_, new_n288_, new_n289_ );
or g185 ( new_n291_, new_n290_, new_n287_ );
and g186 ( new_n292_, new_n286_, new_n291_ );
not g187 ( new_n293_, new_n292_ );
or g188 ( new_n294_, new_n286_, new_n291_ );
and g189 ( new_n295_, new_n293_, new_n294_ );
not g190 ( new_n296_, new_n295_ );
and g191 ( new_n297_, new_n276_, new_n296_ );
and g192 ( new_n298_, new_n275_, new_n295_ );
or g193 ( new_n299_, new_n297_, new_n298_ );
not g194 ( new_n300_, new_n167_ );
and g195 ( new_n301_, new_n300_, keyIn_0_11 );
not g196 ( new_n302_, new_n301_ );
or g197 ( new_n303_, new_n300_, keyIn_0_11 );
and g198 ( new_n304_, new_n302_, new_n303_ );
or g199 ( new_n305_, new_n304_, new_n299_ );
not g200 ( new_n306_, new_n305_ );
and g201 ( new_n307_, new_n306_, new_n266_ );
and g202 ( new_n308_, new_n307_, new_n168_ );
not g203 ( new_n309_, new_n308_ );
or g204 ( new_n310_, new_n307_, new_n168_ );
and g205 ( new_n311_, new_n309_, new_n310_ );
and g206 ( new_n312_, new_n299_, keyIn_0_12 );
and g207 ( new_n313_, new_n312_, new_n236_ );
not g208 ( new_n314_, new_n313_ );
or g209 ( new_n315_, new_n312_, new_n236_ );
not g210 ( new_n316_, new_n265_ );
and g211 ( new_n317_, new_n316_, new_n300_ );
and g212 ( new_n318_, new_n315_, new_n317_ );
and g213 ( new_n319_, new_n318_, new_n314_ );
and g214 ( new_n320_, new_n236_, keyIn_0_13 );
not g215 ( new_n321_, keyIn_0_13 );
and g216 ( new_n322_, new_n237_, new_n321_ );
or g217 ( new_n323_, new_n322_, new_n320_ );
not g218 ( new_n324_, new_n299_ );
and g219 ( new_n325_, new_n316_, new_n167_ );
and g220 ( new_n326_, new_n325_, new_n324_ );
and g221 ( new_n327_, new_n323_, new_n326_ );
or g222 ( new_n328_, new_n319_, new_n327_ );
or g223 ( new_n329_, new_n311_, new_n328_ );
and g224 ( new_n330_, N77, N93 );
and g225 ( new_n331_, new_n128_, new_n113_ );
or g226 ( new_n332_, new_n331_, new_n330_ );
and g227 ( new_n333_, N109, N125 );
and g228 ( new_n334_, new_n171_, new_n201_ );
or g229 ( new_n335_, new_n334_, new_n333_ );
and g230 ( new_n336_, new_n332_, new_n335_ );
not g231 ( new_n337_, new_n336_ );
or g232 ( new_n338_, new_n332_, new_n335_ );
and g233 ( new_n339_, new_n337_, new_n338_ );
not g234 ( new_n340_, keyIn_0_10 );
and g235 ( new_n341_, N49, N53 );
and g236 ( new_n342_, new_n152_, new_n226_ );
or g237 ( new_n343_, new_n342_, new_n341_ );
and g238 ( new_n344_, N57, N61 );
and g239 ( new_n345_, new_n279_, new_n255_ );
or g240 ( new_n346_, new_n345_, new_n344_ );
and g241 ( new_n347_, new_n343_, new_n346_ );
not g242 ( new_n348_, new_n347_ );
or g243 ( new_n349_, new_n343_, new_n346_ );
and g244 ( new_n350_, new_n348_, new_n349_ );
not g245 ( new_n351_, keyIn_0_0 );
and g246 ( new_n352_, N17, N21 );
and g247 ( new_n353_, new_n145_, new_n221_ );
or g248 ( new_n354_, new_n353_, new_n352_ );
or g249 ( new_n355_, new_n354_, new_n351_ );
not g250 ( new_n356_, new_n352_ );
or g251 ( new_n357_, N17, N21 );
and g252 ( new_n358_, new_n356_, new_n357_ );
or g253 ( new_n359_, new_n358_, keyIn_0_0 );
and g254 ( new_n360_, new_n355_, new_n359_ );
and g255 ( new_n361_, N25, N29 );
and g256 ( new_n362_, new_n289_, new_n250_ );
or g257 ( new_n363_, new_n362_, new_n361_ );
not g258 ( new_n364_, new_n363_ );
or g259 ( new_n365_, new_n360_, new_n364_ );
and g260 ( new_n366_, new_n358_, keyIn_0_0 );
and g261 ( new_n367_, new_n354_, new_n351_ );
or g262 ( new_n368_, new_n367_, new_n366_ );
or g263 ( new_n369_, new_n368_, new_n363_ );
and g264 ( new_n370_, new_n369_, new_n365_ );
or g265 ( new_n371_, new_n370_, new_n350_ );
not g266 ( new_n372_, new_n350_ );
and g267 ( new_n373_, new_n368_, new_n363_ );
and g268 ( new_n374_, new_n360_, new_n364_ );
or g269 ( new_n375_, new_n373_, new_n374_ );
or g270 ( new_n376_, new_n375_, new_n372_ );
and g271 ( new_n377_, new_n376_, new_n371_ );
and g272 ( new_n378_, N136, N137 );
or g273 ( new_n379_, new_n377_, new_n378_ );
and g274 ( new_n380_, new_n375_, new_n372_ );
and g275 ( new_n381_, new_n370_, new_n350_ );
or g276 ( new_n382_, new_n380_, new_n381_ );
not g277 ( new_n383_, new_n378_ );
or g278 ( new_n384_, new_n382_, new_n383_ );
and g279 ( new_n385_, new_n384_, new_n379_ );
or g280 ( new_n386_, new_n385_, new_n340_ );
and g281 ( new_n387_, new_n382_, new_n383_ );
and g282 ( new_n388_, new_n377_, new_n378_ );
or g283 ( new_n389_, new_n387_, new_n388_ );
or g284 ( new_n390_, new_n389_, keyIn_0_10 );
and g285 ( new_n391_, new_n390_, new_n386_ );
or g286 ( new_n392_, new_n391_, new_n339_ );
not g287 ( new_n393_, new_n339_ );
and g288 ( new_n394_, new_n389_, keyIn_0_10 );
and g289 ( new_n395_, new_n385_, new_n340_ );
or g290 ( new_n396_, new_n394_, new_n395_ );
or g291 ( new_n397_, new_n396_, new_n393_ );
and g292 ( new_n398_, new_n397_, new_n392_ );
and g293 ( new_n399_, new_n398_, keyIn_0_15 );
not g294 ( new_n400_, new_n399_ );
and g295 ( new_n401_, N1, N5 );
and g296 ( new_n402_, new_n147_, new_n220_ );
or g297 ( new_n403_, new_n402_, new_n401_ );
and g298 ( new_n404_, N9, N13 );
and g299 ( new_n405_, new_n288_, new_n249_ );
or g300 ( new_n406_, new_n405_, new_n404_ );
not g301 ( new_n407_, new_n406_ );
and g302 ( new_n408_, new_n407_, new_n403_ );
not g303 ( new_n409_, new_n408_ );
or g304 ( new_n410_, new_n407_, new_n403_ );
and g305 ( new_n411_, new_n409_, new_n410_ );
and g306 ( new_n412_, new_n375_, new_n411_ );
not g307 ( new_n413_, new_n411_ );
and g308 ( new_n414_, new_n370_, new_n413_ );
or g309 ( new_n415_, new_n412_, new_n414_ );
and g310 ( new_n416_, N133, N137 );
not g311 ( new_n417_, new_n416_ );
and g312 ( new_n418_, new_n415_, new_n417_ );
not g313 ( new_n419_, new_n418_ );
or g314 ( new_n420_, new_n415_, new_n417_ );
and g315 ( new_n421_, new_n419_, new_n420_ );
not g316 ( new_n422_, new_n421_ );
and g317 ( new_n423_, N65, N81 );
and g318 ( new_n424_, new_n123_, new_n108_ );
or g319 ( new_n425_, new_n424_, new_n423_ );
and g320 ( new_n426_, N97, N113 );
and g321 ( new_n427_, new_n180_, new_n190_ );
or g322 ( new_n428_, new_n427_, new_n426_ );
and g323 ( new_n429_, new_n425_, new_n428_ );
not g324 ( new_n430_, new_n429_ );
or g325 ( new_n431_, new_n425_, new_n428_ );
and g326 ( new_n432_, new_n430_, new_n431_ );
not g327 ( new_n433_, new_n432_ );
and g328 ( new_n434_, new_n422_, new_n433_ );
and g329 ( new_n435_, new_n421_, new_n432_ );
or g330 ( new_n436_, new_n434_, new_n435_ );
not g331 ( new_n437_, keyIn_0_5 );
and g332 ( new_n438_, N135, N137 );
or g333 ( new_n439_, new_n438_, new_n437_ );
and g334 ( new_n440_, new_n438_, new_n437_ );
not g335 ( new_n441_, new_n440_ );
and g336 ( new_n442_, new_n441_, new_n439_ );
not g337 ( new_n443_, new_n442_ );
and g338 ( new_n444_, new_n225_, N33 );
and g339 ( new_n445_, new_n151_, N37 );
or g340 ( new_n446_, new_n444_, new_n445_ );
or g341 ( new_n447_, new_n446_, keyIn_0_1 );
not g342 ( new_n448_, keyIn_0_1 );
or g343 ( new_n449_, new_n151_, N37 );
or g344 ( new_n450_, new_n225_, N33 );
and g345 ( new_n451_, new_n449_, new_n450_ );
or g346 ( new_n452_, new_n451_, new_n448_ );
and g347 ( new_n453_, new_n447_, new_n452_ );
and g348 ( new_n454_, N41, N45 );
not g349 ( new_n455_, new_n454_ );
or g350 ( new_n456_, N41, N45 );
and g351 ( new_n457_, new_n455_, new_n456_ );
or g352 ( new_n458_, new_n457_, keyIn_0_2 );
not g353 ( new_n459_, keyIn_0_2 );
and g354 ( new_n460_, new_n278_, new_n254_ );
or g355 ( new_n461_, new_n460_, new_n454_ );
or g356 ( new_n462_, new_n461_, new_n459_ );
and g357 ( new_n463_, new_n462_, new_n458_ );
or g358 ( new_n464_, new_n453_, new_n463_ );
and g359 ( new_n465_, new_n451_, new_n448_ );
and g360 ( new_n466_, new_n446_, keyIn_0_1 );
or g361 ( new_n467_, new_n466_, new_n465_ );
and g362 ( new_n468_, new_n461_, new_n459_ );
and g363 ( new_n469_, new_n457_, keyIn_0_2 );
or g364 ( new_n470_, new_n468_, new_n469_ );
or g365 ( new_n471_, new_n467_, new_n470_ );
and g366 ( new_n472_, new_n471_, new_n464_ );
or g367 ( new_n473_, new_n472_, keyIn_0_8 );
not g368 ( new_n474_, keyIn_0_8 );
and g369 ( new_n475_, new_n467_, new_n470_ );
and g370 ( new_n476_, new_n453_, new_n463_ );
or g371 ( new_n477_, new_n475_, new_n476_ );
or g372 ( new_n478_, new_n477_, new_n474_ );
and g373 ( new_n479_, new_n478_, new_n473_ );
or g374 ( new_n480_, new_n479_, new_n413_ );
and g375 ( new_n481_, new_n477_, new_n474_ );
and g376 ( new_n482_, new_n464_, keyIn_0_8 );
and g377 ( new_n483_, new_n482_, new_n471_ );
or g378 ( new_n484_, new_n481_, new_n483_ );
or g379 ( new_n485_, new_n484_, new_n411_ );
and g380 ( new_n486_, new_n485_, new_n480_ );
or g381 ( new_n487_, new_n486_, new_n443_ );
and g382 ( new_n488_, new_n484_, new_n411_ );
or g383 ( new_n489_, new_n475_, new_n474_ );
or g384 ( new_n490_, new_n489_, new_n476_ );
and g385 ( new_n491_, new_n473_, new_n490_ );
and g386 ( new_n492_, new_n491_, new_n413_ );
or g387 ( new_n493_, new_n492_, new_n442_ );
or g388 ( new_n494_, new_n493_, new_n488_ );
and g389 ( new_n495_, new_n487_, new_n494_ );
and g390 ( new_n496_, N105, N121 );
and g391 ( new_n497_, new_n170_, new_n200_ );
or g392 ( new_n498_, new_n497_, new_n496_ );
and g393 ( new_n499_, new_n498_, keyIn_0_7 );
not g394 ( new_n500_, new_n499_ );
or g395 ( new_n501_, new_n498_, keyIn_0_7 );
and g396 ( new_n502_, new_n500_, new_n501_ );
not g397 ( new_n503_, new_n502_ );
and g398 ( new_n504_, N73, N89 );
and g399 ( new_n505_, new_n127_, new_n112_ );
or g400 ( new_n506_, new_n505_, new_n504_ );
and g401 ( new_n507_, new_n503_, new_n506_ );
not g402 ( new_n508_, new_n507_ );
or g403 ( new_n509_, new_n503_, new_n506_ );
and g404 ( new_n510_, new_n508_, new_n509_ );
not g405 ( new_n511_, new_n510_ );
or g406 ( new_n512_, new_n495_, new_n511_ );
and g407 ( new_n513_, new_n472_, keyIn_0_8 );
or g408 ( new_n514_, new_n481_, new_n513_ );
and g409 ( new_n515_, new_n514_, new_n411_ );
or g410 ( new_n516_, new_n515_, new_n492_ );
and g411 ( new_n517_, new_n516_, new_n442_ );
not g412 ( new_n518_, new_n488_ );
and g413 ( new_n519_, new_n485_, new_n443_ );
and g414 ( new_n520_, new_n519_, new_n518_ );
or g415 ( new_n521_, new_n517_, new_n520_ );
or g416 ( new_n522_, new_n521_, new_n510_ );
and g417 ( new_n523_, new_n522_, new_n512_ );
and g418 ( new_n524_, new_n523_, new_n436_ );
and g419 ( new_n525_, new_n400_, new_n524_ );
and g420 ( new_n526_, N69, N85 );
and g421 ( new_n527_, new_n121_, new_n106_ );
or g422 ( new_n528_, new_n527_, new_n526_ );
and g423 ( new_n529_, N101, N117 );
and g424 ( new_n530_, new_n178_, new_n191_ );
or g425 ( new_n531_, new_n530_, new_n529_ );
and g426 ( new_n532_, new_n528_, new_n531_ );
not g427 ( new_n533_, new_n532_ );
or g428 ( new_n534_, new_n528_, new_n531_ );
and g429 ( new_n535_, new_n533_, new_n534_ );
and g430 ( new_n536_, N134, N137 );
and g431 ( new_n537_, new_n491_, new_n372_ );
and g432 ( new_n538_, new_n484_, new_n350_ );
or g433 ( new_n539_, new_n538_, new_n537_ );
and g434 ( new_n540_, new_n539_, new_n536_ );
not g435 ( new_n541_, new_n536_ );
or g436 ( new_n542_, new_n491_, new_n372_ );
or g437 ( new_n543_, new_n514_, new_n350_ );
and g438 ( new_n544_, new_n543_, new_n542_ );
and g439 ( new_n545_, new_n544_, new_n541_ );
or g440 ( new_n546_, new_n540_, new_n545_ );
or g441 ( new_n547_, new_n546_, new_n535_ );
not g442 ( new_n548_, new_n535_ );
or g443 ( new_n549_, new_n484_, new_n350_ );
and g444 ( new_n550_, new_n549_, new_n542_ );
or g445 ( new_n551_, new_n550_, new_n541_ );
and g446 ( new_n552_, new_n479_, new_n372_ );
or g447 ( new_n553_, new_n538_, new_n552_ );
or g448 ( new_n554_, new_n553_, new_n536_ );
and g449 ( new_n555_, new_n554_, new_n551_ );
or g450 ( new_n556_, new_n555_, new_n548_ );
and g451 ( new_n557_, new_n547_, new_n556_ );
and g452 ( new_n558_, new_n557_, keyIn_0_14 );
not g453 ( new_n559_, new_n558_ );
or g454 ( new_n560_, new_n544_, new_n541_ );
and g455 ( new_n561_, new_n554_, new_n560_ );
or g456 ( new_n562_, new_n561_, new_n548_ );
and g457 ( new_n563_, new_n547_, new_n562_ );
or g458 ( new_n564_, new_n563_, keyIn_0_14 );
or g459 ( new_n565_, new_n398_, keyIn_0_15 );
and g460 ( new_n566_, new_n564_, new_n565_ );
and g461 ( new_n567_, new_n566_, new_n559_ );
and g462 ( new_n568_, new_n567_, new_n525_ );
and g463 ( new_n569_, new_n329_, new_n568_ );
or g464 ( new_n570_, new_n569_, keyIn_0_24 );
and g465 ( new_n571_, new_n569_, keyIn_0_24 );
not g466 ( new_n572_, new_n571_ );
and g467 ( new_n573_, new_n572_, new_n570_ );
and g468 ( new_n574_, new_n573_, new_n167_ );
not g469 ( new_n575_, new_n574_ );
and g470 ( new_n576_, new_n575_, N1 );
and g471 ( new_n577_, new_n574_, new_n147_ );
or g472 ( N724, new_n576_, new_n577_ );
and g473 ( new_n579_, new_n573_, new_n236_ );
not g474 ( new_n580_, new_n579_ );
and g475 ( new_n581_, new_n580_, N5 );
and g476 ( new_n582_, new_n579_, new_n220_ );
or g477 ( N725, new_n581_, new_n582_ );
not g478 ( new_n584_, keyIn_0_24 );
not g479 ( new_n585_, new_n310_ );
or g480 ( new_n586_, new_n585_, new_n308_ );
not g481 ( new_n587_, new_n328_ );
and g482 ( new_n588_, new_n586_, new_n587_ );
not g483 ( new_n589_, new_n568_ );
or g484 ( new_n590_, new_n588_, new_n589_ );
and g485 ( new_n591_, new_n590_, new_n584_ );
or g486 ( new_n592_, new_n591_, new_n571_ );
or g487 ( new_n593_, new_n592_, new_n324_ );
and g488 ( new_n594_, new_n593_, N9 );
and g489 ( new_n595_, new_n573_, new_n299_ );
and g490 ( new_n596_, new_n595_, new_n288_ );
or g491 ( new_n597_, new_n596_, new_n594_ );
and g492 ( new_n598_, new_n597_, keyIn_0_30 );
not g493 ( new_n599_, keyIn_0_30 );
or g494 ( new_n600_, new_n595_, new_n288_ );
or g495 ( new_n601_, new_n593_, N9 );
and g496 ( new_n602_, new_n600_, new_n601_ );
and g497 ( new_n603_, new_n602_, new_n599_ );
or g498 ( N726, new_n598_, new_n603_ );
or g499 ( new_n605_, new_n592_, new_n316_ );
and g500 ( new_n606_, new_n605_, N13 );
and g501 ( new_n607_, new_n573_, new_n265_ );
and g502 ( new_n608_, new_n607_, new_n249_ );
or g503 ( new_n609_, new_n608_, new_n606_ );
and g504 ( new_n610_, new_n609_, keyIn_0_31 );
not g505 ( new_n611_, keyIn_0_31 );
or g506 ( new_n612_, new_n607_, new_n249_ );
or g507 ( new_n613_, new_n605_, N13 );
and g508 ( new_n614_, new_n612_, new_n613_ );
and g509 ( new_n615_, new_n614_, new_n611_ );
or g510 ( N727, new_n610_, new_n615_ );
and g511 ( new_n617_, new_n555_, new_n548_ );
and g512 ( new_n618_, new_n553_, new_n536_ );
or g513 ( new_n619_, new_n618_, new_n545_ );
and g514 ( new_n620_, new_n619_, new_n535_ );
or g515 ( new_n621_, new_n620_, new_n617_ );
and g516 ( new_n622_, new_n621_, new_n436_ );
and g517 ( new_n623_, new_n521_, new_n510_ );
and g518 ( new_n624_, new_n495_, new_n511_ );
or g519 ( new_n625_, new_n623_, new_n624_ );
and g520 ( new_n626_, new_n625_, new_n398_ );
and g521 ( new_n627_, new_n622_, new_n626_ );
and g522 ( new_n628_, new_n329_, new_n627_ );
and g523 ( new_n629_, new_n628_, new_n167_ );
not g524 ( new_n630_, new_n629_ );
and g525 ( new_n631_, new_n630_, N17 );
and g526 ( new_n632_, new_n629_, new_n145_ );
or g527 ( N728, new_n631_, new_n632_ );
and g528 ( new_n634_, new_n628_, new_n236_ );
not g529 ( new_n635_, new_n634_ );
and g530 ( new_n636_, new_n635_, N21 );
and g531 ( new_n637_, new_n634_, new_n221_ );
or g532 ( N729, new_n636_, new_n637_ );
not g533 ( new_n639_, keyIn_0_25 );
and g534 ( new_n640_, new_n628_, new_n299_ );
not g535 ( new_n641_, new_n640_ );
and g536 ( new_n642_, new_n641_, new_n639_ );
and g537 ( new_n643_, new_n640_, keyIn_0_25 );
or g538 ( new_n644_, new_n642_, new_n643_ );
and g539 ( new_n645_, new_n644_, N25 );
not g540 ( new_n646_, new_n644_ );
and g541 ( new_n647_, new_n646_, new_n289_ );
or g542 ( N730, new_n647_, new_n645_ );
and g543 ( new_n649_, new_n628_, new_n265_ );
not g544 ( new_n650_, new_n649_ );
and g545 ( new_n651_, new_n650_, keyIn_0_26 );
not g546 ( new_n652_, new_n651_ );
or g547 ( new_n653_, new_n650_, keyIn_0_26 );
and g548 ( new_n654_, new_n652_, new_n653_ );
not g549 ( new_n655_, new_n654_ );
and g550 ( new_n656_, new_n655_, N29 );
and g551 ( new_n657_, new_n654_, new_n250_ );
or g552 ( N731, new_n656_, new_n657_ );
and g553 ( new_n659_, new_n329_, new_n557_ );
not g554 ( new_n660_, keyIn_0_16 );
and g555 ( new_n661_, new_n436_, new_n660_ );
not g556 ( new_n662_, new_n436_ );
and g557 ( new_n663_, new_n662_, keyIn_0_16 );
or g558 ( new_n664_, new_n663_, new_n661_ );
and g559 ( new_n665_, new_n396_, new_n393_ );
and g560 ( new_n666_, new_n391_, new_n339_ );
or g561 ( new_n667_, new_n665_, new_n666_ );
and g562 ( new_n668_, new_n667_, new_n523_ );
and g563 ( new_n669_, new_n664_, new_n668_ );
and g564 ( new_n670_, new_n659_, new_n669_ );
and g565 ( new_n671_, new_n670_, new_n167_ );
and g566 ( new_n672_, new_n671_, new_n151_ );
not g567 ( new_n673_, new_n671_ );
and g568 ( new_n674_, new_n673_, N33 );
or g569 ( N732, new_n674_, new_n672_ );
and g570 ( new_n676_, new_n670_, new_n236_ );
and g571 ( new_n677_, new_n676_, new_n225_ );
not g572 ( new_n678_, new_n676_ );
and g573 ( new_n679_, new_n678_, N37 );
or g574 ( N733, new_n679_, new_n677_ );
and g575 ( new_n681_, new_n670_, new_n299_ );
and g576 ( new_n682_, new_n681_, new_n278_ );
not g577 ( new_n683_, new_n681_ );
and g578 ( new_n684_, new_n683_, N41 );
or g579 ( N734, new_n684_, new_n682_ );
and g580 ( new_n686_, new_n670_, new_n265_ );
and g581 ( new_n687_, new_n686_, new_n254_ );
not g582 ( new_n688_, new_n686_ );
and g583 ( new_n689_, new_n688_, N45 );
or g584 ( N735, new_n689_, new_n687_ );
or g585 ( new_n691_, new_n667_, new_n523_ );
not g586 ( new_n692_, keyIn_0_17 );
and g587 ( new_n693_, new_n436_, new_n692_ );
and g588 ( new_n694_, new_n662_, keyIn_0_17 );
or g589 ( new_n695_, new_n694_, new_n693_ );
or g590 ( new_n696_, new_n691_, new_n695_ );
not g591 ( new_n697_, new_n696_ );
and g592 ( new_n698_, new_n659_, new_n697_ );
and g593 ( new_n699_, new_n698_, new_n167_ );
not g594 ( new_n700_, new_n699_ );
and g595 ( new_n701_, new_n700_, N49 );
and g596 ( new_n702_, new_n699_, new_n152_ );
or g597 ( N736, new_n701_, new_n702_ );
and g598 ( new_n704_, new_n698_, new_n236_ );
not g599 ( new_n705_, new_n704_ );
and g600 ( new_n706_, new_n705_, N53 );
and g601 ( new_n707_, new_n704_, new_n226_ );
or g602 ( N737, new_n706_, new_n707_ );
and g603 ( new_n709_, new_n698_, new_n299_ );
not g604 ( new_n710_, new_n709_ );
and g605 ( new_n711_, new_n710_, N57 );
and g606 ( new_n712_, new_n709_, new_n279_ );
or g607 ( N738, new_n711_, new_n712_ );
and g608 ( new_n714_, new_n698_, new_n265_ );
not g609 ( new_n715_, new_n714_ );
and g610 ( new_n716_, new_n715_, N61 );
and g611 ( new_n717_, new_n714_, new_n255_ );
or g612 ( N739, new_n716_, new_n717_ );
and g613 ( new_n719_, new_n546_, new_n535_ );
or g614 ( new_n720_, new_n719_, new_n617_ );
and g615 ( new_n721_, new_n720_, new_n662_ );
and g616 ( new_n722_, new_n721_, new_n626_ );
or g617 ( new_n723_, new_n722_, keyIn_0_20 );
or g618 ( new_n724_, new_n563_, new_n662_ );
or g619 ( new_n725_, new_n724_, new_n398_ );
and g620 ( new_n726_, new_n523_, keyIn_0_18 );
not g621 ( new_n727_, keyIn_0_18 );
and g622 ( new_n728_, new_n625_, new_n727_ );
or g623 ( new_n729_, new_n728_, new_n726_ );
or g624 ( new_n730_, new_n725_, new_n729_ );
and g625 ( new_n731_, new_n621_, new_n662_ );
and g626 ( new_n732_, new_n731_, new_n626_ );
and g627 ( new_n733_, new_n732_, keyIn_0_20 );
not g628 ( new_n734_, new_n733_ );
and g629 ( new_n735_, new_n734_, new_n730_ );
and g630 ( new_n736_, new_n735_, new_n723_ );
or g631 ( new_n737_, new_n398_, new_n436_ );
or g632 ( new_n738_, new_n621_, new_n523_ );
or g633 ( new_n739_, new_n738_, new_n737_ );
and g634 ( new_n740_, new_n739_, keyIn_0_22 );
not g635 ( new_n741_, keyIn_0_22 );
and g636 ( new_n742_, new_n667_, new_n662_ );
and g637 ( new_n743_, new_n563_, new_n625_ );
and g638 ( new_n744_, new_n743_, new_n742_ );
and g639 ( new_n745_, new_n744_, new_n741_ );
or g640 ( new_n746_, new_n740_, new_n745_ );
and g641 ( new_n747_, new_n731_, new_n668_ );
and g642 ( new_n748_, new_n747_, keyIn_0_21 );
not g643 ( new_n749_, new_n748_ );
and g644 ( new_n750_, new_n721_, new_n668_ );
or g645 ( new_n751_, new_n750_, keyIn_0_21 );
and g646 ( new_n752_, new_n749_, new_n751_ );
and g647 ( new_n753_, new_n752_, new_n746_ );
and g648 ( new_n754_, new_n736_, new_n753_ );
and g649 ( new_n755_, new_n754_, keyIn_0_23 );
not g650 ( new_n756_, keyIn_0_23 );
not g651 ( new_n757_, new_n723_ );
and g652 ( new_n758_, new_n622_, new_n667_ );
or g653 ( new_n759_, new_n625_, new_n727_ );
or g654 ( new_n760_, new_n523_, keyIn_0_18 );
and g655 ( new_n761_, new_n759_, new_n760_ );
and g656 ( new_n762_, new_n761_, new_n758_ );
or g657 ( new_n763_, new_n762_, new_n733_ );
or g658 ( new_n764_, new_n763_, new_n757_ );
or g659 ( new_n765_, new_n744_, new_n741_ );
or g660 ( new_n766_, new_n739_, keyIn_0_22 );
and g661 ( new_n767_, new_n766_, new_n765_ );
not g662 ( new_n768_, keyIn_0_21 );
or g663 ( new_n769_, new_n625_, new_n398_ );
or g664 ( new_n770_, new_n557_, new_n436_ );
or g665 ( new_n771_, new_n769_, new_n770_ );
and g666 ( new_n772_, new_n771_, new_n768_ );
or g667 ( new_n773_, new_n772_, new_n748_ );
or g668 ( new_n774_, new_n773_, new_n767_ );
or g669 ( new_n775_, new_n774_, new_n764_ );
and g670 ( new_n776_, new_n775_, new_n756_ );
or g671 ( new_n777_, new_n776_, new_n755_ );
or g672 ( new_n778_, new_n777_, new_n662_ );
and g673 ( new_n779_, new_n237_, new_n299_ );
and g674 ( new_n780_, new_n779_, new_n325_ );
not g675 ( new_n781_, new_n780_ );
or g676 ( new_n782_, new_n778_, new_n781_ );
and g677 ( new_n783_, new_n782_, N65 );
not g678 ( new_n784_, new_n782_ );
and g679 ( new_n785_, new_n784_, new_n123_ );
or g680 ( N740, new_n785_, new_n783_ );
or g681 ( new_n787_, new_n777_, new_n720_ );
or g682 ( new_n788_, new_n787_, new_n781_ );
and g683 ( new_n789_, new_n788_, N69 );
not g684 ( new_n790_, new_n788_ );
and g685 ( new_n791_, new_n790_, new_n121_ );
or g686 ( N741, new_n791_, new_n789_ );
or g687 ( new_n793_, new_n777_, new_n625_ );
or g688 ( new_n794_, new_n793_, new_n781_ );
and g689 ( new_n795_, new_n794_, N73 );
not g690 ( new_n796_, new_n794_ );
and g691 ( new_n797_, new_n796_, new_n127_ );
or g692 ( N742, new_n797_, new_n795_ );
or g693 ( new_n799_, new_n777_, new_n667_ );
or g694 ( new_n800_, new_n799_, new_n781_ );
and g695 ( new_n801_, new_n800_, N77 );
not g696 ( new_n802_, new_n800_ );
and g697 ( new_n803_, new_n802_, new_n128_ );
or g698 ( N743, new_n803_, new_n801_ );
and g699 ( new_n805_, new_n324_, new_n167_ );
and g700 ( new_n806_, new_n266_, new_n805_ );
not g701 ( new_n807_, new_n806_ );
or g702 ( new_n808_, new_n778_, new_n807_ );
and g703 ( new_n809_, new_n808_, N81 );
not g704 ( new_n810_, new_n808_ );
and g705 ( new_n811_, new_n810_, new_n108_ );
or g706 ( N744, new_n811_, new_n809_ );
or g707 ( new_n813_, new_n787_, new_n807_ );
and g708 ( new_n814_, keyIn_0_27, N85 );
not g709 ( new_n815_, new_n814_ );
or g710 ( new_n816_, keyIn_0_27, N85 );
and g711 ( new_n817_, new_n815_, new_n816_ );
not g712 ( new_n818_, new_n817_ );
and g713 ( new_n819_, new_n813_, new_n818_ );
not g714 ( new_n820_, new_n813_ );
and g715 ( new_n821_, new_n820_, new_n817_ );
or g716 ( N745, new_n821_, new_n819_ );
or g717 ( new_n823_, new_n793_, new_n807_ );
and g718 ( new_n824_, new_n823_, N89 );
not g719 ( new_n825_, new_n823_ );
and g720 ( new_n826_, new_n825_, new_n112_ );
or g721 ( N746, new_n826_, new_n824_ );
or g722 ( new_n828_, new_n799_, new_n807_ );
and g723 ( new_n829_, new_n828_, N93 );
not g724 ( new_n830_, new_n828_ );
and g725 ( new_n831_, new_n830_, new_n113_ );
or g726 ( N747, new_n831_, new_n829_ );
and g727 ( new_n833_, new_n236_, new_n299_ );
and g728 ( new_n834_, new_n317_, new_n833_ );
not g729 ( new_n835_, new_n834_ );
or g730 ( new_n836_, new_n778_, new_n835_ );
and g731 ( new_n837_, new_n836_, N97 );
not g732 ( new_n838_, new_n836_ );
and g733 ( new_n839_, new_n838_, new_n180_ );
or g734 ( N748, new_n839_, new_n837_ );
or g735 ( new_n841_, new_n787_, new_n835_ );
and g736 ( new_n842_, new_n841_, N101 );
not g737 ( new_n843_, new_n841_ );
and g738 ( new_n844_, new_n843_, new_n178_ );
or g739 ( N749, new_n844_, new_n842_ );
or g740 ( new_n846_, new_n793_, new_n835_ );
and g741 ( new_n847_, new_n846_, N105 );
not g742 ( new_n848_, new_n846_ );
and g743 ( new_n849_, new_n848_, new_n170_ );
or g744 ( N750, new_n849_, new_n847_ );
or g745 ( new_n851_, new_n799_, new_n835_ );
and g746 ( new_n852_, new_n171_, keyIn_0_28 );
not g747 ( new_n853_, new_n852_ );
or g748 ( new_n854_, new_n171_, keyIn_0_28 );
and g749 ( new_n855_, new_n853_, new_n854_ );
not g750 ( new_n856_, new_n855_ );
and g751 ( new_n857_, new_n851_, new_n856_ );
not g752 ( new_n858_, new_n851_ );
and g753 ( new_n859_, new_n858_, new_n855_ );
or g754 ( N751, new_n859_, new_n857_ );
and g755 ( new_n861_, new_n236_, new_n300_ );
and g756 ( new_n862_, new_n265_, new_n324_ );
and g757 ( new_n863_, new_n862_, new_n861_ );
not g758 ( new_n864_, new_n863_ );
or g759 ( new_n865_, new_n778_, new_n864_ );
and g760 ( new_n866_, new_n865_, N113 );
not g761 ( new_n867_, new_n865_ );
and g762 ( new_n868_, new_n867_, new_n190_ );
or g763 ( N752, new_n868_, new_n866_ );
or g764 ( new_n870_, new_n787_, new_n864_ );
and g765 ( new_n871_, new_n870_, keyIn_0_29 );
not g766 ( new_n872_, keyIn_0_29 );
not g767 ( new_n873_, new_n776_ );
not g768 ( new_n874_, keyIn_0_20 );
or g769 ( new_n875_, new_n563_, new_n436_ );
or g770 ( new_n876_, new_n691_, new_n875_ );
and g771 ( new_n877_, new_n876_, new_n874_ );
or g772 ( new_n878_, new_n769_, new_n875_ );
and g773 ( new_n879_, new_n878_, new_n768_ );
or g774 ( new_n880_, new_n877_, new_n879_ );
or g775 ( new_n881_, new_n880_, new_n763_ );
not g776 ( new_n882_, new_n881_ );
and g777 ( new_n883_, new_n749_, keyIn_0_23 );
and g778 ( new_n884_, new_n883_, new_n746_ );
and g779 ( new_n885_, new_n882_, new_n884_ );
not g780 ( new_n886_, new_n885_ );
and g781 ( new_n887_, new_n863_, new_n563_ );
and g782 ( new_n888_, new_n886_, new_n887_ );
and g783 ( new_n889_, new_n888_, new_n873_ );
and g784 ( new_n890_, new_n889_, new_n872_ );
or g785 ( new_n891_, new_n871_, new_n890_ );
and g786 ( new_n892_, new_n891_, N117 );
or g787 ( new_n893_, new_n889_, new_n872_ );
not g788 ( new_n894_, new_n890_ );
and g789 ( new_n895_, new_n894_, new_n191_ );
and g790 ( new_n896_, new_n895_, new_n893_ );
or g791 ( N753, new_n892_, new_n896_ );
or g792 ( new_n898_, new_n793_, new_n864_ );
and g793 ( new_n899_, new_n898_, N121 );
not g794 ( new_n900_, new_n898_ );
and g795 ( new_n901_, new_n900_, new_n200_ );
or g796 ( N754, new_n901_, new_n899_ );
or g797 ( new_n903_, new_n799_, new_n864_ );
and g798 ( new_n904_, new_n903_, N125 );
not g799 ( new_n905_, new_n903_ );
and g800 ( new_n906_, new_n905_, new_n201_ );
or g801 ( N755, new_n906_, new_n904_ );
endmodule