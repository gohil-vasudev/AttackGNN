module add_mul_mix_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        c_0_, c_1_, c_2_, c_3_, d_0_, d_1_, d_2_, d_3_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, c_0_, c_1_, c_2_, c_3_,
         d_0_, d_1_, d_2_, d_3_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208;

  INV_X1 U108 ( .A(n101), .ZN(Result_7_) );
  XNOR2_X1 U109 ( .A(n102), .B(n103), .ZN(Result_6_) );
  NAND2_X1 U110 ( .A1(n104), .A2(n105), .ZN(n102) );
  XNOR2_X1 U111 ( .A(n106), .B(n107), .ZN(Result_5_) );
  NAND2_X1 U112 ( .A1(n108), .A2(n109), .ZN(n106) );
  XNOR2_X1 U113 ( .A(n110), .B(n111), .ZN(Result_4_) );
  XOR2_X1 U114 ( .A(n112), .B(n113), .Z(n111) );
  NAND2_X1 U115 ( .A1(n114), .A2(n105), .ZN(n113) );
  XOR2_X1 U116 ( .A(n115), .B(n116), .Z(Result_3_) );
  XOR2_X1 U117 ( .A(n117), .B(n118), .Z(Result_2_) );
  XNOR2_X1 U118 ( .A(n119), .B(n120), .ZN(Result_1_) );
  NAND2_X1 U119 ( .A1(n121), .A2(n122), .ZN(n120) );
  NAND3_X1 U120 ( .A1(n123), .A2(n121), .A3(n124), .ZN(Result_0_) );
  NAND2_X1 U121 ( .A1(n114), .A2(n125), .ZN(n124) );
  NAND4_X1 U122 ( .A1(n126), .A2(n127), .A3(n114), .A4(n128), .ZN(n121) );
  NOR2_X1 U123 ( .A1(n129), .A2(n125), .ZN(n128) );
  NAND2_X1 U124 ( .A1(n119), .A2(n122), .ZN(n123) );
  NAND3_X1 U125 ( .A1(n130), .A2(n131), .A3(n132), .ZN(n122) );
  NAND2_X1 U126 ( .A1(n133), .A2(n127), .ZN(n132) );
  OR2_X1 U127 ( .A1(n114), .A2(n134), .ZN(n131) );
  NAND3_X1 U128 ( .A1(n114), .A2(n126), .A3(n134), .ZN(n130) );
  INV_X1 U129 ( .A(n125), .ZN(n134) );
  NAND2_X1 U130 ( .A1(n135), .A2(n136), .ZN(n125) );
  NAND2_X1 U131 ( .A1(n126), .A2(n137), .ZN(n136) );
  NAND2_X1 U132 ( .A1(n138), .A2(n139), .ZN(n137) );
  NAND2_X1 U133 ( .A1(n140), .A2(n141), .ZN(n139) );
  NAND2_X1 U134 ( .A1(n142), .A2(n114), .ZN(n138) );
  AND2_X1 U135 ( .A1(n118), .A2(n117), .ZN(n119) );
  XOR2_X1 U136 ( .A(n127), .B(n133), .Z(n117) );
  INV_X1 U137 ( .A(n129), .ZN(n133) );
  XOR2_X1 U138 ( .A(n143), .B(n144), .Z(n129) );
  AND2_X1 U139 ( .A1(n126), .A2(n140), .ZN(n144) );
  NAND2_X1 U140 ( .A1(n135), .A2(n145), .ZN(n143) );
  NAND2_X1 U141 ( .A1(n146), .A2(n147), .ZN(n145) );
  NAND2_X1 U142 ( .A1(n148), .A2(n114), .ZN(n147) );
  INV_X1 U143 ( .A(n141), .ZN(n146) );
  NAND2_X1 U144 ( .A1(n114), .A2(n141), .ZN(n135) );
  NAND2_X1 U145 ( .A1(n149), .A2(n150), .ZN(n141) );
  NAND2_X1 U146 ( .A1(n151), .A2(n152), .ZN(n127) );
  NAND2_X1 U147 ( .A1(n153), .A2(n154), .ZN(n152) );
  AND2_X1 U148 ( .A1(n116), .A2(n115), .ZN(n118) );
  NAND2_X1 U149 ( .A1(n155), .A2(n156), .ZN(n115) );
  NAND3_X1 U150 ( .A1(n105), .A2(n157), .A3(n114), .ZN(n156) );
  OR2_X1 U151 ( .A1(n110), .A2(n112), .ZN(n157) );
  NAND2_X1 U152 ( .A1(n110), .A2(n112), .ZN(n155) );
  NAND2_X1 U153 ( .A1(n108), .A2(n158), .ZN(n112) );
  NAND2_X1 U154 ( .A1(n107), .A2(n109), .ZN(n158) );
  NAND2_X1 U155 ( .A1(n159), .A2(n160), .ZN(n109) );
  NAND2_X1 U156 ( .A1(n140), .A2(n105), .ZN(n160) );
  INV_X1 U157 ( .A(n161), .ZN(n159) );
  XNOR2_X1 U158 ( .A(n162), .B(n163), .ZN(n107) );
  AND2_X1 U159 ( .A1(n164), .A2(n148), .ZN(n163) );
  NAND2_X1 U160 ( .A1(n161), .A2(n140), .ZN(n108) );
  NOR2_X1 U161 ( .A1(n101), .A2(n162), .ZN(n161) );
  NAND2_X1 U162 ( .A1(n165), .A2(n104), .ZN(n162) );
  NAND2_X1 U163 ( .A1(n105), .A2(n164), .ZN(n101) );
  XOR2_X1 U164 ( .A(c_3_), .B(d_3_), .Z(n105) );
  XOR2_X1 U165 ( .A(n166), .B(n167), .Z(n110) );
  XNOR2_X1 U166 ( .A(n168), .B(n169), .ZN(n167) );
  NAND2_X1 U167 ( .A1(n140), .A2(n165), .ZN(n169) );
  XNOR2_X1 U168 ( .A(n170), .B(n153), .ZN(n116) );
  XOR2_X1 U169 ( .A(n171), .B(n149), .Z(n153) );
  NAND2_X1 U170 ( .A1(n172), .A2(n173), .ZN(n149) );
  NAND2_X1 U171 ( .A1(n150), .A2(n174), .ZN(n171) );
  NAND2_X1 U172 ( .A1(n175), .A2(n176), .ZN(n174) );
  NAND2_X1 U173 ( .A1(n126), .A2(n104), .ZN(n175) );
  NAND3_X1 U174 ( .A1(n126), .A2(n104), .A3(n142), .ZN(n150) );
  INV_X1 U175 ( .A(n176), .ZN(n142) );
  NAND2_X1 U176 ( .A1(n148), .A2(n140), .ZN(n176) );
  NAND2_X1 U177 ( .A1(n151), .A2(n154), .ZN(n170) );
  NAND2_X1 U178 ( .A1(n177), .A2(n178), .ZN(n154) );
  NAND2_X1 U179 ( .A1(n114), .A2(n165), .ZN(n178) );
  INV_X1 U180 ( .A(n179), .ZN(n177) );
  NAND2_X1 U181 ( .A1(n114), .A2(n179), .ZN(n151) );
  NAND2_X1 U182 ( .A1(n180), .A2(n181), .ZN(n179) );
  NAND3_X1 U183 ( .A1(n165), .A2(n182), .A3(n140), .ZN(n181) );
  XOR2_X1 U184 ( .A(n183), .B(n184), .Z(n140) );
  XOR2_X1 U185 ( .A(b_1_), .B(a_1_), .Z(n184) );
  OR2_X1 U186 ( .A1(n166), .A2(n168), .ZN(n182) );
  NAND2_X1 U187 ( .A1(n168), .A2(n166), .ZN(n180) );
  XOR2_X1 U188 ( .A(n172), .B(n173), .Z(n166) );
  AND2_X1 U189 ( .A1(n126), .A2(n164), .ZN(n172) );
  XNOR2_X1 U190 ( .A(n185), .B(n186), .ZN(n126) );
  XOR2_X1 U191 ( .A(d_0_), .B(c_0_), .Z(n186) );
  NAND2_X1 U192 ( .A1(n187), .A2(n188), .ZN(n185) );
  NAND2_X1 U193 ( .A1(n189), .A2(n190), .ZN(n188) );
  INV_X1 U194 ( .A(d_1_), .ZN(n190) );
  NAND2_X1 U195 ( .A1(c_1_), .A2(n191), .ZN(n189) );
  OR2_X1 U196 ( .A1(n191), .A2(c_1_), .ZN(n187) );
  AND2_X1 U197 ( .A1(n173), .A2(n103), .ZN(n168) );
  AND2_X1 U198 ( .A1(n165), .A2(n164), .ZN(n103) );
  XOR2_X1 U199 ( .A(a_3_), .B(b_3_), .Z(n164) );
  XNOR2_X1 U200 ( .A(n192), .B(n193), .ZN(n165) );
  XOR2_X1 U201 ( .A(d_2_), .B(c_2_), .Z(n193) );
  NAND2_X1 U202 ( .A1(c_3_), .A2(d_3_), .ZN(n192) );
  AND2_X1 U203 ( .A1(n148), .A2(n104), .ZN(n173) );
  XNOR2_X1 U204 ( .A(n194), .B(n195), .ZN(n104) );
  XOR2_X1 U205 ( .A(b_2_), .B(a_2_), .Z(n195) );
  NAND2_X1 U206 ( .A1(a_3_), .A2(b_3_), .ZN(n194) );
  XOR2_X1 U207 ( .A(n191), .B(n196), .Z(n148) );
  XOR2_X1 U208 ( .A(d_1_), .B(c_1_), .Z(n196) );
  NAND2_X1 U209 ( .A1(n197), .A2(n198), .ZN(n191) );
  NAND3_X1 U210 ( .A1(d_3_), .A2(n199), .A3(c_3_), .ZN(n198) );
  OR2_X1 U211 ( .A1(d_2_), .A2(c_2_), .ZN(n199) );
  NAND2_X1 U212 ( .A1(c_2_), .A2(d_2_), .ZN(n197) );
  XNOR2_X1 U213 ( .A(n200), .B(n201), .ZN(n114) );
  XOR2_X1 U214 ( .A(b_0_), .B(a_0_), .Z(n201) );
  NAND2_X1 U215 ( .A1(n202), .A2(n203), .ZN(n200) );
  NAND2_X1 U216 ( .A1(n204), .A2(n205), .ZN(n203) );
  INV_X1 U217 ( .A(b_1_), .ZN(n205) );
  NAND2_X1 U218 ( .A1(a_1_), .A2(n183), .ZN(n204) );
  OR2_X1 U219 ( .A1(n183), .A2(a_1_), .ZN(n202) );
  NAND2_X1 U220 ( .A1(n206), .A2(n207), .ZN(n183) );
  NAND3_X1 U221 ( .A1(b_3_), .A2(n208), .A3(a_3_), .ZN(n207) );
  OR2_X1 U222 ( .A1(b_2_), .A2(a_2_), .ZN(n208) );
  NAND2_X1 U223 ( .A1(a_2_), .A2(b_2_), .ZN(n206) );
endmodule

