module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n556_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n451_, new_n489_, new_n424_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n462_, new_n564_, new_n500_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n449_, new_n364_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n350_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n137_, new_n183_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n180_, new_n530_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n314_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n562_, new_n485_, new_n525_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n570_, new_n143_, new_n520_, new_n125_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n507_, new_n182_, new_n407_, new_n480_, new_n151_, new_n513_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n522_, new_n428_, new_n199_, new_n487_, new_n360_, new_n546_, new_n302_, new_n191_, new_n225_, new_n544_, new_n476_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n440_, new_n531_, new_n252_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n134_, new_n433_, new_n435_, new_n265_, new_n370_, new_n278_, new_n304_, new_n523_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n412_, new_n327_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n195_, new_n567_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n322_, new_n228_, new_n545_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

nand g000 ( new_n119_, N29, N42, N75 );
not g001 ( N388, new_n119_ );
nand g002 ( new_n121_, N29, N36, N80 );
not g003 ( N389, new_n121_ );
nand g004 ( new_n123_, N29, N36, N42 );
not g005 ( N390, new_n123_ );
nand g006 ( new_n125_, N85, N86 );
not g007 ( N391, new_n125_ );
nand g008 ( new_n127_, N1, N8 );
not g009 ( new_n128_, new_n127_ );
nand g010 ( new_n129_, new_n128_, N13, N17 );
not g011 ( N418, new_n129_ );
not g012 ( new_n131_, keyIn_0_0 );
nand g013 ( new_n132_, N390, new_n131_ );
nand g014 ( new_n133_, new_n123_, keyIn_0_0 );
nand g015 ( new_n134_, new_n132_, new_n133_ );
not g016 ( new_n135_, N13 );
not g017 ( new_n136_, N17 );
nand g018 ( new_n137_, N1, N26 );
nor g019 ( new_n138_, new_n137_, new_n135_, new_n136_ );
nand g020 ( N419, new_n134_, new_n138_ );
nand g021 ( N420, N59, N75, N80 );
nand g022 ( N421, N36, N59, N80 );
nand g023 ( N422, N36, N42, N59 );
not g024 ( new_n143_, N90 );
nor g025 ( new_n144_, N87, N88 );
nor g026 ( N423, new_n144_, new_n143_ );
nand g027 ( N446, new_n132_, new_n133_, new_n138_ );
nand g028 ( new_n147_, N1, N26, N51 );
not g029 ( N447, new_n147_ );
nand g030 ( new_n149_, new_n128_, N13, N55 );
nand g031 ( new_n150_, N29, N68 );
nor g032 ( new_n151_, new_n150_, keyIn_0_1 );
nand g033 ( new_n152_, new_n150_, keyIn_0_1 );
not g034 ( new_n153_, new_n152_ );
nor g035 ( N448, new_n149_, new_n153_, new_n151_ );
not g036 ( new_n155_, N74 );
nand g037 ( new_n156_, N59, N68 );
nor g038 ( N449, new_n149_, new_n155_, new_n156_ );
not g039 ( new_n158_, N89 );
nor g040 ( N450, new_n144_, new_n158_ );
not g041 ( new_n160_, keyIn_0_2 );
nand g042 ( new_n161_, N101, N106 );
nand g043 ( new_n162_, new_n161_, new_n160_ );
nand g044 ( new_n163_, keyIn_0_2, N101, N106 );
nand g045 ( new_n164_, new_n162_, new_n163_ );
not g046 ( new_n165_, N101 );
not g047 ( new_n166_, N106 );
nand g048 ( new_n167_, new_n165_, new_n166_ );
nand g049 ( new_n168_, new_n164_, new_n167_ );
not g050 ( new_n169_, new_n168_ );
nand g051 ( new_n170_, N91, N96 );
not g052 ( new_n171_, new_n170_ );
nor g053 ( new_n172_, N91, N96 );
nor g054 ( new_n173_, new_n171_, new_n172_ );
nand g055 ( new_n174_, new_n169_, keyIn_0_7, new_n173_ );
not g056 ( new_n175_, new_n173_ );
nand g057 ( new_n176_, new_n168_, new_n175_ );
not g058 ( new_n177_, keyIn_0_7 );
nand g059 ( new_n178_, new_n169_, new_n173_ );
nand g060 ( new_n179_, new_n178_, new_n177_ );
nand g061 ( new_n180_, new_n179_, N130, new_n174_, new_n176_ );
nand g062 ( new_n181_, new_n180_, keyIn_0_9 );
not g063 ( new_n182_, new_n181_ );
nor g064 ( new_n183_, new_n180_, keyIn_0_9 );
nor g065 ( new_n184_, new_n182_, new_n183_ );
not g066 ( new_n185_, new_n184_ );
not g067 ( new_n186_, keyIn_0_10 );
not g068 ( new_n187_, N130 );
nand g069 ( new_n188_, new_n179_, new_n174_, new_n176_ );
nand g070 ( new_n189_, new_n188_, new_n187_ );
nand g071 ( new_n190_, new_n189_, new_n186_ );
nand g072 ( new_n191_, new_n188_, keyIn_0_10, new_n187_ );
nand g073 ( new_n192_, new_n185_, new_n190_, new_n191_ );
not g074 ( new_n193_, new_n192_ );
not g075 ( new_n194_, N135 );
not g076 ( new_n195_, N111 );
not g077 ( new_n196_, N116 );
nand g078 ( new_n197_, new_n195_, new_n196_ );
nand g079 ( new_n198_, N111, N116 );
nand g080 ( new_n199_, new_n197_, new_n198_ );
not g081 ( new_n200_, N121 );
not g082 ( new_n201_, N126 );
nand g083 ( new_n202_, new_n200_, new_n201_ );
nand g084 ( new_n203_, N121, N126 );
nand g085 ( new_n204_, new_n202_, new_n203_ );
nand g086 ( new_n205_, new_n199_, new_n204_ );
nand g087 ( new_n206_, new_n197_, new_n202_, new_n198_, new_n203_ );
nand g088 ( new_n207_, new_n205_, new_n206_ );
nand g089 ( new_n208_, new_n207_, new_n194_ );
nand g090 ( new_n209_, new_n205_, N135, new_n206_ );
nand g091 ( new_n210_, new_n208_, new_n209_ );
not g092 ( new_n211_, new_n210_ );
nor g093 ( new_n212_, new_n193_, new_n211_ );
nor g094 ( new_n213_, new_n192_, new_n210_ );
nor g095 ( N767, new_n212_, new_n213_ );
not g096 ( new_n215_, keyIn_0_5 );
nand g097 ( new_n216_, N183, N189 );
not g098 ( new_n217_, new_n216_ );
nor g099 ( new_n218_, N183, N189 );
nor g100 ( new_n219_, new_n217_, new_n218_ );
not g101 ( new_n220_, new_n219_ );
nand g102 ( new_n221_, new_n220_, new_n215_ );
nand g103 ( new_n222_, new_n221_, keyIn_0_6 );
nand g104 ( new_n223_, N195, N201 );
not g105 ( new_n224_, new_n223_ );
nor g106 ( new_n225_, N195, N201 );
nor g107 ( new_n226_, new_n224_, new_n225_ );
nand g108 ( new_n227_, new_n222_, new_n226_ );
not g109 ( new_n228_, new_n226_ );
nand g110 ( new_n229_, new_n228_, keyIn_0_6 );
nand g111 ( new_n230_, new_n229_, new_n215_ );
nand g112 ( new_n231_, new_n230_, new_n219_ );
nand g113 ( new_n232_, new_n227_, new_n231_ );
nand g114 ( new_n233_, new_n232_, N207 );
not g115 ( new_n234_, N207 );
nand g116 ( new_n235_, new_n227_, new_n231_, new_n234_ );
nand g117 ( new_n236_, new_n233_, new_n235_ );
not g118 ( new_n237_, N159 );
not g119 ( new_n238_, N165 );
nand g120 ( new_n239_, new_n237_, new_n238_ );
nand g121 ( new_n240_, N159, N165 );
nand g122 ( new_n241_, new_n239_, new_n240_ );
not g123 ( new_n242_, N171 );
not g124 ( new_n243_, N177 );
nand g125 ( new_n244_, new_n242_, new_n243_ );
nand g126 ( new_n245_, N171, N177 );
nand g127 ( new_n246_, new_n244_, new_n245_ );
nand g128 ( new_n247_, new_n241_, new_n246_ );
nand g129 ( new_n248_, new_n239_, new_n244_, new_n240_, new_n245_ );
nand g130 ( new_n249_, new_n247_, new_n248_ );
nand g131 ( new_n250_, new_n249_, keyIn_0_12, new_n187_ );
not g132 ( new_n251_, keyIn_0_12 );
nand g133 ( new_n252_, new_n249_, new_n187_ );
nand g134 ( new_n253_, new_n252_, new_n251_ );
not g135 ( new_n254_, keyIn_0_15 );
nand g136 ( new_n255_, new_n247_, N130, new_n248_ );
nand g137 ( new_n256_, new_n255_, new_n254_ );
not g138 ( new_n257_, new_n256_ );
nand g139 ( new_n258_, new_n257_, new_n253_, new_n250_ );
not g140 ( new_n259_, new_n258_ );
nand g141 ( new_n260_, new_n236_, new_n259_ );
nand g142 ( new_n261_, new_n233_, new_n235_, new_n258_ );
nand g143 ( N768, new_n260_, new_n261_ );
not g144 ( new_n263_, keyIn_0_11 );
nand g145 ( new_n264_, N59, N156 );
not g146 ( new_n265_, new_n264_ );
nand g147 ( new_n266_, N17, N42 );
not g148 ( new_n267_, N42 );
nand g149 ( new_n268_, new_n136_, new_n267_ );
nand g150 ( new_n269_, N447, new_n265_, new_n268_, new_n266_ );
not g151 ( new_n270_, keyIn_0_4 );
nand g152 ( new_n271_, N1, N8, N17, N51 );
nand g153 ( new_n272_, new_n271_, new_n270_ );
nand g154 ( new_n273_, N17, N51 );
not g155 ( new_n274_, new_n273_ );
nand g156 ( new_n275_, new_n128_, new_n274_, keyIn_0_4 );
nand g157 ( new_n276_, N42, N59, N75 );
nand g158 ( new_n277_, new_n275_, new_n272_, new_n276_ );
nand g159 ( new_n278_, new_n277_, new_n269_ );
nand g160 ( new_n279_, new_n278_, N126 );
nand g161 ( new_n280_, new_n279_, new_n263_ );
nand g162 ( new_n281_, new_n278_, keyIn_0_11, N126 );
nand g163 ( new_n282_, new_n280_, new_n281_ );
not g164 ( new_n283_, N153 );
not g165 ( new_n284_, N1 );
nor g166 ( new_n285_, new_n265_, new_n147_, new_n136_ );
nor g167 ( new_n286_, new_n285_, new_n284_ );
nor g168 ( new_n287_, new_n286_, new_n283_ );
nand g169 ( new_n288_, N447, N55 );
not g170 ( new_n289_, N268 );
nand g171 ( new_n290_, new_n289_, N29, N75, N80 );
nor g172 ( new_n291_, new_n288_, new_n290_ );
nor g173 ( new_n292_, new_n287_, new_n291_ );
nand g174 ( new_n293_, new_n282_, new_n292_ );
nand g175 ( new_n294_, new_n293_, N201 );
not g176 ( new_n295_, N201 );
nand g177 ( new_n296_, new_n282_, new_n295_, new_n292_ );
nand g178 ( new_n297_, new_n294_, new_n296_ );
not g179 ( new_n298_, new_n297_ );
nand g180 ( new_n299_, new_n298_, N261 );
not g181 ( new_n300_, N261 );
nand g182 ( new_n301_, new_n297_, new_n300_ );
nand g183 ( new_n302_, new_n299_, N219, new_n301_ );
nand g184 ( new_n303_, new_n293_, N246 );
nand g185 ( new_n304_, N255, N267 );
nand g186 ( new_n305_, new_n303_, new_n304_ );
nand g187 ( new_n306_, new_n305_, keyIn_0_19 );
nand g188 ( new_n307_, new_n293_, N201, N237 );
nand g189 ( new_n308_, N121, N210 );
nand g190 ( new_n309_, N42, N72, N73 );
nor g191 ( new_n310_, new_n149_, new_n309_, new_n156_ );
nand g192 ( new_n311_, new_n310_, N201 );
nand g193 ( new_n312_, new_n306_, new_n307_, new_n308_, new_n311_ );
not g194 ( new_n313_, new_n312_ );
nand g195 ( new_n314_, new_n298_, N228 );
not g196 ( new_n315_, keyIn_0_19 );
nand g197 ( new_n316_, new_n303_, new_n315_, new_n304_ );
nand g198 ( N850, new_n313_, new_n302_, new_n314_, new_n316_ );
not g199 ( new_n318_, keyIn_0_24 );
not g200 ( new_n319_, N189 );
not g201 ( new_n320_, keyIn_0_13 );
not g202 ( new_n321_, new_n291_ );
nand g203 ( new_n322_, new_n278_, N116 );
not g204 ( new_n323_, new_n286_ );
nand g205 ( new_n324_, new_n323_, N146 );
nand g206 ( new_n325_, new_n322_, new_n324_, new_n321_ );
nand g207 ( new_n326_, new_n325_, new_n320_ );
nand g208 ( new_n327_, new_n322_, new_n324_, keyIn_0_13, new_n321_ );
nand g209 ( new_n328_, new_n326_, new_n319_, new_n327_ );
nand g210 ( new_n329_, new_n296_, N261 );
nand g211 ( new_n330_, new_n329_, new_n294_ );
not g212 ( new_n331_, N195 );
not g213 ( new_n332_, keyIn_0_14 );
nand g214 ( new_n333_, new_n278_, N121 );
nand g215 ( new_n334_, new_n323_, N149 );
nand g216 ( new_n335_, new_n333_, new_n334_, new_n321_ );
nand g217 ( new_n336_, new_n335_, new_n332_ );
nand g218 ( new_n337_, new_n333_, new_n334_, keyIn_0_14, new_n321_ );
nand g219 ( new_n338_, new_n336_, new_n337_ );
nand g220 ( new_n339_, new_n338_, new_n331_ );
nand g221 ( new_n340_, new_n330_, new_n328_, new_n339_ );
not g222 ( new_n341_, keyIn_0_22 );
nand g223 ( new_n342_, new_n326_, new_n327_ );
nand g224 ( new_n343_, new_n342_, N189 );
not g225 ( new_n344_, new_n343_ );
nand g226 ( new_n345_, new_n344_, new_n341_ );
nand g227 ( new_n346_, new_n343_, keyIn_0_22 );
not g228 ( new_n347_, new_n338_ );
nand g229 ( new_n348_, new_n347_, N195, new_n328_ );
nand g230 ( new_n349_, new_n340_, new_n345_, new_n346_, new_n348_ );
nand g231 ( new_n350_, new_n349_, new_n318_ );
nand g232 ( new_n351_, new_n348_, new_n346_ );
not g233 ( new_n352_, new_n351_ );
nand g234 ( new_n353_, new_n352_, keyIn_0_24, new_n340_, new_n345_ );
nand g235 ( new_n354_, new_n350_, new_n353_ );
not g236 ( new_n355_, keyIn_0_17 );
not g237 ( new_n356_, N183 );
nand g238 ( new_n357_, new_n278_, N111 );
not g239 ( new_n358_, new_n357_ );
not g240 ( new_n359_, N143 );
nor g241 ( new_n360_, new_n286_, new_n359_ );
nor g242 ( new_n361_, new_n358_, new_n291_, new_n360_ );
nand g243 ( new_n362_, new_n361_, new_n356_ );
nand g244 ( new_n363_, new_n362_, new_n355_ );
nand g245 ( new_n364_, new_n361_, keyIn_0_17, new_n356_ );
nand g246 ( new_n365_, new_n363_, new_n364_ );
not g247 ( new_n366_, new_n365_ );
not g248 ( new_n367_, new_n361_ );
nand g249 ( new_n368_, new_n367_, N183 );
nand g250 ( new_n369_, new_n366_, new_n368_ );
nand g251 ( new_n370_, new_n354_, new_n369_ );
not g252 ( new_n371_, new_n369_ );
nand g253 ( new_n372_, new_n350_, new_n353_, new_n371_ );
nand g254 ( new_n373_, new_n370_, N219, new_n372_ );
nand g255 ( new_n374_, new_n371_, N228 );
not g256 ( new_n375_, keyIn_0_18 );
nand g257 ( new_n376_, new_n368_, new_n375_ );
nand g258 ( new_n377_, new_n367_, keyIn_0_18, N183 );
nand g259 ( new_n378_, new_n376_, N237, new_n377_ );
nand g260 ( new_n379_, new_n367_, N246 );
nand g261 ( new_n380_, new_n310_, N183 );
nand g262 ( new_n381_, N106, N210 );
nand g263 ( new_n382_, new_n381_, keyIn_0_3 );
not g264 ( new_n383_, keyIn_0_3 );
nand g265 ( new_n384_, new_n383_, N106, N210 );
nand g266 ( new_n385_, new_n379_, new_n380_, new_n382_, new_n384_ );
not g267 ( new_n386_, new_n385_ );
nand g268 ( N863, new_n373_, new_n374_, new_n378_, new_n386_ );
not g269 ( new_n388_, keyIn_0_27 );
nand g270 ( new_n389_, new_n330_, new_n339_ );
nand g271 ( new_n390_, new_n347_, N195 );
nand g272 ( new_n391_, new_n389_, new_n390_ );
nand g273 ( new_n392_, new_n343_, new_n328_ );
not g274 ( new_n393_, new_n392_ );
nand g275 ( new_n394_, new_n391_, new_n393_ );
nand g276 ( new_n395_, new_n389_, new_n390_, new_n392_ );
nand g277 ( new_n396_, new_n394_, N219, new_n395_ );
nand g278 ( new_n397_, new_n393_, N228 );
not g279 ( new_n398_, new_n397_ );
nand g280 ( new_n399_, new_n344_, N237 );
not g281 ( new_n400_, new_n399_ );
nand g282 ( new_n401_, new_n342_, N246 );
nand g283 ( new_n402_, new_n310_, N189 );
nand g284 ( new_n403_, N111, N210 );
nand g285 ( new_n404_, N255, N259 );
nand g286 ( new_n405_, new_n401_, new_n402_, new_n403_, new_n404_ );
nor g287 ( new_n406_, new_n398_, new_n400_, new_n405_ );
nand g288 ( new_n407_, new_n406_, new_n396_ );
nand g289 ( new_n408_, new_n407_, new_n388_ );
nand g290 ( new_n409_, new_n406_, new_n396_, keyIn_0_27 );
nand g291 ( new_n410_, new_n408_, new_n409_ );
not g292 ( N864, new_n410_ );
not g293 ( new_n412_, keyIn_0_28 );
not g294 ( new_n413_, new_n330_ );
nand g295 ( new_n414_, new_n390_, new_n339_ );
nor g296 ( new_n415_, new_n414_, new_n413_ );
not g297 ( new_n416_, new_n415_ );
nand g298 ( new_n417_, new_n416_, keyIn_0_25 );
not g299 ( new_n418_, keyIn_0_25 );
nand g300 ( new_n419_, new_n415_, new_n418_ );
nand g301 ( new_n420_, new_n417_, new_n419_ );
nand g302 ( new_n421_, new_n414_, new_n413_ );
nand g303 ( new_n422_, new_n420_, N219, new_n421_ );
nand g304 ( new_n423_, new_n390_, N228, new_n339_ );
not g305 ( new_n424_, new_n423_ );
nand g306 ( new_n425_, new_n347_, N195, N237 );
not g307 ( new_n426_, new_n425_ );
nand g308 ( new_n427_, new_n347_, N246 );
nand g309 ( new_n428_, new_n310_, N195 );
nand g310 ( new_n429_, N116, N210 );
nand g311 ( new_n430_, N255, N260 );
nand g312 ( new_n431_, new_n427_, new_n428_, new_n429_, new_n430_ );
nor g313 ( new_n432_, new_n424_, new_n426_, new_n431_ );
nand g314 ( new_n433_, new_n422_, new_n432_ );
nand g315 ( new_n434_, new_n433_, new_n412_ );
nand g316 ( new_n435_, new_n422_, keyIn_0_28, new_n432_ );
nand g317 ( new_n436_, new_n434_, new_n435_ );
not g318 ( N865, new_n436_ );
nand g319 ( new_n438_, new_n376_, new_n377_ );
nand g320 ( new_n439_, new_n350_, new_n353_, new_n366_ );
nand g321 ( new_n440_, new_n439_, new_n438_ );
nand g322 ( new_n441_, new_n278_, N106 );
nand g323 ( new_n442_, N447, N55, new_n264_ );
nor g324 ( new_n443_, new_n442_, new_n283_ );
nor g325 ( new_n444_, new_n290_, new_n136_, new_n147_ );
nand g326 ( new_n445_, N138, N152 );
not g327 ( new_n446_, new_n445_ );
nor g328 ( new_n447_, new_n443_, new_n444_, new_n446_ );
nand g329 ( new_n448_, new_n441_, new_n447_, new_n243_ );
nand g330 ( new_n449_, new_n440_, new_n448_ );
nand g331 ( new_n450_, new_n441_, new_n447_ );
nand g332 ( new_n451_, new_n450_, N177 );
nand g333 ( new_n452_, new_n449_, new_n451_ );
nand g334 ( new_n453_, new_n278_, N101 );
not g335 ( new_n454_, N149 );
nor g336 ( new_n455_, new_n442_, new_n454_ );
nand g337 ( new_n456_, N17, N138 );
not g338 ( new_n457_, new_n456_ );
nor g339 ( new_n458_, new_n455_, new_n444_, new_n457_ );
nand g340 ( new_n459_, new_n453_, new_n458_, new_n242_ );
nand g341 ( new_n460_, new_n452_, new_n459_ );
nand g342 ( new_n461_, new_n453_, new_n458_ );
nand g343 ( new_n462_, new_n461_, N171 );
nand g344 ( new_n463_, new_n460_, new_n462_ );
nand g345 ( new_n464_, new_n278_, N96 );
not g346 ( new_n465_, N146 );
nor g347 ( new_n466_, new_n442_, new_n465_ );
nand g348 ( new_n467_, N51, N138 );
not g349 ( new_n468_, new_n467_ );
nor g350 ( new_n469_, new_n466_, new_n444_, new_n468_ );
nand g351 ( new_n470_, new_n464_, new_n469_, new_n238_ );
nand g352 ( new_n471_, new_n463_, new_n470_ );
nand g353 ( new_n472_, new_n464_, new_n469_ );
nand g354 ( new_n473_, new_n472_, N165 );
nand g355 ( new_n474_, new_n473_, keyIn_0_16 );
not g356 ( new_n475_, keyIn_0_16 );
nand g357 ( new_n476_, new_n472_, new_n475_, N165 );
nand g358 ( new_n477_, new_n474_, new_n476_ );
not g359 ( new_n478_, new_n477_ );
nand g360 ( new_n479_, new_n471_, new_n478_ );
nand g361 ( new_n480_, new_n278_, N91 );
not g362 ( new_n481_, new_n444_ );
nand g363 ( new_n482_, new_n481_, keyIn_0_8 );
not g364 ( new_n483_, keyIn_0_8 );
nand g365 ( new_n484_, new_n444_, new_n483_ );
nand g366 ( new_n485_, new_n482_, new_n484_ );
nor g367 ( new_n486_, new_n442_, new_n359_ );
nand g368 ( new_n487_, N8, N138 );
not g369 ( new_n488_, new_n487_ );
nor g370 ( new_n489_, new_n486_, new_n488_ );
nand g371 ( new_n490_, new_n485_, new_n480_, new_n237_, new_n489_ );
nand g372 ( new_n491_, new_n479_, new_n490_ );
nand g373 ( new_n492_, new_n485_, new_n480_, new_n489_ );
nand g374 ( new_n493_, new_n492_, N159 );
nand g375 ( N866, new_n491_, new_n493_ );
nand g376 ( new_n495_, new_n451_, new_n448_ );
not g377 ( new_n496_, new_n495_ );
nand g378 ( new_n497_, new_n440_, new_n496_ );
nand g379 ( new_n498_, new_n439_, new_n438_, new_n495_ );
nand g380 ( new_n499_, new_n497_, N219, new_n498_ );
not g381 ( new_n500_, keyIn_0_23 );
nand g382 ( new_n501_, new_n496_, N228 );
nand g383 ( new_n502_, new_n450_, N177, N237 );
nand g384 ( new_n503_, new_n501_, new_n500_, new_n502_ );
nand g385 ( new_n504_, new_n501_, new_n502_ );
nand g386 ( new_n505_, new_n504_, keyIn_0_23 );
nand g387 ( new_n506_, new_n450_, N246 );
nand g388 ( new_n507_, N101, N210 );
nand g389 ( new_n508_, new_n310_, N177 );
nand g390 ( new_n509_, new_n506_, new_n507_, new_n508_ );
not g391 ( new_n510_, new_n509_ );
nand g392 ( N874, new_n499_, new_n503_, new_n505_, new_n510_ );
not g393 ( new_n512_, keyIn_0_31 );
nand g394 ( new_n513_, new_n493_, new_n490_ );
not g395 ( new_n514_, new_n513_ );
nand g396 ( new_n515_, new_n479_, new_n514_ );
nand g397 ( new_n516_, new_n471_, new_n478_, new_n513_ );
nand g398 ( new_n517_, new_n515_, N219, new_n516_ );
not g399 ( new_n518_, keyIn_0_20 );
nand g400 ( new_n519_, new_n514_, new_n518_, N228 );
nand g401 ( new_n520_, new_n514_, N228 );
nand g402 ( new_n521_, new_n520_, keyIn_0_20 );
nand g403 ( new_n522_, new_n492_, N159, N237 );
nand g404 ( new_n523_, new_n492_, N246 );
nand g405 ( new_n524_, N210, N268 );
nand g406 ( new_n525_, new_n310_, N159 );
nand g407 ( new_n526_, new_n522_, new_n523_, new_n524_, new_n525_ );
not g408 ( new_n527_, new_n526_ );
nand g409 ( new_n528_, new_n521_, new_n519_, new_n527_ );
not g410 ( new_n529_, new_n528_ );
nand g411 ( new_n530_, new_n517_, new_n529_ );
nand g412 ( new_n531_, new_n530_, new_n512_ );
nand g413 ( new_n532_, new_n517_, keyIn_0_31, new_n529_ );
nand g414 ( new_n533_, new_n531_, new_n532_ );
not g415 ( N878, new_n533_ );
not g416 ( new_n535_, keyIn_0_29 );
nand g417 ( new_n536_, new_n478_, new_n470_ );
not g418 ( new_n537_, new_n536_ );
nand g419 ( new_n538_, new_n463_, new_n537_ );
nand g420 ( new_n539_, new_n460_, new_n462_, new_n536_ );
nand g421 ( new_n540_, new_n538_, new_n535_, N219, new_n539_ );
nand g422 ( new_n541_, new_n538_, N219, new_n539_ );
nand g423 ( new_n542_, new_n541_, keyIn_0_29 );
not g424 ( new_n543_, keyIn_0_21 );
nand g425 ( new_n544_, new_n537_, N228 );
nand g426 ( new_n545_, new_n544_, new_n543_ );
nor g427 ( new_n546_, new_n544_, new_n543_ );
nand g428 ( new_n547_, new_n477_, N237 );
nand g429 ( new_n548_, new_n472_, N246 );
nand g430 ( new_n549_, N91, N210 );
nand g431 ( new_n550_, new_n310_, N165 );
nand g432 ( new_n551_, new_n547_, new_n548_, new_n549_, new_n550_ );
nor g433 ( new_n552_, new_n546_, new_n551_ );
nand g434 ( N879, new_n542_, new_n540_, new_n545_, new_n552_ );
not g435 ( new_n554_, keyIn_0_30 );
nand g436 ( new_n555_, new_n462_, new_n459_ );
not g437 ( new_n556_, new_n555_ );
nand g438 ( new_n557_, new_n452_, new_n556_ );
nand g439 ( new_n558_, new_n449_, new_n451_, new_n555_ );
nand g440 ( new_n559_, new_n557_, keyIn_0_26, new_n558_ );
not g441 ( new_n560_, keyIn_0_26 );
nand g442 ( new_n561_, new_n557_, new_n558_ );
nand g443 ( new_n562_, new_n561_, new_n560_ );
nand g444 ( new_n563_, new_n562_, N219, new_n559_ );
nand g445 ( new_n564_, new_n556_, N228 );
not g446 ( new_n565_, new_n564_ );
nand g447 ( new_n566_, new_n461_, N171, N237 );
nand g448 ( new_n567_, new_n461_, N246 );
nand g449 ( new_n568_, N96, N210 );
nand g450 ( new_n569_, new_n310_, N171 );
nand g451 ( new_n570_, new_n566_, new_n567_, new_n568_, new_n569_ );
nor g452 ( new_n571_, new_n565_, new_n570_ );
nand g453 ( new_n572_, new_n563_, new_n571_ );
nand g454 ( new_n573_, new_n572_, new_n554_ );
nand g455 ( new_n574_, new_n563_, keyIn_0_30, new_n571_ );
nand g456 ( new_n575_, new_n573_, new_n574_ );
not g457 ( N880, new_n575_ );
endmodule