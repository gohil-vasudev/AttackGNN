module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n155_, new_n384_, new_n595_, new_n410_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n543_, new_n250_, new_n501_, new_n288_, new_n371_, new_n509_, new_n454_, new_n421_, new_n202_, new_n296_, new_n308_, new_n620_, new_n232_, new_n258_, new_n439_, new_n176_, new_n283_, new_n223_, new_n390_, new_n306_, new_n494_, new_n366_, new_n291_, new_n261_, new_n241_, new_n309_, new_n566_, new_n186_, new_n339_, new_n365_, new_n616_, new_n197_, new_n529_, new_n386_, new_n323_, new_n401_, new_n389_, new_n259_, new_n362_, new_n514_, new_n601_, new_n604_, new_n556_, new_n227_, new_n416_, new_n222_, new_n456_, new_n170_, new_n246_, new_n571_, new_n400_, new_n328_, new_n460_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n130_, new_n505_, new_n619_, new_n419_, new_n471_, new_n268_, new_n374_, new_n577_, new_n534_, new_n376_, new_n380_, new_n214_, new_n451_, new_n489_, new_n424_, new_n138_, new_n310_, new_n602_, new_n144_, new_n275_, new_n188_, new_n240_, new_n413_, new_n526_, new_n352_, new_n442_, new_n575_, new_n525_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n578_, new_n462_, new_n603_, new_n564_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n500_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n317_, new_n344_, new_n143_, new_n520_, new_n125_, new_n253_, new_n504_, new_n403_, new_n475_, new_n237_, new_n427_, new_n234_, new_n532_, new_n472_, new_n557_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n411_, new_n215_, new_n507_, new_n152_, new_n605_, new_n157_, new_n182_, new_n407_, new_n480_, new_n133_, new_n257_, new_n481_, new_n212_, new_n151_, new_n513_, new_n592_, new_n364_, new_n449_, new_n580_, new_n484_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n272_, new_n282_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n487_, new_n360_, new_n546_, new_n612_, new_n315_, new_n302_, new_n191_, new_n326_, new_n554_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n387_, new_n606_, new_n544_, new_n476_, new_n615_, new_n589_, new_n248_, new_n350_, new_n415_, new_n167_, new_n537_, new_n221_, new_n385_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n478_, new_n461_, new_n459_, new_n569_, new_n555_, new_n174_, new_n297_, new_n361_, new_n565_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n340_, new_n147_, new_n510_, new_n285_, new_n502_, new_n613_, new_n351_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n517_, new_n325_, new_n609_, new_n591_, new_n515_, new_n530_, new_n332_, new_n318_, new_n622_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n531_, new_n593_, new_n158_, new_n252_, new_n585_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n312_, new_n271_, new_n535_, new_n274_, new_n372_, new_n242_, new_n503_, new_n527_, new_n218_, new_n497_, new_n307_, new_n190_, new_n305_, new_n420_, new_n568_, new_n597_, new_n408_, new_n470_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n213_, new_n433_, new_n435_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n265_, new_n506_, new_n370_, new_n256_, new_n584_, new_n452_, new_n278_, new_n304_, new_n381_, new_n523_, new_n388_, new_n550_, new_n217_, new_n269_, new_n508_, new_n512_, new_n194_, new_n483_, new_n394_, new_n299_, new_n129_, new_n599_, new_n314_, new_n582_, new_n363_, new_n412_, new_n607_, new_n165_, new_n441_, new_n477_, new_n327_, new_n216_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n280_, new_n574_, new_n426_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n338_, new_n207_, new_n267_, new_n473_, new_n140_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n587_, new_n465_, new_n195_, new_n567_, new_n263_, new_n334_, new_n331_, new_n576_, new_n341_, new_n378_, new_n621_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n245_, new_n402_, new_n474_, new_n579_, new_n467_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n490_, new_n560_, new_n346_, new_n396_, new_n198_, new_n438_, new_n358_, new_n208_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n528_, new_n179_, new_n572_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n185_, new_n399_, new_n596_, new_n373_, new_n559_, new_n540_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n233_, new_n136_, new_n469_, new_n284_, new_n119_, new_n391_, new_n293_, new_n178_, new_n437_, new_n551_, new_n168_, new_n279_, new_n455_, new_n295_, new_n359_, new_n132_, new_n618_, new_n120_, new_n521_, new_n166_, new_n409_, new_n457_, new_n161_, new_n553_, new_n406_, new_n356_, new_n333_, new_n229_, new_n536_, new_n290_, new_n464_, new_n204_, new_n369_, new_n181_, new_n135_, new_n448_, new_n573_, new_n276_, new_n405_;

not g000 ( new_n119_, N75 );
nand g001 ( new_n120_, N29, N42 );
nor g002 ( N388, new_n120_, new_n119_ );
not g003 ( new_n122_, N80 );
nand g004 ( new_n123_, N29, N36 );
nor g005 ( N389, new_n123_, new_n122_ );
not g006 ( new_n125_, N42 );
nor g007 ( N390, new_n123_, new_n125_ );
nand g008 ( new_n127_, N85, N86 );
not g009 ( N391, new_n127_ );
not g010 ( new_n129_, N17 );
not g011 ( new_n130_, N13 );
nand g012 ( new_n131_, N1, N8 );
nor g013 ( new_n132_, new_n131_, new_n130_ );
not g014 ( new_n133_, new_n132_ );
nor g015 ( N418, new_n133_, new_n129_ );
not g016 ( new_n135_, N390 );
nand g017 ( new_n136_, N1, N26 );
nand g018 ( new_n137_, N13, N17 );
nor g019 ( new_n138_, new_n136_, new_n137_ );
nand g020 ( N419, new_n135_, new_n138_ );
nand g021 ( new_n140_, N59, N75 );
not g022 ( new_n141_, new_n140_ );
nand g023 ( N420, new_n141_, N80 );
nand g024 ( new_n143_, N36, N59 );
not g025 ( new_n144_, new_n143_ );
nand g026 ( N421, new_n144_, N80 );
nand g027 ( N422, new_n144_, N42 );
not g028 ( new_n147_, N90 );
nor g029 ( new_n148_, N87, N88 );
nor g030 ( N423, new_n148_, new_n147_ );
nand g031 ( N446, new_n138_, N390 );
not g032 ( new_n151_, N51 );
nor g033 ( new_n152_, new_n136_, new_n151_ );
xnor g034 ( N447, new_n152_, keyIn_0_0 );
nand g035 ( new_n154_, new_n132_, N55 );
nand g036 ( new_n155_, N29, N68 );
nor g037 ( N448, new_n154_, new_n155_ );
nand g038 ( new_n157_, N59, N68 );
not g039 ( new_n158_, new_n157_ );
nand g040 ( new_n159_, new_n158_, N74 );
nor g041 ( N449, new_n154_, new_n159_ );
not g042 ( new_n161_, N89 );
nor g043 ( N450, new_n148_, new_n161_ );
xor g044 ( new_n163_, N111, N116 );
xnor g045 ( new_n164_, N121, N126 );
xnor g046 ( new_n165_, new_n163_, new_n164_ );
xnor g047 ( new_n166_, new_n165_, N135 );
xnor g048 ( new_n167_, N91, N96 );
xnor g049 ( new_n168_, N101, N106 );
xnor g050 ( new_n169_, new_n167_, new_n168_ );
xnor g051 ( new_n170_, new_n169_, N130 );
xnor g052 ( N767, new_n166_, new_n170_ );
xor g053 ( new_n172_, N183, N189 );
xnor g054 ( new_n173_, N195, N201 );
xnor g055 ( new_n174_, new_n172_, new_n173_ );
xnor g056 ( new_n175_, new_n174_, N207 );
xnor g057 ( new_n176_, N159, N165 );
xnor g058 ( new_n177_, N171, N177 );
xnor g059 ( new_n178_, new_n176_, new_n177_ );
xnor g060 ( new_n179_, new_n178_, N130 );
xnor g061 ( N768, new_n175_, new_n179_ );
not g062 ( new_n181_, N201 );
not g063 ( new_n182_, N126 );
not g064 ( new_n183_, keyIn_0_5 );
nand g065 ( new_n184_, N17, N51 );
nor g066 ( new_n185_, new_n131_, new_n184_ );
xnor g067 ( new_n186_, new_n185_, keyIn_0_1 );
nor g068 ( new_n187_, new_n186_, new_n183_ );
nand g069 ( new_n188_, new_n186_, new_n183_ );
nand g070 ( new_n189_, new_n141_, N42 );
nand g071 ( new_n190_, new_n188_, new_n189_ );
nor g072 ( new_n191_, new_n190_, new_n187_ );
xnor g073 ( new_n192_, new_n191_, keyIn_0_8 );
not g074 ( new_n193_, new_n136_ );
nand g075 ( new_n194_, new_n193_, N51 );
nand g076 ( new_n195_, new_n194_, keyIn_0_0 );
not g077 ( new_n196_, keyIn_0_0 );
nand g078 ( new_n197_, new_n152_, new_n196_ );
nand g079 ( new_n198_, new_n195_, new_n197_ );
xnor g080 ( new_n199_, new_n198_, keyIn_0_4 );
nand g081 ( new_n200_, new_n199_, keyIn_0_7 );
not g082 ( new_n201_, keyIn_0_7 );
not g083 ( new_n202_, keyIn_0_4 );
nand g084 ( new_n203_, new_n198_, new_n202_ );
nand g085 ( new_n204_, N447, keyIn_0_4 );
nand g086 ( new_n205_, new_n204_, new_n203_ );
nand g087 ( new_n206_, new_n205_, new_n201_ );
nand g088 ( new_n207_, new_n200_, new_n206_ );
not g089 ( new_n208_, keyIn_0_6 );
nand g090 ( new_n209_, keyIn_0_3, N17 );
not g091 ( new_n210_, new_n209_ );
nand g092 ( new_n211_, new_n210_, N42 );
not g093 ( new_n212_, keyIn_0_3 );
nand g094 ( new_n213_, N17, N42 );
nand g095 ( new_n214_, new_n213_, new_n212_ );
nand g096 ( new_n215_, new_n211_, new_n214_ );
nand g097 ( new_n216_, new_n129_, new_n125_ );
xnor g098 ( new_n217_, new_n216_, keyIn_0_2 );
nand g099 ( new_n218_, new_n217_, new_n215_ );
nor g100 ( new_n219_, new_n218_, new_n208_ );
nand g101 ( new_n220_, new_n218_, new_n208_ );
nand g102 ( new_n221_, N59, N156 );
not g103 ( new_n222_, new_n221_ );
nand g104 ( new_n223_, new_n220_, new_n222_ );
nor g105 ( new_n224_, new_n223_, new_n219_ );
nand g106 ( new_n225_, new_n207_, new_n224_ );
xnor g107 ( new_n226_, new_n225_, keyIn_0_9 );
nor g108 ( new_n227_, new_n226_, new_n192_ );
nand g109 ( new_n228_, new_n227_, keyIn_0_10 );
not g110 ( new_n229_, keyIn_0_10 );
not g111 ( new_n230_, new_n192_ );
not g112 ( new_n231_, keyIn_0_9 );
xnor g113 ( new_n232_, new_n225_, new_n231_ );
nand g114 ( new_n233_, new_n232_, new_n230_ );
nand g115 ( new_n234_, new_n233_, new_n229_ );
nand g116 ( new_n235_, new_n228_, new_n234_ );
not g117 ( new_n236_, new_n235_ );
nor g118 ( new_n237_, new_n236_, new_n182_ );
not g119 ( new_n238_, N153 );
not g120 ( new_n239_, N1 );
nand g121 ( new_n240_, new_n207_, new_n221_ );
nor g122 ( new_n241_, new_n240_, new_n129_ );
nor g123 ( new_n242_, new_n241_, new_n239_ );
nor g124 ( new_n243_, new_n242_, new_n238_ );
nand g125 ( new_n244_, N29, N75 );
nor g126 ( new_n245_, new_n244_, new_n122_ );
nand g127 ( new_n246_, new_n207_, new_n245_ );
not g128 ( new_n247_, new_n246_ );
not g129 ( new_n248_, N55 );
nor g130 ( new_n249_, new_n248_, N268 );
nand g131 ( new_n250_, new_n247_, new_n249_ );
not g132 ( new_n251_, new_n250_ );
nor g133 ( new_n252_, new_n243_, new_n251_ );
not g134 ( new_n253_, new_n252_ );
nor g135 ( new_n254_, new_n237_, new_n253_ );
nand g136 ( new_n255_, new_n254_, new_n181_ );
not g137 ( new_n256_, new_n255_ );
not g138 ( new_n257_, new_n254_ );
nand g139 ( new_n258_, new_n257_, N201 );
not g140 ( new_n259_, new_n258_ );
nor g141 ( new_n260_, new_n259_, new_n256_ );
nand g142 ( new_n261_, new_n260_, N261 );
not g143 ( new_n262_, N219 );
nor g144 ( new_n263_, new_n260_, N261 );
nor g145 ( new_n264_, new_n263_, new_n262_ );
nand g146 ( new_n265_, new_n264_, new_n261_ );
not g147 ( new_n266_, N228 );
not g148 ( new_n267_, new_n260_ );
nor g149 ( new_n268_, new_n267_, new_n266_ );
nand g150 ( new_n269_, new_n259_, N237 );
nand g151 ( new_n270_, new_n257_, N246 );
not g152 ( new_n271_, N73 );
nand g153 ( new_n272_, N42, N72 );
nor g154 ( new_n273_, new_n272_, new_n271_ );
nand g155 ( new_n274_, new_n273_, new_n158_ );
nor g156 ( new_n275_, new_n154_, new_n274_ );
nand g157 ( new_n276_, new_n275_, N201 );
nand g158 ( new_n277_, N121, N210 );
nand g159 ( new_n278_, N255, N267 );
nand g160 ( new_n279_, new_n277_, new_n278_ );
not g161 ( new_n280_, new_n279_ );
nand g162 ( new_n281_, new_n276_, new_n280_ );
not g163 ( new_n282_, new_n281_ );
nand g164 ( new_n283_, new_n270_, new_n282_ );
not g165 ( new_n284_, new_n283_ );
nand g166 ( new_n285_, new_n269_, new_n284_ );
nor g167 ( new_n286_, new_n268_, new_n285_ );
nand g168 ( N850, new_n265_, new_n286_ );
not g169 ( new_n288_, keyIn_0_13 );
not g170 ( new_n289_, keyIn_0_11 );
nand g171 ( new_n290_, new_n235_, N111 );
nor g172 ( new_n291_, new_n290_, new_n289_ );
nand g173 ( new_n292_, new_n290_, new_n289_ );
not g174 ( new_n293_, new_n242_ );
nand g175 ( new_n294_, new_n293_, N143 );
nand g176 ( new_n295_, new_n292_, new_n294_ );
nor g177 ( new_n296_, new_n295_, new_n291_ );
nand g178 ( new_n297_, new_n296_, keyIn_0_12 );
not g179 ( new_n298_, new_n297_ );
not g180 ( new_n299_, keyIn_0_12 );
not g181 ( new_n300_, new_n291_ );
not g182 ( new_n301_, new_n295_ );
nand g183 ( new_n302_, new_n301_, new_n300_ );
nand g184 ( new_n303_, new_n302_, new_n299_ );
nand g185 ( new_n304_, new_n303_, new_n250_ );
nor g186 ( new_n305_, new_n304_, new_n298_ );
nand g187 ( new_n306_, new_n305_, new_n288_ );
nor g188 ( new_n307_, new_n296_, keyIn_0_12 );
nor g189 ( new_n308_, new_n307_, new_n251_ );
nand g190 ( new_n309_, new_n308_, new_n297_ );
nand g191 ( new_n310_, new_n309_, keyIn_0_13 );
nand g192 ( new_n311_, new_n306_, new_n310_ );
nand g193 ( new_n312_, new_n311_, N183 );
xnor g194 ( new_n313_, new_n312_, keyIn_0_14 );
not g195 ( new_n314_, keyIn_0_15 );
nor g196 ( new_n315_, new_n311_, N183 );
nand g197 ( new_n316_, new_n315_, new_n314_ );
not g198 ( new_n317_, N183 );
xnor g199 ( new_n318_, new_n309_, new_n288_ );
nand g200 ( new_n319_, new_n318_, new_n317_ );
nand g201 ( new_n320_, new_n319_, keyIn_0_15 );
nand g202 ( new_n321_, new_n320_, new_n316_ );
nand g203 ( new_n322_, new_n313_, new_n321_ );
nand g204 ( new_n323_, new_n235_, N121 );
not g205 ( new_n324_, N149 );
nor g206 ( new_n325_, new_n242_, new_n324_ );
nor g207 ( new_n326_, new_n325_, new_n251_ );
nand g208 ( new_n327_, new_n323_, new_n326_ );
nor g209 ( new_n328_, new_n327_, N195 );
xor g210 ( new_n329_, new_n328_, keyIn_0_16 );
nand g211 ( new_n330_, new_n329_, new_n259_ );
nand g212 ( new_n331_, new_n327_, N195 );
nand g213 ( new_n332_, new_n330_, new_n331_ );
nand g214 ( new_n333_, new_n235_, N116 );
not g215 ( new_n334_, N146 );
nor g216 ( new_n335_, new_n242_, new_n334_ );
nor g217 ( new_n336_, new_n335_, new_n251_ );
nand g218 ( new_n337_, new_n333_, new_n336_ );
nor g219 ( new_n338_, new_n337_, N189 );
not g220 ( new_n339_, new_n338_ );
nand g221 ( new_n340_, new_n332_, new_n339_ );
nand g222 ( new_n341_, new_n255_, N261 );
nor g223 ( new_n342_, new_n341_, new_n338_ );
nand g224 ( new_n343_, new_n342_, new_n329_ );
nor g225 ( new_n344_, new_n343_, keyIn_0_18 );
nand g226 ( new_n345_, new_n337_, N189 );
nand g227 ( new_n346_, new_n343_, keyIn_0_18 );
nand g228 ( new_n347_, new_n346_, new_n345_ );
nor g229 ( new_n348_, new_n347_, new_n344_ );
nand g230 ( new_n349_, new_n348_, new_n340_ );
not g231 ( new_n350_, new_n349_ );
nand g232 ( new_n351_, new_n322_, new_n350_ );
nor g233 ( new_n352_, new_n322_, new_n350_ );
nor g234 ( new_n353_, new_n352_, new_n262_ );
nand g235 ( new_n354_, new_n353_, new_n351_ );
not g236 ( new_n355_, N237 );
xnor g237 ( new_n356_, new_n313_, keyIn_0_17 );
nor g238 ( new_n357_, new_n356_, new_n355_ );
not g239 ( new_n358_, new_n322_ );
nand g240 ( new_n359_, new_n358_, N228 );
not g241 ( new_n360_, N246 );
nor g242 ( new_n361_, new_n318_, new_n360_ );
nand g243 ( new_n362_, new_n275_, N183 );
nand g244 ( new_n363_, N106, N210 );
nand g245 ( new_n364_, new_n362_, new_n363_ );
nor g246 ( new_n365_, new_n361_, new_n364_ );
nand g247 ( new_n366_, new_n359_, new_n365_ );
nor g248 ( new_n367_, new_n357_, new_n366_ );
nand g249 ( N863, new_n367_, new_n354_ );
nand g250 ( new_n369_, new_n341_, new_n258_ );
nand g251 ( new_n370_, new_n329_, new_n369_ );
nand g252 ( new_n371_, new_n370_, new_n331_ );
not g253 ( new_n372_, new_n345_ );
nor g254 ( new_n373_, new_n372_, new_n338_ );
nand g255 ( new_n374_, new_n371_, new_n373_ );
nor g256 ( new_n375_, new_n371_, new_n373_ );
nor g257 ( new_n376_, new_n375_, new_n262_ );
nand g258 ( new_n377_, new_n376_, new_n374_ );
not g259 ( new_n378_, new_n373_ );
nor g260 ( new_n379_, new_n378_, new_n266_ );
nand g261 ( new_n380_, new_n372_, N237 );
nand g262 ( new_n381_, new_n337_, N246 );
nand g263 ( new_n382_, new_n275_, N189 );
nand g264 ( new_n383_, N111, N210 );
nand g265 ( new_n384_, N255, N259 );
nand g266 ( new_n385_, new_n383_, new_n384_ );
not g267 ( new_n386_, new_n385_ );
nand g268 ( new_n387_, new_n382_, new_n386_ );
not g269 ( new_n388_, new_n387_ );
nand g270 ( new_n389_, new_n381_, new_n388_ );
not g271 ( new_n390_, new_n389_ );
nand g272 ( new_n391_, new_n380_, new_n390_ );
nor g273 ( new_n392_, new_n379_, new_n391_ );
nand g274 ( N864, new_n377_, new_n392_ );
nand g275 ( new_n394_, new_n329_, new_n331_ );
not g276 ( new_n395_, new_n394_ );
nand g277 ( new_n396_, new_n395_, new_n369_ );
not g278 ( new_n397_, new_n369_ );
nand g279 ( new_n398_, new_n394_, new_n397_ );
nand g280 ( new_n399_, new_n398_, N219 );
not g281 ( new_n400_, new_n399_ );
nand g282 ( new_n401_, new_n400_, new_n396_ );
nor g283 ( new_n402_, new_n394_, new_n266_ );
not g284 ( new_n403_, new_n331_ );
nand g285 ( new_n404_, new_n403_, N237 );
nand g286 ( new_n405_, new_n327_, N246 );
nand g287 ( new_n406_, new_n275_, N195 );
nand g288 ( new_n407_, N116, N210 );
nand g289 ( new_n408_, N255, N260 );
nand g290 ( new_n409_, new_n407_, new_n408_ );
not g291 ( new_n410_, new_n409_ );
nand g292 ( new_n411_, new_n406_, new_n410_ );
not g293 ( new_n412_, new_n411_ );
nand g294 ( new_n413_, new_n405_, new_n412_ );
not g295 ( new_n414_, new_n413_ );
nand g296 ( new_n415_, new_n404_, new_n414_ );
nor g297 ( new_n416_, new_n402_, new_n415_ );
nand g298 ( N865, new_n401_, new_n416_ );
not g299 ( new_n418_, keyIn_0_21 );
not g300 ( new_n419_, keyIn_0_17 );
nand g301 ( new_n420_, new_n313_, new_n419_ );
not g302 ( new_n421_, keyIn_0_14 );
xnor g303 ( new_n422_, new_n312_, new_n421_ );
nand g304 ( new_n423_, new_n422_, keyIn_0_17 );
nand g305 ( new_n424_, new_n420_, new_n423_ );
nor g306 ( new_n425_, new_n424_, new_n418_ );
not g307 ( new_n426_, keyIn_0_22 );
nand g308 ( new_n427_, new_n321_, new_n349_ );
xnor g309 ( new_n428_, new_n427_, new_n426_ );
nand g310 ( new_n429_, new_n424_, new_n418_ );
nand g311 ( new_n430_, new_n428_, new_n429_ );
nor g312 ( new_n431_, new_n430_, new_n425_ );
xnor g313 ( new_n432_, new_n431_, keyIn_0_23 );
nand g314 ( new_n433_, new_n235_, N106 );
nor g315 ( new_n434_, new_n240_, new_n248_ );
not g316 ( new_n435_, new_n434_ );
nor g317 ( new_n436_, new_n435_, new_n238_ );
nor g318 ( new_n437_, new_n129_, N268 );
nand g319 ( new_n438_, new_n247_, new_n437_ );
nand g320 ( new_n439_, N138, N152 );
nand g321 ( new_n440_, new_n438_, new_n439_ );
nor g322 ( new_n441_, new_n436_, new_n440_ );
nand g323 ( new_n442_, new_n433_, new_n441_ );
nor g324 ( new_n443_, new_n442_, N177 );
nor g325 ( new_n444_, new_n432_, new_n443_ );
nand g326 ( new_n445_, new_n442_, N177 );
not g327 ( new_n446_, new_n445_ );
nor g328 ( new_n447_, new_n444_, new_n446_ );
not g329 ( new_n448_, new_n447_ );
not g330 ( new_n449_, N171 );
nand g331 ( new_n450_, new_n235_, N101 );
nor g332 ( new_n451_, new_n435_, new_n324_ );
nand g333 ( new_n452_, N17, N138 );
nand g334 ( new_n453_, new_n438_, new_n452_ );
nor g335 ( new_n454_, new_n451_, new_n453_ );
nand g336 ( new_n455_, new_n450_, new_n454_ );
not g337 ( new_n456_, new_n455_ );
nand g338 ( new_n457_, new_n456_, new_n449_ );
nand g339 ( new_n458_, new_n448_, new_n457_ );
nand g340 ( new_n459_, new_n455_, N171 );
nand g341 ( new_n460_, new_n458_, new_n459_ );
not g342 ( new_n461_, N165 );
nand g343 ( new_n462_, new_n235_, N96 );
nor g344 ( new_n463_, new_n435_, new_n334_ );
nand g345 ( new_n464_, N51, N138 );
nand g346 ( new_n465_, new_n438_, new_n464_ );
nor g347 ( new_n466_, new_n463_, new_n465_ );
nand g348 ( new_n467_, new_n462_, new_n466_ );
not g349 ( new_n468_, new_n467_ );
nand g350 ( new_n469_, new_n468_, new_n461_ );
nand g351 ( new_n470_, new_n460_, new_n469_ );
nand g352 ( new_n471_, new_n467_, N165 );
nand g353 ( new_n472_, new_n470_, new_n471_ );
not g354 ( new_n473_, N159 );
nand g355 ( new_n474_, new_n235_, N91 );
nand g356 ( new_n475_, new_n434_, N143 );
not g357 ( new_n476_, new_n475_ );
nand g358 ( new_n477_, N8, N138 );
nand g359 ( new_n478_, new_n438_, new_n477_ );
nor g360 ( new_n479_, new_n476_, new_n478_ );
nand g361 ( new_n480_, new_n474_, new_n479_ );
not g362 ( new_n481_, new_n480_ );
nand g363 ( new_n482_, new_n481_, new_n473_ );
nand g364 ( new_n483_, new_n472_, new_n482_ );
nand g365 ( new_n484_, new_n480_, N159 );
nand g366 ( N866, new_n483_, new_n484_ );
not g367 ( new_n486_, keyIn_0_30 );
not g368 ( new_n487_, keyIn_0_28 );
not g369 ( new_n488_, keyIn_0_24 );
not g370 ( new_n489_, new_n425_ );
xnor g371 ( new_n490_, new_n427_, keyIn_0_22 );
nor g372 ( new_n491_, new_n356_, keyIn_0_21 );
nor g373 ( new_n492_, new_n491_, new_n490_ );
nand g374 ( new_n493_, new_n492_, new_n489_ );
nand g375 ( new_n494_, new_n493_, keyIn_0_23 );
not g376 ( new_n495_, keyIn_0_23 );
nand g377 ( new_n496_, new_n431_, new_n495_ );
nand g378 ( new_n497_, new_n494_, new_n496_ );
nor g379 ( new_n498_, new_n446_, new_n443_ );
nor g380 ( new_n499_, new_n497_, new_n498_ );
nand g381 ( new_n500_, new_n499_, new_n488_ );
not g382 ( new_n501_, new_n498_ );
nand g383 ( new_n502_, new_n432_, new_n501_ );
nand g384 ( new_n503_, new_n502_, keyIn_0_24 );
nand g385 ( new_n504_, new_n500_, new_n503_ );
not g386 ( new_n505_, keyIn_0_25 );
nand g387 ( new_n506_, new_n497_, new_n498_ );
nand g388 ( new_n507_, new_n506_, new_n505_ );
nor g389 ( new_n508_, new_n432_, new_n501_ );
nand g390 ( new_n509_, new_n508_, keyIn_0_25 );
nand g391 ( new_n510_, new_n509_, new_n507_ );
nand g392 ( new_n511_, new_n510_, new_n504_ );
nor g393 ( new_n512_, new_n511_, keyIn_0_26 );
not g394 ( new_n513_, new_n512_ );
nand g395 ( new_n514_, new_n511_, keyIn_0_26 );
nand g396 ( new_n515_, new_n514_, N219 );
not g397 ( new_n516_, new_n515_ );
nand g398 ( new_n517_, new_n516_, new_n513_ );
nor g399 ( new_n518_, new_n517_, keyIn_0_27 );
not g400 ( new_n519_, new_n518_ );
not g401 ( new_n520_, keyIn_0_27 );
nor g402 ( new_n521_, new_n515_, new_n512_ );
nor g403 ( new_n522_, new_n521_, new_n520_ );
nand g404 ( new_n523_, N101, N210 );
not g405 ( new_n524_, new_n523_ );
nor g406 ( new_n525_, new_n522_, new_n524_ );
nand g407 ( new_n526_, new_n519_, new_n525_ );
nor g408 ( new_n527_, new_n526_, new_n487_ );
not g409 ( new_n528_, new_n527_ );
nand g410 ( new_n529_, new_n517_, keyIn_0_27 );
nand g411 ( new_n530_, new_n529_, new_n523_ );
nor g412 ( new_n531_, new_n530_, new_n518_ );
nor g413 ( new_n532_, new_n531_, keyIn_0_28 );
nor g414 ( new_n533_, new_n501_, new_n266_ );
not g415 ( new_n534_, new_n533_ );
nor g416 ( new_n535_, new_n534_, keyIn_0_20 );
nand g417 ( new_n536_, new_n534_, keyIn_0_20 );
nor g418 ( new_n537_, new_n445_, new_n355_ );
nand g419 ( new_n538_, new_n442_, N246 );
nand g420 ( new_n539_, new_n275_, N177 );
nand g421 ( new_n540_, new_n538_, new_n539_ );
nor g422 ( new_n541_, new_n537_, new_n540_ );
nand g423 ( new_n542_, new_n536_, new_n541_ );
nor g424 ( new_n543_, new_n542_, new_n535_ );
not g425 ( new_n544_, new_n543_ );
nor g426 ( new_n545_, new_n532_, new_n544_ );
nand g427 ( new_n546_, new_n545_, new_n528_ );
nand g428 ( new_n547_, new_n546_, keyIn_0_29 );
not g429 ( new_n548_, keyIn_0_29 );
nand g430 ( new_n549_, new_n526_, new_n487_ );
nand g431 ( new_n550_, new_n549_, new_n543_ );
nor g432 ( new_n551_, new_n550_, new_n527_ );
nand g433 ( new_n552_, new_n551_, new_n548_ );
nand g434 ( new_n553_, new_n547_, new_n552_ );
nand g435 ( new_n554_, new_n553_, new_n486_ );
xnor g436 ( new_n555_, new_n551_, keyIn_0_29 );
nand g437 ( new_n556_, new_n555_, keyIn_0_30 );
nand g438 ( new_n557_, new_n556_, new_n554_ );
nand g439 ( new_n558_, new_n557_, keyIn_0_31 );
not g440 ( new_n559_, keyIn_0_31 );
xnor g441 ( new_n560_, new_n553_, keyIn_0_30 );
nand g442 ( new_n561_, new_n560_, new_n559_ );
nand g443 ( N874, new_n561_, new_n558_ );
nand g444 ( new_n563_, new_n482_, new_n484_ );
not g445 ( new_n564_, new_n563_ );
nand g446 ( new_n565_, new_n472_, new_n564_ );
nor g447 ( new_n566_, new_n472_, new_n564_ );
nor g448 ( new_n567_, new_n566_, new_n262_ );
nand g449 ( new_n568_, new_n567_, new_n565_ );
nor g450 ( new_n569_, new_n563_, new_n266_ );
not g451 ( new_n570_, new_n484_ );
nand g452 ( new_n571_, new_n570_, N237 );
nand g453 ( new_n572_, new_n480_, N246 );
nand g454 ( new_n573_, new_n275_, N159 );
nand g455 ( new_n574_, N210, N268 );
nand g456 ( new_n575_, new_n573_, new_n574_ );
not g457 ( new_n576_, new_n575_ );
nand g458 ( new_n577_, new_n572_, new_n576_ );
not g459 ( new_n578_, new_n577_ );
nand g460 ( new_n579_, new_n571_, new_n578_ );
nor g461 ( new_n580_, new_n569_, new_n579_ );
nand g462 ( N878, new_n568_, new_n580_ );
nand g463 ( new_n582_, new_n469_, new_n471_ );
not g464 ( new_n583_, new_n582_ );
nand g465 ( new_n584_, new_n460_, new_n583_ );
nor g466 ( new_n585_, new_n460_, new_n583_ );
nor g467 ( new_n586_, new_n585_, new_n262_ );
nand g468 ( new_n587_, new_n586_, new_n584_ );
nor g469 ( new_n588_, new_n582_, new_n266_ );
not g470 ( new_n589_, new_n471_ );
nand g471 ( new_n590_, new_n589_, N237 );
nand g472 ( new_n591_, new_n467_, N246 );
nand g473 ( new_n592_, new_n275_, N165 );
nand g474 ( new_n593_, N91, N210 );
nand g475 ( new_n594_, new_n592_, new_n593_ );
not g476 ( new_n595_, new_n594_ );
nand g477 ( new_n596_, new_n591_, new_n595_ );
not g478 ( new_n597_, new_n596_ );
nand g479 ( new_n598_, new_n590_, new_n597_ );
nor g480 ( new_n599_, new_n588_, new_n598_ );
nand g481 ( N879, new_n587_, new_n599_ );
nand g482 ( new_n601_, new_n457_, new_n459_ );
nand g483 ( new_n602_, new_n447_, new_n601_ );
not g484 ( new_n603_, new_n601_ );
nand g485 ( new_n604_, new_n448_, new_n603_ );
nand g486 ( new_n605_, new_n604_, N219 );
not g487 ( new_n606_, new_n605_ );
nand g488 ( new_n607_, new_n606_, new_n602_ );
not g489 ( new_n608_, keyIn_0_19 );
nor g490 ( new_n609_, new_n459_, new_n355_ );
nand g491 ( new_n610_, new_n609_, new_n608_ );
nand g492 ( new_n611_, new_n455_, N246 );
nand g493 ( new_n612_, new_n275_, N171 );
nand g494 ( new_n613_, N96, N210 );
nand g495 ( new_n614_, new_n612_, new_n613_ );
not g496 ( new_n615_, new_n614_ );
nand g497 ( new_n616_, new_n611_, new_n615_ );
not g498 ( new_n617_, new_n616_ );
nand g499 ( new_n618_, new_n610_, new_n617_ );
not g500 ( new_n619_, new_n609_ );
nand g501 ( new_n620_, new_n619_, keyIn_0_19 );
nand g502 ( new_n621_, new_n603_, N228 );
nand g503 ( new_n622_, new_n621_, new_n620_ );
nor g504 ( new_n623_, new_n622_, new_n618_ );
nand g505 ( N880, new_n607_, new_n623_ );
endmodule