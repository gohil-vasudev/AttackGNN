module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n1668_, new_n1359_, new_n595_, new_n1233_, new_n2051_, new_n1839_, new_n445_, new_n1009_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n1743_, new_n501_, new_n1157_, new_n2086_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1988_, new_n1433_, new_n1517_, new_n1575_, new_n1472_, new_n1048_, new_n1785_, new_n885_, new_n439_, new_n1532_, new_n1808_, new_n390_, new_n1910_, new_n743_, new_n1962_, new_n1327_, new_n1535_, new_n2041_, new_n1922_, new_n566_, new_n641_, new_n1849_, new_n386_, new_n767_, new_n389_, new_n514_, new_n1865_, new_n1351_, new_n556_, new_n636_, new_n1899_, new_n691_, new_n1024_, new_n670_, new_n456_, new_n1125_, new_n1590_, new_n2095_, new_n1881_, new_n911_, new_n679_, new_n937_, new_n667_, new_n2099_, new_n1879_, new_n1237_, new_n2054_, new_n2026_, new_n1837_, new_n1568_, new_n728_, new_n1479_, new_n1071_, new_n1294_, new_n894_, new_n853_, new_n695_, new_n660_, new_n2038_, new_n1311_, new_n526_, new_n908_, new_n1886_, new_n2023_, new_n552_, new_n678_, new_n1662_, new_n706_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n2063_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n2033_, new_n1163_, new_n786_, new_n2045_, new_n1769_, new_n1103_, new_n1188_, new_n1415_, new_n1390_, new_n721_, new_n504_, new_n1414_, new_n742_, new_n892_, new_n1368_, new_n472_, new_n873_, new_n1919_, new_n1985_, new_n1768_, new_n1167_, new_n1530_, new_n1300_, new_n2070_, new_n1898_, new_n1490_, new_n774_, new_n1777_, new_n792_, new_n1620_, new_n953_, new_n1786_, new_n1946_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n1580_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n1973_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n1851_, new_n1447_, new_n635_, new_n1774_, new_n685_, new_n648_, new_n903_, new_n1595_, new_n1803_, new_n983_, new_n822_, new_n1406_, new_n1990_, new_n1082_, new_n1760_, new_n1018_, new_n1884_, new_n1864_, new_n606_, new_n796_, new_n1054_, new_n655_, new_n1288_, new_n630_, new_n1717_, new_n385_, new_n1670_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n1979_, new_n1196_, new_n1366_, new_n1984_, new_n511_, new_n1714_, new_n2034_, new_n1640_, new_n1285_, new_n1031_, new_n1733_, new_n1216_, new_n1632_, new_n1889_, new_n1987_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1911_, new_n1005_, new_n999_, new_n1647_, new_n1816_, new_n1713_, new_n960_, new_n1377_, new_n1522_, new_n549_, new_n491_, new_n676_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n2072_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n1753_, new_n1678_, new_n568_, new_n420_, new_n876_, new_n1894_, new_n1900_, new_n1950_, new_n1936_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n2032_, new_n1463_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1424_, new_n1062_, new_n680_, new_n981_, new_n506_, new_n872_, new_n1527_, new_n1275_, new_n1277_, new_n1800_, new_n1198_, new_n1428_, new_n1440_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n2012_, new_n483_, new_n1004_, new_n1152_, new_n1558_, new_n394_, new_n935_, new_n1972_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1735_, new_n1113_, new_n785_, new_n1501_, new_n441_, new_n477_, new_n664_, new_n1752_, new_n600_, new_n1737_, new_n1930_, new_n1041_, new_n1657_, new_n1989_, new_n1797_, new_n426_, new_n1036_, new_n1562_, new_n1939_, new_n1953_, new_n398_, new_n1576_, new_n1718_, new_n1333_, new_n395_, new_n1132_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n1740_, new_n1395_, new_n473_, new_n1624_, new_n1147_, new_n1682_, new_n1795_, new_n1373_, new_n1229_, new_n1827_, new_n1422_, new_n1523_, new_n1698_, new_n1468_, new_n1679_, new_n969_, new_n835_, new_n1234_, new_n1360_, new_n378_, new_n1574_, new_n1614_, new_n621_, new_n1423_, new_n1637_, new_n1732_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1798_, new_n1321_, new_n1690_, new_n1209_, new_n1709_, new_n347_, new_n2084_, new_n2100_, new_n659_, new_n700_, new_n1419_, new_n921_, new_n346_, new_n396_, new_n1954_, new_n1315_, new_n1003_, new_n696_, new_n1868_, new_n1039_, new_n1507_, new_n1439_, new_n1658_, new_n1952_, new_n1671_, new_n1239_, new_n1365_, new_n528_, new_n952_, new_n1870_, new_n1158_, new_n1667_, new_n729_, new_n1111_, new_n1413_, new_n1218_, new_n1385_, new_n1346_, new_n1201_, new_n559_, new_n1282_, new_n1630_, new_n762_, new_n1349_, new_n1193_, new_n1547_, new_n1780_, new_n1994_, new_n1437_, new_n1598_, new_n1187_, new_n1205_, new_n1966_, new_n1154_, new_n1253_, new_n1546_, new_n1453_, new_n1256_, new_n1850_, new_n628_, new_n1513_, new_n409_, new_n1090_, new_n1669_, new_n1489_, new_n553_, new_n745_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n834_, new_n1991_, new_n1573_, new_n1781_, new_n1738_, new_n369_, new_n1693_, new_n1171_, new_n867_, new_n954_, new_n1591_, new_n1626_, new_n1032_, new_n1545_, new_n901_, new_n1757_, new_n688_, new_n1255_, new_n1704_, new_n985_, new_n2074_, new_n1995_, new_n851_, new_n1518_, new_n932_, new_n878_, new_n1981_, new_n543_, new_n1943_, new_n1975_, new_n886_, new_n371_, new_n1712_, new_n509_, new_n1761_, new_n2058_, new_n2075_, new_n661_, new_n797_, new_n1358_, new_n724_, new_n1070_, new_n1686_, new_n1416_, new_n1109_, new_n1496_, new_n672_, new_n1269_, new_n616_, new_n1653_, new_n529_, new_n884_, new_n914_, new_n1875_, new_n938_, new_n362_, new_n1600_, new_n1592_, new_n809_, new_n1631_, new_n1142_, new_n1623_, new_n604_, new_n1104_, new_n1703_, new_n1771_, new_n1511_, new_n571_, new_n1859_, new_n1504_, new_n758_, new_n1802_, new_n460_, new_n1267_, new_n2015_, new_n1794_, new_n1705_, new_n2090_, new_n1466_, new_n1707_, new_n1716_, new_n1516_, new_n1299_, new_n380_, new_n1477_, new_n1079_, new_n861_, new_n1564_, new_n1656_, new_n1252_, new_n1993_, new_n1804_, new_n1553_, new_n931_, new_n575_, new_n1493_, new_n562_, new_n1593_, new_n944_, new_n1929_, new_n1638_, new_n1542_, new_n1064_, new_n1949_, new_n1065_, new_n1118_, new_n1645_, new_n493_, new_n547_, new_n1480_, new_n1934_, new_n1745_, new_n1860_, new_n379_, new_n1825_, new_n963_, new_n586_, new_n1481_, new_n1325_, new_n993_, new_n1625_, new_n1357_, new_n1191_, new_n1931_, new_n824_, new_n1628_, new_n717_, new_n1455_, new_n403_, new_n868_, new_n1242_, new_n475_, new_n858_, new_n1612_, new_n1384_, new_n1343_, new_n936_, new_n1459_, new_n1434_, new_n1438_, new_n1016_, new_n411_, new_n673_, new_n1766_, new_n1904_, new_n1144_, new_n2025_, new_n1465_, new_n2082_, new_n666_, new_n1290_, new_n2065_, new_n407_, new_n1897_, new_n1833_, new_n1519_, new_n1407_, new_n1692_, new_n1726_, new_n879_, new_n1417_, new_n1700_, new_n736_, new_n513_, new_n1903_, new_n558_, new_n382_, new_n1370_, new_n718_, new_n2093_, new_n1310_, new_n2042_, new_n1710_, new_n1398_, new_n1126_, new_n2047_, new_n546_, new_n612_, new_n1015_, new_n919_, new_n755_, new_n2017_, new_n1040_, new_n1635_, new_n1509_, new_n1559_, new_n1789_, new_n544_, new_n615_, new_n722_, new_n1941_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n2068_, new_n2066_, new_n499_, new_n533_, new_n1130_, new_n2064_, new_n795_, new_n459_, new_n1441_, new_n1122_, new_n1728_, new_n1185_, new_n1240_, new_n2031_, new_n1510_, new_n354_, new_n1174_, new_n968_, new_n2001_, new_n2055_, new_n1655_, new_n1464_, new_n613_, new_n1508_, new_n1195_, new_n417_, new_n658_, new_n837_, new_n591_, new_n801_, new_n2039_, new_n1458_, new_n2091_, new_n631_, new_n453_, new_n1723_, new_n1818_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1521_, new_n1334_, new_n2044_, new_n531_, new_n1826_, new_n1675_, new_n593_, new_n1543_, new_n974_, new_n1907_, new_n1565_, new_n1248_, new_n1812_, new_n751_, new_n1978_, new_n1038_, new_n372_, new_n1758_, new_n852_, new_n1454_, new_n1474_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n1430_, new_n470_, new_n769_, new_n1660_, new_n433_, new_n871_, new_n2096_, new_n1956_, new_n1450_, new_n992_, new_n1098_, new_n1729_, new_n2069_, new_n732_, new_n1832_, new_n689_, new_n933_, new_n584_, new_n815_, new_n1608_, new_n1492_, new_n1619_, new_n1052_, new_n1425_, new_n1980_, new_n857_, new_n1828_, new_n1379_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n1853_, new_n512_, new_n1471_, new_n1673_, new_n1220_, new_n989_, new_n1741_, new_n1117_, new_n1421_, new_n644_, new_n1594_, new_n836_, new_n1856_, new_n1116_, new_n1684_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n913_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n1427_, new_n818_, new_n881_, new_n1815_, new_n1268_, new_n2052_, new_n1376_, new_n1381_, new_n1876_, new_n1566_, new_n2092_, new_n1534_, new_n684_, new_n640_, new_n1274_, new_n1893_, new_n1665_, new_n754_, new_n1787_, new_n653_, new_n1659_, new_n905_, new_n1258_, new_n1539_, new_n1643_, new_n375_, new_n1958_, new_n962_, new_n1841_, new_n760_, new_n627_, new_n1391_, new_n1724_, new_n1436_, new_n1986_, new_n567_, new_n1353_, new_n1033_, new_n576_, new_n831_, new_n791_, new_n2050_, new_n1153_, new_n1339_, new_n1784_, new_n1970_, new_n984_, new_n780_, new_n1183_, new_n643_, new_n1316_, new_n1194_, new_n1338_, new_n1460_, new_n1878_, new_n1230_, new_n1602_, new_n1027_, new_n610_, new_n1369_, new_n1694_, new_n843_, new_n703_, new_n698_, new_n1639_, new_n1165_, new_n1401_, new_n1259_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n1942_, new_n709_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1928_, new_n1066_, new_n1861_, new_n434_, new_n2021_, new_n422_, new_n1944_, new_n581_, new_n1664_, new_n686_, new_n934_, new_n1567_, new_n1651_, new_n770_, new_n1389_, new_n1400_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n1597_, new_n356_, new_n647_, new_n889_, new_n536_, new_n2083_, new_n1616_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n1806_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n1405_, new_n1249_, new_n1354_, new_n955_, new_n1895_, new_n847_, new_n888_, new_n1505_, new_n1340_, new_n798_, new_n1180_, new_n1926_, new_n1969_, new_n1948_, new_n817_, new_n720_, new_n1801_, new_n753_, new_n620_, new_n368_, new_n1361_, new_n941_, new_n1410_, new_n738_, new_n2073_, new_n827_, new_n1356_, new_n1363_, new_n1747_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n1211_, new_n1412_, new_n1207_, new_n1176_, new_n1374_, new_n1799_, new_n601_, new_n842_, new_n1552_, new_n1057_, new_n1644_, new_n1677_, new_n682_, new_n1075_, new_n1790_, new_n812_, new_n2030_, new_n1563_, new_n821_, new_n1937_, new_n542_, new_n548_, new_n669_, new_n1397_, new_n1402_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n1603_, new_n1971_, new_n451_, new_n489_, new_n804_, new_n1342_, new_n424_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n413_, new_n1906_, new_n1544_, new_n1382_, new_n1896_, new_n442_, new_n677_, new_n1843_, new_n1487_, new_n1646_, new_n642_, new_n1418_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n1814_, new_n1871_, new_n761_, new_n2027_, new_n735_, new_n840_, new_n1283_, new_n1913_, new_n1873_, new_n898_, new_n1734_, new_n799_, new_n1304_, new_n1537_, new_n946_, new_n1764_, new_n1834_, new_n344_, new_n1977_, new_n1108_, new_n1901_, new_n1469_, new_n862_, new_n1749_, new_n1606_, new_n1838_, new_n427_, new_n532_, new_n1739_, new_n393_, new_n1617_, new_n418_, new_n746_, new_n1221_, new_n1585_, new_n1587_, new_n1264_, new_n1319_, new_n626_, new_n1680_, new_n1473_, new_n959_, new_n990_, new_n1629_, new_n2005_, new_n716_, new_n701_, new_n1238_, new_n2062_, new_n1676_, new_n1058_, new_n2037_, new_n1880_, new_n1162_, new_n1730_, new_n2018_, new_n2003_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n1996_, new_n1696_, new_n414_, new_n2028_, new_n1968_, new_n1101_, new_n1250_, new_n2011_, new_n1681_, new_n1482_, new_n1050_, new_n554_, new_n1151_, new_n844_, new_n1302_, new_n2094_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n1083_, new_n759_, new_n1297_, new_n1959_, new_n829_, new_n1257_, new_n1306_, new_n1720_, new_n988_, new_n1858_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n1486_, new_n361_, new_n764_, new_n906_, new_n683_, new_n2081_, new_n1409_, new_n2007_, new_n1429_, new_n1955_, new_n463_, new_n1683_, new_n1372_, new_n510_, new_n966_, new_n1685_, new_n1721_, new_n351_, new_n1877_, new_n1184_, new_n1960_, new_n1292_, new_n1426_, new_n2036_, new_n609_, new_n517_, new_n2077_, new_n1759_, new_n961_, new_n530_, new_n890_, new_n1992_, new_n1006_, new_n1836_, new_n622_, new_n1706_, new_n2006_, new_n702_, new_n2014_, new_n833_, new_n1560_, new_n1701_, new_n1905_, new_n811_, new_n1445_, new_n1371_, new_n443_, new_n1086_, new_n1902_, new_n956_, new_n763_, new_n1622_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n1618_, new_n1652_, new_n1847_, new_n2057_, new_n1170_, new_n845_, new_n768_, new_n1691_, new_n773_, new_n1452_, new_n1051_, new_n899_, new_n1053_, new_n1540_, new_n1611_, new_n1823_, new_n1708_, new_n492_, new_n1200_, new_n1533_, new_n650_, new_n750_, new_n1754_, new_n1750_, new_n1767_, new_n887_, new_n355_, new_n926_, new_n432_, new_n925_, new_n2060_, new_n875_, new_n2040_, new_n1226_, new_n1940_, new_n778_, new_n452_, new_n1727_, new_n381_, new_n1483_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n820_, new_n1386_, new_n771_, new_n979_, new_n1819_, new_n508_, new_n1435_, new_n1844_, new_n714_, new_n1748_, new_n1280_, new_n1007_, new_n1613_, new_n1241_, new_n882_, new_n1145_, new_n1557_, new_n929_, new_n1159_, new_n1584_, new_n1337_, new_n1782_, new_n1348_, new_n917_, new_n2071_, new_n1555_, new_n1636_, new_n1322_, new_n1751_, new_n1133_, new_n1822_, new_n1887_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n2019_, new_n541_, new_n447_, new_n1967_, new_n1388_, new_n1550_, new_n790_, new_n1081_, new_n587_, new_n1247_, new_n1411_, new_n465_, new_n783_, new_n1380_, new_n2016_, new_n2000_, new_n739_, new_n996_, new_n2080_, new_n1601_, new_n1318_, new_n2088_, new_n846_, new_n915_, new_n488_, new_n524_, new_n349_, new_n848_, new_n1921_, new_n1725_, new_n1245_, new_n1772_, new_n663_, new_n1499_, new_n1497_, new_n579_, new_n1791_, new_n2035_, new_n1375_, new_n1908_, new_n1711_, new_n1254_, new_n1689_, new_n438_, new_n1344_, new_n1857_, new_n939_, new_n1393_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n1514_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n1526_, new_n397_, new_n1446_, new_n975_, new_n1199_, new_n399_, new_n1581_, new_n596_, new_n945_, new_n870_, new_n805_, new_n1420_, new_n1882_, new_n1115_, new_n1846_, new_n1403_, new_n1866_, new_n1383_, new_n1231_, new_n948_, new_n1520_, new_n1055_, new_n2043_, new_n1431_, new_n838_, new_n1609_, new_n923_, new_n1755_, new_n1674_, new_n469_, new_n437_, new_n1085_, new_n1633_, new_n1607_, new_n359_, new_n794_, new_n2098_, new_n1924_, new_n457_, new_n1852_, new_n1301_, new_n1999_, new_n1128_, new_n1582_, new_n2056_, new_n1002_, new_n2009_, new_n1169_, new_n1702_, new_n1909_, new_n1810_, new_n448_, new_n1932_, new_n384_, new_n900_, new_n1722_, new_n1824_, new_n1329_, new_n1161_, new_n1788_, new_n1648_, new_n1914_, new_n924_, new_n775_, new_n1867_, new_n454_, new_n1034_, new_n1872_, new_n1124_, new_n1957_, new_n1663_, new_n1000_, new_n1947_, new_n633_, new_n784_, new_n1273_, new_n1396_, new_n1491_, new_n1554_, new_n1923_, new_n2013_, new_n860_, new_n494_, new_n1160_, new_n1166_, new_n1536_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n1920_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n1272_, new_n693_, new_n1287_, new_n1485_, new_n505_, new_n1462_, new_n619_, new_n1890_, new_n471_, new_n967_, new_n577_, new_n1135_, new_n376_, new_n1538_, new_n1579_, new_n1289_, new_n1561_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n1095_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n1776_, new_n1621_, new_n839_, new_n1030_, new_n2078_, new_n485_, new_n578_, new_n525_, new_n1695_, new_n918_, new_n1586_, new_n1805_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n1572_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n1387_, new_n719_, new_n869_, new_n1178_, new_n1775_, new_n1525_, new_n570_, new_n598_, new_n893_, new_n1935_, new_n1063_, new_n520_, new_n1347_, new_n1001_, new_n1917_, new_n825_, new_n1627_, new_n557_, new_n1642_, new_n1807_, new_n1503_, new_n1742_, new_n507_, new_n741_, new_n806_, new_n1699_, new_n605_, new_n1224_, new_n2008_, new_n748_, new_n1074_, new_n1137_, new_n1286_, new_n1551_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n1650_, new_n807_, new_n1326_, new_n592_, new_n1820_, new_n726_, new_n1763_, new_n1263_, new_n1123_, new_n2020_, new_n1080_, new_n583_, new_n617_, new_n1279_, new_n1467_, new_n522_, new_n588_, new_n1762_, new_n1997_, new_n916_, new_n781_, new_n1014_, new_n428_, new_n1855_, new_n487_, new_n675_, new_n1155_, new_n360_, new_n1186_, new_n1915_, new_n1596_, new_n1848_, new_n1261_, new_n2022_, new_n2002_, new_n1863_, new_n1246_, new_n1488_, new_n2024_, new_n922_, new_n2029_, new_n387_, new_n476_, new_n987_, new_n1641_, new_n1951_, new_n949_, new_n2048_, new_n450_, new_n1394_, new_n1179_, new_n1088_, new_n1148_, new_n1146_, new_n1756_, new_n569_, new_n555_, new_n468_, new_n977_, new_n2049_, new_n1139_, new_n782_, new_n1793_, new_n444_, new_n392_, new_n518_, new_n950_, new_n1845_, new_n737_, new_n1022_, new_n692_, new_n502_, new_n1821_, new_n1888_, new_n623_, new_n446_, new_n2089_, new_n590_, new_n826_, new_n2079_, new_n789_, new_n1476_, new_n515_, new_n1854_, new_n972_, new_n1634_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n1835_, new_n1916_, new_n2046_, new_n733_, new_n1983_, new_n1021_, new_n1076_, new_n585_, new_n2076_, new_n1350_, new_n535_, new_n1976_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n1736_, new_n1945_, new_n1378_, new_n1478_, new_n1181_, new_n1093_, new_n597_, new_n1451_, new_n1092_, new_n1783_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1779_, new_n1869_, new_n1296_, new_n435_, new_n1891_, new_n1719_, new_n1883_, new_n1309_, new_n1796_, new_n1010_, new_n776_, new_n1830_, new_n2053_, new_n1885_, new_n687_, new_n1029_, new_n1649_, new_n1862_, new_n1654_, new_n1515_, new_n1746_, new_n638_, new_n523_, new_n909_, new_n1840_, new_n1688_, new_n1963_, new_n1571_, new_n1773_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1610_, new_n1470_, new_n1112_, new_n1715_, new_n1156_, new_n711_, new_n1938_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1475_, new_n1604_, new_n1260_, new_n973_, new_n1529_, new_n607_, new_n1731_, new_n1541_, new_n645_, new_n1087_, new_n1096_, new_n723_, new_n1599_, new_n756_, new_n823_, new_n1549_, new_n1933_, new_n1577_, new_n574_, new_n1500_, new_n928_, new_n1548_, new_n1578_, new_n1008_, new_n2059_, new_n1687_, new_n1661_, new_n1615_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n1291_, new_n539_, new_n1399_, new_n803_, new_n1817_, new_n727_, new_n1531_, new_n1672_, new_n1927_, new_n1589_, new_n2061_, new_n1792_, new_n1965_, new_n1295_, new_n1173_, new_n704_, new_n2087_, new_n1809_, new_n1432_, new_n1570_, new_n1811_, new_n2004_, new_n1189_, new_n1197_, new_n1312_, new_n1502_, new_n1778_, new_n1874_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n467_, new_n404_, new_n1243_, new_n1077_, new_n2067_, new_n490_, new_n560_, new_n1100_, new_n1666_, new_n865_, new_n1744_, new_n358_, new_n877_, new_n1506_, new_n1583_, new_n2085_, new_n1697_, new_n545_, new_n611_, new_n1998_, new_n1011_, new_n425_, new_n896_, new_n1831_, new_n802_, new_n1925_, new_n1236_, new_n1829_, new_n1770_, new_n866_, new_n1556_, new_n947_, new_n994_, new_n1813_, new_n982_, new_n1494_, new_n1449_, new_n964_, new_n1078_, new_n1961_, new_n551_, new_n1408_, new_n455_, new_n1982_, new_n1569_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n1918_, new_n1605_, new_n464_, new_n1498_, new_n2097_, new_n1588_, new_n1974_, new_n573_, new_n765_, new_n1964_, new_n1314_, new_n1892_;

not g0000 ( new_n343_, N75 );
nand g0001 ( new_n344_, N29, N42 );
nor g0002 ( N388, new_n344_, new_n343_ );
not g0003 ( new_n346_, N80 );
nand g0004 ( new_n347_, N29, N36 );
nor g0005 ( N389, new_n347_, new_n346_ );
not g0006 ( new_n349_, N42 );
nor g0007 ( N390, new_n347_, new_n349_ );
nand g0008 ( new_n351_, N85, N86 );
not g0009 ( N391, new_n351_ );
not g0010 ( new_n353_, N17 );
nand g0011 ( new_n354_, N1, N8 );
not g0012 ( new_n355_, new_n354_ );
nand g0013 ( new_n356_, new_n355_, N13 );
nor g0014 ( N418, new_n356_, new_n353_ );
nand g0015 ( new_n358_, N1, N26 );
nand g0016 ( new_n359_, N13, N17 );
nor g0017 ( new_n360_, new_n358_, new_n359_ );
not g0018 ( new_n361_, new_n360_ );
nor g0019 ( new_n362_, new_n361_, N390 );
not g0020 ( new_n363_, new_n362_ );
nand g0021 ( new_n364_, new_n363_, keyIn_0_8 );
not g0022 ( new_n365_, keyIn_0_8 );
nand g0023 ( new_n366_, new_n362_, new_n365_ );
nand g0024 ( N419, new_n364_, new_n366_ );
nand g0025 ( new_n368_, N59, N75 );
not g0026 ( new_n369_, new_n368_ );
nand g0027 ( N420, new_n369_, N80 );
nand g0028 ( new_n371_, N36, N59 );
not g0029 ( new_n372_, new_n371_ );
nand g0030 ( N421, new_n372_, N80 );
nand g0031 ( N422, new_n372_, N42 );
not g0032 ( new_n375_, N90 );
nor g0033 ( new_n376_, N87, N88 );
nor g0034 ( N423, new_n376_, new_n375_ );
nand g0035 ( new_n378_, new_n360_, N390 );
nand g0036 ( new_n379_, new_n378_, keyIn_0_25 );
not g0037 ( new_n380_, keyIn_0_25 );
not g0038 ( new_n381_, new_n378_ );
nand g0039 ( new_n382_, new_n381_, new_n380_ );
nand g0040 ( N446, new_n382_, new_n379_ );
not g0041 ( new_n384_, keyIn_0_0 );
not g0042 ( new_n385_, N51 );
nor g0043 ( new_n386_, new_n358_, new_n385_ );
nor g0044 ( new_n387_, new_n386_, new_n384_ );
not g0045 ( new_n388_, new_n358_ );
nand g0046 ( new_n389_, new_n388_, N51 );
nor g0047 ( new_n390_, new_n389_, keyIn_0_0 );
nor g0048 ( N447, new_n390_, new_n387_ );
not g0049 ( new_n392_, N55 );
nor g0050 ( new_n393_, new_n356_, new_n392_ );
not g0051 ( new_n394_, new_n393_ );
nand g0052 ( new_n395_, N29, N68 );
nor g0053 ( new_n396_, new_n394_, new_n395_ );
not g0054 ( new_n397_, new_n396_ );
nand g0055 ( new_n398_, new_n397_, keyIn_0_12 );
not g0056 ( new_n399_, keyIn_0_12 );
nand g0057 ( new_n400_, new_n396_, new_n399_ );
nand g0058 ( N448, new_n398_, new_n400_ );
not g0059 ( new_n402_, N74 );
nand g0060 ( new_n403_, N59, N68 );
nor g0061 ( new_n404_, new_n403_, new_n402_ );
nand g0062 ( new_n405_, new_n393_, new_n404_ );
nand g0063 ( new_n406_, new_n405_, keyIn_0_13 );
not g0064 ( new_n407_, keyIn_0_13 );
not g0065 ( new_n408_, new_n405_ );
nand g0066 ( new_n409_, new_n408_, new_n407_ );
nand g0067 ( N449, new_n409_, new_n406_ );
not g0068 ( new_n411_, N89 );
nor g0069 ( N450, new_n376_, new_n411_ );
not g0070 ( new_n413_, keyIn_0_139 );
not g0071 ( new_n414_, keyIn_0_106 );
not g0072 ( new_n415_, keyIn_0_95 );
not g0073 ( new_n416_, keyIn_0_73 );
not g0074 ( new_n417_, keyIn_0_53 );
not g0075 ( new_n418_, keyIn_0_43 );
not g0076 ( new_n419_, keyIn_0_32 );
nor g0077 ( new_n420_, N121, N126 );
nand g0078 ( new_n421_, N121, N126 );
not g0079 ( new_n422_, new_n421_ );
nor g0080 ( new_n423_, new_n422_, new_n420_ );
not g0081 ( new_n424_, new_n423_ );
nor g0082 ( new_n425_, new_n424_, keyIn_0_18 );
nand g0083 ( new_n426_, new_n424_, keyIn_0_18 );
not g0084 ( new_n427_, new_n426_ );
nor g0085 ( new_n428_, new_n427_, new_n425_ );
not g0086 ( new_n429_, new_n428_ );
nor g0087 ( new_n430_, new_n429_, new_n419_ );
nor g0088 ( new_n431_, new_n428_, keyIn_0_32 );
nor g0089 ( new_n432_, new_n430_, new_n431_ );
not g0090 ( new_n433_, keyIn_0_31 );
not g0091 ( new_n434_, N111 );
nor g0092 ( new_n435_, new_n434_, N116 );
not g0093 ( new_n436_, N116 );
nor g0094 ( new_n437_, new_n436_, N111 );
nor g0095 ( new_n438_, new_n435_, new_n437_ );
not g0096 ( new_n439_, new_n438_ );
nand g0097 ( new_n440_, new_n439_, keyIn_0_17 );
not g0098 ( new_n441_, new_n440_ );
nor g0099 ( new_n442_, new_n439_, keyIn_0_17 );
nor g0100 ( new_n443_, new_n441_, new_n442_ );
not g0101 ( new_n444_, new_n443_ );
nor g0102 ( new_n445_, new_n444_, new_n433_ );
nor g0103 ( new_n446_, new_n443_, keyIn_0_31 );
nor g0104 ( new_n447_, new_n445_, new_n446_ );
nor g0105 ( new_n448_, new_n447_, new_n432_ );
not g0106 ( new_n449_, new_n448_ );
nand g0107 ( new_n450_, new_n449_, new_n418_ );
not g0108 ( new_n451_, new_n450_ );
nor g0109 ( new_n452_, new_n449_, new_n418_ );
nor g0110 ( new_n453_, new_n451_, new_n452_ );
not g0111 ( new_n454_, keyIn_0_33 );
nor g0112 ( new_n455_, new_n443_, new_n428_ );
not g0113 ( new_n456_, new_n455_ );
nand g0114 ( new_n457_, new_n456_, new_n454_ );
not g0115 ( new_n458_, new_n457_ );
nor g0116 ( new_n459_, new_n456_, new_n454_ );
nor g0117 ( new_n460_, new_n458_, new_n459_ );
nor g0118 ( new_n461_, new_n453_, new_n460_ );
not g0119 ( new_n462_, new_n461_ );
nor g0120 ( new_n463_, new_n462_, new_n417_ );
nor g0121 ( new_n464_, new_n461_, keyIn_0_53 );
nor g0122 ( new_n465_, new_n463_, new_n464_ );
not g0123 ( new_n466_, new_n465_ );
nor g0124 ( new_n467_, new_n466_, N135 );
nor g0125 ( new_n468_, new_n467_, new_n416_ );
nand g0126 ( new_n469_, new_n467_, new_n416_ );
not g0127 ( new_n470_, new_n469_ );
nor g0128 ( new_n471_, new_n470_, new_n468_ );
nand g0129 ( new_n472_, new_n466_, N135 );
nand g0130 ( new_n473_, new_n472_, keyIn_0_72 );
not g0131 ( new_n474_, new_n473_ );
nor g0132 ( new_n475_, new_n472_, keyIn_0_72 );
nor g0133 ( new_n476_, new_n474_, new_n475_ );
nor g0134 ( new_n477_, new_n471_, new_n476_ );
not g0135 ( new_n478_, new_n477_ );
nand g0136 ( new_n479_, new_n478_, new_n415_ );
not g0137 ( new_n480_, new_n479_ );
nor g0138 ( new_n481_, new_n478_, new_n415_ );
nor g0139 ( new_n482_, new_n480_, new_n481_ );
not g0140 ( new_n483_, keyIn_0_71 );
not g0141 ( new_n484_, keyIn_0_52 );
not g0142 ( new_n485_, keyIn_0_28 );
nor g0143 ( new_n486_, N91, N96 );
nand g0144 ( new_n487_, N91, N96 );
not g0145 ( new_n488_, new_n487_ );
nor g0146 ( new_n489_, new_n488_, new_n486_ );
not g0147 ( new_n490_, new_n489_ );
nor g0148 ( new_n491_, new_n490_, keyIn_0_15 );
nand g0149 ( new_n492_, new_n490_, keyIn_0_15 );
not g0150 ( new_n493_, new_n492_ );
nor g0151 ( new_n494_, new_n493_, new_n491_ );
not g0152 ( new_n495_, new_n494_ );
nor g0153 ( new_n496_, new_n495_, new_n485_ );
nor g0154 ( new_n497_, new_n494_, keyIn_0_28 );
nor g0155 ( new_n498_, new_n496_, new_n497_ );
not g0156 ( new_n499_, keyIn_0_29 );
not g0157 ( new_n500_, N101 );
nor g0158 ( new_n501_, new_n500_, N106 );
not g0159 ( new_n502_, N106 );
nor g0160 ( new_n503_, new_n502_, N101 );
nor g0161 ( new_n504_, new_n501_, new_n503_ );
not g0162 ( new_n505_, new_n504_ );
nand g0163 ( new_n506_, new_n505_, keyIn_0_16 );
not g0164 ( new_n507_, new_n506_ );
nor g0165 ( new_n508_, new_n505_, keyIn_0_16 );
nor g0166 ( new_n509_, new_n507_, new_n508_ );
not g0167 ( new_n510_, new_n509_ );
nor g0168 ( new_n511_, new_n510_, new_n499_ );
nor g0169 ( new_n512_, new_n509_, keyIn_0_29 );
nor g0170 ( new_n513_, new_n511_, new_n512_ );
nor g0171 ( new_n514_, new_n513_, new_n498_ );
not g0172 ( new_n515_, new_n514_ );
nor g0173 ( new_n516_, new_n515_, keyIn_0_42 );
nand g0174 ( new_n517_, new_n515_, keyIn_0_42 );
not g0175 ( new_n518_, keyIn_0_30 );
nand g0176 ( new_n519_, new_n510_, new_n495_ );
nor g0177 ( new_n520_, new_n519_, new_n518_ );
nand g0178 ( new_n521_, new_n519_, new_n518_ );
not g0179 ( new_n522_, new_n521_ );
nor g0180 ( new_n523_, new_n522_, new_n520_ );
nand g0181 ( new_n524_, new_n517_, new_n523_ );
nor g0182 ( new_n525_, new_n524_, new_n516_ );
nor g0183 ( new_n526_, new_n525_, new_n484_ );
nand g0184 ( new_n527_, new_n525_, new_n484_ );
not g0185 ( new_n528_, new_n527_ );
nor g0186 ( new_n529_, new_n528_, new_n526_ );
not g0187 ( new_n530_, new_n529_ );
nor g0188 ( new_n531_, new_n530_, N130 );
nor g0189 ( new_n532_, new_n531_, new_n483_ );
nand g0190 ( new_n533_, new_n531_, new_n483_ );
not g0191 ( new_n534_, new_n533_ );
nor g0192 ( new_n535_, new_n534_, new_n532_ );
not g0193 ( new_n536_, keyIn_0_70 );
not g0194 ( new_n537_, N130 );
nor g0195 ( new_n538_, new_n529_, new_n537_ );
not g0196 ( new_n539_, new_n538_ );
nand g0197 ( new_n540_, new_n539_, new_n536_ );
not g0198 ( new_n541_, new_n540_ );
nor g0199 ( new_n542_, new_n539_, new_n536_ );
nor g0200 ( new_n543_, new_n541_, new_n542_ );
nor g0201 ( new_n544_, new_n543_, new_n535_ );
not g0202 ( new_n545_, new_n544_ );
nand g0203 ( new_n546_, new_n545_, keyIn_0_94 );
not g0204 ( new_n547_, new_n546_ );
nor g0205 ( new_n548_, new_n545_, keyIn_0_94 );
nor g0206 ( new_n549_, new_n547_, new_n548_ );
nor g0207 ( new_n550_, new_n482_, new_n549_ );
not g0208 ( new_n551_, new_n550_ );
nand g0209 ( new_n552_, new_n551_, new_n414_ );
nand g0210 ( new_n553_, new_n550_, keyIn_0_106 );
nand g0211 ( new_n554_, new_n552_, new_n553_ );
not g0212 ( new_n555_, keyIn_0_116 );
nand g0213 ( new_n556_, new_n482_, new_n549_ );
not g0214 ( new_n557_, new_n556_ );
nand g0215 ( new_n558_, new_n557_, new_n555_ );
nand g0216 ( new_n559_, new_n556_, keyIn_0_116 );
nand g0217 ( new_n560_, new_n558_, new_n559_ );
nand g0218 ( new_n561_, new_n554_, new_n560_ );
not g0219 ( new_n562_, new_n561_ );
nand g0220 ( new_n563_, new_n562_, new_n413_ );
nand g0221 ( new_n564_, new_n561_, keyIn_0_139 );
nand g0222 ( N767, new_n563_, new_n564_ );
not g0223 ( new_n566_, keyIn_0_140 );
not g0224 ( new_n567_, keyIn_0_91 );
not g0225 ( new_n568_, keyIn_0_36 );
nor g0226 ( new_n569_, N171, N177 );
nand g0227 ( new_n570_, N171, N177 );
not g0228 ( new_n571_, new_n570_ );
nor g0229 ( new_n572_, new_n571_, new_n569_ );
not g0230 ( new_n573_, new_n572_ );
nor g0231 ( new_n574_, new_n573_, keyIn_0_22 );
nand g0232 ( new_n575_, new_n573_, keyIn_0_22 );
not g0233 ( new_n576_, new_n575_ );
nor g0234 ( new_n577_, new_n576_, new_n574_ );
not g0235 ( new_n578_, new_n577_ );
nor g0236 ( new_n579_, new_n578_, new_n568_ );
nor g0237 ( new_n580_, new_n577_, keyIn_0_36 );
nor g0238 ( new_n581_, new_n579_, new_n580_ );
not g0239 ( new_n582_, keyIn_0_35 );
not g0240 ( new_n583_, N159 );
nor g0241 ( new_n584_, new_n583_, N165 );
not g0242 ( new_n585_, N165 );
nor g0243 ( new_n586_, new_n585_, N159 );
nor g0244 ( new_n587_, new_n584_, new_n586_ );
not g0245 ( new_n588_, new_n587_ );
nand g0246 ( new_n589_, new_n588_, keyIn_0_21 );
not g0247 ( new_n590_, new_n589_ );
nor g0248 ( new_n591_, new_n588_, keyIn_0_21 );
nor g0249 ( new_n592_, new_n590_, new_n591_ );
not g0250 ( new_n593_, new_n592_ );
nor g0251 ( new_n594_, new_n593_, new_n582_ );
nor g0252 ( new_n595_, new_n592_, keyIn_0_35 );
nor g0253 ( new_n596_, new_n594_, new_n595_ );
nor g0254 ( new_n597_, new_n596_, new_n581_ );
not g0255 ( new_n598_, new_n597_ );
nand g0256 ( new_n599_, new_n598_, keyIn_0_49 );
not g0257 ( new_n600_, new_n599_ );
nor g0258 ( new_n601_, new_n598_, keyIn_0_49 );
nor g0259 ( new_n602_, new_n600_, new_n601_ );
not g0260 ( new_n603_, keyIn_0_37 );
nor g0261 ( new_n604_, new_n592_, new_n577_ );
not g0262 ( new_n605_, new_n604_ );
nand g0263 ( new_n606_, new_n605_, new_n603_ );
not g0264 ( new_n607_, new_n606_ );
nor g0265 ( new_n608_, new_n605_, new_n603_ );
nor g0266 ( new_n609_, new_n607_, new_n608_ );
nor g0267 ( new_n610_, new_n602_, new_n609_ );
not g0268 ( new_n611_, new_n610_ );
nor g0269 ( new_n612_, new_n611_, keyIn_0_68 );
nand g0270 ( new_n613_, new_n611_, keyIn_0_68 );
not g0271 ( new_n614_, new_n613_ );
nor g0272 ( new_n615_, new_n614_, new_n612_ );
not g0273 ( new_n616_, new_n615_ );
nor g0274 ( new_n617_, new_n616_, N130 );
nor g0275 ( new_n618_, new_n617_, new_n567_ );
nand g0276 ( new_n619_, new_n617_, new_n567_ );
not g0277 ( new_n620_, new_n619_ );
nor g0278 ( new_n621_, new_n620_, new_n618_ );
nor g0279 ( new_n622_, new_n615_, new_n537_ );
not g0280 ( new_n623_, new_n622_ );
nand g0281 ( new_n624_, new_n623_, keyIn_0_90 );
not g0282 ( new_n625_, new_n624_ );
nor g0283 ( new_n626_, new_n623_, keyIn_0_90 );
nor g0284 ( new_n627_, new_n625_, new_n626_ );
nor g0285 ( new_n628_, new_n627_, new_n621_ );
not g0286 ( new_n629_, new_n628_ );
nand g0287 ( new_n630_, new_n629_, keyIn_0_104 );
not g0288 ( new_n631_, new_n630_ );
nor g0289 ( new_n632_, new_n629_, keyIn_0_104 );
nor g0290 ( new_n633_, new_n631_, new_n632_ );
not g0291 ( new_n634_, keyIn_0_105 );
not g0292 ( new_n635_, keyIn_0_93 );
not g0293 ( new_n636_, keyIn_0_69 );
not g0294 ( new_n637_, N183 );
nor g0295 ( new_n638_, new_n637_, N189 );
not g0296 ( new_n639_, N189 );
nor g0297 ( new_n640_, new_n639_, N183 );
nor g0298 ( new_n641_, new_n638_, new_n640_ );
not g0299 ( new_n642_, new_n641_ );
nand g0300 ( new_n643_, new_n642_, keyIn_0_23 );
not g0301 ( new_n644_, new_n643_ );
nor g0302 ( new_n645_, new_n642_, keyIn_0_23 );
nor g0303 ( new_n646_, new_n644_, new_n645_ );
not g0304 ( new_n647_, new_n646_ );
nand g0305 ( new_n648_, new_n647_, keyIn_0_38 );
not g0306 ( new_n649_, keyIn_0_38 );
nand g0307 ( new_n650_, new_n646_, new_n649_ );
nand g0308 ( new_n651_, new_n648_, new_n650_ );
not g0309 ( new_n652_, N195 );
nor g0310 ( new_n653_, new_n652_, N201 );
not g0311 ( new_n654_, N201 );
nor g0312 ( new_n655_, new_n654_, N195 );
nor g0313 ( new_n656_, new_n653_, new_n655_ );
not g0314 ( new_n657_, new_n656_ );
nand g0315 ( new_n658_, new_n657_, keyIn_0_24 );
not g0316 ( new_n659_, new_n658_ );
nor g0317 ( new_n660_, new_n657_, keyIn_0_24 );
nor g0318 ( new_n661_, new_n659_, new_n660_ );
not g0319 ( new_n662_, new_n661_ );
nand g0320 ( new_n663_, new_n662_, keyIn_0_39 );
not g0321 ( new_n664_, keyIn_0_39 );
nand g0322 ( new_n665_, new_n661_, new_n664_ );
nand g0323 ( new_n666_, new_n663_, new_n665_ );
nand g0324 ( new_n667_, new_n651_, new_n666_ );
nand g0325 ( new_n668_, new_n667_, keyIn_0_50 );
nor g0326 ( new_n669_, new_n646_, new_n661_ );
not g0327 ( new_n670_, new_n669_ );
nand g0328 ( new_n671_, new_n670_, keyIn_0_40 );
not g0329 ( new_n672_, new_n671_ );
nor g0330 ( new_n673_, new_n670_, keyIn_0_40 );
nor g0331 ( new_n674_, new_n672_, new_n673_ );
nor g0332 ( new_n675_, new_n667_, keyIn_0_50 );
nor g0333 ( new_n676_, new_n674_, new_n675_ );
nand g0334 ( new_n677_, new_n676_, new_n668_ );
nor g0335 ( new_n678_, new_n677_, new_n636_ );
nand g0336 ( new_n679_, new_n677_, new_n636_ );
not g0337 ( new_n680_, new_n679_ );
nor g0338 ( new_n681_, new_n680_, new_n678_ );
nor g0339 ( new_n682_, new_n681_, N207 );
not g0340 ( new_n683_, new_n682_ );
nand g0341 ( new_n684_, new_n683_, new_n635_ );
not g0342 ( new_n685_, new_n684_ );
nor g0343 ( new_n686_, new_n683_, new_n635_ );
nor g0344 ( new_n687_, new_n685_, new_n686_ );
nand g0345 ( new_n688_, new_n681_, N207 );
nor g0346 ( new_n689_, new_n688_, keyIn_0_92 );
nand g0347 ( new_n690_, new_n688_, keyIn_0_92 );
not g0348 ( new_n691_, new_n690_ );
nor g0349 ( new_n692_, new_n691_, new_n689_ );
nor g0350 ( new_n693_, new_n687_, new_n692_ );
not g0351 ( new_n694_, new_n693_ );
nand g0352 ( new_n695_, new_n694_, new_n634_ );
not g0353 ( new_n696_, new_n695_ );
nor g0354 ( new_n697_, new_n694_, new_n634_ );
nor g0355 ( new_n698_, new_n696_, new_n697_ );
nor g0356 ( new_n699_, new_n633_, new_n698_ );
not g0357 ( new_n700_, new_n699_ );
nand g0358 ( new_n701_, new_n700_, keyIn_0_115 );
not g0359 ( new_n702_, keyIn_0_115 );
nand g0360 ( new_n703_, new_n699_, new_n702_ );
nand g0361 ( new_n704_, new_n701_, new_n703_ );
not g0362 ( new_n705_, keyIn_0_117 );
nand g0363 ( new_n706_, new_n633_, new_n698_ );
not g0364 ( new_n707_, new_n706_ );
nand g0365 ( new_n708_, new_n707_, new_n705_ );
nand g0366 ( new_n709_, new_n706_, keyIn_0_117 );
nand g0367 ( new_n710_, new_n708_, new_n709_ );
nand g0368 ( new_n711_, new_n704_, new_n710_ );
not g0369 ( new_n712_, new_n711_ );
nand g0370 ( new_n713_, new_n712_, new_n566_ );
nand g0371 ( new_n714_, new_n711_, keyIn_0_140 );
nand g0372 ( N768, new_n713_, new_n714_ );
not g0373 ( new_n716_, keyIn_0_210 );
not g0374 ( new_n717_, keyIn_0_202 );
not g0375 ( new_n718_, keyIn_0_163 );
not g0376 ( new_n719_, keyIn_0_114 );
not g0377 ( new_n720_, keyIn_0_103 );
not g0378 ( new_n721_, keyIn_0_88 );
not g0379 ( new_n722_, keyIn_0_5 );
nand g0380 ( new_n723_, N59, N156 );
nor g0381 ( new_n724_, new_n723_, new_n722_ );
nand g0382 ( new_n725_, new_n723_, new_n722_ );
not g0383 ( new_n726_, new_n725_ );
nor g0384 ( new_n727_, new_n726_, new_n724_ );
not g0385 ( new_n728_, keyIn_0_26 );
nor g0386 ( new_n729_, N447, keyIn_0_9 );
not g0387 ( new_n730_, keyIn_0_9 );
nand g0388 ( new_n731_, new_n389_, keyIn_0_0 );
nand g0389 ( new_n732_, new_n386_, new_n384_ );
nand g0390 ( new_n733_, new_n731_, new_n732_ );
nor g0391 ( new_n734_, new_n733_, new_n730_ );
nor g0392 ( new_n735_, new_n729_, new_n734_ );
nor g0393 ( new_n736_, new_n735_, new_n728_ );
nand g0394 ( new_n737_, new_n733_, new_n730_ );
nand g0395 ( new_n738_, N447, keyIn_0_9 );
nand g0396 ( new_n739_, new_n738_, new_n737_ );
nor g0397 ( new_n740_, new_n739_, keyIn_0_26 );
nor g0398 ( new_n741_, new_n736_, new_n740_ );
nor g0399 ( new_n742_, new_n741_, new_n353_ );
nand g0400 ( new_n743_, new_n742_, new_n727_ );
nand g0401 ( new_n744_, new_n743_, keyIn_0_48 );
not g0402 ( new_n745_, keyIn_0_48 );
not g0403 ( new_n746_, new_n727_ );
nand g0404 ( new_n747_, new_n739_, keyIn_0_26 );
nand g0405 ( new_n748_, new_n735_, new_n728_ );
nand g0406 ( new_n749_, new_n748_, new_n747_ );
nand g0407 ( new_n750_, new_n749_, N17 );
nor g0408 ( new_n751_, new_n750_, new_n746_ );
nand g0409 ( new_n752_, new_n751_, new_n745_ );
nand g0410 ( new_n753_, new_n744_, new_n752_ );
nand g0411 ( new_n754_, new_n753_, N1 );
nor g0412 ( new_n755_, new_n754_, keyIn_0_63 );
nand g0413 ( new_n756_, new_n754_, keyIn_0_63 );
nand g0414 ( new_n757_, new_n756_, N153 );
nor g0415 ( new_n758_, new_n757_, new_n755_ );
nand g0416 ( new_n759_, new_n758_, new_n721_ );
not g0417 ( new_n760_, new_n755_ );
not g0418 ( new_n761_, new_n757_ );
nand g0419 ( new_n762_, new_n761_, new_n760_ );
nand g0420 ( new_n763_, new_n762_, keyIn_0_88 );
nand g0421 ( new_n764_, new_n763_, new_n759_ );
not g0422 ( new_n765_, keyIn_0_89 );
not g0423 ( new_n766_, keyIn_0_54 );
not g0424 ( new_n767_, keyIn_0_20 );
nand g0425 ( new_n768_, N17, N42 );
not g0426 ( new_n769_, new_n768_ );
nand g0427 ( new_n770_, new_n769_, keyIn_0_7 );
not g0428 ( new_n771_, keyIn_0_7 );
nand g0429 ( new_n772_, new_n768_, new_n771_ );
nand g0430 ( new_n773_, new_n770_, new_n772_ );
nor g0431 ( new_n774_, N17, N42 );
nor g0432 ( new_n775_, new_n774_, keyIn_0_6 );
not g0433 ( new_n776_, keyIn_0_6 );
not g0434 ( new_n777_, new_n774_ );
nor g0435 ( new_n778_, new_n777_, new_n776_ );
nor g0436 ( new_n779_, new_n778_, new_n775_ );
nand g0437 ( new_n780_, new_n779_, new_n773_ );
nor g0438 ( new_n781_, new_n780_, new_n767_ );
not g0439 ( new_n782_, new_n723_ );
nand g0440 ( new_n783_, new_n780_, new_n767_ );
nand g0441 ( new_n784_, new_n783_, new_n782_ );
nor g0442 ( new_n785_, new_n784_, new_n781_ );
nand g0443 ( new_n786_, new_n749_, new_n785_ );
nor g0444 ( new_n787_, new_n786_, keyIn_0_47 );
nand g0445 ( new_n788_, new_n786_, keyIn_0_47 );
not g0446 ( new_n789_, keyIn_0_34 );
not g0447 ( new_n790_, keyIn_0_3 );
nand g0448 ( new_n791_, N42, N59 );
nor g0449 ( new_n792_, new_n791_, new_n343_ );
not g0450 ( new_n793_, new_n792_ );
nor g0451 ( new_n794_, new_n793_, new_n790_ );
nor g0452 ( new_n795_, new_n792_, keyIn_0_3 );
nor g0453 ( new_n796_, new_n794_, new_n795_ );
not g0454 ( new_n797_, new_n796_ );
nand g0455 ( new_n798_, new_n797_, keyIn_0_14 );
not g0456 ( new_n799_, keyIn_0_14 );
nand g0457 ( new_n800_, new_n796_, new_n799_ );
nand g0458 ( new_n801_, new_n798_, new_n800_ );
nand g0459 ( new_n802_, N17, N51 );
nor g0460 ( new_n803_, new_n354_, new_n802_ );
nor g0461 ( new_n804_, new_n803_, keyIn_0_1 );
nand g0462 ( new_n805_, new_n803_, keyIn_0_1 );
not g0463 ( new_n806_, new_n805_ );
nor g0464 ( new_n807_, new_n806_, new_n804_ );
not g0465 ( new_n808_, new_n807_ );
nand g0466 ( new_n809_, new_n808_, keyIn_0_10 );
not g0467 ( new_n810_, keyIn_0_10 );
nand g0468 ( new_n811_, new_n807_, new_n810_ );
nand g0469 ( new_n812_, new_n809_, new_n811_ );
nand g0470 ( new_n813_, new_n801_, new_n812_ );
nor g0471 ( new_n814_, new_n813_, new_n789_ );
nand g0472 ( new_n815_, new_n813_, new_n789_ );
not g0473 ( new_n816_, new_n815_ );
nor g0474 ( new_n817_, new_n816_, new_n814_ );
nand g0475 ( new_n818_, new_n817_, new_n788_ );
nor g0476 ( new_n819_, new_n818_, new_n787_ );
nand g0477 ( new_n820_, new_n819_, new_n766_ );
not g0478 ( new_n821_, new_n820_ );
nor g0479 ( new_n822_, new_n819_, new_n766_ );
nor g0480 ( new_n823_, new_n821_, new_n822_ );
nand g0481 ( new_n824_, new_n823_, N126 );
nand g0482 ( new_n825_, new_n824_, new_n765_ );
not g0483 ( new_n826_, N126 );
not g0484 ( new_n827_, new_n819_ );
nand g0485 ( new_n828_, new_n827_, keyIn_0_54 );
nand g0486 ( new_n829_, new_n828_, new_n820_ );
nor g0487 ( new_n830_, new_n829_, new_n826_ );
nand g0488 ( new_n831_, new_n830_, keyIn_0_89 );
nand g0489 ( new_n832_, new_n825_, new_n831_ );
nand g0490 ( new_n833_, new_n764_, new_n832_ );
nand g0491 ( new_n834_, new_n833_, new_n720_ );
not g0492 ( new_n835_, keyIn_0_67 );
nor g0493 ( new_n836_, new_n741_, new_n392_ );
not g0494 ( new_n837_, new_n836_ );
nand g0495 ( new_n838_, N29, N75 );
nor g0496 ( new_n839_, new_n838_, new_n346_ );
not g0497 ( new_n840_, new_n839_ );
nor g0498 ( new_n841_, new_n840_, keyIn_0_2 );
nand g0499 ( new_n842_, new_n840_, keyIn_0_2 );
not g0500 ( new_n843_, new_n842_ );
nor g0501 ( new_n844_, new_n843_, new_n841_ );
not g0502 ( new_n845_, new_n844_ );
nor g0503 ( new_n846_, new_n837_, new_n845_ );
not g0504 ( new_n847_, new_n846_ );
nor g0505 ( new_n848_, new_n847_, keyIn_0_46 );
not g0506 ( new_n849_, keyIn_0_19 );
nand g0507 ( new_n850_, keyIn_0_4, N268 );
not g0508 ( new_n851_, new_n850_ );
nor g0509 ( new_n852_, keyIn_0_4, N268 );
nor g0510 ( new_n853_, new_n851_, new_n852_ );
not g0511 ( new_n854_, new_n853_ );
nor g0512 ( new_n855_, new_n854_, new_n849_ );
nor g0513 ( new_n856_, new_n853_, keyIn_0_19 );
nor g0514 ( new_n857_, new_n855_, new_n856_ );
nand g0515 ( new_n858_, new_n847_, keyIn_0_46 );
nand g0516 ( new_n859_, new_n858_, new_n857_ );
nor g0517 ( new_n860_, new_n859_, new_n848_ );
nor g0518 ( new_n861_, new_n860_, new_n835_ );
not g0519 ( new_n862_, new_n860_ );
nor g0520 ( new_n863_, new_n862_, keyIn_0_67 );
nor g0521 ( new_n864_, new_n863_, new_n861_ );
nor g0522 ( new_n865_, new_n833_, new_n720_ );
nor g0523 ( new_n866_, new_n865_, new_n864_ );
nand g0524 ( new_n867_, new_n866_, new_n834_ );
nand g0525 ( new_n868_, new_n867_, new_n719_ );
not g0526 ( new_n869_, new_n834_ );
not g0527 ( new_n870_, new_n864_ );
not g0528 ( new_n871_, new_n759_ );
nor g0529 ( new_n872_, new_n758_, new_n721_ );
nor g0530 ( new_n873_, new_n871_, new_n872_ );
not g0531 ( new_n874_, new_n832_ );
nor g0532 ( new_n875_, new_n873_, new_n874_ );
nand g0533 ( new_n876_, new_n875_, keyIn_0_103 );
nand g0534 ( new_n877_, new_n876_, new_n870_ );
nor g0535 ( new_n878_, new_n877_, new_n869_ );
nand g0536 ( new_n879_, new_n878_, keyIn_0_114 );
nand g0537 ( new_n880_, new_n879_, new_n868_ );
nor g0538 ( new_n881_, new_n880_, N201 );
nor g0539 ( new_n882_, new_n881_, keyIn_0_138 );
not g0540 ( new_n883_, keyIn_0_138 );
nor g0541 ( new_n884_, new_n878_, keyIn_0_114 );
nor g0542 ( new_n885_, new_n867_, new_n719_ );
nor g0543 ( new_n886_, new_n884_, new_n885_ );
nand g0544 ( new_n887_, new_n886_, new_n654_ );
nor g0545 ( new_n888_, new_n887_, new_n883_ );
nor g0546 ( new_n889_, new_n888_, new_n882_ );
nand g0547 ( new_n890_, new_n880_, N201 );
nor g0548 ( new_n891_, new_n890_, keyIn_0_137 );
nand g0549 ( new_n892_, new_n890_, keyIn_0_137 );
not g0550 ( new_n893_, new_n892_ );
nor g0551 ( new_n894_, new_n893_, new_n891_ );
nor g0552 ( new_n895_, new_n894_, new_n889_ );
not g0553 ( new_n896_, new_n895_ );
nand g0554 ( new_n897_, new_n896_, new_n718_ );
not g0555 ( new_n898_, new_n897_ );
nor g0556 ( new_n899_, new_n896_, new_n718_ );
nor g0557 ( new_n900_, new_n898_, new_n899_ );
not g0558 ( new_n901_, new_n900_ );
nor g0559 ( new_n902_, new_n901_, N261 );
not g0560 ( new_n903_, new_n902_ );
nand g0561 ( new_n904_, new_n903_, keyIn_0_184 );
not g0562 ( new_n905_, keyIn_0_184 );
nand g0563 ( new_n906_, new_n902_, new_n905_ );
nand g0564 ( new_n907_, new_n904_, new_n906_ );
not g0565 ( new_n908_, keyIn_0_185 );
not g0566 ( new_n909_, N261 );
nor g0567 ( new_n910_, new_n900_, new_n909_ );
not g0568 ( new_n911_, new_n910_ );
nand g0569 ( new_n912_, new_n911_, new_n908_ );
nand g0570 ( new_n913_, new_n910_, keyIn_0_185 );
nand g0571 ( new_n914_, new_n912_, new_n913_ );
nand g0572 ( new_n915_, new_n907_, new_n914_ );
nor g0573 ( new_n916_, new_n915_, new_n717_ );
nand g0574 ( new_n917_, new_n915_, new_n717_ );
nand g0575 ( new_n918_, new_n917_, N219 );
nor g0576 ( new_n919_, new_n918_, new_n916_ );
nor g0577 ( new_n920_, new_n919_, new_n716_ );
nand g0578 ( new_n921_, new_n919_, new_n716_ );
not g0579 ( new_n922_, new_n921_ );
nor g0580 ( new_n923_, new_n922_, new_n920_ );
nand g0581 ( new_n924_, N121, N210 );
not g0582 ( new_n925_, new_n924_ );
nor g0583 ( new_n926_, new_n923_, new_n925_ );
not g0584 ( new_n927_, new_n926_ );
nor g0585 ( new_n928_, new_n927_, keyIn_0_216 );
nand g0586 ( new_n929_, new_n927_, keyIn_0_216 );
not g0587 ( new_n930_, keyIn_0_203 );
nand g0588 ( new_n931_, new_n901_, N228 );
nand g0589 ( new_n932_, new_n894_, keyIn_0_162 );
not g0590 ( new_n933_, keyIn_0_162 );
not g0591 ( new_n934_, new_n891_ );
nand g0592 ( new_n935_, new_n934_, new_n892_ );
nand g0593 ( new_n936_, new_n935_, new_n933_ );
nand g0594 ( new_n937_, new_n932_, new_n936_ );
nand g0595 ( new_n938_, new_n937_, N237 );
nand g0596 ( new_n939_, new_n931_, new_n938_ );
nand g0597 ( new_n940_, new_n939_, new_n930_ );
not g0598 ( new_n941_, new_n940_ );
not g0599 ( new_n942_, new_n939_ );
nand g0600 ( new_n943_, new_n942_, keyIn_0_203 );
not g0601 ( new_n944_, keyIn_0_164 );
nand g0602 ( new_n945_, new_n880_, N246 );
nand g0603 ( new_n946_, N255, N267 );
nand g0604 ( new_n947_, new_n945_, new_n946_ );
nor g0605 ( new_n948_, new_n947_, new_n944_ );
not g0606 ( new_n949_, keyIn_0_51 );
not g0607 ( new_n950_, N73 );
not g0608 ( new_n951_, keyIn_0_11 );
nand g0609 ( new_n952_, N68, N72 );
nor g0610 ( new_n953_, new_n791_, new_n952_ );
nand g0611 ( new_n954_, new_n393_, new_n953_ );
nor g0612 ( new_n955_, new_n954_, new_n951_ );
nand g0613 ( new_n956_, new_n954_, new_n951_ );
not g0614 ( new_n957_, new_n956_ );
nor g0615 ( new_n958_, new_n957_, new_n955_ );
nor g0616 ( new_n959_, new_n958_, new_n950_ );
not g0617 ( new_n960_, new_n959_ );
nand g0618 ( new_n961_, new_n960_, keyIn_0_27 );
not g0619 ( new_n962_, new_n961_ );
nor g0620 ( new_n963_, new_n960_, keyIn_0_27 );
nor g0621 ( new_n964_, new_n962_, new_n963_ );
not g0622 ( new_n965_, new_n964_ );
nor g0623 ( new_n966_, new_n965_, keyIn_0_41 );
nand g0624 ( new_n967_, new_n965_, keyIn_0_41 );
not g0625 ( new_n968_, new_n967_ );
nor g0626 ( new_n969_, new_n968_, new_n966_ );
not g0627 ( new_n970_, new_n969_ );
nor g0628 ( new_n971_, new_n970_, new_n949_ );
nor g0629 ( new_n972_, new_n969_, keyIn_0_51 );
nor g0630 ( new_n973_, new_n971_, new_n972_ );
nand g0631 ( new_n974_, new_n973_, N201 );
nand g0632 ( new_n975_, new_n947_, new_n944_ );
nand g0633 ( new_n976_, new_n975_, new_n974_ );
nor g0634 ( new_n977_, new_n976_, new_n948_ );
nand g0635 ( new_n978_, new_n943_, new_n977_ );
nor g0636 ( new_n979_, new_n978_, new_n941_ );
nand g0637 ( new_n980_, new_n929_, new_n979_ );
nor g0638 ( new_n981_, new_n980_, new_n928_ );
not g0639 ( new_n982_, new_n981_ );
nand g0640 ( new_n983_, new_n982_, keyIn_0_222 );
not g0641 ( new_n984_, keyIn_0_222 );
nand g0642 ( new_n985_, new_n981_, new_n984_ );
nand g0643 ( N850, new_n983_, new_n985_ );
not g0644 ( new_n987_, keyIn_0_219 );
not g0645 ( new_n988_, N219 );
not g0646 ( new_n989_, keyIn_0_100 );
not g0647 ( new_n990_, keyIn_0_82 );
nand g0648 ( new_n991_, new_n756_, N143 );
nor g0649 ( new_n992_, new_n991_, new_n755_ );
nor g0650 ( new_n993_, new_n992_, new_n990_ );
nand g0651 ( new_n994_, new_n992_, new_n990_ );
nor g0652 ( new_n995_, new_n829_, new_n434_ );
nand g0653 ( new_n996_, new_n995_, keyIn_0_83 );
not g0654 ( new_n997_, keyIn_0_83 );
not g0655 ( new_n998_, new_n995_ );
nand g0656 ( new_n999_, new_n998_, new_n997_ );
nand g0657 ( new_n1000_, new_n999_, new_n996_ );
nand g0658 ( new_n1001_, new_n1000_, new_n994_ );
nor g0659 ( new_n1002_, new_n1001_, new_n993_ );
not g0660 ( new_n1003_, new_n1002_ );
nor g0661 ( new_n1004_, new_n1003_, new_n989_ );
nor g0662 ( new_n1005_, new_n1002_, keyIn_0_100 );
nor g0663 ( new_n1006_, new_n1004_, new_n1005_ );
not g0664 ( new_n1007_, keyIn_0_64 );
nor g0665 ( new_n1008_, new_n860_, new_n1007_ );
nor g0666 ( new_n1009_, new_n862_, keyIn_0_64 );
nor g0667 ( new_n1010_, new_n1009_, new_n1008_ );
nor g0668 ( new_n1011_, new_n1006_, new_n1010_ );
not g0669 ( new_n1012_, new_n1011_ );
nand g0670 ( new_n1013_, new_n1012_, keyIn_0_111 );
not g0671 ( new_n1014_, new_n1013_ );
nor g0672 ( new_n1015_, new_n1012_, keyIn_0_111 );
nor g0673 ( new_n1016_, new_n1014_, new_n1015_ );
nor g0674 ( new_n1017_, new_n1016_, new_n637_ );
not g0675 ( new_n1018_, new_n1017_ );
nor g0676 ( new_n1019_, new_n1018_, keyIn_0_130 );
nand g0677 ( new_n1020_, new_n1018_, keyIn_0_130 );
not g0678 ( new_n1021_, new_n1020_ );
nor g0679 ( new_n1022_, new_n1021_, new_n1019_ );
not g0680 ( new_n1023_, new_n1016_ );
nor g0681 ( new_n1024_, new_n1023_, N183 );
not g0682 ( new_n1025_, new_n1024_ );
nor g0683 ( new_n1026_, new_n1025_, keyIn_0_131 );
nand g0684 ( new_n1027_, new_n1025_, keyIn_0_131 );
not g0685 ( new_n1028_, new_n1027_ );
nor g0686 ( new_n1029_, new_n1028_, new_n1026_ );
not g0687 ( new_n1030_, new_n1029_ );
nor g0688 ( new_n1031_, new_n1030_, new_n1022_ );
not g0689 ( new_n1032_, new_n1031_ );
nor g0690 ( new_n1033_, new_n1032_, keyIn_0_154 );
nand g0691 ( new_n1034_, new_n1032_, keyIn_0_154 );
not g0692 ( new_n1035_, new_n1034_ );
nor g0693 ( new_n1036_, new_n1035_, new_n1033_ );
not g0694 ( new_n1037_, keyIn_0_187 );
not g0695 ( new_n1038_, keyIn_0_159 );
not g0696 ( new_n1039_, keyIn_0_113 );
not g0697 ( new_n1040_, keyIn_0_102 );
nand g0698 ( new_n1041_, new_n756_, N149 );
nor g0699 ( new_n1042_, new_n1041_, new_n755_ );
nor g0700 ( new_n1043_, new_n1042_, keyIn_0_86 );
not g0701 ( new_n1044_, new_n1043_ );
nand g0702 ( new_n1045_, new_n1042_, keyIn_0_86 );
nand g0703 ( new_n1046_, new_n1044_, new_n1045_ );
nand g0704 ( new_n1047_, new_n823_, N121 );
not g0705 ( new_n1048_, new_n1047_ );
nand g0706 ( new_n1049_, new_n1048_, keyIn_0_87 );
not g0707 ( new_n1050_, keyIn_0_87 );
nand g0708 ( new_n1051_, new_n1047_, new_n1050_ );
nand g0709 ( new_n1052_, new_n1049_, new_n1051_ );
nand g0710 ( new_n1053_, new_n1046_, new_n1052_ );
nor g0711 ( new_n1054_, new_n1053_, new_n1040_ );
not g0712 ( new_n1055_, new_n1054_ );
nand g0713 ( new_n1056_, new_n1053_, new_n1040_ );
nor g0714 ( new_n1057_, new_n860_, keyIn_0_66 );
not g0715 ( new_n1058_, keyIn_0_66 );
nor g0716 ( new_n1059_, new_n862_, new_n1058_ );
nor g0717 ( new_n1060_, new_n1059_, new_n1057_ );
nand g0718 ( new_n1061_, new_n1056_, new_n1060_ );
not g0719 ( new_n1062_, new_n1061_ );
nand g0720 ( new_n1063_, new_n1062_, new_n1055_ );
nand g0721 ( new_n1064_, new_n1063_, new_n1039_ );
nor g0722 ( new_n1065_, new_n1061_, new_n1054_ );
nand g0723 ( new_n1066_, new_n1065_, keyIn_0_113 );
nand g0724 ( new_n1067_, new_n1064_, new_n1066_ );
nand g0725 ( new_n1068_, new_n1067_, N195 );
nand g0726 ( new_n1069_, new_n1068_, keyIn_0_135 );
nor g0727 ( new_n1070_, new_n1068_, keyIn_0_135 );
not g0728 ( new_n1071_, new_n1070_ );
nand g0729 ( new_n1072_, new_n1071_, new_n1069_ );
nand g0730 ( new_n1073_, new_n1072_, new_n1038_ );
not g0731 ( new_n1074_, new_n1069_ );
nor g0732 ( new_n1075_, new_n1074_, new_n1070_ );
nand g0733 ( new_n1076_, new_n1075_, keyIn_0_159 );
nand g0734 ( new_n1077_, new_n1076_, new_n1073_ );
not g0735 ( new_n1078_, keyIn_0_134 );
nand g0736 ( new_n1079_, new_n756_, N146 );
not g0737 ( new_n1080_, new_n1079_ );
nand g0738 ( new_n1081_, new_n1080_, new_n760_ );
nand g0739 ( new_n1082_, new_n1081_, keyIn_0_84 );
not g0740 ( new_n1083_, keyIn_0_84 );
nor g0741 ( new_n1084_, new_n1079_, new_n755_ );
nand g0742 ( new_n1085_, new_n1084_, new_n1083_ );
nand g0743 ( new_n1086_, new_n1082_, new_n1085_ );
not g0744 ( new_n1087_, keyIn_0_85 );
nand g0745 ( new_n1088_, new_n823_, N116 );
nand g0746 ( new_n1089_, new_n1088_, new_n1087_ );
nor g0747 ( new_n1090_, new_n829_, new_n436_ );
nand g0748 ( new_n1091_, new_n1090_, keyIn_0_85 );
nand g0749 ( new_n1092_, new_n1089_, new_n1091_ );
nand g0750 ( new_n1093_, new_n1086_, new_n1092_ );
nor g0751 ( new_n1094_, new_n1093_, keyIn_0_101 );
nand g0752 ( new_n1095_, new_n862_, keyIn_0_65 );
not g0753 ( new_n1096_, keyIn_0_65 );
nand g0754 ( new_n1097_, new_n860_, new_n1096_ );
nand g0755 ( new_n1098_, new_n1095_, new_n1097_ );
nand g0756 ( new_n1099_, new_n1093_, keyIn_0_101 );
nand g0757 ( new_n1100_, new_n1099_, new_n1098_ );
nor g0758 ( new_n1101_, new_n1100_, new_n1094_ );
nand g0759 ( new_n1102_, new_n1101_, keyIn_0_112 );
not g0760 ( new_n1103_, keyIn_0_112 );
not g0761 ( new_n1104_, new_n1094_ );
not g0762 ( new_n1105_, new_n1100_ );
nand g0763 ( new_n1106_, new_n1105_, new_n1104_ );
nand g0764 ( new_n1107_, new_n1106_, new_n1103_ );
nand g0765 ( new_n1108_, new_n1107_, new_n1102_ );
nor g0766 ( new_n1109_, new_n1108_, N189 );
nor g0767 ( new_n1110_, new_n1109_, new_n1078_ );
nand g0768 ( new_n1111_, new_n1109_, new_n1078_ );
not g0769 ( new_n1112_, new_n1111_ );
nor g0770 ( new_n1113_, new_n1112_, new_n1110_ );
not g0771 ( new_n1114_, new_n1113_ );
nand g0772 ( new_n1115_, new_n1077_, new_n1114_ );
nand g0773 ( new_n1116_, new_n1115_, new_n1037_ );
not g0774 ( new_n1117_, new_n1115_ );
nand g0775 ( new_n1118_, new_n1117_, keyIn_0_187 );
nand g0776 ( new_n1119_, new_n1118_, new_n1116_ );
not g0777 ( new_n1120_, keyIn_0_188 );
nor g0778 ( new_n1121_, new_n1067_, N195 );
nor g0779 ( new_n1122_, new_n1121_, keyIn_0_136 );
nand g0780 ( new_n1123_, new_n1121_, keyIn_0_136 );
not g0781 ( new_n1124_, new_n1123_ );
nor g0782 ( new_n1125_, new_n1124_, new_n1122_ );
nand g0783 ( new_n1126_, new_n937_, new_n1125_ );
nor g0784 ( new_n1127_, new_n1126_, new_n1113_ );
nor g0785 ( new_n1128_, new_n1127_, new_n1120_ );
not g0786 ( new_n1129_, new_n1128_ );
nand g0787 ( new_n1130_, new_n1129_, new_n1119_ );
nand g0788 ( new_n1131_, new_n1127_, new_n1120_ );
not g0789 ( new_n1132_, new_n1122_ );
nand g0790 ( new_n1133_, new_n1132_, new_n1123_ );
nand g0791 ( new_n1134_, new_n887_, new_n883_ );
nand g0792 ( new_n1135_, new_n881_, keyIn_0_138 );
nand g0793 ( new_n1136_, new_n1134_, new_n1135_ );
nand g0794 ( new_n1137_, new_n1136_, N261 );
nor g0795 ( new_n1138_, new_n1133_, new_n1137_ );
nand g0796 ( new_n1139_, new_n1138_, new_n1114_ );
nand g0797 ( new_n1140_, new_n1139_, keyIn_0_167 );
not g0798 ( new_n1141_, new_n1140_ );
not g0799 ( new_n1142_, keyIn_0_156 );
not g0800 ( new_n1143_, keyIn_0_133 );
nand g0801 ( new_n1144_, new_n1108_, N189 );
nand g0802 ( new_n1145_, new_n1144_, new_n1143_ );
not g0803 ( new_n1146_, new_n1144_ );
nand g0804 ( new_n1147_, new_n1146_, keyIn_0_133 );
nand g0805 ( new_n1148_, new_n1147_, new_n1145_ );
nand g0806 ( new_n1149_, new_n1148_, new_n1142_ );
not g0807 ( new_n1150_, new_n1145_ );
nor g0808 ( new_n1151_, new_n1144_, new_n1143_ );
nor g0809 ( new_n1152_, new_n1150_, new_n1151_ );
nand g0810 ( new_n1153_, new_n1152_, keyIn_0_156 );
nand g0811 ( new_n1154_, new_n1153_, new_n1149_ );
nand g0812 ( new_n1155_, new_n1154_, keyIn_0_177 );
not g0813 ( new_n1156_, keyIn_0_177 );
nor g0814 ( new_n1157_, new_n1152_, keyIn_0_156 );
nor g0815 ( new_n1158_, new_n1148_, new_n1142_ );
nor g0816 ( new_n1159_, new_n1157_, new_n1158_ );
nand g0817 ( new_n1160_, new_n1159_, new_n1156_ );
nand g0818 ( new_n1161_, new_n1160_, new_n1155_ );
not g0819 ( new_n1162_, keyIn_0_167 );
nor g0820 ( new_n1163_, new_n889_, new_n909_ );
nand g0821 ( new_n1164_, new_n1163_, new_n1125_ );
nor g0822 ( new_n1165_, new_n1164_, new_n1113_ );
nand g0823 ( new_n1166_, new_n1165_, new_n1162_ );
nand g0824 ( new_n1167_, new_n1166_, new_n1161_ );
nor g0825 ( new_n1168_, new_n1167_, new_n1141_ );
nand g0826 ( new_n1169_, new_n1168_, new_n1131_ );
nor g0827 ( new_n1170_, new_n1169_, new_n1130_ );
nor g0828 ( new_n1171_, new_n1170_, keyIn_0_196 );
not g0829 ( new_n1172_, new_n1116_ );
nor g0830 ( new_n1173_, new_n1115_, new_n1037_ );
nor g0831 ( new_n1174_, new_n1172_, new_n1173_ );
nor g0832 ( new_n1175_, new_n1174_, new_n1128_ );
nand g0833 ( new_n1176_, new_n1175_, keyIn_0_196 );
nor g0834 ( new_n1177_, new_n1176_, new_n1169_ );
nor g0835 ( new_n1178_, new_n1171_, new_n1177_ );
nor g0836 ( new_n1179_, new_n1178_, new_n1036_ );
not g0837 ( new_n1180_, new_n1179_ );
nand g0838 ( new_n1181_, new_n1180_, keyIn_0_204 );
not g0839 ( new_n1182_, keyIn_0_204 );
nand g0840 ( new_n1183_, new_n1179_, new_n1182_ );
nand g0841 ( new_n1184_, new_n1181_, new_n1183_ );
not g0842 ( new_n1185_, new_n1036_ );
not g0843 ( new_n1186_, keyIn_0_196 );
not g0844 ( new_n1187_, new_n1131_ );
nor g0845 ( new_n1188_, new_n1159_, new_n1156_ );
nor g0846 ( new_n1189_, new_n1154_, keyIn_0_177 );
nor g0847 ( new_n1190_, new_n1188_, new_n1189_ );
nor g0848 ( new_n1191_, new_n1139_, keyIn_0_167 );
nor g0849 ( new_n1192_, new_n1190_, new_n1191_ );
nand g0850 ( new_n1193_, new_n1192_, new_n1140_ );
nor g0851 ( new_n1194_, new_n1193_, new_n1187_ );
nand g0852 ( new_n1195_, new_n1194_, new_n1175_ );
nand g0853 ( new_n1196_, new_n1195_, new_n1186_ );
nor g0854 ( new_n1197_, new_n1130_, new_n1186_ );
nand g0855 ( new_n1198_, new_n1197_, new_n1194_ );
nand g0856 ( new_n1199_, new_n1196_, new_n1198_ );
nor g0857 ( new_n1200_, new_n1185_, new_n1199_ );
nand g0858 ( new_n1201_, new_n1200_, keyIn_0_205 );
not g0859 ( new_n1202_, keyIn_0_205 );
not g0860 ( new_n1203_, new_n1200_ );
nand g0861 ( new_n1204_, new_n1203_, new_n1202_ );
nand g0862 ( new_n1205_, new_n1204_, new_n1201_ );
nand g0863 ( new_n1206_, new_n1205_, new_n1184_ );
nand g0864 ( new_n1207_, new_n1206_, keyIn_0_213 );
not g0865 ( new_n1208_, new_n1207_ );
nor g0866 ( new_n1209_, new_n1206_, keyIn_0_213 );
nor g0867 ( new_n1210_, new_n1208_, new_n1209_ );
nor g0868 ( new_n1211_, new_n1210_, new_n988_ );
nor g0869 ( new_n1212_, new_n1211_, new_n987_ );
nand g0870 ( new_n1213_, new_n1211_, new_n987_ );
not g0871 ( new_n1214_, new_n1213_ );
nor g0872 ( new_n1215_, new_n1214_, new_n1212_ );
nand g0873 ( new_n1216_, N106, N210 );
not g0874 ( new_n1217_, new_n1216_ );
nor g0875 ( new_n1218_, new_n1215_, new_n1217_ );
not g0876 ( new_n1219_, new_n1218_ );
nand g0877 ( new_n1220_, new_n1219_, keyIn_0_230 );
nor g0878 ( new_n1221_, new_n1219_, keyIn_0_230 );
not g0879 ( new_n1222_, keyIn_0_197 );
not g0880 ( new_n1223_, N228 );
nor g0881 ( new_n1224_, new_n1185_, new_n1223_ );
not g0882 ( new_n1225_, new_n1224_ );
nor g0883 ( new_n1226_, new_n1225_, keyIn_0_175 );
nand g0884 ( new_n1227_, new_n1225_, keyIn_0_175 );
not g0885 ( new_n1228_, new_n1227_ );
nor g0886 ( new_n1229_, new_n1228_, new_n1226_ );
not g0887 ( new_n1230_, N237 );
not g0888 ( new_n1231_, keyIn_0_153 );
not g0889 ( new_n1232_, new_n1022_ );
nor g0890 ( new_n1233_, new_n1232_, new_n1231_ );
nor g0891 ( new_n1234_, new_n1022_, keyIn_0_153 );
nor g0892 ( new_n1235_, new_n1233_, new_n1234_ );
nor g0893 ( new_n1236_, new_n1235_, new_n1230_ );
not g0894 ( new_n1237_, new_n1236_ );
nand g0895 ( new_n1238_, new_n1237_, keyIn_0_176 );
not g0896 ( new_n1239_, new_n1238_ );
nor g0897 ( new_n1240_, new_n1237_, keyIn_0_176 );
nor g0898 ( new_n1241_, new_n1239_, new_n1240_ );
nor g0899 ( new_n1242_, new_n1229_, new_n1241_ );
not g0900 ( new_n1243_, new_n1242_ );
nand g0901 ( new_n1244_, new_n1243_, new_n1222_ );
nor g0902 ( new_n1245_, new_n1243_, new_n1222_ );
not g0903 ( new_n1246_, keyIn_0_155 );
not g0904 ( new_n1247_, N246 );
nor g0905 ( new_n1248_, new_n1016_, new_n1247_ );
nor g0906 ( new_n1249_, new_n1248_, keyIn_0_132 );
not g0907 ( new_n1250_, new_n973_ );
nor g0908 ( new_n1251_, new_n1250_, new_n637_ );
nand g0909 ( new_n1252_, new_n1248_, keyIn_0_132 );
not g0910 ( new_n1253_, new_n1252_ );
nor g0911 ( new_n1254_, new_n1253_, new_n1251_ );
not g0912 ( new_n1255_, new_n1254_ );
nor g0913 ( new_n1256_, new_n1255_, new_n1249_ );
nor g0914 ( new_n1257_, new_n1256_, new_n1246_ );
nand g0915 ( new_n1258_, new_n1256_, new_n1246_ );
not g0916 ( new_n1259_, new_n1258_ );
nor g0917 ( new_n1260_, new_n1259_, new_n1257_ );
not g0918 ( new_n1261_, new_n1260_ );
nor g0919 ( new_n1262_, new_n1245_, new_n1261_ );
nand g0920 ( new_n1263_, new_n1262_, new_n1244_ );
nor g0921 ( new_n1264_, new_n1221_, new_n1263_ );
nand g0922 ( new_n1265_, new_n1264_, new_n1220_ );
not g0923 ( new_n1266_, new_n1265_ );
nand g0924 ( new_n1267_, new_n1266_, keyIn_0_240 );
not g0925 ( new_n1268_, keyIn_0_240 );
nand g0926 ( new_n1269_, new_n1265_, new_n1268_ );
nand g0927 ( N863, new_n1267_, new_n1269_ );
not g0928 ( new_n1271_, keyIn_0_214 );
not g0929 ( new_n1272_, keyIn_0_206 );
nor g0930 ( new_n1273_, new_n1113_, new_n1152_ );
not g0931 ( new_n1274_, new_n1273_ );
nand g0932 ( new_n1275_, new_n1274_, keyIn_0_157 );
not g0933 ( new_n1276_, new_n1275_ );
nor g0934 ( new_n1277_, new_n1274_, keyIn_0_157 );
nor g0935 ( new_n1278_, new_n1276_, new_n1277_ );
not g0936 ( new_n1279_, new_n1278_ );
not g0937 ( new_n1280_, keyIn_0_186 );
nand g0938 ( new_n1281_, new_n1126_, new_n1280_ );
not g0939 ( new_n1282_, new_n1281_ );
nor g0940 ( new_n1283_, new_n1126_, new_n1280_ );
nor g0941 ( new_n1284_, new_n1282_, new_n1283_ );
nor g0942 ( new_n1285_, new_n1077_, keyIn_0_180 );
nor g0943 ( new_n1286_, new_n1164_, keyIn_0_166 );
nor g0944 ( new_n1287_, new_n1285_, new_n1286_ );
not g0945 ( new_n1288_, new_n1287_ );
nand g0946 ( new_n1289_, new_n1077_, keyIn_0_180 );
nand g0947 ( new_n1290_, new_n1164_, keyIn_0_166 );
nand g0948 ( new_n1291_, new_n1289_, new_n1290_ );
nor g0949 ( new_n1292_, new_n1288_, new_n1291_ );
not g0950 ( new_n1293_, new_n1292_ );
nor g0951 ( new_n1294_, new_n1293_, new_n1284_ );
nor g0952 ( new_n1295_, new_n1294_, keyIn_0_198 );
nand g0953 ( new_n1296_, new_n1294_, keyIn_0_198 );
not g0954 ( new_n1297_, new_n1296_ );
nor g0955 ( new_n1298_, new_n1297_, new_n1295_ );
not g0956 ( new_n1299_, new_n1298_ );
nor g0957 ( new_n1300_, new_n1299_, new_n1279_ );
not g0958 ( new_n1301_, new_n1300_ );
nor g0959 ( new_n1302_, new_n1301_, new_n1272_ );
nor g0960 ( new_n1303_, new_n1300_, keyIn_0_206 );
nor g0961 ( new_n1304_, new_n1302_, new_n1303_ );
nor g0962 ( new_n1305_, new_n1298_, new_n1278_ );
not g0963 ( new_n1306_, new_n1305_ );
nand g0964 ( new_n1307_, new_n1306_, keyIn_0_207 );
not g0965 ( new_n1308_, new_n1307_ );
nor g0966 ( new_n1309_, new_n1306_, keyIn_0_207 );
nor g0967 ( new_n1310_, new_n1308_, new_n1309_ );
nor g0968 ( new_n1311_, new_n1304_, new_n1310_ );
not g0969 ( new_n1312_, new_n1311_ );
nand g0970 ( new_n1313_, new_n1312_, new_n1271_ );
not g0971 ( new_n1314_, new_n1313_ );
nor g0972 ( new_n1315_, new_n1312_, new_n1271_ );
nor g0973 ( new_n1316_, new_n1314_, new_n1315_ );
nor g0974 ( new_n1317_, new_n1316_, new_n988_ );
not g0975 ( new_n1318_, new_n1317_ );
nand g0976 ( new_n1319_, new_n1318_, keyIn_0_220 );
not g0977 ( new_n1320_, new_n1319_ );
nor g0978 ( new_n1321_, new_n1318_, keyIn_0_220 );
nor g0979 ( new_n1322_, new_n1320_, new_n1321_ );
nand g0980 ( new_n1323_, N111, N210 );
not g0981 ( new_n1324_, new_n1323_ );
nor g0982 ( new_n1325_, new_n1322_, new_n1324_ );
not g0983 ( new_n1326_, new_n1325_ );
nand g0984 ( new_n1327_, new_n1326_, keyIn_0_231 );
nor g0985 ( new_n1328_, new_n1326_, keyIn_0_231 );
not g0986 ( new_n1329_, keyIn_0_199 );
not g0987 ( new_n1330_, keyIn_0_178 );
nor g0988 ( new_n1331_, new_n1278_, new_n1223_ );
not g0989 ( new_n1332_, new_n1331_ );
nand g0990 ( new_n1333_, new_n1332_, new_n1330_ );
not g0991 ( new_n1334_, new_n1333_ );
nor g0992 ( new_n1335_, new_n1332_, new_n1330_ );
nor g0993 ( new_n1336_, new_n1334_, new_n1335_ );
not g0994 ( new_n1337_, keyIn_0_179 );
nor g0995 ( new_n1338_, new_n1154_, new_n1230_ );
not g0996 ( new_n1339_, new_n1338_ );
nor g0997 ( new_n1340_, new_n1339_, new_n1337_ );
nor g0998 ( new_n1341_, new_n1338_, keyIn_0_179 );
nor g0999 ( new_n1342_, new_n1340_, new_n1341_ );
nor g1000 ( new_n1343_, new_n1336_, new_n1342_ );
not g1001 ( new_n1344_, new_n1343_ );
nor g1002 ( new_n1345_, new_n1344_, new_n1329_ );
nand g1003 ( new_n1346_, new_n1344_, new_n1329_ );
nand g1004 ( new_n1347_, new_n1108_, N246 );
nand g1005 ( new_n1348_, N255, N259 );
nand g1006 ( new_n1349_, new_n1347_, new_n1348_ );
nand g1007 ( new_n1350_, new_n1349_, keyIn_0_158 );
not g1008 ( new_n1351_, new_n1350_ );
nand g1009 ( new_n1352_, new_n973_, N189 );
not g1010 ( new_n1353_, keyIn_0_158 );
not g1011 ( new_n1354_, new_n1349_ );
nand g1012 ( new_n1355_, new_n1354_, new_n1353_ );
nand g1013 ( new_n1356_, new_n1355_, new_n1352_ );
nor g1014 ( new_n1357_, new_n1356_, new_n1351_ );
nand g1015 ( new_n1358_, new_n1346_, new_n1357_ );
nor g1016 ( new_n1359_, new_n1358_, new_n1345_ );
not g1017 ( new_n1360_, new_n1359_ );
nor g1018 ( new_n1361_, new_n1328_, new_n1360_ );
nand g1019 ( new_n1362_, new_n1361_, new_n1327_ );
not g1020 ( new_n1363_, new_n1362_ );
nand g1021 ( new_n1364_, new_n1363_, keyIn_0_241 );
not g1022 ( new_n1365_, keyIn_0_241 );
nand g1023 ( new_n1366_, new_n1362_, new_n1365_ );
nand g1024 ( N864, new_n1364_, new_n1366_ );
not g1025 ( new_n1368_, keyIn_0_232 );
not g1026 ( new_n1369_, keyIn_0_221 );
not g1027 ( new_n1370_, keyIn_0_215 );
not g1028 ( new_n1371_, keyIn_0_209 );
not g1029 ( new_n1372_, keyIn_0_160 );
nor g1030 ( new_n1373_, new_n1133_, new_n1075_ );
not g1031 ( new_n1374_, new_n1373_ );
nor g1032 ( new_n1375_, new_n1374_, new_n1372_ );
nor g1033 ( new_n1376_, new_n1373_, keyIn_0_160 );
nor g1034 ( new_n1377_, new_n1375_, new_n1376_ );
not g1035 ( new_n1378_, keyIn_0_200 );
not g1036 ( new_n1379_, keyIn_0_183 );
not g1037 ( new_n1380_, new_n937_ );
nor g1038 ( new_n1381_, new_n1380_, new_n1379_ );
nor g1039 ( new_n1382_, new_n937_, keyIn_0_183 );
nor g1040 ( new_n1383_, new_n1381_, new_n1382_ );
nand g1041 ( new_n1384_, new_n1137_, keyIn_0_165 );
not g1042 ( new_n1385_, new_n1384_ );
nor g1043 ( new_n1386_, new_n1137_, keyIn_0_165 );
nor g1044 ( new_n1387_, new_n1385_, new_n1386_ );
nor g1045 ( new_n1388_, new_n1383_, new_n1387_ );
not g1046 ( new_n1389_, new_n1388_ );
nand g1047 ( new_n1390_, new_n1389_, new_n1378_ );
not g1048 ( new_n1391_, new_n1390_ );
nor g1049 ( new_n1392_, new_n1389_, new_n1378_ );
nor g1050 ( new_n1393_, new_n1391_, new_n1392_ );
nor g1051 ( new_n1394_, new_n1393_, new_n1377_ );
not g1052 ( new_n1395_, new_n1394_ );
nand g1053 ( new_n1396_, new_n1395_, new_n1371_ );
nand g1054 ( new_n1397_, new_n1394_, keyIn_0_209 );
nand g1055 ( new_n1398_, new_n1396_, new_n1397_ );
nand g1056 ( new_n1399_, new_n1393_, new_n1377_ );
not g1057 ( new_n1400_, new_n1399_ );
nand g1058 ( new_n1401_, new_n1400_, keyIn_0_208 );
not g1059 ( new_n1402_, keyIn_0_208 );
nand g1060 ( new_n1403_, new_n1399_, new_n1402_ );
nand g1061 ( new_n1404_, new_n1401_, new_n1403_ );
nand g1062 ( new_n1405_, new_n1398_, new_n1404_ );
nor g1063 ( new_n1406_, new_n1405_, new_n1370_ );
nand g1064 ( new_n1407_, new_n1405_, new_n1370_ );
nand g1065 ( new_n1408_, new_n1407_, N219 );
nor g1066 ( new_n1409_, new_n1408_, new_n1406_ );
not g1067 ( new_n1410_, new_n1409_ );
nor g1068 ( new_n1411_, new_n1410_, new_n1369_ );
nor g1069 ( new_n1412_, new_n1409_, keyIn_0_221 );
nor g1070 ( new_n1413_, new_n1411_, new_n1412_ );
nand g1071 ( new_n1414_, N116, N210 );
not g1072 ( new_n1415_, new_n1414_ );
nor g1073 ( new_n1416_, new_n1413_, new_n1415_ );
not g1074 ( new_n1417_, new_n1416_ );
nor g1075 ( new_n1418_, new_n1417_, new_n1368_ );
nand g1076 ( new_n1419_, new_n1417_, new_n1368_ );
not g1077 ( new_n1420_, keyIn_0_181 );
nor g1078 ( new_n1421_, new_n1377_, new_n1223_ );
not g1079 ( new_n1422_, new_n1421_ );
nand g1080 ( new_n1423_, new_n1422_, new_n1420_ );
not g1081 ( new_n1424_, new_n1423_ );
nor g1082 ( new_n1425_, new_n1422_, new_n1420_ );
nor g1083 ( new_n1426_, new_n1424_, new_n1425_ );
not g1084 ( new_n1427_, keyIn_0_182 );
nor g1085 ( new_n1428_, new_n1075_, keyIn_0_159 );
nor g1086 ( new_n1429_, new_n1072_, new_n1038_ );
nor g1087 ( new_n1430_, new_n1428_, new_n1429_ );
nor g1088 ( new_n1431_, new_n1430_, new_n1230_ );
not g1089 ( new_n1432_, new_n1431_ );
nand g1090 ( new_n1433_, new_n1432_, new_n1427_ );
not g1091 ( new_n1434_, new_n1433_ );
nor g1092 ( new_n1435_, new_n1432_, new_n1427_ );
nor g1093 ( new_n1436_, new_n1434_, new_n1435_ );
nor g1094 ( new_n1437_, new_n1426_, new_n1436_ );
not g1095 ( new_n1438_, new_n1437_ );
nor g1096 ( new_n1439_, new_n1438_, keyIn_0_201 );
not g1097 ( new_n1440_, keyIn_0_201 );
nor g1098 ( new_n1441_, new_n1437_, new_n1440_ );
nor g1099 ( new_n1442_, new_n1439_, new_n1441_ );
not g1100 ( new_n1443_, keyIn_0_161 );
nand g1101 ( new_n1444_, new_n1067_, N246 );
nand g1102 ( new_n1445_, N255, N260 );
nand g1103 ( new_n1446_, new_n1444_, new_n1445_ );
not g1104 ( new_n1447_, new_n1446_ );
nand g1105 ( new_n1448_, new_n1447_, new_n1443_ );
nand g1106 ( new_n1449_, new_n973_, N195 );
nand g1107 ( new_n1450_, new_n1446_, keyIn_0_161 );
nand g1108 ( new_n1451_, new_n1450_, new_n1449_ );
not g1109 ( new_n1452_, new_n1451_ );
nand g1110 ( new_n1453_, new_n1452_, new_n1448_ );
nor g1111 ( new_n1454_, new_n1442_, new_n1453_ );
nand g1112 ( new_n1455_, new_n1419_, new_n1454_ );
nor g1113 ( new_n1456_, new_n1455_, new_n1418_ );
nand g1114 ( new_n1457_, new_n1456_, keyIn_0_242 );
not g1115 ( new_n1458_, keyIn_0_242 );
not g1116 ( new_n1459_, new_n1456_ );
nand g1117 ( new_n1460_, new_n1459_, new_n1458_ );
nand g1118 ( N865, new_n1460_, new_n1457_ );
not g1119 ( new_n1462_, keyIn_0_248 );
not g1120 ( new_n1463_, keyIn_0_225 );
not g1121 ( new_n1464_, keyIn_0_122 );
not g1122 ( new_n1465_, keyIn_0_97 );
not g1123 ( new_n1466_, keyIn_0_76 );
nand g1124 ( new_n1467_, new_n823_, N96 );
nor g1125 ( new_n1468_, new_n1467_, new_n1466_ );
nand g1126 ( new_n1469_, new_n1467_, new_n1466_ );
not g1127 ( new_n1470_, new_n1469_ );
nor g1128 ( new_n1471_, new_n1470_, new_n1468_ );
nand g1129 ( new_n1472_, N51, N138 );
not g1130 ( new_n1473_, new_n1472_ );
nor g1131 ( new_n1474_, new_n1471_, new_n1473_ );
not g1132 ( new_n1475_, new_n1474_ );
nand g1133 ( new_n1476_, new_n1475_, new_n1465_ );
not g1134 ( new_n1477_, new_n1476_ );
nor g1135 ( new_n1478_, new_n1475_, new_n1465_ );
nor g1136 ( new_n1479_, new_n1477_, new_n1478_ );
not g1137 ( new_n1480_, keyIn_0_77 );
not g1138 ( new_n1481_, keyIn_0_57 );
not g1139 ( new_n1482_, keyIn_0_44 );
nor g1140 ( new_n1483_, new_n837_, new_n746_ );
not g1141 ( new_n1484_, new_n1483_ );
nor g1142 ( new_n1485_, new_n1484_, new_n1482_ );
nor g1143 ( new_n1486_, new_n1483_, keyIn_0_44 );
nor g1144 ( new_n1487_, new_n1485_, new_n1486_ );
not g1145 ( new_n1488_, new_n1487_ );
nand g1146 ( new_n1489_, new_n1488_, N146 );
nand g1147 ( new_n1490_, new_n1489_, new_n1481_ );
not g1148 ( new_n1491_, new_n1490_ );
nor g1149 ( new_n1492_, new_n1489_, new_n1481_ );
nor g1150 ( new_n1493_, new_n1491_, new_n1492_ );
not g1151 ( new_n1494_, keyIn_0_58 );
nor g1152 ( new_n1495_, new_n750_, new_n845_ );
not g1153 ( new_n1496_, new_n1495_ );
nor g1154 ( new_n1497_, new_n1496_, keyIn_0_45 );
nand g1155 ( new_n1498_, new_n1496_, keyIn_0_45 );
nand g1156 ( new_n1499_, new_n1498_, new_n853_ );
nor g1157 ( new_n1500_, new_n1499_, new_n1497_ );
not g1158 ( new_n1501_, new_n1500_ );
nor g1159 ( new_n1502_, new_n1501_, new_n1494_ );
nor g1160 ( new_n1503_, new_n1500_, keyIn_0_58 );
nor g1161 ( new_n1504_, new_n1502_, new_n1503_ );
nor g1162 ( new_n1505_, new_n1493_, new_n1504_ );
not g1163 ( new_n1506_, new_n1505_ );
nor g1164 ( new_n1507_, new_n1506_, new_n1480_ );
nor g1165 ( new_n1508_, new_n1505_, keyIn_0_77 );
nor g1166 ( new_n1509_, new_n1507_, new_n1508_ );
nor g1167 ( new_n1510_, new_n1479_, new_n1509_ );
not g1168 ( new_n1511_, new_n1510_ );
nor g1169 ( new_n1512_, new_n1511_, keyIn_0_108 );
nand g1170 ( new_n1513_, new_n1511_, keyIn_0_108 );
not g1171 ( new_n1514_, new_n1513_ );
nor g1172 ( new_n1515_, new_n1514_, new_n1512_ );
not g1173 ( new_n1516_, new_n1515_ );
nor g1174 ( new_n1517_, new_n1516_, N165 );
not g1175 ( new_n1518_, new_n1517_ );
nor g1176 ( new_n1519_, new_n1518_, new_n1464_ );
nor g1177 ( new_n1520_, new_n1517_, keyIn_0_122 );
nor g1178 ( new_n1521_, new_n1519_, new_n1520_ );
not g1179 ( new_n1522_, new_n1521_ );
not g1180 ( new_n1523_, keyIn_0_109 );
not g1181 ( new_n1524_, keyIn_0_79 );
nand g1182 ( new_n1525_, new_n1488_, N149 );
nand g1183 ( new_n1526_, new_n1525_, keyIn_0_59 );
not g1184 ( new_n1527_, new_n1526_ );
nor g1185 ( new_n1528_, new_n1525_, keyIn_0_59 );
nor g1186 ( new_n1529_, new_n1527_, new_n1528_ );
not g1187 ( new_n1530_, keyIn_0_60 );
nor g1188 ( new_n1531_, new_n1501_, new_n1530_ );
nor g1189 ( new_n1532_, new_n1500_, keyIn_0_60 );
nor g1190 ( new_n1533_, new_n1531_, new_n1532_ );
nor g1191 ( new_n1534_, new_n1529_, new_n1533_ );
not g1192 ( new_n1535_, new_n1534_ );
nor g1193 ( new_n1536_, new_n1535_, new_n1524_ );
nor g1194 ( new_n1537_, new_n1534_, keyIn_0_79 );
nor g1195 ( new_n1538_, new_n1536_, new_n1537_ );
not g1196 ( new_n1539_, keyIn_0_78 );
nor g1197 ( new_n1540_, new_n829_, new_n500_ );
not g1198 ( new_n1541_, new_n1540_ );
nor g1199 ( new_n1542_, new_n1541_, new_n1539_ );
nor g1200 ( new_n1543_, new_n1540_, keyIn_0_78 );
nor g1201 ( new_n1544_, new_n1542_, new_n1543_ );
nand g1202 ( new_n1545_, N17, N138 );
not g1203 ( new_n1546_, new_n1545_ );
nor g1204 ( new_n1547_, new_n1544_, new_n1546_ );
not g1205 ( new_n1548_, new_n1547_ );
nand g1206 ( new_n1549_, new_n1548_, keyIn_0_98 );
not g1207 ( new_n1550_, new_n1549_ );
nor g1208 ( new_n1551_, new_n1548_, keyIn_0_98 );
nor g1209 ( new_n1552_, new_n1550_, new_n1551_ );
nor g1210 ( new_n1553_, new_n1552_, new_n1538_ );
not g1211 ( new_n1554_, new_n1553_ );
nor g1212 ( new_n1555_, new_n1554_, new_n1523_ );
nor g1213 ( new_n1556_, new_n1553_, keyIn_0_109 );
nor g1214 ( new_n1557_, new_n1555_, new_n1556_ );
not g1215 ( new_n1558_, new_n1557_ );
nor g1216 ( new_n1559_, new_n1558_, N171 );
not g1217 ( new_n1560_, new_n1559_ );
nor g1218 ( new_n1561_, new_n1560_, keyIn_0_125 );
nand g1219 ( new_n1562_, new_n1560_, keyIn_0_125 );
not g1220 ( new_n1563_, new_n1562_ );
nor g1221 ( new_n1564_, new_n1563_, new_n1561_ );
not g1222 ( new_n1565_, new_n1564_ );
nor g1223 ( new_n1566_, new_n1565_, new_n1522_ );
not g1224 ( new_n1567_, new_n1566_ );
nand g1225 ( new_n1568_, new_n1178_, new_n1029_ );
nand g1226 ( new_n1569_, new_n1568_, keyIn_0_211 );
not g1227 ( new_n1570_, keyIn_0_211 );
nor g1228 ( new_n1571_, new_n1199_, new_n1030_ );
nand g1229 ( new_n1572_, new_n1571_, new_n1570_ );
nand g1230 ( new_n1573_, new_n1572_, new_n1569_ );
not g1231 ( new_n1574_, keyIn_0_174 );
nor g1232 ( new_n1575_, new_n1235_, new_n1574_ );
not g1233 ( new_n1576_, new_n1235_ );
nor g1234 ( new_n1577_, new_n1576_, keyIn_0_174 );
nor g1235 ( new_n1578_, new_n1577_, new_n1575_ );
nand g1236 ( new_n1579_, new_n1573_, new_n1578_ );
nand g1237 ( new_n1580_, new_n1579_, keyIn_0_212 );
not g1238 ( new_n1581_, keyIn_0_212 );
not g1239 ( new_n1582_, new_n1579_ );
nand g1240 ( new_n1583_, new_n1582_, new_n1581_ );
nand g1241 ( new_n1584_, new_n1583_, new_n1580_ );
not g1242 ( new_n1585_, keyIn_0_128 );
not g1243 ( new_n1586_, keyIn_0_110 );
nor g1244 ( new_n1587_, new_n829_, new_n502_ );
not g1245 ( new_n1588_, new_n1587_ );
nor g1246 ( new_n1589_, new_n1588_, keyIn_0_80 );
nand g1247 ( new_n1590_, N138, N152 );
nand g1248 ( new_n1591_, new_n1588_, keyIn_0_80 );
nand g1249 ( new_n1592_, new_n1591_, new_n1590_ );
nor g1250 ( new_n1593_, new_n1592_, new_n1589_ );
nor g1251 ( new_n1594_, new_n1593_, keyIn_0_99 );
nand g1252 ( new_n1595_, new_n1593_, keyIn_0_99 );
not g1253 ( new_n1596_, new_n1595_ );
nand g1254 ( new_n1597_, new_n1488_, N153 );
nand g1255 ( new_n1598_, new_n1597_, keyIn_0_61 );
not g1256 ( new_n1599_, new_n1598_ );
nor g1257 ( new_n1600_, new_n1597_, keyIn_0_61 );
nor g1258 ( new_n1601_, new_n1599_, new_n1600_ );
not g1259 ( new_n1602_, keyIn_0_62 );
nor g1260 ( new_n1603_, new_n1501_, new_n1602_ );
nor g1261 ( new_n1604_, new_n1500_, keyIn_0_62 );
nor g1262 ( new_n1605_, new_n1603_, new_n1604_ );
nor g1263 ( new_n1606_, new_n1601_, new_n1605_ );
not g1264 ( new_n1607_, new_n1606_ );
nor g1265 ( new_n1608_, new_n1607_, keyIn_0_81 );
nand g1266 ( new_n1609_, new_n1607_, keyIn_0_81 );
not g1267 ( new_n1610_, new_n1609_ );
nor g1268 ( new_n1611_, new_n1610_, new_n1608_ );
nor g1269 ( new_n1612_, new_n1611_, new_n1596_ );
not g1270 ( new_n1613_, new_n1612_ );
nor g1271 ( new_n1614_, new_n1613_, new_n1594_ );
not g1272 ( new_n1615_, new_n1614_ );
nor g1273 ( new_n1616_, new_n1615_, new_n1586_ );
nor g1274 ( new_n1617_, new_n1614_, keyIn_0_110 );
nor g1275 ( new_n1618_, new_n1616_, new_n1617_ );
nor g1276 ( new_n1619_, new_n1618_, N177 );
not g1277 ( new_n1620_, new_n1619_ );
nand g1278 ( new_n1621_, new_n1620_, new_n1585_ );
not g1279 ( new_n1622_, new_n1621_ );
nor g1280 ( new_n1623_, new_n1620_, new_n1585_ );
nor g1281 ( new_n1624_, new_n1622_, new_n1623_ );
not g1282 ( new_n1625_, new_n1624_ );
nand g1283 ( new_n1626_, new_n1584_, new_n1625_ );
nor g1284 ( new_n1627_, new_n1626_, new_n1567_ );
nor g1285 ( new_n1628_, new_n1627_, new_n1463_ );
nand g1286 ( new_n1629_, new_n1627_, new_n1463_ );
not g1287 ( new_n1630_, keyIn_0_190 );
not g1288 ( new_n1631_, keyIn_0_147 );
not g1289 ( new_n1632_, keyIn_0_124 );
nand g1290 ( new_n1633_, new_n1558_, N171 );
nand g1291 ( new_n1634_, new_n1633_, new_n1632_ );
not g1292 ( new_n1635_, new_n1634_ );
nor g1293 ( new_n1636_, new_n1633_, new_n1632_ );
nor g1294 ( new_n1637_, new_n1635_, new_n1636_ );
not g1295 ( new_n1638_, new_n1637_ );
nor g1296 ( new_n1639_, new_n1638_, new_n1631_ );
nor g1297 ( new_n1640_, new_n1637_, keyIn_0_147 );
nor g1298 ( new_n1641_, new_n1639_, new_n1640_ );
not g1299 ( new_n1642_, new_n1641_ );
nor g1300 ( new_n1643_, new_n1642_, new_n1522_ );
not g1301 ( new_n1644_, new_n1643_ );
nor g1302 ( new_n1645_, new_n1644_, new_n1630_ );
not g1303 ( new_n1646_, keyIn_0_144 );
nor g1304 ( new_n1647_, new_n1515_, new_n585_ );
not g1305 ( new_n1648_, new_n1647_ );
nand g1306 ( new_n1649_, new_n1648_, keyIn_0_121 );
not g1307 ( new_n1650_, new_n1649_ );
nor g1308 ( new_n1651_, new_n1648_, keyIn_0_121 );
nor g1309 ( new_n1652_, new_n1650_, new_n1651_ );
not g1310 ( new_n1653_, new_n1652_ );
nor g1311 ( new_n1654_, new_n1653_, new_n1646_ );
nor g1312 ( new_n1655_, new_n1652_, keyIn_0_144 );
nor g1313 ( new_n1656_, new_n1654_, new_n1655_ );
nor g1314 ( new_n1657_, new_n1656_, keyIn_0_168 );
nand g1315 ( new_n1658_, new_n1656_, keyIn_0_168 );
not g1316 ( new_n1659_, new_n1658_ );
nor g1317 ( new_n1660_, new_n1659_, new_n1657_ );
nor g1318 ( new_n1661_, new_n1645_, new_n1660_ );
not g1319 ( new_n1662_, new_n1661_ );
not g1320 ( new_n1663_, keyIn_0_191 );
not g1321 ( new_n1664_, keyIn_0_150 );
not g1322 ( new_n1665_, keyIn_0_127 );
not g1323 ( new_n1666_, N177 );
not g1324 ( new_n1667_, new_n1618_ );
nor g1325 ( new_n1668_, new_n1667_, new_n1666_ );
not g1326 ( new_n1669_, new_n1668_ );
nor g1327 ( new_n1670_, new_n1669_, new_n1665_ );
nor g1328 ( new_n1671_, new_n1668_, keyIn_0_127 );
nor g1329 ( new_n1672_, new_n1670_, new_n1671_ );
not g1330 ( new_n1673_, new_n1672_ );
nor g1331 ( new_n1674_, new_n1673_, new_n1664_ );
nor g1332 ( new_n1675_, new_n1672_, keyIn_0_150 );
nor g1333 ( new_n1676_, new_n1674_, new_n1675_ );
nor g1334 ( new_n1677_, new_n1676_, new_n1567_ );
not g1335 ( new_n1678_, new_n1677_ );
nand g1336 ( new_n1679_, new_n1678_, new_n1663_ );
nor g1337 ( new_n1680_, new_n1643_, keyIn_0_190 );
nor g1338 ( new_n1681_, new_n1678_, new_n1663_ );
nor g1339 ( new_n1682_, new_n1681_, new_n1680_ );
nand g1340 ( new_n1683_, new_n1682_, new_n1679_ );
nor g1341 ( new_n1684_, new_n1683_, new_n1662_ );
nand g1342 ( new_n1685_, new_n1629_, new_n1684_ );
nor g1343 ( new_n1686_, new_n1685_, new_n1628_ );
nor g1344 ( new_n1687_, new_n1686_, keyIn_0_226 );
not g1345 ( new_n1688_, keyIn_0_226 );
not g1346 ( new_n1689_, new_n1628_ );
not g1347 ( new_n1690_, new_n1580_ );
nor g1348 ( new_n1691_, new_n1579_, keyIn_0_212 );
nor g1349 ( new_n1692_, new_n1690_, new_n1691_ );
nor g1350 ( new_n1693_, new_n1692_, new_n1624_ );
nand g1351 ( new_n1694_, new_n1693_, new_n1566_ );
nor g1352 ( new_n1695_, new_n1694_, keyIn_0_225 );
not g1353 ( new_n1696_, new_n1684_ );
nor g1354 ( new_n1697_, new_n1695_, new_n1696_ );
nand g1355 ( new_n1698_, new_n1697_, new_n1689_ );
nor g1356 ( new_n1699_, new_n1698_, new_n1688_ );
nor g1357 ( new_n1700_, new_n1699_, new_n1687_ );
not g1358 ( new_n1701_, keyIn_0_74 );
nand g1359 ( new_n1702_, new_n823_, N91 );
nor g1360 ( new_n1703_, new_n1702_, new_n1701_ );
nand g1361 ( new_n1704_, new_n1702_, new_n1701_ );
not g1362 ( new_n1705_, new_n1704_ );
nor g1363 ( new_n1706_, new_n1705_, new_n1703_ );
nand g1364 ( new_n1707_, N8, N138 );
not g1365 ( new_n1708_, new_n1707_ );
nor g1366 ( new_n1709_, new_n1706_, new_n1708_ );
not g1367 ( new_n1710_, new_n1709_ );
nor g1368 ( new_n1711_, new_n1710_, keyIn_0_96 );
nand g1369 ( new_n1712_, new_n1710_, keyIn_0_96 );
not g1370 ( new_n1713_, keyIn_0_75 );
not g1371 ( new_n1714_, keyIn_0_55 );
nand g1372 ( new_n1715_, new_n1488_, N143 );
nand g1373 ( new_n1716_, new_n1715_, new_n1714_ );
not g1374 ( new_n1717_, new_n1716_ );
nor g1375 ( new_n1718_, new_n1715_, new_n1714_ );
nor g1376 ( new_n1719_, new_n1717_, new_n1718_ );
not g1377 ( new_n1720_, keyIn_0_56 );
nor g1378 ( new_n1721_, new_n1501_, new_n1720_ );
nor g1379 ( new_n1722_, new_n1500_, keyIn_0_56 );
nor g1380 ( new_n1723_, new_n1721_, new_n1722_ );
nor g1381 ( new_n1724_, new_n1719_, new_n1723_ );
not g1382 ( new_n1725_, new_n1724_ );
nand g1383 ( new_n1726_, new_n1725_, new_n1713_ );
nand g1384 ( new_n1727_, new_n1724_, keyIn_0_75 );
nand g1385 ( new_n1728_, new_n1726_, new_n1727_ );
nand g1386 ( new_n1729_, new_n1728_, new_n1712_ );
nor g1387 ( new_n1730_, new_n1729_, new_n1711_ );
not g1388 ( new_n1731_, new_n1730_ );
nor g1389 ( new_n1732_, new_n1731_, keyIn_0_107 );
nand g1390 ( new_n1733_, new_n1731_, keyIn_0_107 );
not g1391 ( new_n1734_, new_n1733_ );
nor g1392 ( new_n1735_, new_n1734_, new_n1732_ );
not g1393 ( new_n1736_, new_n1735_ );
nor g1394 ( new_n1737_, new_n1736_, N159 );
not g1395 ( new_n1738_, new_n1737_ );
nor g1396 ( new_n1739_, new_n1738_, keyIn_0_119 );
nand g1397 ( new_n1740_, new_n1738_, keyIn_0_119 );
not g1398 ( new_n1741_, new_n1740_ );
nor g1399 ( new_n1742_, new_n1741_, new_n1739_ );
not g1400 ( new_n1743_, new_n1742_ );
nor g1401 ( new_n1744_, new_n1700_, new_n1743_ );
not g1402 ( new_n1745_, new_n1744_ );
nand g1403 ( new_n1746_, new_n1745_, keyIn_0_243 );
not g1404 ( new_n1747_, keyIn_0_141 );
nor g1405 ( new_n1748_, new_n1735_, new_n583_ );
not g1406 ( new_n1749_, new_n1748_ );
nand g1407 ( new_n1750_, new_n1749_, keyIn_0_118 );
not g1408 ( new_n1751_, new_n1750_ );
nor g1409 ( new_n1752_, new_n1749_, keyIn_0_118 );
nor g1410 ( new_n1753_, new_n1751_, new_n1752_ );
nor g1411 ( new_n1754_, new_n1753_, new_n1747_ );
not g1412 ( new_n1755_, new_n1753_ );
nor g1413 ( new_n1756_, new_n1755_, keyIn_0_141 );
nor g1414 ( new_n1757_, new_n1756_, new_n1754_ );
not g1415 ( new_n1758_, new_n1757_ );
nor g1416 ( new_n1759_, new_n1745_, keyIn_0_243 );
nor g1417 ( new_n1760_, new_n1759_, new_n1758_ );
nand g1418 ( new_n1761_, new_n1760_, new_n1746_ );
nand g1419 ( new_n1762_, new_n1761_, new_n1462_ );
not g1420 ( new_n1763_, new_n1761_ );
nand g1421 ( new_n1764_, new_n1763_, keyIn_0_248 );
nand g1422 ( N866, new_n1764_, new_n1762_ );
not g1423 ( new_n1766_, keyIn_0_247 );
not g1424 ( new_n1767_, keyIn_0_239 );
nor g1425 ( new_n1768_, new_n1672_, new_n1624_ );
not g1426 ( new_n1769_, new_n1768_ );
nor g1427 ( new_n1770_, new_n1769_, keyIn_0_151 );
nand g1428 ( new_n1771_, new_n1769_, keyIn_0_151 );
not g1429 ( new_n1772_, new_n1771_ );
nor g1430 ( new_n1773_, new_n1772_, new_n1770_ );
not g1431 ( new_n1774_, new_n1773_ );
nor g1432 ( new_n1775_, new_n1584_, new_n1774_ );
not g1433 ( new_n1776_, new_n1775_ );
nand g1434 ( new_n1777_, new_n1776_, keyIn_0_217 );
not g1435 ( new_n1778_, keyIn_0_217 );
nand g1436 ( new_n1779_, new_n1775_, new_n1778_ );
nand g1437 ( new_n1780_, new_n1777_, new_n1779_ );
not g1438 ( new_n1781_, keyIn_0_218 );
nor g1439 ( new_n1782_, new_n1692_, new_n1773_ );
nand g1440 ( new_n1783_, new_n1782_, new_n1781_ );
not g1441 ( new_n1784_, new_n1782_ );
nand g1442 ( new_n1785_, new_n1784_, keyIn_0_218 );
nand g1443 ( new_n1786_, new_n1785_, new_n1783_ );
nand g1444 ( new_n1787_, new_n1786_, new_n1780_ );
nand g1445 ( new_n1788_, new_n1787_, keyIn_0_229 );
nor g1446 ( new_n1789_, new_n1787_, keyIn_0_229 );
nor g1447 ( new_n1790_, new_n1789_, new_n988_ );
nand g1448 ( new_n1791_, new_n1790_, new_n1788_ );
not g1449 ( new_n1792_, new_n1791_ );
nor g1450 ( new_n1793_, new_n1792_, new_n1767_ );
nor g1451 ( new_n1794_, new_n1791_, keyIn_0_239 );
nor g1452 ( new_n1795_, new_n1793_, new_n1794_ );
nand g1453 ( new_n1796_, N101, N210 );
not g1454 ( new_n1797_, new_n1796_ );
nor g1455 ( new_n1798_, new_n1795_, new_n1797_ );
not g1456 ( new_n1799_, new_n1798_ );
nand g1457 ( new_n1800_, new_n1799_, new_n1766_ );
not g1458 ( new_n1801_, new_n1800_ );
nor g1459 ( new_n1802_, new_n1799_, new_n1766_ );
nor g1460 ( new_n1803_, new_n1801_, new_n1802_ );
nor g1461 ( new_n1804_, new_n1773_, new_n1223_ );
not g1462 ( new_n1805_, new_n1804_ );
nand g1463 ( new_n1806_, new_n1805_, keyIn_0_172 );
not g1464 ( new_n1807_, new_n1806_ );
nor g1465 ( new_n1808_, new_n1805_, keyIn_0_172 );
nor g1466 ( new_n1809_, new_n1807_, new_n1808_ );
not g1467 ( new_n1810_, keyIn_0_173 );
nor g1468 ( new_n1811_, new_n1676_, new_n1230_ );
not g1469 ( new_n1812_, new_n1811_ );
nand g1470 ( new_n1813_, new_n1812_, new_n1810_ );
not g1471 ( new_n1814_, new_n1813_ );
nor g1472 ( new_n1815_, new_n1812_, new_n1810_ );
nor g1473 ( new_n1816_, new_n1814_, new_n1815_ );
nor g1474 ( new_n1817_, new_n1809_, new_n1816_ );
not g1475 ( new_n1818_, new_n1817_ );
nand g1476 ( new_n1819_, new_n1818_, keyIn_0_195 );
nor g1477 ( new_n1820_, new_n1667_, new_n1247_ );
not g1478 ( new_n1821_, new_n1820_ );
nor g1479 ( new_n1822_, new_n1821_, keyIn_0_129 );
nor g1480 ( new_n1823_, new_n1250_, new_n1666_ );
nand g1481 ( new_n1824_, new_n1821_, keyIn_0_129 );
not g1482 ( new_n1825_, new_n1824_ );
nor g1483 ( new_n1826_, new_n1825_, new_n1823_ );
not g1484 ( new_n1827_, new_n1826_ );
nor g1485 ( new_n1828_, new_n1827_, new_n1822_ );
not g1486 ( new_n1829_, new_n1828_ );
nor g1487 ( new_n1830_, new_n1829_, keyIn_0_152 );
nand g1488 ( new_n1831_, new_n1829_, keyIn_0_152 );
not g1489 ( new_n1832_, new_n1831_ );
nor g1490 ( new_n1833_, new_n1832_, new_n1830_ );
nor g1491 ( new_n1834_, new_n1818_, keyIn_0_195 );
nor g1492 ( new_n1835_, new_n1834_, new_n1833_ );
nand g1493 ( new_n1836_, new_n1835_, new_n1819_ );
nor g1494 ( new_n1837_, new_n1803_, new_n1836_ );
not g1495 ( new_n1838_, new_n1837_ );
nand g1496 ( new_n1839_, new_n1838_, keyIn_0_249 );
not g1497 ( new_n1840_, keyIn_0_249 );
nand g1498 ( new_n1841_, new_n1837_, new_n1840_ );
nand g1499 ( N874, new_n1839_, new_n1841_ );
not g1500 ( new_n1843_, keyIn_0_244 );
nand g1501 ( new_n1844_, new_n1698_, new_n1688_ );
nand g1502 ( new_n1845_, new_n1686_, keyIn_0_226 );
nand g1503 ( new_n1846_, new_n1844_, new_n1845_ );
not g1504 ( new_n1847_, keyIn_0_142 );
nor g1505 ( new_n1848_, new_n1743_, new_n1753_ );
not g1506 ( new_n1849_, new_n1848_ );
nor g1507 ( new_n1850_, new_n1849_, new_n1847_ );
nor g1508 ( new_n1851_, new_n1848_, keyIn_0_142 );
nor g1509 ( new_n1852_, new_n1850_, new_n1851_ );
not g1510 ( new_n1853_, new_n1852_ );
nand g1511 ( new_n1854_, new_n1846_, new_n1853_ );
nand g1512 ( new_n1855_, new_n1854_, keyIn_0_234 );
not g1513 ( new_n1856_, keyIn_0_234 );
nor g1514 ( new_n1857_, new_n1700_, new_n1852_ );
nand g1515 ( new_n1858_, new_n1857_, new_n1856_ );
nand g1516 ( new_n1859_, new_n1858_, new_n1855_ );
nand g1517 ( new_n1860_, new_n1700_, new_n1852_ );
nand g1518 ( new_n1861_, new_n1860_, keyIn_0_233 );
not g1519 ( new_n1862_, keyIn_0_233 );
nor g1520 ( new_n1863_, new_n1846_, new_n1853_ );
nand g1521 ( new_n1864_, new_n1863_, new_n1862_ );
nand g1522 ( new_n1865_, new_n1861_, new_n1864_ );
nand g1523 ( new_n1866_, new_n1859_, new_n1865_ );
nor g1524 ( new_n1867_, new_n1866_, new_n1843_ );
not g1525 ( new_n1868_, new_n1867_ );
nand g1526 ( new_n1869_, new_n1866_, new_n1843_ );
nand g1527 ( new_n1870_, new_n1869_, N219 );
not g1528 ( new_n1871_, new_n1870_ );
nand g1529 ( new_n1872_, new_n1871_, new_n1868_ );
not g1530 ( new_n1873_, N210 );
nor g1531 ( new_n1874_, new_n857_, new_n1873_ );
not g1532 ( new_n1875_, new_n1874_ );
nand g1533 ( new_n1876_, new_n1872_, new_n1875_ );
nand g1534 ( new_n1877_, new_n1876_, keyIn_0_250 );
not g1535 ( new_n1878_, keyIn_0_250 );
nor g1536 ( new_n1879_, new_n1870_, new_n1867_ );
nor g1537 ( new_n1880_, new_n1879_, new_n1874_ );
nand g1538 ( new_n1881_, new_n1880_, new_n1878_ );
nand g1539 ( new_n1882_, new_n1877_, new_n1881_ );
nand g1540 ( new_n1883_, new_n1853_, N228 );
nand g1541 ( new_n1884_, new_n1758_, N237 );
nand g1542 ( new_n1885_, new_n1883_, new_n1884_ );
nand g1543 ( new_n1886_, new_n1885_, keyIn_0_192 );
not g1544 ( new_n1887_, keyIn_0_120 );
nor g1545 ( new_n1888_, new_n1735_, new_n1247_ );
not g1546 ( new_n1889_, new_n1888_ );
nand g1547 ( new_n1890_, new_n1889_, new_n1887_ );
not g1548 ( new_n1891_, new_n1890_ );
nor g1549 ( new_n1892_, new_n1889_, new_n1887_ );
nor g1550 ( new_n1893_, new_n1891_, new_n1892_ );
nor g1551 ( new_n1894_, new_n1250_, new_n583_ );
nor g1552 ( new_n1895_, new_n1893_, new_n1894_ );
nor g1553 ( new_n1896_, new_n1895_, keyIn_0_143 );
nand g1554 ( new_n1897_, new_n1895_, keyIn_0_143 );
not g1555 ( new_n1898_, new_n1897_ );
nor g1556 ( new_n1899_, new_n1898_, new_n1896_ );
nor g1557 ( new_n1900_, new_n1885_, keyIn_0_192 );
nor g1558 ( new_n1901_, new_n1900_, new_n1899_ );
nand g1559 ( new_n1902_, new_n1901_, new_n1886_ );
not g1560 ( new_n1903_, new_n1902_ );
nand g1561 ( new_n1904_, new_n1882_, new_n1903_ );
nand g1562 ( new_n1905_, new_n1904_, keyIn_0_253 );
not g1563 ( new_n1906_, keyIn_0_253 );
nor g1564 ( new_n1907_, new_n1880_, new_n1878_ );
nor g1565 ( new_n1908_, new_n1876_, keyIn_0_250 );
nor g1566 ( new_n1909_, new_n1908_, new_n1907_ );
nor g1567 ( new_n1910_, new_n1909_, new_n1902_ );
nand g1568 ( new_n1911_, new_n1910_, new_n1906_ );
nand g1569 ( N878, new_n1911_, new_n1905_ );
not g1570 ( new_n1913_, keyIn_0_254 );
not g1571 ( new_n1914_, keyIn_0_251 );
not g1572 ( new_n1915_, keyIn_0_236 );
not g1573 ( new_n1916_, keyIn_0_224 );
nand g1574 ( new_n1917_, new_n1693_, new_n1564_ );
nand g1575 ( new_n1918_, new_n1917_, new_n1916_ );
nor g1576 ( new_n1919_, new_n1626_, new_n1565_ );
nand g1577 ( new_n1920_, new_n1919_, keyIn_0_224 );
nand g1578 ( new_n1921_, new_n1918_, new_n1920_ );
not g1579 ( new_n1922_, keyIn_0_189 );
nor g1580 ( new_n1923_, new_n1676_, new_n1565_ );
not g1581 ( new_n1924_, new_n1923_ );
nor g1582 ( new_n1925_, new_n1924_, new_n1922_ );
nand g1583 ( new_n1926_, new_n1924_, new_n1922_ );
not g1584 ( new_n1927_, new_n1926_ );
not g1585 ( new_n1928_, keyIn_0_169 );
nor g1586 ( new_n1929_, new_n1642_, new_n1928_ );
nor g1587 ( new_n1930_, new_n1641_, keyIn_0_169 );
nor g1588 ( new_n1931_, new_n1929_, new_n1930_ );
nor g1589 ( new_n1932_, new_n1927_, new_n1931_ );
not g1590 ( new_n1933_, new_n1932_ );
nor g1591 ( new_n1934_, new_n1933_, new_n1925_ );
nand g1592 ( new_n1935_, new_n1921_, new_n1934_ );
nand g1593 ( new_n1936_, new_n1935_, keyIn_0_227 );
not g1594 ( new_n1937_, keyIn_0_227 );
nor g1595 ( new_n1938_, new_n1919_, keyIn_0_224 );
nor g1596 ( new_n1939_, new_n1917_, new_n1916_ );
nor g1597 ( new_n1940_, new_n1939_, new_n1938_ );
not g1598 ( new_n1941_, new_n1934_ );
nor g1599 ( new_n1942_, new_n1940_, new_n1941_ );
nand g1600 ( new_n1943_, new_n1942_, new_n1937_ );
nand g1601 ( new_n1944_, new_n1943_, new_n1936_ );
not g1602 ( new_n1945_, keyIn_0_145 );
nor g1603 ( new_n1946_, new_n1522_, new_n1652_ );
not g1604 ( new_n1947_, new_n1946_ );
nor g1605 ( new_n1948_, new_n1947_, new_n1945_ );
nor g1606 ( new_n1949_, new_n1946_, keyIn_0_145 );
nor g1607 ( new_n1950_, new_n1948_, new_n1949_ );
not g1608 ( new_n1951_, new_n1950_ );
nand g1609 ( new_n1952_, new_n1944_, new_n1951_ );
nand g1610 ( new_n1953_, new_n1952_, new_n1915_ );
not g1611 ( new_n1954_, new_n1936_ );
nor g1612 ( new_n1955_, new_n1935_, keyIn_0_227 );
nor g1613 ( new_n1956_, new_n1954_, new_n1955_ );
nor g1614 ( new_n1957_, new_n1956_, new_n1950_ );
nand g1615 ( new_n1958_, new_n1957_, keyIn_0_236 );
nand g1616 ( new_n1959_, new_n1958_, new_n1953_ );
nand g1617 ( new_n1960_, new_n1956_, new_n1950_ );
nand g1618 ( new_n1961_, new_n1960_, keyIn_0_235 );
not g1619 ( new_n1962_, keyIn_0_235 );
nor g1620 ( new_n1963_, new_n1944_, new_n1951_ );
nand g1621 ( new_n1964_, new_n1963_, new_n1962_ );
nand g1622 ( new_n1965_, new_n1961_, new_n1964_ );
nand g1623 ( new_n1966_, new_n1959_, new_n1965_ );
nor g1624 ( new_n1967_, new_n1966_, keyIn_0_245 );
not g1625 ( new_n1968_, new_n1967_ );
nand g1626 ( new_n1969_, new_n1966_, keyIn_0_245 );
nand g1627 ( new_n1970_, new_n1969_, N219 );
not g1628 ( new_n1971_, new_n1970_ );
nand g1629 ( new_n1972_, new_n1971_, new_n1968_ );
nand g1630 ( new_n1973_, N91, N210 );
nand g1631 ( new_n1974_, new_n1972_, new_n1973_ );
nand g1632 ( new_n1975_, new_n1974_, new_n1914_ );
nor g1633 ( new_n1976_, new_n1970_, new_n1967_ );
not g1634 ( new_n1977_, new_n1973_ );
nor g1635 ( new_n1978_, new_n1976_, new_n1977_ );
nand g1636 ( new_n1979_, new_n1978_, keyIn_0_251 );
nand g1637 ( new_n1980_, new_n1975_, new_n1979_ );
nand g1638 ( new_n1981_, new_n1951_, N228 );
not g1639 ( new_n1982_, new_n1656_ );
nand g1640 ( new_n1983_, new_n1982_, N237 );
nand g1641 ( new_n1984_, new_n1981_, new_n1983_ );
nand g1642 ( new_n1985_, new_n1984_, keyIn_0_193 );
not g1643 ( new_n1986_, keyIn_0_146 );
nor g1644 ( new_n1987_, new_n1515_, new_n1247_ );
not g1645 ( new_n1988_, new_n1987_ );
nand g1646 ( new_n1989_, new_n1988_, keyIn_0_123 );
not g1647 ( new_n1990_, new_n1989_ );
nor g1648 ( new_n1991_, new_n1988_, keyIn_0_123 );
nor g1649 ( new_n1992_, new_n1990_, new_n1991_ );
nor g1650 ( new_n1993_, new_n1250_, new_n585_ );
nor g1651 ( new_n1994_, new_n1992_, new_n1993_ );
nor g1652 ( new_n1995_, new_n1994_, new_n1986_ );
nand g1653 ( new_n1996_, new_n1994_, new_n1986_ );
not g1654 ( new_n1997_, new_n1996_ );
nor g1655 ( new_n1998_, new_n1997_, new_n1995_ );
nor g1656 ( new_n1999_, new_n1984_, keyIn_0_193 );
nor g1657 ( new_n2000_, new_n1999_, new_n1998_ );
nand g1658 ( new_n2001_, new_n2000_, new_n1985_ );
not g1659 ( new_n2002_, new_n2001_ );
nand g1660 ( new_n2003_, new_n1980_, new_n2002_ );
nand g1661 ( new_n2004_, new_n2003_, new_n1913_ );
nor g1662 ( new_n2005_, new_n1978_, keyIn_0_251 );
nor g1663 ( new_n2006_, new_n1974_, new_n1914_ );
nor g1664 ( new_n2007_, new_n2006_, new_n2005_ );
nor g1665 ( new_n2008_, new_n2007_, new_n2001_ );
nand g1666 ( new_n2009_, new_n2008_, keyIn_0_254 );
nand g1667 ( N879, new_n2009_, new_n2004_ );
not g1668 ( new_n2011_, keyIn_0_252 );
nor g1669 ( new_n2012_, new_n1565_, new_n1637_ );
not g1670 ( new_n2013_, new_n2012_ );
nor g1671 ( new_n2014_, new_n2013_, keyIn_0_148 );
nand g1672 ( new_n2015_, new_n2013_, keyIn_0_148 );
not g1673 ( new_n2016_, new_n2015_ );
nor g1674 ( new_n2017_, new_n2016_, new_n2014_ );
not g1675 ( new_n2018_, keyIn_0_228 );
not g1676 ( new_n2019_, keyIn_0_223 );
nor g1677 ( new_n2020_, new_n1693_, new_n2019_ );
not g1678 ( new_n2021_, new_n2020_ );
nor g1679 ( new_n2022_, new_n1626_, keyIn_0_223 );
not g1680 ( new_n2023_, keyIn_0_171 );
nor g1681 ( new_n2024_, new_n1676_, new_n2023_ );
nand g1682 ( new_n2025_, new_n1676_, new_n2023_ );
not g1683 ( new_n2026_, new_n2025_ );
nor g1684 ( new_n2027_, new_n2026_, new_n2024_ );
not g1685 ( new_n2028_, new_n2027_ );
nor g1686 ( new_n2029_, new_n2022_, new_n2028_ );
nand g1687 ( new_n2030_, new_n2029_, new_n2021_ );
nor g1688 ( new_n2031_, new_n2030_, new_n2018_ );
not g1689 ( new_n2032_, new_n2031_ );
nand g1690 ( new_n2033_, new_n2030_, new_n2018_ );
nand g1691 ( new_n2034_, new_n2032_, new_n2033_ );
nand g1692 ( new_n2035_, new_n2034_, new_n2017_ );
nor g1693 ( new_n2036_, new_n2035_, keyIn_0_237 );
not g1694 ( new_n2037_, new_n2036_ );
nand g1695 ( new_n2038_, new_n2035_, keyIn_0_237 );
nand g1696 ( new_n2039_, new_n2037_, new_n2038_ );
nor g1697 ( new_n2040_, new_n2034_, new_n2017_ );
nor g1698 ( new_n2041_, new_n2040_, keyIn_0_238 );
not g1699 ( new_n2042_, new_n2041_ );
nand g1700 ( new_n2043_, new_n2040_, keyIn_0_238 );
nand g1701 ( new_n2044_, new_n2042_, new_n2043_ );
nand g1702 ( new_n2045_, new_n2044_, new_n2039_ );
nand g1703 ( new_n2046_, new_n2045_, keyIn_0_246 );
nor g1704 ( new_n2047_, new_n2045_, keyIn_0_246 );
nor g1705 ( new_n2048_, new_n2047_, new_n988_ );
nand g1706 ( new_n2049_, new_n2048_, new_n2046_ );
nand g1707 ( new_n2050_, N96, N210 );
nand g1708 ( new_n2051_, new_n2049_, new_n2050_ );
nand g1709 ( new_n2052_, new_n2051_, new_n2011_ );
nor g1710 ( new_n2053_, new_n2051_, new_n2011_ );
not g1711 ( new_n2054_, keyIn_0_170 );
nor g1712 ( new_n2055_, new_n1642_, new_n1230_ );
nor g1713 ( new_n2056_, new_n2055_, new_n2054_ );
nand g1714 ( new_n2057_, new_n2055_, new_n2054_ );
not g1715 ( new_n2058_, new_n2057_ );
nor g1716 ( new_n2059_, new_n2058_, new_n2056_ );
nor g1717 ( new_n2060_, new_n2017_, new_n1223_ );
nor g1718 ( new_n2061_, new_n2059_, new_n2060_ );
not g1719 ( new_n2062_, new_n2061_ );
nand g1720 ( new_n2063_, new_n2062_, keyIn_0_194 );
not g1721 ( new_n2064_, keyIn_0_126 );
nor g1722 ( new_n2065_, new_n1557_, new_n1247_ );
not g1723 ( new_n2066_, new_n2065_ );
nor g1724 ( new_n2067_, new_n2066_, new_n2064_ );
nand g1725 ( new_n2068_, new_n973_, N171 );
nand g1726 ( new_n2069_, new_n2066_, new_n2064_ );
nand g1727 ( new_n2070_, new_n2069_, new_n2068_ );
nor g1728 ( new_n2071_, new_n2070_, new_n2067_ );
nor g1729 ( new_n2072_, new_n2071_, keyIn_0_149 );
nand g1730 ( new_n2073_, new_n2071_, keyIn_0_149 );
not g1731 ( new_n2074_, new_n2073_ );
nor g1732 ( new_n2075_, new_n2074_, new_n2072_ );
nor g1733 ( new_n2076_, new_n2062_, keyIn_0_194 );
nor g1734 ( new_n2077_, new_n2076_, new_n2075_ );
nand g1735 ( new_n2078_, new_n2077_, new_n2063_ );
nor g1736 ( new_n2079_, new_n2053_, new_n2078_ );
nand g1737 ( new_n2080_, new_n2079_, new_n2052_ );
nand g1738 ( new_n2081_, new_n2080_, keyIn_0_255 );
not g1739 ( new_n2082_, keyIn_0_255 );
not g1740 ( new_n2083_, new_n2052_ );
not g1741 ( new_n2084_, new_n2046_ );
not g1742 ( new_n2085_, keyIn_0_246 );
not g1743 ( new_n2086_, new_n2038_ );
nor g1744 ( new_n2087_, new_n2086_, new_n2036_ );
not g1745 ( new_n2088_, new_n2043_ );
nor g1746 ( new_n2089_, new_n2088_, new_n2041_ );
nor g1747 ( new_n2090_, new_n2089_, new_n2087_ );
nand g1748 ( new_n2091_, new_n2090_, new_n2085_ );
nand g1749 ( new_n2092_, new_n2091_, N219 );
nor g1750 ( new_n2093_, new_n2092_, new_n2084_ );
not g1751 ( new_n2094_, new_n2050_ );
nor g1752 ( new_n2095_, new_n2093_, new_n2094_ );
nand g1753 ( new_n2096_, new_n2095_, keyIn_0_252 );
not g1754 ( new_n2097_, new_n2078_ );
nand g1755 ( new_n2098_, new_n2096_, new_n2097_ );
nor g1756 ( new_n2099_, new_n2098_, new_n2083_ );
nand g1757 ( new_n2100_, new_n2099_, new_n2082_ );
nand g1758 ( N880, new_n2100_, new_n2081_ );
endmodule