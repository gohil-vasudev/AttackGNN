module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n288_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n246_, new_n170_, new_n266_, new_n367_, new_n173_, new_n220_, new_n419_, new_n214_, new_n451_, new_n489_, new_n424_, new_n114_, new_n188_, new_n240_, new_n413_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n462_, new_n317_, new_n287_, new_n234_, new_n472_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n212_, new_n364_, new_n449_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n110_, new_n315_, new_n124_, new_n326_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n350_, new_n117_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n150_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n351_, new_n325_, new_n180_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n205_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n256_, new_n452_, new_n381_, new_n388_, new_n194_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n165_, new_n441_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n140_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n488_, new_n277_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n436_, new_n397_, new_n399_, new_n233_, new_n469_, new_n391_, new_n178_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n113_, new_n371_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n130_, new_n268_, new_n374_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n126_, new_n177_, new_n493_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n125_, new_n145_, new_n253_, new_n403_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n107_, new_n182_, new_n480_, new_n151_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n428_, new_n199_, new_n146_, new_n302_, new_n191_, new_n225_, new_n387_, new_n476_, new_n112_, new_n121_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n459_, new_n174_, new_n354_, new_n392_, new_n444_, new_n340_, new_n147_, new_n285_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n332_, new_n453_, new_n163_, new_n148_, new_n440_, new_n122_, new_n111_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n115_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n134_, new_n109_, new_n265_, new_n370_, new_n278_, new_n304_, new_n217_, new_n269_, new_n129_, new_n412_, new_n327_, new_n495_, new_n196_, new_n319_, new_n338_, new_n336_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n128_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n455_, new_n120_, new_n406_, new_n356_, new_n229_, new_n204_, new_n181_, new_n135_, new_n405_;

xor g000 ( new_n106_, N65, N69 );
xnor g001 ( new_n107_, N73, N77 );
xnor g002 ( new_n108_, new_n106_, new_n107_ );
xor g003 ( new_n109_, N81, N85 );
xnor g004 ( new_n110_, N89, N93 );
xnor g005 ( new_n111_, new_n109_, new_n110_ );
xor g006 ( new_n112_, new_n108_, new_n111_ );
nand g007 ( new_n113_, N129, N137 );
xnor g008 ( new_n114_, new_n112_, new_n113_ );
xnor g009 ( new_n115_, N1, N17 );
xnor g010 ( new_n116_, N33, N49 );
xnor g011 ( new_n117_, new_n115_, new_n116_ );
xnor g012 ( new_n118_, new_n114_, new_n117_ );
not g013 ( new_n119_, keyIn_0_9 );
xnor g014 ( new_n120_, N41, N45 );
xnor g015 ( new_n121_, new_n120_, keyIn_0_3 );
not g016 ( new_n122_, keyIn_0_2 );
xor g017 ( new_n123_, N33, N37 );
nand g018 ( new_n124_, new_n123_, new_n122_ );
xnor g019 ( new_n125_, N33, N37 );
nand g020 ( new_n126_, new_n125_, keyIn_0_2 );
nand g021 ( new_n127_, new_n124_, new_n126_ );
nand g022 ( new_n128_, new_n121_, new_n127_ );
not g023 ( new_n129_, keyIn_0_3 );
xnor g024 ( new_n130_, new_n120_, new_n129_ );
xnor g025 ( new_n131_, new_n125_, new_n122_ );
nand g026 ( new_n132_, new_n130_, new_n131_ );
nand g027 ( new_n133_, new_n132_, new_n128_ );
xnor g028 ( new_n134_, new_n133_, keyIn_0_7 );
not g029 ( new_n135_, keyIn_0_5 );
xnor g030 ( new_n136_, N57, N61 );
xnor g031 ( new_n137_, new_n136_, new_n135_ );
not g032 ( new_n138_, keyIn_0_4 );
nand g033 ( new_n139_, N49, N53 );
not g034 ( new_n140_, new_n139_ );
nor g035 ( new_n141_, N49, N53 );
nor g036 ( new_n142_, new_n140_, new_n141_ );
nand g037 ( new_n143_, new_n142_, new_n138_ );
xnor g038 ( new_n144_, N49, N53 );
nand g039 ( new_n145_, new_n144_, keyIn_0_4 );
nand g040 ( new_n146_, new_n143_, new_n145_ );
nand g041 ( new_n147_, new_n137_, new_n146_ );
nand g042 ( new_n148_, new_n136_, keyIn_0_5 );
xor g043 ( new_n149_, N57, N61 );
nand g044 ( new_n150_, new_n149_, new_n135_ );
nand g045 ( new_n151_, new_n150_, new_n148_ );
xnor g046 ( new_n152_, new_n144_, new_n138_ );
nand g047 ( new_n153_, new_n152_, new_n151_ );
nand g048 ( new_n154_, new_n153_, new_n147_ );
nand g049 ( new_n155_, new_n154_, keyIn_0_8 );
not g050 ( new_n156_, keyIn_0_8 );
xnor g051 ( new_n157_, new_n151_, new_n146_ );
nand g052 ( new_n158_, new_n157_, new_n156_ );
nand g053 ( new_n159_, new_n158_, new_n155_ );
nand g054 ( new_n160_, new_n134_, new_n159_ );
not g055 ( new_n161_, keyIn_0_7 );
xnor g056 ( new_n162_, new_n133_, new_n161_ );
xnor g057 ( new_n163_, new_n154_, new_n156_ );
nand g058 ( new_n164_, new_n162_, new_n163_ );
nand g059 ( new_n165_, new_n164_, new_n160_ );
nand g060 ( new_n166_, new_n165_, new_n119_ );
xnor g061 ( new_n167_, new_n162_, new_n159_ );
nand g062 ( new_n168_, new_n167_, keyIn_0_9 );
nand g063 ( new_n169_, new_n168_, new_n166_ );
nand g064 ( new_n170_, N134, N137 );
not g065 ( new_n171_, new_n170_ );
nand g066 ( new_n172_, new_n169_, new_n171_ );
xnor g067 ( new_n173_, new_n165_, keyIn_0_9 );
nand g068 ( new_n174_, new_n173_, new_n170_ );
nand g069 ( new_n175_, new_n174_, new_n172_ );
nand g070 ( new_n176_, new_n175_, keyIn_0_11 );
not g071 ( new_n177_, keyIn_0_11 );
xnor g072 ( new_n178_, new_n169_, new_n170_ );
nand g073 ( new_n179_, new_n178_, new_n177_ );
nand g074 ( new_n180_, new_n179_, new_n176_ );
xnor g075 ( new_n181_, N69, N85 );
xnor g076 ( new_n182_, N101, N117 );
xnor g077 ( new_n183_, new_n181_, new_n182_ );
not g078 ( new_n184_, new_n183_ );
nand g079 ( new_n185_, new_n180_, new_n184_ );
xnor g080 ( new_n186_, new_n175_, new_n177_ );
nand g081 ( new_n187_, new_n186_, new_n183_ );
nand g082 ( new_n188_, new_n187_, new_n185_ );
nand g083 ( new_n189_, new_n188_, keyIn_0_13 );
not g084 ( new_n190_, keyIn_0_13 );
xnor g085 ( new_n191_, new_n180_, new_n183_ );
nand g086 ( new_n192_, new_n191_, new_n190_ );
nand g087 ( new_n193_, new_n192_, new_n189_ );
nand g088 ( new_n194_, new_n193_, keyIn_0_15 );
not g089 ( new_n195_, keyIn_0_15 );
xnor g090 ( new_n196_, new_n188_, new_n190_ );
nand g091 ( new_n197_, new_n196_, new_n195_ );
nand g092 ( new_n198_, new_n197_, new_n194_ );
not g093 ( new_n199_, keyIn_0_12 );
not g094 ( new_n200_, keyIn_0_6 );
xnor g095 ( new_n201_, N9, N13 );
xnor g096 ( new_n202_, new_n201_, keyIn_0_1 );
not g097 ( new_n203_, keyIn_0_0 );
nand g098 ( new_n204_, N1, N5 );
not g099 ( new_n205_, new_n204_ );
nor g100 ( new_n206_, N1, N5 );
nor g101 ( new_n207_, new_n205_, new_n206_ );
nand g102 ( new_n208_, new_n207_, new_n203_ );
xnor g103 ( new_n209_, N1, N5 );
nand g104 ( new_n210_, new_n209_, keyIn_0_0 );
nand g105 ( new_n211_, new_n208_, new_n210_ );
xnor g106 ( new_n212_, new_n202_, new_n211_ );
nand g107 ( new_n213_, new_n212_, new_n200_ );
not g108 ( new_n214_, keyIn_0_1 );
xnor g109 ( new_n215_, new_n201_, new_n214_ );
nand g110 ( new_n216_, new_n215_, new_n211_ );
xnor g111 ( new_n217_, new_n209_, new_n203_ );
nand g112 ( new_n218_, new_n202_, new_n217_ );
nand g113 ( new_n219_, new_n218_, new_n216_ );
nand g114 ( new_n220_, new_n219_, keyIn_0_6 );
nand g115 ( new_n221_, new_n213_, new_n220_ );
xnor g116 ( new_n222_, new_n162_, new_n221_ );
nand g117 ( new_n223_, new_n222_, keyIn_0_10 );
not g118 ( new_n224_, keyIn_0_10 );
nand g119 ( new_n225_, new_n134_, new_n221_ );
xnor g120 ( new_n226_, new_n219_, new_n200_ );
nand g121 ( new_n227_, new_n162_, new_n226_ );
nand g122 ( new_n228_, new_n227_, new_n225_ );
nand g123 ( new_n229_, new_n228_, new_n224_ );
nand g124 ( new_n230_, new_n223_, new_n229_ );
nand g125 ( new_n231_, N135, N137 );
not g126 ( new_n232_, new_n231_ );
xnor g127 ( new_n233_, new_n230_, new_n232_ );
nand g128 ( new_n234_, new_n233_, new_n199_ );
nand g129 ( new_n235_, new_n230_, new_n231_ );
xnor g130 ( new_n236_, new_n228_, keyIn_0_10 );
nand g131 ( new_n237_, new_n236_, new_n232_ );
nand g132 ( new_n238_, new_n237_, new_n235_ );
nand g133 ( new_n239_, new_n238_, keyIn_0_12 );
nand g134 ( new_n240_, new_n234_, new_n239_ );
xnor g135 ( new_n241_, N73, N89 );
xnor g136 ( new_n242_, N105, N121 );
xnor g137 ( new_n243_, new_n241_, new_n242_ );
nand g138 ( new_n244_, new_n240_, new_n243_ );
xnor g139 ( new_n245_, new_n238_, new_n199_ );
not g140 ( new_n246_, new_n243_ );
nand g141 ( new_n247_, new_n245_, new_n246_ );
nand g142 ( new_n248_, new_n247_, new_n244_ );
nand g143 ( new_n249_, new_n248_, keyIn_0_14 );
not g144 ( new_n250_, keyIn_0_14 );
xnor g145 ( new_n251_, new_n240_, new_n246_ );
nand g146 ( new_n252_, new_n251_, new_n250_ );
nand g147 ( new_n253_, new_n252_, new_n249_ );
xor g148 ( new_n254_, N17, N21 );
xnor g149 ( new_n255_, N25, N29 );
xnor g150 ( new_n256_, new_n254_, new_n255_ );
xnor g151 ( new_n257_, new_n159_, new_n256_ );
nand g152 ( new_n258_, N136, N137 );
xnor g153 ( new_n259_, new_n257_, new_n258_ );
xnor g154 ( new_n260_, N77, N93 );
xnor g155 ( new_n261_, N109, N125 );
xnor g156 ( new_n262_, new_n260_, new_n261_ );
xnor g157 ( new_n263_, new_n259_, new_n262_ );
not g158 ( new_n264_, new_n263_ );
nand g159 ( new_n265_, new_n253_, new_n264_ );
not g160 ( new_n266_, new_n118_ );
xnor g161 ( new_n267_, N113, N117 );
xnor g162 ( new_n268_, N121, N125 );
xnor g163 ( new_n269_, new_n267_, new_n268_ );
xnor g164 ( new_n270_, N97, N101 );
xnor g165 ( new_n271_, N105, N109 );
xnor g166 ( new_n272_, new_n270_, new_n271_ );
xor g167 ( new_n273_, new_n269_, new_n272_ );
nand g168 ( new_n274_, N130, N137 );
xnor g169 ( new_n275_, new_n273_, new_n274_ );
xnor g170 ( new_n276_, N5, N21 );
xnor g171 ( new_n277_, N37, N53 );
xnor g172 ( new_n278_, new_n276_, new_n277_ );
xnor g173 ( new_n279_, new_n275_, new_n278_ );
nor g174 ( new_n280_, new_n266_, new_n279_ );
xnor g175 ( new_n281_, new_n108_, new_n272_ );
nand g176 ( new_n282_, N131, N137 );
xnor g177 ( new_n283_, new_n281_, new_n282_ );
xnor g178 ( new_n284_, N9, N25 );
xnor g179 ( new_n285_, N41, N57 );
xnor g180 ( new_n286_, new_n284_, new_n285_ );
xor g181 ( new_n287_, new_n283_, new_n286_ );
nand g182 ( new_n288_, new_n280_, new_n287_ );
not g183 ( new_n289_, new_n279_ );
nor g184 ( new_n290_, new_n289_, new_n118_ );
nand g185 ( new_n291_, new_n290_, new_n287_ );
nand g186 ( new_n292_, new_n288_, new_n291_ );
xnor g187 ( new_n293_, new_n111_, new_n269_ );
nand g188 ( new_n294_, N132, N137 );
xnor g189 ( new_n295_, new_n293_, new_n294_ );
xor g190 ( new_n296_, N13, N29 );
xnor g191 ( new_n297_, N45, N61 );
xnor g192 ( new_n298_, new_n296_, new_n297_ );
xor g193 ( new_n299_, new_n295_, new_n298_ );
not g194 ( new_n300_, new_n299_ );
nand g195 ( new_n301_, new_n292_, new_n300_ );
xnor g196 ( new_n302_, new_n287_, new_n299_ );
nor g197 ( new_n303_, new_n118_, new_n279_ );
nand g198 ( new_n304_, new_n302_, new_n303_ );
nand g199 ( new_n305_, new_n301_, new_n304_ );
xnor g200 ( new_n306_, new_n305_, keyIn_0_17 );
xnor g201 ( new_n307_, new_n226_, new_n256_ );
nand g202 ( new_n308_, N133, N137 );
xnor g203 ( new_n309_, new_n307_, new_n308_ );
xor g204 ( new_n310_, N65, N81 );
xnor g205 ( new_n311_, N97, N113 );
xnor g206 ( new_n312_, new_n310_, new_n311_ );
xnor g207 ( new_n313_, new_n309_, new_n312_ );
not g208 ( new_n314_, new_n313_ );
nand g209 ( new_n315_, new_n306_, new_n314_ );
nor g210 ( new_n316_, new_n265_, new_n315_ );
nand g211 ( new_n317_, new_n316_, new_n198_ );
xnor g212 ( new_n318_, new_n317_, keyIn_0_18 );
nand g213 ( new_n319_, new_n318_, new_n118_ );
nand g214 ( new_n320_, new_n319_, keyIn_0_20 );
not g215 ( new_n321_, keyIn_0_20 );
xnor g216 ( new_n322_, new_n193_, new_n195_ );
xnor g217 ( new_n323_, new_n248_, new_n250_ );
nor g218 ( new_n324_, new_n323_, new_n263_ );
not g219 ( new_n325_, new_n315_ );
nand g220 ( new_n326_, new_n324_, new_n325_ );
nor g221 ( new_n327_, new_n322_, new_n326_ );
nand g222 ( new_n328_, new_n327_, keyIn_0_18 );
not g223 ( new_n329_, keyIn_0_18 );
nand g224 ( new_n330_, new_n317_, new_n329_ );
nand g225 ( new_n331_, new_n328_, new_n330_ );
nor g226 ( new_n332_, new_n331_, new_n266_ );
nand g227 ( new_n333_, new_n332_, new_n321_ );
nand g228 ( new_n334_, new_n333_, new_n320_ );
xnor g229 ( new_n335_, new_n334_, N1 );
nand g230 ( new_n336_, new_n335_, keyIn_0_26 );
not g231 ( new_n337_, keyIn_0_26 );
not g232 ( new_n338_, N1 );
nand g233 ( new_n339_, new_n334_, new_n338_ );
xnor g234 ( new_n340_, new_n319_, new_n321_ );
nand g235 ( new_n341_, new_n340_, N1 );
nand g236 ( new_n342_, new_n341_, new_n339_ );
nand g237 ( new_n343_, new_n342_, new_n337_ );
nand g238 ( N724, new_n336_, new_n343_ );
not g239 ( new_n345_, N5 );
nand g240 ( new_n346_, new_n318_, new_n279_ );
nand g241 ( new_n347_, new_n346_, keyIn_0_21 );
not g242 ( new_n348_, keyIn_0_21 );
nor g243 ( new_n349_, new_n331_, new_n289_ );
nand g244 ( new_n350_, new_n349_, new_n348_ );
nand g245 ( new_n351_, new_n350_, new_n347_ );
xnor g246 ( new_n352_, new_n351_, new_n345_ );
nand g247 ( new_n353_, new_n352_, keyIn_0_27 );
not g248 ( new_n354_, keyIn_0_27 );
nand g249 ( new_n355_, new_n351_, N5 );
xnor g250 ( new_n356_, new_n346_, new_n348_ );
nand g251 ( new_n357_, new_n356_, new_n345_ );
nand g252 ( new_n358_, new_n357_, new_n355_ );
nand g253 ( new_n359_, new_n358_, new_n354_ );
nand g254 ( N725, new_n353_, new_n359_ );
not g255 ( new_n361_, keyIn_0_28 );
not g256 ( new_n362_, new_n287_ );
nand g257 ( new_n363_, new_n318_, new_n362_ );
nand g258 ( new_n364_, new_n363_, keyIn_0_22 );
not g259 ( new_n365_, keyIn_0_22 );
nor g260 ( new_n366_, new_n331_, new_n287_ );
nand g261 ( new_n367_, new_n366_, new_n365_ );
nand g262 ( new_n368_, new_n367_, new_n364_ );
xnor g263 ( new_n369_, new_n368_, N9 );
nand g264 ( new_n370_, new_n369_, new_n361_ );
not g265 ( new_n371_, N9 );
nand g266 ( new_n372_, new_n368_, new_n371_ );
xnor g267 ( new_n373_, new_n363_, new_n365_ );
nand g268 ( new_n374_, new_n373_, N9 );
nand g269 ( new_n375_, new_n374_, new_n372_ );
nand g270 ( new_n376_, new_n375_, keyIn_0_28 );
nand g271 ( N726, new_n370_, new_n376_ );
nand g272 ( new_n378_, new_n318_, new_n299_ );
nand g273 ( new_n379_, new_n378_, keyIn_0_23 );
not g274 ( new_n380_, keyIn_0_23 );
nor g275 ( new_n381_, new_n331_, new_n300_ );
nand g276 ( new_n382_, new_n381_, new_n380_ );
nand g277 ( new_n383_, new_n382_, new_n379_ );
xnor g278 ( new_n384_, new_n383_, N13 );
nand g279 ( new_n385_, new_n384_, keyIn_0_29 );
not g280 ( new_n386_, keyIn_0_29 );
not g281 ( new_n387_, N13 );
nand g282 ( new_n388_, new_n383_, new_n387_ );
xnor g283 ( new_n389_, new_n378_, new_n380_ );
nand g284 ( new_n390_, new_n389_, N13 );
nand g285 ( new_n391_, new_n390_, new_n388_ );
nand g286 ( new_n392_, new_n391_, new_n386_ );
nand g287 ( N727, new_n385_, new_n392_ );
nor g288 ( new_n394_, new_n193_, new_n313_ );
nand g289 ( new_n395_, new_n306_, new_n263_ );
nor g290 ( new_n396_, new_n395_, new_n253_ );
nand g291 ( new_n397_, new_n396_, new_n394_ );
nor g292 ( new_n398_, new_n397_, keyIn_0_19 );
nand g293 ( new_n399_, new_n397_, keyIn_0_19 );
nand g294 ( new_n400_, new_n399_, new_n118_ );
nor g295 ( new_n401_, new_n400_, new_n398_ );
xor g296 ( N728, new_n401_, N17 );
nand g297 ( new_n403_, new_n399_, new_n279_ );
nor g298 ( new_n404_, new_n403_, new_n398_ );
xnor g299 ( new_n405_, new_n404_, keyIn_0_24 );
xnor g300 ( new_n406_, new_n405_, N21 );
xnor g301 ( N729, new_n406_, keyIn_0_30 );
nand g302 ( new_n408_, new_n399_, new_n362_ );
nor g303 ( new_n409_, new_n408_, new_n398_ );
xor g304 ( N730, new_n409_, N25 );
nand g305 ( new_n411_, new_n399_, new_n299_ );
nor g306 ( new_n412_, new_n411_, new_n398_ );
xnor g307 ( new_n413_, new_n412_, keyIn_0_25 );
xnor g308 ( new_n414_, new_n413_, N29 );
xnor g309 ( N731, new_n414_, keyIn_0_31 );
nor g310 ( new_n416_, new_n196_, new_n314_ );
not g311 ( new_n417_, new_n306_ );
nor g312 ( new_n418_, new_n265_, new_n417_ );
nand g313 ( new_n419_, new_n418_, new_n416_ );
nor g314 ( new_n420_, new_n419_, new_n266_ );
xor g315 ( N732, new_n420_, N33 );
nor g316 ( new_n422_, new_n419_, new_n289_ );
xor g317 ( N733, new_n422_, N37 );
nor g318 ( new_n424_, new_n419_, new_n287_ );
xor g319 ( N734, new_n424_, N41 );
nor g320 ( new_n426_, new_n419_, new_n300_ );
xor g321 ( N735, new_n426_, N45 );
nand g322 ( new_n428_, new_n416_, new_n323_ );
nor g323 ( new_n429_, new_n428_, new_n395_ );
nand g324 ( new_n430_, new_n429_, new_n118_ );
xnor g325 ( N736, new_n430_, N49 );
nand g326 ( new_n432_, new_n429_, new_n279_ );
xnor g327 ( N737, new_n432_, N53 );
nand g328 ( new_n434_, new_n429_, new_n362_ );
xnor g329 ( N738, new_n434_, N57 );
nand g330 ( new_n436_, new_n429_, new_n299_ );
xnor g331 ( N739, new_n436_, N61 );
nand g332 ( new_n438_, new_n253_, keyIn_0_16 );
not g333 ( new_n439_, new_n394_ );
nor g334 ( new_n440_, new_n253_, keyIn_0_16 );
nor g335 ( new_n441_, new_n439_, new_n440_ );
nand g336 ( new_n442_, new_n441_, new_n438_ );
nand g337 ( new_n443_, new_n442_, new_n428_ );
nand g338 ( new_n444_, new_n443_, new_n264_ );
nand g339 ( new_n445_, new_n323_, new_n263_ );
nand g340 ( new_n446_, new_n445_, new_n265_ );
nor g341 ( new_n447_, new_n193_, new_n314_ );
nand g342 ( new_n448_, new_n446_, new_n447_ );
nand g343 ( new_n449_, new_n444_, new_n448_ );
nand g344 ( new_n450_, new_n449_, new_n314_ );
not g345 ( new_n451_, new_n450_ );
not g346 ( new_n452_, new_n280_ );
nand g347 ( new_n453_, new_n362_, new_n300_ );
nor g348 ( new_n454_, new_n452_, new_n453_ );
nand g349 ( new_n455_, new_n451_, new_n454_ );
xnor g350 ( N740, new_n455_, N65 );
nand g351 ( new_n457_, new_n449_, new_n193_ );
not g352 ( new_n458_, new_n457_ );
nand g353 ( new_n459_, new_n458_, new_n454_ );
xnor g354 ( N741, new_n459_, N69 );
nand g355 ( new_n461_, new_n449_, new_n253_ );
not g356 ( new_n462_, new_n461_ );
nand g357 ( new_n463_, new_n462_, new_n454_ );
xnor g358 ( N742, new_n463_, N73 );
nand g359 ( new_n465_, new_n449_, new_n263_ );
not g360 ( new_n466_, new_n465_ );
nand g361 ( new_n467_, new_n466_, new_n454_ );
xnor g362 ( N743, new_n467_, N77 );
nor g363 ( new_n469_, new_n288_, new_n300_ );
nand g364 ( new_n470_, new_n451_, new_n469_ );
xnor g365 ( N744, new_n470_, N81 );
nand g366 ( new_n472_, new_n458_, new_n469_ );
xnor g367 ( N745, new_n472_, N85 );
nand g368 ( new_n474_, new_n462_, new_n469_ );
xnor g369 ( N746, new_n474_, N89 );
nand g370 ( new_n476_, new_n466_, new_n469_ );
xnor g371 ( N747, new_n476_, N93 );
not g372 ( new_n478_, new_n290_ );
nor g373 ( new_n479_, new_n478_, new_n453_ );
nand g374 ( new_n480_, new_n451_, new_n479_ );
xnor g375 ( N748, new_n480_, N97 );
nand g376 ( new_n482_, new_n458_, new_n479_ );
xnor g377 ( N749, new_n482_, N101 );
nand g378 ( new_n484_, new_n462_, new_n479_ );
xnor g379 ( N750, new_n484_, N105 );
nand g380 ( new_n486_, new_n466_, new_n479_ );
xnor g381 ( N751, new_n486_, N109 );
nor g382 ( new_n488_, new_n291_, new_n300_ );
nand g383 ( new_n489_, new_n451_, new_n488_ );
xnor g384 ( N752, new_n489_, N113 );
nand g385 ( new_n491_, new_n458_, new_n488_ );
xnor g386 ( N753, new_n491_, N117 );
nand g387 ( new_n493_, new_n462_, new_n488_ );
xnor g388 ( N754, new_n493_, N121 );
nand g389 ( new_n495_, new_n466_, new_n488_ );
xnor g390 ( N755, new_n495_, N125 );
endmodule